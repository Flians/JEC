/*

c432:
	jxor: 1
	jspl: 84
	jspl3: 38
	jnot: 50
	jcb: 96
	jdff: 691
	jand: 92

Summary:
	jxor: 1
	jspl: 84
	jspl3: 38
	jnot: 50
	jcb: 96
	jdff: 691
	jand: 92
*/

module golden_c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G4gat_0;
	wire [2:0] w_G8gat_0;
	wire [1:0] w_G11gat_0;
	wire [1:0] w_G14gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G21gat_0;
	wire [2:0] w_G24gat_0;
	wire [1:0] w_G27gat_0;
	wire [2:0] w_G30gat_0;
	wire [2:0] w_G34gat_0;
	wire [1:0] w_G37gat_0;
	wire [2:0] w_G40gat_0;
	wire [2:0] w_G43gat_0;
	wire [1:0] w_G47gat_0;
	wire [2:0] w_G50gat_0;
	wire [1:0] w_G53gat_0;
	wire [2:0] w_G56gat_0;
	wire [2:0] w_G60gat_0;
	wire [1:0] w_G63gat_0;
	wire [1:0] w_G66gat_0;
	wire [2:0] w_G69gat_0;
	wire [1:0] w_G73gat_0;
	wire [1:0] w_G76gat_0;
	wire [1:0] w_G79gat_0;
	wire [2:0] w_G82gat_0;
	wire [2:0] w_G86gat_0;
	wire [2:0] w_G89gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G95gat_0;
	wire [2:0] w_G99gat_0;
	wire [1:0] w_G102gat_0;
	wire [1:0] w_G105gat_0;
	wire [1:0] w_G112gat_0;
	wire [1:0] w_G115gat_0;
	wire [2:0] w_G223gat_0;
	wire [2:0] w_G223gat_1;
	wire [2:0] w_G223gat_2;
	wire [1:0] w_G223gat_3;
	wire G223gat_fa_;
	wire [2:0] w_G329gat_0;
	wire [2:0] w_G329gat_1;
	wire [2:0] w_G329gat_2;
	wire [2:0] w_G329gat_3;
	wire w_G329gat_4;
	wire G329gat_fa_;
	wire [2:0] w_G370gat_0;
	wire [2:0] w_G370gat_1;
	wire w_G370gat_2;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire [1:0] w_n44_0;
	wire [1:0] w_n46_0;
	wire [1:0] w_n48_0;
	wire [1:0] w_n49_0;
	wire [1:0] w_n51_0;
	wire [1:0] w_n54_0;
	wire [1:0] w_n57_0;
	wire [1:0] w_n60_0;
	wire [1:0] w_n61_0;
	wire [1:0] w_n63_0;
	wire [1:0] w_n65_0;
	wire [1:0] w_n73_0;
	wire [1:0] w_n75_0;
	wire [1:0] w_n80_0;
	wire [1:0] w_n81_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n86_0;
	wire [2:0] w_n91_0;
	wire [2:0] w_n91_1;
	wire [2:0] w_n91_2;
	wire [1:0] w_n91_3;
	wire [1:0] w_n93_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n100_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n105_0;
	wire [1:0] w_n110_0;
	wire [1:0] w_n112_0;
	wire [1:0] w_n114_0;
	wire [1:0] w_n116_0;
	wire [1:0] w_n122_0;
	wire [1:0] w_n123_0;
	wire [1:0] w_n128_0;
	wire [1:0] w_n130_0;
	wire [1:0] w_n137_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n142_0;
	wire [1:0] w_n146_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n155_0;
	wire [1:0] w_n161_0;
	wire [1:0] w_n164_0;
	wire [2:0] w_n169_0;
	wire [2:0] w_n169_1;
	wire [1:0] w_n175_0;
	wire [1:0] w_n179_0;
	wire [1:0] w_n182_0;
	wire [1:0] w_n188_0;
	wire [1:0] w_n189_0;
	wire [1:0] w_n192_0;
	wire [1:0] w_n195_0;
	wire [1:0] w_n197_0;
	wire [1:0] w_n201_0;
	wire [1:0] w_n202_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n209_0;
	wire [1:0] w_n218_0;
	wire [1:0] w_n222_0;
	wire [1:0] w_n225_0;
	wire [1:0] w_n226_0;
	wire [2:0] w_n230_0;
	wire [2:0] w_n230_1;
	wire [2:0] w_n230_2;
	wire [1:0] w_n232_0;
	wire [1:0] w_n234_0;
	wire [1:0] w_n235_0;
	wire [1:0] w_n240_0;
	wire [1:0] w_n243_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n257_0;
	wire [1:0] w_n270_0;
	wire [1:0] w_n272_0;
	wire [1:0] w_n274_0;
	wire w_dff_B_e5alEDkm0_1;
	wire w_dff_B_zc14q3Ww4_0;
	wire w_dff_B_Rr9P4l8Q2_1;
	wire w_dff_B_EKguxQvI2_1;
	wire w_dff_B_0Q6AgxcI3_1;
	wire w_dff_B_hLwXVtbl0_1;
	wire w_dff_B_ygjXYEtf8_1;
	wire w_dff_B_0XZKHc2f5_1;
	wire w_dff_B_smGAGvqp0_1;
	wire w_dff_B_JeATEhhI8_1;
	wire w_dff_B_CdWLwGFg8_1;
	wire w_dff_B_LYVkKKH96_1;
	wire w_dff_B_lq94nuYA8_1;
	wire w_dff_B_0hwomlzi0_1;
	wire w_dff_B_dhJsoA2W5_1;
	wire w_dff_B_sEHsiY7T2_1;
	wire w_dff_B_n4zCBecB6_1;
	wire w_dff_B_mQ8whF5V8_1;
	wire w_dff_B_RnLAEkNG5_1;
	wire w_dff_B_KwMrbmoV3_1;
	wire w_dff_B_BdTi0qlL0_1;
	wire w_dff_A_8GoXyrJa8_1;
	wire w_dff_A_Na4phgtn5_1;
	wire w_dff_A_N54RAZRq8_0;
	wire w_dff_A_jj7v4i1G9_0;
	wire w_dff_A_cqO6S9JU5_1;
	wire w_dff_B_rayBSws80_1;
	wire w_dff_B_WkD10pJW1_1;
	wire w_dff_B_yz9qbQe82_1;
	wire w_dff_B_SIWxHZAL7_1;
	wire w_dff_B_fb5mko2J9_1;
	wire w_dff_B_MHJ9DvKA6_1;
	wire w_dff_B_KChWfxvy8_1;
	wire w_dff_B_EIxEtQhj8_1;
	wire w_dff_B_p1F4fnSJ6_1;
	wire w_dff_B_Xvud4s3Z8_1;
	wire w_dff_B_uREUa1EU9_1;
	wire w_dff_B_XE8vKwi15_1;
	wire w_dff_B_0cZ7qe8m5_1;
	wire w_dff_B_K8ntdtot9_1;
	wire w_dff_B_jkiZY0gw8_1;
	wire w_dff_B_frvgF7bQ7_1;
	wire w_dff_B_AKIuBdTm8_1;
	wire w_dff_B_FdGKqCue2_1;
	wire w_dff_B_EAwqKOMd2_1;
	wire w_dff_A_3iAJhNi49_0;
	wire w_dff_A_iVlygmfK3_0;
	wire w_dff_B_V5i3A9gs7_1;
	wire w_dff_B_XG3Vyga20_1;
	wire w_dff_B_IkpjPyrw7_1;
	wire w_dff_B_ingOgbsg1_1;
	wire w_dff_B_lBrJComX7_1;
	wire w_dff_B_qnaFo5Ee6_1;
	wire w_dff_B_YMdibU7c0_1;
	wire w_dff_B_LQCtmshq1_1;
	wire w_dff_B_Xpm6vzuh9_1;
	wire w_dff_B_GuTKXBH69_1;
	wire w_dff_B_1fx2u2iR2_1;
	wire w_dff_B_RuyKfXgE7_1;
	wire w_dff_B_cdGn0N916_1;
	wire w_dff_B_iPGAxZSf9_1;
	wire w_dff_B_Ii23Vlge6_1;
	wire w_dff_B_Ue4UedO57_1;
	wire w_dff_B_AfHVPBWM0_1;
	wire w_dff_B_qMH1XlYV7_1;
	wire w_dff_B_9PVZRrRo0_1;
	wire w_dff_B_luoa8u5s2_1;
	wire w_dff_B_HGx1crMw7_1;
	wire w_dff_B_isDjTFWc8_1;
	wire w_dff_B_G8pYIdzQ9_1;
	wire w_dff_B_qM6LeDhA0_1;
	wire w_dff_B_942GQbZg7_1;
	wire w_dff_B_KrePHkWA2_1;
	wire w_dff_B_LHgrEym81_1;
	wire w_dff_B_m7Ms08W15_1;
	wire w_dff_B_3qwx3fib2_1;
	wire w_dff_B_hOBeDdU87_1;
	wire w_dff_B_xuEOVQNx2_1;
	wire w_dff_B_O7GXZBuc5_1;
	wire w_dff_B_85UE8Pjn3_1;
	wire w_dff_B_elEKzFxD0_1;
	wire w_dff_B_7Q0HnyIn1_1;
	wire w_dff_B_RRNJMLFZ9_1;
	wire w_dff_B_WTRgCdbs0_1;
	wire w_dff_B_YKhgEew84_1;
	wire w_dff_A_GE2OFhcu2_0;
	wire w_dff_B_PVwqqQDq9_0;
	wire w_dff_B_ruU0o0Zw5_0;
	wire w_dff_B_8KuuX9pm7_0;
	wire w_dff_B_M9k5CzIM1_0;
	wire w_dff_B_yHQjgJuJ2_0;
	wire w_dff_A_ReIXFZ3E4_0;
	wire w_dff_A_n1HDuIrX2_0;
	wire w_dff_A_nCbuYFbF4_0;
	wire w_dff_A_lxuzfnML8_0;
	wire w_dff_A_XVDMd2Qt9_0;
	wire w_dff_A_xkJXqYtU3_0;
	wire w_dff_A_ShDyOuw69_0;
	wire w_dff_B_2ZtFWut93_0;
	wire w_dff_B_oo0lapOU4_0;
	wire w_dff_B_69rNmGGs0_0;
	wire w_dff_B_aQmgpujQ6_0;
	wire w_dff_B_tbSrLAWP7_0;
	wire w_dff_B_LZvlM0IF3_0;
	wire w_dff_B_KD1KIA7h3_0;
	wire w_dff_B_YG4D7ggH7_1;
	wire w_dff_A_PZkuwsVW8_0;
	wire w_dff_A_K4uxcDgn9_0;
	wire w_dff_A_NBc9thxJ3_0;
	wire w_dff_A_AqEWRHx37_0;
	wire w_dff_A_YqZae1nT9_0;
	wire w_dff_A_8AbjdZxs4_0;
	wire w_dff_A_k9U9pe132_0;
	wire w_dff_A_91Cc5cyW2_0;
	wire w_dff_A_8muuYSL54_0;
	wire w_dff_A_fsD8wDjC9_0;
	wire w_dff_A_DhUZeLp19_0;
	wire w_dff_A_PwgyT2Fz5_0;
	wire w_dff_A_WZUhTPdu1_0;
	wire w_dff_A_RQFR3mYA8_0;
	wire w_dff_A_gw2UTSY54_0;
	wire w_dff_A_HLs4KfFJ8_0;
	wire w_dff_A_UP7wXcvy4_0;
	wire w_dff_A_RBu1l1Gf3_0;
	wire w_dff_A_mujE1H1o5_0;
	wire w_dff_A_94zoQHuY9_0;
	wire w_dff_B_68N1zJpU2_0;
	wire w_dff_B_xtkQa4946_0;
	wire w_dff_A_6yfuLoDF4_1;
	wire w_dff_A_ieizIOyX8_1;
	wire w_dff_A_xy0oMfl79_1;
	wire w_dff_A_hAehK1Cs4_1;
	wire w_dff_A_lQHK98mN4_1;
	wire w_dff_A_zELgvyFN6_1;
	wire w_dff_A_McLi8ER78_1;
	wire w_dff_A_BZSrONRL7_1;
	wire w_dff_A_Vgh3MVZc3_1;
	wire w_dff_A_JoDMAQsU7_1;
	wire w_dff_A_8RULKxWV0_1;
	wire w_dff_A_CRsJpwR56_1;
	wire w_dff_A_Q92DefhQ6_1;
	wire w_dff_A_xq92GEQy6_1;
	wire w_dff_A_vyQkkCnx5_1;
	wire w_dff_A_nzXcZcit6_0;
	wire w_dff_A_UnTZFBYV3_0;
	wire w_dff_A_KP6Pf0ls0_0;
	wire w_dff_B_UGFk8mY89_1;
	wire w_dff_B_mJ4HpQ7e4_1;
	wire w_dff_B_cbneefmY0_1;
	wire w_dff_B_ktXJQKyJ8_1;
	wire w_dff_B_28ySflHm4_1;
	wire w_dff_B_r2GEpJMO4_1;
	wire w_dff_B_5GlQwz315_1;
	wire w_dff_B_XbRR5KLx1_1;
	wire w_dff_B_byLwmGvx2_1;
	wire w_dff_B_rVkOIyrO2_1;
	wire w_dff_B_MJYhPC8g8_1;
	wire w_dff_A_4yx1vEpq6_0;
	wire w_dff_A_9wHwzcwr9_0;
	wire w_dff_A_ZIdL7NhX7_0;
	wire w_dff_A_sPeF0eZf4_0;
	wire w_dff_A_YTtw4F179_0;
	wire w_dff_A_GvdEzcgx3_0;
	wire w_dff_A_2efNFSLi2_0;
	wire w_dff_A_7kLnfmXa8_0;
	wire w_dff_A_TJYPW7SA8_0;
	wire w_dff_A_Uc3CZSEp6_0;
	wire w_dff_A_rWyCF3Mx5_0;
	wire w_dff_A_dR0YlQd23_0;
	wire w_dff_A_vsUmunHW1_0;
	wire w_dff_A_yqAPWQ7j5_0;
	wire w_dff_A_E3aw4bMf4_0;
	wire w_dff_A_BnZcShms0_0;
	wire w_dff_A_8dErt7Uh6_0;
	wire w_dff_A_6TmgDA501_0;
	wire w_dff_B_XeoHgJba5_2;
	wire w_dff_B_GCytSAJh7_2;
	wire w_dff_B_2BS1ZbFY3_2;
	wire w_dff_B_iYUb8tV98_2;
	wire w_dff_B_LiqyjzZT8_2;
	wire w_dff_B_byhoR8gJ7_2;
	wire w_dff_B_XRDK1Pva7_2;
	wire w_dff_B_UuBqLHac4_2;
	wire w_dff_B_EU06pYH15_2;
	wire w_dff_B_o8r2mS3D1_2;
	wire w_dff_B_jOeKJE9G9_2;
	wire w_dff_A_5MIIGepJ3_0;
	wire w_dff_A_uvbPFJi35_0;
	wire w_dff_A_Li8I2X4j0_0;
	wire w_dff_A_QI6UNgV19_0;
	wire w_dff_A_CsTHdnFB4_0;
	wire w_dff_A_W2VpZEpB3_0;
	wire w_dff_A_E2fhySV26_0;
	wire w_dff_A_Sgzihm8T1_0;
	wire w_dff_A_tS1vBQgN2_0;
	wire w_dff_A_w2Gc8ey23_0;
	wire w_dff_A_YvMlf2Pl8_0;
	wire w_dff_A_aEGAr0Tv2_0;
	wire w_dff_A_aoQOdcg27_0;
	wire w_dff_A_wxXA6H3I1_0;
	wire w_dff_A_yS8gKoul0_0;
	wire w_dff_A_w8nMvLQ22_1;
	wire w_dff_A_mLWRzPG60_1;
	wire w_dff_A_UIu5GpSN2_1;
	wire w_dff_A_isKyIbqO3_1;
	wire w_dff_A_FyDsKn3i2_1;
	wire w_dff_A_rcjvKEdG1_1;
	wire w_dff_A_RxegrnXh8_1;
	wire w_dff_A_5SZFa6fs4_1;
	wire w_dff_A_tYJmetl42_1;
	wire w_dff_B_VmHWFZ5U6_0;
	wire w_dff_B_HDPAEKzA6_0;
	wire w_dff_B_U6hfzyHL4_0;
	wire w_dff_A_ojvFAyzI4_0;
	wire w_dff_A_WGyhBl7F5_0;
	wire w_dff_A_GzaeScc69_0;
	wire w_dff_A_ldma2cIp4_0;
	wire w_dff_A_EjkXA34m6_0;
	wire w_dff_A_L6DoBOc54_0;
	wire w_dff_A_atlUkYPM4_0;
	wire w_dff_A_Oiq5S9mx3_0;
	wire w_dff_B_ifLLn9bo9_2;
	wire w_dff_B_a9k85SDt9_2;
	wire w_dff_B_LcB3bNJq6_2;
	wire w_dff_B_SGpQRxIW2_2;
	wire w_dff_B_vmMr3mZX0_2;
	wire w_dff_B_oOjS4uHz8_2;
	wire w_dff_A_LjKIH6Ya0_0;
	wire w_dff_A_5Cq5ZEri1_0;
	wire w_dff_A_JaZGIrAh4_0;
	wire w_dff_A_dKayZWHU3_0;
	wire w_dff_A_7uakt8qp7_0;
	wire w_dff_A_2afSD2El5_0;
	wire w_dff_A_iP8barNH1_0;
	wire w_dff_A_GEdCW9EV8_0;
	wire w_dff_A_u3Rvaf0U0_0;
	wire w_dff_A_EMuH6fZS8_0;
	wire w_dff_A_HgpdXnc60_0;
	wire w_dff_A_e10ykomm2_0;
	wire w_dff_A_judq4vel5_0;
	wire w_dff_A_KPJ9DGpu2_0;
	wire w_dff_A_BerntqP88_0;
	wire w_dff_B_yd1ok6pc7_1;
	wire w_dff_B_1PuDcvmp9_1;
	wire w_dff_B_ODrf1TBp8_1;
	wire w_dff_B_stWsCTyc4_1;
	wire w_dff_B_mIss7T1O5_1;
	wire w_dff_B_ZQio1wDY4_1;
	wire w_dff_B_rqcJEdQT1_1;
	wire w_dff_B_E6Nltixk5_1;
	wire w_dff_B_ATBLh0m31_1;
	wire w_dff_B_gvt5VaHr4_1;
	wire w_dff_B_g91zQXQd2_1;
	wire w_dff_A_Ov4Q1z1y4_0;
	wire w_dff_A_CvHOYBHq4_0;
	wire w_dff_A_0yLVUsEt2_0;
	wire w_dff_A_iN07iLxl3_0;
	wire w_dff_A_yM4uPf3c8_0;
	wire w_dff_A_r9uPBkP90_0;
	wire w_dff_A_TbzDJM6C6_0;
	wire w_dff_A_0MstNCHM3_0;
	wire w_dff_A_ECgu0i0u9_0;
	wire w_dff_A_Ke94OlAN3_0;
	wire w_dff_A_Kwz5zZVd7_0;
	wire w_dff_A_c4I3kAog5_0;
	wire w_dff_A_gL4pC2X05_0;
	wire w_dff_A_9cCOg7SE5_0;
	wire w_dff_A_LKzdN1yI2_0;
	wire w_dff_A_m2r5LI4g3_1;
	wire w_dff_A_RhCgGiEP4_1;
	wire w_dff_A_GtfoIOcj3_1;
	wire w_dff_A_IDgJycOp3_1;
	wire w_dff_A_Dx5Cydes3_1;
	wire w_dff_A_h5yox54O9_1;
	wire w_dff_A_G22iVq2z4_1;
	wire w_dff_A_81gjq9Pq9_1;
	wire w_dff_A_61v04UO43_1;
	wire w_dff_B_xl0nsL2C9_0;
	wire w_dff_B_RncHQkKu0_0;
	wire w_dff_B_HQsFRl0s9_0;
	wire w_dff_B_zBaBPsNS7_1;
	wire w_dff_B_Yh1HPGxF1_1;
	wire w_dff_A_EKbmkh4Y2_1;
	wire w_dff_A_ixCgi5V25_1;
	wire w_dff_A_HISKe9X16_1;
	wire w_dff_A_v550qsGB8_1;
	wire w_dff_A_gBfxMIlS5_1;
	wire w_dff_A_GQIGf68I0_1;
	wire w_dff_A_E3VEHWhc4_1;
	wire w_dff_A_aEstPw1q1_1;
	wire w_dff_A_KLXF1nLE7_1;
	wire w_dff_A_uDNfJlIO6_1;
	wire w_dff_A_Un7fl79t1_1;
	wire w_dff_A_g0R80RuZ0_1;
	wire w_dff_A_bkIhgypG9_1;
	wire w_dff_A_pWNaMWyj8_1;
	wire w_dff_A_dSLAO5fQ6_1;
	wire w_dff_A_DNa8Zykm6_1;
	wire w_dff_A_iXkBClZk6_1;
	wire w_dff_A_jkf4lP8S1_1;
	wire w_dff_B_v9KblQxF4_1;
	wire w_dff_B_ja6GFkp55_1;
	wire w_dff_B_PKRTrW9k6_1;
	wire w_dff_B_qchdsOK64_1;
	wire w_dff_B_0eTdbLvy9_1;
	wire w_dff_B_4admQqlc7_1;
	wire w_dff_B_lCZrej0r6_1;
	wire w_dff_B_xArl4hZ86_1;
	wire w_dff_B_ZsflEea39_0;
	wire w_dff_B_B0uRk8bE6_0;
	wire w_dff_B_Dr7YYBEp1_0;
	wire w_dff_B_ekWoYZaN3_0;
	wire w_dff_A_6AUVUaT74_0;
	wire w_dff_A_GPKoMvTx2_0;
	wire w_dff_A_e6Vpsc8Y2_0;
	wire w_dff_A_RHIhLvQ85_0;
	wire w_dff_A_EvJ7Vh3W1_0;
	wire w_dff_A_rOnrJ9g02_0;
	wire w_dff_A_6APx0r583_0;
	wire w_dff_A_JcoH8Tot4_0;
	wire w_dff_A_DspAH3ge2_0;
	wire w_dff_A_2yC9AYMb3_0;
	wire w_dff_A_Iz7S5QaJ7_0;
	wire w_dff_A_VdyfJxk62_0;
	wire w_dff_A_M5ir2P5r5_0;
	wire w_dff_A_Ks7F7ZGn3_0;
	wire w_dff_A_LclFNCTp1_0;
	wire w_dff_A_aW0Pg6av4_0;
	wire w_dff_A_sU6PWbBk3_0;
	wire w_dff_A_F5CDsX0C8_0;
	wire w_dff_B_ZMk9tluA8_1;
	wire w_dff_B_whZGNrI84_1;
	wire w_dff_A_qcDIukFr1_0;
	wire w_dff_A_CBrLCcUq5_0;
	wire w_dff_A_UGzJx2Bv7_0;
	wire w_dff_A_qzvYOYxS1_0;
	wire w_dff_A_pI12VvBE9_0;
	wire w_dff_A_gM7zOEJQ0_0;
	wire w_dff_B_ehbpL0nn8_1;
	wire w_dff_B_J9UvRJ9I9_1;
	wire w_dff_A_oKx4W6Og0_0;
	wire w_dff_A_EaE462m80_0;
	wire w_dff_A_8pYhuuVD5_0;
	wire w_dff_B_bp6EqDuX6_2;
	wire w_dff_B_MRMhKywC7_2;
	wire w_dff_B_qkAUPKKp2_2;
	wire w_dff_B_mGAm7GE30_2;
	wire w_dff_B_SXsvtxlY5_2;
	wire w_dff_B_MQJwHhR13_2;
	wire w_dff_B_X3IFIq1E5_2;
	wire w_dff_B_BMfeVFkL4_2;
	wire w_dff_B_6Iq6BaXp3_2;
	wire w_dff_B_VAejou2l3_2;
	wire w_dff_B_rIMAXny88_2;
	wire w_dff_B_iw6PA2gg1_2;
	wire w_dff_A_dZlt55fP7_0;
	wire w_dff_A_EEO3t36o4_0;
	wire w_dff_A_3132Il2W8_0;
	wire w_dff_A_7MulR8yy0_0;
	wire w_dff_B_egok4NA54_2;
	wire w_dff_B_b1pIRL3U3_2;
	wire w_dff_B_WR30poUH6_2;
	wire w_dff_A_TNod6VTT8_1;
	wire w_dff_A_NEG1lOOz2_1;
	wire w_dff_A_dztB5kxU4_1;
	wire w_dff_A_AbIXbCDW2_1;
	wire w_dff_A_CdACMHy80_1;
	wire w_dff_A_XaNgq4Wh4_1;
	wire w_dff_A_mUeoM9Ob8_1;
	wire w_dff_A_r9qhEyp54_1;
	wire w_dff_A_32tvPrji5_1;
	wire w_dff_A_G3h19LpY7_1;
	wire w_dff_A_bzor4PHd8_1;
	wire w_dff_A_7bQosZHH0_1;
	wire w_dff_A_U1zaGshL6_1;
	wire w_dff_A_FWVp66n37_1;
	wire w_dff_A_CnWadUpS6_1;
	wire w_dff_A_eRHnONse6_1;
	wire w_dff_A_yddNCP299_0;
	wire w_dff_A_GX7VCkeK6_0;
	wire w_dff_A_CRZgAs995_0;
	wire w_dff_A_gmlFuxkv7_0;
	wire w_dff_A_ybgnrxKl4_0;
	wire w_dff_A_9qGbqOMD3_0;
	wire w_dff_A_SVFC7uqp2_0;
	wire w_dff_B_elRkFYIP3_0;
	wire w_dff_A_jr1oo0Bk8_0;
	wire w_dff_A_JzKVPRA03_0;
	wire w_dff_A_OxTkNlyu5_0;
	wire w_dff_A_e01KYA1J0_0;
	wire w_dff_A_iJcbkrHa8_0;
	wire w_dff_A_Yg723xQ76_0;
	wire w_dff_A_x56y1hzt5_0;
	wire w_dff_A_rKzxqIcD0_0;
	wire w_dff_A_cGOhxaoR0_0;
	wire w_dff_A_5Rh6wsVC1_0;
	wire w_dff_B_r3dWirN96_2;
	wire w_dff_B_LUhpJFK08_2;
	wire w_dff_B_O78DKDEn3_2;
	wire w_dff_B_70Yd7APk8_2;
	wire w_dff_B_Zq05Emy40_2;
	wire w_dff_A_zAA0bolL9_0;
	wire w_dff_A_JVtt5KWv5_0;
	wire w_dff_A_rIbykblP1_0;
	wire w_dff_A_AkIkxJsz1_0;
	wire w_dff_A_4IsB3gGg3_0;
	wire w_dff_A_HY3LHZsc6_0;
	wire w_dff_A_5S7pVowj7_0;
	wire w_dff_A_2IOI8oZH0_0;
	wire w_dff_A_4rivU3b73_1;
	wire w_dff_A_ONgI4wLQ4_1;
	wire w_dff_A_8VHJ7YhU7_1;
	wire w_dff_B_MKzUcZ2u5_1;
	wire w_dff_B_T1RyiQcr6_1;
	wire w_dff_B_4YMeAVOs6_1;
	wire w_dff_B_QxgWOeCq5_1;
	wire w_dff_B_yqZGaAPC1_1;
	wire w_dff_A_x0cHKmOc7_0;
	wire w_dff_A_xhtGRUz96_0;
	wire w_dff_A_5vld24Jq3_0;
	wire w_dff_A_OBS4fSpo0_0;
	wire w_dff_A_vSfKcLNB9_0;
	wire w_dff_A_cdwrfuQp7_0;
	wire w_dff_A_TGiIRNbj6_0;
	wire w_dff_A_vyxp6Eid2_0;
	wire w_dff_A_ca0oEeB29_1;
	wire w_dff_A_JEyxBdAt4_1;
	wire w_dff_A_tRoBYtPN0_1;
	wire w_dff_B_9XlDlqN57_1;
	wire w_dff_B_fDBYCPLl7_1;
	wire w_dff_B_IgVYzbtI3_1;
	wire w_dff_B_9uIeXScz6_1;
	wire w_dff_B_YmnvNTO67_1;
	wire w_dff_A_iFzmUClZ2_0;
	wire w_dff_A_Rtsu1nPa4_0;
	wire w_dff_A_SLRSDd8X8_0;
	wire w_dff_A_TfTh3ZeS9_0;
	wire w_dff_A_2M3cQGbu2_0;
	wire w_dff_A_G1e9RZwv5_0;
	wire w_dff_A_CEPNZffk8_0;
	wire w_dff_A_uC2MoJHC9_0;
	wire w_dff_A_MiHGDkhu9_0;
	wire w_dff_A_n4B4x9c09_0;
	wire w_dff_A_a13WHX4j7_0;
	wire w_dff_A_icucMoCM1_0;
	wire w_dff_A_lrvoPlfa9_0;
	wire w_dff_A_ANjHGxGf8_0;
	wire w_dff_A_FwTY1rTi7_0;
	wire w_dff_A_eCiT5ni34_0;
	wire w_dff_A_ukKvqtB41_0;
	wire w_dff_A_OUBJK5dB4_0;
	wire w_dff_B_7ACDJUSU9_2;
	wire w_dff_B_JxN8MC734_2;
	wire w_dff_B_6EjmAgtR4_2;
	wire w_dff_B_rq4XUosw7_2;
	wire w_dff_B_GZI4eWWi3_2;
	wire w_dff_A_j3XIiRRK8_0;
	wire w_dff_A_dPiO0LtP4_0;
	wire w_dff_A_yin4GHKJ1_0;
	wire w_dff_A_F264yvlv0_0;
	wire w_dff_A_Zvw3Jmy07_0;
	wire w_dff_A_GXzQ2Qv23_0;
	wire w_dff_A_nbwRWgXO1_0;
	wire w_dff_A_CNjBBjIk4_0;
	wire w_dff_A_BdrKwSXp0_1;
	wire w_dff_A_zcxX3cwF7_1;
	wire w_dff_A_jIh8pKnM9_1;
	wire w_dff_A_3xsKJLd08_0;
	wire w_dff_A_RX6PzHag1_0;
	wire w_dff_A_YwlIeDW40_0;
	wire w_dff_A_1U80RyWS9_0;
	wire w_dff_A_kRjQN2Aa7_0;
	wire w_dff_A_c2egbizS7_0;
	wire w_dff_A_As2HewtW1_0;
	wire w_dff_A_9BCtItK83_0;
	wire w_dff_A_Exk40fx50_0;
	wire w_dff_A_TYl7dF2w3_0;
	wire w_dff_B_V8hG2G8G4_2;
	wire w_dff_B_CzZGeQ8i5_2;
	wire w_dff_B_v0sDIqxd3_2;
	wire w_dff_B_8SX2Digw1_2;
	wire w_dff_B_HmDgpTZ25_2;
	wire w_dff_A_dkeOH2Ow1_0;
	wire w_dff_A_JUSfIm3S8_0;
	wire w_dff_A_S9xMJYHP2_0;
	wire w_dff_A_wU5caEIS7_0;
	wire w_dff_A_y0bfCXbb4_0;
	wire w_dff_A_DwLkY97D5_0;
	wire w_dff_A_mINrjOlD6_0;
	wire w_dff_A_JCeut76T7_0;
	wire w_dff_A_xRuxKaBe1_1;
	wire w_dff_A_pN0jcjOr6_1;
	wire w_dff_A_tqGg37gq2_1;
	wire w_dff_A_SdRqIHRY4_0;
	wire w_dff_A_Oiv6w4kd5_0;
	wire w_dff_A_M23sTneE8_0;
	wire w_dff_A_iYp5DQIc1_0;
	wire w_dff_A_IGLEGmrh9_0;
	wire w_dff_B_jvnGzxqi9_2;
	wire w_dff_B_VVqurd5k9_2;
	wire w_dff_B_mSkxwXQh3_2;
	wire w_dff_B_t3CuSTtI6_2;
	wire w_dff_B_AmzplG4U7_2;
	wire w_dff_A_9Oywq3Cy4_0;
	wire w_dff_A_qYC8OLbf3_0;
	wire w_dff_A_y5FkzdAj6_0;
	wire w_dff_A_MpICS6oG9_1;
	wire w_dff_A_i3PKVHDZ8_1;
	wire w_dff_A_QLE8tMgA9_1;
	wire w_dff_A_PWpSrhra2_1;
	wire w_dff_A_3iguwmxU7_1;
	wire w_dff_A_XHiXL1vT3_1;
	wire w_dff_A_7szbMaJP7_1;
	wire w_dff_A_nIaoEFj81_1;
	wire w_dff_A_Fn5wJJxq9_0;
	wire w_dff_A_yk1twS921_0;
	wire w_dff_A_r7uKwLKa2_0;
	wire w_dff_A_m7iU58na4_0;
	wire w_dff_A_D4DlJhkB5_0;
	wire w_dff_B_wbf1ntPr9_2;
	wire w_dff_B_bK0v1cy11_2;
	wire w_dff_B_NqZ5Jgx63_2;
	wire w_dff_B_DWRYHzfE4_2;
	wire w_dff_B_vSYbKYBY4_2;
	wire w_dff_A_FKtEcpHY6_0;
	wire w_dff_A_adsLzTVN6_0;
	wire w_dff_A_d7sPam9L9_0;
	wire w_dff_A_iHxyBWcY6_0;
	wire w_dff_A_5wssdGa09_0;
	wire w_dff_A_7xa6gGTi5_0;
	wire w_dff_A_QF3EaDNk1_0;
	wire w_dff_A_LWwWd2XP2_0;
	wire w_dff_A_nPHp5ejD7_1;
	wire w_dff_A_mKSXXTUt3_1;
	wire w_dff_A_GHQIdJ3A2_1;
	wire w_dff_B_1Dqoumz57_0;
	wire w_dff_B_cbdoMM8D3_0;
	wire w_dff_B_Uk8EdMHU4_0;
	wire w_dff_B_nGVCPjFW1_1;
	wire w_dff_B_sggIiMAn0_1;
	wire w_dff_B_zObk1IBb7_1;
	wire w_dff_A_Fy60x3P36_0;
	wire w_dff_A_Yi5W6JXN6_0;
	wire w_dff_A_soVg1WKJ3_0;
	wire w_dff_A_IQMaiIy48_0;
	wire w_dff_A_SBG7leFx0_0;
	wire w_dff_A_K04cbamz3_0;
	wire w_dff_A_W326EnfZ9_2;
	wire w_dff_A_99OEwyVj8_0;
	wire w_dff_A_TO0pI6pW4_0;
	wire w_dff_A_uVAAnEkd7_0;
	wire w_dff_A_TQqw1IkZ8_0;
	wire w_dff_A_mVDjpnBy0_0;
	wire w_dff_A_lDalHZ6U6_0;
	wire w_dff_A_rtpVrcs98_0;
	wire w_dff_A_gbQT9wQ18_0;
	wire w_dff_B_Cm1a5uJJ0_1;
	wire w_dff_B_BEEiQtjO1_1;
	wire w_dff_B_b1qlV9oy7_1;
	wire w_dff_B_lGP9RFp44_1;
	wire w_dff_B_OhC3PUo71_1;
	wire w_dff_B_gX41heb25_1;
	wire w_dff_B_1xpyi4966_1;
	wire w_dff_A_MbQKfbsk6_0;
	wire w_dff_A_rqzoA0Ia7_0;
	wire w_dff_A_yHkvwQj01_0;
	wire w_dff_A_2K2yrrM81_0;
	wire w_dff_A_nrNMB1Qw2_0;
	wire w_dff_A_UkW8ZDk14_0;
	wire w_dff_A_SEUXUfo07_0;
	wire w_dff_A_uMW9eypZ3_0;
	wire w_dff_A_FZXMCCaU2_0;
	wire w_dff_A_8D4StsrM8_0;
	wire w_dff_A_7ScH9M6S5_0;
	wire w_dff_A_zQPleNJo0_0;
	wire w_dff_A_mzmXnC9F9_0;
	wire w_dff_A_vDActhM91_0;
	wire w_dff_A_P2mQQYsi8_0;
	wire w_dff_A_hiserwzi4_0;
	wire w_dff_A_t1cFit3B7_0;
	wire w_dff_A_baWLntZs7_0;
	wire w_dff_A_8xi9B3wd0_0;
	wire w_dff_A_tA2X8DgX2_0;
	wire w_dff_A_pisgjtVx6_0;
	wire w_dff_A_FvT8uCGY0_0;
	wire w_dff_A_K44bNDl21_0;
	wire w_dff_A_SR1ejsZM8_0;
	wire w_dff_A_JYgXQKqk1_0;
	wire w_dff_A_Nz4sdyYA2_0;
	wire w_dff_A_GcwJnUIe9_0;
	wire w_dff_A_sNF0DQIE1_0;
	wire w_dff_A_EAGYtwR70_2;
	wire w_dff_A_1nWO7iXq1_0;
	wire w_dff_A_W0uqm6yX6_0;
	wire w_dff_A_JrjeQhYS0_0;
	wire w_dff_A_ieyc2s8R4_0;
	wire w_dff_A_Oy1yKkZC3_0;
	wire w_dff_A_iQYLfxpb5_0;
	wire w_dff_A_ZYoviDPY0_1;
	wire w_dff_A_FlQoilbD1_0;
	wire w_dff_A_SPW8OOyW2_0;
	wire w_dff_A_9hkp6sgQ4_0;
	wire w_dff_A_0YvkzvW76_0;
	wire w_dff_A_4PQy5beG8_0;
	wire w_dff_A_Cr2ZkKXQ4_0;
	wire w_dff_A_yt9M3IUb6_1;
	wire w_dff_A_pfh2nmvF3_0;
	wire w_dff_A_V7Khcg9C9_0;
	wire w_dff_A_7RPd38vW4_0;
	wire w_dff_A_58oV52wE8_0;
	wire w_dff_B_afx5LJw82_2;
	wire w_dff_A_oSmuBXq48_0;
	wire w_dff_A_UuzPBemQ3_0;
	wire w_dff_A_Nufseag98_0;
	wire w_dff_A_82RAgkJH2_0;
	wire w_dff_A_krz4KfgE3_0;
	wire w_dff_A_I7kKsBev3_0;
	wire w_dff_A_LYsOicH60_0;
	wire w_dff_A_GsuKMg6o3_0;
	wire w_dff_A_GEAeV8tI5_0;
	wire w_dff_A_0SWsR2jh0_2;
	wire w_dff_A_beQQhK370_0;
	wire w_dff_A_E34v5w1D8_0;
	wire w_dff_A_bH46gdET4_0;
	wire w_dff_A_XWRn0zpj8_0;
	wire w_dff_A_w0s2IWhd5_0;
	wire w_dff_A_s7ajoNiA4_0;
	wire w_dff_A_waCCqaoY2_2;
	wire w_dff_A_CZRt8b9D0_0;
	wire w_dff_A_nSpv3FJ57_0;
	wire w_dff_A_KDP78WSH1_0;
	wire w_dff_A_xpJgvIew4_0;
	wire w_dff_A_kLmahsAr0_0;
	wire w_dff_A_HuGCCWpH6_0;
	wire w_dff_A_irsMUWDd8_0;
	wire w_dff_A_KIvKVHvM3_0;
	wire w_dff_A_GYjoS2KM5_0;
	wire w_dff_A_ON2lZaPN2_0;
	wire w_dff_A_dZMPz4bJ0_2;
	wire w_dff_A_1JuT8rBx3_0;
	wire w_dff_A_XRbHuvV03_0;
	wire w_dff_A_ouUnLuhN5_0;
	wire w_dff_A_q1Qym2jm8_0;
	wire w_dff_A_ag0BdDFt3_0;
	wire w_dff_A_vBRpqx6P4_0;
	wire w_dff_A_AFfuu5bo6_1;
	wire w_dff_A_Jlef4EEs7_0;
	wire w_dff_A_0PV6cdnB5_0;
	wire w_dff_A_FOJ7HYgQ0_0;
	wire w_dff_A_8VPOe6SL6_0;
	wire w_dff_A_GtpHoEfs6_0;
	wire w_dff_A_nIt0Sw2C8_2;
	wire w_dff_A_oxqdqFdH8_0;
	wire w_dff_A_A0zQVHCd9_0;
	wire w_dff_A_HAJ8INlW8_0;
	wire w_dff_A_AFXSpOTL0_0;
	wire w_dff_A_gNpeiWC76_0;
	wire w_dff_A_X04574qT0_0;
	wire w_dff_A_bCzKI3Ty9_1;
	wire w_dff_A_iV4VKlYT5_1;
	wire w_dff_A_AQlHL5dX4_1;
	wire w_dff_A_3MH6jBP51_1;
	wire w_dff_A_gHkb2n0z4_1;
	wire w_dff_A_mbmiBSyX7_1;
	wire w_dff_A_VzTadzja5_2;
	wire w_dff_A_rrsSLf0g5_0;
	wire w_dff_A_lR29XX9a3_0;
	wire w_dff_A_dDBMv6kV5_0;
	wire w_dff_A_YICBIYUR5_0;
	wire w_dff_A_O8hs6JXi2_0;
	wire w_dff_A_A5gMHVGY8_0;
	wire w_dff_A_ABan4mVc1_1;
	wire w_dff_A_6tTDm9QE1_1;
	wire w_dff_A_p4a7zD0u7_1;
	wire w_dff_A_FiuEEm6L9_1;
	wire w_dff_A_TrwZZhQ47_1;
	wire w_dff_A_XnK8trYj6_2;
	wire w_dff_A_BdAAYCsi3_0;
	wire w_dff_A_MWyuzg3i9_0;
	wire w_dff_A_Bl61cQJR4_0;
	wire w_dff_A_DNklI1Sz2_0;
	wire w_dff_A_HIO2QXR52_0;
	wire w_dff_A_UEOo2iVB1_0;
	wire w_dff_A_rGuLBSJD8_0;
	wire w_dff_A_VmNbwtX40_0;
	wire w_dff_A_WSKhU4EA2_0;
	wire w_dff_A_Vr58FxO11_0;
	wire w_dff_A_5uny8MAX6_0;
	wire w_dff_A_kXDw8aob9_0;
	wire w_dff_A_jouY31xd5_0;
	wire w_dff_A_l0ipPEzk1_2;
	jnot g000(.din(w_G11gat_0[1]),.dout(n44),.clk(gclk));
	jand g001(.dina(w_G17gat_0[2]),.dinb(w_n44_0[1]),.dout(n45),.clk(gclk));
	jnot g002(.din(w_G76gat_0[1]),.dout(n46),.clk(gclk));
	jand g003(.dina(w_G82gat_0[2]),.dinb(w_n46_0[1]),.dout(n47),.clk(gclk));
	jcb g004(.dina(n47),.dinb(n45),.dout(n48));
	jnot g005(.din(w_G50gat_0[2]),.dout(n49),.clk(gclk));
	jand g006(.dina(w_G56gat_0[2]),.dinb(w_n49_0[1]),.dout(n50),.clk(gclk));
	jnot g007(.din(w_G89gat_0[2]),.dout(n51),.clk(gclk));
	jand g008(.dina(w_G95gat_0[2]),.dinb(w_n51_0[1]),.dout(n52),.clk(gclk));
	jcb g009(.dina(n52),.dinb(n50),.dout(n53));
	jnot g010(.din(w_G63gat_0[1]),.dout(n54),.clk(gclk));
	jand g011(.dina(w_G69gat_0[2]),.dinb(w_n54_0[1]),.dout(n55),.clk(gclk));
	jnot g012(.din(w_G37gat_0[1]),.dout(n56),.clk(gclk));
	jand g013(.dina(w_G43gat_0[2]),.dinb(n56),.dout(n57),.clk(gclk));
	jcb g014(.dina(w_n57_0[1]),.dinb(n55),.dout(n58));
	jcb g015(.dina(n58),.dinb(n53),.dout(n59));
	jnot g016(.din(G108gat),.dout(n60),.clk(gclk));
	jcb g017(.dina(w_n60_0[1]),.dinb(w_G102gat_0[1]),.dout(n61));
	jnot g018(.din(w_n61_0[1]),.dout(n62),.clk(gclk));
	jnot g019(.din(w_G24gat_0[2]),.dout(n63),.clk(gclk));
	jand g020(.dina(w_G30gat_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jnot g021(.din(w_G1gat_0[2]),.dout(n65),.clk(gclk));
	jand g022(.dina(w_G4gat_0[2]),.dinb(w_n65_0[1]),.dout(n66),.clk(gclk));
	jcb g023(.dina(n66),.dinb(n64),.dout(n67));
	jcb g024(.dina(n67),.dinb(n62),.dout(n68));
	jcb g025(.dina(n68),.dinb(n59),.dout(n69));
	jcb g026(.dina(n69),.dinb(w_n48_0[1]),.dout(G223gat_fa_));
	jnot g027(.din(w_G47gat_0[1]),.dout(n71),.clk(gclk));
	jnot g028(.din(w_n48_0[0]),.dout(n72),.clk(gclk));
	jnot g029(.din(w_G56gat_0[1]),.dout(n73),.clk(gclk));
	jcb g030(.dina(w_n73_0[1]),.dinb(w_G50gat_0[1]),.dout(n74));
	jnot g031(.din(w_G95gat_0[1]),.dout(n75),.clk(gclk));
	jcb g032(.dina(w_n75_0[1]),.dinb(w_G89gat_0[1]),.dout(n76));
	jand g033(.dina(n76),.dinb(n74),.dout(n77),.clk(gclk));
	jnot g034(.din(w_G69gat_0[1]),.dout(n78),.clk(gclk));
	jcb g035(.dina(n78),.dinb(w_G63gat_0[0]),.dout(n79));
	jnot g036(.din(w_G43gat_0[1]),.dout(n80),.clk(gclk));
	jcb g037(.dina(w_n80_0[1]),.dinb(w_G37gat_0[0]),.dout(n81));
	jand g038(.dina(w_n81_0[1]),.dinb(n79),.dout(n82),.clk(gclk));
	jand g039(.dina(n82),.dinb(n77),.dout(n83),.clk(gclk));
	jnot g040(.din(w_G30gat_0[1]),.dout(n84),.clk(gclk));
	jcb g041(.dina(w_n84_0[1]),.dinb(w_G24gat_0[1]),.dout(n85));
	jnot g042(.din(w_G4gat_0[1]),.dout(n86),.clk(gclk));
	jcb g043(.dina(w_n86_0[1]),.dinb(w_G1gat_0[1]),.dout(n87));
	jand g044(.dina(n87),.dinb(n85),.dout(n88),.clk(gclk));
	jand g045(.dina(n88),.dinb(w_n61_0[0]),.dout(n89),.clk(gclk));
	jand g046(.dina(n89),.dinb(n83),.dout(n90),.clk(gclk));
	jand g047(.dina(n90),.dinb(w_dff_B_1xpyi4966_1),.dout(n91),.clk(gclk));
	jxor g048(.dina(w_n91_3[1]),.dinb(w_n57_0[0]),.dout(n92),.clk(gclk));
	jand g049(.dina(n92),.dinb(w_G43gat_0[0]),.dout(n93),.clk(gclk));
	jand g050(.dina(w_n93_0[1]),.dinb(w_dff_B_gX41heb25_1),.dout(n94),.clk(gclk));
	jnot g051(.din(w_G112gat_0[1]),.dout(n95),.clk(gclk));
	jand g052(.dina(w_G223gat_3[1]),.dinb(w_G102gat_0[0]),.dout(n96),.clk(gclk));
	jcb g053(.dina(n96),.dinb(w_n60_0[0]),.dout(n97));
	jnot g054(.din(w_n97_0[1]),.dout(n98),.clk(gclk));
	jand g055(.dina(n98),.dinb(w_dff_B_zObk1IBb7_1),.dout(n99),.clk(gclk));
	jcb g056(.dina(w_dff_B_Uk8EdMHU4_0),.dinb(n94),.dout(n100));
	jnot g057(.din(w_G21gat_0[2]),.dout(n101),.clk(gclk));
	jcb g058(.dina(w_n91_3[0]),.dinb(w_n44_0[0]),.dout(n102));
	jand g059(.dina(n102),.dinb(w_G17gat_0[1]),.dout(n103),.clk(gclk));
	jand g060(.dina(n103),.dinb(w_n101_0[1]),.dout(n104),.clk(gclk));
	jnot g061(.din(w_G8gat_0[2]),.dout(n105),.clk(gclk));
	jcb g062(.dina(w_n91_2[2]),.dinb(w_n65_0[0]),.dout(n106));
	jand g063(.dina(n106),.dinb(w_G4gat_0[0]),.dout(n107),.clk(gclk));
	jand g064(.dina(n107),.dinb(w_n105_0[1]),.dout(n108),.clk(gclk));
	jcb g065(.dina(n108),.dinb(n104),.dout(n109));
	jnot g066(.din(w_G34gat_0[2]),.dout(n110),.clk(gclk));
	jcb g067(.dina(w_n91_2[1]),.dinb(w_n63_0[0]),.dout(n111));
	jand g068(.dina(n111),.dinb(w_G30gat_0[0]),.dout(n112),.clk(gclk));
	jand g069(.dina(w_n112_0[1]),.dinb(w_n110_0[1]),.dout(n113),.clk(gclk));
	jnot g070(.din(w_G86gat_0[2]),.dout(n114),.clk(gclk));
	jcb g071(.dina(w_n91_2[0]),.dinb(w_n46_0[0]),.dout(n115));
	jand g072(.dina(n115),.dinb(w_G82gat_0[1]),.dout(n116),.clk(gclk));
	jand g073(.dina(w_n116_0[1]),.dinb(w_n114_0[1]),.dout(n117),.clk(gclk));
	jcb g074(.dina(n117),.dinb(n113),.dout(n118));
	jcb g075(.dina(n118),.dinb(n109),.dout(n119));
	jnot g076(.din(w_G73gat_0[1]),.dout(n120),.clk(gclk));
	jcb g077(.dina(w_n91_1[2]),.dinb(w_n54_0[0]),.dout(n121));
	jand g078(.dina(n121),.dinb(w_G69gat_0[0]),.dout(n122),.clk(gclk));
	jand g079(.dina(w_n122_0[1]),.dinb(w_dff_B_YmnvNTO67_1),.dout(n123),.clk(gclk));
	jnot g080(.din(w_G99gat_0[2]),.dout(n124),.clk(gclk));
	jcb g081(.dina(w_n91_1[1]),.dinb(w_n51_0[0]),.dout(n125));
	jand g082(.dina(n125),.dinb(w_G95gat_0[0]),.dout(n126),.clk(gclk));
	jand g083(.dina(n126),.dinb(w_dff_B_yqZGaAPC1_1),.dout(n127),.clk(gclk));
	jnot g084(.din(w_G60gat_0[2]),.dout(n128),.clk(gclk));
	jcb g085(.dina(w_n91_1[0]),.dinb(w_n49_0[0]),.dout(n129));
	jand g086(.dina(n129),.dinb(w_G56gat_0[0]),.dout(n130),.clk(gclk));
	jand g087(.dina(w_n130_0[1]),.dinb(w_n128_0[1]),.dout(n131),.clk(gclk));
	jcb g088(.dina(n131),.dinb(n127),.dout(n132));
	jcb g089(.dina(n132),.dinb(w_n123_0[1]),.dout(n133));
	jcb g090(.dina(n133),.dinb(n119),.dout(n134));
	jcb g091(.dina(w_dff_B_elRkFYIP3_0),.dinb(w_n100_0[1]),.dout(G329gat_fa_));
	jand g092(.dina(w_G329gat_4),.dinb(w_G112gat_0[0]),.dout(n136),.clk(gclk));
	jcb g093(.dina(n136),.dinb(w_n97_0[0]),.dout(n137));
	jcb g094(.dina(w_n137_0[1]),.dinb(w_G115gat_0[1]),.dout(n138));
	jand g095(.dina(w_G223gat_3[0]),.dinb(w_G1gat_0[0]),.dout(n139),.clk(gclk));
	jcb g096(.dina(n139),.dinb(w_n86_0[0]),.dout(n140));
	jand g097(.dina(w_G329gat_3[2]),.dinb(w_G8gat_0[1]),.dout(n141),.clk(gclk));
	jcb g098(.dina(n141),.dinb(w_n140_0[1]),.dout(n142));
	jnot g099(.din(w_n100_0[0]),.dout(n143),.clk(gclk));
	jnot g100(.din(w_G17gat_0[0]),.dout(n144),.clk(gclk));
	jand g101(.dina(w_G223gat_2[2]),.dinb(w_G11gat_0[0]),.dout(n145),.clk(gclk));
	jcb g102(.dina(n145),.dinb(w_dff_B_J9UvRJ9I9_1),.dout(n146));
	jcb g103(.dina(w_n146_0[1]),.dinb(w_G21gat_0[1]),.dout(n147));
	jcb g104(.dina(w_n140_0[0]),.dinb(w_G8gat_0[0]),.dout(n148));
	jand g105(.dina(n148),.dinb(n147),.dout(n149),.clk(gclk));
	jand g106(.dina(w_G223gat_2[1]),.dinb(w_G24gat_0[0]),.dout(n150),.clk(gclk));
	jcb g107(.dina(n150),.dinb(w_n84_0[0]),.dout(n151));
	jcb g108(.dina(w_n151_0[1]),.dinb(w_G34gat_0[1]),.dout(n152));
	jnot g109(.din(w_G82gat_0[0]),.dout(n153),.clk(gclk));
	jand g110(.dina(w_G223gat_2[0]),.dinb(w_G76gat_0[0]),.dout(n154),.clk(gclk));
	jcb g111(.dina(n154),.dinb(w_dff_B_whZGNrI84_1),.dout(n155));
	jcb g112(.dina(w_n155_0[1]),.dinb(w_G86gat_0[1]),.dout(n156));
	jand g113(.dina(n156),.dinb(n152),.dout(n157),.clk(gclk));
	jand g114(.dina(n157),.dinb(n149),.dout(n158),.clk(gclk));
	jnot g115(.din(w_n123_0[0]),.dout(n159),.clk(gclk));
	jand g116(.dina(w_G223gat_1[2]),.dinb(w_G89gat_0[0]),.dout(n160),.clk(gclk));
	jcb g117(.dina(n160),.dinb(w_n75_0[0]),.dout(n161));
	jcb g118(.dina(w_n161_0[1]),.dinb(w_G99gat_0[1]),.dout(n162));
	jand g119(.dina(w_G223gat_1[1]),.dinb(w_G50gat_0[0]),.dout(n163),.clk(gclk));
	jcb g120(.dina(n163),.dinb(w_n73_0[0]),.dout(n164));
	jcb g121(.dina(w_n164_0[1]),.dinb(w_G60gat_0[1]),.dout(n165));
	jand g122(.dina(n165),.dinb(n162),.dout(n166),.clk(gclk));
	jand g123(.dina(w_dff_B_ekWoYZaN3_0),.dinb(n159),.dout(n167),.clk(gclk));
	jand g124(.dina(n167),.dinb(w_dff_B_xArl4hZ86_1),.dout(n168),.clk(gclk));
	jand g125(.dina(n168),.dinb(w_dff_B_qchdsOK64_1),.dout(n169),.clk(gclk));
	jand g126(.dina(w_n169_1[2]),.dinb(w_n105_0[0]),.dout(n170),.clk(gclk));
	jcb g127(.dina(n170),.dinb(w_G14gat_0[1]),.dout(n171));
	jcb g128(.dina(n171),.dinb(w_n142_0[1]),.dout(n172));
	jand g129(.dina(n172),.dinb(w_dff_B_PKRTrW9k6_1),.dout(n173),.clk(gclk));
	jand g130(.dina(w_G329gat_3[1]),.dinb(w_G99gat_0[0]),.dout(n174),.clk(gclk));
	jcb g131(.dina(n174),.dinb(w_n161_0[0]),.dout(n175));
	jcb g132(.dina(w_n175_0[1]),.dinb(w_G105gat_0[1]),.dout(n176));
	jnot g133(.din(w_n122_0[0]),.dout(n177),.clk(gclk));
	jand g134(.dina(w_G329gat_3[0]),.dinb(w_G73gat_0[0]),.dout(n178),.clk(gclk));
	jcb g135(.dina(n178),.dinb(w_dff_B_Yh1HPGxF1_1),.dout(n179));
	jcb g136(.dina(w_n179_0[1]),.dinb(w_G79gat_0[1]),.dout(n180));
	jand g137(.dina(n180),.dinb(n176),.dout(n181),.clk(gclk));
	jand g138(.dina(w_dff_B_HQsFRl0s9_0),.dinb(n173),.dout(n182),.clk(gclk));
	jnot g139(.din(w_n182_0[1]),.dout(n183),.clk(gclk));
	jnot g140(.din(w_G92gat_0[2]),.dout(n184),.clk(gclk));
	jcb g141(.dina(w_n169_1[1]),.dinb(w_n114_0[0]),.dout(n185));
	jand g142(.dina(n185),.dinb(w_n116_0[0]),.dout(n186),.clk(gclk));
	jand g143(.dina(n186),.dinb(w_dff_B_g91zQXQd2_1),.dout(n187),.clk(gclk));
	jand g144(.dina(w_G329gat_2[2]),.dinb(w_G47gat_0[0]),.dout(n188),.clk(gclk));
	jnot g145(.din(w_G53gat_0[1]),.dout(n189),.clk(gclk));
	jand g146(.dina(w_n93_0[0]),.dinb(w_n189_0[1]),.dout(n190),.clk(gclk));
	jnot g147(.din(n190),.dout(n191),.clk(gclk));
	jcb g148(.dina(n191),.dinb(w_n188_0[1]),.dout(n192));
	jnot g149(.din(w_n192_0[1]),.dout(n193),.clk(gclk));
	jcb g150(.dina(w_dff_B_U6hfzyHL4_0),.dinb(n187),.dout(n194));
	jnot g151(.din(w_G40gat_0[2]),.dout(n195),.clk(gclk));
	jcb g152(.dina(w_n169_1[0]),.dinb(w_n110_0[0]),.dout(n196));
	jand g153(.dina(n196),.dinb(w_n112_0[0]),.dout(n197),.clk(gclk));
	jand g154(.dina(w_n197_0[1]),.dinb(w_n195_0[1]),.dout(n198),.clk(gclk));
	jnot g155(.din(w_G66gat_0[1]),.dout(n199),.clk(gclk));
	jcb g156(.dina(w_n169_0[2]),.dinb(w_n128_0[0]),.dout(n200));
	jand g157(.dina(n200),.dinb(w_n130_0[0]),.dout(n201),.clk(gclk));
	jand g158(.dina(w_n201_0[1]),.dinb(w_dff_B_MJYhPC8g8_1),.dout(n202),.clk(gclk));
	jcb g159(.dina(w_n202_0[1]),.dinb(n198),.dout(n203));
	jcb g160(.dina(n203),.dinb(n194),.dout(n204));
	jand g161(.dina(w_n169_0[1]),.dinb(w_n101_0[0]),.dout(n205),.clk(gclk));
	jand g162(.dina(w_G329gat_2[1]),.dinb(w_G21gat_0[0]),.dout(n206),.clk(gclk));
	jcb g163(.dina(n206),.dinb(w_n146_0[0]),.dout(n207));
	jcb g164(.dina(w_n207_0[1]),.dinb(n205),.dout(n208));
	jcb g165(.dina(n208),.dinb(w_G27gat_0[1]),.dout(n209));
	jnot g166(.din(w_n209_0[1]),.dout(n210),.clk(gclk));
	jcb g167(.dina(n210),.dinb(n204),.dout(n211));
	jcb g168(.dina(w_dff_B_xtkQa4946_0),.dinb(n183),.dout(G370gat_fa_));
	jand g169(.dina(w_G370gat_2),.dinb(w_G14gat_0[0]),.dout(n213),.clk(gclk));
	jcb g170(.dina(n213),.dinb(w_n142_0[0]),.dout(n214));
	jnot g171(.din(w_n179_0[0]),.dout(n215),.clk(gclk));
	jnot g172(.din(w_G79gat_0[0]),.dout(n216),.clk(gclk));
	jand g173(.dina(w_G329gat_2[0]),.dinb(w_G86gat_0[0]),.dout(n217),.clk(gclk));
	jcb g174(.dina(n217),.dinb(w_n155_0[0]),.dout(n218));
	jcb g175(.dina(w_n218_0[1]),.dinb(w_G92gat_0[1]),.dout(n219));
	jand g176(.dina(w_n192_0[0]),.dinb(n219),.dout(n220),.clk(gclk));
	jand g177(.dina(w_G329gat_1[2]),.dinb(w_G34gat_0[0]),.dout(n221),.clk(gclk));
	jcb g178(.dina(n221),.dinb(w_n151_0[0]),.dout(n222));
	jcb g179(.dina(w_n222_0[1]),.dinb(w_G40gat_0[1]),.dout(n223));
	jand g180(.dina(w_G329gat_1[1]),.dinb(w_G60gat_0[0]),.dout(n224),.clk(gclk));
	jcb g181(.dina(n224),.dinb(w_n164_0[0]),.dout(n225));
	jcb g182(.dina(w_n225_0[1]),.dinb(w_G66gat_0[0]),.dout(n226));
	jand g183(.dina(w_n226_0[1]),.dinb(n223),.dout(n227),.clk(gclk));
	jand g184(.dina(n227),.dinb(n220),.dout(n228),.clk(gclk));
	jand g185(.dina(w_n209_0[0]),.dinb(w_dff_B_YG4D7ggH7_1),.dout(n229),.clk(gclk));
	jand g186(.dina(w_dff_B_KD1KIA7h3_0),.dinb(w_n182_0[0]),.dout(n230),.clk(gclk));
	jcb g187(.dina(w_n230_2[2]),.dinb(w_dff_B_EAwqKOMd2_1),.dout(n231));
	jand g188(.dina(n231),.dinb(w_dff_B_fb5mko2J9_1),.dout(n232),.clk(gclk));
	jand g189(.dina(w_G370gat_1[2]),.dinb(w_G92gat_0[0]),.dout(n233),.clk(gclk));
	jcb g190(.dina(n233),.dinb(w_n218_0[0]),.dout(n234));
	jnot g191(.din(w_n234_0[1]),.dout(n235),.clk(gclk));
	jcb g192(.dina(w_n235_0[1]),.dinb(w_n232_0[1]),.dout(n236));
	jnot g193(.din(w_n207_0[0]),.dout(n237),.clk(gclk));
	jnot g194(.din(w_G27gat_0[0]),.dout(n238),.clk(gclk));
	jcb g195(.dina(w_n230_2[1]),.dinb(w_dff_B_9PVZRrRo0_1),.dout(n239));
	jand g196(.dina(n239),.dinb(w_dff_B_lBrJComX7_1),.dout(n240),.clk(gclk));
	jcb g197(.dina(w_n230_2[0]),.dinb(w_n195_0[0]),.dout(n241));
	jand g198(.dina(n241),.dinb(w_n197_0[0]),.dout(n242),.clk(gclk));
	jcb g199(.dina(n242),.dinb(w_n240_0[1]),.dout(n243));
	jcb g200(.dina(w_n230_1[2]),.dinb(w_n189_0[0]),.dout(n244));
	jand g201(.dina(w_G223gat_1[0]),.dinb(w_n81_0[0]),.dout(n245),.clk(gclk));
	jcb g202(.dina(n245),.dinb(w_n80_0[0]),.dout(n246));
	jcb g203(.dina(w_dff_B_LZvlM0IF3_0),.dinb(w_n188_0[0]),.dout(n247));
	jnot g204(.din(w_n247_0[1]),.dout(n248),.clk(gclk));
	jand g205(.dina(w_dff_B_yHQjgJuJ2_0),.dinb(n244),.dout(n249),.clk(gclk));
	jand g206(.dina(w_n230_1[1]),.dinb(w_n201_0[0]),.dout(n250),.clk(gclk));
	jcb g207(.dina(n250),.dinb(w_n202_0[0]),.dout(n251));
	jcb g208(.dina(n251),.dinb(w_n249_0[1]),.dout(n252));
	jcb g209(.dina(n252),.dinb(w_n243_0[1]),.dout(G430gat_fa_));
	jnot g210(.din(w_n175_0[0]),.dout(n254),.clk(gclk));
	jnot g211(.din(w_G105gat_0[0]),.dout(n255),.clk(gclk));
	jcb g212(.dina(w_n230_1[0]),.dinb(w_dff_B_YKhgEew84_1),.dout(n256));
	jand g213(.dina(n256),.dinb(w_dff_B_qM6LeDhA0_1),.dout(n257),.clk(gclk));
	jnot g214(.din(w_n137_0[0]),.dout(n258),.clk(gclk));
	jnot g215(.din(w_G115gat_0[0]),.dout(n259),.clk(gclk));
	jcb g216(.dina(w_n230_0[2]),.dinb(w_dff_B_BdTi0qlL0_1),.dout(n260));
	jand g217(.dina(n260),.dinb(w_dff_B_ygjXYEtf8_1),.dout(n261),.clk(gclk));
	jcb g218(.dina(n261),.dinb(w_n257_0[1]),.dout(n262));
	jcb g219(.dina(n262),.dinb(w_G430gat_0),.dout(n263));
	jcb g220(.dina(w_dff_B_zc14q3Ww4_0),.dinb(n236),.dout(n264));
	jand g221(.dina(n264),.dinb(w_dff_B_e5alEDkm0_1),.dout(G421gat),.clk(gclk));
	jand g222(.dina(w_G370gat_1[1]),.dinb(w_G53gat_0[0]),.dout(n266),.clk(gclk));
	jcb g223(.dina(w_n247_0[0]),.dinb(n266),.dout(n267));
	jcb g224(.dina(w_G370gat_1[0]),.dinb(w_n225_0[0]),.dout(n268));
	jand g225(.dina(n268),.dinb(w_n226_0[0]),.dout(n269),.clk(gclk));
	jand g226(.dina(n269),.dinb(n267),.dout(n270),.clk(gclk));
	jand g227(.dina(w_G370gat_0[2]),.dinb(w_G40gat_0[0]),.dout(n271),.clk(gclk));
	jcb g228(.dina(n271),.dinb(w_n222_0[0]),.dout(n272));
	jand g229(.dina(w_n272_0[1]),.dinb(w_n232_0[0]),.dout(n273),.clk(gclk));
	jand g230(.dina(n273),.dinb(w_n270_0[1]),.dout(n274),.clk(gclk));
	jand g231(.dina(w_n270_0[0]),.dinb(w_n235_0[0]),.dout(n275),.clk(gclk));
	jcb g232(.dina(n275),.dinb(w_n243_0[0]),.dout(n276));
	jcb g233(.dina(n276),.dinb(w_n274_0[1]),.dout(G431gat));
	jand g234(.dina(w_n257_0[0]),.dinb(w_n234_0[0]),.dout(n278),.clk(gclk));
	jcb g235(.dina(n278),.dinb(w_n249_0[0]),.dout(n279));
	jand g236(.dina(n279),.dinb(w_n272_0[0]),.dout(n280),.clk(gclk));
	jcb g237(.dina(w_n274_0[0]),.dinb(w_n240_0[0]),.dout(n281));
	jcb g238(.dina(n281),.dinb(n280),.dout(G432gat));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_iQYLfxpb5_0),.doutb(w_dff_A_ZYoviDPY0_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_dff_A_sNF0DQIE1_0),.doutb(w_G4gat_0[1]),.doutc(w_dff_A_EAGYtwR70_2),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_y5FkzdAj6_0),.doutb(w_dff_A_nIaoEFj81_1),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl jspl_w_G11gat_0(.douta(w_dff_A_UEOo2iVB1_0),.doutb(w_G11gat_0[1]),.din(G11gat));
	jspl jspl_w_G14gat_0(.douta(w_dff_A_8pYhuuVD5_0),.doutb(w_G14gat_0[1]),.din(w_dff_B_iw6PA2gg1_2));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_dff_A_TrwZZhQ47_1),.doutc(w_dff_A_XnK8trYj6_2),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_dff_A_LWwWd2XP2_0),.doutb(w_dff_A_GHQIdJ3A2_1),.doutc(w_G21gat_0[2]),.din(G21gat));
	jspl3 jspl3_w_G24gat_0(.douta(w_dff_A_Cr2ZkKXQ4_0),.doutb(w_dff_A_yt9M3IUb6_1),.doutc(w_G24gat_0[2]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_G27gat_0[0]),.doutb(w_dff_A_vyQkkCnx5_1),.din(G27gat));
	jspl3 jspl3_w_G30gat_0(.douta(w_dff_A_jouY31xd5_0),.doutb(w_G30gat_0[1]),.doutc(w_dff_A_l0ipPEzk1_2),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_dff_A_JCeut76T7_0),.doutb(w_dff_A_tqGg37gq2_1),.doutc(w_G34gat_0[2]),.din(G34gat));
	jspl jspl_w_G37gat_0(.douta(w_dff_A_beQQhK370_0),.doutb(w_G37gat_0[1]),.din(G37gat));
	jspl3 jspl3_w_G40gat_0(.douta(w_dff_A_yS8gKoul0_0),.doutb(w_dff_A_tYJmetl42_1),.doutc(w_G40gat_0[2]),.din(G40gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_dff_A_GEAeV8tI5_0),.doutb(w_G43gat_0[1]),.doutc(w_dff_A_0SWsR2jh0_2),.din(G43gat));
	jspl jspl_w_G47gat_0(.douta(w_dff_A_t1cFit3B7_0),.doutb(w_G47gat_0[1]),.din(G47gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_dff_A_X04574qT0_0),.doutb(w_dff_A_bCzKI3Ty9_1),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_dff_A_BerntqP88_0),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_dff_A_GtpHoEfs6_0),.doutb(w_G56gat_0[1]),.doutc(w_dff_A_nIt0Sw2C8_2),.din(G56gat));
	jspl3 jspl3_w_G60gat_0(.douta(w_dff_A_2IOI8oZH0_0),.doutb(w_dff_A_8VHJ7YhU7_1),.doutc(w_G60gat_0[2]),.din(G60gat));
	jspl jspl_w_G63gat_0(.douta(w_dff_A_kLmahsAr0_0),.doutb(w_G63gat_0[1]),.din(G63gat));
	jspl jspl_w_G66gat_0(.douta(w_dff_A_dR0YlQd23_0),.doutb(w_G66gat_0[1]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_dff_A_s7ajoNiA4_0),.doutb(w_G69gat_0[1]),.doutc(w_dff_A_waCCqaoY2_2),.din(G69gat));
	jspl jspl_w_G73gat_0(.douta(w_dff_A_uC2MoJHC9_0),.doutb(w_G73gat_0[1]),.din(G73gat));
	jspl jspl_w_G76gat_0(.douta(w_dff_A_A5gMHVGY8_0),.doutb(w_G76gat_0[1]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_G79gat_0[0]),.doutb(w_dff_A_KLXF1nLE7_1),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_G82gat_0[0]),.doutb(w_dff_A_mbmiBSyX7_1),.doutc(w_dff_A_VzTadzja5_2),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_dff_A_CNjBBjIk4_0),.doutb(w_dff_A_jIh8pKnM9_1),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G89gat_0(.douta(w_dff_A_vBRpqx6P4_0),.doutb(w_dff_A_AFfuu5bo6_1),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_LKzdN1yI2_0),.doutb(w_dff_A_61v04UO43_1),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_dff_A_ON2lZaPN2_0),.doutb(w_G95gat_0[1]),.doutc(w_dff_A_dZMPz4bJ0_2),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_vyxp6Eid2_0),.doutb(w_dff_A_tRoBYtPN0_1),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl jspl_w_G102gat_0(.douta(w_dff_A_58oV52wE8_0),.doutb(w_G102gat_0[1]),.din(w_dff_B_afx5LJw82_2));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_dff_A_jkf4lP8S1_1),.din(G105gat));
	jspl jspl_w_G112gat_0(.douta(w_dff_A_gbQT9wQ18_0),.doutb(w_G112gat_0[1]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_G115gat_0[0]),.doutb(w_dff_A_eRHnONse6_1),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(w_dff_A_W326EnfZ9_2),.din(w_G223gat_0[2]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl jspl_w_G329gat_4(.douta(w_G329gat_4),.doutb(w_dff_A_mUeoM9Ob8_1),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_G370gat_1[2]),.din(w_G370gat_0[0]));
	jspl jspl_w_G370gat_2(.douta(w_G370gat_2),.doutb(w_dff_A_8GoXyrJa8_1),.din(w_G370gat_0[1]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(w_dff_A_Na4phgtn5_1),.din(G430gat_fa_));
	jspl jspl_w_n44_0(.douta(w_dff_A_DNklI1Sz2_0),.doutb(w_n44_0[1]),.din(n44));
	jspl jspl_w_n46_0(.douta(w_dff_A_YICBIYUR5_0),.doutb(w_n46_0[1]),.din(n46));
	jspl jspl_w_n48_0(.douta(w_n48_0[0]),.doutb(w_n48_0[1]),.din(n48));
	jspl jspl_w_n49_0(.douta(w_dff_A_AFXSpOTL0_0),.doutb(w_n49_0[1]),.din(n49));
	jspl jspl_w_n51_0(.douta(w_dff_A_q1Qym2jm8_0),.doutb(w_n51_0[1]),.din(n51));
	jspl jspl_w_n54_0(.douta(w_dff_A_xpJgvIew4_0),.doutb(w_n54_0[1]),.din(n54));
	jspl jspl_w_n57_0(.douta(w_dff_A_Nufseag98_0),.doutb(w_n57_0[1]),.din(n57));
	jspl jspl_w_n60_0(.douta(w_dff_A_7RPd38vW4_0),.doutb(w_n60_0[1]),.din(n60));
	jspl jspl_w_n61_0(.douta(w_dff_A_pfh2nmvF3_0),.doutb(w_n61_0[1]),.din(n61));
	jspl jspl_w_n63_0(.douta(w_dff_A_0YvkzvW76_0),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n65_0(.douta(w_dff_A_ieyc2s8R4_0),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n73_0(.douta(w_dff_A_FZXMCCaU2_0),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n75_0(.douta(w_dff_A_SEUXUfo07_0),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n80_0(.douta(w_dff_A_nrNMB1Qw2_0),.doutb(w_n80_0[1]),.din(n80));
	jspl jspl_w_n81_0(.douta(w_dff_A_yHkvwQj01_0),.doutb(w_n81_0[1]),.din(n81));
	jspl jspl_w_n84_0(.douta(w_dff_A_VmNbwtX40_0),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_dff_A_rqzoA0Ia7_0),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.doutc(w_n91_0[2]),.din(n91));
	jspl3 jspl3_w_n91_1(.douta(w_n91_1[0]),.doutb(w_n91_1[1]),.doutc(w_n91_1[2]),.din(w_n91_0[0]));
	jspl3 jspl3_w_n91_2(.douta(w_n91_2[0]),.doutb(w_n91_2[1]),.doutc(w_n91_2[2]),.din(w_n91_0[1]));
	jspl jspl_w_n91_3(.douta(w_n91_3[0]),.doutb(w_n91_3[1]),.din(w_n91_0[2]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n97_0(.douta(w_dff_A_K04cbamz3_0),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n100_0(.douta(w_n100_0[0]),.doutb(w_n100_0[1]),.din(n100));
	jspl jspl_w_n101_0(.douta(w_dff_A_D4DlJhkB5_0),.doutb(w_n101_0[1]),.din(w_dff_B_vSYbKYBY4_2));
	jspl jspl_w_n105_0(.douta(w_dff_A_IGLEGmrh9_0),.doutb(w_n105_0[1]),.din(w_dff_B_AmzplG4U7_2));
	jspl jspl_w_n110_0(.douta(w_dff_A_TYl7dF2w3_0),.doutb(w_n110_0[1]),.din(w_dff_B_HmDgpTZ25_2));
	jspl jspl_w_n112_0(.douta(w_dff_A_kRjQN2Aa7_0),.doutb(w_n112_0[1]),.din(n112));
	jspl jspl_w_n114_0(.douta(w_dff_A_OUBJK5dB4_0),.doutb(w_n114_0[1]),.din(w_dff_B_GZI4eWWi3_2));
	jspl jspl_w_n116_0(.douta(w_dff_A_lrvoPlfa9_0),.doutb(w_n116_0[1]),.din(n116));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.din(n122));
	jspl jspl_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n128_0(.douta(w_dff_A_5Rh6wsVC1_0),.doutb(w_n128_0[1]),.din(w_dff_B_Zq05Emy40_2));
	jspl jspl_w_n130_0(.douta(w_dff_A_iJcbkrHa8_0),.doutb(w_n130_0[1]),.din(n130));
	jspl jspl_w_n137_0(.douta(w_n137_0[0]),.doutb(w_n137_0[1]),.din(n137));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_dff_A_XaNgq4Wh4_1),.din(n140));
	jspl jspl_w_n142_0(.douta(w_dff_A_7MulR8yy0_0),.doutb(w_n142_0[1]),.din(w_dff_B_WR30poUH6_2));
	jspl jspl_w_n146_0(.douta(w_dff_A_gM7zOEJQ0_0),.doutb(w_n146_0[1]),.din(n146));
	jspl jspl_w_n151_0(.douta(w_dff_A_K44bNDl21_0),.doutb(w_n151_0[1]),.din(n151));
	jspl jspl_w_n155_0(.douta(w_dff_A_F5CDsX0C8_0),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n161_0(.douta(w_dff_A_VdyfJxk62_0),.doutb(w_n161_0[1]),.din(n161));
	jspl jspl_w_n164_0(.douta(w_dff_A_rOnrJ9g02_0),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.doutc(w_n169_0[2]),.din(n169));
	jspl3 jspl3_w_n169_1(.douta(w_n169_1[0]),.doutb(w_n169_1[1]),.doutc(w_n169_1[2]),.din(w_n169_0[0]));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n179_0(.douta(w_n179_0[0]),.doutb(w_n179_0[1]),.din(n179));
	jspl jspl_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.din(n182));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_dff_A_Oiq5S9mx3_0),.doutb(w_n189_0[1]),.din(w_dff_B_oOjS4uHz8_2));
	jspl jspl_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.din(n192));
	jspl jspl_w_n195_0(.douta(w_dff_A_6TmgDA501_0),.doutb(w_n195_0[1]),.din(w_dff_B_jOeKJE9G9_2));
	jspl jspl_w_n197_0(.douta(w_dff_A_E3aw4bMf4_0),.doutb(w_n197_0[1]),.din(n197));
	jspl jspl_w_n201_0(.douta(w_dff_A_ZIdL7NhX7_0),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n202_0(.douta(w_dff_A_KP6Pf0ls0_0),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_dff_A_xy0oMfl79_1),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.din(n209));
	jspl jspl_w_n218_0(.douta(w_dff_A_mujE1H1o5_0),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n222_0(.douta(w_dff_A_SVFC7uqp2_0),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n225_0(.douta(w_dff_A_PwgyT2Fz5_0),.doutb(w_n225_0[1]),.din(n225));
	jspl jspl_w_n226_0(.douta(w_dff_A_8AbjdZxs4_0),.doutb(w_n226_0[1]),.din(n226));
	jspl3 jspl3_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.doutc(w_n230_0[2]),.din(n230));
	jspl3 jspl3_w_n230_1(.douta(w_n230_1[0]),.doutb(w_n230_1[1]),.doutc(w_n230_1[2]),.din(w_n230_0[0]));
	jspl3 jspl3_w_n230_2(.douta(w_n230_2[0]),.doutb(w_n230_2[1]),.doutc(w_n230_2[2]),.din(w_n230_0[1]));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_dff_A_cqO6S9JU5_1),.din(n232));
	jspl jspl_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.din(n234));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_n235_0[1]),.din(n235));
	jspl jspl_w_n240_0(.douta(w_dff_A_iVlygmfK3_0),.doutb(w_n240_0[1]),.din(n240));
	jspl jspl_w_n243_0(.douta(w_dff_A_jj7v4i1G9_0),.doutb(w_n243_0[1]),.din(n243));
	jspl jspl_w_n247_0(.douta(w_dff_A_ShDyOuw69_0),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_dff_A_GE2OFhcu2_0),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.din(n270));
	jspl jspl_w_n272_0(.douta(w_dff_A_94zoQHuY9_0),.doutb(w_n272_0[1]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jdff dff_B_e5alEDkm0_1(.din(n214),.dout(w_dff_B_e5alEDkm0_1),.clk(gclk));
	jdff dff_B_zc14q3Ww4_0(.din(n263),.dout(w_dff_B_zc14q3Ww4_0),.clk(gclk));
	jdff dff_B_Rr9P4l8Q2_1(.din(n258),.dout(w_dff_B_Rr9P4l8Q2_1),.clk(gclk));
	jdff dff_B_EKguxQvI2_1(.din(w_dff_B_Rr9P4l8Q2_1),.dout(w_dff_B_EKguxQvI2_1),.clk(gclk));
	jdff dff_B_0Q6AgxcI3_1(.din(w_dff_B_EKguxQvI2_1),.dout(w_dff_B_0Q6AgxcI3_1),.clk(gclk));
	jdff dff_B_hLwXVtbl0_1(.din(w_dff_B_0Q6AgxcI3_1),.dout(w_dff_B_hLwXVtbl0_1),.clk(gclk));
	jdff dff_B_ygjXYEtf8_1(.din(w_dff_B_hLwXVtbl0_1),.dout(w_dff_B_ygjXYEtf8_1),.clk(gclk));
	jdff dff_B_0XZKHc2f5_1(.din(n259),.dout(w_dff_B_0XZKHc2f5_1),.clk(gclk));
	jdff dff_B_smGAGvqp0_1(.din(w_dff_B_0XZKHc2f5_1),.dout(w_dff_B_smGAGvqp0_1),.clk(gclk));
	jdff dff_B_JeATEhhI8_1(.din(w_dff_B_smGAGvqp0_1),.dout(w_dff_B_JeATEhhI8_1),.clk(gclk));
	jdff dff_B_CdWLwGFg8_1(.din(w_dff_B_JeATEhhI8_1),.dout(w_dff_B_CdWLwGFg8_1),.clk(gclk));
	jdff dff_B_LYVkKKH96_1(.din(w_dff_B_CdWLwGFg8_1),.dout(w_dff_B_LYVkKKH96_1),.clk(gclk));
	jdff dff_B_lq94nuYA8_1(.din(w_dff_B_LYVkKKH96_1),.dout(w_dff_B_lq94nuYA8_1),.clk(gclk));
	jdff dff_B_0hwomlzi0_1(.din(w_dff_B_lq94nuYA8_1),.dout(w_dff_B_0hwomlzi0_1),.clk(gclk));
	jdff dff_B_dhJsoA2W5_1(.din(w_dff_B_0hwomlzi0_1),.dout(w_dff_B_dhJsoA2W5_1),.clk(gclk));
	jdff dff_B_sEHsiY7T2_1(.din(w_dff_B_dhJsoA2W5_1),.dout(w_dff_B_sEHsiY7T2_1),.clk(gclk));
	jdff dff_B_n4zCBecB6_1(.din(w_dff_B_sEHsiY7T2_1),.dout(w_dff_B_n4zCBecB6_1),.clk(gclk));
	jdff dff_B_mQ8whF5V8_1(.din(w_dff_B_n4zCBecB6_1),.dout(w_dff_B_mQ8whF5V8_1),.clk(gclk));
	jdff dff_B_RnLAEkNG5_1(.din(w_dff_B_mQ8whF5V8_1),.dout(w_dff_B_RnLAEkNG5_1),.clk(gclk));
	jdff dff_B_KwMrbmoV3_1(.din(w_dff_B_RnLAEkNG5_1),.dout(w_dff_B_KwMrbmoV3_1),.clk(gclk));
	jdff dff_B_BdTi0qlL0_1(.din(w_dff_B_KwMrbmoV3_1),.dout(w_dff_B_BdTi0qlL0_1),.clk(gclk));
	jdff dff_A_8GoXyrJa8_1(.dout(G370gat),.din(w_dff_A_8GoXyrJa8_1),.clk(gclk));
	jdff dff_A_Na4phgtn5_1(.dout(G430gat),.din(w_dff_A_Na4phgtn5_1),.clk(gclk));
	jdff dff_A_N54RAZRq8_0(.dout(w_n243_0[0]),.din(w_dff_A_N54RAZRq8_0),.clk(gclk));
	jdff dff_A_jj7v4i1G9_0(.dout(w_dff_A_N54RAZRq8_0),.din(w_dff_A_jj7v4i1G9_0),.clk(gclk));
	jdff dff_A_cqO6S9JU5_1(.dout(w_n232_0[1]),.din(w_dff_A_cqO6S9JU5_1),.clk(gclk));
	jdff dff_B_rayBSws80_1(.din(n215),.dout(w_dff_B_rayBSws80_1),.clk(gclk));
	jdff dff_B_WkD10pJW1_1(.din(w_dff_B_rayBSws80_1),.dout(w_dff_B_WkD10pJW1_1),.clk(gclk));
	jdff dff_B_yz9qbQe82_1(.din(w_dff_B_WkD10pJW1_1),.dout(w_dff_B_yz9qbQe82_1),.clk(gclk));
	jdff dff_B_SIWxHZAL7_1(.din(w_dff_B_yz9qbQe82_1),.dout(w_dff_B_SIWxHZAL7_1),.clk(gclk));
	jdff dff_B_fb5mko2J9_1(.din(w_dff_B_SIWxHZAL7_1),.dout(w_dff_B_fb5mko2J9_1),.clk(gclk));
	jdff dff_B_MHJ9DvKA6_1(.din(n216),.dout(w_dff_B_MHJ9DvKA6_1),.clk(gclk));
	jdff dff_B_KChWfxvy8_1(.din(w_dff_B_MHJ9DvKA6_1),.dout(w_dff_B_KChWfxvy8_1),.clk(gclk));
	jdff dff_B_EIxEtQhj8_1(.din(w_dff_B_KChWfxvy8_1),.dout(w_dff_B_EIxEtQhj8_1),.clk(gclk));
	jdff dff_B_p1F4fnSJ6_1(.din(w_dff_B_EIxEtQhj8_1),.dout(w_dff_B_p1F4fnSJ6_1),.clk(gclk));
	jdff dff_B_Xvud4s3Z8_1(.din(w_dff_B_p1F4fnSJ6_1),.dout(w_dff_B_Xvud4s3Z8_1),.clk(gclk));
	jdff dff_B_uREUa1EU9_1(.din(w_dff_B_Xvud4s3Z8_1),.dout(w_dff_B_uREUa1EU9_1),.clk(gclk));
	jdff dff_B_XE8vKwi15_1(.din(w_dff_B_uREUa1EU9_1),.dout(w_dff_B_XE8vKwi15_1),.clk(gclk));
	jdff dff_B_0cZ7qe8m5_1(.din(w_dff_B_XE8vKwi15_1),.dout(w_dff_B_0cZ7qe8m5_1),.clk(gclk));
	jdff dff_B_K8ntdtot9_1(.din(w_dff_B_0cZ7qe8m5_1),.dout(w_dff_B_K8ntdtot9_1),.clk(gclk));
	jdff dff_B_jkiZY0gw8_1(.din(w_dff_B_K8ntdtot9_1),.dout(w_dff_B_jkiZY0gw8_1),.clk(gclk));
	jdff dff_B_frvgF7bQ7_1(.din(w_dff_B_jkiZY0gw8_1),.dout(w_dff_B_frvgF7bQ7_1),.clk(gclk));
	jdff dff_B_AKIuBdTm8_1(.din(w_dff_B_frvgF7bQ7_1),.dout(w_dff_B_AKIuBdTm8_1),.clk(gclk));
	jdff dff_B_FdGKqCue2_1(.din(w_dff_B_AKIuBdTm8_1),.dout(w_dff_B_FdGKqCue2_1),.clk(gclk));
	jdff dff_B_EAwqKOMd2_1(.din(w_dff_B_FdGKqCue2_1),.dout(w_dff_B_EAwqKOMd2_1),.clk(gclk));
	jdff dff_A_3iAJhNi49_0(.dout(w_n240_0[0]),.din(w_dff_A_3iAJhNi49_0),.clk(gclk));
	jdff dff_A_iVlygmfK3_0(.dout(w_dff_A_3iAJhNi49_0),.din(w_dff_A_iVlygmfK3_0),.clk(gclk));
	jdff dff_B_V5i3A9gs7_1(.din(n237),.dout(w_dff_B_V5i3A9gs7_1),.clk(gclk));
	jdff dff_B_XG3Vyga20_1(.din(w_dff_B_V5i3A9gs7_1),.dout(w_dff_B_XG3Vyga20_1),.clk(gclk));
	jdff dff_B_IkpjPyrw7_1(.din(w_dff_B_XG3Vyga20_1),.dout(w_dff_B_IkpjPyrw7_1),.clk(gclk));
	jdff dff_B_ingOgbsg1_1(.din(w_dff_B_IkpjPyrw7_1),.dout(w_dff_B_ingOgbsg1_1),.clk(gclk));
	jdff dff_B_lBrJComX7_1(.din(w_dff_B_ingOgbsg1_1),.dout(w_dff_B_lBrJComX7_1),.clk(gclk));
	jdff dff_B_qnaFo5Ee6_1(.din(n238),.dout(w_dff_B_qnaFo5Ee6_1),.clk(gclk));
	jdff dff_B_YMdibU7c0_1(.din(w_dff_B_qnaFo5Ee6_1),.dout(w_dff_B_YMdibU7c0_1),.clk(gclk));
	jdff dff_B_LQCtmshq1_1(.din(w_dff_B_YMdibU7c0_1),.dout(w_dff_B_LQCtmshq1_1),.clk(gclk));
	jdff dff_B_Xpm6vzuh9_1(.din(w_dff_B_LQCtmshq1_1),.dout(w_dff_B_Xpm6vzuh9_1),.clk(gclk));
	jdff dff_B_GuTKXBH69_1(.din(w_dff_B_Xpm6vzuh9_1),.dout(w_dff_B_GuTKXBH69_1),.clk(gclk));
	jdff dff_B_1fx2u2iR2_1(.din(w_dff_B_GuTKXBH69_1),.dout(w_dff_B_1fx2u2iR2_1),.clk(gclk));
	jdff dff_B_RuyKfXgE7_1(.din(w_dff_B_1fx2u2iR2_1),.dout(w_dff_B_RuyKfXgE7_1),.clk(gclk));
	jdff dff_B_cdGn0N916_1(.din(w_dff_B_RuyKfXgE7_1),.dout(w_dff_B_cdGn0N916_1),.clk(gclk));
	jdff dff_B_iPGAxZSf9_1(.din(w_dff_B_cdGn0N916_1),.dout(w_dff_B_iPGAxZSf9_1),.clk(gclk));
	jdff dff_B_Ii23Vlge6_1(.din(w_dff_B_iPGAxZSf9_1),.dout(w_dff_B_Ii23Vlge6_1),.clk(gclk));
	jdff dff_B_Ue4UedO57_1(.din(w_dff_B_Ii23Vlge6_1),.dout(w_dff_B_Ue4UedO57_1),.clk(gclk));
	jdff dff_B_AfHVPBWM0_1(.din(w_dff_B_Ue4UedO57_1),.dout(w_dff_B_AfHVPBWM0_1),.clk(gclk));
	jdff dff_B_qMH1XlYV7_1(.din(w_dff_B_AfHVPBWM0_1),.dout(w_dff_B_qMH1XlYV7_1),.clk(gclk));
	jdff dff_B_9PVZRrRo0_1(.din(w_dff_B_qMH1XlYV7_1),.dout(w_dff_B_9PVZRrRo0_1),.clk(gclk));
	jdff dff_B_luoa8u5s2_1(.din(n254),.dout(w_dff_B_luoa8u5s2_1),.clk(gclk));
	jdff dff_B_HGx1crMw7_1(.din(w_dff_B_luoa8u5s2_1),.dout(w_dff_B_HGx1crMw7_1),.clk(gclk));
	jdff dff_B_isDjTFWc8_1(.din(w_dff_B_HGx1crMw7_1),.dout(w_dff_B_isDjTFWc8_1),.clk(gclk));
	jdff dff_B_G8pYIdzQ9_1(.din(w_dff_B_isDjTFWc8_1),.dout(w_dff_B_G8pYIdzQ9_1),.clk(gclk));
	jdff dff_B_qM6LeDhA0_1(.din(w_dff_B_G8pYIdzQ9_1),.dout(w_dff_B_qM6LeDhA0_1),.clk(gclk));
	jdff dff_B_942GQbZg7_1(.din(n255),.dout(w_dff_B_942GQbZg7_1),.clk(gclk));
	jdff dff_B_KrePHkWA2_1(.din(w_dff_B_942GQbZg7_1),.dout(w_dff_B_KrePHkWA2_1),.clk(gclk));
	jdff dff_B_LHgrEym81_1(.din(w_dff_B_KrePHkWA2_1),.dout(w_dff_B_LHgrEym81_1),.clk(gclk));
	jdff dff_B_m7Ms08W15_1(.din(w_dff_B_LHgrEym81_1),.dout(w_dff_B_m7Ms08W15_1),.clk(gclk));
	jdff dff_B_3qwx3fib2_1(.din(w_dff_B_m7Ms08W15_1),.dout(w_dff_B_3qwx3fib2_1),.clk(gclk));
	jdff dff_B_hOBeDdU87_1(.din(w_dff_B_3qwx3fib2_1),.dout(w_dff_B_hOBeDdU87_1),.clk(gclk));
	jdff dff_B_xuEOVQNx2_1(.din(w_dff_B_hOBeDdU87_1),.dout(w_dff_B_xuEOVQNx2_1),.clk(gclk));
	jdff dff_B_O7GXZBuc5_1(.din(w_dff_B_xuEOVQNx2_1),.dout(w_dff_B_O7GXZBuc5_1),.clk(gclk));
	jdff dff_B_85UE8Pjn3_1(.din(w_dff_B_O7GXZBuc5_1),.dout(w_dff_B_85UE8Pjn3_1),.clk(gclk));
	jdff dff_B_elEKzFxD0_1(.din(w_dff_B_85UE8Pjn3_1),.dout(w_dff_B_elEKzFxD0_1),.clk(gclk));
	jdff dff_B_7Q0HnyIn1_1(.din(w_dff_B_elEKzFxD0_1),.dout(w_dff_B_7Q0HnyIn1_1),.clk(gclk));
	jdff dff_B_RRNJMLFZ9_1(.din(w_dff_B_7Q0HnyIn1_1),.dout(w_dff_B_RRNJMLFZ9_1),.clk(gclk));
	jdff dff_B_WTRgCdbs0_1(.din(w_dff_B_RRNJMLFZ9_1),.dout(w_dff_B_WTRgCdbs0_1),.clk(gclk));
	jdff dff_B_YKhgEew84_1(.din(w_dff_B_WTRgCdbs0_1),.dout(w_dff_B_YKhgEew84_1),.clk(gclk));
	jdff dff_A_GE2OFhcu2_0(.dout(w_n249_0[0]),.din(w_dff_A_GE2OFhcu2_0),.clk(gclk));
	jdff dff_B_PVwqqQDq9_0(.din(n248),.dout(w_dff_B_PVwqqQDq9_0),.clk(gclk));
	jdff dff_B_ruU0o0Zw5_0(.din(w_dff_B_PVwqqQDq9_0),.dout(w_dff_B_ruU0o0Zw5_0),.clk(gclk));
	jdff dff_B_8KuuX9pm7_0(.din(w_dff_B_ruU0o0Zw5_0),.dout(w_dff_B_8KuuX9pm7_0),.clk(gclk));
	jdff dff_B_M9k5CzIM1_0(.din(w_dff_B_8KuuX9pm7_0),.dout(w_dff_B_M9k5CzIM1_0),.clk(gclk));
	jdff dff_B_yHQjgJuJ2_0(.din(w_dff_B_M9k5CzIM1_0),.dout(w_dff_B_yHQjgJuJ2_0),.clk(gclk));
	jdff dff_A_ReIXFZ3E4_0(.dout(w_n247_0[0]),.din(w_dff_A_ReIXFZ3E4_0),.clk(gclk));
	jdff dff_A_n1HDuIrX2_0(.dout(w_dff_A_ReIXFZ3E4_0),.din(w_dff_A_n1HDuIrX2_0),.clk(gclk));
	jdff dff_A_nCbuYFbF4_0(.dout(w_dff_A_n1HDuIrX2_0),.din(w_dff_A_nCbuYFbF4_0),.clk(gclk));
	jdff dff_A_lxuzfnML8_0(.dout(w_dff_A_nCbuYFbF4_0),.din(w_dff_A_lxuzfnML8_0),.clk(gclk));
	jdff dff_A_XVDMd2Qt9_0(.dout(w_dff_A_lxuzfnML8_0),.din(w_dff_A_XVDMd2Qt9_0),.clk(gclk));
	jdff dff_A_xkJXqYtU3_0(.dout(w_dff_A_XVDMd2Qt9_0),.din(w_dff_A_xkJXqYtU3_0),.clk(gclk));
	jdff dff_A_ShDyOuw69_0(.dout(w_dff_A_xkJXqYtU3_0),.din(w_dff_A_ShDyOuw69_0),.clk(gclk));
	jdff dff_B_2ZtFWut93_0(.din(n246),.dout(w_dff_B_2ZtFWut93_0),.clk(gclk));
	jdff dff_B_oo0lapOU4_0(.din(w_dff_B_2ZtFWut93_0),.dout(w_dff_B_oo0lapOU4_0),.clk(gclk));
	jdff dff_B_69rNmGGs0_0(.din(w_dff_B_oo0lapOU4_0),.dout(w_dff_B_69rNmGGs0_0),.clk(gclk));
	jdff dff_B_aQmgpujQ6_0(.din(w_dff_B_69rNmGGs0_0),.dout(w_dff_B_aQmgpujQ6_0),.clk(gclk));
	jdff dff_B_tbSrLAWP7_0(.din(w_dff_B_aQmgpujQ6_0),.dout(w_dff_B_tbSrLAWP7_0),.clk(gclk));
	jdff dff_B_LZvlM0IF3_0(.din(w_dff_B_tbSrLAWP7_0),.dout(w_dff_B_LZvlM0IF3_0),.clk(gclk));
	jdff dff_B_KD1KIA7h3_0(.din(n229),.dout(w_dff_B_KD1KIA7h3_0),.clk(gclk));
	jdff dff_B_YG4D7ggH7_1(.din(n228),.dout(w_dff_B_YG4D7ggH7_1),.clk(gclk));
	jdff dff_A_PZkuwsVW8_0(.dout(w_n226_0[0]),.din(w_dff_A_PZkuwsVW8_0),.clk(gclk));
	jdff dff_A_K4uxcDgn9_0(.dout(w_dff_A_PZkuwsVW8_0),.din(w_dff_A_K4uxcDgn9_0),.clk(gclk));
	jdff dff_A_NBc9thxJ3_0(.dout(w_dff_A_K4uxcDgn9_0),.din(w_dff_A_NBc9thxJ3_0),.clk(gclk));
	jdff dff_A_AqEWRHx37_0(.dout(w_dff_A_NBc9thxJ3_0),.din(w_dff_A_AqEWRHx37_0),.clk(gclk));
	jdff dff_A_YqZae1nT9_0(.dout(w_dff_A_AqEWRHx37_0),.din(w_dff_A_YqZae1nT9_0),.clk(gclk));
	jdff dff_A_8AbjdZxs4_0(.dout(w_dff_A_YqZae1nT9_0),.din(w_dff_A_8AbjdZxs4_0),.clk(gclk));
	jdff dff_A_k9U9pe132_0(.dout(w_n225_0[0]),.din(w_dff_A_k9U9pe132_0),.clk(gclk));
	jdff dff_A_91Cc5cyW2_0(.dout(w_dff_A_k9U9pe132_0),.din(w_dff_A_91Cc5cyW2_0),.clk(gclk));
	jdff dff_A_8muuYSL54_0(.dout(w_dff_A_91Cc5cyW2_0),.din(w_dff_A_8muuYSL54_0),.clk(gclk));
	jdff dff_A_fsD8wDjC9_0(.dout(w_dff_A_8muuYSL54_0),.din(w_dff_A_fsD8wDjC9_0),.clk(gclk));
	jdff dff_A_DhUZeLp19_0(.dout(w_dff_A_fsD8wDjC9_0),.din(w_dff_A_DhUZeLp19_0),.clk(gclk));
	jdff dff_A_PwgyT2Fz5_0(.dout(w_dff_A_DhUZeLp19_0),.din(w_dff_A_PwgyT2Fz5_0),.clk(gclk));
	jdff dff_A_WZUhTPdu1_0(.dout(w_n218_0[0]),.din(w_dff_A_WZUhTPdu1_0),.clk(gclk));
	jdff dff_A_RQFR3mYA8_0(.dout(w_dff_A_WZUhTPdu1_0),.din(w_dff_A_RQFR3mYA8_0),.clk(gclk));
	jdff dff_A_gw2UTSY54_0(.dout(w_dff_A_RQFR3mYA8_0),.din(w_dff_A_gw2UTSY54_0),.clk(gclk));
	jdff dff_A_HLs4KfFJ8_0(.dout(w_dff_A_gw2UTSY54_0),.din(w_dff_A_HLs4KfFJ8_0),.clk(gclk));
	jdff dff_A_UP7wXcvy4_0(.dout(w_dff_A_HLs4KfFJ8_0),.din(w_dff_A_UP7wXcvy4_0),.clk(gclk));
	jdff dff_A_RBu1l1Gf3_0(.dout(w_dff_A_UP7wXcvy4_0),.din(w_dff_A_RBu1l1Gf3_0),.clk(gclk));
	jdff dff_A_mujE1H1o5_0(.dout(w_dff_A_RBu1l1Gf3_0),.din(w_dff_A_mujE1H1o5_0),.clk(gclk));
	jdff dff_A_94zoQHuY9_0(.dout(w_n272_0[0]),.din(w_dff_A_94zoQHuY9_0),.clk(gclk));
	jdff dff_B_68N1zJpU2_0(.din(n211),.dout(w_dff_B_68N1zJpU2_0),.clk(gclk));
	jdff dff_B_xtkQa4946_0(.din(w_dff_B_68N1zJpU2_0),.dout(w_dff_B_xtkQa4946_0),.clk(gclk));
	jdff dff_A_6yfuLoDF4_1(.dout(w_n207_0[1]),.din(w_dff_A_6yfuLoDF4_1),.clk(gclk));
	jdff dff_A_ieizIOyX8_1(.dout(w_dff_A_6yfuLoDF4_1),.din(w_dff_A_ieizIOyX8_1),.clk(gclk));
	jdff dff_A_xy0oMfl79_1(.dout(w_dff_A_ieizIOyX8_1),.din(w_dff_A_xy0oMfl79_1),.clk(gclk));
	jdff dff_A_hAehK1Cs4_1(.dout(w_G27gat_0[1]),.din(w_dff_A_hAehK1Cs4_1),.clk(gclk));
	jdff dff_A_lQHK98mN4_1(.dout(w_dff_A_hAehK1Cs4_1),.din(w_dff_A_lQHK98mN4_1),.clk(gclk));
	jdff dff_A_zELgvyFN6_1(.dout(w_dff_A_lQHK98mN4_1),.din(w_dff_A_zELgvyFN6_1),.clk(gclk));
	jdff dff_A_McLi8ER78_1(.dout(w_dff_A_zELgvyFN6_1),.din(w_dff_A_McLi8ER78_1),.clk(gclk));
	jdff dff_A_BZSrONRL7_1(.dout(w_dff_A_McLi8ER78_1),.din(w_dff_A_BZSrONRL7_1),.clk(gclk));
	jdff dff_A_Vgh3MVZc3_1(.dout(w_dff_A_BZSrONRL7_1),.din(w_dff_A_Vgh3MVZc3_1),.clk(gclk));
	jdff dff_A_JoDMAQsU7_1(.dout(w_dff_A_Vgh3MVZc3_1),.din(w_dff_A_JoDMAQsU7_1),.clk(gclk));
	jdff dff_A_8RULKxWV0_1(.dout(w_dff_A_JoDMAQsU7_1),.din(w_dff_A_8RULKxWV0_1),.clk(gclk));
	jdff dff_A_CRsJpwR56_1(.dout(w_dff_A_8RULKxWV0_1),.din(w_dff_A_CRsJpwR56_1),.clk(gclk));
	jdff dff_A_Q92DefhQ6_1(.dout(w_dff_A_CRsJpwR56_1),.din(w_dff_A_Q92DefhQ6_1),.clk(gclk));
	jdff dff_A_xq92GEQy6_1(.dout(w_dff_A_Q92DefhQ6_1),.din(w_dff_A_xq92GEQy6_1),.clk(gclk));
	jdff dff_A_vyQkkCnx5_1(.dout(w_dff_A_xq92GEQy6_1),.din(w_dff_A_vyQkkCnx5_1),.clk(gclk));
	jdff dff_A_nzXcZcit6_0(.dout(w_n202_0[0]),.din(w_dff_A_nzXcZcit6_0),.clk(gclk));
	jdff dff_A_UnTZFBYV3_0(.dout(w_dff_A_nzXcZcit6_0),.din(w_dff_A_UnTZFBYV3_0),.clk(gclk));
	jdff dff_A_KP6Pf0ls0_0(.dout(w_dff_A_UnTZFBYV3_0),.din(w_dff_A_KP6Pf0ls0_0),.clk(gclk));
	jdff dff_B_UGFk8mY89_1(.din(n199),.dout(w_dff_B_UGFk8mY89_1),.clk(gclk));
	jdff dff_B_mJ4HpQ7e4_1(.din(w_dff_B_UGFk8mY89_1),.dout(w_dff_B_mJ4HpQ7e4_1),.clk(gclk));
	jdff dff_B_cbneefmY0_1(.din(w_dff_B_mJ4HpQ7e4_1),.dout(w_dff_B_cbneefmY0_1),.clk(gclk));
	jdff dff_B_ktXJQKyJ8_1(.din(w_dff_B_cbneefmY0_1),.dout(w_dff_B_ktXJQKyJ8_1),.clk(gclk));
	jdff dff_B_28ySflHm4_1(.din(w_dff_B_ktXJQKyJ8_1),.dout(w_dff_B_28ySflHm4_1),.clk(gclk));
	jdff dff_B_r2GEpJMO4_1(.din(w_dff_B_28ySflHm4_1),.dout(w_dff_B_r2GEpJMO4_1),.clk(gclk));
	jdff dff_B_5GlQwz315_1(.din(w_dff_B_r2GEpJMO4_1),.dout(w_dff_B_5GlQwz315_1),.clk(gclk));
	jdff dff_B_XbRR5KLx1_1(.din(w_dff_B_5GlQwz315_1),.dout(w_dff_B_XbRR5KLx1_1),.clk(gclk));
	jdff dff_B_byLwmGvx2_1(.din(w_dff_B_XbRR5KLx1_1),.dout(w_dff_B_byLwmGvx2_1),.clk(gclk));
	jdff dff_B_rVkOIyrO2_1(.din(w_dff_B_byLwmGvx2_1),.dout(w_dff_B_rVkOIyrO2_1),.clk(gclk));
	jdff dff_B_MJYhPC8g8_1(.din(w_dff_B_rVkOIyrO2_1),.dout(w_dff_B_MJYhPC8g8_1),.clk(gclk));
	jdff dff_A_4yx1vEpq6_0(.dout(w_n201_0[0]),.din(w_dff_A_4yx1vEpq6_0),.clk(gclk));
	jdff dff_A_9wHwzcwr9_0(.dout(w_dff_A_4yx1vEpq6_0),.din(w_dff_A_9wHwzcwr9_0),.clk(gclk));
	jdff dff_A_ZIdL7NhX7_0(.dout(w_dff_A_9wHwzcwr9_0),.din(w_dff_A_ZIdL7NhX7_0),.clk(gclk));
	jdff dff_A_sPeF0eZf4_0(.dout(w_G66gat_0[0]),.din(w_dff_A_sPeF0eZf4_0),.clk(gclk));
	jdff dff_A_YTtw4F179_0(.dout(w_dff_A_sPeF0eZf4_0),.din(w_dff_A_YTtw4F179_0),.clk(gclk));
	jdff dff_A_GvdEzcgx3_0(.dout(w_dff_A_YTtw4F179_0),.din(w_dff_A_GvdEzcgx3_0),.clk(gclk));
	jdff dff_A_2efNFSLi2_0(.dout(w_dff_A_GvdEzcgx3_0),.din(w_dff_A_2efNFSLi2_0),.clk(gclk));
	jdff dff_A_7kLnfmXa8_0(.dout(w_dff_A_2efNFSLi2_0),.din(w_dff_A_7kLnfmXa8_0),.clk(gclk));
	jdff dff_A_TJYPW7SA8_0(.dout(w_dff_A_7kLnfmXa8_0),.din(w_dff_A_TJYPW7SA8_0),.clk(gclk));
	jdff dff_A_Uc3CZSEp6_0(.dout(w_dff_A_TJYPW7SA8_0),.din(w_dff_A_Uc3CZSEp6_0),.clk(gclk));
	jdff dff_A_rWyCF3Mx5_0(.dout(w_dff_A_Uc3CZSEp6_0),.din(w_dff_A_rWyCF3Mx5_0),.clk(gclk));
	jdff dff_A_dR0YlQd23_0(.dout(w_dff_A_rWyCF3Mx5_0),.din(w_dff_A_dR0YlQd23_0),.clk(gclk));
	jdff dff_A_vsUmunHW1_0(.dout(w_n197_0[0]),.din(w_dff_A_vsUmunHW1_0),.clk(gclk));
	jdff dff_A_yqAPWQ7j5_0(.dout(w_dff_A_vsUmunHW1_0),.din(w_dff_A_yqAPWQ7j5_0),.clk(gclk));
	jdff dff_A_E3aw4bMf4_0(.dout(w_dff_A_yqAPWQ7j5_0),.din(w_dff_A_E3aw4bMf4_0),.clk(gclk));
	jdff dff_A_BnZcShms0_0(.dout(w_n195_0[0]),.din(w_dff_A_BnZcShms0_0),.clk(gclk));
	jdff dff_A_8dErt7Uh6_0(.dout(w_dff_A_BnZcShms0_0),.din(w_dff_A_8dErt7Uh6_0),.clk(gclk));
	jdff dff_A_6TmgDA501_0(.dout(w_dff_A_8dErt7Uh6_0),.din(w_dff_A_6TmgDA501_0),.clk(gclk));
	jdff dff_B_XeoHgJba5_2(.din(n195),.dout(w_dff_B_XeoHgJba5_2),.clk(gclk));
	jdff dff_B_GCytSAJh7_2(.din(w_dff_B_XeoHgJba5_2),.dout(w_dff_B_GCytSAJh7_2),.clk(gclk));
	jdff dff_B_2BS1ZbFY3_2(.din(w_dff_B_GCytSAJh7_2),.dout(w_dff_B_2BS1ZbFY3_2),.clk(gclk));
	jdff dff_B_iYUb8tV98_2(.din(w_dff_B_2BS1ZbFY3_2),.dout(w_dff_B_iYUb8tV98_2),.clk(gclk));
	jdff dff_B_LiqyjzZT8_2(.din(w_dff_B_iYUb8tV98_2),.dout(w_dff_B_LiqyjzZT8_2),.clk(gclk));
	jdff dff_B_byhoR8gJ7_2(.din(w_dff_B_LiqyjzZT8_2),.dout(w_dff_B_byhoR8gJ7_2),.clk(gclk));
	jdff dff_B_XRDK1Pva7_2(.din(w_dff_B_byhoR8gJ7_2),.dout(w_dff_B_XRDK1Pva7_2),.clk(gclk));
	jdff dff_B_UuBqLHac4_2(.din(w_dff_B_XRDK1Pva7_2),.dout(w_dff_B_UuBqLHac4_2),.clk(gclk));
	jdff dff_B_EU06pYH15_2(.din(w_dff_B_UuBqLHac4_2),.dout(w_dff_B_EU06pYH15_2),.clk(gclk));
	jdff dff_B_o8r2mS3D1_2(.din(w_dff_B_EU06pYH15_2),.dout(w_dff_B_o8r2mS3D1_2),.clk(gclk));
	jdff dff_B_jOeKJE9G9_2(.din(w_dff_B_o8r2mS3D1_2),.dout(w_dff_B_jOeKJE9G9_2),.clk(gclk));
	jdff dff_A_5MIIGepJ3_0(.dout(w_G40gat_0[0]),.din(w_dff_A_5MIIGepJ3_0),.clk(gclk));
	jdff dff_A_uvbPFJi35_0(.dout(w_dff_A_5MIIGepJ3_0),.din(w_dff_A_uvbPFJi35_0),.clk(gclk));
	jdff dff_A_Li8I2X4j0_0(.dout(w_dff_A_uvbPFJi35_0),.din(w_dff_A_Li8I2X4j0_0),.clk(gclk));
	jdff dff_A_QI6UNgV19_0(.dout(w_dff_A_Li8I2X4j0_0),.din(w_dff_A_QI6UNgV19_0),.clk(gclk));
	jdff dff_A_CsTHdnFB4_0(.dout(w_dff_A_QI6UNgV19_0),.din(w_dff_A_CsTHdnFB4_0),.clk(gclk));
	jdff dff_A_W2VpZEpB3_0(.dout(w_dff_A_CsTHdnFB4_0),.din(w_dff_A_W2VpZEpB3_0),.clk(gclk));
	jdff dff_A_E2fhySV26_0(.dout(w_dff_A_W2VpZEpB3_0),.din(w_dff_A_E2fhySV26_0),.clk(gclk));
	jdff dff_A_Sgzihm8T1_0(.dout(w_dff_A_E2fhySV26_0),.din(w_dff_A_Sgzihm8T1_0),.clk(gclk));
	jdff dff_A_tS1vBQgN2_0(.dout(w_dff_A_Sgzihm8T1_0),.din(w_dff_A_tS1vBQgN2_0),.clk(gclk));
	jdff dff_A_w2Gc8ey23_0(.dout(w_dff_A_tS1vBQgN2_0),.din(w_dff_A_w2Gc8ey23_0),.clk(gclk));
	jdff dff_A_YvMlf2Pl8_0(.dout(w_dff_A_w2Gc8ey23_0),.din(w_dff_A_YvMlf2Pl8_0),.clk(gclk));
	jdff dff_A_aEGAr0Tv2_0(.dout(w_dff_A_YvMlf2Pl8_0),.din(w_dff_A_aEGAr0Tv2_0),.clk(gclk));
	jdff dff_A_aoQOdcg27_0(.dout(w_dff_A_aEGAr0Tv2_0),.din(w_dff_A_aoQOdcg27_0),.clk(gclk));
	jdff dff_A_wxXA6H3I1_0(.dout(w_dff_A_aoQOdcg27_0),.din(w_dff_A_wxXA6H3I1_0),.clk(gclk));
	jdff dff_A_yS8gKoul0_0(.dout(w_dff_A_wxXA6H3I1_0),.din(w_dff_A_yS8gKoul0_0),.clk(gclk));
	jdff dff_A_w8nMvLQ22_1(.dout(w_G40gat_0[1]),.din(w_dff_A_w8nMvLQ22_1),.clk(gclk));
	jdff dff_A_mLWRzPG60_1(.dout(w_dff_A_w8nMvLQ22_1),.din(w_dff_A_mLWRzPG60_1),.clk(gclk));
	jdff dff_A_UIu5GpSN2_1(.dout(w_dff_A_mLWRzPG60_1),.din(w_dff_A_UIu5GpSN2_1),.clk(gclk));
	jdff dff_A_isKyIbqO3_1(.dout(w_dff_A_UIu5GpSN2_1),.din(w_dff_A_isKyIbqO3_1),.clk(gclk));
	jdff dff_A_FyDsKn3i2_1(.dout(w_dff_A_isKyIbqO3_1),.din(w_dff_A_FyDsKn3i2_1),.clk(gclk));
	jdff dff_A_rcjvKEdG1_1(.dout(w_dff_A_FyDsKn3i2_1),.din(w_dff_A_rcjvKEdG1_1),.clk(gclk));
	jdff dff_A_RxegrnXh8_1(.dout(w_dff_A_rcjvKEdG1_1),.din(w_dff_A_RxegrnXh8_1),.clk(gclk));
	jdff dff_A_5SZFa6fs4_1(.dout(w_dff_A_RxegrnXh8_1),.din(w_dff_A_5SZFa6fs4_1),.clk(gclk));
	jdff dff_A_tYJmetl42_1(.dout(w_dff_A_5SZFa6fs4_1),.din(w_dff_A_tYJmetl42_1),.clk(gclk));
	jdff dff_B_VmHWFZ5U6_0(.din(n193),.dout(w_dff_B_VmHWFZ5U6_0),.clk(gclk));
	jdff dff_B_HDPAEKzA6_0(.din(w_dff_B_VmHWFZ5U6_0),.dout(w_dff_B_HDPAEKzA6_0),.clk(gclk));
	jdff dff_B_U6hfzyHL4_0(.din(w_dff_B_HDPAEKzA6_0),.dout(w_dff_B_U6hfzyHL4_0),.clk(gclk));
	jdff dff_A_ojvFAyzI4_0(.dout(w_n189_0[0]),.din(w_dff_A_ojvFAyzI4_0),.clk(gclk));
	jdff dff_A_WGyhBl7F5_0(.dout(w_dff_A_ojvFAyzI4_0),.din(w_dff_A_WGyhBl7F5_0),.clk(gclk));
	jdff dff_A_GzaeScc69_0(.dout(w_dff_A_WGyhBl7F5_0),.din(w_dff_A_GzaeScc69_0),.clk(gclk));
	jdff dff_A_ldma2cIp4_0(.dout(w_dff_A_GzaeScc69_0),.din(w_dff_A_ldma2cIp4_0),.clk(gclk));
	jdff dff_A_EjkXA34m6_0(.dout(w_dff_A_ldma2cIp4_0),.din(w_dff_A_EjkXA34m6_0),.clk(gclk));
	jdff dff_A_L6DoBOc54_0(.dout(w_dff_A_EjkXA34m6_0),.din(w_dff_A_L6DoBOc54_0),.clk(gclk));
	jdff dff_A_atlUkYPM4_0(.dout(w_dff_A_L6DoBOc54_0),.din(w_dff_A_atlUkYPM4_0),.clk(gclk));
	jdff dff_A_Oiq5S9mx3_0(.dout(w_dff_A_atlUkYPM4_0),.din(w_dff_A_Oiq5S9mx3_0),.clk(gclk));
	jdff dff_B_ifLLn9bo9_2(.din(n189),.dout(w_dff_B_ifLLn9bo9_2),.clk(gclk));
	jdff dff_B_a9k85SDt9_2(.din(w_dff_B_ifLLn9bo9_2),.dout(w_dff_B_a9k85SDt9_2),.clk(gclk));
	jdff dff_B_LcB3bNJq6_2(.din(w_dff_B_a9k85SDt9_2),.dout(w_dff_B_LcB3bNJq6_2),.clk(gclk));
	jdff dff_B_SGpQRxIW2_2(.din(w_dff_B_LcB3bNJq6_2),.dout(w_dff_B_SGpQRxIW2_2),.clk(gclk));
	jdff dff_B_vmMr3mZX0_2(.din(w_dff_B_SGpQRxIW2_2),.dout(w_dff_B_vmMr3mZX0_2),.clk(gclk));
	jdff dff_B_oOjS4uHz8_2(.din(w_dff_B_vmMr3mZX0_2),.dout(w_dff_B_oOjS4uHz8_2),.clk(gclk));
	jdff dff_A_LjKIH6Ya0_0(.dout(w_G53gat_0[0]),.din(w_dff_A_LjKIH6Ya0_0),.clk(gclk));
	jdff dff_A_5Cq5ZEri1_0(.dout(w_dff_A_LjKIH6Ya0_0),.din(w_dff_A_5Cq5ZEri1_0),.clk(gclk));
	jdff dff_A_JaZGIrAh4_0(.dout(w_dff_A_5Cq5ZEri1_0),.din(w_dff_A_JaZGIrAh4_0),.clk(gclk));
	jdff dff_A_dKayZWHU3_0(.dout(w_dff_A_JaZGIrAh4_0),.din(w_dff_A_dKayZWHU3_0),.clk(gclk));
	jdff dff_A_7uakt8qp7_0(.dout(w_dff_A_dKayZWHU3_0),.din(w_dff_A_7uakt8qp7_0),.clk(gclk));
	jdff dff_A_2afSD2El5_0(.dout(w_dff_A_7uakt8qp7_0),.din(w_dff_A_2afSD2El5_0),.clk(gclk));
	jdff dff_A_iP8barNH1_0(.dout(w_dff_A_2afSD2El5_0),.din(w_dff_A_iP8barNH1_0),.clk(gclk));
	jdff dff_A_GEdCW9EV8_0(.dout(w_dff_A_iP8barNH1_0),.din(w_dff_A_GEdCW9EV8_0),.clk(gclk));
	jdff dff_A_u3Rvaf0U0_0(.dout(w_dff_A_GEdCW9EV8_0),.din(w_dff_A_u3Rvaf0U0_0),.clk(gclk));
	jdff dff_A_EMuH6fZS8_0(.dout(w_dff_A_u3Rvaf0U0_0),.din(w_dff_A_EMuH6fZS8_0),.clk(gclk));
	jdff dff_A_HgpdXnc60_0(.dout(w_dff_A_EMuH6fZS8_0),.din(w_dff_A_HgpdXnc60_0),.clk(gclk));
	jdff dff_A_e10ykomm2_0(.dout(w_dff_A_HgpdXnc60_0),.din(w_dff_A_e10ykomm2_0),.clk(gclk));
	jdff dff_A_judq4vel5_0(.dout(w_dff_A_e10ykomm2_0),.din(w_dff_A_judq4vel5_0),.clk(gclk));
	jdff dff_A_KPJ9DGpu2_0(.dout(w_dff_A_judq4vel5_0),.din(w_dff_A_KPJ9DGpu2_0),.clk(gclk));
	jdff dff_A_BerntqP88_0(.dout(w_dff_A_KPJ9DGpu2_0),.din(w_dff_A_BerntqP88_0),.clk(gclk));
	jdff dff_B_yd1ok6pc7_1(.din(n184),.dout(w_dff_B_yd1ok6pc7_1),.clk(gclk));
	jdff dff_B_1PuDcvmp9_1(.din(w_dff_B_yd1ok6pc7_1),.dout(w_dff_B_1PuDcvmp9_1),.clk(gclk));
	jdff dff_B_ODrf1TBp8_1(.din(w_dff_B_1PuDcvmp9_1),.dout(w_dff_B_ODrf1TBp8_1),.clk(gclk));
	jdff dff_B_stWsCTyc4_1(.din(w_dff_B_ODrf1TBp8_1),.dout(w_dff_B_stWsCTyc4_1),.clk(gclk));
	jdff dff_B_mIss7T1O5_1(.din(w_dff_B_stWsCTyc4_1),.dout(w_dff_B_mIss7T1O5_1),.clk(gclk));
	jdff dff_B_ZQio1wDY4_1(.din(w_dff_B_mIss7T1O5_1),.dout(w_dff_B_ZQio1wDY4_1),.clk(gclk));
	jdff dff_B_rqcJEdQT1_1(.din(w_dff_B_ZQio1wDY4_1),.dout(w_dff_B_rqcJEdQT1_1),.clk(gclk));
	jdff dff_B_E6Nltixk5_1(.din(w_dff_B_rqcJEdQT1_1),.dout(w_dff_B_E6Nltixk5_1),.clk(gclk));
	jdff dff_B_ATBLh0m31_1(.din(w_dff_B_E6Nltixk5_1),.dout(w_dff_B_ATBLh0m31_1),.clk(gclk));
	jdff dff_B_gvt5VaHr4_1(.din(w_dff_B_ATBLh0m31_1),.dout(w_dff_B_gvt5VaHr4_1),.clk(gclk));
	jdff dff_B_g91zQXQd2_1(.din(w_dff_B_gvt5VaHr4_1),.dout(w_dff_B_g91zQXQd2_1),.clk(gclk));
	jdff dff_A_Ov4Q1z1y4_0(.dout(w_G92gat_0[0]),.din(w_dff_A_Ov4Q1z1y4_0),.clk(gclk));
	jdff dff_A_CvHOYBHq4_0(.dout(w_dff_A_Ov4Q1z1y4_0),.din(w_dff_A_CvHOYBHq4_0),.clk(gclk));
	jdff dff_A_0yLVUsEt2_0(.dout(w_dff_A_CvHOYBHq4_0),.din(w_dff_A_0yLVUsEt2_0),.clk(gclk));
	jdff dff_A_iN07iLxl3_0(.dout(w_dff_A_0yLVUsEt2_0),.din(w_dff_A_iN07iLxl3_0),.clk(gclk));
	jdff dff_A_yM4uPf3c8_0(.dout(w_dff_A_iN07iLxl3_0),.din(w_dff_A_yM4uPf3c8_0),.clk(gclk));
	jdff dff_A_r9uPBkP90_0(.dout(w_dff_A_yM4uPf3c8_0),.din(w_dff_A_r9uPBkP90_0),.clk(gclk));
	jdff dff_A_TbzDJM6C6_0(.dout(w_dff_A_r9uPBkP90_0),.din(w_dff_A_TbzDJM6C6_0),.clk(gclk));
	jdff dff_A_0MstNCHM3_0(.dout(w_dff_A_TbzDJM6C6_0),.din(w_dff_A_0MstNCHM3_0),.clk(gclk));
	jdff dff_A_ECgu0i0u9_0(.dout(w_dff_A_0MstNCHM3_0),.din(w_dff_A_ECgu0i0u9_0),.clk(gclk));
	jdff dff_A_Ke94OlAN3_0(.dout(w_dff_A_ECgu0i0u9_0),.din(w_dff_A_Ke94OlAN3_0),.clk(gclk));
	jdff dff_A_Kwz5zZVd7_0(.dout(w_dff_A_Ke94OlAN3_0),.din(w_dff_A_Kwz5zZVd7_0),.clk(gclk));
	jdff dff_A_c4I3kAog5_0(.dout(w_dff_A_Kwz5zZVd7_0),.din(w_dff_A_c4I3kAog5_0),.clk(gclk));
	jdff dff_A_gL4pC2X05_0(.dout(w_dff_A_c4I3kAog5_0),.din(w_dff_A_gL4pC2X05_0),.clk(gclk));
	jdff dff_A_9cCOg7SE5_0(.dout(w_dff_A_gL4pC2X05_0),.din(w_dff_A_9cCOg7SE5_0),.clk(gclk));
	jdff dff_A_LKzdN1yI2_0(.dout(w_dff_A_9cCOg7SE5_0),.din(w_dff_A_LKzdN1yI2_0),.clk(gclk));
	jdff dff_A_m2r5LI4g3_1(.dout(w_G92gat_0[1]),.din(w_dff_A_m2r5LI4g3_1),.clk(gclk));
	jdff dff_A_RhCgGiEP4_1(.dout(w_dff_A_m2r5LI4g3_1),.din(w_dff_A_RhCgGiEP4_1),.clk(gclk));
	jdff dff_A_GtfoIOcj3_1(.dout(w_dff_A_RhCgGiEP4_1),.din(w_dff_A_GtfoIOcj3_1),.clk(gclk));
	jdff dff_A_IDgJycOp3_1(.dout(w_dff_A_GtfoIOcj3_1),.din(w_dff_A_IDgJycOp3_1),.clk(gclk));
	jdff dff_A_Dx5Cydes3_1(.dout(w_dff_A_IDgJycOp3_1),.din(w_dff_A_Dx5Cydes3_1),.clk(gclk));
	jdff dff_A_h5yox54O9_1(.dout(w_dff_A_Dx5Cydes3_1),.din(w_dff_A_h5yox54O9_1),.clk(gclk));
	jdff dff_A_G22iVq2z4_1(.dout(w_dff_A_h5yox54O9_1),.din(w_dff_A_G22iVq2z4_1),.clk(gclk));
	jdff dff_A_81gjq9Pq9_1(.dout(w_dff_A_G22iVq2z4_1),.din(w_dff_A_81gjq9Pq9_1),.clk(gclk));
	jdff dff_A_61v04UO43_1(.dout(w_dff_A_81gjq9Pq9_1),.din(w_dff_A_61v04UO43_1),.clk(gclk));
	jdff dff_B_xl0nsL2C9_0(.din(n181),.dout(w_dff_B_xl0nsL2C9_0),.clk(gclk));
	jdff dff_B_RncHQkKu0_0(.din(w_dff_B_xl0nsL2C9_0),.dout(w_dff_B_RncHQkKu0_0),.clk(gclk));
	jdff dff_B_HQsFRl0s9_0(.din(w_dff_B_RncHQkKu0_0),.dout(w_dff_B_HQsFRl0s9_0),.clk(gclk));
	jdff dff_B_zBaBPsNS7_1(.din(n177),.dout(w_dff_B_zBaBPsNS7_1),.clk(gclk));
	jdff dff_B_Yh1HPGxF1_1(.din(w_dff_B_zBaBPsNS7_1),.dout(w_dff_B_Yh1HPGxF1_1),.clk(gclk));
	jdff dff_A_EKbmkh4Y2_1(.dout(w_G79gat_0[1]),.din(w_dff_A_EKbmkh4Y2_1),.clk(gclk));
	jdff dff_A_ixCgi5V25_1(.dout(w_dff_A_EKbmkh4Y2_1),.din(w_dff_A_ixCgi5V25_1),.clk(gclk));
	jdff dff_A_HISKe9X16_1(.dout(w_dff_A_ixCgi5V25_1),.din(w_dff_A_HISKe9X16_1),.clk(gclk));
	jdff dff_A_v550qsGB8_1(.dout(w_dff_A_HISKe9X16_1),.din(w_dff_A_v550qsGB8_1),.clk(gclk));
	jdff dff_A_gBfxMIlS5_1(.dout(w_dff_A_v550qsGB8_1),.din(w_dff_A_gBfxMIlS5_1),.clk(gclk));
	jdff dff_A_GQIGf68I0_1(.dout(w_dff_A_gBfxMIlS5_1),.din(w_dff_A_GQIGf68I0_1),.clk(gclk));
	jdff dff_A_E3VEHWhc4_1(.dout(w_dff_A_GQIGf68I0_1),.din(w_dff_A_E3VEHWhc4_1),.clk(gclk));
	jdff dff_A_aEstPw1q1_1(.dout(w_dff_A_E3VEHWhc4_1),.din(w_dff_A_aEstPw1q1_1),.clk(gclk));
	jdff dff_A_KLXF1nLE7_1(.dout(w_dff_A_aEstPw1q1_1),.din(w_dff_A_KLXF1nLE7_1),.clk(gclk));
	jdff dff_A_uDNfJlIO6_1(.dout(w_G105gat_0[1]),.din(w_dff_A_uDNfJlIO6_1),.clk(gclk));
	jdff dff_A_Un7fl79t1_1(.dout(w_dff_A_uDNfJlIO6_1),.din(w_dff_A_Un7fl79t1_1),.clk(gclk));
	jdff dff_A_g0R80RuZ0_1(.dout(w_dff_A_Un7fl79t1_1),.din(w_dff_A_g0R80RuZ0_1),.clk(gclk));
	jdff dff_A_bkIhgypG9_1(.dout(w_dff_A_g0R80RuZ0_1),.din(w_dff_A_bkIhgypG9_1),.clk(gclk));
	jdff dff_A_pWNaMWyj8_1(.dout(w_dff_A_bkIhgypG9_1),.din(w_dff_A_pWNaMWyj8_1),.clk(gclk));
	jdff dff_A_dSLAO5fQ6_1(.dout(w_dff_A_pWNaMWyj8_1),.din(w_dff_A_dSLAO5fQ6_1),.clk(gclk));
	jdff dff_A_DNa8Zykm6_1(.dout(w_dff_A_dSLAO5fQ6_1),.din(w_dff_A_DNa8Zykm6_1),.clk(gclk));
	jdff dff_A_iXkBClZk6_1(.dout(w_dff_A_DNa8Zykm6_1),.din(w_dff_A_iXkBClZk6_1),.clk(gclk));
	jdff dff_A_jkf4lP8S1_1(.dout(w_dff_A_iXkBClZk6_1),.din(w_dff_A_jkf4lP8S1_1),.clk(gclk));
	jdff dff_B_v9KblQxF4_1(.din(n138),.dout(w_dff_B_v9KblQxF4_1),.clk(gclk));
	jdff dff_B_ja6GFkp55_1(.din(w_dff_B_v9KblQxF4_1),.dout(w_dff_B_ja6GFkp55_1),.clk(gclk));
	jdff dff_B_PKRTrW9k6_1(.din(w_dff_B_ja6GFkp55_1),.dout(w_dff_B_PKRTrW9k6_1),.clk(gclk));
	jdff dff_B_qchdsOK64_1(.din(n143),.dout(w_dff_B_qchdsOK64_1),.clk(gclk));
	jdff dff_B_0eTdbLvy9_1(.din(n158),.dout(w_dff_B_0eTdbLvy9_1),.clk(gclk));
	jdff dff_B_4admQqlc7_1(.din(w_dff_B_0eTdbLvy9_1),.dout(w_dff_B_4admQqlc7_1),.clk(gclk));
	jdff dff_B_lCZrej0r6_1(.din(w_dff_B_4admQqlc7_1),.dout(w_dff_B_lCZrej0r6_1),.clk(gclk));
	jdff dff_B_xArl4hZ86_1(.din(w_dff_B_lCZrej0r6_1),.dout(w_dff_B_xArl4hZ86_1),.clk(gclk));
	jdff dff_B_ZsflEea39_0(.din(n166),.dout(w_dff_B_ZsflEea39_0),.clk(gclk));
	jdff dff_B_B0uRk8bE6_0(.din(w_dff_B_ZsflEea39_0),.dout(w_dff_B_B0uRk8bE6_0),.clk(gclk));
	jdff dff_B_Dr7YYBEp1_0(.din(w_dff_B_B0uRk8bE6_0),.dout(w_dff_B_Dr7YYBEp1_0),.clk(gclk));
	jdff dff_B_ekWoYZaN3_0(.din(w_dff_B_Dr7YYBEp1_0),.dout(w_dff_B_ekWoYZaN3_0),.clk(gclk));
	jdff dff_A_6AUVUaT74_0(.dout(w_n164_0[0]),.din(w_dff_A_6AUVUaT74_0),.clk(gclk));
	jdff dff_A_GPKoMvTx2_0(.dout(w_dff_A_6AUVUaT74_0),.din(w_dff_A_GPKoMvTx2_0),.clk(gclk));
	jdff dff_A_e6Vpsc8Y2_0(.dout(w_dff_A_GPKoMvTx2_0),.din(w_dff_A_e6Vpsc8Y2_0),.clk(gclk));
	jdff dff_A_RHIhLvQ85_0(.dout(w_dff_A_e6Vpsc8Y2_0),.din(w_dff_A_RHIhLvQ85_0),.clk(gclk));
	jdff dff_A_EvJ7Vh3W1_0(.dout(w_dff_A_RHIhLvQ85_0),.din(w_dff_A_EvJ7Vh3W1_0),.clk(gclk));
	jdff dff_A_rOnrJ9g02_0(.dout(w_dff_A_EvJ7Vh3W1_0),.din(w_dff_A_rOnrJ9g02_0),.clk(gclk));
	jdff dff_A_6APx0r583_0(.dout(w_n161_0[0]),.din(w_dff_A_6APx0r583_0),.clk(gclk));
	jdff dff_A_JcoH8Tot4_0(.dout(w_dff_A_6APx0r583_0),.din(w_dff_A_JcoH8Tot4_0),.clk(gclk));
	jdff dff_A_DspAH3ge2_0(.dout(w_dff_A_JcoH8Tot4_0),.din(w_dff_A_DspAH3ge2_0),.clk(gclk));
	jdff dff_A_2yC9AYMb3_0(.dout(w_dff_A_DspAH3ge2_0),.din(w_dff_A_2yC9AYMb3_0),.clk(gclk));
	jdff dff_A_Iz7S5QaJ7_0(.dout(w_dff_A_2yC9AYMb3_0),.din(w_dff_A_Iz7S5QaJ7_0),.clk(gclk));
	jdff dff_A_VdyfJxk62_0(.dout(w_dff_A_Iz7S5QaJ7_0),.din(w_dff_A_VdyfJxk62_0),.clk(gclk));
	jdff dff_A_M5ir2P5r5_0(.dout(w_n155_0[0]),.din(w_dff_A_M5ir2P5r5_0),.clk(gclk));
	jdff dff_A_Ks7F7ZGn3_0(.dout(w_dff_A_M5ir2P5r5_0),.din(w_dff_A_Ks7F7ZGn3_0),.clk(gclk));
	jdff dff_A_LclFNCTp1_0(.dout(w_dff_A_Ks7F7ZGn3_0),.din(w_dff_A_LclFNCTp1_0),.clk(gclk));
	jdff dff_A_aW0Pg6av4_0(.dout(w_dff_A_LclFNCTp1_0),.din(w_dff_A_aW0Pg6av4_0),.clk(gclk));
	jdff dff_A_sU6PWbBk3_0(.dout(w_dff_A_aW0Pg6av4_0),.din(w_dff_A_sU6PWbBk3_0),.clk(gclk));
	jdff dff_A_F5CDsX0C8_0(.dout(w_dff_A_sU6PWbBk3_0),.din(w_dff_A_F5CDsX0C8_0),.clk(gclk));
	jdff dff_B_ZMk9tluA8_1(.din(n153),.dout(w_dff_B_ZMk9tluA8_1),.clk(gclk));
	jdff dff_B_whZGNrI84_1(.din(w_dff_B_ZMk9tluA8_1),.dout(w_dff_B_whZGNrI84_1),.clk(gclk));
	jdff dff_A_qcDIukFr1_0(.dout(w_n146_0[0]),.din(w_dff_A_qcDIukFr1_0),.clk(gclk));
	jdff dff_A_CBrLCcUq5_0(.dout(w_dff_A_qcDIukFr1_0),.din(w_dff_A_CBrLCcUq5_0),.clk(gclk));
	jdff dff_A_UGzJx2Bv7_0(.dout(w_dff_A_CBrLCcUq5_0),.din(w_dff_A_UGzJx2Bv7_0),.clk(gclk));
	jdff dff_A_qzvYOYxS1_0(.dout(w_dff_A_UGzJx2Bv7_0),.din(w_dff_A_qzvYOYxS1_0),.clk(gclk));
	jdff dff_A_pI12VvBE9_0(.dout(w_dff_A_qzvYOYxS1_0),.din(w_dff_A_pI12VvBE9_0),.clk(gclk));
	jdff dff_A_gM7zOEJQ0_0(.dout(w_dff_A_pI12VvBE9_0),.din(w_dff_A_gM7zOEJQ0_0),.clk(gclk));
	jdff dff_B_ehbpL0nn8_1(.din(n144),.dout(w_dff_B_ehbpL0nn8_1),.clk(gclk));
	jdff dff_B_J9UvRJ9I9_1(.din(w_dff_B_ehbpL0nn8_1),.dout(w_dff_B_J9UvRJ9I9_1),.clk(gclk));
	jdff dff_A_oKx4W6Og0_0(.dout(w_G14gat_0[0]),.din(w_dff_A_oKx4W6Og0_0),.clk(gclk));
	jdff dff_A_EaE462m80_0(.dout(w_dff_A_oKx4W6Og0_0),.din(w_dff_A_EaE462m80_0),.clk(gclk));
	jdff dff_A_8pYhuuVD5_0(.dout(w_dff_A_EaE462m80_0),.din(w_dff_A_8pYhuuVD5_0),.clk(gclk));
	jdff dff_B_bp6EqDuX6_2(.din(G14gat),.dout(w_dff_B_bp6EqDuX6_2),.clk(gclk));
	jdff dff_B_MRMhKywC7_2(.din(w_dff_B_bp6EqDuX6_2),.dout(w_dff_B_MRMhKywC7_2),.clk(gclk));
	jdff dff_B_qkAUPKKp2_2(.din(w_dff_B_MRMhKywC7_2),.dout(w_dff_B_qkAUPKKp2_2),.clk(gclk));
	jdff dff_B_mGAm7GE30_2(.din(w_dff_B_qkAUPKKp2_2),.dout(w_dff_B_mGAm7GE30_2),.clk(gclk));
	jdff dff_B_SXsvtxlY5_2(.din(w_dff_B_mGAm7GE30_2),.dout(w_dff_B_SXsvtxlY5_2),.clk(gclk));
	jdff dff_B_MQJwHhR13_2(.din(w_dff_B_SXsvtxlY5_2),.dout(w_dff_B_MQJwHhR13_2),.clk(gclk));
	jdff dff_B_X3IFIq1E5_2(.din(w_dff_B_MQJwHhR13_2),.dout(w_dff_B_X3IFIq1E5_2),.clk(gclk));
	jdff dff_B_BMfeVFkL4_2(.din(w_dff_B_X3IFIq1E5_2),.dout(w_dff_B_BMfeVFkL4_2),.clk(gclk));
	jdff dff_B_6Iq6BaXp3_2(.din(w_dff_B_BMfeVFkL4_2),.dout(w_dff_B_6Iq6BaXp3_2),.clk(gclk));
	jdff dff_B_VAejou2l3_2(.din(w_dff_B_6Iq6BaXp3_2),.dout(w_dff_B_VAejou2l3_2),.clk(gclk));
	jdff dff_B_rIMAXny88_2(.din(w_dff_B_VAejou2l3_2),.dout(w_dff_B_rIMAXny88_2),.clk(gclk));
	jdff dff_B_iw6PA2gg1_2(.din(w_dff_B_rIMAXny88_2),.dout(w_dff_B_iw6PA2gg1_2),.clk(gclk));
	jdff dff_A_dZlt55fP7_0(.dout(w_n142_0[0]),.din(w_dff_A_dZlt55fP7_0),.clk(gclk));
	jdff dff_A_EEO3t36o4_0(.dout(w_dff_A_dZlt55fP7_0),.din(w_dff_A_EEO3t36o4_0),.clk(gclk));
	jdff dff_A_3132Il2W8_0(.dout(w_dff_A_EEO3t36o4_0),.din(w_dff_A_3132Il2W8_0),.clk(gclk));
	jdff dff_A_7MulR8yy0_0(.dout(w_dff_A_3132Il2W8_0),.din(w_dff_A_7MulR8yy0_0),.clk(gclk));
	jdff dff_B_egok4NA54_2(.din(n142),.dout(w_dff_B_egok4NA54_2),.clk(gclk));
	jdff dff_B_b1pIRL3U3_2(.din(w_dff_B_egok4NA54_2),.dout(w_dff_B_b1pIRL3U3_2),.clk(gclk));
	jdff dff_B_WR30poUH6_2(.din(w_dff_B_b1pIRL3U3_2),.dout(w_dff_B_WR30poUH6_2),.clk(gclk));
	jdff dff_A_TNod6VTT8_1(.dout(w_n140_0[1]),.din(w_dff_A_TNod6VTT8_1),.clk(gclk));
	jdff dff_A_NEG1lOOz2_1(.dout(w_dff_A_TNod6VTT8_1),.din(w_dff_A_NEG1lOOz2_1),.clk(gclk));
	jdff dff_A_dztB5kxU4_1(.dout(w_dff_A_NEG1lOOz2_1),.din(w_dff_A_dztB5kxU4_1),.clk(gclk));
	jdff dff_A_AbIXbCDW2_1(.dout(w_dff_A_dztB5kxU4_1),.din(w_dff_A_AbIXbCDW2_1),.clk(gclk));
	jdff dff_A_CdACMHy80_1(.dout(w_dff_A_AbIXbCDW2_1),.din(w_dff_A_CdACMHy80_1),.clk(gclk));
	jdff dff_A_XaNgq4Wh4_1(.dout(w_dff_A_CdACMHy80_1),.din(w_dff_A_XaNgq4Wh4_1),.clk(gclk));
	jdff dff_A_mUeoM9Ob8_1(.dout(G329gat),.din(w_dff_A_mUeoM9Ob8_1),.clk(gclk));
	jdff dff_A_r9qhEyp54_1(.dout(w_G115gat_0[1]),.din(w_dff_A_r9qhEyp54_1),.clk(gclk));
	jdff dff_A_32tvPrji5_1(.dout(w_dff_A_r9qhEyp54_1),.din(w_dff_A_32tvPrji5_1),.clk(gclk));
	jdff dff_A_G3h19LpY7_1(.dout(w_dff_A_32tvPrji5_1),.din(w_dff_A_G3h19LpY7_1),.clk(gclk));
	jdff dff_A_bzor4PHd8_1(.dout(w_dff_A_G3h19LpY7_1),.din(w_dff_A_bzor4PHd8_1),.clk(gclk));
	jdff dff_A_7bQosZHH0_1(.dout(w_dff_A_bzor4PHd8_1),.din(w_dff_A_7bQosZHH0_1),.clk(gclk));
	jdff dff_A_U1zaGshL6_1(.dout(w_dff_A_7bQosZHH0_1),.din(w_dff_A_U1zaGshL6_1),.clk(gclk));
	jdff dff_A_FWVp66n37_1(.dout(w_dff_A_U1zaGshL6_1),.din(w_dff_A_FWVp66n37_1),.clk(gclk));
	jdff dff_A_CnWadUpS6_1(.dout(w_dff_A_FWVp66n37_1),.din(w_dff_A_CnWadUpS6_1),.clk(gclk));
	jdff dff_A_eRHnONse6_1(.dout(w_dff_A_CnWadUpS6_1),.din(w_dff_A_eRHnONse6_1),.clk(gclk));
	jdff dff_A_yddNCP299_0(.dout(w_n222_0[0]),.din(w_dff_A_yddNCP299_0),.clk(gclk));
	jdff dff_A_GX7VCkeK6_0(.dout(w_dff_A_yddNCP299_0),.din(w_dff_A_GX7VCkeK6_0),.clk(gclk));
	jdff dff_A_CRZgAs995_0(.dout(w_dff_A_GX7VCkeK6_0),.din(w_dff_A_CRZgAs995_0),.clk(gclk));
	jdff dff_A_gmlFuxkv7_0(.dout(w_dff_A_CRZgAs995_0),.din(w_dff_A_gmlFuxkv7_0),.clk(gclk));
	jdff dff_A_ybgnrxKl4_0(.dout(w_dff_A_gmlFuxkv7_0),.din(w_dff_A_ybgnrxKl4_0),.clk(gclk));
	jdff dff_A_9qGbqOMD3_0(.dout(w_dff_A_ybgnrxKl4_0),.din(w_dff_A_9qGbqOMD3_0),.clk(gclk));
	jdff dff_A_SVFC7uqp2_0(.dout(w_dff_A_9qGbqOMD3_0),.din(w_dff_A_SVFC7uqp2_0),.clk(gclk));
	jdff dff_B_elRkFYIP3_0(.din(n134),.dout(w_dff_B_elRkFYIP3_0),.clk(gclk));
	jdff dff_A_jr1oo0Bk8_0(.dout(w_n130_0[0]),.din(w_dff_A_jr1oo0Bk8_0),.clk(gclk));
	jdff dff_A_JzKVPRA03_0(.dout(w_dff_A_jr1oo0Bk8_0),.din(w_dff_A_JzKVPRA03_0),.clk(gclk));
	jdff dff_A_OxTkNlyu5_0(.dout(w_dff_A_JzKVPRA03_0),.din(w_dff_A_OxTkNlyu5_0),.clk(gclk));
	jdff dff_A_e01KYA1J0_0(.dout(w_dff_A_OxTkNlyu5_0),.din(w_dff_A_e01KYA1J0_0),.clk(gclk));
	jdff dff_A_iJcbkrHa8_0(.dout(w_dff_A_e01KYA1J0_0),.din(w_dff_A_iJcbkrHa8_0),.clk(gclk));
	jdff dff_A_Yg723xQ76_0(.dout(w_n128_0[0]),.din(w_dff_A_Yg723xQ76_0),.clk(gclk));
	jdff dff_A_x56y1hzt5_0(.dout(w_dff_A_Yg723xQ76_0),.din(w_dff_A_x56y1hzt5_0),.clk(gclk));
	jdff dff_A_rKzxqIcD0_0(.dout(w_dff_A_x56y1hzt5_0),.din(w_dff_A_rKzxqIcD0_0),.clk(gclk));
	jdff dff_A_cGOhxaoR0_0(.dout(w_dff_A_rKzxqIcD0_0),.din(w_dff_A_cGOhxaoR0_0),.clk(gclk));
	jdff dff_A_5Rh6wsVC1_0(.dout(w_dff_A_cGOhxaoR0_0),.din(w_dff_A_5Rh6wsVC1_0),.clk(gclk));
	jdff dff_B_r3dWirN96_2(.din(n128),.dout(w_dff_B_r3dWirN96_2),.clk(gclk));
	jdff dff_B_LUhpJFK08_2(.din(w_dff_B_r3dWirN96_2),.dout(w_dff_B_LUhpJFK08_2),.clk(gclk));
	jdff dff_B_O78DKDEn3_2(.din(w_dff_B_LUhpJFK08_2),.dout(w_dff_B_O78DKDEn3_2),.clk(gclk));
	jdff dff_B_70Yd7APk8_2(.din(w_dff_B_O78DKDEn3_2),.dout(w_dff_B_70Yd7APk8_2),.clk(gclk));
	jdff dff_B_Zq05Emy40_2(.din(w_dff_B_70Yd7APk8_2),.dout(w_dff_B_Zq05Emy40_2),.clk(gclk));
	jdff dff_A_zAA0bolL9_0(.dout(w_G60gat_0[0]),.din(w_dff_A_zAA0bolL9_0),.clk(gclk));
	jdff dff_A_JVtt5KWv5_0(.dout(w_dff_A_zAA0bolL9_0),.din(w_dff_A_JVtt5KWv5_0),.clk(gclk));
	jdff dff_A_rIbykblP1_0(.dout(w_dff_A_JVtt5KWv5_0),.din(w_dff_A_rIbykblP1_0),.clk(gclk));
	jdff dff_A_AkIkxJsz1_0(.dout(w_dff_A_rIbykblP1_0),.din(w_dff_A_AkIkxJsz1_0),.clk(gclk));
	jdff dff_A_4IsB3gGg3_0(.dout(w_dff_A_AkIkxJsz1_0),.din(w_dff_A_4IsB3gGg3_0),.clk(gclk));
	jdff dff_A_HY3LHZsc6_0(.dout(w_dff_A_4IsB3gGg3_0),.din(w_dff_A_HY3LHZsc6_0),.clk(gclk));
	jdff dff_A_5S7pVowj7_0(.dout(w_dff_A_HY3LHZsc6_0),.din(w_dff_A_5S7pVowj7_0),.clk(gclk));
	jdff dff_A_2IOI8oZH0_0(.dout(w_dff_A_5S7pVowj7_0),.din(w_dff_A_2IOI8oZH0_0),.clk(gclk));
	jdff dff_A_4rivU3b73_1(.dout(w_G60gat_0[1]),.din(w_dff_A_4rivU3b73_1),.clk(gclk));
	jdff dff_A_ONgI4wLQ4_1(.dout(w_dff_A_4rivU3b73_1),.din(w_dff_A_ONgI4wLQ4_1),.clk(gclk));
	jdff dff_A_8VHJ7YhU7_1(.dout(w_dff_A_ONgI4wLQ4_1),.din(w_dff_A_8VHJ7YhU7_1),.clk(gclk));
	jdff dff_B_MKzUcZ2u5_1(.din(n124),.dout(w_dff_B_MKzUcZ2u5_1),.clk(gclk));
	jdff dff_B_T1RyiQcr6_1(.din(w_dff_B_MKzUcZ2u5_1),.dout(w_dff_B_T1RyiQcr6_1),.clk(gclk));
	jdff dff_B_4YMeAVOs6_1(.din(w_dff_B_T1RyiQcr6_1),.dout(w_dff_B_4YMeAVOs6_1),.clk(gclk));
	jdff dff_B_QxgWOeCq5_1(.din(w_dff_B_4YMeAVOs6_1),.dout(w_dff_B_QxgWOeCq5_1),.clk(gclk));
	jdff dff_B_yqZGaAPC1_1(.din(w_dff_B_QxgWOeCq5_1),.dout(w_dff_B_yqZGaAPC1_1),.clk(gclk));
	jdff dff_A_x0cHKmOc7_0(.dout(w_G99gat_0[0]),.din(w_dff_A_x0cHKmOc7_0),.clk(gclk));
	jdff dff_A_xhtGRUz96_0(.dout(w_dff_A_x0cHKmOc7_0),.din(w_dff_A_xhtGRUz96_0),.clk(gclk));
	jdff dff_A_5vld24Jq3_0(.dout(w_dff_A_xhtGRUz96_0),.din(w_dff_A_5vld24Jq3_0),.clk(gclk));
	jdff dff_A_OBS4fSpo0_0(.dout(w_dff_A_5vld24Jq3_0),.din(w_dff_A_OBS4fSpo0_0),.clk(gclk));
	jdff dff_A_vSfKcLNB9_0(.dout(w_dff_A_OBS4fSpo0_0),.din(w_dff_A_vSfKcLNB9_0),.clk(gclk));
	jdff dff_A_cdwrfuQp7_0(.dout(w_dff_A_vSfKcLNB9_0),.din(w_dff_A_cdwrfuQp7_0),.clk(gclk));
	jdff dff_A_TGiIRNbj6_0(.dout(w_dff_A_cdwrfuQp7_0),.din(w_dff_A_TGiIRNbj6_0),.clk(gclk));
	jdff dff_A_vyxp6Eid2_0(.dout(w_dff_A_TGiIRNbj6_0),.din(w_dff_A_vyxp6Eid2_0),.clk(gclk));
	jdff dff_A_ca0oEeB29_1(.dout(w_G99gat_0[1]),.din(w_dff_A_ca0oEeB29_1),.clk(gclk));
	jdff dff_A_JEyxBdAt4_1(.dout(w_dff_A_ca0oEeB29_1),.din(w_dff_A_JEyxBdAt4_1),.clk(gclk));
	jdff dff_A_tRoBYtPN0_1(.dout(w_dff_A_JEyxBdAt4_1),.din(w_dff_A_tRoBYtPN0_1),.clk(gclk));
	jdff dff_B_9XlDlqN57_1(.din(n120),.dout(w_dff_B_9XlDlqN57_1),.clk(gclk));
	jdff dff_B_fDBYCPLl7_1(.din(w_dff_B_9XlDlqN57_1),.dout(w_dff_B_fDBYCPLl7_1),.clk(gclk));
	jdff dff_B_IgVYzbtI3_1(.din(w_dff_B_fDBYCPLl7_1),.dout(w_dff_B_IgVYzbtI3_1),.clk(gclk));
	jdff dff_B_9uIeXScz6_1(.din(w_dff_B_IgVYzbtI3_1),.dout(w_dff_B_9uIeXScz6_1),.clk(gclk));
	jdff dff_B_YmnvNTO67_1(.din(w_dff_B_9uIeXScz6_1),.dout(w_dff_B_YmnvNTO67_1),.clk(gclk));
	jdff dff_A_iFzmUClZ2_0(.dout(w_G73gat_0[0]),.din(w_dff_A_iFzmUClZ2_0),.clk(gclk));
	jdff dff_A_Rtsu1nPa4_0(.dout(w_dff_A_iFzmUClZ2_0),.din(w_dff_A_Rtsu1nPa4_0),.clk(gclk));
	jdff dff_A_SLRSDd8X8_0(.dout(w_dff_A_Rtsu1nPa4_0),.din(w_dff_A_SLRSDd8X8_0),.clk(gclk));
	jdff dff_A_TfTh3ZeS9_0(.dout(w_dff_A_SLRSDd8X8_0),.din(w_dff_A_TfTh3ZeS9_0),.clk(gclk));
	jdff dff_A_2M3cQGbu2_0(.dout(w_dff_A_TfTh3ZeS9_0),.din(w_dff_A_2M3cQGbu2_0),.clk(gclk));
	jdff dff_A_G1e9RZwv5_0(.dout(w_dff_A_2M3cQGbu2_0),.din(w_dff_A_G1e9RZwv5_0),.clk(gclk));
	jdff dff_A_CEPNZffk8_0(.dout(w_dff_A_G1e9RZwv5_0),.din(w_dff_A_CEPNZffk8_0),.clk(gclk));
	jdff dff_A_uC2MoJHC9_0(.dout(w_dff_A_CEPNZffk8_0),.din(w_dff_A_uC2MoJHC9_0),.clk(gclk));
	jdff dff_A_MiHGDkhu9_0(.dout(w_n116_0[0]),.din(w_dff_A_MiHGDkhu9_0),.clk(gclk));
	jdff dff_A_n4B4x9c09_0(.dout(w_dff_A_MiHGDkhu9_0),.din(w_dff_A_n4B4x9c09_0),.clk(gclk));
	jdff dff_A_a13WHX4j7_0(.dout(w_dff_A_n4B4x9c09_0),.din(w_dff_A_a13WHX4j7_0),.clk(gclk));
	jdff dff_A_icucMoCM1_0(.dout(w_dff_A_a13WHX4j7_0),.din(w_dff_A_icucMoCM1_0),.clk(gclk));
	jdff dff_A_lrvoPlfa9_0(.dout(w_dff_A_icucMoCM1_0),.din(w_dff_A_lrvoPlfa9_0),.clk(gclk));
	jdff dff_A_ANjHGxGf8_0(.dout(w_n114_0[0]),.din(w_dff_A_ANjHGxGf8_0),.clk(gclk));
	jdff dff_A_FwTY1rTi7_0(.dout(w_dff_A_ANjHGxGf8_0),.din(w_dff_A_FwTY1rTi7_0),.clk(gclk));
	jdff dff_A_eCiT5ni34_0(.dout(w_dff_A_FwTY1rTi7_0),.din(w_dff_A_eCiT5ni34_0),.clk(gclk));
	jdff dff_A_ukKvqtB41_0(.dout(w_dff_A_eCiT5ni34_0),.din(w_dff_A_ukKvqtB41_0),.clk(gclk));
	jdff dff_A_OUBJK5dB4_0(.dout(w_dff_A_ukKvqtB41_0),.din(w_dff_A_OUBJK5dB4_0),.clk(gclk));
	jdff dff_B_7ACDJUSU9_2(.din(n114),.dout(w_dff_B_7ACDJUSU9_2),.clk(gclk));
	jdff dff_B_JxN8MC734_2(.din(w_dff_B_7ACDJUSU9_2),.dout(w_dff_B_JxN8MC734_2),.clk(gclk));
	jdff dff_B_6EjmAgtR4_2(.din(w_dff_B_JxN8MC734_2),.dout(w_dff_B_6EjmAgtR4_2),.clk(gclk));
	jdff dff_B_rq4XUosw7_2(.din(w_dff_B_6EjmAgtR4_2),.dout(w_dff_B_rq4XUosw7_2),.clk(gclk));
	jdff dff_B_GZI4eWWi3_2(.din(w_dff_B_rq4XUosw7_2),.dout(w_dff_B_GZI4eWWi3_2),.clk(gclk));
	jdff dff_A_j3XIiRRK8_0(.dout(w_G86gat_0[0]),.din(w_dff_A_j3XIiRRK8_0),.clk(gclk));
	jdff dff_A_dPiO0LtP4_0(.dout(w_dff_A_j3XIiRRK8_0),.din(w_dff_A_dPiO0LtP4_0),.clk(gclk));
	jdff dff_A_yin4GHKJ1_0(.dout(w_dff_A_dPiO0LtP4_0),.din(w_dff_A_yin4GHKJ1_0),.clk(gclk));
	jdff dff_A_F264yvlv0_0(.dout(w_dff_A_yin4GHKJ1_0),.din(w_dff_A_F264yvlv0_0),.clk(gclk));
	jdff dff_A_Zvw3Jmy07_0(.dout(w_dff_A_F264yvlv0_0),.din(w_dff_A_Zvw3Jmy07_0),.clk(gclk));
	jdff dff_A_GXzQ2Qv23_0(.dout(w_dff_A_Zvw3Jmy07_0),.din(w_dff_A_GXzQ2Qv23_0),.clk(gclk));
	jdff dff_A_nbwRWgXO1_0(.dout(w_dff_A_GXzQ2Qv23_0),.din(w_dff_A_nbwRWgXO1_0),.clk(gclk));
	jdff dff_A_CNjBBjIk4_0(.dout(w_dff_A_nbwRWgXO1_0),.din(w_dff_A_CNjBBjIk4_0),.clk(gclk));
	jdff dff_A_BdrKwSXp0_1(.dout(w_G86gat_0[1]),.din(w_dff_A_BdrKwSXp0_1),.clk(gclk));
	jdff dff_A_zcxX3cwF7_1(.dout(w_dff_A_BdrKwSXp0_1),.din(w_dff_A_zcxX3cwF7_1),.clk(gclk));
	jdff dff_A_jIh8pKnM9_1(.dout(w_dff_A_zcxX3cwF7_1),.din(w_dff_A_jIh8pKnM9_1),.clk(gclk));
	jdff dff_A_3xsKJLd08_0(.dout(w_n112_0[0]),.din(w_dff_A_3xsKJLd08_0),.clk(gclk));
	jdff dff_A_RX6PzHag1_0(.dout(w_dff_A_3xsKJLd08_0),.din(w_dff_A_RX6PzHag1_0),.clk(gclk));
	jdff dff_A_YwlIeDW40_0(.dout(w_dff_A_RX6PzHag1_0),.din(w_dff_A_YwlIeDW40_0),.clk(gclk));
	jdff dff_A_1U80RyWS9_0(.dout(w_dff_A_YwlIeDW40_0),.din(w_dff_A_1U80RyWS9_0),.clk(gclk));
	jdff dff_A_kRjQN2Aa7_0(.dout(w_dff_A_1U80RyWS9_0),.din(w_dff_A_kRjQN2Aa7_0),.clk(gclk));
	jdff dff_A_c2egbizS7_0(.dout(w_n110_0[0]),.din(w_dff_A_c2egbizS7_0),.clk(gclk));
	jdff dff_A_As2HewtW1_0(.dout(w_dff_A_c2egbizS7_0),.din(w_dff_A_As2HewtW1_0),.clk(gclk));
	jdff dff_A_9BCtItK83_0(.dout(w_dff_A_As2HewtW1_0),.din(w_dff_A_9BCtItK83_0),.clk(gclk));
	jdff dff_A_Exk40fx50_0(.dout(w_dff_A_9BCtItK83_0),.din(w_dff_A_Exk40fx50_0),.clk(gclk));
	jdff dff_A_TYl7dF2w3_0(.dout(w_dff_A_Exk40fx50_0),.din(w_dff_A_TYl7dF2w3_0),.clk(gclk));
	jdff dff_B_V8hG2G8G4_2(.din(n110),.dout(w_dff_B_V8hG2G8G4_2),.clk(gclk));
	jdff dff_B_CzZGeQ8i5_2(.din(w_dff_B_V8hG2G8G4_2),.dout(w_dff_B_CzZGeQ8i5_2),.clk(gclk));
	jdff dff_B_v0sDIqxd3_2(.din(w_dff_B_CzZGeQ8i5_2),.dout(w_dff_B_v0sDIqxd3_2),.clk(gclk));
	jdff dff_B_8SX2Digw1_2(.din(w_dff_B_v0sDIqxd3_2),.dout(w_dff_B_8SX2Digw1_2),.clk(gclk));
	jdff dff_B_HmDgpTZ25_2(.din(w_dff_B_8SX2Digw1_2),.dout(w_dff_B_HmDgpTZ25_2),.clk(gclk));
	jdff dff_A_dkeOH2Ow1_0(.dout(w_G34gat_0[0]),.din(w_dff_A_dkeOH2Ow1_0),.clk(gclk));
	jdff dff_A_JUSfIm3S8_0(.dout(w_dff_A_dkeOH2Ow1_0),.din(w_dff_A_JUSfIm3S8_0),.clk(gclk));
	jdff dff_A_S9xMJYHP2_0(.dout(w_dff_A_JUSfIm3S8_0),.din(w_dff_A_S9xMJYHP2_0),.clk(gclk));
	jdff dff_A_wU5caEIS7_0(.dout(w_dff_A_S9xMJYHP2_0),.din(w_dff_A_wU5caEIS7_0),.clk(gclk));
	jdff dff_A_y0bfCXbb4_0(.dout(w_dff_A_wU5caEIS7_0),.din(w_dff_A_y0bfCXbb4_0),.clk(gclk));
	jdff dff_A_DwLkY97D5_0(.dout(w_dff_A_y0bfCXbb4_0),.din(w_dff_A_DwLkY97D5_0),.clk(gclk));
	jdff dff_A_mINrjOlD6_0(.dout(w_dff_A_DwLkY97D5_0),.din(w_dff_A_mINrjOlD6_0),.clk(gclk));
	jdff dff_A_JCeut76T7_0(.dout(w_dff_A_mINrjOlD6_0),.din(w_dff_A_JCeut76T7_0),.clk(gclk));
	jdff dff_A_xRuxKaBe1_1(.dout(w_G34gat_0[1]),.din(w_dff_A_xRuxKaBe1_1),.clk(gclk));
	jdff dff_A_pN0jcjOr6_1(.dout(w_dff_A_xRuxKaBe1_1),.din(w_dff_A_pN0jcjOr6_1),.clk(gclk));
	jdff dff_A_tqGg37gq2_1(.dout(w_dff_A_pN0jcjOr6_1),.din(w_dff_A_tqGg37gq2_1),.clk(gclk));
	jdff dff_A_SdRqIHRY4_0(.dout(w_n105_0[0]),.din(w_dff_A_SdRqIHRY4_0),.clk(gclk));
	jdff dff_A_Oiv6w4kd5_0(.dout(w_dff_A_SdRqIHRY4_0),.din(w_dff_A_Oiv6w4kd5_0),.clk(gclk));
	jdff dff_A_M23sTneE8_0(.dout(w_dff_A_Oiv6w4kd5_0),.din(w_dff_A_M23sTneE8_0),.clk(gclk));
	jdff dff_A_iYp5DQIc1_0(.dout(w_dff_A_M23sTneE8_0),.din(w_dff_A_iYp5DQIc1_0),.clk(gclk));
	jdff dff_A_IGLEGmrh9_0(.dout(w_dff_A_iYp5DQIc1_0),.din(w_dff_A_IGLEGmrh9_0),.clk(gclk));
	jdff dff_B_jvnGzxqi9_2(.din(n105),.dout(w_dff_B_jvnGzxqi9_2),.clk(gclk));
	jdff dff_B_VVqurd5k9_2(.din(w_dff_B_jvnGzxqi9_2),.dout(w_dff_B_VVqurd5k9_2),.clk(gclk));
	jdff dff_B_mSkxwXQh3_2(.din(w_dff_B_VVqurd5k9_2),.dout(w_dff_B_mSkxwXQh3_2),.clk(gclk));
	jdff dff_B_t3CuSTtI6_2(.din(w_dff_B_mSkxwXQh3_2),.dout(w_dff_B_t3CuSTtI6_2),.clk(gclk));
	jdff dff_B_AmzplG4U7_2(.din(w_dff_B_t3CuSTtI6_2),.dout(w_dff_B_AmzplG4U7_2),.clk(gclk));
	jdff dff_A_9Oywq3Cy4_0(.dout(w_G8gat_0[0]),.din(w_dff_A_9Oywq3Cy4_0),.clk(gclk));
	jdff dff_A_qYC8OLbf3_0(.dout(w_dff_A_9Oywq3Cy4_0),.din(w_dff_A_qYC8OLbf3_0),.clk(gclk));
	jdff dff_A_y5FkzdAj6_0(.dout(w_dff_A_qYC8OLbf3_0),.din(w_dff_A_y5FkzdAj6_0),.clk(gclk));
	jdff dff_A_MpICS6oG9_1(.dout(w_G8gat_0[1]),.din(w_dff_A_MpICS6oG9_1),.clk(gclk));
	jdff dff_A_i3PKVHDZ8_1(.dout(w_dff_A_MpICS6oG9_1),.din(w_dff_A_i3PKVHDZ8_1),.clk(gclk));
	jdff dff_A_QLE8tMgA9_1(.dout(w_dff_A_i3PKVHDZ8_1),.din(w_dff_A_QLE8tMgA9_1),.clk(gclk));
	jdff dff_A_PWpSrhra2_1(.dout(w_dff_A_QLE8tMgA9_1),.din(w_dff_A_PWpSrhra2_1),.clk(gclk));
	jdff dff_A_3iguwmxU7_1(.dout(w_dff_A_PWpSrhra2_1),.din(w_dff_A_3iguwmxU7_1),.clk(gclk));
	jdff dff_A_XHiXL1vT3_1(.dout(w_dff_A_3iguwmxU7_1),.din(w_dff_A_XHiXL1vT3_1),.clk(gclk));
	jdff dff_A_7szbMaJP7_1(.dout(w_dff_A_XHiXL1vT3_1),.din(w_dff_A_7szbMaJP7_1),.clk(gclk));
	jdff dff_A_nIaoEFj81_1(.dout(w_dff_A_7szbMaJP7_1),.din(w_dff_A_nIaoEFj81_1),.clk(gclk));
	jdff dff_A_Fn5wJJxq9_0(.dout(w_n101_0[0]),.din(w_dff_A_Fn5wJJxq9_0),.clk(gclk));
	jdff dff_A_yk1twS921_0(.dout(w_dff_A_Fn5wJJxq9_0),.din(w_dff_A_yk1twS921_0),.clk(gclk));
	jdff dff_A_r7uKwLKa2_0(.dout(w_dff_A_yk1twS921_0),.din(w_dff_A_r7uKwLKa2_0),.clk(gclk));
	jdff dff_A_m7iU58na4_0(.dout(w_dff_A_r7uKwLKa2_0),.din(w_dff_A_m7iU58na4_0),.clk(gclk));
	jdff dff_A_D4DlJhkB5_0(.dout(w_dff_A_m7iU58na4_0),.din(w_dff_A_D4DlJhkB5_0),.clk(gclk));
	jdff dff_B_wbf1ntPr9_2(.din(n101),.dout(w_dff_B_wbf1ntPr9_2),.clk(gclk));
	jdff dff_B_bK0v1cy11_2(.din(w_dff_B_wbf1ntPr9_2),.dout(w_dff_B_bK0v1cy11_2),.clk(gclk));
	jdff dff_B_NqZ5Jgx63_2(.din(w_dff_B_bK0v1cy11_2),.dout(w_dff_B_NqZ5Jgx63_2),.clk(gclk));
	jdff dff_B_DWRYHzfE4_2(.din(w_dff_B_NqZ5Jgx63_2),.dout(w_dff_B_DWRYHzfE4_2),.clk(gclk));
	jdff dff_B_vSYbKYBY4_2(.din(w_dff_B_DWRYHzfE4_2),.dout(w_dff_B_vSYbKYBY4_2),.clk(gclk));
	jdff dff_A_FKtEcpHY6_0(.dout(w_G21gat_0[0]),.din(w_dff_A_FKtEcpHY6_0),.clk(gclk));
	jdff dff_A_adsLzTVN6_0(.dout(w_dff_A_FKtEcpHY6_0),.din(w_dff_A_adsLzTVN6_0),.clk(gclk));
	jdff dff_A_d7sPam9L9_0(.dout(w_dff_A_adsLzTVN6_0),.din(w_dff_A_d7sPam9L9_0),.clk(gclk));
	jdff dff_A_iHxyBWcY6_0(.dout(w_dff_A_d7sPam9L9_0),.din(w_dff_A_iHxyBWcY6_0),.clk(gclk));
	jdff dff_A_5wssdGa09_0(.dout(w_dff_A_iHxyBWcY6_0),.din(w_dff_A_5wssdGa09_0),.clk(gclk));
	jdff dff_A_7xa6gGTi5_0(.dout(w_dff_A_5wssdGa09_0),.din(w_dff_A_7xa6gGTi5_0),.clk(gclk));
	jdff dff_A_QF3EaDNk1_0(.dout(w_dff_A_7xa6gGTi5_0),.din(w_dff_A_QF3EaDNk1_0),.clk(gclk));
	jdff dff_A_LWwWd2XP2_0(.dout(w_dff_A_QF3EaDNk1_0),.din(w_dff_A_LWwWd2XP2_0),.clk(gclk));
	jdff dff_A_nPHp5ejD7_1(.dout(w_G21gat_0[1]),.din(w_dff_A_nPHp5ejD7_1),.clk(gclk));
	jdff dff_A_mKSXXTUt3_1(.dout(w_dff_A_nPHp5ejD7_1),.din(w_dff_A_mKSXXTUt3_1),.clk(gclk));
	jdff dff_A_GHQIdJ3A2_1(.dout(w_dff_A_mKSXXTUt3_1),.din(w_dff_A_GHQIdJ3A2_1),.clk(gclk));
	jdff dff_B_1Dqoumz57_0(.din(n99),.dout(w_dff_B_1Dqoumz57_0),.clk(gclk));
	jdff dff_B_cbdoMM8D3_0(.din(w_dff_B_1Dqoumz57_0),.dout(w_dff_B_cbdoMM8D3_0),.clk(gclk));
	jdff dff_B_Uk8EdMHU4_0(.din(w_dff_B_cbdoMM8D3_0),.dout(w_dff_B_Uk8EdMHU4_0),.clk(gclk));
	jdff dff_B_nGVCPjFW1_1(.din(n95),.dout(w_dff_B_nGVCPjFW1_1),.clk(gclk));
	jdff dff_B_sggIiMAn0_1(.din(w_dff_B_nGVCPjFW1_1),.dout(w_dff_B_sggIiMAn0_1),.clk(gclk));
	jdff dff_B_zObk1IBb7_1(.din(w_dff_B_sggIiMAn0_1),.dout(w_dff_B_zObk1IBb7_1),.clk(gclk));
	jdff dff_A_Fy60x3P36_0(.dout(w_n97_0[0]),.din(w_dff_A_Fy60x3P36_0),.clk(gclk));
	jdff dff_A_Yi5W6JXN6_0(.dout(w_dff_A_Fy60x3P36_0),.din(w_dff_A_Yi5W6JXN6_0),.clk(gclk));
	jdff dff_A_soVg1WKJ3_0(.dout(w_dff_A_Yi5W6JXN6_0),.din(w_dff_A_soVg1WKJ3_0),.clk(gclk));
	jdff dff_A_IQMaiIy48_0(.dout(w_dff_A_soVg1WKJ3_0),.din(w_dff_A_IQMaiIy48_0),.clk(gclk));
	jdff dff_A_SBG7leFx0_0(.dout(w_dff_A_IQMaiIy48_0),.din(w_dff_A_SBG7leFx0_0),.clk(gclk));
	jdff dff_A_K04cbamz3_0(.dout(w_dff_A_SBG7leFx0_0),.din(w_dff_A_K04cbamz3_0),.clk(gclk));
	jdff dff_A_W326EnfZ9_2(.dout(G223gat),.din(w_dff_A_W326EnfZ9_2),.clk(gclk));
	jdff dff_A_99OEwyVj8_0(.dout(w_G112gat_0[0]),.din(w_dff_A_99OEwyVj8_0),.clk(gclk));
	jdff dff_A_TO0pI6pW4_0(.dout(w_dff_A_99OEwyVj8_0),.din(w_dff_A_TO0pI6pW4_0),.clk(gclk));
	jdff dff_A_uVAAnEkd7_0(.dout(w_dff_A_TO0pI6pW4_0),.din(w_dff_A_uVAAnEkd7_0),.clk(gclk));
	jdff dff_A_TQqw1IkZ8_0(.dout(w_dff_A_uVAAnEkd7_0),.din(w_dff_A_TQqw1IkZ8_0),.clk(gclk));
	jdff dff_A_mVDjpnBy0_0(.dout(w_dff_A_TQqw1IkZ8_0),.din(w_dff_A_mVDjpnBy0_0),.clk(gclk));
	jdff dff_A_lDalHZ6U6_0(.dout(w_dff_A_mVDjpnBy0_0),.din(w_dff_A_lDalHZ6U6_0),.clk(gclk));
	jdff dff_A_rtpVrcs98_0(.dout(w_dff_A_lDalHZ6U6_0),.din(w_dff_A_rtpVrcs98_0),.clk(gclk));
	jdff dff_A_gbQT9wQ18_0(.dout(w_dff_A_rtpVrcs98_0),.din(w_dff_A_gbQT9wQ18_0),.clk(gclk));
	jdff dff_B_Cm1a5uJJ0_1(.din(n71),.dout(w_dff_B_Cm1a5uJJ0_1),.clk(gclk));
	jdff dff_B_BEEiQtjO1_1(.din(w_dff_B_Cm1a5uJJ0_1),.dout(w_dff_B_BEEiQtjO1_1),.clk(gclk));
	jdff dff_B_b1qlV9oy7_1(.din(w_dff_B_BEEiQtjO1_1),.dout(w_dff_B_b1qlV9oy7_1),.clk(gclk));
	jdff dff_B_lGP9RFp44_1(.din(w_dff_B_b1qlV9oy7_1),.dout(w_dff_B_lGP9RFp44_1),.clk(gclk));
	jdff dff_B_OhC3PUo71_1(.din(w_dff_B_lGP9RFp44_1),.dout(w_dff_B_OhC3PUo71_1),.clk(gclk));
	jdff dff_B_gX41heb25_1(.din(w_dff_B_OhC3PUo71_1),.dout(w_dff_B_gX41heb25_1),.clk(gclk));
	jdff dff_B_1xpyi4966_1(.din(n72),.dout(w_dff_B_1xpyi4966_1),.clk(gclk));
	jdff dff_A_MbQKfbsk6_0(.dout(w_n86_0[0]),.din(w_dff_A_MbQKfbsk6_0),.clk(gclk));
	jdff dff_A_rqzoA0Ia7_0(.dout(w_dff_A_MbQKfbsk6_0),.din(w_dff_A_rqzoA0Ia7_0),.clk(gclk));
	jdff dff_A_yHkvwQj01_0(.dout(w_n81_0[0]),.din(w_dff_A_yHkvwQj01_0),.clk(gclk));
	jdff dff_A_2K2yrrM81_0(.dout(w_n80_0[0]),.din(w_dff_A_2K2yrrM81_0),.clk(gclk));
	jdff dff_A_nrNMB1Qw2_0(.dout(w_dff_A_2K2yrrM81_0),.din(w_dff_A_nrNMB1Qw2_0),.clk(gclk));
	jdff dff_A_UkW8ZDk14_0(.dout(w_n75_0[0]),.din(w_dff_A_UkW8ZDk14_0),.clk(gclk));
	jdff dff_A_SEUXUfo07_0(.dout(w_dff_A_UkW8ZDk14_0),.din(w_dff_A_SEUXUfo07_0),.clk(gclk));
	jdff dff_A_uMW9eypZ3_0(.dout(w_n73_0[0]),.din(w_dff_A_uMW9eypZ3_0),.clk(gclk));
	jdff dff_A_FZXMCCaU2_0(.dout(w_dff_A_uMW9eypZ3_0),.din(w_dff_A_FZXMCCaU2_0),.clk(gclk));
	jdff dff_A_8D4StsrM8_0(.dout(w_G47gat_0[0]),.din(w_dff_A_8D4StsrM8_0),.clk(gclk));
	jdff dff_A_7ScH9M6S5_0(.dout(w_dff_A_8D4StsrM8_0),.din(w_dff_A_7ScH9M6S5_0),.clk(gclk));
	jdff dff_A_zQPleNJo0_0(.dout(w_dff_A_7ScH9M6S5_0),.din(w_dff_A_zQPleNJo0_0),.clk(gclk));
	jdff dff_A_mzmXnC9F9_0(.dout(w_dff_A_zQPleNJo0_0),.din(w_dff_A_mzmXnC9F9_0),.clk(gclk));
	jdff dff_A_vDActhM91_0(.dout(w_dff_A_mzmXnC9F9_0),.din(w_dff_A_vDActhM91_0),.clk(gclk));
	jdff dff_A_P2mQQYsi8_0(.dout(w_dff_A_vDActhM91_0),.din(w_dff_A_P2mQQYsi8_0),.clk(gclk));
	jdff dff_A_hiserwzi4_0(.dout(w_dff_A_P2mQQYsi8_0),.din(w_dff_A_hiserwzi4_0),.clk(gclk));
	jdff dff_A_t1cFit3B7_0(.dout(w_dff_A_hiserwzi4_0),.din(w_dff_A_t1cFit3B7_0),.clk(gclk));
	jdff dff_A_baWLntZs7_0(.dout(w_n151_0[0]),.din(w_dff_A_baWLntZs7_0),.clk(gclk));
	jdff dff_A_8xi9B3wd0_0(.dout(w_dff_A_baWLntZs7_0),.din(w_dff_A_8xi9B3wd0_0),.clk(gclk));
	jdff dff_A_tA2X8DgX2_0(.dout(w_dff_A_8xi9B3wd0_0),.din(w_dff_A_tA2X8DgX2_0),.clk(gclk));
	jdff dff_A_pisgjtVx6_0(.dout(w_dff_A_tA2X8DgX2_0),.din(w_dff_A_pisgjtVx6_0),.clk(gclk));
	jdff dff_A_FvT8uCGY0_0(.dout(w_dff_A_pisgjtVx6_0),.din(w_dff_A_FvT8uCGY0_0),.clk(gclk));
	jdff dff_A_K44bNDl21_0(.dout(w_dff_A_FvT8uCGY0_0),.din(w_dff_A_K44bNDl21_0),.clk(gclk));
	jdff dff_A_SR1ejsZM8_0(.dout(w_G4gat_0[0]),.din(w_dff_A_SR1ejsZM8_0),.clk(gclk));
	jdff dff_A_JYgXQKqk1_0(.dout(w_dff_A_SR1ejsZM8_0),.din(w_dff_A_JYgXQKqk1_0),.clk(gclk));
	jdff dff_A_Nz4sdyYA2_0(.dout(w_dff_A_JYgXQKqk1_0),.din(w_dff_A_Nz4sdyYA2_0),.clk(gclk));
	jdff dff_A_GcwJnUIe9_0(.dout(w_dff_A_Nz4sdyYA2_0),.din(w_dff_A_GcwJnUIe9_0),.clk(gclk));
	jdff dff_A_sNF0DQIE1_0(.dout(w_dff_A_GcwJnUIe9_0),.din(w_dff_A_sNF0DQIE1_0),.clk(gclk));
	jdff dff_A_EAGYtwR70_2(.dout(w_G4gat_0[2]),.din(w_dff_A_EAGYtwR70_2),.clk(gclk));
	jdff dff_A_1nWO7iXq1_0(.dout(w_n65_0[0]),.din(w_dff_A_1nWO7iXq1_0),.clk(gclk));
	jdff dff_A_W0uqm6yX6_0(.dout(w_dff_A_1nWO7iXq1_0),.din(w_dff_A_W0uqm6yX6_0),.clk(gclk));
	jdff dff_A_JrjeQhYS0_0(.dout(w_dff_A_W0uqm6yX6_0),.din(w_dff_A_JrjeQhYS0_0),.clk(gclk));
	jdff dff_A_ieyc2s8R4_0(.dout(w_dff_A_JrjeQhYS0_0),.din(w_dff_A_ieyc2s8R4_0),.clk(gclk));
	jdff dff_A_Oy1yKkZC3_0(.dout(w_G1gat_0[0]),.din(w_dff_A_Oy1yKkZC3_0),.clk(gclk));
	jdff dff_A_iQYLfxpb5_0(.dout(w_dff_A_Oy1yKkZC3_0),.din(w_dff_A_iQYLfxpb5_0),.clk(gclk));
	jdff dff_A_ZYoviDPY0_1(.dout(w_G1gat_0[1]),.din(w_dff_A_ZYoviDPY0_1),.clk(gclk));
	jdff dff_A_FlQoilbD1_0(.dout(w_n63_0[0]),.din(w_dff_A_FlQoilbD1_0),.clk(gclk));
	jdff dff_A_SPW8OOyW2_0(.dout(w_dff_A_FlQoilbD1_0),.din(w_dff_A_SPW8OOyW2_0),.clk(gclk));
	jdff dff_A_9hkp6sgQ4_0(.dout(w_dff_A_SPW8OOyW2_0),.din(w_dff_A_9hkp6sgQ4_0),.clk(gclk));
	jdff dff_A_0YvkzvW76_0(.dout(w_dff_A_9hkp6sgQ4_0),.din(w_dff_A_0YvkzvW76_0),.clk(gclk));
	jdff dff_A_4PQy5beG8_0(.dout(w_G24gat_0[0]),.din(w_dff_A_4PQy5beG8_0),.clk(gclk));
	jdff dff_A_Cr2ZkKXQ4_0(.dout(w_dff_A_4PQy5beG8_0),.din(w_dff_A_Cr2ZkKXQ4_0),.clk(gclk));
	jdff dff_A_yt9M3IUb6_1(.dout(w_G24gat_0[1]),.din(w_dff_A_yt9M3IUb6_1),.clk(gclk));
	jdff dff_A_pfh2nmvF3_0(.dout(w_n61_0[0]),.din(w_dff_A_pfh2nmvF3_0),.clk(gclk));
	jdff dff_A_V7Khcg9C9_0(.dout(w_n60_0[0]),.din(w_dff_A_V7Khcg9C9_0),.clk(gclk));
	jdff dff_A_7RPd38vW4_0(.dout(w_dff_A_V7Khcg9C9_0),.din(w_dff_A_7RPd38vW4_0),.clk(gclk));
	jdff dff_A_58oV52wE8_0(.dout(w_G102gat_0[0]),.din(w_dff_A_58oV52wE8_0),.clk(gclk));
	jdff dff_B_afx5LJw82_2(.din(G102gat),.dout(w_dff_B_afx5LJw82_2),.clk(gclk));
	jdff dff_A_oSmuBXq48_0(.dout(w_n57_0[0]),.din(w_dff_A_oSmuBXq48_0),.clk(gclk));
	jdff dff_A_UuzPBemQ3_0(.dout(w_dff_A_oSmuBXq48_0),.din(w_dff_A_UuzPBemQ3_0),.clk(gclk));
	jdff dff_A_Nufseag98_0(.dout(w_dff_A_UuzPBemQ3_0),.din(w_dff_A_Nufseag98_0),.clk(gclk));
	jdff dff_A_82RAgkJH2_0(.dout(w_G43gat_0[0]),.din(w_dff_A_82RAgkJH2_0),.clk(gclk));
	jdff dff_A_krz4KfgE3_0(.dout(w_dff_A_82RAgkJH2_0),.din(w_dff_A_krz4KfgE3_0),.clk(gclk));
	jdff dff_A_I7kKsBev3_0(.dout(w_dff_A_krz4KfgE3_0),.din(w_dff_A_I7kKsBev3_0),.clk(gclk));
	jdff dff_A_LYsOicH60_0(.dout(w_dff_A_I7kKsBev3_0),.din(w_dff_A_LYsOicH60_0),.clk(gclk));
	jdff dff_A_GsuKMg6o3_0(.dout(w_dff_A_LYsOicH60_0),.din(w_dff_A_GsuKMg6o3_0),.clk(gclk));
	jdff dff_A_GEAeV8tI5_0(.dout(w_dff_A_GsuKMg6o3_0),.din(w_dff_A_GEAeV8tI5_0),.clk(gclk));
	jdff dff_A_0SWsR2jh0_2(.dout(w_G43gat_0[2]),.din(w_dff_A_0SWsR2jh0_2),.clk(gclk));
	jdff dff_A_beQQhK370_0(.dout(w_G37gat_0[0]),.din(w_dff_A_beQQhK370_0),.clk(gclk));
	jdff dff_A_E34v5w1D8_0(.dout(w_G69gat_0[0]),.din(w_dff_A_E34v5w1D8_0),.clk(gclk));
	jdff dff_A_bH46gdET4_0(.dout(w_dff_A_E34v5w1D8_0),.din(w_dff_A_bH46gdET4_0),.clk(gclk));
	jdff dff_A_XWRn0zpj8_0(.dout(w_dff_A_bH46gdET4_0),.din(w_dff_A_XWRn0zpj8_0),.clk(gclk));
	jdff dff_A_w0s2IWhd5_0(.dout(w_dff_A_XWRn0zpj8_0),.din(w_dff_A_w0s2IWhd5_0),.clk(gclk));
	jdff dff_A_s7ajoNiA4_0(.dout(w_dff_A_w0s2IWhd5_0),.din(w_dff_A_s7ajoNiA4_0),.clk(gclk));
	jdff dff_A_waCCqaoY2_2(.dout(w_G69gat_0[2]),.din(w_dff_A_waCCqaoY2_2),.clk(gclk));
	jdff dff_A_CZRt8b9D0_0(.dout(w_n54_0[0]),.din(w_dff_A_CZRt8b9D0_0),.clk(gclk));
	jdff dff_A_nSpv3FJ57_0(.dout(w_dff_A_CZRt8b9D0_0),.din(w_dff_A_nSpv3FJ57_0),.clk(gclk));
	jdff dff_A_KDP78WSH1_0(.dout(w_dff_A_nSpv3FJ57_0),.din(w_dff_A_KDP78WSH1_0),.clk(gclk));
	jdff dff_A_xpJgvIew4_0(.dout(w_dff_A_KDP78WSH1_0),.din(w_dff_A_xpJgvIew4_0),.clk(gclk));
	jdff dff_A_kLmahsAr0_0(.dout(w_G63gat_0[0]),.din(w_dff_A_kLmahsAr0_0),.clk(gclk));
	jdff dff_A_HuGCCWpH6_0(.dout(w_G95gat_0[0]),.din(w_dff_A_HuGCCWpH6_0),.clk(gclk));
	jdff dff_A_irsMUWDd8_0(.dout(w_dff_A_HuGCCWpH6_0),.din(w_dff_A_irsMUWDd8_0),.clk(gclk));
	jdff dff_A_KIvKVHvM3_0(.dout(w_dff_A_irsMUWDd8_0),.din(w_dff_A_KIvKVHvM3_0),.clk(gclk));
	jdff dff_A_GYjoS2KM5_0(.dout(w_dff_A_KIvKVHvM3_0),.din(w_dff_A_GYjoS2KM5_0),.clk(gclk));
	jdff dff_A_ON2lZaPN2_0(.dout(w_dff_A_GYjoS2KM5_0),.din(w_dff_A_ON2lZaPN2_0),.clk(gclk));
	jdff dff_A_dZMPz4bJ0_2(.dout(w_G95gat_0[2]),.din(w_dff_A_dZMPz4bJ0_2),.clk(gclk));
	jdff dff_A_1JuT8rBx3_0(.dout(w_n51_0[0]),.din(w_dff_A_1JuT8rBx3_0),.clk(gclk));
	jdff dff_A_XRbHuvV03_0(.dout(w_dff_A_1JuT8rBx3_0),.din(w_dff_A_XRbHuvV03_0),.clk(gclk));
	jdff dff_A_ouUnLuhN5_0(.dout(w_dff_A_XRbHuvV03_0),.din(w_dff_A_ouUnLuhN5_0),.clk(gclk));
	jdff dff_A_q1Qym2jm8_0(.dout(w_dff_A_ouUnLuhN5_0),.din(w_dff_A_q1Qym2jm8_0),.clk(gclk));
	jdff dff_A_ag0BdDFt3_0(.dout(w_G89gat_0[0]),.din(w_dff_A_ag0BdDFt3_0),.clk(gclk));
	jdff dff_A_vBRpqx6P4_0(.dout(w_dff_A_ag0BdDFt3_0),.din(w_dff_A_vBRpqx6P4_0),.clk(gclk));
	jdff dff_A_AFfuu5bo6_1(.dout(w_G89gat_0[1]),.din(w_dff_A_AFfuu5bo6_1),.clk(gclk));
	jdff dff_A_Jlef4EEs7_0(.dout(w_G56gat_0[0]),.din(w_dff_A_Jlef4EEs7_0),.clk(gclk));
	jdff dff_A_0PV6cdnB5_0(.dout(w_dff_A_Jlef4EEs7_0),.din(w_dff_A_0PV6cdnB5_0),.clk(gclk));
	jdff dff_A_FOJ7HYgQ0_0(.dout(w_dff_A_0PV6cdnB5_0),.din(w_dff_A_FOJ7HYgQ0_0),.clk(gclk));
	jdff dff_A_8VPOe6SL6_0(.dout(w_dff_A_FOJ7HYgQ0_0),.din(w_dff_A_8VPOe6SL6_0),.clk(gclk));
	jdff dff_A_GtpHoEfs6_0(.dout(w_dff_A_8VPOe6SL6_0),.din(w_dff_A_GtpHoEfs6_0),.clk(gclk));
	jdff dff_A_nIt0Sw2C8_2(.dout(w_G56gat_0[2]),.din(w_dff_A_nIt0Sw2C8_2),.clk(gclk));
	jdff dff_A_oxqdqFdH8_0(.dout(w_n49_0[0]),.din(w_dff_A_oxqdqFdH8_0),.clk(gclk));
	jdff dff_A_A0zQVHCd9_0(.dout(w_dff_A_oxqdqFdH8_0),.din(w_dff_A_A0zQVHCd9_0),.clk(gclk));
	jdff dff_A_HAJ8INlW8_0(.dout(w_dff_A_A0zQVHCd9_0),.din(w_dff_A_HAJ8INlW8_0),.clk(gclk));
	jdff dff_A_AFXSpOTL0_0(.dout(w_dff_A_HAJ8INlW8_0),.din(w_dff_A_AFXSpOTL0_0),.clk(gclk));
	jdff dff_A_gNpeiWC76_0(.dout(w_G50gat_0[0]),.din(w_dff_A_gNpeiWC76_0),.clk(gclk));
	jdff dff_A_X04574qT0_0(.dout(w_dff_A_gNpeiWC76_0),.din(w_dff_A_X04574qT0_0),.clk(gclk));
	jdff dff_A_bCzKI3Ty9_1(.dout(w_G50gat_0[1]),.din(w_dff_A_bCzKI3Ty9_1),.clk(gclk));
	jdff dff_A_iV4VKlYT5_1(.dout(w_G82gat_0[1]),.din(w_dff_A_iV4VKlYT5_1),.clk(gclk));
	jdff dff_A_AQlHL5dX4_1(.dout(w_dff_A_iV4VKlYT5_1),.din(w_dff_A_AQlHL5dX4_1),.clk(gclk));
	jdff dff_A_3MH6jBP51_1(.dout(w_dff_A_AQlHL5dX4_1),.din(w_dff_A_3MH6jBP51_1),.clk(gclk));
	jdff dff_A_gHkb2n0z4_1(.dout(w_dff_A_3MH6jBP51_1),.din(w_dff_A_gHkb2n0z4_1),.clk(gclk));
	jdff dff_A_mbmiBSyX7_1(.dout(w_dff_A_gHkb2n0z4_1),.din(w_dff_A_mbmiBSyX7_1),.clk(gclk));
	jdff dff_A_VzTadzja5_2(.dout(w_G82gat_0[2]),.din(w_dff_A_VzTadzja5_2),.clk(gclk));
	jdff dff_A_rrsSLf0g5_0(.dout(w_n46_0[0]),.din(w_dff_A_rrsSLf0g5_0),.clk(gclk));
	jdff dff_A_lR29XX9a3_0(.dout(w_dff_A_rrsSLf0g5_0),.din(w_dff_A_lR29XX9a3_0),.clk(gclk));
	jdff dff_A_dDBMv6kV5_0(.dout(w_dff_A_lR29XX9a3_0),.din(w_dff_A_dDBMv6kV5_0),.clk(gclk));
	jdff dff_A_YICBIYUR5_0(.dout(w_dff_A_dDBMv6kV5_0),.din(w_dff_A_YICBIYUR5_0),.clk(gclk));
	jdff dff_A_O8hs6JXi2_0(.dout(w_G76gat_0[0]),.din(w_dff_A_O8hs6JXi2_0),.clk(gclk));
	jdff dff_A_A5gMHVGY8_0(.dout(w_dff_A_O8hs6JXi2_0),.din(w_dff_A_A5gMHVGY8_0),.clk(gclk));
	jdff dff_A_ABan4mVc1_1(.dout(w_G17gat_0[1]),.din(w_dff_A_ABan4mVc1_1),.clk(gclk));
	jdff dff_A_6tTDm9QE1_1(.dout(w_dff_A_ABan4mVc1_1),.din(w_dff_A_6tTDm9QE1_1),.clk(gclk));
	jdff dff_A_p4a7zD0u7_1(.dout(w_dff_A_6tTDm9QE1_1),.din(w_dff_A_p4a7zD0u7_1),.clk(gclk));
	jdff dff_A_FiuEEm6L9_1(.dout(w_dff_A_p4a7zD0u7_1),.din(w_dff_A_FiuEEm6L9_1),.clk(gclk));
	jdff dff_A_TrwZZhQ47_1(.dout(w_dff_A_FiuEEm6L9_1),.din(w_dff_A_TrwZZhQ47_1),.clk(gclk));
	jdff dff_A_XnK8trYj6_2(.dout(w_G17gat_0[2]),.din(w_dff_A_XnK8trYj6_2),.clk(gclk));
	jdff dff_A_BdAAYCsi3_0(.dout(w_n44_0[0]),.din(w_dff_A_BdAAYCsi3_0),.clk(gclk));
	jdff dff_A_MWyuzg3i9_0(.dout(w_dff_A_BdAAYCsi3_0),.din(w_dff_A_MWyuzg3i9_0),.clk(gclk));
	jdff dff_A_Bl61cQJR4_0(.dout(w_dff_A_MWyuzg3i9_0),.din(w_dff_A_Bl61cQJR4_0),.clk(gclk));
	jdff dff_A_DNklI1Sz2_0(.dout(w_dff_A_Bl61cQJR4_0),.din(w_dff_A_DNklI1Sz2_0),.clk(gclk));
	jdff dff_A_HIO2QXR52_0(.dout(w_G11gat_0[0]),.din(w_dff_A_HIO2QXR52_0),.clk(gclk));
	jdff dff_A_UEOo2iVB1_0(.dout(w_dff_A_HIO2QXR52_0),.din(w_dff_A_UEOo2iVB1_0),.clk(gclk));
	jdff dff_A_rGuLBSJD8_0(.dout(w_n84_0[0]),.din(w_dff_A_rGuLBSJD8_0),.clk(gclk));
	jdff dff_A_VmNbwtX40_0(.dout(w_dff_A_rGuLBSJD8_0),.din(w_dff_A_VmNbwtX40_0),.clk(gclk));
	jdff dff_A_WSKhU4EA2_0(.dout(w_G30gat_0[0]),.din(w_dff_A_WSKhU4EA2_0),.clk(gclk));
	jdff dff_A_Vr58FxO11_0(.dout(w_dff_A_WSKhU4EA2_0),.din(w_dff_A_Vr58FxO11_0),.clk(gclk));
	jdff dff_A_5uny8MAX6_0(.dout(w_dff_A_Vr58FxO11_0),.din(w_dff_A_5uny8MAX6_0),.clk(gclk));
	jdff dff_A_kXDw8aob9_0(.dout(w_dff_A_5uny8MAX6_0),.din(w_dff_A_kXDw8aob9_0),.clk(gclk));
	jdff dff_A_jouY31xd5_0(.dout(w_dff_A_kXDw8aob9_0),.din(w_dff_A_jouY31xd5_0),.clk(gclk));
	jdff dff_A_l0ipPEzk1_2(.dout(w_G30gat_0[2]),.din(w_dff_A_l0ipPEzk1_2),.clk(gclk));
endmodule

