module rf_c5315(G4115, G4092, G4089, G4087, G3724, G3550, G3548, G3546, G2824, G2358, G1694, G1690, G1689, G562, G552, G545, G534, G468, G435, G4091, G479, G422, G3173, G411, G556, G400, G523, G386, G373, G369, G366, G361, G348, G254, G127, G121, G119, G167, G114, G191, G112, G164, G389, G106, G103, G152, G117, G242, G100, G161, G118, G87, G97, G88, G146, G86, G83, G549, G82, G307, G3717, G46, G245, G358, G265, G11, G27, G123, G54, G116, G374, G43, G26, G31, G1497, G332, G218, G299, G372, G1, G128, G73, G14, G3552, G122, G248, G120, G109, G4, G23, G113, G76, G145, G34, G91, G49, G225, G64, G131, G351, G126, G37, G94, G149, G81, G226, G1691, G61, G80, G79, G280, G20, G67, G308, G503, G241, G70, G130, G200, G559, G132, G135, G188, G206, G209, G335, G136, G137, G141, G140, G197, G490, G155, G185, G158, G315, G170, G129, G17, G173, G176, G179, G182, G273, G293, G194, G210, G457, G53, G233, G234, G251, G289, G257, G514, G264, G288, G2174, G292, G302, G4090, G25, G316, G4088, G272, G323, G24, G203, G40, G324, G52, G331, G446, G281, G217, G338, G115, G341, G658, G807, G843, G685, G679, G654, G651, G648, G645, G742, G727, G869, G712, G854, G782, G826, G882, G818, G702, G813, G699, G696, G824, G670, G792, G762, G752, G693, G661, G1000, G998, G877, G873, G664, G871, G859, G834, G606, G787, G921, G828, G973, G939, G867, G851, G850, G865, G715, G757, G612, G849, G623, G634, G777, G772, G861, G603, G656, G767, G848, G875, G845, G747, G298, G636, G591, G601, G887, G599, G926, G688, G810, G600, G642, G809, G836, G611, G585, G949, G604, G667, G923, G144, G602, G832, G993, G594, G889, G1004, G892, G838, G802, G575, G1002, G978, G797, G593, G704, G717, G820, G737, G639, G732, G847, G673, G863, G707, G830, G632, G690, G598, G610, G682, G676, G588, G621, G615, G629, G626, G722, G815, G618, G822);
    input G4115, G4092, G4089, G4087, G3724, G3550, G3548, G3546, G2824, G2358, G1694, G1690, G1689, G562, G552, G545, G534, G468, G435, G4091, G479, G422, G3173, G411, G556, G400, G523, G386, G373, G369, G366, G361, G348, G254, G127, G121, G119, G167, G114, G191, G112, G164, G389, G106, G103, G152, G117, G242, G100, G161, G118, G87, G97, G88, G146, G86, G83, G549, G82, G307, G3717, G46, G245, G358, G265, G11, G27, G123, G54, G116, G374, G43, G26, G31, G1497, G332, G218, G299, G372, G1, G128, G73, G14, G3552, G122, G248, G120, G109, G4, G23, G113, G76, G145, G34, G91, G49, G225, G64, G131, G351, G126, G37, G94, G149, G81, G226, G1691, G61, G80, G79, G280, G20, G67, G308, G503, G241, G70, G130, G200, G559, G132, G135, G188, G206, G209, G335, G136, G137, G141, G140, G197, G490, G155, G185, G158, G315, G170, G129, G17, G173, G176, G179, G182, G273, G293, G194, G210, G457, G53, G233, G234, G251, G289, G257, G514, G264, G288, G2174, G292, G302, G4090, G25, G316, G4088, G272, G323, G24, G203, G40, G324, G52, G331, G446, G281, G217, G338, G115, G341;
    output G658, G807, G843, G685, G679, G654, G651, G648, G645, G742, G727, G869, G712, G854, G782, G826, G882, G818, G702, G813, G699, G696, G824, G670, G792, G762, G752, G693, G661, G1000, G998, G877, G873, G664, G871, G859, G834, G606, G787, G921, G828, G973, G939, G867, G851, G850, G865, G715, G757, G612, G849, G623, G634, G777, G772, G861, G603, G656, G767, G848, G875, G845, G747, G298, G636, G591, G601, G887, G599, G926, G688, G810, G600, G642, G809, G836, G611, G585, G949, G604, G667, G923, G144, G602, G832, G993, G594, G889, G1004, G892, G838, G802, G575, G1002, G978, G797, G593, G704, G717, G820, G737, G639, G732, G847, G673, G863, G707, G830, G632, G690, G598, G610, G682, G676, G588, G621, G615, G629, G626, G722, G815, G618, G822;
    wire n303;
    wire n306;
    wire n309;
    wire n313;
    wire n316;
    wire n319;
    wire n322;
    wire n326;
    wire n329;
    wire n332;
    wire n335;
    wire n338;
    wire n342;
    wire n345;
    wire n349;
    wire n352;
    wire n356;
    wire n360;
    wire n363;
    wire n366;
    wire n369;
    wire n373;
    wire n377;
    wire n380;
    wire n383;
    wire n386;
    wire n390;
    wire n393;
    wire n397;
    wire n401;
    wire n405;
    wire n408;
    wire n412;
    wire n415;
    wire n419;
    wire n423;
    wire n427;
    wire n430;
    wire n434;
    wire n438;
    wire n442;
    wire n446;
    wire n450;
    wire n454;
    wire n458;
    wire n462;
    wire n466;
    wire n470;
    wire n474;
    wire n478;
    wire n482;
    wire n486;
    wire n490;
    wire n494;
    wire n498;
    wire n502;
    wire n506;
    wire n510;
    wire n514;
    wire n517;
    wire n521;
    wire n524;
    wire n528;
    wire n532;
    wire n536;
    wire n539;
    wire n543;
    wire n546;
    wire n550;
    wire n554;
    wire n558;
    wire n562;
    wire n565;
    wire n569;
    wire n572;
    wire n576;
    wire n580;
    wire n584;
    wire n588;
    wire n592;
    wire n596;
    wire n600;
    wire n604;
    wire n608;
    wire n611;
    wire n614;
    wire n618;
    wire n621;
    wire n624;
    wire n628;
    wire n632;
    wire n636;
    wire n640;
    wire n644;
    wire n648;
    wire n652;
    wire n656;
    wire n659;
    wire n663;
    wire n667;
    wire n671;
    wire n674;
    wire n677;
    wire n681;
    wire n684;
    wire n688;
    wire n692;
    wire n695;
    wire n699;
    wire n702;
    wire n705;
    wire n709;
    wire n713;
    wire n717;
    wire n720;
    wire n723;
    wire n727;
    wire n731;
    wire n735;
    wire n738;
    wire n742;
    wire n746;
    wire n750;
    wire n753;
    wire n757;
    wire n760;
    wire n764;
    wire n768;
    wire n772;
    wire n776;
    wire n780;
    wire n784;
    wire n788;
    wire n792;
    wire n795;
    wire n799;
    wire n802;
    wire n806;
    wire n810;
    wire n814;
    wire n818;
    wire n822;
    wire n826;
    wire n830;
    wire n834;
    wire n838;
    wire n842;
    wire n846;
    wire n849;
    wire n853;
    wire n856;
    wire n860;
    wire n864;
    wire n868;
    wire n872;
    wire n876;
    wire n880;
    wire n884;
    wire n888;
    wire n891;
    wire n895;
    wire n898;
    wire n902;
    wire n906;
    wire n910;
    wire n914;
    wire n918;
    wire n922;
    wire n926;
    wire n930;
    wire n933;
    wire n937;
    wire n940;
    wire n944;
    wire n948;
    wire n952;
    wire n956;
    wire n960;
    wire n964;
    wire n968;
    wire n972;
    wire n976;
    wire n980;
    wire n983;
    wire n987;
    wire n990;
    wire n994;
    wire n998;
    wire n1002;
    wire n1006;
    wire n1010;
    wire n1014;
    wire n1018;
    wire n1022;
    wire n1025;
    wire n1029;
    wire n1032;
    wire n1036;
    wire n1040;
    wire n1044;
    wire n1048;
    wire n1052;
    wire n1056;
    wire n1060;
    wire n1064;
    wire n1068;
    wire n1071;
    wire n1075;
    wire n1078;
    wire n1082;
    wire n1086;
    wire n1090;
    wire n1094;
    wire n1098;
    wire n1102;
    wire n1106;
    wire n1110;
    wire n1113;
    wire n1117;
    wire n1120;
    wire n1124;
    wire n1128;
    wire n1132;
    wire n1136;
    wire n1140;
    wire n1144;
    wire n1148;
    wire n1152;
    wire n1156;
    wire n1159;
    wire n1163;
    wire n1166;
    wire n1170;
    wire n1174;
    wire n1178;
    wire n1182;
    wire n1186;
    wire n1190;
    wire n1194;
    wire n1198;
    wire n1201;
    wire n1205;
    wire n1208;
    wire n1212;
    wire n1216;
    wire n1220;
    wire n1224;
    wire n1228;
    wire n1232;
    wire n1236;
    wire n1240;
    wire n1244;
    wire n1248;
    wire n1252;
    wire n1256;
    wire n1259;
    wire n1263;
    wire n1267;
    wire n1270;
    wire n1274;
    wire n1278;
    wire n1281;
    wire n1284;
    wire n1288;
    wire n1292;
    wire n1296;
    wire n1300;
    wire n1304;
    wire n1308;
    wire n1312;
    wire n1316;
    wire n1319;
    wire n1323;
    wire n1326;
    wire n1330;
    wire n1334;
    wire n1338;
    wire n1342;
    wire n1345;
    wire n1349;
    wire n1353;
    wire n1357;
    wire n1361;
    wire n1365;
    wire n1369;
    wire n1373;
    wire n1376;
    wire n1380;
    wire n1384;
    wire n1388;
    wire n1392;
    wire n1396;
    wire n1400;
    wire n1403;
    wire n1407;
    wire n1411;
    wire n1415;
    wire n1419;
    wire n1423;
    wire n1427;
    wire n1431;
    wire n1435;
    wire n1439;
    wire n1443;
    wire n1447;
    wire n1451;
    wire n1455;
    wire n1459;
    wire n1462;
    wire n1466;
    wire n1470;
    wire n1473;
    wire n1477;
    wire n1481;
    wire n1485;
    wire n1489;
    wire n1493;
    wire n1497;
    wire n1501;
    wire n1505;
    wire n1509;
    wire n1512;
    wire n1516;
    wire n1520;
    wire n1524;
    wire n1528;
    wire n1532;
    wire n1536;
    wire n1540;
    wire n1544;
    wire n1548;
    wire n1551;
    wire n1555;
    wire n1559;
    wire n1563;
    wire n1567;
    wire n1571;
    wire n1575;
    wire n1578;
    wire n1582;
    wire n1585;
    wire n1589;
    wire n1593;
    wire n1597;
    wire n1601;
    wire n1605;
    wire n1609;
    wire n1613;
    wire n1617;
    wire n1621;
    wire n1625;
    wire n1629;
    wire n1633;
    wire n1637;
    wire n1641;
    wire n1645;
    wire n1649;
    wire n1653;
    wire n1657;
    wire n1661;
    wire n1665;
    wire n1668;
    wire n1672;
    wire n1676;
    wire n1680;
    wire n1684;
    wire n1688;
    wire n1692;
    wire n1696;
    wire n1700;
    wire n1704;
    wire n1707;
    wire n1710;
    wire n1714;
    wire n1717;
    wire n1721;
    wire n1724;
    wire n1728;
    wire n1732;
    wire n1736;
    wire n1740;
    wire n1744;
    wire n1747;
    wire n1751;
    wire n1754;
    wire n1758;
    wire n1762;
    wire n1766;
    wire n1770;
    wire n1774;
    wire n1778;
    wire n1782;
    wire n1786;
    wire n1789;
    wire n1793;
    wire n1797;
    wire n1801;
    wire n1805;
    wire n1809;
    wire n1813;
    wire n1817;
    wire n1821;
    wire n1825;
    wire n1829;
    wire n1833;
    wire n1837;
    wire n1841;
    wire n1845;
    wire n1849;
    wire n1853;
    wire n1857;
    wire n1861;
    wire n1865;
    wire n1869;
    wire n1873;
    wire n1877;
    wire n1881;
    wire n1885;
    wire n1889;
    wire n1893;
    wire n1897;
    wire n1901;
    wire n1905;
    wire n1909;
    wire n1913;
    wire n1917;
    wire n1921;
    wire n1925;
    wire n1929;
    wire n1932;
    wire n1936;
    wire n1940;
    wire n1944;
    wire n1947;
    wire n1950;
    wire n1954;
    wire n1957;
    wire n1961;
    wire n1965;
    wire n1969;
    wire n1973;
    wire n1977;
    wire n1981;
    wire n1984;
    wire n1988;
    wire n1991;
    wire n1995;
    wire n1998;
    wire n2002;
    wire n2005;
    wire n2009;
    wire n2013;
    wire n2017;
    wire n2021;
    wire n2025;
    wire n2028;
    wire n2032;
    wire n2035;
    wire n2039;
    wire n2042;
    wire n2046;
    wire n2050;
    wire n2054;
    wire n2058;
    wire n2061;
    wire n2065;
    wire n2069;
    wire n2072;
    wire n2076;
    wire n2080;
    wire n2084;
    wire n2088;
    wire n2091;
    wire n2095;
    wire n2099;
    wire n2102;
    wire n2106;
    wire n2110;
    wire n2113;
    wire n2117;
    wire n2121;
    wire n2125;
    wire n2129;
    wire n2132;
    wire n2136;
    wire n2140;
    wire n2143;
    wire n2147;
    wire n2151;
    wire n2154;
    wire n2157;
    wire n2160;
    wire n2164;
    wire n2168;
    wire n2171;
    wire n2174;
    wire n2178;
    wire n2182;
    wire n2186;
    wire n2190;
    wire n2194;
    wire n2198;
    wire n2202;
    wire n2206;
    wire n2210;
    wire n2214;
    wire n2218;
    wire n2222;
    wire n2226;
    wire n2230;
    wire n2234;
    wire n2238;
    wire n2241;
    wire n2245;
    wire n2249;
    wire n2252;
    wire n2256;
    wire n2260;
    wire n2264;
    wire n2268;
    wire n2272;
    wire n2276;
    wire n2280;
    wire n2284;
    wire n2288;
    wire n2291;
    wire n2295;
    wire n2299;
    wire n2303;
    wire n2307;
    wire n2311;
    wire n2315;
    wire n2319;
    wire n2323;
    wire n2327;
    wire n2330;
    wire n2334;
    wire n2338;
    wire n2341;
    wire n2345;
    wire n2349;
    wire n2352;
    wire n2356;
    wire n2360;
    wire n2364;
    wire n2368;
    wire n2372;
    wire n2376;
    wire n2380;
    wire n2384;
    wire n2388;
    wire n2391;
    wire n2394;
    wire n2398;
    wire n2402;
    wire n2405;
    wire n2408;
    wire n2412;
    wire n2416;
    wire n2420;
    wire n2424;
    wire n2428;
    wire n2432;
    wire n2436;
    wire n2440;
    wire n2443;
    wire n2447;
    wire n2451;
    wire n2455;
    wire n2459;
    wire n2463;
    wire n2467;
    wire n2470;
    wire n2474;
    wire n2478;
    wire n2482;
    wire n2485;
    wire n2489;
    wire n2493;
    wire n2497;
    wire n2501;
    wire n2505;
    wire n2508;
    wire n2512;
    wire n2516;
    wire n2519;
    wire n2523;
    wire n2527;
    wire n2531;
    wire n2535;
    wire n2538;
    wire n2542;
    wire n2546;
    wire n2549;
    wire n2553;
    wire n2557;
    wire n2560;
    wire n2564;
    wire n2568;
    wire n2572;
    wire n2576;
    wire n2580;
    wire n2584;
    wire n2588;
    wire n2592;
    wire n2596;
    wire n2600;
    wire n2603;
    wire n2607;
    wire n2610;
    wire n2614;
    wire n2618;
    wire n2622;
    wire n2626;
    wire n2629;
    wire n2633;
    wire n2637;
    wire n2641;
    wire n2645;
    wire n2649;
    wire n2653;
    wire n2657;
    wire n2661;
    wire n2665;
    wire n2669;
    wire n2673;
    wire n2677;
    wire n2680;
    wire n2683;
    wire n2686;
    wire n2689;
    wire n2692;
    wire n2695;
    wire n2699;
    wire n2702;
    wire n2706;
    wire n2710;
    wire n2714;
    wire n2718;
    wire n2722;
    wire n2726;
    wire n2729;
    wire n2732;
    wire n2735;
    wire n2739;
    wire n2743;
    wire n2746;
    wire n2750;
    wire n2753;
    wire n2756;
    wire n2760;
    wire n2764;
    wire n2768;
    wire n2772;
    wire n2775;
    wire n2778;
    wire n2781;
    wire n2784;
    wire n2788;
    wire n2792;
    wire n2796;
    wire n2800;
    wire n2804;
    wire n2808;
    wire n2812;
    wire n2816;
    wire n2819;
    wire n2823;
    wire n2827;
    wire n2831;
    wire n2835;
    wire n2839;
    wire n2843;
    wire n2846;
    wire n2850;
    wire n2854;
    wire n2858;
    wire n2862;
    wire n2866;
    wire n2870;
    wire n2874;
    wire n2878;
    wire n2882;
    wire n2885;
    wire n2889;
    wire n2893;
    wire n2896;
    wire n2900;
    wire n2904;
    wire n2908;
    wire n2912;
    wire n2916;
    wire n2920;
    wire n2924;
    wire n2928;
    wire n2932;
    wire n2936;
    wire n2939;
    wire n2943;
    wire n2947;
    wire n2950;
    wire n2954;
    wire n2958;
    wire n2962;
    wire n2966;
    wire n2970;
    wire n2974;
    wire n2978;
    wire n2982;
    wire n2986;
    wire n2990;
    wire n2993;
    wire n2997;
    wire n3000;
    wire n3004;
    wire n3008;
    wire n3012;
    wire n3016;
    wire n3020;
    wire n3024;
    wire n3027;
    wire n3031;
    wire n3034;
    wire n3038;
    wire n3042;
    wire n3046;
    wire n3050;
    wire n3054;
    wire n3058;
    wire n3061;
    wire n3065;
    wire n3068;
    wire n3072;
    wire n3076;
    wire n3080;
    wire n3084;
    wire n3088;
    wire n3092;
    wire n3095;
    wire n3099;
    wire n3102;
    wire n3106;
    wire n3110;
    wire n3114;
    wire n3118;
    wire n3122;
    wire n3126;
    wire n3130;
    wire n3134;
    wire n3138;
    wire n3142;
    wire n3146;
    wire n3150;
    wire n3154;
    wire n3158;
    wire n3162;
    wire n3166;
    wire n3170;
    wire n3174;
    wire n3178;
    wire n3182;
    wire n3186;
    wire n3190;
    wire n3194;
    wire n3198;
    wire n3202;
    wire n3206;
    wire n3210;
    wire n3214;
    wire n3218;
    wire n3222;
    wire n3226;
    wire n3230;
    wire n3234;
    wire n3238;
    wire n3242;
    wire n3246;
    wire n3250;
    wire n3254;
    wire n3258;
    wire n3262;
    wire n3266;
    wire n3270;
    wire n3274;
    wire n3278;
    wire n3282;
    wire n3286;
    wire n3290;
    wire n3294;
    wire n3298;
    wire n3302;
    wire n3306;
    wire n3310;
    wire n3314;
    wire n3318;
    wire n3322;
    wire n3326;
    wire n3330;
    wire n3334;
    wire n3338;
    wire n3342;
    wire n3346;
    wire n3350;
    wire n3354;
    wire n3358;
    wire n3362;
    wire n3366;
    wire n3370;
    wire n3374;
    wire n3378;
    wire n3382;
    wire n3386;
    wire n3390;
    wire n3394;
    wire n3398;
    wire n3402;
    wire n3406;
    wire n3410;
    wire n3414;
    wire n3418;
    wire n3422;
    wire n3426;
    wire n3430;
    wire n3434;
    wire n3438;
    wire n3442;
    wire n3446;
    wire n3450;
    wire n3454;
    wire n3458;
    wire n3462;
    wire n3466;
    wire n3470;
    wire n3474;
    wire n3478;
    wire n3482;
    wire n3486;
    wire n3490;
    wire n3494;
    wire n3498;
    wire n3501;
    wire n3504;
    wire n3508;
    wire n3512;
    wire n3516;
    wire n3519;
    wire n3522;
    wire n3526;
    wire n3530;
    wire n3534;
    wire n3537;
    wire n3541;
    wire n3545;
    wire n3549;
    wire n3553;
    wire n3557;
    wire n3561;
    wire n3565;
    wire n3569;
    wire n3573;
    wire n3577;
    wire n3581;
    wire n3585;
    wire n3588;
    wire n3592;
    wire n3596;
    wire n3600;
    wire n3604;
    wire n3607;
    wire n3611;
    wire n3615;
    wire n3619;
    wire n3623;
    wire n3626;
    wire n3630;
    wire n3634;
    wire n3638;
    wire n3641;
    wire n3645;
    wire n3649;
    wire n3652;
    wire n3656;
    wire n3660;
    wire n3663;
    wire n3667;
    wire n3671;
    wire n3675;
    wire n3679;
    wire n3683;
    wire n3687;
    wire n3691;
    wire n3695;
    wire n3698;
    wire n3702;
    wire n3706;
    wire n3710;
    wire n3714;
    wire n3717;
    wire n3721;
    wire n3725;
    wire n3729;
    wire n3732;
    wire n3736;
    wire n3739;
    wire n3743;
    wire n3746;
    wire n3750;
    wire n3754;
    wire n3758;
    wire n3761;
    wire n3765;
    wire n3769;
    wire n3773;
    wire n3776;
    wire n3780;
    wire n3784;
    wire n3787;
    wire n3791;
    wire n3795;
    wire n3799;
    wire n3803;
    wire n3807;
    wire n3811;
    wire n3815;
    wire n3819;
    wire n3823;
    wire n3827;
    wire n3831;
    wire n3835;
    wire n3839;
    wire n3843;
    wire n3847;
    wire n3851;
    wire n3855;
    wire n3858;
    wire n3862;
    wire n3866;
    wire n3870;
    wire n3874;
    wire n3878;
    wire n3882;
    wire n3885;
    wire n3889;
    wire n3892;
    wire n3896;
    wire n3900;
    wire n3904;
    wire n3908;
    wire n3912;
    wire n3916;
    wire n3919;
    wire n3923;
    wire n3926;
    wire n3930;
    wire n3934;
    wire n3938;
    wire n3942;
    wire n3946;
    wire n3950;
    wire n3954;
    wire n3958;
    wire n3962;
    wire n3966;
    wire n3970;
    wire n3974;
    wire n3978;
    wire n3982;
    wire n3986;
    wire n3990;
    wire n3994;
    wire n3998;
    wire n4002;
    wire n4006;
    wire n4010;
    wire n4014;
    wire n4018;
    wire n4022;
    wire n4026;
    wire n4030;
    wire n4034;
    wire n4038;
    wire n4042;
    wire n4046;
    wire n4050;
    wire n4054;
    wire n4058;
    wire n4062;
    wire n4066;
    wire n4070;
    wire n4074;
    wire n4078;
    wire n4082;
    wire n4086;
    wire n4090;
    wire n4094;
    wire n4098;
    wire n4102;
    wire n4106;
    wire n4110;
    wire n4114;
    wire n4118;
    wire n4122;
    wire n4126;
    wire n4130;
    wire n4134;
    wire n4138;
    wire n4142;
    wire n4146;
    wire n4150;
    wire n4154;
    wire n4158;
    wire n4162;
    wire n4166;
    wire n4170;
    wire n4174;
    wire n4178;
    wire n4182;
    wire n4186;
    wire n4190;
    wire n4194;
    wire n4198;
    wire n4202;
    wire n4206;
    wire n4210;
    wire n4214;
    wire n4218;
    wire n4222;
    wire n4226;
    wire n4230;
    wire n4234;
    wire n4238;
    wire n4242;
    wire n4246;
    wire n4250;
    wire n4254;
    wire n4258;
    wire n4262;
    wire n4266;
    wire n4270;
    wire n4274;
    wire n4278;
    wire n4282;
    wire n4286;
    wire n4290;
    wire n4294;
    wire n4298;
    wire n4302;
    wire n4306;
    wire n4310;
    wire n4314;
    wire n4318;
    wire n4322;
    wire n4326;
    wire n4330;
    wire n4334;
    wire n4338;
    wire n4342;
    wire n4346;
    wire n4349;
    wire n4353;
    wire n4357;
    wire n4361;
    wire n4365;
    wire n4369;
    wire n4373;
    wire n4377;
    wire n4381;
    wire n4385;
    wire n4389;
    wire n4393;
    wire n4397;
    wire n4401;
    wire n4405;
    wire n4409;
    wire n4413;
    wire n4417;
    wire n4421;
    wire n4425;
    wire n4429;
    wire n4433;
    wire n4437;
    wire n4441;
    wire n4445;
    wire n4448;
    wire n4452;
    wire n4456;
    wire n4460;
    wire n4464;
    wire n4468;
    wire n4472;
    wire n4475;
    wire n4479;
    wire n4483;
    wire n4487;
    wire n4491;
    wire n4495;
    wire n4499;
    wire n4502;
    wire n4506;
    wire n4509;
    wire n4513;
    wire n4517;
    wire n4521;
    wire n4525;
    wire n4528;
    wire n4532;
    wire n4536;
    wire n4540;
    wire n4543;
    wire n4547;
    wire n4550;
    wire n4554;
    wire n4557;
    wire n4560;
    wire n4564;
    wire n4568;
    wire n4572;
    wire n4576;
    wire n4580;
    wire n4584;
    wire n4587;
    wire n4591;
    wire n4595;
    wire n4599;
    wire n4603;
    wire n4607;
    wire n4610;
    wire n4614;
    wire n4618;
    wire n4622;
    wire n4626;
    wire n4630;
    wire n4634;
    wire n4637;
    wire n4641;
    wire n4645;
    wire n4649;
    wire n4653;
    wire n4656;
    wire n4660;
    wire n4664;
    wire n4668;
    wire n4672;
    wire n4676;
    wire n4680;
    wire n4684;
    wire n4688;
    wire n4692;
    wire n4696;
    wire n4700;
    wire n4704;
    wire n4708;
    wire n4712;
    wire n4716;
    wire n4720;
    wire n4724;
    wire n4728;
    wire n4732;
    wire n4736;
    wire n4740;
    wire n4744;
    wire n4748;
    wire n4752;
    wire n4756;
    wire n4760;
    wire n4764;
    wire n4768;
    wire n4772;
    wire n4776;
    wire n4780;
    wire n4784;
    wire n4788;
    wire n4792;
    wire n4796;
    wire n4800;
    wire n4804;
    wire n4808;
    wire n4812;
    wire n4816;
    wire n4820;
    wire n4824;
    wire n4828;
    wire n4832;
    wire n4836;
    wire n4840;
    wire n4844;
    wire n4848;
    wire n4852;
    wire n4856;
    wire n4860;
    wire n4864;
    wire n4868;
    wire n4872;
    wire n4876;
    wire n4880;
    wire n4884;
    wire n4888;
    wire n4892;
    wire n4896;
    wire n4900;
    wire n4904;
    wire n4908;
    wire n4912;
    wire n4916;
    wire n4920;
    wire n4924;
    wire n4928;
    wire n4932;
    wire n4936;
    wire n4940;
    wire n4944;
    wire n4948;
    wire n4952;
    wire n4956;
    wire n4960;
    wire n4964;
    wire n4968;
    wire n4972;
    wire n4976;
    wire n4980;
    wire n4984;
    wire n4988;
    wire n4992;
    wire n4996;
    wire n5000;
    wire n5004;
    wire n5008;
    wire n5012;
    wire n5016;
    wire n5020;
    wire n5024;
    wire n5028;
    wire n5032;
    wire n5035;
    wire n5039;
    wire n5043;
    wire n5047;
    wire n5051;
    wire n5055;
    wire n5059;
    wire n5063;
    wire n5066;
    wire n5070;
    wire n5074;
    wire n5077;
    wire n5081;
    wire n5085;
    wire n5089;
    wire n5093;
    wire n5097;
    wire n5101;
    wire n5105;
    wire n5109;
    wire n5113;
    wire n5116;
    wire n5120;
    wire n5124;
    wire n5128;
    wire n5132;
    wire n5136;
    wire n5139;
    wire n5143;
    wire n5147;
    wire n5151;
    wire n5155;
    wire n5158;
    wire n5162;
    wire n5166;
    wire n5170;
    wire n5174;
    wire n5178;
    wire n5182;
    wire n5186;
    wire n5190;
    wire n5194;
    wire n5198;
    wire n5202;
    wire n5206;
    wire n5210;
    wire n5213;
    wire n5217;
    wire n5221;
    wire n5225;
    wire n5229;
    wire n5233;
    wire n5237;
    wire n5241;
    wire n5245;
    wire n5249;
    wire n5253;
    wire n5257;
    wire n5260;
    wire n5264;
    wire n5268;
    wire n5272;
    wire n5276;
    wire n5280;
    wire n5284;
    wire n5287;
    wire n5291;
    wire n5294;
    wire n5298;
    wire n5301;
    wire n5305;
    wire n5309;
    wire n5313;
    wire n5317;
    wire n5321;
    wire n5325;
    wire n5329;
    wire n5333;
    wire n5337;
    wire n5341;
    wire n5345;
    wire n5349;
    wire n5353;
    wire n5357;
    wire n5361;
    wire n5365;
    wire n5369;
    wire n5373;
    wire n5377;
    wire n5380;
    wire n5383;
    wire n5387;
    wire n5390;
    wire n5393;
    wire n5397;
    wire n5401;
    wire n5404;
    wire n5407;
    wire n5411;
    wire n5414;
    wire n5417;
    wire n5421;
    wire n5425;
    wire n5429;
    wire n5433;
    wire n5440;
    wire n5444;
    wire n5447;
    wire n5451;
    wire n5454;
    wire n5458;
    wire n5461;
    wire n5465;
    wire n5469;
    wire n5473;
    wire n5477;
    wire n5484;
    wire n5487;
    wire n5490;
    wire n5493;
    wire n5496;
    wire n5499;
    wire n5502;
    wire n5505;
    wire n5508;
    wire n5511;
    wire n5514;
    wire n5517;
    wire n5520;
    wire n5523;
    wire n5526;
    wire n5529;
    wire n5533;
    wire n5537;
    wire n5541;
    wire n5545;
    wire n5549;
    wire n8016;
    wire n8019;
    wire n8022;
    wire n8025;
    wire n8028;
    wire n8031;
    wire n8034;
    wire n8037;
    wire n8040;
    wire n8043;
    wire n8046;
    wire n8049;
    wire n8051;
    wire n8054;
    wire n8057;
    wire n8060;
    wire n8063;
    wire n8066;
    wire n8069;
    wire n8072;
    wire n8076;
    wire n8079;
    wire n8082;
    wire n8085;
    wire n8088;
    wire n8091;
    wire n8093;
    wire n8096;
    wire n8099;
    wire n8102;
    wire n8105;
    wire n8108;
    wire n8111;
    wire n8114;
    wire n8117;
    wire n8120;
    wire n8124;
    wire n8127;
    wire n8130;
    wire n8133;
    wire n8136;
    wire n8139;
    wire n8142;
    wire n8145;
    wire n8148;
    wire n8151;
    wire n8154;
    wire n8157;
    wire n8160;
    wire n8163;
    wire n8166;
    wire n8169;
    wire n8171;
    wire n8174;
    wire n8178;
    wire n8181;
    wire n8184;
    wire n8187;
    wire n8190;
    wire n8193;
    wire n8196;
    wire n8199;
    wire n8202;
    wire n8204;
    wire n8207;
    wire n8210;
    wire n8213;
    wire n8216;
    wire n8219;
    wire n8223;
    wire n8226;
    wire n8229;
    wire n8232;
    wire n8235;
    wire n8238;
    wire n8241;
    wire n8244;
    wire n8247;
    wire n8250;
    wire n8253;
    wire n8256;
    wire n8259;
    wire n8262;
    wire n8265;
    wire n8268;
    wire n8271;
    wire n8274;
    wire n8277;
    wire n8280;
    wire n8283;
    wire n8286;
    wire n8289;
    wire n8292;
    wire n8295;
    wire n8298;
    wire n8301;
    wire n8304;
    wire n8307;
    wire n8310;
    wire n8313;
    wire n8316;
    wire n8319;
    wire n8322;
    wire n8325;
    wire n8328;
    wire n8331;
    wire n8334;
    wire n8337;
    wire n8340;
    wire n8343;
    wire n8346;
    wire n8349;
    wire n8352;
    wire n8355;
    wire n8358;
    wire n8361;
    wire n8364;
    wire n8367;
    wire n8370;
    wire n8373;
    wire n8376;
    wire n8379;
    wire n8382;
    wire n8385;
    wire n8388;
    wire n8391;
    wire n8394;
    wire n8397;
    wire n8400;
    wire n8403;
    wire n8406;
    wire n8409;
    wire n8412;
    wire n8415;
    wire n8418;
    wire n8421;
    wire n8423;
    wire n8426;
    wire n8429;
    wire n8432;
    wire n8435;
    wire n8438;
    wire n8441;
    wire n8444;
    wire n8447;
    wire n8450;
    wire n8453;
    wire n8456;
    wire n8459;
    wire n8462;
    wire n8465;
    wire n8469;
    wire n8472;
    wire n8475;
    wire n8478;
    wire n8481;
    wire n8484;
    wire n8487;
    wire n8490;
    wire n8493;
    wire n8496;
    wire n8499;
    wire n8502;
    wire n8505;
    wire n8508;
    wire n8511;
    wire n8514;
    wire n8517;
    wire n8520;
    wire n8523;
    wire n8526;
    wire n8529;
    wire n8532;
    wire n8535;
    wire n8538;
    wire n8541;
    wire n8544;
    wire n8547;
    wire n8550;
    wire n8553;
    wire n8556;
    wire n8559;
    wire n8562;
    wire n8565;
    wire n8567;
    wire n8570;
    wire n8573;
    wire n8576;
    wire n8579;
    wire n8582;
    wire n8585;
    wire n8588;
    wire n8591;
    wire n8595;
    wire n8598;
    wire n8601;
    wire n8604;
    wire n8607;
    wire n8610;
    wire n8613;
    wire n8616;
    wire n8619;
    wire n8622;
    wire n8625;
    wire n8628;
    wire n8631;
    wire n8634;
    wire n8637;
    wire n8640;
    wire n8643;
    wire n8645;
    wire n8648;
    wire n8651;
    wire n8654;
    wire n8657;
    wire n8660;
    wire n8663;
    wire n8666;
    wire n8669;
    wire n8672;
    wire n8675;
    wire n8678;
    wire n8681;
    wire n8684;
    wire n8687;
    wire n8691;
    wire n8694;
    wire n8697;
    wire n8700;
    wire n8703;
    wire n8706;
    wire n8709;
    wire n8712;
    wire n8715;
    wire n8718;
    wire n8721;
    wire n8724;
    wire n8727;
    wire n8730;
    wire n8733;
    wire n8736;
    wire n8739;
    wire n8742;
    wire n8745;
    wire n8748;
    wire n8751;
    wire n8754;
    wire n8757;
    wire n8760;
    wire n8763;
    wire n8766;
    wire n8769;
    wire n8772;
    wire n8775;
    wire n8778;
    wire n8781;
    wire n8784;
    wire n8787;
    wire n8790;
    wire n8793;
    wire n8796;
    wire n8799;
    wire n8802;
    wire n8805;
    wire n8808;
    wire n8811;
    wire n8814;
    wire n8816;
    wire n8819;
    wire n8822;
    wire n8825;
    wire n8828;
    wire n8831;
    wire n8834;
    wire n8837;
    wire n8840;
    wire n8844;
    wire n8847;
    wire n8850;
    wire n8853;
    wire n8856;
    wire n8859;
    wire n8862;
    wire n8865;
    wire n8868;
    wire n8871;
    wire n8874;
    wire n8877;
    wire n8880;
    wire n8883;
    wire n8885;
    wire n8888;
    wire n8891;
    wire n8894;
    wire n8897;
    wire n8900;
    wire n8903;
    wire n8906;
    wire n8909;
    wire n8912;
    wire n8915;
    wire n8918;
    wire n8921;
    wire n8924;
    wire n8927;
    wire n8931;
    wire n8934;
    wire n8937;
    wire n8940;
    wire n8943;
    wire n8946;
    wire n8949;
    wire n8952;
    wire n8955;
    wire n8958;
    wire n8961;
    wire n8964;
    wire n8967;
    wire n8970;
    wire n8973;
    wire n8976;
    wire n8979;
    wire n8982;
    wire n8985;
    wire n8988;
    wire n8991;
    wire n8993;
    wire n8996;
    wire n8999;
    wire n9002;
    wire n9005;
    wire n9009;
    wire n9012;
    wire n9015;
    wire n9018;
    wire n9021;
    wire n9024;
    wire n9027;
    wire n9030;
    wire n9033;
    wire n9036;
    wire n9039;
    wire n9042;
    wire n9044;
    wire n9047;
    wire n9050;
    wire n9053;
    wire n9056;
    wire n9059;
    wire n9062;
    wire n9065;
    wire n9068;
    wire n9072;
    wire n9075;
    wire n9078;
    wire n9081;
    wire n9084;
    wire n9087;
    wire n9090;
    wire n9093;
    wire n9096;
    wire n9099;
    wire n9102;
    wire n9105;
    wire n9108;
    wire n9111;
    wire n9114;
    wire n9117;
    wire n9120;
    wire n9122;
    wire n9125;
    wire n9128;
    wire n9131;
    wire n9134;
    wire n9137;
    wire n9140;
    wire n9144;
    wire n9147;
    wire n9150;
    wire n9153;
    wire n9156;
    wire n9159;
    wire n9162;
    wire n9165;
    wire n9168;
    wire n9171;
    wire n9174;
    wire n9177;
    wire n9179;
    wire n9182;
    wire n9185;
    wire n9188;
    wire n9191;
    wire n9194;
    wire n9197;
    wire n9200;
    wire n9204;
    wire n9207;
    wire n9210;
    wire n9213;
    wire n9216;
    wire n9219;
    wire n9222;
    wire n9225;
    wire n9228;
    wire n9231;
    wire n9234;
    wire n9237;
    wire n9240;
    wire n9243;
    wire n9246;
    wire n9249;
    wire n9252;
    wire n9255;
    wire n9258;
    wire n9261;
    wire n9264;
    wire n9267;
    wire n9270;
    wire n9273;
    wire n9276;
    wire n9279;
    wire n9282;
    wire n9285;
    wire n9288;
    wire n9291;
    wire n9294;
    wire n9297;
    wire n9300;
    wire n9303;
    wire n9306;
    wire n9309;
    wire n9312;
    wire n9314;
    wire n9318;
    wire n9321;
    wire n9323;
    wire n9327;
    wire n9330;
    wire n9333;
    wire n9336;
    wire n9339;
    wire n9342;
    wire n9345;
    wire n9348;
    wire n9351;
    wire n9354;
    wire n9357;
    wire n9359;
    wire n9362;
    wire n9365;
    wire n9368;
    wire n9371;
    wire n9374;
    wire n9377;
    wire n9380;
    wire n9383;
    wire n9386;
    wire n9389;
    wire n9392;
    wire n9395;
    wire n9398;
    wire n9402;
    wire n9405;
    wire n9408;
    wire n9411;
    wire n9414;
    wire n9417;
    wire n9420;
    wire n9423;
    wire n9426;
    wire n9429;
    wire n9432;
    wire n9435;
    wire n9438;
    wire n9441;
    wire n9444;
    wire n9447;
    wire n9450;
    wire n9453;
    wire n9456;
    wire n9459;
    wire n9462;
    wire n9465;
    wire n9467;
    wire n9470;
    wire n9473;
    wire n9476;
    wire n9479;
    wire n9482;
    wire n9486;
    wire n9489;
    wire n9492;
    wire n9495;
    wire n9498;
    wire n9501;
    wire n9504;
    wire n9507;
    wire n9510;
    wire n9512;
    wire n9516;
    wire n9519;
    wire n9522;
    wire n9525;
    wire n9528;
    wire n9531;
    wire n9534;
    wire n9537;
    wire n9540;
    wire n9543;
    wire n9546;
    wire n9549;
    wire n9552;
    wire n9555;
    wire n9558;
    wire n9561;
    wire n9564;
    wire n9566;
    wire n9569;
    wire n9572;
    wire n9575;
    wire n9578;
    wire n9581;
    wire n9585;
    wire n9588;
    wire n9591;
    wire n9594;
    wire n9597;
    wire n9600;
    wire n9603;
    wire n9606;
    wire n9609;
    wire n9612;
    wire n9615;
    wire n9618;
    wire n9621;
    wire n9624;
    wire n9626;
    wire n9629;
    wire n9632;
    wire n9635;
    wire n9639;
    wire n9642;
    wire n9644;
    wire n9647;
    wire n9650;
    wire n9653;
    wire n9656;
    wire n9659;
    wire n9662;
    wire n9665;
    wire n9668;
    wire n9672;
    wire n9675;
    wire n9678;
    wire n9681;
    wire n9684;
    wire n9687;
    wire n9690;
    wire n9693;
    wire n9696;
    wire n9699;
    wire n9702;
    wire n9705;
    wire n9708;
    wire n9710;
    wire n9713;
    wire n9716;
    wire n9719;
    wire n9723;
    wire n9726;
    wire n9729;
    wire n9732;
    wire n9735;
    wire n9738;
    wire n9741;
    wire n9744;
    wire n9747;
    wire n9750;
    wire n9753;
    wire n9756;
    wire n9759;
    wire n9762;
    wire n9765;
    wire n9768;
    wire n9771;
    wire n9774;
    wire n9777;
    wire n9780;
    wire n9783;
    wire n9786;
    wire n9789;
    wire n9792;
    wire n9795;
    wire n9798;
    wire n9801;
    wire n9804;
    wire n9807;
    wire n9810;
    wire n9813;
    wire n9816;
    wire n9819;
    wire n9822;
    wire n9825;
    wire n9827;
    wire n9830;
    wire n9833;
    wire n9836;
    wire n9839;
    wire n9842;
    wire n9845;
    wire n9848;
    wire n9851;
    wire n9854;
    wire n9857;
    wire n9860;
    wire n9863;
    wire n9866;
    wire n9869;
    wire n9872;
    wire n9875;
    wire n9878;
    wire n9881;
    wire n9884;
    wire n9887;
    wire n9890;
    wire n9893;
    wire n9896;
    wire n9899;
    wire n9902;
    wire n9905;
    wire n9908;
    wire n9911;
    wire n9914;
    wire n9917;
    wire n9920;
    wire n9923;
    wire n9926;
    wire n9929;
    wire n9932;
    wire n9935;
    wire n9938;
    wire n9941;
    wire n9944;
    wire n9947;
    wire n9950;
    wire n9953;
    wire n9957;
    wire n9960;
    wire n9963;
    wire n9966;
    wire n9969;
    wire n9972;
    wire n9975;
    wire n9977;
    wire n9981;
    wire n9983;
    wire n9987;
    wire n9990;
    wire n9993;
    wire n9996;
    wire n9999;
    wire n10002;
    wire n10005;
    wire n10007;
    wire n10010;
    wire n10013;
    wire n10016;
    wire n10020;
    wire n10022;
    wire n10026;
    wire n10029;
    wire n10032;
    wire n10035;
    wire n10038;
    wire n10041;
    wire n10044;
    wire n10047;
    wire n10050;
    wire n10053;
    wire n10056;
    wire n10059;
    wire n10062;
    wire n10065;
    wire n10068;
    wire n10071;
    wire n10074;
    wire n10077;
    wire n10080;
    wire n10083;
    wire n10086;
    wire n10089;
    wire n10092;
    wire n10095;
    wire n10098;
    wire n10101;
    wire n10104;
    wire n10107;
    wire n10110;
    wire n10113;
    wire n10116;
    wire n10119;
    wire n10122;
    wire n10125;
    wire n10128;
    wire n10131;
    wire n10134;
    wire n10137;
    wire n10140;
    wire n10143;
    wire n10146;
    wire n10149;
    wire n10152;
    wire n10155;
    wire n10158;
    wire n10161;
    wire n10164;
    wire n10167;
    wire n10170;
    wire n10173;
    wire n10176;
    wire n10179;
    wire n10182;
    wire n10185;
    wire n10188;
    wire n10191;
    wire n10194;
    wire n10197;
    wire n10200;
    wire n10203;
    wire n10206;
    wire n10209;
    wire n10212;
    wire n10215;
    wire n10218;
    wire n10221;
    wire n10224;
    wire n10227;
    wire n10230;
    wire n10233;
    wire n10236;
    wire n10239;
    wire n10242;
    wire n10244;
    wire n10247;
    wire n10251;
    wire n10254;
    wire n10257;
    wire n10260;
    wire n10263;
    wire n10266;
    wire n10269;
    wire n10272;
    wire n10275;
    wire n10278;
    wire n10281;
    wire n10284;
    wire n10287;
    wire n10290;
    wire n10293;
    wire n10296;
    wire n10299;
    wire n10302;
    wire n10305;
    wire n10308;
    wire n10311;
    wire n10314;
    wire n10317;
    wire n10320;
    wire n10323;
    wire n10326;
    wire n10329;
    wire n10332;
    wire n10335;
    wire n10338;
    wire n10341;
    wire n10344;
    wire n10347;
    wire n10350;
    wire n10353;
    wire n10356;
    wire n10359;
    wire n10362;
    wire n10365;
    wire n10368;
    wire n10371;
    wire n10374;
    wire n10377;
    wire n10380;
    wire n10383;
    wire n10386;
    wire n10389;
    wire n10392;
    wire n10395;
    wire n10398;
    wire n10401;
    wire n10404;
    wire n10407;
    wire n10410;
    wire n10413;
    wire n10416;
    wire n10418;
    wire n10421;
    wire n10425;
    wire n10428;
    wire n10431;
    wire n10434;
    wire n10437;
    wire n10440;
    wire n10443;
    wire n10446;
    wire n10449;
    wire n10452;
    wire n10455;
    wire n10458;
    wire n10461;
    wire n10464;
    wire n10467;
    wire n10470;
    wire n10473;
    wire n10476;
    wire n10479;
    wire n10482;
    wire n10485;
    wire n10488;
    wire n10491;
    wire n10494;
    wire n10497;
    wire n10500;
    wire n10503;
    wire n10506;
    wire n10509;
    wire n10512;
    wire n10515;
    wire n10518;
    wire n10521;
    wire n10524;
    wire n10527;
    wire n10529;
    wire n10532;
    wire n10535;
    wire n10538;
    wire n10541;
    wire n10544;
    wire n10548;
    wire n10551;
    wire n10554;
    wire n10557;
    wire n10560;
    wire n10563;
    wire n10566;
    wire n10569;
    wire n10572;
    wire n10575;
    wire n10578;
    wire n10581;
    wire n10584;
    wire n10587;
    wire n10590;
    wire n10593;
    wire n10596;
    wire n10599;
    wire n10602;
    wire n10605;
    wire n10608;
    wire n10611;
    wire n10614;
    wire n10617;
    wire n10620;
    wire n10623;
    wire n10626;
    wire n10629;
    wire n10632;
    wire n10635;
    wire n10638;
    wire n10641;
    wire n10644;
    wire n10647;
    wire n10649;
    wire n10652;
    wire n10655;
    wire n10658;
    wire n10662;
    wire n10665;
    wire n10668;
    wire n10671;
    wire n10674;
    wire n10677;
    wire n10680;
    wire n10683;
    wire n10686;
    wire n10689;
    wire n10692;
    wire n10695;
    wire n10698;
    wire n10701;
    wire n10704;
    wire n10707;
    wire n10710;
    wire n10713;
    wire n10715;
    wire n10719;
    wire n10722;
    wire n10725;
    wire n10728;
    wire n10731;
    wire n10734;
    wire n10737;
    wire n10740;
    wire n10743;
    wire n10746;
    wire n10749;
    wire n10752;
    wire n10755;
    wire n10758;
    wire n10761;
    wire n10764;
    wire n10767;
    wire n10770;
    wire n10773;
    wire n10776;
    wire n10779;
    wire n10782;
    wire n10785;
    wire n10788;
    wire n10791;
    wire n10794;
    wire n10797;
    wire n10800;
    wire n10803;
    wire n10806;
    wire n10809;
    wire n10812;
    wire n10815;
    wire n10818;
    wire n10821;
    wire n10824;
    wire n10827;
    wire n10830;
    wire n10833;
    wire n10836;
    wire n10839;
    wire n10842;
    wire n10845;
    wire n10848;
    wire n10851;
    wire n10854;
    wire n10857;
    wire n10860;
    wire n10863;
    wire n10866;
    wire n10869;
    wire n10872;
    wire n10875;
    wire n10878;
    wire n10881;
    wire n10884;
    wire n10887;
    wire n10890;
    wire n10893;
    wire n10896;
    wire n10899;
    wire n10902;
    wire n10905;
    wire n10908;
    wire n10911;
    wire n10914;
    wire n10917;
    wire n10920;
    wire n10923;
    wire n10926;
    wire n10929;
    wire n10932;
    wire n10935;
    wire n10938;
    wire n10941;
    wire n10944;
    wire n10947;
    wire n10950;
    wire n10953;
    wire n10956;
    wire n10959;
    wire n10962;
    wire n10964;
    wire n10968;
    wire n10971;
    wire n10974;
    wire n10977;
    wire n10980;
    wire n10983;
    wire n10986;
    wire n10989;
    wire n10992;
    wire n10995;
    wire n10998;
    wire n11001;
    wire n11004;
    wire n11007;
    wire n11010;
    wire n11013;
    wire n11016;
    wire n11019;
    wire n11022;
    wire n11025;
    wire n11028;
    wire n11031;
    wire n11034;
    wire n11037;
    wire n11040;
    wire n11043;
    wire n11046;
    wire n11049;
    wire n11052;
    wire n11055;
    wire n11058;
    wire n11061;
    wire n11064;
    wire n11067;
    wire n11070;
    wire n11073;
    wire n11076;
    wire n11079;
    wire n11082;
    wire n11085;
    wire n11088;
    wire n11091;
    wire n11094;
    wire n11097;
    wire n11100;
    wire n11103;
    wire n11105;
    wire n11108;
    wire n11111;
    wire n11114;
    wire n11117;
    wire n11120;
    wire n11123;
    wire n11126;
    wire n11129;
    wire n11132;
    wire n11135;
    wire n11138;
    wire n11141;
    wire n11144;
    wire n11147;
    wire n11150;
    wire n11153;
    wire n11156;
    wire n11159;
    wire n11162;
    wire n11165;
    wire n11168;
    wire n11171;
    wire n11174;
    wire n11177;
    wire n11181;
    wire n11184;
    wire n11187;
    wire n11190;
    wire n11193;
    wire n11196;
    wire n11199;
    wire n11202;
    wire n11205;
    wire n11208;
    wire n11211;
    wire n11214;
    wire n11217;
    wire n11220;
    wire n11223;
    wire n11226;
    wire n11229;
    wire n11232;
    wire n11235;
    wire n11238;
    wire n11241;
    wire n11244;
    wire n11247;
    wire n11250;
    wire n11253;
    wire n11256;
    wire n11259;
    wire n11262;
    wire n11265;
    wire n11268;
    wire n11271;
    wire n11274;
    wire n11277;
    wire n11280;
    wire n11282;
    wire n11285;
    wire n11288;
    wire n11291;
    wire n11294;
    wire n11297;
    wire n11300;
    wire n11303;
    wire n11306;
    wire n11309;
    wire n11312;
    wire n11315;
    wire n11318;
    wire n11321;
    wire n11324;
    wire n11327;
    wire n11330;
    wire n11333;
    wire n11337;
    wire n11339;
    wire n11342;
    wire n11345;
    wire n11348;
    wire n11351;
    wire n11354;
    wire n11357;
    wire n11360;
    wire n11363;
    wire n11366;
    wire n11369;
    wire n11372;
    wire n11375;
    wire n11379;
    wire n11382;
    wire n11385;
    wire n11388;
    wire n11391;
    wire n11394;
    wire n11397;
    wire n11400;
    wire n11403;
    wire n11406;
    wire n11409;
    wire n11412;
    wire n11415;
    wire n11418;
    wire n11421;
    wire n11424;
    wire n11427;
    wire n11429;
    wire n11433;
    wire n11436;
    wire n11439;
    wire n11441;
    wire n11444;
    wire n11447;
    wire n11450;
    wire n11453;
    wire n11456;
    wire n11459;
    wire n11462;
    wire n11465;
    wire n11468;
    wire n11471;
    wire n11474;
    wire n11477;
    wire n11480;
    wire n11483;
    wire n11487;
    wire n11490;
    wire n11493;
    wire n11496;
    wire n11499;
    wire n11502;
    wire n11505;
    wire n11508;
    wire n11511;
    wire n11514;
    wire n11517;
    wire n11520;
    wire n11523;
    wire n11526;
    wire n11529;
    wire n11532;
    wire n11535;
    wire n11538;
    wire n11541;
    wire n11544;
    wire n11547;
    wire n11550;
    wire n11553;
    wire n11556;
    wire n11559;
    wire n11562;
    wire n11565;
    wire n11568;
    wire n11571;
    wire n11574;
    wire n11577;
    wire n11580;
    wire n11583;
    wire n11586;
    wire n11589;
    wire n11592;
    wire n11594;
    wire n11597;
    wire n11601;
    wire n11604;
    wire n11607;
    wire n11610;
    wire n11613;
    wire n11615;
    wire n11618;
    wire n11621;
    wire n11624;
    wire n11627;
    wire n11630;
    wire n11633;
    wire n11636;
    wire n11639;
    wire n11642;
    wire n11645;
    wire n11648;
    wire n11651;
    wire n11654;
    wire n11657;
    wire n11660;
    wire n11663;
    wire n11666;
    wire n11669;
    wire n11672;
    wire n11675;
    wire n11678;
    wire n11681;
    wire n11684;
    wire n11687;
    wire n11690;
    wire n11693;
    wire n11696;
    wire n11699;
    wire n11703;
    wire n11706;
    wire n11709;
    wire n11712;
    wire n11715;
    wire n11718;
    wire n11721;
    wire n11724;
    wire n11727;
    wire n11730;
    wire n11733;
    wire n11736;
    wire n11739;
    wire n11742;
    wire n11745;
    wire n11748;
    wire n11751;
    wire n11754;
    wire n11756;
    wire n11759;
    wire n11762;
    wire n11765;
    wire n11768;
    wire n11772;
    wire n11775;
    wire n11778;
    wire n11781;
    wire n11784;
    wire n11787;
    wire n11790;
    wire n11793;
    wire n11796;
    wire n11799;
    wire n11802;
    wire n11805;
    wire n11808;
    wire n11811;
    wire n11814;
    wire n11817;
    wire n11820;
    wire n11823;
    wire n11826;
    wire n11828;
    wire n11831;
    wire n11834;
    wire n11837;
    wire n11840;
    wire n11843;
    wire n11847;
    wire n11850;
    wire n11853;
    wire n11856;
    wire n11859;
    wire n11862;
    wire n11865;
    wire n11868;
    wire n11871;
    wire n11874;
    wire n11877;
    wire n11880;
    wire n11883;
    wire n11885;
    wire n11888;
    wire n11891;
    wire n11894;
    wire n11897;
    wire n11900;
    wire n11903;
    wire n11906;
    wire n11909;
    wire n11912;
    wire n11915;
    wire n11918;
    wire n11921;
    wire n11924;
    wire n11927;
    wire n11930;
    wire n11933;
    wire n11936;
    wire n11939;
    wire n11942;
    wire n11945;
    wire n11948;
    wire n11951;
    wire n11954;
    wire n11957;
    wire n11960;
    wire n11963;
    wire n11967;
    wire n11970;
    wire n11973;
    wire n11976;
    wire n11979;
    wire n11982;
    wire n11985;
    wire n11988;
    wire n11991;
    wire n11994;
    wire n11997;
    wire n12000;
    wire n12003;
    wire n12006;
    wire n12009;
    wire n12012;
    wire n12015;
    wire n12018;
    wire n12021;
    wire n12024;
    wire n12027;
    wire n12030;
    wire n12033;
    wire n12036;
    wire n12039;
    wire n12042;
    wire n12045;
    wire n12048;
    wire n12051;
    wire n12054;
    wire n12057;
    wire n12060;
    wire n12063;
    wire n12066;
    wire n12069;
    wire n12072;
    wire n12075;
    wire n12078;
    wire n12081;
    wire n12084;
    wire n12087;
    wire n12090;
    wire n12093;
    wire n12096;
    wire n12099;
    wire n12102;
    wire n12105;
    wire n12108;
    wire n12111;
    wire n12114;
    wire n12117;
    wire n12120;
    wire n12123;
    wire n12126;
    wire n12129;
    wire n12132;
    wire n12135;
    wire n12138;
    wire n12140;
    wire n12143;
    wire n12146;
    wire n12149;
    wire n12152;
    wire n12155;
    wire n12158;
    wire n12161;
    wire n12164;
    wire n12167;
    wire n12170;
    wire n12173;
    wire n12176;
    wire n12179;
    wire n12182;
    wire n12185;
    wire n12188;
    wire n12191;
    wire n12194;
    wire n12197;
    wire n12200;
    wire n12203;
    wire n12206;
    wire n12209;
    wire n12212;
    wire n12215;
    wire n12218;
    wire n12221;
    wire n12224;
    wire n12227;
    wire n12230;
    wire n12233;
    wire n12236;
    wire n12239;
    wire n12242;
    wire n12245;
    wire n12249;
    wire n12252;
    wire n12255;
    wire n12258;
    wire n12261;
    wire n12264;
    wire n12266;
    wire n12269;
    wire n12272;
    wire n12275;
    wire n12278;
    wire n12281;
    wire n12284;
    wire n12287;
    wire n12290;
    wire n12293;
    wire n12296;
    wire n12299;
    wire n12302;
    wire n12305;
    wire n12308;
    wire n12311;
    wire n12314;
    wire n12317;
    wire n12320;
    wire n12323;
    wire n12326;
    wire n12329;
    wire n12332;
    wire n12335;
    wire n12338;
    wire n12341;
    wire n12344;
    wire n12347;
    wire n12350;
    wire n12353;
    wire n12356;
    wire n12359;
    wire n12362;
    wire n12365;
    wire n12368;
    wire n12371;
    wire n12374;
    wire n12377;
    wire n12380;
    wire n12384;
    wire n12387;
    wire n12390;
    wire n12393;
    wire n12396;
    wire n12399;
    wire n12402;
    wire n12404;
    wire n12407;
    wire n12411;
    wire n12414;
    wire n12417;
    wire n12420;
    wire n12423;
    wire n12426;
    wire n12429;
    wire n12432;
    wire n12435;
    wire n12438;
    wire n12441;
    wire n12444;
    wire n12447;
    wire n12450;
    wire n12453;
    wire n12456;
    wire n12459;
    wire n12462;
    wire n12465;
    wire n12468;
    wire n12471;
    wire n12474;
    wire n12477;
    wire n12479;
    wire n12482;
    wire n12485;
    wire n12488;
    wire n12491;
    wire n12494;
    wire n12497;
    wire n12500;
    wire n12503;
    wire n12506;
    wire n12509;
    wire n12512;
    wire n12515;
    wire n12518;
    wire n12521;
    wire n12524;
    wire n12527;
    wire n12530;
    wire n12533;
    wire n12536;
    wire n12539;
    wire n12542;
    wire n12545;
    wire n12548;
    wire n12551;
    wire n12554;
    wire n12557;
    wire n12560;
    wire n12563;
    wire n12566;
    wire n12569;
    wire n12572;
    wire n12575;
    wire n12578;
    wire n12581;
    wire n12584;
    wire n12588;
    wire n12591;
    wire n12594;
    wire n12597;
    wire n12600;
    wire n12603;
    wire n12605;
    wire n12608;
    wire n12611;
    wire n12614;
    wire n12617;
    wire n12620;
    wire n12623;
    wire n12626;
    wire n12629;
    wire n12632;
    wire n12635;
    wire n12638;
    wire n12641;
    wire n12644;
    wire n12647;
    wire n12650;
    wire n12653;
    wire n12656;
    wire n12659;
    wire n12662;
    wire n12665;
    wire n12668;
    wire n12671;
    wire n12674;
    wire n12677;
    wire n12680;
    wire n12683;
    wire n12686;
    wire n12689;
    wire n12692;
    wire n12695;
    wire n12698;
    wire n12701;
    wire n12704;
    wire n12707;
    wire n12710;
    wire n12713;
    wire n12716;
    wire n12719;
    wire n12723;
    wire n12726;
    wire n12729;
    wire n12732;
    wire n12735;
    wire n12738;
    wire n12741;
    wire n12743;
    wire n12746;
    wire n12750;
    wire n12753;
    wire n12756;
    wire n12759;
    wire n12762;
    wire n12765;
    wire n12768;
    wire n12771;
    wire n12774;
    wire n12777;
    wire n12780;
    wire n12783;
    wire n12786;
    wire n12789;
    wire n12792;
    wire n12795;
    wire n12798;
    wire n12801;
    wire n12804;
    wire n12807;
    wire n12810;
    wire n12813;
    wire n12816;
    wire n12819;
    wire n12822;
    wire n12825;
    wire n12828;
    wire n12831;
    wire n12834;
    wire n12837;
    wire n12840;
    wire n12843;
    wire n12846;
    wire n12849;
    wire n12852;
    wire n12855;
    wire n12858;
    wire n12861;
    wire n12864;
    wire n12866;
    wire n12869;
    wire n12872;
    wire n12875;
    wire n12878;
    wire n12881;
    wire n12884;
    wire n12887;
    wire n12890;
    wire n12893;
    wire n12896;
    wire n12899;
    wire n12902;
    wire n12905;
    wire n12908;
    wire n12911;
    wire n12914;
    wire n12917;
    wire n12920;
    wire n12923;
    wire n12926;
    wire n12929;
    wire n12932;
    wire n12935;
    wire n12938;
    wire n12941;
    wire n12944;
    wire n12947;
    wire n12950;
    wire n12953;
    wire n12956;
    wire n12959;
    wire n12962;
    wire n12965;
    wire n12968;
    wire n12971;
    wire n12974;
    wire n12977;
    wire n12980;
    wire n12983;
    wire n12986;
    wire n12989;
    wire n12992;
    wire n12995;
    wire n12998;
    wire n13001;
    wire n13004;
    wire n13008;
    wire n13011;
    wire n13014;
    wire n13017;
    wire n13020;
    wire n13023;
    wire n13026;
    wire n13029;
    wire n13032;
    wire n13035;
    wire n13038;
    wire n13041;
    wire n13044;
    wire n13047;
    wire n13050;
    wire n13053;
    wire n13056;
    wire n13059;
    wire n13062;
    wire n13064;
    wire n13067;
    wire n13070;
    wire n13073;
    wire n13076;
    wire n13079;
    wire n13082;
    wire n13085;
    wire n13088;
    wire n13091;
    wire n13094;
    wire n13097;
    wire n13100;
    wire n13103;
    wire n13106;
    wire n13109;
    wire n13112;
    wire n13115;
    wire n13118;
    wire n13121;
    wire n13124;
    wire n13127;
    wire n13130;
    wire n13133;
    wire n13136;
    wire n13139;
    wire n13142;
    wire n13145;
    wire n13148;
    wire n13151;
    wire n13154;
    wire n13157;
    wire n13160;
    wire n13163;
    wire n13166;
    wire n13169;
    wire n13172;
    wire n13175;
    wire n13178;
    wire n13181;
    wire n13184;
    wire n13187;
    wire n13190;
    wire n13193;
    wire n13196;
    wire n13199;
    wire n13202;
    wire n13205;
    wire n13208;
    wire n13211;
    wire n13214;
    wire n13217;
    wire n13220;
    wire n13223;
    wire n13226;
    wire n13229;
    wire n13233;
    wire n13236;
    wire n13239;
    wire n13242;
    wire n13245;
    wire n13248;
    wire n13251;
    wire n13254;
    wire n13257;
    wire n13260;
    wire n13263;
    wire n13266;
    wire n13269;
    wire n13272;
    wire n13275;
    wire n13278;
    wire n13281;
    wire n13284;
    wire n13287;
    wire n13290;
    wire n13293;
    wire n13296;
    wire n13299;
    wire n13302;
    wire n13305;
    wire n13308;
    wire n13311;
    wire n13314;
    wire n13317;
    wire n13320;
    wire n13323;
    wire n13326;
    wire n13329;
    wire n13332;
    wire n13335;
    wire n13338;
    wire n13341;
    wire n13344;
    wire n13347;
    wire n13350;
    wire n13353;
    wire n13356;
    wire n13359;
    wire n13362;
    wire n13365;
    wire n13368;
    wire n13371;
    wire n13374;
    wire n13377;
    wire n13380;
    wire n13383;
    wire n13386;
    wire n13389;
    wire n13392;
    wire n13395;
    wire n13398;
    wire n13401;
    wire n13404;
    wire n13407;
    wire n13410;
    wire n13413;
    wire n13415;
    wire n13418;
    wire n13421;
    wire n13424;
    wire n13427;
    wire n13430;
    wire n13433;
    wire n13436;
    wire n13439;
    wire n13442;
    wire n13445;
    wire n13448;
    wire n13451;
    wire n13454;
    wire n13457;
    wire n13460;
    wire n13463;
    wire n13466;
    wire n13469;
    wire n13472;
    wire n13476;
    wire n13479;
    wire n13482;
    wire n13485;
    wire n13488;
    wire n13491;
    wire n13493;
    wire n13497;
    wire n13500;
    wire n13503;
    wire n13506;
    wire n13509;
    wire n13512;
    wire n13515;
    wire n13518;
    wire n13521;
    wire n13524;
    wire n13527;
    wire n13530;
    wire n13532;
    wire n13535;
    wire n13538;
    wire n13542;
    wire n13545;
    wire n13548;
    wire n13551;
    wire n13554;
    wire n13557;
    wire n13560;
    wire n13563;
    wire n13566;
    wire n13569;
    wire n13572;
    wire n13575;
    wire n13578;
    wire n13581;
    wire n13584;
    wire n13587;
    wire n13590;
    wire n13593;
    wire n13596;
    wire n13598;
    wire n13601;
    wire n13604;
    wire n13608;
    wire n13610;
    wire n13613;
    wire n13616;
    wire n13619;
    wire n13622;
    wire n13625;
    wire n13628;
    wire n13631;
    wire n13634;
    wire n13637;
    wire n13640;
    wire n13643;
    wire n13646;
    wire n13649;
    wire n13652;
    wire n13655;
    wire n13658;
    wire n13661;
    wire n13664;
    wire n13667;
    wire n13671;
    wire n13674;
    wire n13677;
    wire n13680;
    wire n13683;
    wire n13686;
    wire n13689;
    wire n13692;
    wire n13695;
    wire n13697;
    wire n13700;
    wire n13703;
    wire n13706;
    wire n13709;
    wire n13712;
    wire n13715;
    wire n13718;
    wire n13721;
    wire n13724;
    wire n13727;
    wire n13730;
    wire n13733;
    wire n13736;
    wire n13739;
    wire n13742;
    wire n13745;
    wire n13748;
    wire n13751;
    wire n13754;
    wire n13757;
    wire n13760;
    wire n13763;
    wire n13766;
    wire n13769;
    wire n13772;
    wire n13775;
    wire n13779;
    wire n13782;
    wire n13785;
    wire n13788;
    wire n13791;
    wire n13793;
    wire n13796;
    wire n13799;
    wire n13802;
    wire n13805;
    wire n13809;
    wire n13812;
    wire n13815;
    wire n13818;
    wire n13821;
    wire n13824;
    wire n13827;
    wire n13830;
    wire n13833;
    wire n13836;
    wire n13838;
    wire n13841;
    wire n13844;
    wire n13847;
    wire n13850;
    wire n13853;
    wire n13856;
    wire n13859;
    wire n13862;
    wire n13865;
    wire n13869;
    wire n13871;
    wire n13874;
    wire n13877;
    wire n13880;
    wire n13883;
    wire n13886;
    wire n13889;
    wire n13892;
    wire n13895;
    wire n13899;
    wire n13901;
    wire n13904;
    wire n13907;
    wire n13910;
    wire n13913;
    wire n13916;
    wire n13919;
    wire n13922;
    wire n13925;
    wire n13928;
    wire n13931;
    wire n13934;
    wire n13937;
    wire n13940;
    wire n13943;
    wire n13946;
    wire n13950;
    wire n13953;
    wire n13955;
    wire n13958;
    wire n13961;
    wire n13964;
    wire n13967;
    wire n13970;
    wire n13973;
    wire n13976;
    wire n13979;
    wire n13982;
    wire n13985;
    wire n13988;
    wire n13991;
    wire n13995;
    wire n13998;
    wire n14000;
    wire n14003;
    wire n14006;
    wire n14009;
    wire n14012;
    wire n14015;
    wire n14018;
    wire n14021;
    wire n14024;
    wire n14027;
    wire n14030;
    wire n14033;
    wire n14037;
    wire n14040;
    wire n14043;
    wire n14046;
    wire n14049;
    wire n14051;
    wire n14054;
    wire n14057;
    wire n14060;
    wire n14063;
    wire n14066;
    wire n14069;
    wire n14073;
    wire n14075;
    wire n14078;
    wire n14081;
    wire n14085;
    wire n14087;
    wire n14090;
    wire n14093;
    wire n14096;
    wire n14099;
    wire n14102;
    wire n14105;
    wire n14108;
    wire n14111;
    wire n14114;
    wire n14117;
    wire n14120;
    wire n14123;
    wire n14126;
    wire n14129;
    wire n14132;
    wire n14135;
    wire n14138;
    wire n14141;
    wire n14145;
    wire n14148;
    wire n14151;
    wire n14154;
    wire n14157;
    wire n14160;
    wire n14163;
    wire n14166;
    wire n14169;
    wire n14172;
    wire n14175;
    wire n14178;
    wire n14181;
    wire n14184;
    wire n14187;
    wire n14189;
    wire n14192;
    wire n14195;
    wire n14198;
    wire n14201;
    wire n14204;
    wire n14207;
    wire n14210;
    wire n14213;
    wire n14216;
    wire n14219;
    wire n14222;
    wire n14225;
    wire n14228;
    wire n14231;
    wire n14234;
    wire n14237;
    wire n14240;
    wire n14243;
    wire n14246;
    wire n14249;
    wire n14252;
    wire n14255;
    wire n14258;
    wire n14261;
    wire n14264;
    wire n14267;
    wire n14270;
    wire n14273;
    wire n14276;
    wire n14279;
    wire n14282;
    wire n14286;
    wire n14288;
    wire n14291;
    wire n14294;
    wire n14297;
    wire n14300;
    wire n14303;
    wire n14306;
    wire n14309;
    wire n14312;
    wire n14315;
    wire n14319;
    wire n14322;
    wire n14324;
    wire n14327;
    wire n14330;
    wire n14333;
    wire n14336;
    wire n14339;
    wire n14342;
    wire n14345;
    wire n14348;
    wire n14351;
    wire n14354;
    wire n14357;
    wire n14360;
    wire n14363;
    wire n14366;
    wire n14369;
    wire n14372;
    wire n14375;
    wire n14378;
    wire n14381;
    wire n14384;
    wire n14387;
    wire n14390;
    wire n14393;
    wire n14396;
    wire n14399;
    wire n14402;
    wire n14405;
    wire n14408;
    wire n14411;
    wire n14415;
    wire n14418;
    wire n14421;
    wire n14424;
    wire n14426;
    wire n14429;
    wire n14432;
    wire n14435;
    wire n14438;
    wire n14441;
    wire n14444;
    wire n14447;
    wire n14450;
    wire n14453;
    wire n14456;
    wire n14459;
    wire n14462;
    wire n14465;
    wire n14469;
    wire n14472;
    wire n14474;
    wire n14478;
    wire n14480;
    wire n14483;
    wire n14486;
    wire n14489;
    wire n14493;
    wire n14495;
    wire n14498;
    wire n14501;
    wire n14504;
    wire n14507;
    wire n14510;
    wire n14513;
    wire n14516;
    wire n14519;
    wire n14522;
    wire n14525;
    wire n14528;
    wire n14532;
    wire n14535;
    wire n14538;
    wire n14541;
    wire n14544;
    wire n14546;
    wire n14549;
    wire n14552;
    wire n14555;
    wire n14558;
    wire n14561;
    wire n14564;
    wire n14567;
    wire n14570;
    wire n14573;
    wire n14576;
    wire n14579;
    wire n14583;
    wire n14586;
    wire n14588;
    wire n14591;
    wire n14594;
    wire n14597;
    wire n14600;
    wire n14603;
    wire n14606;
    wire n14609;
    wire n14612;
    wire n14615;
    wire n14618;
    wire n14621;
    wire n14624;
    wire n14627;
    wire n14630;
    wire n14633;
    wire n14636;
    wire n14640;
    wire n14643;
    wire n14645;
    wire n14648;
    wire n14651;
    wire n14654;
    wire n14657;
    wire n14660;
    wire n14663;
    wire n14666;
    wire n14669;
    wire n14672;
    wire n14675;
    wire n14678;
    wire n14681;
    wire n14684;
    wire n14687;
    wire n14690;
    wire n14693;
    wire n14696;
    wire n14699;
    wire n14702;
    wire n14705;
    wire n14708;
    wire n14711;
    wire n14714;
    wire n14717;
    wire n14720;
    wire n14723;
    wire n14726;
    wire n14729;
    wire n14732;
    wire n14735;
    wire n14738;
    wire n14741;
    wire n14744;
    wire n14747;
    wire n14750;
    wire n14753;
    wire n14756;
    wire n14759;
    wire n14762;
    wire n14765;
    wire n14768;
    wire n14771;
    wire n14774;
    wire n14777;
    wire n14780;
    wire n14783;
    wire n14786;
    wire n14789;
    wire n14792;
    wire n14795;
    wire n14798;
    wire n14801;
    wire n14804;
    wire n14807;
    wire n14810;
    wire n14813;
    wire n14816;
    wire n14819;
    wire n14822;
    wire n14825;
    wire n14828;
    wire n14831;
    wire n14834;
    wire n14837;
    wire n14840;
    wire n14843;
    wire n14846;
    wire n14849;
    wire n14853;
    wire n14856;
    wire n14859;
    wire n14862;
    wire n14865;
    wire n14868;
    wire n14871;
    wire n14874;
    wire n14877;
    wire n14880;
    wire n14883;
    wire n14886;
    wire n14889;
    wire n14892;
    wire n14895;
    wire n14898;
    wire n14901;
    wire n14904;
    wire n14907;
    wire n14910;
    wire n14913;
    wire n14916;
    wire n14919;
    wire n14922;
    wire n14925;
    wire n14928;
    wire n14931;
    wire n14934;
    wire n14937;
    wire n14940;
    wire n14943;
    wire n14946;
    wire n14949;
    wire n14952;
    wire n14955;
    wire n14958;
    wire n14961;
    wire n14964;
    wire n14967;
    wire n14970;
    wire n14973;
    wire n14976;
    wire n14979;
    wire n14982;
    wire n14985;
    wire n14988;
    wire n14991;
    wire n14994;
    wire n14997;
    wire n15000;
    wire n15003;
    wire n15006;
    wire n15009;
    wire n15012;
    wire n15015;
    wire n15018;
    wire n15021;
    wire n15024;
    wire n15027;
    wire n15030;
    wire n15033;
    wire n15036;
    wire n15039;
    wire n15042;
    wire n15045;
    wire n15048;
    wire n15051;
    wire n15054;
    wire n15057;
    wire n15060;
    wire n15063;
    wire n15066;
    wire n15069;
    wire n15072;
    wire n15075;
    wire n15078;
    wire n15080;
    wire n15083;
    wire n15087;
    wire n15090;
    wire n15093;
    wire n15096;
    wire n15098;
    wire n15101;
    wire n15104;
    wire n15107;
    wire n15110;
    wire n15113;
    wire n15117;
    wire n15120;
    wire n15123;
    wire n15125;
    wire n15128;
    wire n15132;
    wire n15135;
    wire n15138;
    wire n15141;
    wire n15144;
    wire n15147;
    wire n15150;
    wire n15153;
    wire n15156;
    wire n15159;
    wire n15162;
    wire n15165;
    wire n15168;
    wire n15171;
    wire n15173;
    wire n15176;
    wire n15179;
    wire n15182;
    wire n15185;
    wire n15188;
    wire n15191;
    wire n15194;
    wire n15197;
    wire n15200;
    wire n15203;
    wire n15206;
    wire n15209;
    wire n15212;
    wire n15215;
    wire n15218;
    wire n15221;
    wire n15224;
    wire n15227;
    wire n15230;
    wire n15233;
    wire n15236;
    wire n15239;
    wire n15242;
    wire n15245;
    wire n15248;
    wire n15251;
    wire n15254;
    wire n15257;
    wire n15260;
    wire n15264;
    wire n15267;
    wire n15269;
    wire n15272;
    wire n15275;
    wire n15278;
    wire n15282;
    wire n15285;
    wire n15288;
    wire n15291;
    wire n15294;
    wire n15296;
    wire n15300;
    wire n15303;
    wire n15305;
    wire n15308;
    wire n15311;
    wire n15314;
    wire n15317;
    wire n15320;
    wire n15323;
    wire n15326;
    wire n15329;
    wire n15333;
    wire n15336;
    wire n15339;
    wire n15341;
    wire n15344;
    wire n15347;
    wire n15350;
    wire n15353;
    wire n15357;
    wire n15360;
    wire n15363;
    wire n15365;
    wire n15369;
    wire n15372;
    wire n15374;
    wire n15377;
    wire n15380;
    wire n15383;
    wire n15386;
    wire n15389;
    wire n15392;
    wire n15395;
    wire n15398;
    wire n15401;
    wire n15404;
    wire n15407;
    wire n15410;
    wire n15413;
    wire n15416;
    wire n15419;
    wire n15422;
    wire n15426;
    wire n15429;
    wire n15431;
    wire n15434;
    wire n15437;
    wire n15440;
    wire n15443;
    wire n15446;
    wire n15449;
    wire n15452;
    wire n15455;
    wire n15458;
    wire n15461;
    wire n15464;
    wire n15467;
    wire n15470;
    wire n15473;
    wire n15476;
    wire n15479;
    wire n15482;
    wire n15485;
    wire n15488;
    wire n15491;
    wire n15494;
    wire n15497;
    wire n15500;
    wire n15503;
    wire n15506;
    wire n15510;
    wire n15513;
    wire n15516;
    wire n15519;
    wire n15522;
    wire n15525;
    wire n15528;
    wire n15531;
    wire n15534;
    wire n15536;
    wire n15539;
    wire n15542;
    wire n15545;
    wire n15548;
    wire n15551;
    wire n15554;
    wire n15557;
    wire n15560;
    wire n15563;
    wire n15566;
    wire n15569;
    wire n15572;
    wire n15575;
    wire n15578;
    wire n15581;
    wire n15585;
    wire n15587;
    wire n15590;
    wire n15593;
    wire n15596;
    wire n15599;
    wire n15602;
    wire n15606;
    wire n15609;
    wire n15612;
    wire n15615;
    wire n15618;
    wire n15621;
    wire n15624;
    wire n15627;
    wire n15630;
    wire n15633;
    wire n15636;
    wire n15639;
    wire n15641;
    wire n15644;
    wire n15647;
    wire n15650;
    wire n15653;
    wire n15656;
    wire n15659;
    wire n15662;
    wire n15665;
    wire n15668;
    wire n15671;
    wire n15674;
    wire n15678;
    wire n15680;
    wire n15684;
    wire n15686;
    wire n15689;
    wire n15692;
    wire n15695;
    wire n15698;
    wire n15701;
    wire n15704;
    wire n15707;
    wire n15710;
    wire n15713;
    wire n15716;
    wire n15719;
    wire n15722;
    wire n15725;
    wire n15728;
    wire n15731;
    wire n15734;
    wire n15737;
    wire n15741;
    wire n15744;
    wire n15746;
    wire n15749;
    wire n15752;
    wire n15755;
    wire n15758;
    wire n15761;
    wire n15764;
    wire n15767;
    wire n15770;
    wire n15773;
    wire n15776;
    wire n15779;
    wire n15782;
    wire n15785;
    wire n15788;
    wire n15791;
    wire n15794;
    wire n15797;
    wire n15800;
    wire n15803;
    wire n15806;
    wire n15809;
    wire n15812;
    wire n15815;
    wire n15818;
    wire n15821;
    wire n15824;
    wire n15827;
    wire n15830;
    wire n15833;
    wire n15836;
    wire n15839;
    wire n15842;
    wire n15845;
    wire n15848;
    wire n15851;
    wire n15854;
    wire n15857;
    wire n15860;
    wire n15863;
    wire n15866;
    wire n15869;
    wire n15872;
    wire n15875;
    wire n15878;
    wire n15881;
    wire n15885;
    wire n15888;
    wire n15891;
    wire n15893;
    wire n15896;
    wire n15899;
    wire n15902;
    wire n15905;
    wire n15908;
    wire n15911;
    wire n15914;
    wire n15918;
    wire n15921;
    wire n15923;
    wire n15926;
    wire n15930;
    wire n15933;
    wire n15935;
    wire n15938;
    wire n15941;
    wire n15944;
    wire n15947;
    wire n15951;
    wire n15954;
    wire n15956;
    wire n15959;
    wire n15962;
    wire n15965;
    wire n15968;
    wire n15971;
    wire n15974;
    wire n15977;
    wire n15980;
    wire n15983;
    wire n15986;
    wire n15990;
    wire n15993;
    wire n15995;
    wire n15998;
    wire n16001;
    wire n16004;
    wire n16007;
    wire n16010;
    wire n16013;
    wire n16016;
    wire n16020;
    wire n16023;
    wire n16026;
    wire n16029;
    wire n16031;
    wire n16034;
    wire n16037;
    wire n16040;
    wire n16043;
    wire n16046;
    wire n16049;
    wire n16052;
    wire n16055;
    wire n16058;
    wire n16062;
    wire n16065;
    wire n16068;
    wire n16070;
    wire n16073;
    wire n16076;
    wire n16079;
    wire n16083;
    wire n16085;
    wire n16088;
    wire n16091;
    wire n16094;
    wire n16097;
    wire n16100;
    wire n16103;
    wire n16107;
    wire n16110;
    wire n16113;
    wire n16115;
    wire n16119;
    wire n16121;
    wire n16124;
    wire n16127;
    wire n16130;
    wire n16133;
    wire n16136;
    wire n16139;
    wire n16142;
    wire n16145;
    wire n16148;
    wire n16151;
    wire n16155;
    wire n16158;
    wire n16160;
    wire n16163;
    wire n16166;
    wire n16169;
    wire n16172;
    wire n16175;
    wire n16178;
    wire n16181;
    wire n16184;
    wire n16187;
    wire n16190;
    wire n16193;
    wire n16196;
    wire n16199;
    wire n16202;
    wire n16206;
    wire n16209;
    wire n16211;
    wire n16214;
    wire n16217;
    wire n16220;
    wire n16223;
    wire n16226;
    wire n16229;
    wire n16232;
    wire n16235;
    wire n16238;
    wire n16241;
    wire n16244;
    wire n16247;
    wire n16250;
    wire n16253;
    wire n16256;
    wire n16259;
    wire n16262;
    wire n16265;
    wire n16268;
    wire n16271;
    wire n16274;
    wire n16277;
    wire n16280;
    wire n16283;
    wire n16286;
    wire n16289;
    wire n16292;
    wire n16295;
    wire n16298;
    wire n16301;
    wire n16304;
    wire n16307;
    wire n16310;
    wire n16313;
    wire n16316;
    wire n16319;
    wire n16322;
    wire n16325;
    wire n16328;
    wire n16331;
    wire n16334;
    wire n16337;
    wire n16340;
    wire n16343;
    wire n16346;
    wire n16349;
    wire n16352;
    wire n16355;
    wire n16358;
    wire n16361;
    wire n16364;
    wire n16367;
    wire n16370;
    wire n16373;
    wire n16376;
    wire n16379;
    wire n16382;
    wire n16385;
    wire n16388;
    wire n16391;
    wire n16394;
    wire n16397;
    wire n16400;
    wire n16403;
    wire n16406;
    wire n16409;
    wire n16412;
    wire n16415;
    wire n16418;
    wire n16421;
    wire n16424;
    wire n16427;
    wire n16430;
    wire n16433;
    wire n16436;
    wire n16439;
    wire n16442;
    wire n16445;
    wire n16448;
    wire n16451;
    wire n16454;
    wire n16457;
    wire n16460;
    wire n16463;
    wire n16466;
    wire n16469;
    wire n16472;
    wire n16475;
    wire n16478;
    wire n16481;
    wire n16484;
    wire n16487;
    wire n16491;
    wire n16494;
    wire n16497;
    wire n16500;
    wire n16503;
    wire n16506;
    wire n16509;
    wire n16512;
    wire n16515;
    wire n16518;
    wire n16521;
    wire n16524;
    wire n16527;
    wire n16530;
    wire n16533;
    wire n16536;
    wire n16539;
    wire n16542;
    wire n16545;
    wire n16548;
    wire n16551;
    wire n16554;
    wire n16557;
    wire n16560;
    wire n16562;
    wire n16565;
    wire n16568;
    wire n16571;
    wire n16574;
    wire n16577;
    wire n16580;
    wire n16583;
    wire n16586;
    wire n16589;
    wire n16592;
    wire n16595;
    wire n16598;
    wire n16601;
    wire n16604;
    wire n16607;
    wire n16610;
    wire n16613;
    wire n16616;
    wire n16619;
    wire n16622;
    wire n16625;
    wire n16628;
    wire n16631;
    wire n16634;
    wire n16637;
    wire n16640;
    wire n16643;
    wire n16646;
    wire n16649;
    wire n16652;
    wire n16655;
    wire n16658;
    wire n16661;
    wire n16664;
    wire n16667;
    wire n16670;
    wire n16673;
    wire n16676;
    wire n16679;
    wire n16682;
    wire n16685;
    wire n16688;
    wire n16691;
    wire n16694;
    wire n16697;
    wire n16700;
    wire n16703;
    wire n16706;
    wire n16709;
    wire n16712;
    wire n16715;
    wire n16718;
    wire n16721;
    wire n16724;
    wire n16727;
    wire n16730;
    wire n16733;
    wire n16736;
    wire n16739;
    wire n16742;
    wire n16745;
    wire n16748;
    wire n16751;
    wire n16754;
    wire n16757;
    wire n16760;
    wire n16763;
    wire n16766;
    wire n16769;
    wire n16772;
    wire n16775;
    wire n16778;
    wire n16781;
    wire n16787;
    wire n16790;
    wire n16793;
    wire n16796;
    wire n16799;
    wire n16802;
    wire n16805;
    wire n16808;
    wire n16811;
    wire n16814;
    wire n16817;
    wire n16820;
    wire n16823;
    wire n16826;
    wire n16829;
    wire n16832;
    wire n16835;
    wire n16838;
    wire n16841;
    wire n16844;
    wire n16847;
    wire n16850;
    wire n16853;
    wire n16856;
    wire n16862;
    wire n16865;
    wire n16868;
    wire n16871;
    wire n16874;
    wire n16877;
    wire n16880;
    wire n16883;
    wire n16886;
    wire n16889;
    wire n16892;
    wire n16895;
    wire n16898;
    wire n16901;
    wire n16904;
    wire n16907;
    wire n16910;
    wire n16913;
    wire n16916;
    wire n16919;
    wire n16922;
    wire n16925;
    wire n16928;
    wire n16931;
    wire n16937;
    wire n16940;
    wire n16943;
    wire n16946;
    wire n16949;
    wire n16952;
    wire n16955;
    wire n16958;
    wire n16961;
    wire n16964;
    wire n16967;
    wire n16970;
    wire n16973;
    wire n16976;
    wire n16979;
    wire n16982;
    wire n16985;
    wire n16988;
    wire n16991;
    wire n16994;
    wire n16997;
    wire n17000;
    wire n17003;
    wire n17006;
    wire n17012;
    wire n17015;
    wire n17018;
    wire n17021;
    wire n17024;
    wire n17027;
    wire n17030;
    wire n17033;
    wire n17036;
    wire n17039;
    wire n17042;
    wire n17045;
    wire n17048;
    wire n17051;
    wire n17054;
    wire n17057;
    wire n17060;
    wire n17063;
    wire n17066;
    wire n17069;
    wire n17072;
    wire n17075;
    wire n17078;
    wire n17081;
    wire n17087;
    wire n17090;
    wire n17093;
    wire n17096;
    wire n17099;
    wire n17102;
    wire n17105;
    wire n17108;
    wire n17111;
    wire n17114;
    wire n17117;
    wire n17120;
    wire n17123;
    wire n17126;
    wire n17129;
    wire n17132;
    wire n17135;
    wire n17138;
    wire n17141;
    wire n17144;
    wire n17147;
    wire n17150;
    wire n17153;
    wire n17156;
    wire n17162;
    wire n17165;
    wire n17168;
    wire n17171;
    wire n17174;
    wire n17177;
    wire n17180;
    wire n17183;
    wire n17186;
    wire n17189;
    wire n17192;
    wire n17195;
    wire n17198;
    wire n17201;
    wire n17204;
    wire n17207;
    wire n17210;
    wire n17213;
    wire n17216;
    wire n17219;
    wire n17222;
    wire n17225;
    wire n17228;
    wire n17231;
    wire n17237;
    wire n17240;
    wire n17243;
    wire n17246;
    wire n17249;
    wire n17252;
    wire n17255;
    wire n17258;
    wire n17261;
    wire n17264;
    wire n17267;
    wire n17270;
    wire n17273;
    wire n17276;
    wire n17279;
    wire n17282;
    wire n17285;
    wire n17288;
    wire n17291;
    wire n17294;
    wire n17297;
    wire n17300;
    wire n17303;
    wire n17306;
    wire n17312;
    wire n17315;
    wire n17318;
    wire n17321;
    wire n17324;
    wire n17327;
    wire n17330;
    wire n17333;
    wire n17336;
    wire n17339;
    wire n17342;
    wire n17345;
    wire n17348;
    wire n17351;
    wire n17354;
    wire n17357;
    wire n17360;
    wire n17363;
    wire n17366;
    wire n17369;
    wire n17372;
    wire n17375;
    wire n17378;
    wire n17381;
    wire n17387;
    wire n17390;
    wire n17393;
    wire n17396;
    wire n17399;
    wire n17402;
    wire n17405;
    wire n17408;
    wire n17411;
    wire n17414;
    wire n17417;
    wire n17420;
    wire n17423;
    wire n17426;
    wire n17429;
    wire n17432;
    wire n17435;
    wire n17438;
    wire n17441;
    wire n17444;
    wire n17447;
    wire n17450;
    wire n17453;
    wire n17456;
    wire n17462;
    wire n17465;
    wire n17468;
    wire n17471;
    wire n17474;
    wire n17477;
    wire n17480;
    wire n17483;
    wire n17486;
    wire n17489;
    wire n17492;
    wire n17495;
    wire n17498;
    wire n17501;
    wire n17504;
    wire n17507;
    wire n17510;
    wire n17513;
    wire n17516;
    wire n17519;
    wire n17522;
    wire n17525;
    wire n17528;
    wire n17531;
    wire n17537;
    wire n17540;
    wire n17543;
    wire n17546;
    wire n17549;
    wire n17552;
    wire n17555;
    wire n17558;
    wire n17561;
    wire n17564;
    wire n17567;
    wire n17570;
    wire n17573;
    wire n17576;
    wire n17579;
    wire n17582;
    wire n17585;
    wire n17588;
    wire n17591;
    wire n17594;
    wire n17597;
    wire n17600;
    wire n17603;
    wire n17606;
    wire n17612;
    wire n17615;
    wire n17618;
    wire n17621;
    wire n17624;
    wire n17627;
    wire n17630;
    wire n17633;
    wire n17636;
    wire n17639;
    wire n17642;
    wire n17645;
    wire n17648;
    wire n17651;
    wire n17654;
    wire n17657;
    wire n17660;
    wire n17663;
    wire n17666;
    wire n17669;
    wire n17672;
    wire n17675;
    wire n17678;
    wire n17681;
    wire n17687;
    wire n17690;
    wire n17693;
    wire n17696;
    wire n17699;
    wire n17702;
    wire n17705;
    wire n17708;
    wire n17711;
    wire n17714;
    wire n17717;
    wire n17720;
    wire n17723;
    wire n17726;
    wire n17729;
    wire n17732;
    wire n17735;
    wire n17738;
    wire n17741;
    wire n17744;
    wire n17747;
    wire n17750;
    wire n17753;
    wire n17756;
    wire n17762;
    wire n17765;
    wire n17768;
    wire n17771;
    wire n17774;
    wire n17777;
    wire n17780;
    wire n17783;
    wire n17786;
    wire n17789;
    wire n17792;
    wire n17795;
    wire n17798;
    wire n17801;
    wire n17804;
    wire n17807;
    wire n17810;
    wire n17813;
    wire n17816;
    wire n17819;
    wire n17822;
    wire n17825;
    wire n17828;
    wire n17831;
    wire n17837;
    wire n17840;
    wire n17843;
    wire n17846;
    wire n17849;
    wire n17852;
    wire n17855;
    wire n17858;
    wire n17861;
    wire n17864;
    wire n17867;
    wire n17870;
    wire n17873;
    wire n17876;
    wire n17879;
    wire n17882;
    wire n17885;
    wire n17888;
    wire n17891;
    wire n17894;
    wire n17897;
    wire n17900;
    wire n17903;
    wire n17906;
    wire n17912;
    wire n17915;
    wire n17918;
    wire n17921;
    wire n17924;
    wire n17927;
    wire n17930;
    wire n17933;
    wire n17936;
    wire n17939;
    wire n17942;
    wire n17945;
    wire n17948;
    wire n17951;
    wire n17954;
    wire n17957;
    wire n17960;
    wire n17963;
    wire n17966;
    wire n17969;
    wire n17972;
    wire n17975;
    wire n17978;
    wire n17981;
    wire n17987;
    wire n17990;
    wire n17993;
    wire n17996;
    wire n17999;
    wire n18002;
    wire n18005;
    wire n18008;
    wire n18011;
    wire n18014;
    wire n18017;
    wire n18020;
    wire n18023;
    wire n18026;
    wire n18029;
    wire n18032;
    wire n18035;
    wire n18038;
    wire n18041;
    wire n18044;
    wire n18047;
    wire n18050;
    wire n18053;
    wire n18056;
    wire n18062;
    wire n18065;
    wire n18068;
    wire n18071;
    wire n18074;
    wire n18077;
    wire n18080;
    wire n18083;
    wire n18086;
    wire n18089;
    wire n18092;
    wire n18095;
    wire n18098;
    wire n18101;
    wire n18104;
    wire n18107;
    wire n18110;
    wire n18113;
    wire n18116;
    wire n18119;
    wire n18122;
    wire n18125;
    wire n18128;
    wire n18134;
    wire n18137;
    wire n18140;
    wire n18143;
    wire n18146;
    wire n18149;
    wire n18152;
    wire n18155;
    wire n18158;
    wire n18161;
    wire n18164;
    wire n18167;
    wire n18170;
    wire n18173;
    wire n18176;
    wire n18179;
    wire n18182;
    wire n18185;
    wire n18188;
    wire n18191;
    wire n18194;
    wire n18197;
    wire n18200;
    wire n18206;
    wire n18209;
    wire n18212;
    wire n18215;
    wire n18218;
    wire n18221;
    wire n18224;
    wire n18227;
    wire n18230;
    wire n18233;
    wire n18236;
    wire n18239;
    wire n18242;
    wire n18245;
    wire n18248;
    wire n18251;
    wire n18254;
    wire n18257;
    wire n18260;
    wire n18263;
    wire n18266;
    wire n18269;
    wire n18272;
    wire n18278;
    wire n18281;
    wire n18284;
    wire n18287;
    wire n18290;
    wire n18293;
    wire n18296;
    wire n18299;
    wire n18302;
    wire n18305;
    wire n18308;
    wire n18311;
    wire n18314;
    wire n18317;
    wire n18320;
    wire n18323;
    wire n18326;
    wire n18329;
    wire n18332;
    wire n18335;
    wire n18338;
    wire n18341;
    wire n18344;
    wire n18347;
    wire n18353;
    wire n18356;
    wire n18359;
    wire n18362;
    wire n18365;
    wire n18368;
    wire n18371;
    wire n18374;
    wire n18377;
    wire n18380;
    wire n18383;
    wire n18386;
    wire n18389;
    wire n18392;
    wire n18395;
    wire n18398;
    wire n18401;
    wire n18404;
    wire n18407;
    wire n18410;
    wire n18413;
    wire n18416;
    wire n18419;
    wire n18422;
    wire n18428;
    wire n18431;
    wire n18434;
    wire n18437;
    wire n18440;
    wire n18443;
    wire n18446;
    wire n18449;
    wire n18452;
    wire n18455;
    wire n18458;
    wire n18461;
    wire n18464;
    wire n18467;
    wire n18470;
    wire n18473;
    wire n18476;
    wire n18479;
    wire n18482;
    wire n18485;
    wire n18488;
    wire n18491;
    wire n18494;
    wire n18497;
    wire n18503;
    wire n18506;
    wire n18509;
    wire n18512;
    wire n18515;
    wire n18518;
    wire n18521;
    wire n18524;
    wire n18527;
    wire n18530;
    wire n18533;
    wire n18536;
    wire n18539;
    wire n18542;
    wire n18545;
    wire n18548;
    wire n18551;
    wire n18554;
    wire n18557;
    wire n18560;
    wire n18563;
    wire n18566;
    wire n18569;
    wire n18572;
    wire n18578;
    wire n18581;
    wire n18584;
    wire n18587;
    wire n18590;
    wire n18593;
    wire n18596;
    wire n18599;
    wire n18602;
    wire n18605;
    wire n18608;
    wire n18611;
    wire n18614;
    wire n18617;
    wire n18620;
    wire n18623;
    wire n18626;
    wire n18629;
    wire n18632;
    wire n18635;
    wire n18638;
    wire n18641;
    wire n18644;
    wire n18647;
    wire n18653;
    wire n18656;
    wire n18659;
    wire n18662;
    wire n18665;
    wire n18668;
    wire n18671;
    wire n18674;
    wire n18677;
    wire n18680;
    wire n18683;
    wire n18686;
    wire n18689;
    wire n18692;
    wire n18695;
    wire n18698;
    wire n18701;
    wire n18704;
    wire n18707;
    wire n18710;
    wire n18713;
    wire n18716;
    wire n18719;
    wire n18722;
    wire n18728;
    wire n18731;
    wire n18734;
    wire n18737;
    wire n18740;
    wire n18743;
    wire n18746;
    wire n18749;
    wire n18752;
    wire n18755;
    wire n18758;
    wire n18761;
    wire n18764;
    wire n18767;
    wire n18770;
    wire n18773;
    wire n18776;
    wire n18779;
    wire n18782;
    wire n18785;
    wire n18788;
    wire n18791;
    wire n18797;
    wire n18800;
    wire n18803;
    wire n18806;
    wire n18809;
    wire n18812;
    wire n18815;
    wire n18818;
    wire n18821;
    wire n18824;
    wire n18827;
    wire n18830;
    wire n18833;
    wire n18836;
    wire n18839;
    wire n18842;
    wire n18845;
    wire n18848;
    wire n18851;
    wire n18854;
    wire n18857;
    wire n18860;
    wire n18863;
    wire n18869;
    wire n18872;
    wire n18875;
    wire n18878;
    wire n18881;
    wire n18884;
    wire n18887;
    wire n18890;
    wire n18893;
    wire n18896;
    wire n18899;
    wire n18902;
    wire n18905;
    wire n18908;
    wire n18911;
    wire n18914;
    wire n18917;
    wire n18920;
    wire n18923;
    wire n18926;
    wire n18929;
    wire n18932;
    wire n18935;
    wire n18938;
    wire n18944;
    wire n18947;
    wire n18950;
    wire n18953;
    wire n18956;
    wire n18959;
    wire n18962;
    wire n18965;
    wire n18968;
    wire n18971;
    wire n18974;
    wire n18977;
    wire n18980;
    wire n18983;
    wire n18986;
    wire n18989;
    wire n18992;
    wire n18995;
    wire n18998;
    wire n19001;
    wire n19004;
    wire n19007;
    wire n19010;
    wire n19013;
    wire n19019;
    wire n19022;
    wire n19025;
    wire n19028;
    wire n19031;
    wire n19034;
    wire n19037;
    wire n19040;
    wire n19043;
    wire n19046;
    wire n19049;
    wire n19052;
    wire n19055;
    wire n19058;
    wire n19061;
    wire n19064;
    wire n19067;
    wire n19070;
    wire n19073;
    wire n19076;
    wire n19079;
    wire n19082;
    wire n19085;
    wire n19088;
    wire n19094;
    wire n19097;
    wire n19100;
    wire n19103;
    wire n19106;
    wire n19109;
    wire n19112;
    wire n19115;
    wire n19118;
    wire n19121;
    wire n19124;
    wire n19127;
    wire n19130;
    wire n19133;
    wire n19136;
    wire n19139;
    wire n19142;
    wire n19145;
    wire n19148;
    wire n19151;
    wire n19154;
    wire n19157;
    wire n19160;
    wire n19163;
    wire n19169;
    wire n19172;
    wire n19175;
    wire n19178;
    wire n19181;
    wire n19184;
    wire n19187;
    wire n19190;
    wire n19193;
    wire n19196;
    wire n19199;
    wire n19202;
    wire n19205;
    wire n19208;
    wire n19211;
    wire n19214;
    wire n19217;
    wire n19220;
    wire n19223;
    wire n19226;
    wire n19229;
    wire n19232;
    wire n19235;
    wire n19238;
    wire n19244;
    wire n19247;
    wire n19250;
    wire n19253;
    wire n19256;
    wire n19259;
    wire n19262;
    wire n19265;
    wire n19268;
    wire n19271;
    wire n19274;
    wire n19277;
    wire n19280;
    wire n19283;
    wire n19286;
    wire n19289;
    wire n19292;
    wire n19295;
    wire n19298;
    wire n19301;
    wire n19304;
    wire n19307;
    wire n19310;
    wire n19313;
    wire n19319;
    wire n19322;
    wire n19325;
    wire n19328;
    wire n19331;
    wire n19334;
    wire n19337;
    wire n19340;
    wire n19343;
    wire n19346;
    wire n19349;
    wire n19352;
    wire n19355;
    wire n19358;
    wire n19361;
    wire n19364;
    wire n19367;
    wire n19370;
    wire n19373;
    wire n19376;
    wire n19379;
    wire n19385;
    wire n19388;
    wire n19391;
    wire n19394;
    wire n19397;
    wire n19400;
    wire n19403;
    wire n19406;
    wire n19409;
    wire n19412;
    wire n19415;
    wire n19418;
    wire n19421;
    wire n19424;
    wire n19427;
    wire n19430;
    wire n19433;
    wire n19436;
    wire n19439;
    wire n19442;
    wire n19445;
    wire n19451;
    wire n19454;
    wire n19457;
    wire n19460;
    wire n19463;
    wire n19466;
    wire n19469;
    wire n19472;
    wire n19475;
    wire n19478;
    wire n19481;
    wire n19484;
    wire n19487;
    wire n19490;
    wire n19493;
    wire n19496;
    wire n19499;
    wire n19502;
    wire n19505;
    wire n19508;
    wire n19511;
    wire n19517;
    wire n19520;
    wire n19523;
    wire n19526;
    wire n19529;
    wire n19532;
    wire n19535;
    wire n19538;
    wire n19541;
    wire n19544;
    wire n19547;
    wire n19550;
    wire n19553;
    wire n19556;
    wire n19559;
    wire n19562;
    wire n19565;
    wire n19568;
    wire n19571;
    wire n19574;
    wire n19577;
    wire n19580;
    wire n19586;
    wire n19589;
    wire n19592;
    wire n19595;
    wire n19598;
    wire n19601;
    wire n19604;
    wire n19607;
    wire n19610;
    wire n19613;
    wire n19616;
    wire n19619;
    wire n19622;
    wire n19625;
    wire n19628;
    wire n19631;
    wire n19634;
    wire n19637;
    wire n19640;
    wire n19643;
    wire n19649;
    wire n19652;
    wire n19655;
    wire n19658;
    wire n19661;
    wire n19664;
    wire n19667;
    wire n19670;
    wire n19673;
    wire n19676;
    wire n19679;
    wire n19682;
    wire n19685;
    wire n19688;
    wire n19691;
    wire n19694;
    wire n19697;
    wire n19700;
    wire n19703;
    wire n19706;
    wire n19712;
    wire n19715;
    wire n19718;
    wire n19721;
    wire n19724;
    wire n19727;
    wire n19730;
    wire n19733;
    wire n19736;
    wire n19739;
    wire n19742;
    wire n19745;
    wire n19748;
    wire n19751;
    wire n19754;
    wire n19757;
    wire n19760;
    wire n19763;
    wire n19766;
    wire n19769;
    wire n19775;
    wire n19778;
    wire n19781;
    wire n19784;
    wire n19787;
    wire n19790;
    wire n19793;
    wire n19796;
    wire n19799;
    wire n19802;
    wire n19805;
    wire n19808;
    wire n19811;
    wire n19814;
    wire n19817;
    wire n19820;
    wire n19823;
    wire n19826;
    wire n19829;
    wire n19832;
    wire n19838;
    wire n19841;
    wire n19844;
    wire n19847;
    wire n19850;
    wire n19853;
    wire n19856;
    wire n19859;
    wire n19862;
    wire n19865;
    wire n19868;
    wire n19871;
    wire n19874;
    wire n19877;
    wire n19880;
    wire n19883;
    wire n19889;
    wire n19892;
    wire n19895;
    wire n19898;
    wire n19901;
    wire n19904;
    wire n19907;
    wire n19910;
    wire n19913;
    wire n19916;
    wire n19919;
    wire n19922;
    wire n19925;
    wire n19928;
    wire n19931;
    wire n19934;
    wire n19940;
    wire n19943;
    wire n19946;
    wire n19949;
    wire n19952;
    wire n19955;
    wire n19958;
    wire n19961;
    wire n19964;
    wire n19967;
    wire n19970;
    wire n19973;
    wire n19976;
    wire n19979;
    wire n19985;
    wire n19988;
    wire n19991;
    wire n19994;
    wire n19997;
    wire n20000;
    wire n20003;
    wire n20006;
    wire n20009;
    wire n20012;
    wire n20015;
    wire n20018;
    wire n20021;
    wire n20024;
    wire n20027;
    wire n20030;
    wire n20036;
    wire n20039;
    wire n20042;
    wire n20045;
    wire n20048;
    wire n20051;
    wire n20054;
    wire n20057;
    wire n20060;
    wire n20063;
    wire n20066;
    wire n20069;
    wire n20072;
    wire n20075;
    wire n20078;
    wire n20081;
    wire n20087;
    wire n20090;
    wire n20093;
    wire n20096;
    wire n20099;
    wire n20102;
    wire n20105;
    wire n20108;
    wire n20111;
    wire n20114;
    wire n20117;
    wire n20120;
    wire n20123;
    wire n20126;
    wire n20132;
    wire n20135;
    wire n20138;
    wire n20141;
    wire n20144;
    wire n20147;
    wire n20150;
    wire n20153;
    wire n20156;
    wire n20159;
    wire n20162;
    wire n20165;
    wire n20168;
    wire n20171;
    wire n20174;
    wire n20177;
    wire n20180;
    wire n20183;
    wire n20186;
    wire n20189;
    wire n20195;
    wire n20198;
    wire n20201;
    wire n20204;
    wire n20207;
    wire n20210;
    wire n20213;
    wire n20216;
    wire n20219;
    wire n20222;
    wire n20225;
    wire n20228;
    wire n20231;
    wire n20234;
    wire n20237;
    wire n20240;
    wire n20243;
    wire n20246;
    wire n20249;
    wire n20252;
    wire n20258;
    wire n20261;
    wire n20264;
    wire n20267;
    wire n20270;
    wire n20273;
    wire n20276;
    wire n20279;
    wire n20282;
    wire n20285;
    wire n20288;
    wire n20294;
    wire n20297;
    wire n20300;
    wire n20303;
    wire n20306;
    wire n20309;
    wire n20312;
    wire n20315;
    wire n20318;
    wire n20321;
    wire n20324;
    wire n20330;
    wire n20333;
    wire n20336;
    wire n20339;
    wire n20342;
    wire n20345;
    wire n20348;
    wire n20351;
    wire n20354;
    wire n20357;
    wire n20360;
    wire n20366;
    wire n20369;
    wire n20372;
    wire n20375;
    wire n20378;
    wire n20381;
    wire n20384;
    wire n20387;
    wire n20390;
    wire n20393;
    wire n20396;
    wire n20402;
    wire n20405;
    wire n20408;
    wire n20411;
    wire n20414;
    wire n20417;
    wire n20420;
    wire n20423;
    wire n20426;
    wire n20429;
    wire n20432;
    wire n20435;
    wire n20438;
    wire n20441;
    wire n20444;
    wire n20447;
    wire n20450;
    wire n20453;
    wire n20459;
    wire n20462;
    wire n20465;
    wire n20468;
    wire n20471;
    wire n20474;
    wire n20477;
    wire n20480;
    wire n20483;
    wire n20486;
    wire n20489;
    wire n20492;
    wire n20495;
    wire n20498;
    wire n20501;
    wire n20504;
    wire n20507;
    wire n20513;
    wire n20516;
    wire n20519;
    wire n20522;
    wire n20525;
    wire n20528;
    wire n20531;
    wire n20534;
    wire n20537;
    wire n20540;
    wire n20543;
    wire n20546;
    wire n20549;
    wire n20552;
    wire n20555;
    wire n20558;
    wire n20561;
    wire n20567;
    wire n20570;
    wire n20573;
    wire n20576;
    wire n20579;
    wire n20582;
    wire n20588;
    wire n20591;
    wire n20594;
    wire n20597;
    wire n20600;
    wire n20603;
    wire n20606;
    wire n20609;
    wire n20612;
    wire n20615;
    wire n20618;
    wire n20621;
    wire n20624;
    wire n20627;
    wire n20633;
    wire n20636;
    wire n20639;
    wire n20642;
    wire n20645;
    wire n20648;
    wire n20651;
    wire n20654;
    wire n20657;
    wire n20660;
    wire n20663;
    wire n20669;
    wire n20672;
    wire n20675;
    wire n20678;
    wire n20681;
    wire n20684;
    wire n20687;
    wire n20690;
    wire n20693;
    wire n20696;
    wire n20699;
    wire n20702;
    wire n20705;
    wire n20711;
    wire n20714;
    wire n20717;
    wire n20720;
    wire n20723;
    wire n20726;
    wire n20729;
    wire n20732;
    wire n20735;
    wire n20738;
    wire n20741;
    wire n20744;
    wire n20747;
    wire n20750;
    wire n20753;
    wire n20759;
    wire n20762;
    wire n20765;
    wire n20768;
    wire n20771;
    wire n20774;
    wire n20777;
    wire n20780;
    wire n20783;
    wire n20786;
    wire n20789;
    wire n20792;
    wire n20795;
    wire n20798;
    wire n20804;
    wire n20807;
    wire n20810;
    wire n20813;
    wire n20816;
    wire n20819;
    wire n20822;
    wire n20825;
    wire n20828;
    wire n20834;
    wire n20837;
    wire n20840;
    wire n20843;
    wire n20846;
    wire n20849;
    wire n20852;
    wire n20855;
    wire n20858;
    wire n20861;
    wire n20864;
    wire n20870;
    wire n20873;
    wire n20876;
    wire n20879;
    wire n20882;
    wire n20885;
    wire n20888;
    wire n20891;
    wire n20894;
    wire n20897;
    wire n20900;
    wire n20903;
    wire n20909;
    wire n20912;
    wire n20915;
    wire n20918;
    wire n20921;
    wire n20924;
    wire n20927;
    wire n20930;
    wire n20933;
    wire n20936;
    wire n20939;
    wire n20942;
    wire n20945;
    wire n20951;
    wire n20954;
    wire n20957;
    wire n20960;
    wire n20963;
    wire n20966;
    wire n20969;
    wire n20972;
    wire n20975;
    wire n20978;
    wire n20981;
    wire n20984;
    wire n20987;
    wire n20990;
    wire n20993;
    wire n20996;
    wire n21002;
    wire n21005;
    wire n21008;
    wire n21011;
    wire n21014;
    wire n21017;
    wire n21020;
    wire n21023;
    wire n21026;
    wire n21029;
    wire n21032;
    wire n21035;
    wire n21038;
    wire n21041;
    wire n21044;
    wire n21047;
    wire n21050;
    wire n21053;
    wire n21059;
    wire n21062;
    wire n21065;
    wire n21068;
    wire n21074;
    wire n21077;
    wire n21080;
    wire n21083;
    wire n21086;
    wire n21089;
    wire n21092;
    wire n21098;
    wire n21101;
    wire n21104;
    wire n21107;
    wire n21110;
    wire n21113;
    wire n21116;
    wire n21119;
    wire n21122;
    wire n21125;
    wire n21128;
    wire n21131;
    wire n21134;
    wire n21140;
    wire n21143;
    wire n21146;
    wire n21149;
    wire n21152;
    wire n21155;
    wire n21158;
    wire n21161;
    wire n21164;
    wire n21167;
    wire n21170;
    wire n21173;
    wire n21176;
    wire n21182;
    wire n21185;
    wire n21188;
    wire n21191;
    wire n21194;
    wire n21197;
    wire n21203;
    wire n21206;
    wire n21209;
    wire n21212;
    wire n21215;
    wire n21218;
    wire n21221;
    wire n21224;
    wire n21230;
    wire n21233;
    wire n21236;
    wire n21239;
    wire n21242;
    wire n21245;
    wire n21248;
    wire n21251;
    wire n21254;
    wire n21260;
    wire n21263;
    wire n21266;
    wire n21269;
    wire n21272;
    wire n21275;
    wire n21278;
    wire n21281;
    wire n21284;
    wire n21287;
    wire n21293;
    wire n21296;
    wire n21299;
    wire n21302;
    wire n21305;
    wire n21308;
    wire n21314;
    wire n21317;
    wire n21320;
    wire n21323;
    wire n21326;
    wire n21329;
    wire n21332;
    wire n21335;
    wire n21341;
    wire n21344;
    wire n21347;
    wire n21350;
    wire n21353;
    wire n21356;
    wire n21359;
    wire n21362;
    wire n21365;
    wire n21371;
    wire n21374;
    wire n21377;
    wire n21380;
    wire n21383;
    wire n21386;
    wire n21389;
    wire n21392;
    wire n21395;
    wire n21398;
    wire n21404;
    wire n21407;
    wire n21410;
    wire n21413;
    wire n21416;
    wire n21422;
    wire n21425;
    wire n21428;
    wire n21431;
    wire n21434;
    wire n21437;
    wire n21440;
    wire n21443;
    wire n21446;
    wire n21452;
    wire n21455;
    wire n21458;
    wire n21461;
    wire n21464;
    wire n21467;
    wire n21470;
    wire n21473;
    wire n21479;
    wire n21482;
    wire n21485;
    wire n21488;
    wire n21491;
    wire n21494;
    wire n21497;
    wire n21503;
    wire n21506;
    wire n21509;
    wire n21512;
    wire n21515;
    wire n21521;
    wire n21524;
    wire n21527;
    wire n21530;
    wire n21533;
    wire n21536;
    wire n21539;
    wire n21542;
    wire n21545;
    wire n21551;
    wire n21554;
    wire n21557;
    wire n21560;
    wire n21563;
    wire n21566;
    wire n21569;
    wire n21572;
    wire n21578;
    wire n21581;
    wire n21584;
    wire n21587;
    wire n21590;
    wire n21593;
    wire n21596;
    wire n21602;
    wire n21605;
    wire n21608;
    wire n21611;
    wire n21617;
    wire n21620;
    wire n21623;
    wire n21626;
    wire n21629;
    wire n21632;
    wire n21635;
    wire n21638;
    wire n21644;
    wire n21647;
    wire n21650;
    wire n21653;
    wire n21659;
    wire n21662;
    wire n21665;
    wire n21668;
    wire n21671;
    wire n21674;
    wire n21677;
    wire n21683;
    wire n21686;
    wire n21689;
    wire n21692;
    wire n21695;
    wire n21698;
    wire n21701;
    wire n21707;
    wire n21710;
    wire n21713;
    wire n21716;
    wire n21719;
    wire n21722;
    wire n21725;
    wire n21728;
    wire n21734;
    wire n21737;
    wire n21740;
    wire n21743;
    wire n21746;
    wire n21749;
    wire n21752;
    wire n21755;
    wire n21758;
    wire n21761;
    wire n21764;
    wire n21767;
    wire n21770;
    wire n21773;
    wire n21776;
    wire n21782;
    wire n21785;
    wire n21788;
    wire n21794;
    wire n21797;
    wire n21800;
    wire n21803;
    wire n21809;
    wire n21812;
    wire n21815;
    wire n21818;
    wire n21821;
    wire n21824;
    wire n21830;
    wire n21833;
    wire n21836;
    wire n21839;
    wire n21842;
    wire n21845;
    wire n21848;
    wire n21854;
    wire n21857;
    wire n21863;
    wire n21866;
    wire n21872;
    wire n21875;
    wire n21878;
    wire n21884;
    wire n21887;
    wire n21890;
    wire n21896;
    wire n21899;
    wire n21902;
    wire n21905;
    wire n21911;
    wire n21914;
    wire n21917;
    wire n21923;
    wire n21926;
    wire n21929;
    wire n21935;
    wire n21938;
    wire n21941;
    wire n21944;
    wire n21950;
    wire n21953;
    wire n21956;
    wire n21962;
    wire n21965;
    wire n21971;
    wire n21974;
    wire n21980;
    wire n21986;
    wire n21989;
    wire n21992;
    wire n21998;
    wire n22001;
    wire n22007;
    wire n22010;
    wire n22016;
    wire n22022;
    wire n22025;
    wire n22028;
    wire n22034;
    wire n22037;
    wire n22040;
    jnot g0000(.din(G545), .dout(n303));
    jnot g0001(.din(G348), .dout(n306));
    jnot g0002(.din(G366), .dout(n309));
    jand g0003(.dinb(G552), .dina(G562), .dout(n313));
    jnot g0004(.din(G549), .dout(n316));
    jdff g0005(.din(G338), .dout(n319));
    jnot g0006(.din(G358), .dout(n322));
    jand g0007(.dinb(G141), .dina(G145), .dout(n326));
    jnot g0008(.din(G245), .dout(n329));
    jnot g0009(.din(G552), .dout(n332));
    jnot g0010(.din(G562), .dout(n335));
    jnot g0011(.din(G559), .dout(n338));
    jor g0012(.dinb(G1), .dina(G373), .dout(n342));
    jnot g0013(.din(G3173), .dout(n345));
    jand g0014(.dinb(n8016), .dina(n345), .dout(n349));
    jnot g0015(.din(G27), .dout(n352));
    jor g0016(.dinb(n352), .dina(n8019), .dout(n356));
    jand g0017(.dinb(G386), .dina(G556), .dout(n360));
    jnot g0018(.din(n360), .dout(n363));
    jnot g0019(.din(G140), .dout(n366));
    jnot g0020(.din(G31), .dout(n369));
    jor g0021(.dinb(n352), .dina(n369), .dout(n373));
    jor g0022(.dinb(n8022), .dina(n373), .dout(n377));
    jnot g0023(.din(G299), .dout(n380));
    jnot g0024(.din(G86), .dout(n383));
    jnot g0025(.din(G2358), .dout(n386));
    jand g0026(.dinb(n383), .dina(n386), .dout(n390));
    jnot g0027(.din(G87), .dout(n393));
    jand g0028(.dinb(n393), .dina(n8096), .dout(n397));
    jor g0029(.dinb(n373), .dina(n397), .dout(n401));
    jor g0030(.dinb(n8025), .dina(n401), .dout(n405));
    jnot g0031(.din(G88), .dout(n408));
    jand g0032(.dinb(n408), .dina(n386), .dout(n412));
    jnot g0033(.din(G34), .dout(n415));
    jand g0034(.dinb(n415), .dina(n8093), .dout(n419));
    jor g0035(.dinb(n373), .dina(n419), .dout(n423));
    jor g0036(.dinb(n8028), .dina(n423), .dout(n427));
    jnot g0037(.din(G83), .dout(n430));
    jor g0038(.dinb(n8031), .dina(n373), .dout(n434));
    jand g0039(.dinb(n8040), .dina(n386), .dout(n438));
    jand g0040(.dinb(G25), .dina(G2358), .dout(n442));
    jor g0041(.dinb(n373), .dina(n8037), .dout(n446));
    jor g0042(.dinb(n8034), .dina(n446), .dout(n450));
    jand g0043(.dinb(n8063), .dina(n450), .dout(n454));
    jand g0044(.dinb(n8049), .dina(n386), .dout(n458));
    jand g0045(.dinb(G81), .dina(G2358), .dout(n462));
    jor g0046(.dinb(n373), .dina(n8046), .dout(n466));
    jor g0047(.dinb(n8043), .dina(n466), .dout(n470));
    jand g0048(.dinb(n8051), .dina(n470), .dout(n474));
    jand g0049(.dinb(n8082), .dina(n386), .dout(n478));
    jand g0050(.dinb(G23), .dina(G2358), .dout(n482));
    jor g0051(.dinb(n373), .dina(n8079), .dout(n486));
    jor g0052(.dinb(n8076), .dina(n486), .dout(n490));
    jand g0053(.dinb(n8111), .dina(n490), .dout(n494));
    jand g0054(.dinb(n8091), .dina(n386), .dout(n498));
    jand g0055(.dinb(G80), .dina(G2358), .dout(n502));
    jor g0056(.dinb(n373), .dina(n8088), .dout(n506));
    jor g0057(.dinb(n8085), .dina(n506), .dout(n510));
    jand g0058(.dinb(n8099), .dina(n510), .dout(n514));
    jnot g0059(.din(G308), .dout(n517));
    jand g0060(.dinb(n16142), .dina(n517), .dout(n521));
    jnot g0061(.din(G479), .dout(n524));
    jand g0062(.dinb(G248), .dina(G308), .dout(n528));
    jor g0063(.dinb(n524), .dina(n528), .dout(n532));
    jor g0064(.dinb(n521), .dina(n532), .dout(n536));
    jnot g0065(.din(G254), .dout(n539));
    jand g0066(.dinb(n539), .dina(n517), .dout(n543));
    jnot g0067(.din(G242), .dout(n546));
    jand g0068(.dinb(n546), .dina(n14621), .dout(n550));
    jor g0069(.dinb(n14597), .dina(n550), .dout(n554));
    jor g0070(.dinb(n14586), .dina(n554), .dout(n558));
    jand g0071(.dinb(n14583), .dina(n558), .dout(n562));
    jnot g0072(.din(G316), .dout(n565));
    jand g0073(.dinb(n16139), .dina(n565), .dout(n569));
    jnot g0074(.din(G490), .dout(n572));
    jand g0075(.dinb(G248), .dina(G316), .dout(n576));
    jor g0076(.dinb(n572), .dina(n576), .dout(n580));
    jor g0077(.dinb(n569), .dina(n580), .dout(n584));
    jand g0078(.dinb(n539), .dina(n565), .dout(n588));
    jand g0079(.dinb(n546), .dina(n14579), .dout(n592));
    jor g0080(.dinb(n14555), .dina(n592), .dout(n596));
    jor g0081(.dinb(n14544), .dina(n596), .dout(n600));
    jand g0082(.dinb(n14541), .dina(n600), .dout(n604));
    jand g0083(.dinb(n562), .dina(n604), .dout(n608));
    jnot g0084(.din(G351), .dout(n611));
    jnot g0085(.din(G3550), .dout(n614));
    jand g0086(.dinb(n611), .dina(n614), .dout(n618));
    jnot g0087(.din(G534), .dout(n621));
    jnot g0088(.din(G3552), .dout(n624));
    jand g0089(.dinb(n14495), .dina(n624), .dout(n628));
    jor g0090(.dinb(n14478), .dina(n628), .dout(n632));
    jor g0091(.dinb(n9321), .dina(n632), .dout(n636));
    jand g0092(.dinb(n611), .dina(n11436), .dout(n640));
    jand g0093(.dinb(G351), .dina(G3546), .dout(n644));
    jor g0094(.dinb(n14489), .dina(n644), .dout(n648));
    jor g0095(.dinb(n640), .dina(n648), .dout(n652));
    jand g0096(.dinb(n636), .dina(n9318), .dout(n656));
    jnot g0097(.din(G293), .dout(n659));
    jand g0098(.dinb(n539), .dina(n659), .dout(n663));
    jand g0099(.dinb(n546), .dina(n14636), .dout(n667));
    jor g0100(.dinb(n663), .dina(n667), .dout(n671));
    jnot g0101(.din(G251), .dout(n674));
    jnot g0102(.din(G302), .dout(n677));
    jand g0103(.dinb(n674), .dina(n677), .dout(n681));
    jnot g0104(.din(G248), .dout(n684));
    jand g0105(.dinb(n684), .dina(n14627), .dout(n688));
    jor g0106(.dinb(n681), .dina(n688), .dout(n692));
    jnot g0107(.din(n692), .dout(n695));
    jand g0108(.dinb(n14633), .dina(n695), .dout(n699));
    jnot g0109(.din(G514), .dout(n702));
    jnot g0110(.din(G3546), .dout(n705));
    jand g0111(.dinb(n702), .dina(n705), .dout(n709));
    jand g0112(.dinb(G514), .dina(G3552), .dout(n713));
    jor g0113(.dinb(n709), .dina(n9609), .dout(n717));
    jnot g0114(.din(n717), .dout(n720));
    jnot g0115(.din(G361), .dout(n723));
    jand g0116(.dinb(n674), .dina(n723), .dout(n727));
    jand g0117(.dinb(n684), .dina(n14528), .dout(n731));
    jor g0118(.dinb(n727), .dina(n731), .dout(n735));
    jnot g0119(.din(n735), .dout(n738));
    jand g0120(.dinb(n720), .dina(n738), .dout(n742));
    jand g0121(.dinb(n699), .dina(n742), .dout(n746));
    jand g0122(.dinb(n9314), .dina(n746), .dout(n750));
    jnot g0123(.din(G324), .dout(n753));
    jand g0124(.dinb(n753), .dina(n614), .dout(n757));
    jnot g0125(.din(G503), .dout(n760));
    jand g0126(.dinb(n14462), .dina(n624), .dout(n764));
    jor g0127(.dinb(n14426), .dina(n764), .dout(n768));
    jor g0128(.dinb(n9177), .dina(n768), .dout(n772));
    jand g0129(.dinb(n753), .dina(n11436), .dout(n776));
    jand g0130(.dinb(G324), .dina(G3546), .dout(n780));
    jor g0131(.dinb(n14441), .dina(n780), .dout(n784));
    jor g0132(.dinb(n776), .dina(n784), .dout(n788));
    jand g0133(.dinb(n772), .dina(n9174), .dout(n792));
    jnot g0134(.din(G341), .dout(n795));
    jand g0135(.dinb(n795), .dina(n614), .dout(n799));
    jnot g0136(.din(G523), .dout(n802));
    jand g0137(.dinb(n14672), .dina(n624), .dout(n806));
    jor g0138(.dinb(n14645), .dina(n806), .dout(n810));
    jor g0139(.dinb(n9465), .dina(n810), .dout(n814));
    jand g0140(.dinb(n795), .dina(n11436), .dout(n818));
    jand g0141(.dinb(G341), .dina(G3546), .dout(n822));
    jor g0142(.dinb(n14654), .dina(n822), .dout(n826));
    jor g0143(.dinb(n818), .dina(n826), .dout(n830));
    jand g0144(.dinb(n814), .dina(n9462), .dout(n834));
    jand g0145(.dinb(n792), .dina(n834), .dout(n838));
    jand g0146(.dinb(n750), .dina(n8130), .dout(n842));
    jand g0147(.dinb(n8127), .dina(n842), .dout(n846));
    jnot g0148(.din(G265), .dout(n849));
    jand g0149(.dinb(n849), .dina(n614), .dout(n853));
    jnot g0150(.din(G400), .dout(n856));
    jand g0151(.dinb(n15983), .dina(n624), .dout(n860));
    jor g0152(.dinb(n15956), .dina(n860), .dout(n864));
    jor g0153(.dinb(n9519), .dina(n864), .dout(n868));
    jand g0154(.dinb(n849), .dina(n11436), .dout(n872));
    jand g0155(.dinb(G265), .dina(G3546), .dout(n876));
    jor g0156(.dinb(n15965), .dina(n876), .dout(n880));
    jor g0157(.dinb(n872), .dina(n880), .dout(n884));
    jand g0158(.dinb(n868), .dina(n9516), .dout(n888));
    jnot g0159(.din(G234), .dout(n891));
    jand g0160(.dinb(n891), .dina(n614), .dout(n895));
    jnot g0161(.din(G435), .dout(n898));
    jand g0162(.dinb(n16280), .dina(n624), .dout(n902));
    jor g0163(.dinb(n16238), .dina(n902), .dout(n906));
    jor g0164(.dinb(n9243), .dina(n906), .dout(n910));
    jand g0165(.dinb(n891), .dina(n11436), .dout(n914));
    jand g0166(.dinb(G234), .dina(G3546), .dout(n918));
    jor g0167(.dinb(n16253), .dina(n918), .dout(n922));
    jor g0168(.dinb(n914), .dina(n922), .dout(n926));
    jand g0169(.dinb(n910), .dina(n9240), .dout(n930));
    jnot g0170(.din(G257), .dout(n933));
    jand g0171(.dinb(n933), .dina(n614), .dout(n937));
    jnot g0172(.din(G389), .dout(n940));
    jand g0173(.dinb(n15935), .dina(n624), .dout(n944));
    jor g0174(.dinb(n15930), .dina(n944), .dout(n948));
    jor g0175(.dinb(n9705), .dina(n948), .dout(n952));
    jand g0176(.dinb(n933), .dina(n11436), .dout(n956));
    jand g0177(.dinb(G257), .dina(G3546), .dout(n960));
    jor g0178(.dinb(n15944), .dina(n960), .dout(n964));
    jor g0179(.dinb(n956), .dina(n964), .dout(n968));
    jand g0180(.dinb(n952), .dina(n9702), .dout(n972));
    jand g0181(.dinb(n930), .dina(n972), .dout(n976));
    jand g0182(.dinb(n9512), .dina(n976), .dout(n980));
    jnot g0183(.din(G273), .dout(n983));
    jand g0184(.dinb(n983), .dina(n614), .dout(n987));
    jnot g0185(.din(G411), .dout(n990));
    jand g0186(.dinb(n15911), .dina(n624), .dout(n994));
    jor g0187(.dinb(n15893), .dina(n994), .dout(n998));
    jor g0188(.dinb(n9354), .dina(n998), .dout(n1002));
    jand g0189(.dinb(n983), .dina(n11436), .dout(n1006));
    jand g0190(.dinb(G273), .dina(G3546), .dout(n1010));
    jor g0191(.dinb(n15908), .dina(n1010), .dout(n1014));
    jor g0192(.dinb(n1006), .dina(n1014), .dout(n1018));
    jand g0193(.dinb(n1002), .dina(n9351), .dout(n1022));
    jnot g0194(.din(G281), .dout(n1025));
    jand g0195(.dinb(n1025), .dina(n614), .dout(n1029));
    jnot g0196(.din(G374), .dout(n1032));
    jand g0197(.dinb(n16013), .dina(n624), .dout(n1036));
    jor g0198(.dinb(n15995), .dina(n1036), .dout(n1040));
    jor g0199(.dinb(n8379), .dina(n1040), .dout(n1044));
    jand g0200(.dinb(n1025), .dina(n11436), .dout(n1048));
    jand g0201(.dinb(G281), .dina(G3546), .dout(n1052));
    jor g0202(.dinb(n16010), .dina(n1052), .dout(n1056));
    jor g0203(.dinb(n1048), .dina(n1056), .dout(n1060));
    jand g0204(.dinb(n1044), .dina(n8376), .dout(n1064));
    jand g0205(.dinb(n1022), .dina(n1064), .dout(n1068));
    jnot g0206(.din(G218), .dout(n1071));
    jand g0207(.dinb(n1071), .dina(n614), .dout(n1075));
    jnot g0208(.din(G468), .dout(n1078));
    jand g0209(.dinb(n16085), .dina(n624), .dout(n1082));
    jor g0210(.dinb(n16068), .dina(n1082), .dout(n1086));
    jor g0211(.dinb(n11046), .dina(n1086), .dout(n1090));
    jand g0212(.dinb(n1071), .dina(n11436), .dout(n1094));
    jand g0213(.dinb(G218), .dina(G3546), .dout(n1098));
    jor g0214(.dinb(n16079), .dina(n1098), .dout(n1102));
    jor g0215(.dinb(n1094), .dina(n1102), .dout(n1106));
    jand g0216(.dinb(n1090), .dina(n11043), .dout(n1110));
    jnot g0217(.din(G206), .dout(n1113));
    jand g0218(.dinb(n1113), .dina(n16277), .dout(n1117));
    jnot g0219(.din(G446), .dout(n1120));
    jand g0220(.dinb(G206), .dina(G248), .dout(n1124));
    jor g0221(.dinb(n1120), .dina(n1124), .dout(n1128));
    jor g0222(.dinb(n1117), .dina(n1128), .dout(n1132));
    jand g0223(.dinb(n1113), .dina(n539), .dout(n1136));
    jand g0224(.dinb(n16202), .dina(n546), .dout(n1140));
    jor g0225(.dinb(n16172), .dina(n1140), .dout(n1144));
    jor g0226(.dinb(n16158), .dina(n1144), .dout(n1148));
    jand g0227(.dinb(n16155), .dina(n1148), .dout(n1152));
    jand g0228(.dinb(n1110), .dina(n1152), .dout(n1156));
    jnot g0229(.din(G226), .dout(n1159));
    jand g0230(.dinb(n1159), .dina(n614), .dout(n1163));
    jnot g0231(.din(G422), .dout(n1166));
    jand g0232(.dinb(n16121), .dina(n624), .dout(n1170));
    jor g0233(.dinb(n16113), .dina(n1170), .dout(n1174));
    jor g0234(.dinb(n10860), .dina(n1174), .dout(n1178));
    jand g0235(.dinb(n1159), .dina(n11436), .dout(n1182));
    jand g0236(.dinb(G226), .dina(G3546), .dout(n1186));
    jor g0237(.dinb(n16115), .dina(n1186), .dout(n1190));
    jor g0238(.dinb(n1182), .dina(n1190), .dout(n1194));
    jand g0239(.dinb(n1178), .dina(n10857), .dout(n1198));
    jnot g0240(.din(G210), .dout(n1201));
    jand g0241(.dinb(n1201), .dina(n614), .dout(n1205));
    jnot g0242(.din(G457), .dout(n1208));
    jand g0243(.dinb(n16055), .dina(n624), .dout(n1212));
    jor g0244(.dinb(n16034), .dina(n1212), .dout(n1216));
    jor g0245(.dinb(n11439), .dina(n1216), .dout(n1220));
    jand g0246(.dinb(n1201), .dina(n11436), .dout(n1224));
    jand g0247(.dinb(G210), .dina(G3546), .dout(n1228));
    jor g0248(.dinb(n16037), .dina(n1228), .dout(n1232));
    jor g0249(.dinb(n1224), .dina(n1232), .dout(n1236));
    jand g0250(.dinb(n1220), .dina(n11433), .dout(n1240));
    jand g0251(.dinb(n1198), .dina(n1240), .dout(n1244));
    jand g0252(.dinb(n1156), .dina(n1244), .dout(n1248));
    jand g0253(.dinb(n8136), .dina(n1248), .dout(n1252));
    jand g0254(.dinb(n8133), .dina(n1252), .dout(n1256));
    jnot g0255(.din(G335), .dout(n1259));
    jor g0256(.dinb(n15609), .dina(n1259), .dout(n1263));
    jand g0257(.dinb(n891), .dina(n1259), .dout(n1267));
    jnot g0258(.din(n1267), .dout(n1270));
    jand g0259(.dinb(n15606), .dina(n1270), .dout(n1274));
    jxor g0260(.dinb(n16241), .dina(n1274), .dout(n1278));
    jnot g0261(.din(n1278), .dout(n1281));
    jnot g0262(.din(G288), .dout(n1284));
    jand g0263(.dinb(n1284), .dina(n15746), .dout(n1288));
    jand g0264(.dinb(n1025), .dina(n1259), .dout(n1292));
    jor g0265(.dinb(n1288), .dina(n1292), .dout(n1296));
    jxor g0266(.dinb(n15407), .dina(n1296), .dout(n1300));
    jor g0267(.dinb(n15569), .dina(n1259), .dout(n1304));
    jor g0268(.dinb(G273), .dina(G335), .dout(n1308));
    jand g0269(.dinb(n1304), .dina(n15566), .dout(n1312));
    jxor g0270(.dinb(n15572), .dina(n1312), .dout(n1316));
    jnot g0271(.din(n1316), .dout(n1319));
    jand g0272(.dinb(n15395), .dina(n1319), .dout(n1323));
    jnot g0273(.din(n1323), .dout(n1326));
    jor g0274(.dinb(n15684), .dina(n1259), .dout(n1330));
    jor g0275(.dinb(G257), .dina(G335), .dout(n1334));
    jand g0276(.dinb(n1330), .dina(n15678), .dout(n1338));
    jxor g0277(.dinb(n15692), .dina(n1338), .dout(n1342));
    jnot g0278(.din(G272), .dout(n1345));
    jand g0279(.dinb(n1345), .dina(n15680), .dout(n1349));
    jand g0280(.dinb(n849), .dina(n1259), .dout(n1353));
    jor g0281(.dinb(n1349), .dina(n1353), .dout(n1357));
    jxor g0282(.dinb(n15974), .dina(n1357), .dout(n1361));
    jor g0283(.dinb(n1342), .dina(n1361), .dout(n1365));
    jor g0284(.dinb(n1326), .dina(n15372), .dout(n1369));
    jor g0285(.dinb(n15429), .dina(n1369), .dout(n1373));
    jnot g0286(.din(n1373), .dout(n1376));
    jor g0287(.dinb(n15744), .dina(n1259), .dout(n1380));
    jor g0288(.dinb(G210), .dina(G335), .dout(n1384));
    jand g0289(.dinb(n1380), .dina(n15741), .dout(n1388));
    jxor g0290(.dinb(n16040), .dina(n1388), .dout(n1392));
    jor g0291(.dinb(n15360), .dina(n1259), .dout(n1396));
    jand g0292(.dinb(n1113), .dina(n1259), .dout(n1400));
    jnot g0293(.din(n1400), .dout(n1403));
    jand g0294(.dinb(n15357), .dina(n1403), .dout(n1407));
    jxor g0295(.dinb(n16160), .dina(n1407), .dout(n1411));
    jand g0296(.dinb(n15731), .dina(n1411), .dout(n1415));
    jor g0297(.dinb(n15291), .dina(n1259), .dout(n1419));
    jor g0298(.dinb(G226), .dina(G335), .dout(n1423));
    jand g0299(.dinb(n1419), .dina(n15288), .dout(n1427));
    jxor g0300(.dinb(n16124), .dina(n1427), .dout(n1431));
    jor g0301(.dinb(n15303), .dina(n1259), .dout(n1435));
    jor g0302(.dinb(G218), .dina(G335), .dout(n1439));
    jand g0303(.dinb(n1435), .dina(n15300), .dout(n1443));
    jxor g0304(.dinb(n16070), .dina(n1443), .dout(n1447));
    jand g0305(.dinb(n1431), .dina(n1447), .dout(n1451));
    jand g0306(.dinb(n1415), .dina(n8187), .dout(n1455));
    jand g0307(.dinb(n1376), .dina(n8184), .dout(n1459));
    jnot g0308(.din(G332), .dout(n1462));
    jor g0309(.dinb(n14294), .dina(n1462), .dout(n1466));
    jand g0310(.dinb(n753), .dina(n1462), .dout(n1470));
    jnot g0311(.din(n1470), .dout(n1473));
    jand g0312(.dinb(n14286), .dina(n1473), .dout(n1477));
    jxor g0313(.dinb(n14429), .dina(n1477), .dout(n1481));
    jor g0314(.dinb(n1462), .dina(n14213), .dout(n1485));
    jor g0315(.dinb(G332), .dina(G351), .dout(n1489));
    jand g0316(.dinb(n1485), .dina(n14085), .dout(n1493));
    jxor g0317(.dinb(n14219), .dina(n1493), .dout(n1497));
    jand g0318(.dinb(n14288), .dina(n309), .dout(n1501));
    jand g0319(.dinb(n1462), .dina(n723), .dout(n1505));
    jor g0320(.dinb(n1501), .dina(n1505), .dout(n1509));
    jnot g0321(.din(n1509), .dout(n1512));
    jor g0322(.dinb(n1497), .dina(n1512), .dout(n1516));
    jand g0323(.dinb(n14252), .dina(n319), .dout(n1520));
    jxor g0324(.dinb(n14522), .dina(n1520), .dout(n1524));
    jor g0325(.dinb(n1462), .dina(n14237), .dout(n1528));
    jor g0326(.dinb(G332), .dina(G341), .dout(n1532));
    jand g0327(.dinb(n1528), .dina(n14073), .dout(n1536));
    jxor g0328(.dinb(n14246), .dina(n1536), .dout(n1540));
    jor g0329(.dinb(n14078), .dina(n1540), .dout(n1544));
    jor g0330(.dinb(n1516), .dina(n1544), .dout(n1548));
    jnot g0331(.din(n1548), .dout(n1551));
    jand g0332(.dinb(n14267), .dina(n1551), .dout(n1555));
    jand g0333(.dinb(n380), .dina(n14249), .dout(n1559));
    jand g0334(.dinb(n659), .dina(n1462), .dout(n1563));
    jor g0335(.dinb(n1559), .dina(n1563), .dout(n1567));
    jor g0336(.dinb(n14040), .dina(n1462), .dout(n1571));
    jand g0337(.dinb(n677), .dina(n1462), .dout(n1575));
    jnot g0338(.din(n1575), .dout(n1578));
    jand g0339(.dinb(n14037), .dina(n1578), .dout(n1582));
    jnot g0340(.din(n1582), .dout(n1585));
    jand g0341(.dinb(n13733), .dina(n1585), .dout(n1589));
    jor g0342(.dinb(n13998), .dina(n1462), .dout(n1593));
    jor g0343(.dinb(G308), .dina(G332), .dout(n1597));
    jand g0344(.dinb(n1593), .dina(n13995), .dout(n1601));
    jxor g0345(.dinb(n14612), .dina(n1601), .dout(n1605));
    jor g0346(.dinb(n13953), .dina(n1462), .dout(n1609));
    jor g0347(.dinb(G316), .dina(G332), .dout(n1613));
    jand g0348(.dinb(n1609), .dina(n13950), .dout(n1617));
    jxor g0349(.dinb(n14546), .dina(n1617), .dout(n1621));
    jand g0350(.dinb(n1605), .dina(n1621), .dout(n1625));
    jand g0351(.dinb(n1589), .dina(n13869), .dout(n1629));
    jand g0352(.dinb(n1555), .dina(n8139), .dout(n1633));
    jxor g0353(.dinb(G308), .dina(G316), .dout(n1637));
    jxor g0354(.dinb(G341), .dina(G351), .dout(n1641));
    jxor g0355(.dinb(n1637), .dina(n1641), .dout(n1645));
    jxor g0356(.dinb(G361), .dina(G369), .dout(n1649));
    jxor g0357(.dinb(n753), .dina(n1649), .dout(n1653));
    jxor g0358(.dinb(n659), .dina(n14624), .dout(n1657));
    jxor g0359(.dinb(n1653), .dina(n1657), .dout(n1661));
    jxor g0360(.dinb(n9981), .dina(n1661), .dout(n1665));
    jnot g0361(.din(n1665), .dout(n1668));
    jxor g0362(.dinb(G218), .dina(G226), .dout(n1672));
    jxor g0363(.dinb(G265), .dina(G273), .dout(n1676));
    jxor g0364(.dinb(n1672), .dina(n1676), .dout(n1680));
    jxor g0365(.dinb(G281), .dina(G289), .dout(n1684));
    jxor g0366(.dinb(G234), .dina(G257), .dout(n1688));
    jxor g0367(.dinb(n1684), .dina(n1688), .dout(n1692));
    jxor g0368(.dinb(n1113), .dina(n16031), .dout(n1696));
    jxor g0369(.dinb(n1692), .dina(n1696), .dout(n1700));
    jxor g0370(.dinb(n9987), .dina(n1700), .dout(n1704));
    jnot g0371(.din(n1704), .dout(n1707));
    jnot g0372(.din(n1274), .dout(n1710));
    jand g0373(.dinb(n16226), .dina(n1710), .dout(n1714));
    jnot g0374(.din(n1714), .dout(n1717));
    jand g0375(.dinb(n16262), .dina(n1274), .dout(n1721));
    jnot g0376(.din(n1338), .dout(n1724));
    jand g0377(.dinb(n15686), .dina(n1724), .dout(n1728));
    jor g0378(.dinb(n15923), .dina(n1724), .dout(n1732));
    jand g0379(.dinb(n15587), .dina(n1357), .dout(n1736));
    jor g0380(.dinb(n15998), .dina(n1296), .dout(n1740));
    jor g0381(.dinb(n1740), .dina(n1316), .dout(n1744));
    jnot g0382(.din(G280), .dout(n1747));
    jand g0383(.dinb(n1747), .dina(n15749), .dout(n1751));
    jnot g0384(.din(n1308), .dout(n1754));
    jor g0385(.dinb(n1751), .dina(n1754), .dout(n1758));
    jor g0386(.dinb(n15896), .dina(n1758), .dout(n1762));
    jor g0387(.dinb(n15959), .dina(n1357), .dout(n1766));
    jand g0388(.dinb(n1762), .dina(n1766), .dout(n1770));
    jand g0389(.dinb(n1744), .dina(n1770), .dout(n1774));
    jor g0390(.dinb(n15581), .dina(n1774), .dout(n1778));
    jand g0391(.dinb(n15590), .dina(n1778), .dout(n1782));
    jor g0392(.dinb(n15596), .dina(n1782), .dout(n1786));
    jnot g0393(.din(n1786), .dout(n1789));
    jor g0394(.dinb(n15534), .dina(n1789), .dout(n1793));
    jand g0395(.dinb(n15519), .dina(n1793), .dout(n1797));
    jand g0396(.dinb(n8171), .dina(n1797), .dout(n1801));
    jand g0397(.dinb(n16190), .dina(n1407), .dout(n1805));
    jor g0398(.dinb(n16178), .dina(n1407), .dout(n1809));
    jor g0399(.dinb(n16040), .dina(n1388), .dout(n1813));
    jand g0400(.dinb(n16040), .dina(n1388), .dout(n1817));
    jand g0401(.dinb(n16094), .dina(n1443), .dout(n1821));
    jand g0402(.dinb(n16124), .dina(n1427), .dout(n1825));
    jand g0403(.dinb(n1825), .dina(n1447), .dout(n1829));
    jor g0404(.dinb(n15294), .dina(n1829), .dout(n1833));
    jor g0405(.dinb(n15285), .dina(n1833), .dout(n1837));
    jand g0406(.dinb(n15269), .dina(n1837), .dout(n1841));
    jand g0407(.dinb(n8169), .dina(n1841), .dout(n1845));
    jor g0408(.dinb(n8160), .dina(n1845), .dout(n1849));
    jor g0409(.dinb(n1801), .dina(n8148), .dout(n1853));
    jand g0410(.dinb(n14450), .dina(n1477), .dout(n1857));
    jor g0411(.dinb(n14255), .dina(n1520), .dout(n1861));
    jand g0412(.dinb(n14516), .dina(n1520), .dout(n1865));
    jand g0413(.dinb(n14240), .dina(n306), .dout(n1869));
    jand g0414(.dinb(n1462), .dina(n795), .dout(n1873));
    jor g0415(.dinb(n1869), .dina(n1873), .dout(n1877));
    jand g0416(.dinb(n14243), .dina(n1877), .dout(n1881));
    jand g0417(.dinb(n14291), .dina(n322), .dout(n1885));
    jand g0418(.dinb(n1462), .dina(n611), .dout(n1889));
    jor g0419(.dinb(n1885), .dina(n1889), .dout(n1893));
    jand g0420(.dinb(n14216), .dina(n1893), .dout(n1897));
    jor g0421(.dinb(n1897), .dina(n14192), .dout(n1901));
    jor g0422(.dinb(n14474), .dina(n1893), .dout(n1905));
    jor g0423(.dinb(n14648), .dina(n1877), .dout(n1909));
    jand g0424(.dinb(n1905), .dina(n1909), .dout(n1913));
    jand g0425(.dinb(n1901), .dina(n1913), .dout(n1917));
    jor g0426(.dinb(n14231), .dina(n1917), .dout(n1921));
    jor g0427(.dinb(n14187), .dina(n1921), .dout(n1925));
    jand g0428(.dinb(n14175), .dina(n1925), .dout(n1929));
    jnot g0429(.din(n1929), .dout(n1932));
    jand g0430(.dinb(n14258), .dina(n1932), .dout(n1936));
    jor g0431(.dinb(n14160), .dina(n1936), .dout(n1940));
    jand g0432(.dinb(n8204), .dina(n1940), .dout(n1944));
    jnot g0433(.din(n1589), .dout(n1947));
    jnot g0434(.din(n1601), .dout(n1950));
    jand g0435(.dinb(n14588), .dina(n1950), .dout(n1954));
    jnot g0436(.din(n1954), .dout(n1957));
    jand g0437(.dinb(n14603), .dina(n1601), .dout(n1961));
    jand g0438(.dinb(n14570), .dina(n1617), .dout(n1965));
    jor g0439(.dinb(n1961), .dina(n1965), .dout(n1969));
    jand g0440(.dinb(n1957), .dina(n13901), .dout(n1973));
    jor g0441(.dinb(n1947), .dina(n1973), .dout(n1977));
    jor g0442(.dinb(n1944), .dina(n8202), .dout(n1981));
    jnot g0443(.din(G54), .dout(n1984));
    jxor g0444(.dinb(n9642), .dina(n1509), .dout(n1988));
    jnot g0445(.din(G4092), .dout(n1991));
    jand g0446(.dinb(n15827), .dina(n1991), .dout(n1995));
    jnot g0447(.din(n1995), .dout(n1998));
    jor g0448(.dinb(n1988), .dina(n11337), .dout(n2002));
    jnot g0449(.din(G4091), .dout(n2005));
    jand g0450(.dinb(n2005), .dina(n1991), .dout(n2009));
    jand g0451(.dinb(n735), .dina(n11429), .dout(n2013));
    jand g0452(.dinb(n2005), .dina(n16319), .dout(n2017));
    jand g0453(.dinb(n8361), .dina(n2017), .dout(n2021));
    jor g0454(.dinb(n2013), .dina(n8355), .dout(n2025));
    jnot g0455(.din(n2025), .dout(n2028));
    jand g0456(.dinb(n8352), .dina(n2028), .dout(n2032));
    jnot g0457(.din(n1497), .dout(n2035));
    jand g0458(.dinb(n9642), .dina(n1509), .dout(n2039));
    jnot g0459(.din(n2039), .dout(n2042));
    jand g0460(.dinb(n2035), .dina(n2042), .dout(n2046));
    jand g0461(.dinb(n1497), .dina(n2039), .dout(n2050));
    jor g0462(.dinb(n9323), .dina(n2050), .dout(n2054));
    jor g0463(.dinb(n2046), .dina(n2054), .dout(n2058));
    jnot g0464(.din(n2009), .dout(n2061));
    jor g0465(.dinb(n656), .dina(n11427), .dout(n2065));
    jand g0466(.dinb(n9312), .dina(n2017), .dout(n2069));
    jnot g0467(.din(n2069), .dout(n2072));
    jand g0468(.dinb(n2065), .dina(n9306), .dout(n2076));
    jand g0469(.dinb(n2058), .dina(n2076), .dout(n2080));
    jxor g0470(.dinb(n11856), .dina(n1300), .dout(n2084));
    jand g0471(.dinb(n11363), .dina(n2084), .dout(n2088));
    jnot g0472(.din(n2088), .dout(n2091));
    jor g0473(.dinb(n1064), .dina(n11427), .dout(n2095));
    jand g0474(.dinb(n8373), .dina(n2017), .dout(n2099));
    jnot g0475(.din(n2099), .dout(n2102));
    jand g0476(.dinb(n2095), .dina(n8367), .dout(n2106));
    jand g0477(.dinb(n2091), .dina(n2106), .dout(n2110));
    jnot g0478(.din(n1567), .dout(n2113));
    jand g0479(.dinb(n11615), .dina(n1555), .dout(n2117));
    jor g0480(.dinb(n1940), .dina(n11613), .dout(n2121));
    jand g0481(.dinb(n13847), .dina(n2121), .dout(n2125));
    jor g0482(.dinb(n11639), .dina(n2125), .dout(n2129));
    jnot g0483(.din(n2129), .dout(n2132));
    jor g0484(.dinb(n13697), .dina(n2132), .dout(n2136));
    jxor g0485(.dinb(n2113), .dina(n1582), .dout(n2140));
    jnot g0486(.din(n2140), .dout(n2143));
    jor g0487(.dinb(n2129), .dina(n13695), .dout(n2147));
    jand g0488(.dinb(n2136), .dina(n11604), .dout(n2151));
    jnot g0489(.din(n2151), .dout(n2154));
    jnot g0490(.din(n2110), .dout(n2157));
    jnot g0491(.din(G4087), .dout(n2160));
    jand g0492(.dinb(n2160), .dina(n12404), .dout(n2164));
    jand g0493(.dinb(n2157), .dina(n12402), .dout(n2168));
    jnot g0494(.din(n2032), .dout(n2171));
    jnot g0495(.din(G4088), .dout(n2174));
    jand g0496(.dinb(n2160), .dina(n2174), .dout(n2178));
    jand g0497(.dinb(n2171), .dina(n12264), .dout(n2182));
    jand g0498(.dinb(n12407), .dina(n2174), .dout(n2186));
    jand g0499(.dinb(n8265), .dina(n2186), .dout(n2190));
    jand g0500(.dinb(G4087), .dina(G4088), .dout(n2194));
    jand g0501(.dinb(n8259), .dina(n2194), .dout(n2198));
    jor g0502(.dinb(n2190), .dina(n8238), .dout(n2202));
    jor g0503(.dinb(n2182), .dina(n8235), .dout(n2206));
    jor g0504(.dinb(n2168), .dina(n2206), .dout(n2210));
    jand g0505(.dinb(n14051), .dina(n1929), .dout(n2214));
    jand g0506(.dinb(n9467), .dina(n1929), .dout(n2218));
    jor g0507(.dinb(n2214), .dina(n2218), .dout(n2222));
    jxor g0508(.dinb(n13628), .dina(n2222), .dout(n2226));
    jor g0509(.dinb(n9650), .dina(n2226), .dout(n2230));
    jor g0510(.dinb(n792), .dina(n11427), .dout(n2234));
    jand g0511(.dinb(n9171), .dina(n2017), .dout(n2238));
    jnot g0512(.din(n2238), .dout(n2241));
    jand g0513(.dinb(n2234), .dina(n9165), .dout(n2245));
    jand g0514(.dinb(n2230), .dina(n9159), .dout(n2249));
    jnot g0515(.din(n1524), .dout(n2252));
    jand g0516(.dinb(n9626), .dina(n1921), .dout(n2256));
    jand g0517(.dinb(n14081), .dina(n1917), .dout(n2260));
    jor g0518(.dinb(n14222), .dina(n2260), .dout(n2264));
    jor g0519(.dinb(n2256), .dina(n2264), .dout(n2268));
    jxor g0520(.dinb(n9624), .dina(n2268), .dout(n2272));
    jor g0521(.dinb(n9644), .dina(n2272), .dout(n2276));
    jand g0522(.dinb(n717), .dina(n11756), .dout(n2280));
    jand g0523(.dinb(n9606), .dina(n2017), .dout(n2284));
    jor g0524(.dinb(n2280), .dina(n9600), .dout(n2288));
    jnot g0525(.din(n2288), .dout(n2291));
    jand g0526(.dinb(n2276), .dina(n9597), .dout(n2295));
    jor g0527(.dinb(n14480), .dina(n1493), .dout(n2299));
    jand g0528(.dinb(n14504), .dina(n1493), .dout(n2303));
    jor g0529(.dinb(n13610), .dina(n2042), .dout(n2307));
    jand g0530(.dinb(n13664), .dina(n2307), .dout(n2311));
    jxor g0531(.dinb(n14060), .dina(n2311), .dout(n2315));
    jor g0532(.dinb(n11324), .dina(n2315), .dout(n2319));
    jor g0533(.dinb(n834), .dina(n11427), .dout(n2323));
    jand g0534(.dinb(n9459), .dina(n2017), .dout(n2327));
    jnot g0535(.din(n2327), .dout(n2330));
    jand g0536(.dinb(n2323), .dina(n9453), .dout(n2334));
    jand g0537(.dinb(n2319), .dina(n9447), .dout(n2338));
    jnot g0538(.din(G4090), .dout(n2341));
    jand g0539(.dinb(n12746), .dina(n2341), .dout(n2345));
    jand g0540(.dinb(n2157), .dina(n12741), .dout(n2349));
    jnot g0541(.din(G4089), .dout(n2352));
    jand g0542(.dinb(n2352), .dina(n2341), .dout(n2356));
    jand g0543(.dinb(n2171), .dina(n12603), .dout(n2360));
    jand g0544(.dinb(n2352), .dina(n12743), .dout(n2364));
    jand g0545(.dinb(n8265), .dina(n2364), .dout(n2368));
    jand g0546(.dinb(G4089), .dina(G4090), .dout(n2372));
    jand g0547(.dinb(n8259), .dina(n2372), .dout(n2376));
    jor g0548(.dinb(n2368), .dina(n8256), .dout(n2380));
    jor g0549(.dinb(n2360), .dina(n8253), .dout(n2384));
    jor g0550(.dinb(n2349), .dina(n2384), .dout(n2388));
    jnot g0551(.din(n1728), .dout(n2391));
    jnot g0552(.din(n1732), .dout(n2394));
    jor g0553(.dinb(n1326), .dina(n15374), .dout(n2398));
    jand g0554(.dinb(n15536), .dina(n2398), .dout(n2402));
    jnot g0555(.din(n2402), .dout(n2405));
    jnot g0556(.din(n1778), .dout(n2408));
    jor g0557(.dinb(n9710), .dina(n2408), .dout(n2412));
    jand g0558(.dinb(n2405), .dina(n9708), .dout(n2416));
    jor g0559(.dinb(n15083), .dina(n2416), .dout(n2420));
    jand g0560(.dinb(n9261), .dina(n2420), .dout(n2424));
    jxor g0561(.dinb(n15410), .dina(n2424), .dout(n2428));
    jor g0562(.dinb(n11294), .dina(n2428), .dout(n2432));
    jor g0563(.dinb(n930), .dina(n11427), .dout(n2436));
    jand g0564(.dinb(n9237), .dina(n2017), .dout(n2440));
    jnot g0565(.din(n2440), .dout(n2443));
    jand g0566(.dinb(n2436), .dina(n9231), .dout(n2447));
    jand g0567(.dinb(n2432), .dina(n9225), .dout(n2451));
    jxor g0568(.dinb(n15656), .dina(n2416), .dout(n2455));
    jor g0569(.dinb(n11300), .dina(n2455), .dout(n2459));
    jor g0570(.dinb(n972), .dina(n11427), .dout(n2463));
    jand g0571(.dinb(n9699), .dina(n2017), .dout(n2467));
    jnot g0572(.din(n2467), .dout(n2470));
    jand g0573(.dinb(n2463), .dina(n9693), .dout(n2474));
    jand g0574(.dinb(n2459), .dina(n9687), .dout(n2478));
    jand g0575(.dinb(n11856), .dina(n1300), .dout(n2482));
    jnot g0576(.din(n2482), .dout(n2485));
    jand g0577(.dinb(n15575), .dina(n2485), .dout(n2489));
    jor g0578(.dinb(n15557), .dina(n2489), .dout(n2493));
    jand g0579(.dinb(n15545), .dina(n2493), .dout(n2497));
    jxor g0580(.dinb(n15641), .dina(n2497), .dout(n2501));
    jand g0581(.dinb(n11339), .dina(n2501), .dout(n2505));
    jnot g0582(.din(n2505), .dout(n2508));
    jor g0583(.dinb(n888), .dina(n11427), .dout(n2512));
    jand g0584(.dinb(n9510), .dina(n2017), .dout(n2516));
    jnot g0585(.din(n2516), .dout(n2519));
    jand g0586(.dinb(n2512), .dina(n9504), .dout(n2523));
    jand g0587(.dinb(n2508), .dina(n9498), .dout(n2527));
    jand g0588(.dinb(n1740), .dina(n1316), .dout(n2531));
    jand g0589(.dinb(n2485), .dina(n9357), .dout(n2535));
    jnot g0590(.din(n2535), .dout(n2538));
    jand g0591(.dinb(n2493), .dina(n2538), .dout(n2542));
    jand g0592(.dinb(n11945), .dina(n2542), .dout(n2546));
    jnot g0593(.din(n2546), .dout(n2549));
    jor g0594(.dinb(n1022), .dina(n11427), .dout(n2553));
    jand g0595(.dinb(n9348), .dina(n2017), .dout(n2557));
    jnot g0596(.din(n2557), .dout(n2560));
    jand g0597(.dinb(n2553), .dina(n9342), .dout(n2564));
    jand g0598(.dinb(n2549), .dina(n9336), .dout(n2568));
    jxor g0599(.dinb(n1950), .dina(n13946), .dout(n2572));
    jxor g0600(.dinb(n2140), .dina(n2572), .dout(n2576));
    jxor g0601(.dinb(n10010), .dina(n2576), .dout(n2580));
    jand g0602(.dinb(n1462), .dina(n10007), .dout(n2584));
    jand g0603(.dinb(G332), .dina(G372), .dout(n2588));
    jor g0604(.dinb(n2584), .dina(n10005), .dout(n2592));
    jxor g0605(.dinb(n1493), .dina(n2592), .dout(n2596));
    jxor g0606(.dinb(n14069), .dina(n2596), .dout(n2600));
    jnot g0607(.din(G331), .dout(n2603));
    jand g0608(.dinb(n10002), .dina(n1520), .dout(n2607));
    jnot g0609(.din(n1520), .dout(n2610));
    jand g0610(.dinb(n1477), .dina(n9999), .dout(n2614));
    jor g0611(.dinb(n9996), .dina(n2614), .dout(n2618));
    jxor g0612(.dinb(n9990), .dina(n2618), .dout(n2622));
    jxor g0613(.dinb(n2580), .dina(n2622), .dout(n2626));
    jnot g0614(.din(n2626), .dout(n2629));
    jxor g0615(.dinb(n1296), .dina(n1338), .dout(n2633));
    jxor g0616(.dinb(n1312), .dina(n1357), .dout(n2637));
    jxor g0617(.dinb(n2633), .dina(n2637), .dout(n2641));
    jxor g0618(.dinb(n15734), .dina(n2641), .dout(n2645));
    jand g0619(.dinb(n10022), .dina(n1259), .dout(n2649));
    jand g0620(.dinb(G292), .dina(G335), .dout(n2653));
    jor g0621(.dinb(n2649), .dina(n10020), .dout(n2657));
    jxor g0622(.dinb(n1427), .dina(n2657), .dout(n2661));
    jxor g0623(.dinb(n1274), .dina(n2661), .dout(n2665));
    jxor g0624(.dinb(n1407), .dina(n15296), .dout(n2669));
    jxor g0625(.dinb(n2665), .dina(n2669), .dout(n2673));
    jxor g0626(.dinb(n2645), .dina(n2673), .dout(n2677));
    jnot g0627(.din(n1411), .dout(n2680));
    jnot g0628(.din(n1841), .dout(n2683));
    jnot g0629(.din(n1813), .dout(n2686));
    jnot g0630(.din(n1447), .dout(n2689));
    jnot g0631(.din(n1431), .dout(n2692));
    jnot g0632(.din(n1797), .dout(n2695));
    jand g0633(.dinb(n11828), .dina(n1376), .dout(n2699));
    jnot g0634(.din(n2699), .dout(n2702));
    jand g0635(.dinb(n2695), .dina(n11826), .dout(n2706));
    jor g0636(.dinb(n11883), .dina(n2706), .dout(n2710));
    jor g0637(.dinb(n11823), .dina(n2710), .dout(n2714));
    jor g0638(.dinb(n15236), .dina(n2714), .dout(n2718));
    jand g0639(.dinb(n11793), .dina(n2718), .dout(n2722));
    jxor g0640(.dinb(n15305), .dina(n2722), .dout(n2726));
    jnot g0641(.din(n2726), .dout(n2729));
    jnot g0642(.din(n1392), .dout(n2732));
    jnot g0643(.din(n1833), .dout(n2735));
    jand g0644(.dinb(n15209), .dina(n2714), .dout(n2739));
    jxor g0645(.dinb(n15695), .dina(n2739), .dout(n2743));
    jnot g0646(.din(n2743), .dout(n2746));
    jor g0647(.dinb(n16124), .dina(n1427), .dout(n2750));
    jnot g0648(.din(n2750), .dout(n2753));
    jnot g0649(.din(n1825), .dout(n2756));
    jand g0650(.dinb(n11103), .dina(n2706), .dout(n2760));
    jor g0651(.dinb(n11076), .dina(n2760), .dout(n2764));
    jxor g0652(.dinb(n15173), .dina(n2764), .dout(n2768));
    jxor g0653(.dinb(n11883), .dina(n2706), .dout(n2772));
    jnot g0654(.din(n2772), .dout(n2775));
    jnot g0655(.din(n2501), .dout(n2778));
    jnot g0656(.din(n2084), .dout(n2781));
    jnot g0657(.din(n2542), .dout(n2784));
    jand g0658(.dinb(n8286), .dina(n2784), .dout(n2788));
    jand g0659(.dinb(n2778), .dina(n2788), .dout(n2792));
    jand g0660(.dinb(n2455), .dina(n2792), .dout(n2796));
    jand g0661(.dinb(n2428), .dina(n8274), .dout(n2800));
    jand g0662(.dinb(n2775), .dina(n8271), .dout(n2804));
    jand g0663(.dinb(n2768), .dina(n2804), .dout(n2808));
    jand g0664(.dinb(n2746), .dina(n8268), .dout(n2812));
    jand g0665(.dinb(n2729), .dina(n2812), .dout(n2816));
    jnot g0666(.din(n1605), .dout(n2819));
    jor g0667(.dinb(n14561), .dina(n1617), .dout(n2823));
    jor g0668(.dinb(n13904), .dina(n2121), .dout(n2827));
    jand g0669(.dinb(n13793), .dina(n2827), .dout(n2831));
    jxor g0670(.dinb(n10995), .dina(n2831), .dout(n2835));
    jxor g0671(.dinb(n13955), .dina(n2129), .dout(n2839));
    jxor g0672(.dinb(n13871), .dina(n2121), .dout(n2843));
    jnot g0673(.din(n2843), .dout(n2846));
    jor g0674(.dinb(n9642), .dina(n1509), .dout(n2850));
    jand g0675(.dinb(n13739), .dina(n2850), .dout(n2854));
    jand g0676(.dinb(n2046), .dina(n8304), .dout(n2858));
    jand g0677(.dinb(n2315), .dina(n8301), .dout(n2862));
    jand g0678(.dinb(n2272), .dina(n8298), .dout(n2866));
    jand g0679(.dinb(n2226), .dina(n8295), .dout(n2870));
    jand g0680(.dinb(n2846), .dina(n8292), .dout(n2874));
    jand g0681(.dinb(n2839), .dina(n2874), .dout(n2878));
    jand g0682(.dinb(n10964), .dina(n2878), .dout(n2882));
    jnot g0683(.din(G1690), .dout(n2885));
    jand g0684(.dinb(n13229), .dina(n2885), .dout(n2889));
    jand g0685(.dinb(n2157), .dina(n13064), .dout(n2893));
    jnot g0686(.din(G1689), .dout(n2896));
    jand g0687(.dinb(n2896), .dina(n2885), .dout(n2900));
    jand g0688(.dinb(n2171), .dina(n12866), .dout(n2904));
    jand g0689(.dinb(n2896), .dina(n13226), .dout(n2908));
    jand g0690(.dinb(n8349), .dina(n2908), .dout(n2912));
    jand g0691(.dinb(G1689), .dina(G1690), .dout(n2916));
    jand g0692(.dinb(n8343), .dina(n2916), .dout(n2920));
    jor g0693(.dinb(n2912), .dina(n8322), .dout(n2924));
    jor g0694(.dinb(n2904), .dina(n8319), .dout(n2928));
    jor g0695(.dinb(n2893), .dina(n2928), .dout(n2932));
    jand g0696(.dinb(n16679), .dina(n2932), .dout(n2936));
    jnot g0697(.din(G1694), .dout(n2939));
    jand g0698(.dinb(n16487), .dina(n2939), .dout(n2943));
    jand g0699(.dinb(n2157), .dina(n16322), .dout(n2947));
    jnot g0700(.din(G1691), .dout(n2950));
    jand g0701(.dinb(n2950), .dina(n2939), .dout(n2954));
    jand g0702(.dinb(n2171), .dina(n14711), .dout(n2958));
    jand g0703(.dinb(n2950), .dina(n16484), .dout(n2962));
    jand g0704(.dinb(n8349), .dina(n2962), .dout(n2966));
    jand g0705(.dinb(G1691), .dina(G1694), .dout(n2970));
    jand g0706(.dinb(n8343), .dina(n2970), .dout(n2974));
    jor g0707(.dinb(n2966), .dina(n8340), .dout(n2978));
    jor g0708(.dinb(n2958), .dina(n8337), .dout(n2982));
    jor g0709(.dinb(n2947), .dina(n2982), .dout(n2986));
    jand g0710(.dinb(n16679), .dina(n2986), .dout(n2990));
    jnot g0711(.din(n2451), .dout(n2993));
    jand g0712(.dinb(n8444), .dina(n2993), .dout(n2997));
    jnot g0713(.din(n2249), .dout(n3000));
    jand g0714(.dinb(n8423), .dina(n3000), .dout(n3004));
    jand g0715(.dinb(n8643), .dina(n2186), .dout(n3008));
    jand g0716(.dinb(n8637), .dina(n2194), .dout(n3012));
    jor g0717(.dinb(n3008), .dina(n8421), .dout(n3016));
    jor g0718(.dinb(n3004), .dina(n8418), .dout(n3020));
    jor g0719(.dinb(n2997), .dina(n8382), .dout(n3024));
    jnot g0720(.din(n2478), .dout(n3027));
    jand g0721(.dinb(n8588), .dina(n3027), .dout(n3031));
    jnot g0722(.din(n2295), .dout(n3034));
    jand g0723(.dinb(n8573), .dina(n3034), .dout(n3038));
    jand g0724(.dinb(n8733), .dina(n2186), .dout(n3042));
    jand g0725(.dinb(n8727), .dina(n2194), .dout(n3046));
    jor g0726(.dinb(n3042), .dina(n8502), .dout(n3050));
    jor g0727(.dinb(n3038), .dina(n8499), .dout(n3054));
    jor g0728(.dinb(n3031), .dina(n8469), .dout(n3058));
    jnot g0729(.din(n2527), .dout(n3061));
    jand g0730(.dinb(n8585), .dina(n3061), .dout(n3065));
    jnot g0731(.din(n2338), .dout(n3068));
    jand g0732(.dinb(n8567), .dina(n3068), .dout(n3072));
    jand g0733(.dinb(n8775), .dina(n2186), .dout(n3076));
    jand g0734(.dinb(n8769), .dina(n2194), .dout(n3080));
    jor g0735(.dinb(n3076), .dina(n8535), .dout(n3084));
    jor g0736(.dinb(n3072), .dina(n8532), .dout(n3088));
    jor g0737(.dinb(n3065), .dina(n8508), .dout(n3092));
    jnot g0738(.din(n2568), .dout(n3095));
    jand g0739(.dinb(n12371), .dina(n3095), .dout(n3099));
    jnot g0740(.din(n2080), .dout(n3102));
    jand g0741(.dinb(n3102), .dina(n12245), .dout(n3106));
    jand g0742(.dinb(n8814), .dina(n2186), .dout(n3110));
    jand g0743(.dinb(n8808), .dina(n2194), .dout(n3114));
    jor g0744(.dinb(n3110), .dina(n8565), .dout(n3118));
    jor g0745(.dinb(n3106), .dina(n8562), .dout(n3122));
    jor g0746(.dinb(n3099), .dina(n8544), .dout(n3126));
    jand g0747(.dinb(n8666), .dina(n2993), .dout(n3130));
    jand g0748(.dinb(n3000), .dina(n8645), .dout(n3134));
    jand g0749(.dinb(n8643), .dina(n2364), .dout(n3138));
    jand g0750(.dinb(n8637), .dina(n2372), .dout(n3142));
    jor g0751(.dinb(n3138), .dina(n8634), .dout(n3146));
    jor g0752(.dinb(n3134), .dina(n8631), .dout(n3150));
    jor g0753(.dinb(n3130), .dina(n8595), .dout(n3154));
    jand g0754(.dinb(n8837), .dina(n3027), .dout(n3158));
    jand g0755(.dinb(n3034), .dina(n8822), .dout(n3162));
    jand g0756(.dinb(n8733), .dina(n2364), .dout(n3166));
    jand g0757(.dinb(n8727), .dina(n2372), .dout(n3170));
    jor g0758(.dinb(n3166), .dina(n8724), .dout(n3174));
    jor g0759(.dinb(n3162), .dina(n8721), .dout(n3178));
    jor g0760(.dinb(n3158), .dina(n8691), .dout(n3182));
    jand g0761(.dinb(n8834), .dina(n3061), .dout(n3186));
    jand g0762(.dinb(n3068), .dina(n8816), .dout(n3190));
    jand g0763(.dinb(n8775), .dina(n2364), .dout(n3194));
    jand g0764(.dinb(n8769), .dina(n2372), .dout(n3198));
    jor g0765(.dinb(n3194), .dina(n8766), .dout(n3202));
    jor g0766(.dinb(n3190), .dina(n8763), .dout(n3206));
    jor g0767(.dinb(n3186), .dina(n8739), .dout(n3210));
    jand g0768(.dinb(n12710), .dina(n3095), .dout(n3214));
    jand g0769(.dinb(n3102), .dina(n12584), .dout(n3218));
    jand g0770(.dinb(n8814), .dina(n2364), .dout(n3222));
    jand g0771(.dinb(n8808), .dina(n2372), .dout(n3226));
    jor g0772(.dinb(n3222), .dina(n8805), .dout(n3230));
    jor g0773(.dinb(n3218), .dina(n8802), .dout(n3234));
    jor g0774(.dinb(n3214), .dina(n8784), .dout(n3238));
    jand g0775(.dinb(n2993), .dina(n8906), .dout(n3242));
    jand g0776(.dinb(n3000), .dina(n8885), .dout(n3246));
    jand g0777(.dinb(n9120), .dina(n2908), .dout(n3250));
    jand g0778(.dinb(n9114), .dina(n2916), .dout(n3254));
    jor g0779(.dinb(n3250), .dina(n8883), .dout(n3258));
    jor g0780(.dinb(n3246), .dina(n8880), .dout(n3262));
    jor g0781(.dinb(n3242), .dina(n8844), .dout(n3266));
    jand g0782(.dinb(n8996), .dina(n3266), .dout(n3270));
    jand g0783(.dinb(n3095), .dina(n13193), .dout(n3274));
    jand g0784(.dinb(n3102), .dina(n12986), .dout(n3278));
    jand g0785(.dinb(n9300), .dina(n2908), .dout(n3282));
    jand g0786(.dinb(n9294), .dina(n2916), .dout(n3286));
    jor g0787(.dinb(n3282), .dina(n8958), .dout(n3290));
    jor g0788(.dinb(n3278), .dina(n8955), .dout(n3294));
    jor g0789(.dinb(n3274), .dina(n8937), .dout(n3298));
    jand g0790(.dinb(n9389), .dina(n3298), .dout(n3302));
    jand g0791(.dinb(n3061), .dina(n9068), .dout(n3306));
    jand g0792(.dinb(n3068), .dina(n9056), .dout(n3310));
    jand g0793(.dinb(n9441), .dina(n2908), .dout(n3314));
    jand g0794(.dinb(n9435), .dina(n2916), .dout(n3318));
    jor g0795(.dinb(n3314), .dina(n8991), .dout(n3322));
    jor g0796(.dinb(n3310), .dina(n8988), .dout(n3326));
    jor g0797(.dinb(n3306), .dina(n8964), .dout(n3330));
    jand g0798(.dinb(n8993), .dina(n3330), .dout(n3334));
    jand g0799(.dinb(n3027), .dina(n9062), .dout(n3338));
    jand g0800(.dinb(n3034), .dina(n9044), .dout(n3342));
    jand g0801(.dinb(n9564), .dina(n2908), .dout(n3346));
    jand g0802(.dinb(n9558), .dina(n2916), .dout(n3350));
    jor g0803(.dinb(n3346), .dina(n9042), .dout(n3354));
    jor g0804(.dinb(n3342), .dina(n9039), .dout(n3358));
    jor g0805(.dinb(n3338), .dina(n9009), .dout(n3362));
    jand g0806(.dinb(n9371), .dina(n3362), .dout(n3366));
    jand g0807(.dinb(n2993), .dina(n9179), .dout(n3370));
    jand g0808(.dinb(n3000), .dina(n9122), .dout(n3374));
    jand g0809(.dinb(n9120), .dina(n2962), .dout(n3378));
    jand g0810(.dinb(n9114), .dina(n2970), .dout(n3382));
    jor g0811(.dinb(n3378), .dina(n9111), .dout(n3386));
    jor g0812(.dinb(n3374), .dina(n9108), .dout(n3390));
    jor g0813(.dinb(n3370), .dina(n9072), .dout(n3394));
    jand g0814(.dinb(n9359), .dina(n3394), .dout(n3398));
    jand g0815(.dinb(n3095), .dina(n16451), .dout(n3402));
    jand g0816(.dinb(n3102), .dina(n14831), .dout(n3406));
    jand g0817(.dinb(n9300), .dina(n2962), .dout(n3410));
    jand g0818(.dinb(n9294), .dina(n2970), .dout(n3414));
    jor g0819(.dinb(n3410), .dina(n9291), .dout(n3418));
    jor g0820(.dinb(n3406), .dina(n9288), .dout(n3422));
    jor g0821(.dinb(n3402), .dina(n9270), .dout(n3426));
    jand g0822(.dinb(n9377), .dina(n3426), .dout(n3430));
    jand g0823(.dinb(n3061), .dina(n9668), .dout(n3434));
    jand g0824(.dinb(n3068), .dina(n9578), .dout(n3438));
    jand g0825(.dinb(n9441), .dina(n2962), .dout(n3442));
    jand g0826(.dinb(n9435), .dina(n2970), .dout(n3446));
    jor g0827(.dinb(n3442), .dina(n9432), .dout(n3450));
    jor g0828(.dinb(n3438), .dina(n9429), .dout(n3454));
    jor g0829(.dinb(n3434), .dina(n9405), .dout(n3458));
    jand g0830(.dinb(n16631), .dina(n3458), .dout(n3462));
    jand g0831(.dinb(n3027), .dina(n9662), .dout(n3466));
    jand g0832(.dinb(n3034), .dina(n9566), .dout(n3470));
    jand g0833(.dinb(n9564), .dina(n2962), .dout(n3474));
    jand g0834(.dinb(n9558), .dina(n2970), .dout(n3478));
    jor g0835(.dinb(n3474), .dina(n9555), .dout(n3482));
    jor g0836(.dinb(n3470), .dina(n9552), .dout(n3486));
    jor g0837(.dinb(n3466), .dina(n9522), .dout(n3490));
    jand g0838(.dinb(n10544), .dina(n3490), .dout(n3494));
    jand g0839(.dinb(n9863), .dina(n2151), .dout(n3498));
    jnot g0840(.din(G3717), .dout(n3501));
    jnot g0841(.din(G3724), .dout(n3504));
    jand g0842(.dinb(n11601), .dina(n3504), .dout(n3508));
    jor g0843(.dinb(n9825), .dina(n3508), .dout(n3512));
    jor g0844(.dinb(n3498), .dina(n9822), .dout(n3516));
    jnot g0845(.din(G135), .dout(n3519));
    jnot g0846(.din(G4115), .dout(n3522));
    jor g0847(.dinb(n3519), .dina(n3522), .dout(n3526));
    jxor g0848(.dinb(n9963), .dina(n1567), .dout(n3530));
    jand g0849(.dinb(n9851), .dina(n3530), .dout(n3534));
    jnot g0850(.din(n671), .dout(n3537));
    jand g0851(.dinb(n9827), .dina(n3537), .dout(n3541));
    jor g0852(.dinb(n9836), .dina(n3541), .dout(n3545));
    jor g0853(.dinb(n9774), .dina(n3545), .dout(n3549));
    jand g0854(.dinb(n9771), .dina(n3549), .dout(n3553));
    jand g0855(.dinb(n3516), .dina(n9756), .dout(n3557));
    jor g0856(.dinb(n14003), .dina(n2129), .dout(n3561));
    jxor g0857(.dinb(n9917), .dina(n3561), .dout(n3565));
    jand g0858(.dinb(n11675), .dina(n2151), .dout(n3569));
    jand g0859(.dinb(n11597), .dina(n2017), .dout(n3573));
    jand g0860(.dinb(n3537), .dina(n11594), .dout(n3577));
    jor g0861(.dinb(n11592), .dina(n3577), .dout(n3581));
    jor g0862(.dinb(n3569), .dina(n11586), .dout(n3585));
    jnot g0863(.din(n3585), .dout(n3588));
    jor g0864(.dinb(n11282), .dina(n2839), .dout(n3592));
    jand g0865(.dinb(n692), .dina(n11756), .dout(n3596));
    jand g0866(.dinb(n11280), .dina(n2017), .dout(n3600));
    jor g0867(.dinb(n3596), .dina(n11274), .dout(n3604));
    jnot g0868(.din(n3604), .dout(n3607));
    jand g0869(.dinb(n3592), .dina(n11271), .dout(n3611));
    jor g0870(.dinb(n11144), .dina(n2835), .dout(n3615));
    jor g0871(.dinb(n562), .dina(n11427), .dout(n3619));
    jand g0872(.dinb(n10962), .dina(n2017), .dout(n3623));
    jnot g0873(.din(n3623), .dout(n3626));
    jand g0874(.dinb(n3619), .dina(n10956), .dout(n3630));
    jand g0875(.dinb(n3615), .dina(n10950), .dout(n3634));
    jand g0876(.dinb(n11660), .dina(n2843), .dout(n3638));
    jnot g0877(.din(n3638), .dout(n3641));
    jor g0878(.dinb(n604), .dina(n11427), .dout(n3645));
    jand g0879(.dinb(n10812), .dina(n2017), .dout(n3649));
    jnot g0880(.din(n3649), .dout(n3652));
    jand g0881(.dinb(n3645), .dina(n10806), .dout(n3656));
    jand g0882(.dinb(n3641), .dina(n10800), .dout(n3660));
    jnot g0883(.din(n2677), .dout(n3663));
    jand g0884(.dinb(G245), .dina(G559), .dout(n3667));
    jand g0885(.dinb(n360), .dina(n3667), .dout(n3671));
    jand g0886(.dinb(n9977), .dina(n3671), .dout(n3675));
    jand g0887(.dinb(n1665), .dina(n9975), .dout(n3679));
    jand g0888(.dinb(n9983), .dina(n3679), .dout(n3683));
    jand g0889(.dinb(n2626), .dina(n9972), .dout(n3687));
    jand g0890(.dinb(n9966), .dina(n3687), .dout(n3691));
    jand g0891(.dinb(n11894), .dina(n2726), .dout(n3695));
    jnot g0892(.din(n1152), .dout(n3698));
    jand g0893(.dinb(n3698), .dina(n11759), .dout(n3702));
    jand g0894(.dinb(n11754), .dina(n2017), .dout(n3706));
    jor g0895(.dinb(n3702), .dina(n11748), .dout(n3710));
    jor g0896(.dinb(n3695), .dina(n11736), .dout(n3714));
    jnot g0897(.din(n3714), .dout(n3717));
    jand g0898(.dinb(n11885), .dina(n2743), .dout(n3721));
    jor g0899(.dinb(n1240), .dina(n11427), .dout(n3725));
    jand g0900(.dinb(n11421), .dina(n2017), .dout(n3729));
    jnot g0901(.din(n3729), .dout(n3732));
    jand g0902(.dinb(n3725), .dina(n11415), .dout(n3736));
    jnot g0903(.din(n3736), .dout(n3739));
    jor g0904(.dinb(n3721), .dina(n11409), .dout(n3743));
    jnot g0905(.din(n3743), .dout(n3746));
    jor g0906(.dinb(n11105), .dina(n2768), .dout(n3750));
    jor g0907(.dinb(n1110), .dina(n11427), .dout(n3754));
    jand g0908(.dinb(n11040), .dina(n2017), .dout(n3758));
    jnot g0909(.din(n3758), .dout(n3761));
    jand g0910(.dinb(n3754), .dina(n11034), .dout(n3765));
    jand g0911(.dinb(n3750), .dina(n11028), .dout(n3769));
    jand g0912(.dinb(n11906), .dina(n2772), .dout(n3773));
    jnot g0913(.din(n3773), .dout(n3776));
    jor g0914(.dinb(n1198), .dina(n11427), .dout(n3780));
    jand g0915(.dinb(n10854), .dina(n2017), .dout(n3784));
    jnot g0916(.din(n3784), .dout(n3787));
    jand g0917(.dinb(n3780), .dina(n10848), .dout(n3791));
    jand g0918(.dinb(n3776), .dina(n10842), .dout(n3795));
    jand g0919(.dinb(n10421), .dina(n3714), .dout(n3799));
    jand g0920(.dinb(n10418), .dina(n3585), .dout(n3803));
    jand g0921(.dinb(n10140), .dina(n2364), .dout(n3807));
    jand g0922(.dinb(n10134), .dina(n2372), .dout(n3811));
    jor g0923(.dinb(n3807), .dina(n10077), .dout(n3815));
    jor g0924(.dinb(n3803), .dina(n10074), .dout(n3819));
    jor g0925(.dinb(n3799), .dina(n3819), .dout(n3823));
    jand g0926(.dinb(n10247), .dina(n3714), .dout(n3827));
    jand g0927(.dinb(n10244), .dina(n3585), .dout(n3831));
    jand g0928(.dinb(n10140), .dina(n2186), .dout(n3835));
    jand g0929(.dinb(n10134), .dina(n2194), .dout(n3839));
    jor g0930(.dinb(n3835), .dina(n10131), .dout(n3843));
    jor g0931(.dinb(n3831), .dina(n10128), .dout(n3847));
    jor g0932(.dinb(n3827), .dina(n3847), .dout(n3851));
    jand g0933(.dinb(n12338), .dina(n3743), .dout(n3855));
    jnot g0934(.din(n3611), .dout(n3858));
    jand g0935(.dinb(n12212), .dina(n3858), .dout(n3862));
    jand g0936(.dinb(n10356), .dina(n2186), .dout(n3866));
    jand g0937(.dinb(n10350), .dina(n2194), .dout(n3870));
    jor g0938(.dinb(n3866), .dina(n10191), .dout(n3874));
    jor g0939(.dinb(n3862), .dina(n10188), .dout(n3878));
    jor g0940(.dinb(n3855), .dina(n3878), .dout(n3882));
    jnot g0941(.din(n3769), .dout(n3885));
    jand g0942(.dinb(n12338), .dina(n3885), .dout(n3889));
    jnot g0943(.din(n3634), .dout(n3892));
    jand g0944(.dinb(n12212), .dina(n3892), .dout(n3896));
    jand g0945(.dinb(n10416), .dina(n2186), .dout(n3900));
    jand g0946(.dinb(n10410), .dina(n2194), .dout(n3904));
    jor g0947(.dinb(n3900), .dina(n10242), .dout(n3908));
    jor g0948(.dinb(n3896), .dina(n10239), .dout(n3912));
    jor g0949(.dinb(n3889), .dina(n3912), .dout(n3916));
    jnot g0950(.din(n3795), .dout(n3919));
    jand g0951(.dinb(n12308), .dina(n3919), .dout(n3923));
    jnot g0952(.din(n3660), .dout(n3926));
    jand g0953(.dinb(n12182), .dina(n3926), .dout(n3930));
    jand g0954(.dinb(n10479), .dina(n2186), .dout(n3934));
    jand g0955(.dinb(n10473), .dina(n2194), .dout(n3938));
    jor g0956(.dinb(n3934), .dina(n10296), .dout(n3942));
    jor g0957(.dinb(n3930), .dina(n10293), .dout(n3946));
    jor g0958(.dinb(n3923), .dina(n3946), .dout(n3950));
    jand g0959(.dinb(n12677), .dina(n3743), .dout(n3954));
    jand g0960(.dinb(n12551), .dina(n3858), .dout(n3958));
    jand g0961(.dinb(n10356), .dina(n2364), .dout(n3962));
    jand g0962(.dinb(n10350), .dina(n2372), .dout(n3966));
    jor g0963(.dinb(n3962), .dina(n10347), .dout(n3970));
    jor g0964(.dinb(n3958), .dina(n10344), .dout(n3974));
    jor g0965(.dinb(n3954), .dina(n3974), .dout(n3978));
    jand g0966(.dinb(n12677), .dina(n3885), .dout(n3982));
    jand g0967(.dinb(n12551), .dina(n3892), .dout(n3986));
    jand g0968(.dinb(n10416), .dina(n2364), .dout(n3990));
    jand g0969(.dinb(n10410), .dina(n2372), .dout(n3994));
    jor g0970(.dinb(n3990), .dina(n10407), .dout(n3998));
    jor g0971(.dinb(n3986), .dina(n10404), .dout(n4002));
    jor g0972(.dinb(n3982), .dina(n4002), .dout(n4006));
    jand g0973(.dinb(n12647), .dina(n3919), .dout(n4010));
    jand g0974(.dinb(n12521), .dina(n3926), .dout(n4014));
    jand g0975(.dinb(n10479), .dina(n2364), .dout(n4018));
    jand g0976(.dinb(n10473), .dina(n2372), .dout(n4022));
    jor g0977(.dinb(n4018), .dina(n10470), .dout(n4026));
    jor g0978(.dinb(n4014), .dina(n10467), .dout(n4030));
    jor g0979(.dinb(n4010), .dina(n4030), .dout(n4034));
    jand g0980(.dinb(n13142), .dina(n3919), .dout(n4038));
    jand g0981(.dinb(n12938), .dina(n3926), .dout(n4042));
    jand g0982(.dinb(n10773), .dina(n2908), .dout(n4046));
    jand g0983(.dinb(n10767), .dina(n2916), .dout(n4050));
    jor g0984(.dinb(n4046), .dina(n10527), .dout(n4054));
    jor g0985(.dinb(n4042), .dina(n10524), .dout(n4058));
    jor g0986(.dinb(n4038), .dina(n4058), .dout(n4062));
    jand g0987(.dinb(n10529), .dina(n4062), .dout(n4066));
    jand g0988(.dinb(n10658), .dina(n3885), .dout(n4070));
    jand g0989(.dinb(n10652), .dina(n3892), .dout(n4074));
    jand g0990(.dinb(n10920), .dina(n2908), .dout(n4078));
    jand g0991(.dinb(n10914), .dina(n2916), .dout(n4082));
    jor g0992(.dinb(n4078), .dina(n10596), .dout(n4086));
    jor g0993(.dinb(n4074), .dina(n10593), .dout(n4090));
    jor g0994(.dinb(n4070), .dina(n4090), .dout(n4094));
    jand g0995(.dinb(n11468), .dina(n4094), .dout(n4098));
    jand g0996(.dinb(n10655), .dina(n3743), .dout(n4102));
    jand g0997(.dinb(n10649), .dina(n3858), .dout(n4106));
    jand g0998(.dinb(n11238), .dina(n2908), .dout(n4110));
    jand g0999(.dinb(n11232), .dina(n2916), .dout(n4114));
    jor g1000(.dinb(n4110), .dina(n10647), .dout(n4118));
    jor g1001(.dinb(n4106), .dina(n10644), .dout(n4122));
    jor g1002(.dinb(n4102), .dina(n4122), .dout(n4126));
    jand g1003(.dinb(n11468), .dina(n4126), .dout(n4130));
    jand g1004(.dinb(n13085), .dina(n3714), .dout(n4134));
    jand g1005(.dinb(n12884), .dina(n3585), .dout(n4138));
    jand g1006(.dinb(n11547), .dina(n2908), .dout(n4142));
    jand g1007(.dinb(n11541), .dina(n2916), .dout(n4146));
    jor g1008(.dinb(n4142), .dina(n10713), .dout(n4150));
    jor g1009(.dinb(n4138), .dina(n10710), .dout(n4154));
    jor g1010(.dinb(n4134), .dina(n4154), .dout(n4158));
    jand g1011(.dinb(n10715), .dina(n4158), .dout(n4162));
    jand g1012(.dinb(n16400), .dina(n3919), .dout(n4166));
    jand g1013(.dinb(n14783), .dina(n3926), .dout(n4170));
    jand g1014(.dinb(n10773), .dina(n2962), .dout(n4174));
    jand g1015(.dinb(n10767), .dina(n2970), .dout(n4178));
    jor g1016(.dinb(n4174), .dina(n10764), .dout(n4182));
    jor g1017(.dinb(n4170), .dina(n10761), .dout(n4186));
    jor g1018(.dinb(n4166), .dina(n4186), .dout(n4190));
    jand g1019(.dinb(n11453), .dina(n4190), .dout(n4194));
    jand g1020(.dinb(n11444), .dina(n3885), .dout(n4198));
    jand g1021(.dinb(n11375), .dina(n3892), .dout(n4202));
    jand g1022(.dinb(n10920), .dina(n2962), .dout(n4206));
    jand g1023(.dinb(n10914), .dina(n2970), .dout(n4210));
    jor g1024(.dinb(n4206), .dina(n10911), .dout(n4214));
    jor g1025(.dinb(n4202), .dina(n10908), .dout(n4218));
    jor g1026(.dinb(n4198), .dina(n4218), .dout(n4222));
    jand g1027(.dinb(n11450), .dina(n4222), .dout(n4226));
    jand g1028(.dinb(n11441), .dina(n3743), .dout(n4230));
    jand g1029(.dinb(n11372), .dina(n3858), .dout(n4234));
    jand g1030(.dinb(n11238), .dina(n2962), .dout(n4238));
    jand g1031(.dinb(n11232), .dina(n2970), .dout(n4242));
    jor g1032(.dinb(n4238), .dina(n11229), .dout(n4246));
    jor g1033(.dinb(n4234), .dina(n11226), .dout(n4250));
    jor g1034(.dinb(n4230), .dina(n4250), .dout(n4254));
    jand g1035(.dinb(n11447), .dina(n4254), .dout(n4258));
    jand g1036(.dinb(n16343), .dina(n3714), .dout(n4262));
    jand g1037(.dinb(n14729), .dina(n3585), .dout(n4266));
    jand g1038(.dinb(n11547), .dina(n2962), .dout(n4270));
    jand g1039(.dinb(n11541), .dina(n2970), .dout(n4274));
    jor g1040(.dinb(n4270), .dina(n11538), .dout(n4278));
    jor g1041(.dinb(n4266), .dina(n11535), .dout(n4282));
    jor g1042(.dinb(n4262), .dina(n4282), .dout(n4286));
    jand g1043(.dinb(n16562), .dina(n4286), .dout(n4290));
    jor g1044(.dinb(G120), .dina(G4091), .dout(n4294));
    jand g1045(.dinb(n16277), .dina(n795), .dout(n4298));
    jand g1046(.dinb(G248), .dina(G341), .dout(n4302));
    jor g1047(.dinb(n802), .dina(n4302), .dout(n4306));
    jor g1048(.dinb(n4298), .dina(n4306), .dout(n4310));
    jand g1049(.dinb(n539), .dina(n795), .dout(n4314));
    jand g1050(.dinb(n546), .dina(n14675), .dout(n4318));
    jor g1051(.dinb(n14666), .dina(n4318), .dout(n4322));
    jor g1052(.dinb(n14643), .dina(n4322), .dout(n4326));
    jand g1053(.dinb(n14640), .dina(n4326), .dout(n4330));
    jxor g1054(.dinb(n14630), .dina(n695), .dout(n4334));
    jxor g1055(.dinb(n562), .dina(n604), .dout(n4338));
    jxor g1056(.dinb(n14538), .dina(n4338), .dout(n4342));
    jxor g1057(.dinb(n14535), .dina(n4342), .dout(n4346));
    jnot g1058(.din(n4346), .dout(n4349));
    jor g1059(.dinb(n16223), .dina(n702), .dout(n4353));
    jor g1060(.dinb(n546), .dina(n14519), .dout(n4357));
    jand g1061(.dinb(n4353), .dina(n4357), .dout(n4361));
    jxor g1062(.dinb(n735), .dina(n4361), .dout(n4365));
    jor g1063(.dinb(n674), .dina(n14513), .dout(n4369));
    jor g1064(.dinb(n684), .dina(n611), .dout(n4373));
    jand g1065(.dinb(n14498), .dina(n4373), .dout(n4377));
    jand g1066(.dinb(n14493), .dina(n4377), .dout(n4381));
    jor g1067(.dinb(G254), .dina(G351), .dout(n4385));
    jor g1068(.dinb(n16214), .dina(n611), .dout(n4389));
    jand g1069(.dinb(n14478), .dina(n4389), .dout(n4393));
    jand g1070(.dinb(n14472), .dina(n4393), .dout(n4397));
    jor g1071(.dinb(n4381), .dina(n4397), .dout(n4401));
    jand g1072(.dinb(n16277), .dina(n753), .dout(n4405));
    jand g1073(.dinb(G248), .dina(G324), .dout(n4409));
    jor g1074(.dinb(n760), .dina(n4409), .dout(n4413));
    jor g1075(.dinb(n4405), .dina(n4413), .dout(n4417));
    jand g1076(.dinb(n539), .dina(n753), .dout(n4421));
    jand g1077(.dinb(n546), .dina(n14465), .dout(n4425));
    jor g1078(.dinb(n14444), .dina(n4425), .dout(n4429));
    jor g1079(.dinb(n14424), .dina(n4429), .dout(n4433));
    jand g1080(.dinb(n14421), .dina(n4433), .dout(n4437));
    jxor g1081(.dinb(n4401), .dina(n4437), .dout(n4441));
    jxor g1082(.dinb(n14418), .dina(n4441), .dout(n4445));
    jnot g1083(.din(n4445), .dout(n4448));
    jand g1084(.dinb(n4349), .dina(n14408), .dout(n4452));
    jor g1085(.dinb(n14378), .dina(n4452), .dout(n4456));
    jor g1086(.dinb(n1991), .dina(n4294), .dout(n4460));
    jand g1087(.dinb(n4346), .dina(n4448), .dout(n4464));
    jor g1088(.dinb(n14322), .dina(n4456), .dout(n4468));
    jand g1089(.dinb(n14678), .dina(n4468), .dout(n4472));
    jnot g1090(.din(n4472), .dout(n4475));
    jand g1091(.dinb(n14120), .dina(n1555), .dout(n4479));
    jor g1092(.dinb(n1940), .dina(n14049), .dout(n4483));
    jand g1093(.dinb(n14000), .dina(n1954), .dout(n4487));
    jor g1094(.dinb(n1585), .dina(n1969), .dout(n4491));
    jand g1095(.dinb(n13988), .dina(n4491), .dout(n4495));
    jor g1096(.dinb(n13899), .dina(n4495), .dout(n4499));
    jnot g1097(.din(n4499), .dout(n4502));
    jand g1098(.dinb(n13931), .dina(n4502), .dout(n4506));
    jnot g1099(.din(n1965), .dout(n4509));
    jand g1100(.dinb(n13836), .dina(n4499), .dout(n4513));
    jor g1101(.dinb(n13838), .dina(n4513), .dout(n4517));
    jor g1102(.dinb(n4506), .dina(n4517), .dout(n4521));
    jand g1103(.dinb(n4483), .dina(n13827), .dout(n4525));
    jnot g1104(.din(n4483), .dout(n4528));
    jxor g1105(.dinb(n13821), .dina(n4502), .dout(n4532));
    jand g1106(.dinb(n4528), .dina(n13791), .dout(n4536));
    jor g1107(.dinb(n13779), .dina(n4536), .dout(n4540));
    jnot g1108(.din(n4540), .dout(n4543));
    jxor g1109(.dinb(n14075), .dina(n1540), .dout(n4547));
    jnot g1110(.din(n4547), .dout(n4550));
    jxor g1111(.dinb(n13646), .dina(n2214), .dout(n4554));
    jnot g1112(.din(n1481), .dout(n4557));
    jnot g1113(.din(n1881), .dout(n4560));
    jand g1114(.dinb(n2299), .dina(n1512), .dout(n4564));
    jand g1115(.dinb(n14657), .dina(n1536), .dout(n4568));
    jor g1116(.dinb(n2303), .dina(n4568), .dout(n4572));
    jor g1117(.dinb(n4564), .dina(n4572), .dout(n4576));
    jand g1118(.dinb(n13608), .dina(n4576), .dout(n4580));
    jxor g1119(.dinb(n1497), .dina(n1512), .dout(n4584));
    jnot g1120(.din(n4584), .dout(n4587));
    jor g1121(.dinb(n4580), .dina(n13596), .dout(n4591));
    jor g1122(.dinb(n2264), .dina(n13598), .dout(n4595));
    jand g1123(.dinb(n13593), .dina(n4595), .dout(n4599));
    jxor g1124(.dinb(n13590), .dina(n4599), .dout(n4603));
    jand g1125(.dinb(n4554), .dina(n4603), .dout(n4607));
    jnot g1126(.din(G2174), .dout(n4610));
    jxor g1127(.dinb(n14195), .dina(n2214), .dout(n4614));
    jxor g1128(.dinb(n13613), .dina(n4599), .dout(n4618));
    jand g1129(.dinb(n4614), .dina(n4618), .dout(n4622));
    jor g1130(.dinb(n13578), .dina(n4622), .dout(n4626));
    jor g1131(.dinb(n13545), .dina(n4626), .dout(n4630));
    jxor g1132(.dinb(n14273), .dina(n1929), .dout(n4634));
    jnot g1133(.din(n4634), .dout(n4637));
    jor g1134(.dinb(n1897), .dina(n1512), .dout(n4641));
    jand g1135(.dinb(n14189), .dina(n4641), .dout(n4645));
    jxor g1136(.dinb(n1921), .dina(n13542), .dout(n4649));
    jand g1137(.dinb(n4637), .dina(n13532), .dout(n4653));
    jnot g1138(.din(n4649), .dout(n4656));
    jand g1139(.dinb(n4634), .dina(n13530), .dout(n4660));
    jor g1140(.dinb(n14087), .dina(n4660), .dout(n4664));
    jor g1141(.dinb(n4653), .dina(n4664), .dout(n4668));
    jand g1142(.dinb(n4630), .dina(n13527), .dout(n4672));
    jxor g1143(.dinb(n13695), .dina(n4672), .dout(n4676));
    jxor g1144(.dinb(n13524), .dina(n4676), .dout(n4680));
    jor g1145(.dinb(n4543), .dina(n4680), .dout(n4684));
    jxor g1146(.dinb(n13742), .dina(n4676), .dout(n4688));
    jor g1147(.dinb(n13775), .dina(n4688), .dout(n4692));
    jand g1148(.dinb(n14324), .dina(n4692), .dout(n4696));
    jand g1149(.dinb(n13493), .dina(n4696), .dout(n4700));
    jor g1150(.dinb(n13491), .dina(n4700), .dout(n4704));
    jand g1151(.dinb(n12021), .dina(n4704), .dout(n4708));
    jor g1152(.dinb(G118), .dina(G4091), .dout(n4712));
    jand g1153(.dinb(n891), .dina(n16274), .dout(n4716));
    jand g1154(.dinb(G234), .dina(G248), .dout(n4720));
    jor g1155(.dinb(n898), .dina(n4720), .dout(n4724));
    jor g1156(.dinb(n4716), .dina(n4724), .dout(n4728));
    jand g1157(.dinb(n891), .dina(n539), .dout(n4732));
    jand g1158(.dinb(n16283), .dina(n546), .dout(n4736));
    jor g1159(.dinb(n16256), .dina(n4736), .dout(n4740));
    jor g1160(.dinb(n16209), .dina(n4740), .dout(n4744));
    jand g1161(.dinb(n16206), .dina(n4744), .dout(n4748));
    jor g1162(.dinb(n16151), .dina(n674), .dout(n4752));
    jor g1163(.dinb(n1159), .dina(n684), .dout(n4756));
    jand g1164(.dinb(n16133), .dina(n4756), .dout(n4760));
    jand g1165(.dinb(n16119), .dina(n4760), .dout(n4764));
    jor g1166(.dinb(G226), .dina(G254), .dout(n4768));
    jor g1167(.dinb(n1159), .dina(n16211), .dout(n4772));
    jand g1168(.dinb(n16113), .dina(n4772), .dout(n4776));
    jand g1169(.dinb(n16110), .dina(n4776), .dout(n4780));
    jor g1170(.dinb(n4764), .dina(n4780), .dout(n4784));
    jxor g1171(.dinb(n1152), .dina(n4784), .dout(n4788));
    jor g1172(.dinb(n16103), .dina(n674), .dout(n4792));
    jor g1173(.dinb(n1071), .dina(n684), .dout(n4796));
    jand g1174(.dinb(n16088), .dina(n4796), .dout(n4800));
    jand g1175(.dinb(n16083), .dina(n4800), .dout(n4804));
    jor g1176(.dinb(G218), .dina(G254), .dout(n4808));
    jor g1177(.dinb(n1071), .dina(n16220), .dout(n4812));
    jand g1178(.dinb(n16068), .dina(n4812), .dout(n4816));
    jand g1179(.dinb(n16065), .dina(n4816), .dout(n4820));
    jor g1180(.dinb(n4804), .dina(n4820), .dout(n4824));
    jand g1181(.dinb(n1201), .dina(n16274), .dout(n4828));
    jand g1182(.dinb(G210), .dina(G248), .dout(n4832));
    jor g1183(.dinb(n1208), .dina(n4832), .dout(n4836));
    jor g1184(.dinb(n4828), .dina(n4836), .dout(n4840));
    jand g1185(.dinb(n1201), .dina(n539), .dout(n4844));
    jand g1186(.dinb(n16058), .dina(n546), .dout(n4848));
    jor g1187(.dinb(n16049), .dina(n4848), .dout(n4852));
    jor g1188(.dinb(n16029), .dina(n4852), .dout(n4856));
    jand g1189(.dinb(n16026), .dina(n4856), .dout(n4860));
    jxor g1190(.dinb(n4824), .dina(n4860), .dout(n4864));
    jxor g1191(.dinb(n4788), .dina(n4864), .dout(n4868));
    jxor g1192(.dinb(n16023), .dina(n4868), .dout(n4872));
    jand g1193(.dinb(n16274), .dina(n1025), .dout(n4876));
    jand g1194(.dinb(G248), .dina(G281), .dout(n4880));
    jor g1195(.dinb(n1032), .dina(n4880), .dout(n4884));
    jor g1196(.dinb(n4876), .dina(n4884), .dout(n4888));
    jand g1197(.dinb(n539), .dina(n1025), .dout(n4892));
    jand g1198(.dinb(n546), .dina(n16016), .dout(n4896));
    jor g1199(.dinb(n16004), .dina(n4896), .dout(n4900));
    jor g1200(.dinb(n15993), .dina(n4900), .dout(n4904));
    jand g1201(.dinb(n15990), .dina(n4904), .dout(n4908));
    jand g1202(.dinb(n16148), .dina(n849), .dout(n4912));
    jand g1203(.dinb(G248), .dina(G265), .dout(n4916));
    jor g1204(.dinb(n856), .dina(n4916), .dout(n4920));
    jor g1205(.dinb(n4912), .dina(n4920), .dout(n4924));
    jand g1206(.dinb(n539), .dina(n849), .dout(n4928));
    jand g1207(.dinb(n546), .dina(n15986), .dout(n4932));
    jor g1208(.dinb(n15968), .dina(n4932), .dout(n4936));
    jor g1209(.dinb(n15954), .dina(n4936), .dout(n4940));
    jand g1210(.dinb(n15951), .dina(n4940), .dout(n4944));
    jxor g1211(.dinb(n4908), .dina(n4944), .dout(n4948));
    jor g1212(.dinb(n674), .dina(n15947), .dout(n4952));
    jor g1213(.dinb(n684), .dina(n933), .dout(n4956));
    jand g1214(.dinb(n15938), .dina(n4956), .dout(n4960));
    jand g1215(.dinb(n15933), .dina(n4960), .dout(n4964));
    jor g1216(.dinb(G254), .dina(G257), .dout(n4968));
    jor g1217(.dinb(n16217), .dina(n933), .dout(n4972));
    jand g1218(.dinb(n15930), .dina(n4972), .dout(n4976));
    jand g1219(.dinb(n15921), .dina(n4976), .dout(n4980));
    jor g1220(.dinb(n4964), .dina(n4980), .dout(n4984));
    jand g1221(.dinb(n16145), .dina(n983), .dout(n4988));
    jand g1222(.dinb(G248), .dina(G273), .dout(n4992));
    jor g1223(.dinb(n990), .dina(n4992), .dout(n4996));
    jor g1224(.dinb(n4988), .dina(n4996), .dout(n5000));
    jand g1225(.dinb(n539), .dina(n983), .dout(n5004));
    jand g1226(.dinb(n546), .dina(n15914), .dout(n5008));
    jor g1227(.dinb(n15902), .dina(n5008), .dout(n5012));
    jor g1228(.dinb(n15891), .dina(n5012), .dout(n5016));
    jand g1229(.dinb(n15888), .dina(n5016), .dout(n5020));
    jxor g1230(.dinb(n4984), .dina(n5020), .dout(n5024));
    jxor g1231(.dinb(n4948), .dina(n5024), .dout(n5028));
    jand g1232(.dinb(n4872), .dina(n15885), .dout(n5032));
    jnot g1233(.din(n5032), .dout(n5035));
    jor g1234(.dinb(n4872), .dina(n15885), .dout(n5039));
    jand g1235(.dinb(n15803), .dina(n5039), .dout(n5043));
    jand g1236(.dinb(n5035), .dina(n5043), .dout(n5047));
    jor g1237(.dinb(n1991), .dina(n4712), .dout(n5051));
    jor g1238(.dinb(n16286), .dina(n5047), .dout(n5055));
    jxor g1239(.dinb(n1342), .dina(n1361), .dout(n5059));
    jxor g1240(.dinb(n2732), .dina(n5059), .dout(n5063));
    jnot g1241(.din(n5063), .dout(n5066));
    jand g1242(.dinb(n15479), .dina(n1376), .dout(n5070));
    jor g1243(.dinb(n1797), .dina(n15363), .dout(n5074));
    jnot g1244(.din(n5074), .dout(n5077));
    jor g1245(.dinb(n15267), .dina(n2735), .dout(n5081));
    jand g1246(.dinb(n15278), .dina(n5081), .dout(n5085));
    jxor g1247(.dinb(n15339), .dina(n5085), .dout(n5089));
    jxor g1248(.dinb(n2750), .dina(n1447), .dout(n5093));
    jxor g1249(.dinb(n5089), .dina(n15171), .dout(n5097));
    jand g1250(.dinb(n5077), .dina(n15156), .dout(n5101));
    jxor g1251(.dinb(n1825), .dina(n1447), .dout(n5105));
    jand g1252(.dinb(n2750), .dina(n1447), .dout(n5109));
    jor g1253(.dinb(n15294), .dina(n5109), .dout(n5113));
    jnot g1254(.din(n5113), .dout(n5116));
    jor g1255(.dinb(n15267), .dina(n5116), .dout(n5120));
    jor g1256(.dinb(n1841), .dina(n15125), .dout(n5124));
    jand g1257(.dinb(n15123), .dina(n5124), .dout(n5128));
    jxor g1258(.dinb(n15341), .dina(n5128), .dout(n5132));
    jand g1259(.dinb(n15147), .dina(n5132), .dout(n5136));
    jnot g1260(.din(n5136), .dout(n5139));
    jor g1261(.dinb(n15147), .dina(n5132), .dout(n5143));
    jand g1262(.dinb(n5074), .dina(n15120), .dout(n5147));
    jand g1263(.dinb(n15117), .dina(n5147), .dout(n5151));
    jor g1264(.dinb(n5101), .dina(n5151), .dout(n5155));
    jnot g1265(.din(G1497), .dout(n5158));
    jand g1266(.dinb(n15542), .dina(n1744), .dout(n5162));
    jand g1267(.dinb(n1326), .dina(n15113), .dout(n5166));
    jxor g1268(.dinb(n15434), .dina(n5166), .dout(n5170));
    jxor g1269(.dinb(n15110), .dina(n1319), .dout(n5174));
    jor g1270(.dinb(n15096), .dina(n2405), .dout(n5178));
    jand g1271(.dinb(n15365), .dina(n1786), .dout(n5182));
    jor g1272(.dinb(n15080), .dina(n5182), .dout(n5186));
    jand g1273(.dinb(n5178), .dina(n5186), .dout(n5190));
    jxor g1274(.dinb(n15078), .dina(n5190), .dout(n5194));
    jxor g1275(.dinb(n15060), .dina(n5194), .dout(n5198));
    jor g1276(.dinb(n15048), .dina(n5198), .dout(n5202));
    jxor g1277(.dinb(n15383), .dina(n1786), .dout(n5206));
    jor g1278(.dinb(n15098), .dina(n2408), .dout(n5210));
    jnot g1279(.din(n1740), .dout(n5213));
    jor g1280(.dinb(n5213), .dina(n15585), .dout(n5217));
    jor g1281(.dinb(n15539), .dina(n5217), .dout(n5221));
    jxor g1282(.dinb(n15398), .dina(n5221), .dout(n5225));
    jand g1283(.dinb(n5210), .dina(n15009), .dout(n5229));
    jxor g1284(.dinb(n15431), .dina(n5162), .dout(n5233));
    jxor g1285(.dinb(n5229), .dina(n15006), .dout(n5237));
    jxor g1286(.dinb(n14997), .dina(n5237), .dout(n5241));
    jor g1287(.dinb(n15443), .dina(n5241), .dout(n5245));
    jand g1288(.dinb(n5202), .dina(n14994), .dout(n5249));
    jxor g1289(.dinb(n5155), .dina(n5249), .dout(n5253));
    jand g1290(.dinb(n15639), .dina(n5253), .dout(n5257));
    jnot g1291(.din(n5257), .dout(n5260));
    jor g1292(.dinb(n15639), .dina(n5253), .dout(n5264));
    jand g1293(.dinb(n15830), .dina(n5264), .dout(n5268));
    jand g1294(.dinb(n5260), .dina(n5268), .dout(n5272));
    jor g1295(.dinb(n14988), .dina(n5272), .dout(n5276));
    jand g1296(.dinb(n12078), .dina(n5276), .dout(n5280));
    jand g1297(.dinb(G97), .dina(G4092), .dout(n5284));
    jnot g1298(.din(n5284), .dout(n5287));
    jand g1299(.dinb(n5276), .dina(n14964), .dout(n5291));
    jnot g1300(.din(n5291), .dout(n5294));
    jand g1301(.dinb(n12266), .dina(n5294), .dout(n5298));
    jnot g1302(.din(n4684), .dout(n5301));
    jand g1303(.dinb(n4543), .dina(n4680), .dout(n5305));
    jor g1304(.dinb(n15752), .dina(n5305), .dout(n5309));
    jor g1305(.dinb(n5301), .dina(n5309), .dout(n5313));
    jand g1306(.dinb(n14297), .dina(n5313), .dout(n5317));
    jand g1307(.dinb(G94), .dina(G4092), .dout(n5321));
    jor g1308(.dinb(n5317), .dina(n13415), .dout(n5325));
    jand g1309(.dinb(n12140), .dina(n5325), .dout(n5329));
    jand g1310(.dinb(n12477), .dina(n2186), .dout(n5333));
    jand g1311(.dinb(n12471), .dina(n2194), .dout(n5337));
    jor g1312(.dinb(n5333), .dina(n12138), .dout(n5341));
    jor g1313(.dinb(n5329), .dina(n12135), .dout(n5345));
    jor g1314(.dinb(n5298), .dina(n5345), .dout(n5349));
    jand g1315(.dinb(n12605), .dina(n5294), .dout(n5353));
    jand g1316(.dinb(n12479), .dina(n5325), .dout(n5357));
    jand g1317(.dinb(n12477), .dina(n2364), .dout(n5361));
    jand g1318(.dinb(n12471), .dina(n2372), .dout(n5365));
    jor g1319(.dinb(n5361), .dina(n12468), .dout(n5369));
    jor g1320(.dinb(n5357), .dina(n12465), .dout(n5373));
    jor g1321(.dinb(n5353), .dina(n5373), .dout(n5377));
    jnot g1322(.din(G137), .dout(n5380));
    jnot g1323(.din(n2889), .dout(n5383));
    jor g1324(.dinb(n13062), .dina(n5291), .dout(n5387));
    jnot g1325(.din(n2900), .dout(n5390));
    jnot g1326(.din(n5321), .dout(n5393));
    jand g1327(.dinb(n4704), .dina(n13413), .dout(n5397));
    jor g1328(.dinb(n12864), .dina(n5397), .dout(n5401));
    jnot g1329(.din(G179), .dout(n5404));
    jnot g1330(.din(n2916), .dout(n5407));
    jor g1331(.dinb(n13299), .dina(n5407), .dout(n5411));
    jnot g1332(.din(G176), .dout(n5414));
    jnot g1333(.din(n2908), .dout(n5417));
    jor g1334(.dinb(n13296), .dina(n5417), .dout(n5421));
    jand g1335(.dinb(n12807), .dina(n5421), .dout(n5425));
    jand g1336(.dinb(n5401), .dina(n12804), .dout(n5429));
    jand g1337(.dinb(n12750), .dina(n5429), .dout(n5433));
    jor g1338(.dinb(n16560), .dina(n5433), .dout(G658));
    jnot g1339(.din(n2943), .dout(n5440));
    jor g1340(.dinb(n14907), .dina(n5291), .dout(n5444));
    jnot g1341(.din(n2954), .dout(n5447));
    jor g1342(.dinb(n13356), .dina(n5397), .dout(n5451));
    jnot g1343(.din(n2970), .dout(n5454));
    jor g1344(.dinb(n13299), .dina(n5454), .dout(n5458));
    jnot g1345(.din(n2962), .dout(n5461));
    jor g1346(.dinb(n13296), .dina(n5461), .dout(n5465));
    jand g1347(.dinb(n13290), .dina(n5465), .dout(n5469));
    jand g1348(.dinb(n5451), .dina(n13287), .dout(n5473));
    jand g1349(.dinb(n13233), .dina(n5473), .dout(n5477));
    jor g1350(.dinb(n16560), .dina(n5477), .dout(G690));
    jdff g1351(.din(G141), .dout(n5484));
    jdff g1352(.din(G293), .dout(n5487));
    jdff g1353(.din(G3173), .dout(n5490));
    jnot g1354(.din(G545), .dout(n5493));
    jnot g1355(.din(G545), .dout(n5496));
    jdff g1356(.din(G137), .dout(n5499));
    jdff g1357(.din(G141), .dout(n5502));
    jdff g1358(.din(G1), .dout(n5505));
    jdff g1359(.din(G549), .dout(n5508));
    jdff g1360(.din(G299), .dout(n5511));
    jnot g1361(.din(G549), .dout(n5514));
    jdff g1362(.din(G1), .dout(n5517));
    jdff g1363(.din(G1), .dout(n5520));
    jdff g1364(.din(G1), .dout(n5523));
    jdff g1365(.din(G1), .dout(n5526));
    jdff g1366(.din(G299), .dout(n5529));
    jor g1367(.dinb(n8028), .dina(n423), .dout(n5533));
    jand g1368(.dinb(n1555), .dina(n8139), .dout(n5537));
    jand g1369(.dinb(n1376), .dina(n8184), .dout(n5541));
    jor g1370(.dinb(n1801), .dina(n8148), .dout(n5545));
    jor g1371(.dinb(n1944), .dina(n8202), .dout(n5549));
    jdff dff_A_1hgo6KA25_2(.din(n5377), .dout(G807));
    jdff dff_A_jKaG1UkO8_2(.din(n5349), .dout(G767));
    jdff dff_A_B66RrRug7_0(.din(n22040), .dout(G882));
    jdff dff_A_Gb01iVMQ7_0(.din(n22037), .dout(n22040));
    jdff dff_A_YDRa4Cqv9_0(.din(n22034), .dout(n22037));
    jdff dff_A_uG8smKgl3_2(.din(n5280), .dout(n22034));
    jdff dff_A_pNCoGSMR1_0(.din(n22028), .dout(G843));
    jdff dff_A_IphPcu077_0(.din(n22025), .dout(n22028));
    jdff dff_A_5JQSpGdh3_0(.din(n22022), .dout(n22025));
    jdff dff_A_SURhQcVE9_2(.din(n4708), .dout(n22022));
    jdff dff_A_83ihCwOD9_0(.din(n22016), .dout(G688));
    jdff dff_A_8T6yUygj4_2(.din(n4290), .dout(n22016));
    jdff dff_A_tBzr0fGn3_0(.din(n22010), .dout(G685));
    jdff dff_A_gk80YyZu3_0(.din(n22007), .dout(n22010));
    jdff dff_A_R1XS5Ihe0_2(.din(n4258), .dout(n22007));
    jdff dff_A_gRXC4Tr85_0(.din(n22001), .dout(G682));
    jdff dff_A_uRcD19pB1_0(.din(n21998), .dout(n22001));
    jdff dff_A_pBwC6pVv9_2(.din(n4226), .dout(n21998));
    jdff dff_A_TAD277UN8_0(.din(n21992), .dout(G679));
    jdff dff_A_gmRVeP8O9_0(.din(n21989), .dout(n21992));
    jdff dff_A_2UHCS21P1_0(.din(n21986), .dout(n21989));
    jdff dff_A_Koy1Jatt2_2(.din(n4194), .dout(n21986));
    jdff dff_A_3cv1kEqb2_0(.din(n21980), .dout(G654));
    jdff dff_A_GDUy23aV8_2(.din(n4162), .dout(n21980));
    jdff dff_A_wNH9s7Zb0_0(.din(n21974), .dout(G651));
    jdff dff_A_HJOc8wDx5_0(.din(n21971), .dout(n21974));
    jdff dff_A_yqoRBsWS7_2(.din(n4130), .dout(n21971));
    jdff dff_A_9HeNAnN46_0(.din(n21965), .dout(G648));
    jdff dff_A_0phmmXY59_0(.din(n21962), .dout(n21965));
    jdff dff_A_1QlhlnXk4_2(.din(n4098), .dout(n21962));
    jdff dff_A_R2caKM6X3_0(.din(n21956), .dout(G645));
    jdff dff_A_DlsGPHEV0_0(.din(n21953), .dout(n21956));
    jdff dff_A_oMhcGBxd0_0(.din(n21950), .dout(n21953));
    jdff dff_A_FMg1FwX22_2(.din(n4066), .dout(n21950));
    jdff dff_A_TCsuykfJ9_0(.din(n21944), .dout(G782));
    jdff dff_A_mtX3FGsz2_0(.din(n21941), .dout(n21944));
    jdff dff_A_Uh9DHK8c5_0(.din(n21938), .dout(n21941));
    jdff dff_A_p4Z6OHCa9_0(.din(n21935), .dout(n21938));
    jdff dff_A_W3LY4oTh8_2(.din(n4034), .dout(n21935));
    jdff dff_A_2oSbqiNS6_0(.din(n21929), .dout(G777));
    jdff dff_A_AYIiujB36_0(.din(n21926), .dout(n21929));
    jdff dff_A_USWGTGjs0_0(.din(n21923), .dout(n21926));
    jdff dff_A_Jc6Rpzbn3_2(.din(n4006), .dout(n21923));
    jdff dff_A_4jrRbgWU5_0(.din(n21917), .dout(G772));
    jdff dff_A_YB3NsWiX5_0(.din(n21914), .dout(n21917));
    jdff dff_A_ngOjbvSY8_0(.din(n21911), .dout(n21914));
    jdff dff_A_zLFP5pWE0_2(.din(n3978), .dout(n21911));
    jdff dff_A_EWnvNPoH7_0(.din(n21905), .dout(G742));
    jdff dff_A_u65Zf4pJ9_0(.din(n21902), .dout(n21905));
    jdff dff_A_WO8lGLWg1_0(.din(n21899), .dout(n21902));
    jdff dff_A_sD9RiPX72_0(.din(n21896), .dout(n21899));
    jdff dff_A_PIldz9RX9_2(.din(n3950), .dout(n21896));
    jdff dff_A_nF3iWpjD1_0(.din(n21890), .dout(G737));
    jdff dff_A_AqPdayHI6_0(.din(n21887), .dout(n21890));
    jdff dff_A_tWlDItD29_0(.din(n21884), .dout(n21887));
    jdff dff_A_8UD0c5Ru2_2(.din(n3916), .dout(n21884));
    jdff dff_A_Wh7K7oZ84_0(.din(n21878), .dout(G732));
    jdff dff_A_3mGJs6Ph6_0(.din(n21875), .dout(n21878));
    jdff dff_A_DUQ5RHt73_0(.din(n21872), .dout(n21875));
    jdff dff_A_zT3XBVAo1_2(.din(n3882), .dout(n21872));
    jdff dff_A_vkSUaR3g5_0(.din(n21866), .dout(G727));
    jdff dff_A_DkB9eyZc1_0(.din(n21863), .dout(n21866));
    jdff dff_A_cpxnTtkT7_2(.din(n3851), .dout(n21863));
    jdff dff_A_fWRL19Y44_0(.din(n21857), .dout(G712));
    jdff dff_A_TXy3L1NG6_0(.din(n21854), .dout(n21857));
    jdff dff_A_UTwmXiJV5_2(.din(n3823), .dout(n21854));
    jdff dff_A_rCo1GP2Y6_0(.din(n21848), .dout(G869));
    jdff dff_A_6yUTm2Ws8_0(.din(n21845), .dout(n21848));
    jdff dff_A_NjzqUsoA9_0(.din(n21842), .dout(n21845));
    jdff dff_A_3jeAbU1w5_0(.din(n21839), .dout(n21842));
    jdff dff_A_xdEoz0CS8_0(.din(n21836), .dout(n21839));
    jdff dff_A_1rSdnZCe4_0(.din(n21833), .dout(n21836));
    jdff dff_A_kyD7zK7U1_0(.din(n21830), .dout(n21833));
    jdff dff_A_Y9DXbQ481_1(.din(n3795), .dout(n21830));
    jdff dff_A_2JE9l8j69_0(.din(n21824), .dout(G867));
    jdff dff_A_0s4VnOCC6_0(.din(n21821), .dout(n21824));
    jdff dff_A_DN5dca3V1_0(.din(n21818), .dout(n21821));
    jdff dff_A_clG1kHoL9_0(.din(n21815), .dout(n21818));
    jdff dff_A_8YV8pcFe0_0(.din(n21812), .dout(n21815));
    jdff dff_A_2MU3zQs79_0(.din(n21809), .dout(n21812));
    jdff dff_A_0gsqbsOX9_1(.din(n3769), .dout(n21809));
    jdff dff_A_UTqRB3JZ8_0(.din(n21803), .dout(G865));
    jdff dff_A_1vfEAqKj1_0(.din(n21800), .dout(n21803));
    jdff dff_A_ZKR4KOu15_0(.din(n21797), .dout(n21800));
    jdff dff_A_9HLefwsM7_0(.din(n21794), .dout(n21797));
    jdff dff_A_Xvirj3x92_1(.din(n3746), .dout(n21794));
    jdff dff_A_ybX7Iq9q0_0(.din(n21788), .dout(G863));
    jdff dff_A_ve4s6jcr8_0(.din(n21785), .dout(n21788));
    jdff dff_A_0yPptQX48_0(.din(n21782), .dout(n21785));
    jdff dff_A_Db0Se1s10_1(.din(n3717), .dout(n21782));
    jdff dff_A_G2xREmvo6_0(.din(n21776), .dout(G854));
    jdff dff_A_zEGDd7WI3_0(.din(n21773), .dout(n21776));
    jdff dff_A_vLnah9Nh3_0(.din(n21770), .dout(n21773));
    jdff dff_A_fBGxTbSY1_0(.din(n21767), .dout(n21770));
    jdff dff_A_a2gz8XBV4_0(.din(n21764), .dout(n21767));
    jdff dff_A_JuBUJKWv1_0(.din(n21761), .dout(n21764));
    jdff dff_A_qiqBJ46L3_0(.din(n21758), .dout(n21761));
    jdff dff_A_zwbI27Zl7_0(.din(n21755), .dout(n21758));
    jdff dff_A_OIHn8raU3_0(.din(n21752), .dout(n21755));
    jdff dff_A_K4h0biQT9_0(.din(n21749), .dout(n21752));
    jdff dff_A_7HfiSwIN0_0(.din(n21746), .dout(n21749));
    jdff dff_A_FQcx36GC3_0(.din(n21743), .dout(n21746));
    jdff dff_A_0kZnrD8X5_0(.din(n21740), .dout(n21743));
    jdff dff_A_NHzDBLZ10_0(.din(n21737), .dout(n21740));
    jdff dff_A_CJc1MQX59_0(.din(n21734), .dout(n21737));
    jdff dff_A_kppvDxAs8_2(.din(n3691), .dout(n21734));
    jdff dff_A_vkIbfGlh2_0(.din(n21728), .dout(G830));
    jdff dff_A_CGCd2iDo0_0(.din(n21725), .dout(n21728));
    jdff dff_A_oW4Mql2N5_0(.din(n21722), .dout(n21725));
    jdff dff_A_hqvWELcf9_0(.din(n21719), .dout(n21722));
    jdff dff_A_eJEjRJto9_0(.din(n21716), .dout(n21719));
    jdff dff_A_aqjkUbL88_0(.din(n21713), .dout(n21716));
    jdff dff_A_nTf3kGoq3_0(.din(n21710), .dout(n21713));
    jdff dff_A_Qi12p23v0_0(.din(n21707), .dout(n21710));
    jdff dff_A_FIVSn6jT5_1(.din(n3660), .dout(n21707));
    jdff dff_A_IEdhuDou6_0(.din(n21701), .dout(G828));
    jdff dff_A_IPO3asO77_0(.din(n21698), .dout(n21701));
    jdff dff_A_QdSxRkTV5_0(.din(n21695), .dout(n21698));
    jdff dff_A_EC7USFKY8_0(.din(n21692), .dout(n21695));
    jdff dff_A_XlDDOS1I0_0(.din(n21689), .dout(n21692));
    jdff dff_A_AZMS5jDx8_0(.din(n21686), .dout(n21689));
    jdff dff_A_U8enSGN17_0(.din(n21683), .dout(n21686));
    jdff dff_A_Bmlo6mAl5_1(.din(n3634), .dout(n21683));
    jdff dff_A_5aEQ9g5v0_0(.din(n21677), .dout(G826));
    jdff dff_A_ju0hEPEo9_0(.din(n21674), .dout(n21677));
    jdff dff_A_AR8ckWXU8_0(.din(n21671), .dout(n21674));
    jdff dff_A_SjK7TBBe2_0(.din(n21668), .dout(n21671));
    jdff dff_A_wEHEWSJm2_0(.din(n21665), .dout(n21668));
    jdff dff_A_bDH0qyyM4_0(.din(n21662), .dout(n21665));
    jdff dff_A_YL4vOG652_0(.din(n21659), .dout(n21662));
    jdff dff_A_G7R4DQMb4_1(.din(n3611), .dout(n21659));
    jdff dff_A_BS2SFMqn9_0(.din(n21653), .dout(G824));
    jdff dff_A_ll0iwTxF4_0(.din(n21650), .dout(n21653));
    jdff dff_A_s63tS9o31_0(.din(n21647), .dout(n21650));
    jdff dff_A_sXU9p2Em6_0(.din(n21644), .dout(n21647));
    jdff dff_A_H9l19U0M7_1(.din(n3588), .dout(n21644));
    jdff dff_A_r5dLtpmm2_0(.din(n21638), .dout(G813));
    jdff dff_A_KEmcbVxm3_0(.din(n21635), .dout(n21638));
    jdff dff_A_Fc2CDHyE3_0(.din(n21632), .dout(n21635));
    jdff dff_A_MgBElAsh9_0(.din(n21629), .dout(n21632));
    jdff dff_A_pWQMjWgi5_0(.din(n21626), .dout(n21629));
    jdff dff_A_osVvMOyj5_0(.din(n21623), .dout(n21626));
    jdff dff_A_2MfCMQnB8_0(.din(n21620), .dout(n21623));
    jdff dff_A_xgw7p0Rd0_0(.din(n21617), .dout(n21620));
    jdff dff_A_wjwk8NfH6_2(.din(n3565), .dout(n21617));
    jdff dff_A_0pY5zyR49_0(.din(n21611), .dout(G818));
    jdff dff_A_Nmyz9r8A8_0(.din(n21608), .dout(n21611));
    jdff dff_A_irnvtUxB4_0(.din(n21605), .dout(n21608));
    jdff dff_A_u6EqJ3Cf5_0(.din(n21602), .dout(n21605));
    jdff dff_A_PL0nReCd3_2(.din(n3557), .dout(n21602));
    jdff dff_A_NbP1wXAe0_0(.din(n21596), .dout(G702));
    jdff dff_A_ShpImyfo3_0(.din(n21593), .dout(n21596));
    jdff dff_A_q0FWV8NW2_0(.din(n21590), .dout(n21593));
    jdff dff_A_Ny37ee9D9_0(.din(n21587), .dout(n21590));
    jdff dff_A_W0P9SmEA4_0(.din(n21584), .dout(n21587));
    jdff dff_A_VIbBDNCn6_0(.din(n21581), .dout(n21584));
    jdff dff_A_PD7GVt7w3_0(.din(n21578), .dout(n21581));
    jdff dff_A_pI4UzbjX7_2(.din(n3494), .dout(n21578));
    jdff dff_A_74UZtK6D7_0(.din(n21572), .dout(G699));
    jdff dff_A_w0wt9ylw3_0(.din(n21569), .dout(n21572));
    jdff dff_A_VEesDnjg3_0(.din(n21566), .dout(n21569));
    jdff dff_A_1fEYA2CO0_0(.din(n21563), .dout(n21566));
    jdff dff_A_5DR4MYjN6_0(.din(n21560), .dout(n21563));
    jdff dff_A_60WASzlJ6_0(.din(n21557), .dout(n21560));
    jdff dff_A_DLSBcTjB7_0(.din(n21554), .dout(n21557));
    jdff dff_A_JGwoNHNd1_0(.din(n21551), .dout(n21554));
    jdff dff_A_AX6UZEQe8_2(.din(n3462), .dout(n21551));
    jdff dff_A_RYqammxv7_0(.din(n21545), .dout(G696));
    jdff dff_A_jOZEJrWW1_0(.din(n21542), .dout(n21545));
    jdff dff_A_Pgb2sB8L8_0(.din(n21539), .dout(n21542));
    jdff dff_A_H303VnPt9_0(.din(n21536), .dout(n21539));
    jdff dff_A_LhURLAYy2_0(.din(n21533), .dout(n21536));
    jdff dff_A_I4j4iM1L0_0(.din(n21530), .dout(n21533));
    jdff dff_A_Ei7LzMha6_0(.din(n21527), .dout(n21530));
    jdff dff_A_KosG7yld5_0(.din(n21524), .dout(n21527));
    jdff dff_A_8PyI6sKE1_0(.din(n21521), .dout(n21524));
    jdff dff_A_MqQBwMxU9_2(.din(n3430), .dout(n21521));
    jdff dff_A_t38XyCSz3_0(.din(n21515), .dout(G676));
    jdff dff_A_Wbt5YpQd5_0(.din(n21512), .dout(n21515));
    jdff dff_A_HRPcuduB5_0(.din(n21509), .dout(n21512));
    jdff dff_A_01xYAUnS3_0(.din(n21506), .dout(n21509));
    jdff dff_A_X8y2MPUc5_0(.din(n21503), .dout(n21506));
    jdff dff_A_Dt6jwWtM8_2(.din(n3398), .dout(n21503));
    jdff dff_A_4ZYvl2q66_0(.din(n21497), .dout(G670));
    jdff dff_A_c9VTKL0p0_0(.din(n21494), .dout(n21497));
    jdff dff_A_F4PkPkyH6_0(.din(n21491), .dout(n21494));
    jdff dff_A_EAuFQQyb3_0(.din(n21488), .dout(n21491));
    jdff dff_A_ZpX5zIOT4_0(.din(n21485), .dout(n21488));
    jdff dff_A_0rAlDyUm2_0(.din(n21482), .dout(n21485));
    jdff dff_A_4tbiLbgq2_0(.din(n21479), .dout(n21482));
    jdff dff_A_BCHA1aqF8_2(.din(n3366), .dout(n21479));
    jdff dff_A_NK31XUtu1_0(.din(n21473), .dout(G667));
    jdff dff_A_zsBSBdfK1_0(.din(n21470), .dout(n21473));
    jdff dff_A_T2bI25Oj5_0(.din(n21467), .dout(n21470));
    jdff dff_A_yJUKYI1N5_0(.din(n21464), .dout(n21467));
    jdff dff_A_pNUKCvzA0_0(.din(n21461), .dout(n21464));
    jdff dff_A_CdPWBX9T4_0(.din(n21458), .dout(n21461));
    jdff dff_A_Cy3dTs2N4_0(.din(n21455), .dout(n21458));
    jdff dff_A_vRwhH48E3_0(.din(n21452), .dout(n21455));
    jdff dff_A_3hWNAct47_2(.din(n3334), .dout(n21452));
    jdff dff_A_pTC26Tiz3_0(.din(n21446), .dout(G664));
    jdff dff_A_inf7Of335_0(.din(n21443), .dout(n21446));
    jdff dff_A_yZQ2yunU8_0(.din(n21440), .dout(n21443));
    jdff dff_A_cW0sIP7H9_0(.din(n21437), .dout(n21440));
    jdff dff_A_6Ux2QBei0_0(.din(n21434), .dout(n21437));
    jdff dff_A_5tssc9dj5_0(.din(n21431), .dout(n21434));
    jdff dff_A_ndU0ew5q3_0(.din(n21428), .dout(n21431));
    jdff dff_A_cJNFi75R8_0(.din(n21425), .dout(n21428));
    jdff dff_A_GRR10IgP0_0(.din(n21422), .dout(n21425));
    jdff dff_A_8re8Z0rV0_2(.din(n3302), .dout(n21422));
    jdff dff_A_utYL87sS2_0(.din(n21416), .dout(G642));
    jdff dff_A_cSrNiilW2_0(.din(n21413), .dout(n21416));
    jdff dff_A_yawDQFw12_0(.din(n21410), .dout(n21413));
    jdff dff_A_KyNOtPHU3_0(.din(n21407), .dout(n21410));
    jdff dff_A_z17Rcdpv0_0(.din(n21404), .dout(n21407));
    jdff dff_A_6rpt8BSf5_2(.din(n3270), .dout(n21404));
    jdff dff_A_aQZEqZ2H8_0(.din(n21398), .dout(G802));
    jdff dff_A_CYnA1xGP9_0(.din(n21395), .dout(n21398));
    jdff dff_A_l9nTWXBB3_0(.din(n21392), .dout(n21395));
    jdff dff_A_89UOq2Qy0_0(.din(n21389), .dout(n21392));
    jdff dff_A_OUTDsZUk6_0(.din(n21386), .dout(n21389));
    jdff dff_A_1Zb7RLc86_0(.din(n21383), .dout(n21386));
    jdff dff_A_FiW4QVMn3_0(.din(n21380), .dout(n21383));
    jdff dff_A_r8CcTp2v1_0(.din(n21377), .dout(n21380));
    jdff dff_A_nlQVr92Q0_0(.din(n21374), .dout(n21377));
    jdff dff_A_6qTWw12u7_0(.din(n21371), .dout(n21374));
    jdff dff_A_axuI5cBD5_2(.din(n3238), .dout(n21371));
    jdff dff_A_NQrAO3Rv3_0(.din(n21365), .dout(G797));
    jdff dff_A_AGcDh32s5_0(.din(n21362), .dout(n21365));
    jdff dff_A_7cTf1T4i3_0(.din(n21359), .dout(n21362));
    jdff dff_A_8xqp0GbX0_0(.din(n21356), .dout(n21359));
    jdff dff_A_XDTDN5YN7_0(.din(n21353), .dout(n21356));
    jdff dff_A_IqxEx9ys7_0(.din(n21350), .dout(n21353));
    jdff dff_A_7onYI73d0_0(.din(n21347), .dout(n21350));
    jdff dff_A_WyJvKw7E0_0(.din(n21344), .dout(n21347));
    jdff dff_A_vNqj2az50_0(.din(n21341), .dout(n21344));
    jdff dff_A_7sYsf6TN1_2(.din(n3210), .dout(n21341));
    jdff dff_A_P7pf4Vfe9_0(.din(n21335), .dout(G792));
    jdff dff_A_ICfuHqFr6_0(.din(n21332), .dout(n21335));
    jdff dff_A_HUolGx9D6_0(.din(n21329), .dout(n21332));
    jdff dff_A_WJQibS2G0_0(.din(n21326), .dout(n21329));
    jdff dff_A_pGhyNCH50_0(.din(n21323), .dout(n21326));
    jdff dff_A_e658WdM31_0(.din(n21320), .dout(n21323));
    jdff dff_A_SU6dX10N2_0(.din(n21317), .dout(n21320));
    jdff dff_A_uz6TL8Fv8_0(.din(n21314), .dout(n21317));
    jdff dff_A_oRgwlr2S2_2(.din(n3182), .dout(n21314));
    jdff dff_A_HNL4anZJ1_0(.din(n21308), .dout(G787));
    jdff dff_A_jIVTXgdV8_0(.din(n21305), .dout(n21308));
    jdff dff_A_ccbMY84v3_0(.din(n21302), .dout(n21305));
    jdff dff_A_j2MpnEKC7_0(.din(n21299), .dout(n21302));
    jdff dff_A_CDNEXem76_0(.din(n21296), .dout(n21299));
    jdff dff_A_Ex4eapIB2_0(.din(n21293), .dout(n21296));
    jdff dff_A_cPQHNv5B9_2(.din(n3154), .dout(n21293));
    jdff dff_A_psBQKyDZ2_0(.din(n21287), .dout(G762));
    jdff dff_A_EuGEL2YL8_0(.din(n21284), .dout(n21287));
    jdff dff_A_XblsMeDR1_0(.din(n21281), .dout(n21284));
    jdff dff_A_bC9aoJ696_0(.din(n21278), .dout(n21281));
    jdff dff_A_eEZWHRGO0_0(.din(n21275), .dout(n21278));
    jdff dff_A_BJ3sBhf47_0(.din(n21272), .dout(n21275));
    jdff dff_A_7BkNzJCb6_0(.din(n21269), .dout(n21272));
    jdff dff_A_FvOsX6rh2_0(.din(n21266), .dout(n21269));
    jdff dff_A_Q4LeZp0o5_0(.din(n21263), .dout(n21266));
    jdff dff_A_WpKOQMgU6_0(.din(n21260), .dout(n21263));
    jdff dff_A_V5IgNeJF5_2(.din(n3126), .dout(n21260));
    jdff dff_A_yHFZUxf10_0(.din(n21254), .dout(G757));
    jdff dff_A_2YYotMmc5_0(.din(n21251), .dout(n21254));
    jdff dff_A_ltxeGomy7_0(.din(n21248), .dout(n21251));
    jdff dff_A_xDSaxUyy4_0(.din(n21245), .dout(n21248));
    jdff dff_A_njL2hrF09_0(.din(n21242), .dout(n21245));
    jdff dff_A_QWdDj9Qn7_0(.din(n21239), .dout(n21242));
    jdff dff_A_aPagkDPs1_0(.din(n21236), .dout(n21239));
    jdff dff_A_1Y3wWmRJ0_0(.din(n21233), .dout(n21236));
    jdff dff_A_ksAJL9kY7_0(.din(n21230), .dout(n21233));
    jdff dff_A_m9mvQOBB9_2(.din(n3092), .dout(n21230));
    jdff dff_A_E9glpBty5_0(.din(n21224), .dout(G752));
    jdff dff_A_CWPC1Hao1_0(.din(n21221), .dout(n21224));
    jdff dff_A_q1ZP4Ju71_0(.din(n21218), .dout(n21221));
    jdff dff_A_Ec8wgNHe0_0(.din(n21215), .dout(n21218));
    jdff dff_A_ADLXexMg5_0(.din(n21212), .dout(n21215));
    jdff dff_A_jeVaUGCm4_0(.din(n21209), .dout(n21212));
    jdff dff_A_M8Yz6tkD9_0(.din(n21206), .dout(n21209));
    jdff dff_A_lwtRUbdz2_0(.din(n21203), .dout(n21206));
    jdff dff_A_g0IwlMxo1_2(.din(n3058), .dout(n21203));
    jdff dff_A_UcorWion6_0(.din(n21197), .dout(G747));
    jdff dff_A_pP2OPXy75_0(.din(n21194), .dout(n21197));
    jdff dff_A_VhQuBeBX9_0(.din(n21191), .dout(n21194));
    jdff dff_A_bKoO846w1_0(.din(n21188), .dout(n21191));
    jdff dff_A_s48iNXK05_0(.din(n21185), .dout(n21188));
    jdff dff_A_W2BFYOlt5_0(.din(n21182), .dout(n21185));
    jdff dff_A_xNgk3bJf2_2(.din(n3024), .dout(n21182));
    jdff dff_A_MjH02BQJ1_0(.din(n21176), .dout(G693));
    jdff dff_A_3h2XP5c53_0(.din(n21173), .dout(n21176));
    jdff dff_A_fTI4crZ25_0(.din(n21170), .dout(n21173));
    jdff dff_A_7dbf1h419_0(.din(n21167), .dout(n21170));
    jdff dff_A_dHBnbEgv2_0(.din(n21164), .dout(n21167));
    jdff dff_A_I7zMWBsM7_0(.din(n21161), .dout(n21164));
    jdff dff_A_ncsfzng79_0(.din(n21158), .dout(n21161));
    jdff dff_A_8IpmZLyl1_0(.din(n21155), .dout(n21158));
    jdff dff_A_I4WTF1c89_0(.din(n21152), .dout(n21155));
    jdff dff_A_KkGM2XdS9_0(.din(n21149), .dout(n21152));
    jdff dff_A_1ej4X1Vz2_0(.din(n21146), .dout(n21149));
    jdff dff_A_TNXH6GIs1_0(.din(n21143), .dout(n21146));
    jdff dff_A_mZ8pUlFz5_0(.din(n21140), .dout(n21143));
    jdff dff_A_T2PMMgd24_2(.din(n2990), .dout(n21140));
    jdff dff_A_jjXailx57_0(.din(n21134), .dout(G661));
    jdff dff_A_ONibe0tZ3_0(.din(n21131), .dout(n21134));
    jdff dff_A_Y8i03vy06_0(.din(n21128), .dout(n21131));
    jdff dff_A_gF1yE8Rg5_0(.din(n21125), .dout(n21128));
    jdff dff_A_1sDO05d45_0(.din(n21122), .dout(n21125));
    jdff dff_A_wvNU9kS00_0(.din(n21119), .dout(n21122));
    jdff dff_A_yw6LOFQ46_0(.din(n21116), .dout(n21119));
    jdff dff_A_Qy9pUNkj4_0(.din(n21113), .dout(n21116));
    jdff dff_A_t8fnELcm5_0(.din(n21110), .dout(n21113));
    jdff dff_A_FJ6BLk6H5_0(.din(n21107), .dout(n21110));
    jdff dff_A_PSu94Fp34_0(.din(n21104), .dout(n21107));
    jdff dff_A_Iyon78Eh2_0(.din(n21101), .dout(n21104));
    jdff dff_A_O1uS5i5W7_0(.din(n21098), .dout(n21101));
    jdff dff_A_BjvcmaIf8_2(.din(n2936), .dout(n21098));
    jdff dff_A_FqGrfaly0_0(.din(n21092), .dout(G585));
    jdff dff_A_G63HbYJb4_0(.din(n21089), .dout(n21092));
    jdff dff_A_UbtI2DGo5_0(.din(n21086), .dout(n21089));
    jdff dff_A_1sFFBQuW9_0(.din(n21083), .dout(n21086));
    jdff dff_A_JNkxd2Je5_0(.din(n21080), .dout(n21083));
    jdff dff_A_SYXW0W7J6_0(.din(n21077), .dout(n21080));
    jdff dff_A_1nQkdxS48_0(.din(n21074), .dout(n21077));
    jdff dff_A_aPAHZ5LL4_2(.din(n2882), .dout(n21074));
    jdff dff_A_51s5SvMF4_0(.din(n21068), .dout(G575));
    jdff dff_A_XoYOnOg67_0(.din(n21065), .dout(n21068));
    jdff dff_A_PlH2NXOH3_0(.din(n21062), .dout(n21065));
    jdff dff_A_cx4CKnL32_0(.din(n21059), .dout(n21062));
    jdff dff_A_ZwVSUgu01_2(.din(n2816), .dout(n21059));
    jdff dff_A_UkYV04p32_0(.din(n21053), .dout(G1000));
    jdff dff_A_v6IyGWyY9_0(.din(n21050), .dout(n21053));
    jdff dff_A_WFluOpEp0_0(.din(n21047), .dout(n21050));
    jdff dff_A_TscTtr5T5_0(.din(n21044), .dout(n21047));
    jdff dff_A_lqnMz7y54_0(.din(n21041), .dout(n21044));
    jdff dff_A_P057rDQ20_0(.din(n21038), .dout(n21041));
    jdff dff_A_18nj1Z018_0(.din(n21035), .dout(n21038));
    jdff dff_A_z4QWg72y8_0(.din(n21032), .dout(n21035));
    jdff dff_A_C11h4Fyo7_0(.din(n21029), .dout(n21032));
    jdff dff_A_a52EhNS14_0(.din(n21026), .dout(n21029));
    jdff dff_A_qdLImWtr9_0(.din(n21023), .dout(n21026));
    jdff dff_A_ujXf7ey06_0(.din(n21020), .dout(n21023));
    jdff dff_A_gKKBMyGH2_0(.din(n21017), .dout(n21020));
    jdff dff_A_gpSSDnqP8_0(.din(n21014), .dout(n21017));
    jdff dff_A_txTUDvuk0_0(.din(n21011), .dout(n21014));
    jdff dff_A_o0iOlF0S9_0(.din(n21008), .dout(n21011));
    jdff dff_A_iKEkTV5t6_0(.din(n21005), .dout(n21008));
    jdff dff_A_lol7tGyc9_0(.din(n21002), .dout(n21005));
    jdff dff_A_vxWk0kuz4_1(.din(n2677), .dout(n21002));
    jdff dff_A_xJCTIBfG9_0(.din(n20996), .dout(G998));
    jdff dff_A_Gz5Kq3nn1_0(.din(n20993), .dout(n20996));
    jdff dff_A_PUJJon1W6_0(.din(n20990), .dout(n20993));
    jdff dff_A_3d3sMt6m5_0(.din(n20987), .dout(n20990));
    jdff dff_A_TmORDFHX5_0(.din(n20984), .dout(n20987));
    jdff dff_A_MB8Gfrb67_0(.din(n20981), .dout(n20984));
    jdff dff_A_UlofxvGN3_0(.din(n20978), .dout(n20981));
    jdff dff_A_CAcrCyCy6_0(.din(n20975), .dout(n20978));
    jdff dff_A_x6hpU3qV9_0(.din(n20972), .dout(n20975));
    jdff dff_A_rz5qe9ya3_0(.din(n20969), .dout(n20972));
    jdff dff_A_tMCRbGHo2_0(.din(n20966), .dout(n20969));
    jdff dff_A_Yc6tf6mU9_0(.din(n20963), .dout(n20966));
    jdff dff_A_DBRdP60S9_0(.din(n20960), .dout(n20963));
    jdff dff_A_PtOWfpMy2_0(.din(n20957), .dout(n20960));
    jdff dff_A_ixcoWCSO2_0(.din(n20954), .dout(n20957));
    jdff dff_A_T9asdqcq4_0(.din(n20951), .dout(n20954));
    jdff dff_A_rsHUFwPC0_1(.din(n2629), .dout(n20951));
    jdff dff_A_3QUBX8Qt3_0(.din(n20945), .dout(G877));
    jdff dff_A_ufoCXX3U0_0(.din(n20942), .dout(n20945));
    jdff dff_A_gUT7qUu26_0(.din(n20939), .dout(n20942));
    jdff dff_A_b4ooQjrS2_0(.din(n20936), .dout(n20939));
    jdff dff_A_bMf3h5LL5_0(.din(n20933), .dout(n20936));
    jdff dff_A_IHvtxObP5_0(.din(n20930), .dout(n20933));
    jdff dff_A_JAenVpx02_0(.din(n20927), .dout(n20930));
    jdff dff_A_ODIXZ89F6_0(.din(n20924), .dout(n20927));
    jdff dff_A_k5ZtWuAc5_0(.din(n20921), .dout(n20924));
    jdff dff_A_dBpxepUG6_0(.din(n20918), .dout(n20921));
    jdff dff_A_podGFzGD8_0(.din(n20915), .dout(n20918));
    jdff dff_A_VWi6s1Jw2_0(.din(n20912), .dout(n20915));
    jdff dff_A_4NKiSx5A2_0(.din(n20909), .dout(n20912));
    jdff dff_A_M2r8JevI0_1(.din(n2568), .dout(n20909));
    jdff dff_A_Q01r9AYR6_0(.din(n20903), .dout(G875));
    jdff dff_A_6hDRUkCX4_0(.din(n20900), .dout(n20903));
    jdff dff_A_Zp2sodSg8_0(.din(n20897), .dout(n20900));
    jdff dff_A_Fulb2dLV5_0(.din(n20894), .dout(n20897));
    jdff dff_A_HnAfBtkG4_0(.din(n20891), .dout(n20894));
    jdff dff_A_jwa96Fl75_0(.din(n20888), .dout(n20891));
    jdff dff_A_93DO8Yf21_0(.din(n20885), .dout(n20888));
    jdff dff_A_pgJa7A665_0(.din(n20882), .dout(n20885));
    jdff dff_A_U50f7xEO2_0(.din(n20879), .dout(n20882));
    jdff dff_A_m9DOy8Tk0_0(.din(n20876), .dout(n20879));
    jdff dff_A_RkhlHoH04_0(.din(n20873), .dout(n20876));
    jdff dff_A_VYoBtlWz3_0(.din(n20870), .dout(n20873));
    jdff dff_A_5zsUPBA47_1(.din(n2527), .dout(n20870));
    jdff dff_A_hq6ePeyd7_0(.din(n20864), .dout(G873));
    jdff dff_A_PZOjwCQ04_0(.din(n20861), .dout(n20864));
    jdff dff_A_p11MuTuQ9_0(.din(n20858), .dout(n20861));
    jdff dff_A_ZAVSQPGH8_0(.din(n20855), .dout(n20858));
    jdff dff_A_hYyeh1fV6_0(.din(n20852), .dout(n20855));
    jdff dff_A_A7pY0dpX1_0(.din(n20849), .dout(n20852));
    jdff dff_A_p1vJkx1M8_0(.din(n20846), .dout(n20849));
    jdff dff_A_g94nGanx7_0(.din(n20843), .dout(n20846));
    jdff dff_A_CvZYO3aI0_0(.din(n20840), .dout(n20843));
    jdff dff_A_ypNE6hvh7_0(.din(n20837), .dout(n20840));
    jdff dff_A_c64wwYKJ4_0(.din(n20834), .dout(n20837));
    jdff dff_A_Z21vggDg8_1(.din(n2478), .dout(n20834));
    jdff dff_A_dPMgjU3R7_0(.din(n20828), .dout(G871));
    jdff dff_A_ppkBLltQ7_0(.din(n20825), .dout(n20828));
    jdff dff_A_mFOiPj4c2_0(.din(n20822), .dout(n20825));
    jdff dff_A_Hpj30Ax63_0(.din(n20819), .dout(n20822));
    jdff dff_A_ISZ4NYmR7_0(.din(n20816), .dout(n20819));
    jdff dff_A_RV1WwCaw6_0(.din(n20813), .dout(n20816));
    jdff dff_A_vCOILdJZ5_0(.din(n20810), .dout(n20813));
    jdff dff_A_drEy0vdf7_0(.din(n20807), .dout(n20810));
    jdff dff_A_Uqa9WElK9_0(.din(n20804), .dout(n20807));
    jdff dff_A_N7LHGUu06_1(.din(n2451), .dout(n20804));
    jdff dff_A_1jIKfZT23_0(.din(n20798), .dout(G859));
    jdff dff_A_MuzgbhDl3_0(.din(n20795), .dout(n20798));
    jdff dff_A_pbVMcsM92_0(.din(n20792), .dout(n20795));
    jdff dff_A_h2U5pKVg1_0(.din(n20789), .dout(n20792));
    jdff dff_A_rarOqqIw2_0(.din(n20786), .dout(n20789));
    jdff dff_A_yykVMFx44_0(.din(n20783), .dout(n20786));
    jdff dff_A_BHu1VUKb9_0(.din(n20780), .dout(n20783));
    jdff dff_A_6Etd3qUY3_0(.din(n20777), .dout(n20780));
    jdff dff_A_WFMfEKIz5_0(.din(n20774), .dout(n20777));
    jdff dff_A_cr3jm7j96_0(.din(n20771), .dout(n20774));
    jdff dff_A_WeGYUlUa8_0(.din(n20768), .dout(n20771));
    jdff dff_A_e2k2DRdl7_0(.din(n20765), .dout(n20768));
    jdff dff_A_IYtFxu9W0_0(.din(n20762), .dout(n20765));
    jdff dff_A_ilQmmqJD0_0(.din(n20759), .dout(n20762));
    jdff dff_A_7O2wzkaw1_2(.din(n2388), .dout(n20759));
    jdff dff_A_r7DH87ma9_0(.din(n20753), .dout(G836));
    jdff dff_A_NzPM8eWl4_0(.din(n20750), .dout(n20753));
    jdff dff_A_jPf8QPi70_0(.din(n20747), .dout(n20750));
    jdff dff_A_0ulM0GLY8_0(.din(n20744), .dout(n20747));
    jdff dff_A_SBVJSIm32_0(.din(n20741), .dout(n20744));
    jdff dff_A_LqJlf77v3_0(.din(n20738), .dout(n20741));
    jdff dff_A_oXW4n89S0_0(.din(n20735), .dout(n20738));
    jdff dff_A_2IXg8DsH0_0(.din(n20732), .dout(n20735));
    jdff dff_A_389TtBxd9_0(.din(n20729), .dout(n20732));
    jdff dff_A_18j6Fyyx0_0(.din(n20726), .dout(n20729));
    jdff dff_A_9jv2sYF36_0(.din(n20723), .dout(n20726));
    jdff dff_A_PWBe3cmi9_0(.din(n20720), .dout(n20723));
    jdff dff_A_ybg4YFsM6_0(.din(n20717), .dout(n20720));
    jdff dff_A_Ii5ZwzAM5_0(.din(n20714), .dout(n20717));
    jdff dff_A_qGoG3T8h0_0(.din(n20711), .dout(n20714));
    jdff dff_A_qqGvtkqc6_1(.din(n2338), .dout(n20711));
    jdff dff_A_AA3ph8CU2_0(.din(n20705), .dout(G834));
    jdff dff_A_8MZY8CUr4_0(.din(n20702), .dout(n20705));
    jdff dff_A_DDmMEMTW2_0(.din(n20699), .dout(n20702));
    jdff dff_A_goRRc3wp5_0(.din(n20696), .dout(n20699));
    jdff dff_A_JuZhTEyw5_0(.din(n20693), .dout(n20696));
    jdff dff_A_WcamD9mg6_0(.din(n20690), .dout(n20693));
    jdff dff_A_Jg4vQ9HV2_0(.din(n20687), .dout(n20690));
    jdff dff_A_rAXf54PX9_0(.din(n20684), .dout(n20687));
    jdff dff_A_shiYJbDp9_0(.din(n20681), .dout(n20684));
    jdff dff_A_icOXVjl64_0(.din(n20678), .dout(n20681));
    jdff dff_A_OetBEDxM9_0(.din(n20675), .dout(n20678));
    jdff dff_A_t7z3xsnm6_0(.din(n20672), .dout(n20675));
    jdff dff_A_lMOqQ0rS8_0(.din(n20669), .dout(n20672));
    jdff dff_A_5Xx6TgKH7_1(.din(n2295), .dout(n20669));
    jdff dff_A_FdOzntpk3_0(.din(n20663), .dout(G832));
    jdff dff_A_7WDLAm422_0(.din(n20660), .dout(n20663));
    jdff dff_A_rB5l1Dxt4_0(.din(n20657), .dout(n20660));
    jdff dff_A_bkq4kN653_0(.din(n20654), .dout(n20657));
    jdff dff_A_PSykAM4I7_0(.din(n20651), .dout(n20654));
    jdff dff_A_c2vFd4CO8_0(.din(n20648), .dout(n20651));
    jdff dff_A_bBuWOqqy7_0(.din(n20645), .dout(n20648));
    jdff dff_A_MUGDUylO6_0(.din(n20642), .dout(n20645));
    jdff dff_A_SM2wA2Wy3_0(.din(n20639), .dout(n20642));
    jdff dff_A_og1H0ZN97_0(.din(n20636), .dout(n20639));
    jdff dff_A_XfJEjMF64_0(.din(n20633), .dout(n20636));
    jdff dff_A_wR17c80c2_1(.din(n2249), .dout(n20633));
    jdff dff_A_IbBxoM2o5_0(.din(n20627), .dout(G722));
    jdff dff_A_br8hVELs5_0(.din(n20624), .dout(n20627));
    jdff dff_A_UOiucRSY6_0(.din(n20621), .dout(n20624));
    jdff dff_A_VvWL19su1_0(.din(n20618), .dout(n20621));
    jdff dff_A_CQB6sj5B2_0(.din(n20615), .dout(n20618));
    jdff dff_A_7d04FC6Z1_0(.din(n20612), .dout(n20615));
    jdff dff_A_jMxXD8LX8_0(.din(n20609), .dout(n20612));
    jdff dff_A_cKv4AR9w0_0(.din(n20606), .dout(n20609));
    jdff dff_A_umIRhdYr8_0(.din(n20603), .dout(n20606));
    jdff dff_A_h3ZyZ3hk0_0(.din(n20600), .dout(n20603));
    jdff dff_A_9oNu4w210_0(.din(n20597), .dout(n20600));
    jdff dff_A_UNBiD9eu9_0(.din(n20594), .dout(n20597));
    jdff dff_A_aYgdNbkN9_0(.din(n20591), .dout(n20594));
    jdff dff_A_V4EC7Dd53_0(.din(n20588), .dout(n20591));
    jdff dff_A_ZHMTSP3i6_2(.din(n2210), .dout(n20588));
    jdff dff_A_VkYGSsx51_0(.din(n20582), .dout(G623));
    jdff dff_A_3tpwft3G5_0(.din(n20579), .dout(n20582));
    jdff dff_A_MhaL0zvK2_0(.din(n20576), .dout(n20579));
    jdff dff_A_vGTJbVse1_0(.din(n20573), .dout(n20576));
    jdff dff_A_pEqBSy1B5_0(.din(n20570), .dout(n20573));
    jdff dff_A_dh5p1ikk2_0(.din(n20567), .dout(n20570));
    jdff dff_A_ThmdqykU8_1(.din(n2154), .dout(n20567));
    jdff dff_A_hTLAoxsz8_0(.din(n20561), .dout(G861));
    jdff dff_A_ya5AUVCw8_0(.din(n20558), .dout(n20561));
    jdff dff_A_oOE0Yfsj3_0(.din(n20555), .dout(n20558));
    jdff dff_A_gww8E7655_0(.din(n20552), .dout(n20555));
    jdff dff_A_kXYckNTh4_0(.din(n20549), .dout(n20552));
    jdff dff_A_iTZPwjIH7_0(.din(n20546), .dout(n20549));
    jdff dff_A_ipFZ34Lt1_0(.din(n20543), .dout(n20546));
    jdff dff_A_2WGcBnbR7_0(.din(n20540), .dout(n20543));
    jdff dff_A_v9VaeYR98_0(.din(n20537), .dout(n20540));
    jdff dff_A_JN19R1lq1_0(.din(n20534), .dout(n20537));
    jdff dff_A_Xs2t9kTr4_0(.din(n20531), .dout(n20534));
    jdff dff_A_N1YpechW1_0(.din(n20528), .dout(n20531));
    jdff dff_A_gjHY7BFg2_0(.din(n20525), .dout(n20528));
    jdff dff_A_df8MVVbc5_0(.din(n20522), .dout(n20525));
    jdff dff_A_kqFFAjy18_0(.din(n20519), .dout(n20522));
    jdff dff_A_kldSVPQ84_0(.din(n20516), .dout(n20519));
    jdff dff_A_ZZq4kYo64_0(.din(n20513), .dout(n20516));
    jdff dff_A_ZXolT0V26_1(.din(n2110), .dout(n20513));
    jdff dff_A_wVNaNbx41_0(.din(n20507), .dout(G838));
    jdff dff_A_0NMOQF9m1_0(.din(n20504), .dout(n20507));
    jdff dff_A_k1dgeqFz8_0(.din(n20501), .dout(n20504));
    jdff dff_A_lqf1ogiV1_0(.din(n20498), .dout(n20501));
    jdff dff_A_vOZGE8vc3_0(.din(n20495), .dout(n20498));
    jdff dff_A_kkH6UtBj1_0(.din(n20492), .dout(n20495));
    jdff dff_A_CC1DrSrT2_0(.din(n20489), .dout(n20492));
    jdff dff_A_lO8HBcVh6_0(.din(n20486), .dout(n20489));
    jdff dff_A_E420atvZ0_0(.din(n20483), .dout(n20486));
    jdff dff_A_1vQVqcdV0_0(.din(n20480), .dout(n20483));
    jdff dff_A_E8YSR3hE2_0(.din(n20477), .dout(n20480));
    jdff dff_A_2OaVpKAG8_0(.din(n20474), .dout(n20477));
    jdff dff_A_Uw61XWbZ4_0(.din(n20471), .dout(n20474));
    jdff dff_A_QAWQtNTc2_0(.din(n20468), .dout(n20471));
    jdff dff_A_isKRucTK0_0(.din(n20465), .dout(n20468));
    jdff dff_A_Ybo5zWwy2_0(.din(n20462), .dout(n20465));
    jdff dff_A_Ep3zLD1i4_0(.din(n20459), .dout(n20462));
    jdff dff_A_NU9RSijT7_1(.din(n2080), .dout(n20459));
    jdff dff_A_DEjCMjYR1_0(.din(n20453), .dout(G822));
    jdff dff_A_NoqhdNf00_0(.din(n20450), .dout(n20453));
    jdff dff_A_iRbCYIBv5_0(.din(n20447), .dout(n20450));
    jdff dff_A_VFHKjjf15_0(.din(n20444), .dout(n20447));
    jdff dff_A_q7fYNNpk5_0(.din(n20441), .dout(n20444));
    jdff dff_A_4pz3WHHu2_0(.din(n20438), .dout(n20441));
    jdff dff_A_9tdBiNxn1_0(.din(n20435), .dout(n20438));
    jdff dff_A_7qI3Ea5C9_0(.din(n20432), .dout(n20435));
    jdff dff_A_yASrjxQ85_0(.din(n20429), .dout(n20432));
    jdff dff_A_ao25x0TM2_0(.din(n20426), .dout(n20429));
    jdff dff_A_Y0a6UnnT6_0(.din(n20423), .dout(n20426));
    jdff dff_A_TajhmYGg3_0(.din(n20420), .dout(n20423));
    jdff dff_A_X8V0nYfi7_0(.din(n20417), .dout(n20420));
    jdff dff_A_nz9wzjG16_0(.din(n20414), .dout(n20417));
    jdff dff_A_EMmGKFik4_0(.din(n20411), .dout(n20414));
    jdff dff_A_IOaltbKl6_0(.din(n20408), .dout(n20411));
    jdff dff_A_7cy1O96o3_0(.din(n20405), .dout(n20408));
    jdff dff_A_aq8I2DKO3_0(.din(n20402), .dout(n20405));
    jdff dff_A_snZJi9ST6_1(.din(n2032), .dout(n20402));
    jdff dff_A_cZ9PTVaY6_0(.din(n20396), .dout(G629));
    jdff dff_A_b0E8rjz12_0(.din(n20393), .dout(n20396));
    jdff dff_A_XryDxHHc7_0(.din(n20390), .dout(n20393));
    jdff dff_A_2NiPPrNn4_0(.din(n20387), .dout(n20390));
    jdff dff_A_uPhWfkZE8_0(.din(n20384), .dout(n20387));
    jdff dff_A_sUSzQodi5_0(.din(n20381), .dout(n20384));
    jdff dff_A_c7vrLhPU0_0(.din(n20378), .dout(n20381));
    jdff dff_A_Qvyp2K459_0(.din(n20375), .dout(n20378));
    jdff dff_A_X3xuNiyw9_0(.din(n20372), .dout(n20375));
    jdff dff_A_7Yvj5zxD4_0(.din(n20369), .dout(n20372));
    jdff dff_A_NhrnOveV2_0(.din(n20366), .dout(n20369));
    jdff dff_A_Cy9lkNbV7_2(.din(n5549), .dout(n20366));
    jdff dff_A_YsqjyaXh4_0(.din(n20360), .dout(G621));
    jdff dff_A_YmyiEMt48_0(.din(n20357), .dout(n20360));
    jdff dff_A_PkvviMUt2_0(.din(n20354), .dout(n20357));
    jdff dff_A_i7NRLqUr7_0(.din(n20351), .dout(n20354));
    jdff dff_A_NkyevxkC1_0(.din(n20348), .dout(n20351));
    jdff dff_A_8vHnto142_0(.din(n20345), .dout(n20348));
    jdff dff_A_XVnWRPNy5_0(.din(n20342), .dout(n20345));
    jdff dff_A_x4bT6BTj0_0(.din(n20339), .dout(n20342));
    jdff dff_A_a4yXc90U1_0(.din(n20336), .dout(n20339));
    jdff dff_A_R5rS28be5_0(.din(n20333), .dout(n20336));
    jdff dff_A_d4narGFS4_0(.din(n20330), .dout(n20333));
    jdff dff_A_KD56kTfy9_2(.din(n5545), .dout(n20330));
    jdff dff_A_dVFojz512_0(.din(n20324), .dout(G618));
    jdff dff_A_9YmxPRjd2_0(.din(n20321), .dout(n20324));
    jdff dff_A_g7JJJbif9_0(.din(n20318), .dout(n20321));
    jdff dff_A_3Br8LzRX7_0(.din(n20315), .dout(n20318));
    jdff dff_A_Y6F9dhiL1_0(.din(n20312), .dout(n20315));
    jdff dff_A_mGNG4H3s8_0(.din(n20309), .dout(n20312));
    jdff dff_A_1lDnUSeg9_0(.din(n20306), .dout(n20309));
    jdff dff_A_1TzUogFk7_0(.din(n20303), .dout(n20306));
    jdff dff_A_n1DUMr9q9_0(.din(n20300), .dout(n20303));
    jdff dff_A_k3CyBxZC2_0(.din(n20297), .dout(n20300));
    jdff dff_A_XDTo9of91_0(.din(n20294), .dout(n20297));
    jdff dff_A_dUvFZuI17_2(.din(n1981), .dout(n20294));
    jdff dff_A_7iGFQniU7_0(.din(n20288), .dout(G591));
    jdff dff_A_VCVhWC6d6_0(.din(n20285), .dout(n20288));
    jdff dff_A_DemqSCnw7_0(.din(n20282), .dout(n20285));
    jdff dff_A_g6nfOlMj9_0(.din(n20279), .dout(n20282));
    jdff dff_A_yI5iJGLK9_0(.din(n20276), .dout(n20279));
    jdff dff_A_rG5dGwXV3_0(.din(n20273), .dout(n20276));
    jdff dff_A_ANbg6Wwm2_0(.din(n20270), .dout(n20273));
    jdff dff_A_zGLOD5nD8_0(.din(n20267), .dout(n20270));
    jdff dff_A_ZfCVIXFP5_0(.din(n20264), .dout(n20267));
    jdff dff_A_b14ek91s8_0(.din(n20261), .dout(n20264));
    jdff dff_A_hPhp5Y865_0(.din(n20258), .dout(n20261));
    jdff dff_A_x5Bdeqtt8_2(.din(n1853), .dout(n20258));
    jdff dff_A_JRAIqznC6_0(.din(n20252), .dout(G1004));
    jdff dff_A_2xFGmuuI8_0(.din(n20249), .dout(n20252));
    jdff dff_A_ntWxwqQK1_0(.din(n20246), .dout(n20249));
    jdff dff_A_iqOjJnuo3_0(.din(n20243), .dout(n20246));
    jdff dff_A_hfWDkREK5_0(.din(n20240), .dout(n20243));
    jdff dff_A_4e1Us7Ku2_0(.din(n20237), .dout(n20240));
    jdff dff_A_Q1qsc3s55_0(.din(n20234), .dout(n20237));
    jdff dff_A_dxCAVoLL3_0(.din(n20231), .dout(n20234));
    jdff dff_A_NHS2pa075_0(.din(n20228), .dout(n20231));
    jdff dff_A_UkrFsFir7_0(.din(n20225), .dout(n20228));
    jdff dff_A_ttrUmXIN0_0(.din(n20222), .dout(n20225));
    jdff dff_A_IK7n4Vwj6_0(.din(n20219), .dout(n20222));
    jdff dff_A_ZRANlNYg9_0(.din(n20216), .dout(n20219));
    jdff dff_A_bYF9qzDW2_0(.din(n20213), .dout(n20216));
    jdff dff_A_zseMmEC93_0(.din(n20210), .dout(n20213));
    jdff dff_A_86hg12ZQ9_0(.din(n20207), .dout(n20210));
    jdff dff_A_V1PAS0K72_0(.din(n20204), .dout(n20207));
    jdff dff_A_TkSX4e669_0(.din(n20201), .dout(n20204));
    jdff dff_A_n80DzAQ95_0(.din(n20198), .dout(n20201));
    jdff dff_A_liYurLTQ9_0(.din(n20195), .dout(n20198));
    jdff dff_A_FM7ga7ou8_1(.din(n1707), .dout(n20195));
    jdff dff_A_pheM8mO71_0(.din(n20189), .dout(G1002));
    jdff dff_A_yP86I3PT5_0(.din(n20186), .dout(n20189));
    jdff dff_A_Ez533ZU05_0(.din(n20183), .dout(n20186));
    jdff dff_A_dJA0b8xC9_0(.din(n20180), .dout(n20183));
    jdff dff_A_R3Bi5i7L2_0(.din(n20177), .dout(n20180));
    jdff dff_A_Y9LsZRIZ3_0(.din(n20174), .dout(n20177));
    jdff dff_A_7ZzzLzVy7_0(.din(n20171), .dout(n20174));
    jdff dff_A_hwvb23Lb6_0(.din(n20168), .dout(n20171));
    jdff dff_A_W8pZpPQW0_0(.din(n20165), .dout(n20168));
    jdff dff_A_QK0QUSLo3_0(.din(n20162), .dout(n20165));
    jdff dff_A_2tof4Dml2_0(.din(n20159), .dout(n20162));
    jdff dff_A_JqmkJdmq5_0(.din(n20156), .dout(n20159));
    jdff dff_A_njPV4DTd3_0(.din(n20153), .dout(n20156));
    jdff dff_A_ttc7DjDN3_0(.din(n20150), .dout(n20153));
    jdff dff_A_z7M6r6dH6_0(.din(n20147), .dout(n20150));
    jdff dff_A_G1z6TzYy4_0(.din(n20144), .dout(n20147));
    jdff dff_A_mmWYF7Z63_0(.din(n20141), .dout(n20144));
    jdff dff_A_l0AW4AGy0_0(.din(n20138), .dout(n20141));
    jdff dff_A_Ng0oECXB3_0(.din(n20135), .dout(n20138));
    jdff dff_A_DifVr3Om1_0(.din(n20132), .dout(n20135));
    jdff dff_A_8MThqmXy2_1(.din(n1668), .dout(n20132));
    jdff dff_A_Vto4TfUX5_0(.din(n20126), .dout(G632));
    jdff dff_A_DW0i6k8X9_0(.din(n20123), .dout(n20126));
    jdff dff_A_84XnLP5F1_0(.din(n20120), .dout(n20123));
    jdff dff_A_EPhcu3l71_0(.din(n20117), .dout(n20120));
    jdff dff_A_PF4yy7YQ5_0(.din(n20114), .dout(n20117));
    jdff dff_A_fKGZCOfD7_0(.din(n20111), .dout(n20114));
    jdff dff_A_0ReWyaKS8_0(.din(n20108), .dout(n20111));
    jdff dff_A_fuXWis3a2_0(.din(n20105), .dout(n20108));
    jdff dff_A_2E0x3VZI3_0(.din(n20102), .dout(n20105));
    jdff dff_A_JG0L87Ww6_0(.din(n20099), .dout(n20102));
    jdff dff_A_qBLwA6M94_0(.din(n20096), .dout(n20099));
    jdff dff_A_qxukhu7v4_0(.din(n20093), .dout(n20096));
    jdff dff_A_qKUKWfzu2_0(.din(n20090), .dout(n20093));
    jdff dff_A_XSGwYZJ66_0(.din(n20087), .dout(n20090));
    jdff dff_A_t4OEWpbI4_2(.din(n5541), .dout(n20087));
    jdff dff_A_silvTFXx7_0(.din(n20081), .dout(G626));
    jdff dff_A_zMkrSvUF8_0(.din(n20078), .dout(n20081));
    jdff dff_A_j1vu3Yto4_0(.din(n20075), .dout(n20078));
    jdff dff_A_yW1sngvI9_0(.din(n20072), .dout(n20075));
    jdff dff_A_pU8QpZRt2_0(.din(n20069), .dout(n20072));
    jdff dff_A_jEyBLj9Q6_0(.din(n20066), .dout(n20069));
    jdff dff_A_iDGcRBmp4_0(.din(n20063), .dout(n20066));
    jdff dff_A_0fdM7YKm5_0(.din(n20060), .dout(n20063));
    jdff dff_A_6eBH2sMQ8_0(.din(n20057), .dout(n20060));
    jdff dff_A_vVvcsjH78_0(.din(n20054), .dout(n20057));
    jdff dff_A_3OlaC27m3_0(.din(n20051), .dout(n20054));
    jdff dff_A_QL1opl1b8_0(.din(n20048), .dout(n20051));
    jdff dff_A_x0JF5A1q7_0(.din(n20045), .dout(n20048));
    jdff dff_A_5UvpBk0r5_0(.din(n20042), .dout(n20045));
    jdff dff_A_OGCZ5huo7_0(.din(n20039), .dout(n20042));
    jdff dff_A_qkdo91Fi2_0(.din(n20036), .dout(n20039));
    jdff dff_A_QmKqJRIv2_2(.din(n5537), .dout(n20036));
    jdff dff_A_Qysn4twB7_0(.din(n20030), .dout(G615));
    jdff dff_A_58pnp1Fr3_0(.din(n20027), .dout(n20030));
    jdff dff_A_Svx5lZzP2_0(.din(n20024), .dout(n20027));
    jdff dff_A_KL55QyXJ1_0(.din(n20021), .dout(n20024));
    jdff dff_A_tSL6M70X7_0(.din(n20018), .dout(n20021));
    jdff dff_A_Y3j9diA04_0(.din(n20015), .dout(n20018));
    jdff dff_A_HZi5PSZl0_0(.din(n20012), .dout(n20015));
    jdff dff_A_dNQgYKEB7_0(.din(n20009), .dout(n20012));
    jdff dff_A_igQvbAAg2_0(.din(n20006), .dout(n20009));
    jdff dff_A_Vz2gVHAS2_0(.din(n20003), .dout(n20006));
    jdff dff_A_t0eXidmG0_0(.din(n20000), .dout(n20003));
    jdff dff_A_wzBljx7g8_0(.din(n19997), .dout(n20000));
    jdff dff_A_HCgQiUjK2_0(.din(n19994), .dout(n19997));
    jdff dff_A_35g2JW3m8_0(.din(n19991), .dout(n19994));
    jdff dff_A_8Tk9dvqi4_0(.din(n19988), .dout(n19991));
    jdff dff_A_BC4hp5hS2_0(.din(n19985), .dout(n19988));
    jdff dff_A_n3GGxwow0_2(.din(n1633), .dout(n19985));
    jdff dff_A_LnHzd7tf5_0(.din(n19979), .dout(G588));
    jdff dff_A_IiaX7pO55_0(.din(n19976), .dout(n19979));
    jdff dff_A_KD0XfKV14_0(.din(n19973), .dout(n19976));
    jdff dff_A_aWeCwI952_0(.din(n19970), .dout(n19973));
    jdff dff_B_XssIjf5V0_1(.din(G136), .dout(n8016));
    jdff dff_B_Dal5NXoy4_0(.din(G2824), .dout(n8019));
    jdff dff_B_Mca1lwmy8_1(.din(n366), .dout(n8022));
    jdff dff_B_Fm0mRtxx3_1(.din(n390), .dout(n8025));
    jdff dff_B_D7BgWf7S7_2(.din(n412), .dout(n8028));
    jdff dff_B_S57yGqN83_1(.din(n430), .dout(n8031));
    jdff dff_B_fnTBsdyL9_1(.din(n438), .dout(n8034));
    jdff dff_B_IrVW51x29_0(.din(n442), .dout(n8037));
    jdff dff_B_KSZfTLzP9_1(.din(G24), .dout(n8040));
    jdff dff_B_ODt69OBG6_1(.din(n458), .dout(n8043));
    jdff dff_B_TiA3PYaH3_0(.din(n462), .dout(n8046));
    jdff dff_B_Jfk8n5Ey8_1(.din(G26), .dout(n8049));
    jdff dff_A_WQWmgh6x2_0(.din(n8054), .dout(n8051));
    jdff dff_A_gygGVr8w1_0(.din(n8057), .dout(n8054));
    jdff dff_A_fB1lmueH0_0(.din(n8060), .dout(n8057));
    jdff dff_A_NRmMTPDk0_0(.din(G141), .dout(n8060));
    jdff dff_A_AFxMaLQZ3_1(.din(n8066), .dout(n8063));
    jdff dff_A_9EmKaLaE6_1(.din(n8069), .dout(n8066));
    jdff dff_A_yAeXsPl21_1(.din(n8072), .dout(n8069));
    jdff dff_A_9tMO6vDT1_1(.din(G141), .dout(n8072));
    jdff dff_B_Gkskymn36_1(.din(n478), .dout(n8076));
    jdff dff_B_p9XI6owv5_0(.din(n482), .dout(n8079));
    jdff dff_B_cVsNJJHb0_1(.din(G79), .dout(n8082));
    jdff dff_B_JmCqyBqc5_1(.din(n498), .dout(n8085));
    jdff dff_B_aSvu7Tg51_0(.din(n502), .dout(n8088));
    jdff dff_B_dEkF10QY7_1(.din(G82), .dout(n8091));
    jdff dff_A_ZMRpH7Cm0_0(.din(G2358), .dout(n8093));
    jdff dff_A_bt1O9L7I5_1(.din(G2358), .dout(n8096));
    jdff dff_A_J13aWE4G7_1(.din(n8102), .dout(n8099));
    jdff dff_A_tFnwf5qe7_1(.din(n8105), .dout(n8102));
    jdff dff_A_HybsOoa34_1(.din(n8108), .dout(n8105));
    jdff dff_A_8SuW07jG0_1(.din(G141), .dout(n8108));
    jdff dff_A_ihCZD1qn1_2(.din(n8114), .dout(n8111));
    jdff dff_A_zVDY3vDk9_2(.din(n8117), .dout(n8114));
    jdff dff_A_MJuLq9HB7_2(.din(n8120), .dout(n8117));
    jdff dff_A_a5cZcJOE8_2(.din(G141), .dout(n8120));
    jdff dff_B_WsR53Ip04_1(.din(n608), .dout(n8124));
    jdff dff_B_3CzV9Jej8_1(.din(n8124), .dout(n8127));
    jdff dff_B_Nz0flp8Q2_0(.din(n838), .dout(n8130));
    jdff dff_B_pkjSE7L20_1(.din(n980), .dout(n8133));
    jdff dff_B_kW56YRH88_1(.din(n1068), .dout(n8136));
    jdff dff_B_Ly8y0O7P7_2(.din(n1629), .dout(n8139));
    jdff dff_B_HmIOfsGO3_2(.din(n1849), .dout(n8142));
    jdff dff_B_DEkXRBgq2_2(.din(n8142), .dout(n8145));
    jdff dff_B_giZSAE6j8_2(.din(n8145), .dout(n8148));
    jdff dff_B_8PzF9dIk4_1(.din(n1805), .dout(n8151));
    jdff dff_B_ED7Z7xQZ9_1(.din(n8151), .dout(n8154));
    jdff dff_B_2WzSiiHc7_1(.din(n8154), .dout(n8157));
    jdff dff_B_7XrR9Fu38_1(.din(n8157), .dout(n8160));
    jdff dff_B_ip7ldRLj3_1(.din(n1809), .dout(n8163));
    jdff dff_B_ZcvBg8Sc2_1(.din(n8163), .dout(n8166));
    jdff dff_B_fnflHZ8W5_1(.din(n8166), .dout(n8169));
    jdff dff_A_hrZEm7iI5_1(.din(n8174), .dout(n8171));
    jdff dff_A_bispfRPv1_1(.din(n8184), .dout(n8174));
    jdff dff_B_vZrKh8sv0_3(.din(n1455), .dout(n8178));
    jdff dff_B_yYpi79nI5_3(.din(n8178), .dout(n8181));
    jdff dff_B_NxnJO8Er8_3(.din(n8181), .dout(n8184));
    jdff dff_B_AeDOD12Z9_0(.din(n1451), .dout(n8187));
    jdff dff_B_whth4iwK4_2(.din(n1977), .dout(n8190));
    jdff dff_B_5CtWqWG32_2(.din(n8190), .dout(n8193));
    jdff dff_B_f5WSunBa1_2(.din(n8193), .dout(n8196));
    jdff dff_B_YGtMakNp9_2(.din(n8196), .dout(n8199));
    jdff dff_B_2SZsCcUg8_2(.din(n8199), .dout(n8202));
    jdff dff_A_Z33aOacp4_0(.din(n8207), .dout(n8204));
    jdff dff_A_QHGVysha6_0(.din(n8210), .dout(n8207));
    jdff dff_A_vT0gjAMZ6_0(.din(n8213), .dout(n8210));
    jdff dff_A_JAk0xbai5_0(.din(n8216), .dout(n8213));
    jdff dff_A_IN0CntKv1_0(.din(n8219), .dout(n8216));
    jdff dff_A_KZ6qEmH77_0(.din(n13869), .dout(n8219));
    jdff dff_B_PhzMjzHb8_0(.din(n2202), .dout(n8223));
    jdff dff_B_fBDCGOM50_0(.din(n8223), .dout(n8226));
    jdff dff_B_rGxtK9wi5_0(.din(n8226), .dout(n8229));
    jdff dff_B_ph7LqdJY4_0(.din(n8229), .dout(n8232));
    jdff dff_B_3ewiIPnx2_0(.din(n8232), .dout(n8235));
    jdff dff_B_viMLJl540_0(.din(n2198), .dout(n8238));
    jdff dff_B_b35jbf2Z3_0(.din(n2380), .dout(n8241));
    jdff dff_B_zpGI0mAt6_0(.din(n8241), .dout(n8244));
    jdff dff_B_nQPXoJiJ7_0(.din(n8244), .dout(n8247));
    jdff dff_B_rgBzz1bG1_0(.din(n8247), .dout(n8250));
    jdff dff_B_U2olVBQR0_0(.din(n8250), .dout(n8253));
    jdff dff_B_yMh7HUE44_0(.din(n2376), .dout(n8256));
    jdff dff_B_MZhMwQa67_2(.din(G61), .dout(n8259));
    jdff dff_B_5X48FtVM3_2(.din(G11), .dout(n8262));
    jdff dff_B_CChcr1BA4_2(.din(n8262), .dout(n8265));
    jdff dff_B_bXABOWnN9_0(.din(n2808), .dout(n8268));
    jdff dff_B_W2wYqFAe1_0(.din(n2800), .dout(n8271));
    jdff dff_B_KaCYtSDu2_0(.din(n2796), .dout(n8274));
    jdff dff_B_IrpWIMHD3_1(.din(n2781), .dout(n8277));
    jdff dff_B_EhSDyr2c9_1(.din(n8277), .dout(n8280));
    jdff dff_B_InlKldaq1_1(.din(n8280), .dout(n8283));
    jdff dff_B_3wJGaPeF1_1(.din(n8283), .dout(n8286));
    jdff dff_B_WESzWxWL2_0(.din(n2870), .dout(n8289));
    jdff dff_B_mSFnHuVU1_0(.din(n8289), .dout(n8292));
    jdff dff_B_mAUt7xJU8_0(.din(n2866), .dout(n8295));
    jdff dff_B_tjDkCpYo4_0(.din(n2862), .dout(n8298));
    jdff dff_B_wAe7Cz920_0(.din(n2858), .dout(n8301));
    jdff dff_B_DEajMSUz6_0(.din(n2854), .dout(n8304));
    jdff dff_B_99g6zTEi2_0(.din(n2924), .dout(n8307));
    jdff dff_B_1qYgqFH83_0(.din(n8307), .dout(n8310));
    jdff dff_B_RAli3rd30_0(.din(n8310), .dout(n8313));
    jdff dff_B_0MqjEfGd0_0(.din(n8313), .dout(n8316));
    jdff dff_B_8OjgUUdK4_0(.din(n8316), .dout(n8319));
    jdff dff_B_yzSYTJWf6_0(.din(n2920), .dout(n8322));
    jdff dff_B_R7asPy7h5_0(.din(n2978), .dout(n8325));
    jdff dff_B_M9SHpA5H4_0(.din(n8325), .dout(n8328));
    jdff dff_B_fSRNsPI46_0(.din(n8328), .dout(n8331));
    jdff dff_B_XV3u2wTd0_0(.din(n8331), .dout(n8334));
    jdff dff_B_avY0gwYw0_0(.din(n8334), .dout(n8337));
    jdff dff_B_6TjWitqE6_0(.din(n2974), .dout(n8340));
    jdff dff_B_E8Ow1mSb0_2(.din(G185), .dout(n8343));
    jdff dff_B_mg0MgxRV1_2(.din(G182), .dout(n8346));
    jdff dff_B_uQNPPLHu0_2(.din(n8346), .dout(n8349));
    jdff dff_B_wwrx8AHY9_1(.din(n2002), .dout(n8352));
    jdff dff_B_B227RsBo4_0(.din(n2021), .dout(n8355));
    jdff dff_B_xFtzP4mP1_1(.din(G131), .dout(n8358));
    jdff dff_B_QRg1MG1I3_1(.din(n8358), .dout(n8361));
    jdff dff_B_CzAGbBpC4_0(.din(n2102), .dout(n8364));
    jdff dff_B_33JdFQzd1_0(.din(n8364), .dout(n8367));
    jdff dff_B_plweYquy5_1(.din(G117), .dout(n8370));
    jdff dff_B_gUgiBgL93_1(.din(n8370), .dout(n8373));
    jdff dff_B_qPKMQyte9_0(.din(n1060), .dout(n8376));
    jdff dff_B_KjOV1hzk1_1(.din(n1029), .dout(n8379));
    jdff dff_B_47TbZlIf2_0(.din(n3020), .dout(n8382));
    jdff dff_B_4FPXO9oq2_0(.din(n3016), .dout(n8385));
    jdff dff_B_9do6CGYe5_0(.din(n8385), .dout(n8388));
    jdff dff_B_DK7afoQR6_0(.din(n8388), .dout(n8391));
    jdff dff_B_FWWB7Nqj3_0(.din(n8391), .dout(n8394));
    jdff dff_B_PEUGs7Ix9_0(.din(n8394), .dout(n8397));
    jdff dff_B_CygcLcqT8_0(.din(n8397), .dout(n8400));
    jdff dff_B_piNr54hs0_0(.din(n8400), .dout(n8403));
    jdff dff_B_JYeiFR921_0(.din(n8403), .dout(n8406));
    jdff dff_B_Rv5YJH7z6_0(.din(n8406), .dout(n8409));
    jdff dff_B_vn7svMmu9_0(.din(n8409), .dout(n8412));
    jdff dff_B_BAeuSWTx6_0(.din(n8412), .dout(n8415));
    jdff dff_B_ztWLRg0X4_0(.din(n8415), .dout(n8418));
    jdff dff_B_Ww6v3SSi1_0(.din(n3012), .dout(n8421));
    jdff dff_A_q3zLCPm63_0(.din(n8426), .dout(n8423));
    jdff dff_A_A48mdAmP4_0(.din(n8429), .dout(n8426));
    jdff dff_A_LvF52s4v5_0(.din(n8432), .dout(n8429));
    jdff dff_A_a47M2xaZ7_0(.din(n8435), .dout(n8432));
    jdff dff_A_ZgPCGr6Y6_0(.din(n8438), .dout(n8435));
    jdff dff_A_fcQliiep9_0(.din(n8441), .dout(n8438));
    jdff dff_A_DrEaSfxY2_0(.din(n12264), .dout(n8441));
    jdff dff_A_3dQy5vFe3_0(.din(n8447), .dout(n8444));
    jdff dff_A_xq15hH6Z1_0(.din(n8450), .dout(n8447));
    jdff dff_A_cvnKx47M1_0(.din(n8453), .dout(n8450));
    jdff dff_A_Uwkh47Si4_0(.din(n8456), .dout(n8453));
    jdff dff_A_sJx77pRG2_0(.din(n8459), .dout(n8456));
    jdff dff_A_VC7dsWwV8_0(.din(n8462), .dout(n8459));
    jdff dff_A_m61YsGgv0_0(.din(n8465), .dout(n8462));
    jdff dff_A_pDba1ues0_0(.din(n12402), .dout(n8465));
    jdff dff_B_4QTYj42L0_0(.din(n3054), .dout(n8469));
    jdff dff_B_CYoRH7bO6_0(.din(n3050), .dout(n8472));
    jdff dff_B_8sSrWfTZ6_0(.din(n8472), .dout(n8475));
    jdff dff_B_8w1o0Pwi9_0(.din(n8475), .dout(n8478));
    jdff dff_B_bvSipQJx4_0(.din(n8478), .dout(n8481));
    jdff dff_B_c7m6rXMD7_0(.din(n8481), .dout(n8484));
    jdff dff_B_m58G5xzA9_0(.din(n8484), .dout(n8487));
    jdff dff_B_4fJtjy4U4_0(.din(n8487), .dout(n8490));
    jdff dff_B_CDytwPxH1_0(.din(n8490), .dout(n8493));
    jdff dff_B_rwa9BTLw4_0(.din(n8493), .dout(n8496));
    jdff dff_B_gz8CIbCF7_0(.din(n8496), .dout(n8499));
    jdff dff_B_jHgqreCB4_0(.din(n3046), .dout(n8502));
    jdff dff_B_QIFUOnRh2_0(.din(n3088), .dout(n8505));
    jdff dff_B_syxrlt572_0(.din(n8505), .dout(n8508));
    jdff dff_B_ZkBOZRCt1_0(.din(n3084), .dout(n8511));
    jdff dff_B_Kmqbff6M7_0(.din(n8511), .dout(n8514));
    jdff dff_B_blFGw6jZ5_0(.din(n8514), .dout(n8517));
    jdff dff_B_e5WHWo593_0(.din(n8517), .dout(n8520));
    jdff dff_B_7ZzqMHBu9_0(.din(n8520), .dout(n8523));
    jdff dff_B_XbiAhNVy0_0(.din(n8523), .dout(n8526));
    jdff dff_B_P6BvjMBa8_0(.din(n8526), .dout(n8529));
    jdff dff_B_45NXoFSz2_0(.din(n8529), .dout(n8532));
    jdff dff_B_gOnz1Z622_0(.din(n3080), .dout(n8535));
    jdff dff_B_zng9M7Sd3_0(.din(n3122), .dout(n8538));
    jdff dff_B_KQnOpBxn5_0(.din(n8538), .dout(n8541));
    jdff dff_B_fvPzOQNK9_0(.din(n8541), .dout(n8544));
    jdff dff_B_KLoCxCNO9_0(.din(n3118), .dout(n8547));
    jdff dff_B_5xcSTM5P5_0(.din(n8547), .dout(n8550));
    jdff dff_B_fdVVnm3y2_0(.din(n8550), .dout(n8553));
    jdff dff_B_KEyaKCrz6_0(.din(n8553), .dout(n8556));
    jdff dff_B_MDnUbVep0_0(.din(n8556), .dout(n8559));
    jdff dff_B_zRMVweWr4_0(.din(n8559), .dout(n8562));
    jdff dff_B_04HM0IyZ8_0(.din(n3114), .dout(n8565));
    jdff dff_A_Oc0bOI7p6_1(.din(n8570), .dout(n8567));
    jdff dff_A_Y9bywIRN2_1(.din(n12245), .dout(n8570));
    jdff dff_A_ZwpPDw3o7_2(.din(n8576), .dout(n8573));
    jdff dff_A_5SOsB5WF6_2(.din(n8579), .dout(n8576));
    jdff dff_A_8pRe6LkT2_2(.din(n8582), .dout(n8579));
    jdff dff_A_rTCJRv862_2(.din(n12245), .dout(n8582));
    jdff dff_A_8LEd86GY1_1(.din(n12371), .dout(n8585));
    jdff dff_A_eHXEDivT4_2(.din(n8591), .dout(n8588));
    jdff dff_A_kG0CDKnq1_2(.din(n12371), .dout(n8591));
    jdff dff_B_lpijphA11_0(.din(n3150), .dout(n8595));
    jdff dff_B_GYqsEJOj8_0(.din(n3146), .dout(n8598));
    jdff dff_B_i6JhRNwU6_0(.din(n8598), .dout(n8601));
    jdff dff_B_gmAs5Kix2_0(.din(n8601), .dout(n8604));
    jdff dff_B_jBIxtsFT1_0(.din(n8604), .dout(n8607));
    jdff dff_B_7CYsb0fn5_0(.din(n8607), .dout(n8610));
    jdff dff_B_WgB243ov3_0(.din(n8610), .dout(n8613));
    jdff dff_B_VRcPIPAr5_0(.din(n8613), .dout(n8616));
    jdff dff_B_0IPoP4RU7_0(.din(n8616), .dout(n8619));
    jdff dff_B_gq8X0Bec3_0(.din(n8619), .dout(n8622));
    jdff dff_B_CLUWGzWf2_0(.din(n8622), .dout(n8625));
    jdff dff_B_J9GBjOcs0_0(.din(n8625), .dout(n8628));
    jdff dff_B_IqO4jrNW8_0(.din(n8628), .dout(n8631));
    jdff dff_B_JUusCXk67_0(.din(n3142), .dout(n8634));
    jdff dff_B_S7J5IsmI3_2(.din(G37), .dout(n8637));
    jdff dff_B_Rli16P8U4_2(.din(G43), .dout(n8640));
    jdff dff_B_dxC1OtnG9_2(.din(n8640), .dout(n8643));
    jdff dff_A_H9e2wXoZ0_0(.din(n8648), .dout(n8645));
    jdff dff_A_4VNwIuYC1_0(.din(n8651), .dout(n8648));
    jdff dff_A_mhPKSX9G0_0(.din(n8654), .dout(n8651));
    jdff dff_A_00N8qH0f4_0(.din(n8657), .dout(n8654));
    jdff dff_A_6Rxdd2bt0_0(.din(n8660), .dout(n8657));
    jdff dff_A_P2fmNh136_0(.din(n8663), .dout(n8660));
    jdff dff_A_7Ey6VMuo4_0(.din(n12603), .dout(n8663));
    jdff dff_A_rBWeQVvN4_0(.din(n8669), .dout(n8666));
    jdff dff_A_wE6aJrTb1_0(.din(n8672), .dout(n8669));
    jdff dff_A_h3x6bsEl5_0(.din(n8675), .dout(n8672));
    jdff dff_A_sgNgf0vX6_0(.din(n8678), .dout(n8675));
    jdff dff_A_waHlxvN38_0(.din(n8681), .dout(n8678));
    jdff dff_A_pamI7Pxv1_0(.din(n8684), .dout(n8681));
    jdff dff_A_6f9epyeH3_0(.din(n8687), .dout(n8684));
    jdff dff_A_2YFHNRle2_0(.din(n12741), .dout(n8687));
    jdff dff_B_tm7n7pgN3_0(.din(n3178), .dout(n8691));
    jdff dff_B_spxeXEEB7_0(.din(n3174), .dout(n8694));
    jdff dff_B_B0H0h72i4_0(.din(n8694), .dout(n8697));
    jdff dff_B_StLHkQiI3_0(.din(n8697), .dout(n8700));
    jdff dff_B_3PaLHpKP9_0(.din(n8700), .dout(n8703));
    jdff dff_B_euwC8bRQ4_0(.din(n8703), .dout(n8706));
    jdff dff_B_PJQewawI0_0(.din(n8706), .dout(n8709));
    jdff dff_B_DDX5Fy4I6_0(.din(n8709), .dout(n8712));
    jdff dff_B_NqcF3pch4_0(.din(n8712), .dout(n8715));
    jdff dff_B_Je3HVV2R8_0(.din(n8715), .dout(n8718));
    jdff dff_B_e9AgWHTM3_0(.din(n8718), .dout(n8721));
    jdff dff_B_bMwGzXBW6_0(.din(n3170), .dout(n8724));
    jdff dff_B_ntYLpOYK3_2(.din(G20), .dout(n8727));
    jdff dff_B_K85BdsWi9_2(.din(G76), .dout(n8730));
    jdff dff_B_l3xCiwCo2_2(.din(n8730), .dout(n8733));
    jdff dff_B_XCDHoueb2_0(.din(n3206), .dout(n8736));
    jdff dff_B_TErgr8ko2_0(.din(n8736), .dout(n8739));
    jdff dff_B_unBvVqnu6_0(.din(n3202), .dout(n8742));
    jdff dff_B_D9SjgIIo7_0(.din(n8742), .dout(n8745));
    jdff dff_B_ajTPpUqU0_0(.din(n8745), .dout(n8748));
    jdff dff_B_hQ1ZOIEw6_0(.din(n8748), .dout(n8751));
    jdff dff_B_sgHFWcFo8_0(.din(n8751), .dout(n8754));
    jdff dff_B_JyGP5icQ1_0(.din(n8754), .dout(n8757));
    jdff dff_B_u5lrbKGc5_0(.din(n8757), .dout(n8760));
    jdff dff_B_TKf1DxH57_0(.din(n8760), .dout(n8763));
    jdff dff_B_NwksgsXy5_0(.din(n3198), .dout(n8766));
    jdff dff_B_JPVxV5JX3_2(.din(G17), .dout(n8769));
    jdff dff_B_41uG2RLG8_2(.din(G73), .dout(n8772));
    jdff dff_B_SAJzS6I19_2(.din(n8772), .dout(n8775));
    jdff dff_B_DMJtnIM71_0(.din(n3234), .dout(n8778));
    jdff dff_B_nyxe27eH1_0(.din(n8778), .dout(n8781));
    jdff dff_B_J3jcYmM34_0(.din(n8781), .dout(n8784));
    jdff dff_B_O7THjFWr7_0(.din(n3230), .dout(n8787));
    jdff dff_B_GaElTtFk0_0(.din(n8787), .dout(n8790));
    jdff dff_B_dIDC2yNE2_0(.din(n8790), .dout(n8793));
    jdff dff_B_Mb9koHU65_0(.din(n8793), .dout(n8796));
    jdff dff_B_NBwEMJkl1_0(.din(n8796), .dout(n8799));
    jdff dff_B_QKeZNlHr6_0(.din(n8799), .dout(n8802));
    jdff dff_B_TZ3jdvfl1_0(.din(n3226), .dout(n8805));
    jdff dff_B_gGqDyEHP8_2(.din(G70), .dout(n8808));
    jdff dff_B_tFN5R1Mz9_2(.din(G67), .dout(n8811));
    jdff dff_B_dmDgtYiK5_2(.din(n8811), .dout(n8814));
    jdff dff_A_P2xNaJpc5_1(.din(n8819), .dout(n8816));
    jdff dff_A_np2aySLL9_1(.din(n12584), .dout(n8819));
    jdff dff_A_wHs9jq1k8_2(.din(n8825), .dout(n8822));
    jdff dff_A_4OVrbwy44_2(.din(n8828), .dout(n8825));
    jdff dff_A_oxwMc8g02_2(.din(n8831), .dout(n8828));
    jdff dff_A_ILrysShD0_2(.din(n12584), .dout(n8831));
    jdff dff_A_2SUQv1QZ1_1(.din(n12710), .dout(n8834));
    jdff dff_A_1WNx31T11_2(.din(n8840), .dout(n8837));
    jdff dff_A_GSoiYBCs5_2(.din(n12710), .dout(n8840));
    jdff dff_B_XTnXtpgM8_0(.din(n3262), .dout(n8844));
    jdff dff_B_gtS9rtlA1_0(.din(n3258), .dout(n8847));
    jdff dff_B_a4nihD729_0(.din(n8847), .dout(n8850));
    jdff dff_B_Xh8RYayb9_0(.din(n8850), .dout(n8853));
    jdff dff_B_mCRNHctH2_0(.din(n8853), .dout(n8856));
    jdff dff_B_x8zkF9130_0(.din(n8856), .dout(n8859));
    jdff dff_B_vn3QLHjX3_0(.din(n8859), .dout(n8862));
    jdff dff_B_KW5161zW1_0(.din(n8862), .dout(n8865));
    jdff dff_B_kcz1biqD4_0(.din(n8865), .dout(n8868));
    jdff dff_B_GB4tiu9b0_0(.din(n8868), .dout(n8871));
    jdff dff_B_ay1FvGnp2_0(.din(n8871), .dout(n8874));
    jdff dff_B_DhAD15Lh7_0(.din(n8874), .dout(n8877));
    jdff dff_B_W3ZZw4Cn9_0(.din(n8877), .dout(n8880));
    jdff dff_B_WjCWHaAT4_0(.din(n3254), .dout(n8883));
    jdff dff_A_BxdxAuTy3_0(.din(n8888), .dout(n8885));
    jdff dff_A_QRetefqs5_0(.din(n8891), .dout(n8888));
    jdff dff_A_0rMw0z2f3_0(.din(n8894), .dout(n8891));
    jdff dff_A_fMXsBj9m6_0(.din(n8897), .dout(n8894));
    jdff dff_A_MmLzWgdh3_0(.din(n8900), .dout(n8897));
    jdff dff_A_noo8JoPT4_0(.din(n8903), .dout(n8900));
    jdff dff_A_LzgFPlqJ2_0(.din(n12866), .dout(n8903));
    jdff dff_A_gHzBM0LF5_0(.din(n8909), .dout(n8906));
    jdff dff_A_EysPXUwI6_0(.din(n8912), .dout(n8909));
    jdff dff_A_AyI6GO7f7_0(.din(n8915), .dout(n8912));
    jdff dff_A_guqWhoe00_0(.din(n8918), .dout(n8915));
    jdff dff_A_YiYShXeA3_0(.din(n8921), .dout(n8918));
    jdff dff_A_KRV72M3l8_0(.din(n8924), .dout(n8921));
    jdff dff_A_KyShtKWw0_0(.din(n8927), .dout(n8924));
    jdff dff_A_p7tmQuyS8_0(.din(n13064), .dout(n8927));
    jdff dff_B_FHdlhyxr5_0(.din(n3294), .dout(n8931));
    jdff dff_B_P6gQ9s1P0_0(.din(n8931), .dout(n8934));
    jdff dff_B_T3z170Uf8_0(.din(n8934), .dout(n8937));
    jdff dff_B_gq0Tum2J9_0(.din(n3290), .dout(n8940));
    jdff dff_B_oBnIaTDD1_0(.din(n8940), .dout(n8943));
    jdff dff_B_TWbyM5508_0(.din(n8943), .dout(n8946));
    jdff dff_B_nXtGAaXD7_0(.din(n8946), .dout(n8949));
    jdff dff_B_uSdc2ox50_0(.din(n8949), .dout(n8952));
    jdff dff_B_W18ARSSY5_0(.din(n8952), .dout(n8955));
    jdff dff_B_UroukBto2_0(.din(n3286), .dout(n8958));
    jdff dff_B_EoeafYTF2_0(.din(n3326), .dout(n8961));
    jdff dff_B_KlIGP9566_0(.din(n8961), .dout(n8964));
    jdff dff_B_K7rIN2yn3_0(.din(n3322), .dout(n8967));
    jdff dff_B_62J7ihQl9_0(.din(n8967), .dout(n8970));
    jdff dff_B_1v5WwXJz9_0(.din(n8970), .dout(n8973));
    jdff dff_B_bxUHRyXk9_0(.din(n8973), .dout(n8976));
    jdff dff_B_kriV0NXd8_0(.din(n8976), .dout(n8979));
    jdff dff_B_c7xR3tpJ3_0(.din(n8979), .dout(n8982));
    jdff dff_B_3E2BngQZ8_0(.din(n8982), .dout(n8985));
    jdff dff_B_D7JximM67_0(.din(n8985), .dout(n8988));
    jdff dff_B_0aRS2stc2_0(.din(n3318), .dout(n8991));
    jdff dff_A_1BC24AqY8_0(.din(n9389), .dout(n8993));
    jdff dff_A_gko4YKyK2_2(.din(n8999), .dout(n8996));
    jdff dff_A_px96T8OU9_2(.din(n9002), .dout(n8999));
    jdff dff_A_E9gPA6Lu8_2(.din(n9005), .dout(n9002));
    jdff dff_A_e6UNA8IQ6_2(.din(n9389), .dout(n9005));
    jdff dff_B_BprNyinQ4_0(.din(n3358), .dout(n9009));
    jdff dff_B_OS5ZA7bL9_0(.din(n3354), .dout(n9012));
    jdff dff_B_VEjMUxYL5_0(.din(n9012), .dout(n9015));
    jdff dff_B_no1Xjybo0_0(.din(n9015), .dout(n9018));
    jdff dff_B_EmVfzZRj6_0(.din(n9018), .dout(n9021));
    jdff dff_B_1KUHvEMk1_0(.din(n9021), .dout(n9024));
    jdff dff_B_x8V8CaWD3_0(.din(n9024), .dout(n9027));
    jdff dff_B_u5SYxqAU4_0(.din(n9027), .dout(n9030));
    jdff dff_B_JaNqa41D0_0(.din(n9030), .dout(n9033));
    jdff dff_B_soNc0u147_0(.din(n9033), .dout(n9036));
    jdff dff_B_5qbHPi520_0(.din(n9036), .dout(n9039));
    jdff dff_B_xkoqWe9W8_0(.din(n3350), .dout(n9042));
    jdff dff_A_DyrteZ6p1_0(.din(n9047), .dout(n9044));
    jdff dff_A_HppuP6Js1_0(.din(n9050), .dout(n9047));
    jdff dff_A_DDViaX6f7_0(.din(n9053), .dout(n9050));
    jdff dff_A_dpyfnwzd8_0(.din(n12986), .dout(n9053));
    jdff dff_A_atiftQfm6_1(.din(n9059), .dout(n9056));
    jdff dff_A_SSmOGXFU7_1(.din(n12986), .dout(n9059));
    jdff dff_A_qNjLDCVg7_0(.din(n9065), .dout(n9062));
    jdff dff_A_fCAycZkA0_0(.din(n13193), .dout(n9065));
    jdff dff_A_cN4ywjen3_1(.din(n13193), .dout(n9068));
    jdff dff_B_OgIeoO6B4_0(.din(n3390), .dout(n9072));
    jdff dff_B_En1prRs44_0(.din(n3386), .dout(n9075));
    jdff dff_B_fwlSjpo56_0(.din(n9075), .dout(n9078));
    jdff dff_B_upMTLFBi1_0(.din(n9078), .dout(n9081));
    jdff dff_B_QNvj0gwz1_0(.din(n9081), .dout(n9084));
    jdff dff_B_ZhMkt2bJ3_0(.din(n9084), .dout(n9087));
    jdff dff_B_9dOWhQTQ3_0(.din(n9087), .dout(n9090));
    jdff dff_B_zThJXWQv4_0(.din(n9090), .dout(n9093));
    jdff dff_B_vl0nWUn87_0(.din(n9093), .dout(n9096));
    jdff dff_B_8NuyTHxS8_0(.din(n9096), .dout(n9099));
    jdff dff_B_KanJafkY3_0(.din(n9099), .dout(n9102));
    jdff dff_B_70WijCaP4_0(.din(n9102), .dout(n9105));
    jdff dff_B_GzcXBlx84_0(.din(n9105), .dout(n9108));
    jdff dff_B_5KDeyqNZ2_0(.din(n3382), .dout(n9111));
    jdff dff_B_JcnLwAmB3_2(.din(G170), .dout(n9114));
    jdff dff_B_XcbrhrKy6_2(.din(G200), .dout(n9117));
    jdff dff_B_YbWxK6xW4_2(.din(n9117), .dout(n9120));
    jdff dff_A_9eKJdbRh4_0(.din(n9125), .dout(n9122));
    jdff dff_A_sLqpRWvs9_0(.din(n9128), .dout(n9125));
    jdff dff_A_GgBhcmtO9_0(.din(n9131), .dout(n9128));
    jdff dff_A_47zHNPzp2_0(.din(n9134), .dout(n9131));
    jdff dff_A_deeyw11t2_0(.din(n9137), .dout(n9134));
    jdff dff_A_6Vi4GMIZ8_0(.din(n9140), .dout(n9137));
    jdff dff_A_kMyjH4IQ1_0(.din(n14711), .dout(n9140));
    jdff dff_B_ZpKwYiag7_0(.din(n2245), .dout(n9144));
    jdff dff_B_AP3B4fjv9_0(.din(n9144), .dout(n9147));
    jdff dff_B_BOcGSZIL7_0(.din(n9147), .dout(n9150));
    jdff dff_B_RgcqJiYQ9_0(.din(n9150), .dout(n9153));
    jdff dff_B_COUyQcJW3_0(.din(n9153), .dout(n9156));
    jdff dff_B_6PCInH3y0_0(.din(n9156), .dout(n9159));
    jdff dff_B_eKL3llTz4_0(.din(n2241), .dout(n9162));
    jdff dff_B_FDZowcrK5_0(.din(n9162), .dout(n9165));
    jdff dff_B_MC7EYT0u1_1(.din(G52), .dout(n9168));
    jdff dff_B_TXDqdpuD8_1(.din(n9168), .dout(n9171));
    jdff dff_B_6x1nUjZV6_0(.din(n788), .dout(n9174));
    jdff dff_B_9iNE9XXP0_1(.din(n757), .dout(n9177));
    jdff dff_A_RR97Thn17_0(.din(n9182), .dout(n9179));
    jdff dff_A_7nm7N9su5_0(.din(n9185), .dout(n9182));
    jdff dff_A_3MCc1XmU7_0(.din(n9188), .dout(n9185));
    jdff dff_A_waTVUbUa8_0(.din(n9191), .dout(n9188));
    jdff dff_A_Rr2iFJ0p9_0(.din(n9194), .dout(n9191));
    jdff dff_A_exPsBILN4_0(.din(n9197), .dout(n9194));
    jdff dff_A_mLONIbjn9_0(.din(n9200), .dout(n9197));
    jdff dff_A_a9Qm4DtW7_0(.din(n16322), .dout(n9200));
    jdff dff_B_fq9rhGuf4_0(.din(n2447), .dout(n9204));
    jdff dff_B_PuyzAVSH1_0(.din(n9204), .dout(n9207));
    jdff dff_B_8mQ0XSkc9_0(.din(n9207), .dout(n9210));
    jdff dff_B_R7YEhzvu4_0(.din(n9210), .dout(n9213));
    jdff dff_B_PR0izhPs7_0(.din(n9213), .dout(n9216));
    jdff dff_B_ULeG9tiY5_0(.din(n9216), .dout(n9219));
    jdff dff_B_Vk0JY3u23_0(.din(n9219), .dout(n9222));
    jdff dff_B_94rHWRBM0_0(.din(n9222), .dout(n9225));
    jdff dff_B_1cLKOKWl7_0(.din(n2443), .dout(n9228));
    jdff dff_B_WUOp7OYO9_0(.din(n9228), .dout(n9231));
    jdff dff_B_M89nhxxV1_1(.din(G122), .dout(n9234));
    jdff dff_B_Pvx58Jyu8_1(.din(n9234), .dout(n9237));
    jdff dff_B_FGBLF5RG1_0(.din(n926), .dout(n9240));
    jdff dff_B_4NDoHUfP4_1(.din(n895), .dout(n9243));
    jdff dff_B_iNlZN9jk3_1(.din(n2391), .dout(n9246));
    jdff dff_B_5zist2W43_1(.din(n9246), .dout(n9249));
    jdff dff_B_EmjnAZEq6_1(.din(n9249), .dout(n9252));
    jdff dff_B_pHWzAP7Y9_1(.din(n9252), .dout(n9255));
    jdff dff_B_AuHxWxW40_1(.din(n9255), .dout(n9258));
    jdff dff_B_73bDIewy7_1(.din(n9258), .dout(n9261));
    jdff dff_B_IomaU9x00_0(.din(n3422), .dout(n9264));
    jdff dff_B_b8GBKIl80_0(.din(n9264), .dout(n9267));
    jdff dff_B_CNjIMwUF5_0(.din(n9267), .dout(n9270));
    jdff dff_B_iljtuNsl0_0(.din(n3418), .dout(n9273));
    jdff dff_B_OKBLelgK2_0(.din(n9273), .dout(n9276));
    jdff dff_B_aOxlDQ062_0(.din(n9276), .dout(n9279));
    jdff dff_B_yOorlP4o7_0(.din(n9279), .dout(n9282));
    jdff dff_B_PZcdhNna8_0(.din(n9282), .dout(n9285));
    jdff dff_B_wahLog2R8_0(.din(n9285), .dout(n9288));
    jdff dff_B_Dria40VK9_0(.din(n3414), .dout(n9291));
    jdff dff_B_rhmpJRnq2_2(.din(G158), .dout(n9294));
    jdff dff_B_Kcwo7PKd4_2(.din(G188), .dout(n9297));
    jdff dff_B_oPu1wzDG3_2(.din(n9297), .dout(n9300));
    jdff dff_B_wTdfFCYR9_0(.din(n2072), .dout(n9303));
    jdff dff_B_Dplxahew3_0(.din(n9303), .dout(n9306));
    jdff dff_B_0cZsRaBs4_1(.din(G129), .dout(n9309));
    jdff dff_B_UlMVrDl49_1(.din(n9309), .dout(n9312));
    jdff dff_A_y5ATf2KU7_1(.din(n656), .dout(n9314));
    jdff dff_B_hpRNacob3_0(.din(n652), .dout(n9318));
    jdff dff_B_ME1rjpGW3_1(.din(n618), .dout(n9321));
    jdff dff_A_zE2BDkb14_0(.din(n11337), .dout(n9323));
    jdff dff_B_1cDh0C0P1_0(.din(n2564), .dout(n9327));
    jdff dff_B_e6H0owVM2_0(.din(n9327), .dout(n9330));
    jdff dff_B_XV6f11p15_0(.din(n9330), .dout(n9333));
    jdff dff_B_i7cpOCT88_0(.din(n9333), .dout(n9336));
    jdff dff_B_2NrrkCob0_0(.din(n2560), .dout(n9339));
    jdff dff_B_WEhjN6ji8_0(.din(n9339), .dout(n9342));
    jdff dff_B_HkCz8Ird5_1(.din(G126), .dout(n9345));
    jdff dff_B_mEvSGX876_1(.din(n9345), .dout(n9348));
    jdff dff_B_NznqOe2n0_0(.din(n1018), .dout(n9351));
    jdff dff_B_9BFouGyv7_1(.din(n987), .dout(n9354));
    jdff dff_B_90uOtjj17_0(.din(n2531), .dout(n9357));
    jdff dff_A_Ovfi9hOb9_1(.din(n9362), .dout(n9359));
    jdff dff_A_g0BHYwOQ1_1(.din(n9365), .dout(n9362));
    jdff dff_A_973G9RMs0_1(.din(n9368), .dout(n9365));
    jdff dff_A_Dg47uAWB2_1(.din(n9377), .dout(n9368));
    jdff dff_A_MA2pURe37_2(.din(n9374), .dout(n9371));
    jdff dff_A_srnJSoTh0_2(.din(n9377), .dout(n9374));
    jdff dff_A_Rt3k4Nc34_0(.din(n9380), .dout(n9377));
    jdff dff_A_UZDXURbz1_0(.din(n9383), .dout(n9380));
    jdff dff_A_kZc9yHur4_0(.din(n9386), .dout(n9383));
    jdff dff_A_rYHWvkE08_0(.din(n16679), .dout(n9386));
    jdff dff_A_fGYOpEif8_1(.din(n9392), .dout(n9389));
    jdff dff_A_AHSc45R73_1(.din(n9395), .dout(n9392));
    jdff dff_A_hKm7mnYD0_1(.din(n9398), .dout(n9395));
    jdff dff_A_E3CF4CRp0_1(.din(n16679), .dout(n9398));
    jdff dff_B_joGhvehh8_0(.din(n3454), .dout(n9402));
    jdff dff_B_reDfHA2s8_0(.din(n9402), .dout(n9405));
    jdff dff_B_3ZpPZ9th1_0(.din(n3450), .dout(n9408));
    jdff dff_B_zi3z1JL30_0(.din(n9408), .dout(n9411));
    jdff dff_B_MY3JNuaJ7_0(.din(n9411), .dout(n9414));
    jdff dff_B_PFdWbYIz0_0(.din(n9414), .dout(n9417));
    jdff dff_B_CgAU9tAa9_0(.din(n9417), .dout(n9420));
    jdff dff_B_SIQJrTRL8_0(.din(n9420), .dout(n9423));
    jdff dff_B_t6ibS3ha3_0(.din(n9423), .dout(n9426));
    jdff dff_B_q1U8qdc83_0(.din(n9426), .dout(n9429));
    jdff dff_B_htxaFz5i3_0(.din(n3446), .dout(n9432));
    jdff dff_B_Jwib4FT85_2(.din(G152), .dout(n9435));
    jdff dff_B_nx8Dlb4J8_2(.din(G155), .dout(n9438));
    jdff dff_B_tyClrbYL5_2(.din(n9438), .dout(n9441));
    jdff dff_B_qGUnuodJ7_0(.din(n2334), .dout(n9444));
    jdff dff_B_folb1ScY3_0(.din(n9444), .dout(n9447));
    jdff dff_B_ItJBMpig6_0(.din(n2330), .dout(n9450));
    jdff dff_B_qQWnhljy2_0(.din(n9450), .dout(n9453));
    jdff dff_B_PgOv85E25_1(.din(G119), .dout(n9456));
    jdff dff_B_oO4A8jg59_1(.din(n9456), .dout(n9459));
    jdff dff_B_90sOMuAW5_0(.din(n830), .dout(n9462));
    jdff dff_B_AHuoukWT8_1(.din(n799), .dout(n9465));
    jdff dff_A_wy6D8lKC3_0(.din(n9470), .dout(n9467));
    jdff dff_A_SKuI1rEA3_0(.din(n9473), .dout(n9470));
    jdff dff_A_aaSUKXGg5_0(.din(n9476), .dout(n9473));
    jdff dff_A_sW34QoFa6_0(.din(n9479), .dout(n9476));
    jdff dff_A_J2Ts6Yvv4_0(.din(n9482), .dout(n9479));
    jdff dff_A_9oh8lctW9_0(.din(n9642), .dout(n9482));
    jdff dff_B_Y7QT4HVk9_0(.din(n2523), .dout(n9486));
    jdff dff_B_V597U4Y40_0(.din(n9486), .dout(n9489));
    jdff dff_B_FUXuW4ch9_0(.din(n9489), .dout(n9492));
    jdff dff_B_xfw8lBFP9_0(.din(n9492), .dout(n9495));
    jdff dff_B_UWRP0Y5A5_0(.din(n9495), .dout(n9498));
    jdff dff_B_u9EAxGG46_0(.din(n2519), .dout(n9501));
    jdff dff_B_Y8q27l6j4_0(.din(n9501), .dout(n9504));
    jdff dff_B_cytzVKcL3_1(.din(G127), .dout(n9507));
    jdff dff_B_A0F7fsOW6_1(.din(n9507), .dout(n9510));
    jdff dff_A_8VKltBBU2_1(.din(n888), .dout(n9512));
    jdff dff_B_YwJWY0nX7_0(.din(n884), .dout(n9516));
    jdff dff_B_v0xWcDdw6_1(.din(n853), .dout(n9519));
    jdff dff_B_ZNFHKvU31_0(.din(n3486), .dout(n9522));
    jdff dff_B_6hklEctc2_0(.din(n3482), .dout(n9525));
    jdff dff_B_DuHVaRYy5_0(.din(n9525), .dout(n9528));
    jdff dff_B_WS8OTYFr8_0(.din(n9528), .dout(n9531));
    jdff dff_B_hLJV7IoA7_0(.din(n9531), .dout(n9534));
    jdff dff_B_lgFfUvub0_0(.din(n9534), .dout(n9537));
    jdff dff_B_PhJv75Xw4_0(.din(n9537), .dout(n9540));
    jdff dff_B_wPp1weZE4_0(.din(n9540), .dout(n9543));
    jdff dff_B_hUShEWNF6_0(.din(n9543), .dout(n9546));
    jdff dff_B_y8teBY6p8_0(.din(n9546), .dout(n9549));
    jdff dff_B_tntgAJsr9_0(.din(n9549), .dout(n9552));
    jdff dff_B_1vcrToXD2_0(.din(n3478), .dout(n9555));
    jdff dff_B_Yql3Al7D3_2(.din(G146), .dout(n9558));
    jdff dff_B_eeyDiJgY2_2(.din(G149), .dout(n9561));
    jdff dff_B_uqpvHaIJ6_2(.din(n9561), .dout(n9564));
    jdff dff_A_B0n1OQAi3_0(.din(n9569), .dout(n9566));
    jdff dff_A_63pvQg8h8_0(.din(n9572), .dout(n9569));
    jdff dff_A_BN4vH3IG5_0(.din(n9575), .dout(n9572));
    jdff dff_A_6mb7RBXC1_0(.din(n14831), .dout(n9575));
    jdff dff_A_64erkCvW5_1(.din(n9581), .dout(n9578));
    jdff dff_A_BCAe3P7R0_1(.din(n14831), .dout(n9581));
    jdff dff_B_S2Or8NpQ2_0(.din(n2291), .dout(n9585));
    jdff dff_B_AGGj8wiS0_0(.din(n9585), .dout(n9588));
    jdff dff_B_BAfeW1eF9_0(.din(n9588), .dout(n9591));
    jdff dff_B_35uPWueG1_0(.din(n9591), .dout(n9594));
    jdff dff_B_yl3JbdgC0_0(.din(n9594), .dout(n9597));
    jdff dff_B_J1JxYypK8_0(.din(n2284), .dout(n9600));
    jdff dff_B_AEPhoVEA0_1(.din(G130), .dout(n9603));
    jdff dff_B_eRjeDWEg4_1(.din(n9603), .dout(n9606));
    jdff dff_B_Zz6Hvt2A8_0(.din(n713), .dout(n9609));
    jdff dff_B_33ZGEYC72_1(.din(n2252), .dout(n9612));
    jdff dff_B_6NNxzr0W7_1(.din(n9612), .dout(n9615));
    jdff dff_B_8cbz5lvv5_1(.din(n9615), .dout(n9618));
    jdff dff_B_bjNjYMa54_1(.din(n9618), .dout(n9621));
    jdff dff_B_ltmbQhDK8_1(.din(n9621), .dout(n9624));
    jdff dff_A_hd1Eoys54_2(.din(n9629), .dout(n9626));
    jdff dff_A_GZRNoypF2_2(.din(n9632), .dout(n9629));
    jdff dff_A_4CavtIdX3_2(.din(n9635), .dout(n9632));
    jdff dff_A_wV0klqvI2_2(.din(n9642), .dout(n9635));
    jdff dff_B_Kk0V9Pnr3_3(.din(n1984), .dout(n9639));
    jdff dff_B_4K1igsW85_3(.din(n9639), .dout(n9642));
    jdff dff_A_sS2V6STz4_1(.din(n9647), .dout(n9644));
    jdff dff_A_sHOXtqEZ9_1(.din(n11324), .dout(n9647));
    jdff dff_A_PUPh2Q1J9_2(.din(n9653), .dout(n9650));
    jdff dff_A_bpcWVSnb9_2(.din(n9656), .dout(n9653));
    jdff dff_A_w1Xm0ZBY8_2(.din(n9659), .dout(n9656));
    jdff dff_A_p1fNNdqi8_2(.din(n11324), .dout(n9659));
    jdff dff_A_5Ni3oU0t8_0(.din(n9665), .dout(n9662));
    jdff dff_A_i86dQOnh2_0(.din(n16451), .dout(n9665));
    jdff dff_A_QwZ9RiFX5_1(.din(n16451), .dout(n9668));
    jdff dff_B_0iCX4q2L4_0(.din(n2474), .dout(n9672));
    jdff dff_B_1IUmLE8N8_0(.din(n9672), .dout(n9675));
    jdff dff_B_5MhM0mvX9_0(.din(n9675), .dout(n9678));
    jdff dff_B_PIIXsSd08_0(.din(n9678), .dout(n9681));
    jdff dff_B_yRUs2IVr8_0(.din(n9681), .dout(n9684));
    jdff dff_B_fZP1RiSL2_0(.din(n9684), .dout(n9687));
    jdff dff_B_EcPTGb4R5_0(.din(n2470), .dout(n9690));
    jdff dff_B_wCO12kb00_0(.din(n9690), .dout(n9693));
    jdff dff_B_CXvXgtDY2_1(.din(G128), .dout(n9696));
    jdff dff_B_QJsdoiVI0_1(.din(n9696), .dout(n9699));
    jdff dff_B_twvL3bjd5_0(.din(n968), .dout(n9702));
    jdff dff_B_XnnT7VXe0_1(.din(n937), .dout(n9705));
    jdff dff_B_orm6dmTT0_0(.din(n2412), .dout(n9708));
    jdff dff_A_S3A9iaE13_0(.din(n9713), .dout(n9710));
    jdff dff_A_krEBoHMt1_0(.din(n9716), .dout(n9713));
    jdff dff_A_zbBOPd4Q6_0(.din(n9719), .dout(n9716));
    jdff dff_A_SL3qSCfQ3_0(.din(n11856), .dout(n9719));
    jdff dff_B_rZlufikp0_0(.din(n3553), .dout(n9723));
    jdff dff_B_Z8QgmcpH3_0(.din(n9723), .dout(n9726));
    jdff dff_B_Sx6bZPfX9_0(.din(n9726), .dout(n9729));
    jdff dff_B_tURWSTxm3_0(.din(n9729), .dout(n9732));
    jdff dff_B_EJIcXACC0_0(.din(n9732), .dout(n9735));
    jdff dff_B_RLQnn9YY0_0(.din(n9735), .dout(n9738));
    jdff dff_B_R1vwRNSd9_0(.din(n9738), .dout(n9741));
    jdff dff_B_KkfVonDU0_0(.din(n9741), .dout(n9744));
    jdff dff_B_UydwmAn19_0(.din(n9744), .dout(n9747));
    jdff dff_B_KFyg94CR6_0(.din(n9747), .dout(n9750));
    jdff dff_B_aieW1T711_0(.din(n9750), .dout(n9753));
    jdff dff_B_w7QhIpOV3_0(.din(n9753), .dout(n9756));
    jdff dff_B_JFohs4FV4_1(.din(n3526), .dout(n9759));
    jdff dff_B_b8ZWHRwQ6_1(.din(n9759), .dout(n9762));
    jdff dff_B_i6tiRbtz5_1(.din(n9762), .dout(n9765));
    jdff dff_B_azQH0x1a7_1(.din(n9765), .dout(n9768));
    jdff dff_B_FsbrXkvc7_1(.din(n9768), .dout(n9771));
    jdff dff_B_n1caYDXs8_1(.din(n3534), .dout(n9774));
    jdff dff_B_jOuKGlAG2_0(.din(n3512), .dout(n9777));
    jdff dff_B_XofCy3am5_0(.din(n9777), .dout(n9780));
    jdff dff_B_aYYrDuJW6_0(.din(n9780), .dout(n9783));
    jdff dff_B_PBruMV9M2_0(.din(n9783), .dout(n9786));
    jdff dff_B_HpBSRuLH3_0(.din(n9786), .dout(n9789));
    jdff dff_B_5aYLOKsi5_0(.din(n9789), .dout(n9792));
    jdff dff_B_tIFftIpk1_0(.din(n9792), .dout(n9795));
    jdff dff_B_zNJNcfz89_0(.din(n9795), .dout(n9798));
    jdff dff_B_ICcObu3u6_0(.din(n9798), .dout(n9801));
    jdff dff_B_MojCcEFQ2_0(.din(n9801), .dout(n9804));
    jdff dff_B_1z8FhPUv6_0(.din(n9804), .dout(n9807));
    jdff dff_B_Jp3qyDQ02_0(.din(n9807), .dout(n9810));
    jdff dff_B_5nfTkvUg1_0(.din(n9810), .dout(n9813));
    jdff dff_B_7N6eNxPt9_0(.din(n9813), .dout(n9816));
    jdff dff_B_MWWNPNaA3_0(.din(n9816), .dout(n9819));
    jdff dff_B_FMrwp04V2_0(.din(n9819), .dout(n9822));
    jdff dff_B_J0YdLulo1_1(.din(n3501), .dout(n9825));
    jdff dff_A_K6SzOKp15_0(.din(n9830), .dout(n9827));
    jdff dff_A_qeirXqOk5_0(.din(n9833), .dout(n9830));
    jdff dff_A_osSimo5V6_0(.din(n3504), .dout(n9833));
    jdff dff_A_aKgV9xIY9_0(.din(n9839), .dout(n9836));
    jdff dff_A_sGtT0UpU5_0(.din(n9842), .dout(n9839));
    jdff dff_A_wtCkzWpC0_0(.din(n9845), .dout(n9842));
    jdff dff_A_d2klbvkf6_0(.din(n9848), .dout(n9845));
    jdff dff_A_j4F8Q4Q48_0(.din(G3717), .dout(n9848));
    jdff dff_A_KupFvMek0_0(.din(n9854), .dout(n9851));
    jdff dff_A_YMQddjrZ0_0(.din(n9857), .dout(n9854));
    jdff dff_A_neHuwbZB1_0(.din(n9860), .dout(n9857));
    jdff dff_A_vCMXz4iL1_0(.din(G3724), .dout(n9860));
    jdff dff_A_bkx6wXmx2_2(.din(n9866), .dout(n9863));
    jdff dff_A_INHrCEno2_2(.din(n9869), .dout(n9866));
    jdff dff_A_yAzh50XK3_2(.din(n9872), .dout(n9869));
    jdff dff_A_fRLBZb3v8_2(.din(n9875), .dout(n9872));
    jdff dff_A_HVpc9jXd3_2(.din(n9878), .dout(n9875));
    jdff dff_A_URkEzGnw4_2(.din(n9881), .dout(n9878));
    jdff dff_A_DBvuUKK06_2(.din(n9884), .dout(n9881));
    jdff dff_A_8RgLcLau1_2(.din(n9887), .dout(n9884));
    jdff dff_A_T83pYknB7_2(.din(n9890), .dout(n9887));
    jdff dff_A_8zQhIFMF0_2(.din(n9893), .dout(n9890));
    jdff dff_A_GIzrlDgr3_2(.din(n9896), .dout(n9893));
    jdff dff_A_bbsteKd83_2(.din(n9899), .dout(n9896));
    jdff dff_A_9wEnWf2n6_2(.din(n9902), .dout(n9899));
    jdff dff_A_007DtaO53_2(.din(n9905), .dout(n9902));
    jdff dff_A_afgfJBNd1_2(.din(n9908), .dout(n9905));
    jdff dff_A_awaVXosT6_2(.din(n9911), .dout(n9908));
    jdff dff_A_NZxTyMrq2_2(.din(n9914), .dout(n9911));
    jdff dff_A_Y3km0hto5_2(.din(G3724), .dout(n9914));
    jdff dff_A_CyhbJpPf8_0(.din(n9920), .dout(n9917));
    jdff dff_A_mp7Tnzcw8_0(.din(n9923), .dout(n9920));
    jdff dff_A_gsfJ6xKn8_0(.din(n9926), .dout(n9923));
    jdff dff_A_O9AgyIXz0_0(.din(n9929), .dout(n9926));
    jdff dff_A_oOM8QH7N3_0(.din(n9932), .dout(n9929));
    jdff dff_A_GoffM0QW2_0(.din(n9935), .dout(n9932));
    jdff dff_A_YEkxEUIG5_0(.din(n9938), .dout(n9935));
    jdff dff_A_yt364Pk02_0(.din(n9941), .dout(n9938));
    jdff dff_A_ALYqXm6s4_0(.din(n9944), .dout(n9941));
    jdff dff_A_YzTymrLW3_0(.din(n9947), .dout(n9944));
    jdff dff_A_zzsJyB2j0_0(.din(n9950), .dout(n9947));
    jdff dff_A_ZG2Bd2je4_0(.din(n9953), .dout(n9950));
    jdff dff_A_de4oxTsm6_0(.din(n9963), .dout(n9953));
    jdff dff_B_eXbFNvuK9_2(.din(G132), .dout(n9957));
    jdff dff_B_PQ2AeFZf3_2(.din(n9957), .dout(n9960));
    jdff dff_B_i0Dq756B2_2(.din(n9960), .dout(n9963));
    jdff dff_B_9S8cjbQD0_1(.din(n3663), .dout(n9966));
    jdff dff_B_U0OOsFzQ1_0(.din(n3683), .dout(n9969));
    jdff dff_B_Fk7TrJzz6_0(.din(n9969), .dout(n9972));
    jdff dff_B_NHXjAi4F9_0(.din(n3675), .dout(n9975));
    jdff dff_A_66KJWVwp8_0(.din(n313), .dout(n9977));
    jdff dff_B_UFlG5cKM3_1(.din(n1645), .dout(n9981));
    jdff dff_A_AS70YKql5_0(.din(n1704), .dout(n9983));
    jdff dff_B_QE8FytI96_1(.din(n1680), .dout(n9987));
    jdff dff_B_FhiAzXBB6_1(.din(n2600), .dout(n9990));
    jdff dff_B_g1TD5Row9_1(.din(n2607), .dout(n9993));
    jdff dff_B_JEPeCu9J0_1(.din(n9993), .dout(n9996));
    jdff dff_B_ZG2jwuz38_0(.din(n2610), .dout(n9999));
    jdff dff_B_zQ4MytPc7_1(.din(n2603), .dout(n10002));
    jdff dff_B_jyM7J1ZV9_0(.din(n2588), .dout(n10005));
    jdff dff_A_7RobHvig9_0(.din(G369), .dout(n10007));
    jdff dff_A_jNOtSQy00_0(.din(n10013), .dout(n10010));
    jdff dff_A_3vlUtqyv9_0(.din(n10016), .dout(n10013));
    jdff dff_A_XwwuUsln0_0(.din(n1509), .dout(n10016));
    jdff dff_B_MvjSQb1U2_0(.din(n2653), .dout(n10020));
    jdff dff_A_9cjRjcFv5_0(.din(G289), .dout(n10022));
    jdff dff_B_Ut5Bnd300_0(.din(n3815), .dout(n10026));
    jdff dff_B_bhGgs7uv5_0(.din(n10026), .dout(n10029));
    jdff dff_B_UFJ4mJEx3_0(.din(n10029), .dout(n10032));
    jdff dff_B_z9LDfLam6_0(.din(n10032), .dout(n10035));
    jdff dff_B_pi18C67K0_0(.din(n10035), .dout(n10038));
    jdff dff_B_58hRtFy36_0(.din(n10038), .dout(n10041));
    jdff dff_B_s7n5lhpd8_0(.din(n10041), .dout(n10044));
    jdff dff_B_dtPFA2SD7_0(.din(n10044), .dout(n10047));
    jdff dff_B_9bPkADha1_0(.din(n10047), .dout(n10050));
    jdff dff_B_Yh1o87DF4_0(.din(n10050), .dout(n10053));
    jdff dff_B_q9XTkk1d1_0(.din(n10053), .dout(n10056));
    jdff dff_B_GU6O5mJw0_0(.din(n10056), .dout(n10059));
    jdff dff_B_QNxPHZKg8_0(.din(n10059), .dout(n10062));
    jdff dff_B_Wc5IvLvh3_0(.din(n10062), .dout(n10065));
    jdff dff_B_FlTFRELI9_0(.din(n10065), .dout(n10068));
    jdff dff_B_aEuozjhT5_0(.din(n10068), .dout(n10071));
    jdff dff_B_I2ermMkl7_0(.din(n10071), .dout(n10074));
    jdff dff_B_2C2LaIa98_0(.din(n3811), .dout(n10077));
    jdff dff_B_K8TlxGVZ4_0(.din(n3843), .dout(n10080));
    jdff dff_B_vTLCDkIb0_0(.din(n10080), .dout(n10083));
    jdff dff_B_Gpl903cN2_0(.din(n10083), .dout(n10086));
    jdff dff_B_OtsaWbz08_0(.din(n10086), .dout(n10089));
    jdff dff_B_ZhQRZYta7_0(.din(n10089), .dout(n10092));
    jdff dff_B_ofde5ZOi0_0(.din(n10092), .dout(n10095));
    jdff dff_B_b4G56N331_0(.din(n10095), .dout(n10098));
    jdff dff_B_uPHCEmRC4_0(.din(n10098), .dout(n10101));
    jdff dff_B_F12qWcb15_0(.din(n10101), .dout(n10104));
    jdff dff_B_nU5g4WdW9_0(.din(n10104), .dout(n10107));
    jdff dff_B_X5lc8ERA2_0(.din(n10107), .dout(n10110));
    jdff dff_B_E4BG8Ayw5_0(.din(n10110), .dout(n10113));
    jdff dff_B_IOi2av3N4_0(.din(n10113), .dout(n10116));
    jdff dff_B_DZcULegl0_0(.din(n10116), .dout(n10119));
    jdff dff_B_Qx7oNdWy9_0(.din(n10119), .dout(n10122));
    jdff dff_B_0ztLduFz5_0(.din(n10122), .dout(n10125));
    jdff dff_B_nsPRMNxz1_0(.din(n10125), .dout(n10128));
    jdff dff_B_Ih13jZBk8_0(.din(n3839), .dout(n10131));
    jdff dff_B_skpGvuxw4_2(.din(G106), .dout(n10134));
    jdff dff_B_G5rMUXF48_2(.din(G109), .dout(n10137));
    jdff dff_B_pc46jYw56_2(.din(n10137), .dout(n10140));
    jdff dff_B_xiEtWRdJ3_0(.din(n3874), .dout(n10143));
    jdff dff_B_0QXWl8xb1_0(.din(n10143), .dout(n10146));
    jdff dff_B_axFCVXAq9_0(.din(n10146), .dout(n10149));
    jdff dff_B_q14bpZdM0_0(.din(n10149), .dout(n10152));
    jdff dff_B_xKfuQ16J7_0(.din(n10152), .dout(n10155));
    jdff dff_B_XW5a9qpS3_0(.din(n10155), .dout(n10158));
    jdff dff_B_qoNtuyfN5_0(.din(n10158), .dout(n10161));
    jdff dff_B_lo5eZZYj4_0(.din(n10161), .dout(n10164));
    jdff dff_B_wR7cML9x6_0(.din(n10164), .dout(n10167));
    jdff dff_B_rw2nfGOk0_0(.din(n10167), .dout(n10170));
    jdff dff_B_sZjXSQc00_0(.din(n10170), .dout(n10173));
    jdff dff_B_1MYmZ2Hh8_0(.din(n10173), .dout(n10176));
    jdff dff_B_vZJ4MQiT0_0(.din(n10176), .dout(n10179));
    jdff dff_B_zU4wzDf07_0(.din(n10179), .dout(n10182));
    jdff dff_B_2rdPzQxt5_0(.din(n10182), .dout(n10185));
    jdff dff_B_wsrvTRFU1_0(.din(n10185), .dout(n10188));
    jdff dff_B_bKng4ZYj7_0(.din(n3870), .dout(n10191));
    jdff dff_B_7sDRp8Pe6_0(.din(n3908), .dout(n10194));
    jdff dff_B_jcLLwElZ8_0(.din(n10194), .dout(n10197));
    jdff dff_B_X3W3I4CG0_0(.din(n10197), .dout(n10200));
    jdff dff_B_bxdHV3Tb7_0(.din(n10200), .dout(n10203));
    jdff dff_B_Y7YCJUoX5_0(.din(n10203), .dout(n10206));
    jdff dff_B_qlpAoWjL2_0(.din(n10206), .dout(n10209));
    jdff dff_B_7MN0tEj44_0(.din(n10209), .dout(n10212));
    jdff dff_B_xl0qGUAI6_0(.din(n10212), .dout(n10215));
    jdff dff_B_rM0t2XlX6_0(.din(n10215), .dout(n10218));
    jdff dff_B_FAavZQ1G2_0(.din(n10218), .dout(n10221));
    jdff dff_B_4j68Ncvl4_0(.din(n10221), .dout(n10224));
    jdff dff_B_vwzFit9Q6_0(.din(n10224), .dout(n10227));
    jdff dff_B_Hj7tOlfS8_0(.din(n10227), .dout(n10230));
    jdff dff_B_nBFTz95a8_0(.din(n10230), .dout(n10233));
    jdff dff_B_CiOblOqN6_0(.din(n10233), .dout(n10236));
    jdff dff_B_bOm6xuOr3_0(.din(n10236), .dout(n10239));
    jdff dff_B_uwUSbe004_0(.din(n3904), .dout(n10242));
    jdff dff_A_dkRHlgvt0_2(.din(n12212), .dout(n10244));
    jdff dff_A_ZgzYrzSU2_2(.din(n12338), .dout(n10247));
    jdff dff_B_qYJGFmw80_0(.din(n3942), .dout(n10251));
    jdff dff_B_0xGmt1ef9_0(.din(n10251), .dout(n10254));
    jdff dff_B_WlUJvoLS4_0(.din(n10254), .dout(n10257));
    jdff dff_B_lRZuuHgY9_0(.din(n10257), .dout(n10260));
    jdff dff_B_f1jKh4Xk8_0(.din(n10260), .dout(n10263));
    jdff dff_B_hnUKu0HQ6_0(.din(n10263), .dout(n10266));
    jdff dff_B_jFCmLIkr3_0(.din(n10266), .dout(n10269));
    jdff dff_B_zEnMY9dx2_0(.din(n10269), .dout(n10272));
    jdff dff_B_Tg6LPpdP0_0(.din(n10272), .dout(n10275));
    jdff dff_B_gP81Hn0u5_0(.din(n10275), .dout(n10278));
    jdff dff_B_o0wuvb1b9_0(.din(n10278), .dout(n10281));
    jdff dff_B_IIGwLfn26_0(.din(n10281), .dout(n10284));
    jdff dff_B_ohzHHHUB2_0(.din(n10284), .dout(n10287));
    jdff dff_B_q77aGSrk7_0(.din(n10287), .dout(n10290));
    jdff dff_B_t94d85kX8_0(.din(n10290), .dout(n10293));
    jdff dff_B_5jWzyvJG7_0(.din(n3938), .dout(n10296));
    jdff dff_B_NypKMHDv5_0(.din(n3970), .dout(n10299));
    jdff dff_B_PoebvJ2P8_0(.din(n10299), .dout(n10302));
    jdff dff_B_8fRSbgka8_0(.din(n10302), .dout(n10305));
    jdff dff_B_UmrBnTNH2_0(.din(n10305), .dout(n10308));
    jdff dff_B_v9cFAZLn5_0(.din(n10308), .dout(n10311));
    jdff dff_B_zqDTnKjs4_0(.din(n10311), .dout(n10314));
    jdff dff_B_4vle1Qcn3_0(.din(n10314), .dout(n10317));
    jdff dff_B_k16y28oq0_0(.din(n10317), .dout(n10320));
    jdff dff_B_uv1yIhmW3_0(.din(n10320), .dout(n10323));
    jdff dff_B_2jKjYMzD8_0(.din(n10323), .dout(n10326));
    jdff dff_B_ywD1xsZl0_0(.din(n10326), .dout(n10329));
    jdff dff_B_Z0ns3pPN8_0(.din(n10329), .dout(n10332));
    jdff dff_B_g4KtRWBn3_0(.din(n10332), .dout(n10335));
    jdff dff_B_1DRwYKOB2_0(.din(n10335), .dout(n10338));
    jdff dff_B_77g5Gz7d0_0(.din(n10338), .dout(n10341));
    jdff dff_B_LhUW3Ydi0_0(.din(n10341), .dout(n10344));
    jdff dff_B_Izl0K9OX4_0(.din(n3966), .dout(n10347));
    jdff dff_B_zwPJdQEF4_2(.din(G49), .dout(n10350));
    jdff dff_B_eXvMRe1b0_2(.din(G46), .dout(n10353));
    jdff dff_B_SYbYFckq7_2(.din(n10353), .dout(n10356));
    jdff dff_B_8a1wdmuh6_0(.din(n3998), .dout(n10359));
    jdff dff_B_LcHVNjN99_0(.din(n10359), .dout(n10362));
    jdff dff_B_18MsEnw70_0(.din(n10362), .dout(n10365));
    jdff dff_B_HVS95MvC7_0(.din(n10365), .dout(n10368));
    jdff dff_B_GGddtJoi9_0(.din(n10368), .dout(n10371));
    jdff dff_B_fal9RzBR4_0(.din(n10371), .dout(n10374));
    jdff dff_B_L6FrlyfN6_0(.din(n10374), .dout(n10377));
    jdff dff_B_OxoekeWa1_0(.din(n10377), .dout(n10380));
    jdff dff_B_2Kc6ThxV7_0(.din(n10380), .dout(n10383));
    jdff dff_B_YI2taczn0_0(.din(n10383), .dout(n10386));
    jdff dff_B_Fj3NFwt24_0(.din(n10386), .dout(n10389));
    jdff dff_B_uNgBiU0g9_0(.din(n10389), .dout(n10392));
    jdff dff_B_vRurAE3o3_0(.din(n10392), .dout(n10395));
    jdff dff_B_UrgNl8Ee5_0(.din(n10395), .dout(n10398));
    jdff dff_B_OftxRVgy5_0(.din(n10398), .dout(n10401));
    jdff dff_B_aiw9eHOp9_0(.din(n10401), .dout(n10404));
    jdff dff_B_jlLPp9Vx4_0(.din(n3994), .dout(n10407));
    jdff dff_B_mOQjkljC0_2(.din(G103), .dout(n10410));
    jdff dff_B_zoqcHgRF3_2(.din(G100), .dout(n10413));
    jdff dff_B_0gLVztIc0_2(.din(n10413), .dout(n10416));
    jdff dff_A_YZB8mdmT1_2(.din(n12551), .dout(n10418));
    jdff dff_A_WCC2ZLwE1_2(.din(n12677), .dout(n10421));
    jdff dff_B_pBf9AXCt4_0(.din(n4026), .dout(n10425));
    jdff dff_B_yMNdH2HB6_0(.din(n10425), .dout(n10428));
    jdff dff_B_hjkvwDCd0_0(.din(n10428), .dout(n10431));
    jdff dff_B_AcGrsj9n5_0(.din(n10431), .dout(n10434));
    jdff dff_B_xrmpRsv10_0(.din(n10434), .dout(n10437));
    jdff dff_B_3dgRN1Um7_0(.din(n10437), .dout(n10440));
    jdff dff_B_mWlX1zib4_0(.din(n10440), .dout(n10443));
    jdff dff_B_XBWApV9K6_0(.din(n10443), .dout(n10446));
    jdff dff_B_QfUT9LvJ3_0(.din(n10446), .dout(n10449));
    jdff dff_B_ciLEGZ418_0(.din(n10449), .dout(n10452));
    jdff dff_B_AlFxUvzv6_0(.din(n10452), .dout(n10455));
    jdff dff_B_HeI2mYQu0_0(.din(n10455), .dout(n10458));
    jdff dff_B_MziJslA06_0(.din(n10458), .dout(n10461));
    jdff dff_B_VVs6pJHk9_0(.din(n10461), .dout(n10464));
    jdff dff_B_pcFZ3uXV4_0(.din(n10464), .dout(n10467));
    jdff dff_B_vi4xFXql7_0(.din(n4022), .dout(n10470));
    jdff dff_B_cQ9zOYqq2_2(.din(G40), .dout(n10473));
    jdff dff_B_QWTeqsKZ6_2(.din(G91), .dout(n10476));
    jdff dff_B_jN6unUfh7_2(.din(n10476), .dout(n10479));
    jdff dff_B_Ow9FdZNy8_0(.din(n4054), .dout(n10482));
    jdff dff_B_YGPUoZBU2_0(.din(n10482), .dout(n10485));
    jdff dff_B_rNED4cpP6_0(.din(n10485), .dout(n10488));
    jdff dff_B_ttIkTcL76_0(.din(n10488), .dout(n10491));
    jdff dff_B_83KDtTui9_0(.din(n10491), .dout(n10494));
    jdff dff_B_hUY0udmf3_0(.din(n10494), .dout(n10497));
    jdff dff_B_hEznpjwG7_0(.din(n10497), .dout(n10500));
    jdff dff_B_wcQSsuKc3_0(.din(n10500), .dout(n10503));
    jdff dff_B_RcKiMlGo0_0(.din(n10503), .dout(n10506));
    jdff dff_B_7EqxGuFx2_0(.din(n10506), .dout(n10509));
    jdff dff_B_v6JDwg0L9_0(.din(n10509), .dout(n10512));
    jdff dff_B_OKspzJNu7_0(.din(n10512), .dout(n10515));
    jdff dff_B_APgepRj83_0(.din(n10515), .dout(n10518));
    jdff dff_B_NgUwY59h6_0(.din(n10518), .dout(n10521));
    jdff dff_B_bdxp7AcU3_0(.din(n10521), .dout(n10524));
    jdff dff_B_fis0PEsW9_0(.din(n4050), .dout(n10527));
    jdff dff_A_y1kofuVU5_0(.din(n10532), .dout(n10529));
    jdff dff_A_bZhs7fic4_0(.din(n10535), .dout(n10532));
    jdff dff_A_H5oXzNSF8_0(.din(n10538), .dout(n10535));
    jdff dff_A_H3FSjW8n1_0(.din(n10541), .dout(n10538));
    jdff dff_A_ZlmiawB56_0(.din(n16631), .dout(n10541));
    jdff dff_A_qp4LGAap9_1(.din(n16631), .dout(n10544));
    jdff dff_B_agRsUJDf4_0(.din(n4086), .dout(n10548));
    jdff dff_B_ZKwsOfHf5_0(.din(n10548), .dout(n10551));
    jdff dff_B_V3uCsFml0_0(.din(n10551), .dout(n10554));
    jdff dff_B_SQHPePvO3_0(.din(n10554), .dout(n10557));
    jdff dff_B_TDWBnvTb7_0(.din(n10557), .dout(n10560));
    jdff dff_B_xr8B8iLi1_0(.din(n10560), .dout(n10563));
    jdff dff_B_12MprNB32_0(.din(n10563), .dout(n10566));
    jdff dff_B_5aEKSf3m8_0(.din(n10566), .dout(n10569));
    jdff dff_B_RkBc9UVD7_0(.din(n10569), .dout(n10572));
    jdff dff_B_3hqkoWtI1_0(.din(n10572), .dout(n10575));
    jdff dff_B_sIJUYtiF0_0(.din(n10575), .dout(n10578));
    jdff dff_B_6nGtx7Bc5_0(.din(n10578), .dout(n10581));
    jdff dff_B_7UyEt8Gt1_0(.din(n10581), .dout(n10584));
    jdff dff_B_wjNWKAFj7_0(.din(n10584), .dout(n10587));
    jdff dff_B_EBRwlS4T6_0(.din(n10587), .dout(n10590));
    jdff dff_B_V85onpWG4_0(.din(n10590), .dout(n10593));
    jdff dff_B_294IO92r3_0(.din(n4082), .dout(n10596));
    jdff dff_B_d0YDtxRG3_0(.din(n4118), .dout(n10599));
    jdff dff_B_LAXbZkme6_0(.din(n10599), .dout(n10602));
    jdff dff_B_wMMrjdzF3_0(.din(n10602), .dout(n10605));
    jdff dff_B_Tv3AhgpP7_0(.din(n10605), .dout(n10608));
    jdff dff_B_cbFc7pic9_0(.din(n10608), .dout(n10611));
    jdff dff_B_8GxulXDB4_0(.din(n10611), .dout(n10614));
    jdff dff_B_dM2C0V3V7_0(.din(n10614), .dout(n10617));
    jdff dff_B_g5vUnsM18_0(.din(n10617), .dout(n10620));
    jdff dff_B_KOhDaaUz2_0(.din(n10620), .dout(n10623));
    jdff dff_B_O3LfvDXL3_0(.din(n10623), .dout(n10626));
    jdff dff_B_xyw0L8UL6_0(.din(n10626), .dout(n10629));
    jdff dff_B_AAfTTh1A4_0(.din(n10629), .dout(n10632));
    jdff dff_B_ViAWt65H6_0(.din(n10632), .dout(n10635));
    jdff dff_B_MkvfGRyR6_0(.din(n10635), .dout(n10638));
    jdff dff_B_cssxxx1u9_0(.din(n10638), .dout(n10641));
    jdff dff_B_C1YjVtUI7_0(.din(n10641), .dout(n10644));
    jdff dff_B_FfSLbWuY1_0(.din(n4114), .dout(n10647));
    jdff dff_A_7OW5y9l72_0(.din(n12938), .dout(n10649));
    jdff dff_A_l4jMXvw94_1(.din(n12938), .dout(n10652));
    jdff dff_A_PHBE6jlE2_0(.din(n13142), .dout(n10655));
    jdff dff_A_o45GCSCM4_1(.din(n13142), .dout(n10658));
    jdff dff_B_gVdEtFX19_0(.din(n4150), .dout(n10662));
    jdff dff_B_Ba0686lj8_0(.din(n10662), .dout(n10665));
    jdff dff_B_qsfq8MbL0_0(.din(n10665), .dout(n10668));
    jdff dff_B_KfOZ8Leu1_0(.din(n10668), .dout(n10671));
    jdff dff_B_vj1MW3nq9_0(.din(n10671), .dout(n10674));
    jdff dff_B_uS61SSR74_0(.din(n10674), .dout(n10677));
    jdff dff_B_C9ky7vOl1_0(.din(n10677), .dout(n10680));
    jdff dff_B_R2CeI2Jc3_0(.din(n10680), .dout(n10683));
    jdff dff_B_kMat4lox3_0(.din(n10683), .dout(n10686));
    jdff dff_B_Rdg9HmST9_0(.din(n10686), .dout(n10689));
    jdff dff_B_JhlFtZgN5_0(.din(n10689), .dout(n10692));
    jdff dff_B_3CmVi0QK0_0(.din(n10692), .dout(n10695));
    jdff dff_B_yBsCen7m0_0(.din(n10695), .dout(n10698));
    jdff dff_B_V5ZrAPuN6_0(.din(n10698), .dout(n10701));
    jdff dff_B_xyVYWRYK9_0(.din(n10701), .dout(n10704));
    jdff dff_B_s55vGzNJ3_0(.din(n10704), .dout(n10707));
    jdff dff_B_UhZT5YK20_0(.din(n10707), .dout(n10710));
    jdff dff_B_KImXdIga2_0(.din(n4146), .dout(n10713));
    jdff dff_A_RQQIh7vn0_0(.din(n11468), .dout(n10715));
    jdff dff_B_ZmFCOJy13_0(.din(n4182), .dout(n10719));
    jdff dff_B_JbI7LX1H9_0(.din(n10719), .dout(n10722));
    jdff dff_B_LMESYq2w5_0(.din(n10722), .dout(n10725));
    jdff dff_B_8hAu5rcr9_0(.din(n10725), .dout(n10728));
    jdff dff_B_a35Fo7iV8_0(.din(n10728), .dout(n10731));
    jdff dff_B_t3yeZgE34_0(.din(n10731), .dout(n10734));
    jdff dff_B_4xMKYaLx1_0(.din(n10734), .dout(n10737));
    jdff dff_B_7PEwpT1r2_0(.din(n10737), .dout(n10740));
    jdff dff_B_zu2voKMB9_0(.din(n10740), .dout(n10743));
    jdff dff_B_QUWFna4i9_0(.din(n10743), .dout(n10746));
    jdff dff_B_5Bds0IZW2_0(.din(n10746), .dout(n10749));
    jdff dff_B_CIdUXag39_0(.din(n10749), .dout(n10752));
    jdff dff_B_vmB6lXpv2_0(.din(n10752), .dout(n10755));
    jdff dff_B_SWDiZyBP0_0(.din(n10755), .dout(n10758));
    jdff dff_B_ccTWhB2x9_0(.din(n10758), .dout(n10761));
    jdff dff_B_OKMz4WVo9_0(.din(n4178), .dout(n10764));
    jdff dff_B_SGUhAMb97_2(.din(G173), .dout(n10767));
    jdff dff_B_IFxkz3Y08_2(.din(G203), .dout(n10770));
    jdff dff_B_mLxJD7f59_2(.din(n10770), .dout(n10773));
    jdff dff_B_I9S9Xa0x6_0(.din(n3656), .dout(n10776));
    jdff dff_B_TEtLmidp4_0(.din(n10776), .dout(n10779));
    jdff dff_B_96xzDBIs6_0(.din(n10779), .dout(n10782));
    jdff dff_B_LHpPA1Wf7_0(.din(n10782), .dout(n10785));
    jdff dff_B_cFYJGVhW7_0(.din(n10785), .dout(n10788));
    jdff dff_B_RMXQNnOq9_0(.din(n10788), .dout(n10791));
    jdff dff_B_L4qQWu689_0(.din(n10791), .dout(n10794));
    jdff dff_B_kmG4DrdP9_0(.din(n10794), .dout(n10797));
    jdff dff_B_AQUBKamq2_0(.din(n10797), .dout(n10800));
    jdff dff_B_E1ByTHYL4_0(.din(n3652), .dout(n10803));
    jdff dff_B_62huH6Nq1_0(.din(n10803), .dout(n10806));
    jdff dff_B_3epKLyCT9_1(.din(G112), .dout(n10809));
    jdff dff_B_tYfQVzEI9_1(.din(n10809), .dout(n10812));
    jdff dff_B_17aiqjGc4_0(.din(n3791), .dout(n10815));
    jdff dff_B_dSejLMxx2_0(.din(n10815), .dout(n10818));
    jdff dff_B_nek2bSjm6_0(.din(n10818), .dout(n10821));
    jdff dff_B_IX8EgRQH2_0(.din(n10821), .dout(n10824));
    jdff dff_B_xbHkbq0I8_0(.din(n10824), .dout(n10827));
    jdff dff_B_UnPCY6Db0_0(.din(n10827), .dout(n10830));
    jdff dff_B_dihwUXjS5_0(.din(n10830), .dout(n10833));
    jdff dff_B_gCnKLI5i2_0(.din(n10833), .dout(n10836));
    jdff dff_B_9CBb133i7_0(.din(n10836), .dout(n10839));
    jdff dff_B_jGhB8Mmf3_0(.din(n10839), .dout(n10842));
    jdff dff_B_p23c7erm3_0(.din(n3787), .dout(n10845));
    jdff dff_B_kWzdq82a2_0(.din(n10845), .dout(n10848));
    jdff dff_B_0TVAYJPD2_1(.din(G113), .dout(n10851));
    jdff dff_B_AKDvo7Ba7_1(.din(n10851), .dout(n10854));
    jdff dff_B_2wflkQor3_0(.din(n1194), .dout(n10857));
    jdff dff_B_YdcdSCpG9_1(.din(n1163), .dout(n10860));
    jdff dff_B_09Q8taF07_0(.din(n4214), .dout(n10863));
    jdff dff_B_zEuw58Vs5_0(.din(n10863), .dout(n10866));
    jdff dff_B_qtFTJ7YN5_0(.din(n10866), .dout(n10869));
    jdff dff_B_0rmgxtLS1_0(.din(n10869), .dout(n10872));
    jdff dff_B_dYrKAl9E6_0(.din(n10872), .dout(n10875));
    jdff dff_B_EJQTvFzO7_0(.din(n10875), .dout(n10878));
    jdff dff_B_BiTMPZqi6_0(.din(n10878), .dout(n10881));
    jdff dff_B_dqkJ1ncm3_0(.din(n10881), .dout(n10884));
    jdff dff_B_fmMG05vF3_0(.din(n10884), .dout(n10887));
    jdff dff_B_AtuYmRCA6_0(.din(n10887), .dout(n10890));
    jdff dff_B_IFHSWs6i4_0(.din(n10890), .dout(n10893));
    jdff dff_B_d8G8CC2Z5_0(.din(n10893), .dout(n10896));
    jdff dff_B_aj8h4fjM8_0(.din(n10896), .dout(n10899));
    jdff dff_B_GURgKlrr4_0(.din(n10899), .dout(n10902));
    jdff dff_B_qCbrYods6_0(.din(n10902), .dout(n10905));
    jdff dff_B_lXYnlb5b3_0(.din(n10905), .dout(n10908));
    jdff dff_B_SAWpM6fQ5_0(.din(n4210), .dout(n10911));
    jdff dff_B_MAJmmH5t1_2(.din(G167), .dout(n10914));
    jdff dff_B_50RCKjQP1_2(.din(G197), .dout(n10917));
    jdff dff_B_cFW4n59S5_2(.din(n10917), .dout(n10920));
    jdff dff_B_LIqQJyqB7_0(.din(n3630), .dout(n10923));
    jdff dff_B_154GA88v8_0(.din(n10923), .dout(n10926));
    jdff dff_B_scoLKQWQ0_0(.din(n10926), .dout(n10929));
    jdff dff_B_H5TTfpr02_0(.din(n10929), .dout(n10932));
    jdff dff_B_WVwjElLV1_0(.din(n10932), .dout(n10935));
    jdff dff_B_r8tieEPh9_0(.din(n10935), .dout(n10938));
    jdff dff_B_xGpnWdoj3_0(.din(n10938), .dout(n10941));
    jdff dff_B_fKnP5ZTG4_0(.din(n10941), .dout(n10944));
    jdff dff_B_zpKo9Ccc5_0(.din(n10944), .dout(n10947));
    jdff dff_B_vJHcfLve3_0(.din(n10947), .dout(n10950));
    jdff dff_B_3J5EAi6i6_0(.din(n3626), .dout(n10953));
    jdff dff_B_1QghGSTZ5_0(.din(n10953), .dout(n10956));
    jdff dff_B_odjM5rvn3_1(.din(G116), .dout(n10959));
    jdff dff_B_h2p3nyxB3_1(.din(n10959), .dout(n10962));
    jdff dff_A_sUW6gcWQ9_1(.din(n2835), .dout(n10964));
    jdff dff_B_quMq9nbg5_1(.din(n2819), .dout(n10968));
    jdff dff_B_sQCErxne2_1(.din(n10968), .dout(n10971));
    jdff dff_B_4EsNKvRA1_1(.din(n10971), .dout(n10974));
    jdff dff_B_l8XGactB8_1(.din(n10974), .dout(n10977));
    jdff dff_B_xlzh8Ftl9_1(.din(n10977), .dout(n10980));
    jdff dff_B_c0G0nXkd0_1(.din(n10980), .dout(n10983));
    jdff dff_B_kZeNUo0G9_1(.din(n10983), .dout(n10986));
    jdff dff_B_3nxzTJoj7_1(.din(n10986), .dout(n10989));
    jdff dff_B_kOVmyXKi0_1(.din(n10989), .dout(n10992));
    jdff dff_B_udGqIPxm7_1(.din(n10992), .dout(n10995));
    jdff dff_B_IMe2uchO1_0(.din(n3765), .dout(n10998));
    jdff dff_B_ZReIIt4W8_0(.din(n10998), .dout(n11001));
    jdff dff_B_gw0ZtexQ4_0(.din(n11001), .dout(n11004));
    jdff dff_B_7sCawKEX8_0(.din(n11004), .dout(n11007));
    jdff dff_B_8Ui3d48h8_0(.din(n11007), .dout(n11010));
    jdff dff_B_mSSl9zLJ1_0(.din(n11010), .dout(n11013));
    jdff dff_B_sNTc23mc7_0(.din(n11013), .dout(n11016));
    jdff dff_B_9oJ52C180_0(.din(n11016), .dout(n11019));
    jdff dff_B_MqaT0KJJ5_0(.din(n11019), .dout(n11022));
    jdff dff_B_AQXaAoau3_0(.din(n11022), .dout(n11025));
    jdff dff_B_xAXaJ5Ik2_0(.din(n11025), .dout(n11028));
    jdff dff_B_pxnY8ccd7_0(.din(n3761), .dout(n11031));
    jdff dff_B_7PZywBut2_0(.din(n11031), .dout(n11034));
    jdff dff_B_Nj5vdTif5_1(.din(G53), .dout(n11037));
    jdff dff_B_StV1voEx0_1(.din(n11037), .dout(n11040));
    jdff dff_B_gG2uUQz25_0(.din(n1106), .dout(n11043));
    jdff dff_B_ETgeSkvN4_1(.din(n1075), .dout(n11046));
    jdff dff_B_ixPsF8PX5_1(.din(n2753), .dout(n11049));
    jdff dff_B_4qSErFbZ5_1(.din(n11049), .dout(n11052));
    jdff dff_B_55kHWLt07_1(.din(n11052), .dout(n11055));
    jdff dff_B_PdoLO2ui9_1(.din(n11055), .dout(n11058));
    jdff dff_B_Uo6Ck4sD7_1(.din(n11058), .dout(n11061));
    jdff dff_B_Us86aFVR4_1(.din(n11061), .dout(n11064));
    jdff dff_B_mXczXv536_1(.din(n11064), .dout(n11067));
    jdff dff_B_sf9LzMDB0_1(.din(n11067), .dout(n11070));
    jdff dff_B_c7gxiID30_1(.din(n11070), .dout(n11073));
    jdff dff_B_TffRr9w90_1(.din(n11073), .dout(n11076));
    jdff dff_B_3c94yB1b0_1(.din(n2756), .dout(n11079));
    jdff dff_B_fpTMEgEi4_1(.din(n11079), .dout(n11082));
    jdff dff_B_eeznKk6L0_1(.din(n11082), .dout(n11085));
    jdff dff_B_ConUEDM16_1(.din(n11085), .dout(n11088));
    jdff dff_B_qsOYPMWr4_1(.din(n11088), .dout(n11091));
    jdff dff_B_VbZ4XuZP0_1(.din(n11091), .dout(n11094));
    jdff dff_B_P1WrViCA7_1(.din(n11094), .dout(n11097));
    jdff dff_B_iBWYpPYu7_1(.din(n11097), .dout(n11100));
    jdff dff_B_e5HQDqVp5_1(.din(n11100), .dout(n11103));
    jdff dff_A_sAzoij892_1(.din(n11108), .dout(n11105));
    jdff dff_A_6FYOdVxK6_1(.din(n11111), .dout(n11108));
    jdff dff_A_zNPmARhV5_1(.din(n11114), .dout(n11111));
    jdff dff_A_77DusoA61_1(.din(n11117), .dout(n11114));
    jdff dff_A_aLhqdgZU3_1(.din(n11120), .dout(n11117));
    jdff dff_A_Vgr5vevl1_1(.din(n11123), .dout(n11120));
    jdff dff_A_vb2M1OE24_1(.din(n11126), .dout(n11123));
    jdff dff_A_Ck6oxcC35_1(.din(n11129), .dout(n11126));
    jdff dff_A_RBGRznVJ7_1(.din(n11132), .dout(n11129));
    jdff dff_A_zeRLM1kf4_1(.din(n11135), .dout(n11132));
    jdff dff_A_BmECUsk12_1(.din(n11138), .dout(n11135));
    jdff dff_A_Gu5nNEwY7_1(.din(n11141), .dout(n11138));
    jdff dff_A_FBNMLUe16_1(.din(n11337), .dout(n11141));
    jdff dff_A_nDfkBzeK5_2(.din(n11147), .dout(n11144));
    jdff dff_A_9RebKp3i9_2(.din(n11150), .dout(n11147));
    jdff dff_A_gNbujCMb7_2(.din(n11153), .dout(n11150));
    jdff dff_A_aLH5F6Tt6_2(.din(n11156), .dout(n11153));
    jdff dff_A_Pimr12Am7_2(.din(n11159), .dout(n11156));
    jdff dff_A_ElQe45RG5_2(.din(n11162), .dout(n11159));
    jdff dff_A_2s2YT0uI2_2(.din(n11165), .dout(n11162));
    jdff dff_A_btSBnyTP2_2(.din(n11168), .dout(n11165));
    jdff dff_A_BPkgQXW11_2(.din(n11171), .dout(n11168));
    jdff dff_A_SQAQH26V5_2(.din(n11174), .dout(n11171));
    jdff dff_A_iNS2XPFK1_2(.din(n11177), .dout(n11174));
    jdff dff_A_L5frsO004_2(.din(n11337), .dout(n11177));
    jdff dff_B_9pLJ2O540_0(.din(n4246), .dout(n11181));
    jdff dff_B_cPWzW0kk4_0(.din(n11181), .dout(n11184));
    jdff dff_B_Xe9zhxh66_0(.din(n11184), .dout(n11187));
    jdff dff_B_7iguyQVm5_0(.din(n11187), .dout(n11190));
    jdff dff_B_RNLWmLJJ1_0(.din(n11190), .dout(n11193));
    jdff dff_B_RHF8iTjG5_0(.din(n11193), .dout(n11196));
    jdff dff_B_pQW52dv74_0(.din(n11196), .dout(n11199));
    jdff dff_B_7y1vDWQp2_0(.din(n11199), .dout(n11202));
    jdff dff_B_5vVcP5lv2_0(.din(n11202), .dout(n11205));
    jdff dff_B_Bm4FV72o3_0(.din(n11205), .dout(n11208));
    jdff dff_B_j0If32eX7_0(.din(n11208), .dout(n11211));
    jdff dff_B_CjZodt2l6_0(.din(n11211), .dout(n11214));
    jdff dff_B_DLpxs9L61_0(.din(n11214), .dout(n11217));
    jdff dff_B_yqIm284c6_0(.din(n11217), .dout(n11220));
    jdff dff_B_Bbjyg1EH7_0(.din(n11220), .dout(n11223));
    jdff dff_B_RyyWYobz7_0(.din(n11223), .dout(n11226));
    jdff dff_B_powhZxEO6_0(.din(n4242), .dout(n11229));
    jdff dff_B_TvkVAIn21_2(.din(G164), .dout(n11232));
    jdff dff_B_14vpiaKB5_2(.din(G194), .dout(n11235));
    jdff dff_B_7lMbWqIo5_2(.din(n11235), .dout(n11238));
    jdff dff_B_B84uG7bX8_0(.din(n3607), .dout(n11241));
    jdff dff_B_QjU99fHA3_0(.din(n11241), .dout(n11244));
    jdff dff_B_ucHpOF5h4_0(.din(n11244), .dout(n11247));
    jdff dff_B_Ym1Q9bcb1_0(.din(n11247), .dout(n11250));
    jdff dff_B_ncHijzMR4_0(.din(n11250), .dout(n11253));
    jdff dff_B_y0ZkcAHI7_0(.din(n11253), .dout(n11256));
    jdff dff_B_pY4kvoBt2_0(.din(n11256), .dout(n11259));
    jdff dff_B_TvlAC35e3_0(.din(n11259), .dout(n11262));
    jdff dff_B_Mlmerch91_0(.din(n11262), .dout(n11265));
    jdff dff_B_pehWNw4f6_0(.din(n11265), .dout(n11268));
    jdff dff_B_KrP1yuHQ9_0(.din(n11268), .dout(n11271));
    jdff dff_B_marBBmw55_0(.din(n3600), .dout(n11274));
    jdff dff_B_HXk0kOAM5_1(.din(G121), .dout(n11277));
    jdff dff_B_uKr8CYGs6_1(.din(n11277), .dout(n11280));
    jdff dff_A_aeevJOVS0_0(.din(n11285), .dout(n11282));
    jdff dff_A_vEyg9jp74_0(.din(n11288), .dout(n11285));
    jdff dff_A_X6QMuLAm1_0(.din(n11291), .dout(n11288));
    jdff dff_A_q9i9WFuA3_0(.din(n11300), .dout(n11291));
    jdff dff_A_SBknElrP1_2(.din(n11297), .dout(n11294));
    jdff dff_A_YlD1YxIp1_2(.din(n11300), .dout(n11297));
    jdff dff_A_H1qLvIgG7_1(.din(n11303), .dout(n11300));
    jdff dff_A_xsOeO7oV5_1(.din(n11306), .dout(n11303));
    jdff dff_A_ylCN2lH88_1(.din(n11309), .dout(n11306));
    jdff dff_A_8yOW4PUZ0_1(.din(n11312), .dout(n11309));
    jdff dff_A_y7CO8UH03_1(.din(n11315), .dout(n11312));
    jdff dff_A_qzHdiVqZ7_1(.din(n11318), .dout(n11315));
    jdff dff_A_EnI1yzei1_1(.din(n11321), .dout(n11318));
    jdff dff_A_UQoh7LGe2_1(.din(n11337), .dout(n11321));
    jdff dff_A_wOf1Cfte0_2(.din(n11327), .dout(n11324));
    jdff dff_A_N3h0DbEd0_2(.din(n11330), .dout(n11327));
    jdff dff_A_wRFxOKzz0_2(.din(n11333), .dout(n11330));
    jdff dff_A_a3B1miSq9_2(.din(n11337), .dout(n11333));
    jdff dff_B_qXzrlhWH2_3(.din(n1998), .dout(n11337));
    jdff dff_A_qNY8BP3v7_0(.din(n11342), .dout(n11339));
    jdff dff_A_UXajs5TU9_0(.din(n11345), .dout(n11342));
    jdff dff_A_aPAD6atK6_0(.din(n11348), .dout(n11345));
    jdff dff_A_WBxupp7Q1_0(.din(n11351), .dout(n11348));
    jdff dff_A_n4a7JNKr9_0(.din(n11354), .dout(n11351));
    jdff dff_A_sTj0VN4c4_0(.din(n11357), .dout(n11354));
    jdff dff_A_e0JYmab19_0(.din(n11360), .dout(n11357));
    jdff dff_A_wDe8DPcc0_0(.din(n1995), .dout(n11360));
    jdff dff_A_SqI2yV546_1(.din(n11366), .dout(n11363));
    jdff dff_A_3Vi918I32_1(.din(n11369), .dout(n11366));
    jdff dff_A_gU6XlNYE1_1(.din(n1995), .dout(n11369));
    jdff dff_A_H5bf7n1u2_0(.din(n14783), .dout(n11372));
    jdff dff_A_ITNR949C7_1(.din(n14783), .dout(n11375));
    jdff dff_B_S9J7nqW47_0(.din(n3739), .dout(n11379));
    jdff dff_B_qSC0jK4B7_0(.din(n11379), .dout(n11382));
    jdff dff_B_74MEXcp64_0(.din(n11382), .dout(n11385));
    jdff dff_B_XNwsMo0y7_0(.din(n11385), .dout(n11388));
    jdff dff_B_yNmVYCKB9_0(.din(n11388), .dout(n11391));
    jdff dff_B_9U6ylI2J2_0(.din(n11391), .dout(n11394));
    jdff dff_B_XdZik20e3_0(.din(n11394), .dout(n11397));
    jdff dff_B_vMziX8uU1_0(.din(n11397), .dout(n11400));
    jdff dff_B_r7ZKzvHx2_0(.din(n11400), .dout(n11403));
    jdff dff_B_9DeFJJmY7_0(.din(n11403), .dout(n11406));
    jdff dff_B_WPzhHrAb9_0(.din(n11406), .dout(n11409));
    jdff dff_B_PqJq7Mgt4_0(.din(n3732), .dout(n11412));
    jdff dff_B_XGAPpf743_0(.din(n11412), .dout(n11415));
    jdff dff_B_Nm4EO94P3_1(.din(G114), .dout(n11418));
    jdff dff_B_vNPPy6ed3_1(.din(n11418), .dout(n11421));
    jdff dff_B_jFICK1UL1_3(.din(n2061), .dout(n11424));
    jdff dff_B_rUp8ULsw4_3(.din(n11424), .dout(n11427));
    jdff dff_A_BsgYYTw75_1(.din(n2009), .dout(n11429));
    jdff dff_B_Bb8vETym4_0(.din(n1236), .dout(n11433));
    jdff dff_B_GertBESm2_3(.din(G3548), .dout(n11436));
    jdff dff_B_SCzYglrG4_1(.din(n1205), .dout(n11439));
    jdff dff_A_fYU173FL6_0(.din(n16400), .dout(n11441));
    jdff dff_A_tjHVlKCN6_1(.din(n16400), .dout(n11444));
    jdff dff_A_383ZEy6I1_0(.din(n11453), .dout(n11447));
    jdff dff_A_ju5dP4BX9_1(.din(n11453), .dout(n11450));
    jdff dff_A_y0ZRGQTF0_0(.din(n11456), .dout(n11453));
    jdff dff_A_sKZThTtb6_0(.din(n11459), .dout(n11456));
    jdff dff_A_q4R3ZE6d8_0(.din(n11462), .dout(n11459));
    jdff dff_A_ZCPtQnaG6_0(.din(n11465), .dout(n11462));
    jdff dff_A_so03MYB81_0(.din(n16631), .dout(n11465));
    jdff dff_A_a9J6yTKK2_1(.din(n11471), .dout(n11468));
    jdff dff_A_ZJQjY5Xt2_1(.din(n11474), .dout(n11471));
    jdff dff_A_9IoQ8PG53_1(.din(n11477), .dout(n11474));
    jdff dff_A_HjS9J4X52_1(.din(n11480), .dout(n11477));
    jdff dff_A_Fl8KFQKn2_1(.din(n11483), .dout(n11480));
    jdff dff_A_2NRd1JdT9_1(.din(n16631), .dout(n11483));
    jdff dff_B_n7cutjcq9_0(.din(n4278), .dout(n11487));
    jdff dff_B_yptsFa2p8_0(.din(n11487), .dout(n11490));
    jdff dff_B_JRsmjG7t2_0(.din(n11490), .dout(n11493));
    jdff dff_B_dZSZV8M57_0(.din(n11493), .dout(n11496));
    jdff dff_B_BSzS8LU70_0(.din(n11496), .dout(n11499));
    jdff dff_B_JVHhIBho1_0(.din(n11499), .dout(n11502));
    jdff dff_B_plbfaqeX3_0(.din(n11502), .dout(n11505));
    jdff dff_B_7eWOYkPS2_0(.din(n11505), .dout(n11508));
    jdff dff_B_gKVHduvz1_0(.din(n11508), .dout(n11511));
    jdff dff_B_JV9dXuVZ5_0(.din(n11511), .dout(n11514));
    jdff dff_B_jeGq64yM1_0(.din(n11514), .dout(n11517));
    jdff dff_B_9pGaziJu7_0(.din(n11517), .dout(n11520));
    jdff dff_B_aV5fYulz2_0(.din(n11520), .dout(n11523));
    jdff dff_B_sLKrHYsW7_0(.din(n11523), .dout(n11526));
    jdff dff_B_quMSMqcC0_0(.din(n11526), .dout(n11529));
    jdff dff_B_ZUaMsc4b2_0(.din(n11529), .dout(n11532));
    jdff dff_B_AM3vBMxa2_0(.din(n11532), .dout(n11535));
    jdff dff_B_nXPPc2nM8_0(.din(n4274), .dout(n11538));
    jdff dff_B_wnoB62px8_2(.din(G161), .dout(n11541));
    jdff dff_B_tpfWh4pm0_2(.din(G191), .dout(n11544));
    jdff dff_B_YXrldbBk9_2(.din(n11544), .dout(n11547));
    jdff dff_B_7FRchA6w4_0(.din(n3581), .dout(n11550));
    jdff dff_B_4RhB5ZPW2_0(.din(n11550), .dout(n11553));
    jdff dff_B_7D0ylB5Q9_0(.din(n11553), .dout(n11556));
    jdff dff_B_rEAdzYBT9_0(.din(n11556), .dout(n11559));
    jdff dff_B_AhbaE4kP1_0(.din(n11559), .dout(n11562));
    jdff dff_B_u1HQjpXg7_0(.din(n11562), .dout(n11565));
    jdff dff_B_bmMGZWz43_0(.din(n11565), .dout(n11568));
    jdff dff_B_IQ4cwdyf5_0(.din(n11568), .dout(n11571));
    jdff dff_B_3Of4yyyn8_0(.din(n11571), .dout(n11574));
    jdff dff_B_ZRG9BTvk1_0(.din(n11574), .dout(n11577));
    jdff dff_B_WMfun7bd3_0(.din(n11577), .dout(n11580));
    jdff dff_B_aH6Nh85K3_0(.din(n11580), .dout(n11583));
    jdff dff_B_BWNbPEii0_0(.din(n11583), .dout(n11586));
    jdff dff_B_BKEKWhze3_1(.din(n3573), .dout(n11589));
    jdff dff_B_FE6uwSmS0_1(.din(n11589), .dout(n11592));
    jdff dff_A_7EUgJjEv4_1(.din(n11756), .dout(n11594));
    jdff dff_A_BrrDWsJJ5_0(.din(n11601), .dout(n11597));
    jdff dff_B_k7ccmGjA3_2(.din(G123), .dout(n11601));
    jdff dff_B_BCyhDCpA1_0(.din(n2147), .dout(n11604));
    jdff dff_B_JbPk5Cbw3_0(.din(n2117), .dout(n11607));
    jdff dff_B_t0QenPJK3_0(.din(n11607), .dout(n11610));
    jdff dff_B_enuUWqnO6_0(.din(n11610), .dout(n11613));
    jdff dff_A_FMfDTZPu3_0(.din(n11618), .dout(n11615));
    jdff dff_A_mAXDZyS17_0(.din(n11621), .dout(n11618));
    jdff dff_A_d7HrMQip3_0(.din(n11624), .dout(n11621));
    jdff dff_A_6B2gmyQI5_0(.din(n11627), .dout(n11624));
    jdff dff_A_lCuEXdLn1_0(.din(n11630), .dout(n11627));
    jdff dff_A_LqY3TKdd0_0(.din(n11633), .dout(n11630));
    jdff dff_A_jq7VWQt19_0(.din(n11636), .dout(n11633));
    jdff dff_A_vpdtxn4N0_0(.din(G54), .dout(n11636));
    jdff dff_A_hGTaNu9B9_0(.din(n11642), .dout(n11639));
    jdff dff_A_G8LGNIc74_0(.din(n11645), .dout(n11642));
    jdff dff_A_cDwjwPSq8_0(.din(n11648), .dout(n11645));
    jdff dff_A_NB5iNk0F7_0(.din(n11651), .dout(n11648));
    jdff dff_A_1J23STzd1_0(.din(n11654), .dout(n11651));
    jdff dff_A_sIKpZPM87_0(.din(n11657), .dout(n11654));
    jdff dff_A_xo8iiHrd0_0(.din(n1973), .dout(n11657));
    jdff dff_A_fqc6Redu2_0(.din(n11663), .dout(n11660));
    jdff dff_A_8apAwvBr9_0(.din(n11666), .dout(n11663));
    jdff dff_A_Myua4Nl51_0(.din(n11669), .dout(n11666));
    jdff dff_A_XOvFG1JA5_0(.din(n11672), .dout(n11669));
    jdff dff_A_Zh3Fzkn12_0(.din(n11945), .dout(n11672));
    jdff dff_A_4cCoBgTJ8_1(.din(n11678), .dout(n11675));
    jdff dff_A_q30IOs7B4_1(.din(n11681), .dout(n11678));
    jdff dff_A_0YA5gX3L0_1(.din(n11684), .dout(n11681));
    jdff dff_A_tA6W320N7_1(.din(n11687), .dout(n11684));
    jdff dff_A_G7C3MKLi5_1(.din(n11690), .dout(n11687));
    jdff dff_A_mibvx99g4_1(.din(n11693), .dout(n11690));
    jdff dff_A_B163nOEO9_1(.din(n11696), .dout(n11693));
    jdff dff_A_B6nQ4l5Q2_1(.din(n11699), .dout(n11696));
    jdff dff_A_uvpUTQee1_1(.din(n11945), .dout(n11699));
    jdff dff_B_QB6mvxpj1_0(.din(n3710), .dout(n11703));
    jdff dff_B_bXm5ay248_0(.din(n11703), .dout(n11706));
    jdff dff_B_A0CdZTO27_0(.din(n11706), .dout(n11709));
    jdff dff_B_DMr4WauW9_0(.din(n11709), .dout(n11712));
    jdff dff_B_inQ3U82g4_0(.din(n11712), .dout(n11715));
    jdff dff_B_aYmgZKAm5_0(.din(n11715), .dout(n11718));
    jdff dff_B_KElNYV6G7_0(.din(n11718), .dout(n11721));
    jdff dff_B_DBi65DCa4_0(.din(n11721), .dout(n11724));
    jdff dff_B_VY6FUyUR8_0(.din(n11724), .dout(n11727));
    jdff dff_B_U2snLKEJ8_0(.din(n11727), .dout(n11730));
    jdff dff_B_NxDyucTm8_0(.din(n11730), .dout(n11733));
    jdff dff_B_5R5KWFjg0_0(.din(n11733), .dout(n11736));
    jdff dff_B_JUKEnXWI7_0(.din(n3706), .dout(n11739));
    jdff dff_B_lhXixDxu4_0(.din(n11739), .dout(n11742));
    jdff dff_B_2j8GxOw91_0(.din(n11742), .dout(n11745));
    jdff dff_B_20Y1p8ix0_0(.din(n11745), .dout(n11748));
    jdff dff_B_P1l3ehr71_1(.din(G115), .dout(n11751));
    jdff dff_B_9G85qHLp6_1(.din(n11751), .dout(n11754));
    jdff dff_A_frt58SoM2_0(.din(n2009), .dout(n11756));
    jdff dff_A_OYaMXLGe7_2(.din(n11762), .dout(n11759));
    jdff dff_A_YKKmtzwo8_2(.din(n11765), .dout(n11762));
    jdff dff_A_LGVtW3Qv9_2(.din(n11768), .dout(n11765));
    jdff dff_A_PvOiRHAm7_2(.din(n2009), .dout(n11768));
    jdff dff_B_V0ZC5LCV6_1(.din(n2683), .dout(n11772));
    jdff dff_B_F36k1EPQ8_1(.din(n11772), .dout(n11775));
    jdff dff_B_zTMLTtux5_1(.din(n11775), .dout(n11778));
    jdff dff_B_4RvYDFRq3_1(.din(n11778), .dout(n11781));
    jdff dff_B_Uw8cvXCJ3_1(.din(n11781), .dout(n11784));
    jdff dff_B_KyJLUTO75_1(.din(n11784), .dout(n11787));
    jdff dff_B_thd4XTy23_1(.din(n11787), .dout(n11790));
    jdff dff_B_TG5KVz8b0_1(.din(n11790), .dout(n11793));
    jdff dff_B_Jbi5ZFtY8_1(.din(n2689), .dout(n11796));
    jdff dff_B_ErAA75Sg3_1(.din(n11796), .dout(n11799));
    jdff dff_B_2xvbEX6b6_1(.din(n11799), .dout(n11802));
    jdff dff_B_rBz9tB1n5_1(.din(n11802), .dout(n11805));
    jdff dff_B_xo2Xg6bR2_1(.din(n11805), .dout(n11808));
    jdff dff_B_2TknPHmb6_1(.din(n11808), .dout(n11811));
    jdff dff_B_4BqlQqfc9_1(.din(n11811), .dout(n11814));
    jdff dff_B_5knzVkgt4_1(.din(n11814), .dout(n11817));
    jdff dff_B_nyszu3Qx9_1(.din(n11817), .dout(n11820));
    jdff dff_B_PSye6bXg7_1(.din(n11820), .dout(n11823));
    jdff dff_B_yZEvMHkQ1_0(.din(n2702), .dout(n11826));
    jdff dff_A_bDtXZSfF2_1(.din(n11831), .dout(n11828));
    jdff dff_A_aZsRZRzc4_1(.din(n11834), .dout(n11831));
    jdff dff_A_m6tBuxuy5_1(.din(n11837), .dout(n11834));
    jdff dff_A_LyJqcdhE2_1(.din(n11840), .dout(n11837));
    jdff dff_A_XQ85SI904_1(.din(n11843), .dout(n11840));
    jdff dff_A_KUzeLFZw3_1(.din(n11856), .dout(n11843));
    jdff dff_B_nm6Aqo8B0_3(.din(G4), .dout(n11847));
    jdff dff_B_iP6ndz3S4_3(.din(n11847), .dout(n11850));
    jdff dff_B_CpQk12DH3_3(.din(n11850), .dout(n11853));
    jdff dff_B_3zTcJTIs9_3(.din(n11853), .dout(n11856));
    jdff dff_B_hPJG0ldp5_2(.din(n2692), .dout(n11859));
    jdff dff_B_GP2YH0ms9_2(.din(n11859), .dout(n11862));
    jdff dff_B_mWMwWwPY5_2(.din(n11862), .dout(n11865));
    jdff dff_B_vwcFlwia3_2(.din(n11865), .dout(n11868));
    jdff dff_B_QYKlooOo9_2(.din(n11868), .dout(n11871));
    jdff dff_B_eTDh0uSx2_2(.din(n11871), .dout(n11874));
    jdff dff_B_VN8rMfKo1_2(.din(n11874), .dout(n11877));
    jdff dff_B_RbRQ8xPU8_2(.din(n11877), .dout(n11880));
    jdff dff_B_MVJDqufb2_2(.din(n11880), .dout(n11883));
    jdff dff_A_HLAl1M521_1(.din(n11888), .dout(n11885));
    jdff dff_A_xFXK0hL58_1(.din(n11891), .dout(n11888));
    jdff dff_A_VoHkmlRv2_1(.din(n11906), .dout(n11891));
    jdff dff_A_PssrBKtE0_2(.din(n11897), .dout(n11894));
    jdff dff_A_uE9d4O748_2(.din(n11900), .dout(n11897));
    jdff dff_A_ZDayzo5r4_2(.din(n11903), .dout(n11900));
    jdff dff_A_PRChFjBw1_2(.din(n11906), .dout(n11903));
    jdff dff_A_05wwoAWZ0_0(.din(n11909), .dout(n11906));
    jdff dff_A_CeJleYnU5_0(.din(n11912), .dout(n11909));
    jdff dff_A_KzdNH0DK9_0(.din(n11915), .dout(n11912));
    jdff dff_A_oieLvGfZ1_0(.din(n11918), .dout(n11915));
    jdff dff_A_0FC9zjOJ3_0(.din(n11921), .dout(n11918));
    jdff dff_A_h5iRJ6oW1_0(.din(n11924), .dout(n11921));
    jdff dff_A_rCFMe4uN1_0(.din(n11927), .dout(n11924));
    jdff dff_A_PKfuQANw6_0(.din(n11930), .dout(n11927));
    jdff dff_A_oKPUfezU1_0(.din(n11933), .dout(n11930));
    jdff dff_A_UXYtXNr46_0(.din(n11936), .dout(n11933));
    jdff dff_A_dhsvvXga0_0(.din(n11939), .dout(n11936));
    jdff dff_A_W1gUI3au0_0(.din(n11942), .dout(n11939));
    jdff dff_A_LoCCPFDQ2_0(.din(n1995), .dout(n11942));
    jdff dff_A_njKGqq1g9_1(.din(n11948), .dout(n11945));
    jdff dff_A_bzzNAAMX7_1(.din(n11951), .dout(n11948));
    jdff dff_A_DeQWqwRF8_1(.din(n11954), .dout(n11951));
    jdff dff_A_Hulc4xtm9_1(.din(n11957), .dout(n11954));
    jdff dff_A_vtSH9Vbn1_1(.din(n11960), .dout(n11957));
    jdff dff_A_NWZp0gGh3_1(.din(n11963), .dout(n11960));
    jdff dff_A_Xu5BlIp72_1(.din(n1995), .dout(n11963));
    jdff dff_B_hWyTCKRT3_1(.din(n4460), .dout(n11967));
    jdff dff_B_VDLvyCjj0_1(.din(n11967), .dout(n11970));
    jdff dff_B_sbds70jh7_1(.din(n11970), .dout(n11973));
    jdff dff_B_xVKvmOMW7_1(.din(n11973), .dout(n11976));
    jdff dff_B_NAl70N4K8_1(.din(n11976), .dout(n11979));
    jdff dff_B_5xB1GOzx7_1(.din(n11979), .dout(n11982));
    jdff dff_B_AoYBY6MI2_1(.din(n11982), .dout(n11985));
    jdff dff_B_TtEPmjQ46_1(.din(n11985), .dout(n11988));
    jdff dff_B_clzf3T6G8_1(.din(n11988), .dout(n11991));
    jdff dff_B_cFeYhvnw4_1(.din(n11991), .dout(n11994));
    jdff dff_B_CJ9UndW83_1(.din(n11994), .dout(n11997));
    jdff dff_B_N5MmGJLS4_1(.din(n11997), .dout(n12000));
    jdff dff_B_8DsBHhks9_1(.din(n12000), .dout(n12003));
    jdff dff_B_guLETHEL6_1(.din(n12003), .dout(n12006));
    jdff dff_B_RO1PxrYt8_1(.din(n12006), .dout(n12009));
    jdff dff_B_NlmNpPso8_1(.din(n12009), .dout(n12012));
    jdff dff_B_uTZn3X140_1(.din(n12012), .dout(n12015));
    jdff dff_B_O590Tvgi3_1(.din(n12015), .dout(n12018));
    jdff dff_B_pt4Np9lk0_1(.din(n12018), .dout(n12021));
    jdff dff_B_2fu0Yukz0_1(.din(n5051), .dout(n12024));
    jdff dff_B_XKFhEpvU7_1(.din(n12024), .dout(n12027));
    jdff dff_B_X16GS3k32_1(.din(n12027), .dout(n12030));
    jdff dff_B_lEZqV0FP4_1(.din(n12030), .dout(n12033));
    jdff dff_B_d00V3A903_1(.din(n12033), .dout(n12036));
    jdff dff_B_SiQpf2OB4_1(.din(n12036), .dout(n12039));
    jdff dff_B_37Wt5caT1_1(.din(n12039), .dout(n12042));
    jdff dff_B_isjrsp5R5_1(.din(n12042), .dout(n12045));
    jdff dff_B_3Szipj2D7_1(.din(n12045), .dout(n12048));
    jdff dff_B_2ltHrkJs4_1(.din(n12048), .dout(n12051));
    jdff dff_B_nZ2gg8PF1_1(.din(n12051), .dout(n12054));
    jdff dff_B_AxlY0AT22_1(.din(n12054), .dout(n12057));
    jdff dff_B_sqUS6HAx9_1(.din(n12057), .dout(n12060));
    jdff dff_B_xiX3QdBV9_1(.din(n12060), .dout(n12063));
    jdff dff_B_JpiBi7vB6_1(.din(n12063), .dout(n12066));
    jdff dff_B_LESUyLpb0_1(.din(n12066), .dout(n12069));
    jdff dff_B_9zXaKAsG7_1(.din(n12069), .dout(n12072));
    jdff dff_B_BYPKNXFo4_1(.din(n12072), .dout(n12075));
    jdff dff_B_bUlMydrC4_1(.din(n12075), .dout(n12078));
    jdff dff_B_Oyc7erkj0_0(.din(n5341), .dout(n12081));
    jdff dff_B_3UQXGzYe1_0(.din(n12081), .dout(n12084));
    jdff dff_B_p9iI1GCm6_0(.din(n12084), .dout(n12087));
    jdff dff_B_Fv8oce7b2_0(.din(n12087), .dout(n12090));
    jdff dff_B_xfdXn3gh8_0(.din(n12090), .dout(n12093));
    jdff dff_B_24RTbt2l6_0(.din(n12093), .dout(n12096));
    jdff dff_B_T5QHiW5g4_0(.din(n12096), .dout(n12099));
    jdff dff_B_XUHRBrMY2_0(.din(n12099), .dout(n12102));
    jdff dff_B_rM8hLnGy8_0(.din(n12102), .dout(n12105));
    jdff dff_B_8nFpynAk6_0(.din(n12105), .dout(n12108));
    jdff dff_B_6O0TcsTE8_0(.din(n12108), .dout(n12111));
    jdff dff_B_1ERHSp2e2_0(.din(n12111), .dout(n12114));
    jdff dff_B_KgQ5RStM5_0(.din(n12114), .dout(n12117));
    jdff dff_B_iQkfhazn3_0(.din(n12117), .dout(n12120));
    jdff dff_B_YxjzLB4X2_0(.din(n12120), .dout(n12123));
    jdff dff_B_A6trlIz93_0(.din(n12123), .dout(n12126));
    jdff dff_B_7CFLzJwE9_0(.din(n12126), .dout(n12129));
    jdff dff_B_Acos7NPE2_0(.din(n12129), .dout(n12132));
    jdff dff_B_pn9fF3NJ2_0(.din(n12132), .dout(n12135));
    jdff dff_B_zVkRJpEp9_0(.din(n5337), .dout(n12138));
    jdff dff_A_gDFl44Nf8_1(.din(n12143), .dout(n12140));
    jdff dff_A_QK4tJ5KJ2_1(.din(n12146), .dout(n12143));
    jdff dff_A_WTFoR4Xs3_1(.din(n12149), .dout(n12146));
    jdff dff_A_WnvQZK9R1_1(.din(n12152), .dout(n12149));
    jdff dff_A_YYBwUoaC1_1(.din(n12155), .dout(n12152));
    jdff dff_A_Vv1X4RK16_1(.din(n12158), .dout(n12155));
    jdff dff_A_6t5wCJPH9_1(.din(n12161), .dout(n12158));
    jdff dff_A_nloeYeZH8_1(.din(n12164), .dout(n12161));
    jdff dff_A_Zb1Np2Q13_1(.din(n12167), .dout(n12164));
    jdff dff_A_hOA9568S6_1(.din(n12170), .dout(n12167));
    jdff dff_A_iywbZGbf1_1(.din(n12173), .dout(n12170));
    jdff dff_A_TgEIV9iS0_1(.din(n12176), .dout(n12173));
    jdff dff_A_y3HvpBwO3_1(.din(n12179), .dout(n12176));
    jdff dff_A_wr4dtUjX9_1(.din(n12264), .dout(n12179));
    jdff dff_A_rKVaqn901_2(.din(n12185), .dout(n12182));
    jdff dff_A_ldK5lY4G6_2(.din(n12188), .dout(n12185));
    jdff dff_A_681pEa5P3_2(.din(n12191), .dout(n12188));
    jdff dff_A_XDMjJR8f2_2(.din(n12194), .dout(n12191));
    jdff dff_A_SwdNfqQS8_2(.din(n12197), .dout(n12194));
    jdff dff_A_1IUCxP8Q5_2(.din(n12200), .dout(n12197));
    jdff dff_A_SjRh2TnK2_2(.din(n12203), .dout(n12200));
    jdff dff_A_wffqRqnD2_2(.din(n12206), .dout(n12203));
    jdff dff_A_9b4ItQma5_2(.din(n12209), .dout(n12206));
    jdff dff_A_AJGiieCM9_2(.din(n12264), .dout(n12209));
    jdff dff_A_Zxi2yntb3_1(.din(n12215), .dout(n12212));
    jdff dff_A_iW9kNU8j2_1(.din(n12218), .dout(n12215));
    jdff dff_A_P6fUHoeO5_1(.din(n12221), .dout(n12218));
    jdff dff_A_YyMhI7br9_1(.din(n12224), .dout(n12221));
    jdff dff_A_hFiRqPYe5_1(.din(n12227), .dout(n12224));
    jdff dff_A_9yNuijDT7_1(.din(n12230), .dout(n12227));
    jdff dff_A_J9s8QZEi9_1(.din(n12233), .dout(n12230));
    jdff dff_A_5fop84UG1_1(.din(n12236), .dout(n12233));
    jdff dff_A_ZFi2FESZ2_1(.din(n12239), .dout(n12236));
    jdff dff_A_oRQ7d04F4_1(.din(n12242), .dout(n12239));
    jdff dff_A_MsSSaf845_1(.din(n12264), .dout(n12242));
    jdff dff_A_dsfKY5Mi9_2(.din(n12264), .dout(n12245));
    jdff dff_B_Jj9PwHD67_3(.din(n2178), .dout(n12249));
    jdff dff_B_4yw7WmsD5_3(.din(n12249), .dout(n12252));
    jdff dff_B_z3NZq9r76_3(.din(n12252), .dout(n12255));
    jdff dff_B_i40G09E43_3(.din(n12255), .dout(n12258));
    jdff dff_B_BWtFMQnv4_3(.din(n12258), .dout(n12261));
    jdff dff_B_XABObqKV1_3(.din(n12261), .dout(n12264));
    jdff dff_A_09hrrOSP0_1(.din(n12269), .dout(n12266));
    jdff dff_A_ICxSbAIE1_1(.din(n12272), .dout(n12269));
    jdff dff_A_4bNrqtOu9_1(.din(n12275), .dout(n12272));
    jdff dff_A_56k5cqEv8_1(.din(n12278), .dout(n12275));
    jdff dff_A_zei0RHmK3_1(.din(n12281), .dout(n12278));
    jdff dff_A_rmTAStox6_1(.din(n12284), .dout(n12281));
    jdff dff_A_LIfvZvJn4_1(.din(n12287), .dout(n12284));
    jdff dff_A_AoZXPVz36_1(.din(n12290), .dout(n12287));
    jdff dff_A_6wYzzrQc6_1(.din(n12293), .dout(n12290));
    jdff dff_A_GJPIIFRs0_1(.din(n12296), .dout(n12293));
    jdff dff_A_d3nwqLTE2_1(.din(n12299), .dout(n12296));
    jdff dff_A_AhPdWlgx8_1(.din(n12302), .dout(n12299));
    jdff dff_A_qeOascDE5_1(.din(n12305), .dout(n12302));
    jdff dff_A_xjWfmCDl7_1(.din(n12402), .dout(n12305));
    jdff dff_A_y0oRANoW6_2(.din(n12311), .dout(n12308));
    jdff dff_A_Kzu7LfBS5_2(.din(n12314), .dout(n12311));
    jdff dff_A_ePmZYUO09_2(.din(n12317), .dout(n12314));
    jdff dff_A_6XrdGx970_2(.din(n12320), .dout(n12317));
    jdff dff_A_9HOSXcbI1_2(.din(n12323), .dout(n12320));
    jdff dff_A_v7rzEFQq9_2(.din(n12326), .dout(n12323));
    jdff dff_A_kSD2nT7G3_2(.din(n12329), .dout(n12326));
    jdff dff_A_taAU0pJb7_2(.din(n12332), .dout(n12329));
    jdff dff_A_bktD94j34_2(.din(n12335), .dout(n12332));
    jdff dff_A_S5eA9kuy6_2(.din(n12402), .dout(n12335));
    jdff dff_A_ODzzS0E23_1(.din(n12341), .dout(n12338));
    jdff dff_A_NB3Sle5t5_1(.din(n12344), .dout(n12341));
    jdff dff_A_4yarnEib1_1(.din(n12347), .dout(n12344));
    jdff dff_A_mzgCjKZS7_1(.din(n12350), .dout(n12347));
    jdff dff_A_a1MPQaHw2_1(.din(n12353), .dout(n12350));
    jdff dff_A_vcICGs300_1(.din(n12356), .dout(n12353));
    jdff dff_A_A7zNrVPA7_1(.din(n12359), .dout(n12356));
    jdff dff_A_VzlFDMJE1_1(.din(n12362), .dout(n12359));
    jdff dff_A_60iMxWrC7_1(.din(n12365), .dout(n12362));
    jdff dff_A_NlNYudBi9_1(.din(n12368), .dout(n12365));
    jdff dff_A_rbDetDgH9_1(.din(n12402), .dout(n12368));
    jdff dff_A_SX3MLxt72_2(.din(n12374), .dout(n12371));
    jdff dff_A_02duTM8P5_2(.din(n12377), .dout(n12374));
    jdff dff_A_x3tz2ruC5_2(.din(n12380), .dout(n12377));
    jdff dff_A_4S0qJLoI6_2(.din(n12402), .dout(n12380));
    jdff dff_B_zmntCGcZ5_3(.din(n2164), .dout(n12384));
    jdff dff_B_hc2jIxY07_3(.din(n12384), .dout(n12387));
    jdff dff_B_F7pcUx834_3(.din(n12387), .dout(n12390));
    jdff dff_B_SwKN3pzG4_3(.din(n12390), .dout(n12393));
    jdff dff_B_tAHh98pf8_3(.din(n12393), .dout(n12396));
    jdff dff_B_YW0PqZyk2_3(.din(n12396), .dout(n12399));
    jdff dff_B_dFN2gYon5_3(.din(n12399), .dout(n12402));
    jdff dff_A_Ts5zBysZ3_2(.din(G4088), .dout(n12404));
    jdff dff_A_Jh1PO9Ub9_1(.din(G4087), .dout(n12407));
    jdff dff_B_zaTCGnqh1_0(.din(n5369), .dout(n12411));
    jdff dff_B_PAWhwoeG8_0(.din(n12411), .dout(n12414));
    jdff dff_B_PfRReHWk3_0(.din(n12414), .dout(n12417));
    jdff dff_B_11Gsk3zY7_0(.din(n12417), .dout(n12420));
    jdff dff_B_QYWkJchj3_0(.din(n12420), .dout(n12423));
    jdff dff_B_3vcKBv499_0(.din(n12423), .dout(n12426));
    jdff dff_B_R3xUY0fx2_0(.din(n12426), .dout(n12429));
    jdff dff_B_F1YHIbtk3_0(.din(n12429), .dout(n12432));
    jdff dff_B_MGpcTcz82_0(.din(n12432), .dout(n12435));
    jdff dff_B_wlON81Hb1_0(.din(n12435), .dout(n12438));
    jdff dff_B_9LPqMGjj0_0(.din(n12438), .dout(n12441));
    jdff dff_B_BGfBg8vY1_0(.din(n12441), .dout(n12444));
    jdff dff_B_eT7K70c91_0(.din(n12444), .dout(n12447));
    jdff dff_B_1vmN5luf3_0(.din(n12447), .dout(n12450));
    jdff dff_B_5KAjjyVv9_0(.din(n12450), .dout(n12453));
    jdff dff_B_08wO1yN45_0(.din(n12453), .dout(n12456));
    jdff dff_B_IkqgK7uJ3_0(.din(n12456), .dout(n12459));
    jdff dff_B_Qrk93bQG4_0(.din(n12459), .dout(n12462));
    jdff dff_B_vy2zsUTI4_0(.din(n12462), .dout(n12465));
    jdff dff_B_Iw1JI7LE5_0(.din(n5365), .dout(n12468));
    jdff dff_B_tjMC8laf8_2(.din(G64), .dout(n12471));
    jdff dff_B_R6qd8A5o3_2(.din(G14), .dout(n12474));
    jdff dff_B_UE8GuEbX6_2(.din(n12474), .dout(n12477));
    jdff dff_A_Bw91KRzU6_1(.din(n12482), .dout(n12479));
    jdff dff_A_mFSizQAB5_1(.din(n12485), .dout(n12482));
    jdff dff_A_Tcv2PsEN5_1(.din(n12488), .dout(n12485));
    jdff dff_A_U4ln5SHA2_1(.din(n12491), .dout(n12488));
    jdff dff_A_2Gept2Jo6_1(.din(n12494), .dout(n12491));
    jdff dff_A_KYNLNk6S2_1(.din(n12497), .dout(n12494));
    jdff dff_A_UIvSCv7u3_1(.din(n12500), .dout(n12497));
    jdff dff_A_0f3R6dKC7_1(.din(n12503), .dout(n12500));
    jdff dff_A_rTCv7y8G5_1(.din(n12506), .dout(n12503));
    jdff dff_A_NXzMwWYT0_1(.din(n12509), .dout(n12506));
    jdff dff_A_7Wvx59Ze7_1(.din(n12512), .dout(n12509));
    jdff dff_A_eF1kCpAo5_1(.din(n12515), .dout(n12512));
    jdff dff_A_QMvxRlkL1_1(.din(n12518), .dout(n12515));
    jdff dff_A_WGJbEyxO9_1(.din(n12603), .dout(n12518));
    jdff dff_A_mVjjwKGe3_2(.din(n12524), .dout(n12521));
    jdff dff_A_QV4le3QW2_2(.din(n12527), .dout(n12524));
    jdff dff_A_OpxzFyJB1_2(.din(n12530), .dout(n12527));
    jdff dff_A_77LzJhx87_2(.din(n12533), .dout(n12530));
    jdff dff_A_fTlAtfnV2_2(.din(n12536), .dout(n12533));
    jdff dff_A_XB4NSBmK9_2(.din(n12539), .dout(n12536));
    jdff dff_A_juotzPK26_2(.din(n12542), .dout(n12539));
    jdff dff_A_IZVpXalT3_2(.din(n12545), .dout(n12542));
    jdff dff_A_xS6GkIMI7_2(.din(n12548), .dout(n12545));
    jdff dff_A_Hwmo3KAh3_2(.din(n12603), .dout(n12548));
    jdff dff_A_49N5uduP5_1(.din(n12554), .dout(n12551));
    jdff dff_A_7HfHjDa84_1(.din(n12557), .dout(n12554));
    jdff dff_A_HXCNTPbk8_1(.din(n12560), .dout(n12557));
    jdff dff_A_cQmn4lFP1_1(.din(n12563), .dout(n12560));
    jdff dff_A_pNvcG4Z20_1(.din(n12566), .dout(n12563));
    jdff dff_A_yZz1gfvG6_1(.din(n12569), .dout(n12566));
    jdff dff_A_cv2rVsIN5_1(.din(n12572), .dout(n12569));
    jdff dff_A_4uWKlkDW5_1(.din(n12575), .dout(n12572));
    jdff dff_A_kPq7nZkf0_1(.din(n12578), .dout(n12575));
    jdff dff_A_oo9ebvOe3_1(.din(n12581), .dout(n12578));
    jdff dff_A_kk7zswMP6_1(.din(n12603), .dout(n12581));
    jdff dff_A_ETtXIzyY5_2(.din(n12603), .dout(n12584));
    jdff dff_B_HS0SdTZg8_3(.din(n2356), .dout(n12588));
    jdff dff_B_mhtNTZ0c1_3(.din(n12588), .dout(n12591));
    jdff dff_B_TbCKI1Rc8_3(.din(n12591), .dout(n12594));
    jdff dff_B_E5kYmR2p0_3(.din(n12594), .dout(n12597));
    jdff dff_B_QUibiwm78_3(.din(n12597), .dout(n12600));
    jdff dff_B_YNwcWui00_3(.din(n12600), .dout(n12603));
    jdff dff_A_lQRkkn7L6_1(.din(n12608), .dout(n12605));
    jdff dff_A_A0rPgeOt2_1(.din(n12611), .dout(n12608));
    jdff dff_A_cVR335jI7_1(.din(n12614), .dout(n12611));
    jdff dff_A_ffNL8TsJ5_1(.din(n12617), .dout(n12614));
    jdff dff_A_bxRoYoQg0_1(.din(n12620), .dout(n12617));
    jdff dff_A_A4WVKjca8_1(.din(n12623), .dout(n12620));
    jdff dff_A_8ZmzrnB93_1(.din(n12626), .dout(n12623));
    jdff dff_A_trCIINZ53_1(.din(n12629), .dout(n12626));
    jdff dff_A_RmHbgeXA6_1(.din(n12632), .dout(n12629));
    jdff dff_A_muBslIKH4_1(.din(n12635), .dout(n12632));
    jdff dff_A_DU33Q8n40_1(.din(n12638), .dout(n12635));
    jdff dff_A_kkTUnA3w1_1(.din(n12641), .dout(n12638));
    jdff dff_A_u8b5jmpL2_1(.din(n12644), .dout(n12641));
    jdff dff_A_nLzfCQsM7_1(.din(n12741), .dout(n12644));
    jdff dff_A_VWpPITbl1_2(.din(n12650), .dout(n12647));
    jdff dff_A_VriCAyT59_2(.din(n12653), .dout(n12650));
    jdff dff_A_9veWSEuW6_2(.din(n12656), .dout(n12653));
    jdff dff_A_ESY4zw8P7_2(.din(n12659), .dout(n12656));
    jdff dff_A_WrvQyqRj9_2(.din(n12662), .dout(n12659));
    jdff dff_A_34mx983w1_2(.din(n12665), .dout(n12662));
    jdff dff_A_sj5abWxI0_2(.din(n12668), .dout(n12665));
    jdff dff_A_3ZL6epNk0_2(.din(n12671), .dout(n12668));
    jdff dff_A_ETkTuboE4_2(.din(n12674), .dout(n12671));
    jdff dff_A_8wZX448Z7_2(.din(n12741), .dout(n12674));
    jdff dff_A_xWdDvhNX3_1(.din(n12680), .dout(n12677));
    jdff dff_A_sgeRwZNV6_1(.din(n12683), .dout(n12680));
    jdff dff_A_yd8p5ipB7_1(.din(n12686), .dout(n12683));
    jdff dff_A_TXkCGyfc9_1(.din(n12689), .dout(n12686));
    jdff dff_A_fbiWGzUq3_1(.din(n12692), .dout(n12689));
    jdff dff_A_1ysmOmuF8_1(.din(n12695), .dout(n12692));
    jdff dff_A_MNw5UL0q4_1(.din(n12698), .dout(n12695));
    jdff dff_A_XN9drVBE1_1(.din(n12701), .dout(n12698));
    jdff dff_A_FOjqyKUo7_1(.din(n12704), .dout(n12701));
    jdff dff_A_2QcyE6Bd0_1(.din(n12707), .dout(n12704));
    jdff dff_A_Yw8dhu3K1_1(.din(n12741), .dout(n12707));
    jdff dff_A_MPqETHIJ7_2(.din(n12713), .dout(n12710));
    jdff dff_A_MgUL0Bl02_2(.din(n12716), .dout(n12713));
    jdff dff_A_2s3zZm4n4_2(.din(n12719), .dout(n12716));
    jdff dff_A_1eiEKxGE0_2(.din(n12741), .dout(n12719));
    jdff dff_B_d13xtpX31_3(.din(n2345), .dout(n12723));
    jdff dff_B_46qk7RXw5_3(.din(n12723), .dout(n12726));
    jdff dff_B_wGWUR7wr4_3(.din(n12726), .dout(n12729));
    jdff dff_B_bByIaimR9_3(.din(n12729), .dout(n12732));
    jdff dff_B_7dhOLKPu5_3(.din(n12732), .dout(n12735));
    jdff dff_B_rXjKCc991_3(.din(n12735), .dout(n12738));
    jdff dff_B_ybEFOdHf6_3(.din(n12738), .dout(n12741));
    jdff dff_A_4CRskux41_1(.din(G4090), .dout(n12743));
    jdff dff_A_SGVINllK6_2(.din(G4089), .dout(n12746));
    jdff dff_B_WDSJg6To0_1(.din(n5387), .dout(n12750));
    jdff dff_B_W0VuoQNR9_0(.din(n5425), .dout(n12753));
    jdff dff_B_SJ2s7CJX8_0(.din(n12753), .dout(n12756));
    jdff dff_B_H8iMtuMh1_0(.din(n12756), .dout(n12759));
    jdff dff_B_0PYhF4O05_0(.din(n12759), .dout(n12762));
    jdff dff_B_iEFiicFC9_0(.din(n12762), .dout(n12765));
    jdff dff_B_0qwySIf04_0(.din(n12765), .dout(n12768));
    jdff dff_B_nODTLu8j8_0(.din(n12768), .dout(n12771));
    jdff dff_B_hwZ2QBFM2_0(.din(n12771), .dout(n12774));
    jdff dff_B_cq9WxawO3_0(.din(n12774), .dout(n12777));
    jdff dff_B_guJLuw7V8_0(.din(n12777), .dout(n12780));
    jdff dff_B_ap0gar116_0(.din(n12780), .dout(n12783));
    jdff dff_B_ze3dQJQJ8_0(.din(n12783), .dout(n12786));
    jdff dff_B_N72LmPrQ6_0(.din(n12786), .dout(n12789));
    jdff dff_B_MivFnubg2_0(.din(n12789), .dout(n12792));
    jdff dff_B_eEimXZ8n5_0(.din(n12792), .dout(n12795));
    jdff dff_B_8hT4PvgW8_0(.din(n12795), .dout(n12798));
    jdff dff_B_vLSC3Jhc8_0(.din(n12798), .dout(n12801));
    jdff dff_B_0HFVwDKA1_0(.din(n12801), .dout(n12804));
    jdff dff_B_fNWvu0Ba5_1(.din(n5411), .dout(n12807));
    jdff dff_B_Y8Kz8GFj8_1(.din(n5390), .dout(n12810));
    jdff dff_B_SycmWz7h0_1(.din(n12810), .dout(n12813));
    jdff dff_B_77Z1O1pc6_1(.din(n12813), .dout(n12816));
    jdff dff_B_SLkzalUW6_1(.din(n12816), .dout(n12819));
    jdff dff_B_WmxQRnwC7_1(.din(n12819), .dout(n12822));
    jdff dff_B_Mq51PVmM5_1(.din(n12822), .dout(n12825));
    jdff dff_B_SHf0hWt57_1(.din(n12825), .dout(n12828));
    jdff dff_B_4eLVmgno8_1(.din(n12828), .dout(n12831));
    jdff dff_B_ZJJK44hD6_1(.din(n12831), .dout(n12834));
    jdff dff_B_OZcxFgxD3_1(.din(n12834), .dout(n12837));
    jdff dff_B_S8tdATFH8_1(.din(n12837), .dout(n12840));
    jdff dff_B_RE3od9HI0_1(.din(n12840), .dout(n12843));
    jdff dff_B_ipm9Ljwo2_1(.din(n12843), .dout(n12846));
    jdff dff_B_pq6E21WS5_1(.din(n12846), .dout(n12849));
    jdff dff_B_SZKGjNZO4_1(.din(n12849), .dout(n12852));
    jdff dff_B_f9O6MNGd0_1(.din(n12852), .dout(n12855));
    jdff dff_B_Y58RtSJ29_1(.din(n12855), .dout(n12858));
    jdff dff_B_wotfyTJE5_1(.din(n12858), .dout(n12861));
    jdff dff_B_lU0gpBps2_1(.din(n12861), .dout(n12864));
    jdff dff_A_iHELKUG08_0(.din(n12869), .dout(n12866));
    jdff dff_A_JLMDq7te7_0(.din(n12872), .dout(n12869));
    jdff dff_A_XlXlueqR2_0(.din(n12875), .dout(n12872));
    jdff dff_A_C65bxzey1_0(.din(n12878), .dout(n12875));
    jdff dff_A_jwdxQDeC6_0(.din(n12881), .dout(n12878));
    jdff dff_A_RS3E63ZZ8_0(.din(n2900), .dout(n12881));
    jdff dff_A_zaEMJS5y1_2(.din(n12887), .dout(n12884));
    jdff dff_A_f1Ac9L4z1_2(.din(n12890), .dout(n12887));
    jdff dff_A_4Q7Rqo8r2_2(.din(n12893), .dout(n12890));
    jdff dff_A_5S8BuSF53_2(.din(n12896), .dout(n12893));
    jdff dff_A_n2SQzVNL3_2(.din(n12899), .dout(n12896));
    jdff dff_A_KeYBZipT4_2(.din(n12902), .dout(n12899));
    jdff dff_A_RMdziKXA7_2(.din(n12905), .dout(n12902));
    jdff dff_A_xs8At4Ad5_2(.din(n12908), .dout(n12905));
    jdff dff_A_ssuHvV1x9_2(.din(n12911), .dout(n12908));
    jdff dff_A_YEuyJf9P2_2(.din(n12914), .dout(n12911));
    jdff dff_A_eZyDpLQi3_2(.din(n12917), .dout(n12914));
    jdff dff_A_3d2wZlUO0_2(.din(n12920), .dout(n12917));
    jdff dff_A_XBNuIOju5_2(.din(n12923), .dout(n12920));
    jdff dff_A_wXEszY9E9_2(.din(n12926), .dout(n12923));
    jdff dff_A_Y4SC1a0I0_2(.din(n12929), .dout(n12926));
    jdff dff_A_QLIc4odz2_2(.din(n12932), .dout(n12929));
    jdff dff_A_IkYQX1ya8_2(.din(n12935), .dout(n12932));
    jdff dff_A_WcX8CP5O4_2(.din(n2900), .dout(n12935));
    jdff dff_A_eXFg4IlW1_1(.din(n12941), .dout(n12938));
    jdff dff_A_ScsDh4u38_1(.din(n12944), .dout(n12941));
    jdff dff_A_xhc8N4CO3_1(.din(n12947), .dout(n12944));
    jdff dff_A_V8lgoi8O3_1(.din(n12950), .dout(n12947));
    jdff dff_A_rqzMa1as8_1(.din(n12953), .dout(n12950));
    jdff dff_A_vKmt0qfj2_1(.din(n12956), .dout(n12953));
    jdff dff_A_SBDi12mP8_1(.din(n12959), .dout(n12956));
    jdff dff_A_0n4bZYXa1_1(.din(n12962), .dout(n12959));
    jdff dff_A_wQW1a9xD2_1(.din(n12965), .dout(n12962));
    jdff dff_A_gu81xreD1_1(.din(n12968), .dout(n12965));
    jdff dff_A_OxxtIKWa9_1(.din(n12971), .dout(n12968));
    jdff dff_A_3Vgv66q52_1(.din(n12974), .dout(n12971));
    jdff dff_A_qB07bLz41_1(.din(n12977), .dout(n12974));
    jdff dff_A_JNnxzt9i4_1(.din(n12980), .dout(n12977));
    jdff dff_A_SnYGJwgI1_1(.din(n12983), .dout(n12980));
    jdff dff_A_q74Muz0Z9_1(.din(n2900), .dout(n12983));
    jdff dff_A_FmQcAuyX1_2(.din(n12989), .dout(n12986));
    jdff dff_A_bVDZBFzy6_2(.din(n12992), .dout(n12989));
    jdff dff_A_BJg2IT4b6_2(.din(n12995), .dout(n12992));
    jdff dff_A_PMsPWmz07_2(.din(n12998), .dout(n12995));
    jdff dff_A_JVDka3Zi9_2(.din(n13001), .dout(n12998));
    jdff dff_A_pmBhRDCS4_2(.din(n13004), .dout(n13001));
    jdff dff_A_srwLQ5c40_2(.din(n2900), .dout(n13004));
    jdff dff_B_ADl4x1I67_1(.din(n5383), .dout(n13008));
    jdff dff_B_YIkN63ix3_1(.din(n13008), .dout(n13011));
    jdff dff_B_02i94erj1_1(.din(n13011), .dout(n13014));
    jdff dff_B_1RqGvp9P5_1(.din(n13014), .dout(n13017));
    jdff dff_B_0ZkJsJOg0_1(.din(n13017), .dout(n13020));
    jdff dff_B_xbZwIeDv3_1(.din(n13020), .dout(n13023));
    jdff dff_B_CCf1sQqX0_1(.din(n13023), .dout(n13026));
    jdff dff_B_7i3JhJil5_1(.din(n13026), .dout(n13029));
    jdff dff_B_WdTnOeSQ7_1(.din(n13029), .dout(n13032));
    jdff dff_B_ZILFCqnK7_1(.din(n13032), .dout(n13035));
    jdff dff_B_s0jOnRZr4_1(.din(n13035), .dout(n13038));
    jdff dff_B_T0AZJEkz9_1(.din(n13038), .dout(n13041));
    jdff dff_B_H9PfolCh3_1(.din(n13041), .dout(n13044));
    jdff dff_B_IFzlGp5n3_1(.din(n13044), .dout(n13047));
    jdff dff_B_4dMFw2le9_1(.din(n13047), .dout(n13050));
    jdff dff_B_N973HRmS5_1(.din(n13050), .dout(n13053));
    jdff dff_B_gag6sJdH4_1(.din(n13053), .dout(n13056));
    jdff dff_B_ZhBvSANF8_1(.din(n13056), .dout(n13059));
    jdff dff_B_2TT89mhw0_1(.din(n13059), .dout(n13062));
    jdff dff_A_KaS8Gjmp7_0(.din(n13067), .dout(n13064));
    jdff dff_A_YDSjYdWi1_0(.din(n13070), .dout(n13067));
    jdff dff_A_6sNleYyk2_0(.din(n13073), .dout(n13070));
    jdff dff_A_QeuITl8g9_0(.din(n13076), .dout(n13073));
    jdff dff_A_uopNGU9Q9_0(.din(n13079), .dout(n13076));
    jdff dff_A_A64mu9WC9_0(.din(n13082), .dout(n13079));
    jdff dff_A_Nky4KSlY5_0(.din(n2889), .dout(n13082));
    jdff dff_A_YXbuRvEe6_2(.din(n13088), .dout(n13085));
    jdff dff_A_E8b3whZb0_2(.din(n13091), .dout(n13088));
    jdff dff_A_Z6sV74iU8_2(.din(n13094), .dout(n13091));
    jdff dff_A_ygwnds2u5_2(.din(n13097), .dout(n13094));
    jdff dff_A_BkgepQIr4_2(.din(n13100), .dout(n13097));
    jdff dff_A_EDUFbXmI6_2(.din(n13103), .dout(n13100));
    jdff dff_A_Fqya9Ppc7_2(.din(n13106), .dout(n13103));
    jdff dff_A_bvgAqDQA7_2(.din(n13109), .dout(n13106));
    jdff dff_A_yYPMmlIl2_2(.din(n13112), .dout(n13109));
    jdff dff_A_Yp2IxehB0_2(.din(n13115), .dout(n13112));
    jdff dff_A_Gi0yjUwF7_2(.din(n13118), .dout(n13115));
    jdff dff_A_7LVqeWkA3_2(.din(n13121), .dout(n13118));
    jdff dff_A_OsZUJQAV4_2(.din(n13124), .dout(n13121));
    jdff dff_A_Vf9Gdczv3_2(.din(n13127), .dout(n13124));
    jdff dff_A_LHry1Kob6_2(.din(n13130), .dout(n13127));
    jdff dff_A_yj4xZaDO9_2(.din(n13133), .dout(n13130));
    jdff dff_A_qDdl9PUa3_2(.din(n13136), .dout(n13133));
    jdff dff_A_Gx3srTJB5_2(.din(n13139), .dout(n13136));
    jdff dff_A_9vZJQ24L1_2(.din(n2889), .dout(n13139));
    jdff dff_A_SzmOzkWV1_1(.din(n13145), .dout(n13142));
    jdff dff_A_EawolTbo1_1(.din(n13148), .dout(n13145));
    jdff dff_A_c5kw5qj53_1(.din(n13151), .dout(n13148));
    jdff dff_A_CySUXMTS8_1(.din(n13154), .dout(n13151));
    jdff dff_A_0FhMjHqI6_1(.din(n13157), .dout(n13154));
    jdff dff_A_VUbQvf5T2_1(.din(n13160), .dout(n13157));
    jdff dff_A_KRZJpQur7_1(.din(n13163), .dout(n13160));
    jdff dff_A_VewggG2H4_1(.din(n13166), .dout(n13163));
    jdff dff_A_6QfcUjhk5_1(.din(n13169), .dout(n13166));
    jdff dff_A_qno6efzJ4_1(.din(n13172), .dout(n13169));
    jdff dff_A_foLlheHq1_1(.din(n13175), .dout(n13172));
    jdff dff_A_QOzIT3WG2_1(.din(n13178), .dout(n13175));
    jdff dff_A_DSCTJOUl1_1(.din(n13181), .dout(n13178));
    jdff dff_A_uKVMB4oG5_1(.din(n13184), .dout(n13181));
    jdff dff_A_4G2HRrGl2_1(.din(n13187), .dout(n13184));
    jdff dff_A_EoNtu0H00_1(.din(n13190), .dout(n13187));
    jdff dff_A_RFQeJ0rj8_1(.din(n2889), .dout(n13190));
    jdff dff_A_MN9hvVqO9_2(.din(n13196), .dout(n13193));
    jdff dff_A_zY7AvL4P7_2(.din(n13199), .dout(n13196));
    jdff dff_A_5tARJulS1_2(.din(n13202), .dout(n13199));
    jdff dff_A_iqPyKJ4v2_2(.din(n13205), .dout(n13202));
    jdff dff_A_HPm1gUJ59_2(.din(n13208), .dout(n13205));
    jdff dff_A_DF7xBQUR0_2(.din(n13211), .dout(n13208));
    jdff dff_A_KtPzDrIM2_2(.din(n13214), .dout(n13211));
    jdff dff_A_dwSHW1VY7_2(.din(n13217), .dout(n13214));
    jdff dff_A_TZqrMTYV7_2(.din(n13220), .dout(n13217));
    jdff dff_A_nShUj1GO1_2(.din(n13223), .dout(n13220));
    jdff dff_A_XlHVV9RA6_2(.din(n2889), .dout(n13223));
    jdff dff_A_kWN7fJzX1_1(.din(G1690), .dout(n13226));
    jdff dff_A_shACUS9a7_2(.din(G1689), .dout(n13229));
    jdff dff_B_kO1xlF5h5_1(.din(n5444), .dout(n13233));
    jdff dff_B_LfIV5xTx3_0(.din(n5469), .dout(n13236));
    jdff dff_B_UiMih9lw6_0(.din(n13236), .dout(n13239));
    jdff dff_B_bmXPNjKx8_0(.din(n13239), .dout(n13242));
    jdff dff_B_0XCAjgoC6_0(.din(n13242), .dout(n13245));
    jdff dff_B_7mLXmI0j0_0(.din(n13245), .dout(n13248));
    jdff dff_B_zibivfLm9_0(.din(n13248), .dout(n13251));
    jdff dff_B_rDNdzLCw9_0(.din(n13251), .dout(n13254));
    jdff dff_B_aCpFc6yW1_0(.din(n13254), .dout(n13257));
    jdff dff_B_xG6T76pF6_0(.din(n13257), .dout(n13260));
    jdff dff_B_6ARhtCrO9_0(.din(n13260), .dout(n13263));
    jdff dff_B_nLYEia8J2_0(.din(n13263), .dout(n13266));
    jdff dff_B_sMYYjckc0_0(.din(n13266), .dout(n13269));
    jdff dff_B_lpK4u32E2_0(.din(n13269), .dout(n13272));
    jdff dff_B_Q6TBJCfg7_0(.din(n13272), .dout(n13275));
    jdff dff_B_DenSSNA57_0(.din(n13275), .dout(n13278));
    jdff dff_B_i1VLYggP1_0(.din(n13278), .dout(n13281));
    jdff dff_B_7zETgrhx6_0(.din(n13281), .dout(n13284));
    jdff dff_B_sUjayH6W6_0(.din(n13284), .dout(n13287));
    jdff dff_B_pjxcf6tk2_1(.din(n5458), .dout(n13290));
    jdff dff_B_fnBqcRVL1_2(.din(n5414), .dout(n13293));
    jdff dff_B_9ka1Ae2n2_2(.din(n13293), .dout(n13296));
    jdff dff_B_uXGqDPoi2_2(.din(n5404), .dout(n13299));
    jdff dff_B_5nRWFFqr8_1(.din(n5447), .dout(n13302));
    jdff dff_B_BSIomkER9_1(.din(n13302), .dout(n13305));
    jdff dff_B_mRgcY9Nb7_1(.din(n13305), .dout(n13308));
    jdff dff_B_nCoNP1I53_1(.din(n13308), .dout(n13311));
    jdff dff_B_jSEeUeMY0_1(.din(n13311), .dout(n13314));
    jdff dff_B_DNB5IOhH3_1(.din(n13314), .dout(n13317));
    jdff dff_B_jcYqNVaM4_1(.din(n13317), .dout(n13320));
    jdff dff_B_bsWaEmUV7_1(.din(n13320), .dout(n13323));
    jdff dff_B_nvfFrwUp2_1(.din(n13323), .dout(n13326));
    jdff dff_B_oQwCSowM1_1(.din(n13326), .dout(n13329));
    jdff dff_B_H4yjJnyj3_1(.din(n13329), .dout(n13332));
    jdff dff_B_q7zrlhNy5_1(.din(n13332), .dout(n13335));
    jdff dff_B_IYsRfYYL9_1(.din(n13335), .dout(n13338));
    jdff dff_B_GTWJnPbN0_1(.din(n13338), .dout(n13341));
    jdff dff_B_3YKgXkRR4_1(.din(n13341), .dout(n13344));
    jdff dff_B_whtlgsNr0_1(.din(n13344), .dout(n13347));
    jdff dff_B_iOwKKTv57_1(.din(n13347), .dout(n13350));
    jdff dff_B_Gt6abUR49_1(.din(n13350), .dout(n13353));
    jdff dff_B_QQQYwGwz9_1(.din(n13353), .dout(n13356));
    jdff dff_B_nSyVskDI9_0(.din(n5393), .dout(n13359));
    jdff dff_B_8wF03YzM8_0(.din(n13359), .dout(n13362));
    jdff dff_B_aPuqufsa5_0(.din(n13362), .dout(n13365));
    jdff dff_B_8VUeNZon6_0(.din(n13365), .dout(n13368));
    jdff dff_B_yHoVVJiQ8_0(.din(n13368), .dout(n13371));
    jdff dff_B_WfVGL2fU4_0(.din(n13371), .dout(n13374));
    jdff dff_B_GY4ZbLlM0_0(.din(n13374), .dout(n13377));
    jdff dff_B_ITN3cMfV3_0(.din(n13377), .dout(n13380));
    jdff dff_B_HrHYRHr98_0(.din(n13380), .dout(n13383));
    jdff dff_B_cBe28yCV4_0(.din(n13383), .dout(n13386));
    jdff dff_B_XUgYyT8M9_0(.din(n13386), .dout(n13389));
    jdff dff_B_R9gTmzsv8_0(.din(n13389), .dout(n13392));
    jdff dff_B_AWCXUrGL8_0(.din(n13392), .dout(n13395));
    jdff dff_B_zvaA5D1N9_0(.din(n13395), .dout(n13398));
    jdff dff_B_g8Zkx60P2_0(.din(n13398), .dout(n13401));
    jdff dff_B_5MZ4CJjg4_0(.din(n13401), .dout(n13404));
    jdff dff_B_6rYAchRu8_0(.din(n13404), .dout(n13407));
    jdff dff_B_U9I6NSKP4_0(.din(n13407), .dout(n13410));
    jdff dff_B_VkqJ4JdF2_0(.din(n13410), .dout(n13413));
    jdff dff_A_2qNBQAAz1_1(.din(n13418), .dout(n13415));
    jdff dff_A_KXq6F43g4_1(.din(n13421), .dout(n13418));
    jdff dff_A_M7eigc2J0_1(.din(n13424), .dout(n13421));
    jdff dff_A_mE0bREcL4_1(.din(n13427), .dout(n13424));
    jdff dff_A_e3XV9LNK4_1(.din(n13430), .dout(n13427));
    jdff dff_A_vxnwc74m0_1(.din(n13433), .dout(n13430));
    jdff dff_A_WlQMOzsc4_1(.din(n13436), .dout(n13433));
    jdff dff_A_q6RkgbSP8_1(.din(n13439), .dout(n13436));
    jdff dff_A_XhfRU2u52_1(.din(n13442), .dout(n13439));
    jdff dff_A_0V4Iu1L22_1(.din(n13445), .dout(n13442));
    jdff dff_A_Y90mAvUv5_1(.din(n13448), .dout(n13445));
    jdff dff_A_1iWUyKb64_1(.din(n13451), .dout(n13448));
    jdff dff_A_stdcJoPf5_1(.din(n13454), .dout(n13451));
    jdff dff_A_4erDwzrp7_1(.din(n13457), .dout(n13454));
    jdff dff_A_H93Uu6Zn8_1(.din(n13460), .dout(n13457));
    jdff dff_A_pR8iYj328_1(.din(n13463), .dout(n13460));
    jdff dff_A_EAQwzC245_1(.din(n13466), .dout(n13463));
    jdff dff_A_cKvkMZMF8_1(.din(n13469), .dout(n13466));
    jdff dff_A_a0wee1C72_1(.din(n13472), .dout(n13469));
    jdff dff_A_lOfGrWq38_1(.din(n5321), .dout(n13472));
    jdff dff_B_EiferPjr7_1(.din(n4475), .dout(n13476));
    jdff dff_B_LEYSzV9g6_1(.din(n13476), .dout(n13479));
    jdff dff_B_WDjFJlta3_1(.din(n13479), .dout(n13482));
    jdff dff_B_A5UV8FbO1_1(.din(n13482), .dout(n13485));
    jdff dff_B_vPNP0QHB0_1(.din(n13485), .dout(n13488));
    jdff dff_B_srRKSC302_1(.din(n13488), .dout(n13491));
    jdff dff_A_uP4cssC57_1(.din(n4684), .dout(n13493));
    jdff dff_B_zLvkXYvw7_1(.din(n4550), .dout(n13497));
    jdff dff_B_Ctzvl1pv9_1(.din(n13497), .dout(n13500));
    jdff dff_B_ccoYs86D7_1(.din(n13500), .dout(n13503));
    jdff dff_B_fAtLgESn2_1(.din(n13503), .dout(n13506));
    jdff dff_B_h2h6XhD24_1(.din(n13506), .dout(n13509));
    jdff dff_B_78h5uKli9_1(.din(n13509), .dout(n13512));
    jdff dff_B_y4lPWIZM9_1(.din(n13512), .dout(n13515));
    jdff dff_B_Ycw62p2G9_1(.din(n13515), .dout(n13518));
    jdff dff_B_OKGcimLH4_1(.din(n13518), .dout(n13521));
    jdff dff_B_T5OrYCv76_1(.din(n13521), .dout(n13524));
    jdff dff_B_B8p0AihC4_0(.din(n4668), .dout(n13527));
    jdff dff_B_rYpnkdck4_0(.din(n4656), .dout(n13530));
    jdff dff_A_DAnZjvDa5_1(.din(n13535), .dout(n13532));
    jdff dff_A_RU3PesLf9_1(.din(n13538), .dout(n13535));
    jdff dff_A_i4tnNOao0_1(.din(n4649), .dout(n13538));
    jdff dff_B_JlEetKWX5_0(.din(n4645), .dout(n13542));
    jdff dff_B_93VvCCoL9_1(.din(n4607), .dout(n13545));
    jdff dff_B_fBAZfIPF1_1(.din(n4610), .dout(n13548));
    jdff dff_B_CmMYRjGy6_1(.din(n13548), .dout(n13551));
    jdff dff_B_k8wkP7V45_1(.din(n13551), .dout(n13554));
    jdff dff_B_l5805JJW3_1(.din(n13554), .dout(n13557));
    jdff dff_B_qtoGbi9Q3_1(.din(n13557), .dout(n13560));
    jdff dff_B_DvW9Xmlr0_1(.din(n13560), .dout(n13563));
    jdff dff_B_mn2IDOe53_1(.din(n13563), .dout(n13566));
    jdff dff_B_ImFpiWwF0_1(.din(n13566), .dout(n13569));
    jdff dff_B_6ADLqYUy0_1(.din(n13569), .dout(n13572));
    jdff dff_B_8lN77ZZV8_1(.din(n13572), .dout(n13575));
    jdff dff_B_E8bw2Xc02_1(.din(n13575), .dout(n13578));
    jdff dff_B_5hVWzVVv8_1(.din(n4557), .dout(n13581));
    jdff dff_B_xPpdEmg91_1(.din(n13581), .dout(n13584));
    jdff dff_B_hahaZNaU7_1(.din(n13584), .dout(n13587));
    jdff dff_B_m1reyT1g6_1(.din(n13587), .dout(n13590));
    jdff dff_B_DZsrSaJC9_1(.din(n4591), .dout(n13593));
    jdff dff_B_5XddWEBp3_0(.din(n4587), .dout(n13596));
    jdff dff_A_HcOHyT6M2_0(.din(n13601), .dout(n13598));
    jdff dff_A_X51ckPEc8_0(.din(n13604), .dout(n13601));
    jdff dff_A_dwyuefgZ4_0(.din(n4584), .dout(n13604));
    jdff dff_B_41D4gjXK6_1(.din(n4560), .dout(n13608));
    jdff dff_A_q39Y62Qo9_1(.din(n2303), .dout(n13610));
    jdff dff_A_7U8dAIfM4_0(.din(n13616), .dout(n13613));
    jdff dff_A_Dj08AoB85_0(.din(n13619), .dout(n13616));
    jdff dff_A_3BqQ1vZL7_0(.din(n13622), .dout(n13619));
    jdff dff_A_GRkkIbkc5_0(.din(n13625), .dout(n13622));
    jdff dff_A_yFlhvwaL7_0(.din(n1481), .dout(n13625));
    jdff dff_A_vMZcvEne7_2(.din(n13631), .dout(n13628));
    jdff dff_A_v8ccX43L2_2(.din(n13634), .dout(n13631));
    jdff dff_A_6R0eBoST5_2(.din(n13637), .dout(n13634));
    jdff dff_A_43kEHPEg7_2(.din(n13640), .dout(n13637));
    jdff dff_A_7VdfCcrB8_2(.din(n13643), .dout(n13640));
    jdff dff_A_SfMgCxe87_2(.din(n1481), .dout(n13643));
    jdff dff_A_J6xtzue03_1(.din(n13649), .dout(n13646));
    jdff dff_A_exhrGTRb2_1(.din(n13652), .dout(n13649));
    jdff dff_A_U8cEK5rx7_1(.din(n13655), .dout(n13652));
    jdff dff_A_bsDESXrn1_1(.din(n13658), .dout(n13655));
    jdff dff_A_Llzfcz2D6_1(.din(n13661), .dout(n13658));
    jdff dff_A_9p8FwHgm0_1(.din(n2299), .dout(n13661));
    jdff dff_A_oFlFmqrn6_2(.din(n13667), .dout(n13664));
    jdff dff_A_VZ74eUt02_2(.din(n2299), .dout(n13667));
    jdff dff_B_3haLFshg7_2(.din(n2143), .dout(n13671));
    jdff dff_B_YNCr1ghA7_2(.din(n13671), .dout(n13674));
    jdff dff_B_H8r2rb7a7_2(.din(n13674), .dout(n13677));
    jdff dff_B_qSk3uBpR2_2(.din(n13677), .dout(n13680));
    jdff dff_B_kx3bsKHd9_2(.din(n13680), .dout(n13683));
    jdff dff_B_5c34sflw2_2(.din(n13683), .dout(n13686));
    jdff dff_B_YU7MduXM0_2(.din(n13686), .dout(n13689));
    jdff dff_B_PlWYkjCq5_2(.din(n13689), .dout(n13692));
    jdff dff_B_G0r8g5BP1_2(.din(n13692), .dout(n13695));
    jdff dff_A_p02ZZeyY1_1(.din(n13700), .dout(n13697));
    jdff dff_A_PiutBOKW9_1(.din(n13703), .dout(n13700));
    jdff dff_A_fo7ty2Ig3_1(.din(n13706), .dout(n13703));
    jdff dff_A_vi7fcVaA1_1(.din(n13709), .dout(n13706));
    jdff dff_A_qyJST7g97_1(.din(n13712), .dout(n13709));
    jdff dff_A_T9XOHi6A6_1(.din(n13715), .dout(n13712));
    jdff dff_A_FmJG8Dnv8_1(.din(n13718), .dout(n13715));
    jdff dff_A_19NKEVfM8_1(.din(n13721), .dout(n13718));
    jdff dff_A_zsOTnmHl7_1(.din(n13724), .dout(n13721));
    jdff dff_A_8mvt0AeL9_1(.din(n13727), .dout(n13724));
    jdff dff_A_ZHVBNmEb4_1(.din(n13730), .dout(n13727));
    jdff dff_A_oxz4LApm0_1(.din(n2113), .dout(n13730));
    jdff dff_A_2vLDGwbn1_1(.din(n13736), .dout(n13733));
    jdff dff_A_YybsqF5R9_1(.din(n1567), .dout(n13736));
    jdff dff_A_lDwR0oxZ1_2(.din(n1567), .dout(n13739));
    jdff dff_A_83I4TDbd0_0(.din(n13745), .dout(n13742));
    jdff dff_A_VhoHiYwh2_0(.din(n13748), .dout(n13745));
    jdff dff_A_XEg2A39h3_0(.din(n13751), .dout(n13748));
    jdff dff_A_1MjHR3At8_0(.din(n13754), .dout(n13751));
    jdff dff_A_FKyPYXmF7_0(.din(n13757), .dout(n13754));
    jdff dff_A_CRdPderv7_0(.din(n13760), .dout(n13757));
    jdff dff_A_nQxZ6Apw4_0(.din(n13763), .dout(n13760));
    jdff dff_A_bInQ2ewd0_0(.din(n13766), .dout(n13763));
    jdff dff_A_8aOzhEPB5_0(.din(n13769), .dout(n13766));
    jdff dff_A_9i10deTR1_0(.din(n13772), .dout(n13769));
    jdff dff_A_yQLIJlPF6_0(.din(n4547), .dout(n13772));
    jdff dff_A_07bBmpDT9_0(.din(n4540), .dout(n13775));
    jdff dff_B_jKVjrq5X9_1(.din(n4525), .dout(n13779));
    jdff dff_B_fhLSiVLT7_0(.din(n4532), .dout(n13782));
    jdff dff_B_E6HVoo1T4_0(.din(n13782), .dout(n13785));
    jdff dff_B_TQRLK7av2_0(.din(n13785), .dout(n13788));
    jdff dff_B_0jfqp2Sr6_0(.din(n13788), .dout(n13791));
    jdff dff_A_A7pyJF0q2_1(.din(n13796), .dout(n13793));
    jdff dff_A_GIQAnLri7_1(.din(n13799), .dout(n13796));
    jdff dff_A_c2uT18W97_1(.din(n13802), .dout(n13799));
    jdff dff_A_h1JDWaJA3_1(.din(n13805), .dout(n13802));
    jdff dff_A_qkS26nqD6_1(.din(n13821), .dout(n13805));
    jdff dff_B_M8L1t6OB9_2(.din(n2823), .dout(n13809));
    jdff dff_B_sCZfvn0t7_2(.din(n13809), .dout(n13812));
    jdff dff_B_Ki3Mc9955_2(.din(n13812), .dout(n13815));
    jdff dff_B_p2gEwM9Z5_2(.din(n13815), .dout(n13818));
    jdff dff_B_qYv6NP3V6_2(.din(n13818), .dout(n13821));
    jdff dff_B_246mbD024_0(.din(n4521), .dout(n13824));
    jdff dff_B_IKKyRrnr9_0(.din(n13824), .dout(n13827));
    jdff dff_B_S1s3UIPE3_1(.din(n4509), .dout(n13830));
    jdff dff_B_dh32HErn3_1(.din(n13830), .dout(n13833));
    jdff dff_B_Q5aEoJqx2_1(.din(n13833), .dout(n13836));
    jdff dff_A_qLi9mKAP9_1(.din(n13841), .dout(n13838));
    jdff dff_A_i29xRiPG6_1(.din(n13844), .dout(n13841));
    jdff dff_A_MmFNpZCS8_1(.din(n13869), .dout(n13844));
    jdff dff_A_HmG6Z6ho0_2(.din(n13850), .dout(n13847));
    jdff dff_A_2gdmoAsn9_2(.din(n13853), .dout(n13850));
    jdff dff_A_6tH0pIWo0_2(.din(n13856), .dout(n13853));
    jdff dff_A_RMtnfA0Q2_2(.din(n13859), .dout(n13856));
    jdff dff_A_Cx4XFVwu0_2(.din(n13862), .dout(n13859));
    jdff dff_A_ppNgcQAy5_2(.din(n13865), .dout(n13862));
    jdff dff_A_uonOlQ6T0_2(.din(n13869), .dout(n13865));
    jdff dff_B_5M9btRQs8_3(.din(n1625), .dout(n13869));
    jdff dff_A_l8vT5vQK1_0(.din(n13874), .dout(n13871));
    jdff dff_A_VNLyh4yD4_0(.din(n13877), .dout(n13874));
    jdff dff_A_t9r41Nco3_0(.din(n13880), .dout(n13877));
    jdff dff_A_vw1ZzAog0_0(.din(n13883), .dout(n13880));
    jdff dff_A_kLsYy4kh4_0(.din(n13886), .dout(n13883));
    jdff dff_A_rhwnmWmK9_0(.din(n13889), .dout(n13886));
    jdff dff_A_ohl3pi0p0_0(.din(n13892), .dout(n13889));
    jdff dff_A_nXyAlhw77_0(.din(n13895), .dout(n13892));
    jdff dff_A_KnkyxPvf7_0(.din(n1621), .dout(n13895));
    jdff dff_B_1KEajjX92_1(.din(n4487), .dout(n13899));
    jdff dff_A_kUQDiRdJ1_1(.din(n1969), .dout(n13901));
    jdff dff_A_JlBhJpDg0_0(.din(n13907), .dout(n13904));
    jdff dff_A_d4qRLEDP4_0(.din(n13910), .dout(n13907));
    jdff dff_A_a3SyjLHw4_0(.din(n13913), .dout(n13910));
    jdff dff_A_sutFpcGy7_0(.din(n13916), .dout(n13913));
    jdff dff_A_uCbpn1v40_0(.din(n13919), .dout(n13916));
    jdff dff_A_D8G3IhyY8_0(.din(n13922), .dout(n13919));
    jdff dff_A_ye3YonQl8_0(.din(n13925), .dout(n13922));
    jdff dff_A_wNlLgMxG5_0(.din(n13928), .dout(n13925));
    jdff dff_A_yKP8tZG88_0(.din(n1965), .dout(n13928));
    jdff dff_A_OuggQ7wO4_2(.din(n13934), .dout(n13931));
    jdff dff_A_xoIC4ohq8_2(.din(n13937), .dout(n13934));
    jdff dff_A_cPVSayx24_2(.din(n13940), .dout(n13937));
    jdff dff_A_LSHlXkhS6_2(.din(n13943), .dout(n13940));
    jdff dff_A_FIgmJxWn2_2(.din(n1965), .dout(n13943));
    jdff dff_A_MlFFv0D18_2(.din(n1617), .dout(n13946));
    jdff dff_B_5BaMNZE13_0(.din(n1613), .dout(n13950));
    jdff dff_B_d9S4yyXW1_1(.din(G323), .dout(n13953));
    jdff dff_A_Ah5jx5xq6_0(.din(n13958), .dout(n13955));
    jdff dff_A_5FaKLTAu6_0(.din(n13961), .dout(n13958));
    jdff dff_A_hdHaghVi9_0(.din(n13964), .dout(n13961));
    jdff dff_A_7y3fmF6K9_0(.din(n13967), .dout(n13964));
    jdff dff_A_KMCz86P61_0(.din(n13970), .dout(n13967));
    jdff dff_A_ZHwX3Y8X3_0(.din(n13973), .dout(n13970));
    jdff dff_A_T63qrX6K1_0(.din(n13976), .dout(n13973));
    jdff dff_A_EgHcgpFC8_0(.din(n13979), .dout(n13976));
    jdff dff_A_mB80jkcS5_0(.din(n13982), .dout(n13979));
    jdff dff_A_zpxvzAgL6_0(.din(n13985), .dout(n13982));
    jdff dff_A_OwxKxIKB0_0(.din(n1582), .dout(n13985));
    jdff dff_A_RZPL5dbr7_0(.din(n13991), .dout(n13988));
    jdff dff_A_mdWYaNkU6_0(.din(n1605), .dout(n13991));
    jdff dff_B_kjeHPyV10_0(.din(n1597), .dout(n13995));
    jdff dff_B_Ku26dCwl2_1(.din(G315), .dout(n13998));
    jdff dff_A_7qnZTphL5_1(.din(n1582), .dout(n14000));
    jdff dff_A_BkVAH2ZV8_2(.din(n14006), .dout(n14003));
    jdff dff_A_vwcKKIkE5_2(.din(n14009), .dout(n14006));
    jdff dff_A_VRwsdY0y4_2(.din(n14012), .dout(n14009));
    jdff dff_A_A3OPp8uX3_2(.din(n14015), .dout(n14012));
    jdff dff_A_azJ1Cwza1_2(.din(n14018), .dout(n14015));
    jdff dff_A_6qlwNx9c4_2(.din(n14021), .dout(n14018));
    jdff dff_A_BeDjNIWs3_2(.din(n14024), .dout(n14021));
    jdff dff_A_sp6qozvR2_2(.din(n14027), .dout(n14024));
    jdff dff_A_tAJIxZZM3_2(.din(n14030), .dout(n14027));
    jdff dff_A_zHqaBtl11_2(.din(n14033), .dout(n14030));
    jdff dff_A_m2MJmds47_2(.din(n1582), .dout(n14033));
    jdff dff_B_y2tM4x287_1(.din(n1571), .dout(n14037));
    jdff dff_B_9MSpMEdm3_1(.din(G307), .dout(n14040));
    jdff dff_B_l1rPpzD15_0(.din(n4479), .dout(n14043));
    jdff dff_B_QJtKWBiP2_0(.din(n14043), .dout(n14046));
    jdff dff_B_bavSCnqv8_0(.din(n14046), .dout(n14049));
    jdff dff_A_607vqbmS9_0(.din(n14054), .dout(n14051));
    jdff dff_A_0bob9csf8_0(.din(n14057), .dout(n14054));
    jdff dff_A_HIdUAKGh5_0(.din(n1548), .dout(n14057));
    jdff dff_A_nmDxEz0M2_1(.din(n14063), .dout(n14060));
    jdff dff_A_YPqa7FE77_1(.din(n14066), .dout(n14063));
    jdff dff_A_ArazxxYs6_1(.din(n1540), .dout(n14066));
    jdff dff_A_y078HFsd3_1(.din(n1536), .dout(n14069));
    jdff dff_B_VrYukKn71_0(.din(n1532), .dout(n14073));
    jdff dff_A_PGqWpFTY3_0(.din(n1524), .dout(n14075));
    jdff dff_A_ye7KwXvM9_2(.din(n1524), .dout(n14078));
    jdff dff_A_rPjvbile5_0(.din(n1516), .dout(n14081));
    jdff dff_B_rkiHOKfh7_0(.din(n1489), .dout(n14085));
    jdff dff_A_7yrUm62o8_0(.din(n14090), .dout(n14087));
    jdff dff_A_zm4lqhY66_0(.din(n14093), .dout(n14090));
    jdff dff_A_5Xz5M9m92_0(.din(n14096), .dout(n14093));
    jdff dff_A_ekf3WwRm4_0(.din(n14099), .dout(n14096));
    jdff dff_A_pqviEFAC5_0(.din(n14102), .dout(n14099));
    jdff dff_A_rjfCWH7v3_0(.din(n14105), .dout(n14102));
    jdff dff_A_JZRfTq6S6_0(.din(n14108), .dout(n14105));
    jdff dff_A_IBfCtatM8_0(.din(n14111), .dout(n14108));
    jdff dff_A_tO8jjP8l6_0(.din(n14114), .dout(n14111));
    jdff dff_A_5bV9BeUp6_0(.din(n14117), .dout(n14114));
    jdff dff_A_2PvgxPFn8_0(.din(G2174), .dout(n14117));
    jdff dff_A_J7IMqfUf0_2(.din(n14123), .dout(n14120));
    jdff dff_A_eqOLkfew4_2(.din(n14126), .dout(n14123));
    jdff dff_A_bYIpvWPS6_2(.din(n14129), .dout(n14126));
    jdff dff_A_G1x36azM6_2(.din(n14132), .dout(n14129));
    jdff dff_A_CNIbL2NR6_2(.din(n14135), .dout(n14132));
    jdff dff_A_wKjQFHTu1_2(.din(n14138), .dout(n14135));
    jdff dff_A_ESHT4cdV3_2(.din(n14141), .dout(n14138));
    jdff dff_A_yp2Uiusj4_2(.din(G2174), .dout(n14141));
    jdff dff_B_JGqAcsRr8_1(.din(n1857), .dout(n14145));
    jdff dff_B_GHUFqe1f3_1(.din(n14145), .dout(n14148));
    jdff dff_B_fulIQZQl7_1(.din(n14148), .dout(n14151));
    jdff dff_B_9sooi4Uc8_1(.din(n14151), .dout(n14154));
    jdff dff_B_8kjyRUHx5_1(.din(n14154), .dout(n14157));
    jdff dff_B_UwWcPl1b7_1(.din(n14157), .dout(n14160));
    jdff dff_B_SLHDcqRL3_1(.din(n1861), .dout(n14163));
    jdff dff_B_t1eZh6es9_1(.din(n14163), .dout(n14166));
    jdff dff_B_b1MTaIZk2_1(.din(n14166), .dout(n14169));
    jdff dff_B_LeAwGtZq7_1(.din(n14169), .dout(n14172));
    jdff dff_B_boRSAyMn0_1(.din(n14172), .dout(n14175));
    jdff dff_B_WFuUAlZN4_1(.din(n1865), .dout(n14178));
    jdff dff_B_znUCkEJB4_1(.din(n14178), .dout(n14181));
    jdff dff_B_W4dZU0oB8_1(.din(n14181), .dout(n14184));
    jdff dff_B_J8ZZvl7V7_1(.din(n14184), .dout(n14187));
    jdff dff_A_jDdGjmD57_0(.din(n1905), .dout(n14189));
    jdff dff_A_IFsxbyU17_0(.din(n1509), .dout(n14192));
    jdff dff_A_9v7IrxGW5_1(.din(n14198), .dout(n14195));
    jdff dff_A_xwNgPe5F2_1(.din(n14201), .dout(n14198));
    jdff dff_A_QfJbN9cG1_1(.din(n14204), .dout(n14201));
    jdff dff_A_fZ1P4Zf60_1(.din(n14207), .dout(n14204));
    jdff dff_A_c6KmzTiU9_1(.din(n14210), .dout(n14207));
    jdff dff_A_BlrkuVzQ3_1(.din(n1897), .dout(n14210));
    jdff dff_A_JD0BOWzY6_0(.din(G358), .dout(n14213));
    jdff dff_A_tNKKSYbO1_0(.din(n14478), .dout(n14216));
    jdff dff_A_UvZHh7uC5_1(.din(n14478), .dout(n14219));
    jdff dff_A_6QtFNhGn3_1(.din(n14225), .dout(n14222));
    jdff dff_A_bRFzw5NC2_1(.din(n14228), .dout(n14225));
    jdff dff_A_HKufdfLD0_1(.din(n1881), .dout(n14228));
    jdff dff_A_tGhsZud05_2(.din(n14234), .dout(n14231));
    jdff dff_A_CKr4KLtG9_2(.din(n1881), .dout(n14234));
    jdff dff_A_IcUKXp9b7_0(.din(G348), .dout(n14237));
    jdff dff_A_IDL7tBGd6_0(.din(G332), .dout(n14240));
    jdff dff_A_n0fgwF552_0(.din(n14645), .dout(n14243));
    jdff dff_A_S9nwTBvd1_1(.din(n14645), .dout(n14246));
    jdff dff_A_289YKKsd7_0(.din(G332), .dout(n14249));
    jdff dff_A_5nV0ELg97_2(.din(G332), .dout(n14252));
    jdff dff_A_gHKJPNrq2_0(.din(n702), .dout(n14255));
    jdff dff_A_tX71DhYN1_0(.din(n14261), .dout(n14258));
    jdff dff_A_vjaJejNG5_0(.din(n14264), .dout(n14261));
    jdff dff_A_JWom5X3a3_0(.din(n14267), .dout(n14264));
    jdff dff_A_2HCW811z8_1(.din(n14270), .dout(n14267));
    jdff dff_A_MGTmNajW1_1(.din(n1481), .dout(n14270));
    jdff dff_A_O8HdHmMk5_2(.din(n14276), .dout(n14273));
    jdff dff_A_e2wFTsdm5_2(.din(n14279), .dout(n14276));
    jdff dff_A_sDamZIWu9_2(.din(n14282), .dout(n14279));
    jdff dff_A_HBGiEuX35_2(.din(n1481), .dout(n14282));
    jdff dff_B_rYGqbmNG0_1(.din(n1466), .dout(n14286));
    jdff dff_A_LT5SgMpK3_0(.din(G332), .dout(n14288));
    jdff dff_A_TWNRPvyV2_2(.din(G332), .dout(n14291));
    jdff dff_A_7Eb9Jmja7_1(.din(G331), .dout(n14294));
    jdff dff_A_dWzcPerA0_0(.din(n14300), .dout(n14297));
    jdff dff_A_CaI8okV65_0(.din(n14303), .dout(n14300));
    jdff dff_A_3PmkaxBr7_0(.din(n14306), .dout(n14303));
    jdff dff_A_Sg7RcbN19_0(.din(n14309), .dout(n14306));
    jdff dff_A_rjwvY9S35_0(.din(n14312), .dout(n14309));
    jdff dff_A_ydPM95mj5_0(.din(n14315), .dout(n14312));
    jdff dff_A_2zAA9Umb0_0(.din(n4472), .dout(n14315));
    jdff dff_B_SQxsLgcW7_1(.din(n4464), .dout(n14319));
    jdff dff_B_fwDQ9fKU8_1(.din(n14319), .dout(n14322));
    jdff dff_A_u6mEIkBT1_1(.din(n14327), .dout(n14324));
    jdff dff_A_YprWSQXl2_1(.din(n14330), .dout(n14327));
    jdff dff_A_UQf0Whvu4_1(.din(n14333), .dout(n14330));
    jdff dff_A_8JQLu9eK9_1(.din(n14336), .dout(n14333));
    jdff dff_A_MkKKhlk65_1(.din(n14339), .dout(n14336));
    jdff dff_A_u5EHQxMO5_1(.din(n14342), .dout(n14339));
    jdff dff_A_LNrO9Vr24_1(.din(n14345), .dout(n14342));
    jdff dff_A_dRdZwZm91_1(.din(n14348), .dout(n14345));
    jdff dff_A_sUXL1Gpm1_1(.din(n14351), .dout(n14348));
    jdff dff_A_PSud7I7X4_1(.din(n14354), .dout(n14351));
    jdff dff_A_2nGnnnYf9_1(.din(n14357), .dout(n14354));
    jdff dff_A_nArJsp985_1(.din(n14360), .dout(n14357));
    jdff dff_A_h6TM1nLb0_1(.din(n14363), .dout(n14360));
    jdff dff_A_jl11dvRb3_1(.din(n14366), .dout(n14363));
    jdff dff_A_BuIuQJ7E7_1(.din(n14369), .dout(n14366));
    jdff dff_A_mlFn4RIz5_1(.din(n14372), .dout(n14369));
    jdff dff_A_mJUPKJal7_1(.din(n14375), .dout(n14372));
    jdff dff_A_kLbvHeRq5_1(.din(G4091), .dout(n14375));
    jdff dff_A_WWz6kItk5_2(.din(n14381), .dout(n14378));
    jdff dff_A_yoTy8XiB6_2(.din(n14384), .dout(n14381));
    jdff dff_A_FO2LjoWX8_2(.din(n14387), .dout(n14384));
    jdff dff_A_jRCz178b5_2(.din(n14390), .dout(n14387));
    jdff dff_A_H3iU3qlg3_2(.din(n14393), .dout(n14390));
    jdff dff_A_iDrou3bl9_2(.din(n14396), .dout(n14393));
    jdff dff_A_DVM9SFrA2_2(.din(n14399), .dout(n14396));
    jdff dff_A_bD7SVp1N3_2(.din(n14402), .dout(n14399));
    jdff dff_A_fxY25Nyx7_2(.din(n14405), .dout(n14402));
    jdff dff_A_m8eHBqdZ6_2(.din(G4091), .dout(n14405));
    jdff dff_A_vJ2Onia90_0(.din(n14411), .dout(n14408));
    jdff dff_A_fOBNq5Es2_0(.din(n4445), .dout(n14411));
    jdff dff_B_khmYPcgz9_1(.din(n4365), .dout(n14415));
    jdff dff_B_Cn27TpIJ0_1(.din(n14415), .dout(n14418));
    jdff dff_B_rhIZik0W9_1(.din(n4417), .dout(n14421));
    jdff dff_B_kRJT3wse7_1(.din(n4421), .dout(n14424));
    jdff dff_A_7Lv7AdWl5_1(.din(n760), .dout(n14426));
    jdff dff_A_ddU9OMzw0_0(.din(n14432), .dout(n14429));
    jdff dff_A_VW1wU9Xh5_0(.din(n14435), .dout(n14432));
    jdff dff_A_wK71iNMU8_0(.din(n14438), .dout(n14435));
    jdff dff_A_t8pGFjp86_0(.din(G503), .dout(n14438));
    jdff dff_A_MIQ1Y4FX5_1(.din(G503), .dout(n14441));
    jdff dff_A_THHCLd8W5_1(.din(n14447), .dout(n14444));
    jdff dff_A_uvjxOwaX1_1(.din(G503), .dout(n14447));
    jdff dff_A_C7If0JOz7_2(.din(n14453), .dout(n14450));
    jdff dff_A_y0LvTvBl1_2(.din(n14456), .dout(n14453));
    jdff dff_A_TIFXSPOy5_2(.din(n14459), .dout(n14456));
    jdff dff_A_Pru7XwWy6_2(.din(G503), .dout(n14459));
    jdff dff_A_2TCoX7101_1(.din(G324), .dout(n14462));
    jdff dff_A_o35FUYa91_1(.din(G324), .dout(n14465));
    jdff dff_B_j3XPcoFH2_1(.din(n4385), .dout(n14469));
    jdff dff_B_5XAEIhWx1_1(.din(n14469), .dout(n14472));
    jdff dff_A_x1spk4jM5_2(.din(n14478), .dout(n14474));
    jdff dff_B_Q4dSipxa8_3(.din(n621), .dout(n14478));
    jdff dff_A_5nmcFANn6_0(.din(n14483), .dout(n14480));
    jdff dff_A_gEgy98RR2_0(.din(n14486), .dout(n14483));
    jdff dff_A_hFq9wJpJ8_0(.din(G534), .dout(n14486));
    jdff dff_A_5qhikpfe9_1(.din(G534), .dout(n14489));
    jdff dff_B_aWUAzN4U2_1(.din(n4369), .dout(n14493));
    jdff dff_A_kJ1VNvQG9_1(.din(G351), .dout(n14495));
    jdff dff_A_cvrUomGe6_1(.din(n14501), .dout(n14498));
    jdff dff_A_1OY5sP727_1(.din(G534), .dout(n14501));
    jdff dff_A_VidaYrBB3_2(.din(n14507), .dout(n14504));
    jdff dff_A_xiyzJKe73_2(.din(n14510), .dout(n14507));
    jdff dff_A_0pFK2Ner1_2(.din(G534), .dout(n14510));
    jdff dff_A_OglsVBYO9_0(.din(G351), .dout(n14513));
    jdff dff_A_Rtj5CWw78_2(.din(n702), .dout(n14516));
    jdff dff_A_6st0OpoW4_1(.din(G514), .dout(n14519));
    jdff dff_A_FlZ0ONBZ3_2(.din(n14525), .dout(n14522));
    jdff dff_A_rhNxgrBE4_2(.din(G514), .dout(n14525));
    jdff dff_A_iMsQLFAt3_1(.din(G361), .dout(n14528));
    jdff dff_B_TBo6RMLm5_1(.din(n4330), .dout(n14532));
    jdff dff_B_Ywm0ecfJ3_1(.din(n14532), .dout(n14535));
    jdff dff_B_lAeKIlEP8_1(.din(n4334), .dout(n14538));
    jdff dff_B_Nsmg6kdC0_1(.din(n584), .dout(n14541));
    jdff dff_B_HrGeroVV9_1(.din(n588), .dout(n14544));
    jdff dff_A_T7u7M1HZ3_0(.din(n14549), .dout(n14546));
    jdff dff_A_TiknX4FY5_0(.din(n14552), .dout(n14549));
    jdff dff_A_4rgexoVy5_0(.din(G490), .dout(n14552));
    jdff dff_A_FWhTANMH7_1(.din(n14558), .dout(n14555));
    jdff dff_A_sGs16ISw7_1(.din(G490), .dout(n14558));
    jdff dff_A_yhl7EdmH5_1(.din(n14564), .dout(n14561));
    jdff dff_A_gzcDVFSt0_1(.din(n14567), .dout(n14564));
    jdff dff_A_eREKj2st1_1(.din(G490), .dout(n14567));
    jdff dff_A_LAxhXHmZ7_2(.din(n14573), .dout(n14570));
    jdff dff_A_fTEYH5MJ3_2(.din(n14576), .dout(n14573));
    jdff dff_A_4J7QjujL1_2(.din(G490), .dout(n14576));
    jdff dff_A_msxUPXKl5_0(.din(G316), .dout(n14579));
    jdff dff_B_DYaX8Hgu3_1(.din(n536), .dout(n14583));
    jdff dff_B_Ad7FIs4t6_1(.din(n543), .dout(n14586));
    jdff dff_A_HqRQQ5Dw3_0(.din(n14591), .dout(n14588));
    jdff dff_A_v2PmSzza2_0(.din(n14594), .dout(n14591));
    jdff dff_A_RvHiWXFc7_0(.din(n524), .dout(n14594));
    jdff dff_A_V2gQG1eZ7_0(.din(n14600), .dout(n14597));
    jdff dff_A_MvzDF7Oj4_0(.din(G479), .dout(n14600));
    jdff dff_A_C5PijlUF7_1(.din(n14606), .dout(n14603));
    jdff dff_A_GTBQ4FCe4_1(.din(n14609), .dout(n14606));
    jdff dff_A_1kxmuCHH2_1(.din(G479), .dout(n14609));
    jdff dff_A_DtmHDySL8_2(.din(n14615), .dout(n14612));
    jdff dff_A_swKeyPw01_2(.din(n14618), .dout(n14615));
    jdff dff_A_5hM7wWQg4_2(.din(G479), .dout(n14618));
    jdff dff_A_77KRC1lc4_0(.din(G308), .dout(n14621));
    jdff dff_A_4NWISi2H3_0(.din(G302), .dout(n14624));
    jdff dff_A_j41D3iUL7_1(.din(G302), .dout(n14627));
    jdff dff_A_9RxrP5xD1_0(.din(n671), .dout(n14630));
    jdff dff_A_USqn9juS4_2(.din(n671), .dout(n14633));
    jdff dff_A_rU5hIRg20_1(.din(G293), .dout(n14636));
    jdff dff_B_a2v8VoHg4_1(.din(n4310), .dout(n14640));
    jdff dff_B_nc06qPDF0_1(.din(n4314), .dout(n14643));
    jdff dff_A_X8JEPTvo8_0(.din(n802), .dout(n14645));
    jdff dff_A_SLhPDG6J2_2(.din(n14651), .dout(n14648));
    jdff dff_A_rVsBUueX2_2(.din(n802), .dout(n14651));
    jdff dff_A_QGecVUIb6_0(.din(G523), .dout(n14654));
    jdff dff_A_92YtTzxb0_1(.din(n14660), .dout(n14657));
    jdff dff_A_6KjX17et2_1(.din(n14663), .dout(n14660));
    jdff dff_A_6PiK53K50_1(.din(G523), .dout(n14663));
    jdff dff_A_RDUmUsws8_2(.din(n14669), .dout(n14666));
    jdff dff_A_zDMoByYg7_2(.din(G523), .dout(n14669));
    jdff dff_A_bcnZ5QXg4_1(.din(G341), .dout(n14672));
    jdff dff_A_8Kvxk1sW7_2(.din(G341), .dout(n14675));
    jdff dff_A_aze7x1926_2(.din(n14681), .dout(n14678));
    jdff dff_A_pFPTIqm75_2(.din(n14684), .dout(n14681));
    jdff dff_A_uZpT0iYG7_2(.din(n14687), .dout(n14684));
    jdff dff_A_hvkmYb9T5_2(.din(n14690), .dout(n14687));
    jdff dff_A_W4QeQyRj1_2(.din(n14693), .dout(n14690));
    jdff dff_A_yBmEkHR52_2(.din(n14696), .dout(n14693));
    jdff dff_A_ph5qFrFO9_2(.din(n14699), .dout(n14696));
    jdff dff_A_q9xs8aBf7_2(.din(n14702), .dout(n14699));
    jdff dff_A_IW8s2snX7_2(.din(n14705), .dout(n14702));
    jdff dff_A_rxs8mDsb4_2(.din(n14708), .dout(n14705));
    jdff dff_A_xCoe0Yxo1_2(.din(n1991), .dout(n14708));
    jdff dff_A_NLKlnGtd4_0(.din(n14714), .dout(n14711));
    jdff dff_A_HYLUqFkp4_0(.din(n14717), .dout(n14714));
    jdff dff_A_GYLgjmw42_0(.din(n14720), .dout(n14717));
    jdff dff_A_nm9NQ2Pf3_0(.din(n14723), .dout(n14720));
    jdff dff_A_EfLg9am28_0(.din(n14726), .dout(n14723));
    jdff dff_A_LW7Mt9wV8_0(.din(n2954), .dout(n14726));
    jdff dff_A_7eioFKEk0_2(.din(n14732), .dout(n14729));
    jdff dff_A_ZuuYbSaV3_2(.din(n14735), .dout(n14732));
    jdff dff_A_h1nyXclN6_2(.din(n14738), .dout(n14735));
    jdff dff_A_fdlHF7ir3_2(.din(n14741), .dout(n14738));
    jdff dff_A_HZ5IFSO28_2(.din(n14744), .dout(n14741));
    jdff dff_A_KF45V0xS4_2(.din(n14747), .dout(n14744));
    jdff dff_A_bISymSaK6_2(.din(n14750), .dout(n14747));
    jdff dff_A_taQFjGuE7_2(.din(n14753), .dout(n14750));
    jdff dff_A_Voo3CxCM6_2(.din(n14756), .dout(n14753));
    jdff dff_A_ND6PrY139_2(.din(n14759), .dout(n14756));
    jdff dff_A_Z9p8ucLv1_2(.din(n14762), .dout(n14759));
    jdff dff_A_AIgbrBNr3_2(.din(n14765), .dout(n14762));
    jdff dff_A_xLgZBadQ1_2(.din(n14768), .dout(n14765));
    jdff dff_A_RW3szw4Z4_2(.din(n14771), .dout(n14768));
    jdff dff_A_IjIs24Tj0_2(.din(n14774), .dout(n14771));
    jdff dff_A_kW6BxD995_2(.din(n14777), .dout(n14774));
    jdff dff_A_Ytz3WvXx7_2(.din(n14780), .dout(n14777));
    jdff dff_A_IDxTqGVC1_2(.din(n2954), .dout(n14780));
    jdff dff_A_Deyg2NPH8_1(.din(n14786), .dout(n14783));
    jdff dff_A_RMquG1VH5_1(.din(n14789), .dout(n14786));
    jdff dff_A_qAkVl2KR2_1(.din(n14792), .dout(n14789));
    jdff dff_A_S8Q5VEb37_1(.din(n14795), .dout(n14792));
    jdff dff_A_iGo2aX4h1_1(.din(n14798), .dout(n14795));
    jdff dff_A_QldryrM18_1(.din(n14801), .dout(n14798));
    jdff dff_A_OmHXET6u8_1(.din(n14804), .dout(n14801));
    jdff dff_A_afAF2FrS8_1(.din(n14807), .dout(n14804));
    jdff dff_A_zWIkN5RY2_1(.din(n14810), .dout(n14807));
    jdff dff_A_2CqVssKs0_1(.din(n14813), .dout(n14810));
    jdff dff_A_JreCyYxF9_1(.din(n14816), .dout(n14813));
    jdff dff_A_wYxPPXOo4_1(.din(n14819), .dout(n14816));
    jdff dff_A_7aE8ig800_1(.din(n14822), .dout(n14819));
    jdff dff_A_TH0PPm387_1(.din(n14825), .dout(n14822));
    jdff dff_A_zOfvnnl55_1(.din(n14828), .dout(n14825));
    jdff dff_A_32D0wbyv8_1(.din(n2954), .dout(n14828));
    jdff dff_A_wsDP1bJN1_2(.din(n14834), .dout(n14831));
    jdff dff_A_QRo3H8Pp1_2(.din(n14837), .dout(n14834));
    jdff dff_A_jk0adFD75_2(.din(n14840), .dout(n14837));
    jdff dff_A_FaY6W2PO3_2(.din(n14843), .dout(n14840));
    jdff dff_A_xchrOceB9_2(.din(n14846), .dout(n14843));
    jdff dff_A_SA6K04Ui8_2(.din(n14849), .dout(n14846));
    jdff dff_A_wXW4sHwz1_2(.din(n2954), .dout(n14849));
    jdff dff_B_D0CWybsJ3_1(.din(n5440), .dout(n14853));
    jdff dff_B_E9pVTg2h6_1(.din(n14853), .dout(n14856));
    jdff dff_B_gYfskHur3_1(.din(n14856), .dout(n14859));
    jdff dff_B_iYhTyRRk3_1(.din(n14859), .dout(n14862));
    jdff dff_B_Wik5T94l9_1(.din(n14862), .dout(n14865));
    jdff dff_B_f7yEEDOe6_1(.din(n14865), .dout(n14868));
    jdff dff_B_YNReeq394_1(.din(n14868), .dout(n14871));
    jdff dff_B_266Bsybs0_1(.din(n14871), .dout(n14874));
    jdff dff_B_U7qNGUDw4_1(.din(n14874), .dout(n14877));
    jdff dff_B_w8H034wv6_1(.din(n14877), .dout(n14880));
    jdff dff_B_obFN7baq1_1(.din(n14880), .dout(n14883));
    jdff dff_B_KqzyrakD9_1(.din(n14883), .dout(n14886));
    jdff dff_B_qhIFKDUt1_1(.din(n14886), .dout(n14889));
    jdff dff_B_403AIYZk7_1(.din(n14889), .dout(n14892));
    jdff dff_B_on9cbfOZ0_1(.din(n14892), .dout(n14895));
    jdff dff_B_AvbfHbsE0_1(.din(n14895), .dout(n14898));
    jdff dff_B_3cmqoIzR5_1(.din(n14898), .dout(n14901));
    jdff dff_B_BhU5I1SB5_1(.din(n14901), .dout(n14904));
    jdff dff_B_y6t5PHBq2_1(.din(n14904), .dout(n14907));
    jdff dff_B_m9RvD3KT2_0(.din(n5287), .dout(n14910));
    jdff dff_B_bAjPbLHg5_0(.din(n14910), .dout(n14913));
    jdff dff_B_t283aIEp3_0(.din(n14913), .dout(n14916));
    jdff dff_B_07k7FyeT2_0(.din(n14916), .dout(n14919));
    jdff dff_B_K80B8jMO0_0(.din(n14919), .dout(n14922));
    jdff dff_B_rThIxeqp0_0(.din(n14922), .dout(n14925));
    jdff dff_B_kbljello1_0(.din(n14925), .dout(n14928));
    jdff dff_B_sqNmiUWR4_0(.din(n14928), .dout(n14931));
    jdff dff_B_oeJrBfkf2_0(.din(n14931), .dout(n14934));
    jdff dff_B_dj564phh1_0(.din(n14934), .dout(n14937));
    jdff dff_B_eg3XnDXj7_0(.din(n14937), .dout(n14940));
    jdff dff_B_ruonKnZQ4_0(.din(n14940), .dout(n14943));
    jdff dff_B_jZD2Stwo6_0(.din(n14943), .dout(n14946));
    jdff dff_B_sb0Pk6hN5_0(.din(n14946), .dout(n14949));
    jdff dff_B_55jthq2E1_0(.din(n14949), .dout(n14952));
    jdff dff_B_qSjIQnq75_0(.din(n14952), .dout(n14955));
    jdff dff_B_ZCNmBO4p3_0(.din(n14955), .dout(n14958));
    jdff dff_B_bcAW2MU46_0(.din(n14958), .dout(n14961));
    jdff dff_B_CczamCeA6_0(.din(n14961), .dout(n14964));
    jdff dff_B_y6eSBI4b3_1(.din(n5055), .dout(n14967));
    jdff dff_B_cybQlxok1_1(.din(n14967), .dout(n14970));
    jdff dff_B_71f4yUDK4_1(.din(n14970), .dout(n14973));
    jdff dff_B_cMGm7CZg8_1(.din(n14973), .dout(n14976));
    jdff dff_B_5OhrnJ7w7_1(.din(n14976), .dout(n14979));
    jdff dff_B_cEHmt6JV6_1(.din(n14979), .dout(n14982));
    jdff dff_B_SSdPyBsD3_1(.din(n14982), .dout(n14985));
    jdff dff_B_JxnJFHBJ9_1(.din(n14985), .dout(n14988));
    jdff dff_B_voDq9m3C7_0(.din(n5245), .dout(n14991));
    jdff dff_B_OBkh3hor7_0(.din(n14991), .dout(n14994));
    jdff dff_B_Y0KUzQp49_1(.din(n5206), .dout(n14997));
    jdff dff_B_fDgFNn5p1_0(.din(n5233), .dout(n15000));
    jdff dff_B_HmHRIsmj7_0(.din(n15000), .dout(n15003));
    jdff dff_B_13uFmaH52_0(.din(n15003), .dout(n15006));
    jdff dff_B_8LDZHcFf0_0(.din(n5225), .dout(n15009));
    jdff dff_B_oHymJl9Z4_1(.din(n5158), .dout(n15012));
    jdff dff_B_p0OjHqQ14_1(.din(n15012), .dout(n15015));
    jdff dff_B_Oo98Fwqg2_1(.din(n15015), .dout(n15018));
    jdff dff_B_hvQyuDWe6_1(.din(n15018), .dout(n15021));
    jdff dff_B_kfga65Hg1_1(.din(n15021), .dout(n15024));
    jdff dff_B_oKx2tdWk3_1(.din(n15024), .dout(n15027));
    jdff dff_B_s6FttiPF9_1(.din(n15027), .dout(n15030));
    jdff dff_B_BK8bDYqc8_1(.din(n15030), .dout(n15033));
    jdff dff_B_NRoWvbCT3_1(.din(n15033), .dout(n15036));
    jdff dff_B_zJkuUrqE1_1(.din(n15036), .dout(n15039));
    jdff dff_B_CPYGXWMg6_1(.din(n15039), .dout(n15042));
    jdff dff_B_gm7OfTpl8_1(.din(n15042), .dout(n15045));
    jdff dff_B_KRgvwtkw4_1(.din(n15045), .dout(n15048));
    jdff dff_B_TWtG4G4Q2_1(.din(n5170), .dout(n15051));
    jdff dff_B_m5YzHZ2X8_1(.din(n15051), .dout(n15054));
    jdff dff_B_WWxDy1XO9_1(.din(n15054), .dout(n15057));
    jdff dff_B_ZEHe0Y898_1(.din(n15057), .dout(n15060));
    jdff dff_B_NyEhML011_1(.din(n5174), .dout(n15063));
    jdff dff_B_8v8wTRNY5_1(.din(n15063), .dout(n15066));
    jdff dff_B_PtQ18N2B6_1(.din(n15066), .dout(n15069));
    jdff dff_B_XIfNXhkf4_1(.din(n15069), .dout(n15072));
    jdff dff_B_GIHZRyBw4_1(.din(n15072), .dout(n15075));
    jdff dff_B_LvevyD0u7_1(.din(n15075), .dout(n15078));
    jdff dff_A_hEsPBp8w3_0(.din(n2402), .dout(n15080));
    jdff dff_A_1lupsNG66_1(.din(n15096), .dout(n15083));
    jdff dff_B_MtLqDPHt3_2(.din(n2394), .dout(n15087));
    jdff dff_B_Br1j1YCb7_2(.din(n15087), .dout(n15090));
    jdff dff_B_jurjrizg7_2(.din(n15090), .dout(n15093));
    jdff dff_B_kllcc4En5_2(.din(n15093), .dout(n15096));
    jdff dff_A_QxLJaRx41_0(.din(n15101), .dout(n15098));
    jdff dff_A_9O4EolNm4_0(.din(n15104), .dout(n15101));
    jdff dff_A_srsVW9Af9_0(.din(n15107), .dout(n15104));
    jdff dff_A_j8tzyT2m1_0(.din(n1740), .dout(n15107));
    jdff dff_A_jHm2wTS61_1(.din(n1740), .dout(n15110));
    jdff dff_A_zKmaTsBv8_1(.din(n5162), .dout(n15113));
    jdff dff_B_fiDJVqRi0_1(.din(n5139), .dout(n15117));
    jdff dff_B_9mibG71Y7_0(.din(n5143), .dout(n15120));
    jdff dff_B_IJNya5Rl8_1(.din(n5120), .dout(n15123));
    jdff dff_A_ikduT0UA6_0(.din(n15128), .dout(n15125));
    jdff dff_A_i0edykUa5_0(.din(n5113), .dout(n15128));
    jdff dff_B_LOnslHMK5_2(.din(n5105), .dout(n15132));
    jdff dff_B_KrP6ACxw1_2(.din(n15132), .dout(n15135));
    jdff dff_B_tMwK3bNH7_2(.din(n15135), .dout(n15138));
    jdff dff_B_JjpdH9y39_2(.din(n15138), .dout(n15141));
    jdff dff_B_bsSRZaF56_2(.din(n15141), .dout(n15144));
    jdff dff_B_bK8R2NEB5_2(.din(n15144), .dout(n15147));
    jdff dff_B_3kGxsvzi2_0(.din(n5097), .dout(n15150));
    jdff dff_B_IknBggBW4_0(.din(n15150), .dout(n15153));
    jdff dff_B_wrBjtwS76_0(.din(n15153), .dout(n15156));
    jdff dff_B_CCqndtHG8_0(.din(n5093), .dout(n15159));
    jdff dff_B_7ohlDYPp9_0(.din(n15159), .dout(n15162));
    jdff dff_B_e0AiH9RI4_0(.din(n15162), .dout(n15165));
    jdff dff_B_SCPpuGLX7_0(.din(n15165), .dout(n15168));
    jdff dff_B_3TEKFXjF7_0(.din(n15168), .dout(n15171));
    jdff dff_A_BSIOabYs3_2(.din(n15176), .dout(n15173));
    jdff dff_A_y1EzK1zt2_2(.din(n15179), .dout(n15176));
    jdff dff_A_wJ97G8MC0_2(.din(n15182), .dout(n15179));
    jdff dff_A_aKdImrnP2_2(.din(n15185), .dout(n15182));
    jdff dff_A_SsmDP4dU2_2(.din(n15188), .dout(n15185));
    jdff dff_A_l3KMi0Lf5_2(.din(n15191), .dout(n15188));
    jdff dff_A_YPhObIO37_2(.din(n15194), .dout(n15191));
    jdff dff_A_jWiQ0e9t3_2(.din(n15197), .dout(n15194));
    jdff dff_A_YYDdGiXM6_2(.din(n15200), .dout(n15197));
    jdff dff_A_aTQiV29g7_2(.din(n15203), .dout(n15200));
    jdff dff_A_jLfgwm3B2_2(.din(n15206), .dout(n15203));
    jdff dff_A_vtSVt5Ke4_2(.din(n1447), .dout(n15206));
    jdff dff_A_oxQIZz4S9_1(.din(n15212), .dout(n15209));
    jdff dff_A_GKLhhMUB8_1(.din(n15215), .dout(n15212));
    jdff dff_A_rrWg23Ee9_1(.din(n15218), .dout(n15215));
    jdff dff_A_ogIfQWlc6_1(.din(n15221), .dout(n15218));
    jdff dff_A_1syFJ1BI3_1(.din(n15224), .dout(n15221));
    jdff dff_A_wopdOaqf6_1(.din(n15227), .dout(n15224));
    jdff dff_A_Zw8N9znH7_1(.din(n15230), .dout(n15227));
    jdff dff_A_vvnwE0dB6_1(.din(n15233), .dout(n15230));
    jdff dff_A_JiOFjd856_1(.din(n2735), .dout(n15233));
    jdff dff_A_YA3kvibd3_2(.din(n15239), .dout(n15236));
    jdff dff_A_lcrB65fP0_2(.din(n15242), .dout(n15239));
    jdff dff_A_Dnw3qxl19_2(.din(n15245), .dout(n15242));
    jdff dff_A_HhCA1haI8_2(.din(n15248), .dout(n15245));
    jdff dff_A_myzx6miw8_2(.din(n15251), .dout(n15248));
    jdff dff_A_SuTsqUUz7_2(.din(n15254), .dout(n15251));
    jdff dff_A_lTS9xalW3_2(.din(n15257), .dout(n15254));
    jdff dff_A_xzbAIfva8_2(.din(n15260), .dout(n15257));
    jdff dff_A_DcNViKZO3_2(.din(n15267), .dout(n15260));
    jdff dff_B_8w9SjXgu8_3(.din(n2686), .dout(n15264));
    jdff dff_B_cNCEHzcg0_3(.din(n15264), .dout(n15267));
    jdff dff_A_QPJrCzQ94_1(.din(n15272), .dout(n15269));
    jdff dff_A_uQWcp82E3_1(.din(n15275), .dout(n15272));
    jdff dff_A_HcWZaaDr7_1(.din(n1813), .dout(n15275));
    jdff dff_A_RabxUM5u6_0(.din(n1837), .dout(n15278));
    jdff dff_B_LWfr27by0_1(.din(n1817), .dout(n15282));
    jdff dff_B_zHdUCnVa4_1(.din(n15282), .dout(n15285));
    jdff dff_B_0rl6XDgm3_0(.din(n1423), .dout(n15288));
    jdff dff_B_PV5733b09_1(.din(G233), .dout(n15291));
    jdff dff_B_yJUIuqCl3_2(.din(n1821), .dout(n15294));
    jdff dff_A_d2qPCzLc6_0(.din(n1443), .dout(n15296));
    jdff dff_B_IrYITDwn2_0(.din(n1439), .dout(n15300));
    jdff dff_B_I4f65N7O1_1(.din(G225), .dout(n15303));
    jdff dff_A_BSGd3JMX3_1(.din(n15308), .dout(n15305));
    jdff dff_A_3ESHHXks4_1(.din(n15311), .dout(n15308));
    jdff dff_A_cwv6t5gy6_1(.din(n15314), .dout(n15311));
    jdff dff_A_m14ZmyXb3_1(.din(n15317), .dout(n15314));
    jdff dff_A_SkQ9pSQd8_1(.din(n15320), .dout(n15317));
    jdff dff_A_jEfh31XR7_1(.din(n15323), .dout(n15320));
    jdff dff_A_mLPZdrPX1_1(.din(n15326), .dout(n15323));
    jdff dff_A_ifObSwrm4_1(.din(n15329), .dout(n15326));
    jdff dff_A_pCOCpnTh6_1(.din(n15339), .dout(n15329));
    jdff dff_B_jqKCjf4A8_2(.din(n2680), .dout(n15333));
    jdff dff_B_JLAvMhPP4_2(.din(n15333), .dout(n15336));
    jdff dff_B_tHW24P2b1_2(.din(n15336), .dout(n15339));
    jdff dff_A_0flIumw26_0(.din(n15344), .dout(n15341));
    jdff dff_A_NFa9gf9t3_0(.din(n15347), .dout(n15344));
    jdff dff_A_PfRuB1eH7_0(.din(n15350), .dout(n15347));
    jdff dff_A_S5K49NIm7_0(.din(n15353), .dout(n15350));
    jdff dff_A_09eiEXdN9_0(.din(n1411), .dout(n15353));
    jdff dff_B_p3feOSO34_1(.din(n1396), .dout(n15357));
    jdff dff_B_WCFRpAvJ0_1(.din(G209), .dout(n15360));
    jdff dff_B_6kfQng679_0(.din(n5070), .dout(n15363));
    jdff dff_A_ZUHGbJNA8_0(.din(n1369), .dout(n15365));
    jdff dff_B_CbaEUmP63_0(.din(n1365), .dout(n15369));
    jdff dff_B_SDAncjIu4_0(.din(n15369), .dout(n15372));
    jdff dff_A_7dpqGCjC5_0(.din(n15377), .dout(n15374));
    jdff dff_A_x5NtLHI71_0(.din(n15380), .dout(n15377));
    jdff dff_A_bnNVtO9w5_0(.din(n1361), .dout(n15380));
    jdff dff_A_63KvYAOB7_0(.din(n15386), .dout(n15383));
    jdff dff_A_BPpn6oSc2_0(.din(n15389), .dout(n15386));
    jdff dff_A_JRHCN90s7_0(.din(n15392), .dout(n15389));
    jdff dff_A_EXbfzPrL4_0(.din(n1319), .dout(n15392));
    jdff dff_A_P8xOK5uz1_1(.din(n1300), .dout(n15395));
    jdff dff_A_uK6OIkPM0_1(.din(n15401), .dout(n15398));
    jdff dff_A_wIlEuhuF7_1(.din(n15404), .dout(n15401));
    jdff dff_A_9WJodyuM8_1(.din(n1300), .dout(n15404));
    jdff dff_A_IwN1l2Xb1_0(.din(n15995), .dout(n15407));
    jdff dff_A_fMctWRTU0_0(.din(n15413), .dout(n15410));
    jdff dff_A_92dWOa9m5_0(.din(n15416), .dout(n15413));
    jdff dff_A_zTGz7cTw7_0(.din(n15419), .dout(n15416));
    jdff dff_A_mMMU0x3m6_0(.din(n15422), .dout(n15419));
    jdff dff_A_YLbN2nBA3_0(.din(n15429), .dout(n15422));
    jdff dff_B_Q17ELFLL2_2(.din(n1281), .dout(n15426));
    jdff dff_B_f1SPZpZX8_2(.din(n15426), .dout(n15429));
    jdff dff_A_LT7SfRtI1_0(.din(n1278), .dout(n15431));
    jdff dff_A_QeGAPcQN6_1(.din(n15437), .dout(n15434));
    jdff dff_A_TYKPX5VY6_1(.din(n15440), .dout(n15437));
    jdff dff_A_Q094VyXA8_1(.din(n1278), .dout(n15440));
    jdff dff_A_ZrUszQjG6_0(.din(n15446), .dout(n15443));
    jdff dff_A_5X3yEdkl6_0(.din(n15449), .dout(n15446));
    jdff dff_A_GrRXcfIM7_0(.din(n15452), .dout(n15449));
    jdff dff_A_Bb9lsqzh5_0(.din(n15455), .dout(n15452));
    jdff dff_A_kEMwIXIn5_0(.din(n15458), .dout(n15455));
    jdff dff_A_0Fa8os3z7_0(.din(n15461), .dout(n15458));
    jdff dff_A_FS4Kxid42_0(.din(n15464), .dout(n15461));
    jdff dff_A_oWUaqytK7_0(.din(n15467), .dout(n15464));
    jdff dff_A_dG2Mjsc11_0(.din(n15470), .dout(n15467));
    jdff dff_A_eSrgxN3W7_0(.din(n15473), .dout(n15470));
    jdff dff_A_OYUQNdxS0_0(.din(n15476), .dout(n15473));
    jdff dff_A_JqaM0uqn6_0(.din(G1497), .dout(n15476));
    jdff dff_A_JIsGZ0Ow2_2(.din(n15482), .dout(n15479));
    jdff dff_A_UsYkc8JY3_2(.din(n15485), .dout(n15482));
    jdff dff_A_bFLN5keE7_2(.din(n15488), .dout(n15485));
    jdff dff_A_2PVSg64j2_2(.din(n15491), .dout(n15488));
    jdff dff_A_kdVLLeTI5_2(.din(n15494), .dout(n15491));
    jdff dff_A_t9pvmhFv2_2(.din(n15497), .dout(n15494));
    jdff dff_A_PU2cSZfk8_2(.din(n15500), .dout(n15497));
    jdff dff_A_pMmppbiq0_2(.din(n15503), .dout(n15500));
    jdff dff_A_er9MN6VG4_2(.din(n15506), .dout(n15503));
    jdff dff_A_EWHZ9Osq4_2(.din(G1497), .dout(n15506));
    jdff dff_B_oq0Ywofd2_1(.din(n1717), .dout(n15510));
    jdff dff_B_gZDI64Ns3_1(.din(n15510), .dout(n15513));
    jdff dff_B_7T1LkwOg9_1(.din(n15513), .dout(n15516));
    jdff dff_B_ahsHh9Ol7_1(.din(n15516), .dout(n15519));
    jdff dff_B_CbbG04359_1(.din(n1721), .dout(n15522));
    jdff dff_B_bOYmoYFs5_1(.din(n15522), .dout(n15525));
    jdff dff_B_Xz7zCVNm5_1(.din(n15525), .dout(n15528));
    jdff dff_B_9hso8GXL7_1(.din(n15528), .dout(n15531));
    jdff dff_B_1PaqHFXG2_1(.din(n15531), .dout(n15534));
    jdff dff_A_8v12xvBk6_1(.din(n1778), .dout(n15536));
    jdff dff_A_JOLCGD738_0(.din(n1770), .dout(n15539));
    jdff dff_A_NiKCeGge1_0(.din(n1762), .dout(n15542));
    jdff dff_A_hVs7x4Xo4_1(.din(n15548), .dout(n15545));
    jdff dff_A_qTLdxIJi4_1(.din(n15551), .dout(n15548));
    jdff dff_A_ssmlvYDc9_1(.din(n15554), .dout(n15551));
    jdff dff_A_EvD6p0zS9_1(.din(n1762), .dout(n15554));
    jdff dff_A_VD5hiWkc2_2(.din(n15560), .dout(n15557));
    jdff dff_A_4yccVk0V6_2(.din(n15563), .dout(n15560));
    jdff dff_A_9prX5OOG0_2(.din(n1316), .dout(n15563));
    jdff dff_A_SU22FOku6_1(.din(n1308), .dout(n15566));
    jdff dff_A_dIXvuexv7_1(.din(G280), .dout(n15569));
    jdff dff_A_iqc2tmVP1_0(.din(n15893), .dout(n15572));
    jdff dff_A_pe5x4dCf1_0(.din(n15578), .dout(n15575));
    jdff dff_A_CZu92rYw1_0(.din(n1740), .dout(n15578));
    jdff dff_A_Vpom8c187_1(.din(n15585), .dout(n15581));
    jdff dff_B_97Od1iLj9_2(.din(n1736), .dout(n15585));
    jdff dff_A_rdwYEB797_0(.din(n15956), .dout(n15587));
    jdff dff_A_BUnEjW585_1(.din(n15593), .dout(n15590));
    jdff dff_A_EeOODEu20_1(.din(n1732), .dout(n15593));
    jdff dff_A_LoROC9dG1_1(.din(n15599), .dout(n15596));
    jdff dff_A_6jdQc28D4_1(.din(n15602), .dout(n15599));
    jdff dff_A_cdBdRrEJ6_1(.din(n1728), .dout(n15602));
    jdff dff_B_c5b0SisU2_1(.din(n1263), .dout(n15606));
    jdff dff_B_OdDnxJVz1_1(.din(G241), .dout(n15609));
    jdff dff_B_nYHrPa6X7_2(.din(n5066), .dout(n15612));
    jdff dff_B_NCF2avyc2_2(.din(n15612), .dout(n15615));
    jdff dff_B_70esU5vR8_2(.din(n15615), .dout(n15618));
    jdff dff_B_8sWR1LZ04_2(.din(n15618), .dout(n15621));
    jdff dff_B_MNvJXFBW1_2(.din(n15621), .dout(n15624));
    jdff dff_B_rABvzCqa6_2(.din(n15624), .dout(n15627));
    jdff dff_B_piFvOyF13_2(.din(n15627), .dout(n15630));
    jdff dff_B_FvrOhXZl9_2(.din(n15630), .dout(n15633));
    jdff dff_B_BIDd6ZH78_2(.din(n15633), .dout(n15636));
    jdff dff_B_4ofr7wj29_2(.din(n15636), .dout(n15639));
    jdff dff_A_fAbKqvX35_2(.din(n15644), .dout(n15641));
    jdff dff_A_OQaTlxtk6_2(.din(n15647), .dout(n15644));
    jdff dff_A_uMBcqh5w8_2(.din(n15650), .dout(n15647));
    jdff dff_A_96EIOfti0_2(.din(n15653), .dout(n15650));
    jdff dff_A_OVx7vuIf6_2(.din(n1361), .dout(n15653));
    jdff dff_A_3W9nTXQe8_1(.din(n15659), .dout(n15656));
    jdff dff_A_CZc7oxpZ0_1(.din(n15662), .dout(n15659));
    jdff dff_A_p16N9eAf4_1(.din(n15665), .dout(n15662));
    jdff dff_A_IRvJ5n7H9_1(.din(n15668), .dout(n15665));
    jdff dff_A_mRHePuIw5_1(.din(n15671), .dout(n15668));
    jdff dff_A_ZM6t2rqF7_1(.din(n15674), .dout(n15671));
    jdff dff_A_nLtBEqxt1_1(.din(n1342), .dout(n15674));
    jdff dff_B_y2DrAnYB0_0(.din(n1334), .dout(n15678));
    jdff dff_A_X5VE5Rn87_0(.din(G335), .dout(n15680));
    jdff dff_B_ex8iQiFj3_1(.din(G264), .dout(n15684));
    jdff dff_A_I48WH7cW8_0(.din(n15689), .dout(n15686));
    jdff dff_A_xwueaaXp8_0(.din(n15930), .dout(n15689));
    jdff dff_A_3XYAaoiY3_1(.din(n15930), .dout(n15692));
    jdff dff_A_BBMmeLKm0_1(.din(n15698), .dout(n15695));
    jdff dff_A_rEbBXL8M5_1(.din(n15701), .dout(n15698));
    jdff dff_A_gq866Uyx9_1(.din(n15704), .dout(n15701));
    jdff dff_A_iFiqIPSR9_1(.din(n15707), .dout(n15704));
    jdff dff_A_pTzrZNO72_1(.din(n15710), .dout(n15707));
    jdff dff_A_habZwT1r8_1(.din(n15713), .dout(n15710));
    jdff dff_A_hLTnTAOU5_1(.din(n15716), .dout(n15713));
    jdff dff_A_huzUM75a1_1(.din(n15719), .dout(n15716));
    jdff dff_A_wi0ZbLkl6_1(.din(n15722), .dout(n15719));
    jdff dff_A_n8KaUCZM2_1(.din(n15725), .dout(n15722));
    jdff dff_A_3kVqWks17_1(.din(n15728), .dout(n15725));
    jdff dff_A_rc6cyPT01_1(.din(n2732), .dout(n15728));
    jdff dff_A_nJ2td3iY0_1(.din(n1392), .dout(n15731));
    jdff dff_A_Gt3ZoqjV6_1(.din(n15737), .dout(n15734));
    jdff dff_A_K7sE6wq35_1(.din(n1388), .dout(n15737));
    jdff dff_B_7O06H6yB2_0(.din(n1384), .dout(n15741));
    jdff dff_B_oSc3NJlp1_1(.din(G217), .dout(n15744));
    jdff dff_A_Y0C5iHwL0_0(.din(G335), .dout(n15746));
    jdff dff_A_6CHDTV882_2(.din(G335), .dout(n15749));
    jdff dff_A_SJM3llbf3_1(.din(n15755), .dout(n15752));
    jdff dff_A_u8JSnDQi1_1(.din(n15758), .dout(n15755));
    jdff dff_A_il7T7hol3_1(.din(n15761), .dout(n15758));
    jdff dff_A_IV7T04QO9_1(.din(n15764), .dout(n15761));
    jdff dff_A_NgP28wni9_1(.din(n15767), .dout(n15764));
    jdff dff_A_cuQLzaUW8_1(.din(n15770), .dout(n15767));
    jdff dff_A_bmyElyw24_1(.din(n15773), .dout(n15770));
    jdff dff_A_2ljb2NLh7_1(.din(n15776), .dout(n15773));
    jdff dff_A_1pPdm0Gj8_1(.din(n15779), .dout(n15776));
    jdff dff_A_830R7nnO7_1(.din(n15782), .dout(n15779));
    jdff dff_A_HWW4jZFn9_1(.din(n15785), .dout(n15782));
    jdff dff_A_nFQtPAcr9_1(.din(n15788), .dout(n15785));
    jdff dff_A_8s4z32cf7_1(.din(n15791), .dout(n15788));
    jdff dff_A_zfGaarHY9_1(.din(n15794), .dout(n15791));
    jdff dff_A_EdWZtHnH2_1(.din(n15797), .dout(n15794));
    jdff dff_A_zQQQTv6k9_1(.din(n15800), .dout(n15797));
    jdff dff_A_vGWoQ90w7_1(.din(n2005), .dout(n15800));
    jdff dff_A_HAUkrzKr3_2(.din(n15806), .dout(n15803));
    jdff dff_A_U6v1aeNf5_2(.din(n15809), .dout(n15806));
    jdff dff_A_G3jFXJA17_2(.din(n15812), .dout(n15809));
    jdff dff_A_n6Sv8eHr5_2(.din(n15815), .dout(n15812));
    jdff dff_A_uuHG5Q250_2(.din(n15818), .dout(n15815));
    jdff dff_A_Ru9HNxHt3_2(.din(n15821), .dout(n15818));
    jdff dff_A_uAOJH08I9_2(.din(n15824), .dout(n15821));
    jdff dff_A_NYquPSHS8_2(.din(n2005), .dout(n15824));
    jdff dff_A_5GaXf1406_2(.din(G4091), .dout(n15827));
    jdff dff_A_pMnAPbPy2_2(.din(n15833), .dout(n15830));
    jdff dff_A_fUn5nLBT4_2(.din(n15836), .dout(n15833));
    jdff dff_A_s5nuRzJv2_2(.din(n15839), .dout(n15836));
    jdff dff_A_VThthqik6_2(.din(n15842), .dout(n15839));
    jdff dff_A_zxu4Y6xJ2_2(.din(n15845), .dout(n15842));
    jdff dff_A_2vUuaBgp4_2(.din(n15848), .dout(n15845));
    jdff dff_A_wnUidp9P8_2(.din(n15851), .dout(n15848));
    jdff dff_A_GkHTtTX37_2(.din(n15854), .dout(n15851));
    jdff dff_A_9KWaRm4D7_2(.din(n15857), .dout(n15854));
    jdff dff_A_gV6NFZlV5_2(.din(n15860), .dout(n15857));
    jdff dff_A_vaajNmmr9_2(.din(n15863), .dout(n15860));
    jdff dff_A_xCnhGROG9_2(.din(n15866), .dout(n15863));
    jdff dff_A_ydaMKyjA1_2(.din(n15869), .dout(n15866));
    jdff dff_A_COWnrVOF2_2(.din(n15872), .dout(n15869));
    jdff dff_A_0n8QOOed6_2(.din(n15875), .dout(n15872));
    jdff dff_A_QMHeXJpH0_2(.din(n15878), .dout(n15875));
    jdff dff_A_2K3aXCom4_2(.din(n15881), .dout(n15878));
    jdff dff_A_mDT9zZ7v2_2(.din(G4091), .dout(n15881));
    jdff dff_B_otbjf07u4_2(.din(n5028), .dout(n15885));
    jdff dff_B_m1R52wP16_1(.din(n5000), .dout(n15888));
    jdff dff_B_AJTqV7fd2_1(.din(n5004), .dout(n15891));
    jdff dff_A_1YbHecmV2_0(.din(n990), .dout(n15893));
    jdff dff_A_posRy3dw0_2(.din(n15899), .dout(n15896));
    jdff dff_A_8RSXgteW1_2(.din(n990), .dout(n15899));
    jdff dff_A_d064H4t07_0(.din(n15905), .dout(n15902));
    jdff dff_A_Zw8gwf5R7_0(.din(G411), .dout(n15905));
    jdff dff_A_6BR4DVNt6_1(.din(G411), .dout(n15908));
    jdff dff_A_HlJL891t2_1(.din(G273), .dout(n15911));
    jdff dff_A_rbLJ0fbJ2_2(.din(G273), .dout(n15914));
    jdff dff_B_YIiBl1PT1_1(.din(n4968), .dout(n15918));
    jdff dff_B_pwRFMlrp9_1(.din(n15918), .dout(n15921));
    jdff dff_A_VieoZLRK7_2(.din(n15926), .dout(n15923));
    jdff dff_A_yQsZz6LY3_2(.din(n15930), .dout(n15926));
    jdff dff_B_c5M0faWB5_3(.din(n940), .dout(n15930));
    jdff dff_B_s5CmWdDh1_1(.din(n4952), .dout(n15933));
    jdff dff_A_KFQivGam9_1(.din(G257), .dout(n15935));
    jdff dff_A_PP7ffUZ67_0(.din(n15941), .dout(n15938));
    jdff dff_A_ntbxNQMz8_0(.din(G389), .dout(n15941));
    jdff dff_A_G0yvkdsE8_1(.din(G389), .dout(n15944));
    jdff dff_A_0vmrnqG67_0(.din(G257), .dout(n15947));
    jdff dff_B_8WJiVgDg4_1(.din(n4924), .dout(n15951));
    jdff dff_B_dA7S9O0q4_1(.din(n4928), .dout(n15954));
    jdff dff_A_yzVfqSoE5_0(.din(n856), .dout(n15956));
    jdff dff_A_XPcdGorN6_2(.din(n15962), .dout(n15959));
    jdff dff_A_C9wiUB3i5_2(.din(n856), .dout(n15962));
    jdff dff_A_SQiowSOU1_0(.din(G400), .dout(n15965));
    jdff dff_A_KwfjedKL4_1(.din(n15971), .dout(n15968));
    jdff dff_A_LR4UwY9l0_1(.din(G400), .dout(n15971));
    jdff dff_A_ttdzmNqI7_2(.din(n15977), .dout(n15974));
    jdff dff_A_rSBlSYSC0_2(.din(n15980), .dout(n15977));
    jdff dff_A_bodr78eO0_2(.din(G400), .dout(n15980));
    jdff dff_A_GHf1WuLw3_0(.din(G265), .dout(n15983));
    jdff dff_A_e3JIbNxC8_2(.din(G265), .dout(n15986));
    jdff dff_B_F7dSwWAA2_1(.din(n4888), .dout(n15990));
    jdff dff_B_t4xIJt4T5_1(.din(n4892), .dout(n15993));
    jdff dff_A_CQDvDQIN0_0(.din(n1032), .dout(n15995));
    jdff dff_A_KbGIdVt48_2(.din(n16001), .dout(n15998));
    jdff dff_A_53wdL9Ic4_2(.din(n1032), .dout(n16001));
    jdff dff_A_ZMRooXgA5_0(.din(n16007), .dout(n16004));
    jdff dff_A_jk4Zfurw9_0(.din(G374), .dout(n16007));
    jdff dff_A_rrQKLtgY1_1(.din(G374), .dout(n16010));
    jdff dff_A_zwQWhkLL1_0(.din(G281), .dout(n16013));
    jdff dff_A_Z2ld8Ms42_2(.din(G281), .dout(n16016));
    jdff dff_B_CggUUJyJ9_1(.din(n4748), .dout(n16020));
    jdff dff_B_McPhVsr13_1(.din(n16020), .dout(n16023));
    jdff dff_B_M2BfNANf4_1(.din(n4840), .dout(n16026));
    jdff dff_B_xqQZZMkN9_1(.din(n4844), .dout(n16029));
    jdff dff_A_2Fos1n793_1(.din(G210), .dout(n16031));
    jdff dff_A_K1sSTTDM4_1(.din(n1208), .dout(n16034));
    jdff dff_A_PpQBE0k26_0(.din(G457), .dout(n16037));
    jdff dff_A_ikHJwaSR6_0(.din(n16043), .dout(n16040));
    jdff dff_A_5utZaRT63_0(.din(n16046), .dout(n16043));
    jdff dff_A_kIlLJhno4_0(.din(G457), .dout(n16046));
    jdff dff_A_uzNAGVgL4_2(.din(n16052), .dout(n16049));
    jdff dff_A_NIHaGDVF2_2(.din(G457), .dout(n16052));
    jdff dff_A_Wvhep0ki2_1(.din(G210), .dout(n16055));
    jdff dff_A_W0Bp2O9F7_2(.din(G210), .dout(n16058));
    jdff dff_B_drKLrYsS4_1(.din(n4808), .dout(n16062));
    jdff dff_B_p5kmLarl3_1(.din(n16062), .dout(n16065));
    jdff dff_B_juMTaES87_2(.din(n1078), .dout(n16068));
    jdff dff_A_FCoTUeF00_0(.din(n16073), .dout(n16070));
    jdff dff_A_X5buWeyf0_0(.din(n16076), .dout(n16073));
    jdff dff_A_P62yhVsH3_0(.din(G468), .dout(n16076));
    jdff dff_A_6D3Di4A10_1(.din(G468), .dout(n16079));
    jdff dff_B_rzADqUVV1_1(.din(n4792), .dout(n16083));
    jdff dff_A_sblDCa1a4_1(.din(G218), .dout(n16085));
    jdff dff_A_8XrAwFnq4_1(.din(n16091), .dout(n16088));
    jdff dff_A_IcWadWZz6_1(.din(G468), .dout(n16091));
    jdff dff_A_u3XK0Zs11_2(.din(n16097), .dout(n16094));
    jdff dff_A_KoCm3FHP7_2(.din(n16100), .dout(n16097));
    jdff dff_A_KNLrAf8K1_2(.din(G468), .dout(n16100));
    jdff dff_A_9a9Fd7d06_0(.din(G218), .dout(n16103));
    jdff dff_B_vP9uQ1Iv3_1(.din(n4768), .dout(n16107));
    jdff dff_B_Z0Onc9aE6_1(.din(n16107), .dout(n16110));
    jdff dff_B_E0EfueVk5_2(.din(n1166), .dout(n16113));
    jdff dff_A_dTobYgT19_0(.din(G422), .dout(n16115));
    jdff dff_B_PS8UhcAt3_1(.din(n4752), .dout(n16119));
    jdff dff_A_8jIdLr0h7_1(.din(G226), .dout(n16121));
    jdff dff_A_Hs8KFHmw9_0(.din(n16127), .dout(n16124));
    jdff dff_A_bi0OmC4g3_0(.din(n16130), .dout(n16127));
    jdff dff_A_dQHbuo6n9_0(.din(G422), .dout(n16130));
    jdff dff_A_1yF74THA3_2(.din(n16136), .dout(n16133));
    jdff dff_A_TPUCpvG71_2(.din(G422), .dout(n16136));
    jdff dff_A_g05iV4qr9_1(.din(G251), .dout(n16139));
    jdff dff_A_umsvQfiS2_2(.din(G251), .dout(n16142));
    jdff dff_A_K6d3lJfk5_1(.din(G251), .dout(n16145));
    jdff dff_A_CwMNRSJ39_2(.din(G251), .dout(n16148));
    jdff dff_A_6CZxVukQ2_0(.din(G226), .dout(n16151));
    jdff dff_B_J4fIGD0M8_1(.din(n1132), .dout(n16155));
    jdff dff_B_jPvxMSUl7_1(.din(n1136), .dout(n16158));
    jdff dff_A_a3DYy5kJ1_0(.din(n16163), .dout(n16160));
    jdff dff_A_WDwUZNW40_0(.din(n16166), .dout(n16163));
    jdff dff_A_JOkU9xyp2_0(.din(n16169), .dout(n16166));
    jdff dff_A_5RAOQJeX5_0(.din(G446), .dout(n16169));
    jdff dff_A_RDfsVM6X2_1(.din(n16175), .dout(n16172));
    jdff dff_A_PjIXy07J6_1(.din(G446), .dout(n16175));
    jdff dff_A_L84Mh0M65_1(.din(n16181), .dout(n16178));
    jdff dff_A_1SfBBiXl2_1(.din(n16184), .dout(n16181));
    jdff dff_A_WTBqrzoc1_1(.din(n16187), .dout(n16184));
    jdff dff_A_G6lbEGdA0_1(.din(G446), .dout(n16187));
    jdff dff_A_pJCGRX3l2_2(.din(n16193), .dout(n16190));
    jdff dff_A_WL2r15fE7_2(.din(n16196), .dout(n16193));
    jdff dff_A_yGjiDEl32_2(.din(n16199), .dout(n16196));
    jdff dff_A_jWocplEn0_2(.din(G446), .dout(n16199));
    jdff dff_A_4WsIfzAC9_0(.din(G206), .dout(n16202));
    jdff dff_B_PzdBPeFS4_1(.din(n4728), .dout(n16206));
    jdff dff_B_ESW2Jyin8_1(.din(n4732), .dout(n16209));
    jdff dff_A_cQwm38V27_0(.din(G242), .dout(n16211));
    jdff dff_A_Q5zt9qC28_1(.din(G242), .dout(n16214));
    jdff dff_A_HpUvt8bN7_1(.din(G242), .dout(n16217));
    jdff dff_A_L1bi1yru6_2(.din(G242), .dout(n16220));
    jdff dff_A_iVswdcIQ0_2(.din(G248), .dout(n16223));
    jdff dff_A_zsQn6rAz9_1(.din(n16229), .dout(n16226));
    jdff dff_A_6xE1kp3C5_1(.din(n16232), .dout(n16229));
    jdff dff_A_yPEI7Z7s6_1(.din(n16235), .dout(n16232));
    jdff dff_A_IxdqBATw2_1(.din(n898), .dout(n16235));
    jdff dff_A_CvTLzAgQ6_2(.din(n898), .dout(n16238));
    jdff dff_A_145FCC1R1_0(.din(n16244), .dout(n16241));
    jdff dff_A_E0jDH5bB5_0(.din(n16247), .dout(n16244));
    jdff dff_A_9326LpdF4_0(.din(n16250), .dout(n16247));
    jdff dff_A_BKERlw5H5_0(.din(G435), .dout(n16250));
    jdff dff_A_93DnRBLx5_1(.din(G435), .dout(n16253));
    jdff dff_A_6JXrWEu75_1(.din(n16259), .dout(n16256));
    jdff dff_A_fxjrjCh67_1(.din(G435), .dout(n16259));
    jdff dff_A_jKyhf4HO5_2(.din(n16265), .dout(n16262));
    jdff dff_A_3rQhbg9g1_2(.din(n16268), .dout(n16265));
    jdff dff_A_1AEaBP9I6_2(.din(n16271), .dout(n16268));
    jdff dff_A_93tWPI9q8_2(.din(G435), .dout(n16271));
    jdff dff_A_xBie47Qk2_1(.din(G251), .dout(n16274));
    jdff dff_A_EmzcZY9t8_2(.din(G251), .dout(n16277));
    jdff dff_A_y5HQIe6X9_0(.din(G234), .dout(n16280));
    jdff dff_A_5gdKQzfI4_2(.din(G234), .dout(n16283));
    jdff dff_A_MYR8O7PY4_0(.din(n16289), .dout(n16286));
    jdff dff_A_tBnMUCjT0_0(.din(n16292), .dout(n16289));
    jdff dff_A_ca1oavqp1_0(.din(n16295), .dout(n16292));
    jdff dff_A_gnnwhmDU5_0(.din(n16298), .dout(n16295));
    jdff dff_A_mzXovG4n0_0(.din(n16301), .dout(n16298));
    jdff dff_A_0hup6JtJ1_0(.din(n16304), .dout(n16301));
    jdff dff_A_s8Cwsbp59_0(.din(n16307), .dout(n16304));
    jdff dff_A_9J9gV7LA9_0(.din(n16310), .dout(n16307));
    jdff dff_A_UMSDBrGl4_0(.din(n16313), .dout(n16310));
    jdff dff_A_vPrnZUAq7_0(.din(n16316), .dout(n16313));
    jdff dff_A_c9obuGxY8_0(.din(G4092), .dout(n16316));
    jdff dff_A_zdrI3PDS9_1(.din(G4092), .dout(n16319));
    jdff dff_A_BoMi0olI2_0(.din(n16325), .dout(n16322));
    jdff dff_A_nvTaLphW4_0(.din(n16328), .dout(n16325));
    jdff dff_A_QsJjPFXN5_0(.din(n16331), .dout(n16328));
    jdff dff_A_j3O89ShG0_0(.din(n16334), .dout(n16331));
    jdff dff_A_S0vDBA0J9_0(.din(n16337), .dout(n16334));
    jdff dff_A_iW9HFaD08_0(.din(n16340), .dout(n16337));
    jdff dff_A_rrccWHtp0_0(.din(n2943), .dout(n16340));
    jdff dff_A_Ikjyje7n8_2(.din(n16346), .dout(n16343));
    jdff dff_A_TOXxie9F4_2(.din(n16349), .dout(n16346));
    jdff dff_A_apl4wpDY6_2(.din(n16352), .dout(n16349));
    jdff dff_A_WaRh8NRP3_2(.din(n16355), .dout(n16352));
    jdff dff_A_fYJv7fYP2_2(.din(n16358), .dout(n16355));
    jdff dff_A_lIlX7Wn50_2(.din(n16361), .dout(n16358));
    jdff dff_A_LJliNtAy7_2(.din(n16364), .dout(n16361));
    jdff dff_A_1bp8sStG3_2(.din(n16367), .dout(n16364));
    jdff dff_A_3DLSZKbP5_2(.din(n16370), .dout(n16367));
    jdff dff_A_mYHbTfFD9_2(.din(n16373), .dout(n16370));
    jdff dff_A_szsVc30w8_2(.din(n16376), .dout(n16373));
    jdff dff_A_F3pXSx5e6_2(.din(n16379), .dout(n16376));
    jdff dff_A_MUqtxYMl0_2(.din(n16382), .dout(n16379));
    jdff dff_A_WcsDrtic9_2(.din(n16385), .dout(n16382));
    jdff dff_A_IvX1SISW3_2(.din(n16388), .dout(n16385));
    jdff dff_A_lAQC2soE4_2(.din(n16391), .dout(n16388));
    jdff dff_A_tRXZgcD47_2(.din(n16394), .dout(n16391));
    jdff dff_A_ZKRb0Opf1_2(.din(n16397), .dout(n16394));
    jdff dff_A_A9I8q0GE3_2(.din(n2943), .dout(n16397));
    jdff dff_A_ppyogrIt4_1(.din(n16403), .dout(n16400));
    jdff dff_A_8b3QS6fT7_1(.din(n16406), .dout(n16403));
    jdff dff_A_uJdOCJWZ0_1(.din(n16409), .dout(n16406));
    jdff dff_A_Ie5jSKVK5_1(.din(n16412), .dout(n16409));
    jdff dff_A_b6C8S39j3_1(.din(n16415), .dout(n16412));
    jdff dff_A_ciBTzmfd6_1(.din(n16418), .dout(n16415));
    jdff dff_A_7wqJ9Bsa1_1(.din(n16421), .dout(n16418));
    jdff dff_A_VVDAx3uY1_1(.din(n16424), .dout(n16421));
    jdff dff_A_AD2tdsOF8_1(.din(n16427), .dout(n16424));
    jdff dff_A_4Xvbbywf5_1(.din(n16430), .dout(n16427));
    jdff dff_A_quyEqx870_1(.din(n16433), .dout(n16430));
    jdff dff_A_SJc8o4by1_1(.din(n16436), .dout(n16433));
    jdff dff_A_M7vcgRzt2_1(.din(n16439), .dout(n16436));
    jdff dff_A_oqBQk2bZ4_1(.din(n16442), .dout(n16439));
    jdff dff_A_jXWACblp2_1(.din(n16445), .dout(n16442));
    jdff dff_A_I0qaYEYe2_1(.din(n16448), .dout(n16445));
    jdff dff_A_YkaaOJ3u5_1(.din(n2943), .dout(n16448));
    jdff dff_A_kmY6zEzX4_2(.din(n16454), .dout(n16451));
    jdff dff_A_YSXjvyKU1_2(.din(n16457), .dout(n16454));
    jdff dff_A_WtJarjZg2_2(.din(n16460), .dout(n16457));
    jdff dff_A_puxkd1286_2(.din(n16463), .dout(n16460));
    jdff dff_A_LBmRRY814_2(.din(n16466), .dout(n16463));
    jdff dff_A_VQwgBGOY4_2(.din(n16469), .dout(n16466));
    jdff dff_A_Dhp9Osxv4_2(.din(n16472), .dout(n16469));
    jdff dff_A_i7mXiXBc4_2(.din(n16475), .dout(n16472));
    jdff dff_A_pal6TTlv8_2(.din(n16478), .dout(n16475));
    jdff dff_A_c6gSTUhR6_2(.din(n16481), .dout(n16478));
    jdff dff_A_KgaFGU7S5_2(.din(n2943), .dout(n16481));
    jdff dff_A_UygF6HbI1_1(.din(G1694), .dout(n16484));
    jdff dff_A_T9Chpajb1_2(.din(G1691), .dout(n16487));
    jdff dff_B_7NAwkOja3_2(.din(n5380), .dout(n16491));
    jdff dff_B_RNOSPl9T2_2(.din(n16491), .dout(n16494));
    jdff dff_B_E8goaBHO6_2(.din(n16494), .dout(n16497));
    jdff dff_B_kD7A8Gu39_2(.din(n16497), .dout(n16500));
    jdff dff_B_5VSnKx8E3_2(.din(n16500), .dout(n16503));
    jdff dff_B_4MJXGFq35_2(.din(n16503), .dout(n16506));
    jdff dff_B_IgrxV5K80_2(.din(n16506), .dout(n16509));
    jdff dff_B_SQ4edi7L6_2(.din(n16509), .dout(n16512));
    jdff dff_B_XO2G3nyv7_2(.din(n16512), .dout(n16515));
    jdff dff_B_qrXm9Kl65_2(.din(n16515), .dout(n16518));
    jdff dff_B_0BJ2ic2B4_2(.din(n16518), .dout(n16521));
    jdff dff_B_W6OUSo1Y4_2(.din(n16521), .dout(n16524));
    jdff dff_B_ZCsYp7Y29_2(.din(n16524), .dout(n16527));
    jdff dff_B_myZIM1NK6_2(.din(n16527), .dout(n16530));
    jdff dff_B_vet7eIdY0_2(.din(n16530), .dout(n16533));
    jdff dff_B_xwoFjAZC4_2(.din(n16533), .dout(n16536));
    jdff dff_B_265D6Uep9_2(.din(n16536), .dout(n16539));
    jdff dff_B_ZbQa7PCp5_2(.din(n16539), .dout(n16542));
    jdff dff_B_tzjSzFk76_2(.din(n16542), .dout(n16545));
    jdff dff_B_J7FJ6BEE5_2(.din(n16545), .dout(n16548));
    jdff dff_B_FNrz4wUl8_2(.din(n16548), .dout(n16551));
    jdff dff_B_6IqE0GFm7_2(.din(n16551), .dout(n16554));
    jdff dff_B_jW1C4NRR4_2(.din(n16554), .dout(n16557));
    jdff dff_B_XDizpPKl7_2(.din(n16557), .dout(n16560));
    jdff dff_A_PxRY2uzP1_2(.din(n16565), .dout(n16562));
    jdff dff_A_RDqLBym93_2(.din(n16568), .dout(n16565));
    jdff dff_A_SsyNtHW39_2(.din(n16571), .dout(n16568));
    jdff dff_A_5fuBd4Rc0_2(.din(n16574), .dout(n16571));
    jdff dff_A_2a4lBvd87_2(.din(n16577), .dout(n16574));
    jdff dff_A_lj9TLTIy0_2(.din(n16580), .dout(n16577));
    jdff dff_A_0VuRgy847_2(.din(n16583), .dout(n16580));
    jdff dff_A_YrtCm23Q6_2(.din(n16586), .dout(n16583));
    jdff dff_A_WAFqwUEP9_2(.din(n16589), .dout(n16586));
    jdff dff_A_LD2TpBWz4_2(.din(n16592), .dout(n16589));
    jdff dff_A_k2vTd8Xu7_2(.din(n16595), .dout(n16592));
    jdff dff_A_KA52KHCR6_2(.din(n16598), .dout(n16595));
    jdff dff_A_NGxsdPAI3_2(.din(n16601), .dout(n16598));
    jdff dff_A_UaBDrsHk9_2(.din(n16604), .dout(n16601));
    jdff dff_A_Sz8mgOhv0_2(.din(n16607), .dout(n16604));
    jdff dff_A_dUYkmnTs3_2(.din(n16610), .dout(n16607));
    jdff dff_A_FGNPx9p15_2(.din(n16613), .dout(n16610));
    jdff dff_A_i4GR8iVn4_2(.din(n16616), .dout(n16613));
    jdff dff_A_DUw5Epjj0_2(.din(n16619), .dout(n16616));
    jdff dff_A_hhI9bfnN0_2(.din(n16622), .dout(n16619));
    jdff dff_A_zy1gQ3ov1_2(.din(n16625), .dout(n16622));
    jdff dff_A_Uyj3YvV44_2(.din(n16628), .dout(n16625));
    jdff dff_A_LoVGMRWh5_2(.din(G137), .dout(n16628));
    jdff dff_A_fuRUgZwW6_0(.din(n16634), .dout(n16631));
    jdff dff_A_pHqyWyMF6_0(.din(n16637), .dout(n16634));
    jdff dff_A_BA92vPRz0_0(.din(n16640), .dout(n16637));
    jdff dff_A_bhah2Hxn6_0(.din(n16643), .dout(n16640));
    jdff dff_A_sKt9M6kK5_0(.din(n16646), .dout(n16643));
    jdff dff_A_q9h7freb6_0(.din(n16649), .dout(n16646));
    jdff dff_A_e9Y3whVb1_0(.din(n16652), .dout(n16649));
    jdff dff_A_SscALKln3_0(.din(n16655), .dout(n16652));
    jdff dff_A_mv9Qe9hZ8_0(.din(n16658), .dout(n16655));
    jdff dff_A_5RacaMh79_0(.din(n16661), .dout(n16658));
    jdff dff_A_OhqbPePe9_0(.din(n16664), .dout(n16661));
    jdff dff_A_yfeF5XSX1_0(.din(n16667), .dout(n16664));
    jdff dff_A_hhoDlKC51_0(.din(n16670), .dout(n16667));
    jdff dff_A_cag0b5qf4_0(.din(n16673), .dout(n16670));
    jdff dff_A_PasI4ITh8_0(.din(n16676), .dout(n16673));
    jdff dff_A_Y7lYWyOM7_0(.din(G137), .dout(n16676));
    jdff dff_A_hyar6FWU7_1(.din(n16682), .dout(n16679));
    jdff dff_A_L5vcJehQ6_1(.din(n16685), .dout(n16682));
    jdff dff_A_OCY1RXdO1_1(.din(n16688), .dout(n16685));
    jdff dff_A_jRZYI5ML9_1(.din(n16691), .dout(n16688));
    jdff dff_A_fN4BFm7N2_1(.din(n16694), .dout(n16691));
    jdff dff_A_KRs8Gbmq9_1(.din(n16697), .dout(n16694));
    jdff dff_A_tgGPUvU04_1(.din(n16700), .dout(n16697));
    jdff dff_A_4elJ960V5_1(.din(n16703), .dout(n16700));
    jdff dff_A_SxVrNxLb4_1(.din(n16706), .dout(n16703));
    jdff dff_A_QQuo31aY2_1(.din(n16709), .dout(n16706));
    jdff dff_A_qfPzuRhQ3_1(.din(G137), .dout(n16709));
    jdff dff_A_cb5G565l2_1(.din(n5484), .dout(n16712));
    jdff dff_A_3RHCVIMc4_0(.din(n16712), .dout(n16715));
    jdff dff_A_ISAWvOxo3_0(.din(n16715), .dout(n16718));
    jdff dff_A_9Y9yy8zR4_0(.din(n16718), .dout(n16721));
    jdff dff_A_3irR0KP65_0(.din(n16721), .dout(n16724));
    jdff dff_A_JhPOMwGL6_0(.din(n16724), .dout(n16727));
    jdff dff_A_hYbRxPIL1_0(.din(n16727), .dout(n16730));
    jdff dff_A_mSDgAZtS5_0(.din(n16730), .dout(n16733));
    jdff dff_A_1nelbSrb4_0(.din(n16733), .dout(n16736));
    jdff dff_A_y309zFKo4_0(.din(n16736), .dout(n16739));
    jdff dff_A_B5kI9FwV9_0(.din(n16739), .dout(n16742));
    jdff dff_A_ny7ajQjk6_0(.din(n16742), .dout(n16745));
    jdff dff_A_AJE5QduK8_0(.din(n16745), .dout(n16748));
    jdff dff_A_t07HMYYV8_0(.din(n16748), .dout(n16751));
    jdff dff_A_Vn6bD5F74_0(.din(n16751), .dout(n16754));
    jdff dff_A_sQKv8hqb0_0(.din(n16754), .dout(n16757));
    jdff dff_A_XFJScwnh8_0(.din(n16757), .dout(n16760));
    jdff dff_A_PLWBdEet3_0(.din(n16760), .dout(n16763));
    jdff dff_A_xeKRPcYs3_0(.din(n16763), .dout(n16766));
    jdff dff_A_p16RC3072_0(.din(n16766), .dout(n16769));
    jdff dff_A_oizumvxp6_0(.din(n16769), .dout(n16772));
    jdff dff_A_0HHe19PL3_0(.din(n16772), .dout(n16775));
    jdff dff_A_AstgGGaD1_0(.din(n16775), .dout(n16778));
    jdff dff_A_pCLflLim8_0(.din(n16778), .dout(n16781));
    jdff dff_A_4HYNfnur1_0(.din(n16781), .dout(G144));
    jdff dff_A_HUppY1yx4_1(.din(n5487), .dout(n16787));
    jdff dff_A_JkxxEBys7_0(.din(n16787), .dout(n16790));
    jdff dff_A_q0n3POXW3_0(.din(n16790), .dout(n16793));
    jdff dff_A_cehktUxD0_0(.din(n16793), .dout(n16796));
    jdff dff_A_M44KfxPO4_0(.din(n16796), .dout(n16799));
    jdff dff_A_5bBBem6b8_0(.din(n16799), .dout(n16802));
    jdff dff_A_GPrB7LAM2_0(.din(n16802), .dout(n16805));
    jdff dff_A_TGBFibZw6_0(.din(n16805), .dout(n16808));
    jdff dff_A_apRmpxY45_0(.din(n16808), .dout(n16811));
    jdff dff_A_T89OFW921_0(.din(n16811), .dout(n16814));
    jdff dff_A_8yYH2IQ27_0(.din(n16814), .dout(n16817));
    jdff dff_A_R4kJCjqO1_0(.din(n16817), .dout(n16820));
    jdff dff_A_q9P3EMcU5_0(.din(n16820), .dout(n16823));
    jdff dff_A_PCp7I8GM7_0(.din(n16823), .dout(n16826));
    jdff dff_A_VsAtRIEU7_0(.din(n16826), .dout(n16829));
    jdff dff_A_hIBPr7HU2_0(.din(n16829), .dout(n16832));
    jdff dff_A_0c2WevMi6_0(.din(n16832), .dout(n16835));
    jdff dff_A_x2swy0xC4_0(.din(n16835), .dout(n16838));
    jdff dff_A_Q5s0T84Y1_0(.din(n16838), .dout(n16841));
    jdff dff_A_SZdqoSlS9_0(.din(n16841), .dout(n16844));
    jdff dff_A_Ih4eRD3R7_0(.din(n16844), .dout(n16847));
    jdff dff_A_ViwAE7JN3_0(.din(n16847), .dout(n16850));
    jdff dff_A_wIcM7nXD6_0(.din(n16850), .dout(n16853));
    jdff dff_A_gR3xRhPa6_0(.din(n16853), .dout(n16856));
    jdff dff_A_s7fIBDsj0_0(.din(n16856), .dout(G298));
    jdff dff_A_bgbfZxUg8_1(.din(n5490), .dout(n16862));
    jdff dff_A_3iukpOH64_0(.din(n16862), .dout(n16865));
    jdff dff_A_N2tLGc6e0_0(.din(n16865), .dout(n16868));
    jdff dff_A_382wXYrB6_0(.din(n16868), .dout(n16871));
    jdff dff_A_wognC2Q89_0(.din(n16871), .dout(n16874));
    jdff dff_A_DmT4I2r63_0(.din(n16874), .dout(n16877));
    jdff dff_A_AQZkrOwm2_0(.din(n16877), .dout(n16880));
    jdff dff_A_UTpaR8fz6_0(.din(n16880), .dout(n16883));
    jdff dff_A_wrgdHrHz8_0(.din(n16883), .dout(n16886));
    jdff dff_A_HdUoc6hb0_0(.din(n16886), .dout(n16889));
    jdff dff_A_Zwd2PX9a0_0(.din(n16889), .dout(n16892));
    jdff dff_A_2BwNehvp7_0(.din(n16892), .dout(n16895));
    jdff dff_A_0h2tkLmC1_0(.din(n16895), .dout(n16898));
    jdff dff_A_iXK43Zs41_0(.din(n16898), .dout(n16901));
    jdff dff_A_OmLbW4Iy4_0(.din(n16901), .dout(n16904));
    jdff dff_A_HubVTvWd0_0(.din(n16904), .dout(n16907));
    jdff dff_A_KxWanDai5_0(.din(n16907), .dout(n16910));
    jdff dff_A_hIH32iKu8_0(.din(n16910), .dout(n16913));
    jdff dff_A_4PpY3odB6_0(.din(n16913), .dout(n16916));
    jdff dff_A_qb9watoE0_0(.din(n16916), .dout(n16919));
    jdff dff_A_DDikxFB50_0(.din(n16919), .dout(n16922));
    jdff dff_A_0HXgrLo47_0(.din(n16922), .dout(n16925));
    jdff dff_A_ioyeN63Z6_0(.din(n16925), .dout(n16928));
    jdff dff_A_JN965QCk0_0(.din(n16928), .dout(n16931));
    jdff dff_A_a7Abiasf0_0(.din(n16931), .dout(G973));
    jdff dff_A_xnuHcXtR9_1(.din(n303), .dout(n16937));
    jdff dff_A_Spw7PSBT8_0(.din(n16937), .dout(n16940));
    jdff dff_A_Xd0gO3jg3_0(.din(n16940), .dout(n16943));
    jdff dff_A_dYJW6aHA3_0(.din(n16943), .dout(n16946));
    jdff dff_A_wyOinnPZ9_0(.din(n16946), .dout(n16949));
    jdff dff_A_FAJL4wXN9_0(.din(n16949), .dout(n16952));
    jdff dff_A_UqfFpiUn5_0(.din(n16952), .dout(n16955));
    jdff dff_A_waGytCvG3_0(.din(n16955), .dout(n16958));
    jdff dff_A_d59ubn9F1_0(.din(n16958), .dout(n16961));
    jdff dff_A_NaNrlEHF1_0(.din(n16961), .dout(n16964));
    jdff dff_A_seAYEsp76_0(.din(n16964), .dout(n16967));
    jdff dff_A_T1823c4M5_0(.din(n16967), .dout(n16970));
    jdff dff_A_PHux2mT88_0(.din(n16970), .dout(n16973));
    jdff dff_A_GkeuVsPt3_0(.din(n16973), .dout(n16976));
    jdff dff_A_LXypeAx94_0(.din(n16976), .dout(n16979));
    jdff dff_A_He3iXIhu0_0(.din(n16979), .dout(n16982));
    jdff dff_A_dhrAaJGI9_0(.din(n16982), .dout(n16985));
    jdff dff_A_5jo1I6l73_0(.din(n16985), .dout(n16988));
    jdff dff_A_iVV58X7c6_0(.din(n16988), .dout(n16991));
    jdff dff_A_WSa20qeo2_0(.din(n16991), .dout(n16994));
    jdff dff_A_xkFAl7Fg1_0(.din(n16994), .dout(n16997));
    jdff dff_A_9CD5bB7k9_0(.din(n16997), .dout(n17000));
    jdff dff_A_JVyna9ul2_0(.din(n17000), .dout(n17003));
    jdff dff_A_RPmdp4rG3_0(.din(n17003), .dout(n17006));
    jdff dff_A_S8O1fbJY7_0(.din(n17006), .dout(G594));
    jdff dff_A_ywNt4EiO1_1(.din(n306), .dout(n17012));
    jdff dff_A_VVNM3nxk7_0(.din(n17012), .dout(n17015));
    jdff dff_A_mmjtDoSM2_0(.din(n17015), .dout(n17018));
    jdff dff_A_b2Sh4jsb2_0(.din(n17018), .dout(n17021));
    jdff dff_A_6hYJGPOL7_0(.din(n17021), .dout(n17024));
    jdff dff_A_5umprcy05_0(.din(n17024), .dout(n17027));
    jdff dff_A_D5UXYMnK7_0(.din(n17027), .dout(n17030));
    jdff dff_A_bMwFVns33_0(.din(n17030), .dout(n17033));
    jdff dff_A_40wmxGgT3_0(.din(n17033), .dout(n17036));
    jdff dff_A_fgKMQkj48_0(.din(n17036), .dout(n17039));
    jdff dff_A_0ZQxhR5e9_0(.din(n17039), .dout(n17042));
    jdff dff_A_8dPtbYpI0_0(.din(n17042), .dout(n17045));
    jdff dff_A_Fq3HN0CL1_0(.din(n17045), .dout(n17048));
    jdff dff_A_Bd05Wsy23_0(.din(n17048), .dout(n17051));
    jdff dff_A_ALM58iN24_0(.din(n17051), .dout(n17054));
    jdff dff_A_6t3ZeJx36_0(.din(n17054), .dout(n17057));
    jdff dff_A_g3hPaqWW1_0(.din(n17057), .dout(n17060));
    jdff dff_A_vz1QgAqq4_0(.din(n17060), .dout(n17063));
    jdff dff_A_klPbOt779_0(.din(n17063), .dout(n17066));
    jdff dff_A_XQsxFS3V8_0(.din(n17066), .dout(n17069));
    jdff dff_A_iP1vrYH23_0(.din(n17069), .dout(n17072));
    jdff dff_A_koqwoAFO7_0(.din(n17072), .dout(n17075));
    jdff dff_A_LkXpchdi4_0(.din(n17075), .dout(n17078));
    jdff dff_A_IOYig3dL4_0(.din(n17078), .dout(n17081));
    jdff dff_A_RiPmO5jO7_0(.din(n17081), .dout(G599));
    jdff dff_A_wEbXZwDn0_1(.din(n309), .dout(n17087));
    jdff dff_A_HSvLcFhP5_0(.din(n17087), .dout(n17090));
    jdff dff_A_BCZSTrqm4_0(.din(n17090), .dout(n17093));
    jdff dff_A_311DW8Cb4_0(.din(n17093), .dout(n17096));
    jdff dff_A_EM8T03Ww0_0(.din(n17096), .dout(n17099));
    jdff dff_A_7mfxGjPM5_0(.din(n17099), .dout(n17102));
    jdff dff_A_yGoa4VFG3_0(.din(n17102), .dout(n17105));
    jdff dff_A_BCLyTzPz5_0(.din(n17105), .dout(n17108));
    jdff dff_A_dSxoOqCP5_0(.din(n17108), .dout(n17111));
    jdff dff_A_AaFa3NAg8_0(.din(n17111), .dout(n17114));
    jdff dff_A_onjYlMBl9_0(.din(n17114), .dout(n17117));
    jdff dff_A_XfTgz1Vg6_0(.din(n17117), .dout(n17120));
    jdff dff_A_JncHxJWa5_0(.din(n17120), .dout(n17123));
    jdff dff_A_1g6dkrv70_0(.din(n17123), .dout(n17126));
    jdff dff_A_Yvh6AOlh0_0(.din(n17126), .dout(n17129));
    jdff dff_A_aSNyovvN8_0(.din(n17129), .dout(n17132));
    jdff dff_A_Ev5iRoSw1_0(.din(n17132), .dout(n17135));
    jdff dff_A_ENUbs8W56_0(.din(n17135), .dout(n17138));
    jdff dff_A_Wuoudu227_0(.din(n17138), .dout(n17141));
    jdff dff_A_rJulTKrw4_0(.din(n17141), .dout(n17144));
    jdff dff_A_gOIlfFh00_0(.din(n17144), .dout(n17147));
    jdff dff_A_NwZT58qA1_0(.din(n17147), .dout(n17150));
    jdff dff_A_shR6BZ6X7_0(.din(n17150), .dout(n17153));
    jdff dff_A_YY9zUnjr2_0(.din(n17153), .dout(n17156));
    jdff dff_A_jrqvbr3c8_0(.din(n17156), .dout(G600));
    jdff dff_A_XBKdFEY12_1(.din(n313), .dout(n17162));
    jdff dff_A_W3blJKaT6_0(.din(n17162), .dout(n17165));
    jdff dff_A_m5lxHlBy9_0(.din(n17165), .dout(n17168));
    jdff dff_A_hDxQ0zxn9_0(.din(n17168), .dout(n17171));
    jdff dff_A_Hlx88qOv2_0(.din(n17171), .dout(n17174));
    jdff dff_A_SRZmYHN44_0(.din(n17174), .dout(n17177));
    jdff dff_A_j8WvfXCf3_0(.din(n17177), .dout(n17180));
    jdff dff_A_hGPvJOyA4_0(.din(n17180), .dout(n17183));
    jdff dff_A_1CGvhTYl6_0(.din(n17183), .dout(n17186));
    jdff dff_A_y4T2JSsi1_0(.din(n17186), .dout(n17189));
    jdff dff_A_ghNw8vfW5_0(.din(n17189), .dout(n17192));
    jdff dff_A_lQLqOei06_0(.din(n17192), .dout(n17195));
    jdff dff_A_3un9PmG75_0(.din(n17195), .dout(n17198));
    jdff dff_A_U8ZpNnbz5_0(.din(n17198), .dout(n17201));
    jdff dff_A_CQI7aj3O9_0(.din(n17201), .dout(n17204));
    jdff dff_A_PymAOf9O4_0(.din(n17204), .dout(n17207));
    jdff dff_A_WFBKwnf95_0(.din(n17207), .dout(n17210));
    jdff dff_A_bUgXr9FK0_0(.din(n17210), .dout(n17213));
    jdff dff_A_5ga8yakY1_0(.din(n17213), .dout(n17216));
    jdff dff_A_jyezGBJM0_0(.din(n17216), .dout(n17219));
    jdff dff_A_ADE6YPIK2_0(.din(n17219), .dout(n17222));
    jdff dff_A_ZMSHaKc78_0(.din(n17222), .dout(n17225));
    jdff dff_A_StMOIgqG7_0(.din(n17225), .dout(n17228));
    jdff dff_A_VVPO2BMh9_0(.din(n17228), .dout(n17231));
    jdff dff_A_oe8Go6Nb7_0(.din(n17231), .dout(G601));
    jdff dff_A_5UiApBuf0_1(.din(n316), .dout(n17237));
    jdff dff_A_ZOfNn9lZ0_0(.din(n17237), .dout(n17240));
    jdff dff_A_pCIAjKVy3_0(.din(n17240), .dout(n17243));
    jdff dff_A_lfRHEVvT8_0(.din(n17243), .dout(n17246));
    jdff dff_A_CCsFULqC1_0(.din(n17246), .dout(n17249));
    jdff dff_A_q26Ia2Vz8_0(.din(n17249), .dout(n17252));
    jdff dff_A_txdgd2aV0_0(.din(n17252), .dout(n17255));
    jdff dff_A_Tqyn0PGs2_0(.din(n17255), .dout(n17258));
    jdff dff_A_PupEY9tU4_0(.din(n17258), .dout(n17261));
    jdff dff_A_GulXQyOr1_0(.din(n17261), .dout(n17264));
    jdff dff_A_VwJ7xpip8_0(.din(n17264), .dout(n17267));
    jdff dff_A_JiNepxSR2_0(.din(n17267), .dout(n17270));
    jdff dff_A_fdfoUjCQ8_0(.din(n17270), .dout(n17273));
    jdff dff_A_evjQ1GOQ6_0(.din(n17273), .dout(n17276));
    jdff dff_A_Ai2LZgHB2_0(.din(n17276), .dout(n17279));
    jdff dff_A_qkThCd3n6_0(.din(n17279), .dout(n17282));
    jdff dff_A_wP7OkQIs7_0(.din(n17282), .dout(n17285));
    jdff dff_A_0gh7OFPG4_0(.din(n17285), .dout(n17288));
    jdff dff_A_Bc87HXuD6_0(.din(n17288), .dout(n17291));
    jdff dff_A_IXJSGref9_0(.din(n17291), .dout(n17294));
    jdff dff_A_3RJ4Z2zp8_0(.din(n17294), .dout(n17297));
    jdff dff_A_nZsYqJsJ8_0(.din(n17297), .dout(n17300));
    jdff dff_A_jmvhyzkZ3_0(.din(n17300), .dout(n17303));
    jdff dff_A_TZvXZ9uQ0_0(.din(n17303), .dout(n17306));
    jdff dff_A_uHLArAq26_0(.din(n17306), .dout(G602));
    jdff dff_A_lAjJ6ntN2_1(.din(n5493), .dout(n17312));
    jdff dff_A_gX4l8LdO0_0(.din(n17312), .dout(n17315));
    jdff dff_A_Ez6ANdeV7_0(.din(n17315), .dout(n17318));
    jdff dff_A_0KZsZlnI4_0(.din(n17318), .dout(n17321));
    jdff dff_A_dLJb00FY5_0(.din(n17321), .dout(n17324));
    jdff dff_A_UJcq1LMn1_0(.din(n17324), .dout(n17327));
    jdff dff_A_lD83Iwof9_0(.din(n17327), .dout(n17330));
    jdff dff_A_Nx1kym4p3_0(.din(n17330), .dout(n17333));
    jdff dff_A_QavivzIi6_0(.din(n17333), .dout(n17336));
    jdff dff_A_2t2VTaDi9_0(.din(n17336), .dout(n17339));
    jdff dff_A_CDtK9NDC3_0(.din(n17339), .dout(n17342));
    jdff dff_A_MJ9UoudK5_0(.din(n17342), .dout(n17345));
    jdff dff_A_btQjM91A6_0(.din(n17345), .dout(n17348));
    jdff dff_A_ncjZG1842_0(.din(n17348), .dout(n17351));
    jdff dff_A_BTtIqM3W0_0(.din(n17351), .dout(n17354));
    jdff dff_A_YPsrmVI95_0(.din(n17354), .dout(n17357));
    jdff dff_A_efGUEy068_0(.din(n17357), .dout(n17360));
    jdff dff_A_XMI3Hs1t2_0(.din(n17360), .dout(n17363));
    jdff dff_A_43dXQUqv6_0(.din(n17363), .dout(n17366));
    jdff dff_A_c6UIM3pj6_0(.din(n17366), .dout(n17369));
    jdff dff_A_t6VnbjB46_0(.din(n17369), .dout(n17372));
    jdff dff_A_saPPbtAo1_0(.din(n17372), .dout(n17375));
    jdff dff_A_woxLorAt1_0(.din(n17375), .dout(n17378));
    jdff dff_A_xC83BlN51_0(.din(n17378), .dout(n17381));
    jdff dff_A_yFnvOrBl4_0(.din(n17381), .dout(G603));
    jdff dff_A_0HHr3PS48_1(.din(n5496), .dout(n17387));
    jdff dff_A_Qmt1iINc8_0(.din(n17387), .dout(n17390));
    jdff dff_A_aEUtmnu55_0(.din(n17390), .dout(n17393));
    jdff dff_A_68hFG8kh9_0(.din(n17393), .dout(n17396));
    jdff dff_A_i1ZtKfQ55_0(.din(n17396), .dout(n17399));
    jdff dff_A_02bHml4r6_0(.din(n17399), .dout(n17402));
    jdff dff_A_1D89T5S51_0(.din(n17402), .dout(n17405));
    jdff dff_A_1eccpagy6_0(.din(n17405), .dout(n17408));
    jdff dff_A_69nOebat5_0(.din(n17408), .dout(n17411));
    jdff dff_A_NrxZeAKF7_0(.din(n17411), .dout(n17414));
    jdff dff_A_DhUKxEso9_0(.din(n17414), .dout(n17417));
    jdff dff_A_IhPRGPGP1_0(.din(n17417), .dout(n17420));
    jdff dff_A_RqErZqyq3_0(.din(n17420), .dout(n17423));
    jdff dff_A_mvELn8jo3_0(.din(n17423), .dout(n17426));
    jdff dff_A_XLzwTO640_0(.din(n17426), .dout(n17429));
    jdff dff_A_WbG5VX9j6_0(.din(n17429), .dout(n17432));
    jdff dff_A_PcQC7G1V9_0(.din(n17432), .dout(n17435));
    jdff dff_A_yXkrA4Gj0_0(.din(n17435), .dout(n17438));
    jdff dff_A_lg24CHzt4_0(.din(n17438), .dout(n17441));
    jdff dff_A_U4yiVyUN6_0(.din(n17441), .dout(n17444));
    jdff dff_A_IuxKDhvs7_0(.din(n17444), .dout(n17447));
    jdff dff_A_uJSbDNmw2_0(.din(n17447), .dout(n17450));
    jdff dff_A_9D16R5mB7_0(.din(n17450), .dout(n17453));
    jdff dff_A_nqZkEy4U6_0(.din(n17453), .dout(n17456));
    jdff dff_A_ALW4vH0j8_0(.din(n17456), .dout(G604));
    jdff dff_A_pVw4klAf8_1(.din(n319), .dout(n17462));
    jdff dff_A_QLZW3LF36_0(.din(n17462), .dout(n17465));
    jdff dff_A_U6fvBceE8_0(.din(n17465), .dout(n17468));
    jdff dff_A_j2UNdXJB2_0(.din(n17468), .dout(n17471));
    jdff dff_A_mhqfB2Nq4_0(.din(n17471), .dout(n17474));
    jdff dff_A_lvme9Jct0_0(.din(n17474), .dout(n17477));
    jdff dff_A_jJFicvkV8_0(.din(n17477), .dout(n17480));
    jdff dff_A_6YMLwFrZ2_0(.din(n17480), .dout(n17483));
    jdff dff_A_ja7oAzQ41_0(.din(n17483), .dout(n17486));
    jdff dff_A_nGvgUjE06_0(.din(n17486), .dout(n17489));
    jdff dff_A_24EAdmNA6_0(.din(n17489), .dout(n17492));
    jdff dff_A_GZdqD08q0_0(.din(n17492), .dout(n17495));
    jdff dff_A_4VY4z9Pt4_0(.din(n17495), .dout(n17498));
    jdff dff_A_il4hTyVm3_0(.din(n17498), .dout(n17501));
    jdff dff_A_ZEhDEe0d7_0(.din(n17501), .dout(n17504));
    jdff dff_A_RST6M91K4_0(.din(n17504), .dout(n17507));
    jdff dff_A_NxDDcVaf2_0(.din(n17507), .dout(n17510));
    jdff dff_A_dvmq6JXW8_0(.din(n17510), .dout(n17513));
    jdff dff_A_NQkEYQCw9_0(.din(n17513), .dout(n17516));
    jdff dff_A_BKhPLSCs0_0(.din(n17516), .dout(n17519));
    jdff dff_A_JPzGiUwV2_0(.din(n17519), .dout(n17522));
    jdff dff_A_l2wvO4NR9_0(.din(n17522), .dout(n17525));
    jdff dff_A_W2E9JpJS4_0(.din(n17525), .dout(n17528));
    jdff dff_A_YI2X50pv5_0(.din(n17528), .dout(n17531));
    jdff dff_A_XqTn1v4h0_0(.din(n17531), .dout(G611));
    jdff dff_A_Kl1VYOge1_1(.din(n322), .dout(n17537));
    jdff dff_A_B3EwKRTa9_0(.din(n17537), .dout(n17540));
    jdff dff_A_rbVVryLn6_0(.din(n17540), .dout(n17543));
    jdff dff_A_c6k24Z1B1_0(.din(n17543), .dout(n17546));
    jdff dff_A_2SynLc0q1_0(.din(n17546), .dout(n17549));
    jdff dff_A_O3rLhcNa3_0(.din(n17549), .dout(n17552));
    jdff dff_A_YFCZmZn02_0(.din(n17552), .dout(n17555));
    jdff dff_A_DE6c4i8X6_0(.din(n17555), .dout(n17558));
    jdff dff_A_NeIydeCE1_0(.din(n17558), .dout(n17561));
    jdff dff_A_2Gutarxx1_0(.din(n17561), .dout(n17564));
    jdff dff_A_NuPQ2fAM5_0(.din(n17564), .dout(n17567));
    jdff dff_A_GwN5urio6_0(.din(n17567), .dout(n17570));
    jdff dff_A_k0m57NFn4_0(.din(n17570), .dout(n17573));
    jdff dff_A_MRZmuARF4_0(.din(n17573), .dout(n17576));
    jdff dff_A_veRZFaGf5_0(.din(n17576), .dout(n17579));
    jdff dff_A_EXIBH7FF2_0(.din(n17579), .dout(n17582));
    jdff dff_A_AtIWkV7A8_0(.din(n17582), .dout(n17585));
    jdff dff_A_TFfMWMZO1_0(.din(n17585), .dout(n17588));
    jdff dff_A_iLXbjr3R9_0(.din(n17588), .dout(n17591));
    jdff dff_A_d4aptmOa9_0(.din(n17591), .dout(n17594));
    jdff dff_A_q2MZOYAs3_0(.din(n17594), .dout(n17597));
    jdff dff_A_KMZPdXSE5_0(.din(n17597), .dout(n17600));
    jdff dff_A_BbSM9Wij0_0(.din(n17600), .dout(n17603));
    jdff dff_A_hlhQvUvX2_0(.din(n17603), .dout(n17606));
    jdff dff_A_6NRR88zZ4_0(.din(n17606), .dout(G612));
    jdff dff_A_xWfJIjhY9_2(.din(n326), .dout(n17612));
    jdff dff_A_W4QEECt23_0(.din(n17612), .dout(n17615));
    jdff dff_A_MXJCNFNP1_0(.din(n17615), .dout(n17618));
    jdff dff_A_cSP4Twnl9_0(.din(n17618), .dout(n17621));
    jdff dff_A_iXMe5Czr1_0(.din(n17621), .dout(n17624));
    jdff dff_A_xFIVFouJ1_0(.din(n17624), .dout(n17627));
    jdff dff_A_0gMiaVB54_0(.din(n17627), .dout(n17630));
    jdff dff_A_9jo7rlqd1_0(.din(n17630), .dout(n17633));
    jdff dff_A_3JCQ8Gq22_0(.din(n17633), .dout(n17636));
    jdff dff_A_Ax7jbXJF4_0(.din(n17636), .dout(n17639));
    jdff dff_A_nFmYb7tG1_0(.din(n17639), .dout(n17642));
    jdff dff_A_6VGXosrO9_0(.din(n17642), .dout(n17645));
    jdff dff_A_R0wUTnBv8_0(.din(n17645), .dout(n17648));
    jdff dff_A_qw6D6rlu2_0(.din(n17648), .dout(n17651));
    jdff dff_A_OioMYsVH6_0(.din(n17651), .dout(n17654));
    jdff dff_A_Pfcmgsu95_0(.din(n17654), .dout(n17657));
    jdff dff_A_i8mtKWq51_0(.din(n17657), .dout(n17660));
    jdff dff_A_IsSgKvSD1_0(.din(n17660), .dout(n17663));
    jdff dff_A_uzhGcz4w8_0(.din(n17663), .dout(n17666));
    jdff dff_A_HsMeHz2e6_0(.din(n17666), .dout(n17669));
    jdff dff_A_n5iaUi1I4_0(.din(n17669), .dout(n17672));
    jdff dff_A_TXXm7fNr1_0(.din(n17672), .dout(n17675));
    jdff dff_A_r6nBd33b4_0(.din(n17675), .dout(n17678));
    jdff dff_A_7eHj7Vmb0_0(.din(n17678), .dout(n17681));
    jdff dff_A_aMOluZcQ8_0(.din(n17681), .dout(G810));
    jdff dff_A_DKH03zRr9_1(.din(n329), .dout(n17687));
    jdff dff_A_V9Dl4hlm9_0(.din(n17687), .dout(n17690));
    jdff dff_A_ZevjiADK7_0(.din(n17690), .dout(n17693));
    jdff dff_A_YH5oIzoM3_0(.din(n17693), .dout(n17696));
    jdff dff_A_TYuXSnAM2_0(.din(n17696), .dout(n17699));
    jdff dff_A_ubolZQDz4_0(.din(n17699), .dout(n17702));
    jdff dff_A_J1c3ZeLx1_0(.din(n17702), .dout(n17705));
    jdff dff_A_OCHDOgu56_0(.din(n17705), .dout(n17708));
    jdff dff_A_wU3Gi6uw6_0(.din(n17708), .dout(n17711));
    jdff dff_A_5z0GlFRk3_0(.din(n17711), .dout(n17714));
    jdff dff_A_ISNGNLqq6_0(.din(n17714), .dout(n17717));
    jdff dff_A_itNXrn802_0(.din(n17717), .dout(n17720));
    jdff dff_A_Cjtrg6io1_0(.din(n17720), .dout(n17723));
    jdff dff_A_xtaWXGfw8_0(.din(n17723), .dout(n17726));
    jdff dff_A_SugRY9d51_0(.din(n17726), .dout(n17729));
    jdff dff_A_fXetze8D1_0(.din(n17729), .dout(n17732));
    jdff dff_A_PoTC19mg5_0(.din(n17732), .dout(n17735));
    jdff dff_A_dOIkIvFI4_0(.din(n17735), .dout(n17738));
    jdff dff_A_qYYjo8Di4_0(.din(n17738), .dout(n17741));
    jdff dff_A_50UqEfcW1_0(.din(n17741), .dout(n17744));
    jdff dff_A_enR1XClG3_0(.din(n17744), .dout(n17747));
    jdff dff_A_9S2mwn7J5_0(.din(n17747), .dout(n17750));
    jdff dff_A_RpaTGwKC1_0(.din(n17750), .dout(n17753));
    jdff dff_A_lo72eVtF8_0(.din(n17753), .dout(n17756));
    jdff dff_A_0TcMbMkW1_0(.din(n17756), .dout(G848));
    jdff dff_A_C4E6I9xm8_1(.din(n332), .dout(n17762));
    jdff dff_A_J3wecKfl8_0(.din(n17762), .dout(n17765));
    jdff dff_A_PVdshIEX2_0(.din(n17765), .dout(n17768));
    jdff dff_A_9tqw22TR0_0(.din(n17768), .dout(n17771));
    jdff dff_A_o3O10GqH6_0(.din(n17771), .dout(n17774));
    jdff dff_A_VKsIspZl5_0(.din(n17774), .dout(n17777));
    jdff dff_A_w7nMf7iq6_0(.din(n17777), .dout(n17780));
    jdff dff_A_gD03OdNp1_0(.din(n17780), .dout(n17783));
    jdff dff_A_pWObaypn4_0(.din(n17783), .dout(n17786));
    jdff dff_A_JhTP2HUO8_0(.din(n17786), .dout(n17789));
    jdff dff_A_vNHZzIe48_0(.din(n17789), .dout(n17792));
    jdff dff_A_LcUEyZrV4_0(.din(n17792), .dout(n17795));
    jdff dff_A_tb1jacsR7_0(.din(n17795), .dout(n17798));
    jdff dff_A_KIy3WwXd8_0(.din(n17798), .dout(n17801));
    jdff dff_A_K1ZQVDtw3_0(.din(n17801), .dout(n17804));
    jdff dff_A_JprNTZPk2_0(.din(n17804), .dout(n17807));
    jdff dff_A_QObp4Vzv6_0(.din(n17807), .dout(n17810));
    jdff dff_A_uFxb5Z0a8_0(.din(n17810), .dout(n17813));
    jdff dff_A_mfr59jnh5_0(.din(n17813), .dout(n17816));
    jdff dff_A_hmAAue0G0_0(.din(n17816), .dout(n17819));
    jdff dff_A_KhmX7SqM9_0(.din(n17819), .dout(n17822));
    jdff dff_A_82TbgnjM3_0(.din(n17822), .dout(n17825));
    jdff dff_A_qur3YhbT2_0(.din(n17825), .dout(n17828));
    jdff dff_A_PgAh9jYo8_0(.din(n17828), .dout(n17831));
    jdff dff_A_vJqoAf853_0(.din(n17831), .dout(G849));
    jdff dff_A_IneqafsU3_1(.din(n335), .dout(n17837));
    jdff dff_A_bdp2HV5j4_0(.din(n17837), .dout(n17840));
    jdff dff_A_ZMxhpMte3_0(.din(n17840), .dout(n17843));
    jdff dff_A_T24lEb8t1_0(.din(n17843), .dout(n17846));
    jdff dff_A_zDmCoZu30_0(.din(n17846), .dout(n17849));
    jdff dff_A_woHPVkCV7_0(.din(n17849), .dout(n17852));
    jdff dff_A_s6T66enI5_0(.din(n17852), .dout(n17855));
    jdff dff_A_60S9acg72_0(.din(n17855), .dout(n17858));
    jdff dff_A_IsYTu06N0_0(.din(n17858), .dout(n17861));
    jdff dff_A_CDoPbfqB5_0(.din(n17861), .dout(n17864));
    jdff dff_A_wB8aa1u45_0(.din(n17864), .dout(n17867));
    jdff dff_A_SpKjj8Rh2_0(.din(n17867), .dout(n17870));
    jdff dff_A_FiJF7Unv8_0(.din(n17870), .dout(n17873));
    jdff dff_A_PUkP4kX68_0(.din(n17873), .dout(n17876));
    jdff dff_A_HpCYed7l8_0(.din(n17876), .dout(n17879));
    jdff dff_A_HP3KpLfy3_0(.din(n17879), .dout(n17882));
    jdff dff_A_utArNpwp5_0(.din(n17882), .dout(n17885));
    jdff dff_A_nn2F6oWB8_0(.din(n17885), .dout(n17888));
    jdff dff_A_wFixckNx2_0(.din(n17888), .dout(n17891));
    jdff dff_A_DcnDZqoU9_0(.din(n17891), .dout(n17894));
    jdff dff_A_fnWcAW433_0(.din(n17894), .dout(n17897));
    jdff dff_A_j6BIrdjI5_0(.din(n17897), .dout(n17900));
    jdff dff_A_zF1ysYqI0_0(.din(n17900), .dout(n17903));
    jdff dff_A_JSZIW3jV1_0(.din(n17903), .dout(n17906));
    jdff dff_A_kfRy5ahu9_0(.din(n17906), .dout(G850));
    jdff dff_A_1xSfMYMt0_1(.din(n338), .dout(n17912));
    jdff dff_A_9LKRB3f68_0(.din(n17912), .dout(n17915));
    jdff dff_A_gc0i5aTx3_0(.din(n17915), .dout(n17918));
    jdff dff_A_ZnFsmU7S4_0(.din(n17918), .dout(n17921));
    jdff dff_A_LXhdFnde2_0(.din(n17921), .dout(n17924));
    jdff dff_A_OK9feKSz0_0(.din(n17924), .dout(n17927));
    jdff dff_A_teOyDpbz2_0(.din(n17927), .dout(n17930));
    jdff dff_A_P1SAHPB60_0(.din(n17930), .dout(n17933));
    jdff dff_A_agHq9Vxe8_0(.din(n17933), .dout(n17936));
    jdff dff_A_W6mCaI3z2_0(.din(n17936), .dout(n17939));
    jdff dff_A_8vAThO435_0(.din(n17939), .dout(n17942));
    jdff dff_A_eP8CBvWY0_0(.din(n17942), .dout(n17945));
    jdff dff_A_lJPviwf89_0(.din(n17945), .dout(n17948));
    jdff dff_A_KQClxOC20_0(.din(n17948), .dout(n17951));
    jdff dff_A_xYtiwiq53_0(.din(n17951), .dout(n17954));
    jdff dff_A_jROIc4bY6_0(.din(n17954), .dout(n17957));
    jdff dff_A_V1qaUMme6_0(.din(n17957), .dout(n17960));
    jdff dff_A_jAtJSnBV4_0(.din(n17960), .dout(n17963));
    jdff dff_A_Q4j7EZNm1_0(.din(n17963), .dout(n17966));
    jdff dff_A_dGN7hzBT7_0(.din(n17966), .dout(n17969));
    jdff dff_A_hR5xHatP1_0(.din(n17969), .dout(n17972));
    jdff dff_A_FszJodIF2_0(.din(n17972), .dout(n17975));
    jdff dff_A_mAvnTKmL2_0(.din(n17975), .dout(n17978));
    jdff dff_A_S6IQxkHY2_0(.din(n17978), .dout(n17981));
    jdff dff_A_aqqtuCRt9_0(.din(n17981), .dout(G851));
    jdff dff_A_ZCfZqptZ2_2(.din(n342), .dout(n17987));
    jdff dff_A_AkxK3PXr7_0(.din(n17987), .dout(n17990));
    jdff dff_A_j94OQCS04_0(.din(n17990), .dout(n17993));
    jdff dff_A_cQBw3GLb0_0(.din(n17993), .dout(n17996));
    jdff dff_A_ysenTGml1_0(.din(n17996), .dout(n17999));
    jdff dff_A_AxYT9JZM0_0(.din(n17999), .dout(n18002));
    jdff dff_A_hKYqQDsu7_0(.din(n18002), .dout(n18005));
    jdff dff_A_1r1Xn5aR6_0(.din(n18005), .dout(n18008));
    jdff dff_A_q78m1Ni15_0(.din(n18008), .dout(n18011));
    jdff dff_A_FOJ9xqi72_0(.din(n18011), .dout(n18014));
    jdff dff_A_oWZFgUY55_0(.din(n18014), .dout(n18017));
    jdff dff_A_Zct95VyD4_0(.din(n18017), .dout(n18020));
    jdff dff_A_Yl725GGn9_0(.din(n18020), .dout(n18023));
    jdff dff_A_4vRX5qte9_0(.din(n18023), .dout(n18026));
    jdff dff_A_TzdtOuMs7_0(.din(n18026), .dout(n18029));
    jdff dff_A_ZsjCNNIt6_0(.din(n18029), .dout(n18032));
    jdff dff_A_sNtzgHPm3_0(.din(n18032), .dout(n18035));
    jdff dff_A_W3L6Sddn7_0(.din(n18035), .dout(n18038));
    jdff dff_A_UAHvOLWt6_0(.din(n18038), .dout(n18041));
    jdff dff_A_J7uiRwTk6_0(.din(n18041), .dout(n18044));
    jdff dff_A_l6pT0S5f5_0(.din(n18044), .dout(n18047));
    jdff dff_A_yXpblTTG0_0(.din(n18047), .dout(n18050));
    jdff dff_A_uS9K5RRB1_0(.din(n18050), .dout(n18053));
    jdff dff_A_Xtw3kVUu5_0(.din(n18053), .dout(n18056));
    jdff dff_A_dlMMGcj04_0(.din(n18056), .dout(G634));
    jdff dff_A_85EWI87F1_2(.din(n349), .dout(n18062));
    jdff dff_A_wUlp3ZHb7_0(.din(n18062), .dout(n18065));
    jdff dff_A_CtFMHTU65_0(.din(n18065), .dout(n18068));
    jdff dff_A_VRHQM1D97_0(.din(n18068), .dout(n18071));
    jdff dff_A_vuJDotK36_0(.din(n18071), .dout(n18074));
    jdff dff_A_smtJ0N6p1_0(.din(n18074), .dout(n18077));
    jdff dff_A_nVzTU1wv0_0(.din(n18077), .dout(n18080));
    jdff dff_A_vgYyKTxe5_0(.din(n18080), .dout(n18083));
    jdff dff_A_CbaKDPNt4_0(.din(n18083), .dout(n18086));
    jdff dff_A_NJXZjmGw5_0(.din(n18086), .dout(n18089));
    jdff dff_A_U8hkgIES8_0(.din(n18089), .dout(n18092));
    jdff dff_A_aCh7I36M3_0(.din(n18092), .dout(n18095));
    jdff dff_A_gVs8XcDN0_0(.din(n18095), .dout(n18098));
    jdff dff_A_zkZJzAKK1_0(.din(n18098), .dout(n18101));
    jdff dff_A_2EEfBfON7_0(.din(n18101), .dout(n18104));
    jdff dff_A_m8vJpnEV2_0(.din(n18104), .dout(n18107));
    jdff dff_A_uUKXjEl93_0(.din(n18107), .dout(n18110));
    jdff dff_A_RAsSNRWz7_0(.din(n18110), .dout(n18113));
    jdff dff_A_NTzsG20u9_0(.din(n18113), .dout(n18116));
    jdff dff_A_H8wcQRyh4_0(.din(n18116), .dout(n18119));
    jdff dff_A_L6kVtjQ69_0(.din(n18119), .dout(n18122));
    jdff dff_A_RRt0yPzE5_0(.din(n18122), .dout(n18125));
    jdff dff_A_7o8UcTC54_0(.din(n18125), .dout(n18128));
    jdff dff_A_0ncU4kYV4_0(.din(n18128), .dout(G815));
    jdff dff_A_wbIT1XPG9_2(.din(n356), .dout(n18134));
    jdff dff_A_vgwIbBju5_0(.din(n18134), .dout(n18137));
    jdff dff_A_bkFvrZ5J3_0(.din(n18137), .dout(n18140));
    jdff dff_A_xRcw8JG86_0(.din(n18140), .dout(n18143));
    jdff dff_A_kbBSzTe02_0(.din(n18143), .dout(n18146));
    jdff dff_A_7bH0luB35_0(.din(n18146), .dout(n18149));
    jdff dff_A_zHxniMfJ0_0(.din(n18149), .dout(n18152));
    jdff dff_A_GXJk6YgY3_0(.din(n18152), .dout(n18155));
    jdff dff_A_DklyxYxz6_0(.din(n18155), .dout(n18158));
    jdff dff_A_5J3lHr7j0_0(.din(n18158), .dout(n18161));
    jdff dff_A_gkAYmFWb4_0(.din(n18161), .dout(n18164));
    jdff dff_A_Z9izDOnl8_0(.din(n18164), .dout(n18167));
    jdff dff_A_2UoyOGkc1_0(.din(n18167), .dout(n18170));
    jdff dff_A_besySP5H1_0(.din(n18170), .dout(n18173));
    jdff dff_A_T1cYBKAv7_0(.din(n18173), .dout(n18176));
    jdff dff_A_DWjNw2ar2_0(.din(n18176), .dout(n18179));
    jdff dff_A_yiRhqAu64_0(.din(n18179), .dout(n18182));
    jdff dff_A_3s9vnMc08_0(.din(n18182), .dout(n18185));
    jdff dff_A_1XzhlFWJ2_0(.din(n18185), .dout(n18188));
    jdff dff_A_wSKLq0gu0_0(.din(n18188), .dout(n18191));
    jdff dff_A_BCZp0mBa3_0(.din(n18191), .dout(n18194));
    jdff dff_A_uApHQBbg7_0(.din(n18194), .dout(n18197));
    jdff dff_A_es2KX2yR9_0(.din(n18197), .dout(n18200));
    jdff dff_A_frJMrqSo1_0(.din(n18200), .dout(G845));
    jdff dff_A_baaaIop22_1(.din(n363), .dout(n18206));
    jdff dff_A_qHT3LPmz5_0(.din(n18206), .dout(n18209));
    jdff dff_A_zMglTbSo5_0(.din(n18209), .dout(n18212));
    jdff dff_A_h9dnR1xR0_0(.din(n18212), .dout(n18215));
    jdff dff_A_Wb0DyuPT7_0(.din(n18215), .dout(n18218));
    jdff dff_A_rn7xnLiI9_0(.din(n18218), .dout(n18221));
    jdff dff_A_gpoeS98b4_0(.din(n18221), .dout(n18224));
    jdff dff_A_cJHceGsL9_0(.din(n18224), .dout(n18227));
    jdff dff_A_u3soHglQ8_0(.din(n18227), .dout(n18230));
    jdff dff_A_XrlUDqrv8_0(.din(n18230), .dout(n18233));
    jdff dff_A_3yjouAZG0_0(.din(n18233), .dout(n18236));
    jdff dff_A_jwnGBlz66_0(.din(n18236), .dout(n18239));
    jdff dff_A_NqnhHSnG4_0(.din(n18239), .dout(n18242));
    jdff dff_A_ZzH1PtJZ5_0(.din(n18242), .dout(n18245));
    jdff dff_A_x7LHgaJv8_0(.din(n18245), .dout(n18248));
    jdff dff_A_VZvGSK4Y3_0(.din(n18248), .dout(n18251));
    jdff dff_A_TYHC74x96_0(.din(n18251), .dout(n18254));
    jdff dff_A_23nFjEDI6_0(.din(n18254), .dout(n18257));
    jdff dff_A_ET4TfNhs6_0(.din(n18257), .dout(n18260));
    jdff dff_A_yMhm8xQV2_0(.din(n18260), .dout(n18263));
    jdff dff_A_Pco2ROqo6_0(.din(n18263), .dout(n18266));
    jdff dff_A_pv6D1KCd8_0(.din(n18266), .dout(n18269));
    jdff dff_A_WHxedDe84_0(.din(n18269), .dout(n18272));
    jdff dff_A_Q52y1VST8_0(.din(n18272), .dout(G847));
    jdff dff_A_0NtsHe4k0_1(.din(n5499), .dout(n18278));
    jdff dff_A_z8SEhmuw8_0(.din(n18278), .dout(n18281));
    jdff dff_A_0JW3qpPK1_0(.din(n18281), .dout(n18284));
    jdff dff_A_uZQRpj9u4_0(.din(n18284), .dout(n18287));
    jdff dff_A_UOWIhbIO6_0(.din(n18287), .dout(n18290));
    jdff dff_A_fcI1VUiZ9_0(.din(n18290), .dout(n18293));
    jdff dff_A_BWbThhkX9_0(.din(n18293), .dout(n18296));
    jdff dff_A_4qtfWl6m2_0(.din(n18296), .dout(n18299));
    jdff dff_A_UIUiWn8S4_0(.din(n18299), .dout(n18302));
    jdff dff_A_fvWGtN4H3_0(.din(n18302), .dout(n18305));
    jdff dff_A_VgWcOzhL8_0(.din(n18305), .dout(n18308));
    jdff dff_A_8VCmIRiZ1_0(.din(n18308), .dout(n18311));
    jdff dff_A_aiG5mRhr7_0(.din(n18311), .dout(n18314));
    jdff dff_A_rnff7rdv9_0(.din(n18314), .dout(n18317));
    jdff dff_A_C5fA222u1_0(.din(n18317), .dout(n18320));
    jdff dff_A_in6rFIyp5_0(.din(n18320), .dout(n18323));
    jdff dff_A_xHmOpUZn8_0(.din(n18323), .dout(n18326));
    jdff dff_A_ZO8cscaM6_0(.din(n18326), .dout(n18329));
    jdff dff_A_N8nSplsF6_0(.din(n18329), .dout(n18332));
    jdff dff_A_22FwJYlc0_0(.din(n18332), .dout(n18335));
    jdff dff_A_xbtWDrRh7_0(.din(n18335), .dout(n18338));
    jdff dff_A_JzC9FgC18_0(.din(n18338), .dout(n18341));
    jdff dff_A_DhTOD46w3_0(.din(n18341), .dout(n18344));
    jdff dff_A_0lLBpF6k3_0(.din(n18344), .dout(n18347));
    jdff dff_A_910Pao2f1_0(.din(n18347), .dout(G926));
    jdff dff_A_U6IqrDOA3_1(.din(n5502), .dout(n18353));
    jdff dff_A_JFuCtzja3_0(.din(n18353), .dout(n18356));
    jdff dff_A_gBl0FTYb2_0(.din(n18356), .dout(n18359));
    jdff dff_A_1U6gpGID3_0(.din(n18359), .dout(n18362));
    jdff dff_A_tzfrMzca0_0(.din(n18362), .dout(n18365));
    jdff dff_A_7nS1bCmI1_0(.din(n18365), .dout(n18368));
    jdff dff_A_TxHYNhcK3_0(.din(n18368), .dout(n18371));
    jdff dff_A_6joH87FZ8_0(.din(n18371), .dout(n18374));
    jdff dff_A_Q1vsS2BU7_0(.din(n18374), .dout(n18377));
    jdff dff_A_1lOXF1qY7_0(.din(n18377), .dout(n18380));
    jdff dff_A_QxvhYoBx7_0(.din(n18380), .dout(n18383));
    jdff dff_A_SLCOGf525_0(.din(n18383), .dout(n18386));
    jdff dff_A_4roXJf559_0(.din(n18386), .dout(n18389));
    jdff dff_A_r1zjsBTd8_0(.din(n18389), .dout(n18392));
    jdff dff_A_CLtav2Qi1_0(.din(n18392), .dout(n18395));
    jdff dff_A_WF6cgsK41_0(.din(n18395), .dout(n18398));
    jdff dff_A_dJChjvxg0_0(.din(n18398), .dout(n18401));
    jdff dff_A_8ofXVN961_0(.din(n18401), .dout(n18404));
    jdff dff_A_2WY6iaes8_0(.din(n18404), .dout(n18407));
    jdff dff_A_PhvR06020_0(.din(n18407), .dout(n18410));
    jdff dff_A_gZnyTgn10_0(.din(n18410), .dout(n18413));
    jdff dff_A_OovXxVAL4_0(.din(n18413), .dout(n18416));
    jdff dff_A_XeYo21uv6_0(.din(n18416), .dout(n18419));
    jdff dff_A_EoG4hnUo0_0(.din(n18419), .dout(n18422));
    jdff dff_A_Xe6emeEV6_0(.din(n18422), .dout(G923));
    jdff dff_A_NmT0XjCB0_1(.din(n5505), .dout(n18428));
    jdff dff_A_RZMcr9ml7_0(.din(n18428), .dout(n18431));
    jdff dff_A_n5rXPReW6_0(.din(n18431), .dout(n18434));
    jdff dff_A_ixu9Ajnm3_0(.din(n18434), .dout(n18437));
    jdff dff_A_uawdFRIq5_0(.din(n18437), .dout(n18440));
    jdff dff_A_97KL3mNg1_0(.din(n18440), .dout(n18443));
    jdff dff_A_pms3kupZ5_0(.din(n18443), .dout(n18446));
    jdff dff_A_TRzUWzqA9_0(.din(n18446), .dout(n18449));
    jdff dff_A_4GOOIoBm5_0(.din(n18449), .dout(n18452));
    jdff dff_A_ILzC5j1Y5_0(.din(n18452), .dout(n18455));
    jdff dff_A_2KgoG5uF9_0(.din(n18455), .dout(n18458));
    jdff dff_A_rCHZvA3y5_0(.din(n18458), .dout(n18461));
    jdff dff_A_Q8wagKWl2_0(.din(n18461), .dout(n18464));
    jdff dff_A_vlO09x095_0(.din(n18464), .dout(n18467));
    jdff dff_A_hHuvKOIz6_0(.din(n18467), .dout(n18470));
    jdff dff_A_3HceagY58_0(.din(n18470), .dout(n18473));
    jdff dff_A_SlaJdS6O3_0(.din(n18473), .dout(n18476));
    jdff dff_A_Z0wJn0BU4_0(.din(n18476), .dout(n18479));
    jdff dff_A_PMJ4zAW60_0(.din(n18479), .dout(n18482));
    jdff dff_A_0ZzEXFnr9_0(.din(n18482), .dout(n18485));
    jdff dff_A_MVqRmjUv6_0(.din(n18485), .dout(n18488));
    jdff dff_A_iNYzOTkj1_0(.din(n18488), .dout(n18491));
    jdff dff_A_zC9HvHJF1_0(.din(n18491), .dout(n18494));
    jdff dff_A_yEObtYBs5_0(.din(n18494), .dout(n18497));
    jdff dff_A_2jxIV3B49_0(.din(n18497), .dout(G921));
    jdff dff_A_FwI0aGbj2_1(.din(n5508), .dout(n18503));
    jdff dff_A_XHPaJRCE4_0(.din(n18503), .dout(n18506));
    jdff dff_A_Mhc8ZdV60_0(.din(n18506), .dout(n18509));
    jdff dff_A_InkJaXhL9_0(.din(n18509), .dout(n18512));
    jdff dff_A_3k09P2nw0_0(.din(n18512), .dout(n18515));
    jdff dff_A_ndQSjTAy5_0(.din(n18515), .dout(n18518));
    jdff dff_A_z4Vz3Q9U8_0(.din(n18518), .dout(n18521));
    jdff dff_A_MolwkUZP4_0(.din(n18521), .dout(n18524));
    jdff dff_A_lMu4vz877_0(.din(n18524), .dout(n18527));
    jdff dff_A_1xNYFVuB7_0(.din(n18527), .dout(n18530));
    jdff dff_A_92MBFYl93_0(.din(n18530), .dout(n18533));
    jdff dff_A_A1R43ry02_0(.din(n18533), .dout(n18536));
    jdff dff_A_mi3U7mX09_0(.din(n18536), .dout(n18539));
    jdff dff_A_J4z8VsmN4_0(.din(n18539), .dout(n18542));
    jdff dff_A_cALNuMci9_0(.din(n18542), .dout(n18545));
    jdff dff_A_tHyB8OW05_0(.din(n18545), .dout(n18548));
    jdff dff_A_cjPvDO8B7_0(.din(n18548), .dout(n18551));
    jdff dff_A_1vUF3bQz3_0(.din(n18551), .dout(n18554));
    jdff dff_A_OwwzloIQ9_0(.din(n18554), .dout(n18557));
    jdff dff_A_YYP46nOo1_0(.din(n18557), .dout(n18560));
    jdff dff_A_SuKMQElZ8_0(.din(n18560), .dout(n18563));
    jdff dff_A_SeUcB0pi6_0(.din(n18563), .dout(n18566));
    jdff dff_A_TSnMP6gk0_0(.din(n18566), .dout(n18569));
    jdff dff_A_mIPC2zON9_0(.din(n18569), .dout(n18572));
    jdff dff_A_9Ueuxn9R0_0(.din(n18572), .dout(G892));
    jdff dff_A_IM6ysSsv4_1(.din(n5511), .dout(n18578));
    jdff dff_A_zY63OBZr1_0(.din(n18578), .dout(n18581));
    jdff dff_A_ktX1edDQ1_0(.din(n18581), .dout(n18584));
    jdff dff_A_QJZkZGhW5_0(.din(n18584), .dout(n18587));
    jdff dff_A_WAeZpLlO6_0(.din(n18587), .dout(n18590));
    jdff dff_A_A7bdGS0l1_0(.din(n18590), .dout(n18593));
    jdff dff_A_XlA4f5kQ4_0(.din(n18593), .dout(n18596));
    jdff dff_A_e4AlmKNp9_0(.din(n18596), .dout(n18599));
    jdff dff_A_aKQt76y24_0(.din(n18599), .dout(n18602));
    jdff dff_A_a3EsAeRB6_0(.din(n18602), .dout(n18605));
    jdff dff_A_PoGMbfkG8_0(.din(n18605), .dout(n18608));
    jdff dff_A_QJOSBcQ79_0(.din(n18608), .dout(n18611));
    jdff dff_A_qh2QGmt83_0(.din(n18611), .dout(n18614));
    jdff dff_A_tPJmWqXF3_0(.din(n18614), .dout(n18617));
    jdff dff_A_6j2Kddnx8_0(.din(n18617), .dout(n18620));
    jdff dff_A_VJkgFuuW7_0(.din(n18620), .dout(n18623));
    jdff dff_A_NmESWnZK6_0(.din(n18623), .dout(n18626));
    jdff dff_A_SHBUuRdc2_0(.din(n18626), .dout(n18629));
    jdff dff_A_JV1R3ej42_0(.din(n18629), .dout(n18632));
    jdff dff_A_7uLaISER7_0(.din(n18632), .dout(n18635));
    jdff dff_A_Gl01ovTA0_0(.din(n18635), .dout(n18638));
    jdff dff_A_c9eWRvHJ3_0(.din(n18638), .dout(n18641));
    jdff dff_A_2zS9LLHd5_0(.din(n18641), .dout(n18644));
    jdff dff_A_q7TqjPED9_0(.din(n18644), .dout(n18647));
    jdff dff_A_r9Ba313H0_0(.din(n18647), .dout(G887));
    jdff dff_A_ELUGCjOB6_1(.din(n5514), .dout(n18653));
    jdff dff_A_nCOVKXJW4_0(.din(n18653), .dout(n18656));
    jdff dff_A_gDFQfVk81_0(.din(n18656), .dout(n18659));
    jdff dff_A_x1x58NKi6_0(.din(n18659), .dout(n18662));
    jdff dff_A_DADGKog67_0(.din(n18662), .dout(n18665));
    jdff dff_A_s3y8BDx91_0(.din(n18665), .dout(n18668));
    jdff dff_A_adgIwvf93_0(.din(n18668), .dout(n18671));
    jdff dff_A_uQ4JskQk3_0(.din(n18671), .dout(n18674));
    jdff dff_A_DdINJAaW6_0(.din(n18674), .dout(n18677));
    jdff dff_A_3n3LtgKK4_0(.din(n18677), .dout(n18680));
    jdff dff_A_6ZgYHm3y4_0(.din(n18680), .dout(n18683));
    jdff dff_A_mBmZXUZ80_0(.din(n18683), .dout(n18686));
    jdff dff_A_rsAcAc5H9_0(.din(n18686), .dout(n18689));
    jdff dff_A_XtXrAGbu0_0(.din(n18689), .dout(n18692));
    jdff dff_A_tyukI0qE2_0(.din(n18692), .dout(n18695));
    jdff dff_A_DsSsIf3L7_0(.din(n18695), .dout(n18698));
    jdff dff_A_qHLc86ct6_0(.din(n18698), .dout(n18701));
    jdff dff_A_shdq50ZH0_0(.din(n18701), .dout(n18704));
    jdff dff_A_j5IFX4Zg0_0(.din(n18704), .dout(n18707));
    jdff dff_A_vCy38a642_0(.din(n18707), .dout(n18710));
    jdff dff_A_VD7wn6bm6_0(.din(n18710), .dout(n18713));
    jdff dff_A_TJXtEoKU1_0(.din(n18713), .dout(n18716));
    jdff dff_A_JO5766qF6_0(.din(n18716), .dout(n18719));
    jdff dff_A_4rNpAa2X8_0(.din(n18719), .dout(n18722));
    jdff dff_A_Z42TPgXx5_0(.din(n18722), .dout(G606));
    jdff dff_A_keD9V7g93_2(.din(n377), .dout(n18728));
    jdff dff_A_6No7jZ3l5_0(.din(n18728), .dout(n18731));
    jdff dff_A_YwCOvnJB1_0(.din(n18731), .dout(n18734));
    jdff dff_A_e2Zwj5m62_0(.din(n18734), .dout(n18737));
    jdff dff_A_jj23SIgP4_0(.din(n18737), .dout(n18740));
    jdff dff_A_IpvWiYMh2_0(.din(n18740), .dout(n18743));
    jdff dff_A_RRAU7Feh9_0(.din(n18743), .dout(n18746));
    jdff dff_A_Rs4lQiv80_0(.din(n18746), .dout(n18749));
    jdff dff_A_TaIA0Syt7_0(.din(n18749), .dout(n18752));
    jdff dff_A_Xl2iu4F66_0(.din(n18752), .dout(n18755));
    jdff dff_A_vTMnpaNz6_0(.din(n18755), .dout(n18758));
    jdff dff_A_D9yertSl6_0(.din(n18758), .dout(n18761));
    jdff dff_A_Yb8R0NBp9_0(.din(n18761), .dout(n18764));
    jdff dff_A_zoiV8HqI0_0(.din(n18764), .dout(n18767));
    jdff dff_A_frH1zcVH3_0(.din(n18767), .dout(n18770));
    jdff dff_A_jlSvN7Gi6_0(.din(n18770), .dout(n18773));
    jdff dff_A_l2yUoy9h5_0(.din(n18773), .dout(n18776));
    jdff dff_A_zoYPNHe88_0(.din(n18776), .dout(n18779));
    jdff dff_A_bwEjAIaO7_0(.din(n18779), .dout(n18782));
    jdff dff_A_w7sR6eES9_0(.din(n18782), .dout(n18785));
    jdff dff_A_AsVarqsG3_0(.din(n18785), .dout(n18788));
    jdff dff_A_uJzgPcEF4_0(.din(n18788), .dout(n18791));
    jdff dff_A_PeVg3iqd4_0(.din(n18791), .dout(G656));
    jdff dff_A_x86FEGCI7_2(.din(n373), .dout(n18797));
    jdff dff_A_QZa27yH73_0(.din(n18797), .dout(n18800));
    jdff dff_A_b9fGvEec6_0(.din(n18800), .dout(n18803));
    jdff dff_A_iGk5muXF6_0(.din(n18803), .dout(n18806));
    jdff dff_A_Gh3424E94_0(.din(n18806), .dout(n18809));
    jdff dff_A_LCebUzlT4_0(.din(n18809), .dout(n18812));
    jdff dff_A_PxdHmspX4_0(.din(n18812), .dout(n18815));
    jdff dff_A_TivC2nGk7_0(.din(n18815), .dout(n18818));
    jdff dff_A_u9Lazg1R2_0(.din(n18818), .dout(n18821));
    jdff dff_A_Vsi66rb35_0(.din(n18821), .dout(n18824));
    jdff dff_A_Z1fiM0vR6_0(.din(n18824), .dout(n18827));
    jdff dff_A_3NZ0yDjb3_0(.din(n18827), .dout(n18830));
    jdff dff_A_6SUEWyFS5_0(.din(n18830), .dout(n18833));
    jdff dff_A_YSCxAza49_0(.din(n18833), .dout(n18836));
    jdff dff_A_BlGFREtI4_0(.din(n18836), .dout(n18839));
    jdff dff_A_s5FtIMzv5_0(.din(n18839), .dout(n18842));
    jdff dff_A_00AvwFTZ2_0(.din(n18842), .dout(n18845));
    jdff dff_A_hhMxq2Tc8_0(.din(n18845), .dout(n18848));
    jdff dff_A_fMEkWrrV5_0(.din(n18848), .dout(n18851));
    jdff dff_A_rkNNEXs64_0(.din(n18851), .dout(n18854));
    jdff dff_A_aOJlDXK89_0(.din(n18854), .dout(n18857));
    jdff dff_A_vS5vbLYA1_0(.din(n18857), .dout(n18860));
    jdff dff_A_KofkMd3a9_0(.din(n18860), .dout(n18863));
    jdff dff_A_0g7TGgoS7_0(.din(n18863), .dout(G809));
    jdff dff_A_YeaIpaov7_1(.din(n5517), .dout(n18869));
    jdff dff_A_jiXK9IhC9_0(.din(n18869), .dout(n18872));
    jdff dff_A_0iaZKLE90_0(.din(n18872), .dout(n18875));
    jdff dff_A_o39kVAQT8_0(.din(n18875), .dout(n18878));
    jdff dff_A_BtRLGDEP0_0(.din(n18878), .dout(n18881));
    jdff dff_A_99i7LAPF7_0(.din(n18881), .dout(n18884));
    jdff dff_A_57O3sZWL4_0(.din(n18884), .dout(n18887));
    jdff dff_A_xlNFVysj3_0(.din(n18887), .dout(n18890));
    jdff dff_A_XrLXivbj2_0(.din(n18890), .dout(n18893));
    jdff dff_A_L6iGirEZ7_0(.din(n18893), .dout(n18896));
    jdff dff_A_2JxubHvP6_0(.din(n18896), .dout(n18899));
    jdff dff_A_BZKSH1bR1_0(.din(n18899), .dout(n18902));
    jdff dff_A_o1MoDGsA2_0(.din(n18902), .dout(n18905));
    jdff dff_A_MkJoJj2e9_0(.din(n18905), .dout(n18908));
    jdff dff_A_948uc08y8_0(.din(n18908), .dout(n18911));
    jdff dff_A_zRXXoYv12_0(.din(n18911), .dout(n18914));
    jdff dff_A_Z9DbpMDw3_0(.din(n18914), .dout(n18917));
    jdff dff_A_wFCG80GU4_0(.din(n18917), .dout(n18920));
    jdff dff_A_aygIYzC69_0(.din(n18920), .dout(n18923));
    jdff dff_A_xwJ2ZW0q4_0(.din(n18923), .dout(n18926));
    jdff dff_A_KwXllmL38_0(.din(n18926), .dout(n18929));
    jdff dff_A_Ebnw4n3T0_0(.din(n18929), .dout(n18932));
    jdff dff_A_GLVGhJ037_0(.din(n18932), .dout(n18935));
    jdff dff_A_jcMUFEnB7_0(.din(n18935), .dout(n18938));
    jdff dff_A_TvHVLmIo4_0(.din(n18938), .dout(G993));
    jdff dff_A_SpO2BMhM3_1(.din(n5520), .dout(n18944));
    jdff dff_A_jCo04NMI5_0(.din(n18944), .dout(n18947));
    jdff dff_A_47nucgNw2_0(.din(n18947), .dout(n18950));
    jdff dff_A_kWzdgH5L4_0(.din(n18950), .dout(n18953));
    jdff dff_A_UqajSPWh9_0(.din(n18953), .dout(n18956));
    jdff dff_A_JKzZdKFE9_0(.din(n18956), .dout(n18959));
    jdff dff_A_jJba68X70_0(.din(n18959), .dout(n18962));
    jdff dff_A_4GlW8KNG1_0(.din(n18962), .dout(n18965));
    jdff dff_A_uFgZRCcw0_0(.din(n18965), .dout(n18968));
    jdff dff_A_X5fIxnN13_0(.din(n18968), .dout(n18971));
    jdff dff_A_UXfhf2CA5_0(.din(n18971), .dout(n18974));
    jdff dff_A_nRP8m8mD1_0(.din(n18974), .dout(n18977));
    jdff dff_A_aiFZ5ciw2_0(.din(n18977), .dout(n18980));
    jdff dff_A_qHkjQACn7_0(.din(n18980), .dout(n18983));
    jdff dff_A_qjEkwSO13_0(.din(n18983), .dout(n18986));
    jdff dff_A_s81eWuvH7_0(.din(n18986), .dout(n18989));
    jdff dff_A_Mw9uFUtC9_0(.din(n18989), .dout(n18992));
    jdff dff_A_8PszQ2VZ8_0(.din(n18992), .dout(n18995));
    jdff dff_A_kQXK6ufu9_0(.din(n18995), .dout(n18998));
    jdff dff_A_03d5zdZt4_0(.din(n18998), .dout(n19001));
    jdff dff_A_meMuVMTn9_0(.din(n19001), .dout(n19004));
    jdff dff_A_4VSEAS7z3_0(.din(n19004), .dout(n19007));
    jdff dff_A_OhWZ7Kp21_0(.din(n19007), .dout(n19010));
    jdff dff_A_L5bNWsc53_0(.din(n19010), .dout(n19013));
    jdff dff_A_OtBO3pev2_0(.din(n19013), .dout(G978));
    jdff dff_A_abVhkHvY7_1(.din(n5523), .dout(n19019));
    jdff dff_A_V85JZFxw4_0(.din(n19019), .dout(n19022));
    jdff dff_A_d3Gpi8Jc0_0(.din(n19022), .dout(n19025));
    jdff dff_A_jcmEfclu4_0(.din(n19025), .dout(n19028));
    jdff dff_A_Yb6Nbclj0_0(.din(n19028), .dout(n19031));
    jdff dff_A_R1AK6bSL6_0(.din(n19031), .dout(n19034));
    jdff dff_A_R8FvGvkB6_0(.din(n19034), .dout(n19037));
    jdff dff_A_kcFAIxA96_0(.din(n19037), .dout(n19040));
    jdff dff_A_qZIX0z0i8_0(.din(n19040), .dout(n19043));
    jdff dff_A_famX9DUw0_0(.din(n19043), .dout(n19046));
    jdff dff_A_gNC84Z308_0(.din(n19046), .dout(n19049));
    jdff dff_A_ofIv66Zj4_0(.din(n19049), .dout(n19052));
    jdff dff_A_w6uY1qWn7_0(.din(n19052), .dout(n19055));
    jdff dff_A_6LpPMPaN4_0(.din(n19055), .dout(n19058));
    jdff dff_A_xEfkJmnA8_0(.din(n19058), .dout(n19061));
    jdff dff_A_8G9h2CEO0_0(.din(n19061), .dout(n19064));
    jdff dff_A_XKpVDc3B3_0(.din(n19064), .dout(n19067));
    jdff dff_A_ebKE19mp1_0(.din(n19067), .dout(n19070));
    jdff dff_A_lBxUdizI1_0(.din(n19070), .dout(n19073));
    jdff dff_A_XRZtbF221_0(.din(n19073), .dout(n19076));
    jdff dff_A_FUWpOhri7_0(.din(n19076), .dout(n19079));
    jdff dff_A_eOzo2qa53_0(.din(n19079), .dout(n19082));
    jdff dff_A_jznu23Zk0_0(.din(n19082), .dout(n19085));
    jdff dff_A_9YXdI7EP2_0(.din(n19085), .dout(n19088));
    jdff dff_A_ML9mQqH98_0(.din(n19088), .dout(G949));
    jdff dff_A_qpWbjoOy4_1(.din(n5526), .dout(n19094));
    jdff dff_A_oaFPvoaF5_0(.din(n19094), .dout(n19097));
    jdff dff_A_TrKS8yWm2_0(.din(n19097), .dout(n19100));
    jdff dff_A_E4VJRHTl3_0(.din(n19100), .dout(n19103));
    jdff dff_A_mXSY4zYP5_0(.din(n19103), .dout(n19106));
    jdff dff_A_w9A5TP2H2_0(.din(n19106), .dout(n19109));
    jdff dff_A_VlZUHRa21_0(.din(n19109), .dout(n19112));
    jdff dff_A_IvtZ7P7g1_0(.din(n19112), .dout(n19115));
    jdff dff_A_BfS3k26j9_0(.din(n19115), .dout(n19118));
    jdff dff_A_JOfFvtra7_0(.din(n19118), .dout(n19121));
    jdff dff_A_KvfZLhqi5_0(.din(n19121), .dout(n19124));
    jdff dff_A_9y1c4S6c9_0(.din(n19124), .dout(n19127));
    jdff dff_A_ZojNuHXZ5_0(.din(n19127), .dout(n19130));
    jdff dff_A_xpH9CXJM5_0(.din(n19130), .dout(n19133));
    jdff dff_A_fKaLlKz50_0(.din(n19133), .dout(n19136));
    jdff dff_A_6MgvSZpQ6_0(.din(n19136), .dout(n19139));
    jdff dff_A_AqsUbGqI2_0(.din(n19139), .dout(n19142));
    jdff dff_A_sHrKWhtn6_0(.din(n19142), .dout(n19145));
    jdff dff_A_k4QmlshR7_0(.din(n19145), .dout(n19148));
    jdff dff_A_ptLqqP2h2_0(.din(n19148), .dout(n19151));
    jdff dff_A_TiUNK2D95_0(.din(n19151), .dout(n19154));
    jdff dff_A_uKi4mG2o3_0(.din(n19154), .dout(n19157));
    jdff dff_A_EstgPHQC2_0(.din(n19157), .dout(n19160));
    jdff dff_A_TkpcScS52_0(.din(n19160), .dout(n19163));
    jdff dff_A_wsNhdpVO8_0(.din(n19163), .dout(G939));
    jdff dff_A_lD6XExhc7_1(.din(n5529), .dout(n19169));
    jdff dff_A_Jl4ZNpnA1_0(.din(n19169), .dout(n19172));
    jdff dff_A_YRcS2ikS6_0(.din(n19172), .dout(n19175));
    jdff dff_A_c9n10fjS4_0(.din(n19175), .dout(n19178));
    jdff dff_A_QTjUCbq50_0(.din(n19178), .dout(n19181));
    jdff dff_A_XMibHe3f4_0(.din(n19181), .dout(n19184));
    jdff dff_A_Hgy08DiC8_0(.din(n19184), .dout(n19187));
    jdff dff_A_ty6mWJ6Y6_0(.din(n19187), .dout(n19190));
    jdff dff_A_NcpEUnwM2_0(.din(n19190), .dout(n19193));
    jdff dff_A_zHy5uA2U5_0(.din(n19193), .dout(n19196));
    jdff dff_A_k6LFJOLP7_0(.din(n19196), .dout(n19199));
    jdff dff_A_GQGhDm5G4_0(.din(n19199), .dout(n19202));
    jdff dff_A_iiw7dC0S9_0(.din(n19202), .dout(n19205));
    jdff dff_A_pGv4YvHQ3_0(.din(n19205), .dout(n19208));
    jdff dff_A_ReWdVeme4_0(.din(n19208), .dout(n19211));
    jdff dff_A_IDiLCvME8_0(.din(n19211), .dout(n19214));
    jdff dff_A_ATyGnFjX3_0(.din(n19214), .dout(n19217));
    jdff dff_A_FsvZQZ7i2_0(.din(n19217), .dout(n19220));
    jdff dff_A_RsX6UkSY0_0(.din(n19220), .dout(n19223));
    jdff dff_A_EsQzUZc85_0(.din(n19223), .dout(n19226));
    jdff dff_A_brVQAggx3_0(.din(n19226), .dout(n19229));
    jdff dff_A_cwqWPGr07_0(.din(n19229), .dout(n19232));
    jdff dff_A_dVrG7hGV7_0(.din(n19232), .dout(n19235));
    jdff dff_A_FrYoED5t0_0(.din(n19235), .dout(n19238));
    jdff dff_A_TpleHrMc4_0(.din(n19238), .dout(G889));
    jdff dff_A_4e4EIA5N1_1(.din(n380), .dout(n19244));
    jdff dff_A_NNj3eLVc1_0(.din(n19244), .dout(n19247));
    jdff dff_A_3HlQ2bnD6_0(.din(n19247), .dout(n19250));
    jdff dff_A_K0APsira4_0(.din(n19250), .dout(n19253));
    jdff dff_A_5mirhI067_0(.din(n19253), .dout(n19256));
    jdff dff_A_SgChimeS9_0(.din(n19256), .dout(n19259));
    jdff dff_A_I7tJAHJo4_0(.din(n19259), .dout(n19262));
    jdff dff_A_jEORaBQ79_0(.din(n19262), .dout(n19265));
    jdff dff_A_981HW88k6_0(.din(n19265), .dout(n19268));
    jdff dff_A_rAG8wnC35_0(.din(n19268), .dout(n19271));
    jdff dff_A_yEMSOdVg2_0(.din(n19271), .dout(n19274));
    jdff dff_A_7H2nFOht3_0(.din(n19274), .dout(n19277));
    jdff dff_A_0fRBeq0C1_0(.din(n19277), .dout(n19280));
    jdff dff_A_8X4qeEpt1_0(.din(n19280), .dout(n19283));
    jdff dff_A_ja6OvJz09_0(.din(n19283), .dout(n19286));
    jdff dff_A_FpJLk7TL0_0(.din(n19286), .dout(n19289));
    jdff dff_A_LzWbjckA9_0(.din(n19289), .dout(n19292));
    jdff dff_A_s9R8RfWi8_0(.din(n19292), .dout(n19295));
    jdff dff_A_pqgIY3NN1_0(.din(n19295), .dout(n19298));
    jdff dff_A_26dtetRk3_0(.din(n19298), .dout(n19301));
    jdff dff_A_h3Zg1kjR9_0(.din(n19301), .dout(n19304));
    jdff dff_A_EtvJhjP99_0(.din(n19304), .dout(n19307));
    jdff dff_A_yiqcB09d7_0(.din(n19307), .dout(n19310));
    jdff dff_A_iCRYLmRz2_0(.din(n19310), .dout(n19313));
    jdff dff_A_Uhx4mFUf4_0(.din(n19313), .dout(G593));
    jdff dff_A_5DKWnxSc5_2(.din(n405), .dout(n19319));
    jdff dff_A_xVQWH6Tr1_0(.din(n19319), .dout(n19322));
    jdff dff_A_uI2A11gr1_0(.din(n19322), .dout(n19325));
    jdff dff_A_xr7y9Smy1_0(.din(n19325), .dout(n19328));
    jdff dff_A_E4DmUa6Y8_0(.din(n19328), .dout(n19331));
    jdff dff_A_KCPLWmcP4_0(.din(n19331), .dout(n19334));
    jdff dff_A_6WVWdltR0_0(.din(n19334), .dout(n19337));
    jdff dff_A_ahA86vOb6_0(.din(n19337), .dout(n19340));
    jdff dff_A_6KcVJOQL8_0(.din(n19340), .dout(n19343));
    jdff dff_A_oIjlbJoV5_0(.din(n19343), .dout(n19346));
    jdff dff_A_x57fBEvW9_0(.din(n19346), .dout(n19349));
    jdff dff_A_YwmGE3Am3_0(.din(n19349), .dout(n19352));
    jdff dff_A_pd1p2vGz2_0(.din(n19352), .dout(n19355));
    jdff dff_A_nKTgTCH18_0(.din(n19355), .dout(n19358));
    jdff dff_A_QP5hFykY0_0(.din(n19358), .dout(n19361));
    jdff dff_A_WeoXHbwr4_0(.din(n19361), .dout(n19364));
    jdff dff_A_Ydk4Ner15_0(.din(n19364), .dout(n19367));
    jdff dff_A_uI1fL5E10_0(.din(n19367), .dout(n19370));
    jdff dff_A_NhiN46YI3_0(.din(n19370), .dout(n19373));
    jdff dff_A_BvVZYSyB5_0(.din(n19373), .dout(n19376));
    jdff dff_A_CPpuDR8l0_0(.din(n19376), .dout(n19379));
    jdff dff_A_2AJPeBJv2_0(.din(n19379), .dout(G636));
    jdff dff_A_CXKw5YL30_2(.din(n427), .dout(n19385));
    jdff dff_A_sN8DakQO6_0(.din(n19385), .dout(n19388));
    jdff dff_A_JcOoUIoU0_0(.din(n19388), .dout(n19391));
    jdff dff_A_AMQ9nWoi5_0(.din(n19391), .dout(n19394));
    jdff dff_A_ffv8D3iP0_0(.din(n19394), .dout(n19397));
    jdff dff_A_NLkBdWcm3_0(.din(n19397), .dout(n19400));
    jdff dff_A_rkUBQDy35_0(.din(n19400), .dout(n19403));
    jdff dff_A_gYFtotOP3_0(.din(n19403), .dout(n19406));
    jdff dff_A_WHcSynkR0_0(.din(n19406), .dout(n19409));
    jdff dff_A_lBDItlpU6_0(.din(n19409), .dout(n19412));
    jdff dff_A_07oRUG598_0(.din(n19412), .dout(n19415));
    jdff dff_A_luXZfeUs5_0(.din(n19415), .dout(n19418));
    jdff dff_A_zVtXFOHs9_0(.din(n19418), .dout(n19421));
    jdff dff_A_WGsCsiRH9_0(.din(n19421), .dout(n19424));
    jdff dff_A_NweTt4l64_0(.din(n19424), .dout(n19427));
    jdff dff_A_if2qgv0H6_0(.din(n19427), .dout(n19430));
    jdff dff_A_wAsJxjbj2_0(.din(n19430), .dout(n19433));
    jdff dff_A_9xIy5x3z4_0(.din(n19433), .dout(n19436));
    jdff dff_A_6JOjYtxb7_0(.din(n19436), .dout(n19439));
    jdff dff_A_cRKkT0PC0_0(.din(n19439), .dout(n19442));
    jdff dff_A_aItKAicj2_0(.din(n19442), .dout(n19445));
    jdff dff_A_wTQCLBXD0_0(.din(n19445), .dout(G704));
    jdff dff_A_TR3QSKJ91_2(.din(n5533), .dout(n19451));
    jdff dff_A_RkLtvXpE6_0(.din(n19451), .dout(n19454));
    jdff dff_A_z0TMj8TG3_0(.din(n19454), .dout(n19457));
    jdff dff_A_64wFIkQ95_0(.din(n19457), .dout(n19460));
    jdff dff_A_puWSMKTF7_0(.din(n19460), .dout(n19463));
    jdff dff_A_dk9tfpKv2_0(.din(n19463), .dout(n19466));
    jdff dff_A_8tTZc8Kw2_0(.din(n19466), .dout(n19469));
    jdff dff_A_Xevm6M2H3_0(.din(n19469), .dout(n19472));
    jdff dff_A_FyPeZUxw6_0(.din(n19472), .dout(n19475));
    jdff dff_A_9aTbQNIu4_0(.din(n19475), .dout(n19478));
    jdff dff_A_nzxuVn7x7_0(.din(n19478), .dout(n19481));
    jdff dff_A_gLUPRY4w4_0(.din(n19481), .dout(n19484));
    jdff dff_A_PBKA6CSE2_0(.din(n19484), .dout(n19487));
    jdff dff_A_40L5QOHL3_0(.din(n19487), .dout(n19490));
    jdff dff_A_VDZx6CGd6_0(.din(n19490), .dout(n19493));
    jdff dff_A_wr4CqXl23_0(.din(n19493), .dout(n19496));
    jdff dff_A_TjeCiBd20_0(.din(n19496), .dout(n19499));
    jdff dff_A_jh06xNKB8_0(.din(n19499), .dout(n19502));
    jdff dff_A_xpbmMFm96_0(.din(n19502), .dout(n19505));
    jdff dff_A_3X92xAxM1_0(.din(n19505), .dout(n19508));
    jdff dff_A_3aVTff5Z7_0(.din(n19508), .dout(n19511));
    jdff dff_A_wISkywuW2_0(.din(n19511), .dout(G717));
    jdff dff_A_9yC0VVfO7_2(.din(n434), .dout(n19517));
    jdff dff_A_jFXPlW4o6_0(.din(n19517), .dout(n19520));
    jdff dff_A_xJpXaXBX8_0(.din(n19520), .dout(n19523));
    jdff dff_A_5kSP9aBD0_0(.din(n19523), .dout(n19526));
    jdff dff_A_zNTpmbIP0_0(.din(n19526), .dout(n19529));
    jdff dff_A_a2AJYJZY2_0(.din(n19529), .dout(n19532));
    jdff dff_A_S7QEW4ah1_0(.din(n19532), .dout(n19535));
    jdff dff_A_9NJzThi50_0(.din(n19535), .dout(n19538));
    jdff dff_A_ilQaAq009_0(.din(n19538), .dout(n19541));
    jdff dff_A_I6OnOS4L9_0(.din(n19541), .dout(n19544));
    jdff dff_A_Kqfm5GjQ8_0(.din(n19544), .dout(n19547));
    jdff dff_A_DQQxTDK83_0(.din(n19547), .dout(n19550));
    jdff dff_A_2z7dsrkQ1_0(.din(n19550), .dout(n19553));
    jdff dff_A_7xiub2BF7_0(.din(n19553), .dout(n19556));
    jdff dff_A_pj51po7o9_0(.din(n19556), .dout(n19559));
    jdff dff_A_jekEyZBi1_0(.din(n19559), .dout(n19562));
    jdff dff_A_1mn3SqOD2_0(.din(n19562), .dout(n19565));
    jdff dff_A_A90jU8Hx4_0(.din(n19565), .dout(n19568));
    jdff dff_A_NS9tbqK98_0(.din(n19568), .dout(n19571));
    jdff dff_A_TGZ9z4nW7_0(.din(n19571), .dout(n19574));
    jdff dff_A_ymbLtiM65_0(.din(n19574), .dout(n19577));
    jdff dff_A_D3s1irdO4_0(.din(n19577), .dout(n19580));
    jdff dff_A_lQWDjGuG1_0(.din(n19580), .dout(G820));
    jdff dff_A_rizW0C430_2(.din(n454), .dout(n19586));
    jdff dff_A_KgAAbwuH8_0(.din(n19586), .dout(n19589));
    jdff dff_A_7nnuyk1Q2_0(.din(n19589), .dout(n19592));
    jdff dff_A_vYgPw98P2_0(.din(n19592), .dout(n19595));
    jdff dff_A_GiHiMhTQ7_0(.din(n19595), .dout(n19598));
    jdff dff_A_AUqkSgAN4_0(.din(n19598), .dout(n19601));
    jdff dff_A_aDDEqaYT7_0(.din(n19601), .dout(n19604));
    jdff dff_A_wChBvq3p6_0(.din(n19604), .dout(n19607));
    jdff dff_A_vJm1Pm654_0(.din(n19607), .dout(n19610));
    jdff dff_A_MQroQ7IC1_0(.din(n19610), .dout(n19613));
    jdff dff_A_GiyvZx260_0(.din(n19613), .dout(n19616));
    jdff dff_A_jcrhMJgS8_0(.din(n19616), .dout(n19619));
    jdff dff_A_gs4gCJG75_0(.din(n19619), .dout(n19622));
    jdff dff_A_43PrkEhK8_0(.din(n19622), .dout(n19625));
    jdff dff_A_blgBBLO64_0(.din(n19625), .dout(n19628));
    jdff dff_A_Mn3y9pAO6_0(.din(n19628), .dout(n19631));
    jdff dff_A_OmwUq7pT7_0(.din(n19631), .dout(n19634));
    jdff dff_A_wTIzYJdY3_0(.din(n19634), .dout(n19637));
    jdff dff_A_X6fMt0Zj0_0(.din(n19637), .dout(n19640));
    jdff dff_A_kU02qcPQ1_0(.din(n19640), .dout(n19643));
    jdff dff_A_adtuXUxE0_0(.din(n19643), .dout(G639));
    jdff dff_A_elugQIR87_2(.din(n474), .dout(n19649));
    jdff dff_A_vjOvb3W06_0(.din(n19649), .dout(n19652));
    jdff dff_A_f7oJb32k4_0(.din(n19652), .dout(n19655));
    jdff dff_A_cGLVsDBl2_0(.din(n19655), .dout(n19658));
    jdff dff_A_LAicCfTh9_0(.din(n19658), .dout(n19661));
    jdff dff_A_zPpsueOZ2_0(.din(n19661), .dout(n19664));
    jdff dff_A_ncAURSH36_0(.din(n19664), .dout(n19667));
    jdff dff_A_kCSS4AZq0_0(.din(n19667), .dout(n19670));
    jdff dff_A_NYHD2jE67_0(.din(n19670), .dout(n19673));
    jdff dff_A_oYi4of0D3_0(.din(n19673), .dout(n19676));
    jdff dff_A_Hb4ytExg0_0(.din(n19676), .dout(n19679));
    jdff dff_A_mhiIvyDJ5_0(.din(n19679), .dout(n19682));
    jdff dff_A_GMirbeNl4_0(.din(n19682), .dout(n19685));
    jdff dff_A_6PHqUvff5_0(.din(n19685), .dout(n19688));
    jdff dff_A_NhBUSYdt2_0(.din(n19688), .dout(n19691));
    jdff dff_A_njyrBR860_0(.din(n19691), .dout(n19694));
    jdff dff_A_0fI8E1tn5_0(.din(n19694), .dout(n19697));
    jdff dff_A_LjAQVpdm0_0(.din(n19697), .dout(n19700));
    jdff dff_A_hOjv7GI27_0(.din(n19700), .dout(n19703));
    jdff dff_A_fvRySZuu8_0(.din(n19703), .dout(n19706));
    jdff dff_A_FrydKVP70_0(.din(n19706), .dout(G673));
    jdff dff_A_FaokHENP3_2(.din(n494), .dout(n19712));
    jdff dff_A_0QcR0jCY9_0(.din(n19712), .dout(n19715));
    jdff dff_A_fkXPbOey1_0(.din(n19715), .dout(n19718));
    jdff dff_A_FBlijyyz1_0(.din(n19718), .dout(n19721));
    jdff dff_A_oaAOkGXK3_0(.din(n19721), .dout(n19724));
    jdff dff_A_K7S56rVT4_0(.din(n19724), .dout(n19727));
    jdff dff_A_KCQuRw3E0_0(.din(n19727), .dout(n19730));
    jdff dff_A_fgZNn9MB6_0(.din(n19730), .dout(n19733));
    jdff dff_A_TbSvztVd9_0(.din(n19733), .dout(n19736));
    jdff dff_A_S7lPsxhh1_0(.din(n19736), .dout(n19739));
    jdff dff_A_xOKC3ko35_0(.din(n19739), .dout(n19742));
    jdff dff_A_d3Ip3zeE9_0(.din(n19742), .dout(n19745));
    jdff dff_A_64YrB5C19_0(.din(n19745), .dout(n19748));
    jdff dff_A_iSOwSdHN7_0(.din(n19748), .dout(n19751));
    jdff dff_A_n29ScSW67_0(.din(n19751), .dout(n19754));
    jdff dff_A_xQwsdKbI5_0(.din(n19754), .dout(n19757));
    jdff dff_A_XqEADTOL7_0(.din(n19757), .dout(n19760));
    jdff dff_A_QXQ2Bv1S2_0(.din(n19760), .dout(n19763));
    jdff dff_A_ao6Jk5qP6_0(.din(n19763), .dout(n19766));
    jdff dff_A_xTYZkzUF4_0(.din(n19766), .dout(n19769));
    jdff dff_A_K4tG1aVx5_0(.din(n19769), .dout(G707));
    jdff dff_A_xsbWQ4I27_2(.din(n514), .dout(n19775));
    jdff dff_A_ZmxnlbO75_0(.din(n19775), .dout(n19778));
    jdff dff_A_pGGRNlkO6_0(.din(n19778), .dout(n19781));
    jdff dff_A_vT2fL17A8_0(.din(n19781), .dout(n19784));
    jdff dff_A_HyQ7vQWy2_0(.din(n19784), .dout(n19787));
    jdff dff_A_gUlXqVgu7_0(.din(n19787), .dout(n19790));
    jdff dff_A_mFipyJM54_0(.din(n19790), .dout(n19793));
    jdff dff_A_vnhY7zrE0_0(.din(n19793), .dout(n19796));
    jdff dff_A_zvh8j5m56_0(.din(n19796), .dout(n19799));
    jdff dff_A_NX87CFfs2_0(.din(n19799), .dout(n19802));
    jdff dff_A_bMeo0Xii2_0(.din(n19802), .dout(n19805));
    jdff dff_A_0gDixBLJ5_0(.din(n19805), .dout(n19808));
    jdff dff_A_ShcqrH7E4_0(.din(n19808), .dout(n19811));
    jdff dff_A_uXKUj2lM3_0(.din(n19811), .dout(n19814));
    jdff dff_A_ayzisLxe1_0(.din(n19814), .dout(n19817));
    jdff dff_A_B7C4cCNj4_0(.din(n19817), .dout(n19820));
    jdff dff_A_VyHL6giX3_0(.din(n19820), .dout(n19823));
    jdff dff_A_p7En6qza1_0(.din(n19823), .dout(n19826));
    jdff dff_A_wlaTIjaE6_0(.din(n19826), .dout(n19829));
    jdff dff_A_ASPWIk2T1_0(.din(n19829), .dout(n19832));
    jdff dff_A_6SUGHeB62_0(.din(n19832), .dout(G715));
    jdff dff_A_BEb53Iaq1_2(.din(n846), .dout(n19838));
    jdff dff_A_oloWKfMa0_0(.din(n19838), .dout(n19841));
    jdff dff_A_pqD3GZ3g8_0(.din(n19841), .dout(n19844));
    jdff dff_A_EYGuIKep0_0(.din(n19844), .dout(n19847));
    jdff dff_A_9LMeRw9x6_0(.din(n19847), .dout(n19850));
    jdff dff_A_deNX8pML9_0(.din(n19850), .dout(n19853));
    jdff dff_A_MxDtdVQe0_0(.din(n19853), .dout(n19856));
    jdff dff_A_nl4mcWAu4_0(.din(n19856), .dout(n19859));
    jdff dff_A_ewEv8Ybp9_0(.din(n19859), .dout(n19862));
    jdff dff_A_U6aBBlE37_0(.din(n19862), .dout(n19865));
    jdff dff_A_sgeIN7sc3_0(.din(n19865), .dout(n19868));
    jdff dff_A_P1ICeaaJ8_0(.din(n19868), .dout(n19871));
    jdff dff_A_QA7VTbku3_0(.din(n19871), .dout(n19874));
    jdff dff_A_sgG74Gx40_0(.din(n19874), .dout(n19877));
    jdff dff_A_CUgQ3iz31_0(.din(n19877), .dout(n19880));
    jdff dff_A_aJMDk6zR2_0(.din(n19880), .dout(n19883));
    jdff dff_A_SUtsIFMm6_0(.din(n19883), .dout(G598));
    jdff dff_A_j4efVi3O6_2(.din(n1256), .dout(n19889));
    jdff dff_A_Yq0pu1wW0_0(.din(n19889), .dout(n19892));
    jdff dff_A_GOBiuBFn1_0(.din(n19892), .dout(n19895));
    jdff dff_A_WbbPGbyL9_0(.din(n19895), .dout(n19898));
    jdff dff_A_QUDDyT3N6_0(.din(n19898), .dout(n19901));
    jdff dff_A_SRlVGceg3_0(.din(n19901), .dout(n19904));
    jdff dff_A_uALdLlXS3_0(.din(n19904), .dout(n19907));
    jdff dff_A_5DWrPsbL7_0(.din(n19907), .dout(n19910));
    jdff dff_A_TJ8wjj571_0(.din(n19910), .dout(n19913));
    jdff dff_A_g4gbUWNR7_0(.din(n19913), .dout(n19916));
    jdff dff_A_awoE7okF8_0(.din(n19916), .dout(n19919));
    jdff dff_A_lUxuw5nY6_0(.din(n19919), .dout(n19922));
    jdff dff_A_HON1Q2SL5_0(.din(n19922), .dout(n19925));
    jdff dff_A_VA68RU7z1_0(.din(n19925), .dout(n19928));
    jdff dff_A_iT40JmC66_0(.din(n19928), .dout(n19931));
    jdff dff_A_U5oLsT2f1_0(.din(n19931), .dout(n19934));
    jdff dff_A_I4bktKWu6_0(.din(n19934), .dout(G610));
    jdff dff_A_4Xgg3Wdu6_2(.din(n1459), .dout(n19940));
    jdff dff_A_1M4z8uvC6_0(.din(n19940), .dout(n19943));
    jdff dff_A_5FiHU8d02_0(.din(n19943), .dout(n19946));
    jdff dff_A_tjm3Ww215_0(.din(n19946), .dout(n19949));
    jdff dff_A_71ej5SFX2_0(.din(n19949), .dout(n19952));
    jdff dff_A_TkQReInG0_0(.din(n19952), .dout(n19955));
    jdff dff_A_3Nz5jTUP4_0(.din(n19955), .dout(n19958));
    jdff dff_A_GuaHMZHy1_0(.din(n19958), .dout(n19961));
    jdff dff_A_G3Nt3byh6_0(.din(n19961), .dout(n19964));
    jdff dff_A_CJkqSmBs2_0(.din(n19964), .dout(n19967));
    jdff dff_A_MN2Ias6m6_0(.din(n19967), .dout(n19970));
endmodule

