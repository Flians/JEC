module gf_c880(G268gat, G267gat, G111gat, G87gat, G130gat, G159gat, G261gat, G101gat, G152gat, G86gat, G29gat, G13gat, G106gat, G74gat, G96gat, G91gat, G149gat, G73gat, G80gat, G138gat, G72gat, G90gat, G8gat, G51gat, G143gat, G26gat, G55gat, G36gat, G153gat, G17gat, G246gat, G85gat, G59gat, G116gat, G121gat, G146gat, G126gat, G135gat, G89gat, G219gat, G68gat, G156gat, G165gat, G42gat, G171gat, G177gat, G195gat, G259gat, G183gat, G88gat, G189gat, G210gat, G237gat, G201gat, G75gat, G1gat, G207gat, G228gat, G255gat, G260gat, G879gat, G878gat, G874gat, G865gat, G864gat, G767gat, G450gat, G423gat, G850gat, G389gat, G390gat, G447gat, G880gat, G449gat, G391gat, G418gat, G863gat, G419gat, G768gat, G422gat, G420gat, G421gat, G448gat, G866gat, G388gat, G446gat);
    input G268gat, G267gat, G111gat, G87gat, G130gat, G159gat, G261gat, G101gat, G152gat, G86gat, G29gat, G13gat, G106gat, G74gat, G96gat, G91gat, G149gat, G73gat, G80gat, G138gat, G72gat, G90gat, G8gat, G51gat, G143gat, G26gat, G55gat, G36gat, G153gat, G17gat, G246gat, G85gat, G59gat, G116gat, G121gat, G146gat, G126gat, G135gat, G89gat, G219gat, G68gat, G156gat, G165gat, G42gat, G171gat, G177gat, G195gat, G259gat, G183gat, G88gat, G189gat, G210gat, G237gat, G201gat, G75gat, G1gat, G207gat, G228gat, G255gat, G260gat;
    output G879gat, G878gat, G874gat, G865gat, G864gat, G767gat, G450gat, G423gat, G850gat, G389gat, G390gat, G447gat, G880gat, G449gat, G391gat, G418gat, G863gat, G419gat, G768gat, G422gat, G420gat, G421gat, G448gat, G866gat, G388gat, G446gat;
    wire n89;
    wire n93;
    wire n97;
    wire n101;
    wire n105;
    wire n109;
    wire n113;
    wire n117;
    wire n121;
    wire n124;
    wire n127;
    wire n130;
    wire n133;
    wire n137;
    wire n141;
    wire n145;
    wire n149;
    wire n152;
    wire n156;
    wire n159;
    wire n163;
    wire n166;
    wire n169;
    wire n173;
    wire n177;
    wire n180;
    wire n184;
    wire n188;
    wire n192;
    wire n195;
    wire n199;
    wire n203;
    wire n207;
    wire n211;
    wire n215;
    wire n219;
    wire n223;
    wire n227;
    wire n231;
    wire n235;
    wire n239;
    wire n243;
    wire n247;
    wire n251;
    wire n255;
    wire n259;
    wire n263;
    wire n267;
    wire n271;
    wire n275;
    wire n279;
    wire n283;
    wire n287;
    wire n291;
    wire n295;
    wire n299;
    wire n303;
    wire n307;
    wire n310;
    wire n314;
    wire n318;
    wire n322;
    wire n326;
    wire n330;
    wire n333;
    wire n337;
    wire n341;
    wire n344;
    wire n348;
    wire n352;
    wire n356;
    wire n359;
    wire n363;
    wire n367;
    wire n370;
    wire n374;
    wire n378;
    wire n381;
    wire n385;
    wire n389;
    wire n392;
    wire n396;
    wire n400;
    wire n404;
    wire n408;
    wire n412;
    wire n416;
    wire n420;
    wire n424;
    wire n428;
    wire n432;
    wire n436;
    wire n440;
    wire n444;
    wire n448;
    wire n451;
    wire n454;
    wire n457;
    wire n460;
    wire n464;
    wire n468;
    wire n472;
    wire n476;
    wire n480;
    wire n484;
    wire n487;
    wire n491;
    wire n495;
    wire n499;
    wire n503;
    wire n507;
    wire n511;
    wire n515;
    wire n519;
    wire n523;
    wire n527;
    wire n531;
    wire n535;
    wire n539;
    wire n543;
    wire n547;
    wire n551;
    wire n555;
    wire n558;
    wire n561;
    wire n565;
    wire n569;
    wire n573;
    wire n577;
    wire n581;
    wire n585;
    wire n589;
    wire n593;
    wire n597;
    wire n601;
    wire n605;
    wire n609;
    wire n613;
    wire n617;
    wire n621;
    wire n625;
    wire n629;
    wire n633;
    wire n637;
    wire n641;
    wire n645;
    wire n649;
    wire n653;
    wire n657;
    wire n661;
    wire n665;
    wire n669;
    wire n673;
    wire n677;
    wire n681;
    wire n685;
    wire n689;
    wire n692;
    wire n696;
    wire n700;
    wire n704;
    wire n708;
    wire n712;
    wire n716;
    wire n720;
    wire n723;
    wire n726;
    wire n729;
    wire n732;
    wire n735;
    wire n739;
    wire n743;
    wire n747;
    wire n751;
    wire n755;
    wire n759;
    wire n763;
    wire n767;
    wire n771;
    wire n775;
    wire n779;
    wire n783;
    wire n787;
    wire n791;
    wire n795;
    wire n799;
    wire n803;
    wire n807;
    wire n811;
    wire n815;
    wire n819;
    wire n823;
    wire n827;
    wire n831;
    wire n834;
    wire n838;
    wire n842;
    wire n846;
    wire n850;
    wire n854;
    wire n858;
    wire n862;
    wire n866;
    wire n870;
    wire n874;
    wire n878;
    wire n882;
    wire n886;
    wire n890;
    wire n894;
    wire n898;
    wire n902;
    wire n905;
    wire n909;
    wire n913;
    wire n917;
    wire n921;
    wire n925;
    wire n929;
    wire n933;
    wire n937;
    wire n941;
    wire n945;
    wire n949;
    wire n953;
    wire n957;
    wire n961;
    wire n965;
    wire n969;
    wire n973;
    wire n977;
    wire n981;
    wire n985;
    wire n989;
    wire n993;
    wire n997;
    wire n1001;
    wire n1005;
    wire n1009;
    wire n1013;
    wire n1017;
    wire n1021;
    wire n1025;
    wire n1029;
    wire n1033;
    wire n1037;
    wire n1041;
    wire n1045;
    wire n1049;
    wire n1053;
    wire n1057;
    wire n1060;
    wire n1063;
    wire n1067;
    wire n1070;
    wire n1073;
    wire n1076;
    wire n1080;
    wire n1083;
    wire n1087;
    wire n1091;
    wire n1095;
    wire n1099;
    wire n1103;
    wire n1107;
    wire n1111;
    wire n1115;
    wire n1119;
    wire n1123;
    wire n1127;
    wire n1130;
    wire n1134;
    wire n1138;
    wire n1141;
    wire n1145;
    wire n1149;
    wire n1153;
    wire n1157;
    wire n1161;
    wire n1165;
    wire n1169;
    wire n1173;
    wire n1177;
    wire n1181;
    wire n1185;
    wire n1189;
    wire n1193;
    wire n1197;
    wire n1201;
    wire n1205;
    wire n1209;
    wire n1213;
    wire n1217;
    wire n1221;
    wire n1225;
    wire n1229;
    wire n1233;
    wire n1237;
    wire n1241;
    wire n1244;
    wire n1247;
    wire n1250;
    wire n1253;
    wire n1256;
    wire n1260;
    wire n1264;
    wire n1268;
    wire n1272;
    wire n1276;
    wire n1280;
    wire n1283;
    wire n1287;
    wire n1291;
    wire n1295;
    wire n1303;
    wire n1307;
    wire n1311;
    wire n1315;
    wire n1319;
    wire n1323;
    wire n1327;
    wire n1331;
    wire n1335;
    wire n1339;
    wire n1343;
    wire n1346;
    wire n1350;
    wire n1354;
    wire n1358;
    wire n1362;
    wire n1366;
    wire n1370;
    wire n1374;
    wire n1378;
    wire n1382;
    wire n1386;
    wire n1390;
    wire n1394;
    wire n1398;
    wire n1402;
    wire n1405;
    wire n1409;
    wire n1413;
    wire n1417;
    wire n1421;
    wire n1425;
    wire n2043;
    wire n2046;
    wire n2049;
    wire n2052;
    wire n2054;
    wire n2057;
    wire n2061;
    wire n2064;
    wire n2067;
    wire n2070;
    wire n2073;
    wire n2076;
    wire n2079;
    wire n2081;
    wire n2085;
    wire n2088;
    wire n2091;
    wire n2094;
    wire n2097;
    wire n2100;
    wire n2103;
    wire n2106;
    wire n2109;
    wire n2112;
    wire n2115;
    wire n2118;
    wire n2121;
    wire n2124;
    wire n2127;
    wire n2130;
    wire n2133;
    wire n2136;
    wire n2139;
    wire n2142;
    wire n2144;
    wire n2147;
    wire n2150;
    wire n2153;
    wire n2157;
    wire n2160;
    wire n2163;
    wire n2166;
    wire n2169;
    wire n2172;
    wire n2175;
    wire n2178;
    wire n2181;
    wire n2184;
    wire n2187;
    wire n2190;
    wire n2193;
    wire n2196;
    wire n2199;
    wire n2202;
    wire n2205;
    wire n2208;
    wire n2211;
    wire n2214;
    wire n2217;
    wire n2220;
    wire n2223;
    wire n2226;
    wire n2229;
    wire n2232;
    wire n2235;
    wire n2238;
    wire n2241;
    wire n2243;
    wire n2246;
    wire n2249;
    wire n2252;
    wire n2255;
    wire n2258;
    wire n2261;
    wire n2264;
    wire n2267;
    wire n2270;
    wire n2273;
    wire n2276;
    wire n2279;
    wire n2282;
    wire n2285;
    wire n2288;
    wire n2291;
    wire n2294;
    wire n2297;
    wire n2300;
    wire n2303;
    wire n2306;
    wire n2310;
    wire n2313;
    wire n2316;
    wire n2319;
    wire n2322;
    wire n2325;
    wire n2328;
    wire n2331;
    wire n2334;
    wire n2337;
    wire n2339;
    wire n2342;
    wire n2345;
    wire n2348;
    wire n2351;
    wire n2354;
    wire n2357;
    wire n2360;
    wire n2364;
    wire n2367;
    wire n2370;
    wire n2373;
    wire n2376;
    wire n2379;
    wire n2382;
    wire n2385;
    wire n2388;
    wire n2391;
    wire n2394;
    wire n2397;
    wire n2400;
    wire n2403;
    wire n2406;
    wire n2409;
    wire n2412;
    wire n2415;
    wire n2418;
    wire n2421;
    wire n2424;
    wire n2427;
    wire n2430;
    wire n2432;
    wire n2435;
    wire n2438;
    wire n2441;
    wire n2444;
    wire n2448;
    wire n2451;
    wire n2454;
    wire n2457;
    wire n2460;
    wire n2463;
    wire n2466;
    wire n2469;
    wire n2472;
    wire n2475;
    wire n2478;
    wire n2481;
    wire n2484;
    wire n2487;
    wire n2490;
    wire n2493;
    wire n2496;
    wire n2499;
    wire n2502;
    wire n2505;
    wire n2508;
    wire n2511;
    wire n2514;
    wire n2517;
    wire n2520;
    wire n2523;
    wire n2526;
    wire n2529;
    wire n2532;
    wire n2534;
    wire n2537;
    wire n2540;
    wire n2544;
    wire n2547;
    wire n2550;
    wire n2553;
    wire n2556;
    wire n2559;
    wire n2562;
    wire n2565;
    wire n2568;
    wire n2571;
    wire n2574;
    wire n2577;
    wire n2580;
    wire n2583;
    wire n2586;
    wire n2589;
    wire n2592;
    wire n2595;
    wire n2598;
    wire n2601;
    wire n2604;
    wire n2607;
    wire n2610;
    wire n2613;
    wire n2616;
    wire n2619;
    wire n2622;
    wire n2625;
    wire n2628;
    wire n2630;
    wire n2633;
    wire n2636;
    wire n2639;
    wire n2642;
    wire n2645;
    wire n2648;
    wire n2651;
    wire n2654;
    wire n2657;
    wire n2660;
    wire n2663;
    wire n2666;
    wire n2669;
    wire n2672;
    wire n2675;
    wire n2678;
    wire n2681;
    wire n2685;
    wire n2688;
    wire n2691;
    wire n2694;
    wire n2697;
    wire n2700;
    wire n2703;
    wire n2706;
    wire n2709;
    wire n2712;
    wire n2715;
    wire n2718;
    wire n2721;
    wire n2724;
    wire n2727;
    wire n2730;
    wire n2733;
    wire n2736;
    wire n2739;
    wire n2741;
    wire n2744;
    wire n2747;
    wire n2750;
    wire n2753;
    wire n2756;
    wire n2759;
    wire n2762;
    wire n2765;
    wire n2768;
    wire n2771;
    wire n2774;
    wire n2777;
    wire n2780;
    wire n2783;
    wire n2786;
    wire n2789;
    wire n2792;
    wire n2795;
    wire n2798;
    wire n2801;
    wire n2804;
    wire n2807;
    wire n2810;
    wire n2813;
    wire n2816;
    wire n2819;
    wire n2822;
    wire n2826;
    wire n2829;
    wire n2832;
    wire n2835;
    wire n2838;
    wire n2841;
    wire n2844;
    wire n2847;
    wire n2849;
    wire n2852;
    wire n2855;
    wire n2858;
    wire n2861;
    wire n2864;
    wire n2867;
    wire n2870;
    wire n2873;
    wire n2876;
    wire n2879;
    wire n2882;
    wire n2885;
    wire n2888;
    wire n2891;
    wire n2894;
    wire n2897;
    wire n2900;
    wire n2903;
    wire n2906;
    wire n2910;
    wire n2913;
    wire n2916;
    wire n2919;
    wire n2922;
    wire n2925;
    wire n2928;
    wire n2931;
    wire n2934;
    wire n2937;
    wire n2940;
    wire n2943;
    wire n2946;
    wire n2949;
    wire n2952;
    wire n2955;
    wire n2958;
    wire n2961;
    wire n2964;
    wire n2967;
    wire n2970;
    wire n2973;
    wire n2976;
    wire n2979;
    wire n2982;
    wire n2985;
    wire n2988;
    wire n2991;
    wire n2994;
    wire n2997;
    wire n3000;
    wire n3003;
    wire n3006;
    wire n3009;
    wire n3012;
    wire n3015;
    wire n3018;
    wire n3021;
    wire n3024;
    wire n3027;
    wire n3030;
    wire n3033;
    wire n3036;
    wire n3039;
    wire n3042;
    wire n3045;
    wire n3048;
    wire n3051;
    wire n3054;
    wire n3057;
    wire n3059;
    wire n3062;
    wire n3065;
    wire n3068;
    wire n3071;
    wire n3074;
    wire n3077;
    wire n3080;
    wire n3083;
    wire n3086;
    wire n3089;
    wire n3092;
    wire n3095;
    wire n3098;
    wire n3101;
    wire n3104;
    wire n3107;
    wire n3110;
    wire n3113;
    wire n3116;
    wire n3119;
    wire n3122;
    wire n3125;
    wire n3128;
    wire n3131;
    wire n3134;
    wire n3137;
    wire n3140;
    wire n3143;
    wire n3146;
    wire n3149;
    wire n3152;
    wire n3155;
    wire n3158;
    wire n3161;
    wire n3164;
    wire n3167;
    wire n3170;
    wire n3173;
    wire n3176;
    wire n3179;
    wire n3183;
    wire n3186;
    wire n3189;
    wire n3192;
    wire n3195;
    wire n3198;
    wire n3201;
    wire n3204;
    wire n3207;
    wire n3210;
    wire n3213;
    wire n3216;
    wire n3219;
    wire n3221;
    wire n3224;
    wire n3227;
    wire n3230;
    wire n3233;
    wire n3236;
    wire n3239;
    wire n3242;
    wire n3245;
    wire n3248;
    wire n3251;
    wire n3254;
    wire n3257;
    wire n3260;
    wire n3264;
    wire n3267;
    wire n3270;
    wire n3273;
    wire n3276;
    wire n3279;
    wire n3282;
    wire n3285;
    wire n3287;
    wire n3290;
    wire n3293;
    wire n3296;
    wire n3299;
    wire n3302;
    wire n3305;
    wire n3308;
    wire n3311;
    wire n3314;
    wire n3317;
    wire n3320;
    wire n3323;
    wire n3326;
    wire n3329;
    wire n3332;
    wire n3335;
    wire n3338;
    wire n3341;
    wire n3344;
    wire n3348;
    wire n3351;
    wire n3354;
    wire n3357;
    wire n3360;
    wire n3363;
    wire n3366;
    wire n3369;
    wire n3372;
    wire n3375;
    wire n3378;
    wire n3381;
    wire n3384;
    wire n3387;
    wire n3390;
    wire n3393;
    wire n3396;
    wire n3399;
    wire n3402;
    wire n3405;
    wire n3408;
    wire n3411;
    wire n3414;
    wire n3417;
    wire n3420;
    wire n3423;
    wire n3426;
    wire n3429;
    wire n3432;
    wire n3435;
    wire n3438;
    wire n3441;
    wire n3444;
    wire n3447;
    wire n3450;
    wire n3453;
    wire n3456;
    wire n3459;
    wire n3462;
    wire n3465;
    wire n3468;
    wire n3471;
    wire n3473;
    wire n3476;
    wire n3479;
    wire n3482;
    wire n3485;
    wire n3488;
    wire n3491;
    wire n3494;
    wire n3497;
    wire n3500;
    wire n3503;
    wire n3506;
    wire n3509;
    wire n3512;
    wire n3515;
    wire n3518;
    wire n3521;
    wire n3524;
    wire n3527;
    wire n3530;
    wire n3533;
    wire n3536;
    wire n3539;
    wire n3542;
    wire n3545;
    wire n3548;
    wire n3551;
    wire n3554;
    wire n3557;
    wire n3560;
    wire n3563;
    wire n3566;
    wire n3569;
    wire n3572;
    wire n3575;
    wire n3578;
    wire n3581;
    wire n3584;
    wire n3587;
    wire n3591;
    wire n3594;
    wire n3597;
    wire n3600;
    wire n3603;
    wire n3606;
    wire n3609;
    wire n3612;
    wire n3615;
    wire n3618;
    wire n3621;
    wire n3624;
    wire n3627;
    wire n3629;
    wire n3632;
    wire n3635;
    wire n3638;
    wire n3641;
    wire n3644;
    wire n3647;
    wire n3650;
    wire n3653;
    wire n3656;
    wire n3659;
    wire n3662;
    wire n3665;
    wire n3668;
    wire n3671;
    wire n3674;
    wire n3677;
    wire n3680;
    wire n3684;
    wire n3687;
    wire n3690;
    wire n3693;
    wire n3696;
    wire n3698;
    wire n3701;
    wire n3704;
    wire n3707;
    wire n3710;
    wire n3713;
    wire n3716;
    wire n3719;
    wire n3722;
    wire n3725;
    wire n3728;
    wire n3731;
    wire n3734;
    wire n3737;
    wire n3740;
    wire n3743;
    wire n3746;
    wire n3749;
    wire n3752;
    wire n3755;
    wire n3759;
    wire n3762;
    wire n3765;
    wire n3768;
    wire n3771;
    wire n3774;
    wire n3777;
    wire n3780;
    wire n3783;
    wire n3786;
    wire n3789;
    wire n3792;
    wire n3795;
    wire n3798;
    wire n3801;
    wire n3804;
    wire n3807;
    wire n3810;
    wire n3813;
    wire n3816;
    wire n3819;
    wire n3822;
    wire n3825;
    wire n3827;
    wire n3830;
    wire n3833;
    wire n3836;
    wire n3839;
    wire n3842;
    wire n3845;
    wire n3848;
    wire n3851;
    wire n3854;
    wire n3857;
    wire n3860;
    wire n3863;
    wire n3866;
    wire n3869;
    wire n3872;
    wire n3876;
    wire n3879;
    wire n3882;
    wire n3885;
    wire n3888;
    wire n3891;
    wire n3894;
    wire n3897;
    wire n3900;
    wire n3903;
    wire n3906;
    wire n3909;
    wire n3912;
    wire n3915;
    wire n3918;
    wire n3921;
    wire n3924;
    wire n3927;
    wire n3930;
    wire n3933;
    wire n3936;
    wire n3939;
    wire n3942;
    wire n3945;
    wire n3948;
    wire n3951;
    wire n3954;
    wire n3957;
    wire n3960;
    wire n3963;
    wire n3966;
    wire n3969;
    wire n3972;
    wire n3975;
    wire n3978;
    wire n3981;
    wire n3984;
    wire n3987;
    wire n3990;
    wire n3993;
    wire n3996;
    wire n3999;
    wire n4002;
    wire n4005;
    wire n4008;
    wire n4011;
    wire n4014;
    wire n4017;
    wire n4020;
    wire n4023;
    wire n4025;
    wire n4029;
    wire n4032;
    wire n4035;
    wire n4038;
    wire n4041;
    wire n4044;
    wire n4047;
    wire n4050;
    wire n4053;
    wire n4055;
    wire n4058;
    wire n4061;
    wire n4064;
    wire n4067;
    wire n4070;
    wire n4073;
    wire n4076;
    wire n4079;
    wire n4082;
    wire n4085;
    wire n4088;
    wire n4091;
    wire n4094;
    wire n4097;
    wire n4100;
    wire n4103;
    wire n4106;
    wire n4109;
    wire n4112;
    wire n4115;
    wire n4119;
    wire n4122;
    wire n4125;
    wire n4128;
    wire n4131;
    wire n4134;
    wire n4137;
    wire n4140;
    wire n4143;
    wire n4146;
    wire n4149;
    wire n4152;
    wire n4154;
    wire n4157;
    wire n4160;
    wire n4163;
    wire n4166;
    wire n4169;
    wire n4173;
    wire n4176;
    wire n4179;
    wire n4182;
    wire n4185;
    wire n4188;
    wire n4191;
    wire n4194;
    wire n4196;
    wire n4199;
    wire n4202;
    wire n4205;
    wire n4208;
    wire n4211;
    wire n4214;
    wire n4217;
    wire n4220;
    wire n4223;
    wire n4226;
    wire n4229;
    wire n4232;
    wire n4235;
    wire n4238;
    wire n4241;
    wire n4244;
    wire n4247;
    wire n4250;
    wire n4253;
    wire n4256;
    wire n4259;
    wire n4262;
    wire n4265;
    wire n4268;
    wire n4271;
    wire n4274;
    wire n4277;
    wire n4280;
    wire n4283;
    wire n4286;
    wire n4289;
    wire n4292;
    wire n4295;
    wire n4298;
    wire n4301;
    wire n4304;
    wire n4307;
    wire n4310;
    wire n4313;
    wire n4316;
    wire n4319;
    wire n4322;
    wire n4325;
    wire n4328;
    wire n4331;
    wire n4334;
    wire n4337;
    wire n4340;
    wire n4343;
    wire n4346;
    wire n4349;
    wire n4352;
    wire n4355;
    wire n4358;
    wire n4361;
    wire n4364;
    wire n4367;
    wire n4370;
    wire n4373;
    wire n4376;
    wire n4379;
    wire n4382;
    wire n4385;
    wire n4388;
    wire n4391;
    wire n4394;
    wire n4397;
    wire n4400;
    wire n4403;
    wire n4406;
    wire n4409;
    wire n4412;
    wire n4415;
    wire n4418;
    wire n4421;
    wire n4424;
    wire n4427;
    wire n4431;
    wire n4434;
    wire n4437;
    wire n4440;
    wire n4442;
    wire n4445;
    wire n4448;
    wire n4451;
    wire n4454;
    wire n4457;
    wire n4460;
    wire n4463;
    wire n4466;
    wire n4469;
    wire n4472;
    wire n4475;
    wire n4478;
    wire n4481;
    wire n4484;
    wire n4487;
    wire n4490;
    wire n4493;
    wire n4496;
    wire n4499;
    wire n4502;
    wire n4505;
    wire n4508;
    wire n4511;
    wire n4515;
    wire n4518;
    wire n4521;
    wire n4524;
    wire n4527;
    wire n4530;
    wire n4533;
    wire n4536;
    wire n4538;
    wire n4541;
    wire n4544;
    wire n4547;
    wire n4550;
    wire n4553;
    wire n4556;
    wire n4559;
    wire n4562;
    wire n4565;
    wire n4568;
    wire n4571;
    wire n4575;
    wire n4578;
    wire n4581;
    wire n4584;
    wire n4586;
    wire n4589;
    wire n4592;
    wire n4595;
    wire n4598;
    wire n4601;
    wire n4604;
    wire n4607;
    wire n4610;
    wire n4613;
    wire n4616;
    wire n4619;
    wire n4622;
    wire n4625;
    wire n4628;
    wire n4631;
    wire n4634;
    wire n4637;
    wire n4640;
    wire n4643;
    wire n4646;
    wire n4649;
    wire n4652;
    wire n4656;
    wire n4659;
    wire n4662;
    wire n4665;
    wire n4668;
    wire n4671;
    wire n4674;
    wire n4677;
    wire n4680;
    wire n4682;
    wire n4685;
    wire n4688;
    wire n4691;
    wire n4694;
    wire n4697;
    wire n4700;
    wire n4703;
    wire n4706;
    wire n4710;
    wire n4713;
    wire n4716;
    wire n4719;
    wire n4722;
    wire n4724;
    wire n4727;
    wire n4730;
    wire n4733;
    wire n4736;
    wire n4739;
    wire n4742;
    wire n4745;
    wire n4748;
    wire n4751;
    wire n4754;
    wire n4757;
    wire n4760;
    wire n4763;
    wire n4766;
    wire n4769;
    wire n4772;
    wire n4775;
    wire n4778;
    wire n4781;
    wire n4784;
    wire n4787;
    wire n4790;
    wire n4793;
    wire n4796;
    wire n4799;
    wire n4802;
    wire n4805;
    wire n4808;
    wire n4811;
    wire n4814;
    wire n4817;
    wire n4820;
    wire n4823;
    wire n4826;
    wire n4829;
    wire n4832;
    wire n4836;
    wire n4839;
    wire n4842;
    wire n4844;
    wire n4847;
    wire n4850;
    wire n4853;
    wire n4856;
    wire n4859;
    wire n4862;
    wire n4865;
    wire n4868;
    wire n4871;
    wire n4874;
    wire n4877;
    wire n4880;
    wire n4883;
    wire n4886;
    wire n4890;
    wire n4893;
    wire n4896;
    wire n4899;
    wire n4902;
    wire n4905;
    wire n4908;
    wire n4911;
    wire n4914;
    wire n4917;
    wire n4920;
    wire n4922;
    wire n4925;
    wire n4928;
    wire n4931;
    wire n4934;
    wire n4937;
    wire n4940;
    wire n4943;
    wire n4946;
    wire n4949;
    wire n4952;
    wire n4955;
    wire n4958;
    wire n4961;
    wire n4964;
    wire n4967;
    wire n4970;
    wire n4974;
    wire n4977;
    wire n4980;
    wire n4983;
    wire n4986;
    wire n4989;
    wire n4992;
    wire n4995;
    wire n4998;
    wire n5001;
    wire n5004;
    wire n5007;
    wire n5010;
    wire n5013;
    wire n5015;
    wire n5019;
    wire n5022;
    wire n5025;
    wire n5028;
    wire n5030;
    wire n5034;
    wire n5037;
    wire n5039;
    wire n5042;
    wire n5046;
    wire n5048;
    wire n5051;
    wire n5054;
    wire n5057;
    wire n5060;
    wire n5063;
    wire n5066;
    wire n5069;
    wire n5072;
    wire n5075;
    wire n5078;
    wire n5081;
    wire n5084;
    wire n5087;
    wire n5090;
    wire n5093;
    wire n5096;
    wire n5099;
    wire n5102;
    wire n5105;
    wire n5108;
    wire n5111;
    wire n5114;
    wire n5117;
    wire n5120;
    wire n5123;
    wire n5126;
    wire n5129;
    wire n5132;
    wire n5135;
    wire n5138;
    wire n5141;
    wire n5144;
    wire n5147;
    wire n5150;
    wire n5153;
    wire n5156;
    wire n5159;
    wire n5163;
    wire n5166;
    wire n5169;
    wire n5172;
    wire n5174;
    wire n5177;
    wire n5180;
    wire n5183;
    wire n5186;
    wire n5189;
    wire n5192;
    wire n5195;
    wire n5198;
    wire n5201;
    wire n5204;
    wire n5207;
    wire n5210;
    wire n5213;
    wire n5216;
    wire n5219;
    wire n5222;
    wire n5225;
    wire n5228;
    wire n5231;
    wire n5234;
    wire n5237;
    wire n5240;
    wire n5243;
    wire n5247;
    wire n5249;
    wire n5252;
    wire n5255;
    wire n5258;
    wire n5261;
    wire n5264;
    wire n5267;
    wire n5270;
    wire n5273;
    wire n5276;
    wire n5279;
    wire n5282;
    wire n5285;
    wire n5288;
    wire n5291;
    wire n5294;
    wire n5297;
    wire n5300;
    wire n5304;
    wire n5307;
    wire n5309;
    wire n5312;
    wire n5315;
    wire n5318;
    wire n5321;
    wire n5324;
    wire n5327;
    wire n5330;
    wire n5333;
    wire n5336;
    wire n5339;
    wire n5342;
    wire n5345;
    wire n5348;
    wire n5351;
    wire n5354;
    wire n5357;
    wire n5360;
    wire n5363;
    wire n5366;
    wire n5369;
    wire n5372;
    wire n5375;
    wire n5378;
    wire n5381;
    wire n5384;
    wire n5387;
    wire n5390;
    wire n5393;
    wire n5396;
    wire n5399;
    wire n5402;
    wire n5405;
    wire n5408;
    wire n5411;
    wire n5414;
    wire n5417;
    wire n5420;
    wire n5423;
    wire n5426;
    wire n5429;
    wire n5432;
    wire n5435;
    wire n5438;
    wire n5441;
    wire n5447;
    wire n5450;
    wire n5453;
    wire n5456;
    wire n5459;
    wire n5462;
    wire n5465;
    wire n5468;
    wire n5471;
    wire n5474;
    wire n5477;
    wire n5480;
    wire n5483;
    wire n5486;
    wire n5489;
    wire n5492;
    wire n5495;
    wire n5498;
    wire n5501;
    wire n5504;
    wire n5507;
    wire n5510;
    wire n5513;
    wire n5516;
    wire n5519;
    wire n5525;
    wire n5528;
    wire n5531;
    wire n5534;
    wire n5537;
    wire n5540;
    wire n5543;
    wire n5546;
    wire n5549;
    wire n5552;
    wire n5555;
    wire n5558;
    wire n5561;
    wire n5564;
    wire n5567;
    wire n5570;
    wire n5573;
    wire n5576;
    wire n5579;
    wire n5582;
    wire n5585;
    wire n5588;
    wire n5591;
    wire n5594;
    wire n5597;
    wire n5603;
    wire n5606;
    wire n5609;
    wire n5612;
    wire n5615;
    wire n5618;
    wire n5621;
    wire n5624;
    wire n5627;
    wire n5630;
    wire n5633;
    wire n5636;
    wire n5639;
    wire n5642;
    wire n5645;
    wire n5648;
    wire n5651;
    wire n5654;
    wire n5657;
    wire n5660;
    wire n5663;
    wire n5666;
    wire n5669;
    wire n5672;
    wire n5675;
    wire n5678;
    wire n5684;
    wire n5687;
    wire n5690;
    wire n5693;
    wire n5696;
    wire n5699;
    wire n5702;
    wire n5705;
    wire n5708;
    wire n5711;
    wire n5714;
    wire n5717;
    wire n5720;
    wire n5723;
    wire n5726;
    wire n5729;
    wire n5732;
    wire n5735;
    wire n5738;
    wire n5741;
    wire n5744;
    wire n5747;
    wire n5750;
    wire n5753;
    wire n5759;
    wire n5762;
    wire n5765;
    wire n5768;
    wire n5771;
    wire n5774;
    wire n5777;
    wire n5780;
    wire n5783;
    wire n5786;
    wire n5789;
    wire n5792;
    wire n5795;
    wire n5798;
    wire n5801;
    wire n5804;
    wire n5807;
    wire n5810;
    wire n5813;
    wire n5816;
    wire n5819;
    wire n5822;
    wire n5828;
    wire n5831;
    wire n5834;
    wire n5837;
    wire n5840;
    wire n5843;
    wire n5846;
    wire n5849;
    wire n5852;
    wire n5855;
    wire n5858;
    wire n5861;
    wire n5864;
    wire n5867;
    wire n5870;
    wire n5873;
    wire n5876;
    wire n5879;
    wire n5882;
    wire n5885;
    wire n5888;
    wire n5891;
    wire n5894;
    wire n5897;
    wire n5903;
    wire n5906;
    wire n5909;
    wire n5912;
    wire n5915;
    wire n5918;
    wire n5921;
    wire n5924;
    wire n5927;
    wire n5930;
    wire n5933;
    wire n5936;
    wire n5939;
    wire n5942;
    wire n5945;
    wire n5948;
    wire n5951;
    wire n5954;
    wire n5957;
    wire n5960;
    wire n5963;
    wire n5966;
    wire n5969;
    wire n5972;
    wire n5978;
    wire n5981;
    wire n5984;
    wire n5987;
    wire n5990;
    wire n5993;
    wire n5996;
    wire n5999;
    wire n6002;
    wire n6005;
    wire n6008;
    wire n6011;
    wire n6014;
    wire n6017;
    wire n6020;
    wire n6023;
    wire n6026;
    wire n6029;
    wire n6032;
    wire n6035;
    wire n6038;
    wire n6041;
    wire n6044;
    wire n6047;
    wire n6053;
    wire n6056;
    wire n6059;
    wire n6062;
    wire n6065;
    wire n6068;
    wire n6071;
    wire n6074;
    wire n6077;
    wire n6080;
    wire n6083;
    wire n6086;
    wire n6089;
    wire n6092;
    wire n6095;
    wire n6098;
    wire n6101;
    wire n6104;
    wire n6107;
    wire n6110;
    wire n6113;
    wire n6116;
    wire n6119;
    wire n6122;
    wire n6125;
    wire n6131;
    wire n6134;
    wire n6137;
    wire n6140;
    wire n6143;
    wire n6146;
    wire n6149;
    wire n6152;
    wire n6155;
    wire n6158;
    wire n6161;
    wire n6164;
    wire n6167;
    wire n6170;
    wire n6173;
    wire n6176;
    wire n6179;
    wire n6182;
    wire n6185;
    wire n6188;
    wire n6191;
    wire n6194;
    wire n6200;
    wire n6203;
    wire n6206;
    wire n6209;
    wire n6212;
    wire n6215;
    wire n6218;
    wire n6221;
    wire n6224;
    wire n6227;
    wire n6230;
    wire n6233;
    wire n6236;
    wire n6239;
    wire n6242;
    wire n6245;
    wire n6248;
    wire n6251;
    wire n6254;
    wire n6257;
    wire n6260;
    wire n6263;
    wire n6266;
    wire n6269;
    wire n6272;
    wire n6278;
    wire n6281;
    wire n6284;
    wire n6287;
    wire n6290;
    wire n6293;
    wire n6296;
    wire n6299;
    wire n6302;
    wire n6305;
    wire n6308;
    wire n6311;
    wire n6314;
    wire n6317;
    wire n6320;
    wire n6323;
    wire n6326;
    wire n6329;
    wire n6332;
    wire n6335;
    wire n6338;
    wire n6341;
    wire n6347;
    wire n6350;
    wire n6353;
    wire n6356;
    wire n6359;
    wire n6362;
    wire n6365;
    wire n6368;
    wire n6371;
    wire n6374;
    wire n6377;
    wire n6380;
    wire n6383;
    wire n6386;
    wire n6389;
    wire n6392;
    wire n6395;
    wire n6398;
    wire n6401;
    wire n6404;
    wire n6407;
    wire n6410;
    wire n6416;
    wire n6419;
    wire n6422;
    wire n6425;
    wire n6428;
    wire n6431;
    wire n6434;
    wire n6437;
    wire n6440;
    wire n6443;
    wire n6446;
    wire n6449;
    wire n6452;
    wire n6455;
    wire n6458;
    wire n6461;
    wire n6464;
    wire n6467;
    wire n6470;
    wire n6473;
    wire n6476;
    wire n6479;
    wire n6482;
    wire n6485;
    wire n6488;
    wire n6494;
    wire n6497;
    wire n6500;
    wire n6503;
    wire n6506;
    wire n6509;
    wire n6512;
    wire n6515;
    wire n6518;
    wire n6521;
    wire n6524;
    wire n6527;
    wire n6530;
    wire n6533;
    wire n6536;
    wire n6539;
    wire n6542;
    wire n6545;
    wire n6548;
    wire n6551;
    wire n6554;
    wire n6557;
    wire n6560;
    wire n6566;
    wire n6569;
    wire n6572;
    wire n6575;
    wire n6578;
    wire n6581;
    wire n6584;
    wire n6587;
    wire n6590;
    wire n6593;
    wire n6596;
    wire n6599;
    wire n6602;
    wire n6605;
    wire n6608;
    wire n6611;
    wire n6614;
    wire n6617;
    wire n6620;
    wire n6623;
    wire n6626;
    wire n6629;
    wire n6632;
    wire n6638;
    wire n6641;
    wire n6644;
    wire n6647;
    wire n6650;
    wire n6653;
    wire n6656;
    wire n6659;
    wire n6662;
    wire n6665;
    wire n6668;
    wire n6671;
    wire n6677;
    wire n6680;
    wire n6683;
    wire n6686;
    wire n6689;
    wire n6692;
    wire n6695;
    wire n6701;
    wire n6704;
    wire n6707;
    wire n6710;
    wire n6713;
    wire n6716;
    wire n6719;
    wire n6722;
    wire n6725;
    wire n6731;
    wire n6734;
    wire n6737;
    wire n6740;
    wire n6743;
    wire n6746;
    wire n6749;
    wire n6752;
    wire n6755;
    wire n6758;
    wire n6761;
    wire n6767;
    wire n6773;
    wire n6776;
    wire n6779;
    wire n6782;
    wire n6788;
    wire n6794;
    wire n6797;
    wire n6800;
    jand g000(.dinb(G29gat), .dina(G75gat), .dout(n89));
    jand g001(.dinb(n5270), .dina(n89), .dout(n93));
    jand g002(.dinb(G29gat), .dina(G36gat), .dout(n97));
    jand g003(.dinb(n5123), .dina(n97), .dout(n101));
    jand g004(.dinb(n5270), .dina(n97), .dout(n105));
    jand g005(.dinb(G85gat), .dina(G86gat), .dout(n109));
    jand g006(.dinb(G1gat), .dina(G8gat), .dout(n113));
    jand g007(.dinb(n5291), .dina(n113), .dout(n117));
    jand g008(.dinb(n5075), .dina(n117), .dout(n121));
    jnot g009(.din(G17gat), .dout(n124));
    jnot g010(.din(G13gat), .dout(n127));
    jnot g011(.din(G1gat), .dout(n130));
    jnot g012(.din(G26gat), .dout(n133));
    jor g013(.dinb(n130), .dina(n133), .dout(n137));
    jor g014(.dinb(n2052), .dina(n137), .dout(n141));
    jor g015(.dinb(n5069), .dina(n141), .dout(n145));
    jor g016(.dinb(n2054), .dina(n145), .dout(n149));
    jnot g017(.din(G80gat), .dout(n152));
    jand g018(.dinb(G59gat), .dina(G75gat), .dout(n156));
    jnot g019(.din(n156), .dout(n159));
    jor g020(.dinb(n2043), .dina(n159), .dout(n163));
    jnot g021(.din(G36gat), .dout(n166));
    jnot g022(.din(G59gat), .dout(n169));
    jor g023(.dinb(n166), .dina(n169), .dout(n173));
    jor g024(.dinb(n2043), .dina(n173), .dout(n177));
    jnot g025(.din(G42gat), .dout(n180));
    jor g026(.dinb(n5054), .dina(n173), .dout(n184));
    jor g027(.dinb(G87gat), .dina(G88gat), .dout(n188));
    jand g028(.dinb(n2046), .dina(n188), .dout(n192));
    jnot g029(.din(n105), .dout(n195));
    jor g030(.dinb(n2049), .dina(n145), .dout(n199));
    jand g031(.dinb(G1gat), .dina(G26gat), .dout(n203));
    jand g032(.dinb(n5114), .dina(n203), .dout(n207));
    jand g033(.dinb(n5307), .dina(n117), .dout(n211));
    jand g034(.dinb(n5132), .dina(n211), .dout(n215));
    jand g035(.dinb(n5258), .dina(n215), .dout(n219));
    jand g036(.dinb(G59gat), .dina(G68gat), .dout(n223));
    jand g037(.dinb(n2067), .dina(n211), .dout(n227));
    jand g038(.dinb(n5249), .dina(n227), .dout(n231));
    jand g039(.dinb(n2070), .dina(n188), .dout(n235));
    jxor g040(.dinb(G111gat), .dina(G116gat), .dout(n239));
    jxor g041(.dinb(n2076), .dina(n239), .dout(n243));
    jxor g042(.dinb(G91gat), .dina(G96gat), .dout(n247));
    jxor g043(.dinb(n2081), .dina(n247), .dout(n251));
    jxor g044(.dinb(G101gat), .dina(G106gat), .dout(n255));
    jxor g045(.dinb(G121gat), .dina(G126gat), .dout(n259));
    jxor g046(.dinb(n255), .dina(n259), .dout(n263));
    jxor g047(.dinb(n251), .dina(n263), .dout(n267));
    jxor g048(.dinb(n2073), .dina(n267), .dout(n271));
    jxor g049(.dinb(G183gat), .dina(G189gat), .dout(n275));
    jxor g050(.dinb(n2085), .dina(n275), .dout(n279));
    jxor g051(.dinb(G130gat), .dina(G159gat), .dout(n283));
    jxor g052(.dinb(n3759), .dina(n283), .dout(n287));
    jxor g053(.dinb(G171gat), .dina(G177gat), .dout(n291));
    jxor g054(.dinb(G195gat), .dina(G201gat), .dout(n295));
    jxor g055(.dinb(n291), .dina(n295), .dout(n299));
    jxor g056(.dinb(n287), .dina(n299), .dout(n303));
    jxor g057(.dinb(n2079), .dina(n303), .dout(n307));
    jnot g058(.din(G268gat), .dout(n310));
    jand g059(.dinb(n5117), .dina(n207), .dout(n314));
    jand g060(.dinb(n5126), .dina(n314), .dout(n318));
    jand g061(.dinb(n5297), .dina(n318), .dout(n322));
    jand g062(.dinb(n5172), .dina(n322), .dout(n326));
    jand g063(.dinb(n124), .dina(n180), .dout(n330));
    jnot g064(.din(n330), .dout(n333));
    jand g065(.dinb(G59gat), .dina(G156gat), .dout(n337));
    jand g066(.dinb(G17gat), .dina(G42gat), .dout(n341));
    jnot g067(.din(n341), .dout(n344));
    jand g068(.dinb(n5046), .dina(n344), .dout(n348));
    jand g069(.dinb(n5111), .dina(n348), .dout(n352));
    jand g070(.dinb(n5037), .dina(n352), .dout(n356));
    jnot g071(.din(n113), .dout(n359));
    jand g072(.dinb(n5057), .dina(n156), .dout(n363));
    jand g073(.dinb(G17gat), .dina(G51gat), .dout(n367));
    jnot g074(.din(n367), .dout(n370));
    jor g075(.dinb(n363), .dina(n370), .dout(n374));
    jor g076(.dinb(n5034), .dina(n374), .dout(n378));
    jnot g077(.din(n378), .dout(n381));
    jor g078(.dinb(n356), .dina(n381), .dout(n385));
    jand g079(.dinb(n4154), .dina(n385), .dout(n389));
    jnot g080(.din(G156gat), .dout(n392));
    jor g081(.dinb(n169), .dina(n392), .dout(n396));
    jand g082(.dinb(n207), .dina(n396), .dout(n400));
    jand g083(.dinb(n5153), .dina(n400), .dout(n404));
    jor g084(.dinb(n4562), .dina(n404), .dout(n408));
    jand g085(.dinb(n4736), .dina(n408), .dout(n412));
    jor g086(.dinb(n389), .dina(n3825), .dout(n416));
    jor g087(.dinb(n4586), .dina(n416), .dout(n420));
    jand g088(.dinb(n2243), .dina(n420), .dout(n424));
    jand g089(.dinb(n5273), .dina(n223), .dout(n428));
    jand g090(.dinb(G72gat), .dina(G73gat), .dout(n432));
    jand g091(.dinb(n428), .dina(n5247), .dout(n436));
    jand g092(.dinb(n211), .dina(n436), .dout(n440));
    jand g093(.dinb(n2144), .dina(n440), .dout(n444));
    jor g094(.dinb(n424), .dina(n2142), .dout(n448));
    jnot g095(.din(G201gat), .dout(n451));
    jnot g096(.din(n326), .dout(n454));
    jnot g097(.din(G126gat), .dout(n457));
    jnot g098(.din(G51gat), .dout(n460));
    jor g099(.dinb(n4152), .dina(n137), .dout(n464));
    jor g100(.dinb(n396), .dina(n5039), .dout(n468));
    jor g101(.dinb(n464), .dina(n468), .dout(n472));
    jor g102(.dinb(n5048), .dina(n472), .dout(n476));
    jand g103(.dinb(n476), .dina(n5030), .dout(n480));
    jor g104(.dinb(n4149), .dina(n480), .dout(n484));
    jnot g105(.din(G153gat), .dout(n487));
    jor g106(.dinb(n464), .dina(n5042), .dout(n491));
    jor g107(.dinb(n5060), .dina(n491), .dout(n495));
    jand g108(.dinb(n5276), .dina(n495), .dout(n499));
    jor g109(.dinb(n4134), .dina(n499), .dout(n503));
    jand g110(.dinb(n484), .dina(n503), .dout(n507));
    jand g111(.dinb(n4119), .dina(n507), .dout(n511));
    jxor g112(.dinb(n4194), .dina(n511), .dout(n515));
    jand g113(.dinb(n2306), .dina(n515), .dout(n519));
    jand g114(.dinb(n4196), .dina(n420), .dout(n523));
    jand g115(.dinb(n2246), .dina(n523), .dout(n527));
    jand g116(.dinb(G121gat), .dina(G210gat), .dout(n531));
    jand g117(.dinb(G255gat), .dina(G267gat), .dout(n535));
    jor g118(.dinb(n531), .dina(n535), .dout(n539));
    jor g119(.dinb(n527), .dina(n2127), .dout(n543));
    jor g120(.dinb(n2100), .dina(n543), .dout(n547));
    jor g121(.dinb(n2097), .dina(n547), .dout(n551));
    jor g122(.dinb(n4085), .dina(n515), .dout(n555));
    jnot g123(.din(G261gat), .dout(n558));
    jnot g124(.din(n515), .dout(n561));
    jor g125(.dinb(n4025), .dina(n561), .dout(n565));
    jand g126(.dinb(n3909), .dina(n565), .dout(n569));
    jand g127(.dinb(n2091), .dina(n569), .dout(n573));
    jor g128(.dinb(n551), .dina(n573), .dout(n577));
    jand g129(.dinb(n4592), .dina(n385), .dout(n581));
    jand g130(.dinb(n4571), .dina(n408), .dout(n585));
    jor g131(.dinb(n326), .dina(n585), .dout(n589));
    jor g132(.dinb(n581), .dina(n589), .dout(n593));
    jxor g133(.dinb(n2282), .dina(n593), .dout(n597));
    jand g134(.dinb(n4998), .dina(n597), .dout(n601));
    jand g135(.dinb(n2270), .dina(n440), .dout(n605));
    jand g136(.dinb(n4610), .dina(n593), .dout(n609));
    jand g137(.dinb(n5201), .dina(n609), .dout(n613));
    jand g138(.dinb(n4868), .dina(n593), .dout(n617));
    jand g139(.dinb(G106gat), .dina(G210gat), .dout(n621));
    jor g140(.dinb(n617), .dina(n2241), .dout(n625));
    jor g141(.dinb(n613), .dina(n625), .dout(n629));
    jor g142(.dinb(n2217), .dina(n629), .dout(n633));
    jor g143(.dinb(n2199), .dina(n633), .dout(n637));
    jand g144(.dinb(n4442), .dina(n385), .dout(n641));
    jand g145(.dinb(n4427), .dina(n408), .dout(n645));
    jor g146(.dinb(n326), .dina(n645), .dout(n649));
    jor g147(.dinb(n641), .dina(n649), .dout(n653));
    jand g148(.dinb(n4460), .dina(n653), .dout(n657));
    jor g149(.dinb(n4385), .dina(n653), .dout(n661));
    jand g150(.dinb(n4292), .dina(n385), .dout(n665));
    jand g151(.dinb(n5015), .dina(n408), .dout(n669));
    jor g152(.dinb(n326), .dina(n669), .dout(n673));
    jor g153(.dinb(n665), .dina(n673), .dout(n677));
    jand g154(.dinb(n4310), .dina(n677), .dout(n681));
    jor g155(.dinb(n4256), .dina(n677), .dout(n685));
    jand g156(.dinb(n4194), .dina(n511), .dout(n689));
    jnot g157(.din(n689), .dout(n692));
    jor g158(.dinb(n4055), .dina(n523), .dout(n696));
    jand g159(.dinb(n692), .dina(n696), .dout(n700));
    jand g160(.dinb(n4223), .dina(n700), .dout(n704));
    jor g161(.dinb(n4280), .dina(n704), .dout(n708));
    jand g162(.dinb(n4346), .dina(n708), .dout(n712));
    jor g163(.dinb(n4409), .dina(n712), .dout(n716));
    jor g164(.dinb(n2249), .dina(n716), .dout(n720));
    jnot g165(.din(n597), .dout(n723));
    jnot g166(.din(n657), .dout(n726));
    jnot g167(.din(n661), .dout(n729));
    jnot g168(.din(n681), .dout(n732));
    jnot g169(.din(n685), .dout(n735));
    jor g170(.dinb(n4194), .dina(n511), .dout(n739));
    jand g171(.dinb(n4053), .dina(n739), .dout(n743));
    jor g172(.dinb(n4115), .dina(n743), .dout(n747));
    jor g173(.dinb(n4023), .dina(n747), .dout(n751));
    jand g174(.dinb(n4017), .dina(n751), .dout(n755));
    jor g175(.dinb(n4008), .dina(n755), .dout(n759));
    jand g176(.dinb(n3996), .dina(n759), .dout(n763));
    jor g177(.dinb(n2193), .dina(n763), .dout(n767));
    jand g178(.dinb(n2348), .dina(n767), .dout(n771));
    jand g179(.dinb(n2175), .dina(n771), .dout(n775));
    jor g180(.dinb(n2172), .dina(n775), .dout(n779));
    jxor g181(.dinb(n4361), .dina(n653), .dout(n783));
    jand g182(.dinb(n4998), .dina(n783), .dout(n787));
    jand g183(.dinb(G111gat), .dina(G210gat), .dout(n791));
    jand g184(.dinb(G189gat), .dina(G237gat), .dout(n795));
    jor g185(.dinb(n4890), .dina(n795), .dout(n799));
    jand g186(.dinb(n653), .dina(n2430), .dout(n803));
    jor g187(.dinb(n2412), .dina(n803), .dout(n807));
    jand g188(.dinb(G255gat), .dina(G259gat), .dout(n811));
    jand g189(.dinb(n4484), .dina(n440), .dout(n815));
    jor g190(.dinb(n2388), .dina(n815), .dout(n819));
    jor g191(.dinb(n807), .dina(n2376), .dout(n823));
    jor g192(.dinb(n2364), .dina(n823), .dout(n827));
    jor g193(.dinb(n708), .dina(n2432), .dout(n831));
    jnot g194(.din(n783), .dout(n834));
    jor g195(.dinb(n755), .dina(n2337), .dout(n838));
    jand g196(.dinb(n2339), .dina(n838), .dout(n842));
    jand g197(.dinb(n2325), .dina(n842), .dout(n846));
    jor g198(.dinb(n2322), .dina(n846), .dout(n850));
    jxor g199(.dinb(n4232), .dina(n677), .dout(n854));
    jand g200(.dinb(n4998), .dina(n854), .dout(n858));
    jand g201(.dinb(G116gat), .dina(G210gat), .dout(n862));
    jand g202(.dinb(G195gat), .dina(G237gat), .dout(n866));
    jor g203(.dinb(n4890), .dina(n866), .dout(n870));
    jand g204(.dinb(n677), .dina(n2532), .dout(n874));
    jor g205(.dinb(n2514), .dina(n874), .dout(n878));
    jand g206(.dinb(n4334), .dina(n440), .dout(n882));
    jand g207(.dinb(G255gat), .dina(G260gat), .dout(n886));
    jor g208(.dinb(n882), .dina(n2490), .dout(n890));
    jor g209(.dinb(n878), .dina(n2478), .dout(n894));
    jor g210(.dinb(n2466), .dina(n894), .dout(n898));
    jor g211(.dinb(n700), .dina(n2534), .dout(n902));
    jnot g212(.din(n854), .dout(n905));
    jor g213(.dinb(n747), .dina(n2463), .dout(n909));
    jand g214(.dinb(n3872), .dina(n909), .dout(n913));
    jand g215(.dinb(n2457), .dina(n913), .dout(n917));
    jor g216(.dinb(n2454), .dina(n917), .dout(n921));
    jand g217(.dinb(n5294), .dina(n400), .dout(n925));
    jand g218(.dinb(n4584), .dina(n925), .dout(n929));
    jand g219(.dinb(n5141), .dina(n318), .dout(n933));
    jand g220(.dinb(n5172), .dina(n933), .dout(n937));
    jor g221(.dinb(n3285), .dina(n937), .dout(n941));
    jand g222(.dinb(n3629), .dina(n385), .dout(n945));
    jand g223(.dinb(G8gat), .dina(G138gat), .dout(n949));
    jor g224(.dinb(n945), .dina(n3282), .dout(n953));
    jor g225(.dinb(n3264), .dina(n953), .dout(n957));
    jand g226(.dinb(n2657), .dina(n957), .dout(n961));
    jor g227(.dinb(n2630), .dina(n957), .dout(n965));
    jand g228(.dinb(n4922), .dina(n385), .dout(n969));
    jand g229(.dinb(n4440), .dina(n925), .dout(n973));
    jand g230(.dinb(G51gat), .dina(G138gat), .dout(n977));
    jor g231(.dinb(n973), .dina(n3696), .dout(n981));
    jor g232(.dinb(n969), .dina(n3684), .dout(n985));
    jor g233(.dinb(n3698), .dina(n985), .dout(n989));
    jand g234(.dinb(n3158), .dina(n989), .dout(n993));
    jor g235(.dinb(n3134), .dina(n989), .dout(n997));
    jand g236(.dinb(n5081), .dina(n385), .dout(n1001));
    jand g237(.dinb(n5028), .dina(n925), .dout(n1005));
    jand g238(.dinb(G17gat), .dina(G138gat), .dout(n1009));
    jor g239(.dinb(n1005), .dina(n5013), .dout(n1013));
    jor g240(.dinb(n1001), .dina(n5001), .dout(n1017));
    jor g241(.dinb(n5105), .dina(n1017), .dout(n1021));
    jand g242(.dinb(n3563), .dina(n1021), .dout(n1025));
    jor g243(.dinb(n3536), .dina(n1021), .dout(n1029));
    jand g244(.dinb(n4751), .dina(n385), .dout(n1033));
    jand g245(.dinb(n4724), .dina(n925), .dout(n1037));
    jand g246(.dinb(G138gat), .dina(G152gat), .dout(n1041));
    jor g247(.dinb(n1037), .dina(n4722), .dout(n1045));
    jor g248(.dinb(n1033), .dina(n4710), .dout(n1049));
    jor g249(.dinb(n5099), .dina(n1049), .dout(n1053));
    jand g250(.dinb(n4769), .dina(n1053), .dout(n1057));
    jnot g251(.din(G177gat), .dout(n1060));
    jnot g252(.din(n1053), .dout(n1063));
    jand g253(.dinb(n4680), .dina(n1063), .dout(n1067));
    jnot g254(.din(n1067), .dout(n1070));
    jnot g255(.din(G183gat), .dout(n1073));
    jnot g256(.din(n593), .dout(n1076));
    jand g257(.dinb(n4536), .dina(n1076), .dout(n1080));
    jnot g258(.din(n1080), .dout(n1083));
    jand g259(.dinb(n3822), .dina(n716), .dout(n1087));
    jor g260(.dinb(n4538), .dina(n1087), .dout(n1091));
    jand g261(.dinb(n3807), .dina(n1091), .dout(n1095));
    jor g262(.dinb(n4682), .dina(n1095), .dout(n1099));
    jand g263(.dinb(n3473), .dina(n1099), .dout(n1103));
    jor g264(.dinb(n3503), .dina(n1103), .dout(n1107));
    jand g265(.dinb(n3059), .dina(n1107), .dout(n1111));
    jor g266(.dinb(n3095), .dina(n1111), .dout(n1115));
    jand g267(.dinb(n2628), .dina(n1115), .dout(n1119));
    jor g268(.dinb(n2586), .dina(n1119), .dout(n1123));
    jxor g269(.dinb(n4808), .dina(n1053), .dout(n1127));
    jnot g270(.din(n1127), .dout(n1130));
    jand g271(.dinb(n2864), .dina(n1091), .dout(n1134));
    jand g272(.dinb(n2847), .dina(n1134), .dout(n1138));
    jnot g273(.din(n609), .dout(n1141));
    jor g274(.dinb(n4496), .dina(n763), .dout(n1145));
    jand g275(.dinb(n3981), .dina(n1145), .dout(n1149));
    jand g276(.dinb(n2849), .dina(n1149), .dout(n1153));
    jor g277(.dinb(n2795), .dina(n1153), .dout(n1157));
    jand g278(.dinb(n2879), .dina(n1157), .dout(n1161));
    jand g279(.dinb(n2765), .dina(n1057), .dout(n1165));
    jand g280(.dinb(n2741), .dina(n1053), .dout(n1169));
    jand g281(.dinb(G101gat), .dina(G210gat), .dout(n1173));
    jand g282(.dinb(n4796), .dina(n440), .dout(n1177));
    jor g283(.dinb(n2739), .dina(n1177), .dout(n1181));
    jor g284(.dinb(n1169), .dina(n2727), .dout(n1185));
    jor g285(.dinb(n1165), .dina(n1185), .dout(n1189));
    jor g286(.dinb(n1161), .dina(n2715), .dout(n1193));
    jor g287(.dinb(n2688), .dina(n1193), .dout(n1197));
    jand g288(.dinb(n5174), .dina(n957), .dout(n1201));
    jor g289(.dinb(n5228), .dina(n1201), .dout(n1205));
    jand g290(.dinb(n3314), .dina(n1205), .dout(n1209));
    jxor g291(.dinb(n3287), .dina(n957), .dout(n1213));
    jand g292(.dinb(n4970), .dina(n1213), .dout(n1217));
    jand g293(.dinb(G210gat), .dina(G268gat), .dout(n1221));
    jor g294(.dinb(n1217), .dina(n3219), .dout(n1225));
    jand g295(.dinb(n4844), .dina(n957), .dout(n1229));
    jor g296(.dinb(n1225), .dina(n3189), .dout(n1233));
    jor g297(.dinb(n3183), .dina(n1233), .dout(n1237));
    jor g298(.dinb(n1115), .dina(n3221), .dout(n1241));
    jnot g299(.din(n993), .dout(n1244));
    jnot g300(.din(n997), .dout(n1247));
    jnot g301(.din(n1025), .dout(n1250));
    jnot g302(.din(n1029), .dout(n1253));
    jnot g303(.din(n1057), .dout(n1256));
    jor g304(.dinb(n4634), .dina(n1149), .dout(n1260));
    jand g305(.dinb(n3960), .dina(n1260), .dout(n1264));
    jor g306(.dinb(n3471), .dina(n1264), .dout(n1268));
    jand g307(.dinb(n3444), .dina(n1268), .dout(n1272));
    jor g308(.dinb(n3057), .dina(n1272), .dout(n1276));
    jand g309(.dinb(n3024), .dina(n1276), .dout(n1280));
    jnot g310(.din(n1213), .dout(n1283));
    jor g311(.dinb(n1280), .dina(n2988), .dout(n1287));
    jand g312(.dinb(n3833), .dina(n1287), .dout(n1291));
    jand g313(.dinb(n2949), .dina(n1291), .dout(n1295));
    jor g314(.dinb(n2946), .dina(n1295), .dout(G878gat));
    jand g315(.dinb(n5174), .dina(n989), .dout(n1303));
    jor g316(.dinb(n5228), .dina(n1303), .dout(n1307));
    jand g317(.dinb(n3728), .dina(n1307), .dout(n1311));
    jxor g318(.dinb(n3704), .dina(n989), .dout(n1315));
    jand g319(.dinb(n4970), .dina(n1315), .dout(n1319));
    jand g320(.dinb(G91gat), .dina(G210gat), .dout(n1323));
    jor g321(.dinb(n1319), .dina(n3627), .dout(n1327));
    jand g322(.dinb(n4844), .dina(n989), .dout(n1331));
    jor g323(.dinb(n1327), .dina(n3597), .dout(n1335));
    jor g324(.dinb(n3591), .dina(n1335), .dout(n1339));
    jor g325(.dinb(n1107), .dina(n3647), .dout(n1343));
    jnot g326(.din(n1315), .dout(n1346));
    jor g327(.dinb(n1272), .dina(n3414), .dout(n1350));
    jand g328(.dinb(n3827), .dina(n1350), .dout(n1354));
    jand g329(.dinb(n3381), .dina(n1354), .dout(n1358));
    jor g330(.dinb(n3378), .dina(n1358), .dout(n1362));
    jand g331(.dinb(n5174), .dina(n1021), .dout(n1366));
    jor g332(.dinb(n5228), .dina(n1366), .dout(n1370));
    jand g333(.dinb(n5336), .dina(n1370), .dout(n1374));
    jxor g334(.dinb(n5309), .dina(n1021), .dout(n1378));
    jand g335(.dinb(n4970), .dina(n1378), .dout(n1382));
    jand g336(.dinb(G96gat), .dina(G210gat), .dout(n1386));
    jor g337(.dinb(n1382), .dina(n4920), .dout(n1390));
    jand g338(.dinb(n4844), .dina(n1021), .dout(n1394));
    jor g339(.dinb(n1390), .dina(n4842), .dout(n1398));
    jor g340(.dinb(n4836), .dina(n1398), .dout(n1402));
    jnot g341(.din(n1378), .dout(n1405));
    jor g342(.dinb(n1264), .dina(n3936), .dout(n1409));
    jor g343(.dinb(n1099), .dina(n4940), .dout(n1413));
    jand g344(.dinb(n3845), .dina(n1413), .dout(n1417));
    jand g345(.dinb(n3789), .dina(n1417), .dout(n1421));
    jor g346(.dinb(n3786), .dina(n1421), .dout(n1425));
    jdff dff_A_RrvOc9bb9_0(.din(n6800), .dout(G880gat));
    jdff dff_A_ToHw2GrJ1_0(.din(n6797), .dout(n6800));
    jdff dff_A_hKsJVxjJ0_0(.din(n6794), .dout(n6797));
    jdff dff_A_yvuvlarN9_2(.din(n1425), .dout(n6794));
    jdff dff_A_peHDjjEc4_0(.din(n6788), .dout(G879gat));
    jdff dff_A_j2wVWtWp7_2(.din(n1362), .dout(n6788));
    jdff dff_A_k6q6b7sE7_0(.din(n6782), .dout(G874gat));
    jdff dff_A_t0q54zPC0_0(.din(n6779), .dout(n6782));
    jdff dff_A_Qci0cMBR4_0(.din(n6776), .dout(n6779));
    jdff dff_A_HlFeHme37_0(.din(n6773), .dout(n6776));
    jdff dff_A_59cdx3DS7_2(.din(n1197), .dout(n6773));
    jdff dff_A_TgbimvxW0_0(.din(n6767), .dout(G866gat));
    jdff dff_A_uu90gjxu6_2(.din(n1123), .dout(n6767));
    jdff dff_A_OWy0ZP7R1_0(.din(n6761), .dout(G865gat));
    jdff dff_A_vdT0ciDk9_0(.din(n6758), .dout(n6761));
    jdff dff_A_VdkCCeHd8_0(.din(n6755), .dout(n6758));
    jdff dff_A_OKY0dIbs7_0(.din(n6752), .dout(n6755));
    jdff dff_A_1sEohxXZ4_0(.din(n6749), .dout(n6752));
    jdff dff_A_IulKnn1f1_0(.din(n6746), .dout(n6749));
    jdff dff_A_UxxXG8wq0_0(.din(n6743), .dout(n6746));
    jdff dff_A_xvs9Erk25_0(.din(n6740), .dout(n6743));
    jdff dff_A_nAlhdSUP5_0(.din(n6737), .dout(n6740));
    jdff dff_A_T2UfIs6M5_0(.din(n6734), .dout(n6737));
    jdff dff_A_rvjWJORW9_0(.din(n6731), .dout(n6734));
    jdff dff_A_i7fpZ1qg5_2(.din(n921), .dout(n6731));
    jdff dff_A_a8gxr0EZ7_0(.din(n6725), .dout(G864gat));
    jdff dff_A_CZ2WFe3r6_0(.din(n6722), .dout(n6725));
    jdff dff_A_luZJ4B4N8_0(.din(n6719), .dout(n6722));
    jdff dff_A_8iMkopc76_0(.din(n6716), .dout(n6719));
    jdff dff_A_gWtLxFGp7_0(.din(n6713), .dout(n6716));
    jdff dff_A_pCjPIYbn1_0(.din(n6710), .dout(n6713));
    jdff dff_A_Kl7a5jAB0_0(.din(n6707), .dout(n6710));
    jdff dff_A_rihFLxqu4_0(.din(n6704), .dout(n6707));
    jdff dff_A_Yw8WOXeD3_0(.din(n6701), .dout(n6704));
    jdff dff_A_EaLwtXtj9_2(.din(n850), .dout(n6701));
    jdff dff_A_bfi6CDsu0_0(.din(n6695), .dout(G863gat));
    jdff dff_A_o0Ti0cIn1_0(.din(n6692), .dout(n6695));
    jdff dff_A_FIPprnkS9_0(.din(n6689), .dout(n6692));
    jdff dff_A_iJBFqXoD7_0(.din(n6686), .dout(n6689));
    jdff dff_A_tWQhGJB15_0(.din(n6683), .dout(n6686));
    jdff dff_A_rCvrwCWK4_0(.din(n6680), .dout(n6683));
    jdff dff_A_WifP3QV35_0(.din(n6677), .dout(n6680));
    jdff dff_A_kOlKxf7O4_2(.din(n779), .dout(n6677));
    jdff dff_A_z2UgFbIY1_0(.din(n6671), .dout(G850gat));
    jdff dff_A_zisxz3fN4_0(.din(n6668), .dout(n6671));
    jdff dff_A_Q8RntV027_0(.din(n6665), .dout(n6668));
    jdff dff_A_2TSW3xlc0_0(.din(n6662), .dout(n6665));
    jdff dff_A_SC86Nwwo5_0(.din(n6659), .dout(n6662));
    jdff dff_A_0sjJb1qh1_0(.din(n6656), .dout(n6659));
    jdff dff_A_RDyqs1ny6_0(.din(n6653), .dout(n6656));
    jdff dff_A_BjlvJ0cv9_0(.din(n6650), .dout(n6653));
    jdff dff_A_7AnUinVD1_0(.din(n6647), .dout(n6650));
    jdff dff_A_DDv9Ri6O3_0(.din(n6644), .dout(n6647));
    jdff dff_A_p3rjj3bx0_0(.din(n6641), .dout(n6644));
    jdff dff_A_FW3tNPOQ3_0(.din(n6638), .dout(n6641));
    jdff dff_A_0bei3kWP7_2(.din(n577), .dout(n6638));
    jdff dff_A_154bAPmV3_0(.din(n6632), .dout(G768gat));
    jdff dff_A_MyBrPLSD4_0(.din(n6629), .dout(n6632));
    jdff dff_A_ikFvfpAo1_0(.din(n6626), .dout(n6629));
    jdff dff_A_f6YJmiCl1_0(.din(n6623), .dout(n6626));
    jdff dff_A_Kankvch38_0(.din(n6620), .dout(n6623));
    jdff dff_A_1TKF6j2i2_0(.din(n6617), .dout(n6620));
    jdff dff_A_2vWaFgIl2_0(.din(n6614), .dout(n6617));
    jdff dff_A_uq1pQA367_0(.din(n6611), .dout(n6614));
    jdff dff_A_IJZegaBq5_0(.din(n6608), .dout(n6611));
    jdff dff_A_qRogF6Ix9_0(.din(n6605), .dout(n6608));
    jdff dff_A_rJVwUmKk0_0(.din(n6602), .dout(n6605));
    jdff dff_A_xqnlnMaR6_0(.din(n6599), .dout(n6602));
    jdff dff_A_DyDUDH0p4_0(.din(n6596), .dout(n6599));
    jdff dff_A_kFyR0jOj6_0(.din(n6593), .dout(n6596));
    jdff dff_A_M4Z4rDQt2_0(.din(n6590), .dout(n6593));
    jdff dff_A_xRYGPthN0_0(.din(n6587), .dout(n6590));
    jdff dff_A_R7Y3MG942_0(.din(n6584), .dout(n6587));
    jdff dff_A_pHqeztw50_0(.din(n6581), .dout(n6584));
    jdff dff_A_COMTXygF4_0(.din(n6578), .dout(n6581));
    jdff dff_A_0sGc09mi4_0(.din(n6575), .dout(n6578));
    jdff dff_A_rFqSc2Fp3_0(.din(n6572), .dout(n6575));
    jdff dff_A_4MHuud4Z4_0(.din(n6569), .dout(n6572));
    jdff dff_A_tfJCnvsX0_0(.din(n6566), .dout(n6569));
    jdff dff_A_kFURueqb2_2(.din(n307), .dout(n6566));
    jdff dff_A_GaIMETuo0_0(.din(n6560), .dout(G767gat));
    jdff dff_A_pRnNxhi55_0(.din(n6557), .dout(n6560));
    jdff dff_A_MhpwNvY03_0(.din(n6554), .dout(n6557));
    jdff dff_A_zayDYMAC9_0(.din(n6551), .dout(n6554));
    jdff dff_A_4cghf02G5_0(.din(n6548), .dout(n6551));
    jdff dff_A_lJZCFmRb2_0(.din(n6545), .dout(n6548));
    jdff dff_A_f4YfKqPQ5_0(.din(n6542), .dout(n6545));
    jdff dff_A_nRN3mXyO0_0(.din(n6539), .dout(n6542));
    jdff dff_A_VtjWYBoD7_0(.din(n6536), .dout(n6539));
    jdff dff_A_lKvVqxvf2_0(.din(n6533), .dout(n6536));
    jdff dff_A_M4wox5Ln1_0(.din(n6530), .dout(n6533));
    jdff dff_A_KL22KnRp0_0(.din(n6527), .dout(n6530));
    jdff dff_A_mgNFwFQI6_0(.din(n6524), .dout(n6527));
    jdff dff_A_zCXOxBdL0_0(.din(n6521), .dout(n6524));
    jdff dff_A_l10DnAiv7_0(.din(n6518), .dout(n6521));
    jdff dff_A_oSp4Wycw9_0(.din(n6515), .dout(n6518));
    jdff dff_A_dA3HrudG7_0(.din(n6512), .dout(n6515));
    jdff dff_A_HDSOKIyw3_0(.din(n6509), .dout(n6512));
    jdff dff_A_yrZBHJd72_0(.din(n6506), .dout(n6509));
    jdff dff_A_vXcrQt8P2_0(.din(n6503), .dout(n6506));
    jdff dff_A_2As3Gp9u4_0(.din(n6500), .dout(n6503));
    jdff dff_A_Mz9qLphq2_0(.din(n6497), .dout(n6500));
    jdff dff_A_TM5MgPuX3_0(.din(n6494), .dout(n6497));
    jdff dff_A_U7erAsDQ5_2(.din(n271), .dout(n6494));
    jdff dff_A_vyrLqLGJ4_0(.din(n6488), .dout(G450gat));
    jdff dff_A_D604cKvP7_0(.din(n6485), .dout(n6488));
    jdff dff_A_McwYecOY1_0(.din(n6482), .dout(n6485));
    jdff dff_A_QMKe07Im0_0(.din(n6479), .dout(n6482));
    jdff dff_A_lQ1dH66v6_0(.din(n6476), .dout(n6479));
    jdff dff_A_MdzUCVzI6_0(.din(n6473), .dout(n6476));
    jdff dff_A_YaBG4oSU9_0(.din(n6470), .dout(n6473));
    jdff dff_A_2vQiqEB96_0(.din(n6467), .dout(n6470));
    jdff dff_A_0RQkebOo9_0(.din(n6464), .dout(n6467));
    jdff dff_A_4c9L0DV80_0(.din(n6461), .dout(n6464));
    jdff dff_A_QikJSJ3d1_0(.din(n6458), .dout(n6461));
    jdff dff_A_uISI1WsD5_0(.din(n6455), .dout(n6458));
    jdff dff_A_COVMCks73_0(.din(n6452), .dout(n6455));
    jdff dff_A_hQgmV7lM8_0(.din(n6449), .dout(n6452));
    jdff dff_A_qd0YjtjN5_0(.din(n6446), .dout(n6449));
    jdff dff_A_pgP4yugU0_0(.din(n6443), .dout(n6446));
    jdff dff_A_q6NT3oCv1_0(.din(n6440), .dout(n6443));
    jdff dff_A_Ml5hqJBm4_0(.din(n6437), .dout(n6440));
    jdff dff_A_pkjTEZjv2_0(.din(n6434), .dout(n6437));
    jdff dff_A_8B4y4y9K3_0(.din(n6431), .dout(n6434));
    jdff dff_A_MLGMIGu43_0(.din(n6428), .dout(n6431));
    jdff dff_A_JdOCm0dx1_0(.din(n6425), .dout(n6428));
    jdff dff_A_9jwx3rml7_0(.din(n6422), .dout(n6425));
    jdff dff_A_wgptwsmK8_0(.din(n6419), .dout(n6422));
    jdff dff_A_C0PghwRv6_0(.din(n6416), .dout(n6419));
    jdff dff_A_46oFJh5I3_2(.din(n235), .dout(n6416));
    jdff dff_A_4P6xKnKW5_0(.din(n6410), .dout(G449gat));
    jdff dff_A_Retbe4sH3_0(.din(n6407), .dout(n6410));
    jdff dff_A_AqquzEvy1_0(.din(n6404), .dout(n6407));
    jdff dff_A_4N8IUoXA7_0(.din(n6401), .dout(n6404));
    jdff dff_A_gvAHydQ76_0(.din(n6398), .dout(n6401));
    jdff dff_A_fVFkq9qw8_0(.din(n6395), .dout(n6398));
    jdff dff_A_Vnn3D59h3_0(.din(n6392), .dout(n6395));
    jdff dff_A_rqYgT0Dl0_0(.din(n6389), .dout(n6392));
    jdff dff_A_z9iQBznL7_0(.din(n6386), .dout(n6389));
    jdff dff_A_AggPnzlb1_0(.din(n6383), .dout(n6386));
    jdff dff_A_HFBl8UVZ8_0(.din(n6380), .dout(n6383));
    jdff dff_A_3qJoRJzD0_0(.din(n6377), .dout(n6380));
    jdff dff_A_xuXfIYyy9_0(.din(n6374), .dout(n6377));
    jdff dff_A_ZEsUSQyw7_0(.din(n6371), .dout(n6374));
    jdff dff_A_B5NMwLW42_0(.din(n6368), .dout(n6371));
    jdff dff_A_GvkBVEZY7_0(.din(n6365), .dout(n6368));
    jdff dff_A_HtYxp3CU8_0(.din(n6362), .dout(n6365));
    jdff dff_A_50WfZlRv9_0(.din(n6359), .dout(n6362));
    jdff dff_A_ZwYGWjRz5_0(.din(n6356), .dout(n6359));
    jdff dff_A_wFDivU5a4_0(.din(n6353), .dout(n6356));
    jdff dff_A_Jgo03Sv45_0(.din(n6350), .dout(n6353));
    jdff dff_A_CgoddBim3_0(.din(n6347), .dout(n6350));
    jdff dff_A_VbVzM2jM1_2(.din(n231), .dout(n6347));
    jdff dff_A_eu2X2mip2_0(.din(n6341), .dout(G448gat));
    jdff dff_A_07fLWie52_0(.din(n6338), .dout(n6341));
    jdff dff_A_EJJpLg9J1_0(.din(n6335), .dout(n6338));
    jdff dff_A_Q3xRzlFV7_0(.din(n6332), .dout(n6335));
    jdff dff_A_VdSaoWRT1_0(.din(n6329), .dout(n6332));
    jdff dff_A_um8nsU6v7_0(.din(n6326), .dout(n6329));
    jdff dff_A_U2k9AOlS6_0(.din(n6323), .dout(n6326));
    jdff dff_A_8dZ3D4dc2_0(.din(n6320), .dout(n6323));
    jdff dff_A_KSV1Dyqt8_0(.din(n6317), .dout(n6320));
    jdff dff_A_S4xidspa6_0(.din(n6314), .dout(n6317));
    jdff dff_A_K6ykE9Es0_0(.din(n6311), .dout(n6314));
    jdff dff_A_mdki67i10_0(.din(n6308), .dout(n6311));
    jdff dff_A_3wsZMJIN8_0(.din(n6305), .dout(n6308));
    jdff dff_A_yII40mDR7_0(.din(n6302), .dout(n6305));
    jdff dff_A_Md0LfRkU8_0(.din(n6299), .dout(n6302));
    jdff dff_A_zM3QRekq3_0(.din(n6296), .dout(n6299));
    jdff dff_A_LcxT1DII1_0(.din(n6293), .dout(n6296));
    jdff dff_A_8RtDEWQX2_0(.din(n6290), .dout(n6293));
    jdff dff_A_6PQ7w8RY1_0(.din(n6287), .dout(n6290));
    jdff dff_A_72IKoJsn0_0(.din(n6284), .dout(n6287));
    jdff dff_A_Yl5exmZf3_0(.din(n6281), .dout(n6284));
    jdff dff_A_MhstYeIf3_0(.din(n6278), .dout(n6281));
    jdff dff_B_GSIaywte5_2(.din(n152), .dout(n2043));
    jdff dff_B_tAReGijg0_1(.din(G90gat), .dout(n2046));
    jdff dff_B_zHSEY54C2_1(.din(n195), .dout(n2049));
    jdff dff_B_kiZvJ92o9_1(.din(n127), .dout(n2052));
    jdff dff_A_xHbkrqDb3_1(.din(n2057), .dout(n2054));
    jdff dff_A_6u0KVS2n6_1(.din(n105), .dout(n2057));
    jdff dff_B_p7UUrr9R3_1(.din(G74gat), .dout(n2061));
    jdff dff_B_N3gDhnya0_1(.din(n2061), .dout(n2064));
    jdff dff_B_kggM7kW44_1(.din(n2064), .dout(n2067));
    jdff dff_B_qVLElNTY8_1(.din(G89gat), .dout(n2070));
    jdff dff_B_rs6GoOFe1_1(.din(n243), .dout(n2073));
    jdff dff_B_IYnRNLZA4_1(.din(G135gat), .dout(n2076));
    jdff dff_B_CaTEttEE8_1(.din(n279), .dout(n2079));
    jdff dff_A_VbHs2Mun8_1(.din(G130gat), .dout(n2081));
    jdff dff_B_xZ4cSpAA9_1(.din(G207gat), .dout(n2085));
    jdff dff_B_MsViwyTq7_1(.din(n555), .dout(n2088));
    jdff dff_B_KBWPjDHB7_1(.din(n2088), .dout(n2091));
    jdff dff_B_lBXbOrwb0_1(.din(n448), .dout(n2094));
    jdff dff_B_ZpbdFtNi8_1(.din(n2094), .dout(n2097));
    jdff dff_B_EPAe0jse5_1(.din(n519), .dout(n2100));
    jdff dff_B_yeiXuvcf0_0(.din(n539), .dout(n2103));
    jdff dff_B_UGuoYXmm1_0(.din(n2103), .dout(n2106));
    jdff dff_B_NiLdjS6E0_0(.din(n2106), .dout(n2109));
    jdff dff_B_iODpJsBp4_0(.din(n2109), .dout(n2112));
    jdff dff_B_CqEcUHpB6_0(.din(n2112), .dout(n2115));
    jdff dff_B_13NRcRbk2_0(.din(n2115), .dout(n2118));
    jdff dff_B_PRsgJq3f1_0(.din(n2118), .dout(n2121));
    jdff dff_B_ldYpc67U9_0(.din(n2121), .dout(n2124));
    jdff dff_B_qzjTKzz27_0(.din(n2124), .dout(n2127));
    jdff dff_B_4Awn7C4E9_0(.din(n444), .dout(n2130));
    jdff dff_B_7yALASj83_0(.din(n2130), .dout(n2133));
    jdff dff_B_RU1Eypu97_0(.din(n2133), .dout(n2136));
    jdff dff_B_aDLR7Kvq2_0(.din(n2136), .dout(n2139));
    jdff dff_B_glchsX2h6_0(.din(n2139), .dout(n2142));
    jdff dff_A_lbbwU5MU8_0(.din(n2147), .dout(n2144));
    jdff dff_A_ovymAdQG1_0(.din(n2150), .dout(n2147));
    jdff dff_A_SmruBy2C7_0(.din(n2153), .dout(n2150));
    jdff dff_A_jJiEuFvK4_0(.din(G201gat), .dout(n2153));
    jdff dff_B_KRXK0BIK7_1(.din(n637), .dout(n2157));
    jdff dff_B_JS8AxjnQ2_1(.din(n2157), .dout(n2160));
    jdff dff_B_CcigUWsG8_1(.din(n2160), .dout(n2163));
    jdff dff_B_Y30hR4Xq7_1(.din(n2163), .dout(n2166));
    jdff dff_B_cmC4qDUJ6_1(.din(n2166), .dout(n2169));
    jdff dff_B_4rqCsIZw9_1(.din(n2169), .dout(n2172));
    jdff dff_B_fDhPSzWG5_1(.din(n720), .dout(n2175));
    jdff dff_B_5tPrt5TS0_1(.din(n723), .dout(n2178));
    jdff dff_B_DMUQEEkT6_1(.din(n2178), .dout(n2181));
    jdff dff_B_5RxU2FrA5_1(.din(n2181), .dout(n2184));
    jdff dff_B_dQ96iAXH6_1(.din(n2184), .dout(n2187));
    jdff dff_B_8yNUeOwK7_1(.din(n2187), .dout(n2190));
    jdff dff_B_7UJ5sV2m1_1(.din(n2190), .dout(n2193));
    jdff dff_B_6pSDPMc78_1(.din(n601), .dout(n2196));
    jdff dff_B_7gnwILmQ9_1(.din(n2196), .dout(n2199));
    jdff dff_B_9AMMAbma1_1(.din(n605), .dout(n2202));
    jdff dff_B_RMJa3JFY2_1(.din(n2202), .dout(n2205));
    jdff dff_B_V2HBIQJY9_1(.din(n2205), .dout(n2208));
    jdff dff_B_7TXgyzlL9_1(.din(n2208), .dout(n2211));
    jdff dff_B_jQkrUx4e0_1(.din(n2211), .dout(n2214));
    jdff dff_B_84n8DlGf3_1(.din(n2214), .dout(n2217));
    jdff dff_B_uIXJncuN6_0(.din(n621), .dout(n2220));
    jdff dff_B_oVL95WD29_0(.din(n2220), .dout(n2223));
    jdff dff_B_BEQmc9da3_0(.din(n2223), .dout(n2226));
    jdff dff_B_mzBl8A180_0(.din(n2226), .dout(n2229));
    jdff dff_B_ff64FpwW7_0(.din(n2229), .dout(n2232));
    jdff dff_B_YFBtf0H28_0(.din(n2232), .dout(n2235));
    jdff dff_B_nqqmaY0D9_0(.din(n2235), .dout(n2238));
    jdff dff_B_7PLyaIN99_0(.din(n2238), .dout(n2241));
    jdff dff_A_EAMIyyQt3_1(.din(n4868), .dout(n2243));
    jdff dff_A_CXvq3uDD5_1(.din(n5201), .dout(n2246));
    jdff dff_A_RKnVw1t78_1(.din(n2252), .dout(n2249));
    jdff dff_A_LS30gOEK1_1(.din(n2255), .dout(n2252));
    jdff dff_A_XCbuhe4z0_1(.din(n2258), .dout(n2255));
    jdff dff_A_JtT7Xivj8_1(.din(n2261), .dout(n2258));
    jdff dff_A_YIUMp9I11_1(.din(n2264), .dout(n2261));
    jdff dff_A_qgTNje5x7_1(.din(n2267), .dout(n2264));
    jdff dff_A_HzVUopj19_1(.din(n597), .dout(n2267));
    jdff dff_A_IaniZYls9_0(.din(n2273), .dout(n2270));
    jdff dff_A_o46JxSdL2_0(.din(n2276), .dout(n2273));
    jdff dff_A_8hignWYJ0_0(.din(n2279), .dout(n2276));
    jdff dff_A_SYl1ZTaK7_0(.din(G183gat), .dout(n2279));
    jdff dff_A_foXrpMJg4_1(.din(n2285), .dout(n2282));
    jdff dff_A_QQFj4ndL4_1(.din(n2288), .dout(n2285));
    jdff dff_A_0uaWIG1l7_1(.din(n2291), .dout(n2288));
    jdff dff_A_NLAVdITU2_1(.din(n2294), .dout(n2291));
    jdff dff_A_ODHcvoO50_1(.din(n2297), .dout(n2294));
    jdff dff_A_dGtI2dac5_1(.din(n2300), .dout(n2297));
    jdff dff_A_84Y2JVtx4_1(.din(n2303), .dout(n2300));
    jdff dff_A_0099FcX74_1(.din(G183gat), .dout(n2303));
    jdff dff_A_j14IaQH59_1(.din(n4998), .dout(n2306));
    jdff dff_B_tPIYVKvH9_1(.din(n827), .dout(n2310));
    jdff dff_B_F0f1ClMC4_1(.din(n2310), .dout(n2313));
    jdff dff_B_A932LBmu1_1(.din(n2313), .dout(n2316));
    jdff dff_B_ijtp4fIJ1_1(.din(n2316), .dout(n2319));
    jdff dff_B_lTkxRn4p5_1(.din(n2319), .dout(n2322));
    jdff dff_B_FU6iXRqU8_1(.din(n831), .dout(n2325));
    jdff dff_B_Hu5j9bju6_0(.din(n834), .dout(n2328));
    jdff dff_B_TLrXwqyY7_0(.din(n2328), .dout(n2331));
    jdff dff_B_P7XkTJJ67_0(.din(n2331), .dout(n2334));
    jdff dff_B_JIUTpmJ50_0(.din(n2334), .dout(n2337));
    jdff dff_A_jO3Qq5u22_0(.din(n2342), .dout(n2339));
    jdff dff_A_I47TRL0K7_0(.din(n2345), .dout(n2342));
    jdff dff_A_cswhGIzL9_0(.din(n3909), .dout(n2345));
    jdff dff_A_aF2RwkzK0_1(.din(n2351), .dout(n2348));
    jdff dff_A_PVgGCB742_1(.din(n2354), .dout(n2351));
    jdff dff_A_HcTM1GVX3_1(.din(n2357), .dout(n2354));
    jdff dff_A_kEdOAhc04_1(.din(n2360), .dout(n2357));
    jdff dff_A_jC3o60vi7_1(.din(n3909), .dout(n2360));
    jdff dff_B_s73pqaah1_1(.din(n787), .dout(n2364));
    jdff dff_B_nn6wMOGk0_0(.din(n819), .dout(n2367));
    jdff dff_B_7cjJs6LO5_0(.din(n2367), .dout(n2370));
    jdff dff_B_20CebZ979_0(.din(n2370), .dout(n2373));
    jdff dff_B_6E7KgVIu3_0(.din(n2373), .dout(n2376));
    jdff dff_B_9r22lERW4_1(.din(n811), .dout(n2379));
    jdff dff_B_OmeFB6pZ1_1(.din(n2379), .dout(n2382));
    jdff dff_B_H0zx1ZtW2_1(.din(n2382), .dout(n2385));
    jdff dff_B_3ZMkq8Hj4_1(.din(n2385), .dout(n2388));
    jdff dff_B_x3DtjL5f7_1(.din(n791), .dout(n2391));
    jdff dff_B_1a2TZAgG4_1(.din(n2391), .dout(n2394));
    jdff dff_B_Y1cVy0MP9_1(.din(n2394), .dout(n2397));
    jdff dff_B_D8OM8Dun0_1(.din(n2397), .dout(n2400));
    jdff dff_B_nomCx90E8_1(.din(n2400), .dout(n2403));
    jdff dff_B_rBgMgBtT9_1(.din(n2403), .dout(n2406));
    jdff dff_B_WCr7dEsS6_1(.din(n2406), .dout(n2409));
    jdff dff_B_eALMfTKs8_1(.din(n2409), .dout(n2412));
    jdff dff_B_WS4odQnb5_0(.din(n799), .dout(n2415));
    jdff dff_B_iQF6CmOP3_0(.din(n2415), .dout(n2418));
    jdff dff_B_eNyofXta8_0(.din(n2418), .dout(n2421));
    jdff dff_B_5LYf5VqB1_0(.din(n2421), .dout(n2424));
    jdff dff_B_mXgbvMDp2_0(.din(n2424), .dout(n2427));
    jdff dff_B_XpaDHBzu2_0(.din(n2427), .dout(n2430));
    jdff dff_A_ma28hyni2_1(.din(n2435), .dout(n2432));
    jdff dff_A_ryLF9ho38_1(.din(n2438), .dout(n2435));
    jdff dff_A_MICi2kaS5_1(.din(n2441), .dout(n2438));
    jdff dff_A_oPYePDtu1_1(.din(n2444), .dout(n2441));
    jdff dff_A_Ld9vuEK63_1(.din(n783), .dout(n2444));
    jdff dff_B_sv0h8F5G0_1(.din(n898), .dout(n2448));
    jdff dff_B_doZbIsdq4_1(.din(n2448), .dout(n2451));
    jdff dff_B_quorBJTR4_1(.din(n2451), .dout(n2454));
    jdff dff_B_FdyFEEuq6_1(.din(n902), .dout(n2457));
    jdff dff_B_yFZnzdM23_0(.din(n905), .dout(n2460));
    jdff dff_B_uQCll2v58_0(.din(n2460), .dout(n2463));
    jdff dff_B_uYfs2cxK6_1(.din(n858), .dout(n2466));
    jdff dff_B_hQhrmT7l8_0(.din(n890), .dout(n2469));
    jdff dff_B_vqXqbZSx8_0(.din(n2469), .dout(n2472));
    jdff dff_B_zCUSekvJ1_0(.din(n2472), .dout(n2475));
    jdff dff_B_9QPYehDS4_0(.din(n2475), .dout(n2478));
    jdff dff_B_pfDKVsB08_0(.din(n886), .dout(n2481));
    jdff dff_B_N6L8NkBI2_0(.din(n2481), .dout(n2484));
    jdff dff_B_itdv4hEJ5_0(.din(n2484), .dout(n2487));
    jdff dff_B_pg4cL8EJ9_0(.din(n2487), .dout(n2490));
    jdff dff_B_A16QuiJk1_1(.din(n862), .dout(n2493));
    jdff dff_B_D1GtwHkq2_1(.din(n2493), .dout(n2496));
    jdff dff_B_lbCEY3NP1_1(.din(n2496), .dout(n2499));
    jdff dff_B_TY17PhMk2_1(.din(n2499), .dout(n2502));
    jdff dff_B_BJwEZ6133_1(.din(n2502), .dout(n2505));
    jdff dff_B_dDcipXBN9_1(.din(n2505), .dout(n2508));
    jdff dff_B_6OVoBhBC5_1(.din(n2508), .dout(n2511));
    jdff dff_B_Cx9viwQK4_1(.din(n2511), .dout(n2514));
    jdff dff_B_KKr6Xmht4_0(.din(n870), .dout(n2517));
    jdff dff_B_oFbHHbPU4_0(.din(n2517), .dout(n2520));
    jdff dff_B_IJ1xQlMV2_0(.din(n2520), .dout(n2523));
    jdff dff_B_XSdgvg7a2_0(.din(n2523), .dout(n2526));
    jdff dff_B_WGeQ4lVH4_0(.din(n2526), .dout(n2529));
    jdff dff_B_Cy6GudwD7_0(.din(n2529), .dout(n2532));
    jdff dff_A_A6pBvmPj2_1(.din(n2537), .dout(n2534));
    jdff dff_A_uSC7OrEy1_1(.din(n2540), .dout(n2537));
    jdff dff_A_KWSQz0Ql4_1(.din(n854), .dout(n2540));
    jdff dff_B_Rbgx2vm75_1(.din(n961), .dout(n2544));
    jdff dff_B_3eNKzKk52_1(.din(n2544), .dout(n2547));
    jdff dff_B_AzUGH2hI5_1(.din(n2547), .dout(n2550));
    jdff dff_B_ml8j43294_1(.din(n2550), .dout(n2553));
    jdff dff_B_VakEVg175_1(.din(n2553), .dout(n2556));
    jdff dff_B_20wcC6Ne3_1(.din(n2556), .dout(n2559));
    jdff dff_B_g8o3Zviv8_1(.din(n2559), .dout(n2562));
    jdff dff_B_5cFhrUcq6_1(.din(n2562), .dout(n2565));
    jdff dff_B_QKePrQ611_1(.din(n2565), .dout(n2568));
    jdff dff_B_ghwV2H0S0_1(.din(n2568), .dout(n2571));
    jdff dff_B_eJ50nooN0_1(.din(n2571), .dout(n2574));
    jdff dff_B_HEUlk5BE9_1(.din(n2574), .dout(n2577));
    jdff dff_B_voHXs2Qa4_1(.din(n2577), .dout(n2580));
    jdff dff_B_8r6bEAey5_1(.din(n2580), .dout(n2583));
    jdff dff_B_vSOUwK2N3_1(.din(n2583), .dout(n2586));
    jdff dff_B_efrgUlBb8_1(.din(n965), .dout(n2589));
    jdff dff_B_fFyNbHDS8_1(.din(n2589), .dout(n2592));
    jdff dff_B_LbgnQHev8_1(.din(n2592), .dout(n2595));
    jdff dff_B_P8gRLnd94_1(.din(n2595), .dout(n2598));
    jdff dff_B_JeXEp6s22_1(.din(n2598), .dout(n2601));
    jdff dff_B_cK3e9Z3T8_1(.din(n2601), .dout(n2604));
    jdff dff_B_BUnj0QyW7_1(.din(n2604), .dout(n2607));
    jdff dff_B_0f3GhMrc8_1(.din(n2607), .dout(n2610));
    jdff dff_B_agPU4M1E7_1(.din(n2610), .dout(n2613));
    jdff dff_B_yxqbIcDq2_1(.din(n2613), .dout(n2616));
    jdff dff_B_RmIz27ih2_1(.din(n2616), .dout(n2619));
    jdff dff_B_TCubaHiW8_1(.din(n2619), .dout(n2622));
    jdff dff_B_Crsi5cq54_1(.din(n2622), .dout(n2625));
    jdff dff_B_G5W7pFqL9_1(.din(n2625), .dout(n2628));
    jdff dff_A_xVCbd2lf1_0(.din(n2633), .dout(n2630));
    jdff dff_A_HC0x09Pj9_0(.din(n2636), .dout(n2633));
    jdff dff_A_kR5YIjbe0_0(.din(n2639), .dout(n2636));
    jdff dff_A_ATAq18RA7_0(.din(n2642), .dout(n2639));
    jdff dff_A_568KjyB94_0(.din(n2645), .dout(n2642));
    jdff dff_A_DqioWgSz5_0(.din(n2648), .dout(n2645));
    jdff dff_A_es7kT23C2_0(.din(n2651), .dout(n2648));
    jdff dff_A_1BKxyyK10_0(.din(n2654), .dout(n2651));
    jdff dff_A_O8Vklup97_0(.din(G159gat), .dout(n2654));
    jdff dff_A_DFUfRgTK0_1(.din(n2660), .dout(n2657));
    jdff dff_A_t2TQ3gLM1_1(.din(n2663), .dout(n2660));
    jdff dff_A_ULzcb9f16_1(.din(n2666), .dout(n2663));
    jdff dff_A_Exgb0kkr0_1(.din(n2669), .dout(n2666));
    jdff dff_A_LLlRukt87_1(.din(n2672), .dout(n2669));
    jdff dff_A_gnkWmC5J5_1(.din(n2675), .dout(n2672));
    jdff dff_A_Cz0Cu0aV2_1(.din(n2678), .dout(n2675));
    jdff dff_A_jFhtMyKy5_1(.din(n2681), .dout(n2678));
    jdff dff_A_5rMxZFOJ6_1(.din(G159gat), .dout(n2681));
    jdff dff_B_GPhE9peD1_1(.din(n1138), .dout(n2685));
    jdff dff_B_dDZMWDgu2_1(.din(n2685), .dout(n2688));
    jdff dff_B_FN5MSQz78_0(.din(n1189), .dout(n2691));
    jdff dff_B_JOYH0Xz12_0(.din(n2691), .dout(n2694));
    jdff dff_B_FuOOvbjw1_0(.din(n2694), .dout(n2697));
    jdff dff_B_nhK3TEkx1_0(.din(n2697), .dout(n2700));
    jdff dff_B_YJfwExrU1_0(.din(n2700), .dout(n2703));
    jdff dff_B_1pV9Y5bC2_0(.din(n2703), .dout(n2706));
    jdff dff_B_oM4e1fGD4_0(.din(n2706), .dout(n2709));
    jdff dff_B_oYpqn9Si8_0(.din(n2709), .dout(n2712));
    jdff dff_B_KIQzMffs8_0(.din(n2712), .dout(n2715));
    jdff dff_B_45YLzm8C4_0(.din(n1181), .dout(n2718));
    jdff dff_B_t1lwdvkp9_0(.din(n2718), .dout(n2721));
    jdff dff_B_mCEZtpVI8_0(.din(n2721), .dout(n2724));
    jdff dff_B_3ejL3m9E0_0(.din(n2724), .dout(n2727));
    jdff dff_B_gpVBdfsV2_1(.din(n1173), .dout(n2730));
    jdff dff_B_3nLihxdL9_1(.din(n2730), .dout(n2733));
    jdff dff_B_1r9sycvd2_1(.din(n2733), .dout(n2736));
    jdff dff_B_C2QS22wE8_1(.din(n2736), .dout(n2739));
    jdff dff_A_59789IK71_0(.din(n2744), .dout(n2741));
    jdff dff_A_vxoLuX1Q7_0(.din(n2747), .dout(n2744));
    jdff dff_A_JhfWkjJ38_0(.din(n2750), .dout(n2747));
    jdff dff_A_7VJLBtPY3_0(.din(n2753), .dout(n2750));
    jdff dff_A_sGzLHVee3_0(.din(n2756), .dout(n2753));
    jdff dff_A_g8THXuPB6_0(.din(n2759), .dout(n2756));
    jdff dff_A_tNk60cMu8_0(.din(n2762), .dout(n2759));
    jdff dff_A_h4gHO2iu9_0(.din(n4890), .dout(n2762));
    jdff dff_A_eThL9HM11_0(.din(n2768), .dout(n2765));
    jdff dff_A_gDlbk4Ia6_0(.din(n2771), .dout(n2768));
    jdff dff_A_ch7dmcIp8_0(.din(n2774), .dout(n2771));
    jdff dff_A_2UGetOFz2_0(.din(n2777), .dout(n2774));
    jdff dff_A_u2asBRF63_0(.din(n2780), .dout(n2777));
    jdff dff_A_MSP3JsP91_0(.din(n2783), .dout(n2780));
    jdff dff_A_Fb5zEkqL0_0(.din(n2786), .dout(n2783));
    jdff dff_A_zu6g0c7R2_0(.din(n2789), .dout(n2786));
    jdff dff_A_1LorvZwg6_0(.din(n2792), .dout(n2789));
    jdff dff_A_Gs7sp7nX6_0(.din(G237gat), .dout(n2792));
    jdff dff_A_lBzLUwpW9_0(.din(n2798), .dout(n2795));
    jdff dff_A_G51sbAmz5_0(.din(n2801), .dout(n2798));
    jdff dff_A_nDEMpseI7_0(.din(n2804), .dout(n2801));
    jdff dff_A_BUhkNS0b3_0(.din(n2807), .dout(n2804));
    jdff dff_A_tIFLXirb2_0(.din(n2810), .dout(n2807));
    jdff dff_A_Oe9a0CGt2_0(.din(n2813), .dout(n2810));
    jdff dff_A_REtwFYfb2_0(.din(n2816), .dout(n2813));
    jdff dff_A_XYTdUqX19_0(.din(n2819), .dout(n2816));
    jdff dff_A_W48Xm7nX1_0(.din(n2822), .dout(n2819));
    jdff dff_A_XHTaupih4_0(.din(n4998), .dout(n2822));
    jdff dff_B_n2gwc0Wj5_1(.din(n1130), .dout(n2826));
    jdff dff_B_b8rYDj6P0_1(.din(n2826), .dout(n2829));
    jdff dff_B_3TSyV1bV3_1(.din(n2829), .dout(n2832));
    jdff dff_B_GuAntEwq1_1(.din(n2832), .dout(n2835));
    jdff dff_B_j7SlwgB99_1(.din(n2835), .dout(n2838));
    jdff dff_B_kh9VxO0k5_1(.din(n2838), .dout(n2841));
    jdff dff_B_ndfcPuaT1_1(.din(n2841), .dout(n2844));
    jdff dff_B_bYpKujEX4_1(.din(n2844), .dout(n2847));
    jdff dff_A_bJ3daH7s7_0(.din(n2852), .dout(n2849));
    jdff dff_A_FFFIshbQ3_0(.din(n2855), .dout(n2852));
    jdff dff_A_qtemNoQF6_0(.din(n2858), .dout(n2855));
    jdff dff_A_GArnw1Hh2_0(.din(n2861), .dout(n2858));
    jdff dff_A_veE51J5r6_0(.din(n3872), .dout(n2861));
    jdff dff_A_sidqFTyr6_1(.din(n2867), .dout(n2864));
    jdff dff_A_q8r5PICu7_1(.din(n2870), .dout(n2867));
    jdff dff_A_MoxOgXXi2_1(.din(n2873), .dout(n2870));
    jdff dff_A_5ThYq8HY6_1(.din(n2876), .dout(n2873));
    jdff dff_A_HdP8i38R0_1(.din(n3872), .dout(n2876));
    jdff dff_A_tSxS8ex92_0(.din(n2882), .dout(n2879));
    jdff dff_A_9HdxmpXx7_0(.din(n2885), .dout(n2882));
    jdff dff_A_k2Q75X6R6_0(.din(n2888), .dout(n2885));
    jdff dff_A_7iYUx3bS4_0(.din(n2891), .dout(n2888));
    jdff dff_A_c2ulKy9Q7_0(.din(n2894), .dout(n2891));
    jdff dff_A_zxLR4eFD5_0(.din(n2897), .dout(n2894));
    jdff dff_A_MuNfmDZT5_0(.din(n2900), .dout(n2897));
    jdff dff_A_LCf2uBmQ9_0(.din(n2903), .dout(n2900));
    jdff dff_A_9Z1wnDuS3_0(.din(n2906), .dout(n2903));
    jdff dff_A_WTmwzHhH3_0(.din(n1127), .dout(n2906));
    jdff dff_B_70CWGrjI8_1(.din(n1237), .dout(n2910));
    jdff dff_B_K4KwPQzj4_1(.din(n2910), .dout(n2913));
    jdff dff_B_elh2Lk664_1(.din(n2913), .dout(n2916));
    jdff dff_B_QJXJPvJC7_1(.din(n2916), .dout(n2919));
    jdff dff_B_JcgMogmf8_1(.din(n2919), .dout(n2922));
    jdff dff_B_TAxAW1TE0_1(.din(n2922), .dout(n2925));
    jdff dff_B_p6qSeAFm5_1(.din(n2925), .dout(n2928));
    jdff dff_B_UBdkgCNo1_1(.din(n2928), .dout(n2931));
    jdff dff_B_3TIzWT7q7_1(.din(n2931), .dout(n2934));
    jdff dff_B_jllHzEmu8_1(.din(n2934), .dout(n2937));
    jdff dff_B_dZ8btkFc7_1(.din(n2937), .dout(n2940));
    jdff dff_B_ZJiliUBo6_1(.din(n2940), .dout(n2943));
    jdff dff_B_ijMSrt5x0_1(.din(n2943), .dout(n2946));
    jdff dff_B_mfXSlU7j1_1(.din(n1241), .dout(n2949));
    jdff dff_B_gjEntSGG0_0(.din(n1283), .dout(n2952));
    jdff dff_B_TtY3cPI91_0(.din(n2952), .dout(n2955));
    jdff dff_B_eeKoyiNY8_0(.din(n2955), .dout(n2958));
    jdff dff_B_0UUyqVNO3_0(.din(n2958), .dout(n2961));
    jdff dff_B_nS0kYOT68_0(.din(n2961), .dout(n2964));
    jdff dff_B_LavBUcDn8_0(.din(n2964), .dout(n2967));
    jdff dff_B_x7scORUO7_0(.din(n2967), .dout(n2970));
    jdff dff_B_bnIP7UBA7_0(.din(n2970), .dout(n2973));
    jdff dff_B_dEFVNWWr4_0(.din(n2973), .dout(n2976));
    jdff dff_B_E5dNJnVk6_0(.din(n2976), .dout(n2979));
    jdff dff_B_ekhsX9qf0_0(.din(n2979), .dout(n2982));
    jdff dff_B_zyDzmDZh4_0(.din(n2982), .dout(n2985));
    jdff dff_B_1H8axePV9_0(.din(n2985), .dout(n2988));
    jdff dff_B_fp7LMI6Y1_1(.din(n1244), .dout(n2991));
    jdff dff_B_2NjnirCd9_1(.din(n2991), .dout(n2994));
    jdff dff_B_ecR09ZOB4_1(.din(n2994), .dout(n2997));
    jdff dff_B_bRMTJVsK4_1(.din(n2997), .dout(n3000));
    jdff dff_B_y3lGjh756_1(.din(n3000), .dout(n3003));
    jdff dff_B_jU7pNuAJ5_1(.din(n3003), .dout(n3006));
    jdff dff_B_WFd4YglH5_1(.din(n3006), .dout(n3009));
    jdff dff_B_Di7pQTo20_1(.din(n3009), .dout(n3012));
    jdff dff_B_OBxQareG3_1(.din(n3012), .dout(n3015));
    jdff dff_B_dcIdBJQX2_1(.din(n3015), .dout(n3018));
    jdff dff_B_yueMlWGZ3_1(.din(n3018), .dout(n3021));
    jdff dff_B_YkK2LiLL9_1(.din(n3021), .dout(n3024));
    jdff dff_B_aHvNFreD1_1(.din(n1247), .dout(n3027));
    jdff dff_B_CSXGgycY4_1(.din(n3027), .dout(n3030));
    jdff dff_B_Up8wcUm81_1(.din(n3030), .dout(n3033));
    jdff dff_B_xRKcFhbq1_1(.din(n3033), .dout(n3036));
    jdff dff_B_jubtWu7l6_1(.din(n3036), .dout(n3039));
    jdff dff_B_kSzUQxZW4_1(.din(n3039), .dout(n3042));
    jdff dff_B_O0Co4cgu7_1(.din(n3042), .dout(n3045));
    jdff dff_B_N6UCPSSF5_1(.din(n3045), .dout(n3048));
    jdff dff_B_aKNoyOfg5_1(.din(n3048), .dout(n3051));
    jdff dff_B_eDgVJC478_1(.din(n3051), .dout(n3054));
    jdff dff_B_ORnpkLBA5_1(.din(n3054), .dout(n3057));
    jdff dff_A_SPd4hQoH9_1(.din(n3062), .dout(n3059));
    jdff dff_A_alXJXg7B6_1(.din(n3065), .dout(n3062));
    jdff dff_A_dHrcjvzZ0_1(.din(n3068), .dout(n3065));
    jdff dff_A_5zOnVWgp5_1(.din(n3071), .dout(n3068));
    jdff dff_A_WtDQ0C6I6_1(.din(n3074), .dout(n3071));
    jdff dff_A_MN2wCX0R6_1(.din(n3077), .dout(n3074));
    jdff dff_A_kiWtPUaK0_1(.din(n3080), .dout(n3077));
    jdff dff_A_kDsYcmTD4_1(.din(n3083), .dout(n3080));
    jdff dff_A_S0lkKPoz1_1(.din(n3086), .dout(n3083));
    jdff dff_A_k27b6J7i0_1(.din(n3089), .dout(n3086));
    jdff dff_A_xpGovbfh8_1(.din(n3092), .dout(n3089));
    jdff dff_A_uy3vY4jq6_1(.din(n997), .dout(n3092));
    jdff dff_A_i3iRedDT1_1(.din(n3098), .dout(n3095));
    jdff dff_A_Vtb3yNv80_1(.din(n3101), .dout(n3098));
    jdff dff_A_NB21JOM31_1(.din(n3104), .dout(n3101));
    jdff dff_A_8FnFl0Ka1_1(.din(n3107), .dout(n3104));
    jdff dff_A_Bfh220527_1(.din(n3110), .dout(n3107));
    jdff dff_A_Bd3YpNBu6_1(.din(n3113), .dout(n3110));
    jdff dff_A_L2jm9TSj8_1(.din(n3116), .dout(n3113));
    jdff dff_A_RzrELDkc0_1(.din(n3119), .dout(n3116));
    jdff dff_A_5DNRdYme2_1(.din(n3122), .dout(n3119));
    jdff dff_A_rwqahejY1_1(.din(n3125), .dout(n3122));
    jdff dff_A_Wm0Jxyom7_1(.din(n3128), .dout(n3125));
    jdff dff_A_P7w0ZNjN8_1(.din(n3131), .dout(n3128));
    jdff dff_A_pcKRiF3c5_1(.din(n993), .dout(n3131));
    jdff dff_A_f0Tnz2Rf4_0(.din(n3137), .dout(n3134));
    jdff dff_A_hYU0cSRm4_0(.din(n3140), .dout(n3137));
    jdff dff_A_IKgKATdn5_0(.din(n3143), .dout(n3140));
    jdff dff_A_0392metA6_0(.din(n3146), .dout(n3143));
    jdff dff_A_hfHBCBrd4_0(.din(n3149), .dout(n3146));
    jdff dff_A_mwI5hC6T4_0(.din(n3152), .dout(n3149));
    jdff dff_A_BjfqaBXx3_0(.din(n3155), .dout(n3152));
    jdff dff_A_e8Ofl2I68_0(.din(n3759), .dout(n3155));
    jdff dff_A_C391u25s3_1(.din(n3161), .dout(n3158));
    jdff dff_A_zPqbXuor2_1(.din(n3164), .dout(n3161));
    jdff dff_A_cx3u6k8U7_1(.din(n3167), .dout(n3164));
    jdff dff_A_EZKn2qb88_1(.din(n3170), .dout(n3167));
    jdff dff_A_Rm1vi7Dm2_1(.din(n3173), .dout(n3170));
    jdff dff_A_T6MFeb4P1_1(.din(n3176), .dout(n3173));
    jdff dff_A_Ubtbp1NT0_1(.din(n3179), .dout(n3176));
    jdff dff_A_gCsMnsrE5_1(.din(n3759), .dout(n3179));
    jdff dff_B_TnSxArNL8_1(.din(n1209), .dout(n3183));
    jdff dff_B_KipvtkXk5_0(.din(n1229), .dout(n3186));
    jdff dff_B_dhwGUi4C4_0(.din(n3186), .dout(n3189));
    jdff dff_B_MHrCsJvJ9_0(.din(n1221), .dout(n3192));
    jdff dff_B_CpbJkFt88_0(.din(n3192), .dout(n3195));
    jdff dff_B_HtzshIPQ6_0(.din(n3195), .dout(n3198));
    jdff dff_B_Its1ghR50_0(.din(n3198), .dout(n3201));
    jdff dff_B_qBnUhGcF5_0(.din(n3201), .dout(n3204));
    jdff dff_B_7sJIehnG8_0(.din(n3204), .dout(n3207));
    jdff dff_B_3ohoTttX1_0(.din(n3207), .dout(n3210));
    jdff dff_B_BYWnBMy53_0(.din(n3210), .dout(n3213));
    jdff dff_B_VrBGeUMi8_0(.din(n3213), .dout(n3216));
    jdff dff_B_bwf0huTv8_0(.din(n3216), .dout(n3219));
    jdff dff_A_7ATrk8lA0_1(.din(n3224), .dout(n3221));
    jdff dff_A_fI0k704R3_1(.din(n3227), .dout(n3224));
    jdff dff_A_FTX2Vn1G9_1(.din(n3230), .dout(n3227));
    jdff dff_A_oTX2lA851_1(.din(n3233), .dout(n3230));
    jdff dff_A_6elblald0_1(.din(n3236), .dout(n3233));
    jdff dff_A_wOf0Vs3J2_1(.din(n3239), .dout(n3236));
    jdff dff_A_rEdaWlZD6_1(.din(n3242), .dout(n3239));
    jdff dff_A_wpFhUrYf7_1(.din(n3245), .dout(n3242));
    jdff dff_A_1zoxcUQz6_1(.din(n3248), .dout(n3245));
    jdff dff_A_5uR6ew4C1_1(.din(n3251), .dout(n3248));
    jdff dff_A_PzTRTfC43_1(.din(n3254), .dout(n3251));
    jdff dff_A_QWIExkVG9_1(.din(n3257), .dout(n3254));
    jdff dff_A_xHEuLEKk9_1(.din(n3260), .dout(n3257));
    jdff dff_A_L9BAJdW84_1(.din(n1213), .dout(n3260));
    jdff dff_B_CLxBbHRk0_1(.din(n941), .dout(n3264));
    jdff dff_B_mE57rEnW3_0(.din(n949), .dout(n3267));
    jdff dff_B_JyLV2Q8U5_0(.din(n3267), .dout(n3270));
    jdff dff_B_iqj695lP5_0(.din(n3270), .dout(n3273));
    jdff dff_B_I7u5Bzyw3_0(.din(n3273), .dout(n3276));
    jdff dff_B_hAr2lqVH2_0(.din(n3276), .dout(n3279));
    jdff dff_B_gNuOt0Qh5_0(.din(n3279), .dout(n3282));
    jdff dff_B_mf2zHNDT5_1(.din(n929), .dout(n3285));
    jdff dff_A_RPvBiwtN1_1(.din(n3290), .dout(n3287));
    jdff dff_A_AhNfZjqw4_1(.din(n3293), .dout(n3290));
    jdff dff_A_ii5jO80d8_1(.din(n3296), .dout(n3293));
    jdff dff_A_FRKPHSb78_1(.din(n3299), .dout(n3296));
    jdff dff_A_xfzsnMIv6_1(.din(n3302), .dout(n3299));
    jdff dff_A_BAHIDpAU2_1(.din(n3305), .dout(n3302));
    jdff dff_A_KrKVBosd4_1(.din(n3308), .dout(n3305));
    jdff dff_A_mztmAX8J0_1(.din(n3311), .dout(n3308));
    jdff dff_A_Cdh1RHdS9_1(.din(G159gat), .dout(n3311));
    jdff dff_A_Lq5lGMV70_2(.din(n3317), .dout(n3314));
    jdff dff_A_mS6P4vMk2_2(.din(n3320), .dout(n3317));
    jdff dff_A_zjTxZgD94_2(.din(n3323), .dout(n3320));
    jdff dff_A_D4q2zQEj8_2(.din(n3326), .dout(n3323));
    jdff dff_A_OiQ2ftAf5_2(.din(n3329), .dout(n3326));
    jdff dff_A_LA9QaM5A7_2(.din(n3332), .dout(n3329));
    jdff dff_A_U6k3qrq82_2(.din(n3335), .dout(n3332));
    jdff dff_A_l6nWrpZy7_2(.din(n3338), .dout(n3335));
    jdff dff_A_WIZqdezD2_2(.din(n3341), .dout(n3338));
    jdff dff_A_Gj1DOGlz4_2(.din(n3344), .dout(n3341));
    jdff dff_A_ooxJvQMe3_2(.din(G159gat), .dout(n3344));
    jdff dff_B_IxmWWaaA2_1(.din(n1339), .dout(n3348));
    jdff dff_B_6niYvNzb6_1(.din(n3348), .dout(n3351));
    jdff dff_B_Kpy8p9277_1(.din(n3351), .dout(n3354));
    jdff dff_B_Fr1O2fo07_1(.din(n3354), .dout(n3357));
    jdff dff_B_o3W47Yud8_1(.din(n3357), .dout(n3360));
    jdff dff_B_ZQQbyMHB4_1(.din(n3360), .dout(n3363));
    jdff dff_B_SpTcmguP0_1(.din(n3363), .dout(n3366));
    jdff dff_B_ThYCInlC6_1(.din(n3366), .dout(n3369));
    jdff dff_B_TgmfaMBk4_1(.din(n3369), .dout(n3372));
    jdff dff_B_8fNxos089_1(.din(n3372), .dout(n3375));
    jdff dff_B_b77xlsdY5_1(.din(n3375), .dout(n3378));
    jdff dff_B_mebxrYF86_1(.din(n1343), .dout(n3381));
    jdff dff_B_5sJrgmDu4_0(.din(n1346), .dout(n3384));
    jdff dff_B_1pydwt8Y6_0(.din(n3384), .dout(n3387));
    jdff dff_B_BzkI7QOS5_0(.din(n3387), .dout(n3390));
    jdff dff_B_ObuiwlhG6_0(.din(n3390), .dout(n3393));
    jdff dff_B_uQgBBIEg4_0(.din(n3393), .dout(n3396));
    jdff dff_B_mi3XB9ba4_0(.din(n3396), .dout(n3399));
    jdff dff_B_P6C7vMeD7_0(.din(n3399), .dout(n3402));
    jdff dff_B_VKR7baJS2_0(.din(n3402), .dout(n3405));
    jdff dff_B_D9jll0ar0_0(.din(n3405), .dout(n3408));
    jdff dff_B_6pyf0hvZ3_0(.din(n3408), .dout(n3411));
    jdff dff_B_2CBrTZA57_0(.din(n3411), .dout(n3414));
    jdff dff_B_UZNijE2z1_1(.din(n1250), .dout(n3417));
    jdff dff_B_3LU1e96R4_1(.din(n3417), .dout(n3420));
    jdff dff_B_XRT4DgV51_1(.din(n3420), .dout(n3423));
    jdff dff_B_YLPxsV2m2_1(.din(n3423), .dout(n3426));
    jdff dff_B_eF1gTHkW1_1(.din(n3426), .dout(n3429));
    jdff dff_B_E0dRo7Ap4_1(.din(n3429), .dout(n3432));
    jdff dff_B_pwYc6g3t5_1(.din(n3432), .dout(n3435));
    jdff dff_B_1LJfeufW8_1(.din(n3435), .dout(n3438));
    jdff dff_B_0NfAE29N8_1(.din(n3438), .dout(n3441));
    jdff dff_B_BPEUKfMy0_1(.din(n3441), .dout(n3444));
    jdff dff_B_oEAOUbTH8_1(.din(n1253), .dout(n3447));
    jdff dff_B_gJRVFlMj1_1(.din(n3447), .dout(n3450));
    jdff dff_B_E5vJf1TA7_1(.din(n3450), .dout(n3453));
    jdff dff_B_PQc7fllE3_1(.din(n3453), .dout(n3456));
    jdff dff_B_9ixuTAQ49_1(.din(n3456), .dout(n3459));
    jdff dff_B_UtgkDoeP8_1(.din(n3459), .dout(n3462));
    jdff dff_B_qejEdbeU3_1(.din(n3462), .dout(n3465));
    jdff dff_B_rmn6hfnz2_1(.din(n3465), .dout(n3468));
    jdff dff_B_A3NTip0I7_1(.din(n3468), .dout(n3471));
    jdff dff_A_d2q87DtS4_1(.din(n3476), .dout(n3473));
    jdff dff_A_XFTT5lTa1_1(.din(n3479), .dout(n3476));
    jdff dff_A_DAZQY4LC8_1(.din(n3482), .dout(n3479));
    jdff dff_A_rxU9HR7l9_1(.din(n3485), .dout(n3482));
    jdff dff_A_NFzSnkBu4_1(.din(n3488), .dout(n3485));
    jdff dff_A_hzmtlQNW0_1(.din(n3491), .dout(n3488));
    jdff dff_A_XLbgnOm52_1(.din(n3494), .dout(n3491));
    jdff dff_A_TBEbmUIM3_1(.din(n3497), .dout(n3494));
    jdff dff_A_92L2Is1y1_1(.din(n3500), .dout(n3497));
    jdff dff_A_g1NKNY736_1(.din(n1029), .dout(n3500));
    jdff dff_A_9ojVpIRN3_1(.din(n3506), .dout(n3503));
    jdff dff_A_08R7Lev64_1(.din(n3509), .dout(n3506));
    jdff dff_A_WdjsqJVn3_1(.din(n3512), .dout(n3509));
    jdff dff_A_n8CJ7ICn0_1(.din(n3515), .dout(n3512));
    jdff dff_A_R8Vs0EG03_1(.din(n3518), .dout(n3515));
    jdff dff_A_mV0FOiNZ9_1(.din(n3521), .dout(n3518));
    jdff dff_A_CMxlevNE6_1(.din(n3524), .dout(n3521));
    jdff dff_A_RUTyJ0s48_1(.din(n3527), .dout(n3524));
    jdff dff_A_MM3tbpEL4_1(.din(n3530), .dout(n3527));
    jdff dff_A_l4Ds0gqY9_1(.din(n3533), .dout(n3530));
    jdff dff_A_GAhtxgvl0_1(.din(n1025), .dout(n3533));
    jdff dff_A_yf3Es2g00_0(.din(n3539), .dout(n3536));
    jdff dff_A_USrduznW5_0(.din(n3542), .dout(n3539));
    jdff dff_A_RyCpXcoG7_0(.din(n3545), .dout(n3542));
    jdff dff_A_RlEP8WcD4_0(.din(n3548), .dout(n3545));
    jdff dff_A_19Wqj0xR3_0(.din(n3551), .dout(n3548));
    jdff dff_A_LfoXiNxK0_0(.din(n3554), .dout(n3551));
    jdff dff_A_5l1pAPm48_0(.din(n3557), .dout(n3554));
    jdff dff_A_XRapL5ry9_0(.din(n3560), .dout(n3557));
    jdff dff_A_5UnxKDUu8_0(.din(G171gat), .dout(n3560));
    jdff dff_A_ppOcJGmE8_1(.din(n3566), .dout(n3563));
    jdff dff_A_pioUJZBQ7_1(.din(n3569), .dout(n3566));
    jdff dff_A_JYwpyw1R4_1(.din(n3572), .dout(n3569));
    jdff dff_A_Xyx0mOje4_1(.din(n3575), .dout(n3572));
    jdff dff_A_OzXuUR4n4_1(.din(n3578), .dout(n3575));
    jdff dff_A_4Fo6cjNh2_1(.din(n3581), .dout(n3578));
    jdff dff_A_TS9LzjdN2_1(.din(n3584), .dout(n3581));
    jdff dff_A_yrGGfm964_1(.din(n3587), .dout(n3584));
    jdff dff_A_SDHk0Ayh3_1(.din(G171gat), .dout(n3587));
    jdff dff_B_em656vaO0_1(.din(n1311), .dout(n3591));
    jdff dff_B_LNaa5wLb6_0(.din(n1331), .dout(n3594));
    jdff dff_B_6GQCrwjA3_0(.din(n3594), .dout(n3597));
    jdff dff_B_0VR8D4NB0_0(.din(n1323), .dout(n3600));
    jdff dff_B_LH3CBpk42_0(.din(n3600), .dout(n3603));
    jdff dff_B_Qr1Exhr47_0(.din(n3603), .dout(n3606));
    jdff dff_B_vXtvioYj5_0(.din(n3606), .dout(n3609));
    jdff dff_B_WNAWS9qW8_0(.din(n3609), .dout(n3612));
    jdff dff_B_BWDOHGqr9_0(.din(n3612), .dout(n3615));
    jdff dff_B_LAuNqCAH6_0(.din(n3615), .dout(n3618));
    jdff dff_B_ZlYS1TIf0_0(.din(n3618), .dout(n3621));
    jdff dff_B_8yfsx2nm3_0(.din(n3621), .dout(n3624));
    jdff dff_B_wTQ1267p5_0(.din(n3624), .dout(n3627));
    jdff dff_A_YiYdZcsI5_1(.din(n3632), .dout(n3629));
    jdff dff_A_lIdggpTg7_1(.din(n3635), .dout(n3632));
    jdff dff_A_Bx15hbLn1_1(.din(n3638), .dout(n3635));
    jdff dff_A_z2n6usdp9_1(.din(n3641), .dout(n3638));
    jdff dff_A_hHT4DfCN8_1(.din(n3644), .dout(n3641));
    jdff dff_A_pSUFoYvh7_1(.din(G91gat), .dout(n3644));
    jdff dff_A_BcMDqKgm5_1(.din(n3650), .dout(n3647));
    jdff dff_A_SCgwyVPp8_1(.din(n3653), .dout(n3650));
    jdff dff_A_86jZxEJm1_1(.din(n3656), .dout(n3653));
    jdff dff_A_iFAjw0GP6_1(.din(n3659), .dout(n3656));
    jdff dff_A_BvksVKM82_1(.din(n3662), .dout(n3659));
    jdff dff_A_zHL6klVf2_1(.din(n3665), .dout(n3662));
    jdff dff_A_ogtdX02Z2_1(.din(n3668), .dout(n3665));
    jdff dff_A_f7gAH5oF8_1(.din(n3671), .dout(n3668));
    jdff dff_A_lcXQg14O7_1(.din(n3674), .dout(n3671));
    jdff dff_A_FodcDkDs4_1(.din(n3677), .dout(n3674));
    jdff dff_A_JJoZkWO27_1(.din(n3680), .dout(n3677));
    jdff dff_A_Xa5F2hGi1_1(.din(n1315), .dout(n3680));
    jdff dff_B_py9DwAIB7_0(.din(n981), .dout(n3684));
    jdff dff_B_ME3aqBur3_0(.din(n977), .dout(n3687));
    jdff dff_B_FGhC9g0D4_0(.din(n3687), .dout(n3690));
    jdff dff_B_8IAzCC8t9_0(.din(n3690), .dout(n3693));
    jdff dff_B_sDlKO3YR9_0(.din(n3693), .dout(n3696));
    jdff dff_A_aNQIUORM4_0(.din(n3701), .dout(n3698));
    jdff dff_A_6ZGK6Eos5_0(.din(n937), .dout(n3701));
    jdff dff_A_f16D6L1E6_1(.din(n3707), .dout(n3704));
    jdff dff_A_VMDtzSMh3_1(.din(n3710), .dout(n3707));
    jdff dff_A_2H6Iw6yB7_1(.din(n3713), .dout(n3710));
    jdff dff_A_di2SfrFP5_1(.din(n3716), .dout(n3713));
    jdff dff_A_ugTcDXZo3_1(.din(n3719), .dout(n3716));
    jdff dff_A_ZzoTFIye8_1(.din(n3722), .dout(n3719));
    jdff dff_A_pfeKiM682_1(.din(n3725), .dout(n3722));
    jdff dff_A_D05oNxKZ1_1(.din(n3759), .dout(n3725));
    jdff dff_A_gV8tk6AY7_2(.din(n3731), .dout(n3728));
    jdff dff_A_FCaw76er3_2(.din(n3734), .dout(n3731));
    jdff dff_A_ZTSQR2WJ0_2(.din(n3737), .dout(n3734));
    jdff dff_A_6KPCu3Km9_2(.din(n3740), .dout(n3737));
    jdff dff_A_ItNotLYK3_2(.din(n3743), .dout(n3740));
    jdff dff_A_wwwFtVNb1_2(.din(n3746), .dout(n3743));
    jdff dff_A_38dpMtXr9_2(.din(n3749), .dout(n3746));
    jdff dff_A_md0ncrWr1_2(.din(n3752), .dout(n3749));
    jdff dff_A_BTy1ECCB1_2(.din(n3755), .dout(n3752));
    jdff dff_A_ZuaxcF6B6_2(.din(n3759), .dout(n3755));
    jdff dff_B_epr6vjWz6_3(.din(G165gat), .dout(n3759));
    jdff dff_B_TjZuYqWm5_1(.din(n1402), .dout(n3762));
    jdff dff_B_RQ8n5l5u4_1(.din(n3762), .dout(n3765));
    jdff dff_B_8YmqLXfr9_1(.din(n3765), .dout(n3768));
    jdff dff_B_SsrziKMG3_1(.din(n3768), .dout(n3771));
    jdff dff_B_9DIcCkY60_1(.din(n3771), .dout(n3774));
    jdff dff_B_nUPNL3Do2_1(.din(n3774), .dout(n3777));
    jdff dff_B_7T0nKnwn6_1(.din(n3777), .dout(n3780));
    jdff dff_B_Ypdj6s0X1_1(.din(n3780), .dout(n3783));
    jdff dff_B_lvNTZ2L67_1(.din(n3783), .dout(n3786));
    jdff dff_B_EwFU9vN70_1(.din(n1409), .dout(n3789));
    jdff dff_B_W3z3T0lt7_1(.din(n1070), .dout(n3792));
    jdff dff_B_YvFDfzdB1_1(.din(n3792), .dout(n3795));
    jdff dff_B_OXuQGpJw2_1(.din(n3795), .dout(n3798));
    jdff dff_B_6DpSRe6W7_1(.din(n3798), .dout(n3801));
    jdff dff_B_pcnzQFld0_1(.din(n3801), .dout(n3804));
    jdff dff_B_8Q9L2Ugr5_1(.din(n3804), .dout(n3807));
    jdff dff_B_GmmfPo5h3_1(.din(n1083), .dout(n3810));
    jdff dff_B_EY4aSTkf0_1(.din(n3810), .dout(n3813));
    jdff dff_B_yoby2iPW5_1(.din(n3813), .dout(n3816));
    jdff dff_B_id5kLjQl1_1(.din(n3816), .dout(n3819));
    jdff dff_B_vbu4v1jM8_1(.din(n3819), .dout(n3822));
    jdff dff_B_rl9Vq7JE8_0(.din(n412), .dout(n3825));
    jdff dff_A_rWOHNZkG3_1(.din(n3830), .dout(n3827));
    jdff dff_A_sqprAlgC0_1(.din(n3845), .dout(n3830));
    jdff dff_A_lslrCMJR3_2(.din(n3836), .dout(n3833));
    jdff dff_A_UUauDlHl2_2(.din(n3839), .dout(n3836));
    jdff dff_A_QObBHfh02_2(.din(n3842), .dout(n3839));
    jdff dff_A_4Sd4npID9_2(.din(n3845), .dout(n3842));
    jdff dff_A_O1Lucx3I5_0(.din(n3848), .dout(n3845));
    jdff dff_A_uzqWPfXI1_0(.din(n3851), .dout(n3848));
    jdff dff_A_a1FPNMpL1_0(.din(n3854), .dout(n3851));
    jdff dff_A_asF04T9x1_0(.din(n3857), .dout(n3854));
    jdff dff_A_edw16gTV5_0(.din(n3860), .dout(n3857));
    jdff dff_A_kOUkT3XB5_0(.din(n3863), .dout(n3860));
    jdff dff_A_jtlU4Qz41_0(.din(n3866), .dout(n3863));
    jdff dff_A_yV2b8S5z8_0(.din(n3869), .dout(n3866));
    jdff dff_A_SfnO8thz7_0(.din(n3909), .dout(n3869));
    jdff dff_A_sMiNjPDH1_1(.din(n3909), .dout(n3872));
    jdff dff_B_PLaI4vFA4_3(.din(G219gat), .dout(n3876));
    jdff dff_B_UIDBElnm6_3(.din(n3876), .dout(n3879));
    jdff dff_B_wqnAYARH5_3(.din(n3879), .dout(n3882));
    jdff dff_B_BfeD4erD1_3(.din(n3882), .dout(n3885));
    jdff dff_B_R9hstALJ1_3(.din(n3885), .dout(n3888));
    jdff dff_B_o3Pi5RmB4_3(.din(n3888), .dout(n3891));
    jdff dff_B_ptPcvAMe1_3(.din(n3891), .dout(n3894));
    jdff dff_B_q7NuIUaE4_3(.din(n3894), .dout(n3897));
    jdff dff_B_2xljmZZE0_3(.din(n3897), .dout(n3900));
    jdff dff_B_R3Xi5MM07_3(.din(n3900), .dout(n3903));
    jdff dff_B_cexpfoTi9_3(.din(n3903), .dout(n3906));
    jdff dff_B_kEi3TNjC8_3(.din(n3906), .dout(n3909));
    jdff dff_B_9wLbiQPo5_0(.din(n1405), .dout(n3912));
    jdff dff_B_KjaHok4l3_0(.din(n3912), .dout(n3915));
    jdff dff_B_CgkK8ZDX5_0(.din(n3915), .dout(n3918));
    jdff dff_B_cvEIrjfx2_0(.din(n3918), .dout(n3921));
    jdff dff_B_onPodhm80_0(.din(n3921), .dout(n3924));
    jdff dff_B_csD3o8sT0_0(.din(n3924), .dout(n3927));
    jdff dff_B_TnQ6bYOD9_0(.din(n3927), .dout(n3930));
    jdff dff_B_WB2r8z254_0(.din(n3930), .dout(n3933));
    jdff dff_B_bOfGwb3m3_0(.din(n3933), .dout(n3936));
    jdff dff_B_WSMxIz7D4_1(.din(n1256), .dout(n3939));
    jdff dff_B_xeCAAGe97_1(.din(n3939), .dout(n3942));
    jdff dff_B_wPr6t00I9_1(.din(n3942), .dout(n3945));
    jdff dff_B_oQvKxCeK5_1(.din(n3945), .dout(n3948));
    jdff dff_B_rBwTdNrd7_1(.din(n3948), .dout(n3951));
    jdff dff_B_MIa4ORsT9_1(.din(n3951), .dout(n3954));
    jdff dff_B_eALyMLm19_1(.din(n3954), .dout(n3957));
    jdff dff_B_9YbA9GZ99_1(.din(n3957), .dout(n3960));
    jdff dff_B_2niJCX933_1(.din(n1141), .dout(n3963));
    jdff dff_B_2tdBkyD23_1(.din(n3963), .dout(n3966));
    jdff dff_B_L7mGhCgb8_1(.din(n3966), .dout(n3969));
    jdff dff_B_YBwhKsRa3_1(.din(n3969), .dout(n3972));
    jdff dff_B_NjjmpL1C0_1(.din(n3972), .dout(n3975));
    jdff dff_B_axRcZCmb1_1(.din(n3975), .dout(n3978));
    jdff dff_B_Y9ex9KpT5_1(.din(n3978), .dout(n3981));
    jdff dff_B_qKC3uJD64_1(.din(n726), .dout(n3984));
    jdff dff_B_VXLgkgsg4_1(.din(n3984), .dout(n3987));
    jdff dff_B_IGXkI59T7_1(.din(n3987), .dout(n3990));
    jdff dff_B_ZEdnkMpZ5_1(.din(n3990), .dout(n3993));
    jdff dff_B_XRitnMuY1_1(.din(n3993), .dout(n3996));
    jdff dff_B_BjzQLaOI5_1(.din(n729), .dout(n3999));
    jdff dff_B_YfHJEGy66_1(.din(n3999), .dout(n4002));
    jdff dff_B_EXS4HU1R9_1(.din(n4002), .dout(n4005));
    jdff dff_B_a0X6tw2p1_1(.din(n4005), .dout(n4008));
    jdff dff_B_LVXLDEJp9_1(.din(n732), .dout(n4011));
    jdff dff_B_5z8THAnV5_1(.din(n4011), .dout(n4014));
    jdff dff_B_E84IDsFC6_1(.din(n4014), .dout(n4017));
    jdff dff_B_a8bqaFgB0_1(.din(n735), .dout(n4020));
    jdff dff_B_E40CS4Av2_1(.din(n4020), .dout(n4023));
    jdff dff_A_r3WANGgp2_1(.din(n4053), .dout(n4025));
    jdff dff_B_TcBGh5e38_2(.din(n558), .dout(n4029));
    jdff dff_B_GZI1XtSJ9_2(.din(n4029), .dout(n4032));
    jdff dff_B_qJeypqZ09_2(.din(n4032), .dout(n4035));
    jdff dff_B_GdrfCwyA0_2(.din(n4035), .dout(n4038));
    jdff dff_B_gjPcV6FL6_2(.din(n4038), .dout(n4041));
    jdff dff_B_Od2j9ylF8_2(.din(n4041), .dout(n4044));
    jdff dff_B_hmAaJchv4_2(.din(n4044), .dout(n4047));
    jdff dff_B_yM4KmRWJ9_2(.din(n4047), .dout(n4050));
    jdff dff_B_OnztqHNG8_2(.din(n4050), .dout(n4053));
    jdff dff_A_3MnImfhx0_0(.din(n4058), .dout(n4055));
    jdff dff_A_hbDEDvy40_0(.din(n4061), .dout(n4058));
    jdff dff_A_96Mgs9Aq8_0(.din(n4064), .dout(n4061));
    jdff dff_A_URHxRA7b2_0(.din(n4067), .dout(n4064));
    jdff dff_A_5gUO1yCr0_0(.din(n4070), .dout(n4067));
    jdff dff_A_LAyl2Q3X3_0(.din(n4073), .dout(n4070));
    jdff dff_A_AhYmlxv09_0(.din(n4076), .dout(n4073));
    jdff dff_A_dGt58nX79_0(.din(n4079), .dout(n4076));
    jdff dff_A_GVhlbfMO6_0(.din(n4082), .dout(n4079));
    jdff dff_A_ccCzQTdh6_0(.din(G261gat), .dout(n4082));
    jdff dff_A_xhCMx9Wp1_2(.din(n4088), .dout(n4085));
    jdff dff_A_gQCTnKEc5_2(.din(n4091), .dout(n4088));
    jdff dff_A_Oo3s6GkZ7_2(.din(n4094), .dout(n4091));
    jdff dff_A_Utk7lrqA7_2(.din(n4097), .dout(n4094));
    jdff dff_A_HNm7eEoG8_2(.din(n4100), .dout(n4097));
    jdff dff_A_zV5pQmm24_2(.din(n4103), .dout(n4100));
    jdff dff_A_mPWFUcQR4_2(.din(n4106), .dout(n4103));
    jdff dff_A_QeE2dAfw5_2(.din(n4109), .dout(n4106));
    jdff dff_A_GcNMlFBW8_2(.din(n4112), .dout(n4109));
    jdff dff_A_TBAA5QPO6_2(.din(G261gat), .dout(n4112));
    jdff dff_A_DB211iR03_0(.din(n689), .dout(n4115));
    jdff dff_B_f9PFycb75_1(.din(n454), .dout(n4119));
    jdff dff_B_02REkNbb6_1(.din(n487), .dout(n4122));
    jdff dff_B_y2AXDNAR1_1(.din(n4122), .dout(n4125));
    jdff dff_B_7CUkmzZD5_1(.din(n4125), .dout(n4128));
    jdff dff_B_ObvjXfyc0_1(.din(n4128), .dout(n4131));
    jdff dff_B_kvx6MqsJ7_1(.din(n4131), .dout(n4134));
    jdff dff_B_HnluH0Uh6_1(.din(n457), .dout(n4137));
    jdff dff_B_901NAY6l2_1(.din(n4137), .dout(n4140));
    jdff dff_B_XmavlbES5_1(.din(n4140), .dout(n4143));
    jdff dff_B_hKw61krO9_1(.din(n4143), .dout(n4146));
    jdff dff_B_jn0YtmUD9_1(.din(n4146), .dout(n4149));
    jdff dff_B_BJriCuaR1_1(.din(n460), .dout(n4152));
    jdff dff_A_dU3YKqVA4_1(.din(n4157), .dout(n4154));
    jdff dff_A_7iacd3fw9_1(.din(n4160), .dout(n4157));
    jdff dff_A_HyAzXTRm3_1(.din(n4163), .dout(n4160));
    jdff dff_A_7HQPvZec9_1(.din(n4166), .dout(n4163));
    jdff dff_A_RGLzaIRm5_1(.din(n4169), .dout(n4166));
    jdff dff_A_IxPp00Gn2_1(.din(G126gat), .dout(n4169));
    jdff dff_B_0z4F70Dg9_3(.din(n451), .dout(n4173));
    jdff dff_B_Ythl7dYS6_3(.din(n4173), .dout(n4176));
    jdff dff_B_WZmIcOnv1_3(.din(n4176), .dout(n4179));
    jdff dff_B_xcZpoV7G9_3(.din(n4179), .dout(n4182));
    jdff dff_B_Mh9Rh9t26_3(.din(n4182), .dout(n4185));
    jdff dff_B_AyRVInel9_3(.din(n4185), .dout(n4188));
    jdff dff_B_zrgDDyU05_3(.din(n4188), .dout(n4191));
    jdff dff_B_juyi9VzG8_3(.din(n4191), .dout(n4194));
    jdff dff_A_WAOntSsh3_1(.din(n4199), .dout(n4196));
    jdff dff_A_PKGxXbie3_1(.din(n4202), .dout(n4199));
    jdff dff_A_SnGcm0yV3_1(.din(n4205), .dout(n4202));
    jdff dff_A_eT09wCdN9_1(.din(n4208), .dout(n4205));
    jdff dff_A_lyUuIx8R6_1(.din(n4211), .dout(n4208));
    jdff dff_A_9ZGB39M65_1(.din(n4214), .dout(n4211));
    jdff dff_A_VkU8dekx9_1(.din(n4217), .dout(n4214));
    jdff dff_A_25R4wEmD7_1(.din(n4220), .dout(n4217));
    jdff dff_A_DVUZWOLC3_1(.din(G201gat), .dout(n4220));
    jdff dff_A_ZsvT9tFg9_1(.din(n4226), .dout(n4223));
    jdff dff_A_vnB3XQGd9_1(.din(n4229), .dout(n4226));
    jdff dff_A_HtD9ivyS4_1(.din(n685), .dout(n4229));
    jdff dff_A_X388gADN1_1(.din(n4235), .dout(n4232));
    jdff dff_A_nFZrfz888_1(.din(n4238), .dout(n4235));
    jdff dff_A_75Z0Ttk17_1(.din(n4241), .dout(n4238));
    jdff dff_A_JkpUGZBf2_1(.din(n4244), .dout(n4241));
    jdff dff_A_Piy7sRBc7_1(.din(n4247), .dout(n4244));
    jdff dff_A_bI3C978E9_1(.din(n4250), .dout(n4247));
    jdff dff_A_DZOh1sNt7_1(.din(n4253), .dout(n4250));
    jdff dff_A_TKBNZ3Sl1_1(.din(G195gat), .dout(n4253));
    jdff dff_A_oB8wX8y63_2(.din(n4259), .dout(n4256));
    jdff dff_A_KD6KpCBg7_2(.din(n4262), .dout(n4259));
    jdff dff_A_TyLearqF5_2(.din(n4265), .dout(n4262));
    jdff dff_A_dHwoZXZW7_2(.din(n4268), .dout(n4265));
    jdff dff_A_GldfbQnw1_2(.din(n4271), .dout(n4268));
    jdff dff_A_YhlLimJq7_2(.din(n4274), .dout(n4271));
    jdff dff_A_0L2Xkrqe9_2(.din(n4277), .dout(n4274));
    jdff dff_A_FKwPJQjV2_2(.din(G195gat), .dout(n4277));
    jdff dff_A_RcHTt1r62_1(.din(n4283), .dout(n4280));
    jdff dff_A_Q4NqfTz41_1(.din(n4286), .dout(n4283));
    jdff dff_A_LfhSIsyo9_1(.din(n4289), .dout(n4286));
    jdff dff_A_P4zV80J80_1(.din(n681), .dout(n4289));
    jdff dff_A_zB6Gv0j14_0(.din(n4295), .dout(n4292));
    jdff dff_A_4TbRHPQ64_0(.din(n4298), .dout(n4295));
    jdff dff_A_K2ZbbhQx8_0(.din(n4301), .dout(n4298));
    jdff dff_A_DGPwAcHs4_0(.din(n4304), .dout(n4301));
    jdff dff_A_PdUsLsWK7_0(.din(n4307), .dout(n4304));
    jdff dff_A_2O2Q4pOl4_0(.din(G121gat), .dout(n4307));
    jdff dff_A_4e58sPPQ2_0(.din(n4313), .dout(n4310));
    jdff dff_A_vAJMRL0o8_0(.din(n4316), .dout(n4313));
    jdff dff_A_e8keUhLf1_0(.din(n4319), .dout(n4316));
    jdff dff_A_yBKCEkH24_0(.din(n4322), .dout(n4319));
    jdff dff_A_XjCVYkKl7_0(.din(n4325), .dout(n4322));
    jdff dff_A_SKoyFyBL6_0(.din(n4328), .dout(n4325));
    jdff dff_A_a1EvICEe9_0(.din(n4331), .dout(n4328));
    jdff dff_A_gzSCnwQh6_0(.din(G195gat), .dout(n4331));
    jdff dff_A_58KEmVE42_2(.din(n4337), .dout(n4334));
    jdff dff_A_Gz0ZKhMP3_2(.din(n4340), .dout(n4337));
    jdff dff_A_hsRqyjQF2_2(.din(n4343), .dout(n4340));
    jdff dff_A_7I1OU8ZZ1_2(.din(G195gat), .dout(n4343));
    jdff dff_A_HQIrl6Va9_1(.din(n4349), .dout(n4346));
    jdff dff_A_T7BVjZmB1_1(.din(n4352), .dout(n4349));
    jdff dff_A_KorqsZZp3_1(.din(n4355), .dout(n4352));
    jdff dff_A_KtvHNEcG6_1(.din(n4358), .dout(n4355));
    jdff dff_A_CB2CKF6I5_1(.din(n661), .dout(n4358));
    jdff dff_A_H6T3bKCf7_1(.din(n4364), .dout(n4361));
    jdff dff_A_68Es0FZV4_1(.din(n4367), .dout(n4364));
    jdff dff_A_iIdqfS259_1(.din(n4370), .dout(n4367));
    jdff dff_A_mW1Fgj0O8_1(.din(n4373), .dout(n4370));
    jdff dff_A_panc784W4_1(.din(n4376), .dout(n4373));
    jdff dff_A_mkV3RWMw8_1(.din(n4379), .dout(n4376));
    jdff dff_A_0RWsyMFv1_1(.din(n4382), .dout(n4379));
    jdff dff_A_JQ4JKKZN3_1(.din(G189gat), .dout(n4382));
    jdff dff_A_3kGgvMV84_2(.din(n4388), .dout(n4385));
    jdff dff_A_gFPaDQdq1_2(.din(n4391), .dout(n4388));
    jdff dff_A_zjrh4Zhi9_2(.din(n4394), .dout(n4391));
    jdff dff_A_N1dGASNL1_2(.din(n4397), .dout(n4394));
    jdff dff_A_Qeh2TP0d5_2(.din(n4400), .dout(n4397));
    jdff dff_A_TiRiaqpM7_2(.din(n4403), .dout(n4400));
    jdff dff_A_fJHNsO0G1_2(.din(n4406), .dout(n4403));
    jdff dff_A_BONYvIGV9_2(.din(G189gat), .dout(n4406));
    jdff dff_A_biPzaajY5_1(.din(n4412), .dout(n4409));
    jdff dff_A_CdGEj5VR7_1(.din(n4415), .dout(n4412));
    jdff dff_A_xeuZn17I5_1(.din(n4418), .dout(n4415));
    jdff dff_A_UucWkXq47_1(.din(n4421), .dout(n4418));
    jdff dff_A_3lnmUeB01_1(.din(n4424), .dout(n4421));
    jdff dff_A_k3roUDba9_1(.din(n657), .dout(n4424));
    jdff dff_A_RgrZBGyU8_1(.din(n4440), .dout(n4427));
    jdff dff_B_43DQC57i3_2(.din(G146gat), .dout(n4431));
    jdff dff_B_XqQFUiyg4_2(.din(n4431), .dout(n4434));
    jdff dff_B_dQhxHCWz2_2(.din(n4434), .dout(n4437));
    jdff dff_B_ELVxRGg83_2(.din(n4437), .dout(n4440));
    jdff dff_A_6nBN1ogq9_1(.din(n4445), .dout(n4442));
    jdff dff_A_ROKh5EhK0_1(.din(n4448), .dout(n4445));
    jdff dff_A_1kIFFkiw8_1(.din(n4451), .dout(n4448));
    jdff dff_A_gw22SdBI6_1(.din(n4454), .dout(n4451));
    jdff dff_A_cYPOGd2v4_1(.din(n4457), .dout(n4454));
    jdff dff_A_d6biRXab9_1(.din(G116gat), .dout(n4457));
    jdff dff_A_CRKecSso3_0(.din(n4463), .dout(n4460));
    jdff dff_A_T6ccq5hL7_0(.din(n4466), .dout(n4463));
    jdff dff_A_p5d4la7a7_0(.din(n4469), .dout(n4466));
    jdff dff_A_J9Wi2rGg5_0(.din(n4472), .dout(n4469));
    jdff dff_A_Yf6uo45Z9_0(.din(n4475), .dout(n4472));
    jdff dff_A_xCZKXQlo2_0(.din(n4478), .dout(n4475));
    jdff dff_A_6wM7kc4N2_0(.din(n4481), .dout(n4478));
    jdff dff_A_15PxcqHD1_0(.din(G189gat), .dout(n4481));
    jdff dff_A_zOXzmiA46_2(.din(n4487), .dout(n4484));
    jdff dff_A_ptCLX6vO7_2(.din(n4490), .dout(n4487));
    jdff dff_A_IKVk7OZN7_2(.din(n4493), .dout(n4490));
    jdff dff_A_OWu9GO5M9_2(.din(G189gat), .dout(n4493));
    jdff dff_A_EGJT6SzF8_0(.din(n4499), .dout(n4496));
    jdff dff_A_vpcGVEZ13_0(.din(n4502), .dout(n4499));
    jdff dff_A_zljUsMXi2_0(.din(n4505), .dout(n4502));
    jdff dff_A_DdnYctoD0_0(.din(n4508), .dout(n4505));
    jdff dff_A_wAhB5Dpr9_0(.din(n4511), .dout(n4508));
    jdff dff_A_SfACn2Ng8_0(.din(n1080), .dout(n4511));
    jdff dff_B_17GVwLMI4_1(.din(n1073), .dout(n4515));
    jdff dff_B_NXo4Vcax5_1(.din(n4515), .dout(n4518));
    jdff dff_B_pklLYb6D2_1(.din(n4518), .dout(n4521));
    jdff dff_B_zMH2pYu61_1(.din(n4521), .dout(n4524));
    jdff dff_B_Xnfmz8m85_1(.din(n4524), .dout(n4527));
    jdff dff_B_IsHlgTDw1_1(.din(n4527), .dout(n4530));
    jdff dff_B_rYhg64yR0_1(.din(n4530), .dout(n4533));
    jdff dff_B_THrVAbF30_1(.din(n4533), .dout(n4536));
    jdff dff_A_7s7pj6yq6_1(.din(n4541), .dout(n4538));
    jdff dff_A_4CdHw3xI2_1(.din(n4544), .dout(n4541));
    jdff dff_A_IKaGLcQx4_1(.din(n4547), .dout(n4544));
    jdff dff_A_yX7WiixN2_1(.din(n4550), .dout(n4547));
    jdff dff_A_w0TsZFF95_1(.din(n4553), .dout(n4550));
    jdff dff_A_hFE75WfB3_1(.din(n4556), .dout(n4553));
    jdff dff_A_QCIoRFPs4_1(.din(n4559), .dout(n4556));
    jdff dff_A_uyfWmlS52_1(.din(n609), .dout(n4559));
    jdff dff_A_nQJVdCYi2_0(.din(n4565), .dout(n4562));
    jdff dff_A_QqjlHKmk1_0(.din(n4568), .dout(n4565));
    jdff dff_A_6GAsQtzw5_0(.din(n130), .dout(n4568));
    jdff dff_A_PH8TGeuR4_1(.din(n4584), .dout(n4571));
    jdff dff_B_ckQ37O4F2_2(.din(G143gat), .dout(n4575));
    jdff dff_B_tJWrjoTV0_2(.din(n4575), .dout(n4578));
    jdff dff_B_pvufKJtW7_2(.din(n4578), .dout(n4581));
    jdff dff_B_65QB3twe0_2(.din(n4581), .dout(n4584));
    jdff dff_A_x0AiMJPD2_2(.din(n4589), .dout(n4586));
    jdff dff_A_yVEYHzL20_2(.din(n326), .dout(n4589));
    jdff dff_A_zd94hS645_1(.din(n4595), .dout(n4592));
    jdff dff_A_XFB29Rx80_1(.din(n4598), .dout(n4595));
    jdff dff_A_0ss6Ng1O9_1(.din(n4601), .dout(n4598));
    jdff dff_A_z2blFpm61_1(.din(n4604), .dout(n4601));
    jdff dff_A_bjp8xU1K8_1(.din(n4607), .dout(n4604));
    jdff dff_A_cThWVYcY6_1(.din(G111gat), .dout(n4607));
    jdff dff_A_QqaogmRE3_2(.din(n4613), .dout(n4610));
    jdff dff_A_gRlOYoRF9_2(.din(n4616), .dout(n4613));
    jdff dff_A_0EMUVmRj6_2(.din(n4619), .dout(n4616));
    jdff dff_A_soEfiLC39_2(.din(n4622), .dout(n4619));
    jdff dff_A_RJlScyza6_2(.din(n4625), .dout(n4622));
    jdff dff_A_pOLLdz346_2(.din(n4628), .dout(n4625));
    jdff dff_A_3Cz6OzwJ3_2(.din(n4631), .dout(n4628));
    jdff dff_A_54e5qKsY5_2(.din(G183gat), .dout(n4631));
    jdff dff_A_w73sto869_0(.din(n4637), .dout(n4634));
    jdff dff_A_pwpjSjNC8_0(.din(n4640), .dout(n4637));
    jdff dff_A_paMU3kcr5_0(.din(n4643), .dout(n4640));
    jdff dff_A_DhIYGIoK8_0(.din(n4646), .dout(n4643));
    jdff dff_A_zFIWgomP6_0(.din(n4649), .dout(n4646));
    jdff dff_A_p742Ppg74_0(.din(n4652), .dout(n4649));
    jdff dff_A_lyr1kNRw7_0(.din(n1067), .dout(n4652));
    jdff dff_B_BHrdnGlM6_1(.din(n1060), .dout(n4656));
    jdff dff_B_GWM0xa6L8_1(.din(n4656), .dout(n4659));
    jdff dff_B_T713Ti4e7_1(.din(n4659), .dout(n4662));
    jdff dff_B_2JnXiDwJ0_1(.din(n4662), .dout(n4665));
    jdff dff_B_j8ejU5395_1(.din(n4665), .dout(n4668));
    jdff dff_B_1BnI7T5Q0_1(.din(n4668), .dout(n4671));
    jdff dff_B_TBWOYx9H7_1(.din(n4671), .dout(n4674));
    jdff dff_B_GQdyiRzL9_1(.din(n4674), .dout(n4677));
    jdff dff_B_zRWcyhoV2_1(.din(n4677), .dout(n4680));
    jdff dff_A_iaarpLbz1_2(.din(n4685), .dout(n4682));
    jdff dff_A_aeWtvHSd9_2(.din(n4688), .dout(n4685));
    jdff dff_A_siMNGYZJ1_2(.din(n4691), .dout(n4688));
    jdff dff_A_szMHMi966_2(.din(n4694), .dout(n4691));
    jdff dff_A_j8R3cMdQ2_2(.din(n4697), .dout(n4694));
    jdff dff_A_DPPJxwXO3_2(.din(n4700), .dout(n4697));
    jdff dff_A_qyfsu4mV1_2(.din(n4703), .dout(n4700));
    jdff dff_A_wzlfTpSR4_2(.din(n4706), .dout(n4703));
    jdff dff_A_SexcC3WA1_2(.din(n1057), .dout(n4706));
    jdff dff_B_6GSYaz0e9_0(.din(n1045), .dout(n4710));
    jdff dff_B_XR90HrZC3_0(.din(n1041), .dout(n4713));
    jdff dff_B_eOwpGUK18_0(.din(n4713), .dout(n4716));
    jdff dff_B_4eSsaiJV7_0(.din(n4716), .dout(n4719));
    jdff dff_B_Kn1FYWoV5_0(.din(n4719), .dout(n4722));
    jdff dff_A_X3qLaOM47_0(.din(n4727), .dout(n4724));
    jdff dff_A_2meL8y736_0(.din(n4730), .dout(n4727));
    jdff dff_A_64HgHN3Q9_0(.din(n4733), .dout(n4730));
    jdff dff_A_fWbf8oFC2_0(.din(G153gat), .dout(n4733));
    jdff dff_A_1tJh7omA6_2(.din(n4739), .dout(n4736));
    jdff dff_A_wqRgMnMr2_2(.din(n4742), .dout(n4739));
    jdff dff_A_cKVQ8j5j7_2(.din(n4745), .dout(n4742));
    jdff dff_A_1Sr3NbGH3_2(.din(n4748), .dout(n4745));
    jdff dff_A_kiWkekqw1_2(.din(G153gat), .dout(n4748));
    jdff dff_A_CUbpgPGn2_0(.din(n4754), .dout(n4751));
    jdff dff_A_s3zAHzsd5_0(.din(n4757), .dout(n4754));
    jdff dff_A_eB2W1GEJ3_0(.din(n4760), .dout(n4757));
    jdff dff_A_c2a3JZsZ6_0(.din(n4763), .dout(n4760));
    jdff dff_A_6EYbj9qD5_0(.din(n4766), .dout(n4763));
    jdff dff_A_URmQRko84_0(.din(G106gat), .dout(n4766));
    jdff dff_A_jwCTRDKo0_1(.din(n4772), .dout(n4769));
    jdff dff_A_KHqIG8Ny1_1(.din(n4775), .dout(n4772));
    jdff dff_A_l7HuiG969_1(.din(n4778), .dout(n4775));
    jdff dff_A_1Tv02Wh29_1(.din(n4781), .dout(n4778));
    jdff dff_A_HJjv8p6k1_1(.din(n4784), .dout(n4781));
    jdff dff_A_5rAKIP7Z4_1(.din(n4787), .dout(n4784));
    jdff dff_A_eAq0ZszF3_1(.din(n4790), .dout(n4787));
    jdff dff_A_Tfb3Se8u8_1(.din(n4793), .dout(n4790));
    jdff dff_A_NT7xUXH68_1(.din(G177gat), .dout(n4793));
    jdff dff_A_ST8w2acz9_1(.din(n4799), .dout(n4796));
    jdff dff_A_Zlcc1WBo6_1(.din(n4802), .dout(n4799));
    jdff dff_A_R26fKNaK3_1(.din(n4805), .dout(n4802));
    jdff dff_A_VewlEDL70_1(.din(G177gat), .dout(n4805));
    jdff dff_A_yyUdDatr8_2(.din(n4811), .dout(n4808));
    jdff dff_A_KgHjpYpx2_2(.din(n4814), .dout(n4811));
    jdff dff_A_WLRj8K4X0_2(.din(n4817), .dout(n4814));
    jdff dff_A_h308vyhu8_2(.din(n4820), .dout(n4817));
    jdff dff_A_j7fqDAxq3_2(.din(n4823), .dout(n4820));
    jdff dff_A_C8L4BNUS5_2(.din(n4826), .dout(n4823));
    jdff dff_A_nYV1IXK00_2(.din(n4829), .dout(n4826));
    jdff dff_A_sX7oZQmF4_2(.din(n4832), .dout(n4829));
    jdff dff_A_eyk3KoDE9_2(.din(G177gat), .dout(n4832));
    jdff dff_B_9BWndEVS6_1(.din(n1374), .dout(n4836));
    jdff dff_B_JDVZwhDt8_0(.din(n1394), .dout(n4839));
    jdff dff_B_guRjmfLS2_0(.din(n4839), .dout(n4842));
    jdff dff_A_YoFWnBwt3_0(.din(n4847), .dout(n4844));
    jdff dff_A_d1HhWs9R1_0(.din(n4850), .dout(n4847));
    jdff dff_A_jYjxtVsY3_0(.din(n4853), .dout(n4850));
    jdff dff_A_fIGaozpt2_0(.din(n4856), .dout(n4853));
    jdff dff_A_sv7ef6nn8_0(.din(n4859), .dout(n4856));
    jdff dff_A_uvliav676_0(.din(n4862), .dout(n4859));
    jdff dff_A_Bm7VBKl85_0(.din(n4865), .dout(n4862));
    jdff dff_A_pRmQpTHG9_0(.din(n4890), .dout(n4865));
    jdff dff_A_v2wpW7I60_2(.din(n4871), .dout(n4868));
    jdff dff_A_HYAAvPMU0_2(.din(n4874), .dout(n4871));
    jdff dff_A_q812jhGF1_2(.din(n4877), .dout(n4874));
    jdff dff_A_wYIuQO3E2_2(.din(n4880), .dout(n4877));
    jdff dff_A_6yWhX6pT4_2(.din(n4883), .dout(n4880));
    jdff dff_A_8823zXGq1_2(.din(n4886), .dout(n4883));
    jdff dff_A_zoxLnd2T6_2(.din(n4890), .dout(n4886));
    jdff dff_B_FbsYManE5_3(.din(G246gat), .dout(n4890));
    jdff dff_B_tPbzwCid2_0(.din(n1386), .dout(n4893));
    jdff dff_B_DkZqUcE39_0(.din(n4893), .dout(n4896));
    jdff dff_B_iyOm5jen4_0(.din(n4896), .dout(n4899));
    jdff dff_B_fJz966m29_0(.din(n4899), .dout(n4902));
    jdff dff_B_0xpvP6Sy8_0(.din(n4902), .dout(n4905));
    jdff dff_B_yzzNuLNe8_0(.din(n4905), .dout(n4908));
    jdff dff_B_auaD2fl65_0(.din(n4908), .dout(n4911));
    jdff dff_B_HS5mRapg2_0(.din(n4911), .dout(n4914));
    jdff dff_B_spCLzmLV8_0(.din(n4914), .dout(n4917));
    jdff dff_B_q5Ktwy8s3_0(.din(n4917), .dout(n4920));
    jdff dff_A_SqO57Zob2_1(.din(n4925), .dout(n4922));
    jdff dff_A_sCOXXYkL6_1(.din(n4928), .dout(n4925));
    jdff dff_A_JhEi1HTD5_1(.din(n4931), .dout(n4928));
    jdff dff_A_ENmqCqTt3_1(.din(n4934), .dout(n4931));
    jdff dff_A_6TrxxOM32_1(.din(n4937), .dout(n4934));
    jdff dff_A_i58d2qx50_1(.din(G96gat), .dout(n4937));
    jdff dff_A_WBLbT3Mu9_0(.din(n4943), .dout(n4940));
    jdff dff_A_3b3TYrUP1_0(.din(n4946), .dout(n4943));
    jdff dff_A_jiIgGLHY5_0(.din(n4949), .dout(n4946));
    jdff dff_A_CjbDfE3e9_0(.din(n4952), .dout(n4949));
    jdff dff_A_cODPshmq1_0(.din(n4955), .dout(n4952));
    jdff dff_A_JDBYFYWt7_0(.din(n4958), .dout(n4955));
    jdff dff_A_e6nOEHk31_0(.din(n4961), .dout(n4958));
    jdff dff_A_HOXSNJxj9_0(.din(n4964), .dout(n4961));
    jdff dff_A_oeP4XS5h4_0(.din(n4967), .dout(n4964));
    jdff dff_A_H1gPzLXb4_0(.din(n1378), .dout(n4967));
    jdff dff_A_HlfwhfIe3_0(.din(n4998), .dout(n4970));
    jdff dff_B_WkQ1Z08U2_3(.din(G228gat), .dout(n4974));
    jdff dff_B_yj19BfzW4_3(.din(n4974), .dout(n4977));
    jdff dff_B_jcyjnR323_3(.din(n4977), .dout(n4980));
    jdff dff_B_9P6gXs5P0_3(.din(n4980), .dout(n4983));
    jdff dff_B_Jlkm723F3_3(.din(n4983), .dout(n4986));
    jdff dff_B_vFDnUJ2v2_3(.din(n4986), .dout(n4989));
    jdff dff_B_aw3uN2ng6_3(.din(n4989), .dout(n4992));
    jdff dff_B_MkHlyEnr7_3(.din(n4992), .dout(n4995));
    jdff dff_B_QR0EmBkX8_3(.din(n4995), .dout(n4998));
    jdff dff_B_s45QQpiD1_0(.din(n1013), .dout(n5001));
    jdff dff_B_Uv6o4uxD1_0(.din(n1009), .dout(n5004));
    jdff dff_B_ZJXg71DB7_0(.din(n5004), .dout(n5007));
    jdff dff_B_nqHDBrNL8_0(.din(n5007), .dout(n5010));
    jdff dff_B_QzdtIJtd4_0(.din(n5010), .dout(n5013));
    jdff dff_A_VIBDWbqU0_1(.din(n5028), .dout(n5015));
    jdff dff_B_jGyfQp2c6_2(.din(G149gat), .dout(n5019));
    jdff dff_B_aJ6kLBXZ2_2(.din(n5019), .dout(n5022));
    jdff dff_B_ZvYqvzJP6_2(.din(n5022), .dout(n5025));
    jdff dff_B_rozhVQNP3_2(.din(n5025), .dout(n5028));
    jdff dff_A_3dL30TBv8_0(.din(n378), .dout(n5030));
    jdff dff_B_XXbV3zQw3_1(.din(n359), .dout(n5034));
    jdff dff_B_hMdlKyK58_1(.din(n333), .dout(n5037));
    jdff dff_A_cSLTPijy3_0(.din(n341), .dout(n5039));
    jdff dff_A_srPCK7nJ5_0(.din(n5046), .dout(n5042));
    jdff dff_B_Yh1MOgGx9_2(.din(n337), .dout(n5046));
    jdff dff_A_O39kA17A9_0(.din(n5051), .dout(n5048));
    jdff dff_A_H2GZtF6F1_0(.din(n330), .dout(n5051));
    jdff dff_A_FcRWR8m76_1(.din(n180), .dout(n5054));
    jdff dff_A_7Xsqoc8r5_0(.din(G42gat), .dout(n5057));
    jdff dff_A_vFzjVfJl1_0(.din(n5063), .dout(n5060));
    jdff dff_A_CJ6pJ0Sd6_0(.din(n5066), .dout(n5063));
    jdff dff_A_883qTqWJ8_0(.din(n124), .dout(n5066));
    jdff dff_A_RYpoHz774_2(.din(n5072), .dout(n5069));
    jdff dff_A_SWS8zYQ67_2(.din(n124), .dout(n5072));
    jdff dff_A_BJqiOklz3_2(.din(n5078), .dout(n5075));
    jdff dff_A_uzkzW8UG4_2(.din(G17gat), .dout(n5078));
    jdff dff_A_QNvHU31e7_1(.din(n5084), .dout(n5081));
    jdff dff_A_Q8n0dWw79_1(.din(n5087), .dout(n5084));
    jdff dff_A_7H4wQV9e9_1(.din(n5090), .dout(n5087));
    jdff dff_A_T9ZOG8LW8_1(.din(n5093), .dout(n5090));
    jdff dff_A_AsnBQUSc1_1(.din(n5096), .dout(n5093));
    jdff dff_A_Kq8CvxTw7_1(.din(G101gat), .dout(n5096));
    jdff dff_A_tmgnPL9s8_1(.din(n5102), .dout(n5099));
    jdff dff_A_WZEDCsWq4_1(.din(n937), .dout(n5102));
    jdff dff_A_bYVKdZ3g4_2(.din(n5108), .dout(n5105));
    jdff dff_A_vg7FDJnQ3_2(.din(n937), .dout(n5108));
    jdff dff_A_QRFb94mw6_2(.din(n207), .dout(n5111));
    jdff dff_A_udxixTEL4_1(.din(G51gat), .dout(n5114));
    jdff dff_A_qjh96vI27_0(.din(n5120), .dout(n5117));
    jdff dff_A_fzqXj6HD0_0(.din(G80gat), .dout(n5120));
    jdff dff_A_gsqSXBtL6_2(.din(G80gat), .dout(n5123));
    jdff dff_A_inIXd7Eh8_0(.din(n5129), .dout(n5126));
    jdff dff_A_ChJmihjf4_0(.din(n89), .dout(n5129));
    jdff dff_A_eFGwfiAL1_0(.din(n5135), .dout(n5132));
    jdff dff_A_WzQeFSph6_0(.din(n5138), .dout(n5135));
    jdff dff_A_6lqp49I31_0(.din(G29gat), .dout(n5138));
    jdff dff_A_d0pgtZvo9_0(.din(n5144), .dout(n5141));
    jdff dff_A_6a7MvcJ44_0(.din(n5147), .dout(n5144));
    jdff dff_A_47CLtQ8n0_0(.din(n5150), .dout(n5147));
    jdff dff_A_pLKY32TV0_0(.din(G17gat), .dout(n5150));
    jdff dff_A_9QSAiuJY3_1(.din(n5156), .dout(n5153));
    jdff dff_A_hAcwclaT7_1(.din(n5159), .dout(n5156));
    jdff dff_A_tABhtonR0_1(.din(G17gat), .dout(n5159));
    jdff dff_B_bGky21ci8_2(.din(n310), .dout(n5163));
    jdff dff_B_ZRqV7zKa0_2(.din(n5163), .dout(n5166));
    jdff dff_B_hXi4GvvB5_2(.din(n5166), .dout(n5169));
    jdff dff_B_kzHPPf338_2(.din(n5169), .dout(n5172));
    jdff dff_A_ur5K87AI0_0(.din(n5177), .dout(n5174));
    jdff dff_A_oFPbvM8S9_0(.din(n5180), .dout(n5177));
    jdff dff_A_6s5JWaOQ9_0(.din(n5183), .dout(n5180));
    jdff dff_A_FQ3gAwJT5_0(.din(n5186), .dout(n5183));
    jdff dff_A_1lCmjEwm4_0(.din(n5189), .dout(n5186));
    jdff dff_A_KpHEoisX1_0(.din(n5192), .dout(n5189));
    jdff dff_A_2PZPIQRa0_0(.din(n5195), .dout(n5192));
    jdff dff_A_H81VmuLa9_0(.din(n5198), .dout(n5195));
    jdff dff_A_JCmb31hf1_0(.din(G237gat), .dout(n5198));
    jdff dff_A_4fkzmxwA3_2(.din(n5204), .dout(n5201));
    jdff dff_A_0cSXR2PC0_2(.din(n5207), .dout(n5204));
    jdff dff_A_UmHC5iqM7_2(.din(n5210), .dout(n5207));
    jdff dff_A_epP6TRl44_2(.din(n5213), .dout(n5210));
    jdff dff_A_yZveYZra3_2(.din(n5216), .dout(n5213));
    jdff dff_A_KkiWDRZQ4_2(.din(n5219), .dout(n5216));
    jdff dff_A_xjav24r93_2(.din(n5222), .dout(n5219));
    jdff dff_A_xjJ1q6HZ2_2(.din(n5225), .dout(n5222));
    jdff dff_A_5Xt0KupC1_2(.din(G237gat), .dout(n5225));
    jdff dff_A_BANckRck8_0(.din(n5231), .dout(n5228));
    jdff dff_A_kXUfKTBt6_0(.din(n5234), .dout(n5231));
    jdff dff_A_hZhmGr6N0_0(.din(n5237), .dout(n5234));
    jdff dff_A_yKn7Acjc5_0(.din(n5240), .dout(n5237));
    jdff dff_A_QnxKz3Rl1_0(.din(n5243), .dout(n5240));
    jdff dff_A_nABzgguu0_0(.din(n440), .dout(n5243));
    jdff dff_B_neQ6GObu2_0(.din(n432), .dout(n5247));
    jdff dff_A_qGEjEI2b9_1(.din(n5252), .dout(n5249));
    jdff dff_A_bQ1HpIsw9_1(.din(n5255), .dout(n5252));
    jdff dff_A_QqoOc1Jz9_1(.din(n223), .dout(n5255));
    jdff dff_A_1bJBU0Ea0_1(.din(n5261), .dout(n5258));
    jdff dff_A_CJN7BoNr6_1(.din(n5264), .dout(n5261));
    jdff dff_A_fOOkhVnI6_1(.din(n5267), .dout(n5264));
    jdff dff_A_dADlnIYC6_1(.din(G68gat), .dout(n5267));
    jdff dff_A_fVb50uyJ6_1(.din(G42gat), .dout(n5270));
    jdff dff_A_FaerhiMT4_2(.din(G42gat), .dout(n5273));
    jdff dff_A_T7TLZoUt2_1(.din(n5279), .dout(n5276));
    jdff dff_A_qO7i5XFD5_1(.din(n5282), .dout(n5279));
    jdff dff_A_y1OnYwrt7_1(.din(n5285), .dout(n5282));
    jdff dff_A_Xok89pFc6_1(.din(n5288), .dout(n5285));
    jdff dff_A_Lst0McxJ1_1(.din(G1gat), .dout(n5288));
    jdff dff_A_QxIfccYM2_1(.din(G13gat), .dout(n5291));
    jdff dff_A_egK1zrPp8_0(.din(n5307), .dout(n5294));
    jdff dff_A_rW7uXXy70_1(.din(n5300), .dout(n5297));
    jdff dff_A_5WA9MwRB4_1(.din(n5307), .dout(n5300));
    jdff dff_B_244tRTRv6_3(.din(G55gat), .dout(n5304));
    jdff dff_B_lEMQTvZA9_3(.din(n5304), .dout(n5307));
    jdff dff_A_OrDC34Ke6_1(.din(n5312), .dout(n5309));
    jdff dff_A_sh3SKIBB9_1(.din(n5315), .dout(n5312));
    jdff dff_A_K3NLT9Ak4_1(.din(n5318), .dout(n5315));
    jdff dff_A_k3sAJFMy3_1(.din(n5321), .dout(n5318));
    jdff dff_A_V3aHJn8o0_1(.din(n5324), .dout(n5321));
    jdff dff_A_2f98JMSZ7_1(.din(n5327), .dout(n5324));
    jdff dff_A_foFC6nAh4_1(.din(n5330), .dout(n5327));
    jdff dff_A_6PmdFaOp5_1(.din(n5333), .dout(n5330));
    jdff dff_A_aWmdXhqw4_1(.din(G171gat), .dout(n5333));
    jdff dff_A_vx1IlplW0_2(.din(n5339), .dout(n5336));
    jdff dff_A_UCXNWv1U7_2(.din(n5342), .dout(n5339));
    jdff dff_A_0qBQ3hYR1_2(.din(n5345), .dout(n5342));
    jdff dff_A_2crjAIGA0_2(.din(n5348), .dout(n5345));
    jdff dff_A_IqrXtOF58_2(.din(n5351), .dout(n5348));
    jdff dff_A_IMua5r6F0_2(.din(n5354), .dout(n5351));
    jdff dff_A_M6cJgRvz3_2(.din(n5357), .dout(n5354));
    jdff dff_A_bnf6zr3H2_2(.din(n5360), .dout(n5357));
    jdff dff_A_cyJN6K3q5_2(.din(n5363), .dout(n5360));
    jdff dff_A_MchCa0XT1_2(.din(n5366), .dout(n5363));
    jdff dff_A_YEa8x4XB1_2(.din(G171gat), .dout(n5366));
    jdff dff_A_wF8Cl85X4_2(.din(n93), .dout(n5369));
    jdff dff_A_ClLJEkci1_0(.din(n5369), .dout(n5372));
    jdff dff_A_f6kzESnr4_0(.din(n5372), .dout(n5375));
    jdff dff_A_tKHLe5Cw2_0(.din(n5375), .dout(n5378));
    jdff dff_A_JWwv185I6_0(.din(n5378), .dout(n5381));
    jdff dff_A_FC34CPBS3_0(.din(n5381), .dout(n5384));
    jdff dff_A_QqRuJ6Mz7_0(.din(n5384), .dout(n5387));
    jdff dff_A_hPp50bWJ9_0(.din(n5387), .dout(n5390));
    jdff dff_A_ClnPAPNM7_0(.din(n5390), .dout(n5393));
    jdff dff_A_mFisWiIl3_0(.din(n5393), .dout(n5396));
    jdff dff_A_LQZ9fwxO8_0(.din(n5396), .dout(n5399));
    jdff dff_A_sZJoyY4C3_0(.din(n5399), .dout(n5402));
    jdff dff_A_IK1gHZ8x6_0(.din(n5402), .dout(n5405));
    jdff dff_A_joFkzNBo9_0(.din(n5405), .dout(n5408));
    jdff dff_A_EME01GPk3_0(.din(n5408), .dout(n5411));
    jdff dff_A_2KG3pNHw2_0(.din(n5411), .dout(n5414));
    jdff dff_A_evZ0erhW1_0(.din(n5414), .dout(n5417));
    jdff dff_A_6lm5GJZU3_0(.din(n5417), .dout(n5420));
    jdff dff_A_4RpFJ8NO5_0(.din(n5420), .dout(n5423));
    jdff dff_A_Db8WX77x7_0(.din(n5423), .dout(n5426));
    jdff dff_A_oUv0FQ8Q0_0(.din(n5426), .dout(n5429));
    jdff dff_A_1vk4U44o1_0(.din(n5429), .dout(n5432));
    jdff dff_A_TlymtKvy7_0(.din(n5432), .dout(n5435));
    jdff dff_A_bZ5MyR6O9_0(.din(n5435), .dout(n5438));
    jdff dff_A_6rixA4pP6_0(.din(n5438), .dout(n5441));
    jdff dff_A_HsDIHK2K7_0(.din(n5441), .dout(G388gat));
    jdff dff_A_URn4EI0h7_2(.din(n101), .dout(n5447));
    jdff dff_A_XU4X6X4G4_0(.din(n5447), .dout(n5450));
    jdff dff_A_eN3cOpU68_0(.din(n5450), .dout(n5453));
    jdff dff_A_Phqa3cVI6_0(.din(n5453), .dout(n5456));
    jdff dff_A_WMxX7sO32_0(.din(n5456), .dout(n5459));
    jdff dff_A_VsfHtiiX0_0(.din(n5459), .dout(n5462));
    jdff dff_A_YygaCAQN5_0(.din(n5462), .dout(n5465));
    jdff dff_A_6gY5i48W2_0(.din(n5465), .dout(n5468));
    jdff dff_A_Gfwt14mj8_0(.din(n5468), .dout(n5471));
    jdff dff_A_k34j0FCu9_0(.din(n5471), .dout(n5474));
    jdff dff_A_v20MPbiG9_0(.din(n5474), .dout(n5477));
    jdff dff_A_gjGv3n1a4_0(.din(n5477), .dout(n5480));
    jdff dff_A_g5vGD8Aq1_0(.din(n5480), .dout(n5483));
    jdff dff_A_4ZouqCnj2_0(.din(n5483), .dout(n5486));
    jdff dff_A_1DA1D5Mc6_0(.din(n5486), .dout(n5489));
    jdff dff_A_drPR7nGB2_0(.din(n5489), .dout(n5492));
    jdff dff_A_UKTifiP88_0(.din(n5492), .dout(n5495));
    jdff dff_A_gycEUIEt7_0(.din(n5495), .dout(n5498));
    jdff dff_A_qbSLaw9U7_0(.din(n5498), .dout(n5501));
    jdff dff_A_sRsqK2Np6_0(.din(n5501), .dout(n5504));
    jdff dff_A_2h9Grpbb5_0(.din(n5504), .dout(n5507));
    jdff dff_A_kjPyLyTg1_0(.din(n5507), .dout(n5510));
    jdff dff_A_hqqkMEyB7_0(.din(n5510), .dout(n5513));
    jdff dff_A_j95b8i4I1_0(.din(n5513), .dout(n5516));
    jdff dff_A_MpPJ47RF0_0(.din(n5516), .dout(n5519));
    jdff dff_A_CkOdEVXw9_0(.din(n5519), .dout(G389gat));
    jdff dff_A_DCUnLUjN5_2(.din(n105), .dout(n5525));
    jdff dff_A_LK3B1J3Q0_0(.din(n5525), .dout(n5528));
    jdff dff_A_4UCHGtCy9_0(.din(n5528), .dout(n5531));
    jdff dff_A_L5lWpIQT0_0(.din(n5531), .dout(n5534));
    jdff dff_A_YpNPzlTs9_0(.din(n5534), .dout(n5537));
    jdff dff_A_vvj60zCk8_0(.din(n5537), .dout(n5540));
    jdff dff_A_J9zBqNvc1_0(.din(n5540), .dout(n5543));
    jdff dff_A_VuZSqEM76_0(.din(n5543), .dout(n5546));
    jdff dff_A_ySaquppi4_0(.din(n5546), .dout(n5549));
    jdff dff_A_QOoTBZhk3_0(.din(n5549), .dout(n5552));
    jdff dff_A_4pUseqsY3_0(.din(n5552), .dout(n5555));
    jdff dff_A_vuKy39YH7_0(.din(n5555), .dout(n5558));
    jdff dff_A_O6bLVEVt0_0(.din(n5558), .dout(n5561));
    jdff dff_A_ORTJY1pH6_0(.din(n5561), .dout(n5564));
    jdff dff_A_lQDhlEbv0_0(.din(n5564), .dout(n5567));
    jdff dff_A_Pyv83LjJ3_0(.din(n5567), .dout(n5570));
    jdff dff_A_sQ48iNgC9_0(.din(n5570), .dout(n5573));
    jdff dff_A_6XZ86Acu6_0(.din(n5573), .dout(n5576));
    jdff dff_A_35EwFhGE1_0(.din(n5576), .dout(n5579));
    jdff dff_A_6Yz27eOL3_0(.din(n5579), .dout(n5582));
    jdff dff_A_T5XnaazA0_0(.din(n5582), .dout(n5585));
    jdff dff_A_EPCzY0nk0_0(.din(n5585), .dout(n5588));
    jdff dff_A_ySH44Wtm2_0(.din(n5588), .dout(n5591));
    jdff dff_A_HVtHdww27_0(.din(n5591), .dout(n5594));
    jdff dff_A_XoQZlwbF4_0(.din(n5594), .dout(n5597));
    jdff dff_A_f97qhAPz3_0(.din(n5597), .dout(G390gat));
    jdff dff_A_8pBCiBMs8_2(.din(n109), .dout(n5603));
    jdff dff_A_clRKRtNn5_0(.din(n5603), .dout(n5606));
    jdff dff_A_F1xYbvEk6_0(.din(n5606), .dout(n5609));
    jdff dff_A_mwbhn23q5_0(.din(n5609), .dout(n5612));
    jdff dff_A_F4CG209h0_0(.din(n5612), .dout(n5615));
    jdff dff_A_6SrCwavk3_0(.din(n5615), .dout(n5618));
    jdff dff_A_erjEthf31_0(.din(n5618), .dout(n5621));
    jdff dff_A_a68gOB9j7_0(.din(n5621), .dout(n5624));
    jdff dff_A_WB4HwnZq6_0(.din(n5624), .dout(n5627));
    jdff dff_A_Zxswmoi59_0(.din(n5627), .dout(n5630));
    jdff dff_A_rHv7T4Nd0_0(.din(n5630), .dout(n5633));
    jdff dff_A_2ZAVattz3_0(.din(n5633), .dout(n5636));
    jdff dff_A_p3eZOdir1_0(.din(n5636), .dout(n5639));
    jdff dff_A_o6NAy5RB9_0(.din(n5639), .dout(n5642));
    jdff dff_A_hBWVZAPV9_0(.din(n5642), .dout(n5645));
    jdff dff_A_K71kYyS69_0(.din(n5645), .dout(n5648));
    jdff dff_A_ssp9WvJv0_0(.din(n5648), .dout(n5651));
    jdff dff_A_ZwAROs2J7_0(.din(n5651), .dout(n5654));
    jdff dff_A_Ebv1GTbQ8_0(.din(n5654), .dout(n5657));
    jdff dff_A_S0BYbNXc0_0(.din(n5657), .dout(n5660));
    jdff dff_A_tgchaNDi7_0(.din(n5660), .dout(n5663));
    jdff dff_A_1V4BEQ3z7_0(.din(n5663), .dout(n5666));
    jdff dff_A_8u12CGUO6_0(.din(n5666), .dout(n5669));
    jdff dff_A_KD0GetWJ0_0(.din(n5669), .dout(n5672));
    jdff dff_A_LhUQn7548_0(.din(n5672), .dout(n5675));
    jdff dff_A_04EcVYd20_0(.din(n5675), .dout(n5678));
    jdff dff_A_te6HLR6I3_0(.din(n5678), .dout(G391gat));
    jdff dff_A_h8jo52As9_2(.din(n121), .dout(n5684));
    jdff dff_A_R75aPu7G3_0(.din(n5684), .dout(n5687));
    jdff dff_A_EwHYCa2j3_0(.din(n5687), .dout(n5690));
    jdff dff_A_3hOOZs231_0(.din(n5690), .dout(n5693));
    jdff dff_A_UNaLyMaH6_0(.din(n5693), .dout(n5696));
    jdff dff_A_tNThjERl2_0(.din(n5696), .dout(n5699));
    jdff dff_A_uHLHGbMT5_0(.din(n5699), .dout(n5702));
    jdff dff_A_HTYfIR785_0(.din(n5702), .dout(n5705));
    jdff dff_A_M9YJ3cWh0_0(.din(n5705), .dout(n5708));
    jdff dff_A_8SPFwIRK5_0(.din(n5708), .dout(n5711));
    jdff dff_A_XoWZiUEt3_0(.din(n5711), .dout(n5714));
    jdff dff_A_2uGbiMSz7_0(.din(n5714), .dout(n5717));
    jdff dff_A_XJMQcD9b0_0(.din(n5717), .dout(n5720));
    jdff dff_A_tCtRc8VJ8_0(.din(n5720), .dout(n5723));
    jdff dff_A_UNHayenH9_0(.din(n5723), .dout(n5726));
    jdff dff_A_YRDJ7zfO1_0(.din(n5726), .dout(n5729));
    jdff dff_A_RE4s87sI8_0(.din(n5729), .dout(n5732));
    jdff dff_A_H1e0lKX53_0(.din(n5732), .dout(n5735));
    jdff dff_A_9sVH2EWT8_0(.din(n5735), .dout(n5738));
    jdff dff_A_UJ29qjt87_0(.din(n5738), .dout(n5741));
    jdff dff_A_j6E1AQjs1_0(.din(n5741), .dout(n5744));
    jdff dff_A_ywOoEXd11_0(.din(n5744), .dout(n5747));
    jdff dff_A_rEkvsX6m7_0(.din(n5747), .dout(n5750));
    jdff dff_A_xTDZk3NR1_0(.din(n5750), .dout(n5753));
    jdff dff_A_gyR8xsKb6_0(.din(n5753), .dout(G418gat));
    jdff dff_A_laVyLnLT1_2(.din(n149), .dout(n5759));
    jdff dff_A_DIISTH446_0(.din(n5759), .dout(n5762));
    jdff dff_A_z5pexYFN7_0(.din(n5762), .dout(n5765));
    jdff dff_A_C7NokHXA2_0(.din(n5765), .dout(n5768));
    jdff dff_A_cDGkuiuT6_0(.din(n5768), .dout(n5771));
    jdff dff_A_lopyjr0n8_0(.din(n5771), .dout(n5774));
    jdff dff_A_dHbgcKoN5_0(.din(n5774), .dout(n5777));
    jdff dff_A_YrhhiGQw7_0(.din(n5777), .dout(n5780));
    jdff dff_A_RtdbOFHE2_0(.din(n5780), .dout(n5783));
    jdff dff_A_C6d8BV7I8_0(.din(n5783), .dout(n5786));
    jdff dff_A_qopnCWSg8_0(.din(n5786), .dout(n5789));
    jdff dff_A_C3l1wK7Q2_0(.din(n5789), .dout(n5792));
    jdff dff_A_NPaJ6teP8_0(.din(n5792), .dout(n5795));
    jdff dff_A_lMVnUSQa9_0(.din(n5795), .dout(n5798));
    jdff dff_A_VwATLboz1_0(.din(n5798), .dout(n5801));
    jdff dff_A_Ov7GXoYI1_0(.din(n5801), .dout(n5804));
    jdff dff_A_w1fPEtm99_0(.din(n5804), .dout(n5807));
    jdff dff_A_mMXNLHmQ0_0(.din(n5807), .dout(n5810));
    jdff dff_A_WHGfAUfB5_0(.din(n5810), .dout(n5813));
    jdff dff_A_bePrq1Ae9_0(.din(n5813), .dout(n5816));
    jdff dff_A_gJZmO8AF9_0(.din(n5816), .dout(n5819));
    jdff dff_A_fFKp0A8X8_0(.din(n5819), .dout(n5822));
    jdff dff_A_nBLlvPvN3_0(.din(n5822), .dout(G419gat));
    jdff dff_A_deOSyrnr7_2(.din(n163), .dout(n5828));
    jdff dff_A_a4fwSDdu0_0(.din(n5828), .dout(n5831));
    jdff dff_A_Bjl15bpH7_0(.din(n5831), .dout(n5834));
    jdff dff_A_b8SdHcNp8_0(.din(n5834), .dout(n5837));
    jdff dff_A_Ovob1aRK7_0(.din(n5837), .dout(n5840));
    jdff dff_A_SQXgrj802_0(.din(n5840), .dout(n5843));
    jdff dff_A_gfpiyVsr9_0(.din(n5843), .dout(n5846));
    jdff dff_A_q9RiCr198_0(.din(n5846), .dout(n5849));
    jdff dff_A_6cGXUVLp6_0(.din(n5849), .dout(n5852));
    jdff dff_A_NBR5S5FV9_0(.din(n5852), .dout(n5855));
    jdff dff_A_tgussN988_0(.din(n5855), .dout(n5858));
    jdff dff_A_kLK4FU254_0(.din(n5858), .dout(n5861));
    jdff dff_A_S0tChvUW8_0(.din(n5861), .dout(n5864));
    jdff dff_A_vNXHHIjf9_0(.din(n5864), .dout(n5867));
    jdff dff_A_H937d63b3_0(.din(n5867), .dout(n5870));
    jdff dff_A_EUn111oZ0_0(.din(n5870), .dout(n5873));
    jdff dff_A_ioefZaX57_0(.din(n5873), .dout(n5876));
    jdff dff_A_9H0l3MS87_0(.din(n5876), .dout(n5879));
    jdff dff_A_xBDueBwD2_0(.din(n5879), .dout(n5882));
    jdff dff_A_CuuDcqMy7_0(.din(n5882), .dout(n5885));
    jdff dff_A_b0mAXX6M5_0(.din(n5885), .dout(n5888));
    jdff dff_A_akTJ28XZ2_0(.din(n5888), .dout(n5891));
    jdff dff_A_fVpoRMzG0_0(.din(n5891), .dout(n5894));
    jdff dff_A_QEwcGjuL7_0(.din(n5894), .dout(n5897));
    jdff dff_A_K9G3agmX4_0(.din(n5897), .dout(G420gat));
    jdff dff_A_lrqAObpH1_2(.din(n177), .dout(n5903));
    jdff dff_A_GcKxzyGJ6_0(.din(n5903), .dout(n5906));
    jdff dff_A_GmhPtNCE3_0(.din(n5906), .dout(n5909));
    jdff dff_A_nwps0OYt5_0(.din(n5909), .dout(n5912));
    jdff dff_A_PiJuzgoU7_0(.din(n5912), .dout(n5915));
    jdff dff_A_nLm44Rnf1_0(.din(n5915), .dout(n5918));
    jdff dff_A_IZBxedDW6_0(.din(n5918), .dout(n5921));
    jdff dff_A_yXKPRIBm4_0(.din(n5921), .dout(n5924));
    jdff dff_A_UanwxyNM5_0(.din(n5924), .dout(n5927));
    jdff dff_A_hnWstzmq3_0(.din(n5927), .dout(n5930));
    jdff dff_A_rEqdIL1A6_0(.din(n5930), .dout(n5933));
    jdff dff_A_aDdIWWAw5_0(.din(n5933), .dout(n5936));
    jdff dff_A_nC26oicF6_0(.din(n5936), .dout(n5939));
    jdff dff_A_6uET4wis0_0(.din(n5939), .dout(n5942));
    jdff dff_A_AEDBBR8K6_0(.din(n5942), .dout(n5945));
    jdff dff_A_5eQrw2qB3_0(.din(n5945), .dout(n5948));
    jdff dff_A_i8KaPZQ84_0(.din(n5948), .dout(n5951));
    jdff dff_A_9BbMzB5n3_0(.din(n5951), .dout(n5954));
    jdff dff_A_nTfYHYpn1_0(.din(n5954), .dout(n5957));
    jdff dff_A_glGd2eIY0_0(.din(n5957), .dout(n5960));
    jdff dff_A_kFXj5wby9_0(.din(n5960), .dout(n5963));
    jdff dff_A_FR4YFsJa2_0(.din(n5963), .dout(n5966));
    jdff dff_A_bZpnLv9f9_0(.din(n5966), .dout(n5969));
    jdff dff_A_o90m62D30_0(.din(n5969), .dout(n5972));
    jdff dff_A_vUia2Ft49_0(.din(n5972), .dout(G421gat));
    jdff dff_A_wFW2ch691_2(.din(n184), .dout(n5978));
    jdff dff_A_nUq230zl4_0(.din(n5978), .dout(n5981));
    jdff dff_A_qSwWXXuX5_0(.din(n5981), .dout(n5984));
    jdff dff_A_JYnFWZ4p0_0(.din(n5984), .dout(n5987));
    jdff dff_A_6Tbd5IY18_0(.din(n5987), .dout(n5990));
    jdff dff_A_dFpr3Elq1_0(.din(n5990), .dout(n5993));
    jdff dff_A_RyCOhIiE7_0(.din(n5993), .dout(n5996));
    jdff dff_A_oimxdRd20_0(.din(n5996), .dout(n5999));
    jdff dff_A_eBcUOe005_0(.din(n5999), .dout(n6002));
    jdff dff_A_x3WlSW253_0(.din(n6002), .dout(n6005));
    jdff dff_A_heONL2uT7_0(.din(n6005), .dout(n6008));
    jdff dff_A_EV4S88b56_0(.din(n6008), .dout(n6011));
    jdff dff_A_rgZALcik5_0(.din(n6011), .dout(n6014));
    jdff dff_A_4eWjyWWv5_0(.din(n6014), .dout(n6017));
    jdff dff_A_VNptx7qK4_0(.din(n6017), .dout(n6020));
    jdff dff_A_iUn7dDuR6_0(.din(n6020), .dout(n6023));
    jdff dff_A_Ut4nLxxv1_0(.din(n6023), .dout(n6026));
    jdff dff_A_BJQ5DKvF3_0(.din(n6026), .dout(n6029));
    jdff dff_A_lTPtvgTj5_0(.din(n6029), .dout(n6032));
    jdff dff_A_l0yD8ZRM2_0(.din(n6032), .dout(n6035));
    jdff dff_A_y02V02D96_0(.din(n6035), .dout(n6038));
    jdff dff_A_ycCJAbyC0_0(.din(n6038), .dout(n6041));
    jdff dff_A_8ejQo4jA0_0(.din(n6041), .dout(n6044));
    jdff dff_A_ljXSKrKm8_0(.din(n6044), .dout(n6047));
    jdff dff_A_yAVcfKPP6_0(.din(n6047), .dout(G422gat));
    jdff dff_A_EI1AbcoC2_2(.din(n192), .dout(n6053));
    jdff dff_A_8JD0Pdk98_0(.din(n6053), .dout(n6056));
    jdff dff_A_osCCU1Yc0_0(.din(n6056), .dout(n6059));
    jdff dff_A_QiF03HjA7_0(.din(n6059), .dout(n6062));
    jdff dff_A_Cl8U4e6d0_0(.din(n6062), .dout(n6065));
    jdff dff_A_X0ZFpbfj8_0(.din(n6065), .dout(n6068));
    jdff dff_A_QCHUAAkh1_0(.din(n6068), .dout(n6071));
    jdff dff_A_tNR47FzG2_0(.din(n6071), .dout(n6074));
    jdff dff_A_SEEB3kFx5_0(.din(n6074), .dout(n6077));
    jdff dff_A_Wj5wxuFc3_0(.din(n6077), .dout(n6080));
    jdff dff_A_7dVf7Ssj6_0(.din(n6080), .dout(n6083));
    jdff dff_A_wy33EccP1_0(.din(n6083), .dout(n6086));
    jdff dff_A_vShCL3cO4_0(.din(n6086), .dout(n6089));
    jdff dff_A_oj45jCHk3_0(.din(n6089), .dout(n6092));
    jdff dff_A_GM5B2vaZ3_0(.din(n6092), .dout(n6095));
    jdff dff_A_eonXjgxS2_0(.din(n6095), .dout(n6098));
    jdff dff_A_MxmfaX7b7_0(.din(n6098), .dout(n6101));
    jdff dff_A_PGsUldvm8_0(.din(n6101), .dout(n6104));
    jdff dff_A_iXOBFjoF4_0(.din(n6104), .dout(n6107));
    jdff dff_A_Et2Sl7yz8_0(.din(n6107), .dout(n6110));
    jdff dff_A_gXPrIarz7_0(.din(n6110), .dout(n6113));
    jdff dff_A_yJanGnWa1_0(.din(n6113), .dout(n6116));
    jdff dff_A_JU2DrTmE6_0(.din(n6116), .dout(n6119));
    jdff dff_A_niZrNab53_0(.din(n6119), .dout(n6122));
    jdff dff_A_yjBKcbmZ0_0(.din(n6122), .dout(n6125));
    jdff dff_A_V3bxT7gL2_0(.din(n6125), .dout(G423gat));
    jdff dff_A_O6jn1Gue3_2(.din(n199), .dout(n6131));
    jdff dff_A_kgsD6hKS3_0(.din(n6131), .dout(n6134));
    jdff dff_A_5IvpyKGc3_0(.din(n6134), .dout(n6137));
    jdff dff_A_fu73RqIQ8_0(.din(n6137), .dout(n6140));
    jdff dff_A_X9OVA8s22_0(.din(n6140), .dout(n6143));
    jdff dff_A_EZqJvrRG6_0(.din(n6143), .dout(n6146));
    jdff dff_A_Rps1wixn1_0(.din(n6146), .dout(n6149));
    jdff dff_A_r5whXDcm0_0(.din(n6149), .dout(n6152));
    jdff dff_A_oGwqlfyY7_0(.din(n6152), .dout(n6155));
    jdff dff_A_f0kZlnSr0_0(.din(n6155), .dout(n6158));
    jdff dff_A_lUJL6bqw8_0(.din(n6158), .dout(n6161));
    jdff dff_A_lW3LOW715_0(.din(n6161), .dout(n6164));
    jdff dff_A_cIiEsxtk6_0(.din(n6164), .dout(n6167));
    jdff dff_A_5uFhLSaM2_0(.din(n6167), .dout(n6170));
    jdff dff_A_uqrlZ0w69_0(.din(n6170), .dout(n6173));
    jdff dff_A_aUBDG2uL6_0(.din(n6173), .dout(n6176));
    jdff dff_A_ovWTiWeL1_0(.din(n6176), .dout(n6179));
    jdff dff_A_uDPFbiSV5_0(.din(n6179), .dout(n6182));
    jdff dff_A_PFnYDDsh9_0(.din(n6182), .dout(n6185));
    jdff dff_A_LyxSbZFw9_0(.din(n6185), .dout(n6188));
    jdff dff_A_6auhD7d33_0(.din(n6188), .dout(n6191));
    jdff dff_A_gK4yLJSg5_0(.din(n6191), .dout(n6194));
    jdff dff_A_NFlCp7eI0_0(.din(n6194), .dout(G446gat));
    jdff dff_A_bDsVM3Cz7_1(.din(n207), .dout(n6200));
    jdff dff_A_BEa6ECR94_0(.din(n6200), .dout(n6203));
    jdff dff_A_j8BSzuoO5_0(.din(n6203), .dout(n6206));
    jdff dff_A_wqewGXlq4_0(.din(n6206), .dout(n6209));
    jdff dff_A_Xrjtlo7x2_0(.din(n6209), .dout(n6212));
    jdff dff_A_JygVPBNZ0_0(.din(n6212), .dout(n6215));
    jdff dff_A_4gQ4kPKd2_0(.din(n6215), .dout(n6218));
    jdff dff_A_UjBAK97Z1_0(.din(n6218), .dout(n6221));
    jdff dff_A_v6i9W8d93_0(.din(n6221), .dout(n6224));
    jdff dff_A_dReMKxeq8_0(.din(n6224), .dout(n6227));
    jdff dff_A_hBzNvfgR7_0(.din(n6227), .dout(n6230));
    jdff dff_A_9IfKUUth2_0(.din(n6230), .dout(n6233));
    jdff dff_A_ecr7qeEJ3_0(.din(n6233), .dout(n6236));
    jdff dff_A_vfAaOUuf3_0(.din(n6236), .dout(n6239));
    jdff dff_A_r5YP6lXY8_0(.din(n6239), .dout(n6242));
    jdff dff_A_83NxtOxK1_0(.din(n6242), .dout(n6245));
    jdff dff_A_ee9mZmBx6_0(.din(n6245), .dout(n6248));
    jdff dff_A_QXu8jWsX3_0(.din(n6248), .dout(n6251));
    jdff dff_A_AKZURNN02_0(.din(n6251), .dout(n6254));
    jdff dff_A_WvwA8LiT6_0(.din(n6254), .dout(n6257));
    jdff dff_A_Krl3ZUX24_0(.din(n6257), .dout(n6260));
    jdff dff_A_bPIcYI5T0_0(.din(n6260), .dout(n6263));
    jdff dff_A_6iYzJI2M5_0(.din(n6263), .dout(n6266));
    jdff dff_A_YCHX3iBi0_0(.din(n6266), .dout(n6269));
    jdff dff_A_Ptv9l8jB6_0(.din(n6269), .dout(n6272));
    jdff dff_A_JveD93U55_0(.din(n6272), .dout(G447gat));
    jdff dff_A_d7DwcygA1_2(.din(n219), .dout(n6278));
endmodule

