module gf_c6288(G511gat, G154gat, G222gat, G256gat, G375gat, G137gat, G52gat, G35gat, G171gat, G69gat, G18gat, G86gat, G409gat, G443gat, G188gat, G1gat, G120gat, G494gat, G477gat, G205gat, G307gat, G239gat, G273gat, G290gat, G358gat, G324gat, G528gat, G341gat, G392gat, G426gat, G103gat, G460gat, G6287gat, G6280gat, G5308gat, G4591gat, G2877gat, G4946gat, G3895gat, G3552gat, G6250gat, G3211gat, G2548gat, G6270gat, G1901gat, G6170gat, G1581gat, G4241gat, G545gat, G5672gat, G6160gat, G5971gat, G6123gat, G6200gat, G6288gat, G6150gat, G2223gat, G6260gat, G6180gat, G6190gat, G6220gat, G6230gat, G6210gat, G6240gat);
    input G511gat, G154gat, G222gat, G256gat, G375gat, G137gat, G52gat, G35gat, G171gat, G69gat, G18gat, G86gat, G409gat, G443gat, G188gat, G1gat, G120gat, G494gat, G477gat, G205gat, G307gat, G239gat, G273gat, G290gat, G358gat, G324gat, G528gat, G341gat, G392gat, G426gat, G103gat, G460gat;
    output G6287gat, G6280gat, G5308gat, G4591gat, G2877gat, G4946gat, G3895gat, G3552gat, G6250gat, G3211gat, G2548gat, G6270gat, G1901gat, G6170gat, G1581gat, G4241gat, G545gat, G5672gat, G6160gat, G5971gat, G6123gat, G6200gat, G6288gat, G6150gat, G2223gat, G6260gat, G6180gat, G6190gat, G6220gat, G6230gat, G6210gat, G6240gat;
    wire n67;
    wire n71;
    wire n75;
    wire n78;
    wire n81;
    wire n84;
    wire n88;
    wire n91;
    wire n95;
    wire n99;
    wire n103;
    wire n107;
    wire n110;
    wire n113;
    wire n116;
    wire n120;
    wire n124;
    wire n128;
    wire n132;
    wire n136;
    wire n140;
    wire n144;
    wire n148;
    wire n151;
    wire n155;
    wire n159;
    wire n163;
    wire n167;
    wire n170;
    wire n173;
    wire n177;
    wire n180;
    wire n184;
    wire n188;
    wire n192;
    wire n196;
    wire n200;
    wire n204;
    wire n208;
    wire n212;
    wire n216;
    wire n220;
    wire n224;
    wire n227;
    wire n230;
    wire n234;
    wire n238;
    wire n242;
    wire n246;
    wire n249;
    wire n253;
    wire n257;
    wire n261;
    wire n265;
    wire n269;
    wire n272;
    wire n275;
    wire n279;
    wire n283;
    wire n286;
    wire n290;
    wire n294;
    wire n298;
    wire n302;
    wire n306;
    wire n310;
    wire n313;
    wire n317;
    wire n321;
    wire n325;
    wire n329;
    wire n333;
    wire n336;
    wire n339;
    wire n343;
    wire n347;
    wire n351;
    wire n355;
    wire n358;
    wire n362;
    wire n366;
    wire n370;
    wire n374;
    wire n378;
    wire n381;
    wire n385;
    wire n388;
    wire n392;
    wire n396;
    wire n400;
    wire n403;
    wire n407;
    wire n411;
    wire n414;
    wire n418;
    wire n422;
    wire n426;
    wire n430;
    wire n434;
    wire n438;
    wire n442;
    wire n445;
    wire n449;
    wire n453;
    wire n457;
    wire n461;
    wire n465;
    wire n468;
    wire n471;
    wire n475;
    wire n479;
    wire n483;
    wire n487;
    wire n490;
    wire n494;
    wire n498;
    wire n502;
    wire n506;
    wire n510;
    wire n513;
    wire n517;
    wire n521;
    wire n525;
    wire n529;
    wire n532;
    wire n535;
    wire n539;
    wire n543;
    wire n547;
    wire n551;
    wire n554;
    wire n558;
    wire n562;
    wire n565;
    wire n569;
    wire n573;
    wire n577;
    wire n581;
    wire n585;
    wire n589;
    wire n593;
    wire n597;
    wire n601;
    wire n604;
    wire n608;
    wire n612;
    wire n616;
    wire n620;
    wire n624;
    wire n627;
    wire n630;
    wire n634;
    wire n638;
    wire n642;
    wire n646;
    wire n649;
    wire n653;
    wire n657;
    wire n661;
    wire n665;
    wire n669;
    wire n672;
    wire n676;
    wire n680;
    wire n684;
    wire n688;
    wire n691;
    wire n695;
    wire n699;
    wire n703;
    wire n707;
    wire n710;
    wire n713;
    wire n717;
    wire n721;
    wire n725;
    wire n729;
    wire n732;
    wire n736;
    wire n740;
    wire n743;
    wire n747;
    wire n751;
    wire n755;
    wire n759;
    wire n763;
    wire n767;
    wire n771;
    wire n775;
    wire n779;
    wire n783;
    wire n787;
    wire n790;
    wire n794;
    wire n798;
    wire n802;
    wire n806;
    wire n810;
    wire n813;
    wire n816;
    wire n820;
    wire n824;
    wire n828;
    wire n832;
    wire n835;
    wire n839;
    wire n843;
    wire n847;
    wire n851;
    wire n855;
    wire n858;
    wire n862;
    wire n866;
    wire n870;
    wire n874;
    wire n877;
    wire n881;
    wire n885;
    wire n889;
    wire n893;
    wire n896;
    wire n900;
    wire n904;
    wire n908;
    wire n912;
    wire n915;
    wire n919;
    wire n922;
    wire n926;
    wire n930;
    wire n934;
    wire n937;
    wire n941;
    wire n945;
    wire n948;
    wire n952;
    wire n956;
    wire n960;
    wire n964;
    wire n968;
    wire n972;
    wire n976;
    wire n980;
    wire n984;
    wire n988;
    wire n992;
    wire n996;
    wire n1000;
    wire n1003;
    wire n1007;
    wire n1011;
    wire n1015;
    wire n1019;
    wire n1023;
    wire n1026;
    wire n1029;
    wire n1033;
    wire n1037;
    wire n1041;
    wire n1045;
    wire n1048;
    wire n1052;
    wire n1056;
    wire n1060;
    wire n1064;
    wire n1068;
    wire n1071;
    wire n1075;
    wire n1079;
    wire n1083;
    wire n1087;
    wire n1090;
    wire n1094;
    wire n1098;
    wire n1102;
    wire n1106;
    wire n1109;
    wire n1113;
    wire n1117;
    wire n1121;
    wire n1125;
    wire n1128;
    wire n1132;
    wire n1136;
    wire n1140;
    wire n1144;
    wire n1147;
    wire n1151;
    wire n1154;
    wire n1158;
    wire n1162;
    wire n1166;
    wire n1169;
    wire n1173;
    wire n1177;
    wire n1180;
    wire n1184;
    wire n1188;
    wire n1192;
    wire n1196;
    wire n1200;
    wire n1204;
    wire n1208;
    wire n1212;
    wire n1216;
    wire n1220;
    wire n1224;
    wire n1228;
    wire n1232;
    wire n1236;
    wire n1240;
    wire n1243;
    wire n1247;
    wire n1251;
    wire n1255;
    wire n1259;
    wire n1263;
    wire n1266;
    wire n1269;
    wire n1273;
    wire n1277;
    wire n1281;
    wire n1285;
    wire n1288;
    wire n1292;
    wire n1296;
    wire n1300;
    wire n1304;
    wire n1308;
    wire n1311;
    wire n1315;
    wire n1319;
    wire n1323;
    wire n1327;
    wire n1330;
    wire n1334;
    wire n1338;
    wire n1342;
    wire n1346;
    wire n1349;
    wire n1353;
    wire n1357;
    wire n1361;
    wire n1365;
    wire n1368;
    wire n1372;
    wire n1376;
    wire n1380;
    wire n1384;
    wire n1387;
    wire n1391;
    wire n1395;
    wire n1399;
    wire n1403;
    wire n1406;
    wire n1410;
    wire n1414;
    wire n1417;
    wire n1421;
    wire n1424;
    wire n1428;
    wire n1431;
    wire n1435;
    wire n1439;
    wire n1442;
    wire n1446;
    wire n1450;
    wire n1454;
    wire n1458;
    wire n1462;
    wire n1466;
    wire n1470;
    wire n1474;
    wire n1478;
    wire n1482;
    wire n1486;
    wire n1490;
    wire n1494;
    wire n1498;
    wire n1502;
    wire n1506;
    wire n1510;
    wire n1513;
    wire n1517;
    wire n1521;
    wire n1525;
    wire n1529;
    wire n1533;
    wire n1536;
    wire n1539;
    wire n1543;
    wire n1547;
    wire n1551;
    wire n1555;
    wire n1558;
    wire n1562;
    wire n1566;
    wire n1570;
    wire n1574;
    wire n1578;
    wire n1581;
    wire n1585;
    wire n1589;
    wire n1593;
    wire n1597;
    wire n1600;
    wire n1604;
    wire n1608;
    wire n1612;
    wire n1616;
    wire n1619;
    wire n1623;
    wire n1627;
    wire n1631;
    wire n1635;
    wire n1638;
    wire n1642;
    wire n1646;
    wire n1650;
    wire n1654;
    wire n1657;
    wire n1661;
    wire n1665;
    wire n1669;
    wire n1673;
    wire n1676;
    wire n1680;
    wire n1684;
    wire n1688;
    wire n1692;
    wire n1695;
    wire n1699;
    wire n1703;
    wire n1706;
    wire n1710;
    wire n1713;
    wire n1717;
    wire n1720;
    wire n1724;
    wire n1728;
    wire n1731;
    wire n1735;
    wire n1739;
    wire n1743;
    wire n1747;
    wire n1751;
    wire n1755;
    wire n1759;
    wire n1763;
    wire n1767;
    wire n1771;
    wire n1775;
    wire n1779;
    wire n1783;
    wire n1787;
    wire n1791;
    wire n1795;
    wire n1799;
    wire n1803;
    wire n1807;
    wire n1810;
    wire n1814;
    wire n1818;
    wire n1822;
    wire n1826;
    wire n1830;
    wire n1833;
    wire n1836;
    wire n1840;
    wire n1844;
    wire n1848;
    wire n1852;
    wire n1855;
    wire n1859;
    wire n1863;
    wire n1867;
    wire n1871;
    wire n1875;
    wire n1878;
    wire n1882;
    wire n1886;
    wire n1890;
    wire n1894;
    wire n1897;
    wire n1901;
    wire n1905;
    wire n1909;
    wire n1913;
    wire n1916;
    wire n1920;
    wire n1924;
    wire n1928;
    wire n1932;
    wire n1935;
    wire n1939;
    wire n1943;
    wire n1947;
    wire n1951;
    wire n1954;
    wire n1958;
    wire n1962;
    wire n1966;
    wire n1970;
    wire n1973;
    wire n1977;
    wire n1981;
    wire n1985;
    wire n1989;
    wire n1992;
    wire n1996;
    wire n2000;
    wire n2004;
    wire n2008;
    wire n2011;
    wire n2015;
    wire n2019;
    wire n2022;
    wire n2026;
    wire n2029;
    wire n2033;
    wire n2036;
    wire n2040;
    wire n2044;
    wire n2047;
    wire n2051;
    wire n2055;
    wire n2059;
    wire n2063;
    wire n2067;
    wire n2071;
    wire n2075;
    wire n2079;
    wire n2083;
    wire n2087;
    wire n2091;
    wire n2095;
    wire n2099;
    wire n2103;
    wire n2107;
    wire n2111;
    wire n2115;
    wire n2119;
    wire n2123;
    wire n2127;
    wire n2131;
    wire n2134;
    wire n2138;
    wire n2142;
    wire n2146;
    wire n2150;
    wire n2154;
    wire n2157;
    wire n2160;
    wire n2164;
    wire n2168;
    wire n2172;
    wire n2176;
    wire n2179;
    wire n2183;
    wire n2187;
    wire n2191;
    wire n2195;
    wire n2199;
    wire n2202;
    wire n2206;
    wire n2210;
    wire n2214;
    wire n2218;
    wire n2221;
    wire n2225;
    wire n2229;
    wire n2233;
    wire n2237;
    wire n2240;
    wire n2244;
    wire n2248;
    wire n2252;
    wire n2256;
    wire n2259;
    wire n2263;
    wire n2267;
    wire n2271;
    wire n2275;
    wire n2278;
    wire n2282;
    wire n2286;
    wire n2290;
    wire n2294;
    wire n2297;
    wire n2301;
    wire n2305;
    wire n2309;
    wire n2313;
    wire n2316;
    wire n2320;
    wire n2324;
    wire n2328;
    wire n2332;
    wire n2335;
    wire n2339;
    wire n2343;
    wire n2347;
    wire n2351;
    wire n2354;
    wire n2358;
    wire n2362;
    wire n2365;
    wire n2369;
    wire n2372;
    wire n2376;
    wire n2379;
    wire n2383;
    wire n2387;
    wire n2390;
    wire n2394;
    wire n2398;
    wire n2402;
    wire n2406;
    wire n2410;
    wire n2414;
    wire n2418;
    wire n2422;
    wire n2426;
    wire n2430;
    wire n2434;
    wire n2438;
    wire n2442;
    wire n2446;
    wire n2450;
    wire n2454;
    wire n2458;
    wire n2462;
    wire n2466;
    wire n2470;
    wire n2474;
    wire n2478;
    wire n2482;
    wire n2485;
    wire n2489;
    wire n2493;
    wire n2497;
    wire n2501;
    wire n2505;
    wire n2508;
    wire n2511;
    wire n2515;
    wire n2519;
    wire n2523;
    wire n2527;
    wire n2530;
    wire n2534;
    wire n2538;
    wire n2542;
    wire n2546;
    wire n2550;
    wire n2553;
    wire n2557;
    wire n2561;
    wire n2565;
    wire n2569;
    wire n2572;
    wire n2576;
    wire n2580;
    wire n2584;
    wire n2588;
    wire n2591;
    wire n2595;
    wire n2599;
    wire n2603;
    wire n2607;
    wire n2610;
    wire n2614;
    wire n2618;
    wire n2622;
    wire n2626;
    wire n2629;
    wire n2633;
    wire n2637;
    wire n2641;
    wire n2645;
    wire n2648;
    wire n2652;
    wire n2656;
    wire n2660;
    wire n2664;
    wire n2667;
    wire n2671;
    wire n2675;
    wire n2679;
    wire n2683;
    wire n2686;
    wire n2690;
    wire n2694;
    wire n2698;
    wire n2702;
    wire n2705;
    wire n2709;
    wire n2713;
    wire n2717;
    wire n2721;
    wire n2724;
    wire n2728;
    wire n2732;
    wire n2735;
    wire n2739;
    wire n2742;
    wire n2746;
    wire n2749;
    wire n2753;
    wire n2757;
    wire n2760;
    wire n2764;
    wire n2768;
    wire n2772;
    wire n2776;
    wire n2780;
    wire n2784;
    wire n2788;
    wire n2792;
    wire n2796;
    wire n2800;
    wire n2804;
    wire n2808;
    wire n2812;
    wire n2816;
    wire n2820;
    wire n2824;
    wire n2828;
    wire n2832;
    wire n2836;
    wire n2840;
    wire n2844;
    wire n2848;
    wire n2852;
    wire n2856;
    wire n2860;
    wire n2863;
    wire n2867;
    wire n2871;
    wire n2875;
    wire n2879;
    wire n2883;
    wire n2886;
    wire n2889;
    wire n2893;
    wire n2897;
    wire n2901;
    wire n2905;
    wire n2909;
    wire n2913;
    wire n2917;
    wire n2921;
    wire n2925;
    wire n2928;
    wire n2932;
    wire n2936;
    wire n2940;
    wire n2944;
    wire n2947;
    wire n2951;
    wire n2955;
    wire n2959;
    wire n2963;
    wire n2966;
    wire n2970;
    wire n2974;
    wire n2978;
    wire n2982;
    wire n2985;
    wire n2989;
    wire n2993;
    wire n2997;
    wire n3001;
    wire n3004;
    wire n3008;
    wire n3012;
    wire n3016;
    wire n3020;
    wire n3023;
    wire n3027;
    wire n3031;
    wire n3035;
    wire n3039;
    wire n3042;
    wire n3046;
    wire n3050;
    wire n3054;
    wire n3058;
    wire n3061;
    wire n3065;
    wire n3069;
    wire n3073;
    wire n3077;
    wire n3080;
    wire n3084;
    wire n3088;
    wire n3092;
    wire n3096;
    wire n3099;
    wire n3103;
    wire n3107;
    wire n3111;
    wire n3115;
    wire n3118;
    wire n3122;
    wire n3126;
    wire n3129;
    wire n3133;
    wire n3136;
    wire n3140;
    wire n3143;
    wire n3147;
    wire n3151;
    wire n3155;
    wire n3159;
    wire n3163;
    wire n3167;
    wire n3171;
    wire n3175;
    wire n3179;
    wire n3183;
    wire n3187;
    wire n3191;
    wire n3195;
    wire n3199;
    wire n3203;
    wire n3207;
    wire n3211;
    wire n3215;
    wire n3219;
    wire n3223;
    wire n3227;
    wire n3231;
    wire n3235;
    wire n3239;
    wire n3243;
    wire n3247;
    wire n3251;
    wire n3255;
    wire n3259;
    wire n3263;
    wire n3267;
    wire n3271;
    wire n3274;
    wire n3278;
    wire n3282;
    wire n3286;
    wire n3290;
    wire n3293;
    wire n3297;
    wire n3301;
    wire n3305;
    wire n3309;
    wire n3313;
    wire n3316;
    wire n3319;
    wire n3323;
    wire n3327;
    wire n3331;
    wire n3335;
    wire n3338;
    wire n3342;
    wire n3346;
    wire n3350;
    wire n3354;
    wire n3357;
    wire n3361;
    wire n3365;
    wire n3369;
    wire n3373;
    wire n3376;
    wire n3380;
    wire n3384;
    wire n3388;
    wire n3392;
    wire n3395;
    wire n3399;
    wire n3403;
    wire n3407;
    wire n3411;
    wire n3414;
    wire n3418;
    wire n3422;
    wire n3426;
    wire n3430;
    wire n3433;
    wire n3437;
    wire n3441;
    wire n3445;
    wire n3449;
    wire n3452;
    wire n3456;
    wire n3460;
    wire n3464;
    wire n3468;
    wire n3471;
    wire n3475;
    wire n3479;
    wire n3483;
    wire n3487;
    wire n3490;
    wire n3494;
    wire n3498;
    wire n3502;
    wire n3506;
    wire n3509;
    wire n3513;
    wire n3517;
    wire n3521;
    wire n3525;
    wire n3528;
    wire n3532;
    wire n3535;
    wire n3539;
    wire n3542;
    wire n3545;
    wire n3549;
    wire n3553;
    wire n3556;
    wire n3560;
    wire n3564;
    wire n3568;
    wire n3572;
    wire n3576;
    wire n3580;
    wire n3584;
    wire n3588;
    wire n3592;
    wire n3596;
    wire n3600;
    wire n3604;
    wire n3608;
    wire n3612;
    wire n3616;
    wire n3620;
    wire n3624;
    wire n3628;
    wire n3632;
    wire n3636;
    wire n3640;
    wire n3644;
    wire n3648;
    wire n3652;
    wire n3656;
    wire n3660;
    wire n3663;
    wire n3667;
    wire n3671;
    wire n3675;
    wire n3679;
    wire n3683;
    wire n3687;
    wire n3691;
    wire n3695;
    wire n3699;
    wire n3702;
    wire n3706;
    wire n3710;
    wire n3714;
    wire n3718;
    wire n3722;
    wire n3726;
    wire n3730;
    wire n3734;
    wire n3737;
    wire n3741;
    wire n3745;
    wire n3749;
    wire n3753;
    wire n3756;
    wire n3760;
    wire n3764;
    wire n3768;
    wire n3772;
    wire n3775;
    wire n3779;
    wire n3783;
    wire n3787;
    wire n3791;
    wire n3794;
    wire n3798;
    wire n3802;
    wire n3806;
    wire n3810;
    wire n3813;
    wire n3817;
    wire n3821;
    wire n3825;
    wire n3829;
    wire n3832;
    wire n3836;
    wire n3840;
    wire n3844;
    wire n3848;
    wire n3851;
    wire n3855;
    wire n3859;
    wire n3863;
    wire n3867;
    wire n3870;
    wire n3874;
    wire n3878;
    wire n3882;
    wire n3886;
    wire n3889;
    wire n3893;
    wire n3897;
    wire n3901;
    wire n3905;
    wire n3908;
    wire n3912;
    wire n3916;
    wire n3920;
    wire n3924;
    wire n3928;
    wire n3932;
    wire n3936;
    wire n3940;
    wire n3943;
    wire n3947;
    wire n3951;
    wire n3955;
    wire n3959;
    wire n3963;
    wire n3967;
    wire n3971;
    wire n3975;
    wire n3979;
    wire n3983;
    wire n3987;
    wire n3991;
    wire n3995;
    wire n3999;
    wire n4003;
    wire n4007;
    wire n4011;
    wire n4015;
    wire n4019;
    wire n4023;
    wire n4027;
    wire n4031;
    wire n4034;
    wire n4038;
    wire n4042;
    wire n4046;
    wire n4050;
    wire n4053;
    wire n4057;
    wire n4060;
    wire n4064;
    wire n4068;
    wire n4072;
    wire n4075;
    wire n4079;
    wire n4083;
    wire n4087;
    wire n4091;
    wire n4095;
    wire n4098;
    wire n4102;
    wire n4106;
    wire n4110;
    wire n4113;
    wire n4117;
    wire n4121;
    wire n4125;
    wire n4129;
    wire n4132;
    wire n4136;
    wire n4140;
    wire n4144;
    wire n4148;
    wire n4151;
    wire n4155;
    wire n4159;
    wire n4163;
    wire n4167;
    wire n4170;
    wire n4174;
    wire n4178;
    wire n4182;
    wire n4186;
    wire n4189;
    wire n4193;
    wire n4197;
    wire n4201;
    wire n4205;
    wire n4208;
    wire n4212;
    wire n4216;
    wire n4220;
    wire n4224;
    wire n4227;
    wire n4231;
    wire n4235;
    wire n4239;
    wire n4243;
    wire n4246;
    wire n4250;
    wire n4254;
    wire n4258;
    wire n4262;
    wire n4265;
    wire n4269;
    wire n4273;
    wire n4277;
    wire n4281;
    wire n4284;
    wire n4288;
    wire n4292;
    wire n4296;
    wire n4300;
    wire n4304;
    wire n4308;
    wire n4312;
    wire n4316;
    wire n4320;
    wire n4323;
    wire n4327;
    wire n4331;
    wire n4335;
    wire n4339;
    wire n4343;
    wire n4347;
    wire n4351;
    wire n4355;
    wire n4359;
    wire n4363;
    wire n4367;
    wire n4371;
    wire n4375;
    wire n4379;
    wire n4383;
    wire n4387;
    wire n4391;
    wire n4395;
    wire n4399;
    wire n4403;
    wire n4407;
    wire n4410;
    wire n4414;
    wire n4417;
    wire n4421;
    wire n4425;
    wire n4428;
    wire n4432;
    wire n4435;
    wire n4439;
    wire n4443;
    wire n4447;
    wire n4451;
    wire n4455;
    wire n4459;
    wire n4463;
    wire n4467;
    wire n4471;
    wire n4475;
    wire n4479;
    wire n4482;
    wire n4486;
    wire n4490;
    wire n4494;
    wire n4498;
    wire n4501;
    wire n4505;
    wire n4509;
    wire n4513;
    wire n4517;
    wire n4520;
    wire n4524;
    wire n4528;
    wire n4532;
    wire n4536;
    wire n4539;
    wire n4543;
    wire n4547;
    wire n4551;
    wire n4555;
    wire n4558;
    wire n4562;
    wire n4566;
    wire n4570;
    wire n4574;
    wire n4577;
    wire n4581;
    wire n4585;
    wire n4589;
    wire n4593;
    wire n4596;
    wire n4600;
    wire n4604;
    wire n4608;
    wire n4612;
    wire n4615;
    wire n4619;
    wire n4623;
    wire n4627;
    wire n4631;
    wire n4634;
    wire n4638;
    wire n4642;
    wire n4646;
    wire n4650;
    wire n4654;
    wire n4658;
    wire n4662;
    wire n4666;
    wire n4670;
    wire n4673;
    wire n4677;
    wire n4681;
    wire n4685;
    wire n4689;
    wire n4693;
    wire n4697;
    wire n4701;
    wire n4705;
    wire n4709;
    wire n4713;
    wire n4717;
    wire n4721;
    wire n4725;
    wire n4729;
    wire n4733;
    wire n4737;
    wire n4741;
    wire n4745;
    wire n4749;
    wire n4753;
    wire n4756;
    wire n4760;
    wire n4764;
    wire n4767;
    wire n4771;
    wire n4774;
    wire n4778;
    wire n4782;
    wire n4786;
    wire n4789;
    wire n4792;
    wire n4796;
    wire n4800;
    wire n4804;
    wire n4808;
    wire n4812;
    wire n4816;
    wire n4820;
    wire n4824;
    wire n4827;
    wire n4831;
    wire n4835;
    wire n4839;
    wire n4843;
    wire n4846;
    wire n4850;
    wire n4854;
    wire n4858;
    wire n4862;
    wire n4865;
    wire n4869;
    wire n4873;
    wire n4877;
    wire n4881;
    wire n4884;
    wire n4888;
    wire n4892;
    wire n4896;
    wire n4900;
    wire n4903;
    wire n4907;
    wire n4911;
    wire n4915;
    wire n4919;
    wire n4922;
    wire n4926;
    wire n4930;
    wire n4934;
    wire n4938;
    wire n4941;
    wire n4945;
    wire n4949;
    wire n4953;
    wire n4957;
    wire n4960;
    wire n4964;
    wire n4968;
    wire n4972;
    wire n4976;
    wire n4980;
    wire n4984;
    wire n4988;
    wire n4992;
    wire n4996;
    wire n4999;
    wire n5003;
    wire n5007;
    wire n5011;
    wire n5015;
    wire n5019;
    wire n5023;
    wire n5027;
    wire n5031;
    wire n5035;
    wire n5039;
    wire n5043;
    wire n5047;
    wire n5051;
    wire n5055;
    wire n5059;
    wire n5063;
    wire n5067;
    wire n5071;
    wire n5074;
    wire n5078;
    wire n5081;
    wire n5085;
    wire n5089;
    wire n5093;
    wire n5096;
    wire n5100;
    wire n5104;
    wire n5107;
    wire n5110;
    wire n5114;
    wire n5118;
    wire n5122;
    wire n5126;
    wire n5130;
    wire n5134;
    wire n5138;
    wire n5142;
    wire n5145;
    wire n5149;
    wire n5153;
    wire n5157;
    wire n5161;
    wire n5164;
    wire n5168;
    wire n5172;
    wire n5176;
    wire n5180;
    wire n5183;
    wire n5187;
    wire n5191;
    wire n5195;
    wire n5199;
    wire n5202;
    wire n5206;
    wire n5210;
    wire n5214;
    wire n5218;
    wire n5221;
    wire n5225;
    wire n5229;
    wire n5233;
    wire n5237;
    wire n5240;
    wire n5244;
    wire n5248;
    wire n5252;
    wire n5256;
    wire n5259;
    wire n5263;
    wire n5267;
    wire n5271;
    wire n5275;
    wire n5279;
    wire n5283;
    wire n5287;
    wire n5291;
    wire n5295;
    wire n5298;
    wire n5302;
    wire n5306;
    wire n5310;
    wire n5314;
    wire n5318;
    wire n5322;
    wire n5326;
    wire n5330;
    wire n5334;
    wire n5338;
    wire n5342;
    wire n5346;
    wire n5350;
    wire n5354;
    wire n5358;
    wire n5362;
    wire n5365;
    wire n5369;
    wire n5372;
    wire n5376;
    wire n5380;
    wire n5384;
    wire n5387;
    wire n5391;
    wire n5395;
    wire n5398;
    wire n5401;
    wire n5405;
    wire n5409;
    wire n5413;
    wire n5417;
    wire n5421;
    wire n5425;
    wire n5429;
    wire n5433;
    wire n5436;
    wire n5440;
    wire n5444;
    wire n5448;
    wire n5452;
    wire n5455;
    wire n5459;
    wire n5463;
    wire n5467;
    wire n5471;
    wire n5474;
    wire n5478;
    wire n5482;
    wire n5486;
    wire n5490;
    wire n5493;
    wire n5497;
    wire n5501;
    wire n5505;
    wire n5509;
    wire n5512;
    wire n5516;
    wire n5520;
    wire n5524;
    wire n5528;
    wire n5531;
    wire n5535;
    wire n5539;
    wire n5543;
    wire n5547;
    wire n5551;
    wire n5555;
    wire n5559;
    wire n5563;
    wire n5567;
    wire n5570;
    wire n5574;
    wire n5578;
    wire n5582;
    wire n5586;
    wire n5590;
    wire n5594;
    wire n5598;
    wire n5602;
    wire n5606;
    wire n5610;
    wire n5614;
    wire n5618;
    wire n5622;
    wire n5626;
    wire n5629;
    wire n5633;
    wire n5636;
    wire n5640;
    wire n5644;
    wire n5648;
    wire n5651;
    wire n5655;
    wire n5659;
    wire n5662;
    wire n5665;
    wire n5669;
    wire n5673;
    wire n5677;
    wire n5681;
    wire n5685;
    wire n5689;
    wire n5693;
    wire n5697;
    wire n5700;
    wire n5704;
    wire n5708;
    wire n5712;
    wire n5716;
    wire n5719;
    wire n5723;
    wire n5727;
    wire n5731;
    wire n5735;
    wire n5738;
    wire n5742;
    wire n5746;
    wire n5750;
    wire n5754;
    wire n5757;
    wire n5761;
    wire n5765;
    wire n5769;
    wire n5773;
    wire n5776;
    wire n5780;
    wire n5784;
    wire n5788;
    wire n5792;
    wire n5796;
    wire n5800;
    wire n5804;
    wire n5808;
    wire n5812;
    wire n5815;
    wire n5819;
    wire n5823;
    wire n5827;
    wire n5831;
    wire n5835;
    wire n5839;
    wire n5843;
    wire n5847;
    wire n5851;
    wire n5855;
    wire n5859;
    wire n5863;
    wire n5866;
    wire n5870;
    wire n5873;
    wire n5877;
    wire n5881;
    wire n5885;
    wire n5888;
    wire n5892;
    wire n5896;
    wire n5899;
    wire n5902;
    wire n5906;
    wire n5910;
    wire n5914;
    wire n5918;
    wire n5922;
    wire n5926;
    wire n5930;
    wire n5934;
    wire n5937;
    wire n5941;
    wire n5945;
    wire n5949;
    wire n5953;
    wire n5956;
    wire n5960;
    wire n5964;
    wire n5968;
    wire n5972;
    wire n5975;
    wire n5979;
    wire n5983;
    wire n5987;
    wire n5991;
    wire n5994;
    wire n5998;
    wire n6002;
    wire n6006;
    wire n6010;
    wire n6014;
    wire n6018;
    wire n6022;
    wire n6026;
    wire n6030;
    wire n6033;
    wire n6037;
    wire n6041;
    wire n6045;
    wire n6049;
    wire n6053;
    wire n6057;
    wire n6061;
    wire n6065;
    wire n6069;
    wire n6073;
    wire n6076;
    wire n6080;
    wire n6083;
    wire n6087;
    wire n6091;
    wire n6095;
    wire n6098;
    wire n6102;
    wire n6106;
    wire n6109;
    wire n6112;
    wire n6116;
    wire n6120;
    wire n6124;
    wire n6128;
    wire n6131;
    wire n6135;
    wire n6139;
    wire n6143;
    wire n6147;
    wire n6150;
    wire n6154;
    wire n6158;
    wire n6162;
    wire n6166;
    wire n6169;
    wire n6173;
    wire n6177;
    wire n6181;
    wire n6185;
    wire n6188;
    wire n6192;
    wire n6196;
    wire n6200;
    wire n6204;
    wire n6208;
    wire n6212;
    wire n6216;
    wire n6220;
    wire n6224;
    wire n6227;
    wire n6231;
    wire n6235;
    wire n6239;
    wire n6243;
    wire n6247;
    wire n6251;
    wire n6255;
    wire n6259;
    wire n6263;
    wire n6266;
    wire n6270;
    wire n6274;
    wire n6278;
    wire n6281;
    wire n6285;
    wire n6289;
    wire n6293;
    wire n6297;
    wire n6301;
    wire n6305;
    wire n6308;
    wire n6312;
    wire n6316;
    wire n6320;
    wire n6324;
    wire n6327;
    wire n6331;
    wire n6335;
    wire n6339;
    wire n6343;
    wire n6346;
    wire n6350;
    wire n6354;
    wire n6358;
    wire n6362;
    wire n6366;
    wire n6370;
    wire n6374;
    wire n6378;
    wire n6382;
    wire n6385;
    wire n6389;
    wire n6393;
    wire n6397;
    wire n6401;
    wire n6405;
    wire n6409;
    wire n6413;
    wire n6417;
    wire n6421;
    wire n6424;
    wire n6427;
    wire n6431;
    wire n6434;
    wire n6438;
    wire n6442;
    wire n6446;
    wire n6450;
    wire n6454;
    wire n6458;
    wire n6461;
    wire n6465;
    wire n6469;
    wire n6473;
    wire n6477;
    wire n6480;
    wire n6484;
    wire n6488;
    wire n6492;
    wire n6496;
    wire n6500;
    wire n6504;
    wire n6508;
    wire n6512;
    wire n6516;
    wire n6519;
    wire n6523;
    wire n6527;
    wire n6531;
    wire n6535;
    wire n6539;
    wire n6543;
    wire n6547;
    wire n6550;
    wire n6553;
    wire n6557;
    wire n6560;
    wire n6564;
    wire n6568;
    wire n6572;
    wire n6576;
    wire n6580;
    wire n6584;
    wire n6587;
    wire n6591;
    wire n6595;
    wire n6599;
    wire n6603;
    wire n6607;
    wire n6611;
    wire n6615;
    wire n6619;
    wire n6623;
    wire n6626;
    wire n6630;
    wire n6634;
    wire n6638;
    wire n6642;
    wire n6646;
    wire n6649;
    wire n6652;
    wire n6656;
    wire n6659;
    wire n6663;
    wire n6667;
    wire n6671;
    wire n6675;
    wire n6679;
    wire n6683;
    wire n6687;
    wire n6691;
    wire n6695;
    wire n6699;
    wire n6703;
    wire n6706;
    wire n6710;
    wire n6714;
    wire n6718;
    wire n6722;
    wire n6726;
    wire n6730;
    wire n6734;
    wire n6738;
    wire n6741;
    wire n6744;
    wire n6748;
    wire n6751;
    wire n6755;
    wire n6759;
    wire n6763;
    wire n6766;
    wire n6770;
    wire n6778;
    wire n10593;
    wire n10596;
    wire n10599;
    wire n10602;
    wire n10605;
    wire n10608;
    wire n10611;
    wire n10614;
    wire n10617;
    wire n10620;
    wire n10623;
    wire n10626;
    wire n10629;
    wire n10632;
    wire n10635;
    wire n10638;
    wire n10641;
    wire n10644;
    wire n10647;
    wire n10650;
    wire n10653;
    wire n10656;
    wire n10659;
    wire n10662;
    wire n10665;
    wire n10668;
    wire n10671;
    wire n10674;
    wire n10677;
    wire n10680;
    wire n10683;
    wire n10686;
    wire n10689;
    wire n10692;
    wire n10695;
    wire n10698;
    wire n10701;
    wire n10704;
    wire n10707;
    wire n10710;
    wire n10713;
    wire n10716;
    wire n10719;
    wire n10722;
    wire n10725;
    wire n10728;
    wire n10731;
    wire n10734;
    wire n10737;
    wire n10740;
    wire n10743;
    wire n10746;
    wire n10749;
    wire n10752;
    wire n10755;
    wire n10758;
    wire n10761;
    wire n10764;
    wire n10767;
    wire n10770;
    wire n10773;
    wire n10776;
    wire n10779;
    wire n10782;
    wire n10785;
    wire n10788;
    wire n10791;
    wire n10794;
    wire n10797;
    wire n10800;
    wire n10803;
    wire n10806;
    wire n10809;
    wire n10812;
    wire n10815;
    wire n10818;
    wire n10821;
    wire n10824;
    wire n10827;
    wire n10830;
    wire n10833;
    wire n10836;
    wire n10839;
    wire n10842;
    wire n10845;
    wire n10848;
    wire n10851;
    wire n10854;
    wire n10857;
    wire n10860;
    wire n10863;
    wire n10866;
    wire n10869;
    wire n10872;
    wire n10875;
    wire n10878;
    wire n10881;
    wire n10884;
    wire n10887;
    wire n10890;
    wire n10893;
    wire n10896;
    wire n10899;
    wire n10902;
    wire n10905;
    wire n10908;
    wire n10911;
    wire n10914;
    wire n10917;
    wire n10920;
    wire n10923;
    wire n10926;
    wire n10929;
    wire n10932;
    wire n10935;
    wire n10938;
    wire n10941;
    wire n10944;
    wire n10947;
    wire n10950;
    wire n10953;
    wire n10956;
    wire n10959;
    wire n10962;
    wire n10965;
    wire n10968;
    wire n10971;
    wire n10974;
    wire n10977;
    wire n10980;
    wire n10983;
    wire n10986;
    wire n10989;
    wire n10992;
    wire n10995;
    wire n10998;
    wire n11001;
    wire n11004;
    wire n11007;
    wire n11010;
    wire n11013;
    wire n11016;
    wire n11019;
    wire n11022;
    wire n11025;
    wire n11028;
    wire n11031;
    wire n11034;
    wire n11037;
    wire n11040;
    wire n11043;
    wire n11046;
    wire n11049;
    wire n11052;
    wire n11055;
    wire n11058;
    wire n11061;
    wire n11064;
    wire n11067;
    wire n11070;
    wire n11073;
    wire n11076;
    wire n11079;
    wire n11082;
    wire n11085;
    wire n11088;
    wire n11091;
    wire n11094;
    wire n11097;
    wire n11100;
    wire n11103;
    wire n11106;
    wire n11109;
    wire n11112;
    wire n11115;
    wire n11118;
    wire n11121;
    wire n11124;
    wire n11127;
    wire n11130;
    wire n11133;
    wire n11136;
    wire n11139;
    wire n11142;
    wire n11145;
    wire n11148;
    wire n11151;
    wire n11154;
    wire n11157;
    wire n11160;
    wire n11163;
    wire n11166;
    wire n11169;
    wire n11172;
    wire n11175;
    wire n11178;
    wire n11181;
    wire n11184;
    wire n11187;
    wire n11190;
    wire n11193;
    wire n11196;
    wire n11199;
    wire n11202;
    wire n11205;
    wire n11208;
    wire n11211;
    wire n11214;
    wire n11217;
    wire n11220;
    wire n11223;
    wire n11226;
    wire n11229;
    wire n11232;
    wire n11235;
    wire n11238;
    wire n11241;
    wire n11244;
    wire n11247;
    wire n11250;
    wire n11253;
    wire n11256;
    wire n11259;
    wire n11262;
    wire n11265;
    wire n11268;
    wire n11271;
    wire n11274;
    wire n11277;
    wire n11280;
    wire n11283;
    wire n11286;
    wire n11289;
    wire n11292;
    wire n11295;
    wire n11298;
    wire n11301;
    wire n11304;
    wire n11307;
    wire n11310;
    wire n11313;
    wire n11316;
    wire n11319;
    wire n11322;
    wire n11325;
    wire n11328;
    wire n11331;
    wire n11334;
    wire n11337;
    wire n11340;
    wire n11343;
    wire n11346;
    wire n11349;
    wire n11352;
    wire n11355;
    wire n11358;
    wire n11361;
    wire n11364;
    wire n11367;
    wire n11370;
    wire n11373;
    wire n11376;
    wire n11379;
    wire n11382;
    wire n11385;
    wire n11388;
    wire n11391;
    wire n11394;
    wire n11397;
    wire n11400;
    wire n11403;
    wire n11406;
    wire n11409;
    wire n11412;
    wire n11415;
    wire n11418;
    wire n11421;
    wire n11424;
    wire n11427;
    wire n11430;
    wire n11433;
    wire n11436;
    wire n11439;
    wire n11442;
    wire n11445;
    wire n11448;
    wire n11451;
    wire n11454;
    wire n11457;
    wire n11460;
    wire n11463;
    wire n11466;
    wire n11469;
    wire n11472;
    wire n11475;
    wire n11478;
    wire n11481;
    wire n11484;
    wire n11487;
    wire n11490;
    wire n11493;
    wire n11496;
    wire n11499;
    wire n11502;
    wire n11505;
    wire n11508;
    wire n11511;
    wire n11514;
    wire n11517;
    wire n11520;
    wire n11523;
    wire n11526;
    wire n11529;
    wire n11532;
    wire n11535;
    wire n11538;
    wire n11541;
    wire n11544;
    wire n11547;
    wire n11550;
    wire n11553;
    wire n11556;
    wire n11559;
    wire n11562;
    wire n11565;
    wire n11568;
    wire n11571;
    wire n11574;
    wire n11577;
    wire n11580;
    wire n11583;
    wire n11586;
    wire n11589;
    wire n11592;
    wire n11595;
    wire n11598;
    wire n11601;
    wire n11604;
    wire n11607;
    wire n11610;
    wire n11613;
    wire n11616;
    wire n11619;
    wire n11622;
    wire n11625;
    wire n11628;
    wire n11630;
    wire n11633;
    wire n11636;
    wire n11639;
    wire n11642;
    wire n11645;
    wire n11648;
    wire n11651;
    wire n11654;
    wire n11657;
    wire n11660;
    wire n11663;
    wire n11666;
    wire n11669;
    wire n11673;
    wire n11676;
    wire n11679;
    wire n11682;
    wire n11685;
    wire n11688;
    wire n11691;
    wire n11694;
    wire n11697;
    wire n11700;
    wire n11703;
    wire n11706;
    wire n11709;
    wire n11712;
    wire n11715;
    wire n11718;
    wire n11721;
    wire n11724;
    wire n11727;
    wire n11730;
    wire n11733;
    wire n11736;
    wire n11739;
    wire n11742;
    wire n11745;
    wire n11748;
    wire n11751;
    wire n11754;
    wire n11757;
    wire n11760;
    wire n11763;
    wire n11766;
    wire n11769;
    wire n11772;
    wire n11775;
    wire n11778;
    wire n11781;
    wire n11784;
    wire n11787;
    wire n11790;
    wire n11793;
    wire n11796;
    wire n11799;
    wire n11802;
    wire n11805;
    wire n11808;
    wire n11811;
    wire n11814;
    wire n11817;
    wire n11820;
    wire n11823;
    wire n11826;
    wire n11829;
    wire n11832;
    wire n11835;
    wire n11838;
    wire n11841;
    wire n11844;
    wire n11847;
    wire n11850;
    wire n11853;
    wire n11856;
    wire n11859;
    wire n11862;
    wire n11865;
    wire n11868;
    wire n11871;
    wire n11874;
    wire n11877;
    wire n11880;
    wire n11883;
    wire n11886;
    wire n11889;
    wire n11892;
    wire n11895;
    wire n11898;
    wire n11901;
    wire n11904;
    wire n11907;
    wire n11910;
    wire n11913;
    wire n11916;
    wire n11919;
    wire n11922;
    wire n11924;
    wire n11927;
    wire n11930;
    wire n11933;
    wire n11936;
    wire n11939;
    wire n11942;
    wire n11945;
    wire n11948;
    wire n11951;
    wire n11954;
    wire n11957;
    wire n11960;
    wire n11964;
    wire n11967;
    wire n11970;
    wire n11973;
    wire n11976;
    wire n11979;
    wire n11982;
    wire n11985;
    wire n11988;
    wire n11991;
    wire n11994;
    wire n11997;
    wire n12000;
    wire n12003;
    wire n12006;
    wire n12009;
    wire n12012;
    wire n12015;
    wire n12018;
    wire n12021;
    wire n12024;
    wire n12027;
    wire n12030;
    wire n12033;
    wire n12036;
    wire n12038;
    wire n12041;
    wire n12044;
    wire n12047;
    wire n12050;
    wire n12053;
    wire n12056;
    wire n12059;
    wire n12062;
    wire n12065;
    wire n12068;
    wire n12071;
    wire n12074;
    wire n12078;
    wire n12081;
    wire n12084;
    wire n12087;
    wire n12090;
    wire n12093;
    wire n12096;
    wire n12099;
    wire n12102;
    wire n12105;
    wire n12108;
    wire n12111;
    wire n12114;
    wire n12117;
    wire n12120;
    wire n12123;
    wire n12126;
    wire n12129;
    wire n12132;
    wire n12135;
    wire n12138;
    wire n12141;
    wire n12144;
    wire n12147;
    wire n12150;
    wire n12152;
    wire n12155;
    wire n12158;
    wire n12161;
    wire n12164;
    wire n12167;
    wire n12170;
    wire n12173;
    wire n12176;
    wire n12179;
    wire n12182;
    wire n12185;
    wire n12188;
    wire n12192;
    wire n12195;
    wire n12198;
    wire n12201;
    wire n12204;
    wire n12207;
    wire n12210;
    wire n12213;
    wire n12216;
    wire n12219;
    wire n12222;
    wire n12225;
    wire n12228;
    wire n12231;
    wire n12234;
    wire n12237;
    wire n12240;
    wire n12243;
    wire n12246;
    wire n12249;
    wire n12252;
    wire n12255;
    wire n12258;
    wire n12261;
    wire n12264;
    wire n12266;
    wire n12269;
    wire n12272;
    wire n12275;
    wire n12278;
    wire n12281;
    wire n12284;
    wire n12287;
    wire n12290;
    wire n12293;
    wire n12296;
    wire n12299;
    wire n12302;
    wire n12306;
    wire n12309;
    wire n12312;
    wire n12315;
    wire n12318;
    wire n12321;
    wire n12324;
    wire n12327;
    wire n12330;
    wire n12333;
    wire n12336;
    wire n12339;
    wire n12342;
    wire n12345;
    wire n12348;
    wire n12351;
    wire n12354;
    wire n12357;
    wire n12360;
    wire n12363;
    wire n12366;
    wire n12369;
    wire n12372;
    wire n12375;
    wire n12377;
    wire n12380;
    wire n12383;
    wire n12386;
    wire n12389;
    wire n12392;
    wire n12395;
    wire n12398;
    wire n12401;
    wire n12404;
    wire n12407;
    wire n12410;
    wire n12414;
    wire n12417;
    wire n12420;
    wire n12423;
    wire n12426;
    wire n12429;
    wire n12432;
    wire n12435;
    wire n12438;
    wire n12441;
    wire n12444;
    wire n12447;
    wire n12450;
    wire n12453;
    wire n12456;
    wire n12459;
    wire n12462;
    wire n12465;
    wire n12468;
    wire n12471;
    wire n12474;
    wire n12477;
    wire n12479;
    wire n12482;
    wire n12485;
    wire n12488;
    wire n12491;
    wire n12494;
    wire n12497;
    wire n12500;
    wire n12503;
    wire n12506;
    wire n12509;
    wire n12513;
    wire n12516;
    wire n12519;
    wire n12522;
    wire n12525;
    wire n12528;
    wire n12531;
    wire n12534;
    wire n12537;
    wire n12540;
    wire n12543;
    wire n12546;
    wire n12549;
    wire n12552;
    wire n12555;
    wire n12558;
    wire n12561;
    wire n12564;
    wire n12566;
    wire n12569;
    wire n12572;
    wire n12575;
    wire n12578;
    wire n12581;
    wire n12584;
    wire n12587;
    wire n12590;
    wire n12594;
    wire n12597;
    wire n12600;
    wire n12603;
    wire n12606;
    wire n12609;
    wire n12612;
    wire n12615;
    wire n12618;
    wire n12621;
    wire n12624;
    wire n12627;
    wire n12630;
    wire n12633;
    wire n12635;
    wire n12638;
    wire n12641;
    wire n12644;
    wire n12647;
    wire n12650;
    wire n12653;
    wire n12657;
    wire n12660;
    wire n12663;
    wire n12666;
    wire n12669;
    wire n12672;
    wire n12675;
    wire n12678;
    wire n12681;
    wire n12684;
    wire n12687;
    wire n12690;
    wire n12692;
    wire n12695;
    wire n12698;
    wire n12701;
    wire n12704;
    wire n12707;
    wire n12711;
    wire n12714;
    wire n12717;
    wire n12720;
    wire n12723;
    wire n12726;
    wire n12729;
    wire n12732;
    wire n12735;
    wire n12738;
    wire n12740;
    wire n12743;
    wire n12746;
    wire n12749;
    wire n12752;
    wire n12756;
    wire n12759;
    wire n12762;
    wire n12764;
    wire n12767;
    wire n12771;
    wire n12773;
    wire n12777;
    wire n12779;
    wire n12783;
    wire n12786;
    wire n12788;
    wire n12791;
    wire n12794;
    wire n12797;
    wire n12800;
    wire n12803;
    wire n12806;
    wire n12809;
    wire n12812;
    wire n12815;
    wire n12818;
    wire n12821;
    wire n12824;
    wire n12827;
    wire n12830;
    wire n12833;
    wire n12836;
    wire n12839;
    wire n12842;
    wire n12845;
    wire n12848;
    wire n12851;
    wire n12854;
    wire n12857;
    wire n12860;
    wire n12863;
    wire n12866;
    wire n12869;
    wire n12872;
    wire n12875;
    wire n12878;
    wire n12881;
    wire n12884;
    wire n12887;
    wire n12890;
    wire n12893;
    wire n12896;
    wire n12899;
    wire n12902;
    wire n12905;
    wire n12908;
    wire n12911;
    wire n12914;
    wire n12917;
    wire n12921;
    wire n12923;
    wire n12926;
    wire n12929;
    wire n12932;
    wire n12935;
    wire n12938;
    wire n12941;
    wire n12944;
    wire n12947;
    wire n12950;
    wire n12953;
    wire n12956;
    wire n12959;
    wire n12962;
    wire n12965;
    wire n12968;
    wire n12971;
    wire n12974;
    wire n12977;
    wire n12980;
    wire n12983;
    wire n12986;
    wire n12989;
    wire n12992;
    wire n12995;
    wire n12998;
    wire n13001;
    wire n13004;
    wire n13007;
    wire n13010;
    wire n13013;
    wire n13016;
    wire n13019;
    wire n13022;
    wire n13025;
    wire n13028;
    wire n13031;
    wire n13034;
    wire n13037;
    wire n13040;
    wire n13043;
    wire n13047;
    wire n13050;
    wire n13053;
    wire n13056;
    wire n13059;
    wire n13062;
    wire n13065;
    wire n13068;
    wire n13071;
    wire n13074;
    wire n13077;
    wire n13080;
    wire n13083;
    wire n13086;
    wire n13089;
    wire n13092;
    wire n13095;
    wire n13098;
    wire n13101;
    wire n13104;
    wire n13107;
    wire n13110;
    wire n13113;
    wire n13116;
    wire n13119;
    wire n13122;
    wire n13125;
    wire n13128;
    wire n13131;
    wire n13134;
    wire n13137;
    wire n13140;
    wire n13143;
    wire n13146;
    wire n13149;
    wire n13152;
    wire n13155;
    wire n13157;
    wire n13160;
    wire n13163;
    wire n13166;
    wire n13169;
    wire n13172;
    wire n13175;
    wire n13178;
    wire n13181;
    wire n13184;
    wire n13187;
    wire n13190;
    wire n13193;
    wire n13196;
    wire n13199;
    wire n13202;
    wire n13205;
    wire n13208;
    wire n13211;
    wire n13214;
    wire n13217;
    wire n13220;
    wire n13223;
    wire n13226;
    wire n13229;
    wire n13232;
    wire n13235;
    wire n13238;
    wire n13241;
    wire n13244;
    wire n13247;
    wire n13250;
    wire n13253;
    wire n13256;
    wire n13259;
    wire n13262;
    wire n13265;
    wire n13268;
    wire n13272;
    wire n13275;
    wire n13278;
    wire n13281;
    wire n13284;
    wire n13287;
    wire n13290;
    wire n13293;
    wire n13296;
    wire n13299;
    wire n13302;
    wire n13305;
    wire n13308;
    wire n13311;
    wire n13314;
    wire n13317;
    wire n13320;
    wire n13323;
    wire n13326;
    wire n13329;
    wire n13332;
    wire n13335;
    wire n13338;
    wire n13341;
    wire n13344;
    wire n13347;
    wire n13350;
    wire n13353;
    wire n13356;
    wire n13359;
    wire n13362;
    wire n13365;
    wire n13368;
    wire n13371;
    wire n13373;
    wire n13376;
    wire n13379;
    wire n13382;
    wire n13385;
    wire n13388;
    wire n13391;
    wire n13394;
    wire n13397;
    wire n13400;
    wire n13403;
    wire n13406;
    wire n13409;
    wire n13412;
    wire n13415;
    wire n13418;
    wire n13421;
    wire n13424;
    wire n13427;
    wire n13430;
    wire n13433;
    wire n13436;
    wire n13439;
    wire n13442;
    wire n13445;
    wire n13448;
    wire n13451;
    wire n13454;
    wire n13457;
    wire n13460;
    wire n13463;
    wire n13466;
    wire n13469;
    wire n13472;
    wire n13475;
    wire n13479;
    wire n13482;
    wire n13485;
    wire n13488;
    wire n13491;
    wire n13494;
    wire n13497;
    wire n13500;
    wire n13503;
    wire n13506;
    wire n13509;
    wire n13512;
    wire n13515;
    wire n13518;
    wire n13521;
    wire n13524;
    wire n13527;
    wire n13530;
    wire n13533;
    wire n13536;
    wire n13539;
    wire n13542;
    wire n13545;
    wire n13548;
    wire n13551;
    wire n13554;
    wire n13557;
    wire n13560;
    wire n13563;
    wire n13566;
    wire n13569;
    wire n13571;
    wire n13574;
    wire n13577;
    wire n13580;
    wire n13583;
    wire n13586;
    wire n13589;
    wire n13592;
    wire n13595;
    wire n13598;
    wire n13601;
    wire n13604;
    wire n13607;
    wire n13610;
    wire n13613;
    wire n13616;
    wire n13619;
    wire n13622;
    wire n13625;
    wire n13628;
    wire n13631;
    wire n13634;
    wire n13637;
    wire n13640;
    wire n13643;
    wire n13646;
    wire n13649;
    wire n13652;
    wire n13655;
    wire n13658;
    wire n13661;
    wire n13664;
    wire n13668;
    wire n13671;
    wire n13674;
    wire n13677;
    wire n13680;
    wire n13683;
    wire n13686;
    wire n13689;
    wire n13692;
    wire n13695;
    wire n13698;
    wire n13701;
    wire n13704;
    wire n13707;
    wire n13710;
    wire n13713;
    wire n13716;
    wire n13719;
    wire n13722;
    wire n13725;
    wire n13728;
    wire n13731;
    wire n13734;
    wire n13737;
    wire n13740;
    wire n13743;
    wire n13746;
    wire n13749;
    wire n13751;
    wire n13754;
    wire n13757;
    wire n13760;
    wire n13763;
    wire n13766;
    wire n13769;
    wire n13772;
    wire n13775;
    wire n13778;
    wire n13781;
    wire n13784;
    wire n13787;
    wire n13790;
    wire n13793;
    wire n13796;
    wire n13799;
    wire n13802;
    wire n13805;
    wire n13808;
    wire n13811;
    wire n13814;
    wire n13817;
    wire n13820;
    wire n13823;
    wire n13826;
    wire n13829;
    wire n13832;
    wire n13835;
    wire n13839;
    wire n13842;
    wire n13845;
    wire n13848;
    wire n13851;
    wire n13854;
    wire n13857;
    wire n13860;
    wire n13863;
    wire n13866;
    wire n13869;
    wire n13872;
    wire n13875;
    wire n13878;
    wire n13881;
    wire n13884;
    wire n13887;
    wire n13890;
    wire n13893;
    wire n13896;
    wire n13899;
    wire n13902;
    wire n13905;
    wire n13908;
    wire n13911;
    wire n13913;
    wire n13916;
    wire n13919;
    wire n13922;
    wire n13925;
    wire n13928;
    wire n13931;
    wire n13934;
    wire n13937;
    wire n13940;
    wire n13943;
    wire n13946;
    wire n13949;
    wire n13952;
    wire n13955;
    wire n13958;
    wire n13961;
    wire n13964;
    wire n13967;
    wire n13970;
    wire n13973;
    wire n13976;
    wire n13979;
    wire n13982;
    wire n13985;
    wire n13988;
    wire n13992;
    wire n13995;
    wire n13998;
    wire n14001;
    wire n14004;
    wire n14007;
    wire n14010;
    wire n14013;
    wire n14016;
    wire n14019;
    wire n14022;
    wire n14025;
    wire n14028;
    wire n14031;
    wire n14034;
    wire n14037;
    wire n14040;
    wire n14043;
    wire n14046;
    wire n14049;
    wire n14052;
    wire n14055;
    wire n14057;
    wire n14060;
    wire n14063;
    wire n14066;
    wire n14069;
    wire n14072;
    wire n14075;
    wire n14078;
    wire n14081;
    wire n14084;
    wire n14087;
    wire n14090;
    wire n14093;
    wire n14096;
    wire n14099;
    wire n14102;
    wire n14105;
    wire n14108;
    wire n14111;
    wire n14114;
    wire n14117;
    wire n14120;
    wire n14123;
    wire n14127;
    wire n14130;
    wire n14133;
    wire n14136;
    wire n14139;
    wire n14142;
    wire n14145;
    wire n14148;
    wire n14151;
    wire n14154;
    wire n14157;
    wire n14160;
    wire n14163;
    wire n14166;
    wire n14169;
    wire n14172;
    wire n14175;
    wire n14178;
    wire n14181;
    wire n14183;
    wire n14186;
    wire n14189;
    wire n14192;
    wire n14195;
    wire n14198;
    wire n14201;
    wire n14204;
    wire n14207;
    wire n14210;
    wire n14213;
    wire n14216;
    wire n14219;
    wire n14222;
    wire n14225;
    wire n14228;
    wire n14231;
    wire n14234;
    wire n14237;
    wire n14240;
    wire n14244;
    wire n14247;
    wire n14250;
    wire n14253;
    wire n14256;
    wire n14259;
    wire n14262;
    wire n14265;
    wire n14268;
    wire n14271;
    wire n14274;
    wire n14277;
    wire n14280;
    wire n14283;
    wire n14286;
    wire n14289;
    wire n14291;
    wire n14294;
    wire n14297;
    wire n14300;
    wire n14303;
    wire n14306;
    wire n14309;
    wire n14312;
    wire n14315;
    wire n14318;
    wire n14321;
    wire n14324;
    wire n14327;
    wire n14330;
    wire n14333;
    wire n14336;
    wire n14339;
    wire n14343;
    wire n14346;
    wire n14349;
    wire n14352;
    wire n14355;
    wire n14358;
    wire n14361;
    wire n14364;
    wire n14367;
    wire n14370;
    wire n14373;
    wire n14376;
    wire n14379;
    wire n14381;
    wire n14384;
    wire n14387;
    wire n14390;
    wire n14393;
    wire n14396;
    wire n14399;
    wire n14402;
    wire n14405;
    wire n14408;
    wire n14411;
    wire n14414;
    wire n14417;
    wire n14420;
    wire n14424;
    wire n14427;
    wire n14430;
    wire n14433;
    wire n14436;
    wire n14439;
    wire n14442;
    wire n14445;
    wire n14448;
    wire n14451;
    wire n14453;
    wire n14456;
    wire n14459;
    wire n14462;
    wire n14465;
    wire n14468;
    wire n14471;
    wire n14474;
    wire n14477;
    wire n14480;
    wire n14483;
    wire n14487;
    wire n14490;
    wire n14493;
    wire n14496;
    wire n14499;
    wire n14502;
    wire n14505;
    wire n14507;
    wire n14510;
    wire n14513;
    wire n14516;
    wire n14519;
    wire n14522;
    wire n14525;
    wire n14528;
    wire n14532;
    wire n14535;
    wire n14538;
    wire n14541;
    wire n14544;
    wire n14546;
    wire n14549;
    wire n14552;
    wire n14555;
    wire n14559;
    wire n14561;
    wire n14564;
    wire n14567;
    wire n14571;
    wire n14574;
    wire n14577;
    wire n14580;
    wire n14583;
    wire n14586;
    wire n14589;
    wire n14592;
    wire n14595;
    wire n14598;
    wire n14601;
    wire n14604;
    wire n14607;
    wire n14610;
    wire n14613;
    wire n14616;
    wire n14619;
    wire n14622;
    wire n14625;
    wire n14628;
    wire n14631;
    wire n14634;
    wire n14637;
    wire n14640;
    wire n14643;
    wire n14646;
    wire n14649;
    wire n14652;
    wire n14655;
    wire n14658;
    wire n14661;
    wire n14664;
    wire n14667;
    wire n14670;
    wire n14673;
    wire n14676;
    wire n14679;
    wire n14682;
    wire n14685;
    wire n14688;
    wire n14691;
    wire n14694;
    wire n14697;
    wire n14700;
    wire n14702;
    wire n14706;
    wire n14709;
    wire n14712;
    wire n14715;
    wire n14718;
    wire n14721;
    wire n14724;
    wire n14727;
    wire n14730;
    wire n14733;
    wire n14736;
    wire n14739;
    wire n14742;
    wire n14745;
    wire n14748;
    wire n14751;
    wire n14754;
    wire n14757;
    wire n14760;
    wire n14763;
    wire n14766;
    wire n14769;
    wire n14772;
    wire n14775;
    wire n14778;
    wire n14781;
    wire n14784;
    wire n14787;
    wire n14790;
    wire n14793;
    wire n14796;
    wire n14799;
    wire n14802;
    wire n14805;
    wire n14808;
    wire n14811;
    wire n14814;
    wire n14817;
    wire n14820;
    wire n14823;
    wire n14826;
    wire n14828;
    wire n14832;
    wire n14835;
    wire n14838;
    wire n14841;
    wire n14844;
    wire n14847;
    wire n14850;
    wire n14853;
    wire n14856;
    wire n14859;
    wire n14862;
    wire n14865;
    wire n14868;
    wire n14871;
    wire n14874;
    wire n14877;
    wire n14880;
    wire n14883;
    wire n14886;
    wire n14889;
    wire n14892;
    wire n14895;
    wire n14898;
    wire n14901;
    wire n14904;
    wire n14907;
    wire n14910;
    wire n14913;
    wire n14916;
    wire n14919;
    wire n14922;
    wire n14925;
    wire n14928;
    wire n14931;
    wire n14934;
    wire n14937;
    wire n14940;
    wire n14942;
    wire n14945;
    wire n14948;
    wire n14951;
    wire n14954;
    wire n14957;
    wire n14960;
    wire n14963;
    wire n14966;
    wire n14969;
    wire n14972;
    wire n14975;
    wire n14978;
    wire n14981;
    wire n14984;
    wire n14987;
    wire n14990;
    wire n14993;
    wire n14996;
    wire n14999;
    wire n15002;
    wire n15005;
    wire n15008;
    wire n15011;
    wire n15014;
    wire n15017;
    wire n15020;
    wire n15023;
    wire n15026;
    wire n15029;
    wire n15032;
    wire n15035;
    wire n15038;
    wire n15041;
    wire n15044;
    wire n15047;
    wire n15050;
    wire n15053;
    wire n15057;
    wire n15059;
    wire n15062;
    wire n15065;
    wire n15068;
    wire n15071;
    wire n15074;
    wire n15077;
    wire n15080;
    wire n15083;
    wire n15086;
    wire n15089;
    wire n15092;
    wire n15095;
    wire n15098;
    wire n15101;
    wire n15104;
    wire n15107;
    wire n15110;
    wire n15113;
    wire n15116;
    wire n15119;
    wire n15122;
    wire n15125;
    wire n15128;
    wire n15131;
    wire n15134;
    wire n15137;
    wire n15140;
    wire n15143;
    wire n15146;
    wire n15149;
    wire n15152;
    wire n15155;
    wire n15158;
    wire n15161;
    wire n15165;
    wire n15167;
    wire n15170;
    wire n15173;
    wire n15176;
    wire n15179;
    wire n15182;
    wire n15185;
    wire n15188;
    wire n15191;
    wire n15194;
    wire n15197;
    wire n15200;
    wire n15203;
    wire n15206;
    wire n15209;
    wire n15212;
    wire n15215;
    wire n15218;
    wire n15221;
    wire n15224;
    wire n15227;
    wire n15230;
    wire n15233;
    wire n15236;
    wire n15239;
    wire n15242;
    wire n15245;
    wire n15248;
    wire n15251;
    wire n15254;
    wire n15257;
    wire n15260;
    wire n15264;
    wire n15266;
    wire n15269;
    wire n15272;
    wire n15275;
    wire n15278;
    wire n15281;
    wire n15284;
    wire n15287;
    wire n15290;
    wire n15293;
    wire n15296;
    wire n15299;
    wire n15302;
    wire n15305;
    wire n15308;
    wire n15311;
    wire n15314;
    wire n15317;
    wire n15320;
    wire n15323;
    wire n15326;
    wire n15329;
    wire n15332;
    wire n15335;
    wire n15338;
    wire n15341;
    wire n15344;
    wire n15347;
    wire n15350;
    wire n15354;
    wire n15356;
    wire n15359;
    wire n15362;
    wire n15365;
    wire n15368;
    wire n15371;
    wire n15374;
    wire n15377;
    wire n15380;
    wire n15383;
    wire n15386;
    wire n15389;
    wire n15392;
    wire n15395;
    wire n15398;
    wire n15401;
    wire n15404;
    wire n15407;
    wire n15410;
    wire n15413;
    wire n15416;
    wire n15419;
    wire n15422;
    wire n15425;
    wire n15428;
    wire n15431;
    wire n15435;
    wire n15437;
    wire n15440;
    wire n15443;
    wire n15446;
    wire n15449;
    wire n15452;
    wire n15455;
    wire n15458;
    wire n15461;
    wire n15464;
    wire n15467;
    wire n15470;
    wire n15473;
    wire n15476;
    wire n15479;
    wire n15482;
    wire n15485;
    wire n15488;
    wire n15491;
    wire n15494;
    wire n15497;
    wire n15500;
    wire n15503;
    wire n15507;
    wire n15509;
    wire n15512;
    wire n15515;
    wire n15518;
    wire n15521;
    wire n15524;
    wire n15527;
    wire n15530;
    wire n15533;
    wire n15536;
    wire n15539;
    wire n15542;
    wire n15545;
    wire n15548;
    wire n15551;
    wire n15554;
    wire n15557;
    wire n15560;
    wire n15563;
    wire n15566;
    wire n15570;
    wire n15572;
    wire n15575;
    wire n15578;
    wire n15581;
    wire n15584;
    wire n15587;
    wire n15590;
    wire n15593;
    wire n15596;
    wire n15599;
    wire n15602;
    wire n15605;
    wire n15608;
    wire n15611;
    wire n15614;
    wire n15617;
    wire n15620;
    wire n15624;
    wire n15626;
    wire n15629;
    wire n15632;
    wire n15635;
    wire n15638;
    wire n15641;
    wire n15644;
    wire n15647;
    wire n15650;
    wire n15653;
    wire n15656;
    wire n15659;
    wire n15662;
    wire n15665;
    wire n15669;
    wire n15671;
    wire n15674;
    wire n15677;
    wire n15680;
    wire n15683;
    wire n15686;
    wire n15689;
    wire n15692;
    wire n15695;
    wire n15698;
    wire n15701;
    wire n15705;
    wire n15707;
    wire n15710;
    wire n15713;
    wire n15716;
    wire n15719;
    wire n15722;
    wire n15725;
    wire n15728;
    wire n15732;
    wire n15734;
    wire n15737;
    wire n15740;
    wire n15743;
    wire n15747;
    wire n15749;
    wire n15752;
    wire n15756;
    wire n15759;
    wire n15762;
    wire n15765;
    wire n15768;
    wire n15771;
    wire n15774;
    wire n15777;
    wire n15780;
    wire n15783;
    wire n15786;
    wire n15789;
    wire n15792;
    wire n15795;
    wire n15798;
    wire n15801;
    wire n15804;
    wire n15807;
    wire n15810;
    wire n15813;
    wire n15816;
    wire n15819;
    wire n15822;
    wire n15825;
    wire n15828;
    wire n15831;
    wire n15834;
    wire n15837;
    wire n15840;
    wire n15843;
    wire n15846;
    wire n15849;
    wire n15852;
    wire n15855;
    wire n15858;
    wire n15861;
    wire n15864;
    wire n15867;
    wire n15870;
    wire n15873;
    wire n15876;
    wire n15879;
    wire n15882;
    wire n15885;
    wire n15887;
    wire n15891;
    wire n15894;
    wire n15897;
    wire n15900;
    wire n15903;
    wire n15906;
    wire n15909;
    wire n15912;
    wire n15915;
    wire n15918;
    wire n15921;
    wire n15924;
    wire n15927;
    wire n15930;
    wire n15933;
    wire n15936;
    wire n15939;
    wire n15942;
    wire n15945;
    wire n15948;
    wire n15951;
    wire n15954;
    wire n15957;
    wire n15960;
    wire n15963;
    wire n15966;
    wire n15969;
    wire n15972;
    wire n15975;
    wire n15978;
    wire n15981;
    wire n15984;
    wire n15987;
    wire n15990;
    wire n15993;
    wire n15996;
    wire n15999;
    wire n16002;
    wire n16005;
    wire n16008;
    wire n16011;
    wire n16013;
    wire n16016;
    wire n16019;
    wire n16022;
    wire n16025;
    wire n16028;
    wire n16031;
    wire n16034;
    wire n16037;
    wire n16040;
    wire n16043;
    wire n16046;
    wire n16049;
    wire n16052;
    wire n16055;
    wire n16058;
    wire n16061;
    wire n16064;
    wire n16067;
    wire n16070;
    wire n16073;
    wire n16076;
    wire n16079;
    wire n16082;
    wire n16085;
    wire n16088;
    wire n16091;
    wire n16094;
    wire n16097;
    wire n16100;
    wire n16103;
    wire n16106;
    wire n16109;
    wire n16112;
    wire n16115;
    wire n16118;
    wire n16121;
    wire n16124;
    wire n16127;
    wire n16130;
    wire n16134;
    wire n16137;
    wire n16140;
    wire n16143;
    wire n16146;
    wire n16149;
    wire n16152;
    wire n16155;
    wire n16158;
    wire n16161;
    wire n16164;
    wire n16167;
    wire n16170;
    wire n16173;
    wire n16176;
    wire n16179;
    wire n16182;
    wire n16185;
    wire n16188;
    wire n16191;
    wire n16194;
    wire n16197;
    wire n16200;
    wire n16203;
    wire n16206;
    wire n16209;
    wire n16212;
    wire n16215;
    wire n16218;
    wire n16221;
    wire n16224;
    wire n16227;
    wire n16230;
    wire n16233;
    wire n16236;
    wire n16239;
    wire n16242;
    wire n16245;
    wire n16248;
    wire n16251;
    wire n16254;
    wire n16257;
    wire n16260;
    wire n16263;
    wire n16266;
    wire n16269;
    wire n16272;
    wire n16275;
    wire n16278;
    wire n16281;
    wire n16284;
    wire n16287;
    wire n16290;
    wire n16293;
    wire n16296;
    wire n16299;
    wire n16302;
    wire n16305;
    wire n16308;
    wire n16311;
    wire n16314;
    wire n16317;
    wire n16320;
    wire n16323;
    wire n16326;
    wire n16329;
    wire n16332;
    wire n16335;
    wire n16338;
    wire n16341;
    wire n16344;
    wire n16347;
    wire n16350;
    wire n16353;
    wire n16356;
    wire n16359;
    wire n16362;
    wire n16365;
    wire n16368;
    wire n16371;
    wire n16374;
    wire n16377;
    wire n16380;
    wire n16383;
    wire n16386;
    wire n16389;
    wire n16392;
    wire n16395;
    wire n16398;
    wire n16401;
    wire n16404;
    wire n16407;
    wire n16410;
    wire n16413;
    wire n16416;
    wire n16419;
    wire n16422;
    wire n16425;
    wire n16428;
    wire n16431;
    wire n16434;
    wire n16437;
    wire n16440;
    wire n16443;
    wire n16446;
    wire n16449;
    wire n16452;
    wire n16455;
    wire n16458;
    wire n16461;
    wire n16464;
    wire n16467;
    wire n16470;
    wire n16473;
    wire n16476;
    wire n16479;
    wire n16482;
    wire n16485;
    wire n16488;
    wire n16491;
    wire n16494;
    wire n16497;
    wire n16500;
    wire n16503;
    wire n16506;
    wire n16509;
    wire n16512;
    wire n16515;
    wire n16518;
    wire n16521;
    wire n16524;
    wire n16527;
    wire n16530;
    wire n16533;
    wire n16536;
    wire n16539;
    wire n16542;
    wire n16545;
    wire n16548;
    wire n16551;
    wire n16554;
    wire n16557;
    wire n16560;
    wire n16563;
    wire n16566;
    wire n16569;
    wire n16572;
    wire n16575;
    wire n16578;
    wire n16581;
    wire n16584;
    wire n16587;
    wire n16590;
    wire n16593;
    wire n16596;
    wire n16599;
    wire n16602;
    wire n16605;
    wire n16608;
    wire n16611;
    wire n16614;
    wire n16617;
    wire n16620;
    wire n16623;
    wire n16626;
    wire n16629;
    wire n16632;
    wire n16635;
    wire n16638;
    wire n16641;
    wire n16644;
    wire n16647;
    wire n16650;
    wire n16653;
    wire n16656;
    wire n16659;
    wire n16662;
    wire n16665;
    wire n16668;
    wire n16671;
    wire n16674;
    wire n16677;
    wire n16680;
    wire n16683;
    wire n16686;
    wire n16689;
    wire n16692;
    wire n16695;
    wire n16698;
    wire n16701;
    wire n16704;
    wire n16707;
    wire n16710;
    wire n16713;
    wire n16716;
    wire n16719;
    wire n16722;
    wire n16725;
    wire n16728;
    wire n16731;
    wire n16734;
    wire n16737;
    wire n16740;
    wire n16743;
    wire n16746;
    wire n16749;
    wire n16752;
    wire n16755;
    wire n16758;
    wire n16761;
    wire n16764;
    wire n16767;
    wire n16770;
    wire n16773;
    wire n16776;
    wire n16779;
    wire n16782;
    wire n16785;
    wire n16788;
    wire n16791;
    wire n16793;
    wire n16796;
    wire n16800;
    wire n16803;
    wire n16806;
    wire n16809;
    wire n16812;
    wire n16815;
    wire n16818;
    wire n16821;
    wire n16824;
    wire n16827;
    wire n16830;
    wire n16833;
    wire n16836;
    wire n16839;
    wire n16842;
    wire n16845;
    wire n16848;
    wire n16851;
    wire n16854;
    wire n16857;
    wire n16860;
    wire n16863;
    wire n16866;
    wire n16869;
    wire n16872;
    wire n16875;
    wire n16878;
    wire n16881;
    wire n16884;
    wire n16887;
    wire n16890;
    wire n16893;
    wire n16896;
    wire n16899;
    wire n16902;
    wire n16905;
    wire n16908;
    wire n16911;
    wire n16914;
    wire n16917;
    wire n16920;
    wire n16923;
    wire n16926;
    wire n16929;
    wire n16932;
    wire n16935;
    wire n16938;
    wire n16941;
    wire n16944;
    wire n16947;
    wire n16950;
    wire n16953;
    wire n16956;
    wire n16959;
    wire n16962;
    wire n16965;
    wire n16968;
    wire n16971;
    wire n16974;
    wire n16977;
    wire n16980;
    wire n16983;
    wire n16986;
    wire n16989;
    wire n16992;
    wire n16995;
    wire n16998;
    wire n17001;
    wire n17004;
    wire n17007;
    wire n17010;
    wire n17013;
    wire n17016;
    wire n17019;
    wire n17022;
    wire n17025;
    wire n17028;
    wire n17031;
    wire n17034;
    wire n17037;
    wire n17040;
    wire n17043;
    wire n17046;
    wire n17049;
    wire n17052;
    wire n17055;
    wire n17058;
    wire n17061;
    wire n17064;
    wire n17067;
    wire n17070;
    wire n17073;
    wire n17076;
    wire n17079;
    wire n17082;
    wire n17085;
    wire n17088;
    wire n17091;
    wire n17094;
    wire n17097;
    wire n17100;
    wire n17103;
    wire n17106;
    wire n17109;
    wire n17112;
    wire n17115;
    wire n17118;
    wire n17121;
    wire n17124;
    wire n17127;
    wire n17130;
    wire n17133;
    wire n17136;
    wire n17139;
    wire n17142;
    wire n17145;
    wire n17148;
    wire n17151;
    wire n17154;
    wire n17157;
    wire n17160;
    wire n17163;
    wire n17166;
    wire n17169;
    wire n17172;
    wire n17175;
    wire n17178;
    wire n17181;
    wire n17184;
    wire n17187;
    wire n17190;
    wire n17193;
    wire n17196;
    wire n17199;
    wire n17202;
    wire n17205;
    wire n17208;
    wire n17211;
    wire n17214;
    wire n17217;
    wire n17220;
    wire n17223;
    wire n17226;
    wire n17229;
    wire n17232;
    wire n17235;
    wire n17238;
    wire n17241;
    wire n17244;
    wire n17247;
    wire n17250;
    wire n17253;
    wire n17256;
    wire n17259;
    wire n17262;
    wire n17265;
    wire n17268;
    wire n17271;
    wire n17274;
    wire n17277;
    wire n17280;
    wire n17283;
    wire n17286;
    wire n17289;
    wire n17292;
    wire n17295;
    wire n17298;
    wire n17301;
    wire n17304;
    wire n17307;
    wire n17310;
    wire n17313;
    wire n17316;
    wire n17319;
    wire n17322;
    wire n17325;
    wire n17328;
    wire n17331;
    wire n17334;
    wire n17337;
    wire n17340;
    wire n17343;
    wire n17346;
    wire n17349;
    wire n17352;
    wire n17355;
    wire n17358;
    wire n17361;
    wire n17364;
    wire n17367;
    wire n17370;
    wire n17373;
    wire n17376;
    wire n17379;
    wire n17382;
    wire n17385;
    wire n17388;
    wire n17391;
    wire n17394;
    wire n17397;
    wire n17400;
    wire n17403;
    wire n17406;
    wire n17409;
    wire n17412;
    wire n17415;
    wire n17418;
    wire n17421;
    wire n17424;
    wire n17427;
    wire n17430;
    wire n17433;
    wire n17436;
    wire n17439;
    wire n17442;
    wire n17445;
    wire n17448;
    wire n17451;
    wire n17454;
    wire n17457;
    wire n17460;
    wire n17463;
    wire n17466;
    wire n17469;
    wire n17472;
    wire n17475;
    wire n17478;
    wire n17481;
    wire n17484;
    wire n17487;
    wire n17490;
    wire n17493;
    wire n17496;
    wire n17499;
    wire n17502;
    wire n17505;
    wire n17508;
    wire n17511;
    wire n17514;
    wire n17517;
    wire n17520;
    wire n17523;
    wire n17526;
    wire n17529;
    wire n17532;
    wire n17535;
    wire n17538;
    wire n17541;
    wire n17544;
    wire n17547;
    wire n17550;
    wire n17553;
    wire n17556;
    wire n17559;
    wire n17562;
    wire n17565;
    wire n17568;
    wire n17571;
    wire n17574;
    wire n17577;
    wire n17580;
    wire n17583;
    wire n17586;
    wire n17589;
    wire n17592;
    wire n17595;
    wire n17598;
    wire n17601;
    wire n17604;
    wire n17607;
    wire n17610;
    wire n17613;
    wire n17616;
    wire n17619;
    wire n17622;
    wire n17625;
    wire n17628;
    wire n17631;
    wire n17634;
    wire n17637;
    wire n17640;
    wire n17643;
    wire n17646;
    wire n17649;
    wire n17652;
    wire n17655;
    wire n17658;
    wire n17661;
    wire n17664;
    wire n17667;
    wire n17670;
    wire n17673;
    wire n17676;
    wire n17679;
    wire n17682;
    wire n17685;
    wire n17688;
    wire n17691;
    wire n17694;
    wire n17697;
    wire n17700;
    wire n17703;
    wire n17706;
    wire n17709;
    wire n17712;
    wire n17715;
    wire n17718;
    wire n17721;
    wire n17724;
    wire n17727;
    wire n17730;
    wire n17733;
    wire n17736;
    wire n17739;
    wire n17742;
    wire n17745;
    wire n17748;
    wire n17751;
    wire n17754;
    wire n17757;
    wire n17760;
    wire n17763;
    wire n17766;
    wire n17769;
    wire n17772;
    wire n17775;
    wire n17778;
    wire n17781;
    wire n17784;
    wire n17787;
    wire n17790;
    wire n17793;
    wire n17796;
    wire n17799;
    wire n17802;
    wire n17805;
    wire n17808;
    wire n17811;
    wire n17814;
    wire n17817;
    wire n17820;
    wire n17823;
    wire n17826;
    wire n17829;
    wire n17832;
    wire n17835;
    wire n17838;
    wire n17841;
    wire n17843;
    wire n17846;
    wire n17849;
    wire n17852;
    wire n17856;
    wire n17859;
    wire n17862;
    wire n17865;
    wire n17868;
    wire n17871;
    wire n17874;
    wire n17877;
    wire n17880;
    wire n17883;
    wire n17886;
    wire n17889;
    wire n17892;
    wire n17895;
    wire n17898;
    wire n17901;
    wire n17904;
    wire n17907;
    wire n17910;
    wire n17913;
    wire n17916;
    wire n17919;
    wire n17922;
    wire n17925;
    wire n17928;
    wire n17931;
    wire n17934;
    wire n17937;
    wire n17940;
    wire n17943;
    wire n17946;
    wire n17949;
    wire n17952;
    wire n17955;
    wire n17958;
    wire n17961;
    wire n17964;
    wire n17967;
    wire n17970;
    wire n17973;
    wire n17976;
    wire n17979;
    wire n17982;
    wire n17985;
    wire n17988;
    wire n17991;
    wire n17993;
    wire n17997;
    wire n18000;
    wire n18003;
    wire n18006;
    wire n18009;
    wire n18012;
    wire n18015;
    wire n18018;
    wire n18021;
    wire n18024;
    wire n18027;
    wire n18030;
    wire n18033;
    wire n18036;
    wire n18039;
    wire n18042;
    wire n18045;
    wire n18048;
    wire n18051;
    wire n18054;
    wire n18057;
    wire n18060;
    wire n18063;
    wire n18066;
    wire n18069;
    wire n18072;
    wire n18075;
    wire n18078;
    wire n18081;
    wire n18084;
    wire n18087;
    wire n18090;
    wire n18093;
    wire n18096;
    wire n18099;
    wire n18102;
    wire n18105;
    wire n18108;
    wire n18111;
    wire n18114;
    wire n18117;
    wire n18120;
    wire n18123;
    wire n18126;
    wire n18129;
    wire n18132;
    wire n18135;
    wire n18138;
    wire n18141;
    wire n18144;
    wire n18147;
    wire n18150;
    wire n18153;
    wire n18156;
    wire n18159;
    wire n18162;
    wire n18165;
    wire n18168;
    wire n18171;
    wire n18174;
    wire n18177;
    wire n18180;
    wire n18183;
    wire n18186;
    wire n18189;
    wire n18192;
    wire n18195;
    wire n18198;
    wire n18201;
    wire n18204;
    wire n18207;
    wire n18210;
    wire n18213;
    wire n18216;
    wire n18219;
    wire n18222;
    wire n18225;
    wire n18228;
    wire n18231;
    wire n18234;
    wire n18237;
    wire n18240;
    wire n18243;
    wire n18246;
    wire n18249;
    wire n18252;
    wire n18255;
    wire n18258;
    wire n18261;
    wire n18264;
    wire n18267;
    wire n18270;
    wire n18273;
    wire n18276;
    wire n18279;
    wire n18282;
    wire n18285;
    wire n18288;
    wire n18291;
    wire n18294;
    wire n18297;
    wire n18300;
    wire n18303;
    wire n18306;
    wire n18309;
    wire n18312;
    wire n18315;
    wire n18318;
    wire n18321;
    wire n18324;
    wire n18327;
    wire n18330;
    wire n18333;
    wire n18336;
    wire n18339;
    wire n18342;
    wire n18345;
    wire n18348;
    wire n18351;
    wire n18354;
    wire n18357;
    wire n18360;
    wire n18363;
    wire n18366;
    wire n18369;
    wire n18372;
    wire n18375;
    wire n18378;
    wire n18381;
    wire n18384;
    wire n18387;
    wire n18390;
    wire n18393;
    wire n18396;
    wire n18399;
    wire n18402;
    wire n18405;
    wire n18408;
    wire n18411;
    wire n18414;
    wire n18417;
    wire n18420;
    wire n18423;
    wire n18426;
    wire n18429;
    wire n18432;
    wire n18435;
    wire n18438;
    wire n18441;
    wire n18444;
    wire n18447;
    wire n18450;
    wire n18453;
    wire n18456;
    wire n18459;
    wire n18462;
    wire n18465;
    wire n18468;
    wire n18471;
    wire n18474;
    wire n18477;
    wire n18480;
    wire n18483;
    wire n18486;
    wire n18489;
    wire n18492;
    wire n18495;
    wire n18498;
    wire n18501;
    wire n18504;
    wire n18507;
    wire n18510;
    wire n18513;
    wire n18516;
    wire n18519;
    wire n18522;
    wire n18525;
    wire n18528;
    wire n18531;
    wire n18534;
    wire n18537;
    wire n18540;
    wire n18543;
    wire n18546;
    wire n18549;
    wire n18552;
    wire n18555;
    wire n18558;
    wire n18561;
    wire n18564;
    wire n18567;
    wire n18570;
    wire n18573;
    wire n18576;
    wire n18579;
    wire n18582;
    wire n18585;
    wire n18588;
    wire n18591;
    wire n18594;
    wire n18597;
    wire n18600;
    wire n18603;
    wire n18606;
    wire n18609;
    wire n18612;
    wire n18615;
    wire n18618;
    wire n18621;
    wire n18624;
    wire n18627;
    wire n18630;
    wire n18633;
    wire n18636;
    wire n18639;
    wire n18642;
    wire n18645;
    wire n18648;
    wire n18651;
    wire n18654;
    wire n18657;
    wire n18660;
    wire n18663;
    wire n18666;
    wire n18669;
    wire n18672;
    wire n18675;
    wire n18678;
    wire n18681;
    wire n18684;
    wire n18687;
    wire n18690;
    wire n18693;
    wire n18696;
    wire n18699;
    wire n18702;
    wire n18705;
    wire n18708;
    wire n18711;
    wire n18714;
    wire n18717;
    wire n18720;
    wire n18723;
    wire n18726;
    wire n18729;
    wire n18732;
    wire n18735;
    wire n18738;
    wire n18741;
    wire n18744;
    wire n18747;
    wire n18750;
    wire n18753;
    wire n18756;
    wire n18759;
    wire n18762;
    wire n18765;
    wire n18768;
    wire n18771;
    wire n18774;
    wire n18777;
    wire n18780;
    wire n18783;
    wire n18786;
    wire n18789;
    wire n18792;
    wire n18795;
    wire n18798;
    wire n18801;
    wire n18804;
    wire n18807;
    wire n18810;
    wire n18813;
    wire n18816;
    wire n18819;
    wire n18822;
    wire n18825;
    wire n18828;
    wire n18831;
    wire n18834;
    wire n18837;
    wire n18840;
    wire n18843;
    wire n18846;
    wire n18849;
    wire n18852;
    wire n18855;
    wire n18858;
    wire n18861;
    wire n18864;
    wire n18867;
    wire n18870;
    wire n18873;
    wire n18876;
    wire n18879;
    wire n18882;
    wire n18885;
    wire n18888;
    wire n18890;
    wire n18893;
    wire n18896;
    wire n18899;
    wire n18903;
    wire n18906;
    wire n18909;
    wire n18912;
    wire n18915;
    wire n18918;
    wire n18921;
    wire n18924;
    wire n18927;
    wire n18930;
    wire n18933;
    wire n18936;
    wire n18939;
    wire n18942;
    wire n18945;
    wire n18948;
    wire n18951;
    wire n18954;
    wire n18957;
    wire n18960;
    wire n18963;
    wire n18966;
    wire n18969;
    wire n18972;
    wire n18975;
    wire n18978;
    wire n18981;
    wire n18984;
    wire n18987;
    wire n18990;
    wire n18993;
    wire n18996;
    wire n18999;
    wire n19002;
    wire n19005;
    wire n19008;
    wire n19011;
    wire n19014;
    wire n19017;
    wire n19020;
    wire n19023;
    wire n19026;
    wire n19029;
    wire n19032;
    wire n19035;
    wire n19038;
    wire n19041;
    wire n19044;
    wire n19047;
    wire n19050;
    wire n19053;
    wire n19056;
    wire n19059;
    wire n19062;
    wire n19065;
    wire n19068;
    wire n19071;
    wire n19074;
    wire n19077;
    wire n19080;
    wire n19083;
    wire n19086;
    wire n19089;
    wire n19092;
    wire n19095;
    wire n19098;
    wire n19101;
    wire n19104;
    wire n19107;
    wire n19110;
    wire n19113;
    wire n19116;
    wire n19119;
    wire n19122;
    wire n19125;
    wire n19128;
    wire n19131;
    wire n19134;
    wire n19137;
    wire n19140;
    wire n19143;
    wire n19146;
    wire n19149;
    wire n19152;
    wire n19155;
    wire n19158;
    wire n19161;
    wire n19164;
    wire n19167;
    wire n19170;
    wire n19173;
    wire n19176;
    wire n19179;
    wire n19182;
    wire n19185;
    wire n19188;
    wire n19191;
    wire n19194;
    wire n19197;
    wire n19200;
    wire n19203;
    wire n19206;
    wire n19209;
    wire n19212;
    wire n19215;
    wire n19218;
    wire n19221;
    wire n19224;
    wire n19227;
    wire n19230;
    wire n19233;
    wire n19236;
    wire n19239;
    wire n19242;
    wire n19245;
    wire n19248;
    wire n19251;
    wire n19254;
    wire n19257;
    wire n19260;
    wire n19263;
    wire n19266;
    wire n19269;
    wire n19272;
    wire n19275;
    wire n19278;
    wire n19281;
    wire n19284;
    wire n19287;
    wire n19290;
    wire n19293;
    wire n19296;
    wire n19299;
    wire n19302;
    wire n19305;
    wire n19308;
    wire n19311;
    wire n19314;
    wire n19317;
    wire n19320;
    wire n19323;
    wire n19326;
    wire n19329;
    wire n19332;
    wire n19335;
    wire n19338;
    wire n19341;
    wire n19344;
    wire n19347;
    wire n19350;
    wire n19353;
    wire n19356;
    wire n19359;
    wire n19362;
    wire n19365;
    wire n19368;
    wire n19371;
    wire n19374;
    wire n19377;
    wire n19380;
    wire n19383;
    wire n19386;
    wire n19389;
    wire n19392;
    wire n19395;
    wire n19398;
    wire n19401;
    wire n19404;
    wire n19407;
    wire n19410;
    wire n19413;
    wire n19416;
    wire n19419;
    wire n19422;
    wire n19425;
    wire n19428;
    wire n19431;
    wire n19434;
    wire n19437;
    wire n19440;
    wire n19443;
    wire n19446;
    wire n19449;
    wire n19452;
    wire n19455;
    wire n19458;
    wire n19461;
    wire n19464;
    wire n19467;
    wire n19470;
    wire n19473;
    wire n19476;
    wire n19479;
    wire n19482;
    wire n19485;
    wire n19488;
    wire n19491;
    wire n19494;
    wire n19497;
    wire n19500;
    wire n19503;
    wire n19506;
    wire n19509;
    wire n19512;
    wire n19515;
    wire n19518;
    wire n19521;
    wire n19524;
    wire n19527;
    wire n19530;
    wire n19533;
    wire n19536;
    wire n19539;
    wire n19542;
    wire n19545;
    wire n19548;
    wire n19551;
    wire n19554;
    wire n19557;
    wire n19560;
    wire n19563;
    wire n19566;
    wire n19569;
    wire n19572;
    wire n19575;
    wire n19578;
    wire n19581;
    wire n19584;
    wire n19587;
    wire n19590;
    wire n19593;
    wire n19596;
    wire n19599;
    wire n19602;
    wire n19605;
    wire n19608;
    wire n19611;
    wire n19614;
    wire n19617;
    wire n19620;
    wire n19623;
    wire n19626;
    wire n19629;
    wire n19632;
    wire n19635;
    wire n19638;
    wire n19641;
    wire n19644;
    wire n19647;
    wire n19650;
    wire n19653;
    wire n19656;
    wire n19659;
    wire n19662;
    wire n19665;
    wire n19668;
    wire n19671;
    wire n19674;
    wire n19677;
    wire n19680;
    wire n19683;
    wire n19686;
    wire n19689;
    wire n19692;
    wire n19695;
    wire n19698;
    wire n19701;
    wire n19704;
    wire n19707;
    wire n19710;
    wire n19713;
    wire n19716;
    wire n19719;
    wire n19722;
    wire n19725;
    wire n19728;
    wire n19731;
    wire n19734;
    wire n19737;
    wire n19740;
    wire n19743;
    wire n19746;
    wire n19749;
    wire n19752;
    wire n19755;
    wire n19758;
    wire n19761;
    wire n19764;
    wire n19767;
    wire n19770;
    wire n19773;
    wire n19776;
    wire n19779;
    wire n19782;
    wire n19785;
    wire n19788;
    wire n19791;
    wire n19794;
    wire n19797;
    wire n19800;
    wire n19803;
    wire n19806;
    wire n19809;
    wire n19812;
    wire n19815;
    wire n19818;
    wire n19821;
    wire n19824;
    wire n19827;
    wire n19830;
    wire n19833;
    wire n19836;
    wire n19839;
    wire n19842;
    wire n19845;
    wire n19848;
    wire n19851;
    wire n19854;
    wire n19857;
    wire n19860;
    wire n19863;
    wire n19866;
    wire n19869;
    wire n19872;
    wire n19875;
    wire n19878;
    wire n19881;
    wire n19884;
    wire n19887;
    wire n19890;
    wire n19893;
    wire n19896;
    wire n19899;
    wire n19902;
    wire n19904;
    wire n19907;
    wire n19910;
    wire n19913;
    wire n19917;
    wire n19920;
    wire n19923;
    wire n19926;
    wire n19929;
    wire n19932;
    wire n19935;
    wire n19938;
    wire n19941;
    wire n19944;
    wire n19947;
    wire n19950;
    wire n19953;
    wire n19956;
    wire n19959;
    wire n19962;
    wire n19965;
    wire n19968;
    wire n19971;
    wire n19974;
    wire n19977;
    wire n19980;
    wire n19983;
    wire n19986;
    wire n19989;
    wire n19992;
    wire n19995;
    wire n19998;
    wire n20001;
    wire n20004;
    wire n20007;
    wire n20010;
    wire n20013;
    wire n20016;
    wire n20019;
    wire n20022;
    wire n20025;
    wire n20028;
    wire n20031;
    wire n20034;
    wire n20037;
    wire n20040;
    wire n20043;
    wire n20046;
    wire n20049;
    wire n20052;
    wire n20055;
    wire n20058;
    wire n20061;
    wire n20064;
    wire n20067;
    wire n20070;
    wire n20073;
    wire n20076;
    wire n20079;
    wire n20082;
    wire n20085;
    wire n20088;
    wire n20091;
    wire n20094;
    wire n20097;
    wire n20100;
    wire n20103;
    wire n20106;
    wire n20109;
    wire n20112;
    wire n20115;
    wire n20118;
    wire n20121;
    wire n20124;
    wire n20127;
    wire n20130;
    wire n20133;
    wire n20136;
    wire n20139;
    wire n20142;
    wire n20145;
    wire n20148;
    wire n20151;
    wire n20154;
    wire n20157;
    wire n20160;
    wire n20163;
    wire n20166;
    wire n20169;
    wire n20172;
    wire n20175;
    wire n20178;
    wire n20181;
    wire n20184;
    wire n20187;
    wire n20190;
    wire n20193;
    wire n20196;
    wire n20199;
    wire n20202;
    wire n20205;
    wire n20208;
    wire n20211;
    wire n20214;
    wire n20217;
    wire n20220;
    wire n20223;
    wire n20226;
    wire n20229;
    wire n20232;
    wire n20235;
    wire n20238;
    wire n20241;
    wire n20244;
    wire n20247;
    wire n20250;
    wire n20253;
    wire n20256;
    wire n20259;
    wire n20262;
    wire n20265;
    wire n20268;
    wire n20271;
    wire n20274;
    wire n20277;
    wire n20280;
    wire n20283;
    wire n20286;
    wire n20289;
    wire n20292;
    wire n20295;
    wire n20298;
    wire n20301;
    wire n20304;
    wire n20307;
    wire n20310;
    wire n20313;
    wire n20316;
    wire n20319;
    wire n20322;
    wire n20325;
    wire n20328;
    wire n20331;
    wire n20334;
    wire n20337;
    wire n20340;
    wire n20343;
    wire n20346;
    wire n20349;
    wire n20352;
    wire n20355;
    wire n20358;
    wire n20361;
    wire n20364;
    wire n20367;
    wire n20370;
    wire n20373;
    wire n20376;
    wire n20379;
    wire n20382;
    wire n20385;
    wire n20388;
    wire n20391;
    wire n20394;
    wire n20397;
    wire n20400;
    wire n20403;
    wire n20406;
    wire n20409;
    wire n20412;
    wire n20415;
    wire n20418;
    wire n20421;
    wire n20424;
    wire n20427;
    wire n20430;
    wire n20433;
    wire n20436;
    wire n20439;
    wire n20442;
    wire n20445;
    wire n20448;
    wire n20451;
    wire n20454;
    wire n20457;
    wire n20460;
    wire n20463;
    wire n20466;
    wire n20469;
    wire n20472;
    wire n20475;
    wire n20478;
    wire n20481;
    wire n20484;
    wire n20487;
    wire n20490;
    wire n20493;
    wire n20496;
    wire n20499;
    wire n20502;
    wire n20505;
    wire n20508;
    wire n20511;
    wire n20514;
    wire n20517;
    wire n20520;
    wire n20523;
    wire n20526;
    wire n20529;
    wire n20532;
    wire n20535;
    wire n20538;
    wire n20541;
    wire n20544;
    wire n20547;
    wire n20550;
    wire n20553;
    wire n20556;
    wire n20559;
    wire n20562;
    wire n20565;
    wire n20568;
    wire n20571;
    wire n20574;
    wire n20577;
    wire n20580;
    wire n20583;
    wire n20586;
    wire n20589;
    wire n20592;
    wire n20595;
    wire n20598;
    wire n20601;
    wire n20604;
    wire n20607;
    wire n20610;
    wire n20613;
    wire n20616;
    wire n20619;
    wire n20622;
    wire n20625;
    wire n20628;
    wire n20631;
    wire n20634;
    wire n20637;
    wire n20640;
    wire n20643;
    wire n20646;
    wire n20649;
    wire n20652;
    wire n20655;
    wire n20658;
    wire n20661;
    wire n20664;
    wire n20667;
    wire n20670;
    wire n20673;
    wire n20676;
    wire n20679;
    wire n20682;
    wire n20685;
    wire n20688;
    wire n20691;
    wire n20694;
    wire n20697;
    wire n20700;
    wire n20703;
    wire n20706;
    wire n20709;
    wire n20712;
    wire n20715;
    wire n20718;
    wire n20721;
    wire n20724;
    wire n20727;
    wire n20730;
    wire n20733;
    wire n20736;
    wire n20739;
    wire n20742;
    wire n20745;
    wire n20748;
    wire n20751;
    wire n20754;
    wire n20757;
    wire n20760;
    wire n20763;
    wire n20766;
    wire n20769;
    wire n20772;
    wire n20775;
    wire n20778;
    wire n20781;
    wire n20784;
    wire n20787;
    wire n20790;
    wire n20793;
    wire n20796;
    wire n20799;
    wire n20802;
    wire n20805;
    wire n20808;
    wire n20811;
    wire n20814;
    wire n20817;
    wire n20820;
    wire n20823;
    wire n20826;
    wire n20829;
    wire n20832;
    wire n20835;
    wire n20838;
    wire n20841;
    wire n20844;
    wire n20847;
    wire n20850;
    wire n20853;
    wire n20856;
    wire n20859;
    wire n20862;
    wire n20865;
    wire n20868;
    wire n20871;
    wire n20874;
    wire n20877;
    wire n20880;
    wire n20883;
    wire n20886;
    wire n20889;
    wire n20892;
    wire n20895;
    wire n20898;
    wire n20901;
    wire n20904;
    wire n20907;
    wire n20910;
    wire n20913;
    wire n20916;
    wire n20919;
    wire n20922;
    wire n20925;
    wire n20928;
    wire n20931;
    wire n20934;
    wire n20937;
    wire n20940;
    wire n20943;
    wire n20946;
    wire n20949;
    wire n20952;
    wire n20954;
    wire n20957;
    wire n20960;
    wire n20963;
    wire n20967;
    wire n20970;
    wire n20973;
    wire n20976;
    wire n20979;
    wire n20982;
    wire n20985;
    wire n20988;
    wire n20991;
    wire n20994;
    wire n20997;
    wire n21000;
    wire n21003;
    wire n21006;
    wire n21009;
    wire n21012;
    wire n21015;
    wire n21018;
    wire n21021;
    wire n21024;
    wire n21027;
    wire n21030;
    wire n21033;
    wire n21036;
    wire n21039;
    wire n21042;
    wire n21045;
    wire n21048;
    wire n21051;
    wire n21054;
    wire n21057;
    wire n21060;
    wire n21063;
    wire n21066;
    wire n21069;
    wire n21072;
    wire n21075;
    wire n21078;
    wire n21081;
    wire n21084;
    wire n21087;
    wire n21090;
    wire n21093;
    wire n21096;
    wire n21099;
    wire n21102;
    wire n21105;
    wire n21108;
    wire n21110;
    wire n21114;
    wire n21117;
    wire n21120;
    wire n21123;
    wire n21126;
    wire n21129;
    wire n21132;
    wire n21135;
    wire n21138;
    wire n21141;
    wire n21144;
    wire n21147;
    wire n21150;
    wire n21153;
    wire n21156;
    wire n21159;
    wire n21162;
    wire n21165;
    wire n21168;
    wire n21171;
    wire n21174;
    wire n21177;
    wire n21180;
    wire n21183;
    wire n21186;
    wire n21189;
    wire n21192;
    wire n21195;
    wire n21198;
    wire n21201;
    wire n21204;
    wire n21207;
    wire n21210;
    wire n21213;
    wire n21216;
    wire n21219;
    wire n21222;
    wire n21225;
    wire n21228;
    wire n21231;
    wire n21234;
    wire n21237;
    wire n21240;
    wire n21243;
    wire n21246;
    wire n21249;
    wire n21252;
    wire n21255;
    wire n21258;
    wire n21261;
    wire n21264;
    wire n21267;
    wire n21270;
    wire n21273;
    wire n21276;
    wire n21279;
    wire n21282;
    wire n21285;
    wire n21288;
    wire n21291;
    wire n21294;
    wire n21297;
    wire n21300;
    wire n21303;
    wire n21306;
    wire n21309;
    wire n21312;
    wire n21315;
    wire n21318;
    wire n21321;
    wire n21324;
    wire n21327;
    wire n21330;
    wire n21333;
    wire n21336;
    wire n21339;
    wire n21342;
    wire n21345;
    wire n21348;
    wire n21351;
    wire n21354;
    wire n21357;
    wire n21360;
    wire n21363;
    wire n21366;
    wire n21369;
    wire n21372;
    wire n21375;
    wire n21378;
    wire n21381;
    wire n21384;
    wire n21387;
    wire n21390;
    wire n21393;
    wire n21396;
    wire n21399;
    wire n21402;
    wire n21405;
    wire n21408;
    wire n21411;
    wire n21414;
    wire n21417;
    wire n21420;
    wire n21423;
    wire n21426;
    wire n21429;
    wire n21432;
    wire n21435;
    wire n21438;
    wire n21441;
    wire n21444;
    wire n21447;
    wire n21450;
    wire n21453;
    wire n21456;
    wire n21459;
    wire n21462;
    wire n21465;
    wire n21468;
    wire n21471;
    wire n21474;
    wire n21477;
    wire n21480;
    wire n21483;
    wire n21486;
    wire n21489;
    wire n21492;
    wire n21495;
    wire n21498;
    wire n21501;
    wire n21504;
    wire n21507;
    wire n21510;
    wire n21513;
    wire n21516;
    wire n21519;
    wire n21522;
    wire n21525;
    wire n21528;
    wire n21531;
    wire n21534;
    wire n21537;
    wire n21540;
    wire n21543;
    wire n21546;
    wire n21549;
    wire n21552;
    wire n21555;
    wire n21558;
    wire n21561;
    wire n21564;
    wire n21567;
    wire n21570;
    wire n21573;
    wire n21576;
    wire n21579;
    wire n21582;
    wire n21585;
    wire n21588;
    wire n21591;
    wire n21594;
    wire n21597;
    wire n21600;
    wire n21603;
    wire n21606;
    wire n21609;
    wire n21612;
    wire n21615;
    wire n21618;
    wire n21621;
    wire n21624;
    wire n21627;
    wire n21630;
    wire n21633;
    wire n21636;
    wire n21639;
    wire n21642;
    wire n21645;
    wire n21648;
    wire n21651;
    wire n21654;
    wire n21657;
    wire n21660;
    wire n21663;
    wire n21666;
    wire n21669;
    wire n21672;
    wire n21675;
    wire n21678;
    wire n21681;
    wire n21684;
    wire n21687;
    wire n21690;
    wire n21693;
    wire n21696;
    wire n21699;
    wire n21702;
    wire n21705;
    wire n21708;
    wire n21711;
    wire n21714;
    wire n21717;
    wire n21720;
    wire n21723;
    wire n21726;
    wire n21729;
    wire n21732;
    wire n21735;
    wire n21738;
    wire n21741;
    wire n21744;
    wire n21747;
    wire n21750;
    wire n21753;
    wire n21756;
    wire n21759;
    wire n21762;
    wire n21765;
    wire n21768;
    wire n21771;
    wire n21774;
    wire n21777;
    wire n21780;
    wire n21783;
    wire n21786;
    wire n21789;
    wire n21792;
    wire n21795;
    wire n21798;
    wire n21801;
    wire n21804;
    wire n21807;
    wire n21810;
    wire n21813;
    wire n21816;
    wire n21819;
    wire n21822;
    wire n21825;
    wire n21828;
    wire n21831;
    wire n21834;
    wire n21837;
    wire n21840;
    wire n21843;
    wire n21846;
    wire n21849;
    wire n21852;
    wire n21855;
    wire n21858;
    wire n21861;
    wire n21864;
    wire n21867;
    wire n21870;
    wire n21873;
    wire n21876;
    wire n21879;
    wire n21882;
    wire n21885;
    wire n21888;
    wire n21891;
    wire n21894;
    wire n21897;
    wire n21900;
    wire n21903;
    wire n21906;
    wire n21909;
    wire n21912;
    wire n21915;
    wire n21918;
    wire n21921;
    wire n21924;
    wire n21927;
    wire n21930;
    wire n21933;
    wire n21936;
    wire n21939;
    wire n21942;
    wire n21945;
    wire n21948;
    wire n21951;
    wire n21954;
    wire n21957;
    wire n21960;
    wire n21963;
    wire n21966;
    wire n21969;
    wire n21972;
    wire n21975;
    wire n21978;
    wire n21981;
    wire n21984;
    wire n21987;
    wire n21990;
    wire n21993;
    wire n21996;
    wire n21999;
    wire n22002;
    wire n22005;
    wire n22008;
    wire n22011;
    wire n22014;
    wire n22017;
    wire n22020;
    wire n22023;
    wire n22026;
    wire n22029;
    wire n22032;
    wire n22035;
    wire n22038;
    wire n22041;
    wire n22044;
    wire n22047;
    wire n22050;
    wire n22053;
    wire n22056;
    wire n22059;
    wire n22062;
    wire n22065;
    wire n22068;
    wire n22071;
    wire n22074;
    wire n22077;
    wire n22080;
    wire n22083;
    wire n22086;
    wire n22089;
    wire n22091;
    wire n22094;
    wire n22097;
    wire n22100;
    wire n22104;
    wire n22107;
    wire n22110;
    wire n22113;
    wire n22116;
    wire n22119;
    wire n22122;
    wire n22125;
    wire n22128;
    wire n22131;
    wire n22134;
    wire n22137;
    wire n22140;
    wire n22143;
    wire n22146;
    wire n22149;
    wire n22152;
    wire n22155;
    wire n22158;
    wire n22161;
    wire n22164;
    wire n22167;
    wire n22170;
    wire n22173;
    wire n22176;
    wire n22179;
    wire n22182;
    wire n22185;
    wire n22188;
    wire n22191;
    wire n22194;
    wire n22197;
    wire n22200;
    wire n22203;
    wire n22206;
    wire n22209;
    wire n22212;
    wire n22215;
    wire n22218;
    wire n22221;
    wire n22224;
    wire n22227;
    wire n22230;
    wire n22233;
    wire n22236;
    wire n22239;
    wire n22242;
    wire n22245;
    wire n22247;
    wire n22251;
    wire n22254;
    wire n22257;
    wire n22260;
    wire n22263;
    wire n22266;
    wire n22269;
    wire n22272;
    wire n22275;
    wire n22278;
    wire n22281;
    wire n22284;
    wire n22287;
    wire n22290;
    wire n22293;
    wire n22296;
    wire n22299;
    wire n22302;
    wire n22305;
    wire n22308;
    wire n22311;
    wire n22314;
    wire n22317;
    wire n22320;
    wire n22323;
    wire n22326;
    wire n22329;
    wire n22332;
    wire n22335;
    wire n22338;
    wire n22341;
    wire n22344;
    wire n22347;
    wire n22350;
    wire n22353;
    wire n22356;
    wire n22359;
    wire n22362;
    wire n22365;
    wire n22368;
    wire n22371;
    wire n22374;
    wire n22377;
    wire n22380;
    wire n22383;
    wire n22386;
    wire n22389;
    wire n22392;
    wire n22395;
    wire n22398;
    wire n22401;
    wire n22404;
    wire n22407;
    wire n22410;
    wire n22413;
    wire n22416;
    wire n22419;
    wire n22422;
    wire n22425;
    wire n22428;
    wire n22431;
    wire n22434;
    wire n22437;
    wire n22440;
    wire n22443;
    wire n22446;
    wire n22449;
    wire n22452;
    wire n22455;
    wire n22458;
    wire n22461;
    wire n22464;
    wire n22467;
    wire n22470;
    wire n22473;
    wire n22476;
    wire n22479;
    wire n22482;
    wire n22485;
    wire n22488;
    wire n22491;
    wire n22494;
    wire n22497;
    wire n22500;
    wire n22503;
    wire n22506;
    wire n22509;
    wire n22512;
    wire n22515;
    wire n22518;
    wire n22521;
    wire n22524;
    wire n22527;
    wire n22530;
    wire n22533;
    wire n22536;
    wire n22539;
    wire n22542;
    wire n22545;
    wire n22548;
    wire n22551;
    wire n22554;
    wire n22557;
    wire n22560;
    wire n22563;
    wire n22566;
    wire n22569;
    wire n22572;
    wire n22575;
    wire n22578;
    wire n22581;
    wire n22584;
    wire n22587;
    wire n22590;
    wire n22593;
    wire n22596;
    wire n22599;
    wire n22602;
    wire n22605;
    wire n22608;
    wire n22611;
    wire n22614;
    wire n22617;
    wire n22620;
    wire n22623;
    wire n22626;
    wire n22629;
    wire n22632;
    wire n22635;
    wire n22638;
    wire n22641;
    wire n22644;
    wire n22647;
    wire n22650;
    wire n22653;
    wire n22656;
    wire n22659;
    wire n22662;
    wire n22665;
    wire n22668;
    wire n22671;
    wire n22674;
    wire n22677;
    wire n22680;
    wire n22683;
    wire n22686;
    wire n22689;
    wire n22692;
    wire n22695;
    wire n22698;
    wire n22701;
    wire n22704;
    wire n22707;
    wire n22710;
    wire n22713;
    wire n22716;
    wire n22719;
    wire n22722;
    wire n22725;
    wire n22728;
    wire n22731;
    wire n22734;
    wire n22737;
    wire n22740;
    wire n22743;
    wire n22746;
    wire n22749;
    wire n22752;
    wire n22755;
    wire n22758;
    wire n22761;
    wire n22764;
    wire n22767;
    wire n22770;
    wire n22773;
    wire n22776;
    wire n22779;
    wire n22782;
    wire n22785;
    wire n22788;
    wire n22791;
    wire n22794;
    wire n22797;
    wire n22800;
    wire n22803;
    wire n22806;
    wire n22809;
    wire n22812;
    wire n22815;
    wire n22818;
    wire n22821;
    wire n22824;
    wire n22827;
    wire n22830;
    wire n22833;
    wire n22836;
    wire n22839;
    wire n22842;
    wire n22845;
    wire n22848;
    wire n22851;
    wire n22854;
    wire n22857;
    wire n22860;
    wire n22863;
    wire n22866;
    wire n22869;
    wire n22872;
    wire n22875;
    wire n22878;
    wire n22881;
    wire n22884;
    wire n22887;
    wire n22890;
    wire n22893;
    wire n22896;
    wire n22899;
    wire n22902;
    wire n22905;
    wire n22908;
    wire n22911;
    wire n22914;
    wire n22917;
    wire n22920;
    wire n22923;
    wire n22926;
    wire n22929;
    wire n22932;
    wire n22935;
    wire n22938;
    wire n22941;
    wire n22944;
    wire n22947;
    wire n22950;
    wire n22953;
    wire n22956;
    wire n22959;
    wire n22962;
    wire n22965;
    wire n22968;
    wire n22971;
    wire n22974;
    wire n22977;
    wire n22980;
    wire n22983;
    wire n22986;
    wire n22989;
    wire n22992;
    wire n22995;
    wire n22998;
    wire n23001;
    wire n23004;
    wire n23007;
    wire n23010;
    wire n23013;
    wire n23016;
    wire n23019;
    wire n23022;
    wire n23025;
    wire n23028;
    wire n23031;
    wire n23034;
    wire n23037;
    wire n23040;
    wire n23043;
    wire n23046;
    wire n23049;
    wire n23052;
    wire n23055;
    wire n23058;
    wire n23061;
    wire n23064;
    wire n23067;
    wire n23070;
    wire n23073;
    wire n23076;
    wire n23079;
    wire n23082;
    wire n23085;
    wire n23088;
    wire n23091;
    wire n23094;
    wire n23097;
    wire n23100;
    wire n23103;
    wire n23106;
    wire n23109;
    wire n23112;
    wire n23115;
    wire n23118;
    wire n23121;
    wire n23124;
    wire n23127;
    wire n23130;
    wire n23133;
    wire n23136;
    wire n23139;
    wire n23142;
    wire n23145;
    wire n23148;
    wire n23151;
    wire n23154;
    wire n23157;
    wire n23160;
    wire n23163;
    wire n23166;
    wire n23169;
    wire n23172;
    wire n23175;
    wire n23178;
    wire n23181;
    wire n23184;
    wire n23187;
    wire n23190;
    wire n23193;
    wire n23196;
    wire n23199;
    wire n23202;
    wire n23205;
    wire n23208;
    wire n23211;
    wire n23214;
    wire n23217;
    wire n23220;
    wire n23223;
    wire n23226;
    wire n23228;
    wire n23231;
    wire n23234;
    wire n23237;
    wire n23241;
    wire n23244;
    wire n23247;
    wire n23250;
    wire n23253;
    wire n23256;
    wire n23259;
    wire n23262;
    wire n23265;
    wire n23268;
    wire n23271;
    wire n23274;
    wire n23277;
    wire n23280;
    wire n23283;
    wire n23286;
    wire n23289;
    wire n23292;
    wire n23295;
    wire n23298;
    wire n23301;
    wire n23304;
    wire n23307;
    wire n23310;
    wire n23313;
    wire n23316;
    wire n23319;
    wire n23322;
    wire n23325;
    wire n23328;
    wire n23331;
    wire n23334;
    wire n23337;
    wire n23340;
    wire n23343;
    wire n23346;
    wire n23349;
    wire n23352;
    wire n23355;
    wire n23358;
    wire n23361;
    wire n23364;
    wire n23367;
    wire n23370;
    wire n23373;
    wire n23376;
    wire n23379;
    wire n23382;
    wire n23385;
    wire n23388;
    wire n23391;
    wire n23394;
    wire n23397;
    wire n23400;
    wire n23403;
    wire n23406;
    wire n23409;
    wire n23412;
    wire n23415;
    wire n23418;
    wire n23421;
    wire n23424;
    wire n23427;
    wire n23430;
    wire n23433;
    wire n23436;
    wire n23439;
    wire n23442;
    wire n23445;
    wire n23448;
    wire n23451;
    wire n23454;
    wire n23457;
    wire n23460;
    wire n23463;
    wire n23466;
    wire n23469;
    wire n23472;
    wire n23475;
    wire n23478;
    wire n23481;
    wire n23484;
    wire n23487;
    wire n23490;
    wire n23493;
    wire n23496;
    wire n23499;
    wire n23502;
    wire n23505;
    wire n23508;
    wire n23511;
    wire n23514;
    wire n23517;
    wire n23520;
    wire n23523;
    wire n23526;
    wire n23529;
    wire n23532;
    wire n23535;
    wire n23538;
    wire n23541;
    wire n23544;
    wire n23547;
    wire n23550;
    wire n23553;
    wire n23556;
    wire n23559;
    wire n23562;
    wire n23565;
    wire n23568;
    wire n23571;
    wire n23574;
    wire n23577;
    wire n23580;
    wire n23583;
    wire n23586;
    wire n23589;
    wire n23592;
    wire n23595;
    wire n23598;
    wire n23601;
    wire n23604;
    wire n23607;
    wire n23610;
    wire n23613;
    wire n23616;
    wire n23619;
    wire n23622;
    wire n23625;
    wire n23628;
    wire n23631;
    wire n23634;
    wire n23637;
    wire n23640;
    wire n23643;
    wire n23646;
    wire n23649;
    wire n23652;
    wire n23655;
    wire n23658;
    wire n23661;
    wire n23664;
    wire n23667;
    wire n23670;
    wire n23673;
    wire n23676;
    wire n23679;
    wire n23682;
    wire n23685;
    wire n23688;
    wire n23691;
    wire n23694;
    wire n23697;
    wire n23700;
    wire n23703;
    wire n23706;
    wire n23709;
    wire n23712;
    wire n23715;
    wire n23718;
    wire n23721;
    wire n23724;
    wire n23727;
    wire n23730;
    wire n23733;
    wire n23736;
    wire n23739;
    wire n23742;
    wire n23745;
    wire n23748;
    wire n23751;
    wire n23754;
    wire n23757;
    wire n23760;
    wire n23763;
    wire n23766;
    wire n23769;
    wire n23772;
    wire n23775;
    wire n23778;
    wire n23781;
    wire n23784;
    wire n23787;
    wire n23790;
    wire n23793;
    wire n23796;
    wire n23799;
    wire n23802;
    wire n23805;
    wire n23808;
    wire n23811;
    wire n23814;
    wire n23817;
    wire n23820;
    wire n23823;
    wire n23826;
    wire n23829;
    wire n23832;
    wire n23835;
    wire n23838;
    wire n23841;
    wire n23844;
    wire n23847;
    wire n23850;
    wire n23853;
    wire n23856;
    wire n23859;
    wire n23862;
    wire n23865;
    wire n23868;
    wire n23871;
    wire n23874;
    wire n23877;
    wire n23880;
    wire n23883;
    wire n23886;
    wire n23889;
    wire n23892;
    wire n23895;
    wire n23898;
    wire n23901;
    wire n23904;
    wire n23907;
    wire n23910;
    wire n23913;
    wire n23916;
    wire n23919;
    wire n23922;
    wire n23925;
    wire n23928;
    wire n23931;
    wire n23934;
    wire n23937;
    wire n23940;
    wire n23943;
    wire n23946;
    wire n23949;
    wire n23952;
    wire n23955;
    wire n23958;
    wire n23961;
    wire n23964;
    wire n23967;
    wire n23970;
    wire n23973;
    wire n23976;
    wire n23979;
    wire n23982;
    wire n23985;
    wire n23988;
    wire n23991;
    wire n23994;
    wire n23997;
    wire n24000;
    wire n24003;
    wire n24006;
    wire n24009;
    wire n24012;
    wire n24015;
    wire n24018;
    wire n24021;
    wire n24024;
    wire n24027;
    wire n24030;
    wire n24033;
    wire n24036;
    wire n24039;
    wire n24042;
    wire n24045;
    wire n24048;
    wire n24051;
    wire n24054;
    wire n24057;
    wire n24060;
    wire n24063;
    wire n24066;
    wire n24069;
    wire n24072;
    wire n24075;
    wire n24078;
    wire n24081;
    wire n24084;
    wire n24087;
    wire n24090;
    wire n24093;
    wire n24096;
    wire n24099;
    wire n24102;
    wire n24105;
    wire n24108;
    wire n24111;
    wire n24114;
    wire n24117;
    wire n24120;
    wire n24123;
    wire n24126;
    wire n24129;
    wire n24132;
    wire n24135;
    wire n24138;
    wire n24141;
    wire n24144;
    wire n24147;
    wire n24150;
    wire n24153;
    wire n24156;
    wire n24159;
    wire n24162;
    wire n24165;
    wire n24168;
    wire n24171;
    wire n24174;
    wire n24177;
    wire n24180;
    wire n24183;
    wire n24186;
    wire n24189;
    wire n24192;
    wire n24195;
    wire n24198;
    wire n24201;
    wire n24204;
    wire n24207;
    wire n24210;
    wire n24213;
    wire n24216;
    wire n24219;
    wire n24222;
    wire n24225;
    wire n24228;
    wire n24231;
    wire n24234;
    wire n24237;
    wire n24240;
    wire n24243;
    wire n24246;
    wire n24249;
    wire n24252;
    wire n24255;
    wire n24258;
    wire n24261;
    wire n24264;
    wire n24267;
    wire n24270;
    wire n24273;
    wire n24276;
    wire n24279;
    wire n24282;
    wire n24285;
    wire n24288;
    wire n24291;
    wire n24294;
    wire n24297;
    wire n24300;
    wire n24303;
    wire n24306;
    wire n24309;
    wire n24312;
    wire n24315;
    wire n24318;
    wire n24321;
    wire n24324;
    wire n24327;
    wire n24330;
    wire n24333;
    wire n24336;
    wire n24339;
    wire n24342;
    wire n24345;
    wire n24348;
    wire n24351;
    wire n24354;
    wire n24357;
    wire n24360;
    wire n24362;
    wire n24365;
    wire n24368;
    wire n24371;
    wire n24375;
    wire n24377;
    wire n24381;
    wire n24384;
    wire n24387;
    wire n24390;
    wire n24393;
    wire n24396;
    wire n24399;
    wire n24402;
    wire n24405;
    wire n24408;
    wire n24411;
    wire n24414;
    wire n24417;
    wire n24420;
    wire n24423;
    wire n24426;
    wire n24429;
    wire n24432;
    wire n24435;
    wire n24438;
    wire n24441;
    wire n24444;
    wire n24447;
    wire n24450;
    wire n24453;
    wire n24456;
    wire n24459;
    wire n24462;
    wire n24465;
    wire n24468;
    wire n24471;
    wire n24474;
    wire n24477;
    wire n24480;
    wire n24483;
    wire n24486;
    wire n24489;
    wire n24492;
    wire n24495;
    wire n24498;
    wire n24501;
    wire n24504;
    wire n24507;
    wire n24510;
    wire n24513;
    wire n24516;
    wire n24519;
    wire n24522;
    wire n24525;
    wire n24528;
    wire n24531;
    wire n24534;
    wire n24537;
    wire n24540;
    wire n24543;
    wire n24546;
    wire n24549;
    wire n24552;
    wire n24555;
    wire n24558;
    wire n24561;
    wire n24564;
    wire n24567;
    wire n24570;
    wire n24573;
    wire n24576;
    wire n24579;
    wire n24582;
    wire n24585;
    wire n24588;
    wire n24591;
    wire n24594;
    wire n24597;
    wire n24600;
    wire n24603;
    wire n24606;
    wire n24609;
    wire n24612;
    wire n24615;
    wire n24618;
    wire n24621;
    wire n24624;
    wire n24627;
    wire n24630;
    wire n24633;
    wire n24636;
    wire n24639;
    wire n24642;
    wire n24645;
    wire n24648;
    wire n24651;
    wire n24654;
    wire n24657;
    wire n24660;
    wire n24663;
    wire n24666;
    wire n24669;
    wire n24672;
    wire n24675;
    wire n24678;
    wire n24681;
    wire n24684;
    wire n24687;
    wire n24690;
    wire n24693;
    wire n24696;
    wire n24699;
    wire n24702;
    wire n24705;
    wire n24708;
    wire n24711;
    wire n24714;
    wire n24717;
    wire n24720;
    wire n24723;
    wire n24726;
    wire n24729;
    wire n24732;
    wire n24735;
    wire n24738;
    wire n24741;
    wire n24744;
    wire n24747;
    wire n24750;
    wire n24753;
    wire n24756;
    wire n24759;
    wire n24762;
    wire n24765;
    wire n24768;
    wire n24771;
    wire n24774;
    wire n24777;
    wire n24780;
    wire n24783;
    wire n24786;
    wire n24789;
    wire n24792;
    wire n24795;
    wire n24798;
    wire n24801;
    wire n24804;
    wire n24807;
    wire n24810;
    wire n24813;
    wire n24816;
    wire n24819;
    wire n24822;
    wire n24825;
    wire n24828;
    wire n24831;
    wire n24834;
    wire n24837;
    wire n24840;
    wire n24843;
    wire n24846;
    wire n24849;
    wire n24852;
    wire n24855;
    wire n24858;
    wire n24861;
    wire n24864;
    wire n24867;
    wire n24870;
    wire n24873;
    wire n24876;
    wire n24879;
    wire n24882;
    wire n24885;
    wire n24888;
    wire n24891;
    wire n24894;
    wire n24897;
    wire n24900;
    wire n24903;
    wire n24906;
    wire n24909;
    wire n24912;
    wire n24915;
    wire n24918;
    wire n24921;
    wire n24924;
    wire n24927;
    wire n24930;
    wire n24933;
    wire n24936;
    wire n24939;
    wire n24942;
    wire n24945;
    wire n24948;
    wire n24951;
    wire n24954;
    wire n24957;
    wire n24960;
    wire n24963;
    wire n24966;
    wire n24969;
    wire n24972;
    wire n24975;
    wire n24978;
    wire n24981;
    wire n24984;
    wire n24987;
    wire n24990;
    wire n24993;
    wire n24996;
    wire n24999;
    wire n25002;
    wire n25005;
    wire n25008;
    wire n25011;
    wire n25014;
    wire n25017;
    wire n25020;
    wire n25023;
    wire n25026;
    wire n25029;
    wire n25032;
    wire n25035;
    wire n25038;
    wire n25041;
    wire n25044;
    wire n25047;
    wire n25050;
    wire n25053;
    wire n25056;
    wire n25059;
    wire n25062;
    wire n25065;
    wire n25068;
    wire n25071;
    wire n25074;
    wire n25077;
    wire n25080;
    wire n25083;
    wire n25086;
    wire n25089;
    wire n25092;
    wire n25095;
    wire n25098;
    wire n25101;
    wire n25104;
    wire n25107;
    wire n25110;
    wire n25113;
    wire n25116;
    wire n25119;
    wire n25122;
    wire n25125;
    wire n25128;
    wire n25131;
    wire n25134;
    wire n25137;
    wire n25140;
    wire n25143;
    wire n25146;
    wire n25149;
    wire n25152;
    wire n25155;
    wire n25158;
    wire n25161;
    wire n25164;
    wire n25167;
    wire n25170;
    wire n25173;
    wire n25176;
    wire n25179;
    wire n25182;
    wire n25185;
    wire n25188;
    wire n25191;
    wire n25194;
    wire n25197;
    wire n25200;
    wire n25203;
    wire n25206;
    wire n25209;
    wire n25212;
    wire n25215;
    wire n25218;
    wire n25221;
    wire n25224;
    wire n25227;
    wire n25230;
    wire n25233;
    wire n25236;
    wire n25239;
    wire n25242;
    wire n25245;
    wire n25248;
    wire n25251;
    wire n25254;
    wire n25257;
    wire n25260;
    wire n25263;
    wire n25266;
    wire n25269;
    wire n25272;
    wire n25275;
    wire n25278;
    wire n25281;
    wire n25284;
    wire n25287;
    wire n25290;
    wire n25293;
    wire n25296;
    wire n25299;
    wire n25302;
    wire n25305;
    wire n25308;
    wire n25311;
    wire n25314;
    wire n25317;
    wire n25320;
    wire n25323;
    wire n25326;
    wire n25329;
    wire n25332;
    wire n25335;
    wire n25338;
    wire n25341;
    wire n25344;
    wire n25347;
    wire n25350;
    wire n25353;
    wire n25356;
    wire n25359;
    wire n25362;
    wire n25365;
    wire n25368;
    wire n25371;
    wire n25374;
    wire n25377;
    wire n25380;
    wire n25383;
    wire n25386;
    wire n25389;
    wire n25392;
    wire n25395;
    wire n25398;
    wire n25401;
    wire n25404;
    wire n25407;
    wire n25410;
    wire n25413;
    wire n25416;
    wire n25419;
    wire n25422;
    wire n25425;
    wire n25428;
    wire n25431;
    wire n25434;
    wire n25437;
    wire n25440;
    wire n25443;
    wire n25446;
    wire n25449;
    wire n25452;
    wire n25455;
    wire n25458;
    wire n25461;
    wire n25464;
    wire n25467;
    wire n25470;
    wire n25473;
    wire n25476;
    wire n25479;
    wire n25482;
    wire n25485;
    wire n25488;
    wire n25491;
    wire n25494;
    wire n25497;
    wire n25500;
    wire n25502;
    wire n25505;
    wire n25508;
    wire n25511;
    wire n25515;
    wire n25517;
    wire n25521;
    wire n25524;
    wire n25527;
    wire n25530;
    wire n25533;
    wire n25536;
    wire n25539;
    wire n25542;
    wire n25545;
    wire n25548;
    wire n25551;
    wire n25554;
    wire n25557;
    wire n25560;
    wire n25563;
    wire n25566;
    wire n25569;
    wire n25572;
    wire n25575;
    wire n25578;
    wire n25581;
    wire n25584;
    wire n25587;
    wire n25590;
    wire n25593;
    wire n25596;
    wire n25599;
    wire n25602;
    wire n25605;
    wire n25608;
    wire n25611;
    wire n25614;
    wire n25617;
    wire n25620;
    wire n25623;
    wire n25626;
    wire n25629;
    wire n25632;
    wire n25635;
    wire n25638;
    wire n25641;
    wire n25644;
    wire n25647;
    wire n25650;
    wire n25653;
    wire n25656;
    wire n25659;
    wire n25662;
    wire n25665;
    wire n25668;
    wire n25671;
    wire n25674;
    wire n25677;
    wire n25680;
    wire n25683;
    wire n25686;
    wire n25689;
    wire n25692;
    wire n25695;
    wire n25698;
    wire n25701;
    wire n25704;
    wire n25707;
    wire n25710;
    wire n25713;
    wire n25716;
    wire n25719;
    wire n25722;
    wire n25725;
    wire n25728;
    wire n25731;
    wire n25734;
    wire n25737;
    wire n25740;
    wire n25743;
    wire n25746;
    wire n25749;
    wire n25752;
    wire n25755;
    wire n25758;
    wire n25761;
    wire n25764;
    wire n25767;
    wire n25770;
    wire n25773;
    wire n25776;
    wire n25779;
    wire n25782;
    wire n25785;
    wire n25788;
    wire n25791;
    wire n25794;
    wire n25797;
    wire n25800;
    wire n25803;
    wire n25806;
    wire n25809;
    wire n25812;
    wire n25815;
    wire n25818;
    wire n25821;
    wire n25824;
    wire n25827;
    wire n25830;
    wire n25833;
    wire n25836;
    wire n25839;
    wire n25842;
    wire n25845;
    wire n25848;
    wire n25851;
    wire n25854;
    wire n25857;
    wire n25860;
    wire n25863;
    wire n25866;
    wire n25869;
    wire n25872;
    wire n25875;
    wire n25878;
    wire n25881;
    wire n25884;
    wire n25887;
    wire n25890;
    wire n25893;
    wire n25896;
    wire n25899;
    wire n25902;
    wire n25905;
    wire n25908;
    wire n25911;
    wire n25914;
    wire n25917;
    wire n25920;
    wire n25923;
    wire n25926;
    wire n25929;
    wire n25932;
    wire n25935;
    wire n25938;
    wire n25941;
    wire n25944;
    wire n25947;
    wire n25950;
    wire n25953;
    wire n25956;
    wire n25959;
    wire n25962;
    wire n25965;
    wire n25968;
    wire n25971;
    wire n25974;
    wire n25977;
    wire n25980;
    wire n25983;
    wire n25986;
    wire n25989;
    wire n25992;
    wire n25995;
    wire n25998;
    wire n26001;
    wire n26004;
    wire n26007;
    wire n26010;
    wire n26013;
    wire n26016;
    wire n26019;
    wire n26022;
    wire n26025;
    wire n26028;
    wire n26031;
    wire n26034;
    wire n26037;
    wire n26040;
    wire n26043;
    wire n26046;
    wire n26049;
    wire n26052;
    wire n26055;
    wire n26058;
    wire n26061;
    wire n26064;
    wire n26067;
    wire n26070;
    wire n26073;
    wire n26076;
    wire n26079;
    wire n26082;
    wire n26085;
    wire n26088;
    wire n26091;
    wire n26094;
    wire n26097;
    wire n26100;
    wire n26103;
    wire n26106;
    wire n26109;
    wire n26112;
    wire n26115;
    wire n26118;
    wire n26121;
    wire n26124;
    wire n26127;
    wire n26130;
    wire n26133;
    wire n26136;
    wire n26139;
    wire n26142;
    wire n26145;
    wire n26148;
    wire n26151;
    wire n26154;
    wire n26157;
    wire n26160;
    wire n26163;
    wire n26166;
    wire n26169;
    wire n26172;
    wire n26175;
    wire n26178;
    wire n26181;
    wire n26184;
    wire n26187;
    wire n26190;
    wire n26193;
    wire n26196;
    wire n26199;
    wire n26202;
    wire n26205;
    wire n26208;
    wire n26211;
    wire n26214;
    wire n26217;
    wire n26220;
    wire n26223;
    wire n26226;
    wire n26229;
    wire n26232;
    wire n26235;
    wire n26238;
    wire n26241;
    wire n26244;
    wire n26247;
    wire n26250;
    wire n26253;
    wire n26256;
    wire n26259;
    wire n26262;
    wire n26265;
    wire n26268;
    wire n26271;
    wire n26274;
    wire n26277;
    wire n26280;
    wire n26283;
    wire n26286;
    wire n26289;
    wire n26292;
    wire n26295;
    wire n26298;
    wire n26301;
    wire n26304;
    wire n26307;
    wire n26310;
    wire n26313;
    wire n26316;
    wire n26319;
    wire n26322;
    wire n26325;
    wire n26328;
    wire n26331;
    wire n26334;
    wire n26337;
    wire n26340;
    wire n26343;
    wire n26346;
    wire n26349;
    wire n26352;
    wire n26355;
    wire n26358;
    wire n26361;
    wire n26364;
    wire n26367;
    wire n26370;
    wire n26373;
    wire n26376;
    wire n26379;
    wire n26382;
    wire n26385;
    wire n26388;
    wire n26391;
    wire n26394;
    wire n26397;
    wire n26400;
    wire n26403;
    wire n26406;
    wire n26409;
    wire n26412;
    wire n26415;
    wire n26418;
    wire n26421;
    wire n26424;
    wire n26427;
    wire n26430;
    wire n26433;
    wire n26436;
    wire n26439;
    wire n26442;
    wire n26445;
    wire n26448;
    wire n26451;
    wire n26454;
    wire n26457;
    wire n26460;
    wire n26463;
    wire n26466;
    wire n26469;
    wire n26472;
    wire n26475;
    wire n26478;
    wire n26481;
    wire n26484;
    wire n26487;
    wire n26490;
    wire n26493;
    wire n26496;
    wire n26499;
    wire n26502;
    wire n26505;
    wire n26508;
    wire n26511;
    wire n26514;
    wire n26517;
    wire n26520;
    wire n26523;
    wire n26526;
    wire n26529;
    wire n26532;
    wire n26535;
    wire n26538;
    wire n26541;
    wire n26544;
    wire n26547;
    wire n26550;
    wire n26553;
    wire n26556;
    wire n26559;
    wire n26562;
    wire n26565;
    wire n26568;
    wire n26571;
    wire n26574;
    wire n26577;
    wire n26580;
    wire n26583;
    wire n26586;
    wire n26589;
    wire n26592;
    wire n26595;
    wire n26598;
    wire n26601;
    wire n26604;
    wire n26607;
    wire n26610;
    wire n26613;
    wire n26616;
    wire n26619;
    wire n26622;
    wire n26625;
    wire n26628;
    wire n26631;
    wire n26634;
    wire n26637;
    wire n26640;
    wire n26643;
    wire n26646;
    wire n26649;
    wire n26652;
    wire n26655;
    wire n26658;
    wire n26661;
    wire n26663;
    wire n26666;
    wire n26669;
    wire n26672;
    wire n26676;
    wire n26678;
    wire n26682;
    wire n26685;
    wire n26688;
    wire n26691;
    wire n26694;
    wire n26697;
    wire n26700;
    wire n26703;
    wire n26706;
    wire n26709;
    wire n26712;
    wire n26715;
    wire n26718;
    wire n26721;
    wire n26724;
    wire n26727;
    wire n26730;
    wire n26733;
    wire n26736;
    wire n26739;
    wire n26742;
    wire n26745;
    wire n26748;
    wire n26751;
    wire n26754;
    wire n26757;
    wire n26760;
    wire n26763;
    wire n26766;
    wire n26769;
    wire n26772;
    wire n26775;
    wire n26778;
    wire n26781;
    wire n26784;
    wire n26787;
    wire n26790;
    wire n26793;
    wire n26796;
    wire n26799;
    wire n26802;
    wire n26805;
    wire n26808;
    wire n26811;
    wire n26814;
    wire n26817;
    wire n26820;
    wire n26823;
    wire n26826;
    wire n26829;
    wire n26832;
    wire n26835;
    wire n26838;
    wire n26841;
    wire n26844;
    wire n26847;
    wire n26850;
    wire n26853;
    wire n26856;
    wire n26859;
    wire n26862;
    wire n26865;
    wire n26868;
    wire n26871;
    wire n26874;
    wire n26877;
    wire n26880;
    wire n26883;
    wire n26886;
    wire n26889;
    wire n26892;
    wire n26895;
    wire n26898;
    wire n26901;
    wire n26904;
    wire n26907;
    wire n26910;
    wire n26913;
    wire n26916;
    wire n26919;
    wire n26922;
    wire n26925;
    wire n26928;
    wire n26931;
    wire n26934;
    wire n26937;
    wire n26940;
    wire n26943;
    wire n26946;
    wire n26949;
    wire n26952;
    wire n26955;
    wire n26958;
    wire n26961;
    wire n26964;
    wire n26967;
    wire n26970;
    wire n26973;
    wire n26976;
    wire n26979;
    wire n26982;
    wire n26985;
    wire n26988;
    wire n26991;
    wire n26994;
    wire n26997;
    wire n27000;
    wire n27003;
    wire n27006;
    wire n27009;
    wire n27012;
    wire n27015;
    wire n27018;
    wire n27021;
    wire n27024;
    wire n27027;
    wire n27030;
    wire n27033;
    wire n27036;
    wire n27039;
    wire n27042;
    wire n27045;
    wire n27048;
    wire n27051;
    wire n27054;
    wire n27057;
    wire n27060;
    wire n27063;
    wire n27066;
    wire n27069;
    wire n27072;
    wire n27075;
    wire n27078;
    wire n27081;
    wire n27084;
    wire n27087;
    wire n27090;
    wire n27093;
    wire n27096;
    wire n27099;
    wire n27102;
    wire n27105;
    wire n27108;
    wire n27111;
    wire n27114;
    wire n27117;
    wire n27120;
    wire n27123;
    wire n27126;
    wire n27129;
    wire n27132;
    wire n27135;
    wire n27138;
    wire n27141;
    wire n27144;
    wire n27147;
    wire n27150;
    wire n27153;
    wire n27156;
    wire n27159;
    wire n27162;
    wire n27165;
    wire n27168;
    wire n27171;
    wire n27174;
    wire n27177;
    wire n27180;
    wire n27183;
    wire n27186;
    wire n27189;
    wire n27192;
    wire n27195;
    wire n27198;
    wire n27201;
    wire n27204;
    wire n27207;
    wire n27210;
    wire n27213;
    wire n27216;
    wire n27219;
    wire n27222;
    wire n27225;
    wire n27228;
    wire n27231;
    wire n27234;
    wire n27237;
    wire n27240;
    wire n27243;
    wire n27246;
    wire n27249;
    wire n27252;
    wire n27255;
    wire n27258;
    wire n27261;
    wire n27264;
    wire n27267;
    wire n27270;
    wire n27273;
    wire n27276;
    wire n27279;
    wire n27282;
    wire n27285;
    wire n27288;
    wire n27291;
    wire n27294;
    wire n27297;
    wire n27300;
    wire n27303;
    wire n27306;
    wire n27309;
    wire n27312;
    wire n27315;
    wire n27318;
    wire n27321;
    wire n27324;
    wire n27327;
    wire n27330;
    wire n27333;
    wire n27336;
    wire n27339;
    wire n27342;
    wire n27345;
    wire n27348;
    wire n27351;
    wire n27354;
    wire n27357;
    wire n27360;
    wire n27363;
    wire n27366;
    wire n27369;
    wire n27372;
    wire n27375;
    wire n27378;
    wire n27381;
    wire n27384;
    wire n27387;
    wire n27390;
    wire n27393;
    wire n27396;
    wire n27399;
    wire n27402;
    wire n27405;
    wire n27408;
    wire n27411;
    wire n27414;
    wire n27417;
    wire n27420;
    wire n27423;
    wire n27426;
    wire n27429;
    wire n27432;
    wire n27435;
    wire n27438;
    wire n27441;
    wire n27444;
    wire n27447;
    wire n27450;
    wire n27453;
    wire n27456;
    wire n27459;
    wire n27462;
    wire n27465;
    wire n27468;
    wire n27471;
    wire n27474;
    wire n27477;
    wire n27480;
    wire n27483;
    wire n27486;
    wire n27489;
    wire n27492;
    wire n27495;
    wire n27498;
    wire n27501;
    wire n27504;
    wire n27507;
    wire n27510;
    wire n27513;
    wire n27516;
    wire n27519;
    wire n27522;
    wire n27525;
    wire n27528;
    wire n27531;
    wire n27534;
    wire n27537;
    wire n27540;
    wire n27543;
    wire n27546;
    wire n27549;
    wire n27552;
    wire n27555;
    wire n27558;
    wire n27561;
    wire n27564;
    wire n27567;
    wire n27570;
    wire n27573;
    wire n27576;
    wire n27579;
    wire n27582;
    wire n27585;
    wire n27588;
    wire n27591;
    wire n27594;
    wire n27597;
    wire n27600;
    wire n27603;
    wire n27606;
    wire n27609;
    wire n27612;
    wire n27615;
    wire n27618;
    wire n27621;
    wire n27624;
    wire n27627;
    wire n27630;
    wire n27633;
    wire n27636;
    wire n27639;
    wire n27642;
    wire n27645;
    wire n27648;
    wire n27651;
    wire n27654;
    wire n27657;
    wire n27660;
    wire n27663;
    wire n27666;
    wire n27669;
    wire n27672;
    wire n27675;
    wire n27678;
    wire n27681;
    wire n27684;
    wire n27687;
    wire n27690;
    wire n27693;
    wire n27696;
    wire n27699;
    wire n27702;
    wire n27705;
    wire n27708;
    wire n27711;
    wire n27714;
    wire n27717;
    wire n27720;
    wire n27723;
    wire n27726;
    wire n27729;
    wire n27732;
    wire n27735;
    wire n27738;
    wire n27741;
    wire n27744;
    wire n27747;
    wire n27750;
    wire n27753;
    wire n27756;
    wire n27759;
    wire n27762;
    wire n27765;
    wire n27768;
    wire n27771;
    wire n27774;
    wire n27777;
    wire n27780;
    wire n27783;
    wire n27786;
    wire n27789;
    wire n27792;
    wire n27795;
    wire n27798;
    wire n27801;
    wire n27804;
    wire n27807;
    wire n27810;
    wire n27813;
    wire n27816;
    wire n27819;
    wire n27822;
    wire n27825;
    wire n27828;
    wire n27831;
    wire n27834;
    wire n27837;
    wire n27840;
    wire n27843;
    wire n27846;
    wire n27849;
    wire n27852;
    wire n27855;
    wire n27857;
    wire n27860;
    wire n27863;
    wire n27866;
    wire n27870;
    wire n27873;
    wire n27876;
    wire n27879;
    wire n27882;
    wire n27885;
    wire n27888;
    wire n27891;
    wire n27894;
    wire n27897;
    wire n27900;
    wire n27903;
    wire n27906;
    wire n27909;
    wire n27912;
    wire n27915;
    wire n27918;
    wire n27921;
    wire n27924;
    wire n27927;
    wire n27930;
    wire n27933;
    wire n27936;
    wire n27939;
    wire n27942;
    wire n27945;
    wire n27948;
    wire n27951;
    wire n27954;
    wire n27957;
    wire n27960;
    wire n27963;
    wire n27966;
    wire n27969;
    wire n27972;
    wire n27975;
    wire n27978;
    wire n27981;
    wire n27984;
    wire n27987;
    wire n27990;
    wire n27993;
    wire n27996;
    wire n27999;
    wire n28002;
    wire n28005;
    wire n28008;
    wire n28011;
    wire n28014;
    wire n28017;
    wire n28020;
    wire n28023;
    wire n28026;
    wire n28029;
    wire n28032;
    wire n28035;
    wire n28038;
    wire n28041;
    wire n28044;
    wire n28047;
    wire n28050;
    wire n28053;
    wire n28056;
    wire n28059;
    wire n28062;
    wire n28065;
    wire n28068;
    wire n28071;
    wire n28074;
    wire n28077;
    wire n28080;
    wire n28083;
    wire n28086;
    wire n28089;
    wire n28092;
    wire n28095;
    wire n28098;
    wire n28101;
    wire n28104;
    wire n28107;
    wire n28110;
    wire n28113;
    wire n28116;
    wire n28119;
    wire n28122;
    wire n28125;
    wire n28128;
    wire n28131;
    wire n28134;
    wire n28137;
    wire n28140;
    wire n28143;
    wire n28146;
    wire n28149;
    wire n28152;
    wire n28155;
    wire n28158;
    wire n28161;
    wire n28164;
    wire n28167;
    wire n28170;
    wire n28173;
    wire n28176;
    wire n28179;
    wire n28182;
    wire n28185;
    wire n28188;
    wire n28191;
    wire n28194;
    wire n28197;
    wire n28200;
    wire n28202;
    wire n28206;
    wire n28209;
    wire n28212;
    wire n28215;
    wire n28218;
    wire n28221;
    wire n28224;
    wire n28227;
    wire n28230;
    wire n28233;
    wire n28236;
    wire n28239;
    wire n28242;
    wire n28245;
    wire n28248;
    wire n28251;
    wire n28254;
    wire n28257;
    wire n28260;
    wire n28263;
    wire n28266;
    wire n28269;
    wire n28272;
    wire n28275;
    wire n28278;
    wire n28281;
    wire n28284;
    wire n28287;
    wire n28290;
    wire n28293;
    wire n28296;
    wire n28299;
    wire n28302;
    wire n28305;
    wire n28308;
    wire n28311;
    wire n28314;
    wire n28317;
    wire n28320;
    wire n28323;
    wire n28326;
    wire n28329;
    wire n28332;
    wire n28335;
    wire n28338;
    wire n28341;
    wire n28344;
    wire n28347;
    wire n28350;
    wire n28353;
    wire n28356;
    wire n28359;
    wire n28362;
    wire n28365;
    wire n28368;
    wire n28371;
    wire n28374;
    wire n28377;
    wire n28380;
    wire n28383;
    wire n28386;
    wire n28389;
    wire n28392;
    wire n28395;
    wire n28398;
    wire n28401;
    wire n28404;
    wire n28407;
    wire n28410;
    wire n28413;
    wire n28416;
    wire n28419;
    wire n28422;
    wire n28425;
    wire n28428;
    wire n28431;
    wire n28434;
    wire n28437;
    wire n28440;
    wire n28443;
    wire n28446;
    wire n28449;
    wire n28452;
    wire n28455;
    wire n28458;
    wire n28461;
    wire n28464;
    wire n28467;
    wire n28470;
    wire n28473;
    wire n28476;
    wire n28479;
    wire n28482;
    wire n28485;
    wire n28488;
    wire n28491;
    wire n28494;
    wire n28497;
    wire n28500;
    wire n28503;
    wire n28506;
    wire n28509;
    wire n28512;
    wire n28515;
    wire n28518;
    wire n28521;
    wire n28524;
    wire n28527;
    wire n28530;
    wire n28533;
    wire n28536;
    wire n28539;
    wire n28542;
    wire n28545;
    wire n28548;
    wire n28551;
    wire n28554;
    wire n28557;
    wire n28560;
    wire n28563;
    wire n28566;
    wire n28569;
    wire n28572;
    wire n28575;
    wire n28578;
    wire n28581;
    wire n28584;
    wire n28587;
    wire n28590;
    wire n28593;
    wire n28596;
    wire n28599;
    wire n28602;
    wire n28605;
    wire n28608;
    wire n28611;
    wire n28614;
    wire n28617;
    wire n28620;
    wire n28623;
    wire n28626;
    wire n28629;
    wire n28632;
    wire n28635;
    wire n28638;
    wire n28641;
    wire n28644;
    wire n28647;
    wire n28650;
    wire n28653;
    wire n28656;
    wire n28659;
    wire n28662;
    wire n28665;
    wire n28668;
    wire n28671;
    wire n28674;
    wire n28677;
    wire n28680;
    wire n28683;
    wire n28686;
    wire n28689;
    wire n28692;
    wire n28695;
    wire n28698;
    wire n28701;
    wire n28704;
    wire n28707;
    wire n28710;
    wire n28713;
    wire n28716;
    wire n28719;
    wire n28722;
    wire n28725;
    wire n28728;
    wire n28731;
    wire n28734;
    wire n28737;
    wire n28740;
    wire n28743;
    wire n28746;
    wire n28749;
    wire n28752;
    wire n28755;
    wire n28758;
    wire n28761;
    wire n28764;
    wire n28767;
    wire n28770;
    wire n28773;
    wire n28776;
    wire n28779;
    wire n28782;
    wire n28785;
    wire n28788;
    wire n28791;
    wire n28794;
    wire n28797;
    wire n28800;
    wire n28803;
    wire n28806;
    wire n28809;
    wire n28812;
    wire n28815;
    wire n28818;
    wire n28821;
    wire n28824;
    wire n28827;
    wire n28830;
    wire n28833;
    wire n28836;
    wire n28839;
    wire n28842;
    wire n28845;
    wire n28848;
    wire n28851;
    wire n28854;
    wire n28857;
    wire n28860;
    wire n28863;
    wire n28866;
    wire n28869;
    wire n28872;
    wire n28875;
    wire n28878;
    wire n28881;
    wire n28884;
    wire n28887;
    wire n28890;
    wire n28893;
    wire n28896;
    wire n28899;
    wire n28902;
    wire n28905;
    wire n28908;
    wire n28911;
    wire n28914;
    wire n28917;
    wire n28920;
    wire n28923;
    wire n28926;
    wire n28929;
    wire n28932;
    wire n28935;
    wire n28938;
    wire n28941;
    wire n28944;
    wire n28947;
    wire n28950;
    wire n28953;
    wire n28956;
    wire n28959;
    wire n28962;
    wire n28965;
    wire n28968;
    wire n28971;
    wire n28974;
    wire n28977;
    wire n28980;
    wire n28983;
    wire n28986;
    wire n28989;
    wire n28992;
    wire n28995;
    wire n28998;
    wire n29001;
    wire n29004;
    wire n29007;
    wire n29010;
    wire n29013;
    wire n29016;
    wire n29019;
    wire n29022;
    wire n29025;
    wire n29028;
    wire n29031;
    wire n29034;
    wire n29037;
    wire n29040;
    wire n29043;
    wire n29046;
    wire n29049;
    wire n29052;
    wire n29055;
    wire n29058;
    wire n29061;
    wire n29064;
    wire n29067;
    wire n29070;
    wire n29073;
    wire n29076;
    wire n29079;
    wire n29082;
    wire n29085;
    wire n29088;
    wire n29091;
    wire n29094;
    wire n29097;
    wire n29100;
    wire n29103;
    wire n29106;
    wire n29109;
    wire n29112;
    wire n29115;
    wire n29118;
    wire n29121;
    wire n29124;
    wire n29127;
    wire n29130;
    wire n29133;
    wire n29136;
    wire n29139;
    wire n29142;
    wire n29145;
    wire n29148;
    wire n29151;
    wire n29154;
    wire n29157;
    wire n29160;
    wire n29163;
    wire n29166;
    wire n29169;
    wire n29172;
    wire n29175;
    wire n29178;
    wire n29181;
    wire n29184;
    wire n29187;
    wire n29190;
    wire n29193;
    wire n29196;
    wire n29199;
    wire n29202;
    wire n29205;
    wire n29208;
    wire n29211;
    wire n29214;
    wire n29217;
    wire n29220;
    wire n29223;
    wire n29226;
    wire n29229;
    wire n29232;
    wire n29235;
    wire n29238;
    wire n29241;
    wire n29244;
    wire n29247;
    wire n29250;
    wire n29253;
    wire n29256;
    wire n29259;
    wire n29262;
    wire n29265;
    wire n29268;
    wire n29271;
    wire n29274;
    wire n29277;
    wire n29280;
    wire n29283;
    wire n29286;
    wire n29289;
    wire n29292;
    wire n29295;
    wire n29298;
    wire n29301;
    wire n29304;
    wire n29307;
    wire n29310;
    wire n29313;
    wire n29316;
    wire n29319;
    wire n29322;
    wire n29325;
    wire n29328;
    wire n29331;
    wire n29334;
    wire n29337;
    wire n29340;
    wire n29343;
    wire n29346;
    wire n29349;
    wire n29352;
    wire n29355;
    wire n29358;
    wire n29361;
    wire n29364;
    wire n29367;
    wire n29370;
    wire n29373;
    wire n29376;
    wire n29379;
    wire n29382;
    wire n29385;
    wire n29388;
    wire n29391;
    wire n29394;
    wire n29397;
    wire n29400;
    wire n29403;
    wire n29406;
    wire n29409;
    wire n29412;
    wire n29415;
    wire n29418;
    wire n29421;
    wire n29424;
    wire n29427;
    wire n29430;
    wire n29433;
    wire n29436;
    wire n29439;
    wire n29442;
    wire n29445;
    wire n29448;
    wire n29451;
    wire n29454;
    wire n29457;
    wire n29460;
    wire n29463;
    wire n29466;
    wire n29469;
    wire n29472;
    wire n29475;
    wire n29478;
    wire n29481;
    wire n29484;
    wire n29487;
    wire n29490;
    wire n29493;
    wire n29496;
    wire n29499;
    wire n29502;
    wire n29505;
    wire n29508;
    wire n29511;
    wire n29514;
    wire n29517;
    wire n29520;
    wire n29523;
    wire n29526;
    wire n29529;
    wire n29532;
    wire n29535;
    wire n29538;
    wire n29541;
    wire n29544;
    wire n29547;
    wire n29550;
    wire n29553;
    wire n29556;
    wire n29559;
    wire n29562;
    wire n29565;
    wire n29568;
    wire n29571;
    wire n29574;
    wire n29577;
    wire n29580;
    wire n29583;
    wire n29586;
    wire n29589;
    wire n29592;
    wire n29595;
    wire n29598;
    wire n29601;
    wire n29604;
    wire n29607;
    wire n29610;
    wire n29613;
    wire n29616;
    wire n29619;
    wire n29622;
    wire n29625;
    wire n29628;
    wire n29631;
    wire n29634;
    wire n29637;
    wire n29640;
    wire n29643;
    wire n29646;
    wire n29649;
    wire n29652;
    wire n29655;
    wire n29658;
    wire n29661;
    wire n29664;
    wire n29667;
    wire n29670;
    wire n29673;
    wire n29676;
    wire n29679;
    wire n29682;
    wire n29685;
    wire n29688;
    wire n29691;
    wire n29694;
    wire n29697;
    wire n29700;
    wire n29703;
    wire n29706;
    wire n29709;
    wire n29712;
    wire n29715;
    wire n29718;
    wire n29721;
    wire n29724;
    wire n29727;
    wire n29730;
    wire n29733;
    wire n29736;
    wire n29739;
    wire n29742;
    wire n29745;
    wire n29748;
    wire n29751;
    wire n29754;
    wire n29757;
    wire n29760;
    wire n29763;
    wire n29766;
    wire n29769;
    wire n29772;
    wire n29775;
    wire n29778;
    wire n29781;
    wire n29784;
    wire n29787;
    wire n29790;
    wire n29793;
    wire n29796;
    wire n29799;
    wire n29802;
    wire n29805;
    wire n29808;
    wire n29811;
    wire n29814;
    wire n29817;
    wire n29820;
    wire n29823;
    wire n29826;
    wire n29829;
    wire n29832;
    wire n29835;
    wire n29838;
    wire n29841;
    wire n29844;
    wire n29847;
    wire n29850;
    wire n29853;
    wire n29856;
    wire n29859;
    wire n29862;
    wire n29865;
    wire n29868;
    wire n29871;
    wire n29874;
    wire n29877;
    wire n29880;
    wire n29883;
    wire n29886;
    wire n29889;
    wire n29892;
    wire n29895;
    wire n29898;
    wire n29901;
    wire n29904;
    wire n29907;
    wire n29910;
    wire n29913;
    wire n29916;
    wire n29919;
    wire n29922;
    wire n29925;
    wire n29928;
    wire n29931;
    wire n29934;
    wire n29937;
    wire n29940;
    wire n29943;
    wire n29946;
    wire n29949;
    wire n29952;
    wire n29955;
    wire n29958;
    wire n29961;
    wire n29964;
    wire n29967;
    wire n29970;
    wire n29973;
    wire n29976;
    wire n29979;
    wire n29982;
    wire n29985;
    wire n29988;
    wire n29991;
    wire n29994;
    wire n29997;
    wire n30000;
    wire n30003;
    wire n30006;
    wire n30009;
    wire n30012;
    wire n30015;
    wire n30018;
    wire n30021;
    wire n30024;
    wire n30027;
    wire n30030;
    wire n30033;
    wire n30036;
    wire n30039;
    wire n30042;
    wire n30045;
    wire n30048;
    wire n30051;
    wire n30054;
    wire n30057;
    wire n30060;
    wire n30063;
    wire n30066;
    wire n30069;
    wire n30072;
    wire n30075;
    wire n30078;
    wire n30081;
    wire n30084;
    wire n30087;
    wire n30090;
    wire n30093;
    wire n30096;
    wire n30099;
    wire n30102;
    wire n30105;
    wire n30108;
    wire n30111;
    wire n30114;
    wire n30117;
    wire n30120;
    wire n30123;
    wire n30126;
    wire n30129;
    wire n30132;
    wire n30135;
    wire n30138;
    wire n30141;
    wire n30144;
    wire n30147;
    wire n30150;
    wire n30153;
    wire n30156;
    wire n30159;
    wire n30162;
    wire n30165;
    wire n30168;
    wire n30171;
    wire n30174;
    wire n30177;
    wire n30180;
    wire n30183;
    wire n30186;
    wire n30189;
    wire n30192;
    wire n30195;
    wire n30198;
    wire n30201;
    wire n30204;
    wire n30207;
    wire n30210;
    wire n30213;
    wire n30216;
    wire n30219;
    wire n30222;
    wire n30225;
    wire n30228;
    wire n30231;
    wire n30234;
    wire n30237;
    wire n30240;
    wire n30243;
    wire n30246;
    wire n30249;
    wire n30252;
    wire n30255;
    wire n30258;
    wire n30261;
    wire n30264;
    wire n30267;
    wire n30270;
    wire n30273;
    wire n30276;
    wire n30279;
    wire n30282;
    wire n30285;
    wire n30288;
    wire n30291;
    wire n30294;
    wire n30297;
    wire n30300;
    wire n30303;
    wire n30306;
    wire n30309;
    wire n30312;
    wire n30315;
    wire n30318;
    wire n30321;
    wire n30324;
    wire n30327;
    wire n30330;
    wire n30333;
    wire n30336;
    wire n30339;
    wire n30342;
    wire n30345;
    wire n30348;
    wire n30351;
    wire n30354;
    wire n30357;
    wire n30360;
    wire n30363;
    wire n30366;
    wire n30369;
    wire n30372;
    wire n30375;
    wire n30378;
    wire n30381;
    wire n30384;
    wire n30387;
    wire n30390;
    wire n30393;
    wire n30396;
    wire n30399;
    wire n30402;
    wire n30405;
    wire n30408;
    wire n30411;
    wire n30414;
    wire n30417;
    wire n30420;
    wire n30423;
    wire n30426;
    wire n30429;
    wire n30432;
    wire n30435;
    wire n30438;
    wire n30441;
    wire n30444;
    wire n30447;
    wire n30450;
    wire n30453;
    wire n30456;
    wire n30459;
    wire n30462;
    wire n30465;
    wire n30468;
    wire n30471;
    wire n30474;
    wire n30477;
    wire n30480;
    wire n30483;
    wire n30486;
    wire n30489;
    wire n30492;
    wire n30495;
    wire n30498;
    wire n30501;
    wire n30504;
    wire n30507;
    wire n30510;
    wire n30513;
    wire n30516;
    wire n30519;
    wire n30522;
    wire n30525;
    wire n30528;
    wire n30531;
    wire n30534;
    wire n30537;
    wire n30540;
    wire n30543;
    wire n30546;
    wire n30549;
    wire n30552;
    wire n30555;
    wire n30558;
    wire n30561;
    wire n30564;
    wire n30567;
    wire n30570;
    wire n30573;
    wire n30576;
    wire n30579;
    wire n30582;
    wire n30585;
    wire n30588;
    wire n30591;
    wire n30594;
    wire n30597;
    wire n30600;
    wire n30603;
    wire n30606;
    wire n30609;
    wire n30612;
    wire n30615;
    wire n30618;
    wire n30621;
    wire n30624;
    wire n30627;
    wire n30630;
    wire n30633;
    wire n30636;
    wire n30639;
    wire n30642;
    wire n30645;
    wire n30648;
    wire n30651;
    wire n30654;
    wire n30657;
    wire n30660;
    wire n30663;
    wire n30666;
    wire n30669;
    wire n30672;
    wire n30675;
    wire n30678;
    wire n30681;
    wire n30684;
    wire n30687;
    wire n30690;
    wire n30693;
    wire n30696;
    wire n30699;
    wire n30702;
    wire n30705;
    wire n30708;
    wire n30711;
    wire n30714;
    wire n30717;
    wire n30720;
    wire n30723;
    wire n30726;
    wire n30729;
    wire n30732;
    wire n30735;
    wire n30738;
    wire n30741;
    wire n30744;
    wire n30747;
    wire n30750;
    wire n30753;
    wire n30756;
    wire n30759;
    wire n30762;
    wire n30765;
    wire n30768;
    wire n30771;
    wire n30774;
    wire n30777;
    wire n30780;
    wire n30783;
    wire n30786;
    wire n30789;
    wire n30792;
    wire n30795;
    wire n30798;
    wire n30801;
    wire n30804;
    wire n30807;
    wire n30810;
    wire n30813;
    wire n30816;
    wire n30819;
    wire n30822;
    wire n30825;
    wire n30828;
    wire n30831;
    wire n30834;
    wire n30837;
    wire n30840;
    wire n30843;
    wire n30846;
    wire n30849;
    wire n30852;
    wire n30855;
    wire n30858;
    wire n30861;
    wire n30864;
    wire n30867;
    wire n30870;
    wire n30873;
    wire n30876;
    wire n30879;
    wire n30882;
    wire n30885;
    wire n30888;
    wire n30891;
    wire n30894;
    wire n30897;
    wire n30900;
    wire n30903;
    wire n30906;
    wire n30909;
    wire n30912;
    wire n30915;
    wire n30918;
    wire n30921;
    wire n30924;
    wire n30927;
    wire n30930;
    wire n30933;
    wire n30936;
    wire n30939;
    wire n30942;
    wire n30945;
    wire n30948;
    wire n30951;
    wire n30954;
    wire n30957;
    wire n30960;
    wire n30963;
    wire n30966;
    wire n30969;
    wire n30972;
    wire n30975;
    wire n30978;
    wire n30981;
    wire n30984;
    wire n30987;
    wire n30990;
    wire n30993;
    wire n30996;
    wire n30999;
    wire n31002;
    wire n31005;
    wire n31008;
    wire n31011;
    wire n31014;
    wire n31017;
    wire n31020;
    wire n31023;
    wire n31026;
    wire n31029;
    wire n31032;
    wire n31035;
    wire n31038;
    wire n31041;
    wire n31044;
    wire n31047;
    wire n31050;
    wire n31053;
    wire n31056;
    wire n31059;
    wire n31062;
    wire n31065;
    wire n31068;
    wire n31071;
    wire n31074;
    wire n31077;
    wire n31080;
    wire n31083;
    wire n31086;
    wire n31089;
    wire n31092;
    wire n31095;
    wire n31098;
    wire n31101;
    wire n31104;
    wire n31107;
    wire n31110;
    wire n31113;
    wire n31116;
    wire n31119;
    wire n31122;
    wire n31125;
    wire n31128;
    wire n31131;
    wire n31134;
    wire n31137;
    wire n31140;
    wire n31143;
    wire n31146;
    wire n31149;
    wire n31152;
    wire n31155;
    wire n31158;
    wire n31161;
    wire n31164;
    wire n31167;
    wire n31170;
    wire n31173;
    wire n31176;
    wire n31179;
    wire n31182;
    wire n31185;
    wire n31188;
    wire n31191;
    wire n31194;
    wire n31197;
    wire n31200;
    wire n31203;
    wire n31206;
    wire n31209;
    wire n31212;
    wire n31215;
    wire n31218;
    wire n31221;
    wire n31224;
    wire n31227;
    wire n31230;
    wire n31233;
    wire n31236;
    wire n31239;
    wire n31242;
    wire n31245;
    wire n31248;
    wire n31251;
    wire n31254;
    wire n31257;
    wire n31260;
    wire n31263;
    wire n31266;
    wire n31269;
    wire n31272;
    wire n31275;
    wire n31278;
    wire n31281;
    wire n31284;
    wire n31287;
    wire n31290;
    wire n31293;
    wire n31296;
    wire n31299;
    wire n31302;
    wire n31305;
    wire n31308;
    wire n31311;
    wire n31314;
    wire n31317;
    wire n31320;
    wire n31323;
    wire n31326;
    wire n31329;
    wire n31332;
    wire n31335;
    wire n31338;
    wire n31341;
    wire n31344;
    wire n31347;
    wire n31350;
    wire n31353;
    wire n31356;
    wire n31359;
    wire n31362;
    wire n31365;
    wire n31368;
    wire n31371;
    wire n31374;
    wire n31377;
    wire n31380;
    wire n31383;
    wire n31386;
    wire n31389;
    wire n31392;
    wire n31395;
    wire n31398;
    wire n31401;
    wire n31404;
    wire n31407;
    wire n31410;
    wire n31413;
    wire n31416;
    wire n31419;
    wire n31422;
    wire n31425;
    wire n31428;
    wire n31431;
    wire n31434;
    wire n31437;
    wire n31440;
    wire n31443;
    wire n31446;
    wire n31449;
    wire n31452;
    wire n31455;
    wire n31458;
    wire n31461;
    wire n31464;
    wire n31467;
    wire n31470;
    wire n31473;
    wire n31476;
    wire n31479;
    wire n31482;
    wire n31485;
    wire n31488;
    wire n31491;
    wire n31494;
    wire n31497;
    wire n31500;
    wire n31503;
    wire n31506;
    wire n31509;
    wire n31511;
    wire n31514;
    wire n31517;
    wire n31521;
    wire n31523;
    wire n31526;
    wire n31529;
    wire n31533;
    wire n31535;
    wire n31538;
    wire n31542;
    wire n31545;
    wire n31548;
    wire n31550;
    wire n31553;
    wire n31556;
    wire n31559;
    wire n31562;
    wire n31565;
    wire n31568;
    wire n31571;
    wire n31574;
    wire n31577;
    wire n31580;
    wire n31583;
    wire n31586;
    wire n31589;
    wire n31592;
    wire n31595;
    wire n31598;
    wire n31601;
    wire n31604;
    wire n31607;
    wire n31610;
    wire n31613;
    wire n31616;
    wire n31619;
    wire n31622;
    wire n31625;
    wire n31628;
    wire n31631;
    wire n31634;
    wire n31637;
    wire n31640;
    wire n31643;
    wire n31646;
    wire n31649;
    wire n31652;
    wire n31655;
    wire n31658;
    wire n31661;
    wire n31664;
    wire n31667;
    wire n31670;
    wire n31673;
    wire n31676;
    wire n31679;
    wire n31682;
    wire n31685;
    wire n31688;
    wire n31691;
    wire n31694;
    wire n31697;
    wire n31700;
    wire n31703;
    wire n31706;
    wire n31709;
    wire n31712;
    wire n31715;
    wire n31718;
    wire n31721;
    wire n31724;
    wire n31727;
    wire n31730;
    wire n31733;
    wire n31736;
    wire n31739;
    wire n31742;
    wire n31745;
    wire n31748;
    wire n31751;
    wire n31754;
    wire n31757;
    wire n31760;
    wire n31763;
    wire n31766;
    wire n31772;
    wire n31775;
    wire n31778;
    wire n31781;
    wire n31784;
    wire n31787;
    wire n31790;
    wire n31793;
    wire n31796;
    wire n31799;
    wire n31802;
    wire n31805;
    wire n31808;
    wire n31811;
    wire n31814;
    wire n31817;
    wire n31820;
    wire n31823;
    wire n31826;
    wire n31829;
    wire n31832;
    wire n31835;
    wire n31838;
    wire n31841;
    wire n31844;
    wire n31847;
    wire n31850;
    wire n31853;
    wire n31856;
    wire n31859;
    wire n31862;
    wire n31865;
    wire n31868;
    wire n31871;
    wire n31874;
    wire n31877;
    wire n31880;
    wire n31883;
    wire n31886;
    wire n31889;
    wire n31892;
    wire n31895;
    wire n31898;
    wire n31901;
    wire n31904;
    wire n31907;
    wire n31910;
    wire n31913;
    wire n31916;
    wire n31919;
    wire n31922;
    wire n31925;
    wire n31928;
    wire n31931;
    wire n31934;
    wire n31937;
    wire n31940;
    wire n31943;
    wire n31946;
    wire n31949;
    wire n31952;
    wire n31955;
    wire n31958;
    wire n31961;
    wire n31964;
    wire n31967;
    wire n31970;
    wire n31973;
    wire n31976;
    wire n31982;
    wire n31985;
    wire n31988;
    wire n31991;
    wire n31994;
    wire n31997;
    wire n32000;
    wire n32003;
    wire n32006;
    wire n32009;
    wire n32012;
    wire n32015;
    wire n32018;
    wire n32021;
    wire n32024;
    wire n32027;
    wire n32030;
    wire n32033;
    wire n32036;
    wire n32039;
    wire n32042;
    wire n32045;
    wire n32048;
    wire n32051;
    wire n32054;
    wire n32057;
    wire n32060;
    wire n32063;
    wire n32066;
    wire n32069;
    wire n32072;
    wire n32075;
    wire n32078;
    wire n32081;
    wire n32084;
    wire n32087;
    wire n32090;
    wire n32093;
    wire n32096;
    wire n32099;
    wire n32102;
    wire n32105;
    wire n32108;
    wire n32111;
    wire n32114;
    wire n32117;
    wire n32120;
    wire n32123;
    wire n32126;
    wire n32129;
    wire n32132;
    wire n32135;
    wire n32138;
    wire n32141;
    wire n32144;
    wire n32147;
    wire n32150;
    wire n32153;
    wire n32156;
    wire n32159;
    wire n32162;
    wire n32165;
    wire n32168;
    wire n32171;
    wire n32174;
    wire n32177;
    wire n32180;
    wire n32183;
    wire n32189;
    wire n32192;
    wire n32195;
    wire n32198;
    wire n32201;
    wire n32204;
    wire n32207;
    wire n32210;
    wire n32213;
    wire n32216;
    wire n32219;
    wire n32222;
    wire n32225;
    wire n32228;
    wire n32231;
    wire n32234;
    wire n32237;
    wire n32240;
    wire n32243;
    wire n32246;
    wire n32249;
    wire n32252;
    wire n32255;
    wire n32258;
    wire n32261;
    wire n32264;
    wire n32267;
    wire n32270;
    wire n32273;
    wire n32276;
    wire n32279;
    wire n32282;
    wire n32285;
    wire n32288;
    wire n32291;
    wire n32294;
    wire n32297;
    wire n32300;
    wire n32303;
    wire n32306;
    wire n32309;
    wire n32312;
    wire n32315;
    wire n32318;
    wire n32321;
    wire n32324;
    wire n32327;
    wire n32330;
    wire n32333;
    wire n32336;
    wire n32339;
    wire n32342;
    wire n32345;
    wire n32348;
    wire n32351;
    wire n32354;
    wire n32357;
    wire n32360;
    wire n32363;
    wire n32366;
    wire n32369;
    wire n32372;
    wire n32375;
    wire n32378;
    wire n32381;
    wire n32387;
    wire n32390;
    wire n32393;
    wire n32396;
    wire n32399;
    wire n32402;
    wire n32405;
    wire n32408;
    wire n32411;
    wire n32414;
    wire n32417;
    wire n32420;
    wire n32423;
    wire n32426;
    wire n32429;
    wire n32432;
    wire n32435;
    wire n32438;
    wire n32441;
    wire n32444;
    wire n32447;
    wire n32450;
    wire n32453;
    wire n32456;
    wire n32459;
    wire n32462;
    wire n32465;
    wire n32468;
    wire n32471;
    wire n32474;
    wire n32477;
    wire n32480;
    wire n32483;
    wire n32486;
    wire n32489;
    wire n32492;
    wire n32495;
    wire n32498;
    wire n32501;
    wire n32504;
    wire n32507;
    wire n32510;
    wire n32513;
    wire n32516;
    wire n32519;
    wire n32522;
    wire n32525;
    wire n32528;
    wire n32531;
    wire n32534;
    wire n32537;
    wire n32540;
    wire n32543;
    wire n32546;
    wire n32549;
    wire n32552;
    wire n32555;
    wire n32558;
    wire n32561;
    wire n32564;
    wire n32567;
    wire n32570;
    wire n32576;
    wire n32579;
    wire n32582;
    wire n32585;
    wire n32588;
    wire n32591;
    wire n32594;
    wire n32597;
    wire n32600;
    wire n32603;
    wire n32606;
    wire n32609;
    wire n32612;
    wire n32615;
    wire n32618;
    wire n32621;
    wire n32624;
    wire n32627;
    wire n32630;
    wire n32633;
    wire n32636;
    wire n32639;
    wire n32642;
    wire n32645;
    wire n32648;
    wire n32651;
    wire n32654;
    wire n32657;
    wire n32660;
    wire n32663;
    wire n32666;
    wire n32669;
    wire n32672;
    wire n32675;
    wire n32678;
    wire n32681;
    wire n32684;
    wire n32687;
    wire n32690;
    wire n32693;
    wire n32696;
    wire n32699;
    wire n32702;
    wire n32705;
    wire n32708;
    wire n32711;
    wire n32714;
    wire n32717;
    wire n32720;
    wire n32723;
    wire n32726;
    wire n32729;
    wire n32732;
    wire n32735;
    wire n32738;
    wire n32741;
    wire n32744;
    wire n32747;
    wire n32750;
    wire n32756;
    wire n32759;
    wire n32762;
    wire n32765;
    wire n32768;
    wire n32771;
    wire n32774;
    wire n32777;
    wire n32780;
    wire n32783;
    wire n32786;
    wire n32789;
    wire n32792;
    wire n32795;
    wire n32798;
    wire n32801;
    wire n32804;
    wire n32807;
    wire n32810;
    wire n32813;
    wire n32816;
    wire n32819;
    wire n32822;
    wire n32825;
    wire n32828;
    wire n32831;
    wire n32834;
    wire n32837;
    wire n32840;
    wire n32843;
    wire n32846;
    wire n32849;
    wire n32852;
    wire n32855;
    wire n32858;
    wire n32861;
    wire n32864;
    wire n32867;
    wire n32870;
    wire n32873;
    wire n32876;
    wire n32879;
    wire n32882;
    wire n32885;
    wire n32888;
    wire n32891;
    wire n32894;
    wire n32897;
    wire n32900;
    wire n32903;
    wire n32906;
    wire n32909;
    wire n32912;
    wire n32915;
    wire n32918;
    wire n32921;
    wire n32927;
    wire n32930;
    wire n32933;
    wire n32936;
    wire n32939;
    wire n32942;
    wire n32945;
    wire n32948;
    wire n32951;
    wire n32954;
    wire n32957;
    wire n32960;
    wire n32963;
    wire n32966;
    wire n32969;
    wire n32972;
    wire n32975;
    wire n32978;
    wire n32981;
    wire n32984;
    wire n32987;
    wire n32990;
    wire n32993;
    wire n32996;
    wire n32999;
    wire n33002;
    wire n33005;
    wire n33008;
    wire n33011;
    wire n33014;
    wire n33017;
    wire n33020;
    wire n33023;
    wire n33026;
    wire n33029;
    wire n33032;
    wire n33035;
    wire n33038;
    wire n33041;
    wire n33044;
    wire n33047;
    wire n33050;
    wire n33053;
    wire n33056;
    wire n33059;
    wire n33062;
    wire n33065;
    wire n33068;
    wire n33071;
    wire n33074;
    wire n33077;
    wire n33080;
    wire n33083;
    wire n33089;
    wire n33092;
    wire n33095;
    wire n33098;
    wire n33101;
    wire n33104;
    wire n33107;
    wire n33110;
    wire n33113;
    wire n33116;
    wire n33119;
    wire n33122;
    wire n33125;
    wire n33128;
    wire n33131;
    wire n33134;
    wire n33137;
    wire n33140;
    wire n33143;
    wire n33146;
    wire n33149;
    wire n33152;
    wire n33155;
    wire n33158;
    wire n33161;
    wire n33164;
    wire n33167;
    wire n33170;
    wire n33173;
    wire n33176;
    wire n33179;
    wire n33182;
    wire n33185;
    wire n33188;
    wire n33191;
    wire n33194;
    wire n33197;
    wire n33200;
    wire n33203;
    wire n33206;
    wire n33209;
    wire n33212;
    wire n33215;
    wire n33218;
    wire n33221;
    wire n33224;
    wire n33227;
    wire n33230;
    wire n33233;
    wire n33236;
    wire n33242;
    wire n33245;
    wire n33248;
    wire n33251;
    wire n33254;
    wire n33257;
    wire n33260;
    wire n33263;
    wire n33266;
    wire n33269;
    wire n33272;
    wire n33275;
    wire n33278;
    wire n33281;
    wire n33284;
    wire n33287;
    wire n33290;
    wire n33293;
    wire n33296;
    wire n33299;
    wire n33302;
    wire n33305;
    wire n33308;
    wire n33311;
    wire n33314;
    wire n33317;
    wire n33320;
    wire n33323;
    wire n33326;
    wire n33329;
    wire n33332;
    wire n33335;
    wire n33338;
    wire n33341;
    wire n33344;
    wire n33347;
    wire n33350;
    wire n33353;
    wire n33356;
    wire n33359;
    wire n33362;
    wire n33365;
    wire n33368;
    wire n33371;
    wire n33374;
    wire n33377;
    wire n33380;
    wire n33386;
    wire n33389;
    wire n33392;
    wire n33395;
    wire n33398;
    wire n33401;
    wire n33404;
    wire n33407;
    wire n33410;
    wire n33413;
    wire n33416;
    wire n33419;
    wire n33422;
    wire n33425;
    wire n33428;
    wire n33431;
    wire n33434;
    wire n33437;
    wire n33440;
    wire n33443;
    wire n33446;
    wire n33449;
    wire n33452;
    wire n33455;
    wire n33458;
    wire n33461;
    wire n33464;
    wire n33467;
    wire n33470;
    wire n33473;
    wire n33476;
    wire n33479;
    wire n33482;
    wire n33485;
    wire n33488;
    wire n33491;
    wire n33494;
    wire n33497;
    wire n33500;
    wire n33503;
    wire n33506;
    wire n33509;
    wire n33512;
    wire n33515;
    wire n33521;
    wire n33524;
    wire n33527;
    wire n33530;
    wire n33533;
    wire n33536;
    wire n33539;
    wire n33542;
    wire n33545;
    wire n33548;
    wire n33551;
    wire n33554;
    wire n33557;
    wire n33560;
    wire n33563;
    wire n33566;
    wire n33569;
    wire n33572;
    wire n33575;
    wire n33578;
    wire n33581;
    wire n33584;
    wire n33587;
    wire n33590;
    wire n33593;
    wire n33596;
    wire n33599;
    wire n33602;
    wire n33605;
    wire n33608;
    wire n33611;
    wire n33614;
    wire n33617;
    wire n33620;
    wire n33623;
    wire n33626;
    wire n33629;
    wire n33632;
    wire n33635;
    wire n33638;
    wire n33641;
    wire n33647;
    wire n33650;
    wire n33653;
    wire n33656;
    wire n33659;
    wire n33662;
    wire n33665;
    wire n33668;
    wire n33671;
    wire n33674;
    wire n33677;
    wire n33680;
    wire n33683;
    wire n33686;
    wire n33689;
    wire n33692;
    wire n33695;
    wire n33698;
    wire n33701;
    wire n33704;
    wire n33707;
    wire n33710;
    wire n33713;
    wire n33716;
    wire n33719;
    wire n33722;
    wire n33725;
    wire n33728;
    wire n33731;
    wire n33734;
    wire n33737;
    wire n33740;
    wire n33743;
    wire n33746;
    wire n33749;
    wire n33752;
    wire n33755;
    wire n33758;
    wire n33764;
    wire n33767;
    wire n33770;
    wire n33773;
    wire n33776;
    wire n33779;
    wire n33782;
    wire n33785;
    wire n33788;
    wire n33791;
    wire n33794;
    wire n33797;
    wire n33800;
    wire n33803;
    wire n33806;
    wire n33809;
    wire n33812;
    wire n33815;
    wire n33818;
    wire n33821;
    wire n33824;
    wire n33827;
    wire n33830;
    wire n33833;
    wire n33836;
    wire n33839;
    wire n33842;
    wire n33845;
    wire n33848;
    wire n33851;
    wire n33854;
    wire n33857;
    wire n33860;
    wire n33863;
    wire n33866;
    wire n33872;
    wire n33875;
    wire n33878;
    wire n33881;
    wire n33884;
    wire n33887;
    wire n33890;
    wire n33893;
    wire n33896;
    wire n33899;
    wire n33902;
    wire n33905;
    wire n33908;
    wire n33911;
    wire n33914;
    wire n33917;
    wire n33920;
    wire n33923;
    wire n33926;
    wire n33929;
    wire n33932;
    wire n33935;
    wire n33938;
    wire n33941;
    wire n33944;
    wire n33947;
    wire n33950;
    wire n33953;
    wire n33956;
    wire n33959;
    wire n33962;
    wire n33965;
    wire n33971;
    wire n33974;
    wire n33977;
    wire n33980;
    wire n33983;
    wire n33986;
    wire n33989;
    wire n33992;
    wire n33995;
    wire n33998;
    wire n34001;
    wire n34004;
    wire n34007;
    wire n34010;
    wire n34013;
    wire n34016;
    wire n34019;
    wire n34022;
    wire n34025;
    wire n34028;
    wire n34031;
    wire n34034;
    wire n34037;
    wire n34040;
    wire n34043;
    wire n34046;
    wire n34049;
    wire n34052;
    wire n34055;
    wire n34061;
    wire n34064;
    wire n34067;
    wire n34070;
    wire n34073;
    wire n34076;
    wire n34079;
    wire n34082;
    wire n34085;
    wire n34088;
    wire n34091;
    wire n34094;
    wire n34097;
    wire n34100;
    wire n34103;
    wire n34106;
    wire n34109;
    wire n34112;
    wire n34115;
    wire n34118;
    wire n34121;
    wire n34124;
    wire n34127;
    wire n34130;
    wire n34133;
    wire n34136;
    wire n34139;
    wire n34145;
    wire n34148;
    wire n34151;
    wire n34154;
    wire n34157;
    wire n34160;
    wire n34163;
    wire n34166;
    wire n34169;
    wire n34172;
    wire n34175;
    wire n34178;
    wire n34181;
    wire n34184;
    wire n34187;
    wire n34190;
    wire n34193;
    wire n34196;
    wire n34199;
    wire n34202;
    wire n34205;
    wire n34208;
    wire n34211;
    wire n34214;
    wire n34217;
    wire n34223;
    wire n34226;
    wire n34229;
    wire n34232;
    wire n34235;
    wire n34238;
    wire n34241;
    wire n34244;
    wire n34247;
    wire n34250;
    wire n34253;
    wire n34256;
    wire n34259;
    wire n34262;
    wire n34265;
    wire n34268;
    wire n34271;
    wire n34274;
    wire n34277;
    wire n34280;
    wire n34283;
    wire n34286;
    wire n34289;
    wire n34292;
    wire n34298;
    wire n34301;
    wire n34304;
    wire n34307;
    wire n34310;
    wire n34313;
    wire n34316;
    wire n34319;
    wire n34322;
    wire n34325;
    wire n34328;
    wire n34331;
    wire n34334;
    wire n34337;
    wire n34340;
    wire n34343;
    wire n34346;
    wire n34349;
    wire n34352;
    wire n34355;
    wire n34358;
    wire n34361;
    wire n34367;
    wire n34370;
    wire n34373;
    wire n34376;
    wire n34379;
    wire n34382;
    wire n34385;
    wire n34388;
    wire n34391;
    wire n34394;
    wire n34397;
    wire n34400;
    wire n34403;
    wire n34406;
    wire n34409;
    wire n34412;
    wire n34415;
    wire n34418;
    wire n34421;
    wire n34424;
    wire n34430;
    wire n34433;
    wire n34436;
    wire n34439;
    wire n34442;
    wire n34445;
    wire n34448;
    wire n34451;
    wire n34454;
    wire n34457;
    wire n34460;
    wire n34463;
    wire n34466;
    wire n34469;
    wire n34472;
    wire n34475;
    wire n34478;
    wire n34481;
    wire n34487;
    wire n34490;
    wire n34493;
    wire n34496;
    wire n34499;
    wire n34502;
    wire n34505;
    wire n34508;
    wire n34511;
    wire n34514;
    wire n34517;
    wire n34520;
    wire n34523;
    wire n34526;
    wire n34529;
    wire n34532;
    wire n34538;
    wire n34541;
    wire n34544;
    wire n34547;
    wire n34550;
    wire n34553;
    wire n34556;
    wire n34559;
    wire n34562;
    wire n34565;
    wire n34568;
    wire n34571;
    wire n34574;
    wire n34577;
    wire n34583;
    wire n34586;
    wire n34589;
    wire n34592;
    wire n34595;
    wire n34598;
    wire n34601;
    wire n34604;
    wire n34607;
    wire n34610;
    wire n34613;
    wire n34616;
    wire n34622;
    wire n34625;
    wire n34628;
    wire n34631;
    wire n34634;
    wire n34637;
    wire n34640;
    wire n34643;
    wire n34646;
    wire n34649;
    wire n34655;
    wire n34658;
    wire n34661;
    wire n34664;
    wire n34667;
    wire n34670;
    wire n34673;
    wire n34676;
    wire n34682;
    wire n34685;
    wire n34688;
    wire n34691;
    wire n34694;
    wire n34697;
    wire n34703;
    wire n34706;
    wire n34709;
    wire n34712;
    wire n34718;
    wire n34721;
    jand g0000(.dinb(G1gat), .dina(G273gat), .dout(n67));
    jand g0001(.dinb(G18gat), .dina(G290gat), .dout(n71));
    jand g0002(.dinb(n67), .dina(n71), .dout(n75));
    jnot g0003(.din(n75), .dout(n78));
    jnot g0004(.din(G18gat), .dout(n81));
    jnot g0005(.din(G273gat), .dout(n84));
    jor g0006(.dinb(n81), .dina(n84), .dout(n88));
    jnot g0007(.din(n88), .dout(n91));
    jand g0008(.dinb(G1gat), .dina(G290gat), .dout(n95));
    jor g0009(.dinb(n91), .dina(n10596), .dout(n99));
    jand g0010(.dinb(n14544), .dina(n99), .dout(n103));
    jand g0011(.dinb(G1gat), .dina(G307gat), .dout(n107));
    jnot g0012(.din(n107), .dout(n110));
    jnot g0013(.din(G35gat), .dout(n113));
    jnot g0014(.din(G290gat), .dout(n116));
    jor g0015(.dinb(n113), .dina(n116), .dout(n120));
    jor g0016(.dinb(n88), .dina(n120), .dout(n124));
    jand g0017(.dinb(G35gat), .dina(G273gat), .dout(n128));
    jor g0018(.dinb(n71), .dina(n128), .dout(n132));
    jand g0019(.dinb(n124), .dina(n14559), .dout(n136));
    jxor g0020(.dinb(n14544), .dina(n136), .dout(n140));
    jxor g0021(.dinb(n10605), .dina(n140), .dout(n144));
    jand g0022(.dinb(G1gat), .dina(G324gat), .dout(n148));
    jnot g0023(.din(n148), .dout(n151));
    jor g0024(.dinb(n14561), .dina(n136), .dout(n155));
    jor g0025(.dinb(n14546), .dina(n140), .dout(n159));
    jand g0026(.dinb(n14541), .dina(n159), .dout(n163));
    jand g0027(.dinb(G18gat), .dina(G307gat), .dout(n167));
    jnot g0028(.din(n167), .dout(n170));
    jnot g0029(.din(n124), .dout(n173));
    jor g0030(.dinb(n113), .dina(n84), .dout(n177));
    jnot g0031(.din(G52gat), .dout(n180));
    jor g0032(.dinb(n180), .dina(n116), .dout(n184));
    jor g0033(.dinb(n177), .dina(n184), .dout(n188));
    jand g0034(.dinb(G35gat), .dina(G290gat), .dout(n192));
    jand g0035(.dinb(G52gat), .dina(G273gat), .dout(n196));
    jor g0036(.dinb(n192), .dina(n196), .dout(n200));
    jand g0037(.dinb(n188), .dina(n15747), .dout(n204));
    jxor g0038(.dinb(n173), .dina(n204), .dout(n208));
    jxor g0039(.dinb(n14538), .dina(n208), .dout(n212));
    jxor g0040(.dinb(n163), .dina(n14528), .dout(n216));
    jxor g0041(.dinb(n10623), .dina(n216), .dout(n220));
    jand g0042(.dinb(G1gat), .dina(G341gat), .dout(n224));
    jnot g0043(.din(n224), .dout(n227));
    jnot g0044(.din(n212), .dout(n230));
    jor g0045(.dinb(n163), .dina(n230), .dout(n234));
    jor g0046(.dinb(n14507), .dina(n216), .dout(n238));
    jand g0047(.dinb(n14505), .dina(n238), .dout(n242));
    jand g0048(.dinb(G18gat), .dina(G324gat), .dout(n246));
    jnot g0049(.din(n246), .dout(n249));
    jor g0050(.dinb(n173), .dina(n204), .dout(n253));
    jxor g0051(.dinb(n15749), .dina(n204), .dout(n257));
    jor g0052(.dinb(n15734), .dina(n257), .dout(n261));
    jand g0053(.dinb(n15732), .dina(n261), .dout(n265));
    jand g0054(.dinb(G35gat), .dina(G307gat), .dout(n269));
    jnot g0055(.din(n269), .dout(n272));
    jnot g0056(.din(n188), .dout(n275));
    jand g0057(.dinb(G69gat), .dina(G290gat), .dout(n279));
    jand g0058(.dinb(n196), .dina(n279), .dout(n283));
    jnot g0059(.din(n283), .dout(n286));
    jand g0060(.dinb(G52gat), .dina(G290gat), .dout(n290));
    jand g0061(.dinb(G69gat), .dina(G273gat), .dout(n294));
    jor g0062(.dinb(n290), .dina(n294), .dout(n298));
    jand g0063(.dinb(n286), .dina(n16788), .dout(n302));
    jxor g0064(.dinb(n275), .dina(n302), .dout(n306));
    jxor g0065(.dinb(n16785), .dina(n306), .dout(n310));
    jnot g0066(.din(n310), .dout(n313));
    jxor g0067(.dinb(n265), .dina(n313), .dout(n317));
    jxor g0068(.dinb(n14502), .dina(n317), .dout(n321));
    jxor g0069(.dinb(n242), .dina(n14483), .dout(n325));
    jxor g0070(.dinb(n10650), .dina(n325), .dout(n329));
    jand g0071(.dinb(G1gat), .dina(G358gat), .dout(n333));
    jnot g0072(.din(n333), .dout(n336));
    jnot g0073(.din(n321), .dout(n339));
    jor g0074(.dinb(n242), .dina(n339), .dout(n343));
    jor g0075(.dinb(n14453), .dina(n325), .dout(n347));
    jand g0076(.dinb(n14451), .dina(n347), .dout(n351));
    jand g0077(.dinb(G18gat), .dina(G341gat), .dout(n355));
    jnot g0078(.din(n355), .dout(n358));
    jor g0079(.dinb(n265), .dina(n313), .dout(n362));
    jxor g0080(.dinb(n265), .dina(n15728), .dout(n366));
    jor g0081(.dinb(n15707), .dina(n366), .dout(n370));
    jand g0082(.dinb(n15705), .dina(n370), .dout(n374));
    jand g0083(.dinb(G35gat), .dina(G324gat), .dout(n378));
    jnot g0084(.din(n378), .dout(n381));
    jor g0085(.dinb(n275), .dina(n302), .dout(n385));
    jnot g0086(.din(n385), .dout(n388));
    jand g0087(.dinb(n16785), .dina(n306), .dout(n392));
    jor g0088(.dinb(n388), .dina(n392), .dout(n396));
    jand g0089(.dinb(G52gat), .dina(G307gat), .dout(n400));
    jnot g0090(.din(n400), .dout(n403));
    jand g0091(.dinb(G86gat), .dina(G290gat), .dout(n407));
    jand g0092(.dinb(n294), .dina(n407), .dout(n411));
    jnot g0093(.din(n411), .dout(n414));
    jand g0094(.dinb(G86gat), .dina(G273gat), .dout(n418));
    jor g0095(.dinb(n279), .dina(n418), .dout(n422));
    jand g0096(.dinb(n414), .dina(n17841), .dout(n426));
    jxor g0097(.dinb(n17849), .dina(n426), .dout(n430));
    jxor g0098(.dinb(n17838), .dina(n430), .dout(n434));
    jxor g0099(.dinb(n396), .dina(n16776), .dout(n438));
    jxor g0100(.dinb(n16773), .dina(n438), .dout(n442));
    jnot g0101(.din(n442), .dout(n445));
    jxor g0102(.dinb(n374), .dina(n445), .dout(n449));
    jxor g0103(.dinb(n14448), .dina(n449), .dout(n453));
    jxor g0104(.dinb(n351), .dina(n14420), .dout(n457));
    jxor g0105(.dinb(n10686), .dina(n457), .dout(n461));
    jand g0106(.dinb(G1gat), .dina(G375gat), .dout(n465));
    jnot g0107(.din(n465), .dout(n468));
    jnot g0108(.din(n453), .dout(n471));
    jor g0109(.dinb(n351), .dina(n471), .dout(n475));
    jor g0110(.dinb(n14381), .dina(n457), .dout(n479));
    jand g0111(.dinb(n14379), .dina(n479), .dout(n483));
    jand g0112(.dinb(G18gat), .dina(G358gat), .dout(n487));
    jnot g0113(.din(n487), .dout(n490));
    jor g0114(.dinb(n374), .dina(n445), .dout(n494));
    jxor g0115(.dinb(n374), .dina(n15701), .dout(n498));
    jor g0116(.dinb(n15671), .dina(n498), .dout(n502));
    jand g0117(.dinb(n15669), .dina(n502), .dout(n506));
    jand g0118(.dinb(G35gat), .dina(G341gat), .dout(n510));
    jnot g0119(.din(n510), .dout(n513));
    jand g0120(.dinb(n396), .dina(n16776), .dout(n517));
    jand g0121(.dinb(n16773), .dina(n438), .dout(n521));
    jor g0122(.dinb(n16755), .dina(n521), .dout(n525));
    jand g0123(.dinb(G52gat), .dina(G324gat), .dout(n529));
    jnot g0124(.din(n529), .dout(n532));
    jnot g0125(.din(n426), .dout(n535));
    jand g0126(.dinb(n17843), .dina(n535), .dout(n539));
    jand g0127(.dinb(n17838), .dina(n430), .dout(n543));
    jor g0128(.dinb(n539), .dina(n543), .dout(n547));
    jand g0129(.dinb(G69gat), .dina(G307gat), .dout(n551));
    jnot g0130(.din(n551), .dout(n554));
    jand g0131(.dinb(G103gat), .dina(G290gat), .dout(n558));
    jand g0132(.dinb(n418), .dina(n558), .dout(n562));
    jnot g0133(.din(n562), .dout(n565));
    jand g0134(.dinb(G103gat), .dina(G273gat), .dout(n569));
    jor g0135(.dinb(n407), .dina(n569), .dout(n573));
    jand g0136(.dinb(n565), .dina(n18888), .dout(n577));
    jxor g0137(.dinb(n18896), .dina(n577), .dout(n581));
    jxor g0138(.dinb(n18885), .dina(n581), .dout(n585));
    jxor g0139(.dinb(n547), .dina(n17829), .dout(n589));
    jxor g0140(.dinb(n17826), .dina(n589), .dout(n593));
    jxor g0141(.dinb(n525), .dina(n16752), .dout(n597));
    jxor g0142(.dinb(n16749), .dina(n597), .dout(n601));
    jnot g0143(.din(n601), .dout(n604));
    jxor g0144(.dinb(n506), .dina(n604), .dout(n608));
    jxor g0145(.dinb(n14376), .dina(n608), .dout(n612));
    jxor g0146(.dinb(n483), .dina(n14339), .dout(n616));
    jxor g0147(.dinb(n10731), .dina(n616), .dout(n620));
    jand g0148(.dinb(G1gat), .dina(G392gat), .dout(n624));
    jnot g0149(.din(n624), .dout(n627));
    jnot g0150(.din(n612), .dout(n630));
    jor g0151(.dinb(n483), .dina(n630), .dout(n634));
    jor g0152(.dinb(n14291), .dina(n616), .dout(n638));
    jand g0153(.dinb(n14289), .dina(n638), .dout(n642));
    jand g0154(.dinb(G18gat), .dina(G375gat), .dout(n646));
    jnot g0155(.din(n646), .dout(n649));
    jor g0156(.dinb(n506), .dina(n604), .dout(n653));
    jxor g0157(.dinb(n506), .dina(n15665), .dout(n657));
    jor g0158(.dinb(n15626), .dina(n657), .dout(n661));
    jand g0159(.dinb(n15624), .dina(n661), .dout(n665));
    jand g0160(.dinb(G35gat), .dina(G358gat), .dout(n669));
    jnot g0161(.din(n669), .dout(n672));
    jand g0162(.dinb(n525), .dina(n16752), .dout(n676));
    jand g0163(.dinb(n16749), .dina(n597), .dout(n680));
    jor g0164(.dinb(n16722), .dina(n680), .dout(n684));
    jand g0165(.dinb(G52gat), .dina(G341gat), .dout(n688));
    jnot g0166(.din(n688), .dout(n691));
    jand g0167(.dinb(n547), .dina(n17829), .dout(n695));
    jand g0168(.dinb(n17826), .dina(n589), .dout(n699));
    jor g0169(.dinb(n17808), .dina(n699), .dout(n703));
    jand g0170(.dinb(G69gat), .dina(G324gat), .dout(n707));
    jnot g0171(.din(n707), .dout(n710));
    jnot g0172(.din(n577), .dout(n713));
    jand g0173(.dinb(n18890), .dina(n713), .dout(n717));
    jand g0174(.dinb(n18885), .dina(n581), .dout(n721));
    jor g0175(.dinb(n717), .dina(n721), .dout(n725));
    jand g0176(.dinb(G86gat), .dina(G307gat), .dout(n729));
    jnot g0177(.din(n729), .dout(n732));
    jand g0178(.dinb(G120gat), .dina(G290gat), .dout(n736));
    jand g0179(.dinb(n569), .dina(n736), .dout(n740));
    jnot g0180(.din(n740), .dout(n743));
    jand g0181(.dinb(G120gat), .dina(G273gat), .dout(n747));
    jor g0182(.dinb(n558), .dina(n747), .dout(n751));
    jand g0183(.dinb(n743), .dina(n19902), .dout(n755));
    jxor g0184(.dinb(n19910), .dina(n755), .dout(n759));
    jxor g0185(.dinb(n19899), .dina(n759), .dout(n763));
    jxor g0186(.dinb(n725), .dina(n18876), .dout(n767));
    jxor g0187(.dinb(n18873), .dina(n767), .dout(n771));
    jxor g0188(.dinb(n703), .dina(n17805), .dout(n775));
    jxor g0189(.dinb(n17802), .dina(n775), .dout(n779));
    jxor g0190(.dinb(n684), .dina(n16719), .dout(n783));
    jxor g0191(.dinb(n16716), .dina(n783), .dout(n787));
    jnot g0192(.din(n787), .dout(n790));
    jxor g0193(.dinb(n665), .dina(n790), .dout(n794));
    jxor g0194(.dinb(n14286), .dina(n794), .dout(n798));
    jxor g0195(.dinb(n642), .dina(n14240), .dout(n802));
    jxor g0196(.dinb(n10785), .dina(n802), .dout(n806));
    jand g0197(.dinb(G1gat), .dina(G409gat), .dout(n810));
    jnot g0198(.din(n810), .dout(n813));
    jnot g0199(.din(n798), .dout(n816));
    jor g0200(.dinb(n642), .dina(n816), .dout(n820));
    jor g0201(.dinb(n14183), .dina(n802), .dout(n824));
    jand g0202(.dinb(n14181), .dina(n824), .dout(n828));
    jand g0203(.dinb(G18gat), .dina(G392gat), .dout(n832));
    jnot g0204(.din(n832), .dout(n835));
    jor g0205(.dinb(n665), .dina(n790), .dout(n839));
    jxor g0206(.dinb(n665), .dina(n15620), .dout(n843));
    jor g0207(.dinb(n15572), .dina(n843), .dout(n847));
    jand g0208(.dinb(n15570), .dina(n847), .dout(n851));
    jand g0209(.dinb(G35gat), .dina(G375gat), .dout(n855));
    jnot g0210(.din(n855), .dout(n858));
    jand g0211(.dinb(n684), .dina(n16719), .dout(n862));
    jand g0212(.dinb(n16716), .dina(n783), .dout(n866));
    jor g0213(.dinb(n16680), .dina(n866), .dout(n870));
    jand g0214(.dinb(G52gat), .dina(G358gat), .dout(n874));
    jnot g0215(.din(n874), .dout(n877));
    jand g0216(.dinb(n703), .dina(n17805), .dout(n881));
    jand g0217(.dinb(n17802), .dina(n775), .dout(n885));
    jor g0218(.dinb(n17775), .dina(n885), .dout(n889));
    jand g0219(.dinb(G69gat), .dina(G341gat), .dout(n893));
    jnot g0220(.din(n893), .dout(n896));
    jand g0221(.dinb(n725), .dina(n18876), .dout(n900));
    jand g0222(.dinb(n18873), .dina(n767), .dout(n904));
    jor g0223(.dinb(n18855), .dina(n904), .dout(n908));
    jand g0224(.dinb(G86gat), .dina(G324gat), .dout(n912));
    jnot g0225(.din(n912), .dout(n915));
    jor g0226(.dinb(n19904), .dina(n755), .dout(n919));
    jnot g0227(.din(n919), .dout(n922));
    jand g0228(.dinb(n19899), .dina(n759), .dout(n926));
    jor g0229(.dinb(n922), .dina(n926), .dout(n930));
    jand g0230(.dinb(G103gat), .dina(G307gat), .dout(n934));
    jnot g0231(.din(n934), .dout(n937));
    jand g0232(.dinb(G137gat), .dina(G290gat), .dout(n941));
    jand g0233(.dinb(n747), .dina(n941), .dout(n945));
    jnot g0234(.din(n945), .dout(n948));
    jand g0235(.dinb(G137gat), .dina(G273gat), .dout(n952));
    jor g0236(.dinb(n736), .dina(n952), .dout(n956));
    jand g0237(.dinb(n948), .dina(n20952), .dout(n960));
    jxor g0238(.dinb(n20960), .dina(n960), .dout(n964));
    jxor g0239(.dinb(n20949), .dina(n964), .dout(n968));
    jxor g0240(.dinb(n930), .dina(n19890), .dout(n972));
    jxor g0241(.dinb(n19887), .dina(n972), .dout(n976));
    jxor g0242(.dinb(n908), .dina(n18852), .dout(n980));
    jxor g0243(.dinb(n18849), .dina(n980), .dout(n984));
    jxor g0244(.dinb(n889), .dina(n17772), .dout(n988));
    jxor g0245(.dinb(n17769), .dina(n988), .dout(n992));
    jxor g0246(.dinb(n870), .dina(n16677), .dout(n996));
    jxor g0247(.dinb(n16674), .dina(n996), .dout(n1000));
    jnot g0248(.din(n1000), .dout(n1003));
    jxor g0249(.dinb(n851), .dina(n1003), .dout(n1007));
    jxor g0250(.dinb(n14178), .dina(n1007), .dout(n1011));
    jxor g0251(.dinb(n828), .dina(n14123), .dout(n1015));
    jxor g0252(.dinb(n10848), .dina(n1015), .dout(n1019));
    jand g0253(.dinb(G1gat), .dina(G426gat), .dout(n1023));
    jnot g0254(.din(n1023), .dout(n1026));
    jnot g0255(.din(n1011), .dout(n1029));
    jor g0256(.dinb(n828), .dina(n1029), .dout(n1033));
    jor g0257(.dinb(n14057), .dina(n1015), .dout(n1037));
    jand g0258(.dinb(n14055), .dina(n1037), .dout(n1041));
    jand g0259(.dinb(G18gat), .dina(G409gat), .dout(n1045));
    jnot g0260(.din(n1045), .dout(n1048));
    jor g0261(.dinb(n851), .dina(n1003), .dout(n1052));
    jxor g0262(.dinb(n851), .dina(n15566), .dout(n1056));
    jor g0263(.dinb(n15509), .dina(n1056), .dout(n1060));
    jand g0264(.dinb(n15507), .dina(n1060), .dout(n1064));
    jand g0265(.dinb(G35gat), .dina(G392gat), .dout(n1068));
    jnot g0266(.din(n1068), .dout(n1071));
    jand g0267(.dinb(n870), .dina(n16677), .dout(n1075));
    jand g0268(.dinb(n16674), .dina(n996), .dout(n1079));
    jor g0269(.dinb(n16629), .dina(n1079), .dout(n1083));
    jand g0270(.dinb(G52gat), .dina(G375gat), .dout(n1087));
    jnot g0271(.din(n1087), .dout(n1090));
    jand g0272(.dinb(n889), .dina(n17772), .dout(n1094));
    jand g0273(.dinb(n17769), .dina(n988), .dout(n1098));
    jor g0274(.dinb(n17733), .dina(n1098), .dout(n1102));
    jand g0275(.dinb(G69gat), .dina(G358gat), .dout(n1106));
    jnot g0276(.din(n1106), .dout(n1109));
    jand g0277(.dinb(n908), .dina(n18852), .dout(n1113));
    jand g0278(.dinb(n18849), .dina(n980), .dout(n1117));
    jor g0279(.dinb(n18822), .dina(n1117), .dout(n1121));
    jand g0280(.dinb(G86gat), .dina(G341gat), .dout(n1125));
    jnot g0281(.din(n1125), .dout(n1128));
    jand g0282(.dinb(n930), .dina(n19890), .dout(n1132));
    jand g0283(.dinb(n19887), .dina(n972), .dout(n1136));
    jor g0284(.dinb(n19869), .dina(n1136), .dout(n1140));
    jand g0285(.dinb(G103gat), .dina(G324gat), .dout(n1144));
    jnot g0286(.din(n1144), .dout(n1147));
    jor g0287(.dinb(n20954), .dina(n960), .dout(n1151));
    jnot g0288(.din(n1151), .dout(n1154));
    jand g0289(.dinb(n20949), .dina(n964), .dout(n1158));
    jor g0290(.dinb(n1154), .dina(n1158), .dout(n1162));
    jand g0291(.dinb(G120gat), .dina(G307gat), .dout(n1166));
    jnot g0292(.din(n1166), .dout(n1169));
    jand g0293(.dinb(G154gat), .dina(G290gat), .dout(n1173));
    jand g0294(.dinb(n952), .dina(n1173), .dout(n1177));
    jnot g0295(.din(n1177), .dout(n1180));
    jand g0296(.dinb(G154gat), .dina(G273gat), .dout(n1184));
    jor g0297(.dinb(n941), .dina(n1184), .dout(n1188));
    jand g0298(.dinb(n1180), .dina(n22089), .dout(n1192));
    jxor g0299(.dinb(n22097), .dina(n1192), .dout(n1196));
    jxor g0300(.dinb(n22086), .dina(n1196), .dout(n1200));
    jxor g0301(.dinb(n1162), .dina(n20940), .dout(n1204));
    jxor g0302(.dinb(n20937), .dina(n1204), .dout(n1208));
    jxor g0303(.dinb(n1140), .dina(n19866), .dout(n1212));
    jxor g0304(.dinb(n19863), .dina(n1212), .dout(n1216));
    jxor g0305(.dinb(n1121), .dina(n18819), .dout(n1220));
    jxor g0306(.dinb(n18816), .dina(n1220), .dout(n1224));
    jxor g0307(.dinb(n1102), .dina(n17730), .dout(n1228));
    jxor g0308(.dinb(n17727), .dina(n1228), .dout(n1232));
    jxor g0309(.dinb(n1083), .dina(n16626), .dout(n1236));
    jxor g0310(.dinb(n16623), .dina(n1236), .dout(n1240));
    jnot g0311(.din(n1240), .dout(n1243));
    jxor g0312(.dinb(n1064), .dina(n1243), .dout(n1247));
    jxor g0313(.dinb(n14052), .dina(n1247), .dout(n1251));
    jxor g0314(.dinb(n1041), .dina(n13988), .dout(n1255));
    jxor g0315(.dinb(n10920), .dina(n1255), .dout(n1259));
    jand g0316(.dinb(G1gat), .dina(G443gat), .dout(n1263));
    jnot g0317(.din(n1263), .dout(n1266));
    jnot g0318(.din(n1251), .dout(n1269));
    jor g0319(.dinb(n1041), .dina(n1269), .dout(n1273));
    jor g0320(.dinb(n13913), .dina(n1255), .dout(n1277));
    jand g0321(.dinb(n13911), .dina(n1277), .dout(n1281));
    jand g0322(.dinb(G18gat), .dina(G426gat), .dout(n1285));
    jnot g0323(.din(n1285), .dout(n1288));
    jor g0324(.dinb(n1064), .dina(n1243), .dout(n1292));
    jxor g0325(.dinb(n1064), .dina(n15503), .dout(n1296));
    jor g0326(.dinb(n15437), .dina(n1296), .dout(n1300));
    jand g0327(.dinb(n15435), .dina(n1300), .dout(n1304));
    jand g0328(.dinb(G35gat), .dina(G409gat), .dout(n1308));
    jnot g0329(.din(n1308), .dout(n1311));
    jand g0330(.dinb(n1083), .dina(n16626), .dout(n1315));
    jand g0331(.dinb(n16623), .dina(n1236), .dout(n1319));
    jor g0332(.dinb(n16569), .dina(n1319), .dout(n1323));
    jand g0333(.dinb(G52gat), .dina(G392gat), .dout(n1327));
    jnot g0334(.din(n1327), .dout(n1330));
    jand g0335(.dinb(n1102), .dina(n17730), .dout(n1334));
    jand g0336(.dinb(n17727), .dina(n1228), .dout(n1338));
    jor g0337(.dinb(n17682), .dina(n1338), .dout(n1342));
    jand g0338(.dinb(G69gat), .dina(G375gat), .dout(n1346));
    jnot g0339(.din(n1346), .dout(n1349));
    jand g0340(.dinb(n1121), .dina(n18819), .dout(n1353));
    jand g0341(.dinb(n18816), .dina(n1220), .dout(n1357));
    jor g0342(.dinb(n18780), .dina(n1357), .dout(n1361));
    jand g0343(.dinb(G86gat), .dina(G358gat), .dout(n1365));
    jnot g0344(.din(n1365), .dout(n1368));
    jand g0345(.dinb(n1140), .dina(n19866), .dout(n1372));
    jand g0346(.dinb(n19863), .dina(n1212), .dout(n1376));
    jor g0347(.dinb(n19836), .dina(n1376), .dout(n1380));
    jand g0348(.dinb(G103gat), .dina(G341gat), .dout(n1384));
    jnot g0349(.din(n1384), .dout(n1387));
    jand g0350(.dinb(n1162), .dina(n20940), .dout(n1391));
    jand g0351(.dinb(n20937), .dina(n1204), .dout(n1395));
    jor g0352(.dinb(n20919), .dina(n1395), .dout(n1399));
    jand g0353(.dinb(G120gat), .dina(G324gat), .dout(n1403));
    jnot g0354(.din(n1403), .dout(n1406));
    jor g0355(.dinb(n22091), .dina(n1192), .dout(n1410));
    jand g0356(.dinb(n22086), .dina(n1196), .dout(n1414));
    jnot g0357(.din(n1414), .dout(n1417));
    jand g0358(.dinb(n22077), .dina(n1417), .dout(n1421));
    jnot g0359(.din(n1421), .dout(n1424));
    jand g0360(.dinb(G137gat), .dina(G307gat), .dout(n1428));
    jnot g0361(.din(n1428), .dout(n1431));
    jand g0362(.dinb(G171gat), .dina(G290gat), .dout(n1435));
    jand g0363(.dinb(n1184), .dina(n1435), .dout(n1439));
    jnot g0364(.din(n1439), .dout(n1442));
    jand g0365(.dinb(G171gat), .dina(G273gat), .dout(n1446));
    jor g0366(.dinb(n1173), .dina(n1446), .dout(n1450));
    jand g0367(.dinb(n1442), .dina(n23226), .dout(n1454));
    jxor g0368(.dinb(n23234), .dina(n1454), .dout(n1458));
    jxor g0369(.dinb(n23223), .dina(n1458), .dout(n1462));
    jxor g0370(.dinb(n1424), .dina(n22071), .dout(n1466));
    jxor g0371(.dinb(n22062), .dina(n1466), .dout(n1470));
    jxor g0372(.dinb(n20916), .dina(n1470), .dout(n1474));
    jxor g0373(.dinb(n20913), .dina(n1474), .dout(n1478));
    jxor g0374(.dinb(n1380), .dina(n1478), .dout(n1482));
    jxor g0375(.dinb(n19833), .dina(n1482), .dout(n1486));
    jxor g0376(.dinb(n1361), .dina(n18777), .dout(n1490));
    jxor g0377(.dinb(n18774), .dina(n1490), .dout(n1494));
    jxor g0378(.dinb(n1342), .dina(n17679), .dout(n1498));
    jxor g0379(.dinb(n17676), .dina(n1498), .dout(n1502));
    jxor g0380(.dinb(n1323), .dina(n16566), .dout(n1506));
    jxor g0381(.dinb(n16563), .dina(n1506), .dout(n1510));
    jnot g0382(.din(n1510), .dout(n1513));
    jxor g0383(.dinb(n1304), .dina(n1513), .dout(n1517));
    jxor g0384(.dinb(n13908), .dina(n1517), .dout(n1521));
    jxor g0385(.dinb(n1281), .dina(n13835), .dout(n1525));
    jxor g0386(.dinb(n11001), .dina(n1525), .dout(n1529));
    jand g0387(.dinb(G1gat), .dina(G460gat), .dout(n1533));
    jnot g0388(.din(n1533), .dout(n1536));
    jnot g0389(.din(n1521), .dout(n1539));
    jor g0390(.dinb(n1281), .dina(n1539), .dout(n1543));
    jor g0391(.dinb(n13751), .dina(n1525), .dout(n1547));
    jand g0392(.dinb(n13749), .dina(n1547), .dout(n1551));
    jand g0393(.dinb(G18gat), .dina(G443gat), .dout(n1555));
    jnot g0394(.din(n1555), .dout(n1558));
    jor g0395(.dinb(n1304), .dina(n1513), .dout(n1562));
    jxor g0396(.dinb(n1304), .dina(n15431), .dout(n1566));
    jor g0397(.dinb(n15356), .dina(n1566), .dout(n1570));
    jand g0398(.dinb(n15354), .dina(n1570), .dout(n1574));
    jand g0399(.dinb(G35gat), .dina(G426gat), .dout(n1578));
    jnot g0400(.din(n1578), .dout(n1581));
    jand g0401(.dinb(n1323), .dina(n16566), .dout(n1585));
    jand g0402(.dinb(n16563), .dina(n1506), .dout(n1589));
    jor g0403(.dinb(n16500), .dina(n1589), .dout(n1593));
    jand g0404(.dinb(G52gat), .dina(G409gat), .dout(n1597));
    jnot g0405(.din(n1597), .dout(n1600));
    jand g0406(.dinb(n1342), .dina(n17679), .dout(n1604));
    jand g0407(.dinb(n17676), .dina(n1498), .dout(n1608));
    jor g0408(.dinb(n17622), .dina(n1608), .dout(n1612));
    jand g0409(.dinb(G69gat), .dina(G392gat), .dout(n1616));
    jnot g0410(.din(n1616), .dout(n1619));
    jand g0411(.dinb(n1361), .dina(n18777), .dout(n1623));
    jand g0412(.dinb(n18774), .dina(n1490), .dout(n1627));
    jor g0413(.dinb(n18729), .dina(n1627), .dout(n1631));
    jand g0414(.dinb(G86gat), .dina(G375gat), .dout(n1635));
    jnot g0415(.din(n1635), .dout(n1638));
    jand g0416(.dinb(n1380), .dina(n1478), .dout(n1642));
    jand g0417(.dinb(n19833), .dina(n1482), .dout(n1646));
    jor g0418(.dinb(n19797), .dina(n1646), .dout(n1650));
    jand g0419(.dinb(G103gat), .dina(G358gat), .dout(n1654));
    jnot g0420(.din(n1654), .dout(n1657));
    jand g0421(.dinb(n20916), .dina(n1470), .dout(n1661));
    jand g0422(.dinb(n20913), .dina(n1474), .dout(n1665));
    jor g0423(.dinb(n20883), .dina(n1665), .dout(n1669));
    jand g0424(.dinb(G120gat), .dina(G341gat), .dout(n1673));
    jnot g0425(.din(n1673), .dout(n1676));
    jand g0426(.dinb(n1424), .dina(n22071), .dout(n1680));
    jand g0427(.dinb(n22062), .dina(n1466), .dout(n1684));
    jor g0428(.dinb(n22038), .dina(n1684), .dout(n1688));
    jand g0429(.dinb(G137gat), .dina(G324gat), .dout(n1692));
    jnot g0430(.din(n1692), .dout(n1695));
    jor g0431(.dinb(n23228), .dina(n1454), .dout(n1699));
    jand g0432(.dinb(n23223), .dina(n1458), .dout(n1703));
    jnot g0433(.din(n1703), .dout(n1706));
    jand g0434(.dinb(n23214), .dina(n1706), .dout(n1710));
    jnot g0435(.din(n1710), .dout(n1713));
    jand g0436(.dinb(G154gat), .dina(G307gat), .dout(n1717));
    jnot g0437(.din(n1717), .dout(n1720));
    jand g0438(.dinb(G188gat), .dina(G290gat), .dout(n1724));
    jand g0439(.dinb(n1446), .dina(n1724), .dout(n1728));
    jnot g0440(.din(n1728), .dout(n1731));
    jand g0441(.dinb(G188gat), .dina(G273gat), .dout(n1735));
    jor g0442(.dinb(n1435), .dina(n1735), .dout(n1739));
    jand g0443(.dinb(n1731), .dina(n24360), .dout(n1743));
    jxor g0444(.dinb(n24368), .dina(n1743), .dout(n1747));
    jxor g0445(.dinb(n24357), .dina(n1747), .dout(n1751));
    jxor g0446(.dinb(n1713), .dina(n23208), .dout(n1755));
    jxor g0447(.dinb(n23199), .dina(n1755), .dout(n1759));
    jxor g0448(.dinb(n1688), .dina(n22035), .dout(n1763));
    jxor g0449(.dinb(n22032), .dina(n1763), .dout(n1767));
    jxor g0450(.dinb(n1669), .dina(n1767), .dout(n1771));
    jxor g0451(.dinb(n20880), .dina(n1771), .dout(n1775));
    jxor g0452(.dinb(n1650), .dina(n1775), .dout(n1779));
    jxor g0453(.dinb(n19794), .dina(n1779), .dout(n1783));
    jxor g0454(.dinb(n1631), .dina(n18726), .dout(n1787));
    jxor g0455(.dinb(n18723), .dina(n1787), .dout(n1791));
    jxor g0456(.dinb(n1612), .dina(n17619), .dout(n1795));
    jxor g0457(.dinb(n17616), .dina(n1795), .dout(n1799));
    jxor g0458(.dinb(n1593), .dina(n16497), .dout(n1803));
    jxor g0459(.dinb(n16494), .dina(n1803), .dout(n1807));
    jnot g0460(.din(n1807), .dout(n1810));
    jxor g0461(.dinb(n1574), .dina(n1810), .dout(n1814));
    jxor g0462(.dinb(n13746), .dina(n1814), .dout(n1818));
    jxor g0463(.dinb(n1551), .dina(n13664), .dout(n1822));
    jxor g0464(.dinb(n11091), .dina(n1822), .dout(n1826));
    jand g0465(.dinb(G1gat), .dina(G477gat), .dout(n1830));
    jnot g0466(.din(n1830), .dout(n1833));
    jnot g0467(.din(n1818), .dout(n1836));
    jor g0468(.dinb(n1551), .dina(n1836), .dout(n1840));
    jor g0469(.dinb(n13571), .dina(n1822), .dout(n1844));
    jand g0470(.dinb(n13569), .dina(n1844), .dout(n1848));
    jand g0471(.dinb(G18gat), .dina(G460gat), .dout(n1852));
    jnot g0472(.din(n1852), .dout(n1855));
    jor g0473(.dinb(n1574), .dina(n1810), .dout(n1859));
    jxor g0474(.dinb(n1574), .dina(n15350), .dout(n1863));
    jor g0475(.dinb(n15266), .dina(n1863), .dout(n1867));
    jand g0476(.dinb(n15264), .dina(n1867), .dout(n1871));
    jand g0477(.dinb(G35gat), .dina(G443gat), .dout(n1875));
    jnot g0478(.din(n1875), .dout(n1878));
    jand g0479(.dinb(n1593), .dina(n16497), .dout(n1882));
    jand g0480(.dinb(n16494), .dina(n1803), .dout(n1886));
    jor g0481(.dinb(n16422), .dina(n1886), .dout(n1890));
    jand g0482(.dinb(G52gat), .dina(G426gat), .dout(n1894));
    jnot g0483(.din(n1894), .dout(n1897));
    jand g0484(.dinb(n1612), .dina(n17619), .dout(n1901));
    jand g0485(.dinb(n17616), .dina(n1795), .dout(n1905));
    jor g0486(.dinb(n17553), .dina(n1905), .dout(n1909));
    jand g0487(.dinb(G69gat), .dina(G409gat), .dout(n1913));
    jnot g0488(.din(n1913), .dout(n1916));
    jand g0489(.dinb(n1631), .dina(n18726), .dout(n1920));
    jand g0490(.dinb(n18723), .dina(n1787), .dout(n1924));
    jor g0491(.dinb(n18669), .dina(n1924), .dout(n1928));
    jand g0492(.dinb(G86gat), .dina(G392gat), .dout(n1932));
    jnot g0493(.din(n1932), .dout(n1935));
    jand g0494(.dinb(n1650), .dina(n1775), .dout(n1939));
    jand g0495(.dinb(n19794), .dina(n1779), .dout(n1943));
    jor g0496(.dinb(n19749), .dina(n1943), .dout(n1947));
    jand g0497(.dinb(G103gat), .dina(G375gat), .dout(n1951));
    jnot g0498(.din(n1951), .dout(n1954));
    jand g0499(.dinb(n1669), .dina(n1767), .dout(n1958));
    jand g0500(.dinb(n20880), .dina(n1771), .dout(n1962));
    jor g0501(.dinb(n20841), .dina(n1962), .dout(n1966));
    jand g0502(.dinb(G120gat), .dina(G358gat), .dout(n1970));
    jnot g0503(.din(n1970), .dout(n1973));
    jand g0504(.dinb(n1688), .dina(n22035), .dout(n1977));
    jand g0505(.dinb(n22032), .dina(n1763), .dout(n1981));
    jor g0506(.dinb(n21999), .dina(n1981), .dout(n1985));
    jand g0507(.dinb(G137gat), .dina(G341gat), .dout(n1989));
    jnot g0508(.din(n1989), .dout(n1992));
    jand g0509(.dinb(n1713), .dina(n23208), .dout(n1996));
    jand g0510(.dinb(n23199), .dina(n1755), .dout(n2000));
    jor g0511(.dinb(n23175), .dina(n2000), .dout(n2004));
    jand g0512(.dinb(G154gat), .dina(G324gat), .dout(n2008));
    jnot g0513(.din(n2008), .dout(n2011));
    jor g0514(.dinb(n24362), .dina(n1743), .dout(n2015));
    jand g0515(.dinb(n24357), .dina(n1747), .dout(n2019));
    jnot g0516(.din(n2019), .dout(n2022));
    jand g0517(.dinb(n24348), .dina(n2022), .dout(n2026));
    jnot g0518(.din(n2026), .dout(n2029));
    jand g0519(.dinb(G171gat), .dina(G307gat), .dout(n2033));
    jnot g0520(.din(n2033), .dout(n2036));
    jand g0521(.dinb(G205gat), .dina(G290gat), .dout(n2040));
    jand g0522(.dinb(n1735), .dina(n2040), .dout(n2044));
    jnot g0523(.din(n2044), .dout(n2047));
    jand g0524(.dinb(G205gat), .dina(G273gat), .dout(n2051));
    jor g0525(.dinb(n1724), .dina(n2051), .dout(n2055));
    jand g0526(.dinb(n2047), .dina(n25500), .dout(n2059));
    jxor g0527(.dinb(n25508), .dina(n2059), .dout(n2063));
    jxor g0528(.dinb(n25497), .dina(n2063), .dout(n2067));
    jxor g0529(.dinb(n2029), .dina(n24342), .dout(n2071));
    jxor g0530(.dinb(n24333), .dina(n2071), .dout(n2075));
    jxor g0531(.dinb(n2004), .dina(n23172), .dout(n2079));
    jxor g0532(.dinb(n23169), .dina(n2079), .dout(n2083));
    jxor g0533(.dinb(n1985), .dina(n21996), .dout(n2087));
    jxor g0534(.dinb(n21993), .dina(n2087), .dout(n2091));
    jxor g0535(.dinb(n1966), .dina(n2091), .dout(n2095));
    jxor g0536(.dinb(n20838), .dina(n2095), .dout(n2099));
    jxor g0537(.dinb(n1947), .dina(n2099), .dout(n2103));
    jxor g0538(.dinb(n19746), .dina(n2103), .dout(n2107));
    jxor g0539(.dinb(n1928), .dina(n18666), .dout(n2111));
    jxor g0540(.dinb(n18663), .dina(n2111), .dout(n2115));
    jxor g0541(.dinb(n1909), .dina(n17550), .dout(n2119));
    jxor g0542(.dinb(n17547), .dina(n2119), .dout(n2123));
    jxor g0543(.dinb(n1890), .dina(n16419), .dout(n2127));
    jxor g0544(.dinb(n16416), .dina(n2127), .dout(n2131));
    jnot g0545(.din(n2131), .dout(n2134));
    jxor g0546(.dinb(n1871), .dina(n2134), .dout(n2138));
    jxor g0547(.dinb(n13566), .dina(n2138), .dout(n2142));
    jxor g0548(.dinb(n1848), .dina(n13475), .dout(n2146));
    jxor g0549(.dinb(n11190), .dina(n2146), .dout(n2150));
    jand g0550(.dinb(G1gat), .dina(G494gat), .dout(n2154));
    jnot g0551(.din(n2154), .dout(n2157));
    jnot g0552(.din(n2142), .dout(n2160));
    jor g0553(.dinb(n1848), .dina(n2160), .dout(n2164));
    jor g0554(.dinb(n13373), .dina(n2146), .dout(n2168));
    jand g0555(.dinb(n13371), .dina(n2168), .dout(n2172));
    jand g0556(.dinb(G18gat), .dina(G477gat), .dout(n2176));
    jnot g0557(.din(n2176), .dout(n2179));
    jor g0558(.dinb(n1871), .dina(n2134), .dout(n2183));
    jxor g0559(.dinb(n1871), .dina(n15260), .dout(n2187));
    jor g0560(.dinb(n15167), .dina(n2187), .dout(n2191));
    jand g0561(.dinb(n15165), .dina(n2191), .dout(n2195));
    jand g0562(.dinb(G35gat), .dina(G460gat), .dout(n2199));
    jnot g0563(.din(n2199), .dout(n2202));
    jand g0564(.dinb(n1890), .dina(n16419), .dout(n2206));
    jand g0565(.dinb(n16416), .dina(n2127), .dout(n2210));
    jor g0566(.dinb(n16335), .dina(n2210), .dout(n2214));
    jand g0567(.dinb(G52gat), .dina(G443gat), .dout(n2218));
    jnot g0568(.din(n2218), .dout(n2221));
    jand g0569(.dinb(n1909), .dina(n17550), .dout(n2225));
    jand g0570(.dinb(n17547), .dina(n2119), .dout(n2229));
    jor g0571(.dinb(n17475), .dina(n2229), .dout(n2233));
    jand g0572(.dinb(G69gat), .dina(G426gat), .dout(n2237));
    jnot g0573(.din(n2237), .dout(n2240));
    jand g0574(.dinb(n1928), .dina(n18666), .dout(n2244));
    jand g0575(.dinb(n18663), .dina(n2111), .dout(n2248));
    jor g0576(.dinb(n18600), .dina(n2248), .dout(n2252));
    jand g0577(.dinb(G86gat), .dina(G409gat), .dout(n2256));
    jnot g0578(.din(n2256), .dout(n2259));
    jand g0579(.dinb(n1947), .dina(n2099), .dout(n2263));
    jand g0580(.dinb(n19746), .dina(n2103), .dout(n2267));
    jor g0581(.dinb(n19692), .dina(n2267), .dout(n2271));
    jand g0582(.dinb(G103gat), .dina(G392gat), .dout(n2275));
    jnot g0583(.din(n2275), .dout(n2278));
    jand g0584(.dinb(n1966), .dina(n2091), .dout(n2282));
    jand g0585(.dinb(n20838), .dina(n2095), .dout(n2286));
    jor g0586(.dinb(n20790), .dina(n2286), .dout(n2290));
    jand g0587(.dinb(G120gat), .dina(G375gat), .dout(n2294));
    jnot g0588(.din(n2294), .dout(n2297));
    jand g0589(.dinb(n1985), .dina(n21996), .dout(n2301));
    jand g0590(.dinb(n21993), .dina(n2087), .dout(n2305));
    jor g0591(.dinb(n21951), .dina(n2305), .dout(n2309));
    jand g0592(.dinb(G137gat), .dina(G358gat), .dout(n2313));
    jnot g0593(.din(n2313), .dout(n2316));
    jand g0594(.dinb(n2004), .dina(n23172), .dout(n2320));
    jand g0595(.dinb(n23169), .dina(n2079), .dout(n2324));
    jor g0596(.dinb(n23136), .dina(n2324), .dout(n2328));
    jand g0597(.dinb(G154gat), .dina(G341gat), .dout(n2332));
    jnot g0598(.din(n2332), .dout(n2335));
    jand g0599(.dinb(n2029), .dina(n24342), .dout(n2339));
    jand g0600(.dinb(n24333), .dina(n2071), .dout(n2343));
    jor g0601(.dinb(n24309), .dina(n2343), .dout(n2347));
    jand g0602(.dinb(G171gat), .dina(G324gat), .dout(n2351));
    jnot g0603(.din(n2351), .dout(n2354));
    jor g0604(.dinb(n25502), .dina(n2059), .dout(n2358));
    jand g0605(.dinb(n25497), .dina(n2063), .dout(n2362));
    jnot g0606(.din(n2362), .dout(n2365));
    jand g0607(.dinb(n25488), .dina(n2365), .dout(n2369));
    jnot g0608(.din(n2369), .dout(n2372));
    jand g0609(.dinb(G188gat), .dina(G307gat), .dout(n2376));
    jnot g0610(.din(n2376), .dout(n2379));
    jand g0611(.dinb(G222gat), .dina(G290gat), .dout(n2383));
    jand g0612(.dinb(n2051), .dina(n2383), .dout(n2387));
    jnot g0613(.din(n2387), .dout(n2390));
    jand g0614(.dinb(G222gat), .dina(G273gat), .dout(n2394));
    jor g0615(.dinb(n2040), .dina(n2394), .dout(n2398));
    jand g0616(.dinb(n2390), .dina(n26661), .dout(n2402));
    jxor g0617(.dinb(n26669), .dina(n2402), .dout(n2406));
    jxor g0618(.dinb(n26658), .dina(n2406), .dout(n2410));
    jxor g0619(.dinb(n2372), .dina(n25482), .dout(n2414));
    jxor g0620(.dinb(n25473), .dina(n2414), .dout(n2418));
    jxor g0621(.dinb(n2347), .dina(n24306), .dout(n2422));
    jxor g0622(.dinb(n24303), .dina(n2422), .dout(n2426));
    jxor g0623(.dinb(n2328), .dina(n23133), .dout(n2430));
    jxor g0624(.dinb(n23130), .dina(n2430), .dout(n2434));
    jxor g0625(.dinb(n2309), .dina(n21948), .dout(n2438));
    jxor g0626(.dinb(n21945), .dina(n2438), .dout(n2442));
    jxor g0627(.dinb(n2290), .dina(n2442), .dout(n2446));
    jxor g0628(.dinb(n20787), .dina(n2446), .dout(n2450));
    jxor g0629(.dinb(n2271), .dina(n2450), .dout(n2454));
    jxor g0630(.dinb(n19689), .dina(n2454), .dout(n2458));
    jxor g0631(.dinb(n2252), .dina(n18597), .dout(n2462));
    jxor g0632(.dinb(n18594), .dina(n2462), .dout(n2466));
    jxor g0633(.dinb(n2233), .dina(n17472), .dout(n2470));
    jxor g0634(.dinb(n17469), .dina(n2470), .dout(n2474));
    jxor g0635(.dinb(n2214), .dina(n16332), .dout(n2478));
    jxor g0636(.dinb(n16329), .dina(n2478), .dout(n2482));
    jnot g0637(.din(n2482), .dout(n2485));
    jxor g0638(.dinb(n2195), .dina(n2485), .dout(n2489));
    jxor g0639(.dinb(n13368), .dina(n2489), .dout(n2493));
    jxor g0640(.dinb(n2172), .dina(n13268), .dout(n2497));
    jxor g0641(.dinb(n11298), .dina(n2497), .dout(n2501));
    jand g0642(.dinb(G1gat), .dina(G511gat), .dout(n2505));
    jnot g0643(.din(n2505), .dout(n2508));
    jnot g0644(.din(n2493), .dout(n2511));
    jor g0645(.dinb(n2172), .dina(n2511), .dout(n2515));
    jor g0646(.dinb(n13157), .dina(n2497), .dout(n2519));
    jand g0647(.dinb(n13155), .dina(n2519), .dout(n2523));
    jand g0648(.dinb(G18gat), .dina(G494gat), .dout(n2527));
    jnot g0649(.din(n2527), .dout(n2530));
    jor g0650(.dinb(n2195), .dina(n2485), .dout(n2534));
    jxor g0651(.dinb(n2195), .dina(n15161), .dout(n2538));
    jor g0652(.dinb(n15059), .dina(n2538), .dout(n2542));
    jand g0653(.dinb(n15057), .dina(n2542), .dout(n2546));
    jand g0654(.dinb(G35gat), .dina(G477gat), .dout(n2550));
    jnot g0655(.din(n2550), .dout(n2553));
    jand g0656(.dinb(n2214), .dina(n16332), .dout(n2557));
    jand g0657(.dinb(n16329), .dina(n2478), .dout(n2561));
    jor g0658(.dinb(n16239), .dina(n2561), .dout(n2565));
    jand g0659(.dinb(G52gat), .dina(G460gat), .dout(n2569));
    jnot g0660(.din(n2569), .dout(n2572));
    jand g0661(.dinb(n2233), .dina(n17472), .dout(n2576));
    jand g0662(.dinb(n17469), .dina(n2470), .dout(n2580));
    jor g0663(.dinb(n17388), .dina(n2580), .dout(n2584));
    jand g0664(.dinb(G69gat), .dina(G443gat), .dout(n2588));
    jnot g0665(.din(n2588), .dout(n2591));
    jand g0666(.dinb(n2252), .dina(n18597), .dout(n2595));
    jand g0667(.dinb(n18594), .dina(n2462), .dout(n2599));
    jor g0668(.dinb(n18522), .dina(n2599), .dout(n2603));
    jand g0669(.dinb(G86gat), .dina(G426gat), .dout(n2607));
    jnot g0670(.din(n2607), .dout(n2610));
    jand g0671(.dinb(n2271), .dina(n2450), .dout(n2614));
    jand g0672(.dinb(n19689), .dina(n2454), .dout(n2618));
    jor g0673(.dinb(n19626), .dina(n2618), .dout(n2622));
    jand g0674(.dinb(G103gat), .dina(G409gat), .dout(n2626));
    jnot g0675(.din(n2626), .dout(n2629));
    jand g0676(.dinb(n2290), .dina(n2442), .dout(n2633));
    jand g0677(.dinb(n20787), .dina(n2446), .dout(n2637));
    jor g0678(.dinb(n20730), .dina(n2637), .dout(n2641));
    jand g0679(.dinb(G120gat), .dina(G392gat), .dout(n2645));
    jnot g0680(.din(n2645), .dout(n2648));
    jand g0681(.dinb(n2309), .dina(n21948), .dout(n2652));
    jand g0682(.dinb(n21945), .dina(n2438), .dout(n2656));
    jor g0683(.dinb(n21894), .dina(n2656), .dout(n2660));
    jand g0684(.dinb(G137gat), .dina(G375gat), .dout(n2664));
    jnot g0685(.din(n2664), .dout(n2667));
    jand g0686(.dinb(n2328), .dina(n23133), .dout(n2671));
    jand g0687(.dinb(n23130), .dina(n2430), .dout(n2675));
    jor g0688(.dinb(n23088), .dina(n2675), .dout(n2679));
    jand g0689(.dinb(G154gat), .dina(G358gat), .dout(n2683));
    jnot g0690(.din(n2683), .dout(n2686));
    jand g0691(.dinb(n2347), .dina(n24306), .dout(n2690));
    jand g0692(.dinb(n24303), .dina(n2422), .dout(n2694));
    jor g0693(.dinb(n24270), .dina(n2694), .dout(n2698));
    jand g0694(.dinb(G171gat), .dina(G341gat), .dout(n2702));
    jnot g0695(.din(n2702), .dout(n2705));
    jand g0696(.dinb(n2372), .dina(n25482), .dout(n2709));
    jand g0697(.dinb(n25473), .dina(n2414), .dout(n2713));
    jor g0698(.dinb(n25449), .dina(n2713), .dout(n2717));
    jand g0699(.dinb(G188gat), .dina(G324gat), .dout(n2721));
    jnot g0700(.din(n2721), .dout(n2724));
    jor g0701(.dinb(n26663), .dina(n2402), .dout(n2728));
    jand g0702(.dinb(n26658), .dina(n2406), .dout(n2732));
    jnot g0703(.din(n2732), .dout(n2735));
    jand g0704(.dinb(n26649), .dina(n2735), .dout(n2739));
    jnot g0705(.din(n2739), .dout(n2742));
    jand g0706(.dinb(G205gat), .dina(G307gat), .dout(n2746));
    jnot g0707(.din(n2746), .dout(n2749));
    jand g0708(.dinb(G239gat), .dina(G290gat), .dout(n2753));
    jand g0709(.dinb(n2394), .dina(n2753), .dout(n2757));
    jnot g0710(.din(n2757), .dout(n2760));
    jand g0711(.dinb(G239gat), .dina(G273gat), .dout(n2764));
    jor g0712(.dinb(n2383), .dina(n2764), .dout(n2768));
    jand g0713(.dinb(n2760), .dina(n27855), .dout(n2772));
    jxor g0714(.dinb(n27863), .dina(n2772), .dout(n2776));
    jxor g0715(.dinb(n27852), .dina(n2776), .dout(n2780));
    jxor g0716(.dinb(n2742), .dina(n26643), .dout(n2784));
    jxor g0717(.dinb(n26634), .dina(n2784), .dout(n2788));
    jxor g0718(.dinb(n2717), .dina(n25446), .dout(n2792));
    jxor g0719(.dinb(n25443), .dina(n2792), .dout(n2796));
    jxor g0720(.dinb(n2698), .dina(n24267), .dout(n2800));
    jxor g0721(.dinb(n24264), .dina(n2800), .dout(n2804));
    jxor g0722(.dinb(n2679), .dina(n23085), .dout(n2808));
    jxor g0723(.dinb(n23082), .dina(n2808), .dout(n2812));
    jxor g0724(.dinb(n2660), .dina(n21891), .dout(n2816));
    jxor g0725(.dinb(n21888), .dina(n2816), .dout(n2820));
    jxor g0726(.dinb(n2641), .dina(n2820), .dout(n2824));
    jxor g0727(.dinb(n20727), .dina(n2824), .dout(n2828));
    jxor g0728(.dinb(n2622), .dina(n2828), .dout(n2832));
    jxor g0729(.dinb(n19623), .dina(n2832), .dout(n2836));
    jxor g0730(.dinb(n2603), .dina(n18519), .dout(n2840));
    jxor g0731(.dinb(n18516), .dina(n2840), .dout(n2844));
    jxor g0732(.dinb(n2584), .dina(n17385), .dout(n2848));
    jxor g0733(.dinb(n17382), .dina(n2848), .dout(n2852));
    jxor g0734(.dinb(n2565), .dina(n16236), .dout(n2856));
    jxor g0735(.dinb(n16233), .dina(n2856), .dout(n2860));
    jnot g0736(.din(n2860), .dout(n2863));
    jxor g0737(.dinb(n2546), .dina(n2863), .dout(n2867));
    jxor g0738(.dinb(n13152), .dina(n2867), .dout(n2871));
    jxor g0739(.dinb(n2523), .dina(n13043), .dout(n2875));
    jxor g0740(.dinb(n11415), .dina(n2875), .dout(n2879));
    jand g0741(.dinb(G1gat), .dina(G528gat), .dout(n2883));
    jnot g0742(.din(n2883), .dout(n2886));
    jnot g0743(.din(n2871), .dout(n2889));
    jor g0744(.dinb(n2523), .dina(n2889), .dout(n2893));
    jor g0745(.dinb(n12923), .dina(n2875), .dout(n2897));
    jand g0746(.dinb(n12921), .dina(n2897), .dout(n2901));
    jand g0747(.dinb(G18gat), .dina(G511gat), .dout(n2905));
    jor g0748(.dinb(n2546), .dina(n2863), .dout(n2909));
    jxor g0749(.dinb(n2546), .dina(n15053), .dout(n2913));
    jor g0750(.dinb(n14942), .dina(n2913), .dout(n2917));
    jand g0751(.dinb(n14940), .dina(n2917), .dout(n2921));
    jand g0752(.dinb(G35gat), .dina(G494gat), .dout(n2925));
    jnot g0753(.din(n2925), .dout(n2928));
    jand g0754(.dinb(n2565), .dina(n16236), .dout(n2932));
    jand g0755(.dinb(n16233), .dina(n2856), .dout(n2936));
    jor g0756(.dinb(n16134), .dina(n2936), .dout(n2940));
    jand g0757(.dinb(G52gat), .dina(G477gat), .dout(n2944));
    jnot g0758(.din(n2944), .dout(n2947));
    jand g0759(.dinb(n2584), .dina(n17385), .dout(n2951));
    jand g0760(.dinb(n17382), .dina(n2848), .dout(n2955));
    jor g0761(.dinb(n17292), .dina(n2955), .dout(n2959));
    jand g0762(.dinb(G69gat), .dina(G460gat), .dout(n2963));
    jnot g0763(.din(n2963), .dout(n2966));
    jand g0764(.dinb(n2603), .dina(n18519), .dout(n2970));
    jand g0765(.dinb(n18516), .dina(n2840), .dout(n2974));
    jor g0766(.dinb(n18435), .dina(n2974), .dout(n2978));
    jand g0767(.dinb(G86gat), .dina(G443gat), .dout(n2982));
    jnot g0768(.din(n2982), .dout(n2985));
    jand g0769(.dinb(n2622), .dina(n2828), .dout(n2989));
    jand g0770(.dinb(n19623), .dina(n2832), .dout(n2993));
    jor g0771(.dinb(n19551), .dina(n2993), .dout(n2997));
    jand g0772(.dinb(G103gat), .dina(G426gat), .dout(n3001));
    jnot g0773(.din(n3001), .dout(n3004));
    jand g0774(.dinb(n2641), .dina(n2820), .dout(n3008));
    jand g0775(.dinb(n20727), .dina(n2824), .dout(n3012));
    jor g0776(.dinb(n20661), .dina(n3012), .dout(n3016));
    jand g0777(.dinb(G120gat), .dina(G409gat), .dout(n3020));
    jnot g0778(.din(n3020), .dout(n3023));
    jand g0779(.dinb(n2660), .dina(n21891), .dout(n3027));
    jand g0780(.dinb(n21888), .dina(n2816), .dout(n3031));
    jor g0781(.dinb(n21828), .dina(n3031), .dout(n3035));
    jand g0782(.dinb(G137gat), .dina(G392gat), .dout(n3039));
    jnot g0783(.din(n3039), .dout(n3042));
    jand g0784(.dinb(n2679), .dina(n23085), .dout(n3046));
    jand g0785(.dinb(n23082), .dina(n2808), .dout(n3050));
    jor g0786(.dinb(n23031), .dina(n3050), .dout(n3054));
    jand g0787(.dinb(G154gat), .dina(G375gat), .dout(n3058));
    jnot g0788(.din(n3058), .dout(n3061));
    jand g0789(.dinb(n2698), .dina(n24267), .dout(n3065));
    jand g0790(.dinb(n24264), .dina(n2800), .dout(n3069));
    jor g0791(.dinb(n24222), .dina(n3069), .dout(n3073));
    jand g0792(.dinb(G171gat), .dina(G358gat), .dout(n3077));
    jnot g0793(.din(n3077), .dout(n3080));
    jand g0794(.dinb(n2717), .dina(n25446), .dout(n3084));
    jand g0795(.dinb(n25443), .dina(n2792), .dout(n3088));
    jor g0796(.dinb(n25410), .dina(n3088), .dout(n3092));
    jand g0797(.dinb(G188gat), .dina(G341gat), .dout(n3096));
    jnot g0798(.din(n3096), .dout(n3099));
    jand g0799(.dinb(n2742), .dina(n26643), .dout(n3103));
    jand g0800(.dinb(n26634), .dina(n2784), .dout(n3107));
    jor g0801(.dinb(n26610), .dina(n3107), .dout(n3111));
    jand g0802(.dinb(G205gat), .dina(G324gat), .dout(n3115));
    jnot g0803(.din(n3115), .dout(n3118));
    jor g0804(.dinb(n27857), .dina(n2772), .dout(n3122));
    jand g0805(.dinb(n27852), .dina(n2776), .dout(n3126));
    jnot g0806(.din(n3126), .dout(n3129));
    jand g0807(.dinb(n27843), .dina(n3129), .dout(n3133));
    jnot g0808(.din(n3133), .dout(n3136));
    jand g0809(.dinb(G222gat), .dina(G307gat), .dout(n3140));
    jnot g0810(.din(n3140), .dout(n3143));
    jand g0811(.dinb(G256gat), .dina(G273gat), .dout(n3147));
    jxor g0812(.dinb(n2753), .dina(n3147), .dout(n3151));
    jor g0813(.dinb(n2757), .dina(n3151), .dout(n3155));
    jor g0814(.dinb(n2760), .dina(n31535), .dout(n3159));
    jand g0815(.dinb(n31533), .dina(n3159), .dout(n3163));
    jxor g0816(.dinb(n31548), .dina(n3163), .dout(n3167));
    jxor g0817(.dinb(n3136), .dina(n27837), .dout(n3171));
    jxor g0818(.dinb(n27828), .dina(n3171), .dout(n3175));
    jxor g0819(.dinb(n3111), .dina(n26607), .dout(n3179));
    jxor g0820(.dinb(n26604), .dina(n3179), .dout(n3183));
    jxor g0821(.dinb(n3092), .dina(n25407), .dout(n3187));
    jxor g0822(.dinb(n25404), .dina(n3187), .dout(n3191));
    jxor g0823(.dinb(n3073), .dina(n24219), .dout(n3195));
    jxor g0824(.dinb(n24216), .dina(n3195), .dout(n3199));
    jxor g0825(.dinb(n3054), .dina(n23028), .dout(n3203));
    jxor g0826(.dinb(n23025), .dina(n3203), .dout(n3207));
    jxor g0827(.dinb(n3035), .dina(n21825), .dout(n3211));
    jxor g0828(.dinb(n21822), .dina(n3211), .dout(n3215));
    jxor g0829(.dinb(n3016), .dina(n3215), .dout(n3219));
    jxor g0830(.dinb(n20658), .dina(n3219), .dout(n3223));
    jxor g0831(.dinb(n2997), .dina(n3223), .dout(n3227));
    jxor g0832(.dinb(n19548), .dina(n3227), .dout(n3231));
    jxor g0833(.dinb(n2978), .dina(n18432), .dout(n3235));
    jxor g0834(.dinb(n18429), .dina(n3235), .dout(n3239));
    jxor g0835(.dinb(n2959), .dina(n17289), .dout(n3243));
    jxor g0836(.dinb(n17286), .dina(n3243), .dout(n3247));
    jxor g0837(.dinb(n2940), .dina(n16130), .dout(n3251));
    jxor g0838(.dinb(n14937), .dina(n3251), .dout(n3255));
    jxor g0839(.dinb(n2921), .dina(n14828), .dout(n3259));
    jxor g0840(.dinb(n14826), .dina(n3259), .dout(n3263));
    jxor g0841(.dinb(n2901), .dina(n12917), .dout(n3267));
    jxor g0842(.dinb(n11541), .dina(n3267), .dout(n3271));
    jnot g0843(.din(n3263), .dout(n3274));
    jor g0844(.dinb(n2901), .dina(n3274), .dout(n3278));
    jor g0845(.dinb(n12788), .dina(n3267), .dout(n3282));
    jand g0846(.dinb(n12786), .dina(n3282), .dout(n3286));
    jand g0847(.dinb(G18gat), .dina(G528gat), .dout(n3290));
    jnot g0848(.din(n3255), .dout(n3293));
    jor g0849(.dinb(n2921), .dina(n3293), .dout(n3297));
    jor g0850(.dinb(n14826), .dina(n3259), .dout(n3301));
    jand g0851(.dinb(n14706), .dina(n3301), .dout(n3305));
    jand g0852(.dinb(G35gat), .dina(G511gat), .dout(n3309));
    jand g0853(.dinb(n2940), .dina(n16127), .dout(n3313));
    jnot g0854(.din(n3313), .dout(n3316));
    jnot g0855(.din(n3247), .dout(n3319));
    jxor g0856(.dinb(n2940), .dina(n3319), .dout(n3323));
    jor g0857(.dinb(n16016), .dina(n3323), .dout(n3327));
    jand g0858(.dinb(n3316), .dina(n3327), .dout(n3331));
    jand g0859(.dinb(G52gat), .dina(G494gat), .dout(n3335));
    jnot g0860(.din(n3335), .dout(n3338));
    jand g0861(.dinb(n2959), .dina(n17289), .dout(n3342));
    jand g0862(.dinb(n17286), .dina(n3243), .dout(n3346));
    jor g0863(.dinb(n17187), .dina(n3346), .dout(n3350));
    jand g0864(.dinb(G69gat), .dina(G477gat), .dout(n3354));
    jnot g0865(.din(n3354), .dout(n3357));
    jand g0866(.dinb(n2978), .dina(n18432), .dout(n3361));
    jand g0867(.dinb(n18429), .dina(n3235), .dout(n3365));
    jor g0868(.dinb(n18339), .dina(n3365), .dout(n3369));
    jand g0869(.dinb(G86gat), .dina(G460gat), .dout(n3373));
    jnot g0870(.din(n3373), .dout(n3376));
    jand g0871(.dinb(n2997), .dina(n3223), .dout(n3380));
    jand g0872(.dinb(n19548), .dina(n3227), .dout(n3384));
    jor g0873(.dinb(n19467), .dina(n3384), .dout(n3388));
    jand g0874(.dinb(G103gat), .dina(G443gat), .dout(n3392));
    jnot g0875(.din(n3392), .dout(n3395));
    jand g0876(.dinb(n3016), .dina(n3215), .dout(n3399));
    jand g0877(.dinb(n20658), .dina(n3219), .dout(n3403));
    jor g0878(.dinb(n20583), .dina(n3403), .dout(n3407));
    jand g0879(.dinb(G120gat), .dina(G426gat), .dout(n3411));
    jnot g0880(.din(n3411), .dout(n3414));
    jand g0881(.dinb(n3035), .dina(n21825), .dout(n3418));
    jand g0882(.dinb(n21822), .dina(n3211), .dout(n3422));
    jor g0883(.dinb(n21753), .dina(n3422), .dout(n3426));
    jand g0884(.dinb(G137gat), .dina(G409gat), .dout(n3430));
    jnot g0885(.din(n3430), .dout(n3433));
    jand g0886(.dinb(n3054), .dina(n23028), .dout(n3437));
    jand g0887(.dinb(n23025), .dina(n3203), .dout(n3441));
    jor g0888(.dinb(n22965), .dina(n3441), .dout(n3445));
    jand g0889(.dinb(G154gat), .dina(G392gat), .dout(n3449));
    jnot g0890(.din(n3449), .dout(n3452));
    jand g0891(.dinb(n3073), .dina(n24219), .dout(n3456));
    jand g0892(.dinb(n24216), .dina(n3195), .dout(n3460));
    jor g0893(.dinb(n24165), .dina(n3460), .dout(n3464));
    jand g0894(.dinb(G171gat), .dina(G375gat), .dout(n3468));
    jnot g0895(.din(n3468), .dout(n3471));
    jand g0896(.dinb(n3092), .dina(n25407), .dout(n3475));
    jand g0897(.dinb(n25404), .dina(n3187), .dout(n3479));
    jor g0898(.dinb(n25362), .dina(n3479), .dout(n3483));
    jand g0899(.dinb(G188gat), .dina(G358gat), .dout(n3487));
    jnot g0900(.din(n3487), .dout(n3490));
    jand g0901(.dinb(n3111), .dina(n26607), .dout(n3494));
    jand g0902(.dinb(n26604), .dina(n3179), .dout(n3498));
    jor g0903(.dinb(n26571), .dina(n3498), .dout(n3502));
    jand g0904(.dinb(G205gat), .dina(G341gat), .dout(n3506));
    jnot g0905(.din(n3506), .dout(n3509));
    jand g0906(.dinb(n3136), .dina(n27837), .dout(n3513));
    jand g0907(.dinb(n27828), .dina(n3171), .dout(n3517));
    jor g0908(.dinb(n27804), .dina(n3517), .dout(n3521));
    jand g0909(.dinb(G222gat), .dina(G324gat), .dout(n3525));
    jnot g0910(.din(n3525), .dout(n3528));
    jand g0911(.dinb(n31548), .dina(n3163), .dout(n3532));
    jnot g0912(.din(n3532), .dout(n3535));
    jand g0913(.dinb(n31523), .dina(n3535), .dout(n3539));
    jnot g0914(.din(n3539), .dout(n3542));
    jnot g0915(.din(n2764), .dout(n3545));
    jand g0916(.dinb(G256gat), .dina(G290gat), .dout(n3549));
    jand g0917(.dinb(n3545), .dina(n31521), .dout(n3553));
    jnot g0918(.din(n3553), .dout(n3556));
    jand g0919(.dinb(G239gat), .dina(G307gat), .dout(n3560));
    jxor g0920(.dinb(n3556), .dina(n31509), .dout(n3564));
    jxor g0921(.dinb(n3542), .dina(n31500), .dout(n3568));
    jxor g0922(.dinb(n31488), .dina(n3568), .dout(n3572));
    jxor g0923(.dinb(n3521), .dina(n27801), .dout(n3576));
    jxor g0924(.dinb(n27798), .dina(n3576), .dout(n3580));
    jxor g0925(.dinb(n3502), .dina(n26568), .dout(n3584));
    jxor g0926(.dinb(n26565), .dina(n3584), .dout(n3588));
    jxor g0927(.dinb(n3483), .dina(n25359), .dout(n3592));
    jxor g0928(.dinb(n25356), .dina(n3592), .dout(n3596));
    jxor g0929(.dinb(n3464), .dina(n24162), .dout(n3600));
    jxor g0930(.dinb(n24159), .dina(n3600), .dout(n3604));
    jxor g0931(.dinb(n3445), .dina(n22962), .dout(n3608));
    jxor g0932(.dinb(n22959), .dina(n3608), .dout(n3612));
    jxor g0933(.dinb(n3426), .dina(n21750), .dout(n3616));
    jxor g0934(.dinb(n21747), .dina(n3616), .dout(n3620));
    jxor g0935(.dinb(n3407), .dina(n3620), .dout(n3624));
    jxor g0936(.dinb(n20580), .dina(n3624), .dout(n3628));
    jxor g0937(.dinb(n3388), .dina(n3628), .dout(n3632));
    jxor g0938(.dinb(n19464), .dina(n3632), .dout(n3636));
    jxor g0939(.dinb(n3369), .dina(n18336), .dout(n3640));
    jxor g0940(.dinb(n18333), .dina(n3640), .dout(n3644));
    jxor g0941(.dinb(n3350), .dina(n17184), .dout(n3648));
    jxor g0942(.dinb(n17181), .dina(n3648), .dout(n3652));
    jxor g0943(.dinb(n3331), .dina(n16013), .dout(n3656));
    jxor g0944(.dinb(n16011), .dina(n3656), .dout(n3660));
    jnot g0945(.din(n3660), .dout(n3663));
    jxor g0946(.dinb(n3305), .dina(n3663), .dout(n3667));
    jxor g0947(.dinb(n14700), .dina(n3667), .dout(n3671));
    jxor g0948(.dinb(n3286), .dina(n12783), .dout(n3675));
    jand g0949(.dinb(n3286), .dina(n12783), .dout(n3679));
    jor g0950(.dinb(n3305), .dina(n3663), .dout(n3683));
    jxor g0951(.dinb(n3305), .dina(n14702), .dout(n3687));
    jor g0952(.dinb(n14700), .dina(n3687), .dout(n3691));
    jand g0953(.dinb(n14571), .dina(n3691), .dout(n3695));
    jand g0954(.dinb(G35gat), .dina(G528gat), .dout(n3699));
    jnot g0955(.din(n3652), .dout(n3702));
    jor g0956(.dinb(n3331), .dina(n3702), .dout(n3706));
    jor g0957(.dinb(n16011), .dina(n3656), .dout(n3710));
    jand g0958(.dinb(n15891), .dina(n3710), .dout(n3714));
    jand g0959(.dinb(G52gat), .dina(G511gat), .dout(n3718));
    jand g0960(.dinb(n3350), .dina(n17184), .dout(n3722));
    jand g0961(.dinb(n17181), .dina(n3648), .dout(n3726));
    jor g0962(.dinb(n17073), .dina(n3726), .dout(n3730));
    jand g0963(.dinb(G69gat), .dina(G494gat), .dout(n3734));
    jnot g0964(.din(n3734), .dout(n3737));
    jand g0965(.dinb(n3369), .dina(n18336), .dout(n3741));
    jand g0966(.dinb(n18333), .dina(n3640), .dout(n3745));
    jor g0967(.dinb(n18234), .dina(n3745), .dout(n3749));
    jand g0968(.dinb(G86gat), .dina(G477gat), .dout(n3753));
    jnot g0969(.din(n3753), .dout(n3756));
    jand g0970(.dinb(n3388), .dina(n3628), .dout(n3760));
    jand g0971(.dinb(n19464), .dina(n3632), .dout(n3764));
    jor g0972(.dinb(n19374), .dina(n3764), .dout(n3768));
    jand g0973(.dinb(G103gat), .dina(G460gat), .dout(n3772));
    jnot g0974(.din(n3772), .dout(n3775));
    jand g0975(.dinb(n3407), .dina(n3620), .dout(n3779));
    jand g0976(.dinb(n20580), .dina(n3624), .dout(n3783));
    jor g0977(.dinb(n20496), .dina(n3783), .dout(n3787));
    jand g0978(.dinb(G120gat), .dina(G443gat), .dout(n3791));
    jnot g0979(.din(n3791), .dout(n3794));
    jand g0980(.dinb(n3426), .dina(n21750), .dout(n3798));
    jand g0981(.dinb(n21747), .dina(n3616), .dout(n3802));
    jor g0982(.dinb(n21669), .dina(n3802), .dout(n3806));
    jand g0983(.dinb(G137gat), .dina(G426gat), .dout(n3810));
    jnot g0984(.din(n3810), .dout(n3813));
    jand g0985(.dinb(n3445), .dina(n22962), .dout(n3817));
    jand g0986(.dinb(n22959), .dina(n3608), .dout(n3821));
    jor g0987(.dinb(n22890), .dina(n3821), .dout(n3825));
    jand g0988(.dinb(G154gat), .dina(G409gat), .dout(n3829));
    jnot g0989(.din(n3829), .dout(n3832));
    jand g0990(.dinb(n3464), .dina(n24162), .dout(n3836));
    jand g0991(.dinb(n24159), .dina(n3600), .dout(n3840));
    jor g0992(.dinb(n24099), .dina(n3840), .dout(n3844));
    jand g0993(.dinb(G171gat), .dina(G392gat), .dout(n3848));
    jnot g0994(.din(n3848), .dout(n3851));
    jand g0995(.dinb(n3483), .dina(n25359), .dout(n3855));
    jand g0996(.dinb(n25356), .dina(n3592), .dout(n3859));
    jor g0997(.dinb(n25305), .dina(n3859), .dout(n3863));
    jand g0998(.dinb(G188gat), .dina(G375gat), .dout(n3867));
    jnot g0999(.din(n3867), .dout(n3870));
    jand g1000(.dinb(n3502), .dina(n26568), .dout(n3874));
    jand g1001(.dinb(n26565), .dina(n3584), .dout(n3878));
    jor g1002(.dinb(n26523), .dina(n3878), .dout(n3882));
    jand g1003(.dinb(G205gat), .dina(G358gat), .dout(n3886));
    jnot g1004(.din(n3886), .dout(n3889));
    jand g1005(.dinb(n3521), .dina(n27801), .dout(n3893));
    jand g1006(.dinb(n27798), .dina(n3576), .dout(n3897));
    jor g1007(.dinb(n27765), .dina(n3897), .dout(n3901));
    jand g1008(.dinb(G222gat), .dina(G341gat), .dout(n3905));
    jnot g1009(.din(n3905), .dout(n3908));
    jand g1010(.dinb(n3542), .dina(n31500), .dout(n3912));
    jand g1011(.dinb(n31488), .dina(n3568), .dout(n3916));
    jor g1012(.dinb(n31464), .dina(n3916), .dout(n3920));
    jand g1013(.dinb(G239gat), .dina(G324gat), .dout(n3924));
    jand g1014(.dinb(G256gat), .dina(G307gat), .dout(n3928));
    jor g1015(.dinb(n3556), .dina(n31509), .dout(n3932));
    jand g1016(.dinb(n31511), .dina(n3932), .dout(n3936));
    jxor g1017(.dinb(n31440), .dina(n3936), .dout(n3940));
    jnot g1018(.din(n3940), .dout(n3943));
    jxor g1019(.dinb(n31461), .dina(n3943), .dout(n3947));
    jxor g1020(.dinb(n3920), .dina(n31425), .dout(n3951));
    jxor g1021(.dinb(n31416), .dina(n3951), .dout(n3955));
    jxor g1022(.dinb(n3901), .dina(n27762), .dout(n3959));
    jxor g1023(.dinb(n27759), .dina(n3959), .dout(n3963));
    jxor g1024(.dinb(n3882), .dina(n26520), .dout(n3967));
    jxor g1025(.dinb(n26517), .dina(n3967), .dout(n3971));
    jxor g1026(.dinb(n3863), .dina(n25302), .dout(n3975));
    jxor g1027(.dinb(n25299), .dina(n3975), .dout(n3979));
    jxor g1028(.dinb(n3844), .dina(n24096), .dout(n3983));
    jxor g1029(.dinb(n24093), .dina(n3983), .dout(n3987));
    jxor g1030(.dinb(n3825), .dina(n22887), .dout(n3991));
    jxor g1031(.dinb(n22884), .dina(n3991), .dout(n3995));
    jxor g1032(.dinb(n3806), .dina(n21666), .dout(n3999));
    jxor g1033(.dinb(n21663), .dina(n3999), .dout(n4003));
    jxor g1034(.dinb(n3787), .dina(n4003), .dout(n4007));
    jxor g1035(.dinb(n20493), .dina(n4007), .dout(n4011));
    jxor g1036(.dinb(n3768), .dina(n4011), .dout(n4015));
    jxor g1037(.dinb(n19371), .dina(n4015), .dout(n4019));
    jxor g1038(.dinb(n3749), .dina(n18231), .dout(n4023));
    jxor g1039(.dinb(n18228), .dina(n4023), .dout(n4027));
    jxor g1040(.dinb(n3730), .dina(n17070), .dout(n4031));
    jnot g1041(.din(n4031), .dout(n4034));
    jxor g1042(.dinb(n17067), .dina(n4034), .dout(n4038));
    jxor g1043(.dinb(n3714), .dina(n4038), .dout(n4042));
    jxor g1044(.dinb(n15885), .dina(n4042), .dout(n4046));
    jxor g1045(.dinb(n3695), .dina(n14567), .dout(n4050));
    jnot g1046(.din(n4050), .dout(n4053));
    jxor g1047(.dinb(n12779), .dina(n4053), .dout(n4057));
    jnot g1048(.din(n4046), .dout(n4060));
    jor g1049(.dinb(n3695), .dina(n4060), .dout(n4064));
    jor g1050(.dinb(n3679), .dina(n4050), .dout(n4068));
    jand g1051(.dinb(n12777), .dina(n4068), .dout(n4072));
    jnot g1052(.din(n4038), .dout(n4075));
    jor g1053(.dinb(n15887), .dina(n4075), .dout(n4079));
    jor g1054(.dinb(n15885), .dina(n4042), .dout(n4083));
    jand g1055(.dinb(n4079), .dina(n4083), .dout(n4087));
    jand g1056(.dinb(G52gat), .dina(G528gat), .dout(n4091));
    jand g1057(.dinb(n3730), .dina(n17070), .dout(n4095));
    jnot g1058(.din(n4095), .dout(n4098));
    jor g1059(.dinb(n17067), .dina(n4034), .dout(n4102));
    jand g1060(.dinb(n16944), .dina(n4102), .dout(n4106));
    jand g1061(.dinb(G69gat), .dina(G511gat), .dout(n4110));
    jnot g1062(.din(n4110), .dout(n4113));
    jand g1063(.dinb(n3749), .dina(n18231), .dout(n4117));
    jand g1064(.dinb(n18228), .dina(n4023), .dout(n4121));
    jor g1065(.dinb(n18120), .dina(n4121), .dout(n4125));
    jand g1066(.dinb(G86gat), .dina(G494gat), .dout(n4129));
    jnot g1067(.din(n4129), .dout(n4132));
    jand g1068(.dinb(n3768), .dina(n4011), .dout(n4136));
    jand g1069(.dinb(n19371), .dina(n4015), .dout(n4140));
    jor g1070(.dinb(n19272), .dina(n4140), .dout(n4144));
    jand g1071(.dinb(G103gat), .dina(G477gat), .dout(n4148));
    jnot g1072(.din(n4148), .dout(n4151));
    jand g1073(.dinb(n3787), .dina(n4003), .dout(n4155));
    jand g1074(.dinb(n20493), .dina(n4007), .dout(n4159));
    jor g1075(.dinb(n20400), .dina(n4159), .dout(n4163));
    jand g1076(.dinb(G120gat), .dina(G460gat), .dout(n4167));
    jnot g1077(.din(n4167), .dout(n4170));
    jand g1078(.dinb(n3806), .dina(n21666), .dout(n4174));
    jand g1079(.dinb(n21663), .dina(n3999), .dout(n4178));
    jor g1080(.dinb(n21576), .dina(n4178), .dout(n4182));
    jand g1081(.dinb(G137gat), .dina(G443gat), .dout(n4186));
    jnot g1082(.din(n4186), .dout(n4189));
    jand g1083(.dinb(n3825), .dina(n22887), .dout(n4193));
    jand g1084(.dinb(n22884), .dina(n3991), .dout(n4197));
    jor g1085(.dinb(n22806), .dina(n4197), .dout(n4201));
    jand g1086(.dinb(G154gat), .dina(G426gat), .dout(n4205));
    jnot g1087(.din(n4205), .dout(n4208));
    jand g1088(.dinb(n3844), .dina(n24096), .dout(n4212));
    jand g1089(.dinb(n24093), .dina(n3983), .dout(n4216));
    jor g1090(.dinb(n24024), .dina(n4216), .dout(n4220));
    jand g1091(.dinb(G171gat), .dina(G409gat), .dout(n4224));
    jnot g1092(.din(n4224), .dout(n4227));
    jand g1093(.dinb(n3863), .dina(n25302), .dout(n4231));
    jand g1094(.dinb(n25299), .dina(n3975), .dout(n4235));
    jor g1095(.dinb(n25239), .dina(n4235), .dout(n4239));
    jand g1096(.dinb(G188gat), .dina(G392gat), .dout(n4243));
    jnot g1097(.din(n4243), .dout(n4246));
    jand g1098(.dinb(n3882), .dina(n26520), .dout(n4250));
    jand g1099(.dinb(n26517), .dina(n3967), .dout(n4254));
    jor g1100(.dinb(n26466), .dina(n4254), .dout(n4258));
    jand g1101(.dinb(G205gat), .dina(G375gat), .dout(n4262));
    jnot g1102(.din(n4262), .dout(n4265));
    jand g1103(.dinb(n3901), .dina(n27762), .dout(n4269));
    jand g1104(.dinb(n27759), .dina(n3959), .dout(n4273));
    jor g1105(.dinb(n27717), .dina(n4273), .dout(n4277));
    jand g1106(.dinb(G222gat), .dina(G358gat), .dout(n4281));
    jnot g1107(.din(n4281), .dout(n4284));
    jand g1108(.dinb(n3920), .dina(n31425), .dout(n4288));
    jand g1109(.dinb(n31416), .dina(n3951), .dout(n4292));
    jor g1110(.dinb(n31383), .dina(n4292), .dout(n4296));
    jand g1111(.dinb(G239gat), .dina(G341gat), .dout(n4300));
    jand g1112(.dinb(G256gat), .dina(G324gat), .dout(n4304));
    jor g1113(.dinb(n31440), .dina(n3936), .dout(n4308));
    jor g1114(.dinb(n31461), .dina(n3943), .dout(n4312));
    jand g1115(.dinb(n31320), .dina(n4312), .dout(n4316));
    jxor g1116(.dinb(n31347), .dina(n4316), .dout(n4320));
    jnot g1117(.din(n4320), .dout(n4323));
    jxor g1118(.dinb(n31380), .dina(n4323), .dout(n4327));
    jxor g1119(.dinb(n4296), .dina(n31314), .dout(n4331));
    jxor g1120(.dinb(n31308), .dina(n4331), .dout(n4335));
    jxor g1121(.dinb(n4277), .dina(n27714), .dout(n4339));
    jxor g1122(.dinb(n27711), .dina(n4339), .dout(n4343));
    jxor g1123(.dinb(n4258), .dina(n26463), .dout(n4347));
    jxor g1124(.dinb(n26460), .dina(n4347), .dout(n4351));
    jxor g1125(.dinb(n4239), .dina(n25236), .dout(n4355));
    jxor g1126(.dinb(n25233), .dina(n4355), .dout(n4359));
    jxor g1127(.dinb(n4220), .dina(n24021), .dout(n4363));
    jxor g1128(.dinb(n24018), .dina(n4363), .dout(n4367));
    jxor g1129(.dinb(n4201), .dina(n22803), .dout(n4371));
    jxor g1130(.dinb(n22800), .dina(n4371), .dout(n4375));
    jxor g1131(.dinb(n4182), .dina(n21573), .dout(n4379));
    jxor g1132(.dinb(n21570), .dina(n4379), .dout(n4383));
    jxor g1133(.dinb(n4163), .dina(n4383), .dout(n4387));
    jxor g1134(.dinb(n20397), .dina(n4387), .dout(n4391));
    jxor g1135(.dinb(n4144), .dina(n4391), .dout(n4395));
    jxor g1136(.dinb(n19269), .dina(n4395), .dout(n4399));
    jxor g1137(.dinb(n4125), .dina(n18117), .dout(n4403));
    jxor g1138(.dinb(n18114), .dina(n4403), .dout(n4407));
    jnot g1139(.din(n4407), .dout(n4410));
    jxor g1140(.dinb(n4106), .dina(n16941), .dout(n4414));
    jnot g1141(.din(n4414), .dout(n4417));
    jxor g1142(.dinb(n16938), .dina(n4417), .dout(n4421));
    jxor g1143(.dinb(n15756), .dina(n4421), .dout(n4425));
    jnot g1144(.din(n4425), .dout(n4428));
    jxor g1145(.dinb(n4072), .dina(n4428), .dout(n4432));
    jnot g1146(.din(n4421), .dout(n4435));
    jor g1147(.dinb(n15752), .dina(n4435), .dout(n4439));
    jor g1148(.dinb(n4072), .dina(n12773), .dout(n4443));
    jand g1149(.dinb(n12771), .dina(n4443), .dout(n4447));
    jor g1150(.dinb(n4106), .dina(n16941), .dout(n4451));
    jor g1151(.dinb(n16938), .dina(n4417), .dout(n4455));
    jand g1152(.dinb(n16803), .dina(n4455), .dout(n4459));
    jand g1153(.dinb(G69gat), .dina(G528gat), .dout(n4463));
    jand g1154(.dinb(n4125), .dina(n18117), .dout(n4467));
    jand g1155(.dinb(n18114), .dina(n4403), .dout(n4471));
    jor g1156(.dinb(n17997), .dina(n4471), .dout(n4475));
    jand g1157(.dinb(G86gat), .dina(G511gat), .dout(n4479));
    jnot g1158(.din(n4479), .dout(n4482));
    jand g1159(.dinb(n4144), .dina(n4391), .dout(n4486));
    jand g1160(.dinb(n19269), .dina(n4395), .dout(n4490));
    jor g1161(.dinb(n19161), .dina(n4490), .dout(n4494));
    jand g1162(.dinb(G103gat), .dina(G494gat), .dout(n4498));
    jnot g1163(.din(n4498), .dout(n4501));
    jand g1164(.dinb(n4163), .dina(n4383), .dout(n4505));
    jand g1165(.dinb(n20397), .dina(n4387), .dout(n4509));
    jor g1166(.dinb(n20295), .dina(n4509), .dout(n4513));
    jand g1167(.dinb(G120gat), .dina(G477gat), .dout(n4517));
    jnot g1168(.din(n4517), .dout(n4520));
    jand g1169(.dinb(n4182), .dina(n21573), .dout(n4524));
    jand g1170(.dinb(n21570), .dina(n4379), .dout(n4528));
    jor g1171(.dinb(n21474), .dina(n4528), .dout(n4532));
    jand g1172(.dinb(G137gat), .dina(G460gat), .dout(n4536));
    jnot g1173(.din(n4536), .dout(n4539));
    jand g1174(.dinb(n4201), .dina(n22803), .dout(n4543));
    jand g1175(.dinb(n22800), .dina(n4371), .dout(n4547));
    jor g1176(.dinb(n22713), .dina(n4547), .dout(n4551));
    jand g1177(.dinb(G154gat), .dina(G443gat), .dout(n4555));
    jnot g1178(.din(n4555), .dout(n4558));
    jand g1179(.dinb(n4220), .dina(n24021), .dout(n4562));
    jand g1180(.dinb(n24018), .dina(n4363), .dout(n4566));
    jor g1181(.dinb(n23940), .dina(n4566), .dout(n4570));
    jand g1182(.dinb(G171gat), .dina(G426gat), .dout(n4574));
    jnot g1183(.din(n4574), .dout(n4577));
    jand g1184(.dinb(n4239), .dina(n25236), .dout(n4581));
    jand g1185(.dinb(n25233), .dina(n4355), .dout(n4585));
    jor g1186(.dinb(n25164), .dina(n4585), .dout(n4589));
    jand g1187(.dinb(G188gat), .dina(G409gat), .dout(n4593));
    jnot g1188(.din(n4593), .dout(n4596));
    jand g1189(.dinb(n4258), .dina(n26463), .dout(n4600));
    jand g1190(.dinb(n26460), .dina(n4347), .dout(n4604));
    jor g1191(.dinb(n26400), .dina(n4604), .dout(n4608));
    jand g1192(.dinb(G205gat), .dina(G392gat), .dout(n4612));
    jnot g1193(.din(n4612), .dout(n4615));
    jand g1194(.dinb(n4277), .dina(n27714), .dout(n4619));
    jand g1195(.dinb(n27711), .dina(n4339), .dout(n4623));
    jor g1196(.dinb(n27660), .dina(n4623), .dout(n4627));
    jand g1197(.dinb(G222gat), .dina(G375gat), .dout(n4631));
    jnot g1198(.din(n4631), .dout(n4634));
    jand g1199(.dinb(n4296), .dina(n31314), .dout(n4638));
    jand g1200(.dinb(n31308), .dina(n4331), .dout(n4642));
    jor g1201(.dinb(n31266), .dina(n4642), .dout(n4646));
    jand g1202(.dinb(G239gat), .dina(G358gat), .dout(n4650));
    jand g1203(.dinb(G256gat), .dina(G341gat), .dout(n4654));
    jor g1204(.dinb(n31347), .dina(n4316), .dout(n4658));
    jor g1205(.dinb(n31380), .dina(n4323), .dout(n4662));
    jand g1206(.dinb(n31179), .dina(n4662), .dout(n4666));
    jxor g1207(.dinb(n31218), .dina(n4666), .dout(n4670));
    jnot g1208(.din(n4670), .dout(n4673));
    jxor g1209(.dinb(n31263), .dina(n4673), .dout(n4677));
    jxor g1210(.dinb(n4646), .dina(n31173), .dout(n4681));
    jxor g1211(.dinb(n31170), .dina(n4681), .dout(n4685));
    jxor g1212(.dinb(n4627), .dina(n27657), .dout(n4689));
    jxor g1213(.dinb(n27654), .dina(n4689), .dout(n4693));
    jxor g1214(.dinb(n4608), .dina(n26397), .dout(n4697));
    jxor g1215(.dinb(n26394), .dina(n4697), .dout(n4701));
    jxor g1216(.dinb(n4589), .dina(n25161), .dout(n4705));
    jxor g1217(.dinb(n25158), .dina(n4705), .dout(n4709));
    jxor g1218(.dinb(n4570), .dina(n23937), .dout(n4713));
    jxor g1219(.dinb(n23934), .dina(n4713), .dout(n4717));
    jxor g1220(.dinb(n4551), .dina(n22710), .dout(n4721));
    jxor g1221(.dinb(n22707), .dina(n4721), .dout(n4725));
    jxor g1222(.dinb(n4532), .dina(n21471), .dout(n4729));
    jxor g1223(.dinb(n21468), .dina(n4729), .dout(n4733));
    jxor g1224(.dinb(n4513), .dina(n4733), .dout(n4737));
    jxor g1225(.dinb(n20292), .dina(n4737), .dout(n4741));
    jxor g1226(.dinb(n4494), .dina(n4741), .dout(n4745));
    jxor g1227(.dinb(n19158), .dina(n4745), .dout(n4749));
    jxor g1228(.dinb(n4475), .dina(n17993), .dout(n4753));
    jnot g1229(.din(n4753), .dout(n4756));
    jxor g1230(.dinb(n17988), .dina(n4756), .dout(n4760));
    jxor g1231(.dinb(n4459), .dina(n16793), .dout(n4764));
    jnot g1232(.din(n4764), .dout(n4767));
    jxor g1233(.dinb(n4447), .dina(n11544), .dout(n4771));
    jnot g1234(.din(n4760), .dout(n4774));
    jor g1235(.dinb(n4459), .dina(n16791), .dout(n4778));
    jor g1236(.dinb(n4447), .dina(n12764), .dout(n4782));
    jand g1237(.dinb(n12762), .dina(n4782), .dout(n4786));
    jnot g1238(.din(n4475), .dout(n4789));
    jnot g1239(.din(n4749), .dout(n4792));
    jor g1240(.dinb(n4789), .dina(n17991), .dout(n4796));
    jor g1241(.dinb(n17988), .dina(n4756), .dout(n4800));
    jand g1242(.dinb(n17856), .dina(n4800), .dout(n4804));
    jand g1243(.dinb(G86gat), .dina(G528gat), .dout(n4808));
    jand g1244(.dinb(n4494), .dina(n4741), .dout(n4812));
    jand g1245(.dinb(n19158), .dina(n4745), .dout(n4816));
    jor g1246(.dinb(n19041), .dina(n4816), .dout(n4820));
    jand g1247(.dinb(G103gat), .dina(G511gat), .dout(n4824));
    jnot g1248(.din(n4824), .dout(n4827));
    jand g1249(.dinb(n4513), .dina(n4733), .dout(n4831));
    jand g1250(.dinb(n20292), .dina(n4737), .dout(n4835));
    jor g1251(.dinb(n20181), .dina(n4835), .dout(n4839));
    jand g1252(.dinb(G120gat), .dina(G494gat), .dout(n4843));
    jnot g1253(.din(n4843), .dout(n4846));
    jand g1254(.dinb(n4532), .dina(n21471), .dout(n4850));
    jand g1255(.dinb(n21468), .dina(n4729), .dout(n4854));
    jor g1256(.dinb(n21363), .dina(n4854), .dout(n4858));
    jand g1257(.dinb(G137gat), .dina(G477gat), .dout(n4862));
    jnot g1258(.din(n4862), .dout(n4865));
    jand g1259(.dinb(n4551), .dina(n22710), .dout(n4869));
    jand g1260(.dinb(n22707), .dina(n4721), .dout(n4873));
    jor g1261(.dinb(n22611), .dina(n4873), .dout(n4877));
    jand g1262(.dinb(G154gat), .dina(G460gat), .dout(n4881));
    jnot g1263(.din(n4881), .dout(n4884));
    jand g1264(.dinb(n4570), .dina(n23937), .dout(n4888));
    jand g1265(.dinb(n23934), .dina(n4713), .dout(n4892));
    jor g1266(.dinb(n23847), .dina(n4892), .dout(n4896));
    jand g1267(.dinb(G171gat), .dina(G443gat), .dout(n4900));
    jnot g1268(.din(n4900), .dout(n4903));
    jand g1269(.dinb(n4589), .dina(n25161), .dout(n4907));
    jand g1270(.dinb(n25158), .dina(n4705), .dout(n4911));
    jor g1271(.dinb(n25080), .dina(n4911), .dout(n4915));
    jand g1272(.dinb(G188gat), .dina(G426gat), .dout(n4919));
    jnot g1273(.din(n4919), .dout(n4922));
    jand g1274(.dinb(n4608), .dina(n26397), .dout(n4926));
    jand g1275(.dinb(n26394), .dina(n4697), .dout(n4930));
    jor g1276(.dinb(n26325), .dina(n4930), .dout(n4934));
    jand g1277(.dinb(G205gat), .dina(G409gat), .dout(n4938));
    jnot g1278(.din(n4938), .dout(n4941));
    jand g1279(.dinb(n4627), .dina(n27657), .dout(n4945));
    jand g1280(.dinb(n27654), .dina(n4689), .dout(n4949));
    jor g1281(.dinb(n27594), .dina(n4949), .dout(n4953));
    jand g1282(.dinb(G222gat), .dina(G392gat), .dout(n4957));
    jnot g1283(.din(n4957), .dout(n4960));
    jand g1284(.dinb(n4646), .dina(n31173), .dout(n4964));
    jand g1285(.dinb(n31170), .dina(n4681), .dout(n4968));
    jor g1286(.dinb(n31119), .dina(n4968), .dout(n4972));
    jand g1287(.dinb(G239gat), .dina(G375gat), .dout(n4976));
    jand g1288(.dinb(G256gat), .dina(G358gat), .dout(n4980));
    jor g1289(.dinb(n31218), .dina(n4666), .dout(n4984));
    jor g1290(.dinb(n31263), .dina(n4673), .dout(n4988));
    jand g1291(.dinb(n31008), .dina(n4988), .dout(n4992));
    jxor g1292(.dinb(n31059), .dina(n4992), .dout(n4996));
    jnot g1293(.din(n4996), .dout(n4999));
    jxor g1294(.dinb(n31116), .dina(n4999), .dout(n5003));
    jxor g1295(.dinb(n4972), .dina(n5003), .dout(n5007));
    jxor g1296(.dinb(n31002), .dina(n5007), .dout(n5011));
    jxor g1297(.dinb(n4953), .dina(n27591), .dout(n5015));
    jxor g1298(.dinb(n27588), .dina(n5015), .dout(n5019));
    jxor g1299(.dinb(n4934), .dina(n26322), .dout(n5023));
    jxor g1300(.dinb(n26319), .dina(n5023), .dout(n5027));
    jxor g1301(.dinb(n4915), .dina(n25077), .dout(n5031));
    jxor g1302(.dinb(n25074), .dina(n5031), .dout(n5035));
    jxor g1303(.dinb(n4896), .dina(n23844), .dout(n5039));
    jxor g1304(.dinb(n23841), .dina(n5039), .dout(n5043));
    jxor g1305(.dinb(n4877), .dina(n22608), .dout(n5047));
    jxor g1306(.dinb(n22605), .dina(n5047), .dout(n5051));
    jxor g1307(.dinb(n4858), .dina(n21360), .dout(n5055));
    jxor g1308(.dinb(n21357), .dina(n5055), .dout(n5059));
    jxor g1309(.dinb(n4839), .dina(n5059), .dout(n5063));
    jxor g1310(.dinb(n20178), .dina(n5063), .dout(n5067));
    jxor g1311(.dinb(n4820), .dina(n5067), .dout(n5071));
    jnot g1312(.din(n5071), .dout(n5074));
    jxor g1313(.dinb(n19038), .dina(n5074), .dout(n5078));
    jnot g1314(.din(n5078), .dout(n5081));
    jxor g1315(.dinb(n4804), .dina(n5081), .dout(n5085));
    jxor g1316(.dinb(n4786), .dina(n12740), .dout(n5089));
    jor g1317(.dinb(n4804), .dina(n5081), .dout(n5093));
    jnot g1318(.din(n5085), .dout(n5096));
    jor g1319(.dinb(n4786), .dina(n12738), .dout(n5100));
    jand g1320(.dinb(n12726), .dina(n5100), .dout(n5104));
    jnot g1321(.din(n4820), .dout(n5107));
    jnot g1322(.din(n5067), .dout(n5110));
    jor g1323(.dinb(n5107), .dina(n5110), .dout(n5114));
    jor g1324(.dinb(n19038), .dina(n5074), .dout(n5118));
    jand g1325(.dinb(n18906), .dina(n5118), .dout(n5122));
    jand g1326(.dinb(G103gat), .dina(G528gat), .dout(n5126));
    jand g1327(.dinb(n4839), .dina(n5059), .dout(n5130));
    jand g1328(.dinb(n20178), .dina(n5063), .dout(n5134));
    jor g1329(.dinb(n20058), .dina(n5134), .dout(n5138));
    jand g1330(.dinb(G120gat), .dina(G511gat), .dout(n5142));
    jnot g1331(.din(n5142), .dout(n5145));
    jand g1332(.dinb(n4858), .dina(n21360), .dout(n5149));
    jand g1333(.dinb(n21357), .dina(n5055), .dout(n5153));
    jor g1334(.dinb(n21243), .dina(n5153), .dout(n5157));
    jand g1335(.dinb(G137gat), .dina(G494gat), .dout(n5161));
    jnot g1336(.din(n5161), .dout(n5164));
    jand g1337(.dinb(n4877), .dina(n22608), .dout(n5168));
    jand g1338(.dinb(n22605), .dina(n5047), .dout(n5172));
    jor g1339(.dinb(n22500), .dina(n5172), .dout(n5176));
    jand g1340(.dinb(G154gat), .dina(G477gat), .dout(n5180));
    jnot g1341(.din(n5180), .dout(n5183));
    jand g1342(.dinb(n4896), .dina(n23844), .dout(n5187));
    jand g1343(.dinb(n23841), .dina(n5039), .dout(n5191));
    jor g1344(.dinb(n23745), .dina(n5191), .dout(n5195));
    jand g1345(.dinb(G171gat), .dina(G460gat), .dout(n5199));
    jnot g1346(.din(n5199), .dout(n5202));
    jand g1347(.dinb(n4915), .dina(n25077), .dout(n5206));
    jand g1348(.dinb(n25074), .dina(n5031), .dout(n5210));
    jor g1349(.dinb(n24987), .dina(n5210), .dout(n5214));
    jand g1350(.dinb(G188gat), .dina(G443gat), .dout(n5218));
    jnot g1351(.din(n5218), .dout(n5221));
    jand g1352(.dinb(n4934), .dina(n26322), .dout(n5225));
    jand g1353(.dinb(n26319), .dina(n5023), .dout(n5229));
    jor g1354(.dinb(n26241), .dina(n5229), .dout(n5233));
    jand g1355(.dinb(G205gat), .dina(G426gat), .dout(n5237));
    jnot g1356(.din(n5237), .dout(n5240));
    jand g1357(.dinb(n4953), .dina(n27591), .dout(n5244));
    jand g1358(.dinb(n27588), .dina(n5015), .dout(n5248));
    jor g1359(.dinb(n27519), .dina(n5248), .dout(n5252));
    jand g1360(.dinb(G222gat), .dina(G409gat), .dout(n5256));
    jnot g1361(.din(n5256), .dout(n5259));
    jand g1362(.dinb(n4972), .dina(n5003), .dout(n5263));
    jand g1363(.dinb(n31002), .dina(n5007), .dout(n5267));
    jor g1364(.dinb(n30942), .dina(n5267), .dout(n5271));
    jand g1365(.dinb(G239gat), .dina(G392gat), .dout(n5275));
    jand g1366(.dinb(G256gat), .dina(G375gat), .dout(n5279));
    jor g1367(.dinb(n31059), .dina(n4992), .dout(n5283));
    jor g1368(.dinb(n31116), .dina(n4999), .dout(n5287));
    jand g1369(.dinb(n30804), .dina(n5287), .dout(n5291));
    jxor g1370(.dinb(n30867), .dina(n5291), .dout(n5295));
    jnot g1371(.din(n5295), .dout(n5298));
    jxor g1372(.dinb(n30936), .dina(n5298), .dout(n5302));
    jxor g1373(.dinb(n30939), .dina(n5302), .dout(n5306));
    jxor g1374(.dinb(n30798), .dina(n5306), .dout(n5310));
    jxor g1375(.dinb(n5252), .dina(n5310), .dout(n5314));
    jxor g1376(.dinb(n27516), .dina(n5314), .dout(n5318));
    jxor g1377(.dinb(n5233), .dina(n26238), .dout(n5322));
    jxor g1378(.dinb(n26235), .dina(n5322), .dout(n5326));
    jxor g1379(.dinb(n5214), .dina(n24984), .dout(n5330));
    jxor g1380(.dinb(n24981), .dina(n5330), .dout(n5334));
    jxor g1381(.dinb(n5195), .dina(n23742), .dout(n5338));
    jxor g1382(.dinb(n23739), .dina(n5338), .dout(n5342));
    jxor g1383(.dinb(n5176), .dina(n22497), .dout(n5346));
    jxor g1384(.dinb(n22494), .dina(n5346), .dout(n5350));
    jxor g1385(.dinb(n5157), .dina(n21240), .dout(n5354));
    jxor g1386(.dinb(n21237), .dina(n5354), .dout(n5358));
    jxor g1387(.dinb(n5138), .dina(n5358), .dout(n5362));
    jnot g1388(.din(n5362), .dout(n5365));
    jxor g1389(.dinb(n20055), .dina(n5365), .dout(n5369));
    jnot g1390(.din(n5369), .dout(n5372));
    jxor g1391(.dinb(n18903), .dina(n5372), .dout(n5376));
    jxor g1392(.dinb(n5104), .dina(n12692), .dout(n5380));
    jor g1393(.dinb(n18903), .dina(n5372), .dout(n5384));
    jnot g1394(.din(n5376), .dout(n5387));
    jor g1395(.dinb(n5104), .dina(n12690), .dout(n5391));
    jand g1396(.dinb(n12675), .dina(n5391), .dout(n5395));
    jnot g1397(.din(n5138), .dout(n5398));
    jnot g1398(.din(n5358), .dout(n5401));
    jor g1399(.dinb(n5398), .dina(n5401), .dout(n5405));
    jor g1400(.dinb(n20055), .dina(n5365), .dout(n5409));
    jand g1401(.dinb(n19920), .dina(n5409), .dout(n5413));
    jand g1402(.dinb(G120gat), .dina(G528gat), .dout(n5417));
    jand g1403(.dinb(n5157), .dina(n21240), .dout(n5421));
    jand g1404(.dinb(n21237), .dina(n5354), .dout(n5425));
    jor g1405(.dinb(n21114), .dina(n5425), .dout(n5429));
    jand g1406(.dinb(G137gat), .dina(G511gat), .dout(n5433));
    jnot g1407(.din(n5433), .dout(n5436));
    jand g1408(.dinb(n5176), .dina(n22497), .dout(n5440));
    jand g1409(.dinb(n22494), .dina(n5346), .dout(n5444));
    jor g1410(.dinb(n22380), .dina(n5444), .dout(n5448));
    jand g1411(.dinb(G154gat), .dina(G494gat), .dout(n5452));
    jnot g1412(.din(n5452), .dout(n5455));
    jand g1413(.dinb(n5195), .dina(n23742), .dout(n5459));
    jand g1414(.dinb(n23739), .dina(n5338), .dout(n5463));
    jor g1415(.dinb(n23634), .dina(n5463), .dout(n5467));
    jand g1416(.dinb(G171gat), .dina(G477gat), .dout(n5471));
    jnot g1417(.din(n5471), .dout(n5474));
    jand g1418(.dinb(n5214), .dina(n24984), .dout(n5478));
    jand g1419(.dinb(n24981), .dina(n5330), .dout(n5482));
    jor g1420(.dinb(n24885), .dina(n5482), .dout(n5486));
    jand g1421(.dinb(G188gat), .dina(G460gat), .dout(n5490));
    jnot g1422(.din(n5490), .dout(n5493));
    jand g1423(.dinb(n5233), .dina(n26238), .dout(n5497));
    jand g1424(.dinb(n26235), .dina(n5322), .dout(n5501));
    jor g1425(.dinb(n26148), .dina(n5501), .dout(n5505));
    jand g1426(.dinb(G205gat), .dina(G443gat), .dout(n5509));
    jnot g1427(.din(n5509), .dout(n5512));
    jand g1428(.dinb(n5252), .dina(n5310), .dout(n5516));
    jand g1429(.dinb(n27516), .dina(n5314), .dout(n5520));
    jor g1430(.dinb(n27438), .dina(n5520), .dout(n5524));
    jand g1431(.dinb(G222gat), .dina(G426gat), .dout(n5528));
    jnot g1432(.din(n5528), .dout(n5531));
    jand g1433(.dinb(n30939), .dina(n5302), .dout(n5535));
    jand g1434(.dinb(n30798), .dina(n5306), .dout(n5539));
    jor g1435(.dinb(n30726), .dina(n5539), .dout(n5543));
    jand g1436(.dinb(G239gat), .dina(G409gat), .dout(n5547));
    jand g1437(.dinb(G256gat), .dina(G392gat), .dout(n5551));
    jor g1438(.dinb(n30867), .dina(n5291), .dout(n5555));
    jor g1439(.dinb(n30936), .dina(n5298), .dout(n5559));
    jand g1440(.dinb(n30564), .dina(n5559), .dout(n5563));
    jxor g1441(.dinb(n30639), .dina(n5563), .dout(n5567));
    jnot g1442(.din(n5567), .dout(n5570));
    jxor g1443(.dinb(n30720), .dina(n5570), .dout(n5574));
    jxor g1444(.dinb(n30723), .dina(n5574), .dout(n5578));
    jxor g1445(.dinb(n30558), .dina(n5578), .dout(n5582));
    jxor g1446(.dinb(n27435), .dina(n5582), .dout(n5586));
    jxor g1447(.dinb(n27432), .dina(n5586), .dout(n5590));
    jxor g1448(.dinb(n5505), .dina(n5590), .dout(n5594));
    jxor g1449(.dinb(n26145), .dina(n5594), .dout(n5598));
    jxor g1450(.dinb(n5486), .dina(n24882), .dout(n5602));
    jxor g1451(.dinb(n24879), .dina(n5602), .dout(n5606));
    jxor g1452(.dinb(n5467), .dina(n23631), .dout(n5610));
    jxor g1453(.dinb(n23628), .dina(n5610), .dout(n5614));
    jxor g1454(.dinb(n5448), .dina(n22377), .dout(n5618));
    jxor g1455(.dinb(n22374), .dina(n5618), .dout(n5622));
    jxor g1456(.dinb(n5429), .dina(n21110), .dout(n5626));
    jnot g1457(.din(n5626), .dout(n5629));
    jxor g1458(.dinb(n21105), .dina(n5629), .dout(n5633));
    jnot g1459(.din(n5633), .dout(n5636));
    jxor g1460(.dinb(n19917), .dina(n5636), .dout(n5640));
    jxor g1461(.dinb(n5395), .dina(n12635), .dout(n5644));
    jor g1462(.dinb(n19917), .dina(n5636), .dout(n5648));
    jnot g1463(.din(n5640), .dout(n5651));
    jor g1464(.dinb(n5395), .dina(n12633), .dout(n5655));
    jand g1465(.dinb(n12615), .dina(n5655), .dout(n5659));
    jnot g1466(.din(n5429), .dout(n5662));
    jnot g1467(.din(n5622), .dout(n5665));
    jor g1468(.dinb(n5662), .dina(n21108), .dout(n5669));
    jor g1469(.dinb(n21105), .dina(n5629), .dout(n5673));
    jand g1470(.dinb(n20967), .dina(n5673), .dout(n5677));
    jand g1471(.dinb(G137gat), .dina(G528gat), .dout(n5681));
    jand g1472(.dinb(n5448), .dina(n22377), .dout(n5685));
    jand g1473(.dinb(n22374), .dina(n5618), .dout(n5689));
    jor g1474(.dinb(n22251), .dina(n5689), .dout(n5693));
    jand g1475(.dinb(G154gat), .dina(G511gat), .dout(n5697));
    jnot g1476(.din(n5697), .dout(n5700));
    jand g1477(.dinb(n5467), .dina(n23631), .dout(n5704));
    jand g1478(.dinb(n23628), .dina(n5610), .dout(n5708));
    jor g1479(.dinb(n23514), .dina(n5708), .dout(n5712));
    jand g1480(.dinb(G171gat), .dina(G494gat), .dout(n5716));
    jnot g1481(.din(n5716), .dout(n5719));
    jand g1482(.dinb(n5486), .dina(n24882), .dout(n5723));
    jand g1483(.dinb(n24879), .dina(n5602), .dout(n5727));
    jor g1484(.dinb(n24774), .dina(n5727), .dout(n5731));
    jand g1485(.dinb(G188gat), .dina(G477gat), .dout(n5735));
    jnot g1486(.din(n5735), .dout(n5738));
    jand g1487(.dinb(n5505), .dina(n5590), .dout(n5742));
    jand g1488(.dinb(n26145), .dina(n5594), .dout(n5746));
    jor g1489(.dinb(n26049), .dina(n5746), .dout(n5750));
    jand g1490(.dinb(G205gat), .dina(G460gat), .dout(n5754));
    jnot g1491(.din(n5754), .dout(n5757));
    jand g1492(.dinb(n27435), .dina(n5582), .dout(n5761));
    jand g1493(.dinb(n27432), .dina(n5586), .dout(n5765));
    jor g1494(.dinb(n27342), .dina(n5765), .dout(n5769));
    jand g1495(.dinb(G222gat), .dina(G443gat), .dout(n5773));
    jnot g1496(.din(n5773), .dout(n5776));
    jand g1497(.dinb(n30723), .dina(n5574), .dout(n5780));
    jand g1498(.dinb(n30558), .dina(n5578), .dout(n5784));
    jor g1499(.dinb(n30474), .dina(n5784), .dout(n5788));
    jand g1500(.dinb(G239gat), .dina(G426gat), .dout(n5792));
    jand g1501(.dinb(G256gat), .dina(G409gat), .dout(n5796));
    jor g1502(.dinb(n30639), .dina(n5563), .dout(n5800));
    jor g1503(.dinb(n30720), .dina(n5570), .dout(n5804));
    jand g1504(.dinb(n30288), .dina(n5804), .dout(n5808));
    jxor g1505(.dinb(n30375), .dina(n5808), .dout(n5812));
    jnot g1506(.din(n5812), .dout(n5815));
    jxor g1507(.dinb(n30468), .dina(n5815), .dout(n5819));
    jxor g1508(.dinb(n30471), .dina(n5819), .dout(n5823));
    jxor g1509(.dinb(n30282), .dina(n5823), .dout(n5827));
    jxor g1510(.dinb(n27339), .dina(n5827), .dout(n5831));
    jxor g1511(.dinb(n27336), .dina(n5831), .dout(n5835));
    jxor g1512(.dinb(n26046), .dina(n5835), .dout(n5839));
    jxor g1513(.dinb(n26043), .dina(n5839), .dout(n5843));
    jxor g1514(.dinb(n5731), .dina(n5843), .dout(n5847));
    jxor g1515(.dinb(n24771), .dina(n5847), .dout(n5851));
    jxor g1516(.dinb(n5712), .dina(n23511), .dout(n5855));
    jxor g1517(.dinb(n23508), .dina(n5855), .dout(n5859));
    jxor g1518(.dinb(n5693), .dina(n22247), .dout(n5863));
    jnot g1519(.din(n5863), .dout(n5866));
    jxor g1520(.dinb(n22242), .dina(n5866), .dout(n5870));
    jnot g1521(.din(n5870), .dout(n5873));
    jxor g1522(.dinb(n5677), .dina(n5873), .dout(n5877));
    jxor g1523(.dinb(n5659), .dina(n12566), .dout(n5881));
    jor g1524(.dinb(n5677), .dina(n5873), .dout(n5885));
    jnot g1525(.din(n5877), .dout(n5888));
    jor g1526(.dinb(n5659), .dina(n12564), .dout(n5892));
    jand g1527(.dinb(n12540), .dina(n5892), .dout(n5896));
    jnot g1528(.din(n5693), .dout(n5899));
    jnot g1529(.din(n5859), .dout(n5902));
    jor g1530(.dinb(n5899), .dina(n22245), .dout(n5906));
    jor g1531(.dinb(n22242), .dina(n5866), .dout(n5910));
    jand g1532(.dinb(n22104), .dina(n5910), .dout(n5914));
    jand g1533(.dinb(G154gat), .dina(G528gat), .dout(n5918));
    jand g1534(.dinb(n5712), .dina(n23511), .dout(n5922));
    jand g1535(.dinb(n23508), .dina(n5855), .dout(n5926));
    jor g1536(.dinb(n23385), .dina(n5926), .dout(n5930));
    jand g1537(.dinb(G171gat), .dina(G511gat), .dout(n5934));
    jnot g1538(.din(n5934), .dout(n5937));
    jand g1539(.dinb(n5731), .dina(n5843), .dout(n5941));
    jand g1540(.dinb(n24771), .dina(n5847), .dout(n5945));
    jor g1541(.dinb(n24657), .dina(n5945), .dout(n5949));
    jand g1542(.dinb(G188gat), .dina(G494gat), .dout(n5953));
    jnot g1543(.din(n5953), .dout(n5956));
    jand g1544(.dinb(n26046), .dina(n5835), .dout(n5960));
    jand g1545(.dinb(n26043), .dina(n5839), .dout(n5964));
    jor g1546(.dinb(n25935), .dina(n5964), .dout(n5968));
    jand g1547(.dinb(G205gat), .dina(G477gat), .dout(n5972));
    jnot g1548(.din(n5972), .dout(n5975));
    jand g1549(.dinb(n27339), .dina(n5827), .dout(n5979));
    jand g1550(.dinb(n27336), .dina(n5831), .dout(n5983));
    jor g1551(.dinb(n27234), .dina(n5983), .dout(n5987));
    jand g1552(.dinb(G222gat), .dina(G460gat), .dout(n5991));
    jnot g1553(.din(n5991), .dout(n5994));
    jand g1554(.dinb(n30471), .dina(n5819), .dout(n5998));
    jand g1555(.dinb(n30282), .dina(n5823), .dout(n6002));
    jor g1556(.dinb(n30186), .dina(n6002), .dout(n6006));
    jand g1557(.dinb(G239gat), .dina(G443gat), .dout(n6010));
    jand g1558(.dinb(G256gat), .dina(G426gat), .dout(n6014));
    jor g1559(.dinb(n30375), .dina(n5808), .dout(n6018));
    jor g1560(.dinb(n30468), .dina(n5815), .dout(n6022));
    jand g1561(.dinb(n29976), .dina(n6022), .dout(n6026));
    jxor g1562(.dinb(n30075), .dina(n6026), .dout(n6030));
    jnot g1563(.din(n6030), .dout(n6033));
    jxor g1564(.dinb(n30180), .dina(n6033), .dout(n6037));
    jxor g1565(.dinb(n30183), .dina(n6037), .dout(n6041));
    jxor g1566(.dinb(n29970), .dina(n6041), .dout(n6045));
    jxor g1567(.dinb(n27231), .dina(n6045), .dout(n6049));
    jxor g1568(.dinb(n27228), .dina(n6049), .dout(n6053));
    jxor g1569(.dinb(n25932), .dina(n6053), .dout(n6057));
    jxor g1570(.dinb(n25929), .dina(n6057), .dout(n6061));
    jxor g1571(.dinb(n24654), .dina(n6061), .dout(n6065));
    jxor g1572(.dinb(n24651), .dina(n6065), .dout(n6069));
    jxor g1573(.dinb(n5930), .dina(n6069), .dout(n6073));
    jnot g1574(.din(n6073), .dout(n6076));
    jxor g1575(.dinb(n23382), .dina(n6076), .dout(n6080));
    jnot g1576(.din(n6080), .dout(n6083));
    jxor g1577(.dinb(n5914), .dina(n6083), .dout(n6087));
    jxor g1578(.dinb(n5896), .dina(n12479), .dout(n6091));
    jor g1579(.dinb(n5914), .dina(n6083), .dout(n6095));
    jnot g1580(.din(n6087), .dout(n6098));
    jor g1581(.dinb(n5896), .dina(n12477), .dout(n6102));
    jand g1582(.dinb(n12447), .dina(n6102), .dout(n6106));
    jnot g1583(.din(n5930), .dout(n6109));
    jnot g1584(.din(n6069), .dout(n6112));
    jor g1585(.dinb(n6109), .dina(n6112), .dout(n6116));
    jor g1586(.dinb(n23382), .dina(n6076), .dout(n6120));
    jand g1587(.dinb(n23244), .dina(n6120), .dout(n6124));
    jand g1588(.dinb(G171gat), .dina(G528gat), .dout(n6128));
    jnot g1589(.din(n6128), .dout(n6131));
    jand g1590(.dinb(n24654), .dina(n6061), .dout(n6135));
    jand g1591(.dinb(n24651), .dina(n6065), .dout(n6139));
    jor g1592(.dinb(n24525), .dina(n6139), .dout(n6143));
    jand g1593(.dinb(G188gat), .dina(G511gat), .dout(n6147));
    jnot g1594(.din(n6147), .dout(n6150));
    jand g1595(.dinb(n25932), .dina(n6053), .dout(n6154));
    jand g1596(.dinb(n25929), .dina(n6057), .dout(n6158));
    jor g1597(.dinb(n25809), .dina(n6158), .dout(n6162));
    jand g1598(.dinb(G205gat), .dina(G494gat), .dout(n6166));
    jnot g1599(.din(n6166), .dout(n6169));
    jand g1600(.dinb(n27231), .dina(n6045), .dout(n6173));
    jand g1601(.dinb(n27228), .dina(n6049), .dout(n6177));
    jor g1602(.dinb(n27114), .dina(n6177), .dout(n6181));
    jand g1603(.dinb(G222gat), .dina(G477gat), .dout(n6185));
    jnot g1604(.din(n6185), .dout(n6188));
    jand g1605(.dinb(n30183), .dina(n6037), .dout(n6192));
    jand g1606(.dinb(n29970), .dina(n6041), .dout(n6196));
    jor g1607(.dinb(n29862), .dina(n6196), .dout(n6200));
    jand g1608(.dinb(G239gat), .dina(G460gat), .dout(n6204));
    jand g1609(.dinb(G256gat), .dina(G443gat), .dout(n6208));
    jor g1610(.dinb(n30075), .dina(n6026), .dout(n6212));
    jor g1611(.dinb(n30180), .dina(n6033), .dout(n6216));
    jand g1612(.dinb(n29628), .dina(n6216), .dout(n6220));
    jxor g1613(.dinb(n29739), .dina(n6220), .dout(n6224));
    jnot g1614(.din(n6224), .dout(n6227));
    jxor g1615(.dinb(n29856), .dina(n6227), .dout(n6231));
    jxor g1616(.dinb(n29859), .dina(n6231), .dout(n6235));
    jxor g1617(.dinb(n29622), .dina(n6235), .dout(n6239));
    jxor g1618(.dinb(n27111), .dina(n6239), .dout(n6243));
    jxor g1619(.dinb(n27108), .dina(n6243), .dout(n6247));
    jxor g1620(.dinb(n25806), .dina(n6247), .dout(n6251));
    jxor g1621(.dinb(n25803), .dina(n6251), .dout(n6255));
    jxor g1622(.dinb(n24522), .dina(n6255), .dout(n6259));
    jxor g1623(.dinb(n24519), .dina(n6259), .dout(n6263));
    jnot g1624(.din(n6263), .dout(n6266));
    jxor g1625(.dinb(n23241), .dina(n6266), .dout(n6270));
    jxor g1626(.dinb(n6106), .dina(n12377), .dout(n6274));
    jor g1627(.dinb(n23241), .dina(n6266), .dout(n6278));
    jnot g1628(.din(n6270), .dout(n6281));
    jor g1629(.dinb(n6106), .dina(n12375), .dout(n6285));
    jand g1630(.dinb(n12342), .dina(n6285), .dout(n6289));
    jand g1631(.dinb(n24522), .dina(n6255), .dout(n6293));
    jand g1632(.dinb(n24519), .dina(n6259), .dout(n6297));
    jor g1633(.dinb(n24381), .dina(n6297), .dout(n6301));
    jand g1634(.dinb(G188gat), .dina(G528gat), .dout(n6305));
    jnot g1635(.din(n6305), .dout(n6308));
    jand g1636(.dinb(n25806), .dina(n6247), .dout(n6312));
    jand g1637(.dinb(n25803), .dina(n6251), .dout(n6316));
    jor g1638(.dinb(n25671), .dina(n6316), .dout(n6320));
    jand g1639(.dinb(G205gat), .dina(G511gat), .dout(n6324));
    jnot g1640(.din(n6324), .dout(n6327));
    jand g1641(.dinb(n27111), .dina(n6239), .dout(n6331));
    jand g1642(.dinb(n27108), .dina(n6243), .dout(n6335));
    jor g1643(.dinb(n26982), .dina(n6335), .dout(n6339));
    jand g1644(.dinb(G222gat), .dina(G494gat), .dout(n6343));
    jnot g1645(.din(n6343), .dout(n6346));
    jand g1646(.dinb(n29859), .dina(n6231), .dout(n6350));
    jand g1647(.dinb(n29622), .dina(n6235), .dout(n6354));
    jor g1648(.dinb(n29502), .dina(n6354), .dout(n6358));
    jand g1649(.dinb(G239gat), .dina(G477gat), .dout(n6362));
    jand g1650(.dinb(G256gat), .dina(G460gat), .dout(n6366));
    jor g1651(.dinb(n29739), .dina(n6220), .dout(n6370));
    jor g1652(.dinb(n29856), .dina(n6227), .dout(n6374));
    jand g1653(.dinb(n29244), .dina(n6374), .dout(n6378));
    jxor g1654(.dinb(n29367), .dina(n6378), .dout(n6382));
    jnot g1655(.din(n6382), .dout(n6385));
    jxor g1656(.dinb(n29496), .dina(n6385), .dout(n6389));
    jxor g1657(.dinb(n29499), .dina(n6389), .dout(n6393));
    jxor g1658(.dinb(n29238), .dina(n6393), .dout(n6397));
    jxor g1659(.dinb(n26979), .dina(n6397), .dout(n6401));
    jxor g1660(.dinb(n26976), .dina(n6401), .dout(n6405));
    jxor g1661(.dinb(n25668), .dina(n6405), .dout(n6409));
    jxor g1662(.dinb(n25665), .dina(n6409), .dout(n6413));
    jxor g1663(.dinb(n24377), .dina(n6413), .dout(n6417));
    jxor g1664(.dinb(n6289), .dina(n12266), .dout(n6421));
    jnot g1665(.din(n6301), .dout(n6424));
    jnot g1666(.din(n6413), .dout(n6427));
    jor g1667(.dinb(n24375), .dina(n6427), .dout(n6431));
    jnot g1668(.din(n6417), .dout(n6434));
    jor g1669(.dinb(n6289), .dina(n12264), .dout(n6438));
    jand g1670(.dinb(n12228), .dina(n6438), .dout(n6442));
    jand g1671(.dinb(n25668), .dina(n6405), .dout(n6446));
    jand g1672(.dinb(n25665), .dina(n6409), .dout(n6450));
    jor g1673(.dinb(n25521), .dina(n6450), .dout(n6454));
    jand g1674(.dinb(G205gat), .dina(G528gat), .dout(n6458));
    jnot g1675(.din(n6458), .dout(n6461));
    jand g1676(.dinb(n26979), .dina(n6397), .dout(n6465));
    jand g1677(.dinb(n26976), .dina(n6401), .dout(n6469));
    jor g1678(.dinb(n26838), .dina(n6469), .dout(n6473));
    jand g1679(.dinb(G222gat), .dina(G511gat), .dout(n6477));
    jnot g1680(.din(n6477), .dout(n6480));
    jand g1681(.dinb(n29499), .dina(n6389), .dout(n6484));
    jand g1682(.dinb(n29238), .dina(n6393), .dout(n6488));
    jor g1683(.dinb(n29106), .dina(n6488), .dout(n6492));
    jand g1684(.dinb(G239gat), .dina(G494gat), .dout(n6496));
    jand g1685(.dinb(G256gat), .dina(G477gat), .dout(n6500));
    jor g1686(.dinb(n29367), .dina(n6378), .dout(n6504));
    jor g1687(.dinb(n29496), .dina(n6385), .dout(n6508));
    jand g1688(.dinb(n28824), .dina(n6508), .dout(n6512));
    jxor g1689(.dinb(n28959), .dina(n6512), .dout(n6516));
    jnot g1690(.din(n6516), .dout(n6519));
    jxor g1691(.dinb(n29100), .dina(n6519), .dout(n6523));
    jxor g1692(.dinb(n29103), .dina(n6523), .dout(n6527));
    jxor g1693(.dinb(n28818), .dina(n6527), .dout(n6531));
    jxor g1694(.dinb(n26835), .dina(n6531), .dout(n6535));
    jxor g1695(.dinb(n26832), .dina(n6535), .dout(n6539));
    jxor g1696(.dinb(n25517), .dina(n6539), .dout(n6543));
    jxor g1697(.dinb(n6442), .dina(n12152), .dout(n6547));
    jnot g1698(.din(n6454), .dout(n6550));
    jnot g1699(.din(n6539), .dout(n6553));
    jor g1700(.dinb(n25515), .dina(n6553), .dout(n6557));
    jnot g1701(.din(n6543), .dout(n6560));
    jor g1702(.dinb(n6442), .dina(n12150), .dout(n6564));
    jand g1703(.dinb(n12114), .dina(n6564), .dout(n6568));
    jand g1704(.dinb(n26835), .dina(n6531), .dout(n6572));
    jand g1705(.dinb(n26832), .dina(n6535), .dout(n6576));
    jor g1706(.dinb(n26682), .dina(n6576), .dout(n6580));
    jand g1707(.dinb(G222gat), .dina(G528gat), .dout(n6584));
    jnot g1708(.din(n6584), .dout(n6587));
    jand g1709(.dinb(n29103), .dina(n6523), .dout(n6591));
    jand g1710(.dinb(n28818), .dina(n6527), .dout(n6595));
    jor g1711(.dinb(n28674), .dina(n6595), .dout(n6599));
    jand g1712(.dinb(G239gat), .dina(G511gat), .dout(n6603));
    jand g1713(.dinb(G256gat), .dina(G494gat), .dout(n6607));
    jor g1714(.dinb(n28959), .dina(n6512), .dout(n6611));
    jor g1715(.dinb(n29100), .dina(n6519), .dout(n6615));
    jand g1716(.dinb(n28368), .dina(n6615), .dout(n6619));
    jxor g1717(.dinb(n28515), .dina(n6619), .dout(n6623));
    jnot g1718(.din(n6623), .dout(n6626));
    jxor g1719(.dinb(n28668), .dina(n6626), .dout(n6630));
    jxor g1720(.dinb(n28671), .dina(n6630), .dout(n6634));
    jxor g1721(.dinb(n28362), .dina(n6634), .dout(n6638));
    jxor g1722(.dinb(n26678), .dina(n6638), .dout(n6642));
    jxor g1723(.dinb(n6568), .dina(n12038), .dout(n6646));
    jnot g1724(.din(n6580), .dout(n6649));
    jnot g1725(.din(n6638), .dout(n6652));
    jor g1726(.dinb(n26676), .dina(n6652), .dout(n6656));
    jnot g1727(.din(n6642), .dout(n6659));
    jor g1728(.dinb(n6568), .dina(n12036), .dout(n6663));
    jand g1729(.dinb(n12000), .dina(n6663), .dout(n6667));
    jand g1730(.dinb(n28671), .dina(n6630), .dout(n6671));
    jand g1731(.dinb(n28362), .dina(n6634), .dout(n6675));
    jor g1732(.dinb(n28206), .dina(n6675), .dout(n6679));
    jand g1733(.dinb(G239gat), .dina(G528gat), .dout(n6683));
    jand g1734(.dinb(G256gat), .dina(G511gat), .dout(n6687));
    jor g1735(.dinb(n28515), .dina(n6619), .dout(n6691));
    jor g1736(.dinb(n28668), .dina(n6626), .dout(n6695));
    jand g1737(.dinb(n27876), .dina(n6695), .dout(n6699));
    jxor g1738(.dinb(n28035), .dina(n6699), .dout(n6703));
    jnot g1739(.din(n6703), .dout(n6706));
    jxor g1740(.dinb(n28200), .dina(n6706), .dout(n6710));
    jxor g1741(.dinb(n28202), .dina(n6710), .dout(n6714));
    jxor g1742(.dinb(n6667), .dina(n11924), .dout(n6718));
    jand g1743(.dinb(G256gat), .dina(G528gat), .dout(n6722));
    jor g1744(.dinb(n28035), .dina(n6699), .dout(n6726));
    jor g1745(.dinb(n28200), .dina(n6706), .dout(n6730));
    jand g1746(.dinb(n11676), .dina(n6730), .dout(n6734));
    jor g1747(.dinb(n11847), .dina(n6734), .dout(n6738));
    jnot g1748(.din(n6679), .dout(n6741));
    jnot g1749(.din(n6710), .dout(n6744));
    jor g1750(.dinb(n27870), .dina(n6744), .dout(n6748));
    jnot g1751(.din(n6714), .dout(n6751));
    jor g1752(.dinb(n6667), .dina(n11922), .dout(n6755));
    jand g1753(.dinb(n11886), .dina(n6755), .dout(n6759));
    jxor g1754(.dinb(n11847), .dina(n6734), .dout(n6763));
    jnot g1755(.din(n6763), .dout(n6766));
    jor g1756(.dinb(n6759), .dina(n11628), .dout(n6770));
    jand g1757(.dinb(n11589), .dina(n6770), .dout(G6287gat));
    jxor g1758(.dinb(n6759), .dina(n11630), .dout(n6778));
    jdff dff_A_l6uLDiYR0_2(.din(n6778), .dout(G6288gat));
    jdff dff_A_N2tTzVE14_0(.din(n34721), .dout(G6280gat));
    jdff dff_A_PAyX2J2a8_0(.din(n34718), .dout(n34721));
    jdff dff_A_GvGhDXPx3_2(.din(n6718), .dout(n34718));
    jdff dff_A_j9NUrqag8_0(.din(n34712), .dout(G6270gat));
    jdff dff_A_ZVdSCnXX0_0(.din(n34709), .dout(n34712));
    jdff dff_A_wSRmAakt8_0(.din(n34706), .dout(n34709));
    jdff dff_A_KzyXslny6_0(.din(n34703), .dout(n34706));
    jdff dff_A_MtaWg8ib7_2(.din(n6646), .dout(n34703));
    jdff dff_A_OnBH3vUl3_0(.din(n34697), .dout(G6260gat));
    jdff dff_A_7HV5KXse8_0(.din(n34694), .dout(n34697));
    jdff dff_A_QWaLqLGT0_0(.din(n34691), .dout(n34694));
    jdff dff_A_apui6QwY8_0(.din(n34688), .dout(n34691));
    jdff dff_A_AvJiQkvT6_0(.din(n34685), .dout(n34688));
    jdff dff_A_zgz3aUWA5_0(.din(n34682), .dout(n34685));
    jdff dff_A_cTXjgFSt7_2(.din(n6547), .dout(n34682));
    jdff dff_A_JW9f4wSa2_0(.din(n34676), .dout(G6250gat));
    jdff dff_A_ytZxEyU76_0(.din(n34673), .dout(n34676));
    jdff dff_A_kuq4Pi7Z7_0(.din(n34670), .dout(n34673));
    jdff dff_A_WR9E9Aag2_0(.din(n34667), .dout(n34670));
    jdff dff_A_r3sMAMPb3_0(.din(n34664), .dout(n34667));
    jdff dff_A_AjLI4VpR0_0(.din(n34661), .dout(n34664));
    jdff dff_A_wDfxn7zY6_0(.din(n34658), .dout(n34661));
    jdff dff_A_x8t5Shk49_0(.din(n34655), .dout(n34658));
    jdff dff_A_c6Fm6OCo3_2(.din(n6421), .dout(n34655));
    jdff dff_A_vcl3bDJl7_0(.din(n34649), .dout(G6240gat));
    jdff dff_A_dua3Bi0M8_0(.din(n34646), .dout(n34649));
    jdff dff_A_b1vuRf3a4_0(.din(n34643), .dout(n34646));
    jdff dff_A_4PmcjKeH8_0(.din(n34640), .dout(n34643));
    jdff dff_A_udNx3lHZ0_0(.din(n34637), .dout(n34640));
    jdff dff_A_tBkbXq5g4_0(.din(n34634), .dout(n34637));
    jdff dff_A_Tyex67UV2_0(.din(n34631), .dout(n34634));
    jdff dff_A_bV8WZ6pc6_0(.din(n34628), .dout(n34631));
    jdff dff_A_esA7WomA6_0(.din(n34625), .dout(n34628));
    jdff dff_A_tJmfc1aX8_0(.din(n34622), .dout(n34625));
    jdff dff_A_FgSjYYdM3_2(.din(n6274), .dout(n34622));
    jdff dff_A_ldmD4Pg34_0(.din(n34616), .dout(G6230gat));
    jdff dff_A_PM8G6V623_0(.din(n34613), .dout(n34616));
    jdff dff_A_uD06ZPIu0_0(.din(n34610), .dout(n34613));
    jdff dff_A_Cv8Wk0hu7_0(.din(n34607), .dout(n34610));
    jdff dff_A_DKlpFjiM6_0(.din(n34604), .dout(n34607));
    jdff dff_A_GgkbaN2K3_0(.din(n34601), .dout(n34604));
    jdff dff_A_XTmRmp8A1_0(.din(n34598), .dout(n34601));
    jdff dff_A_P87da74r3_0(.din(n34595), .dout(n34598));
    jdff dff_A_CG92fvNm1_0(.din(n34592), .dout(n34595));
    jdff dff_A_j2EuERaM6_0(.din(n34589), .dout(n34592));
    jdff dff_A_5lHIJwDH5_0(.din(n34586), .dout(n34589));
    jdff dff_A_H03cf2lL9_0(.din(n34583), .dout(n34586));
    jdff dff_A_OWGNsutV7_2(.din(n6091), .dout(n34583));
    jdff dff_A_VtS6o35P7_0(.din(n34577), .dout(G6220gat));
    jdff dff_A_cW4hY6gH8_0(.din(n34574), .dout(n34577));
    jdff dff_A_ZJxOxn1Z9_0(.din(n34571), .dout(n34574));
    jdff dff_A_5CXZnEeV2_0(.din(n34568), .dout(n34571));
    jdff dff_A_EbVELEbw0_0(.din(n34565), .dout(n34568));
    jdff dff_A_MaLPbrWR8_0(.din(n34562), .dout(n34565));
    jdff dff_A_f1KZGQfn5_0(.din(n34559), .dout(n34562));
    jdff dff_A_vM5byLDi9_0(.din(n34556), .dout(n34559));
    jdff dff_A_cfkZlF4D1_0(.din(n34553), .dout(n34556));
    jdff dff_A_9sFUi5mS4_0(.din(n34550), .dout(n34553));
    jdff dff_A_Bi1nK5XC8_0(.din(n34547), .dout(n34550));
    jdff dff_A_CL7wU4204_0(.din(n34544), .dout(n34547));
    jdff dff_A_8al8690v7_0(.din(n34541), .dout(n34544));
    jdff dff_A_9CKZi3AS6_0(.din(n34538), .dout(n34541));
    jdff dff_A_5arqhEZw5_2(.din(n5881), .dout(n34538));
    jdff dff_A_uQFiSjFw0_0(.din(n34532), .dout(G6210gat));
    jdff dff_A_WU8237Lx4_0(.din(n34529), .dout(n34532));
    jdff dff_A_QYdJGrRl3_0(.din(n34526), .dout(n34529));
    jdff dff_A_MSuQjyhW9_0(.din(n34523), .dout(n34526));
    jdff dff_A_HaGpOdSV0_0(.din(n34520), .dout(n34523));
    jdff dff_A_kD5VZRvd3_0(.din(n34517), .dout(n34520));
    jdff dff_A_EAGjHtSv9_0(.din(n34514), .dout(n34517));
    jdff dff_A_Qm70PGdU8_0(.din(n34511), .dout(n34514));
    jdff dff_A_3GSiUFl94_0(.din(n34508), .dout(n34511));
    jdff dff_A_RyDYXRC51_0(.din(n34505), .dout(n34508));
    jdff dff_A_kM1wyV0K5_0(.din(n34502), .dout(n34505));
    jdff dff_A_hkNq3aHH0_0(.din(n34499), .dout(n34502));
    jdff dff_A_JNkMfS620_0(.din(n34496), .dout(n34499));
    jdff dff_A_6ivIQwPA9_0(.din(n34493), .dout(n34496));
    jdff dff_A_jmf8UfBV6_0(.din(n34490), .dout(n34493));
    jdff dff_A_RpX5OA6x2_0(.din(n34487), .dout(n34490));
    jdff dff_A_HN7yDTv85_2(.din(n5644), .dout(n34487));
    jdff dff_A_euOPKNzS4_0(.din(n34481), .dout(G6200gat));
    jdff dff_A_l2BaYcZ29_0(.din(n34478), .dout(n34481));
    jdff dff_A_105n3lWY2_0(.din(n34475), .dout(n34478));
    jdff dff_A_oOspxazI5_0(.din(n34472), .dout(n34475));
    jdff dff_A_XRf37nWQ7_0(.din(n34469), .dout(n34472));
    jdff dff_A_snNeLaxx7_0(.din(n34466), .dout(n34469));
    jdff dff_A_hwvQOeus6_0(.din(n34463), .dout(n34466));
    jdff dff_A_pA2bGjJH7_0(.din(n34460), .dout(n34463));
    jdff dff_A_giftbn219_0(.din(n34457), .dout(n34460));
    jdff dff_A_ENYoDgN90_0(.din(n34454), .dout(n34457));
    jdff dff_A_KDyyAq3I6_0(.din(n34451), .dout(n34454));
    jdff dff_A_z6O5gkmr2_0(.din(n34448), .dout(n34451));
    jdff dff_A_0gGD8cSC0_0(.din(n34445), .dout(n34448));
    jdff dff_A_ZlkLXRqS6_0(.din(n34442), .dout(n34445));
    jdff dff_A_GThilhKC2_0(.din(n34439), .dout(n34442));
    jdff dff_A_zMy2P6rC1_0(.din(n34436), .dout(n34439));
    jdff dff_A_dZ5hM3BL9_0(.din(n34433), .dout(n34436));
    jdff dff_A_YmJQOPXe6_0(.din(n34430), .dout(n34433));
    jdff dff_A_CdP4FEpr4_2(.din(n5380), .dout(n34430));
    jdff dff_A_upFUzfVE3_0(.din(n34424), .dout(G6190gat));
    jdff dff_A_mMZtzphy0_0(.din(n34421), .dout(n34424));
    jdff dff_A_oVAjaGor1_0(.din(n34418), .dout(n34421));
    jdff dff_A_Fkys4IKG2_0(.din(n34415), .dout(n34418));
    jdff dff_A_hz74bhKB2_0(.din(n34412), .dout(n34415));
    jdff dff_A_2gUMQ6Ez8_0(.din(n34409), .dout(n34412));
    jdff dff_A_uK05PgXN7_0(.din(n34406), .dout(n34409));
    jdff dff_A_nvlstr0F3_0(.din(n34403), .dout(n34406));
    jdff dff_A_nmauDiGY8_0(.din(n34400), .dout(n34403));
    jdff dff_A_uXi4uYz30_0(.din(n34397), .dout(n34400));
    jdff dff_A_y3QdUFRR8_0(.din(n34394), .dout(n34397));
    jdff dff_A_wU7Ypb4D1_0(.din(n34391), .dout(n34394));
    jdff dff_A_dv9MIYmE0_0(.din(n34388), .dout(n34391));
    jdff dff_A_EuHGMMbj1_0(.din(n34385), .dout(n34388));
    jdff dff_A_ou10IiEt3_0(.din(n34382), .dout(n34385));
    jdff dff_A_KJIJFdNi3_0(.din(n34379), .dout(n34382));
    jdff dff_A_V1TQ6Yxg8_0(.din(n34376), .dout(n34379));
    jdff dff_A_I70Es19W1_0(.din(n34373), .dout(n34376));
    jdff dff_A_t3iTvneP3_0(.din(n34370), .dout(n34373));
    jdff dff_A_nYyHfqI36_0(.din(n34367), .dout(n34370));
    jdff dff_A_yzVOykgA5_2(.din(n5089), .dout(n34367));
    jdff dff_A_ZzX8KFrT7_0(.din(n34361), .dout(G6180gat));
    jdff dff_A_HeJUNTxn5_0(.din(n34358), .dout(n34361));
    jdff dff_A_5hturpCd7_0(.din(n34355), .dout(n34358));
    jdff dff_A_sezIkoQa5_0(.din(n34352), .dout(n34355));
    jdff dff_A_PKjcF8ZR7_0(.din(n34349), .dout(n34352));
    jdff dff_A_lInS9lwp3_0(.din(n34346), .dout(n34349));
    jdff dff_A_zWlbSlYz7_0(.din(n34343), .dout(n34346));
    jdff dff_A_HIv5fYST7_0(.din(n34340), .dout(n34343));
    jdff dff_A_hSmILgKU8_0(.din(n34337), .dout(n34340));
    jdff dff_A_A4pMx8fq4_0(.din(n34334), .dout(n34337));
    jdff dff_A_dV7twkBH2_0(.din(n34331), .dout(n34334));
    jdff dff_A_QtSPrnah2_0(.din(n34328), .dout(n34331));
    jdff dff_A_Sb09y2jW7_0(.din(n34325), .dout(n34328));
    jdff dff_A_wsZ5ojC10_0(.din(n34322), .dout(n34325));
    jdff dff_A_olkl87Jj3_0(.din(n34319), .dout(n34322));
    jdff dff_A_3sKt7CUo6_0(.din(n34316), .dout(n34319));
    jdff dff_A_1Jc7roqJ1_0(.din(n34313), .dout(n34316));
    jdff dff_A_LEc3BTSR4_0(.din(n34310), .dout(n34313));
    jdff dff_A_dk5s9Qxe5_0(.din(n34307), .dout(n34310));
    jdff dff_A_2oxaerVo3_0(.din(n34304), .dout(n34307));
    jdff dff_A_y9lT7fhQ5_0(.din(n34301), .dout(n34304));
    jdff dff_A_OISVg6qP5_0(.din(n34298), .dout(n34301));
    jdff dff_A_5lkC1ky40_2(.din(n4771), .dout(n34298));
    jdff dff_A_nCWPNuLc1_0(.din(n34292), .dout(G6170gat));
    jdff dff_A_3MmwWSic9_0(.din(n34289), .dout(n34292));
    jdff dff_A_72L7YKCR9_0(.din(n34286), .dout(n34289));
    jdff dff_A_K7faFUhy4_0(.din(n34283), .dout(n34286));
    jdff dff_A_qXI94FpI0_0(.din(n34280), .dout(n34283));
    jdff dff_A_j1s66bpE5_0(.din(n34277), .dout(n34280));
    jdff dff_A_sQEAefrg6_0(.din(n34274), .dout(n34277));
    jdff dff_A_oUED2Fr67_0(.din(n34271), .dout(n34274));
    jdff dff_A_gS5j8tEI6_0(.din(n34268), .dout(n34271));
    jdff dff_A_SE7CBLWH4_0(.din(n34265), .dout(n34268));
    jdff dff_A_T5wClN0H7_0(.din(n34262), .dout(n34265));
    jdff dff_A_JkVAFg4G2_0(.din(n34259), .dout(n34262));
    jdff dff_A_c5N44hHk3_0(.din(n34256), .dout(n34259));
    jdff dff_A_H0X0Wm9v6_0(.din(n34253), .dout(n34256));
    jdff dff_A_N30RBU3j1_0(.din(n34250), .dout(n34253));
    jdff dff_A_a4aepqnD1_0(.din(n34247), .dout(n34250));
    jdff dff_A_7wOeM5Yg7_0(.din(n34244), .dout(n34247));
    jdff dff_A_xvfqY82a2_0(.din(n34241), .dout(n34244));
    jdff dff_A_jGs2LuPI6_0(.din(n34238), .dout(n34241));
    jdff dff_A_NpWq06f96_0(.din(n34235), .dout(n34238));
    jdff dff_A_LZyI69R21_0(.din(n34232), .dout(n34235));
    jdff dff_A_7RC0Upu28_0(.din(n34229), .dout(n34232));
    jdff dff_A_qbNEzUsY4_0(.din(n34226), .dout(n34229));
    jdff dff_A_CLR1cD3l5_0(.din(n34223), .dout(n34226));
    jdff dff_A_UyaYymEo5_2(.din(n4432), .dout(n34223));
    jdff dff_A_nESaPY9Y1_0(.din(n34217), .dout(G6160gat));
    jdff dff_A_QvzwaO3j7_0(.din(n34214), .dout(n34217));
    jdff dff_A_NM6yUNZu4_0(.din(n34211), .dout(n34214));
    jdff dff_A_CnQxLwoq5_0(.din(n34208), .dout(n34211));
    jdff dff_A_2kzLPTvc2_0(.din(n34205), .dout(n34208));
    jdff dff_A_8CQWHjB58_0(.din(n34202), .dout(n34205));
    jdff dff_A_mIDikPEU3_0(.din(n34199), .dout(n34202));
    jdff dff_A_Cpf0AO8S8_0(.din(n34196), .dout(n34199));
    jdff dff_A_yFybcONs6_0(.din(n34193), .dout(n34196));
    jdff dff_A_Cqeo3oVs2_0(.din(n34190), .dout(n34193));
    jdff dff_A_m7XT8p5y2_0(.din(n34187), .dout(n34190));
    jdff dff_A_SZPHObf33_0(.din(n34184), .dout(n34187));
    jdff dff_A_2r97kzzL1_0(.din(n34181), .dout(n34184));
    jdff dff_A_MFUeYaer4_0(.din(n34178), .dout(n34181));
    jdff dff_A_wkmvjhQv7_0(.din(n34175), .dout(n34178));
    jdff dff_A_8RJtbIcx6_0(.din(n34172), .dout(n34175));
    jdff dff_A_t9AJSCtL8_0(.din(n34169), .dout(n34172));
    jdff dff_A_ScY5LJbO9_0(.din(n34166), .dout(n34169));
    jdff dff_A_OXZH8Ev40_0(.din(n34163), .dout(n34166));
    jdff dff_A_cGcdneVv0_0(.din(n34160), .dout(n34163));
    jdff dff_A_EO82gKr26_0(.din(n34157), .dout(n34160));
    jdff dff_A_xWsUKLVc5_0(.din(n34154), .dout(n34157));
    jdff dff_A_Qeapd9vl1_0(.din(n34151), .dout(n34154));
    jdff dff_A_1tBOBIB03_0(.din(n34148), .dout(n34151));
    jdff dff_A_TH0McGuv2_0(.din(n34145), .dout(n34148));
    jdff dff_A_3iIVPtIy0_2(.din(n4057), .dout(n34145));
    jdff dff_A_hT8zARTA3_0(.din(n34139), .dout(G6150gat));
    jdff dff_A_ShKNXAb48_0(.din(n34136), .dout(n34139));
    jdff dff_A_uQZ1sL6C8_0(.din(n34133), .dout(n34136));
    jdff dff_A_TjEhGHcb0_0(.din(n34130), .dout(n34133));
    jdff dff_A_qvypK3uu5_0(.din(n34127), .dout(n34130));
    jdff dff_A_3hJ0cqb57_0(.din(n34124), .dout(n34127));
    jdff dff_A_XenvYTYa7_0(.din(n34121), .dout(n34124));
    jdff dff_A_TjnycSFa1_0(.din(n34118), .dout(n34121));
    jdff dff_A_fhHm3dOI4_0(.din(n34115), .dout(n34118));
    jdff dff_A_d4vweEuQ4_0(.din(n34112), .dout(n34115));
    jdff dff_A_IcRl3GVm5_0(.din(n34109), .dout(n34112));
    jdff dff_A_eMN0Lyhf3_0(.din(n34106), .dout(n34109));
    jdff dff_A_hGO9D4ZK3_0(.din(n34103), .dout(n34106));
    jdff dff_A_Q7M2dmfq1_0(.din(n34100), .dout(n34103));
    jdff dff_A_gfUeqGK95_0(.din(n34097), .dout(n34100));
    jdff dff_A_FORKC9420_0(.din(n34094), .dout(n34097));
    jdff dff_A_oic7v7yG5_0(.din(n34091), .dout(n34094));
    jdff dff_A_eb5JBGlA6_0(.din(n34088), .dout(n34091));
    jdff dff_A_lgumkYTG3_0(.din(n34085), .dout(n34088));
    jdff dff_A_cHwFbjZE0_0(.din(n34082), .dout(n34085));
    jdff dff_A_lRk8e8la5_0(.din(n34079), .dout(n34082));
    jdff dff_A_uNXe2iYU3_0(.din(n34076), .dout(n34079));
    jdff dff_A_vSOF2bZ24_0(.din(n34073), .dout(n34076));
    jdff dff_A_9F7A4NHn8_0(.din(n34070), .dout(n34073));
    jdff dff_A_D4aIypSf1_0(.din(n34067), .dout(n34070));
    jdff dff_A_jqnpxvNa9_0(.din(n34064), .dout(n34067));
    jdff dff_A_mmqCAwQQ0_0(.din(n34061), .dout(n34064));
    jdff dff_A_okMi2w5I6_2(.din(n3675), .dout(n34061));
    jdff dff_A_qTqooJ4g5_0(.din(n34055), .dout(G6123gat));
    jdff dff_A_ClIG4uEj0_0(.din(n34052), .dout(n34055));
    jdff dff_A_mc2ocRHi5_0(.din(n34049), .dout(n34052));
    jdff dff_A_edrMVVhI0_0(.din(n34046), .dout(n34049));
    jdff dff_A_NqQJ7Q9N7_0(.din(n34043), .dout(n34046));
    jdff dff_A_5sxAXsZZ2_0(.din(n34040), .dout(n34043));
    jdff dff_A_cBWohS1Z9_0(.din(n34037), .dout(n34040));
    jdff dff_A_WUnYuut38_0(.din(n34034), .dout(n34037));
    jdff dff_A_02Bq87UL8_0(.din(n34031), .dout(n34034));
    jdff dff_A_m86Z4tSp8_0(.din(n34028), .dout(n34031));
    jdff dff_A_TnokJ5nQ7_0(.din(n34025), .dout(n34028));
    jdff dff_A_hN7dwSJE8_0(.din(n34022), .dout(n34025));
    jdff dff_A_iKGDNwfx3_0(.din(n34019), .dout(n34022));
    jdff dff_A_8UlC83LO4_0(.din(n34016), .dout(n34019));
    jdff dff_A_86whUlow5_0(.din(n34013), .dout(n34016));
    jdff dff_A_kM3AliSJ6_0(.din(n34010), .dout(n34013));
    jdff dff_A_OhTY83Rd8_0(.din(n34007), .dout(n34010));
    jdff dff_A_Q8l7aJsV0_0(.din(n34004), .dout(n34007));
    jdff dff_A_keZsIW5T0_0(.din(n34001), .dout(n34004));
    jdff dff_A_29S28ue60_0(.din(n33998), .dout(n34001));
    jdff dff_A_PLOyHNKq5_0(.din(n33995), .dout(n33998));
    jdff dff_A_72D0u0by4_0(.din(n33992), .dout(n33995));
    jdff dff_A_woTG74pO7_0(.din(n33989), .dout(n33992));
    jdff dff_A_vrhsss888_0(.din(n33986), .dout(n33989));
    jdff dff_A_ieo9pNzn8_0(.din(n33983), .dout(n33986));
    jdff dff_A_ZlJw7U003_0(.din(n33980), .dout(n33983));
    jdff dff_A_zaboybat2_0(.din(n33977), .dout(n33980));
    jdff dff_A_RzkSdMIb4_0(.din(n33974), .dout(n33977));
    jdff dff_A_Xgwsrhnl1_0(.din(n33971), .dout(n33974));
    jdff dff_A_b9xSmEOi6_2(.din(n3271), .dout(n33971));
    jdff dff_A_QAAJOoP98_0(.din(n33965), .dout(G5971gat));
    jdff dff_A_kD19nGPu9_0(.din(n33962), .dout(n33965));
    jdff dff_A_rL6AXHc15_0(.din(n33959), .dout(n33962));
    jdff dff_A_K83xiXkF9_0(.din(n33956), .dout(n33959));
    jdff dff_A_hwYXCZVQ2_0(.din(n33953), .dout(n33956));
    jdff dff_A_B55TaYlr1_0(.din(n33950), .dout(n33953));
    jdff dff_A_nd2IUhhm0_0(.din(n33947), .dout(n33950));
    jdff dff_A_9s0IZ3cU9_0(.din(n33944), .dout(n33947));
    jdff dff_A_gilxwOXP8_0(.din(n33941), .dout(n33944));
    jdff dff_A_dCOIv1RO8_0(.din(n33938), .dout(n33941));
    jdff dff_A_OeX0mVef4_0(.din(n33935), .dout(n33938));
    jdff dff_A_BdpJywMH1_0(.din(n33932), .dout(n33935));
    jdff dff_A_IIEnOhAI5_0(.din(n33929), .dout(n33932));
    jdff dff_A_7m7ZrYDo0_0(.din(n33926), .dout(n33929));
    jdff dff_A_wfeZErTh7_0(.din(n33923), .dout(n33926));
    jdff dff_A_v2uaTy926_0(.din(n33920), .dout(n33923));
    jdff dff_A_fP7OT9lk4_0(.din(n33917), .dout(n33920));
    jdff dff_A_PNOJfyzw4_0(.din(n33914), .dout(n33917));
    jdff dff_A_0To7aDDQ0_0(.din(n33911), .dout(n33914));
    jdff dff_A_ujjTKTyt5_0(.din(n33908), .dout(n33911));
    jdff dff_A_vvzIJkBd2_0(.din(n33905), .dout(n33908));
    jdff dff_A_XwcQiECs5_0(.din(n33902), .dout(n33905));
    jdff dff_A_ztgUPg7q4_0(.din(n33899), .dout(n33902));
    jdff dff_A_w1ApzctC7_0(.din(n33896), .dout(n33899));
    jdff dff_A_tqQXvXDU0_0(.din(n33893), .dout(n33896));
    jdff dff_A_AFM0uJ5l6_0(.din(n33890), .dout(n33893));
    jdff dff_A_8uBpOEXy0_0(.din(n33887), .dout(n33890));
    jdff dff_A_we1nG2fK9_0(.din(n33884), .dout(n33887));
    jdff dff_A_034Fj5gR5_0(.din(n33881), .dout(n33884));
    jdff dff_A_Udra6jHd0_0(.din(n33878), .dout(n33881));
    jdff dff_A_3f80n6Gs2_0(.din(n33875), .dout(n33878));
    jdff dff_A_pqB8Fko46_0(.din(n33872), .dout(n33875));
    jdff dff_A_GrvPvRzD1_2(.din(n2879), .dout(n33872));
    jdff dff_A_6VkxC2es4_0(.din(n33866), .dout(G5672gat));
    jdff dff_A_iKzjfTVX4_0(.din(n33863), .dout(n33866));
    jdff dff_A_tjFBlMny9_0(.din(n33860), .dout(n33863));
    jdff dff_A_EgeqZIwH2_0(.din(n33857), .dout(n33860));
    jdff dff_A_zwpytITb0_0(.din(n33854), .dout(n33857));
    jdff dff_A_w16I4wIA3_0(.din(n33851), .dout(n33854));
    jdff dff_A_cJ2U47NJ9_0(.din(n33848), .dout(n33851));
    jdff dff_A_2CJ6JoJ82_0(.din(n33845), .dout(n33848));
    jdff dff_A_Dg9NJat15_0(.din(n33842), .dout(n33845));
    jdff dff_A_DDAQjcyZ1_0(.din(n33839), .dout(n33842));
    jdff dff_A_SHwyh0c18_0(.din(n33836), .dout(n33839));
    jdff dff_A_vw1RV2NV0_0(.din(n33833), .dout(n33836));
    jdff dff_A_7MN3KpQd6_0(.din(n33830), .dout(n33833));
    jdff dff_A_BphnsUee2_0(.din(n33827), .dout(n33830));
    jdff dff_A_9shebP5b4_0(.din(n33824), .dout(n33827));
    jdff dff_A_s7UaRNx12_0(.din(n33821), .dout(n33824));
    jdff dff_A_9VucbSb85_0(.din(n33818), .dout(n33821));
    jdff dff_A_yxNV3cxa8_0(.din(n33815), .dout(n33818));
    jdff dff_A_JlQ5wT8n6_0(.din(n33812), .dout(n33815));
    jdff dff_A_yy7jIqcN3_0(.din(n33809), .dout(n33812));
    jdff dff_A_bzvuPIrZ7_0(.din(n33806), .dout(n33809));
    jdff dff_A_h2AvVCpa7_0(.din(n33803), .dout(n33806));
    jdff dff_A_Q1tb5loz6_0(.din(n33800), .dout(n33803));
    jdff dff_A_p6E1KrtO2_0(.din(n33797), .dout(n33800));
    jdff dff_A_U4JsR3Uq9_0(.din(n33794), .dout(n33797));
    jdff dff_A_htZXRUfj3_0(.din(n33791), .dout(n33794));
    jdff dff_A_J9I248Jp1_0(.din(n33788), .dout(n33791));
    jdff dff_A_XRjeNN6X4_0(.din(n33785), .dout(n33788));
    jdff dff_A_u2yetZ701_0(.din(n33782), .dout(n33785));
    jdff dff_A_aZpy6ceA4_0(.din(n33779), .dout(n33782));
    jdff dff_A_EopLJP5f8_0(.din(n33776), .dout(n33779));
    jdff dff_A_3Pq8IOer9_0(.din(n33773), .dout(n33776));
    jdff dff_A_p0IlcEKG9_0(.din(n33770), .dout(n33773));
    jdff dff_A_fdPLxgoC7_0(.din(n33767), .dout(n33770));
    jdff dff_A_mdoLfKW24_0(.din(n33764), .dout(n33767));
    jdff dff_A_dSuBmHpc5_2(.din(n2501), .dout(n33764));
    jdff dff_A_IOeZXjCa0_0(.din(n33758), .dout(G5308gat));
    jdff dff_A_J77gEn0R7_0(.din(n33755), .dout(n33758));
    jdff dff_A_zlYlzgot0_0(.din(n33752), .dout(n33755));
    jdff dff_A_5JzA5IOY5_0(.din(n33749), .dout(n33752));
    jdff dff_A_uYc1LZQA9_0(.din(n33746), .dout(n33749));
    jdff dff_A_JfbYWNPY1_0(.din(n33743), .dout(n33746));
    jdff dff_A_CYdXihWS8_0(.din(n33740), .dout(n33743));
    jdff dff_A_BPTIuZLw0_0(.din(n33737), .dout(n33740));
    jdff dff_A_T5g9g3CF7_0(.din(n33734), .dout(n33737));
    jdff dff_A_EGGfkYTS7_0(.din(n33731), .dout(n33734));
    jdff dff_A_Hb5cXusa5_0(.din(n33728), .dout(n33731));
    jdff dff_A_dYamHiU94_0(.din(n33725), .dout(n33728));
    jdff dff_A_4k8yGm471_0(.din(n33722), .dout(n33725));
    jdff dff_A_wRVKJ3jY9_0(.din(n33719), .dout(n33722));
    jdff dff_A_KI8nbasE7_0(.din(n33716), .dout(n33719));
    jdff dff_A_jCTNTG1a6_0(.din(n33713), .dout(n33716));
    jdff dff_A_1QWCMiNR1_0(.din(n33710), .dout(n33713));
    jdff dff_A_GawTFX1o1_0(.din(n33707), .dout(n33710));
    jdff dff_A_8Kb0HGMS8_0(.din(n33704), .dout(n33707));
    jdff dff_A_fwwJw1VS2_0(.din(n33701), .dout(n33704));
    jdff dff_A_zowmw9a57_0(.din(n33698), .dout(n33701));
    jdff dff_A_AC60Ks0n6_0(.din(n33695), .dout(n33698));
    jdff dff_A_qZU0jvS74_0(.din(n33692), .dout(n33695));
    jdff dff_A_AbD197dt4_0(.din(n33689), .dout(n33692));
    jdff dff_A_phchnPF09_0(.din(n33686), .dout(n33689));
    jdff dff_A_ARnkUL2z7_0(.din(n33683), .dout(n33686));
    jdff dff_A_fBj8Bayd6_0(.din(n33680), .dout(n33683));
    jdff dff_A_7z4bE0cu6_0(.din(n33677), .dout(n33680));
    jdff dff_A_sSoUT4GB2_0(.din(n33674), .dout(n33677));
    jdff dff_A_Ifjcdlbu3_0(.din(n33671), .dout(n33674));
    jdff dff_A_GlRNSy3p5_0(.din(n33668), .dout(n33671));
    jdff dff_A_yw5RLx8R4_0(.din(n33665), .dout(n33668));
    jdff dff_A_hV3B999W1_0(.din(n33662), .dout(n33665));
    jdff dff_A_WA9QuyfT8_0(.din(n33659), .dout(n33662));
    jdff dff_A_42z0BhHr9_0(.din(n33656), .dout(n33659));
    jdff dff_A_JrxqGUmX7_0(.din(n33653), .dout(n33656));
    jdff dff_A_MjSvTIG88_0(.din(n33650), .dout(n33653));
    jdff dff_A_HZt5ri3T9_0(.din(n33647), .dout(n33650));
    jdff dff_A_Whz6y90z4_2(.din(n2150), .dout(n33647));
    jdff dff_A_akbihhF17_0(.din(n33641), .dout(G4946gat));
    jdff dff_A_CXuqsHmV8_0(.din(n33638), .dout(n33641));
    jdff dff_A_0SptStsj3_0(.din(n33635), .dout(n33638));
    jdff dff_A_J58U6LNq4_0(.din(n33632), .dout(n33635));
    jdff dff_A_JODvmQXA8_0(.din(n33629), .dout(n33632));
    jdff dff_A_DOBWTF6i9_0(.din(n33626), .dout(n33629));
    jdff dff_A_77moib451_0(.din(n33623), .dout(n33626));
    jdff dff_A_8zV5OEf07_0(.din(n33620), .dout(n33623));
    jdff dff_A_GmhKQyBS2_0(.din(n33617), .dout(n33620));
    jdff dff_A_Lw05cSSz2_0(.din(n33614), .dout(n33617));
    jdff dff_A_sbxqpdEo3_0(.din(n33611), .dout(n33614));
    jdff dff_A_iervmNT84_0(.din(n33608), .dout(n33611));
    jdff dff_A_RwfZcAnT6_0(.din(n33605), .dout(n33608));
    jdff dff_A_WoDYBINQ3_0(.din(n33602), .dout(n33605));
    jdff dff_A_V4m9BGio9_0(.din(n33599), .dout(n33602));
    jdff dff_A_l2OkezNQ1_0(.din(n33596), .dout(n33599));
    jdff dff_A_fgwJtztX6_0(.din(n33593), .dout(n33596));
    jdff dff_A_gc1VAXFE5_0(.din(n33590), .dout(n33593));
    jdff dff_A_HePwnezM4_0(.din(n33587), .dout(n33590));
    jdff dff_A_buRSM4VA9_0(.din(n33584), .dout(n33587));
    jdff dff_A_Nda5H63m0_0(.din(n33581), .dout(n33584));
    jdff dff_A_bsshSqi58_0(.din(n33578), .dout(n33581));
    jdff dff_A_D0caj4ux5_0(.din(n33575), .dout(n33578));
    jdff dff_A_Ov99oSIH4_0(.din(n33572), .dout(n33575));
    jdff dff_A_9lcWTbCJ1_0(.din(n33569), .dout(n33572));
    jdff dff_A_YzZJmEw44_0(.din(n33566), .dout(n33569));
    jdff dff_A_lpelPjES3_0(.din(n33563), .dout(n33566));
    jdff dff_A_S9hkccD34_0(.din(n33560), .dout(n33563));
    jdff dff_A_n7I5sYsL8_0(.din(n33557), .dout(n33560));
    jdff dff_A_J2rQYll28_0(.din(n33554), .dout(n33557));
    jdff dff_A_QcnA24mZ2_0(.din(n33551), .dout(n33554));
    jdff dff_A_Hrg1rnYa5_0(.din(n33548), .dout(n33551));
    jdff dff_A_5VnNimcs2_0(.din(n33545), .dout(n33548));
    jdff dff_A_UrPv5nGB4_0(.din(n33542), .dout(n33545));
    jdff dff_A_ljf05tGS0_0(.din(n33539), .dout(n33542));
    jdff dff_A_6aVrzrep2_0(.din(n33536), .dout(n33539));
    jdff dff_A_VZNs2JDX5_0(.din(n33533), .dout(n33536));
    jdff dff_A_XnWeIXQY3_0(.din(n33530), .dout(n33533));
    jdff dff_A_u11dQkLr8_0(.din(n33527), .dout(n33530));
    jdff dff_A_XL6evCQi0_0(.din(n33524), .dout(n33527));
    jdff dff_A_Aglkn81E6_0(.din(n33521), .dout(n33524));
    jdff dff_A_k3iKXLIe4_2(.din(n1826), .dout(n33521));
    jdff dff_A_sCnUazWe3_0(.din(n33515), .dout(G4591gat));
    jdff dff_A_uHFALARi1_0(.din(n33512), .dout(n33515));
    jdff dff_A_pIiXC78S0_0(.din(n33509), .dout(n33512));
    jdff dff_A_KlfMuHA29_0(.din(n33506), .dout(n33509));
    jdff dff_A_J7KP6UIZ4_0(.din(n33503), .dout(n33506));
    jdff dff_A_B3kiD3K41_0(.din(n33500), .dout(n33503));
    jdff dff_A_9vqiQXsy9_0(.din(n33497), .dout(n33500));
    jdff dff_A_ATFtiSAo6_0(.din(n33494), .dout(n33497));
    jdff dff_A_uMQoYzc75_0(.din(n33491), .dout(n33494));
    jdff dff_A_YZlIMUAR2_0(.din(n33488), .dout(n33491));
    jdff dff_A_y0kfxqN95_0(.din(n33485), .dout(n33488));
    jdff dff_A_RIlCVX171_0(.din(n33482), .dout(n33485));
    jdff dff_A_Z1MctO2O6_0(.din(n33479), .dout(n33482));
    jdff dff_A_tcKMdUFV7_0(.din(n33476), .dout(n33479));
    jdff dff_A_Sid51fXI9_0(.din(n33473), .dout(n33476));
    jdff dff_A_FySOt3Ij6_0(.din(n33470), .dout(n33473));
    jdff dff_A_IM87GUaO0_0(.din(n33467), .dout(n33470));
    jdff dff_A_T5LinO5h6_0(.din(n33464), .dout(n33467));
    jdff dff_A_SN8bqs2Q8_0(.din(n33461), .dout(n33464));
    jdff dff_A_nSqJEH3d4_0(.din(n33458), .dout(n33461));
    jdff dff_A_TECjVfwv6_0(.din(n33455), .dout(n33458));
    jdff dff_A_2UBEBqK12_0(.din(n33452), .dout(n33455));
    jdff dff_A_jgkdZ4zw3_0(.din(n33449), .dout(n33452));
    jdff dff_A_fQm5pxXj3_0(.din(n33446), .dout(n33449));
    jdff dff_A_JQlLSURC0_0(.din(n33443), .dout(n33446));
    jdff dff_A_9K9WqwCv8_0(.din(n33440), .dout(n33443));
    jdff dff_A_lhRRBONw1_0(.din(n33437), .dout(n33440));
    jdff dff_A_e9OojFyN1_0(.din(n33434), .dout(n33437));
    jdff dff_A_tsng1w7b9_0(.din(n33431), .dout(n33434));
    jdff dff_A_3Gxy1OxP4_0(.din(n33428), .dout(n33431));
    jdff dff_A_Ahq83ELf3_0(.din(n33425), .dout(n33428));
    jdff dff_A_gPMwZevJ4_0(.din(n33422), .dout(n33425));
    jdff dff_A_G3oFA62V3_0(.din(n33419), .dout(n33422));
    jdff dff_A_rC9QR0lC5_0(.din(n33416), .dout(n33419));
    jdff dff_A_obzNNO2M9_0(.din(n33413), .dout(n33416));
    jdff dff_A_GL7PML9S7_0(.din(n33410), .dout(n33413));
    jdff dff_A_aS2bhrfJ1_0(.din(n33407), .dout(n33410));
    jdff dff_A_h0g5HjaA9_0(.din(n33404), .dout(n33407));
    jdff dff_A_fLjFoE160_0(.din(n33401), .dout(n33404));
    jdff dff_A_jHmMc3Ki1_0(.din(n33398), .dout(n33401));
    jdff dff_A_fM681KaE7_0(.din(n33395), .dout(n33398));
    jdff dff_A_r8okHQLl2_0(.din(n33392), .dout(n33395));
    jdff dff_A_jTOenI3v4_0(.din(n33389), .dout(n33392));
    jdff dff_A_pXTROB3q9_0(.din(n33386), .dout(n33389));
    jdff dff_A_xANsDdVz6_2(.din(n1529), .dout(n33386));
    jdff dff_A_HLXQTx3j8_0(.din(n33380), .dout(G4241gat));
    jdff dff_A_YFPYsXl46_0(.din(n33377), .dout(n33380));
    jdff dff_A_LXNOeWHW9_0(.din(n33374), .dout(n33377));
    jdff dff_A_KXkzmyTm3_0(.din(n33371), .dout(n33374));
    jdff dff_A_yFAQckSv6_0(.din(n33368), .dout(n33371));
    jdff dff_A_v0BdXfzU6_0(.din(n33365), .dout(n33368));
    jdff dff_A_jWvUl0xN3_0(.din(n33362), .dout(n33365));
    jdff dff_A_1OeTwyEH9_0(.din(n33359), .dout(n33362));
    jdff dff_A_wuCqWLwH1_0(.din(n33356), .dout(n33359));
    jdff dff_A_SitAz65p3_0(.din(n33353), .dout(n33356));
    jdff dff_A_ahm8CCsf0_0(.din(n33350), .dout(n33353));
    jdff dff_A_46sTgkrF7_0(.din(n33347), .dout(n33350));
    jdff dff_A_hBewRon32_0(.din(n33344), .dout(n33347));
    jdff dff_A_HcBfl0mh6_0(.din(n33341), .dout(n33344));
    jdff dff_A_fioCgruU3_0(.din(n33338), .dout(n33341));
    jdff dff_A_fnJRMVzh6_0(.din(n33335), .dout(n33338));
    jdff dff_A_jVvIQzwF0_0(.din(n33332), .dout(n33335));
    jdff dff_A_ftGxvHZw6_0(.din(n33329), .dout(n33332));
    jdff dff_A_VXlBulOn1_0(.din(n33326), .dout(n33329));
    jdff dff_A_el1TYYkf6_0(.din(n33323), .dout(n33326));
    jdff dff_A_ffaHNuvX1_0(.din(n33320), .dout(n33323));
    jdff dff_A_HtpdOZjk3_0(.din(n33317), .dout(n33320));
    jdff dff_A_kIFd3SPK5_0(.din(n33314), .dout(n33317));
    jdff dff_A_ZcDslSaE2_0(.din(n33311), .dout(n33314));
    jdff dff_A_t339kxfb7_0(.din(n33308), .dout(n33311));
    jdff dff_A_ueVP981F2_0(.din(n33305), .dout(n33308));
    jdff dff_A_OWnu9flQ8_0(.din(n33302), .dout(n33305));
    jdff dff_A_sfwro9XK1_0(.din(n33299), .dout(n33302));
    jdff dff_A_lTAA7f5n6_0(.din(n33296), .dout(n33299));
    jdff dff_A_3R3qCcjJ9_0(.din(n33293), .dout(n33296));
    jdff dff_A_Rz9JcqBr3_0(.din(n33290), .dout(n33293));
    jdff dff_A_AdmSjIPk7_0(.din(n33287), .dout(n33290));
    jdff dff_A_S5XawaYp1_0(.din(n33284), .dout(n33287));
    jdff dff_A_T2pNZOI31_0(.din(n33281), .dout(n33284));
    jdff dff_A_BtXZHzpo6_0(.din(n33278), .dout(n33281));
    jdff dff_A_p8WJsDxe2_0(.din(n33275), .dout(n33278));
    jdff dff_A_Lerj2lpD7_0(.din(n33272), .dout(n33275));
    jdff dff_A_2eYmAzvl3_0(.din(n33269), .dout(n33272));
    jdff dff_A_WJWPnB9Q8_0(.din(n33266), .dout(n33269));
    jdff dff_A_H1MTa1pn2_0(.din(n33263), .dout(n33266));
    jdff dff_A_HYrZCvr05_0(.din(n33260), .dout(n33263));
    jdff dff_A_YZwxnTFa8_0(.din(n33257), .dout(n33260));
    jdff dff_A_liYaWvap4_0(.din(n33254), .dout(n33257));
    jdff dff_A_nE69rSCD7_0(.din(n33251), .dout(n33254));
    jdff dff_A_kG6bMXmL9_0(.din(n33248), .dout(n33251));
    jdff dff_A_f8dCr8qN6_0(.din(n33245), .dout(n33248));
    jdff dff_A_wCy1wkOG8_0(.din(n33242), .dout(n33245));
    jdff dff_A_rFD3ruyP8_2(.din(n1259), .dout(n33242));
    jdff dff_A_pWkdBPgJ1_0(.din(n33236), .dout(G3895gat));
    jdff dff_A_yKbQ2N8Z4_0(.din(n33233), .dout(n33236));
    jdff dff_A_cd5jhFgd7_0(.din(n33230), .dout(n33233));
    jdff dff_A_nbbZbNnd3_0(.din(n33227), .dout(n33230));
    jdff dff_A_ksiK7KtB0_0(.din(n33224), .dout(n33227));
    jdff dff_A_IBHNEwXx5_0(.din(n33221), .dout(n33224));
    jdff dff_A_PzDEvjIy5_0(.din(n33218), .dout(n33221));
    jdff dff_A_2Jk1u5j47_0(.din(n33215), .dout(n33218));
    jdff dff_A_q1dML4Pk2_0(.din(n33212), .dout(n33215));
    jdff dff_A_JaRRQPGI6_0(.din(n33209), .dout(n33212));
    jdff dff_A_fum6iNeP8_0(.din(n33206), .dout(n33209));
    jdff dff_A_IBxT8tdI5_0(.din(n33203), .dout(n33206));
    jdff dff_A_ppQja7TY5_0(.din(n33200), .dout(n33203));
    jdff dff_A_EmEDWUDA7_0(.din(n33197), .dout(n33200));
    jdff dff_A_IcrTRLzk1_0(.din(n33194), .dout(n33197));
    jdff dff_A_emgBjAc66_0(.din(n33191), .dout(n33194));
    jdff dff_A_d4PDu5js1_0(.din(n33188), .dout(n33191));
    jdff dff_A_fvZktCYV2_0(.din(n33185), .dout(n33188));
    jdff dff_A_0W8NKevD2_0(.din(n33182), .dout(n33185));
    jdff dff_A_8aYcfREe7_0(.din(n33179), .dout(n33182));
    jdff dff_A_dbNCtryU3_0(.din(n33176), .dout(n33179));
    jdff dff_A_HcoYOmkU1_0(.din(n33173), .dout(n33176));
    jdff dff_A_c87I8tIR1_0(.din(n33170), .dout(n33173));
    jdff dff_A_jyS6FEhA3_0(.din(n33167), .dout(n33170));
    jdff dff_A_Q3yKlTyM2_0(.din(n33164), .dout(n33167));
    jdff dff_A_FciaFmtN9_0(.din(n33161), .dout(n33164));
    jdff dff_A_h48HmMfn9_0(.din(n33158), .dout(n33161));
    jdff dff_A_pqKVAr1L2_0(.din(n33155), .dout(n33158));
    jdff dff_A_EDcfrQLi4_0(.din(n33152), .dout(n33155));
    jdff dff_A_MQ0iiGvh3_0(.din(n33149), .dout(n33152));
    jdff dff_A_UvrOH25s6_0(.din(n33146), .dout(n33149));
    jdff dff_A_5g1JbNwe1_0(.din(n33143), .dout(n33146));
    jdff dff_A_MvOEAy0u1_0(.din(n33140), .dout(n33143));
    jdff dff_A_UMl2PSNY9_0(.din(n33137), .dout(n33140));
    jdff dff_A_AYNaDx281_0(.din(n33134), .dout(n33137));
    jdff dff_A_EoZBtHPh3_0(.din(n33131), .dout(n33134));
    jdff dff_A_EGwqlcHe5_0(.din(n33128), .dout(n33131));
    jdff dff_A_KD3YEOd65_0(.din(n33125), .dout(n33128));
    jdff dff_A_pYQCQtA32_0(.din(n33122), .dout(n33125));
    jdff dff_A_PNytZXnZ6_0(.din(n33119), .dout(n33122));
    jdff dff_A_o7mc7g1c8_0(.din(n33116), .dout(n33119));
    jdff dff_A_7nhZJRs75_0(.din(n33113), .dout(n33116));
    jdff dff_A_19AlYVxb6_0(.din(n33110), .dout(n33113));
    jdff dff_A_ubCCc7Ut7_0(.din(n33107), .dout(n33110));
    jdff dff_A_46XjdZOD8_0(.din(n33104), .dout(n33107));
    jdff dff_A_ztwIVD195_0(.din(n33101), .dout(n33104));
    jdff dff_A_zBD61QgE5_0(.din(n33098), .dout(n33101));
    jdff dff_A_76c5jxDK0_0(.din(n33095), .dout(n33098));
    jdff dff_A_tEARLD7D6_0(.din(n33092), .dout(n33095));
    jdff dff_A_D1ljxla53_0(.din(n33089), .dout(n33092));
    jdff dff_A_fdK3GZD42_2(.din(n1019), .dout(n33089));
    jdff dff_A_uZFEBlv00_0(.din(n33083), .dout(G3552gat));
    jdff dff_A_RaSdH8Ma7_0(.din(n33080), .dout(n33083));
    jdff dff_A_N1CbjniU6_0(.din(n33077), .dout(n33080));
    jdff dff_A_0NeDqDHN7_0(.din(n33074), .dout(n33077));
    jdff dff_A_c2T70DH62_0(.din(n33071), .dout(n33074));
    jdff dff_A_7uhaWb3b0_0(.din(n33068), .dout(n33071));
    jdff dff_A_Xhq0SttG8_0(.din(n33065), .dout(n33068));
    jdff dff_A_KJnPgomu6_0(.din(n33062), .dout(n33065));
    jdff dff_A_mhy64e4S5_0(.din(n33059), .dout(n33062));
    jdff dff_A_IAwfR51o0_0(.din(n33056), .dout(n33059));
    jdff dff_A_nCyqUpG01_0(.din(n33053), .dout(n33056));
    jdff dff_A_cTzWC01n7_0(.din(n33050), .dout(n33053));
    jdff dff_A_CI30zncL7_0(.din(n33047), .dout(n33050));
    jdff dff_A_XzN1SUH75_0(.din(n33044), .dout(n33047));
    jdff dff_A_BTqd9MWm2_0(.din(n33041), .dout(n33044));
    jdff dff_A_7gmrsr0L6_0(.din(n33038), .dout(n33041));
    jdff dff_A_2EloxUDu8_0(.din(n33035), .dout(n33038));
    jdff dff_A_Mo7K6gIZ5_0(.din(n33032), .dout(n33035));
    jdff dff_A_48kgtEq73_0(.din(n33029), .dout(n33032));
    jdff dff_A_ubRN5I0d2_0(.din(n33026), .dout(n33029));
    jdff dff_A_5xZ55Ezy0_0(.din(n33023), .dout(n33026));
    jdff dff_A_DFFZ0xWL5_0(.din(n33020), .dout(n33023));
    jdff dff_A_btiNppzx2_0(.din(n33017), .dout(n33020));
    jdff dff_A_DRa0OLxR4_0(.din(n33014), .dout(n33017));
    jdff dff_A_Wc3AONrK4_0(.din(n33011), .dout(n33014));
    jdff dff_A_GLZ5Xeui5_0(.din(n33008), .dout(n33011));
    jdff dff_A_J0AoCJDc7_0(.din(n33005), .dout(n33008));
    jdff dff_A_w36IsMES2_0(.din(n33002), .dout(n33005));
    jdff dff_A_vnxznyvI0_0(.din(n32999), .dout(n33002));
    jdff dff_A_8kmJIDCC6_0(.din(n32996), .dout(n32999));
    jdff dff_A_rfc8MkMO1_0(.din(n32993), .dout(n32996));
    jdff dff_A_UAPm7bfk6_0(.din(n32990), .dout(n32993));
    jdff dff_A_RN94JaGJ7_0(.din(n32987), .dout(n32990));
    jdff dff_A_1QJpCATX3_0(.din(n32984), .dout(n32987));
    jdff dff_A_swYR5ZIm2_0(.din(n32981), .dout(n32984));
    jdff dff_A_V79hsKxC5_0(.din(n32978), .dout(n32981));
    jdff dff_A_2gmMJMzL1_0(.din(n32975), .dout(n32978));
    jdff dff_A_zgdFauPo1_0(.din(n32972), .dout(n32975));
    jdff dff_A_dFA43SZV8_0(.din(n32969), .dout(n32972));
    jdff dff_A_ONKKmu3q0_0(.din(n32966), .dout(n32969));
    jdff dff_A_vspatCTH4_0(.din(n32963), .dout(n32966));
    jdff dff_A_V3wRKQ6T0_0(.din(n32960), .dout(n32963));
    jdff dff_A_C6QyKAcU4_0(.din(n32957), .dout(n32960));
    jdff dff_A_pln3Ak7p8_0(.din(n32954), .dout(n32957));
    jdff dff_A_88CXVLny9_0(.din(n32951), .dout(n32954));
    jdff dff_A_kPlYeg6T3_0(.din(n32948), .dout(n32951));
    jdff dff_A_QqVaIVsn3_0(.din(n32945), .dout(n32948));
    jdff dff_A_hahDbAXu3_0(.din(n32942), .dout(n32945));
    jdff dff_A_TEWSREFY8_0(.din(n32939), .dout(n32942));
    jdff dff_A_NkTNLiv69_0(.din(n32936), .dout(n32939));
    jdff dff_A_yV6upp311_0(.din(n32933), .dout(n32936));
    jdff dff_A_WC9m3MTH6_0(.din(n32930), .dout(n32933));
    jdff dff_A_HPUO8x400_0(.din(n32927), .dout(n32930));
    jdff dff_A_1S7EK9uC0_2(.din(n806), .dout(n32927));
    jdff dff_A_68phYQ4d9_0(.din(n32921), .dout(G3211gat));
    jdff dff_A_9mk7is8K3_0(.din(n32918), .dout(n32921));
    jdff dff_A_DcnzQsiz7_0(.din(n32915), .dout(n32918));
    jdff dff_A_r47pQr0d3_0(.din(n32912), .dout(n32915));
    jdff dff_A_i15bLFzL8_0(.din(n32909), .dout(n32912));
    jdff dff_A_Aj89iEXp0_0(.din(n32906), .dout(n32909));
    jdff dff_A_S5aMvSkZ1_0(.din(n32903), .dout(n32906));
    jdff dff_A_tTPD9ViQ9_0(.din(n32900), .dout(n32903));
    jdff dff_A_ySqeQT9u0_0(.din(n32897), .dout(n32900));
    jdff dff_A_uAUxLrQH5_0(.din(n32894), .dout(n32897));
    jdff dff_A_yjXakVSd2_0(.din(n32891), .dout(n32894));
    jdff dff_A_zOl2rtiz9_0(.din(n32888), .dout(n32891));
    jdff dff_A_3Wp3jCBv0_0(.din(n32885), .dout(n32888));
    jdff dff_A_BfQIop7N9_0(.din(n32882), .dout(n32885));
    jdff dff_A_PfzGn3X40_0(.din(n32879), .dout(n32882));
    jdff dff_A_Pwa9WOzs5_0(.din(n32876), .dout(n32879));
    jdff dff_A_XuZzfXVF6_0(.din(n32873), .dout(n32876));
    jdff dff_A_8oG1HlPz7_0(.din(n32870), .dout(n32873));
    jdff dff_A_SxpUWssj6_0(.din(n32867), .dout(n32870));
    jdff dff_A_Q3nwZ8B10_0(.din(n32864), .dout(n32867));
    jdff dff_A_v1i21oW54_0(.din(n32861), .dout(n32864));
    jdff dff_A_Xxxmtu9M9_0(.din(n32858), .dout(n32861));
    jdff dff_A_pDxQtBqK4_0(.din(n32855), .dout(n32858));
    jdff dff_A_Z8m1LNur4_0(.din(n32852), .dout(n32855));
    jdff dff_A_TiiRIfM07_0(.din(n32849), .dout(n32852));
    jdff dff_A_zW3StyU38_0(.din(n32846), .dout(n32849));
    jdff dff_A_PYTHsVSV6_0(.din(n32843), .dout(n32846));
    jdff dff_A_EqIcwaNl4_0(.din(n32840), .dout(n32843));
    jdff dff_A_cMnCFvqz6_0(.din(n32837), .dout(n32840));
    jdff dff_A_rTm3ETE66_0(.din(n32834), .dout(n32837));
    jdff dff_A_wRWZrKDl9_0(.din(n32831), .dout(n32834));
    jdff dff_A_VnGbh9Xj3_0(.din(n32828), .dout(n32831));
    jdff dff_A_94PULiMl6_0(.din(n32825), .dout(n32828));
    jdff dff_A_Y45WbqMa1_0(.din(n32822), .dout(n32825));
    jdff dff_A_d9dXtT5D1_0(.din(n32819), .dout(n32822));
    jdff dff_A_6Klz3CAM9_0(.din(n32816), .dout(n32819));
    jdff dff_A_3GNKu7tj4_0(.din(n32813), .dout(n32816));
    jdff dff_A_ocPFOu4n9_0(.din(n32810), .dout(n32813));
    jdff dff_A_uXKjIZUZ8_0(.din(n32807), .dout(n32810));
    jdff dff_A_dlri9R6W5_0(.din(n32804), .dout(n32807));
    jdff dff_A_R16Af9wA2_0(.din(n32801), .dout(n32804));
    jdff dff_A_8NgEBRJE8_0(.din(n32798), .dout(n32801));
    jdff dff_A_2KUCl9DI3_0(.din(n32795), .dout(n32798));
    jdff dff_A_EAgXLHIO1_0(.din(n32792), .dout(n32795));
    jdff dff_A_KINI6req8_0(.din(n32789), .dout(n32792));
    jdff dff_A_AGXvGq6D7_0(.din(n32786), .dout(n32789));
    jdff dff_A_vxA7COBK1_0(.din(n32783), .dout(n32786));
    jdff dff_A_bSzpXqiR9_0(.din(n32780), .dout(n32783));
    jdff dff_A_gKZFgW2Y3_0(.din(n32777), .dout(n32780));
    jdff dff_A_1nyx4VDY1_0(.din(n32774), .dout(n32777));
    jdff dff_A_OOkiQ2DN0_0(.din(n32771), .dout(n32774));
    jdff dff_A_RMJAOgWq7_0(.din(n32768), .dout(n32771));
    jdff dff_A_ijIFejDa8_0(.din(n32765), .dout(n32768));
    jdff dff_A_22qSoX7d0_0(.din(n32762), .dout(n32765));
    jdff dff_A_m3ufP3LF0_0(.din(n32759), .dout(n32762));
    jdff dff_A_6iTRBODh0_0(.din(n32756), .dout(n32759));
    jdff dff_A_fzty24Fg7_2(.din(n620), .dout(n32756));
    jdff dff_A_V5ARinu60_0(.din(n32750), .dout(G2877gat));
    jdff dff_A_PIQxSxvV7_0(.din(n32747), .dout(n32750));
    jdff dff_A_jMtAlfG86_0(.din(n32744), .dout(n32747));
    jdff dff_A_gffDqlbO2_0(.din(n32741), .dout(n32744));
    jdff dff_A_ZcD82bRK2_0(.din(n32738), .dout(n32741));
    jdff dff_A_D67H8ryT4_0(.din(n32735), .dout(n32738));
    jdff dff_A_VDOZAGKJ3_0(.din(n32732), .dout(n32735));
    jdff dff_A_33pAvLiG4_0(.din(n32729), .dout(n32732));
    jdff dff_A_IRQLmgfl1_0(.din(n32726), .dout(n32729));
    jdff dff_A_C3F1ytOH2_0(.din(n32723), .dout(n32726));
    jdff dff_A_2stJmJAI3_0(.din(n32720), .dout(n32723));
    jdff dff_A_X2xmfMcN5_0(.din(n32717), .dout(n32720));
    jdff dff_A_Ah9bIosR8_0(.din(n32714), .dout(n32717));
    jdff dff_A_diZSij045_0(.din(n32711), .dout(n32714));
    jdff dff_A_q5LOD2tg7_0(.din(n32708), .dout(n32711));
    jdff dff_A_XSaSblFD4_0(.din(n32705), .dout(n32708));
    jdff dff_A_UbCLgaYO7_0(.din(n32702), .dout(n32705));
    jdff dff_A_gajrwyFc3_0(.din(n32699), .dout(n32702));
    jdff dff_A_pajuTJ4l9_0(.din(n32696), .dout(n32699));
    jdff dff_A_LcacxyjB4_0(.din(n32693), .dout(n32696));
    jdff dff_A_lzbFtxis8_0(.din(n32690), .dout(n32693));
    jdff dff_A_wWWm1iD94_0(.din(n32687), .dout(n32690));
    jdff dff_A_mKHUZWye9_0(.din(n32684), .dout(n32687));
    jdff dff_A_XMy9xEqY6_0(.din(n32681), .dout(n32684));
    jdff dff_A_0UJhvR7F7_0(.din(n32678), .dout(n32681));
    jdff dff_A_So9rCyCz4_0(.din(n32675), .dout(n32678));
    jdff dff_A_X3aSuwpr7_0(.din(n32672), .dout(n32675));
    jdff dff_A_lIMMJ4mF0_0(.din(n32669), .dout(n32672));
    jdff dff_A_dQW0Y0CM0_0(.din(n32666), .dout(n32669));
    jdff dff_A_8ctyCZPs9_0(.din(n32663), .dout(n32666));
    jdff dff_A_JpKvjN0Q8_0(.din(n32660), .dout(n32663));
    jdff dff_A_3ohWSRwp6_0(.din(n32657), .dout(n32660));
    jdff dff_A_MDG60FCl4_0(.din(n32654), .dout(n32657));
    jdff dff_A_vCbl7ueO9_0(.din(n32651), .dout(n32654));
    jdff dff_A_xRpkV9632_0(.din(n32648), .dout(n32651));
    jdff dff_A_pqHE9Al20_0(.din(n32645), .dout(n32648));
    jdff dff_A_lEqnh4SU5_0(.din(n32642), .dout(n32645));
    jdff dff_A_npCZH30I8_0(.din(n32639), .dout(n32642));
    jdff dff_A_15wk6lWG7_0(.din(n32636), .dout(n32639));
    jdff dff_A_bLq4l5x63_0(.din(n32633), .dout(n32636));
    jdff dff_A_6S5w8DWx4_0(.din(n32630), .dout(n32633));
    jdff dff_A_NSmRaWpA6_0(.din(n32627), .dout(n32630));
    jdff dff_A_BXAf8yXK6_0(.din(n32624), .dout(n32627));
    jdff dff_A_2MQGX1sc5_0(.din(n32621), .dout(n32624));
    jdff dff_A_K7xAnZbI1_0(.din(n32618), .dout(n32621));
    jdff dff_A_AH7xB5E76_0(.din(n32615), .dout(n32618));
    jdff dff_A_7tYKSSNk7_0(.din(n32612), .dout(n32615));
    jdff dff_A_CIi0AJt59_0(.din(n32609), .dout(n32612));
    jdff dff_A_05M9lXxp1_0(.din(n32606), .dout(n32609));
    jdff dff_A_hmCun4bB8_0(.din(n32603), .dout(n32606));
    jdff dff_A_0B793M7y4_0(.din(n32600), .dout(n32603));
    jdff dff_A_alVAfPKn5_0(.din(n32597), .dout(n32600));
    jdff dff_A_bo9Idjg63_0(.din(n32594), .dout(n32597));
    jdff dff_A_FF4UYeuX9_0(.din(n32591), .dout(n32594));
    jdff dff_A_CQnTGkZN9_0(.din(n32588), .dout(n32591));
    jdff dff_A_QwIXjRXM8_0(.din(n32585), .dout(n32588));
    jdff dff_A_zwrkMT7A1_0(.din(n32582), .dout(n32585));
    jdff dff_A_QQtvKVR79_0(.din(n32579), .dout(n32582));
    jdff dff_A_nscWjhLV4_0(.din(n32576), .dout(n32579));
    jdff dff_A_4JhpDJQk1_2(.din(n461), .dout(n32576));
    jdff dff_A_YIn3qLDg7_0(.din(n32570), .dout(G2548gat));
    jdff dff_A_x5RKSedm6_0(.din(n32567), .dout(n32570));
    jdff dff_A_Z8lnYFP37_0(.din(n32564), .dout(n32567));
    jdff dff_A_8ZFaHYJb2_0(.din(n32561), .dout(n32564));
    jdff dff_A_IgrKJTUo6_0(.din(n32558), .dout(n32561));
    jdff dff_A_7WfemrKq0_0(.din(n32555), .dout(n32558));
    jdff dff_A_iVSpAhTK7_0(.din(n32552), .dout(n32555));
    jdff dff_A_v01lq88z1_0(.din(n32549), .dout(n32552));
    jdff dff_A_aODrlKhT3_0(.din(n32546), .dout(n32549));
    jdff dff_A_wtIb7jUO1_0(.din(n32543), .dout(n32546));
    jdff dff_A_dbq52p2K5_0(.din(n32540), .dout(n32543));
    jdff dff_A_vGJVRWXF6_0(.din(n32537), .dout(n32540));
    jdff dff_A_zQLlC5Jg5_0(.din(n32534), .dout(n32537));
    jdff dff_A_ej3NMY796_0(.din(n32531), .dout(n32534));
    jdff dff_A_MiTYFQNb2_0(.din(n32528), .dout(n32531));
    jdff dff_A_Hy0Ia5YF8_0(.din(n32525), .dout(n32528));
    jdff dff_A_xLl8ZBKx4_0(.din(n32522), .dout(n32525));
    jdff dff_A_cKcQoA330_0(.din(n32519), .dout(n32522));
    jdff dff_A_UaAQEaEB1_0(.din(n32516), .dout(n32519));
    jdff dff_A_EDJQ5LCw3_0(.din(n32513), .dout(n32516));
    jdff dff_A_KHz6G9TZ1_0(.din(n32510), .dout(n32513));
    jdff dff_A_I40QanF71_0(.din(n32507), .dout(n32510));
    jdff dff_A_fbPW6fY64_0(.din(n32504), .dout(n32507));
    jdff dff_A_WdTMREwU5_0(.din(n32501), .dout(n32504));
    jdff dff_A_kQuEI4zD7_0(.din(n32498), .dout(n32501));
    jdff dff_A_fK22dD7y6_0(.din(n32495), .dout(n32498));
    jdff dff_A_tExBP91x7_0(.din(n32492), .dout(n32495));
    jdff dff_A_NJuuxCSy0_0(.din(n32489), .dout(n32492));
    jdff dff_A_8ObDaeqV8_0(.din(n32486), .dout(n32489));
    jdff dff_A_IS1vNVL88_0(.din(n32483), .dout(n32486));
    jdff dff_A_rV90dYuF4_0(.din(n32480), .dout(n32483));
    jdff dff_A_fcy7mX9L5_0(.din(n32477), .dout(n32480));
    jdff dff_A_cYohB2Ig3_0(.din(n32474), .dout(n32477));
    jdff dff_A_nValV1yi1_0(.din(n32471), .dout(n32474));
    jdff dff_A_IOKbtvmm5_0(.din(n32468), .dout(n32471));
    jdff dff_A_vi7yjqHw6_0(.din(n32465), .dout(n32468));
    jdff dff_A_2XcVAt7h1_0(.din(n32462), .dout(n32465));
    jdff dff_A_aVzL60u73_0(.din(n32459), .dout(n32462));
    jdff dff_A_Zuq8soWV9_0(.din(n32456), .dout(n32459));
    jdff dff_A_KPqNtckk9_0(.din(n32453), .dout(n32456));
    jdff dff_A_UJpwuqi06_0(.din(n32450), .dout(n32453));
    jdff dff_A_X8hL8fkt7_0(.din(n32447), .dout(n32450));
    jdff dff_A_KwVgtCfR3_0(.din(n32444), .dout(n32447));
    jdff dff_A_O1FQhSMu2_0(.din(n32441), .dout(n32444));
    jdff dff_A_xY2YEdT17_0(.din(n32438), .dout(n32441));
    jdff dff_A_vDpKBRS55_0(.din(n32435), .dout(n32438));
    jdff dff_A_5n9ZpK7C5_0(.din(n32432), .dout(n32435));
    jdff dff_A_EErckhbs1_0(.din(n32429), .dout(n32432));
    jdff dff_A_BHdxHAt01_0(.din(n32426), .dout(n32429));
    jdff dff_A_kTaoyh0S4_0(.din(n32423), .dout(n32426));
    jdff dff_A_yIzZqKfb5_0(.din(n32420), .dout(n32423));
    jdff dff_A_w4Aj6XlB2_0(.din(n32417), .dout(n32420));
    jdff dff_A_pFZUHEKQ7_0(.din(n32414), .dout(n32417));
    jdff dff_A_ABzoDVs39_0(.din(n32411), .dout(n32414));
    jdff dff_A_pRcNIFEJ4_0(.din(n32408), .dout(n32411));
    jdff dff_A_U5OLYsr97_0(.din(n32405), .dout(n32408));
    jdff dff_A_9QY3BGhr5_0(.din(n32402), .dout(n32405));
    jdff dff_A_5waJCCo93_0(.din(n32399), .dout(n32402));
    jdff dff_A_oTtkERGX3_0(.din(n32396), .dout(n32399));
    jdff dff_A_qRfJJhsW8_0(.din(n32393), .dout(n32396));
    jdff dff_A_yy540UXo8_0(.din(n32390), .dout(n32393));
    jdff dff_A_DWMixp4U9_0(.din(n32387), .dout(n32390));
    jdff dff_A_gefk1wav5_2(.din(n329), .dout(n32387));
    jdff dff_A_7yE0NEGK3_0(.din(n32381), .dout(G2223gat));
    jdff dff_A_O6hg4Dry9_0(.din(n32378), .dout(n32381));
    jdff dff_A_vjiFzC1H3_0(.din(n32375), .dout(n32378));
    jdff dff_A_SbpdLbA98_0(.din(n32372), .dout(n32375));
    jdff dff_A_D98vrOpP9_0(.din(n32369), .dout(n32372));
    jdff dff_A_HXAkp2Hr2_0(.din(n32366), .dout(n32369));
    jdff dff_A_48zxiKJh3_0(.din(n32363), .dout(n32366));
    jdff dff_A_XNimF5mI3_0(.din(n32360), .dout(n32363));
    jdff dff_A_Lo4r26GP1_0(.din(n32357), .dout(n32360));
    jdff dff_A_RZtG7oBe2_0(.din(n32354), .dout(n32357));
    jdff dff_A_LS7bFTju7_0(.din(n32351), .dout(n32354));
    jdff dff_A_sqbHbFPC4_0(.din(n32348), .dout(n32351));
    jdff dff_A_MZG1aCZA7_0(.din(n32345), .dout(n32348));
    jdff dff_A_waG2YfAb8_0(.din(n32342), .dout(n32345));
    jdff dff_A_8WYA2Jd19_0(.din(n32339), .dout(n32342));
    jdff dff_A_6Ljx9aGY4_0(.din(n32336), .dout(n32339));
    jdff dff_A_i29UEyo96_0(.din(n32333), .dout(n32336));
    jdff dff_A_merpgjMT5_0(.din(n32330), .dout(n32333));
    jdff dff_A_C84v9WI28_0(.din(n32327), .dout(n32330));
    jdff dff_A_KPVd0E3G7_0(.din(n32324), .dout(n32327));
    jdff dff_A_7ao35V7m9_0(.din(n32321), .dout(n32324));
    jdff dff_A_vL4YCkmB6_0(.din(n32318), .dout(n32321));
    jdff dff_A_YsSHIPp28_0(.din(n32315), .dout(n32318));
    jdff dff_A_urcuM0of9_0(.din(n32312), .dout(n32315));
    jdff dff_A_pBRyccUm1_0(.din(n32309), .dout(n32312));
    jdff dff_A_XvVgFn9P0_0(.din(n32306), .dout(n32309));
    jdff dff_A_yWsc2FG58_0(.din(n32303), .dout(n32306));
    jdff dff_A_79qyOkIc4_0(.din(n32300), .dout(n32303));
    jdff dff_A_adCT9SwV1_0(.din(n32297), .dout(n32300));
    jdff dff_A_Sr626VtM9_0(.din(n32294), .dout(n32297));
    jdff dff_A_y9xN8TYu4_0(.din(n32291), .dout(n32294));
    jdff dff_A_u0gJUiq52_0(.din(n32288), .dout(n32291));
    jdff dff_A_mSmIWK7j9_0(.din(n32285), .dout(n32288));
    jdff dff_A_OO8pCVS49_0(.din(n32282), .dout(n32285));
    jdff dff_A_mpJjQPkg4_0(.din(n32279), .dout(n32282));
    jdff dff_A_6VIPgpEI3_0(.din(n32276), .dout(n32279));
    jdff dff_A_htM5lZks8_0(.din(n32273), .dout(n32276));
    jdff dff_A_i74p85CP1_0(.din(n32270), .dout(n32273));
    jdff dff_A_shQg4kMP0_0(.din(n32267), .dout(n32270));
    jdff dff_A_0VBGkh5x9_0(.din(n32264), .dout(n32267));
    jdff dff_A_iSUWP2vl4_0(.din(n32261), .dout(n32264));
    jdff dff_A_liEFXoqg6_0(.din(n32258), .dout(n32261));
    jdff dff_A_Lp23YidW0_0(.din(n32255), .dout(n32258));
    jdff dff_A_jIfjbs3p4_0(.din(n32252), .dout(n32255));
    jdff dff_A_qez06FdT3_0(.din(n32249), .dout(n32252));
    jdff dff_A_65S7st0f9_0(.din(n32246), .dout(n32249));
    jdff dff_A_44b5Za3q0_0(.din(n32243), .dout(n32246));
    jdff dff_A_LkTXmiTN2_0(.din(n32240), .dout(n32243));
    jdff dff_A_R5d8JNCG8_0(.din(n32237), .dout(n32240));
    jdff dff_A_VoeJeHDR0_0(.din(n32234), .dout(n32237));
    jdff dff_A_sANRdrOi4_0(.din(n32231), .dout(n32234));
    jdff dff_A_n0dU0Hwf3_0(.din(n32228), .dout(n32231));
    jdff dff_A_mEgezkWX4_0(.din(n32225), .dout(n32228));
    jdff dff_A_Ytp4l8vM7_0(.din(n32222), .dout(n32225));
    jdff dff_A_3ho92WB04_0(.din(n32219), .dout(n32222));
    jdff dff_A_0sdC5CQt8_0(.din(n32216), .dout(n32219));
    jdff dff_A_hmRtgyuR3_0(.din(n32213), .dout(n32216));
    jdff dff_A_T7K3CaY87_0(.din(n32210), .dout(n32213));
    jdff dff_A_M7REda1w2_0(.din(n32207), .dout(n32210));
    jdff dff_A_DL4jujl76_0(.din(n32204), .dout(n32207));
    jdff dff_A_DJaz2nfu9_0(.din(n32201), .dout(n32204));
    jdff dff_A_KceAzcYC0_0(.din(n32198), .dout(n32201));
    jdff dff_A_ItSyCivU4_0(.din(n32195), .dout(n32198));
    jdff dff_A_aAxv4qMc1_0(.din(n32192), .dout(n32195));
    jdff dff_A_w7Qg4Ogm6_0(.din(n32189), .dout(n32192));
    jdff dff_A_dMBLpPmk9_2(.din(n220), .dout(n32189));
    jdff dff_A_5QNzbAT64_0(.din(n32183), .dout(G1901gat));
    jdff dff_A_vUbw6a1X3_0(.din(n32180), .dout(n32183));
    jdff dff_A_yyGiPMnY0_0(.din(n32177), .dout(n32180));
    jdff dff_A_yKS96IHA5_0(.din(n32174), .dout(n32177));
    jdff dff_A_DHpCUB6Q1_0(.din(n32171), .dout(n32174));
    jdff dff_A_ZI9Vowwm3_0(.din(n32168), .dout(n32171));
    jdff dff_A_U6lDBDTs0_0(.din(n32165), .dout(n32168));
    jdff dff_A_wGpiu0r74_0(.din(n32162), .dout(n32165));
    jdff dff_A_c4TVz89o2_0(.din(n32159), .dout(n32162));
    jdff dff_A_paKgfGkd1_0(.din(n32156), .dout(n32159));
    jdff dff_A_MdHWVO2B3_0(.din(n32153), .dout(n32156));
    jdff dff_A_O0SO8ROF3_0(.din(n32150), .dout(n32153));
    jdff dff_A_zlcWMyib6_0(.din(n32147), .dout(n32150));
    jdff dff_A_w8sKohNk5_0(.din(n32144), .dout(n32147));
    jdff dff_A_UI1R9Le08_0(.din(n32141), .dout(n32144));
    jdff dff_A_cMcUBohz8_0(.din(n32138), .dout(n32141));
    jdff dff_A_GnMpStnz1_0(.din(n32135), .dout(n32138));
    jdff dff_A_6wZbilJl2_0(.din(n32132), .dout(n32135));
    jdff dff_A_rp2XgVWh3_0(.din(n32129), .dout(n32132));
    jdff dff_A_6zutFgaU6_0(.din(n32126), .dout(n32129));
    jdff dff_A_JBUAY8Fw0_0(.din(n32123), .dout(n32126));
    jdff dff_A_l8jeQ4254_0(.din(n32120), .dout(n32123));
    jdff dff_A_Gr02eWPc5_0(.din(n32117), .dout(n32120));
    jdff dff_A_LmlYMnMJ8_0(.din(n32114), .dout(n32117));
    jdff dff_A_jBE172ew3_0(.din(n32111), .dout(n32114));
    jdff dff_A_OLAfH0io7_0(.din(n32108), .dout(n32111));
    jdff dff_A_1YDCgfkD9_0(.din(n32105), .dout(n32108));
    jdff dff_A_WpnxNDUE8_0(.din(n32102), .dout(n32105));
    jdff dff_A_Vw5fECnz2_0(.din(n32099), .dout(n32102));
    jdff dff_A_IGxYFOR93_0(.din(n32096), .dout(n32099));
    jdff dff_A_CoeC1kwg1_0(.din(n32093), .dout(n32096));
    jdff dff_A_mAfEbpZI0_0(.din(n32090), .dout(n32093));
    jdff dff_A_hdGFVPii0_0(.din(n32087), .dout(n32090));
    jdff dff_A_kyvCI4jS6_0(.din(n32084), .dout(n32087));
    jdff dff_A_R7C45UMu6_0(.din(n32081), .dout(n32084));
    jdff dff_A_Tyj5oO2W9_0(.din(n32078), .dout(n32081));
    jdff dff_A_gz1GsxHp5_0(.din(n32075), .dout(n32078));
    jdff dff_A_CqixKKVX0_0(.din(n32072), .dout(n32075));
    jdff dff_A_XvhIP3zA9_0(.din(n32069), .dout(n32072));
    jdff dff_A_seEZ09Bf8_0(.din(n32066), .dout(n32069));
    jdff dff_A_FMlrkncn3_0(.din(n32063), .dout(n32066));
    jdff dff_A_fIYMeOPI7_0(.din(n32060), .dout(n32063));
    jdff dff_A_nv6ZFavq7_0(.din(n32057), .dout(n32060));
    jdff dff_A_AARyv2OZ4_0(.din(n32054), .dout(n32057));
    jdff dff_A_AhkEpVkb3_0(.din(n32051), .dout(n32054));
    jdff dff_A_lySbVBV65_0(.din(n32048), .dout(n32051));
    jdff dff_A_NsfJuRvx0_0(.din(n32045), .dout(n32048));
    jdff dff_A_7hQEarXC6_0(.din(n32042), .dout(n32045));
    jdff dff_A_kW8m9Uc21_0(.din(n32039), .dout(n32042));
    jdff dff_A_rmuaJVc84_0(.din(n32036), .dout(n32039));
    jdff dff_A_Ie2YxNOe9_0(.din(n32033), .dout(n32036));
    jdff dff_A_57ZLz1p54_0(.din(n32030), .dout(n32033));
    jdff dff_A_g0eAg3Co1_0(.din(n32027), .dout(n32030));
    jdff dff_A_WijUF9467_0(.din(n32024), .dout(n32027));
    jdff dff_A_zbTTgX4P1_0(.din(n32021), .dout(n32024));
    jdff dff_A_kwZ2gT2t5_0(.din(n32018), .dout(n32021));
    jdff dff_A_IScTT8RI7_0(.din(n32015), .dout(n32018));
    jdff dff_A_smRvgRlM3_0(.din(n32012), .dout(n32015));
    jdff dff_A_95RTOtd64_0(.din(n32009), .dout(n32012));
    jdff dff_A_7Q7l75KR3_0(.din(n32006), .dout(n32009));
    jdff dff_A_NBJwJOM78_0(.din(n32003), .dout(n32006));
    jdff dff_A_X7s0jOUv1_0(.din(n32000), .dout(n32003));
    jdff dff_A_WOiBWxin6_0(.din(n31997), .dout(n32000));
    jdff dff_A_WaoXTjPl0_0(.din(n31994), .dout(n31997));
    jdff dff_A_JBM5vqQf6_0(.din(n31991), .dout(n31994));
    jdff dff_A_G7Yi1Tj75_0(.din(n31988), .dout(n31991));
    jdff dff_A_poLHy51T9_0(.din(n31985), .dout(n31988));
    jdff dff_A_TXQDmXQu9_0(.din(n31982), .dout(n31985));
    jdff dff_A_buo4FdL10_2(.din(n144), .dout(n31982));
    jdff dff_A_blGfFtq53_0(.din(n31976), .dout(G1581gat));
    jdff dff_A_lamaJPT51_0(.din(n31973), .dout(n31976));
    jdff dff_A_q6O0bSP29_0(.din(n31970), .dout(n31973));
    jdff dff_A_vRK7OhD86_0(.din(n31967), .dout(n31970));
    jdff dff_A_0Lq0JNAS8_0(.din(n31964), .dout(n31967));
    jdff dff_A_WLCOgiXJ7_0(.din(n31961), .dout(n31964));
    jdff dff_A_81v8lyms0_0(.din(n31958), .dout(n31961));
    jdff dff_A_vwszhUu81_0(.din(n31955), .dout(n31958));
    jdff dff_A_AL20DwRz2_0(.din(n31952), .dout(n31955));
    jdff dff_A_CPjkiGVQ2_0(.din(n31949), .dout(n31952));
    jdff dff_A_rOO9VspZ6_0(.din(n31946), .dout(n31949));
    jdff dff_A_VBddhrBH2_0(.din(n31943), .dout(n31946));
    jdff dff_A_rOD5n1Y23_0(.din(n31940), .dout(n31943));
    jdff dff_A_EEkZZj2h4_0(.din(n31937), .dout(n31940));
    jdff dff_A_T0mmnZeG6_0(.din(n31934), .dout(n31937));
    jdff dff_A_UXcMNORi3_0(.din(n31931), .dout(n31934));
    jdff dff_A_SShDmPL80_0(.din(n31928), .dout(n31931));
    jdff dff_A_zs9xhk1c1_0(.din(n31925), .dout(n31928));
    jdff dff_A_EsqYMR8O7_0(.din(n31922), .dout(n31925));
    jdff dff_A_epFCYmGl7_0(.din(n31919), .dout(n31922));
    jdff dff_A_2tnSaPAX0_0(.din(n31916), .dout(n31919));
    jdff dff_A_INDGoFkg3_0(.din(n31913), .dout(n31916));
    jdff dff_A_tBVi5mJQ8_0(.din(n31910), .dout(n31913));
    jdff dff_A_dbATNVWm6_0(.din(n31907), .dout(n31910));
    jdff dff_A_BdaQd5Rb9_0(.din(n31904), .dout(n31907));
    jdff dff_A_7gBGe5ps6_0(.din(n31901), .dout(n31904));
    jdff dff_A_lAIycoQE7_0(.din(n31898), .dout(n31901));
    jdff dff_A_RS0rcUYA9_0(.din(n31895), .dout(n31898));
    jdff dff_A_KUtIuPcF4_0(.din(n31892), .dout(n31895));
    jdff dff_A_K5RERxYj4_0(.din(n31889), .dout(n31892));
    jdff dff_A_Eb114fix2_0(.din(n31886), .dout(n31889));
    jdff dff_A_mniHZ3B98_0(.din(n31883), .dout(n31886));
    jdff dff_A_1EVHpBAP4_0(.din(n31880), .dout(n31883));
    jdff dff_A_D6UvXoZM2_0(.din(n31877), .dout(n31880));
    jdff dff_A_Fv68ae0f3_0(.din(n31874), .dout(n31877));
    jdff dff_A_sMZeNh7a9_0(.din(n31871), .dout(n31874));
    jdff dff_A_PhEvehmV8_0(.din(n31868), .dout(n31871));
    jdff dff_A_htP9gWyX3_0(.din(n31865), .dout(n31868));
    jdff dff_A_20HUvyKL2_0(.din(n31862), .dout(n31865));
    jdff dff_A_CkV3fprj9_0(.din(n31859), .dout(n31862));
    jdff dff_A_W1dEsIh73_0(.din(n31856), .dout(n31859));
    jdff dff_A_V3EB6ZcX4_0(.din(n31853), .dout(n31856));
    jdff dff_A_GtoYfMj76_0(.din(n31850), .dout(n31853));
    jdff dff_A_HJyifzUq5_0(.din(n31847), .dout(n31850));
    jdff dff_A_P4W3ewrv5_0(.din(n31844), .dout(n31847));
    jdff dff_A_0ExLSiUF7_0(.din(n31841), .dout(n31844));
    jdff dff_A_tuzudz8Y8_0(.din(n31838), .dout(n31841));
    jdff dff_A_AiXJQjp85_0(.din(n31835), .dout(n31838));
    jdff dff_A_F6cmjWKV8_0(.din(n31832), .dout(n31835));
    jdff dff_A_Evb8SzQx3_0(.din(n31829), .dout(n31832));
    jdff dff_A_csbgERdT2_0(.din(n31826), .dout(n31829));
    jdff dff_A_ke1r9i094_0(.din(n31823), .dout(n31826));
    jdff dff_A_ZwjQEB1m5_0(.din(n31820), .dout(n31823));
    jdff dff_A_7HqJiyOl4_0(.din(n31817), .dout(n31820));
    jdff dff_A_tew7kQNq2_0(.din(n31814), .dout(n31817));
    jdff dff_A_jSaQJkPg7_0(.din(n31811), .dout(n31814));
    jdff dff_A_unkegTzu8_0(.din(n31808), .dout(n31811));
    jdff dff_A_cszTkADn4_0(.din(n31805), .dout(n31808));
    jdff dff_A_NAQK3TVa0_0(.din(n31802), .dout(n31805));
    jdff dff_A_T1wKX3wU2_0(.din(n31799), .dout(n31802));
    jdff dff_A_NWvETIUF0_0(.din(n31796), .dout(n31799));
    jdff dff_A_2TrdDXiy6_0(.din(n31793), .dout(n31796));
    jdff dff_A_KQCOlCla5_0(.din(n31790), .dout(n31793));
    jdff dff_A_Sbe3YF118_0(.din(n31787), .dout(n31790));
    jdff dff_A_6hyZpext7_0(.din(n31784), .dout(n31787));
    jdff dff_A_rw9zDxdR1_0(.din(n31781), .dout(n31784));
    jdff dff_A_yFw1wAaJ8_0(.din(n31778), .dout(n31781));
    jdff dff_A_C73LlL5J4_0(.din(n31775), .dout(n31778));
    jdff dff_A_vRJlwoKH4_0(.din(n31772), .dout(n31775));
    jdff dff_A_TXpAQk9U3_2(.din(n103), .dout(n31772));
    jdff dff_A_tJS67BLc6_0(.din(n31766), .dout(G545gat));
    jdff dff_A_JVsAVccg2_0(.din(n31763), .dout(n31766));
    jdff dff_A_ohbgeCYa9_0(.din(n31760), .dout(n31763));
    jdff dff_A_ooBTxhM42_0(.din(n31757), .dout(n31760));
    jdff dff_A_5GQGx5pO5_0(.din(n31754), .dout(n31757));
    jdff dff_A_rDYz4CU07_0(.din(n31751), .dout(n31754));
    jdff dff_A_890P4iKA2_0(.din(n31748), .dout(n31751));
    jdff dff_A_PRlghX754_0(.din(n31745), .dout(n31748));
    jdff dff_A_WHkIXC9S7_0(.din(n31742), .dout(n31745));
    jdff dff_A_SXdZkzCK8_0(.din(n31739), .dout(n31742));
    jdff dff_A_h5p1L6Im0_0(.din(n31736), .dout(n31739));
    jdff dff_A_pw8NBRHb1_0(.din(n31733), .dout(n31736));
    jdff dff_A_y0Lfbng75_0(.din(n31730), .dout(n31733));
    jdff dff_A_oOvTVNbi6_0(.din(n31727), .dout(n31730));
    jdff dff_A_15MuG5kP2_0(.din(n31724), .dout(n31727));
    jdff dff_A_MKLHHGtO8_0(.din(n31721), .dout(n31724));
    jdff dff_A_xIqktCFN7_0(.din(n31718), .dout(n31721));
    jdff dff_A_AsbJXWKL8_0(.din(n31715), .dout(n31718));
    jdff dff_A_WxxUDhz89_0(.din(n31712), .dout(n31715));
    jdff dff_A_6ntCjEA50_0(.din(n31709), .dout(n31712));
    jdff dff_A_er8aXkTg5_0(.din(n31706), .dout(n31709));
    jdff dff_A_DxGRfkrQ7_0(.din(n31703), .dout(n31706));
    jdff dff_A_RBtRBIYw7_0(.din(n31700), .dout(n31703));
    jdff dff_A_IsojOi9V4_0(.din(n31697), .dout(n31700));
    jdff dff_A_0vxVuywM2_0(.din(n31694), .dout(n31697));
    jdff dff_A_PJj3rKIH7_0(.din(n31691), .dout(n31694));
    jdff dff_A_GkZLiVdJ6_0(.din(n31688), .dout(n31691));
    jdff dff_A_IhD23cpZ7_0(.din(n31685), .dout(n31688));
    jdff dff_A_lJavKu555_0(.din(n31682), .dout(n31685));
    jdff dff_A_80IDQ1SK6_0(.din(n31679), .dout(n31682));
    jdff dff_A_wn67Koel0_0(.din(n31676), .dout(n31679));
    jdff dff_A_JoN3L7Ym8_0(.din(n31673), .dout(n31676));
    jdff dff_A_u9QVAb9v2_0(.din(n31670), .dout(n31673));
    jdff dff_A_LD4LPZq52_0(.din(n31667), .dout(n31670));
    jdff dff_A_OW6khchs0_0(.din(n31664), .dout(n31667));
    jdff dff_A_MWZThVTg6_0(.din(n31661), .dout(n31664));
    jdff dff_A_p8qqB4hC7_0(.din(n31658), .dout(n31661));
    jdff dff_A_BvpnkpUv4_0(.din(n31655), .dout(n31658));
    jdff dff_A_3aywD2BY3_0(.din(n31652), .dout(n31655));
    jdff dff_A_Lq5pI89p4_0(.din(n31649), .dout(n31652));
    jdff dff_A_fzMSTGnW4_0(.din(n31646), .dout(n31649));
    jdff dff_A_0GuCBN7h6_0(.din(n31643), .dout(n31646));
    jdff dff_A_XFPGfoyo9_0(.din(n31640), .dout(n31643));
    jdff dff_A_vttlEuDG3_0(.din(n31637), .dout(n31640));
    jdff dff_A_dd4IHaLo4_0(.din(n31634), .dout(n31637));
    jdff dff_A_Fj4mPkYJ5_0(.din(n31631), .dout(n31634));
    jdff dff_A_OlotAoqD8_0(.din(n31628), .dout(n31631));
    jdff dff_A_xhkOA6d50_0(.din(n31625), .dout(n31628));
    jdff dff_A_6VIoMdNo0_0(.din(n31622), .dout(n31625));
    jdff dff_A_1otuXqZt4_0(.din(n31619), .dout(n31622));
    jdff dff_A_9Eor3Hjo5_0(.din(n31616), .dout(n31619));
    jdff dff_A_y7Vu8jfj0_0(.din(n31613), .dout(n31616));
    jdff dff_A_3n7Q4p9d4_0(.din(n31610), .dout(n31613));
    jdff dff_A_8rg70ohz8_0(.din(n31607), .dout(n31610));
    jdff dff_A_vQku3r5r0_0(.din(n31604), .dout(n31607));
    jdff dff_A_vb3okClZ5_0(.din(n31601), .dout(n31604));
    jdff dff_A_8G0ZVXKd4_0(.din(n31598), .dout(n31601));
    jdff dff_A_tltlAlJX5_0(.din(n31595), .dout(n31598));
    jdff dff_A_IcvCZ8672_0(.din(n31592), .dout(n31595));
    jdff dff_A_nhrO4Cok2_0(.din(n31589), .dout(n31592));
    jdff dff_A_kBEVpuim4_0(.din(n31586), .dout(n31589));
    jdff dff_A_vDxG6o7n8_0(.din(n31583), .dout(n31586));
    jdff dff_A_OiAZEN2v0_0(.din(n31580), .dout(n31583));
    jdff dff_A_QYQci1fk0_0(.din(n31577), .dout(n31580));
    jdff dff_A_zo0549vH2_0(.din(n31574), .dout(n31577));
    jdff dff_A_iPlPA2Ip5_0(.din(n31571), .dout(n31574));
    jdff dff_A_7Y8JO7ZJ2_0(.din(n31568), .dout(n31571));
    jdff dff_A_YeHL9aIy8_0(.din(n31565), .dout(n31568));
    jdff dff_A_LljHSyni0_0(.din(n31562), .dout(n31565));
    jdff dff_A_PdpyK4ry0_0(.din(n31559), .dout(n31562));
    jdff dff_A_eI17mUKL4_0(.din(n31556), .dout(n31559));
    jdff dff_A_pPQigq9M5_0(.din(n31553), .dout(n31556));
    jdff dff_A_4gQ9ZUKu3_0(.din(n31550), .dout(n31553));
    jdff dff_A_SBHDbXIx1_1(.din(n67), .dout(n31550));
    jdff dff_B_6xdhJ48v5_2(.din(n31545), .dout(n31548));
    jdff dff_B_iwILiT0Z8_2(.din(n31542), .dout(n31545));
    jdff dff_B_rJjPETkF3_2(.din(n3143), .dout(n31542));
    jdff dff_A_ZGZ8rWrU5_0(.din(n3147), .dout(n31538));
    jdff dff_A_cIGZ47B76_0(.din(n31538), .dout(n31535));
    jdff dff_B_4DEEQ4gN5_2(.din(n3155), .dout(n31533));
    jdff dff_A_kM3WLGk62_0(.din(n31533), .dout(n31529));
    jdff dff_A_MSQpi08P7_0(.din(n31529), .dout(n31526));
    jdff dff_A_UzGkmPuH7_0(.din(n31526), .dout(n31523));
    jdff dff_B_pWjCZ7xu6_2(.din(n3549), .dout(n31521));
    jdff dff_A_CQ0L2kB03_0(.din(n31521), .dout(n31517));
    jdff dff_A_4HSIEWTC5_0(.din(n31517), .dout(n31514));
    jdff dff_A_FudOx7h20_0(.din(n31514), .dout(n31511));
    jdff dff_B_lQTeKuBM6_2(.din(n31506), .dout(n31509));
    jdff dff_B_4QMQO2HH8_2(.din(n31503), .dout(n31506));
    jdff dff_B_zSwb67hh5_2(.din(n3560), .dout(n31503));
    jdff dff_B_uSkMMjTT2_2(.din(n31497), .dout(n31500));
    jdff dff_B_P1VSDqeu3_2(.din(n31494), .dout(n31497));
    jdff dff_B_pUoWxrfk5_2(.din(n31491), .dout(n31494));
    jdff dff_B_PuzwdCvi4_2(.din(n3564), .dout(n31491));
    jdff dff_B_rHluWfOf0_2(.din(n31485), .dout(n31488));
    jdff dff_B_WfJUC5Th7_2(.din(n31482), .dout(n31485));
    jdff dff_B_XFWsS37N1_2(.din(n31479), .dout(n31482));
    jdff dff_B_jomUdwLt9_2(.din(n31476), .dout(n31479));
    jdff dff_B_5JAcsR253_2(.din(n31473), .dout(n31476));
    jdff dff_B_VUMyWcSP6_2(.din(n31470), .dout(n31473));
    jdff dff_B_mkivJK7r1_2(.din(n31467), .dout(n31470));
    jdff dff_B_b7VkWaVq0_2(.din(n3528), .dout(n31467));
    jdff dff_B_Kvu2NZ8E1_1(.din(n3912), .dout(n31464));
    jdff dff_B_nWASdzTi0_2(.din(n31458), .dout(n31461));
    jdff dff_B_9AOZzDh31_2(.din(n31455), .dout(n31458));
    jdff dff_B_w1LqP5Ba0_2(.din(n31452), .dout(n31455));
    jdff dff_B_dj0bbnkz3_2(.din(n31449), .dout(n31452));
    jdff dff_B_Hs3Qj9xI6_2(.din(n31446), .dout(n31449));
    jdff dff_B_UIoTEzfY3_2(.din(n31443), .dout(n31446));
    jdff dff_B_NO34ytKQ1_2(.din(n3924), .dout(n31443));
    jdff dff_B_PJgaHfRU1_2(.din(n31437), .dout(n31440));
    jdff dff_B_k7SHEqls8_2(.din(n31434), .dout(n31437));
    jdff dff_B_VHvBBpfl8_2(.din(n31431), .dout(n31434));
    jdff dff_B_SmC5t9hb1_2(.din(n31428), .dout(n31431));
    jdff dff_B_xBcfH5Hk6_2(.din(n3928), .dout(n31428));
    jdff dff_B_gbsWdu792_2(.din(n31422), .dout(n31425));
    jdff dff_B_RbHQ6WDG5_2(.din(n31419), .dout(n31422));
    jdff dff_B_1KLaqIJr5_2(.din(n3947), .dout(n31419));
    jdff dff_B_dsSb6e5W5_2(.din(n31413), .dout(n31416));
    jdff dff_B_lBt4bscN8_2(.din(n31410), .dout(n31413));
    jdff dff_B_LoTTiBbr1_2(.din(n31407), .dout(n31410));
    jdff dff_B_gN1PgTyV2_2(.din(n31404), .dout(n31407));
    jdff dff_B_pdwwQ1TC8_2(.din(n31401), .dout(n31404));
    jdff dff_B_JOJvbckc7_2(.din(n31398), .dout(n31401));
    jdff dff_B_aCqy50DP1_2(.din(n31395), .dout(n31398));
    jdff dff_B_UF2C35uT0_2(.din(n31392), .dout(n31395));
    jdff dff_B_N2I7r5sW2_2(.din(n31389), .dout(n31392));
    jdff dff_B_7r0mPeHX4_2(.din(n31386), .dout(n31389));
    jdff dff_B_wsTcT6Du0_2(.din(n3908), .dout(n31386));
    jdff dff_B_5fzawKms6_1(.din(n4288), .dout(n31383));
    jdff dff_B_VjTNHORE0_2(.din(n31377), .dout(n31380));
    jdff dff_B_QVDCbL2V2_2(.din(n31374), .dout(n31377));
    jdff dff_B_qGvxvP9i8_2(.din(n31371), .dout(n31374));
    jdff dff_B_R6DVXZaE2_2(.din(n31368), .dout(n31371));
    jdff dff_B_ucHTXldm6_2(.din(n31365), .dout(n31368));
    jdff dff_B_yr5QtQdn2_2(.din(n31362), .dout(n31365));
    jdff dff_B_CIjp0FNg9_2(.din(n31359), .dout(n31362));
    jdff dff_B_APs3vc0s8_2(.din(n31356), .dout(n31359));
    jdff dff_B_7IvXLYJf4_2(.din(n31353), .dout(n31356));
    jdff dff_B_HvS5g1lJ0_2(.din(n31350), .dout(n31353));
    jdff dff_B_mPD3MaaR6_2(.din(n4300), .dout(n31350));
    jdff dff_B_0k8pGfeg4_2(.din(n31344), .dout(n31347));
    jdff dff_B_TbL9iLmj7_2(.din(n31341), .dout(n31344));
    jdff dff_B_2KlZSCcS2_2(.din(n31338), .dout(n31341));
    jdff dff_B_37Ba0chz7_2(.din(n31335), .dout(n31338));
    jdff dff_B_7bXp8v1W7_2(.din(n31332), .dout(n31335));
    jdff dff_B_OX3vOu7t7_2(.din(n31329), .dout(n31332));
    jdff dff_B_J7EFGDsQ1_2(.din(n31326), .dout(n31329));
    jdff dff_B_bpSmEV1q8_2(.din(n31323), .dout(n31326));
    jdff dff_B_QaLurC0e0_2(.din(n4304), .dout(n31323));
    jdff dff_B_SD9sF0Cs1_1(.din(n31317), .dout(n31320));
    jdff dff_B_OFzGlZfO7_1(.din(n4308), .dout(n31317));
    jdff dff_B_OJa5jAA83_2(.din(n31311), .dout(n31314));
    jdff dff_B_vLBFI7kX2_2(.din(n4327), .dout(n31311));
    jdff dff_B_DnRcI9J06_2(.din(n31305), .dout(n31308));
    jdff dff_B_u6FExlep8_2(.din(n31302), .dout(n31305));
    jdff dff_B_LU2xYyHE0_2(.din(n31299), .dout(n31302));
    jdff dff_B_PMHAVfwd9_2(.din(n31296), .dout(n31299));
    jdff dff_B_ruSHOu9E3_2(.din(n31293), .dout(n31296));
    jdff dff_B_vpbQY6bd2_2(.din(n31290), .dout(n31293));
    jdff dff_B_gK4EYb8k8_2(.din(n31287), .dout(n31290));
    jdff dff_B_oY9Nxm7D8_2(.din(n31284), .dout(n31287));
    jdff dff_B_mLmBGkIA4_2(.din(n31281), .dout(n31284));
    jdff dff_B_zejx364E6_2(.din(n31278), .dout(n31281));
    jdff dff_B_4vgmQj8H5_2(.din(n31275), .dout(n31278));
    jdff dff_B_iij9tUrU4_2(.din(n31272), .dout(n31275));
    jdff dff_B_0ZlW6rUd3_2(.din(n31269), .dout(n31272));
    jdff dff_B_gz4ugIcs0_2(.din(n4284), .dout(n31269));
    jdff dff_B_aeNosS844_1(.din(n4638), .dout(n31266));
    jdff dff_B_BP1LWsrF9_2(.din(n31260), .dout(n31263));
    jdff dff_B_Iu5vrsMQ1_2(.din(n31257), .dout(n31260));
    jdff dff_B_tYLlUs1z0_2(.din(n31254), .dout(n31257));
    jdff dff_B_WpxNynRH4_2(.din(n31251), .dout(n31254));
    jdff dff_B_GHJChAcJ6_2(.din(n31248), .dout(n31251));
    jdff dff_B_rpMtXSaV3_2(.din(n31245), .dout(n31248));
    jdff dff_B_Zaa1qRCy2_2(.din(n31242), .dout(n31245));
    jdff dff_B_BNAFJrX09_2(.din(n31239), .dout(n31242));
    jdff dff_B_GJtcJ5q20_2(.din(n31236), .dout(n31239));
    jdff dff_B_JlVxxxPi2_2(.din(n31233), .dout(n31236));
    jdff dff_B_q5f0g6KW4_2(.din(n31230), .dout(n31233));
    jdff dff_B_pgm5CIOg2_2(.din(n31227), .dout(n31230));
    jdff dff_B_XquK6lfj3_2(.din(n31224), .dout(n31227));
    jdff dff_B_BxPtfmVg5_2(.din(n31221), .dout(n31224));
    jdff dff_B_tkPmTYjn8_2(.din(n4650), .dout(n31221));
    jdff dff_B_HYsBGq0B0_2(.din(n31215), .dout(n31218));
    jdff dff_B_kHxt7nel9_2(.din(n31212), .dout(n31215));
    jdff dff_B_jOZ1XtX40_2(.din(n31209), .dout(n31212));
    jdff dff_B_siqKQiPV5_2(.din(n31206), .dout(n31209));
    jdff dff_B_ZRGZ9G752_2(.din(n31203), .dout(n31206));
    jdff dff_B_vAaQu0rq1_2(.din(n31200), .dout(n31203));
    jdff dff_B_nbQo6sYz5_2(.din(n31197), .dout(n31200));
    jdff dff_B_24l28blo8_2(.din(n31194), .dout(n31197));
    jdff dff_B_eLLo6tPw3_2(.din(n31191), .dout(n31194));
    jdff dff_B_EZgn3QZ04_2(.din(n31188), .dout(n31191));
    jdff dff_B_BtC00bdT3_2(.din(n31185), .dout(n31188));
    jdff dff_B_IUVelolb2_2(.din(n31182), .dout(n31185));
    jdff dff_B_S7miAAlE2_2(.din(n4654), .dout(n31182));
    jdff dff_B_DIHpMLGD7_1(.din(n31176), .dout(n31179));
    jdff dff_B_w3UW7JaH0_1(.din(n4658), .dout(n31176));
    jdff dff_B_PgfjzkDW5_2(.din(n4677), .dout(n31173));
    jdff dff_B_YDaxvvi08_2(.din(n31167), .dout(n31170));
    jdff dff_B_CQzbtU104_0(.din(n95), .dout(n10593));
    jdff dff_B_lEuxbv5F0_0(.din(n10593), .dout(n10596));
    jdff dff_B_m2YFsOFD9_1(.din(n110), .dout(n10599));
    jdff dff_B_b2YnYtSV1_1(.din(n10599), .dout(n10602));
    jdff dff_B_5LuDeCfj3_1(.din(n10602), .dout(n10605));
    jdff dff_B_WFVxcR7l8_1(.din(n151), .dout(n10608));
    jdff dff_B_A4lZUm4M2_1(.din(n10608), .dout(n10611));
    jdff dff_B_6FQXuesw2_1(.din(n10611), .dout(n10614));
    jdff dff_B_0gcEPcrz3_1(.din(n10614), .dout(n10617));
    jdff dff_B_KvMrhP0T4_1(.din(n10617), .dout(n10620));
    jdff dff_B_HfeP3lcw0_1(.din(n10620), .dout(n10623));
    jdff dff_B_i8xu0OGh6_1(.din(n227), .dout(n10626));
    jdff dff_B_OQQcgr6h1_1(.din(n10626), .dout(n10629));
    jdff dff_B_q9eLr02q1_1(.din(n10629), .dout(n10632));
    jdff dff_B_I3Ru0P1g5_1(.din(n10632), .dout(n10635));
    jdff dff_B_7YBUKEnd7_1(.din(n10635), .dout(n10638));
    jdff dff_B_Zkre0t9S8_1(.din(n10638), .dout(n10641));
    jdff dff_B_QCM5rOcm5_1(.din(n10641), .dout(n10644));
    jdff dff_B_vmjV8cet6_1(.din(n10644), .dout(n10647));
    jdff dff_B_k71p4s1n3_1(.din(n10647), .dout(n10650));
    jdff dff_B_HH8HPvVI0_1(.din(n336), .dout(n10653));
    jdff dff_B_QqQK8s0U3_1(.din(n10653), .dout(n10656));
    jdff dff_B_kCeu8XBG1_1(.din(n10656), .dout(n10659));
    jdff dff_B_dxQzISG90_1(.din(n10659), .dout(n10662));
    jdff dff_B_FGCQnwCp5_1(.din(n10662), .dout(n10665));
    jdff dff_B_1CSPJc2a0_1(.din(n10665), .dout(n10668));
    jdff dff_B_uPvNFZ5c1_1(.din(n10668), .dout(n10671));
    jdff dff_B_BNbxdmAq4_1(.din(n10671), .dout(n10674));
    jdff dff_B_tBwCKQwe8_1(.din(n10674), .dout(n10677));
    jdff dff_B_DPQZ5tvD5_1(.din(n10677), .dout(n10680));
    jdff dff_B_fqpEbCij6_1(.din(n10680), .dout(n10683));
    jdff dff_B_PcDM2u6M1_1(.din(n10683), .dout(n10686));
    jdff dff_B_yAJYlebs5_1(.din(n468), .dout(n10689));
    jdff dff_B_L9zoaLbS3_1(.din(n10689), .dout(n10692));
    jdff dff_B_ZF4KR1sm0_1(.din(n10692), .dout(n10695));
    jdff dff_B_IUAIBhO16_1(.din(n10695), .dout(n10698));
    jdff dff_B_zZlEm5fz8_1(.din(n10698), .dout(n10701));
    jdff dff_B_vjaNgyfC6_1(.din(n10701), .dout(n10704));
    jdff dff_B_U7jcckH96_1(.din(n10704), .dout(n10707));
    jdff dff_B_kWtxciCH1_1(.din(n10707), .dout(n10710));
    jdff dff_B_cL18KVjY0_1(.din(n10710), .dout(n10713));
    jdff dff_B_5OBCqHq93_1(.din(n10713), .dout(n10716));
    jdff dff_B_SFJx1Xso7_1(.din(n10716), .dout(n10719));
    jdff dff_B_Kja5SFmP6_1(.din(n10719), .dout(n10722));
    jdff dff_B_tYDsVwD79_1(.din(n10722), .dout(n10725));
    jdff dff_B_r7koO1Cd2_1(.din(n10725), .dout(n10728));
    jdff dff_B_5lzuWr6g6_1(.din(n10728), .dout(n10731));
    jdff dff_B_rvQUMrX54_1(.din(n627), .dout(n10734));
    jdff dff_B_lXCG7Vdi4_1(.din(n10734), .dout(n10737));
    jdff dff_B_QcjPscN71_1(.din(n10737), .dout(n10740));
    jdff dff_B_8Z8mEQet0_1(.din(n10740), .dout(n10743));
    jdff dff_B_vqGt22TA8_1(.din(n10743), .dout(n10746));
    jdff dff_B_buYVPwG02_1(.din(n10746), .dout(n10749));
    jdff dff_B_axfIYrza8_1(.din(n10749), .dout(n10752));
    jdff dff_B_GcG9iY9w2_1(.din(n10752), .dout(n10755));
    jdff dff_B_bOkHvbh19_1(.din(n10755), .dout(n10758));
    jdff dff_B_DVNXvqNt3_1(.din(n10758), .dout(n10761));
    jdff dff_B_HqbXxAvh1_1(.din(n10761), .dout(n10764));
    jdff dff_B_OAhj6Tw48_1(.din(n10764), .dout(n10767));
    jdff dff_B_aRs7Cx5P3_1(.din(n10767), .dout(n10770));
    jdff dff_B_wZ0tyaKd6_1(.din(n10770), .dout(n10773));
    jdff dff_B_ZY3QDktq1_1(.din(n10773), .dout(n10776));
    jdff dff_B_9qnEvK782_1(.din(n10776), .dout(n10779));
    jdff dff_B_gPfvKI8H1_1(.din(n10779), .dout(n10782));
    jdff dff_B_so7U7eC87_1(.din(n10782), .dout(n10785));
    jdff dff_B_BUyvwPbb1_1(.din(n813), .dout(n10788));
    jdff dff_B_elVOzZ7q4_1(.din(n10788), .dout(n10791));
    jdff dff_B_Vh7Y9NNi4_1(.din(n10791), .dout(n10794));
    jdff dff_B_JULEhToh9_1(.din(n10794), .dout(n10797));
    jdff dff_B_ZH3oGxlj7_1(.din(n10797), .dout(n10800));
    jdff dff_B_xsy6icMC9_1(.din(n10800), .dout(n10803));
    jdff dff_B_WTuFu6Cv4_1(.din(n10803), .dout(n10806));
    jdff dff_B_cRFxGYkK1_1(.din(n10806), .dout(n10809));
    jdff dff_B_AgMqf6K30_1(.din(n10809), .dout(n10812));
    jdff dff_B_XYW3L56N0_1(.din(n10812), .dout(n10815));
    jdff dff_B_lQf1FyrY4_1(.din(n10815), .dout(n10818));
    jdff dff_B_CLGPZbuj3_1(.din(n10818), .dout(n10821));
    jdff dff_B_4CV3vP6I7_1(.din(n10821), .dout(n10824));
    jdff dff_B_RUUqzdH85_1(.din(n10824), .dout(n10827));
    jdff dff_B_A4zxo8ba5_1(.din(n10827), .dout(n10830));
    jdff dff_B_PkSuJ1jH0_1(.din(n10830), .dout(n10833));
    jdff dff_B_IwnpOftq1_1(.din(n10833), .dout(n10836));
    jdff dff_B_rgS15Ok66_1(.din(n10836), .dout(n10839));
    jdff dff_B_EpuBHSCh7_1(.din(n10839), .dout(n10842));
    jdff dff_B_0esQzCRK8_1(.din(n10842), .dout(n10845));
    jdff dff_B_m3PEL1Gm3_1(.din(n10845), .dout(n10848));
    jdff dff_B_om5yi6oo6_1(.din(n1026), .dout(n10851));
    jdff dff_B_RNaMrRvH6_1(.din(n10851), .dout(n10854));
    jdff dff_B_SENSpIqz4_1(.din(n10854), .dout(n10857));
    jdff dff_B_P9Uq7ySz0_1(.din(n10857), .dout(n10860));
    jdff dff_B_gGLWvwHE0_1(.din(n10860), .dout(n10863));
    jdff dff_B_5xawmo587_1(.din(n10863), .dout(n10866));
    jdff dff_B_HF85Sorq0_1(.din(n10866), .dout(n10869));
    jdff dff_B_McV18ixf3_1(.din(n10869), .dout(n10872));
    jdff dff_B_tspBcsNe5_1(.din(n10872), .dout(n10875));
    jdff dff_B_8KvmIXAE4_1(.din(n10875), .dout(n10878));
    jdff dff_B_1PlvDrQ21_1(.din(n10878), .dout(n10881));
    jdff dff_B_RRqtvSfw5_1(.din(n10881), .dout(n10884));
    jdff dff_B_nSHEtc8K3_1(.din(n10884), .dout(n10887));
    jdff dff_B_p4kuG29k6_1(.din(n10887), .dout(n10890));
    jdff dff_B_dd5qWz7c1_1(.din(n10890), .dout(n10893));
    jdff dff_B_G8juxv5v1_1(.din(n10893), .dout(n10896));
    jdff dff_B_s2YN9vxX1_1(.din(n10896), .dout(n10899));
    jdff dff_B_5YcMWnSx7_1(.din(n10899), .dout(n10902));
    jdff dff_B_GfcNu1Pm8_1(.din(n10902), .dout(n10905));
    jdff dff_B_Q0U8vNiJ5_1(.din(n10905), .dout(n10908));
    jdff dff_B_RTNinQqY8_1(.din(n10908), .dout(n10911));
    jdff dff_B_xgb81Vz88_1(.din(n10911), .dout(n10914));
    jdff dff_B_RoA3tBvL4_1(.din(n10914), .dout(n10917));
    jdff dff_B_vGQOMZBB4_1(.din(n10917), .dout(n10920));
    jdff dff_B_1thrLE4J6_1(.din(n1266), .dout(n10923));
    jdff dff_B_d6xtxwtY7_1(.din(n10923), .dout(n10926));
    jdff dff_B_pBJyrQGT0_1(.din(n10926), .dout(n10929));
    jdff dff_B_zfMrTPdX8_1(.din(n10929), .dout(n10932));
    jdff dff_B_rqsZCN590_1(.din(n10932), .dout(n10935));
    jdff dff_B_RgPVaUv77_1(.din(n10935), .dout(n10938));
    jdff dff_B_2YqoXrLH1_1(.din(n10938), .dout(n10941));
    jdff dff_B_oRoaPbra3_1(.din(n10941), .dout(n10944));
    jdff dff_B_xaVLPsu49_1(.din(n10944), .dout(n10947));
    jdff dff_B_wQlgNhLa9_1(.din(n10947), .dout(n10950));
    jdff dff_B_WrfQEx1C9_1(.din(n10950), .dout(n10953));
    jdff dff_B_Sd5vFueX7_1(.din(n10953), .dout(n10956));
    jdff dff_B_SN7GOMXW4_1(.din(n10956), .dout(n10959));
    jdff dff_B_fK4bgWEk7_1(.din(n10959), .dout(n10962));
    jdff dff_B_fW7d0Ilt6_1(.din(n10962), .dout(n10965));
    jdff dff_B_Uq6KDSWv2_1(.din(n10965), .dout(n10968));
    jdff dff_B_JW9BKxOH9_1(.din(n10968), .dout(n10971));
    jdff dff_B_JV781Cy01_1(.din(n10971), .dout(n10974));
    jdff dff_B_bY10uaJ73_1(.din(n10974), .dout(n10977));
    jdff dff_B_sgIQiEtB3_1(.din(n10977), .dout(n10980));
    jdff dff_B_C2SNLFqJ7_1(.din(n10980), .dout(n10983));
    jdff dff_B_ahZNrPcM3_1(.din(n10983), .dout(n10986));
    jdff dff_B_PRVmNAZi2_1(.din(n10986), .dout(n10989));
    jdff dff_B_JoZcubzt1_1(.din(n10989), .dout(n10992));
    jdff dff_B_n3g5oXJa5_1(.din(n10992), .dout(n10995));
    jdff dff_B_BznF3FIb6_1(.din(n10995), .dout(n10998));
    jdff dff_B_0X766xLg1_1(.din(n10998), .dout(n11001));
    jdff dff_B_Ohaxnjpv1_1(.din(n1536), .dout(n11004));
    jdff dff_B_Wv2zYr603_1(.din(n11004), .dout(n11007));
    jdff dff_B_qCibCRSU7_1(.din(n11007), .dout(n11010));
    jdff dff_B_esUgqMcf7_1(.din(n11010), .dout(n11013));
    jdff dff_B_g5YFE9H99_1(.din(n11013), .dout(n11016));
    jdff dff_B_QQv9vc7A3_1(.din(n11016), .dout(n11019));
    jdff dff_B_QcL6UJab8_1(.din(n11019), .dout(n11022));
    jdff dff_B_TSTDwVwp3_1(.din(n11022), .dout(n11025));
    jdff dff_B_Uf0UaQSc9_1(.din(n11025), .dout(n11028));
    jdff dff_B_xKDbCvj80_1(.din(n11028), .dout(n11031));
    jdff dff_B_a9NgOcio2_1(.din(n11031), .dout(n11034));
    jdff dff_B_HcrrAszy4_1(.din(n11034), .dout(n11037));
    jdff dff_B_BX3Q1osR8_1(.din(n11037), .dout(n11040));
    jdff dff_B_b7YPd1iR0_1(.din(n11040), .dout(n11043));
    jdff dff_B_mKgddXPJ7_1(.din(n11043), .dout(n11046));
    jdff dff_B_Ul9xBQiK3_1(.din(n11046), .dout(n11049));
    jdff dff_B_TpvobFwx6_1(.din(n11049), .dout(n11052));
    jdff dff_B_lpnll1dX3_1(.din(n11052), .dout(n11055));
    jdff dff_B_RYRal4Ol3_1(.din(n11055), .dout(n11058));
    jdff dff_B_hHpZTndD7_1(.din(n11058), .dout(n11061));
    jdff dff_B_3B7n4IN74_1(.din(n11061), .dout(n11064));
    jdff dff_B_x8QwSilg4_1(.din(n11064), .dout(n11067));
    jdff dff_B_apnd5IDr9_1(.din(n11067), .dout(n11070));
    jdff dff_B_IHiiTo3O6_1(.din(n11070), .dout(n11073));
    jdff dff_B_sIpOpXkx0_1(.din(n11073), .dout(n11076));
    jdff dff_B_s83mAJLg8_1(.din(n11076), .dout(n11079));
    jdff dff_B_yeVQDdmo1_1(.din(n11079), .dout(n11082));
    jdff dff_B_zfGdRU5l7_1(.din(n11082), .dout(n11085));
    jdff dff_B_67DesMrR9_1(.din(n11085), .dout(n11088));
    jdff dff_B_1Aoe1Zp02_1(.din(n11088), .dout(n11091));
    jdff dff_B_KJ8ERTgx0_1(.din(n1833), .dout(n11094));
    jdff dff_B_t6pgtpSN5_1(.din(n11094), .dout(n11097));
    jdff dff_B_0wvmjINJ5_1(.din(n11097), .dout(n11100));
    jdff dff_B_c1bT9x5k3_1(.din(n11100), .dout(n11103));
    jdff dff_B_4LN2QOOh6_1(.din(n11103), .dout(n11106));
    jdff dff_B_OfhxVnc54_1(.din(n11106), .dout(n11109));
    jdff dff_B_tiIEoovw4_1(.din(n11109), .dout(n11112));
    jdff dff_B_b53M9FKu8_1(.din(n11112), .dout(n11115));
    jdff dff_B_XxgO3fsy4_1(.din(n11115), .dout(n11118));
    jdff dff_B_Xlc5vSBR1_1(.din(n11118), .dout(n11121));
    jdff dff_B_aoAsfADC9_1(.din(n11121), .dout(n11124));
    jdff dff_B_2Mb77foR9_1(.din(n11124), .dout(n11127));
    jdff dff_B_5WwukQxC4_1(.din(n11127), .dout(n11130));
    jdff dff_B_RQ5xwhgu3_1(.din(n11130), .dout(n11133));
    jdff dff_B_bYMdPLlh5_1(.din(n11133), .dout(n11136));
    jdff dff_B_iwxCcSjO6_1(.din(n11136), .dout(n11139));
    jdff dff_B_fQfxNQOK0_1(.din(n11139), .dout(n11142));
    jdff dff_B_s8kfIGKo6_1(.din(n11142), .dout(n11145));
    jdff dff_B_tyYRCZIO8_1(.din(n11145), .dout(n11148));
    jdff dff_B_OEb6m1KX0_1(.din(n11148), .dout(n11151));
    jdff dff_B_Vo9cFIp64_1(.din(n11151), .dout(n11154));
    jdff dff_B_8y9R6sCY2_1(.din(n11154), .dout(n11157));
    jdff dff_B_tmAYfzY61_1(.din(n11157), .dout(n11160));
    jdff dff_B_LL1POgVB0_1(.din(n11160), .dout(n11163));
    jdff dff_B_1ywzHM0E6_1(.din(n11163), .dout(n11166));
    jdff dff_B_G2YRkX784_1(.din(n11166), .dout(n11169));
    jdff dff_B_euuIZCO06_1(.din(n11169), .dout(n11172));
    jdff dff_B_AOLl8XXU4_1(.din(n11172), .dout(n11175));
    jdff dff_B_3tJ6Ru2z1_1(.din(n11175), .dout(n11178));
    jdff dff_B_1xWW39aW4_1(.din(n11178), .dout(n11181));
    jdff dff_B_igPDpLnN4_1(.din(n11181), .dout(n11184));
    jdff dff_B_BQUck8pw6_1(.din(n11184), .dout(n11187));
    jdff dff_B_EMXdE2Dp7_1(.din(n11187), .dout(n11190));
    jdff dff_B_o5KyN9Av8_1(.din(n2157), .dout(n11193));
    jdff dff_B_iRKRjkPD3_1(.din(n11193), .dout(n11196));
    jdff dff_B_bNiXRNEt7_1(.din(n11196), .dout(n11199));
    jdff dff_B_VEZuYu6E5_1(.din(n11199), .dout(n11202));
    jdff dff_B_b0yhfW5y1_1(.din(n11202), .dout(n11205));
    jdff dff_B_XmdeWYy09_1(.din(n11205), .dout(n11208));
    jdff dff_B_RvcMJutV0_1(.din(n11208), .dout(n11211));
    jdff dff_B_q54efvMt6_1(.din(n11211), .dout(n11214));
    jdff dff_B_LZfvazFs7_1(.din(n11214), .dout(n11217));
    jdff dff_B_zkdoqCH55_1(.din(n11217), .dout(n11220));
    jdff dff_B_ldcZC9kl6_1(.din(n11220), .dout(n11223));
    jdff dff_B_zyZGnLg48_1(.din(n11223), .dout(n11226));
    jdff dff_B_6PCwuYHb9_1(.din(n11226), .dout(n11229));
    jdff dff_B_KO4JF4GX2_1(.din(n11229), .dout(n11232));
    jdff dff_B_xlK0L1Ug7_1(.din(n11232), .dout(n11235));
    jdff dff_B_wJjdlrfB6_1(.din(n11235), .dout(n11238));
    jdff dff_B_3Ji2gMQm7_1(.din(n11238), .dout(n11241));
    jdff dff_B_PfB9bUjh7_1(.din(n11241), .dout(n11244));
    jdff dff_B_dC8IHqIJ1_1(.din(n11244), .dout(n11247));
    jdff dff_B_HBS5AwK51_1(.din(n11247), .dout(n11250));
    jdff dff_B_EouPxaki8_1(.din(n11250), .dout(n11253));
    jdff dff_B_RrulAtdA1_1(.din(n11253), .dout(n11256));
    jdff dff_B_pF2aKIxn5_1(.din(n11256), .dout(n11259));
    jdff dff_B_MU30OuBi8_1(.din(n11259), .dout(n11262));
    jdff dff_B_2OfEKHBX4_1(.din(n11262), .dout(n11265));
    jdff dff_B_LS0Nnnbe9_1(.din(n11265), .dout(n11268));
    jdff dff_B_UI1ALbJ59_1(.din(n11268), .dout(n11271));
    jdff dff_B_i2YItJvF0_1(.din(n11271), .dout(n11274));
    jdff dff_B_u8OfvAuj2_1(.din(n11274), .dout(n11277));
    jdff dff_B_46lwCQV27_1(.din(n11277), .dout(n11280));
    jdff dff_B_ieZy9wnn7_1(.din(n11280), .dout(n11283));
    jdff dff_B_UM2IZ2TQ9_1(.din(n11283), .dout(n11286));
    jdff dff_B_G7fpRx6n5_1(.din(n11286), .dout(n11289));
    jdff dff_B_lWOX5vnu7_1(.din(n11289), .dout(n11292));
    jdff dff_B_w8mdgQxL8_1(.din(n11292), .dout(n11295));
    jdff dff_B_g0rjQRyU7_1(.din(n11295), .dout(n11298));
    jdff dff_B_mSkAwcO57_1(.din(n2508), .dout(n11301));
    jdff dff_B_8aKZDA7T4_1(.din(n11301), .dout(n11304));
    jdff dff_B_qiYe6hHG4_1(.din(n11304), .dout(n11307));
    jdff dff_B_p2oC7vdN4_1(.din(n11307), .dout(n11310));
    jdff dff_B_JbZNPpgs7_1(.din(n11310), .dout(n11313));
    jdff dff_B_HaaH6aMG8_1(.din(n11313), .dout(n11316));
    jdff dff_B_J7folQdM4_1(.din(n11316), .dout(n11319));
    jdff dff_B_yizmqqar9_1(.din(n11319), .dout(n11322));
    jdff dff_B_35aKkuzV0_1(.din(n11322), .dout(n11325));
    jdff dff_B_EHn5wVSy5_1(.din(n11325), .dout(n11328));
    jdff dff_B_JFgDmkrW3_1(.din(n11328), .dout(n11331));
    jdff dff_B_uXi9tDhs3_1(.din(n11331), .dout(n11334));
    jdff dff_B_vdqwhCzo3_1(.din(n11334), .dout(n11337));
    jdff dff_B_FqzXHXep2_1(.din(n11337), .dout(n11340));
    jdff dff_B_5UKeuiYK9_1(.din(n11340), .dout(n11343));
    jdff dff_B_qvxQFtuE9_1(.din(n11343), .dout(n11346));
    jdff dff_B_bXpVsNP53_1(.din(n11346), .dout(n11349));
    jdff dff_B_0fmmWaq16_1(.din(n11349), .dout(n11352));
    jdff dff_B_OeStJnji3_1(.din(n11352), .dout(n11355));
    jdff dff_B_LDuQEcWd1_1(.din(n11355), .dout(n11358));
    jdff dff_B_xifPqPjM2_1(.din(n11358), .dout(n11361));
    jdff dff_B_tXSItKuV4_1(.din(n11361), .dout(n11364));
    jdff dff_B_i0Qc3n010_1(.din(n11364), .dout(n11367));
    jdff dff_B_4Qc3BT602_1(.din(n11367), .dout(n11370));
    jdff dff_B_oKhZ9Px72_1(.din(n11370), .dout(n11373));
    jdff dff_B_r7Cgy82A9_1(.din(n11373), .dout(n11376));
    jdff dff_B_azoRYASO7_1(.din(n11376), .dout(n11379));
    jdff dff_B_5LPQTviR3_1(.din(n11379), .dout(n11382));
    jdff dff_B_oalh4PKc8_1(.din(n11382), .dout(n11385));
    jdff dff_B_VSJ31bKI6_1(.din(n11385), .dout(n11388));
    jdff dff_B_ERF1bee34_1(.din(n11388), .dout(n11391));
    jdff dff_B_GjShUze15_1(.din(n11391), .dout(n11394));
    jdff dff_B_xBN9sYd73_1(.din(n11394), .dout(n11397));
    jdff dff_B_TrtEvN463_1(.din(n11397), .dout(n11400));
    jdff dff_B_Dto28vYA0_1(.din(n11400), .dout(n11403));
    jdff dff_B_Wd6tI4do1_1(.din(n11403), .dout(n11406));
    jdff dff_B_nrI87EEZ2_1(.din(n11406), .dout(n11409));
    jdff dff_B_WuR5d0mp4_1(.din(n11409), .dout(n11412));
    jdff dff_B_R5ONn5iw7_1(.din(n11412), .dout(n11415));
    jdff dff_B_PP0smkJr0_1(.din(n2886), .dout(n11418));
    jdff dff_B_Z6uSNpOy7_1(.din(n11418), .dout(n11421));
    jdff dff_B_FkH7Nsub6_1(.din(n11421), .dout(n11424));
    jdff dff_B_bMddaBju1_1(.din(n11424), .dout(n11427));
    jdff dff_B_aNQnMqfL8_1(.din(n11427), .dout(n11430));
    jdff dff_B_cfoY5vZH4_1(.din(n11430), .dout(n11433));
    jdff dff_B_D1TEAkdy4_1(.din(n11433), .dout(n11436));
    jdff dff_B_nYixf4ck7_1(.din(n11436), .dout(n11439));
    jdff dff_B_E7GihjsA6_1(.din(n11439), .dout(n11442));
    jdff dff_B_OsmL041d6_1(.din(n11442), .dout(n11445));
    jdff dff_B_H0AYqXlV5_1(.din(n11445), .dout(n11448));
    jdff dff_B_AqCS8Wmr0_1(.din(n11448), .dout(n11451));
    jdff dff_B_5E5N8fbG7_1(.din(n11451), .dout(n11454));
    jdff dff_B_mbyGOUyK7_1(.din(n11454), .dout(n11457));
    jdff dff_B_NE2Esbso4_1(.din(n11457), .dout(n11460));
    jdff dff_B_hKZQVC1B9_1(.din(n11460), .dout(n11463));
    jdff dff_B_OaZI88vZ2_1(.din(n11463), .dout(n11466));
    jdff dff_B_QS0AaBq25_1(.din(n11466), .dout(n11469));
    jdff dff_B_nR662HS23_1(.din(n11469), .dout(n11472));
    jdff dff_B_fCejSuMv7_1(.din(n11472), .dout(n11475));
    jdff dff_B_fAWzTRaQ1_1(.din(n11475), .dout(n11478));
    jdff dff_B_yOrbzuPC5_1(.din(n11478), .dout(n11481));
    jdff dff_B_pzsHEBWb6_1(.din(n11481), .dout(n11484));
    jdff dff_B_Zn469Bwc7_1(.din(n11484), .dout(n11487));
    jdff dff_B_VLtRZy4v3_1(.din(n11487), .dout(n11490));
    jdff dff_B_ptQ25fex8_1(.din(n11490), .dout(n11493));
    jdff dff_B_jVX8F6Xl3_1(.din(n11493), .dout(n11496));
    jdff dff_B_CawEFLW32_1(.din(n11496), .dout(n11499));
    jdff dff_B_6Uk0kY1J5_1(.din(n11499), .dout(n11502));
    jdff dff_B_bbrhRmbf2_1(.din(n11502), .dout(n11505));
    jdff dff_B_Z3OEavTf6_1(.din(n11505), .dout(n11508));
    jdff dff_B_igpowbij3_1(.din(n11508), .dout(n11511));
    jdff dff_B_olWfDcaN6_1(.din(n11511), .dout(n11514));
    jdff dff_B_YXhLdMks0_1(.din(n11514), .dout(n11517));
    jdff dff_B_NQAj0qbZ9_1(.din(n11517), .dout(n11520));
    jdff dff_B_ngqDtuqD7_1(.din(n11520), .dout(n11523));
    jdff dff_B_kNPbp8J69_1(.din(n11523), .dout(n11526));
    jdff dff_B_8VV8Qc1M7_1(.din(n11526), .dout(n11529));
    jdff dff_B_ttafBy0w3_1(.din(n11529), .dout(n11532));
    jdff dff_B_bHVB0p1Z3_1(.din(n11532), .dout(n11535));
    jdff dff_B_AiGyld9I4_1(.din(n11535), .dout(n11538));
    jdff dff_B_6y3Mt8UG5_1(.din(n11538), .dout(n11541));
    jdff dff_B_z8w0zcKB8_0(.din(n4767), .dout(n11544));
    jdff dff_B_hV2wI3hE3_1(.din(n6738), .dout(n11547));
    jdff dff_B_tPuf6rMo7_1(.din(n11547), .dout(n11550));
    jdff dff_B_NK12tZbp3_1(.din(n11550), .dout(n11553));
    jdff dff_B_SKk71p9z7_1(.din(n11553), .dout(n11556));
    jdff dff_B_GiwqYT4t5_1(.din(n11556), .dout(n11559));
    jdff dff_B_gzxu1Q299_1(.din(n11559), .dout(n11562));
    jdff dff_B_7eVcSRTQ8_1(.din(n11562), .dout(n11565));
    jdff dff_B_DQvoTz455_1(.din(n11565), .dout(n11568));
    jdff dff_B_6cc3BkZ72_1(.din(n11568), .dout(n11571));
    jdff dff_B_IkXUt7xC5_1(.din(n11571), .dout(n11574));
    jdff dff_B_B10s512I5_1(.din(n11574), .dout(n11577));
    jdff dff_B_US89lrvl8_1(.din(n11577), .dout(n11580));
    jdff dff_B_hSmZqu2u0_1(.din(n11580), .dout(n11583));
    jdff dff_B_bJ7asy1c2_1(.din(n11583), .dout(n11586));
    jdff dff_B_huyM6Sbm7_1(.din(n11586), .dout(n11589));
    jdff dff_B_Zzjqdy094_0(.din(n6766), .dout(n11592));
    jdff dff_B_Lx8y4Qgd1_0(.din(n11592), .dout(n11595));
    jdff dff_B_n1DYH6Eu0_0(.din(n11595), .dout(n11598));
    jdff dff_B_BbkwgzEX7_0(.din(n11598), .dout(n11601));
    jdff dff_B_AnWxIQvn7_0(.din(n11601), .dout(n11604));
    jdff dff_B_Cu2zUTVv4_0(.din(n11604), .dout(n11607));
    jdff dff_B_fCzsxwc23_0(.din(n11607), .dout(n11610));
    jdff dff_B_hC0stYPe2_0(.din(n11610), .dout(n11613));
    jdff dff_B_xDjbwjZR5_0(.din(n11613), .dout(n11616));
    jdff dff_B_22CDTs6g3_0(.din(n11616), .dout(n11619));
    jdff dff_B_y0h7Pa8r2_0(.din(n11619), .dout(n11622));
    jdff dff_B_nUH4L31U6_0(.din(n11622), .dout(n11625));
    jdff dff_B_sQArDvcX8_0(.din(n11625), .dout(n11628));
    jdff dff_A_zNSE46Vu5_0(.din(n11633), .dout(n11630));
    jdff dff_A_V2Fsx7BU9_0(.din(n11636), .dout(n11633));
    jdff dff_A_bvULOijl7_0(.din(n11639), .dout(n11636));
    jdff dff_A_YY2plMGm3_0(.din(n11642), .dout(n11639));
    jdff dff_A_ccwjmVMm4_0(.din(n11645), .dout(n11642));
    jdff dff_A_AmWwTINm2_0(.din(n11648), .dout(n11645));
    jdff dff_A_jj2KitXd6_0(.din(n11651), .dout(n11648));
    jdff dff_A_0QE3QVJE9_0(.din(n11654), .dout(n11651));
    jdff dff_A_rZ7ONRVB7_0(.din(n11657), .dout(n11654));
    jdff dff_A_WEIV3QYS9_0(.din(n11660), .dout(n11657));
    jdff dff_A_rErx2SLH9_0(.din(n11663), .dout(n11660));
    jdff dff_A_gxGqzSXs2_0(.din(n11666), .dout(n11663));
    jdff dff_A_pgjsqp0w8_0(.din(n11669), .dout(n11666));
    jdff dff_A_L8ueDPvO2_0(.din(n6763), .dout(n11669));
    jdff dff_B_CwRSeIak2_1(.din(n6726), .dout(n11673));
    jdff dff_B_JdEVAEq01_1(.din(n11673), .dout(n11676));
    jdff dff_B_9c9ST8518_2(.din(n6722), .dout(n11679));
    jdff dff_B_MdcDDMGE5_2(.din(n11679), .dout(n11682));
    jdff dff_B_oGKanOkl0_2(.din(n11682), .dout(n11685));
    jdff dff_B_NgeIEH9P2_2(.din(n11685), .dout(n11688));
    jdff dff_B_DzNTginG5_2(.din(n11688), .dout(n11691));
    jdff dff_B_eKoW9Bcr7_2(.din(n11691), .dout(n11694));
    jdff dff_B_xKfx4z0l9_2(.din(n11694), .dout(n11697));
    jdff dff_B_47pJCbFJ9_2(.din(n11697), .dout(n11700));
    jdff dff_B_md9S7CLo4_2(.din(n11700), .dout(n11703));
    jdff dff_B_Wug8SRLh9_2(.din(n11703), .dout(n11706));
    jdff dff_B_c5thFNV69_2(.din(n11706), .dout(n11709));
    jdff dff_B_avL0NWVT2_2(.din(n11709), .dout(n11712));
    jdff dff_B_yldM4uHr4_2(.din(n11712), .dout(n11715));
    jdff dff_B_yyCtVycQ4_2(.din(n11715), .dout(n11718));
    jdff dff_B_Fb5PdAwy2_2(.din(n11718), .dout(n11721));
    jdff dff_B_4XwPFce52_2(.din(n11721), .dout(n11724));
    jdff dff_B_SPLC5CPS6_2(.din(n11724), .dout(n11727));
    jdff dff_B_HaKW4JTM6_2(.din(n11727), .dout(n11730));
    jdff dff_B_88C9hQyN6_2(.din(n11730), .dout(n11733));
    jdff dff_B_gda2oCd96_2(.din(n11733), .dout(n11736));
    jdff dff_B_QoPMMl6n7_2(.din(n11736), .dout(n11739));
    jdff dff_B_1DjAqkbo8_2(.din(n11739), .dout(n11742));
    jdff dff_B_EaUyJfyk4_2(.din(n11742), .dout(n11745));
    jdff dff_B_4p0V0LEh8_2(.din(n11745), .dout(n11748));
    jdff dff_B_GwtcKxKR3_2(.din(n11748), .dout(n11751));
    jdff dff_B_8dBBk3Rk7_2(.din(n11751), .dout(n11754));
    jdff dff_B_PMIi69VZ4_2(.din(n11754), .dout(n11757));
    jdff dff_B_GMkvc1yV0_2(.din(n11757), .dout(n11760));
    jdff dff_B_jO2yocm39_2(.din(n11760), .dout(n11763));
    jdff dff_B_Tv2aRw1p4_2(.din(n11763), .dout(n11766));
    jdff dff_B_6g1LHoz31_2(.din(n11766), .dout(n11769));
    jdff dff_B_dEqZoGSd7_2(.din(n11769), .dout(n11772));
    jdff dff_B_hQI3iIFS4_2(.din(n11772), .dout(n11775));
    jdff dff_B_WO3SNvig4_2(.din(n11775), .dout(n11778));
    jdff dff_B_p620AGEX3_2(.din(n11778), .dout(n11781));
    jdff dff_B_UDwP52Ud7_2(.din(n11781), .dout(n11784));
    jdff dff_B_wsO7XN0l8_2(.din(n11784), .dout(n11787));
    jdff dff_B_TSTtLijB6_2(.din(n11787), .dout(n11790));
    jdff dff_B_ijDm1qaW2_2(.din(n11790), .dout(n11793));
    jdff dff_B_0EXD4U4H2_2(.din(n11793), .dout(n11796));
    jdff dff_B_ia58TNRU7_2(.din(n11796), .dout(n11799));
    jdff dff_B_xNE0itga9_2(.din(n11799), .dout(n11802));
    jdff dff_B_KIGMbyhU2_2(.din(n11802), .dout(n11805));
    jdff dff_B_TrggROkz2_2(.din(n11805), .dout(n11808));
    jdff dff_B_mPZEw0Sx3_2(.din(n11808), .dout(n11811));
    jdff dff_B_2wUTUvBm1_2(.din(n11811), .dout(n11814));
    jdff dff_B_Zbsd94kw5_2(.din(n11814), .dout(n11817));
    jdff dff_B_qUOymOHe4_2(.din(n11817), .dout(n11820));
    jdff dff_B_bPgX9GmS9_2(.din(n11820), .dout(n11823));
    jdff dff_B_9eiVS16e5_2(.din(n11823), .dout(n11826));
    jdff dff_B_gdKuuyar9_2(.din(n11826), .dout(n11829));
    jdff dff_B_iT1HOUD15_2(.din(n11829), .dout(n11832));
    jdff dff_B_pls9ok3V1_2(.din(n11832), .dout(n11835));
    jdff dff_B_Ao8U18wJ8_2(.din(n11835), .dout(n11838));
    jdff dff_B_vA60CrKa1_2(.din(n11838), .dout(n11841));
    jdff dff_B_ulT9deez7_2(.din(n11841), .dout(n11844));
    jdff dff_B_TnNJYkFP3_2(.din(n11844), .dout(n11847));
    jdff dff_B_7cLve7654_1(.din(n6748), .dout(n11850));
    jdff dff_B_B7AqmFwC0_1(.din(n11850), .dout(n11853));
    jdff dff_B_ZBDtyjBf7_1(.din(n11853), .dout(n11856));
    jdff dff_B_nfKhVY6U7_1(.din(n11856), .dout(n11859));
    jdff dff_B_s2zwTIMK9_1(.din(n11859), .dout(n11862));
    jdff dff_B_fH90MPwb5_1(.din(n11862), .dout(n11865));
    jdff dff_B_yYdbQXdC5_1(.din(n11865), .dout(n11868));
    jdff dff_B_kcXlAPcu8_1(.din(n11868), .dout(n11871));
    jdff dff_B_hl3AyHsE8_1(.din(n11871), .dout(n11874));
    jdff dff_B_lViDSS2w3_1(.din(n11874), .dout(n11877));
    jdff dff_B_TIDP2gBH7_1(.din(n11877), .dout(n11880));
    jdff dff_B_Jif6Ryib0_1(.din(n11880), .dout(n11883));
    jdff dff_B_rKvz3qNj9_1(.din(n11883), .dout(n11886));
    jdff dff_B_NTsVBm794_0(.din(n6751), .dout(n11889));
    jdff dff_B_X3m0Mhqr1_0(.din(n11889), .dout(n11892));
    jdff dff_B_JJsjNdCn2_0(.din(n11892), .dout(n11895));
    jdff dff_B_xpjB9u8B6_0(.din(n11895), .dout(n11898));
    jdff dff_B_fMFD8vZA7_0(.din(n11898), .dout(n11901));
    jdff dff_B_XbszIEMB1_0(.din(n11901), .dout(n11904));
    jdff dff_B_pdpPE8Ce2_0(.din(n11904), .dout(n11907));
    jdff dff_B_uFpunoN25_0(.din(n11907), .dout(n11910));
    jdff dff_B_Bz1ltoA82_0(.din(n11910), .dout(n11913));
    jdff dff_B_1vNNiMQ23_0(.din(n11913), .dout(n11916));
    jdff dff_B_oT7xWidf7_0(.din(n11916), .dout(n11919));
    jdff dff_B_uG0G052K0_0(.din(n11919), .dout(n11922));
    jdff dff_A_WPGvsqm03_1(.din(n11927), .dout(n11924));
    jdff dff_A_hETNtujh0_1(.din(n11930), .dout(n11927));
    jdff dff_A_78BxAME50_1(.din(n11933), .dout(n11930));
    jdff dff_A_KFoJGfPx5_1(.din(n11936), .dout(n11933));
    jdff dff_A_TzyQriov7_1(.din(n11939), .dout(n11936));
    jdff dff_A_SczVSiE31_1(.din(n11942), .dout(n11939));
    jdff dff_A_DqlTu6MF6_1(.din(n11945), .dout(n11942));
    jdff dff_A_MSz7eijY0_1(.din(n11948), .dout(n11945));
    jdff dff_A_yQFGxJ9h3_1(.din(n11951), .dout(n11948));
    jdff dff_A_Mgt8YJNu3_1(.din(n11954), .dout(n11951));
    jdff dff_A_hP7rHZ7F3_1(.din(n11957), .dout(n11954));
    jdff dff_A_rstKqXmV5_1(.din(n11960), .dout(n11957));
    jdff dff_A_bKLg2vTL0_1(.din(n6714), .dout(n11960));
    jdff dff_B_YmazJ7807_1(.din(n6656), .dout(n11964));
    jdff dff_B_bGUZDYX04_1(.din(n11964), .dout(n11967));
    jdff dff_B_LjhZY2LC8_1(.din(n11967), .dout(n11970));
    jdff dff_B_LrYV5Ntu7_1(.din(n11970), .dout(n11973));
    jdff dff_B_oawRA7Kw5_1(.din(n11973), .dout(n11976));
    jdff dff_B_8vfzK27C1_1(.din(n11976), .dout(n11979));
    jdff dff_B_aKUpKm3y4_1(.din(n11979), .dout(n11982));
    jdff dff_B_RFLUSRNx9_1(.din(n11982), .dout(n11985));
    jdff dff_B_iDbRK6Ty8_1(.din(n11985), .dout(n11988));
    jdff dff_B_ix4VJOmh3_1(.din(n11988), .dout(n11991));
    jdff dff_B_JpgOkr6L9_1(.din(n11991), .dout(n11994));
    jdff dff_B_mwwiw5lE1_1(.din(n11994), .dout(n11997));
    jdff dff_B_yRWuqKkw5_1(.din(n11997), .dout(n12000));
    jdff dff_B_GnbcdT6s3_0(.din(n6659), .dout(n12003));
    jdff dff_B_PQTROi1O5_0(.din(n12003), .dout(n12006));
    jdff dff_B_fXrwwZH15_0(.din(n12006), .dout(n12009));
    jdff dff_B_2Mux3wgO2_0(.din(n12009), .dout(n12012));
    jdff dff_B_pwpySj0Q4_0(.din(n12012), .dout(n12015));
    jdff dff_B_Ys9Lr5Gk2_0(.din(n12015), .dout(n12018));
    jdff dff_B_YKptjCab5_0(.din(n12018), .dout(n12021));
    jdff dff_B_8sy3xX1L0_0(.din(n12021), .dout(n12024));
    jdff dff_B_7XPHU3ij2_0(.din(n12024), .dout(n12027));
    jdff dff_B_6MQAk3Jk8_0(.din(n12027), .dout(n12030));
    jdff dff_B_Ue28N7Wt2_0(.din(n12030), .dout(n12033));
    jdff dff_B_ZeYPt54T0_0(.din(n12033), .dout(n12036));
    jdff dff_A_DRe20etP5_1(.din(n12041), .dout(n12038));
    jdff dff_A_Payo0NRM4_1(.din(n12044), .dout(n12041));
    jdff dff_A_NCnB7HKx1_1(.din(n12047), .dout(n12044));
    jdff dff_A_xtky17vQ9_1(.din(n12050), .dout(n12047));
    jdff dff_A_76v08Zms2_1(.din(n12053), .dout(n12050));
    jdff dff_A_GHVd2Zyw9_1(.din(n12056), .dout(n12053));
    jdff dff_A_J7RdBkdz0_1(.din(n12059), .dout(n12056));
    jdff dff_A_r3anLi1b9_1(.din(n12062), .dout(n12059));
    jdff dff_A_1l4xKHte9_1(.din(n12065), .dout(n12062));
    jdff dff_A_BzNfuLlh3_1(.din(n12068), .dout(n12065));
    jdff dff_A_9SNYp1wM0_1(.din(n12071), .dout(n12068));
    jdff dff_A_Rjsuyn4I3_1(.din(n12074), .dout(n12071));
    jdff dff_A_7qFQCJai5_1(.din(n6642), .dout(n12074));
    jdff dff_B_eNlUkgVG5_1(.din(n6557), .dout(n12078));
    jdff dff_B_YWAHMO8q9_1(.din(n12078), .dout(n12081));
    jdff dff_B_dtiGdofG0_1(.din(n12081), .dout(n12084));
    jdff dff_B_4duU7BmE7_1(.din(n12084), .dout(n12087));
    jdff dff_B_Z8govWyO5_1(.din(n12087), .dout(n12090));
    jdff dff_B_HzdqHQ8b1_1(.din(n12090), .dout(n12093));
    jdff dff_B_49hZUSiv5_1(.din(n12093), .dout(n12096));
    jdff dff_B_yBNeNkrt9_1(.din(n12096), .dout(n12099));
    jdff dff_B_NV8Mmotu3_1(.din(n12099), .dout(n12102));
    jdff dff_B_UfNvOxqL0_1(.din(n12102), .dout(n12105));
    jdff dff_B_DuRBjKw84_1(.din(n12105), .dout(n12108));
    jdff dff_B_JQXNLPIO4_1(.din(n12108), .dout(n12111));
    jdff dff_B_7RvKsDtP2_1(.din(n12111), .dout(n12114));
    jdff dff_B_amPhIF7z0_0(.din(n6560), .dout(n12117));
    jdff dff_B_0jufnKom3_0(.din(n12117), .dout(n12120));
    jdff dff_B_FhmQjCn73_0(.din(n12120), .dout(n12123));
    jdff dff_B_HT2msORh7_0(.din(n12123), .dout(n12126));
    jdff dff_B_RkqyehRP2_0(.din(n12126), .dout(n12129));
    jdff dff_B_NSVuilWk4_0(.din(n12129), .dout(n12132));
    jdff dff_B_RNWkcmDE6_0(.din(n12132), .dout(n12135));
    jdff dff_B_mRCXoC721_0(.din(n12135), .dout(n12138));
    jdff dff_B_P1j5d9o49_0(.din(n12138), .dout(n12141));
    jdff dff_B_gmYC9GAI3_0(.din(n12141), .dout(n12144));
    jdff dff_B_DpBUIqX74_0(.din(n12144), .dout(n12147));
    jdff dff_B_uwUQSseo9_0(.din(n12147), .dout(n12150));
    jdff dff_A_tVT1kRa81_1(.din(n12155), .dout(n12152));
    jdff dff_A_m27y9gzO1_1(.din(n12158), .dout(n12155));
    jdff dff_A_xd4Zz27l4_1(.din(n12161), .dout(n12158));
    jdff dff_A_Kc73B2Dy1_1(.din(n12164), .dout(n12161));
    jdff dff_A_Imk16Ha12_1(.din(n12167), .dout(n12164));
    jdff dff_A_rcnkaNm23_1(.din(n12170), .dout(n12167));
    jdff dff_A_iChtqyvu4_1(.din(n12173), .dout(n12170));
    jdff dff_A_ThzbdRSI1_1(.din(n12176), .dout(n12173));
    jdff dff_A_jm8Lkqrz0_1(.din(n12179), .dout(n12176));
    jdff dff_A_e6Ndbnko0_1(.din(n12182), .dout(n12179));
    jdff dff_A_kMsrLRUe9_1(.din(n12185), .dout(n12182));
    jdff dff_A_oPgmPD5s8_1(.din(n12188), .dout(n12185));
    jdff dff_A_RXQQeR0j4_1(.din(n6543), .dout(n12188));
    jdff dff_B_Nxv2lKfY3_1(.din(n6431), .dout(n12192));
    jdff dff_B_Svgiq7dL8_1(.din(n12192), .dout(n12195));
    jdff dff_B_90TNmHwt5_1(.din(n12195), .dout(n12198));
    jdff dff_B_FrOJXGS59_1(.din(n12198), .dout(n12201));
    jdff dff_B_sxy5MF9o5_1(.din(n12201), .dout(n12204));
    jdff dff_B_Nq6ZbYhD8_1(.din(n12204), .dout(n12207));
    jdff dff_B_hj7KsYkM8_1(.din(n12207), .dout(n12210));
    jdff dff_B_EuXoRDHk3_1(.din(n12210), .dout(n12213));
    jdff dff_B_SD6C0Zyb9_1(.din(n12213), .dout(n12216));
    jdff dff_B_N8NeO2o61_1(.din(n12216), .dout(n12219));
    jdff dff_B_GRBTspeu4_1(.din(n12219), .dout(n12222));
    jdff dff_B_mLqofTnu3_1(.din(n12222), .dout(n12225));
    jdff dff_B_gEpp6YSE9_1(.din(n12225), .dout(n12228));
    jdff dff_B_5xmx5qGV8_0(.din(n6434), .dout(n12231));
    jdff dff_B_eLSVE3a04_0(.din(n12231), .dout(n12234));
    jdff dff_B_gncrlQUf1_0(.din(n12234), .dout(n12237));
    jdff dff_B_uOqhqrZZ5_0(.din(n12237), .dout(n12240));
    jdff dff_B_Uh3br8OP1_0(.din(n12240), .dout(n12243));
    jdff dff_B_sNHTtnzO9_0(.din(n12243), .dout(n12246));
    jdff dff_B_BzJNnD1D7_0(.din(n12246), .dout(n12249));
    jdff dff_B_BH4Of6eP9_0(.din(n12249), .dout(n12252));
    jdff dff_B_aVgAbiVL2_0(.din(n12252), .dout(n12255));
    jdff dff_B_A9IBnHUG1_0(.din(n12255), .dout(n12258));
    jdff dff_B_CZSJDSlp4_0(.din(n12258), .dout(n12261));
    jdff dff_B_CZ6KcnlD1_0(.din(n12261), .dout(n12264));
    jdff dff_A_Xqu6oyos0_1(.din(n12269), .dout(n12266));
    jdff dff_A_FZsRS98w9_1(.din(n12272), .dout(n12269));
    jdff dff_A_c2ocHHsM0_1(.din(n12275), .dout(n12272));
    jdff dff_A_4hJbz2qi8_1(.din(n12278), .dout(n12275));
    jdff dff_A_UMsmR2nH5_1(.din(n12281), .dout(n12278));
    jdff dff_A_XA7goTYL7_1(.din(n12284), .dout(n12281));
    jdff dff_A_zak9b8nx1_1(.din(n12287), .dout(n12284));
    jdff dff_A_6AwDm7zx1_1(.din(n12290), .dout(n12287));
    jdff dff_A_ZVsb9R9N5_1(.din(n12293), .dout(n12290));
    jdff dff_A_3MqrD0346_1(.din(n12296), .dout(n12293));
    jdff dff_A_y6QKNNti8_1(.din(n12299), .dout(n12296));
    jdff dff_A_9f82srkK4_1(.din(n12302), .dout(n12299));
    jdff dff_A_5HE7nm6i7_1(.din(n6417), .dout(n12302));
    jdff dff_B_NiDVM0IL5_1(.din(n6278), .dout(n12306));
    jdff dff_B_THVXFYeH5_1(.din(n12306), .dout(n12309));
    jdff dff_B_7I4s2tqs1_1(.din(n12309), .dout(n12312));
    jdff dff_B_RMbF241J6_1(.din(n12312), .dout(n12315));
    jdff dff_B_BmFgoTeU9_1(.din(n12315), .dout(n12318));
    jdff dff_B_DTPtxRqV5_1(.din(n12318), .dout(n12321));
    jdff dff_B_U4l6Lo1O8_1(.din(n12321), .dout(n12324));
    jdff dff_B_opdsPIUC0_1(.din(n12324), .dout(n12327));
    jdff dff_B_R2IaWWdf9_1(.din(n12327), .dout(n12330));
    jdff dff_B_CfiCXOBP8_1(.din(n12330), .dout(n12333));
    jdff dff_B_d17h1mHL1_1(.din(n12333), .dout(n12336));
    jdff dff_B_mKcOYGMj2_1(.din(n12336), .dout(n12339));
    jdff dff_B_BJyvovda8_1(.din(n12339), .dout(n12342));
    jdff dff_B_PHS5PLeG6_0(.din(n6281), .dout(n12345));
    jdff dff_B_JIpurjGO8_0(.din(n12345), .dout(n12348));
    jdff dff_B_sG6rwZFY1_0(.din(n12348), .dout(n12351));
    jdff dff_B_oBhBHtF84_0(.din(n12351), .dout(n12354));
    jdff dff_B_OdtYtcLg4_0(.din(n12354), .dout(n12357));
    jdff dff_B_xsNTFTtr1_0(.din(n12357), .dout(n12360));
    jdff dff_B_WNGqTnbW3_0(.din(n12360), .dout(n12363));
    jdff dff_B_FKsoa0ir1_0(.din(n12363), .dout(n12366));
    jdff dff_B_RQHNHvPB1_0(.din(n12366), .dout(n12369));
    jdff dff_B_hxzfebwW3_0(.din(n12369), .dout(n12372));
    jdff dff_B_OfOjkk3r2_0(.din(n12372), .dout(n12375));
    jdff dff_A_vpGPPpDK3_1(.din(n12380), .dout(n12377));
    jdff dff_A_pSKzezHl3_1(.din(n12383), .dout(n12380));
    jdff dff_A_Rusjejt27_1(.din(n12386), .dout(n12383));
    jdff dff_A_M9euufRg3_1(.din(n12389), .dout(n12386));
    jdff dff_A_eRHyMjoD2_1(.din(n12392), .dout(n12389));
    jdff dff_A_PVXk5nwi7_1(.din(n12395), .dout(n12392));
    jdff dff_A_MfpC0Ifo4_1(.din(n12398), .dout(n12395));
    jdff dff_A_hMwGH2CM1_1(.din(n12401), .dout(n12398));
    jdff dff_A_Ybb0AtZm0_1(.din(n12404), .dout(n12401));
    jdff dff_A_aXTdrMCm9_1(.din(n12407), .dout(n12404));
    jdff dff_A_S3s5DZjn4_1(.din(n12410), .dout(n12407));
    jdff dff_A_tcFSoMZz5_1(.din(n6270), .dout(n12410));
    jdff dff_B_e3ghwwLt7_1(.din(n6095), .dout(n12414));
    jdff dff_B_L9j5KGTg7_1(.din(n12414), .dout(n12417));
    jdff dff_B_2GY2a0XT6_1(.din(n12417), .dout(n12420));
    jdff dff_B_HVPxgTXN8_1(.din(n12420), .dout(n12423));
    jdff dff_B_mJSyy9Rn2_1(.din(n12423), .dout(n12426));
    jdff dff_B_Aigm1sfF2_1(.din(n12426), .dout(n12429));
    jdff dff_B_s606KOLh5_1(.din(n12429), .dout(n12432));
    jdff dff_B_OF9NdZiU4_1(.din(n12432), .dout(n12435));
    jdff dff_B_xoSSOig16_1(.din(n12435), .dout(n12438));
    jdff dff_B_m1bmlMH42_1(.din(n12438), .dout(n12441));
    jdff dff_B_s8cq0cag8_1(.din(n12441), .dout(n12444));
    jdff dff_B_Dr5rfgtG5_1(.din(n12444), .dout(n12447));
    jdff dff_B_D1a7pTL46_0(.din(n6098), .dout(n12450));
    jdff dff_B_OyFgyPyf2_0(.din(n12450), .dout(n12453));
    jdff dff_B_3Ws6aF4L7_0(.din(n12453), .dout(n12456));
    jdff dff_B_ymzlpt8I1_0(.din(n12456), .dout(n12459));
    jdff dff_B_OnHE1AtY9_0(.din(n12459), .dout(n12462));
    jdff dff_B_1oA95bXm2_0(.din(n12462), .dout(n12465));
    jdff dff_B_dgtYZbqV3_0(.din(n12465), .dout(n12468));
    jdff dff_B_Jo74UEam3_0(.din(n12468), .dout(n12471));
    jdff dff_B_0nBRYLJG4_0(.din(n12471), .dout(n12474));
    jdff dff_B_Dmfo7PaF5_0(.din(n12474), .dout(n12477));
    jdff dff_A_4gYtos4m5_1(.din(n12482), .dout(n12479));
    jdff dff_A_FV8rHZS99_1(.din(n12485), .dout(n12482));
    jdff dff_A_ydxLPViJ9_1(.din(n12488), .dout(n12485));
    jdff dff_A_dhhiH5bd2_1(.din(n12491), .dout(n12488));
    jdff dff_A_Vcc0JimF0_1(.din(n12494), .dout(n12491));
    jdff dff_A_V8eDVjaH6_1(.din(n12497), .dout(n12494));
    jdff dff_A_GwGo1QBI6_1(.din(n12500), .dout(n12497));
    jdff dff_A_njHiTBld0_1(.din(n12503), .dout(n12500));
    jdff dff_A_S8IsL0Ib0_1(.din(n12506), .dout(n12503));
    jdff dff_A_DhK7EMWn8_1(.din(n12509), .dout(n12506));
    jdff dff_A_0iecNvAh2_1(.din(n6087), .dout(n12509));
    jdff dff_B_LJJlWnk41_1(.din(n5885), .dout(n12513));
    jdff dff_B_3piuALWv7_1(.din(n12513), .dout(n12516));
    jdff dff_B_oTDNCRoU0_1(.din(n12516), .dout(n12519));
    jdff dff_B_9Cz1FamL9_1(.din(n12519), .dout(n12522));
    jdff dff_B_Ag025cPL1_1(.din(n12522), .dout(n12525));
    jdff dff_B_lk0hO8Yq2_1(.din(n12525), .dout(n12528));
    jdff dff_B_Z6oXm97H1_1(.din(n12528), .dout(n12531));
    jdff dff_B_WQEF9ekj2_1(.din(n12531), .dout(n12534));
    jdff dff_B_hmfNt6b79_1(.din(n12534), .dout(n12537));
    jdff dff_B_fPT3ph2e2_1(.din(n12537), .dout(n12540));
    jdff dff_B_lxy4xvBU3_0(.din(n5888), .dout(n12543));
    jdff dff_B_zpgqweIC2_0(.din(n12543), .dout(n12546));
    jdff dff_B_PrMF6BJ27_0(.din(n12546), .dout(n12549));
    jdff dff_B_dNHn36ia0_0(.din(n12549), .dout(n12552));
    jdff dff_B_dMpuQB7g0_0(.din(n12552), .dout(n12555));
    jdff dff_B_vyKnG3id5_0(.din(n12555), .dout(n12558));
    jdff dff_B_FU2qZ6LP7_0(.din(n12558), .dout(n12561));
    jdff dff_B_7MkU68A62_0(.din(n12561), .dout(n12564));
    jdff dff_A_MRcvc1uA4_1(.din(n12569), .dout(n12566));
    jdff dff_A_yu7UUQFT7_1(.din(n12572), .dout(n12569));
    jdff dff_A_OthvHi1X1_1(.din(n12575), .dout(n12572));
    jdff dff_A_bF84zSeK2_1(.din(n12578), .dout(n12575));
    jdff dff_A_ENBa59xu0_1(.din(n12581), .dout(n12578));
    jdff dff_A_1h5GEteT0_1(.din(n12584), .dout(n12581));
    jdff dff_A_Usz5I9JG5_1(.din(n12587), .dout(n12584));
    jdff dff_A_2sHKpfZJ6_1(.din(n12590), .dout(n12587));
    jdff dff_A_xuraak5w1_1(.din(n5877), .dout(n12590));
    jdff dff_B_ufxgNgqS8_1(.din(n5648), .dout(n12594));
    jdff dff_B_ztb9utD51_1(.din(n12594), .dout(n12597));
    jdff dff_B_kKiGYkkF8_1(.din(n12597), .dout(n12600));
    jdff dff_B_FLJ4YpMp7_1(.din(n12600), .dout(n12603));
    jdff dff_B_sDoBt1Vb4_1(.din(n12603), .dout(n12606));
    jdff dff_B_pgsVoisl2_1(.din(n12606), .dout(n12609));
    jdff dff_B_wJdjq6UD9_1(.din(n12609), .dout(n12612));
    jdff dff_B_la4C7ecR3_1(.din(n12612), .dout(n12615));
    jdff dff_B_dWAYz2Rc7_0(.din(n5651), .dout(n12618));
    jdff dff_B_1epMpAng0_0(.din(n12618), .dout(n12621));
    jdff dff_B_Bz65Kcuo5_0(.din(n12621), .dout(n12624));
    jdff dff_B_98FrXcK27_0(.din(n12624), .dout(n12627));
    jdff dff_B_5zVSnA2z6_0(.din(n12627), .dout(n12630));
    jdff dff_B_NW2B2g9Z9_0(.din(n12630), .dout(n12633));
    jdff dff_A_XFDpb1RG5_1(.din(n12638), .dout(n12635));
    jdff dff_A_3JmpqIru4_1(.din(n12641), .dout(n12638));
    jdff dff_A_xbN7cE4m9_1(.din(n12644), .dout(n12641));
    jdff dff_A_AGCUTb3e5_1(.din(n12647), .dout(n12644));
    jdff dff_A_o1mjaOtS0_1(.din(n12650), .dout(n12647));
    jdff dff_A_CzaZjN317_1(.din(n12653), .dout(n12650));
    jdff dff_A_G45fXfk25_1(.din(n5640), .dout(n12653));
    jdff dff_B_99jEtv879_1(.din(n5384), .dout(n12657));
    jdff dff_B_RwJTWK5E1_1(.din(n12657), .dout(n12660));
    jdff dff_B_D62o8hER1_1(.din(n12660), .dout(n12663));
    jdff dff_B_JohTtuWZ5_1(.din(n12663), .dout(n12666));
    jdff dff_B_zctOC7Yx2_1(.din(n12666), .dout(n12669));
    jdff dff_B_u2wEuWIl8_1(.din(n12669), .dout(n12672));
    jdff dff_B_6M8TUMrb7_1(.din(n12672), .dout(n12675));
    jdff dff_B_uzcjNXjC1_0(.din(n5387), .dout(n12678));
    jdff dff_B_zq4uOzPE2_0(.din(n12678), .dout(n12681));
    jdff dff_B_7hI0vCHj9_0(.din(n12681), .dout(n12684));
    jdff dff_B_HrYEjpWa5_0(.din(n12684), .dout(n12687));
    jdff dff_B_HRfc0iEy8_0(.din(n12687), .dout(n12690));
    jdff dff_A_Lrjqb8Q71_1(.din(n12695), .dout(n12692));
    jdff dff_A_ggzCto9m0_1(.din(n12698), .dout(n12695));
    jdff dff_A_VVPVeflc3_1(.din(n12701), .dout(n12698));
    jdff dff_A_6UoLyPy62_1(.din(n12704), .dout(n12701));
    jdff dff_A_ajr6RC2b0_1(.din(n12707), .dout(n12704));
    jdff dff_A_vTJCgUqr5_1(.din(n5376), .dout(n12707));
    jdff dff_B_DtWOtbt48_1(.din(n5093), .dout(n12711));
    jdff dff_B_x6YGrWCP2_1(.din(n12711), .dout(n12714));
    jdff dff_B_cgKo1uKb5_1(.din(n12714), .dout(n12717));
    jdff dff_B_sNmOolNm6_1(.din(n12717), .dout(n12720));
    jdff dff_B_Ly4X3evK3_1(.din(n12720), .dout(n12723));
    jdff dff_B_5Qqva24S8_1(.din(n12723), .dout(n12726));
    jdff dff_B_0BX5uYEF9_0(.din(n5096), .dout(n12729));
    jdff dff_B_b6oP3IBR6_0(.din(n12729), .dout(n12732));
    jdff dff_B_2pCn1TmJ8_0(.din(n12732), .dout(n12735));
    jdff dff_B_ZlZ6Nbus7_0(.din(n12735), .dout(n12738));
    jdff dff_A_4ONEt3wy6_1(.din(n12743), .dout(n12740));
    jdff dff_A_2j2h0TO31_1(.din(n12746), .dout(n12743));
    jdff dff_A_LPtiH6V44_1(.din(n12749), .dout(n12746));
    jdff dff_A_ytACUHtR0_1(.din(n12752), .dout(n12749));
    jdff dff_A_eCoR4Xyq0_1(.din(n5085), .dout(n12752));
    jdff dff_B_ciEhE5oa1_1(.din(n4778), .dout(n12756));
    jdff dff_B_CwNbjt9l7_1(.din(n12756), .dout(n12759));
    jdff dff_B_kUkGjYFU6_1(.din(n12759), .dout(n12762));
    jdff dff_A_LFIfuljK0_0(.din(n12767), .dout(n12764));
    jdff dff_A_HSElSoIF5_0(.din(n4764), .dout(n12767));
    jdff dff_B_4lbaaL8i8_1(.din(n4439), .dout(n12771));
    jdff dff_A_PYphhLrQ4_0(.din(n4425), .dout(n12773));
    jdff dff_B_RwNnqVnb6_1(.din(n4064), .dout(n12777));
    jdff dff_A_0ILHXRq21_1(.din(n3679), .dout(n12779));
    jdff dff_B_T4lBY7sl2_2(.din(n3671), .dout(n12783));
    jdff dff_B_4xi7J29C7_1(.din(n3278), .dout(n12786));
    jdff dff_A_7wZHuWQL2_0(.din(n12791), .dout(n12788));
    jdff dff_A_6cJ0fW5k2_0(.din(n12794), .dout(n12791));
    jdff dff_A_uhSwwA6H0_0(.din(n12797), .dout(n12794));
    jdff dff_A_f0TEMAuq8_0(.din(n12800), .dout(n12797));
    jdff dff_A_h7EAVs6D4_0(.din(n12803), .dout(n12800));
    jdff dff_A_rq093ssw9_0(.din(n12806), .dout(n12803));
    jdff dff_A_tdctkbOV7_0(.din(n12809), .dout(n12806));
    jdff dff_A_IRIJoYKg8_0(.din(n12812), .dout(n12809));
    jdff dff_A_x3REjARl0_0(.din(n12815), .dout(n12812));
    jdff dff_A_BnG97WkD2_0(.din(n12818), .dout(n12815));
    jdff dff_A_519OxtWA7_0(.din(n12821), .dout(n12818));
    jdff dff_A_GUR3HTEq2_0(.din(n12824), .dout(n12821));
    jdff dff_A_Ol7f7Yt26_0(.din(n12827), .dout(n12824));
    jdff dff_A_qEkqeOYb4_0(.din(n12830), .dout(n12827));
    jdff dff_A_p7tFtE577_0(.din(n12833), .dout(n12830));
    jdff dff_A_ZBV2MSCJ5_0(.din(n12836), .dout(n12833));
    jdff dff_A_Ye1uCfar5_0(.din(n12839), .dout(n12836));
    jdff dff_A_U3V8u78H4_0(.din(n12842), .dout(n12839));
    jdff dff_A_pvdl4QGc7_0(.din(n12845), .dout(n12842));
    jdff dff_A_hJ8zBZk38_0(.din(n12848), .dout(n12845));
    jdff dff_A_UAq6hRJH3_0(.din(n12851), .dout(n12848));
    jdff dff_A_NGo2YtPo8_0(.din(n12854), .dout(n12851));
    jdff dff_A_2sVv8gC40_0(.din(n12857), .dout(n12854));
    jdff dff_A_G5Ho0abw3_0(.din(n12860), .dout(n12857));
    jdff dff_A_zQaSjH4w4_0(.din(n12863), .dout(n12860));
    jdff dff_A_6vw6P3qt7_0(.din(n12866), .dout(n12863));
    jdff dff_A_fSUzXhIk9_0(.din(n12869), .dout(n12866));
    jdff dff_A_5ulZx8a16_0(.din(n12872), .dout(n12869));
    jdff dff_A_VItp2do45_0(.din(n12875), .dout(n12872));
    jdff dff_A_xLxnb5Pd4_0(.din(n12878), .dout(n12875));
    jdff dff_A_mADrcsg95_0(.din(n12881), .dout(n12878));
    jdff dff_A_gL54cPH75_0(.din(n12884), .dout(n12881));
    jdff dff_A_IORHVl6G9_0(.din(n12887), .dout(n12884));
    jdff dff_A_TyhxclkV9_0(.din(n12890), .dout(n12887));
    jdff dff_A_3vCRfo9D2_0(.din(n12893), .dout(n12890));
    jdff dff_A_DWvgFadZ6_0(.din(n12896), .dout(n12893));
    jdff dff_A_yC5md7O78_0(.din(n12899), .dout(n12896));
    jdff dff_A_Pamahlte9_0(.din(n12902), .dout(n12899));
    jdff dff_A_SlVhe1Ga5_0(.din(n12905), .dout(n12902));
    jdff dff_A_ozVsdxvV6_0(.din(n12908), .dout(n12905));
    jdff dff_A_2j9truBF6_0(.din(n12911), .dout(n12908));
    jdff dff_A_nCOFFhXa2_0(.din(n12914), .dout(n12911));
    jdff dff_A_fOMSH2Sk7_0(.din(n2883), .dout(n12914));
    jdff dff_A_ra8b89sL4_1(.din(n3263), .dout(n12917));
    jdff dff_B_fUgsaO6R2_1(.din(n2893), .dout(n12921));
    jdff dff_A_9MiIiI5w5_0(.din(n12926), .dout(n12923));
    jdff dff_A_waEKkhjf6_0(.din(n12929), .dout(n12926));
    jdff dff_A_69ytUQ3A2_0(.din(n12932), .dout(n12929));
    jdff dff_A_cricFCtc1_0(.din(n12935), .dout(n12932));
    jdff dff_A_FqntZ5Tl4_0(.din(n12938), .dout(n12935));
    jdff dff_A_BDf71oEe9_0(.din(n12941), .dout(n12938));
    jdff dff_A_VV4S4COs5_0(.din(n12944), .dout(n12941));
    jdff dff_A_iEuW9GLf4_0(.din(n12947), .dout(n12944));
    jdff dff_A_wGF92iH39_0(.din(n12950), .dout(n12947));
    jdff dff_A_0cM9jCbq7_0(.din(n12953), .dout(n12950));
    jdff dff_A_1RFis5Qd1_0(.din(n12956), .dout(n12953));
    jdff dff_A_M7FYKQnL0_0(.din(n12959), .dout(n12956));
    jdff dff_A_ZuQNXriM2_0(.din(n12962), .dout(n12959));
    jdff dff_A_A8vXEfk04_0(.din(n12965), .dout(n12962));
    jdff dff_A_fHoQzASn9_0(.din(n12968), .dout(n12965));
    jdff dff_A_q3L2bRJV4_0(.din(n12971), .dout(n12968));
    jdff dff_A_BHblP0pF8_0(.din(n12974), .dout(n12971));
    jdff dff_A_80Ax4HiU1_0(.din(n12977), .dout(n12974));
    jdff dff_A_a7bQXuza9_0(.din(n12980), .dout(n12977));
    jdff dff_A_d3Gl7lLy4_0(.din(n12983), .dout(n12980));
    jdff dff_A_meFxOqsl9_0(.din(n12986), .dout(n12983));
    jdff dff_A_S2lwdrPZ8_0(.din(n12989), .dout(n12986));
    jdff dff_A_y5gs4Hco1_0(.din(n12992), .dout(n12989));
    jdff dff_A_2QmPDKaM1_0(.din(n12995), .dout(n12992));
    jdff dff_A_82jbZI446_0(.din(n12998), .dout(n12995));
    jdff dff_A_rK3tfZIg7_0(.din(n13001), .dout(n12998));
    jdff dff_A_UAWSx7hy1_0(.din(n13004), .dout(n13001));
    jdff dff_A_Ko96IlfN0_0(.din(n13007), .dout(n13004));
    jdff dff_A_j9RYdZ2H2_0(.din(n13010), .dout(n13007));
    jdff dff_A_Q0cTpnbQ8_0(.din(n13013), .dout(n13010));
    jdff dff_A_wNsxdpsx3_0(.din(n13016), .dout(n13013));
    jdff dff_A_avqQY4bb2_0(.din(n13019), .dout(n13016));
    jdff dff_A_infK8D7j8_0(.din(n13022), .dout(n13019));
    jdff dff_A_pbCOyc8h0_0(.din(n13025), .dout(n13022));
    jdff dff_A_DtMsdpwU6_0(.din(n13028), .dout(n13025));
    jdff dff_A_A5FpTrrD7_0(.din(n13031), .dout(n13028));
    jdff dff_A_CVFsShbn7_0(.din(n13034), .dout(n13031));
    jdff dff_A_75sGKR2N7_0(.din(n13037), .dout(n13034));
    jdff dff_A_juJ0YWCi8_0(.din(n13040), .dout(n13037));
    jdff dff_A_Evzuf2IR8_0(.din(n2505), .dout(n13040));
    jdff dff_A_8ocpneNJ7_1(.din(n2871), .dout(n13043));
    jdff dff_B_f2s8ll5S7_1(.din(n2530), .dout(n13047));
    jdff dff_B_7zUKubWB6_1(.din(n13047), .dout(n13050));
    jdff dff_B_g3NAIaP19_1(.din(n13050), .dout(n13053));
    jdff dff_B_zKyZ22v46_1(.din(n13053), .dout(n13056));
    jdff dff_B_mpMOliPw9_1(.din(n13056), .dout(n13059));
    jdff dff_B_bcE9CSpy9_1(.din(n13059), .dout(n13062));
    jdff dff_B_dlzDynoQ1_1(.din(n13062), .dout(n13065));
    jdff dff_B_j0tIeTl78_1(.din(n13065), .dout(n13068));
    jdff dff_B_pLlDu1QI6_1(.din(n13068), .dout(n13071));
    jdff dff_B_IPAGpyNa0_1(.din(n13071), .dout(n13074));
    jdff dff_B_u30lyc8x6_1(.din(n13074), .dout(n13077));
    jdff dff_B_g9Bj4mR33_1(.din(n13077), .dout(n13080));
    jdff dff_B_nKzF8pWz9_1(.din(n13080), .dout(n13083));
    jdff dff_B_TEq6th2s5_1(.din(n13083), .dout(n13086));
    jdff dff_B_nKuV32Vx8_1(.din(n13086), .dout(n13089));
    jdff dff_B_h6kLfVcb0_1(.din(n13089), .dout(n13092));
    jdff dff_B_RiyIr1VH1_1(.din(n13092), .dout(n13095));
    jdff dff_B_Gympt39G8_1(.din(n13095), .dout(n13098));
    jdff dff_B_auS0WcJ65_1(.din(n13098), .dout(n13101));
    jdff dff_B_uHsCIQpA1_1(.din(n13101), .dout(n13104));
    jdff dff_B_pOAFj4aZ1_1(.din(n13104), .dout(n13107));
    jdff dff_B_aYxePEI51_1(.din(n13107), .dout(n13110));
    jdff dff_B_KW18rf0u3_1(.din(n13110), .dout(n13113));
    jdff dff_B_hygbpTQG2_1(.din(n13113), .dout(n13116));
    jdff dff_B_l2DXJUKw7_1(.din(n13116), .dout(n13119));
    jdff dff_B_bpVekJAE0_1(.din(n13119), .dout(n13122));
    jdff dff_B_P0Vt5Ayd2_1(.din(n13122), .dout(n13125));
    jdff dff_B_whaAqAAA6_1(.din(n13125), .dout(n13128));
    jdff dff_B_CGGRfG9D1_1(.din(n13128), .dout(n13131));
    jdff dff_B_jqOp89Qm7_1(.din(n13131), .dout(n13134));
    jdff dff_B_cPDyFdle6_1(.din(n13134), .dout(n13137));
    jdff dff_B_vWgwoJ0C9_1(.din(n13137), .dout(n13140));
    jdff dff_B_WcWjvEIU6_1(.din(n13140), .dout(n13143));
    jdff dff_B_gumcnGAx1_1(.din(n13143), .dout(n13146));
    jdff dff_B_nBj5gObl3_1(.din(n13146), .dout(n13149));
    jdff dff_B_BYWga9r30_1(.din(n13149), .dout(n13152));
    jdff dff_B_fCo7Mjhw4_1(.din(n2515), .dout(n13155));
    jdff dff_A_ZJqsWTE38_0(.din(n13160), .dout(n13157));
    jdff dff_A_DCweRg5G9_0(.din(n13163), .dout(n13160));
    jdff dff_A_hX73WQSW0_0(.din(n13166), .dout(n13163));
    jdff dff_A_USYjXc4M0_0(.din(n13169), .dout(n13166));
    jdff dff_A_ixLA7BGJ6_0(.din(n13172), .dout(n13169));
    jdff dff_A_wxoBXF8s7_0(.din(n13175), .dout(n13172));
    jdff dff_A_qEHhoYL80_0(.din(n13178), .dout(n13175));
    jdff dff_A_cX3KY70c8_0(.din(n13181), .dout(n13178));
    jdff dff_A_ijblW0et0_0(.din(n13184), .dout(n13181));
    jdff dff_A_O56tFSYs1_0(.din(n13187), .dout(n13184));
    jdff dff_A_0qlK8UcB2_0(.din(n13190), .dout(n13187));
    jdff dff_A_0ai6Xu861_0(.din(n13193), .dout(n13190));
    jdff dff_A_c7qtzy478_0(.din(n13196), .dout(n13193));
    jdff dff_A_WcqWStd04_0(.din(n13199), .dout(n13196));
    jdff dff_A_fdY2wFf83_0(.din(n13202), .dout(n13199));
    jdff dff_A_iYs6F8116_0(.din(n13205), .dout(n13202));
    jdff dff_A_T5gWcaLG1_0(.din(n13208), .dout(n13205));
    jdff dff_A_JudO6DsY1_0(.din(n13211), .dout(n13208));
    jdff dff_A_poqCqyYs2_0(.din(n13214), .dout(n13211));
    jdff dff_A_su1z9E7p4_0(.din(n13217), .dout(n13214));
    jdff dff_A_fSXXNJlq9_0(.din(n13220), .dout(n13217));
    jdff dff_A_wEsTfLSH6_0(.din(n13223), .dout(n13220));
    jdff dff_A_xCLZBxnn9_0(.din(n13226), .dout(n13223));
    jdff dff_A_ZGgbvMH67_0(.din(n13229), .dout(n13226));
    jdff dff_A_Sej4oIN88_0(.din(n13232), .dout(n13229));
    jdff dff_A_oyV8gBJ34_0(.din(n13235), .dout(n13232));
    jdff dff_A_l7rrKOUt6_0(.din(n13238), .dout(n13235));
    jdff dff_A_IM9QaROx9_0(.din(n13241), .dout(n13238));
    jdff dff_A_g2VpbbBh7_0(.din(n13244), .dout(n13241));
    jdff dff_A_cx1u4WQ89_0(.din(n13247), .dout(n13244));
    jdff dff_A_e7tTKAds4_0(.din(n13250), .dout(n13247));
    jdff dff_A_XqkBEqQ31_0(.din(n13253), .dout(n13250));
    jdff dff_A_PWjDeHci6_0(.din(n13256), .dout(n13253));
    jdff dff_A_dY0r4lcd6_0(.din(n13259), .dout(n13256));
    jdff dff_A_5BRhJD7N1_0(.din(n13262), .dout(n13259));
    jdff dff_A_vAxDeasC0_0(.din(n13265), .dout(n13262));
    jdff dff_A_QDiMJm2D6_0(.din(n2154), .dout(n13265));
    jdff dff_A_iUY45Q7M8_1(.din(n2493), .dout(n13268));
    jdff dff_B_A9VAm78q2_1(.din(n2179), .dout(n13272));
    jdff dff_B_LzmwLakx0_1(.din(n13272), .dout(n13275));
    jdff dff_B_ZSyUTwRc7_1(.din(n13275), .dout(n13278));
    jdff dff_B_42Ahjxve6_1(.din(n13278), .dout(n13281));
    jdff dff_B_WlzyMSi54_1(.din(n13281), .dout(n13284));
    jdff dff_B_2rCRDrJq6_1(.din(n13284), .dout(n13287));
    jdff dff_B_L977e37d9_1(.din(n13287), .dout(n13290));
    jdff dff_B_6CTHGhie9_1(.din(n13290), .dout(n13293));
    jdff dff_B_cZeONxXS9_1(.din(n13293), .dout(n13296));
    jdff dff_B_JNLUcxS15_1(.din(n13296), .dout(n13299));
    jdff dff_B_LogmgIUp3_1(.din(n13299), .dout(n13302));
    jdff dff_B_mgBfWcrG7_1(.din(n13302), .dout(n13305));
    jdff dff_B_EumMpXXp3_1(.din(n13305), .dout(n13308));
    jdff dff_B_7qv4UN6Y2_1(.din(n13308), .dout(n13311));
    jdff dff_B_gnVaiatE6_1(.din(n13311), .dout(n13314));
    jdff dff_B_mECXKtel3_1(.din(n13314), .dout(n13317));
    jdff dff_B_MIaqtrIC0_1(.din(n13317), .dout(n13320));
    jdff dff_B_3oUq2jOq1_1(.din(n13320), .dout(n13323));
    jdff dff_B_zgz4uphr2_1(.din(n13323), .dout(n13326));
    jdff dff_B_rd9DjhPC2_1(.din(n13326), .dout(n13329));
    jdff dff_B_7AHnIwJO3_1(.din(n13329), .dout(n13332));
    jdff dff_B_V2fvPVmd2_1(.din(n13332), .dout(n13335));
    jdff dff_B_vCZDwaJ74_1(.din(n13335), .dout(n13338));
    jdff dff_B_qLM4d4355_1(.din(n13338), .dout(n13341));
    jdff dff_B_DwxN9Yr58_1(.din(n13341), .dout(n13344));
    jdff dff_B_00rLh3e55_1(.din(n13344), .dout(n13347));
    jdff dff_B_fYR1K5me0_1(.din(n13347), .dout(n13350));
    jdff dff_B_KKRx64nL9_1(.din(n13350), .dout(n13353));
    jdff dff_B_eEHalRt61_1(.din(n13353), .dout(n13356));
    jdff dff_B_vuomH4Em3_1(.din(n13356), .dout(n13359));
    jdff dff_B_m0uvBwCu9_1(.din(n13359), .dout(n13362));
    jdff dff_B_SoQs1uK54_1(.din(n13362), .dout(n13365));
    jdff dff_B_0W0p7jUR3_1(.din(n13365), .dout(n13368));
    jdff dff_B_ZVITaAWb1_1(.din(n2164), .dout(n13371));
    jdff dff_A_nhDvlxFe4_0(.din(n13376), .dout(n13373));
    jdff dff_A_hEzlDyid1_0(.din(n13379), .dout(n13376));
    jdff dff_A_LMN6QWFi3_0(.din(n13382), .dout(n13379));
    jdff dff_A_zdwR896X3_0(.din(n13385), .dout(n13382));
    jdff dff_A_Cmglstuh2_0(.din(n13388), .dout(n13385));
    jdff dff_A_Nl0zI5LZ5_0(.din(n13391), .dout(n13388));
    jdff dff_A_RSNCOae38_0(.din(n13394), .dout(n13391));
    jdff dff_A_N1FfJhoA5_0(.din(n13397), .dout(n13394));
    jdff dff_A_HYh079cz5_0(.din(n13400), .dout(n13397));
    jdff dff_A_tZljyAks7_0(.din(n13403), .dout(n13400));
    jdff dff_A_8X8Jhouy3_0(.din(n13406), .dout(n13403));
    jdff dff_A_Gie4ZqOK9_0(.din(n13409), .dout(n13406));
    jdff dff_A_xgNC3I4N5_0(.din(n13412), .dout(n13409));
    jdff dff_A_iSccoqyV6_0(.din(n13415), .dout(n13412));
    jdff dff_A_boqlekLb4_0(.din(n13418), .dout(n13415));
    jdff dff_A_nOoTvesv8_0(.din(n13421), .dout(n13418));
    jdff dff_A_OuPDWl9o5_0(.din(n13424), .dout(n13421));
    jdff dff_A_IFEyOzj68_0(.din(n13427), .dout(n13424));
    jdff dff_A_hu77U5f90_0(.din(n13430), .dout(n13427));
    jdff dff_A_lIkyySYt0_0(.din(n13433), .dout(n13430));
    jdff dff_A_atsADPc67_0(.din(n13436), .dout(n13433));
    jdff dff_A_6ZuKJLlt6_0(.din(n13439), .dout(n13436));
    jdff dff_A_w7li6z5p6_0(.din(n13442), .dout(n13439));
    jdff dff_A_DmifbVad4_0(.din(n13445), .dout(n13442));
    jdff dff_A_PCxv85Wy7_0(.din(n13448), .dout(n13445));
    jdff dff_A_31BEGkBD1_0(.din(n13451), .dout(n13448));
    jdff dff_A_CFjU7RDm6_0(.din(n13454), .dout(n13451));
    jdff dff_A_2drIfCX83_0(.din(n13457), .dout(n13454));
    jdff dff_A_ek3ulER84_0(.din(n13460), .dout(n13457));
    jdff dff_A_IItxrOUx2_0(.din(n13463), .dout(n13460));
    jdff dff_A_AMAesH8T0_0(.din(n13466), .dout(n13463));
    jdff dff_A_vIpGoxcf1_0(.din(n13469), .dout(n13466));
    jdff dff_A_qHCW8PGe7_0(.din(n13472), .dout(n13469));
    jdff dff_A_bu9jZuxo2_0(.din(n1830), .dout(n13472));
    jdff dff_A_tWZbizCL0_1(.din(n2142), .dout(n13475));
    jdff dff_B_kCHBFrzY0_1(.din(n1855), .dout(n13479));
    jdff dff_B_Rd8TzzGj5_1(.din(n13479), .dout(n13482));
    jdff dff_B_tENXyBbO8_1(.din(n13482), .dout(n13485));
    jdff dff_B_g6xqOmz25_1(.din(n13485), .dout(n13488));
    jdff dff_B_hrUXolzj6_1(.din(n13488), .dout(n13491));
    jdff dff_B_ugocssaZ4_1(.din(n13491), .dout(n13494));
    jdff dff_B_CSr6RIpv1_1(.din(n13494), .dout(n13497));
    jdff dff_B_iBwWptcJ3_1(.din(n13497), .dout(n13500));
    jdff dff_B_Fj0Pwj9V7_1(.din(n13500), .dout(n13503));
    jdff dff_B_ER53Vsgq1_1(.din(n13503), .dout(n13506));
    jdff dff_B_uXHMzpMj3_1(.din(n13506), .dout(n13509));
    jdff dff_B_i2aGU7eZ7_1(.din(n13509), .dout(n13512));
    jdff dff_B_Ko8H580d3_1(.din(n13512), .dout(n13515));
    jdff dff_B_qqmrnoyj5_1(.din(n13515), .dout(n13518));
    jdff dff_B_M5TtD4UT8_1(.din(n13518), .dout(n13521));
    jdff dff_B_gEHEpSTY6_1(.din(n13521), .dout(n13524));
    jdff dff_B_p8LGoybh8_1(.din(n13524), .dout(n13527));
    jdff dff_B_V5hUxEtK1_1(.din(n13527), .dout(n13530));
    jdff dff_B_25lRxmGI1_1(.din(n13530), .dout(n13533));
    jdff dff_B_IyNrAS8v8_1(.din(n13533), .dout(n13536));
    jdff dff_B_y8CD5oan6_1(.din(n13536), .dout(n13539));
    jdff dff_B_748Wehi27_1(.din(n13539), .dout(n13542));
    jdff dff_B_kh3cpPPq2_1(.din(n13542), .dout(n13545));
    jdff dff_B_yOohTYGP9_1(.din(n13545), .dout(n13548));
    jdff dff_B_FEgnCTD95_1(.din(n13548), .dout(n13551));
    jdff dff_B_AnnayLHC9_1(.din(n13551), .dout(n13554));
    jdff dff_B_Uyh8CFlP1_1(.din(n13554), .dout(n13557));
    jdff dff_B_fq7cDSzQ7_1(.din(n13557), .dout(n13560));
    jdff dff_B_9mT4DgtD6_1(.din(n13560), .dout(n13563));
    jdff dff_B_vR0plZ4L4_1(.din(n13563), .dout(n13566));
    jdff dff_B_VXK70yMo3_1(.din(n1840), .dout(n13569));
    jdff dff_A_OTZF4ZFo9_0(.din(n13574), .dout(n13571));
    jdff dff_A_Cb8ck3cf5_0(.din(n13577), .dout(n13574));
    jdff dff_A_N3kcUESC7_0(.din(n13580), .dout(n13577));
    jdff dff_A_fBeDrGu99_0(.din(n13583), .dout(n13580));
    jdff dff_A_hHwR3u782_0(.din(n13586), .dout(n13583));
    jdff dff_A_AUvVvqXm5_0(.din(n13589), .dout(n13586));
    jdff dff_A_OSAg4mRU4_0(.din(n13592), .dout(n13589));
    jdff dff_A_hSXfgab13_0(.din(n13595), .dout(n13592));
    jdff dff_A_aVSZUbVy0_0(.din(n13598), .dout(n13595));
    jdff dff_A_tZZZ0Cgd1_0(.din(n13601), .dout(n13598));
    jdff dff_A_a4zs17Eo1_0(.din(n13604), .dout(n13601));
    jdff dff_A_GcPPHrYn8_0(.din(n13607), .dout(n13604));
    jdff dff_A_vJB0qnwq9_0(.din(n13610), .dout(n13607));
    jdff dff_A_pfhOpkfR0_0(.din(n13613), .dout(n13610));
    jdff dff_A_2QKP8nLj5_0(.din(n13616), .dout(n13613));
    jdff dff_A_lhi8bUCk6_0(.din(n13619), .dout(n13616));
    jdff dff_A_n9iK2LAY2_0(.din(n13622), .dout(n13619));
    jdff dff_A_pCPGAd0k0_0(.din(n13625), .dout(n13622));
    jdff dff_A_AdIacxm98_0(.din(n13628), .dout(n13625));
    jdff dff_A_wi5K90kP1_0(.din(n13631), .dout(n13628));
    jdff dff_A_OzyeiJQp1_0(.din(n13634), .dout(n13631));
    jdff dff_A_IzGg7SBo5_0(.din(n13637), .dout(n13634));
    jdff dff_A_1tXWoT3N0_0(.din(n13640), .dout(n13637));
    jdff dff_A_Yhmi73pX0_0(.din(n13643), .dout(n13640));
    jdff dff_A_HW5x8sja4_0(.din(n13646), .dout(n13643));
    jdff dff_A_JCaxpzaX2_0(.din(n13649), .dout(n13646));
    jdff dff_A_79MTMddy7_0(.din(n13652), .dout(n13649));
    jdff dff_A_bvmvRzxa6_0(.din(n13655), .dout(n13652));
    jdff dff_A_56tZM1Q22_0(.din(n13658), .dout(n13655));
    jdff dff_A_90ofgxfk4_0(.din(n13661), .dout(n13658));
    jdff dff_A_ERRIE9kX2_0(.din(n1533), .dout(n13661));
    jdff dff_A_kiwmOoXQ4_1(.din(n1818), .dout(n13664));
    jdff dff_B_zBMuKWgD3_1(.din(n1558), .dout(n13668));
    jdff dff_B_DnZAdYla3_1(.din(n13668), .dout(n13671));
    jdff dff_B_R4Ar9KN49_1(.din(n13671), .dout(n13674));
    jdff dff_B_KcFTeE4h5_1(.din(n13674), .dout(n13677));
    jdff dff_B_RXR5pRJ54_1(.din(n13677), .dout(n13680));
    jdff dff_B_G6ai8QNX2_1(.din(n13680), .dout(n13683));
    jdff dff_B_LTqYmLE73_1(.din(n13683), .dout(n13686));
    jdff dff_B_c7cHTrDQ1_1(.din(n13686), .dout(n13689));
    jdff dff_B_vwTbbMfu9_1(.din(n13689), .dout(n13692));
    jdff dff_B_qzxyu0aN4_1(.din(n13692), .dout(n13695));
    jdff dff_B_HIYPKxAn3_1(.din(n13695), .dout(n13698));
    jdff dff_B_jU9d4w7i2_1(.din(n13698), .dout(n13701));
    jdff dff_B_4z6oZ8he6_1(.din(n13701), .dout(n13704));
    jdff dff_B_XvF1Glm41_1(.din(n13704), .dout(n13707));
    jdff dff_B_zXNSOptH7_1(.din(n13707), .dout(n13710));
    jdff dff_B_otfm0FSw6_1(.din(n13710), .dout(n13713));
    jdff dff_B_8O76r0r17_1(.din(n13713), .dout(n13716));
    jdff dff_B_UUJVWsuS2_1(.din(n13716), .dout(n13719));
    jdff dff_B_FF4VzAs23_1(.din(n13719), .dout(n13722));
    jdff dff_B_WsWMziBW5_1(.din(n13722), .dout(n13725));
    jdff dff_B_Hwa1W5oB3_1(.din(n13725), .dout(n13728));
    jdff dff_B_uyrPcFlQ2_1(.din(n13728), .dout(n13731));
    jdff dff_B_ODTl2ZlX6_1(.din(n13731), .dout(n13734));
    jdff dff_B_Ak0VIRh19_1(.din(n13734), .dout(n13737));
    jdff dff_B_YezfJTEd4_1(.din(n13737), .dout(n13740));
    jdff dff_B_YrzUY8kt2_1(.din(n13740), .dout(n13743));
    jdff dff_B_YUvxqxm79_1(.din(n13743), .dout(n13746));
    jdff dff_B_LJWEIvt20_1(.din(n1543), .dout(n13749));
    jdff dff_A_xFbdq81z3_0(.din(n13754), .dout(n13751));
    jdff dff_A_FCQ7mtkf0_0(.din(n13757), .dout(n13754));
    jdff dff_A_FEfsb2Wf5_0(.din(n13760), .dout(n13757));
    jdff dff_A_Ri2JnhyP2_0(.din(n13763), .dout(n13760));
    jdff dff_A_RVueaT9M4_0(.din(n13766), .dout(n13763));
    jdff dff_A_6peDFwnx9_0(.din(n13769), .dout(n13766));
    jdff dff_A_4aofisUd7_0(.din(n13772), .dout(n13769));
    jdff dff_A_7GCzgXLn8_0(.din(n13775), .dout(n13772));
    jdff dff_A_SRM2ThGz5_0(.din(n13778), .dout(n13775));
    jdff dff_A_Gqg9NpGL7_0(.din(n13781), .dout(n13778));
    jdff dff_A_TpbmBRl95_0(.din(n13784), .dout(n13781));
    jdff dff_A_Nmm34HsN3_0(.din(n13787), .dout(n13784));
    jdff dff_A_qz0O7cJg1_0(.din(n13790), .dout(n13787));
    jdff dff_A_t4KNzypt8_0(.din(n13793), .dout(n13790));
    jdff dff_A_HYwUUR276_0(.din(n13796), .dout(n13793));
    jdff dff_A_UADPqvIj5_0(.din(n13799), .dout(n13796));
    jdff dff_A_RzRk2Cvz2_0(.din(n13802), .dout(n13799));
    jdff dff_A_TulId1XP1_0(.din(n13805), .dout(n13802));
    jdff dff_A_z1uLUdZy3_0(.din(n13808), .dout(n13805));
    jdff dff_A_kiJJroz33_0(.din(n13811), .dout(n13808));
    jdff dff_A_niUUt0470_0(.din(n13814), .dout(n13811));
    jdff dff_A_G00qHLd81_0(.din(n13817), .dout(n13814));
    jdff dff_A_X0F482pz5_0(.din(n13820), .dout(n13817));
    jdff dff_A_MCwLeiD24_0(.din(n13823), .dout(n13820));
    jdff dff_A_7H8fdpvx4_0(.din(n13826), .dout(n13823));
    jdff dff_A_QCgajTaP8_0(.din(n13829), .dout(n13826));
    jdff dff_A_Cffrl4qT1_0(.din(n13832), .dout(n13829));
    jdff dff_A_mhHgcLc15_0(.din(n1263), .dout(n13832));
    jdff dff_A_RSzIhc3H1_1(.din(n1521), .dout(n13835));
    jdff dff_B_8IzsM0oD3_1(.din(n1288), .dout(n13839));
    jdff dff_B_jL7slHTw7_1(.din(n13839), .dout(n13842));
    jdff dff_B_MxMOhbsl4_1(.din(n13842), .dout(n13845));
    jdff dff_B_kYRKIEJe8_1(.din(n13845), .dout(n13848));
    jdff dff_B_AzhsXSAm8_1(.din(n13848), .dout(n13851));
    jdff dff_B_l27U4c4U9_1(.din(n13851), .dout(n13854));
    jdff dff_B_Y2BR2rwX8_1(.din(n13854), .dout(n13857));
    jdff dff_B_dQ7RhL0j2_1(.din(n13857), .dout(n13860));
    jdff dff_B_M3EBURiR6_1(.din(n13860), .dout(n13863));
    jdff dff_B_wBDy8Uej1_1(.din(n13863), .dout(n13866));
    jdff dff_B_DVoJ7zCR3_1(.din(n13866), .dout(n13869));
    jdff dff_B_S9ZaIGoN3_1(.din(n13869), .dout(n13872));
    jdff dff_B_mc7YIRdA1_1(.din(n13872), .dout(n13875));
    jdff dff_B_ci266ybB5_1(.din(n13875), .dout(n13878));
    jdff dff_B_UWT8ro7g5_1(.din(n13878), .dout(n13881));
    jdff dff_B_QskdNfw20_1(.din(n13881), .dout(n13884));
    jdff dff_B_75B13Y7W2_1(.din(n13884), .dout(n13887));
    jdff dff_B_Ag1D4aU29_1(.din(n13887), .dout(n13890));
    jdff dff_B_15cdKQOx4_1(.din(n13890), .dout(n13893));
    jdff dff_B_5Sw6A1Cq3_1(.din(n13893), .dout(n13896));
    jdff dff_B_7SAOGW3R3_1(.din(n13896), .dout(n13899));
    jdff dff_B_vMg1hHGn4_1(.din(n13899), .dout(n13902));
    jdff dff_B_BGqwVxJj0_1(.din(n13902), .dout(n13905));
    jdff dff_B_o39bPTKi1_1(.din(n13905), .dout(n13908));
    jdff dff_B_qUFUEihJ6_1(.din(n1273), .dout(n13911));
    jdff dff_A_6OLEzaXf3_0(.din(n13916), .dout(n13913));
    jdff dff_A_eY119YXw3_0(.din(n13919), .dout(n13916));
    jdff dff_A_n9av7IQb4_0(.din(n13922), .dout(n13919));
    jdff dff_A_auMVzTH99_0(.din(n13925), .dout(n13922));
    jdff dff_A_XrQEAPYG6_0(.din(n13928), .dout(n13925));
    jdff dff_A_0nzDlDOa0_0(.din(n13931), .dout(n13928));
    jdff dff_A_eSBgJxCX8_0(.din(n13934), .dout(n13931));
    jdff dff_A_Ila1lE2m4_0(.din(n13937), .dout(n13934));
    jdff dff_A_WKUXKNJR6_0(.din(n13940), .dout(n13937));
    jdff dff_A_8xVbUGRS1_0(.din(n13943), .dout(n13940));
    jdff dff_A_MJZC7UVW9_0(.din(n13946), .dout(n13943));
    jdff dff_A_P7rHvVYo6_0(.din(n13949), .dout(n13946));
    jdff dff_A_c9UHDsyl7_0(.din(n13952), .dout(n13949));
    jdff dff_A_ERqEylzL4_0(.din(n13955), .dout(n13952));
    jdff dff_A_MJGTWWdj1_0(.din(n13958), .dout(n13955));
    jdff dff_A_U95dLSqh6_0(.din(n13961), .dout(n13958));
    jdff dff_A_G2zgbwfV5_0(.din(n13964), .dout(n13961));
    jdff dff_A_o2RSMPzA4_0(.din(n13967), .dout(n13964));
    jdff dff_A_RXOCSMT92_0(.din(n13970), .dout(n13967));
    jdff dff_A_WtEesyWf0_0(.din(n13973), .dout(n13970));
    jdff dff_A_vDLIzGEw7_0(.din(n13976), .dout(n13973));
    jdff dff_A_WCsDVMnX1_0(.din(n13979), .dout(n13976));
    jdff dff_A_6vSefmfV5_0(.din(n13982), .dout(n13979));
    jdff dff_A_7HWt21FX3_0(.din(n13985), .dout(n13982));
    jdff dff_A_k1BBpuyE8_0(.din(n1023), .dout(n13985));
    jdff dff_A_Bovu7nZx1_1(.din(n1251), .dout(n13988));
    jdff dff_B_e8GjJcCW9_1(.din(n1048), .dout(n13992));
    jdff dff_B_BuGj6LmC7_1(.din(n13992), .dout(n13995));
    jdff dff_B_RqGqG74g8_1(.din(n13995), .dout(n13998));
    jdff dff_B_WImsQgUi5_1(.din(n13998), .dout(n14001));
    jdff dff_B_vF7Lls0q3_1(.din(n14001), .dout(n14004));
    jdff dff_B_Gy6lrtYG3_1(.din(n14004), .dout(n14007));
    jdff dff_B_eKfU6hzp1_1(.din(n14007), .dout(n14010));
    jdff dff_B_yndFDEJi3_1(.din(n14010), .dout(n14013));
    jdff dff_B_sbJdPLQ23_1(.din(n14013), .dout(n14016));
    jdff dff_B_ibPIAYSx6_1(.din(n14016), .dout(n14019));
    jdff dff_B_feS9UsVx4_1(.din(n14019), .dout(n14022));
    jdff dff_B_FurDQtN38_1(.din(n14022), .dout(n14025));
    jdff dff_B_5HMl790y2_1(.din(n14025), .dout(n14028));
    jdff dff_B_jyvY51ll4_1(.din(n14028), .dout(n14031));
    jdff dff_B_td2FHD193_1(.din(n14031), .dout(n14034));
    jdff dff_B_KbefJUfY2_1(.din(n14034), .dout(n14037));
    jdff dff_B_eBGwZBbY3_1(.din(n14037), .dout(n14040));
    jdff dff_B_WzNbvo4m5_1(.din(n14040), .dout(n14043));
    jdff dff_B_1d3JgBps1_1(.din(n14043), .dout(n14046));
    jdff dff_B_oEH0J9py3_1(.din(n14046), .dout(n14049));
    jdff dff_B_Y7eTPMcT7_1(.din(n14049), .dout(n14052));
    jdff dff_B_P7NpbNA11_1(.din(n1033), .dout(n14055));
    jdff dff_A_D0Qidzpm9_0(.din(n14060), .dout(n14057));
    jdff dff_A_yMczb0lx9_0(.din(n14063), .dout(n14060));
    jdff dff_A_DMy0DIpY8_0(.din(n14066), .dout(n14063));
    jdff dff_A_oiy70Ye71_0(.din(n14069), .dout(n14066));
    jdff dff_A_V1h4Rjwg7_0(.din(n14072), .dout(n14069));
    jdff dff_A_CWeX05oF3_0(.din(n14075), .dout(n14072));
    jdff dff_A_5qC8yfzW7_0(.din(n14078), .dout(n14075));
    jdff dff_A_13OJlsHp3_0(.din(n14081), .dout(n14078));
    jdff dff_A_h5S33M530_0(.din(n14084), .dout(n14081));
    jdff dff_A_poXiEqOV4_0(.din(n14087), .dout(n14084));
    jdff dff_A_5kNhbh6y7_0(.din(n14090), .dout(n14087));
    jdff dff_A_e8JIFoMd9_0(.din(n14093), .dout(n14090));
    jdff dff_A_9EEJxgeo5_0(.din(n14096), .dout(n14093));
    jdff dff_A_ZOgyuoVn7_0(.din(n14099), .dout(n14096));
    jdff dff_A_Cf2f3QFx5_0(.din(n14102), .dout(n14099));
    jdff dff_A_zvRImTZy9_0(.din(n14105), .dout(n14102));
    jdff dff_A_D6LMTFrW8_0(.din(n14108), .dout(n14105));
    jdff dff_A_k7yBVQ1b5_0(.din(n14111), .dout(n14108));
    jdff dff_A_r7j8Heqh9_0(.din(n14114), .dout(n14111));
    jdff dff_A_Hn8yPNAj3_0(.din(n14117), .dout(n14114));
    jdff dff_A_HRlk4xJI7_0(.din(n14120), .dout(n14117));
    jdff dff_A_MScdtDYV3_0(.din(n810), .dout(n14120));
    jdff dff_A_z1v3IO1U1_1(.din(n1011), .dout(n14123));
    jdff dff_B_OatZHRhl5_1(.din(n835), .dout(n14127));
    jdff dff_B_E2m2I4tc4_1(.din(n14127), .dout(n14130));
    jdff dff_B_chenxPSq4_1(.din(n14130), .dout(n14133));
    jdff dff_B_J1Ave9H68_1(.din(n14133), .dout(n14136));
    jdff dff_B_AnLyatS00_1(.din(n14136), .dout(n14139));
    jdff dff_B_FhbxRMqo2_1(.din(n14139), .dout(n14142));
    jdff dff_B_Nns16vPM0_1(.din(n14142), .dout(n14145));
    jdff dff_B_XjGdVqET9_1(.din(n14145), .dout(n14148));
    jdff dff_B_GfNLBomx2_1(.din(n14148), .dout(n14151));
    jdff dff_B_EwLD71nM2_1(.din(n14151), .dout(n14154));
    jdff dff_B_zMiVHBW53_1(.din(n14154), .dout(n14157));
    jdff dff_B_6Z095BjI0_1(.din(n14157), .dout(n14160));
    jdff dff_B_DZPrepAl3_1(.din(n14160), .dout(n14163));
    jdff dff_B_xkW8tMkH8_1(.din(n14163), .dout(n14166));
    jdff dff_B_ZkP7TBDr9_1(.din(n14166), .dout(n14169));
    jdff dff_B_LQ6f3UFc1_1(.din(n14169), .dout(n14172));
    jdff dff_B_odZ837622_1(.din(n14172), .dout(n14175));
    jdff dff_B_vzXoSk9X4_1(.din(n14175), .dout(n14178));
    jdff dff_B_adsMT2n22_1(.din(n820), .dout(n14181));
    jdff dff_A_k4xenT4h7_0(.din(n14186), .dout(n14183));
    jdff dff_A_a7we9Gva3_0(.din(n14189), .dout(n14186));
    jdff dff_A_I0ImGIF14_0(.din(n14192), .dout(n14189));
    jdff dff_A_13YisptX2_0(.din(n14195), .dout(n14192));
    jdff dff_A_I9Lt9Vzd6_0(.din(n14198), .dout(n14195));
    jdff dff_A_BTmGs1Yk9_0(.din(n14201), .dout(n14198));
    jdff dff_A_tPINrfYB9_0(.din(n14204), .dout(n14201));
    jdff dff_A_BPjLgJLX3_0(.din(n14207), .dout(n14204));
    jdff dff_A_ucfuI76z7_0(.din(n14210), .dout(n14207));
    jdff dff_A_dkBXmf8y8_0(.din(n14213), .dout(n14210));
    jdff dff_A_5HtJrMS99_0(.din(n14216), .dout(n14213));
    jdff dff_A_5zkDC9HT5_0(.din(n14219), .dout(n14216));
    jdff dff_A_YOSbSJAe4_0(.din(n14222), .dout(n14219));
    jdff dff_A_Aw2O2uyB6_0(.din(n14225), .dout(n14222));
    jdff dff_A_2eztFaSA8_0(.din(n14228), .dout(n14225));
    jdff dff_A_6D4g2EIK1_0(.din(n14231), .dout(n14228));
    jdff dff_A_wbKw1Hd12_0(.din(n14234), .dout(n14231));
    jdff dff_A_Z720XUCY7_0(.din(n14237), .dout(n14234));
    jdff dff_A_mzsbKJ0A0_0(.din(n624), .dout(n14237));
    jdff dff_A_mMzflZNv3_1(.din(n798), .dout(n14240));
    jdff dff_B_AdKknkAd7_1(.din(n649), .dout(n14244));
    jdff dff_B_Ym6Vbl3d6_1(.din(n14244), .dout(n14247));
    jdff dff_B_ATfipyHE7_1(.din(n14247), .dout(n14250));
    jdff dff_B_psPElH7X9_1(.din(n14250), .dout(n14253));
    jdff dff_B_o9LOOIpQ2_1(.din(n14253), .dout(n14256));
    jdff dff_B_57Rkjt1g2_1(.din(n14256), .dout(n14259));
    jdff dff_B_oYqScWT52_1(.din(n14259), .dout(n14262));
    jdff dff_B_lV0f9tA09_1(.din(n14262), .dout(n14265));
    jdff dff_B_hVxklnD74_1(.din(n14265), .dout(n14268));
    jdff dff_B_5jGr5oyl7_1(.din(n14268), .dout(n14271));
    jdff dff_B_Dcg3VGSg8_1(.din(n14271), .dout(n14274));
    jdff dff_B_ptQJVMAC3_1(.din(n14274), .dout(n14277));
    jdff dff_B_b6MtkQpX9_1(.din(n14277), .dout(n14280));
    jdff dff_B_rKwLbcEY2_1(.din(n14280), .dout(n14283));
    jdff dff_B_aBcORKe87_1(.din(n14283), .dout(n14286));
    jdff dff_B_e2lxoe595_1(.din(n634), .dout(n14289));
    jdff dff_A_0pDleJ5R5_0(.din(n14294), .dout(n14291));
    jdff dff_A_mHUCRWvC3_0(.din(n14297), .dout(n14294));
    jdff dff_A_KvTRu6M32_0(.din(n14300), .dout(n14297));
    jdff dff_A_NMlXlc5E6_0(.din(n14303), .dout(n14300));
    jdff dff_A_6Vq3yUtu1_0(.din(n14306), .dout(n14303));
    jdff dff_A_EnQjXoip4_0(.din(n14309), .dout(n14306));
    jdff dff_A_Lr4elQOt6_0(.din(n14312), .dout(n14309));
    jdff dff_A_8UBRyQ647_0(.din(n14315), .dout(n14312));
    jdff dff_A_JYv7GULW8_0(.din(n14318), .dout(n14315));
    jdff dff_A_GscKWzc12_0(.din(n14321), .dout(n14318));
    jdff dff_A_guE4PUy30_0(.din(n14324), .dout(n14321));
    jdff dff_A_Ju6eZYVy8_0(.din(n14327), .dout(n14324));
    jdff dff_A_R1jzM2gi9_0(.din(n14330), .dout(n14327));
    jdff dff_A_MElvZuSi2_0(.din(n14333), .dout(n14330));
    jdff dff_A_8MtG78A65_0(.din(n14336), .dout(n14333));
    jdff dff_A_O45etuQo1_0(.din(n465), .dout(n14336));
    jdff dff_A_w1J36y282_1(.din(n612), .dout(n14339));
    jdff dff_B_kMJdIi8X0_1(.din(n490), .dout(n14343));
    jdff dff_B_acniKS1l7_1(.din(n14343), .dout(n14346));
    jdff dff_B_sKMPpX0Y6_1(.din(n14346), .dout(n14349));
    jdff dff_B_lkREedsx8_1(.din(n14349), .dout(n14352));
    jdff dff_B_LuK1vCnM8_1(.din(n14352), .dout(n14355));
    jdff dff_B_7iCANmHr3_1(.din(n14355), .dout(n14358));
    jdff dff_B_5R1v7BSg4_1(.din(n14358), .dout(n14361));
    jdff dff_B_lIklxeFu5_1(.din(n14361), .dout(n14364));
    jdff dff_B_EMIjIBl47_1(.din(n14364), .dout(n14367));
    jdff dff_B_pRj0KyJu7_1(.din(n14367), .dout(n14370));
    jdff dff_B_Zyuwm4wT3_1(.din(n14370), .dout(n14373));
    jdff dff_B_223yyBnc1_1(.din(n14373), .dout(n14376));
    jdff dff_B_mivY9yYO3_1(.din(n475), .dout(n14379));
    jdff dff_A_YghuRqzn2_0(.din(n14384), .dout(n14381));
    jdff dff_A_mCe75unF2_0(.din(n14387), .dout(n14384));
    jdff dff_A_LLBwnret3_0(.din(n14390), .dout(n14387));
    jdff dff_A_A2uk5kT93_0(.din(n14393), .dout(n14390));
    jdff dff_A_GRq9yJjw4_0(.din(n14396), .dout(n14393));
    jdff dff_A_IbVR6JTN4_0(.din(n14399), .dout(n14396));
    jdff dff_A_Kcu7LNBs7_0(.din(n14402), .dout(n14399));
    jdff dff_A_rGT5YZ3j4_0(.din(n14405), .dout(n14402));
    jdff dff_A_ApxXQGR94_0(.din(n14408), .dout(n14405));
    jdff dff_A_V76GR7Iw8_0(.din(n14411), .dout(n14408));
    jdff dff_A_2TC2PRkm0_0(.din(n14414), .dout(n14411));
    jdff dff_A_ItZ3DfJD9_0(.din(n14417), .dout(n14414));
    jdff dff_A_vEHJDhK88_0(.din(n333), .dout(n14417));
    jdff dff_A_RjMD47tF9_1(.din(n453), .dout(n14420));
    jdff dff_B_uW5YyeLi5_1(.din(n358), .dout(n14424));
    jdff dff_B_F8HT6iDB7_1(.din(n14424), .dout(n14427));
    jdff dff_B_spgkFarl1_1(.din(n14427), .dout(n14430));
    jdff dff_B_Cl3PKAn14_1(.din(n14430), .dout(n14433));
    jdff dff_B_H0hHKyTQ3_1(.din(n14433), .dout(n14436));
    jdff dff_B_3NaMh7mf2_1(.din(n14436), .dout(n14439));
    jdff dff_B_8u50gTNV8_1(.din(n14439), .dout(n14442));
    jdff dff_B_U8ykEoTV5_1(.din(n14442), .dout(n14445));
    jdff dff_B_kHBgj2ct0_1(.din(n14445), .dout(n14448));
    jdff dff_B_gf04LRoR5_1(.din(n343), .dout(n14451));
    jdff dff_A_KFtXeObF6_0(.din(n14456), .dout(n14453));
    jdff dff_A_gDAG2uvu0_0(.din(n14459), .dout(n14456));
    jdff dff_A_l3fN9AQo9_0(.din(n14462), .dout(n14459));
    jdff dff_A_zmhu8g9k0_0(.din(n14465), .dout(n14462));
    jdff dff_A_DlyKsRMP4_0(.din(n14468), .dout(n14465));
    jdff dff_A_4nmWnb527_0(.din(n14471), .dout(n14468));
    jdff dff_A_valVlmqL2_0(.din(n14474), .dout(n14471));
    jdff dff_A_gF5BJC1H4_0(.din(n14477), .dout(n14474));
    jdff dff_A_CxuUWjyH7_0(.din(n14480), .dout(n14477));
    jdff dff_A_mRes1rl40_0(.din(n224), .dout(n14480));
    jdff dff_A_WxYnSB6O0_1(.din(n321), .dout(n14483));
    jdff dff_B_IuinFrhh4_1(.din(n249), .dout(n14487));
    jdff dff_B_BQSZpY1a8_1(.din(n14487), .dout(n14490));
    jdff dff_B_PdmuyN320_1(.din(n14490), .dout(n14493));
    jdff dff_B_W36D3cMK6_1(.din(n14493), .dout(n14496));
    jdff dff_B_NGmeOSA00_1(.din(n14496), .dout(n14499));
    jdff dff_B_Su360Bny1_1(.din(n14499), .dout(n14502));
    jdff dff_B_wzAgij7Z4_1(.din(n234), .dout(n14505));
    jdff dff_A_9U95j5xh3_0(.din(n14510), .dout(n14507));
    jdff dff_A_ZP3HyAxE7_0(.din(n14513), .dout(n14510));
    jdff dff_A_uiWKBazU3_0(.din(n14516), .dout(n14513));
    jdff dff_A_kFeW8RfP9_0(.din(n14519), .dout(n14516));
    jdff dff_A_KoVx2Kan5_0(.din(n14522), .dout(n14519));
    jdff dff_A_Ylz2tDqD9_0(.din(n14525), .dout(n14522));
    jdff dff_A_GHg8aXye0_0(.din(n148), .dout(n14525));
    jdff dff_A_GQBtAAG96_1(.din(n212), .dout(n14528));
    jdff dff_B_Uv9ReWOd9_1(.din(n170), .dout(n14532));
    jdff dff_B_NMrMQwpv2_1(.din(n14532), .dout(n14535));
    jdff dff_B_cXBzVoJC3_1(.din(n14535), .dout(n14538));
    jdff dff_B_bRNIW5P95_1(.din(n155), .dout(n14541));
    jdff dff_B_9Vf5Icva4_2(.din(n78), .dout(n14544));
    jdff dff_A_CH6f1AEo0_0(.din(n14549), .dout(n14546));
    jdff dff_A_BfS0jTiv1_0(.din(n14552), .dout(n14549));
    jdff dff_A_HwO8AQJo2_0(.din(n14555), .dout(n14552));
    jdff dff_A_eQtCUR2S4_0(.din(n107), .dout(n14555));
    jdff dff_B_QKLZD07U2_0(.din(n132), .dout(n14559));
    jdff dff_A_HWHyE6Iw3_0(.din(n14564), .dout(n14561));
    jdff dff_A_eAFIM9nI2_0(.din(n75), .dout(n14564));
    jdff dff_A_ezmFXke16_1(.din(n4046), .dout(n14567));
    jdff dff_B_ha1f2K3W5_1(.din(n3683), .dout(n14571));
    jdff dff_B_SVlH4JPV1_2(.din(n3290), .dout(n14574));
    jdff dff_B_1dCmcIVs7_2(.din(n14574), .dout(n14577));
    jdff dff_B_HXwN8Lw13_2(.din(n14577), .dout(n14580));
    jdff dff_B_z04SlnyX3_2(.din(n14580), .dout(n14583));
    jdff dff_B_Yq8ukHI04_2(.din(n14583), .dout(n14586));
    jdff dff_B_NmQc9hKf4_2(.din(n14586), .dout(n14589));
    jdff dff_B_XuNwJZp97_2(.din(n14589), .dout(n14592));
    jdff dff_B_fKhPNZ3o0_2(.din(n14592), .dout(n14595));
    jdff dff_B_13MhYITO2_2(.din(n14595), .dout(n14598));
    jdff dff_B_XFPRGYNU8_2(.din(n14598), .dout(n14601));
    jdff dff_B_buTV6WBg6_2(.din(n14601), .dout(n14604));
    jdff dff_B_UjuXZ5CJ3_2(.din(n14604), .dout(n14607));
    jdff dff_B_05ly3pzf6_2(.din(n14607), .dout(n14610));
    jdff dff_B_1BVgJJ1u8_2(.din(n14610), .dout(n14613));
    jdff dff_B_XLESq5Yo7_2(.din(n14613), .dout(n14616));
    jdff dff_B_bvomDQYL5_2(.din(n14616), .dout(n14619));
    jdff dff_B_q9w15ckF9_2(.din(n14619), .dout(n14622));
    jdff dff_B_hD4v8Ou89_2(.din(n14622), .dout(n14625));
    jdff dff_B_X7ecC6Wd5_2(.din(n14625), .dout(n14628));
    jdff dff_B_QafV0eiG5_2(.din(n14628), .dout(n14631));
    jdff dff_B_RrjQB6hy1_2(.din(n14631), .dout(n14634));
    jdff dff_B_NGJoTSCz3_2(.din(n14634), .dout(n14637));
    jdff dff_B_ayq64um91_2(.din(n14637), .dout(n14640));
    jdff dff_B_19hUALFP2_2(.din(n14640), .dout(n14643));
    jdff dff_B_MGeJWS6N6_2(.din(n14643), .dout(n14646));
    jdff dff_B_S4elgKpK0_2(.din(n14646), .dout(n14649));
    jdff dff_B_NUkd8ZMM3_2(.din(n14649), .dout(n14652));
    jdff dff_B_Pdm31MgI0_2(.din(n14652), .dout(n14655));
    jdff dff_B_ST9919Fo5_2(.din(n14655), .dout(n14658));
    jdff dff_B_rykJtCo34_2(.din(n14658), .dout(n14661));
    jdff dff_B_v9OHv9Jy7_2(.din(n14661), .dout(n14664));
    jdff dff_B_9UDA5jTH7_2(.din(n14664), .dout(n14667));
    jdff dff_B_o96nVqcz0_2(.din(n14667), .dout(n14670));
    jdff dff_B_dsntBdmM9_2(.din(n14670), .dout(n14673));
    jdff dff_B_PGcsK3oM3_2(.din(n14673), .dout(n14676));
    jdff dff_B_DW5CnjLJ6_2(.din(n14676), .dout(n14679));
    jdff dff_B_kPbPoVDA1_2(.din(n14679), .dout(n14682));
    jdff dff_B_U2tUafzD3_2(.din(n14682), .dout(n14685));
    jdff dff_B_eWjOhlCz6_2(.din(n14685), .dout(n14688));
    jdff dff_B_n3CbNZ7m1_2(.din(n14688), .dout(n14691));
    jdff dff_B_h19lBGnf6_2(.din(n14691), .dout(n14694));
    jdff dff_B_YmRQM7ho6_2(.din(n14694), .dout(n14697));
    jdff dff_B_5PjTactY9_2(.din(n14697), .dout(n14700));
    jdff dff_A_2JoOJDSK2_0(.din(n3660), .dout(n14702));
    jdff dff_B_dHhXXkpS5_1(.din(n3297), .dout(n14706));
    jdff dff_B_J4iVVmD45_2(.din(n2905), .dout(n14709));
    jdff dff_B_kRUpxviw3_2(.din(n14709), .dout(n14712));
    jdff dff_B_00tmrzpk5_2(.din(n14712), .dout(n14715));
    jdff dff_B_sX4AHlqn2_2(.din(n14715), .dout(n14718));
    jdff dff_B_XiFH1nWY4_2(.din(n14718), .dout(n14721));
    jdff dff_B_JjgOmFdZ7_2(.din(n14721), .dout(n14724));
    jdff dff_B_xCXM2NdE3_2(.din(n14724), .dout(n14727));
    jdff dff_B_tXtJZLsf3_2(.din(n14727), .dout(n14730));
    jdff dff_B_C68lsUKi6_2(.din(n14730), .dout(n14733));
    jdff dff_B_o8ytgLja9_2(.din(n14733), .dout(n14736));
    jdff dff_B_5maTWP3Q7_2(.din(n14736), .dout(n14739));
    jdff dff_B_EOLkSml62_2(.din(n14739), .dout(n14742));
    jdff dff_B_5J2p2Z6a5_2(.din(n14742), .dout(n14745));
    jdff dff_B_wiSXpisI5_2(.din(n14745), .dout(n14748));
    jdff dff_B_T20hXRdQ5_2(.din(n14748), .dout(n14751));
    jdff dff_B_hyFsdzvO5_2(.din(n14751), .dout(n14754));
    jdff dff_B_ZHpLUpvA3_2(.din(n14754), .dout(n14757));
    jdff dff_B_C6MODavM5_2(.din(n14757), .dout(n14760));
    jdff dff_B_Q4GKMZ6Q8_2(.din(n14760), .dout(n14763));
    jdff dff_B_yBBfHVMM8_2(.din(n14763), .dout(n14766));
    jdff dff_B_6rFDfqKX0_2(.din(n14766), .dout(n14769));
    jdff dff_B_rYoQMKwM4_2(.din(n14769), .dout(n14772));
    jdff dff_B_mC83W5Rc5_2(.din(n14772), .dout(n14775));
    jdff dff_B_uJtnMJem2_2(.din(n14775), .dout(n14778));
    jdff dff_B_QKsNVTjd3_2(.din(n14778), .dout(n14781));
    jdff dff_B_oqvn98nS2_2(.din(n14781), .dout(n14784));
    jdff dff_B_7BcMa4337_2(.din(n14784), .dout(n14787));
    jdff dff_B_8hs0nVhs3_2(.din(n14787), .dout(n14790));
    jdff dff_B_Vc8OozMm0_2(.din(n14790), .dout(n14793));
    jdff dff_B_PYBsMJ9P9_2(.din(n14793), .dout(n14796));
    jdff dff_B_xMXPbBb82_2(.din(n14796), .dout(n14799));
    jdff dff_B_p2nWBI8F7_2(.din(n14799), .dout(n14802));
    jdff dff_B_ddwJvNLP0_2(.din(n14802), .dout(n14805));
    jdff dff_B_KjfHu9ii9_2(.din(n14805), .dout(n14808));
    jdff dff_B_0AxgoCU34_2(.din(n14808), .dout(n14811));
    jdff dff_B_FGlZw0UB6_2(.din(n14811), .dout(n14814));
    jdff dff_B_apCgWL839_2(.din(n14814), .dout(n14817));
    jdff dff_B_AgWRX1l88_2(.din(n14817), .dout(n14820));
    jdff dff_B_WQwPjHer9_2(.din(n14820), .dout(n14823));
    jdff dff_B_hfAiVJWe3_2(.din(n14823), .dout(n14826));
    jdff dff_A_5cOfMQR71_1(.din(n3255), .dout(n14828));
    jdff dff_B_RNAk0Tkx4_1(.din(n2928), .dout(n14832));
    jdff dff_B_PhiVPLAi5_1(.din(n14832), .dout(n14835));
    jdff dff_B_InFZxYzN7_1(.din(n14835), .dout(n14838));
    jdff dff_B_oBaMsv0G5_1(.din(n14838), .dout(n14841));
    jdff dff_B_jMryvljm0_1(.din(n14841), .dout(n14844));
    jdff dff_B_jMceVpjg0_1(.din(n14844), .dout(n14847));
    jdff dff_B_heRGCE8B9_1(.din(n14847), .dout(n14850));
    jdff dff_B_GaBfpLVx4_1(.din(n14850), .dout(n14853));
    jdff dff_B_9uO6NMfn0_1(.din(n14853), .dout(n14856));
    jdff dff_B_x3ieAqcX2_1(.din(n14856), .dout(n14859));
    jdff dff_B_7IiFwS3P8_1(.din(n14859), .dout(n14862));
    jdff dff_B_MMbV8bfs2_1(.din(n14862), .dout(n14865));
    jdff dff_B_EwlDGIH42_1(.din(n14865), .dout(n14868));
    jdff dff_B_cdFzpImB1_1(.din(n14868), .dout(n14871));
    jdff dff_B_dl5NeYNR9_1(.din(n14871), .dout(n14874));
    jdff dff_B_5vqpXoGX5_1(.din(n14874), .dout(n14877));
    jdff dff_B_ZjGfVioi1_1(.din(n14877), .dout(n14880));
    jdff dff_B_0q1L5jKI0_1(.din(n14880), .dout(n14883));
    jdff dff_B_G80Po5kR9_1(.din(n14883), .dout(n14886));
    jdff dff_B_huyKn8U95_1(.din(n14886), .dout(n14889));
    jdff dff_B_VSsqfEtz9_1(.din(n14889), .dout(n14892));
    jdff dff_B_fHp5JBK31_1(.din(n14892), .dout(n14895));
    jdff dff_B_Y50gPpK19_1(.din(n14895), .dout(n14898));
    jdff dff_B_3ivmdiVg8_1(.din(n14898), .dout(n14901));
    jdff dff_B_iX1uKm0m5_1(.din(n14901), .dout(n14904));
    jdff dff_B_SyEwpmjE0_1(.din(n14904), .dout(n14907));
    jdff dff_B_lZFbIdAi7_1(.din(n14907), .dout(n14910));
    jdff dff_B_p6NBbtwH1_1(.din(n14910), .dout(n14913));
    jdff dff_B_yEzUR16l3_1(.din(n14913), .dout(n14916));
    jdff dff_B_BVIuilGA2_1(.din(n14916), .dout(n14919));
    jdff dff_B_9Dp1CswD9_1(.din(n14919), .dout(n14922));
    jdff dff_B_0UZTnRyO1_1(.din(n14922), .dout(n14925));
    jdff dff_B_mGM3q0Vz8_1(.din(n14925), .dout(n14928));
    jdff dff_B_KUOq6v4B6_1(.din(n14928), .dout(n14931));
    jdff dff_B_Ga6U3ZaT1_1(.din(n14931), .dout(n14934));
    jdff dff_B_i87Plare9_1(.din(n14934), .dout(n14937));
    jdff dff_B_Z8LzQloI7_1(.din(n2909), .dout(n14940));
    jdff dff_A_nvzMUPSq9_0(.din(n14945), .dout(n14942));
    jdff dff_A_mFVKxGu34_0(.din(n14948), .dout(n14945));
    jdff dff_A_irLXAV5G9_0(.din(n14951), .dout(n14948));
    jdff dff_A_RyDPdlYE3_0(.din(n14954), .dout(n14951));
    jdff dff_A_cE9ToscC4_0(.din(n14957), .dout(n14954));
    jdff dff_A_E4D3sfKA6_0(.din(n14960), .dout(n14957));
    jdff dff_A_Jk9NLDmv1_0(.din(n14963), .dout(n14960));
    jdff dff_A_MX7Ewhas0_0(.din(n14966), .dout(n14963));
    jdff dff_A_B8nYgEY25_0(.din(n14969), .dout(n14966));
    jdff dff_A_eZzfNJOH7_0(.din(n14972), .dout(n14969));
    jdff dff_A_UsNuXq1X7_0(.din(n14975), .dout(n14972));
    jdff dff_A_MXIAfFn31_0(.din(n14978), .dout(n14975));
    jdff dff_A_yO15gPJr5_0(.din(n14981), .dout(n14978));
    jdff dff_A_vP0gkV1y6_0(.din(n14984), .dout(n14981));
    jdff dff_A_kdFHnUVh3_0(.din(n14987), .dout(n14984));
    jdff dff_A_Lm5Gs0yh8_0(.din(n14990), .dout(n14987));
    jdff dff_A_TOM3HrQ90_0(.din(n14993), .dout(n14990));
    jdff dff_A_dViOtFSk2_0(.din(n14996), .dout(n14993));
    jdff dff_A_AZWB3P7r5_0(.din(n14999), .dout(n14996));
    jdff dff_A_60ukqH3e5_0(.din(n15002), .dout(n14999));
    jdff dff_A_k9uGuW0y1_0(.din(n15005), .dout(n15002));
    jdff dff_A_aJjaHec75_0(.din(n15008), .dout(n15005));
    jdff dff_A_DnOZtxGb6_0(.din(n15011), .dout(n15008));
    jdff dff_A_KYdOX3r87_0(.din(n15014), .dout(n15011));
    jdff dff_A_h8Kp11Vq8_0(.din(n15017), .dout(n15014));
    jdff dff_A_Bt6sxac45_0(.din(n15020), .dout(n15017));
    jdff dff_A_BPXW0qTw3_0(.din(n15023), .dout(n15020));
    jdff dff_A_t55fvk2X7_0(.din(n15026), .dout(n15023));
    jdff dff_A_MaHfv1FW1_0(.din(n15029), .dout(n15026));
    jdff dff_A_Y7GbduvZ9_0(.din(n15032), .dout(n15029));
    jdff dff_A_14xhSJk46_0(.din(n15035), .dout(n15032));
    jdff dff_A_ImEE9lU15_0(.din(n15038), .dout(n15035));
    jdff dff_A_iLKi4kvh6_0(.din(n15041), .dout(n15038));
    jdff dff_A_9KENl70F9_0(.din(n15044), .dout(n15041));
    jdff dff_A_4Rx08WPt0_0(.din(n15047), .dout(n15044));
    jdff dff_A_RF7ZFcvi5_0(.din(n15050), .dout(n15047));
    jdff dff_A_4Ww2YHwk1_0(.din(n2527), .dout(n15050));
    jdff dff_A_CozEEMQj4_0(.din(n2860), .dout(n15053));
    jdff dff_B_BOjcivN93_1(.din(n2534), .dout(n15057));
    jdff dff_A_BxerMc0E2_0(.din(n15062), .dout(n15059));
    jdff dff_A_cimKIYuX4_0(.din(n15065), .dout(n15062));
    jdff dff_A_WayADUjb1_0(.din(n15068), .dout(n15065));
    jdff dff_A_KuDZC9I02_0(.din(n15071), .dout(n15068));
    jdff dff_A_08M9oir51_0(.din(n15074), .dout(n15071));
    jdff dff_A_tL04Z9ZC3_0(.din(n15077), .dout(n15074));
    jdff dff_A_lQBRQG533_0(.din(n15080), .dout(n15077));
    jdff dff_A_yc2Ulbxy7_0(.din(n15083), .dout(n15080));
    jdff dff_A_WALWMKSr5_0(.din(n15086), .dout(n15083));
    jdff dff_A_kTz6nelh8_0(.din(n15089), .dout(n15086));
    jdff dff_A_CBnURHp55_0(.din(n15092), .dout(n15089));
    jdff dff_A_FbDy6Hqa8_0(.din(n15095), .dout(n15092));
    jdff dff_A_wE4lDe5G2_0(.din(n15098), .dout(n15095));
    jdff dff_A_6gPJGe730_0(.din(n15101), .dout(n15098));
    jdff dff_A_VhV8I7eJ5_0(.din(n15104), .dout(n15101));
    jdff dff_A_gzDa1RYH1_0(.din(n15107), .dout(n15104));
    jdff dff_A_nwetkaC47_0(.din(n15110), .dout(n15107));
    jdff dff_A_9EQNKs7y2_0(.din(n15113), .dout(n15110));
    jdff dff_A_0n1Cb1087_0(.din(n15116), .dout(n15113));
    jdff dff_A_0CZJAKpG5_0(.din(n15119), .dout(n15116));
    jdff dff_A_X2SkhwMt9_0(.din(n15122), .dout(n15119));
    jdff dff_A_F5OZ1ssi3_0(.din(n15125), .dout(n15122));
    jdff dff_A_f3oK9d4V5_0(.din(n15128), .dout(n15125));
    jdff dff_A_lOdRId168_0(.din(n15131), .dout(n15128));
    jdff dff_A_SyaBC5oX3_0(.din(n15134), .dout(n15131));
    jdff dff_A_PNUyjw2S6_0(.din(n15137), .dout(n15134));
    jdff dff_A_VHH0K7Fk1_0(.din(n15140), .dout(n15137));
    jdff dff_A_I0vO1TjO2_0(.din(n15143), .dout(n15140));
    jdff dff_A_QcxV2Gco2_0(.din(n15146), .dout(n15143));
    jdff dff_A_Uz29G7AQ7_0(.din(n15149), .dout(n15146));
    jdff dff_A_AALeN3uJ1_0(.din(n15152), .dout(n15149));
    jdff dff_A_VUxJTziZ8_0(.din(n15155), .dout(n15152));
    jdff dff_A_8AzY1BgI9_0(.din(n15158), .dout(n15155));
    jdff dff_A_z3WtrQqV4_0(.din(n2176), .dout(n15158));
    jdff dff_A_UaJP31Zr4_0(.din(n2482), .dout(n15161));
    jdff dff_B_L54OtKa01_1(.din(n2183), .dout(n15165));
    jdff dff_A_j5LpYyAI9_0(.din(n15170), .dout(n15167));
    jdff dff_A_4GuMcs7N8_0(.din(n15173), .dout(n15170));
    jdff dff_A_p0kP9c4r6_0(.din(n15176), .dout(n15173));
    jdff dff_A_za4cIv037_0(.din(n15179), .dout(n15176));
    jdff dff_A_wAJFscVw8_0(.din(n15182), .dout(n15179));
    jdff dff_A_b7g7ZcYN2_0(.din(n15185), .dout(n15182));
    jdff dff_A_z2ZGlGEA4_0(.din(n15188), .dout(n15185));
    jdff dff_A_umsH6zCL8_0(.din(n15191), .dout(n15188));
    jdff dff_A_JLlDFbRd2_0(.din(n15194), .dout(n15191));
    jdff dff_A_x5KzGJFz5_0(.din(n15197), .dout(n15194));
    jdff dff_A_NdGpRJNo7_0(.din(n15200), .dout(n15197));
    jdff dff_A_MvVhzOVP0_0(.din(n15203), .dout(n15200));
    jdff dff_A_mh6JhjAo7_0(.din(n15206), .dout(n15203));
    jdff dff_A_7hFL9iPU2_0(.din(n15209), .dout(n15206));
    jdff dff_A_zEVAQUr66_0(.din(n15212), .dout(n15209));
    jdff dff_A_SnifY13u4_0(.din(n15215), .dout(n15212));
    jdff dff_A_k3fn1NIj1_0(.din(n15218), .dout(n15215));
    jdff dff_A_6zqEzYZu6_0(.din(n15221), .dout(n15218));
    jdff dff_A_7XWCDsIC5_0(.din(n15224), .dout(n15221));
    jdff dff_A_fNutgw799_0(.din(n15227), .dout(n15224));
    jdff dff_A_rUtuXh2z2_0(.din(n15230), .dout(n15227));
    jdff dff_A_X6Mg3W7K6_0(.din(n15233), .dout(n15230));
    jdff dff_A_WuETERNJ9_0(.din(n15236), .dout(n15233));
    jdff dff_A_m8Rt0BIM9_0(.din(n15239), .dout(n15236));
    jdff dff_A_ZhwonHSi7_0(.din(n15242), .dout(n15239));
    jdff dff_A_CULjJBlH4_0(.din(n15245), .dout(n15242));
    jdff dff_A_TdxwIVvD1_0(.din(n15248), .dout(n15245));
    jdff dff_A_HfS7QI0y6_0(.din(n15251), .dout(n15248));
    jdff dff_A_bim36IMe0_0(.din(n15254), .dout(n15251));
    jdff dff_A_PDCWZ8WG3_0(.din(n15257), .dout(n15254));
    jdff dff_A_fuaXEbQU2_0(.din(n1852), .dout(n15257));
    jdff dff_A_tK0LOVYt9_0(.din(n2131), .dout(n15260));
    jdff dff_B_25LyZmhv8_1(.din(n1859), .dout(n15264));
    jdff dff_A_1DTD4n8o4_0(.din(n15269), .dout(n15266));
    jdff dff_A_27Vjn8E55_0(.din(n15272), .dout(n15269));
    jdff dff_A_BliCZHBw1_0(.din(n15275), .dout(n15272));
    jdff dff_A_fXjxcnL24_0(.din(n15278), .dout(n15275));
    jdff dff_A_HOjB8P6M0_0(.din(n15281), .dout(n15278));
    jdff dff_A_1EmnySFl3_0(.din(n15284), .dout(n15281));
    jdff dff_A_FuMXZAhx2_0(.din(n15287), .dout(n15284));
    jdff dff_A_UxwMdAWx5_0(.din(n15290), .dout(n15287));
    jdff dff_A_pWCk4pl57_0(.din(n15293), .dout(n15290));
    jdff dff_A_VAfjNRrt7_0(.din(n15296), .dout(n15293));
    jdff dff_A_fOvk9cU14_0(.din(n15299), .dout(n15296));
    jdff dff_A_wAk2BdGn2_0(.din(n15302), .dout(n15299));
    jdff dff_A_Zz4QNO8u9_0(.din(n15305), .dout(n15302));
    jdff dff_A_kqjg2sC43_0(.din(n15308), .dout(n15305));
    jdff dff_A_bHnznFdG8_0(.din(n15311), .dout(n15308));
    jdff dff_A_aVJMZtkD3_0(.din(n15314), .dout(n15311));
    jdff dff_A_TliCd5nd7_0(.din(n15317), .dout(n15314));
    jdff dff_A_vgzIR9E05_0(.din(n15320), .dout(n15317));
    jdff dff_A_86JmCiBZ5_0(.din(n15323), .dout(n15320));
    jdff dff_A_z9Z0vJC13_0(.din(n15326), .dout(n15323));
    jdff dff_A_bVLbzTMZ9_0(.din(n15329), .dout(n15326));
    jdff dff_A_OanEgcdL1_0(.din(n15332), .dout(n15329));
    jdff dff_A_ZQtBZvJU8_0(.din(n15335), .dout(n15332));
    jdff dff_A_qfSXjFBA6_0(.din(n15338), .dout(n15335));
    jdff dff_A_L6IHRjm13_0(.din(n15341), .dout(n15338));
    jdff dff_A_4Wo6oDnA2_0(.din(n15344), .dout(n15341));
    jdff dff_A_CqY9cvf81_0(.din(n15347), .dout(n15344));
    jdff dff_A_ufPHR4DL3_0(.din(n1555), .dout(n15347));
    jdff dff_A_ZUZuYvs31_0(.din(n1807), .dout(n15350));
    jdff dff_B_n8ulN2hL2_1(.din(n1562), .dout(n15354));
    jdff dff_A_xjivaEHV1_0(.din(n15359), .dout(n15356));
    jdff dff_A_ZvFdidse1_0(.din(n15362), .dout(n15359));
    jdff dff_A_xFCNRFwu0_0(.din(n15365), .dout(n15362));
    jdff dff_A_Kua27kwP5_0(.din(n15368), .dout(n15365));
    jdff dff_A_1FeNvmBt3_0(.din(n15371), .dout(n15368));
    jdff dff_A_IxzFZAqA6_0(.din(n15374), .dout(n15371));
    jdff dff_A_2qGJEOFE4_0(.din(n15377), .dout(n15374));
    jdff dff_A_kaogT0kH7_0(.din(n15380), .dout(n15377));
    jdff dff_A_bKpgsxEn1_0(.din(n15383), .dout(n15380));
    jdff dff_A_NZwXKZmx8_0(.din(n15386), .dout(n15383));
    jdff dff_A_KHPVtjxh0_0(.din(n15389), .dout(n15386));
    jdff dff_A_xrEJUqYf1_0(.din(n15392), .dout(n15389));
    jdff dff_A_jY8NaeET5_0(.din(n15395), .dout(n15392));
    jdff dff_A_POqxp1OC9_0(.din(n15398), .dout(n15395));
    jdff dff_A_cgWZzR0d5_0(.din(n15401), .dout(n15398));
    jdff dff_A_e5NLw3368_0(.din(n15404), .dout(n15401));
    jdff dff_A_L0BiFdBL6_0(.din(n15407), .dout(n15404));
    jdff dff_A_iW3Ri9iE7_0(.din(n15410), .dout(n15407));
    jdff dff_A_xoUAkCg02_0(.din(n15413), .dout(n15410));
    jdff dff_A_K3HezAHJ7_0(.din(n15416), .dout(n15413));
    jdff dff_A_HGeg1hHW6_0(.din(n15419), .dout(n15416));
    jdff dff_A_gL9w6xVe1_0(.din(n15422), .dout(n15419));
    jdff dff_A_w2bfYK5X3_0(.din(n15425), .dout(n15422));
    jdff dff_A_rkplaC5G5_0(.din(n15428), .dout(n15425));
    jdff dff_A_9rwQQ0ko5_0(.din(n1285), .dout(n15428));
    jdff dff_A_WZktrhNT6_0(.din(n1510), .dout(n15431));
    jdff dff_B_XzZDx8md5_1(.din(n1292), .dout(n15435));
    jdff dff_A_S8SNoUsr9_0(.din(n15440), .dout(n15437));
    jdff dff_A_wpuGUwG39_0(.din(n15443), .dout(n15440));
    jdff dff_A_FvzflmIP5_0(.din(n15446), .dout(n15443));
    jdff dff_A_X1Fed3WN2_0(.din(n15449), .dout(n15446));
    jdff dff_A_4EEzFBoY1_0(.din(n15452), .dout(n15449));
    jdff dff_A_4guQfGBD0_0(.din(n15455), .dout(n15452));
    jdff dff_A_wS0E1z5y9_0(.din(n15458), .dout(n15455));
    jdff dff_A_YrXEYsNd4_0(.din(n15461), .dout(n15458));
    jdff dff_A_OjWPk9ni2_0(.din(n15464), .dout(n15461));
    jdff dff_A_YignJEAz3_0(.din(n15467), .dout(n15464));
    jdff dff_A_UPRj53l43_0(.din(n15470), .dout(n15467));
    jdff dff_A_RHGOpSsd7_0(.din(n15473), .dout(n15470));
    jdff dff_A_4aoOijak7_0(.din(n15476), .dout(n15473));
    jdff dff_A_6Ja7ZXuS3_0(.din(n15479), .dout(n15476));
    jdff dff_A_pWKTwEMx6_0(.din(n15482), .dout(n15479));
    jdff dff_A_7gdt2f474_0(.din(n15485), .dout(n15482));
    jdff dff_A_4U1aKAbU6_0(.din(n15488), .dout(n15485));
    jdff dff_A_28mJBR7X3_0(.din(n15491), .dout(n15488));
    jdff dff_A_0vlo5Euv3_0(.din(n15494), .dout(n15491));
    jdff dff_A_b3Uh1PC65_0(.din(n15497), .dout(n15494));
    jdff dff_A_GzMRwxlk0_0(.din(n15500), .dout(n15497));
    jdff dff_A_Y1PZdxHC4_0(.din(n1045), .dout(n15500));
    jdff dff_A_pUfXEeqD8_0(.din(n1240), .dout(n15503));
    jdff dff_B_qxEaHlTH9_1(.din(n1052), .dout(n15507));
    jdff dff_A_TgP2QZxM9_0(.din(n15512), .dout(n15509));
    jdff dff_A_0OEhDnkf8_0(.din(n15515), .dout(n15512));
    jdff dff_A_OZmavzp60_0(.din(n15518), .dout(n15515));
    jdff dff_A_dUy6AJW28_0(.din(n15521), .dout(n15518));
    jdff dff_A_eGm3zfLS4_0(.din(n15524), .dout(n15521));
    jdff dff_A_Z04TkIfy3_0(.din(n15527), .dout(n15524));
    jdff dff_A_we4WEDFt3_0(.din(n15530), .dout(n15527));
    jdff dff_A_KjXsNrp10_0(.din(n15533), .dout(n15530));
    jdff dff_A_rjJE9DLc2_0(.din(n15536), .dout(n15533));
    jdff dff_A_glNc0pJw3_0(.din(n15539), .dout(n15536));
    jdff dff_A_BEOL1gef2_0(.din(n15542), .dout(n15539));
    jdff dff_A_617rBd9v6_0(.din(n15545), .dout(n15542));
    jdff dff_A_gUGhPz4P7_0(.din(n15548), .dout(n15545));
    jdff dff_A_SIE3Puh01_0(.din(n15551), .dout(n15548));
    jdff dff_A_DuFthvhz9_0(.din(n15554), .dout(n15551));
    jdff dff_A_byQnZsMu2_0(.din(n15557), .dout(n15554));
    jdff dff_A_ggmsijOl8_0(.din(n15560), .dout(n15557));
    jdff dff_A_HEERYzqX3_0(.din(n15563), .dout(n15560));
    jdff dff_A_07ryFYOn6_0(.din(n832), .dout(n15563));
    jdff dff_A_9FZh6byn6_0(.din(n1000), .dout(n15566));
    jdff dff_B_r4hNDjzn8_1(.din(n839), .dout(n15570));
    jdff dff_A_I8DUMGoX0_0(.din(n15575), .dout(n15572));
    jdff dff_A_Lq53wyEv9_0(.din(n15578), .dout(n15575));
    jdff dff_A_ZDDJNgU28_0(.din(n15581), .dout(n15578));
    jdff dff_A_lIx0bLKJ0_0(.din(n15584), .dout(n15581));
    jdff dff_A_MfRrB5g66_0(.din(n15587), .dout(n15584));
    jdff dff_A_Y63wSNTp3_0(.din(n15590), .dout(n15587));
    jdff dff_A_iwE2BmLL0_0(.din(n15593), .dout(n15590));
    jdff dff_A_I1qV6Jaa1_0(.din(n15596), .dout(n15593));
    jdff dff_A_yRNag3fp1_0(.din(n15599), .dout(n15596));
    jdff dff_A_RlUYuPSY5_0(.din(n15602), .dout(n15599));
    jdff dff_A_rAoiwxM79_0(.din(n15605), .dout(n15602));
    jdff dff_A_k0fiZLEa3_0(.din(n15608), .dout(n15605));
    jdff dff_A_aFVBh2xO5_0(.din(n15611), .dout(n15608));
    jdff dff_A_9jfXyD3y3_0(.din(n15614), .dout(n15611));
    jdff dff_A_U1tuxpQ13_0(.din(n15617), .dout(n15614));
    jdff dff_A_ZGD17F2e9_0(.din(n646), .dout(n15617));
    jdff dff_A_nhN25l222_0(.din(n787), .dout(n15620));
    jdff dff_B_3vhxBByS6_1(.din(n653), .dout(n15624));
    jdff dff_A_Ps0Tcvho8_0(.din(n15629), .dout(n15626));
    jdff dff_A_25z5P6Bh1_0(.din(n15632), .dout(n15629));
    jdff dff_A_WkQvTt551_0(.din(n15635), .dout(n15632));
    jdff dff_A_npWI4njK8_0(.din(n15638), .dout(n15635));
    jdff dff_A_YRLimjjR8_0(.din(n15641), .dout(n15638));
    jdff dff_A_jBdQNVfI9_0(.din(n15644), .dout(n15641));
    jdff dff_A_7PdzuaE90_0(.din(n15647), .dout(n15644));
    jdff dff_A_nA7dc5BY9_0(.din(n15650), .dout(n15647));
    jdff dff_A_jhRbLA6Q7_0(.din(n15653), .dout(n15650));
    jdff dff_A_4EuBYuut9_0(.din(n15656), .dout(n15653));
    jdff dff_A_yhwUhhM33_0(.din(n15659), .dout(n15656));
    jdff dff_A_m062pSjM0_0(.din(n15662), .dout(n15659));
    jdff dff_A_Usx6TU591_0(.din(n487), .dout(n15662));
    jdff dff_A_xTHqHmzl2_0(.din(n601), .dout(n15665));
    jdff dff_B_HfKmuf415_1(.din(n494), .dout(n15669));
    jdff dff_A_0qNLck1J0_0(.din(n15674), .dout(n15671));
    jdff dff_A_17ZMACWF0_0(.din(n15677), .dout(n15674));
    jdff dff_A_Gc39vKPx9_0(.din(n15680), .dout(n15677));
    jdff dff_A_RtNC1uB15_0(.din(n15683), .dout(n15680));
    jdff dff_A_PV9EYaJr3_0(.din(n15686), .dout(n15683));
    jdff dff_A_OMyJ6xQq8_0(.din(n15689), .dout(n15686));
    jdff dff_A_UFZvJpGt8_0(.din(n15692), .dout(n15689));
    jdff dff_A_E2NoMfwW0_0(.din(n15695), .dout(n15692));
    jdff dff_A_jALWbNxy6_0(.din(n15698), .dout(n15695));
    jdff dff_A_Ub9v0iXs2_0(.din(n355), .dout(n15698));
    jdff dff_A_uGHgRN7S4_0(.din(n442), .dout(n15701));
    jdff dff_B_BZ4iv02w0_1(.din(n362), .dout(n15705));
    jdff dff_A_DMVcyFUf3_0(.din(n15710), .dout(n15707));
    jdff dff_A_mIiBCANF5_0(.din(n15713), .dout(n15710));
    jdff dff_A_oJ5GVM8I1_0(.din(n15716), .dout(n15713));
    jdff dff_A_lfYOIB5d5_0(.din(n15719), .dout(n15716));
    jdff dff_A_3gPfbbnv4_0(.din(n15722), .dout(n15719));
    jdff dff_A_kYqYKoxr2_0(.din(n15725), .dout(n15722));
    jdff dff_A_yz2g5o3T1_0(.din(n246), .dout(n15725));
    jdff dff_A_OcGInJTO8_0(.din(n310), .dout(n15728));
    jdff dff_B_lka824er8_1(.din(n253), .dout(n15732));
    jdff dff_A_ZdyDGYRF6_0(.din(n15737), .dout(n15734));
    jdff dff_A_7RScKASn6_0(.din(n15740), .dout(n15737));
    jdff dff_A_G0LNzcrn8_0(.din(n15743), .dout(n15740));
    jdff dff_A_wyHhALjm2_0(.din(n167), .dout(n15743));
    jdff dff_B_AsRBWcbj0_0(.din(n200), .dout(n15747));
    jdff dff_A_iGsqUyTS8_0(.din(n124), .dout(n15749));
    jdff dff_A_kHDRHVTJ0_0(.din(n15756), .dout(n15752));
    jdff dff_B_cMjIhJEV7_2(.din(n4087), .dout(n15756));
    jdff dff_B_sWP56mRH1_2(.din(n3699), .dout(n15759));
    jdff dff_B_z2gJh9B52_2(.din(n15759), .dout(n15762));
    jdff dff_B_s9MKeXFT0_2(.din(n15762), .dout(n15765));
    jdff dff_B_BlJtStrS9_2(.din(n15765), .dout(n15768));
    jdff dff_B_4ZrApfOc7_2(.din(n15768), .dout(n15771));
    jdff dff_B_8WTIScRC8_2(.din(n15771), .dout(n15774));
    jdff dff_B_aaE8ibXH6_2(.din(n15774), .dout(n15777));
    jdff dff_B_p8XQ9mHl2_2(.din(n15777), .dout(n15780));
    jdff dff_B_rsoZITgZ2_2(.din(n15780), .dout(n15783));
    jdff dff_B_jskZ009W2_2(.din(n15783), .dout(n15786));
    jdff dff_B_xaX5NC4Z6_2(.din(n15786), .dout(n15789));
    jdff dff_B_zVOHL91y4_2(.din(n15789), .dout(n15792));
    jdff dff_B_AoneoiBe9_2(.din(n15792), .dout(n15795));
    jdff dff_B_oa4YAf3i9_2(.din(n15795), .dout(n15798));
    jdff dff_B_JsRxpWHk4_2(.din(n15798), .dout(n15801));
    jdff dff_B_V75BtALJ3_2(.din(n15801), .dout(n15804));
    jdff dff_B_wMJb6RMj2_2(.din(n15804), .dout(n15807));
    jdff dff_B_C2abLtti9_2(.din(n15807), .dout(n15810));
    jdff dff_B_aiyDfmbh1_2(.din(n15810), .dout(n15813));
    jdff dff_B_kFzdtis48_2(.din(n15813), .dout(n15816));
    jdff dff_B_9puinoJx4_2(.din(n15816), .dout(n15819));
    jdff dff_B_PJWfu2Pf8_2(.din(n15819), .dout(n15822));
    jdff dff_B_DYGmZ1rB0_2(.din(n15822), .dout(n15825));
    jdff dff_B_9ImUXCEc7_2(.din(n15825), .dout(n15828));
    jdff dff_B_AqnN7G0m1_2(.din(n15828), .dout(n15831));
    jdff dff_B_AGVbdhUS4_2(.din(n15831), .dout(n15834));
    jdff dff_B_ItjhBvyb7_2(.din(n15834), .dout(n15837));
    jdff dff_B_q11eEC790_2(.din(n15837), .dout(n15840));
    jdff dff_B_GlJLWQMp1_2(.din(n15840), .dout(n15843));
    jdff dff_B_w76aUxrT4_2(.din(n15843), .dout(n15846));
    jdff dff_B_0gDijboI2_2(.din(n15846), .dout(n15849));
    jdff dff_B_jGYKGauk4_2(.din(n15849), .dout(n15852));
    jdff dff_B_rLjNOMb91_2(.din(n15852), .dout(n15855));
    jdff dff_B_zAdSHiSq5_2(.din(n15855), .dout(n15858));
    jdff dff_B_2emaucSo3_2(.din(n15858), .dout(n15861));
    jdff dff_B_Eevua5uk6_2(.din(n15861), .dout(n15864));
    jdff dff_B_shMmYz582_2(.din(n15864), .dout(n15867));
    jdff dff_B_NZ4Gurnf1_2(.din(n15867), .dout(n15870));
    jdff dff_B_htANaIDt2_2(.din(n15870), .dout(n15873));
    jdff dff_B_lJ5FMkbB7_2(.din(n15873), .dout(n15876));
    jdff dff_B_F9pzeo6i8_2(.din(n15876), .dout(n15879));
    jdff dff_B_eu71PbNQ2_2(.din(n15879), .dout(n15882));
    jdff dff_B_SYqhYXJy0_2(.din(n15882), .dout(n15885));
    jdff dff_A_pjjutMCB9_0(.din(n3714), .dout(n15887));
    jdff dff_B_YGBk4d6B0_1(.din(n3706), .dout(n15891));
    jdff dff_B_DNzvvfS67_2(.din(n3309), .dout(n15894));
    jdff dff_B_9PEsjT5o3_2(.din(n15894), .dout(n15897));
    jdff dff_B_F9IZMHeN6_2(.din(n15897), .dout(n15900));
    jdff dff_B_n4xbpcwy0_2(.din(n15900), .dout(n15903));
    jdff dff_B_TX0PA1M27_2(.din(n15903), .dout(n15906));
    jdff dff_B_s0ldgvR69_2(.din(n15906), .dout(n15909));
    jdff dff_B_ufuef6bT3_2(.din(n15909), .dout(n15912));
    jdff dff_B_AWDttdoo6_2(.din(n15912), .dout(n15915));
    jdff dff_B_46xmwMo04_2(.din(n15915), .dout(n15918));
    jdff dff_B_DdNHP23u2_2(.din(n15918), .dout(n15921));
    jdff dff_B_3si6Bylu5_2(.din(n15921), .dout(n15924));
    jdff dff_B_6md3Pfvk6_2(.din(n15924), .dout(n15927));
    jdff dff_B_zMoJKukp6_2(.din(n15927), .dout(n15930));
    jdff dff_B_T7pmnkJE6_2(.din(n15930), .dout(n15933));
    jdff dff_B_pJFDvR551_2(.din(n15933), .dout(n15936));
    jdff dff_B_XdTbbgsw2_2(.din(n15936), .dout(n15939));
    jdff dff_B_3GcBCU8N6_2(.din(n15939), .dout(n15942));
    jdff dff_B_ONcR3NhH2_2(.din(n15942), .dout(n15945));
    jdff dff_B_mKjN1i3f4_2(.din(n15945), .dout(n15948));
    jdff dff_B_bLNxqumJ4_2(.din(n15948), .dout(n15951));
    jdff dff_B_bBPrEfQk3_2(.din(n15951), .dout(n15954));
    jdff dff_B_dfR48Bq79_2(.din(n15954), .dout(n15957));
    jdff dff_B_tkF1pB0Z6_2(.din(n15957), .dout(n15960));
    jdff dff_B_4DlmKAeM9_2(.din(n15960), .dout(n15963));
    jdff dff_B_6oKVEMCU6_2(.din(n15963), .dout(n15966));
    jdff dff_B_EnQPCE8p7_2(.din(n15966), .dout(n15969));
    jdff dff_B_cHf5ylHZ9_2(.din(n15969), .dout(n15972));
    jdff dff_B_BAK4Yd0c4_2(.din(n15972), .dout(n15975));
    jdff dff_B_SlQVWnTe7_2(.din(n15975), .dout(n15978));
    jdff dff_B_S8kf8kxz5_2(.din(n15978), .dout(n15981));
    jdff dff_B_fsWyEvLm5_2(.din(n15981), .dout(n15984));
    jdff dff_B_kvg1jy7G3_2(.din(n15984), .dout(n15987));
    jdff dff_B_zxP7er6f1_2(.din(n15987), .dout(n15990));
    jdff dff_B_lYmcxQpE6_2(.din(n15990), .dout(n15993));
    jdff dff_B_dDExMTO48_2(.din(n15993), .dout(n15996));
    jdff dff_B_vl2mcgNi2_2(.din(n15996), .dout(n15999));
    jdff dff_B_TgsGOfhP3_2(.din(n15999), .dout(n16002));
    jdff dff_B_DyxWsHIf6_2(.din(n16002), .dout(n16005));
    jdff dff_B_aPoveLqF9_2(.din(n16005), .dout(n16008));
    jdff dff_B_h1Ll7FdX5_2(.din(n16008), .dout(n16011));
    jdff dff_A_hK4FPsXJ4_1(.din(n3652), .dout(n16013));
    jdff dff_A_IkfscCdt0_0(.din(n16019), .dout(n16016));
    jdff dff_A_o7mAy3Ez9_0(.din(n16022), .dout(n16019));
    jdff dff_A_0GxAqjJG5_0(.din(n16025), .dout(n16022));
    jdff dff_A_5SACCQAh5_0(.din(n16028), .dout(n16025));
    jdff dff_A_Ik0Oth9e5_0(.din(n16031), .dout(n16028));
    jdff dff_A_nsYC6Hbg7_0(.din(n16034), .dout(n16031));
    jdff dff_A_An1SyVrE2_0(.din(n16037), .dout(n16034));
    jdff dff_A_M7gSdpXs0_0(.din(n16040), .dout(n16037));
    jdff dff_A_5rpS1fqF4_0(.din(n16043), .dout(n16040));
    jdff dff_A_pSdRuKNy8_0(.din(n16046), .dout(n16043));
    jdff dff_A_XKVGVf5W9_0(.din(n16049), .dout(n16046));
    jdff dff_A_VWHnLsL63_0(.din(n16052), .dout(n16049));
    jdff dff_A_WEnicOu88_0(.din(n16055), .dout(n16052));
    jdff dff_A_1zrSoqdJ3_0(.din(n16058), .dout(n16055));
    jdff dff_A_yVQzp8SB4_0(.din(n16061), .dout(n16058));
    jdff dff_A_xslBY8zI0_0(.din(n16064), .dout(n16061));
    jdff dff_A_35C7cfdF6_0(.din(n16067), .dout(n16064));
    jdff dff_A_8cBoGORk7_0(.din(n16070), .dout(n16067));
    jdff dff_A_egw93r2D5_0(.din(n16073), .dout(n16070));
    jdff dff_A_WZxTySWC9_0(.din(n16076), .dout(n16073));
    jdff dff_A_DZBG9ZFJ8_0(.din(n16079), .dout(n16076));
    jdff dff_A_R99VK25B9_0(.din(n16082), .dout(n16079));
    jdff dff_A_wHvWHxvY7_0(.din(n16085), .dout(n16082));
    jdff dff_A_Q1y6kjRc2_0(.din(n16088), .dout(n16085));
    jdff dff_A_JRrZcsmk8_0(.din(n16091), .dout(n16088));
    jdff dff_A_LYjliNrx4_0(.din(n16094), .dout(n16091));
    jdff dff_A_vGqp6JRk5_0(.din(n16097), .dout(n16094));
    jdff dff_A_mR8NV3dy0_0(.din(n16100), .dout(n16097));
    jdff dff_A_lBdYvBH87_0(.din(n16103), .dout(n16100));
    jdff dff_A_RC3CelW55_0(.din(n16106), .dout(n16103));
    jdff dff_A_YHXS3FzX4_0(.din(n16109), .dout(n16106));
    jdff dff_A_WlHj1mDf7_0(.din(n16112), .dout(n16109));
    jdff dff_A_eaK2RJ0m7_0(.din(n16115), .dout(n16112));
    jdff dff_A_uca9syKp0_0(.din(n16118), .dout(n16115));
    jdff dff_A_lio901276_0(.din(n16121), .dout(n16118));
    jdff dff_A_1EnTW8GZ1_0(.din(n16124), .dout(n16121));
    jdff dff_A_4lszyFn33_0(.din(n2925), .dout(n16124));
    jdff dff_A_PaeTrKK39_1(.din(n3247), .dout(n16127));
    jdff dff_A_1ezDC40J1_2(.din(n3247), .dout(n16130));
    jdff dff_B_S4ORdUCC3_1(.din(n2932), .dout(n16134));
    jdff dff_B_OKyzk8Am3_2(.din(n2553), .dout(n16137));
    jdff dff_B_QrOMOxpq3_2(.din(n16137), .dout(n16140));
    jdff dff_B_HQ5mZaLc5_2(.din(n16140), .dout(n16143));
    jdff dff_B_mWzklsGZ8_2(.din(n16143), .dout(n16146));
    jdff dff_B_sPbXZwBI1_2(.din(n16146), .dout(n16149));
    jdff dff_B_Hy6mtHDx0_2(.din(n16149), .dout(n16152));
    jdff dff_B_x3l5EV4w5_2(.din(n16152), .dout(n16155));
    jdff dff_B_4cEYmsvB1_2(.din(n16155), .dout(n16158));
    jdff dff_B_8MIdHzbJ5_2(.din(n16158), .dout(n16161));
    jdff dff_B_kdifOqQd7_2(.din(n16161), .dout(n16164));
    jdff dff_B_vrR4YgeA2_2(.din(n16164), .dout(n16167));
    jdff dff_B_lJIkTdyN4_2(.din(n16167), .dout(n16170));
    jdff dff_B_jDm2Xwa08_2(.din(n16170), .dout(n16173));
    jdff dff_B_RYTP8VTC3_2(.din(n16173), .dout(n16176));
    jdff dff_B_HFKsYVuF3_2(.din(n16176), .dout(n16179));
    jdff dff_B_I4ktasz51_2(.din(n16179), .dout(n16182));
    jdff dff_B_nw3p254o3_2(.din(n16182), .dout(n16185));
    jdff dff_B_QimNdpqH1_2(.din(n16185), .dout(n16188));
    jdff dff_B_mbMrcQet5_2(.din(n16188), .dout(n16191));
    jdff dff_B_dy8Lzjex8_2(.din(n16191), .dout(n16194));
    jdff dff_B_30BLDKRy9_2(.din(n16194), .dout(n16197));
    jdff dff_B_1NGgOigZ9_2(.din(n16197), .dout(n16200));
    jdff dff_B_FN4SjH7s3_2(.din(n16200), .dout(n16203));
    jdff dff_B_Ppqrb9gF4_2(.din(n16203), .dout(n16206));
    jdff dff_B_ikvOKAlh6_2(.din(n16206), .dout(n16209));
    jdff dff_B_3TVZMWGu1_2(.din(n16209), .dout(n16212));
    jdff dff_B_KW8k5q2W6_2(.din(n16212), .dout(n16215));
    jdff dff_B_JAMLgE5S9_2(.din(n16215), .dout(n16218));
    jdff dff_B_xLQ3FboZ2_2(.din(n16218), .dout(n16221));
    jdff dff_B_SuUU2NdK7_2(.din(n16221), .dout(n16224));
    jdff dff_B_6GiWr4pP6_2(.din(n16224), .dout(n16227));
    jdff dff_B_iI2UZcQj6_2(.din(n16227), .dout(n16230));
    jdff dff_B_48MqtL2S3_2(.din(n16230), .dout(n16233));
    jdff dff_B_Ch8v8ZGe5_2(.din(n2852), .dout(n16236));
    jdff dff_B_HgCApr8i9_1(.din(n2557), .dout(n16239));
    jdff dff_B_7rpKxDZC5_2(.din(n2202), .dout(n16242));
    jdff dff_B_PA0FYVIU6_2(.din(n16242), .dout(n16245));
    jdff dff_B_udIlobvs4_2(.din(n16245), .dout(n16248));
    jdff dff_B_4RYQuMem5_2(.din(n16248), .dout(n16251));
    jdff dff_B_CrwMvU7m9_2(.din(n16251), .dout(n16254));
    jdff dff_B_tNMH12mS0_2(.din(n16254), .dout(n16257));
    jdff dff_B_l5jHD8MR4_2(.din(n16257), .dout(n16260));
    jdff dff_B_qePmiZwV4_2(.din(n16260), .dout(n16263));
    jdff dff_B_OLuMQmi39_2(.din(n16263), .dout(n16266));
    jdff dff_B_8KIr8lb44_2(.din(n16266), .dout(n16269));
    jdff dff_B_czveACIn4_2(.din(n16269), .dout(n16272));
    jdff dff_B_hAZy3l651_2(.din(n16272), .dout(n16275));
    jdff dff_B_NQ8nkmsP1_2(.din(n16275), .dout(n16278));
    jdff dff_B_fk6Cz92y8_2(.din(n16278), .dout(n16281));
    jdff dff_B_ZqHVFzJZ2_2(.din(n16281), .dout(n16284));
    jdff dff_B_mTFfpFVL5_2(.din(n16284), .dout(n16287));
    jdff dff_B_GDRo23Pv9_2(.din(n16287), .dout(n16290));
    jdff dff_B_QiA1G6pS1_2(.din(n16290), .dout(n16293));
    jdff dff_B_niBFkt3b7_2(.din(n16293), .dout(n16296));
    jdff dff_B_QKoQBLWg2_2(.din(n16296), .dout(n16299));
    jdff dff_B_HEmFGvd54_2(.din(n16299), .dout(n16302));
    jdff dff_B_mKI4ZSl27_2(.din(n16302), .dout(n16305));
    jdff dff_B_jULFZCLS9_2(.din(n16305), .dout(n16308));
    jdff dff_B_KtQEJS3O6_2(.din(n16308), .dout(n16311));
    jdff dff_B_IYezIVQ78_2(.din(n16311), .dout(n16314));
    jdff dff_B_foWNZZ9p7_2(.din(n16314), .dout(n16317));
    jdff dff_B_UZL6lfpx4_2(.din(n16317), .dout(n16320));
    jdff dff_B_ZPYN26713_2(.din(n16320), .dout(n16323));
    jdff dff_B_ellVHP0T5_2(.din(n16323), .dout(n16326));
    jdff dff_B_QaEcDSuD5_2(.din(n16326), .dout(n16329));
    jdff dff_B_TJA2DPQ43_2(.din(n2474), .dout(n16332));
    jdff dff_B_AAk7rBFR0_1(.din(n2206), .dout(n16335));
    jdff dff_B_ZWLLn9iO4_2(.din(n1878), .dout(n16338));
    jdff dff_B_B5DJdmPx2_2(.din(n16338), .dout(n16341));
    jdff dff_B_B0ltlHbD7_2(.din(n16341), .dout(n16344));
    jdff dff_B_rtksfZyz1_2(.din(n16344), .dout(n16347));
    jdff dff_B_IZqBLimd3_2(.din(n16347), .dout(n16350));
    jdff dff_B_L5uThb3m5_2(.din(n16350), .dout(n16353));
    jdff dff_B_edTWyWv18_2(.din(n16353), .dout(n16356));
    jdff dff_B_oXxetAOU7_2(.din(n16356), .dout(n16359));
    jdff dff_B_buIo5cxD3_2(.din(n16359), .dout(n16362));
    jdff dff_B_OzSw6qXi9_2(.din(n16362), .dout(n16365));
    jdff dff_B_TiI6N7T87_2(.din(n16365), .dout(n16368));
    jdff dff_B_RCrHm3Xz7_2(.din(n16368), .dout(n16371));
    jdff dff_B_it2SQyoQ9_2(.din(n16371), .dout(n16374));
    jdff dff_B_QMs1OM2m9_2(.din(n16374), .dout(n16377));
    jdff dff_B_ybz9E4168_2(.din(n16377), .dout(n16380));
    jdff dff_B_zgUtsPIU0_2(.din(n16380), .dout(n16383));
    jdff dff_B_95oHT9fe1_2(.din(n16383), .dout(n16386));
    jdff dff_B_eRILAvIh6_2(.din(n16386), .dout(n16389));
    jdff dff_B_Md6ppQSk7_2(.din(n16389), .dout(n16392));
    jdff dff_B_etzLcrmj9_2(.din(n16392), .dout(n16395));
    jdff dff_B_SinFgzVt4_2(.din(n16395), .dout(n16398));
    jdff dff_B_SvLkIe8e0_2(.din(n16398), .dout(n16401));
    jdff dff_B_1q12hnRw7_2(.din(n16401), .dout(n16404));
    jdff dff_B_xBntAbYr8_2(.din(n16404), .dout(n16407));
    jdff dff_B_An2QI8fG8_2(.din(n16407), .dout(n16410));
    jdff dff_B_ehX91O2y4_2(.din(n16410), .dout(n16413));
    jdff dff_B_SabJs8jz7_2(.din(n16413), .dout(n16416));
    jdff dff_B_hR5poCbV0_2(.din(n2123), .dout(n16419));
    jdff dff_B_E0zn4wyP8_1(.din(n1882), .dout(n16422));
    jdff dff_B_ZZyPhveW8_2(.din(n1581), .dout(n16425));
    jdff dff_B_MIqa1AyF2_2(.din(n16425), .dout(n16428));
    jdff dff_B_qBmtmQtj2_2(.din(n16428), .dout(n16431));
    jdff dff_B_rd3rvPc38_2(.din(n16431), .dout(n16434));
    jdff dff_B_usGTkVpu1_2(.din(n16434), .dout(n16437));
    jdff dff_B_825KKHae9_2(.din(n16437), .dout(n16440));
    jdff dff_B_N8ROcOzd9_2(.din(n16440), .dout(n16443));
    jdff dff_B_xYtmxULo3_2(.din(n16443), .dout(n16446));
    jdff dff_B_nrQD752S8_2(.din(n16446), .dout(n16449));
    jdff dff_B_EMqMMHyE5_2(.din(n16449), .dout(n16452));
    jdff dff_B_Q106ELUE1_2(.din(n16452), .dout(n16455));
    jdff dff_B_uaLusQio5_2(.din(n16455), .dout(n16458));
    jdff dff_B_q8welTEc0_2(.din(n16458), .dout(n16461));
    jdff dff_B_oDDvjCoj2_2(.din(n16461), .dout(n16464));
    jdff dff_B_8HwWkaG32_2(.din(n16464), .dout(n16467));
    jdff dff_B_MIVvcWb63_2(.din(n16467), .dout(n16470));
    jdff dff_B_B0z1MmyT0_2(.din(n16470), .dout(n16473));
    jdff dff_B_9EBzyWvx7_2(.din(n16473), .dout(n16476));
    jdff dff_B_5monQgmX4_2(.din(n16476), .dout(n16479));
    jdff dff_B_rmr0cjqc3_2(.din(n16479), .dout(n16482));
    jdff dff_B_ULDb7L4G2_2(.din(n16482), .dout(n16485));
    jdff dff_B_TtEmYi327_2(.din(n16485), .dout(n16488));
    jdff dff_B_w0Tkh8XO5_2(.din(n16488), .dout(n16491));
    jdff dff_B_q57hWTjr9_2(.din(n16491), .dout(n16494));
    jdff dff_B_0xyfVBWM7_2(.din(n1799), .dout(n16497));
    jdff dff_B_Jh6lq4521_1(.din(n1585), .dout(n16500));
    jdff dff_B_lANTmmel5_2(.din(n1311), .dout(n16503));
    jdff dff_B_0ZG2LOSb2_2(.din(n16503), .dout(n16506));
    jdff dff_B_c7ztxUz32_2(.din(n16506), .dout(n16509));
    jdff dff_B_sXmtubWl5_2(.din(n16509), .dout(n16512));
    jdff dff_B_yb5GS2Gt2_2(.din(n16512), .dout(n16515));
    jdff dff_B_mtJ3BfXa4_2(.din(n16515), .dout(n16518));
    jdff dff_B_KDc0nzDV6_2(.din(n16518), .dout(n16521));
    jdff dff_B_k8XBaHQ05_2(.din(n16521), .dout(n16524));
    jdff dff_B_lJSoHneo5_2(.din(n16524), .dout(n16527));
    jdff dff_B_NSEFXBjI0_2(.din(n16527), .dout(n16530));
    jdff dff_B_rMwsg27l6_2(.din(n16530), .dout(n16533));
    jdff dff_B_BgW5oD0n5_2(.din(n16533), .dout(n16536));
    jdff dff_B_KZPQY57t3_2(.din(n16536), .dout(n16539));
    jdff dff_B_B70Eamoi1_2(.din(n16539), .dout(n16542));
    jdff dff_B_Jl3RscIH9_2(.din(n16542), .dout(n16545));
    jdff dff_B_LcQSTCgc3_2(.din(n16545), .dout(n16548));
    jdff dff_B_UduQqCAt0_2(.din(n16548), .dout(n16551));
    jdff dff_B_mzj2trgd0_2(.din(n16551), .dout(n16554));
    jdff dff_B_uUV632eO3_2(.din(n16554), .dout(n16557));
    jdff dff_B_KPaKpPg85_2(.din(n16557), .dout(n16560));
    jdff dff_B_TLAx6knM4_2(.din(n16560), .dout(n16563));
    jdff dff_B_1M3mdTob1_2(.din(n1502), .dout(n16566));
    jdff dff_B_ZPrv69rY1_1(.din(n1315), .dout(n16569));
    jdff dff_B_lLyytNMO4_2(.din(n1071), .dout(n16572));
    jdff dff_B_q9Gu2eiS7_2(.din(n16572), .dout(n16575));
    jdff dff_B_Qnk4Z3XI8_2(.din(n16575), .dout(n16578));
    jdff dff_B_JDG4hyvH6_2(.din(n16578), .dout(n16581));
    jdff dff_B_YibEVKDh6_2(.din(n16581), .dout(n16584));
    jdff dff_B_mbI4Fcqw5_2(.din(n16584), .dout(n16587));
    jdff dff_B_TYspeDOi8_2(.din(n16587), .dout(n16590));
    jdff dff_B_I7HuwlUW0_2(.din(n16590), .dout(n16593));
    jdff dff_B_ZJeV8KQq0_2(.din(n16593), .dout(n16596));
    jdff dff_B_UyzBVT2o6_2(.din(n16596), .dout(n16599));
    jdff dff_B_D39Jdf8i9_2(.din(n16599), .dout(n16602));
    jdff dff_B_0ErRhg7G6_2(.din(n16602), .dout(n16605));
    jdff dff_B_V8zmzqOd3_2(.din(n16605), .dout(n16608));
    jdff dff_B_vlvm1FA74_2(.din(n16608), .dout(n16611));
    jdff dff_B_Odve1Lhe6_2(.din(n16611), .dout(n16614));
    jdff dff_B_delXOXpE8_2(.din(n16614), .dout(n16617));
    jdff dff_B_bvDYa1ZN5_2(.din(n16617), .dout(n16620));
    jdff dff_B_ciueZflC7_2(.din(n16620), .dout(n16623));
    jdff dff_B_sqKLcQOC4_2(.din(n1232), .dout(n16626));
    jdff dff_B_TLyREf666_1(.din(n1075), .dout(n16629));
    jdff dff_B_IrrZjGgS5_2(.din(n858), .dout(n16632));
    jdff dff_B_cGe2yHM70_2(.din(n16632), .dout(n16635));
    jdff dff_B_1wgzXjHn1_2(.din(n16635), .dout(n16638));
    jdff dff_B_1jjrzbDi0_2(.din(n16638), .dout(n16641));
    jdff dff_B_heFUKkxg4_2(.din(n16641), .dout(n16644));
    jdff dff_B_1VszxwXr2_2(.din(n16644), .dout(n16647));
    jdff dff_B_csLb90T36_2(.din(n16647), .dout(n16650));
    jdff dff_B_R6PbYK4y9_2(.din(n16650), .dout(n16653));
    jdff dff_B_T7akaYFz9_2(.din(n16653), .dout(n16656));
    jdff dff_B_4HVlGHnt6_2(.din(n16656), .dout(n16659));
    jdff dff_B_IfJ7XFg28_2(.din(n16659), .dout(n16662));
    jdff dff_B_YFvkUf2B4_2(.din(n16662), .dout(n16665));
    jdff dff_B_vQSkTbsO0_2(.din(n16665), .dout(n16668));
    jdff dff_B_gOonVgmw2_2(.din(n16668), .dout(n16671));
    jdff dff_B_DlfQu4jH3_2(.din(n16671), .dout(n16674));
    jdff dff_B_jQbxvzmW2_2(.din(n992), .dout(n16677));
    jdff dff_B_genMed2k6_1(.din(n862), .dout(n16680));
    jdff dff_B_euvDCGwU1_2(.din(n672), .dout(n16683));
    jdff dff_B_jm1HdqEf7_2(.din(n16683), .dout(n16686));
    jdff dff_B_PvityzRU3_2(.din(n16686), .dout(n16689));
    jdff dff_B_fbqMY5Fy7_2(.din(n16689), .dout(n16692));
    jdff dff_B_XlrAH4nN9_2(.din(n16692), .dout(n16695));
    jdff dff_B_VDOgafZk5_2(.din(n16695), .dout(n16698));
    jdff dff_B_yIxQC1JB1_2(.din(n16698), .dout(n16701));
    jdff dff_B_R9KdxMF81_2(.din(n16701), .dout(n16704));
    jdff dff_B_PFtbiEVC2_2(.din(n16704), .dout(n16707));
    jdff dff_B_qmSAHCoo1_2(.din(n16707), .dout(n16710));
    jdff dff_B_YeWPrfTF1_2(.din(n16710), .dout(n16713));
    jdff dff_B_4w5HXiWm6_2(.din(n16713), .dout(n16716));
    jdff dff_B_tnSzTt9L3_2(.din(n779), .dout(n16719));
    jdff dff_B_wrVJX94M6_1(.din(n676), .dout(n16722));
    jdff dff_B_895YVFTo0_2(.din(n513), .dout(n16725));
    jdff dff_B_4s2w8K9Y7_2(.din(n16725), .dout(n16728));
    jdff dff_B_ZI8ipCT06_2(.din(n16728), .dout(n16731));
    jdff dff_B_bX9VQi0l8_2(.din(n16731), .dout(n16734));
    jdff dff_B_3eTLC9ts9_2(.din(n16734), .dout(n16737));
    jdff dff_B_042cQft63_2(.din(n16737), .dout(n16740));
    jdff dff_B_Acj0Q3uf9_2(.din(n16740), .dout(n16743));
    jdff dff_B_Hotdf22T6_2(.din(n16743), .dout(n16746));
    jdff dff_B_e4Sw9TXZ8_2(.din(n16746), .dout(n16749));
    jdff dff_B_ezZqCDx86_2(.din(n593), .dout(n16752));
    jdff dff_B_APnmgULd0_1(.din(n517), .dout(n16755));
    jdff dff_B_4chyMujv4_2(.din(n381), .dout(n16758));
    jdff dff_B_OyqFo2pv3_2(.din(n16758), .dout(n16761));
    jdff dff_B_YlC1PFSL0_2(.din(n16761), .dout(n16764));
    jdff dff_B_hgHBTYbN4_2(.din(n16764), .dout(n16767));
    jdff dff_B_RwhEWNGK6_2(.din(n16767), .dout(n16770));
    jdff dff_B_NaR232Rg3_2(.din(n16770), .dout(n16773));
    jdff dff_B_Z5Otzmzb1_2(.din(n434), .dout(n16776));
    jdff dff_B_577uiCVg7_2(.din(n272), .dout(n16779));
    jdff dff_B_sx2C9rLO4_2(.din(n16779), .dout(n16782));
    jdff dff_B_O43b9nPM6_2(.din(n16782), .dout(n16785));
    jdff dff_B_dzB81Hgh7_0(.din(n298), .dout(n16788));
    jdff dff_B_LoIPBci80_0(.din(n4774), .dout(n16791));
    jdff dff_A_qpxHJBxk7_1(.din(n16796), .dout(n16793));
    jdff dff_A_2JNqYLSr2_1(.din(n4760), .dout(n16796));
    jdff dff_B_1fupoCDN4_1(.din(n4451), .dout(n16800));
    jdff dff_B_bDw6z2Oz2_1(.din(n16800), .dout(n16803));
    jdff dff_B_agULwE7d2_2(.din(n4091), .dout(n16806));
    jdff dff_B_9G69aGdd5_2(.din(n16806), .dout(n16809));
    jdff dff_B_tKOA0cNV7_2(.din(n16809), .dout(n16812));
    jdff dff_B_I8NQoZMb0_2(.din(n16812), .dout(n16815));
    jdff dff_B_3d7BK34F9_2(.din(n16815), .dout(n16818));
    jdff dff_B_Z7r1eV5q3_2(.din(n16818), .dout(n16821));
    jdff dff_B_0Lb0Z4XO1_2(.din(n16821), .dout(n16824));
    jdff dff_B_nQFnVsln3_2(.din(n16824), .dout(n16827));
    jdff dff_B_Kb7Zeb3Y6_2(.din(n16827), .dout(n16830));
    jdff dff_B_2X3IdqpE8_2(.din(n16830), .dout(n16833));
    jdff dff_B_AM3Gsmgg2_2(.din(n16833), .dout(n16836));
    jdff dff_B_js2o9Z0f2_2(.din(n16836), .dout(n16839));
    jdff dff_B_jABkcMLU9_2(.din(n16839), .dout(n16842));
    jdff dff_B_GEq0rs3t1_2(.din(n16842), .dout(n16845));
    jdff dff_B_z3jHJwCv0_2(.din(n16845), .dout(n16848));
    jdff dff_B_OsDbvXug6_2(.din(n16848), .dout(n16851));
    jdff dff_B_yCyNaL3H4_2(.din(n16851), .dout(n16854));
    jdff dff_B_qc7t4wag4_2(.din(n16854), .dout(n16857));
    jdff dff_B_zNShhUgA5_2(.din(n16857), .dout(n16860));
    jdff dff_B_ZfHSKcpl7_2(.din(n16860), .dout(n16863));
    jdff dff_B_4nWPXNbs0_2(.din(n16863), .dout(n16866));
    jdff dff_B_p2gXxWfN5_2(.din(n16866), .dout(n16869));
    jdff dff_B_zJyTFgA67_2(.din(n16869), .dout(n16872));
    jdff dff_B_rz3cbqO80_2(.din(n16872), .dout(n16875));
    jdff dff_B_6zMnba1y1_2(.din(n16875), .dout(n16878));
    jdff dff_B_79eag0Im4_2(.din(n16878), .dout(n16881));
    jdff dff_B_s7YJnI191_2(.din(n16881), .dout(n16884));
    jdff dff_B_QQAIagTG4_2(.din(n16884), .dout(n16887));
    jdff dff_B_1lIRuHz28_2(.din(n16887), .dout(n16890));
    jdff dff_B_IidVnOHl6_2(.din(n16890), .dout(n16893));
    jdff dff_B_Tp1iF3st0_2(.din(n16893), .dout(n16896));
    jdff dff_B_WkK6Jg3g3_2(.din(n16896), .dout(n16899));
    jdff dff_B_lH4z1VnS0_2(.din(n16899), .dout(n16902));
    jdff dff_B_rEbARcMs4_2(.din(n16902), .dout(n16905));
    jdff dff_B_g7WqY3Vk1_2(.din(n16905), .dout(n16908));
    jdff dff_B_NUMWLlKW5_2(.din(n16908), .dout(n16911));
    jdff dff_B_JrUy5QGY1_2(.din(n16911), .dout(n16914));
    jdff dff_B_aPPa0fvm0_2(.din(n16914), .dout(n16917));
    jdff dff_B_7H0YXTN93_2(.din(n16917), .dout(n16920));
    jdff dff_B_1nH08Sja8_2(.din(n16920), .dout(n16923));
    jdff dff_B_XG3sNIfl3_2(.din(n16923), .dout(n16926));
    jdff dff_B_yXpJVcTT4_2(.din(n16926), .dout(n16929));
    jdff dff_B_R2JGXC7W8_2(.din(n16929), .dout(n16932));
    jdff dff_B_Yl0vInWa3_2(.din(n16932), .dout(n16935));
    jdff dff_B_wGGF3adj5_2(.din(n16935), .dout(n16938));
    jdff dff_B_cdwtbpXo2_2(.din(n4410), .dout(n16941));
    jdff dff_B_DqGxwHbC1_1(.din(n4098), .dout(n16944));
    jdff dff_B_VV78izEa9_2(.din(n3718), .dout(n16947));
    jdff dff_B_JMfHh7yQ0_2(.din(n16947), .dout(n16950));
    jdff dff_B_ZYCJzGjH1_2(.din(n16950), .dout(n16953));
    jdff dff_B_wf8qKgqo5_2(.din(n16953), .dout(n16956));
    jdff dff_B_Ob14SXDA6_2(.din(n16956), .dout(n16959));
    jdff dff_B_H8wrZPF16_2(.din(n16959), .dout(n16962));
    jdff dff_B_t6MrAjES9_2(.din(n16962), .dout(n16965));
    jdff dff_B_XnWuqa858_2(.din(n16965), .dout(n16968));
    jdff dff_B_kZDBTZal0_2(.din(n16968), .dout(n16971));
    jdff dff_B_6yvoHXFB8_2(.din(n16971), .dout(n16974));
    jdff dff_B_kmO6vQG50_2(.din(n16974), .dout(n16977));
    jdff dff_B_4k5jc4My3_2(.din(n16977), .dout(n16980));
    jdff dff_B_vr977IGf2_2(.din(n16980), .dout(n16983));
    jdff dff_B_nSYaRnhO1_2(.din(n16983), .dout(n16986));
    jdff dff_B_vJ78mm8x6_2(.din(n16986), .dout(n16989));
    jdff dff_B_RyP6E7gn7_2(.din(n16989), .dout(n16992));
    jdff dff_B_Myshnbe47_2(.din(n16992), .dout(n16995));
    jdff dff_B_qKkLw8Kc0_2(.din(n16995), .dout(n16998));
    jdff dff_B_IisZFHk28_2(.din(n16998), .dout(n17001));
    jdff dff_B_173zE3wI9_2(.din(n17001), .dout(n17004));
    jdff dff_B_iRmfp9v25_2(.din(n17004), .dout(n17007));
    jdff dff_B_Q9WrxAtQ0_2(.din(n17007), .dout(n17010));
    jdff dff_B_IneNu71y8_2(.din(n17010), .dout(n17013));
    jdff dff_B_u2K4lrpV7_2(.din(n17013), .dout(n17016));
    jdff dff_B_gfMryNpa4_2(.din(n17016), .dout(n17019));
    jdff dff_B_fRjP8YWz6_2(.din(n17019), .dout(n17022));
    jdff dff_B_D5pOJyV48_2(.din(n17022), .dout(n17025));
    jdff dff_B_lrRpCMSJ2_2(.din(n17025), .dout(n17028));
    jdff dff_B_Xvy2Y6VW9_2(.din(n17028), .dout(n17031));
    jdff dff_B_kapuTbQO3_2(.din(n17031), .dout(n17034));
    jdff dff_B_XGW6OSEY6_2(.din(n17034), .dout(n17037));
    jdff dff_B_vCc9X8W45_2(.din(n17037), .dout(n17040));
    jdff dff_B_it0Mh74z4_2(.din(n17040), .dout(n17043));
    jdff dff_B_hFTNOiXp8_2(.din(n17043), .dout(n17046));
    jdff dff_B_r37wjaCq0_2(.din(n17046), .dout(n17049));
    jdff dff_B_xdNBrZCi3_2(.din(n17049), .dout(n17052));
    jdff dff_B_hbOlwcAs2_2(.din(n17052), .dout(n17055));
    jdff dff_B_czKOHofc8_2(.din(n17055), .dout(n17058));
    jdff dff_B_ygtjzrFC1_2(.din(n17058), .dout(n17061));
    jdff dff_B_QYiA9Km83_2(.din(n17061), .dout(n17064));
    jdff dff_B_73M7BQO13_2(.din(n17064), .dout(n17067));
    jdff dff_B_falzzeP72_2(.din(n4027), .dout(n17070));
    jdff dff_B_hUWPJ5Ia0_1(.din(n3722), .dout(n17073));
    jdff dff_B_38pXlEXW0_2(.din(n3338), .dout(n17076));
    jdff dff_B_Crpe4JDv4_2(.din(n17076), .dout(n17079));
    jdff dff_B_97xQvbry6_2(.din(n17079), .dout(n17082));
    jdff dff_B_mrqPKc1Z9_2(.din(n17082), .dout(n17085));
    jdff dff_B_jt0FEUrP4_2(.din(n17085), .dout(n17088));
    jdff dff_B_mGJMO9eB6_2(.din(n17088), .dout(n17091));
    jdff dff_B_RT6MvAg04_2(.din(n17091), .dout(n17094));
    jdff dff_B_1LtO1l2e5_2(.din(n17094), .dout(n17097));
    jdff dff_B_Q2eDYiTU0_2(.din(n17097), .dout(n17100));
    jdff dff_B_ezHkWKvm5_2(.din(n17100), .dout(n17103));
    jdff dff_B_M6PcMdri6_2(.din(n17103), .dout(n17106));
    jdff dff_B_P3VgKcs09_2(.din(n17106), .dout(n17109));
    jdff dff_B_yBk1mHDO0_2(.din(n17109), .dout(n17112));
    jdff dff_B_BlxQOUZS7_2(.din(n17112), .dout(n17115));
    jdff dff_B_ltFOv6Vo1_2(.din(n17115), .dout(n17118));
    jdff dff_B_4J8Yf2W26_2(.din(n17118), .dout(n17121));
    jdff dff_B_BYr64GK65_2(.din(n17121), .dout(n17124));
    jdff dff_B_8rB9nKcx1_2(.din(n17124), .dout(n17127));
    jdff dff_B_wqUHvkBj8_2(.din(n17127), .dout(n17130));
    jdff dff_B_ywuXpUg47_2(.din(n17130), .dout(n17133));
    jdff dff_B_8gURS7ci2_2(.din(n17133), .dout(n17136));
    jdff dff_B_7jpLkQnA1_2(.din(n17136), .dout(n17139));
    jdff dff_B_ZxD3NAAN4_2(.din(n17139), .dout(n17142));
    jdff dff_B_V06AWYwM1_2(.din(n17142), .dout(n17145));
    jdff dff_B_9SUaudRb2_2(.din(n17145), .dout(n17148));
    jdff dff_B_VrWv7SJo9_2(.din(n17148), .dout(n17151));
    jdff dff_B_Apnxg2Su3_2(.din(n17151), .dout(n17154));
    jdff dff_B_a4hT12As6_2(.din(n17154), .dout(n17157));
    jdff dff_B_iJMMg6Ci0_2(.din(n17157), .dout(n17160));
    jdff dff_B_udsFMJq63_2(.din(n17160), .dout(n17163));
    jdff dff_B_nh31iq2e9_2(.din(n17163), .dout(n17166));
    jdff dff_B_3OVzZOA39_2(.din(n17166), .dout(n17169));
    jdff dff_B_HTKKiomk7_2(.din(n17169), .dout(n17172));
    jdff dff_B_35qTgeS53_2(.din(n17172), .dout(n17175));
    jdff dff_B_Zn1pUUIV4_2(.din(n17175), .dout(n17178));
    jdff dff_B_TERMiXSN4_2(.din(n17178), .dout(n17181));
    jdff dff_B_0s0TzxQu7_2(.din(n3644), .dout(n17184));
    jdff dff_B_kcbxlRjy9_1(.din(n3342), .dout(n17187));
    jdff dff_B_sXUB0K114_2(.din(n2947), .dout(n17190));
    jdff dff_B_YYgudbEX2_2(.din(n17190), .dout(n17193));
    jdff dff_B_vJXMOotG0_2(.din(n17193), .dout(n17196));
    jdff dff_B_NTZ2dVIL2_2(.din(n17196), .dout(n17199));
    jdff dff_B_X4nHCl4w9_2(.din(n17199), .dout(n17202));
    jdff dff_B_gAE62IgG1_2(.din(n17202), .dout(n17205));
    jdff dff_B_aQZGDkUz8_2(.din(n17205), .dout(n17208));
    jdff dff_B_onVMGKRj3_2(.din(n17208), .dout(n17211));
    jdff dff_B_FgjOxEOF1_2(.din(n17211), .dout(n17214));
    jdff dff_B_bfyIWMSJ1_2(.din(n17214), .dout(n17217));
    jdff dff_B_xDZnBuEW5_2(.din(n17217), .dout(n17220));
    jdff dff_B_GErPVUKH1_2(.din(n17220), .dout(n17223));
    jdff dff_B_Gd7Hg6vj8_2(.din(n17223), .dout(n17226));
    jdff dff_B_pMVFnvOx5_2(.din(n17226), .dout(n17229));
    jdff dff_B_AehMOhl39_2(.din(n17229), .dout(n17232));
    jdff dff_B_TpH9i84D8_2(.din(n17232), .dout(n17235));
    jdff dff_B_AQPdMPZB4_2(.din(n17235), .dout(n17238));
    jdff dff_B_GU4ROdY50_2(.din(n17238), .dout(n17241));
    jdff dff_B_hoyULrMt1_2(.din(n17241), .dout(n17244));
    jdff dff_B_REC2RIuZ3_2(.din(n17244), .dout(n17247));
    jdff dff_B_3WRI4TEW0_2(.din(n17247), .dout(n17250));
    jdff dff_B_AOovrG2I8_2(.din(n17250), .dout(n17253));
    jdff dff_B_iVdF1zSj9_2(.din(n17253), .dout(n17256));
    jdff dff_B_CSJejrr00_2(.din(n17256), .dout(n17259));
    jdff dff_B_TmgQY7aq7_2(.din(n17259), .dout(n17262));
    jdff dff_B_h0FRUO3j1_2(.din(n17262), .dout(n17265));
    jdff dff_B_cxljlFJk5_2(.din(n17265), .dout(n17268));
    jdff dff_B_YT0MdckA4_2(.din(n17268), .dout(n17271));
    jdff dff_B_G4X87IfJ0_2(.din(n17271), .dout(n17274));
    jdff dff_B_CXA7bD8E7_2(.din(n17274), .dout(n17277));
    jdff dff_B_Kr04a6zH7_2(.din(n17277), .dout(n17280));
    jdff dff_B_wiemeGC85_2(.din(n17280), .dout(n17283));
    jdff dff_B_6PAvUIMV1_2(.din(n17283), .dout(n17286));
    jdff dff_B_2oTC1IeI8_2(.din(n3239), .dout(n17289));
    jdff dff_B_ga3xMME42_1(.din(n2951), .dout(n17292));
    jdff dff_B_vTMbvAtu7_2(.din(n2572), .dout(n17295));
    jdff dff_B_G4nAPH1o3_2(.din(n17295), .dout(n17298));
    jdff dff_B_NnmeNfwY3_2(.din(n17298), .dout(n17301));
    jdff dff_B_rfwclIUl9_2(.din(n17301), .dout(n17304));
    jdff dff_B_2qcbZqSG7_2(.din(n17304), .dout(n17307));
    jdff dff_B_Jv9X6WHL8_2(.din(n17307), .dout(n17310));
    jdff dff_B_7tMLKjnG5_2(.din(n17310), .dout(n17313));
    jdff dff_B_7001iSvU5_2(.din(n17313), .dout(n17316));
    jdff dff_B_i7ycTdzN4_2(.din(n17316), .dout(n17319));
    jdff dff_B_IIDlM1ND3_2(.din(n17319), .dout(n17322));
    jdff dff_B_9dRHixW77_2(.din(n17322), .dout(n17325));
    jdff dff_B_PYVcYUhh0_2(.din(n17325), .dout(n17328));
    jdff dff_B_6uRsDfVo0_2(.din(n17328), .dout(n17331));
    jdff dff_B_bIISXcli7_2(.din(n17331), .dout(n17334));
    jdff dff_B_Et2FDZtn3_2(.din(n17334), .dout(n17337));
    jdff dff_B_8qZZ8Nt57_2(.din(n17337), .dout(n17340));
    jdff dff_B_AERnxkmb3_2(.din(n17340), .dout(n17343));
    jdff dff_B_dpix5o353_2(.din(n17343), .dout(n17346));
    jdff dff_B_XSC01LDr4_2(.din(n17346), .dout(n17349));
    jdff dff_B_VzC8j6nj0_2(.din(n17349), .dout(n17352));
    jdff dff_B_rXnnaJ8p2_2(.din(n17352), .dout(n17355));
    jdff dff_B_99nxWuam3_2(.din(n17355), .dout(n17358));
    jdff dff_B_7xjFRmPL5_2(.din(n17358), .dout(n17361));
    jdff dff_B_mRuCOBGJ1_2(.din(n17361), .dout(n17364));
    jdff dff_B_oXeNmgWz7_2(.din(n17364), .dout(n17367));
    jdff dff_B_ycWV6Zts4_2(.din(n17367), .dout(n17370));
    jdff dff_B_fZhepIFF1_2(.din(n17370), .dout(n17373));
    jdff dff_B_5V2BFPIT7_2(.din(n17373), .dout(n17376));
    jdff dff_B_MY9aCvZg6_2(.din(n17376), .dout(n17379));
    jdff dff_B_dn6khCWy1_2(.din(n17379), .dout(n17382));
    jdff dff_B_kQ3pLChE1_2(.din(n2844), .dout(n17385));
    jdff dff_B_72vJHDRm4_1(.din(n2576), .dout(n17388));
    jdff dff_B_WNXECbNp2_2(.din(n2221), .dout(n17391));
    jdff dff_B_6yy8D0MW7_2(.din(n17391), .dout(n17394));
    jdff dff_B_095mUswf9_2(.din(n17394), .dout(n17397));
    jdff dff_B_ra6e7fzJ3_2(.din(n17397), .dout(n17400));
    jdff dff_B_bnGmFO3i5_2(.din(n17400), .dout(n17403));
    jdff dff_B_dIlXzTbE6_2(.din(n17403), .dout(n17406));
    jdff dff_B_ke0Ex4BD3_2(.din(n17406), .dout(n17409));
    jdff dff_B_KAHiQ5MD5_2(.din(n17409), .dout(n17412));
    jdff dff_B_bQJjeAAb6_2(.din(n17412), .dout(n17415));
    jdff dff_B_S8pShqH10_2(.din(n17415), .dout(n17418));
    jdff dff_B_MxzhyBte1_2(.din(n17418), .dout(n17421));
    jdff dff_B_jbY18xuA5_2(.din(n17421), .dout(n17424));
    jdff dff_B_GjZpbovM5_2(.din(n17424), .dout(n17427));
    jdff dff_B_NsfHKnrZ2_2(.din(n17427), .dout(n17430));
    jdff dff_B_WaTfX6FN6_2(.din(n17430), .dout(n17433));
    jdff dff_B_arKz1MVK2_2(.din(n17433), .dout(n17436));
    jdff dff_B_Ud9JqVjp2_2(.din(n17436), .dout(n17439));
    jdff dff_B_wf0MDSsA7_2(.din(n17439), .dout(n17442));
    jdff dff_B_GvL24ZfN1_2(.din(n17442), .dout(n17445));
    jdff dff_B_M83a0Eab1_2(.din(n17445), .dout(n17448));
    jdff dff_B_ME0FJdGH6_2(.din(n17448), .dout(n17451));
    jdff dff_B_mQ5KoUqM3_2(.din(n17451), .dout(n17454));
    jdff dff_B_87p6jvvS3_2(.din(n17454), .dout(n17457));
    jdff dff_B_0HG02Vwh6_2(.din(n17457), .dout(n17460));
    jdff dff_B_UfNS9ONN4_2(.din(n17460), .dout(n17463));
    jdff dff_B_Toz374d67_2(.din(n17463), .dout(n17466));
    jdff dff_B_SVn0Kq5S2_2(.din(n17466), .dout(n17469));
    jdff dff_B_QMXPycXa7_2(.din(n2466), .dout(n17472));
    jdff dff_B_pzUmcCNM8_1(.din(n2225), .dout(n17475));
    jdff dff_B_C42Mg9dF7_2(.din(n1897), .dout(n17478));
    jdff dff_B_pVjvpTb82_2(.din(n17478), .dout(n17481));
    jdff dff_B_QZ5Ergr54_2(.din(n17481), .dout(n17484));
    jdff dff_B_0F1z5oQc6_2(.din(n17484), .dout(n17487));
    jdff dff_B_UeUDiyVH4_2(.din(n17487), .dout(n17490));
    jdff dff_B_LanzuH9v9_2(.din(n17490), .dout(n17493));
    jdff dff_B_z233RMrP0_2(.din(n17493), .dout(n17496));
    jdff dff_B_NqmiiqCc0_2(.din(n17496), .dout(n17499));
    jdff dff_B_FkWLYgRS5_2(.din(n17499), .dout(n17502));
    jdff dff_B_cGomwskl3_2(.din(n17502), .dout(n17505));
    jdff dff_B_hqs1QI3m7_2(.din(n17505), .dout(n17508));
    jdff dff_B_SMA1iwBW7_2(.din(n17508), .dout(n17511));
    jdff dff_B_8CGju51P5_2(.din(n17511), .dout(n17514));
    jdff dff_B_4P63Sk099_2(.din(n17514), .dout(n17517));
    jdff dff_B_8RovYKMb4_2(.din(n17517), .dout(n17520));
    jdff dff_B_fmaC9uC59_2(.din(n17520), .dout(n17523));
    jdff dff_B_lF1rxL5v7_2(.din(n17523), .dout(n17526));
    jdff dff_B_Cwkc5HQG3_2(.din(n17526), .dout(n17529));
    jdff dff_B_aKonAQ029_2(.din(n17529), .dout(n17532));
    jdff dff_B_qCDbyKzR8_2(.din(n17532), .dout(n17535));
    jdff dff_B_tmX8AwQQ1_2(.din(n17535), .dout(n17538));
    jdff dff_B_0YCRTGia0_2(.din(n17538), .dout(n17541));
    jdff dff_B_dLSiwg0c4_2(.din(n17541), .dout(n17544));
    jdff dff_B_uGOp2fnT2_2(.din(n17544), .dout(n17547));
    jdff dff_B_m8OWrTci8_2(.din(n2115), .dout(n17550));
    jdff dff_B_TF5vSIb98_1(.din(n1901), .dout(n17553));
    jdff dff_B_tQ4qXZ1x6_2(.din(n1600), .dout(n17556));
    jdff dff_B_mClwyOzS8_2(.din(n17556), .dout(n17559));
    jdff dff_B_Kxlplazs1_2(.din(n17559), .dout(n17562));
    jdff dff_B_N5a60De67_2(.din(n17562), .dout(n17565));
    jdff dff_B_ektGJC4b7_2(.din(n17565), .dout(n17568));
    jdff dff_B_kUC2MXDG0_2(.din(n17568), .dout(n17571));
    jdff dff_B_BWCi4y7u3_2(.din(n17571), .dout(n17574));
    jdff dff_B_yKfef8Pu0_2(.din(n17574), .dout(n17577));
    jdff dff_B_Fp8V6JlI0_2(.din(n17577), .dout(n17580));
    jdff dff_B_DnZORb424_2(.din(n17580), .dout(n17583));
    jdff dff_B_7p2Mnrod6_2(.din(n17583), .dout(n17586));
    jdff dff_B_NzmfXrmJ6_2(.din(n17586), .dout(n17589));
    jdff dff_B_CkSWZqT83_2(.din(n17589), .dout(n17592));
    jdff dff_B_Gb3iBuFG9_2(.din(n17592), .dout(n17595));
    jdff dff_B_mOkqK3Gg9_2(.din(n17595), .dout(n17598));
    jdff dff_B_JWUZTMPr4_2(.din(n17598), .dout(n17601));
    jdff dff_B_AyP0BeJS5_2(.din(n17601), .dout(n17604));
    jdff dff_B_2AWjIdOv7_2(.din(n17604), .dout(n17607));
    jdff dff_B_oh0qzwZ21_2(.din(n17607), .dout(n17610));
    jdff dff_B_2gms4NKT4_2(.din(n17610), .dout(n17613));
    jdff dff_B_1obje77m9_2(.din(n17613), .dout(n17616));
    jdff dff_B_yR9CiLXM5_2(.din(n1791), .dout(n17619));
    jdff dff_B_dbiXsX4n4_1(.din(n1604), .dout(n17622));
    jdff dff_B_S6ClhJNw1_2(.din(n1330), .dout(n17625));
    jdff dff_B_WSKv8KBR4_2(.din(n17625), .dout(n17628));
    jdff dff_B_xbLX4O0F3_2(.din(n17628), .dout(n17631));
    jdff dff_B_S23IViRA3_2(.din(n17631), .dout(n17634));
    jdff dff_B_W2KmOD0e8_2(.din(n17634), .dout(n17637));
    jdff dff_B_8F2KyJNg0_2(.din(n17637), .dout(n17640));
    jdff dff_B_cCmCpYAe2_2(.din(n17640), .dout(n17643));
    jdff dff_B_4ViM8jpT8_2(.din(n17643), .dout(n17646));
    jdff dff_B_iqCsRr4K0_2(.din(n17646), .dout(n17649));
    jdff dff_B_b3U0LBdv4_2(.din(n17649), .dout(n17652));
    jdff dff_B_GxMsT4im8_2(.din(n17652), .dout(n17655));
    jdff dff_B_esmiuX8b5_2(.din(n17655), .dout(n17658));
    jdff dff_B_3HHKbp6f0_2(.din(n17658), .dout(n17661));
    jdff dff_B_PLmQuOCZ8_2(.din(n17661), .dout(n17664));
    jdff dff_B_mkCIRXr34_2(.din(n17664), .dout(n17667));
    jdff dff_B_iOstxyim7_2(.din(n17667), .dout(n17670));
    jdff dff_B_IV2nnOEA5_2(.din(n17670), .dout(n17673));
    jdff dff_B_0vg8Nkm94_2(.din(n17673), .dout(n17676));
    jdff dff_B_a3vhh17j0_2(.din(n1494), .dout(n17679));
    jdff dff_B_8KXdKmmc6_1(.din(n1334), .dout(n17682));
    jdff dff_B_81DpVl7v2_2(.din(n1090), .dout(n17685));
    jdff dff_B_kAjE0D7I4_2(.din(n17685), .dout(n17688));
    jdff dff_B_RAeSevz53_2(.din(n17688), .dout(n17691));
    jdff dff_B_IuAArMSN9_2(.din(n17691), .dout(n17694));
    jdff dff_B_DgacSUbd6_2(.din(n17694), .dout(n17697));
    jdff dff_B_N6zbtjUG2_2(.din(n17697), .dout(n17700));
    jdff dff_B_87EYA9Y24_2(.din(n17700), .dout(n17703));
    jdff dff_B_j7nDCuoL8_2(.din(n17703), .dout(n17706));
    jdff dff_B_7EixtPTM1_2(.din(n17706), .dout(n17709));
    jdff dff_B_eJVg4sHJ5_2(.din(n17709), .dout(n17712));
    jdff dff_B_VMoPedRs6_2(.din(n17712), .dout(n17715));
    jdff dff_B_01JQ4hfl9_2(.din(n17715), .dout(n17718));
    jdff dff_B_DjleBzKY8_2(.din(n17718), .dout(n17721));
    jdff dff_B_c9L2D4CH9_2(.din(n17721), .dout(n17724));
    jdff dff_B_4GGfpT8Z2_2(.din(n17724), .dout(n17727));
    jdff dff_B_hUuxM9Cj6_2(.din(n1224), .dout(n17730));
    jdff dff_B_npBmo3FI2_1(.din(n1094), .dout(n17733));
    jdff dff_B_RhK0niGN5_2(.din(n877), .dout(n17736));
    jdff dff_B_OEwf7hP66_2(.din(n17736), .dout(n17739));
    jdff dff_B_MtaKCeQ73_2(.din(n17739), .dout(n17742));
    jdff dff_B_cqrkvAVp5_2(.din(n17742), .dout(n17745));
    jdff dff_B_NgYT9d8Q1_2(.din(n17745), .dout(n17748));
    jdff dff_B_K1oAFODJ0_2(.din(n17748), .dout(n17751));
    jdff dff_B_7lGNjVI75_2(.din(n17751), .dout(n17754));
    jdff dff_B_kWvFYJsq6_2(.din(n17754), .dout(n17757));
    jdff dff_B_1vqvDT3b4_2(.din(n17757), .dout(n17760));
    jdff dff_B_4jZlZdKo0_2(.din(n17760), .dout(n17763));
    jdff dff_B_eHDaJjSf8_2(.din(n17763), .dout(n17766));
    jdff dff_B_YuxiLJVP8_2(.din(n17766), .dout(n17769));
    jdff dff_B_FPWiNprk3_2(.din(n984), .dout(n17772));
    jdff dff_B_Y4Mwki8N8_1(.din(n881), .dout(n17775));
    jdff dff_B_buPbW46o2_2(.din(n691), .dout(n17778));
    jdff dff_B_SDqNf5448_2(.din(n17778), .dout(n17781));
    jdff dff_B_jdejU4C27_2(.din(n17781), .dout(n17784));
    jdff dff_B_0AFkGHTD9_2(.din(n17784), .dout(n17787));
    jdff dff_B_NAGmiFYT7_2(.din(n17787), .dout(n17790));
    jdff dff_B_taqlKBRo7_2(.din(n17790), .dout(n17793));
    jdff dff_B_brYJ81LH6_2(.din(n17793), .dout(n17796));
    jdff dff_B_lNswk0dg6_2(.din(n17796), .dout(n17799));
    jdff dff_B_NoOfWuhP6_2(.din(n17799), .dout(n17802));
    jdff dff_B_uVj7vMka2_2(.din(n771), .dout(n17805));
    jdff dff_B_FHDfKqcc2_1(.din(n695), .dout(n17808));
    jdff dff_B_fUk4hqjq2_2(.din(n532), .dout(n17811));
    jdff dff_B_NMJW5qQQ6_2(.din(n17811), .dout(n17814));
    jdff dff_B_p0VVpxOD7_2(.din(n17814), .dout(n17817));
    jdff dff_B_fcmW6xwU6_2(.din(n17817), .dout(n17820));
    jdff dff_B_guLnpw2S4_2(.din(n17820), .dout(n17823));
    jdff dff_B_Z7m1PGz53_2(.din(n17823), .dout(n17826));
    jdff dff_B_9pL1rP5c5_2(.din(n585), .dout(n17829));
    jdff dff_B_2iH3l9Ps9_2(.din(n403), .dout(n17832));
    jdff dff_B_rcPjiLWS1_2(.din(n17832), .dout(n17835));
    jdff dff_B_qFMZlzBN6_2(.din(n17835), .dout(n17838));
    jdff dff_B_p96wqOZf1_0(.din(n422), .dout(n17841));
    jdff dff_A_hn2ihA4X7_0(.din(n17846), .dout(n17843));
    jdff dff_A_uRE18QYz7_0(.din(n286), .dout(n17846));
    jdff dff_A_9DHjInrX5_0(.din(n17852), .dout(n17849));
    jdff dff_A_VnVkTe6E1_0(.din(n283), .dout(n17852));
    jdff dff_B_QzRqY8Wk5_1(.din(n4796), .dout(n17856));
    jdff dff_B_EkBsbp5C6_2(.din(n4463), .dout(n17859));
    jdff dff_B_V9gy66MR8_2(.din(n17859), .dout(n17862));
    jdff dff_B_yvxOb0tX3_2(.din(n17862), .dout(n17865));
    jdff dff_B_0htVR8JQ3_2(.din(n17865), .dout(n17868));
    jdff dff_B_kgx9rspv3_2(.din(n17868), .dout(n17871));
    jdff dff_B_wW5J3Qoh9_2(.din(n17871), .dout(n17874));
    jdff dff_B_soxLtRFc3_2(.din(n17874), .dout(n17877));
    jdff dff_B_FWVnXE4p0_2(.din(n17877), .dout(n17880));
    jdff dff_B_WzvgQYNR4_2(.din(n17880), .dout(n17883));
    jdff dff_B_mAyzAEGv6_2(.din(n17883), .dout(n17886));
    jdff dff_B_5kND4eji3_2(.din(n17886), .dout(n17889));
    jdff dff_B_DbAaB1HS5_2(.din(n17889), .dout(n17892));
    jdff dff_B_e4KXCDof2_2(.din(n17892), .dout(n17895));
    jdff dff_B_49mKgtxF0_2(.din(n17895), .dout(n17898));
    jdff dff_B_9CdU1SOe2_2(.din(n17898), .dout(n17901));
    jdff dff_B_5hYqEvx10_2(.din(n17901), .dout(n17904));
    jdff dff_B_pvutrAiR3_2(.din(n17904), .dout(n17907));
    jdff dff_B_AqLBlfe52_2(.din(n17907), .dout(n17910));
    jdff dff_B_2GA041mq3_2(.din(n17910), .dout(n17913));
    jdff dff_B_C2zU20Io9_2(.din(n17913), .dout(n17916));
    jdff dff_B_rU33edgr0_2(.din(n17916), .dout(n17919));
    jdff dff_B_OjLXyaVm5_2(.din(n17919), .dout(n17922));
    jdff dff_B_81I1jSqI7_2(.din(n17922), .dout(n17925));
    jdff dff_B_U93Whbfi2_2(.din(n17925), .dout(n17928));
    jdff dff_B_OyWiSILw4_2(.din(n17928), .dout(n17931));
    jdff dff_B_4PLsqf2P9_2(.din(n17931), .dout(n17934));
    jdff dff_B_YFt1gIIa4_2(.din(n17934), .dout(n17937));
    jdff dff_B_v7PNWjxa0_2(.din(n17937), .dout(n17940));
    jdff dff_B_z7Ry1QkT6_2(.din(n17940), .dout(n17943));
    jdff dff_B_cDt5Zpe71_2(.din(n17943), .dout(n17946));
    jdff dff_B_OoEpJWQ75_2(.din(n17946), .dout(n17949));
    jdff dff_B_qZ5tv5vY1_2(.din(n17949), .dout(n17952));
    jdff dff_B_kwTMnRty0_2(.din(n17952), .dout(n17955));
    jdff dff_B_1Xdjdf6N3_2(.din(n17955), .dout(n17958));
    jdff dff_B_Pmgh6Obo0_2(.din(n17958), .dout(n17961));
    jdff dff_B_AnrDfWcl1_2(.din(n17961), .dout(n17964));
    jdff dff_B_cROquOB40_2(.din(n17964), .dout(n17967));
    jdff dff_B_8iPXoG4N2_2(.din(n17967), .dout(n17970));
    jdff dff_B_dFmAg3GA4_2(.din(n17970), .dout(n17973));
    jdff dff_B_MBQbCFaM1_2(.din(n17973), .dout(n17976));
    jdff dff_B_r03NUlUN3_2(.din(n17976), .dout(n17979));
    jdff dff_B_XQyldepu8_2(.din(n17979), .dout(n17982));
    jdff dff_B_ihKtn3974_2(.din(n17982), .dout(n17985));
    jdff dff_B_lMmJApGb6_2(.din(n17985), .dout(n17988));
    jdff dff_B_qZbCVfzj9_0(.din(n4792), .dout(n17991));
    jdff dff_A_KSJU7kjs1_1(.din(n4749), .dout(n17993));
    jdff dff_B_PIGqr8be1_1(.din(n4467), .dout(n17997));
    jdff dff_B_Ty8a6ple1_2(.din(n4113), .dout(n18000));
    jdff dff_B_TgjVLXRI8_2(.din(n18000), .dout(n18003));
    jdff dff_B_iX1SIyCK9_2(.din(n18003), .dout(n18006));
    jdff dff_B_Bpbbljzn2_2(.din(n18006), .dout(n18009));
    jdff dff_B_BWbAjSqr9_2(.din(n18009), .dout(n18012));
    jdff dff_B_QiCnsXfR8_2(.din(n18012), .dout(n18015));
    jdff dff_B_ndOyVV2j6_2(.din(n18015), .dout(n18018));
    jdff dff_B_61lASTgb5_2(.din(n18018), .dout(n18021));
    jdff dff_B_5DdOldDp4_2(.din(n18021), .dout(n18024));
    jdff dff_B_MW2rohRv5_2(.din(n18024), .dout(n18027));
    jdff dff_B_vw7WS6Vh2_2(.din(n18027), .dout(n18030));
    jdff dff_B_O72Qgpf74_2(.din(n18030), .dout(n18033));
    jdff dff_B_y1TaDchZ3_2(.din(n18033), .dout(n18036));
    jdff dff_B_tUTWzf819_2(.din(n18036), .dout(n18039));
    jdff dff_B_YFiYT1dE0_2(.din(n18039), .dout(n18042));
    jdff dff_B_zvHLBJFV5_2(.din(n18042), .dout(n18045));
    jdff dff_B_2Mx7iK5f4_2(.din(n18045), .dout(n18048));
    jdff dff_B_bRBWLhek8_2(.din(n18048), .dout(n18051));
    jdff dff_B_otkSlVI13_2(.din(n18051), .dout(n18054));
    jdff dff_B_ENapcN2Q7_2(.din(n18054), .dout(n18057));
    jdff dff_B_wznB5eDK4_2(.din(n18057), .dout(n18060));
    jdff dff_B_3GKlaIZe6_2(.din(n18060), .dout(n18063));
    jdff dff_B_uoHfKMwe3_2(.din(n18063), .dout(n18066));
    jdff dff_B_QUFRqTmT9_2(.din(n18066), .dout(n18069));
    jdff dff_B_DtG11sPz5_2(.din(n18069), .dout(n18072));
    jdff dff_B_XgtGxpl03_2(.din(n18072), .dout(n18075));
    jdff dff_B_1vmPD2DE7_2(.din(n18075), .dout(n18078));
    jdff dff_B_YZQ42WSY0_2(.din(n18078), .dout(n18081));
    jdff dff_B_KYsVBEqh2_2(.din(n18081), .dout(n18084));
    jdff dff_B_sQAQDt9x0_2(.din(n18084), .dout(n18087));
    jdff dff_B_oyWSxQ8s7_2(.din(n18087), .dout(n18090));
    jdff dff_B_VVkazXL08_2(.din(n18090), .dout(n18093));
    jdff dff_B_p14iwy2s5_2(.din(n18093), .dout(n18096));
    jdff dff_B_nWvH51cH1_2(.din(n18096), .dout(n18099));
    jdff dff_B_mXrTqje64_2(.din(n18099), .dout(n18102));
    jdff dff_B_mMzPzBnB3_2(.din(n18102), .dout(n18105));
    jdff dff_B_pDd7DsGf2_2(.din(n18105), .dout(n18108));
    jdff dff_B_7UA23h9k2_2(.din(n18108), .dout(n18111));
    jdff dff_B_b70qJSYz4_2(.din(n18111), .dout(n18114));
    jdff dff_B_5iKIACOp3_2(.din(n4399), .dout(n18117));
    jdff dff_B_sd11iQz02_1(.din(n4117), .dout(n18120));
    jdff dff_B_hEbWQPmX7_2(.din(n3737), .dout(n18123));
    jdff dff_B_iSAHyJDU1_2(.din(n18123), .dout(n18126));
    jdff dff_B_fWquE1lm3_2(.din(n18126), .dout(n18129));
    jdff dff_B_IXoj6phy2_2(.din(n18129), .dout(n18132));
    jdff dff_B_F6nurJeV8_2(.din(n18132), .dout(n18135));
    jdff dff_B_6BhQ51V03_2(.din(n18135), .dout(n18138));
    jdff dff_B_bCwoT1087_2(.din(n18138), .dout(n18141));
    jdff dff_B_63redlre2_2(.din(n18141), .dout(n18144));
    jdff dff_B_KhVip9yp2_2(.din(n18144), .dout(n18147));
    jdff dff_B_9eFEpYFy0_2(.din(n18147), .dout(n18150));
    jdff dff_B_IiLtqin01_2(.din(n18150), .dout(n18153));
    jdff dff_B_p2cgsK5s6_2(.din(n18153), .dout(n18156));
    jdff dff_B_of7gZplG1_2(.din(n18156), .dout(n18159));
    jdff dff_B_bs3hwhOS7_2(.din(n18159), .dout(n18162));
    jdff dff_B_eduZAaEZ4_2(.din(n18162), .dout(n18165));
    jdff dff_B_S0g0nGY06_2(.din(n18165), .dout(n18168));
    jdff dff_B_3MpBENIv7_2(.din(n18168), .dout(n18171));
    jdff dff_B_wtFYxcyM4_2(.din(n18171), .dout(n18174));
    jdff dff_B_AV4j1lCr9_2(.din(n18174), .dout(n18177));
    jdff dff_B_ppbbj4CA7_2(.din(n18177), .dout(n18180));
    jdff dff_B_CgPF2nQd7_2(.din(n18180), .dout(n18183));
    jdff dff_B_zHiCCIu05_2(.din(n18183), .dout(n18186));
    jdff dff_B_LfNVZFHD4_2(.din(n18186), .dout(n18189));
    jdff dff_B_3PL62WaT2_2(.din(n18189), .dout(n18192));
    jdff dff_B_ZSbUGnJW2_2(.din(n18192), .dout(n18195));
    jdff dff_B_pWWTM2Y27_2(.din(n18195), .dout(n18198));
    jdff dff_B_Al4mrGMr3_2(.din(n18198), .dout(n18201));
    jdff dff_B_6nyFcD707_2(.din(n18201), .dout(n18204));
    jdff dff_B_hcK1CvGR3_2(.din(n18204), .dout(n18207));
    jdff dff_B_EzUzla1W5_2(.din(n18207), .dout(n18210));
    jdff dff_B_FmlE7YQ12_2(.din(n18210), .dout(n18213));
    jdff dff_B_zAg5CuoL4_2(.din(n18213), .dout(n18216));
    jdff dff_B_cHCEvE6K0_2(.din(n18216), .dout(n18219));
    jdff dff_B_hiXhoUJe8_2(.din(n18219), .dout(n18222));
    jdff dff_B_GAIlJRWL5_2(.din(n18222), .dout(n18225));
    jdff dff_B_yxORPfpV4_2(.din(n18225), .dout(n18228));
    jdff dff_B_kFtO13Jo8_2(.din(n4019), .dout(n18231));
    jdff dff_B_h5RKjoXL7_1(.din(n3741), .dout(n18234));
    jdff dff_B_NnjAGsoU7_2(.din(n3357), .dout(n18237));
    jdff dff_B_LYVkxd7D5_2(.din(n18237), .dout(n18240));
    jdff dff_B_VmWTAZtv4_2(.din(n18240), .dout(n18243));
    jdff dff_B_tnMALOZq3_2(.din(n18243), .dout(n18246));
    jdff dff_B_d7bR3JMp8_2(.din(n18246), .dout(n18249));
    jdff dff_B_ruUHm3AQ6_2(.din(n18249), .dout(n18252));
    jdff dff_B_TC4EuuNo9_2(.din(n18252), .dout(n18255));
    jdff dff_B_yM2L6Mdt9_2(.din(n18255), .dout(n18258));
    jdff dff_B_0IPI0RnW8_2(.din(n18258), .dout(n18261));
    jdff dff_B_Q3q1zVDc1_2(.din(n18261), .dout(n18264));
    jdff dff_B_bI9xB2bZ9_2(.din(n18264), .dout(n18267));
    jdff dff_B_TjPZ7ovH1_2(.din(n18267), .dout(n18270));
    jdff dff_B_Lm9FGTjR5_2(.din(n18270), .dout(n18273));
    jdff dff_B_tZNQvoH75_2(.din(n18273), .dout(n18276));
    jdff dff_B_4pJm1sHH8_2(.din(n18276), .dout(n18279));
    jdff dff_B_H4pbYAZF2_2(.din(n18279), .dout(n18282));
    jdff dff_B_sVdGHBeJ4_2(.din(n18282), .dout(n18285));
    jdff dff_B_so5KxBVc1_2(.din(n18285), .dout(n18288));
    jdff dff_B_OLx5nN6y6_2(.din(n18288), .dout(n18291));
    jdff dff_B_A6cRI4CC0_2(.din(n18291), .dout(n18294));
    jdff dff_B_H5aKrbt48_2(.din(n18294), .dout(n18297));
    jdff dff_B_tQKB44Qv3_2(.din(n18297), .dout(n18300));
    jdff dff_B_cFMP2liM2_2(.din(n18300), .dout(n18303));
    jdff dff_B_mAIyepEz8_2(.din(n18303), .dout(n18306));
    jdff dff_B_kTr9xOqP9_2(.din(n18306), .dout(n18309));
    jdff dff_B_vCH8Yl6s0_2(.din(n18309), .dout(n18312));
    jdff dff_B_zXluw1Pn2_2(.din(n18312), .dout(n18315));
    jdff dff_B_9colIbKg8_2(.din(n18315), .dout(n18318));
    jdff dff_B_ZAZGKhV92_2(.din(n18318), .dout(n18321));
    jdff dff_B_cPn2rPyx0_2(.din(n18321), .dout(n18324));
    jdff dff_B_cn1O666u4_2(.din(n18324), .dout(n18327));
    jdff dff_B_41p4QyuJ8_2(.din(n18327), .dout(n18330));
    jdff dff_B_uKmEUj662_2(.din(n18330), .dout(n18333));
    jdff dff_B_ZU10pe9H4_2(.din(n3636), .dout(n18336));
    jdff dff_B_btAzBAx92_1(.din(n3361), .dout(n18339));
    jdff dff_B_VfH5eDLA1_2(.din(n2966), .dout(n18342));
    jdff dff_B_oaqYiaht3_2(.din(n18342), .dout(n18345));
    jdff dff_B_0yXjSoOC4_2(.din(n18345), .dout(n18348));
    jdff dff_B_0M9xiurG3_2(.din(n18348), .dout(n18351));
    jdff dff_B_NHpPM4v32_2(.din(n18351), .dout(n18354));
    jdff dff_B_tOnSlKTU0_2(.din(n18354), .dout(n18357));
    jdff dff_B_2ODDkCKI1_2(.din(n18357), .dout(n18360));
    jdff dff_B_joaL3qXE0_2(.din(n18360), .dout(n18363));
    jdff dff_B_CLQvEiQE2_2(.din(n18363), .dout(n18366));
    jdff dff_B_jDHRomNs2_2(.din(n18366), .dout(n18369));
    jdff dff_B_gUogtGF26_2(.din(n18369), .dout(n18372));
    jdff dff_B_OQVanudn7_2(.din(n18372), .dout(n18375));
    jdff dff_B_6SX5KmRQ8_2(.din(n18375), .dout(n18378));
    jdff dff_B_yzV2Or5e4_2(.din(n18378), .dout(n18381));
    jdff dff_B_tvV6kvBu0_2(.din(n18381), .dout(n18384));
    jdff dff_B_5K8zSqgW8_2(.din(n18384), .dout(n18387));
    jdff dff_B_kxCncmAs0_2(.din(n18387), .dout(n18390));
    jdff dff_B_Ag3YV6zH0_2(.din(n18390), .dout(n18393));
    jdff dff_B_PlsJUzfM3_2(.din(n18393), .dout(n18396));
    jdff dff_B_l2dIo4kx2_2(.din(n18396), .dout(n18399));
    jdff dff_B_U0akR9E61_2(.din(n18399), .dout(n18402));
    jdff dff_B_NNCM58xX8_2(.din(n18402), .dout(n18405));
    jdff dff_B_oixyRztc2_2(.din(n18405), .dout(n18408));
    jdff dff_B_OXM9SkIO4_2(.din(n18408), .dout(n18411));
    jdff dff_B_oC5ZLoHu2_2(.din(n18411), .dout(n18414));
    jdff dff_B_mOPvEqd12_2(.din(n18414), .dout(n18417));
    jdff dff_B_zUZlpJFU2_2(.din(n18417), .dout(n18420));
    jdff dff_B_5ICvawnu0_2(.din(n18420), .dout(n18423));
    jdff dff_B_aBYRBPMW7_2(.din(n18423), .dout(n18426));
    jdff dff_B_l0x3636S9_2(.din(n18426), .dout(n18429));
    jdff dff_B_8D3wYtpI7_2(.din(n3231), .dout(n18432));
    jdff dff_B_njc17Ywt8_1(.din(n2970), .dout(n18435));
    jdff dff_B_6cC8yWm12_2(.din(n2591), .dout(n18438));
    jdff dff_B_plZlpx0s6_2(.din(n18438), .dout(n18441));
    jdff dff_B_xb8gVmEt6_2(.din(n18441), .dout(n18444));
    jdff dff_B_w5Xido9G2_2(.din(n18444), .dout(n18447));
    jdff dff_B_HOPuzNZf5_2(.din(n18447), .dout(n18450));
    jdff dff_B_Qvz7TyA18_2(.din(n18450), .dout(n18453));
    jdff dff_B_wuIZJW1W9_2(.din(n18453), .dout(n18456));
    jdff dff_B_bvELdRvx3_2(.din(n18456), .dout(n18459));
    jdff dff_B_ceOTJzh47_2(.din(n18459), .dout(n18462));
    jdff dff_B_TKpfZjDq6_2(.din(n18462), .dout(n18465));
    jdff dff_B_WuACwFQS9_2(.din(n18465), .dout(n18468));
    jdff dff_B_tx0XA0783_2(.din(n18468), .dout(n18471));
    jdff dff_B_NWz40CIk0_2(.din(n18471), .dout(n18474));
    jdff dff_B_vIFXtAW55_2(.din(n18474), .dout(n18477));
    jdff dff_B_bzFWu4ny1_2(.din(n18477), .dout(n18480));
    jdff dff_B_75wCUuzk0_2(.din(n18480), .dout(n18483));
    jdff dff_B_tfdl6AfL5_2(.din(n18483), .dout(n18486));
    jdff dff_B_YZpG7Fea5_2(.din(n18486), .dout(n18489));
    jdff dff_B_LaH0a9xn0_2(.din(n18489), .dout(n18492));
    jdff dff_B_UJ4MCAKo1_2(.din(n18492), .dout(n18495));
    jdff dff_B_fOYjXp3i4_2(.din(n18495), .dout(n18498));
    jdff dff_B_vJoXqYFp8_2(.din(n18498), .dout(n18501));
    jdff dff_B_g2y8LwN22_2(.din(n18501), .dout(n18504));
    jdff dff_B_i2MIQDRW4_2(.din(n18504), .dout(n18507));
    jdff dff_B_NIJGMWC59_2(.din(n18507), .dout(n18510));
    jdff dff_B_51UgwMD87_2(.din(n18510), .dout(n18513));
    jdff dff_B_uISdzOLI9_2(.din(n18513), .dout(n18516));
    jdff dff_B_xUzkRPVC2_2(.din(n2836), .dout(n18519));
    jdff dff_B_xlYWbEmV9_1(.din(n2595), .dout(n18522));
    jdff dff_B_pt8vCAy86_2(.din(n2240), .dout(n18525));
    jdff dff_B_s5txgLny6_2(.din(n18525), .dout(n18528));
    jdff dff_B_t4oyNgGK6_2(.din(n18528), .dout(n18531));
    jdff dff_B_yTAOYG8R6_2(.din(n18531), .dout(n18534));
    jdff dff_B_qt64Ig8W3_2(.din(n18534), .dout(n18537));
    jdff dff_B_2Eme1FDV3_2(.din(n18537), .dout(n18540));
    jdff dff_B_6tjTP7AH4_2(.din(n18540), .dout(n18543));
    jdff dff_B_9RCxY58A2_2(.din(n18543), .dout(n18546));
    jdff dff_B_aTQZ94k94_2(.din(n18546), .dout(n18549));
    jdff dff_B_sJyoePeo2_2(.din(n18549), .dout(n18552));
    jdff dff_B_ImeqOoTv9_2(.din(n18552), .dout(n18555));
    jdff dff_B_1Itl3AOh3_2(.din(n18555), .dout(n18558));
    jdff dff_B_mZbG4vqC8_2(.din(n18558), .dout(n18561));
    jdff dff_B_rSfylnvx7_2(.din(n18561), .dout(n18564));
    jdff dff_B_m61EIGg49_2(.din(n18564), .dout(n18567));
    jdff dff_B_MqoDtEPs3_2(.din(n18567), .dout(n18570));
    jdff dff_B_2MiqQLhx2_2(.din(n18570), .dout(n18573));
    jdff dff_B_1Gyz0rPC4_2(.din(n18573), .dout(n18576));
    jdff dff_B_FiWusDru0_2(.din(n18576), .dout(n18579));
    jdff dff_B_slO8bQ4h7_2(.din(n18579), .dout(n18582));
    jdff dff_B_7A5LtFVb7_2(.din(n18582), .dout(n18585));
    jdff dff_B_rKjJMvQ06_2(.din(n18585), .dout(n18588));
    jdff dff_B_hZEEUm4Y3_2(.din(n18588), .dout(n18591));
    jdff dff_B_5DMS3Dqa4_2(.din(n18591), .dout(n18594));
    jdff dff_B_cHYOWHXB5_2(.din(n2458), .dout(n18597));
    jdff dff_B_zA1fVh209_1(.din(n2244), .dout(n18600));
    jdff dff_B_1TX4ygRy1_2(.din(n1916), .dout(n18603));
    jdff dff_B_2Ap0Oqjh9_2(.din(n18603), .dout(n18606));
    jdff dff_B_fy72smUI6_2(.din(n18606), .dout(n18609));
    jdff dff_B_v6yxoG7W3_2(.din(n18609), .dout(n18612));
    jdff dff_B_9xjHvdEt9_2(.din(n18612), .dout(n18615));
    jdff dff_B_Pcfv2wn50_2(.din(n18615), .dout(n18618));
    jdff dff_B_XPrzWFuJ1_2(.din(n18618), .dout(n18621));
    jdff dff_B_jWl5kXsp0_2(.din(n18621), .dout(n18624));
    jdff dff_B_dgaqfbzw1_2(.din(n18624), .dout(n18627));
    jdff dff_B_moLpdjUd3_2(.din(n18627), .dout(n18630));
    jdff dff_B_yKpLB11R7_2(.din(n18630), .dout(n18633));
    jdff dff_B_Lcg9y8Rs8_2(.din(n18633), .dout(n18636));
    jdff dff_B_dYU88pkw3_2(.din(n18636), .dout(n18639));
    jdff dff_B_jAOlGQVv3_2(.din(n18639), .dout(n18642));
    jdff dff_B_anPlZ8127_2(.din(n18642), .dout(n18645));
    jdff dff_B_GHpfCaqR4_2(.din(n18645), .dout(n18648));
    jdff dff_B_RLwUrAon2_2(.din(n18648), .dout(n18651));
    jdff dff_B_stLmgViI4_2(.din(n18651), .dout(n18654));
    jdff dff_B_N3kdYXo48_2(.din(n18654), .dout(n18657));
    jdff dff_B_MgyIN9sG8_2(.din(n18657), .dout(n18660));
    jdff dff_B_EPOCiutL4_2(.din(n18660), .dout(n18663));
    jdff dff_B_EnMmaieR2_2(.din(n2107), .dout(n18666));
    jdff dff_B_5tQ7JrXv8_1(.din(n1920), .dout(n18669));
    jdff dff_B_unxCXfma1_2(.din(n1619), .dout(n18672));
    jdff dff_B_DP6qr3E65_2(.din(n18672), .dout(n18675));
    jdff dff_B_8WCx9P2a0_2(.din(n18675), .dout(n18678));
    jdff dff_B_s9KaS7nA7_2(.din(n18678), .dout(n18681));
    jdff dff_B_Qk2RJZfU0_2(.din(n18681), .dout(n18684));
    jdff dff_B_HucCc95M5_2(.din(n18684), .dout(n18687));
    jdff dff_B_aEXFm0rz2_2(.din(n18687), .dout(n18690));
    jdff dff_B_8bl8lquq5_2(.din(n18690), .dout(n18693));
    jdff dff_B_Yhzy4Ndu3_2(.din(n18693), .dout(n18696));
    jdff dff_B_njnJNp6A2_2(.din(n18696), .dout(n18699));
    jdff dff_B_cS8zJBEm8_2(.din(n18699), .dout(n18702));
    jdff dff_B_5CUOBbrJ7_2(.din(n18702), .dout(n18705));
    jdff dff_B_HqXxARjb4_2(.din(n18705), .dout(n18708));
    jdff dff_B_xOSps5fC8_2(.din(n18708), .dout(n18711));
    jdff dff_B_iZ8ykPvT0_2(.din(n18711), .dout(n18714));
    jdff dff_B_2ZKYKSsb9_2(.din(n18714), .dout(n18717));
    jdff dff_B_tsuREzKB2_2(.din(n18717), .dout(n18720));
    jdff dff_B_4CxapzYz1_2(.din(n18720), .dout(n18723));
    jdff dff_B_4qBsAPLP7_2(.din(n1783), .dout(n18726));
    jdff dff_B_OJBqW99N0_1(.din(n1623), .dout(n18729));
    jdff dff_B_8TiqfJm83_2(.din(n1349), .dout(n18732));
    jdff dff_B_spq7FsAY6_2(.din(n18732), .dout(n18735));
    jdff dff_B_iU8hxj5e1_2(.din(n18735), .dout(n18738));
    jdff dff_B_PoU6hK8L2_2(.din(n18738), .dout(n18741));
    jdff dff_B_YEs4TTuI8_2(.din(n18741), .dout(n18744));
    jdff dff_B_aKduiEst8_2(.din(n18744), .dout(n18747));
    jdff dff_B_4qvfDN7q2_2(.din(n18747), .dout(n18750));
    jdff dff_B_8hgihRAU9_2(.din(n18750), .dout(n18753));
    jdff dff_B_1GD3gS9O6_2(.din(n18753), .dout(n18756));
    jdff dff_B_EOP7VZoZ8_2(.din(n18756), .dout(n18759));
    jdff dff_B_lovxccja4_2(.din(n18759), .dout(n18762));
    jdff dff_B_itFyY2Vu1_2(.din(n18762), .dout(n18765));
    jdff dff_B_gQntoKex1_2(.din(n18765), .dout(n18768));
    jdff dff_B_9hBpI5fz1_2(.din(n18768), .dout(n18771));
    jdff dff_B_BS4fxE5g2_2(.din(n18771), .dout(n18774));
    jdff dff_B_r0V17XPo8_2(.din(n1486), .dout(n18777));
    jdff dff_B_SU23IKnx1_1(.din(n1353), .dout(n18780));
    jdff dff_B_Qg4SlNPd6_2(.din(n1109), .dout(n18783));
    jdff dff_B_mZfea7FP3_2(.din(n18783), .dout(n18786));
    jdff dff_B_Cq93G2qv7_2(.din(n18786), .dout(n18789));
    jdff dff_B_kpgUEfDk0_2(.din(n18789), .dout(n18792));
    jdff dff_B_Kfx9Yzom1_2(.din(n18792), .dout(n18795));
    jdff dff_B_FE3Gv6zn0_2(.din(n18795), .dout(n18798));
    jdff dff_B_zx2YoD5R1_2(.din(n18798), .dout(n18801));
    jdff dff_B_DxyAWonr9_2(.din(n18801), .dout(n18804));
    jdff dff_B_elgOHi1A7_2(.din(n18804), .dout(n18807));
    jdff dff_B_Hm7V5PC60_2(.din(n18807), .dout(n18810));
    jdff dff_B_cbYwfaWm6_2(.din(n18810), .dout(n18813));
    jdff dff_B_aXqrKbzR6_2(.din(n18813), .dout(n18816));
    jdff dff_B_wdsUzH4j4_2(.din(n1216), .dout(n18819));
    jdff dff_B_7jaHZNBo7_1(.din(n1113), .dout(n18822));
    jdff dff_B_7DToSdmf9_2(.din(n896), .dout(n18825));
    jdff dff_B_M4yhwTvW1_2(.din(n18825), .dout(n18828));
    jdff dff_B_lcqc8b7C2_2(.din(n18828), .dout(n18831));
    jdff dff_B_epfj3P5X7_2(.din(n18831), .dout(n18834));
    jdff dff_B_MansYrIu4_2(.din(n18834), .dout(n18837));
    jdff dff_B_EQiZtGhV6_2(.din(n18837), .dout(n18840));
    jdff dff_B_AdXqyWo67_2(.din(n18840), .dout(n18843));
    jdff dff_B_JKAZmDuY8_2(.din(n18843), .dout(n18846));
    jdff dff_B_vjmx9RdH1_2(.din(n18846), .dout(n18849));
    jdff dff_B_waBKwR1N6_2(.din(n976), .dout(n18852));
    jdff dff_B_bwQLdsF85_1(.din(n900), .dout(n18855));
    jdff dff_B_rWS67cWL3_2(.din(n710), .dout(n18858));
    jdff dff_B_eJtv3WUt9_2(.din(n18858), .dout(n18861));
    jdff dff_B_cYqClYIx4_2(.din(n18861), .dout(n18864));
    jdff dff_B_CV3Uu8y61_2(.din(n18864), .dout(n18867));
    jdff dff_B_atcqW1Xi4_2(.din(n18867), .dout(n18870));
    jdff dff_B_MLy6fGzE4_2(.din(n18870), .dout(n18873));
    jdff dff_B_NTfgZDis7_2(.din(n763), .dout(n18876));
    jdff dff_B_pD4IhY2h2_2(.din(n554), .dout(n18879));
    jdff dff_B_vgbS1Rp80_2(.din(n18879), .dout(n18882));
    jdff dff_B_cj34X8qx6_2(.din(n18882), .dout(n18885));
    jdff dff_B_Bo96JeWH4_0(.din(n573), .dout(n18888));
    jdff dff_A_9FnJfSj86_0(.din(n18893), .dout(n18890));
    jdff dff_A_0Gfv49f07_0(.din(n414), .dout(n18893));
    jdff dff_A_bfPU2Rw02_0(.din(n18899), .dout(n18896));
    jdff dff_A_NFpSeRGc1_0(.din(n411), .dout(n18899));
    jdff dff_B_82kEDmpO3_2(.din(n5122), .dout(n18903));
    jdff dff_B_p8CFYD8r0_1(.din(n5114), .dout(n18906));
    jdff dff_B_HI0qfoCK6_2(.din(n4808), .dout(n18909));
    jdff dff_B_w73QtY3Q9_2(.din(n18909), .dout(n18912));
    jdff dff_B_LNYBxVAH7_2(.din(n18912), .dout(n18915));
    jdff dff_B_lPzsAtnl1_2(.din(n18915), .dout(n18918));
    jdff dff_B_i6rbg7Gh2_2(.din(n18918), .dout(n18921));
    jdff dff_B_H2vf3QHQ9_2(.din(n18921), .dout(n18924));
    jdff dff_B_644zwNW39_2(.din(n18924), .dout(n18927));
    jdff dff_B_AUHmEi0s6_2(.din(n18927), .dout(n18930));
    jdff dff_B_0XDnDoZu7_2(.din(n18930), .dout(n18933));
    jdff dff_B_GWh1cxgr8_2(.din(n18933), .dout(n18936));
    jdff dff_B_Mc1DBr5L5_2(.din(n18936), .dout(n18939));
    jdff dff_B_OaBZf7ZE6_2(.din(n18939), .dout(n18942));
    jdff dff_B_58AJcBXl5_2(.din(n18942), .dout(n18945));
    jdff dff_B_5tmlsUO70_2(.din(n18945), .dout(n18948));
    jdff dff_B_Tmk9yV9w1_2(.din(n18948), .dout(n18951));
    jdff dff_B_WdOXA5mO3_2(.din(n18951), .dout(n18954));
    jdff dff_B_Zs0lAgYe5_2(.din(n18954), .dout(n18957));
    jdff dff_B_ZBSGuona0_2(.din(n18957), .dout(n18960));
    jdff dff_B_DSnE9pEi0_2(.din(n18960), .dout(n18963));
    jdff dff_B_N3MGM5NK5_2(.din(n18963), .dout(n18966));
    jdff dff_B_0QJHOML52_2(.din(n18966), .dout(n18969));
    jdff dff_B_DAQtcvhJ1_2(.din(n18969), .dout(n18972));
    jdff dff_B_JhCNHU203_2(.din(n18972), .dout(n18975));
    jdff dff_B_iPkvAayr1_2(.din(n18975), .dout(n18978));
    jdff dff_B_yIxlhDMw1_2(.din(n18978), .dout(n18981));
    jdff dff_B_ANWPsLnT1_2(.din(n18981), .dout(n18984));
    jdff dff_B_8OEexEgb5_2(.din(n18984), .dout(n18987));
    jdff dff_B_PX4UNlqr5_2(.din(n18987), .dout(n18990));
    jdff dff_B_oa0pRPl03_2(.din(n18990), .dout(n18993));
    jdff dff_B_FibqFtvc0_2(.din(n18993), .dout(n18996));
    jdff dff_B_zzVScD3D7_2(.din(n18996), .dout(n18999));
    jdff dff_B_luxOHkko4_2(.din(n18999), .dout(n19002));
    jdff dff_B_yfR7hewW4_2(.din(n19002), .dout(n19005));
    jdff dff_B_jRtBBDC25_2(.din(n19005), .dout(n19008));
    jdff dff_B_WxJYm7pB9_2(.din(n19008), .dout(n19011));
    jdff dff_B_uMKWbvTc7_2(.din(n19011), .dout(n19014));
    jdff dff_B_CvaJ2SY51_2(.din(n19014), .dout(n19017));
    jdff dff_B_FmLZ3YRa6_2(.din(n19017), .dout(n19020));
    jdff dff_B_obwItojH0_2(.din(n19020), .dout(n19023));
    jdff dff_B_bC6drbKZ5_2(.din(n19023), .dout(n19026));
    jdff dff_B_2xx4hGKK8_2(.din(n19026), .dout(n19029));
    jdff dff_B_78y7PVT11_2(.din(n19029), .dout(n19032));
    jdff dff_B_SmH6ODnO9_2(.din(n19032), .dout(n19035));
    jdff dff_B_RRUhEdFG0_2(.din(n19035), .dout(n19038));
    jdff dff_B_8gNLrgrL5_1(.din(n4812), .dout(n19041));
    jdff dff_B_EGvTs1xQ9_2(.din(n4482), .dout(n19044));
    jdff dff_B_vmsMTtn00_2(.din(n19044), .dout(n19047));
    jdff dff_B_Zzdhxzqe1_2(.din(n19047), .dout(n19050));
    jdff dff_B_r0mzhX8g9_2(.din(n19050), .dout(n19053));
    jdff dff_B_ABwxiugB5_2(.din(n19053), .dout(n19056));
    jdff dff_B_QmTSpFZp3_2(.din(n19056), .dout(n19059));
    jdff dff_B_FWRpa9tG3_2(.din(n19059), .dout(n19062));
    jdff dff_B_CuoKJ7Sx5_2(.din(n19062), .dout(n19065));
    jdff dff_B_WowdH8jj9_2(.din(n19065), .dout(n19068));
    jdff dff_B_fSLnroM98_2(.din(n19068), .dout(n19071));
    jdff dff_B_SDYmAZBe9_2(.din(n19071), .dout(n19074));
    jdff dff_B_CnjXIl4S1_2(.din(n19074), .dout(n19077));
    jdff dff_B_RTL4yCjC8_2(.din(n19077), .dout(n19080));
    jdff dff_B_YEiyUClY1_2(.din(n19080), .dout(n19083));
    jdff dff_B_M6m0kAGz4_2(.din(n19083), .dout(n19086));
    jdff dff_B_RNWrOxw22_2(.din(n19086), .dout(n19089));
    jdff dff_B_VZj7Jbbp9_2(.din(n19089), .dout(n19092));
    jdff dff_B_gL287Ds75_2(.din(n19092), .dout(n19095));
    jdff dff_B_noyylPMX4_2(.din(n19095), .dout(n19098));
    jdff dff_B_GUT3ncYz4_2(.din(n19098), .dout(n19101));
    jdff dff_B_Qye8awiK7_2(.din(n19101), .dout(n19104));
    jdff dff_B_O7kn2KFC2_2(.din(n19104), .dout(n19107));
    jdff dff_B_xaYz8JMU4_2(.din(n19107), .dout(n19110));
    jdff dff_B_QzuES2Gt2_2(.din(n19110), .dout(n19113));
    jdff dff_B_frUWt0if3_2(.din(n19113), .dout(n19116));
    jdff dff_B_gPjMMraJ6_2(.din(n19116), .dout(n19119));
    jdff dff_B_rQAbOnRM8_2(.din(n19119), .dout(n19122));
    jdff dff_B_iTUhyJ955_2(.din(n19122), .dout(n19125));
    jdff dff_B_gO1OiREC7_2(.din(n19125), .dout(n19128));
    jdff dff_B_GI2S4c4N1_2(.din(n19128), .dout(n19131));
    jdff dff_B_PbHefd6e7_2(.din(n19131), .dout(n19134));
    jdff dff_B_20oLcZmG6_2(.din(n19134), .dout(n19137));
    jdff dff_B_xMYI3rRT2_2(.din(n19137), .dout(n19140));
    jdff dff_B_CSBp4CcL0_2(.din(n19140), .dout(n19143));
    jdff dff_B_k0b7nD5x0_2(.din(n19143), .dout(n19146));
    jdff dff_B_odrsetPv7_2(.din(n19146), .dout(n19149));
    jdff dff_B_CWleIVRD5_2(.din(n19149), .dout(n19152));
    jdff dff_B_ZrBCp82e3_2(.din(n19152), .dout(n19155));
    jdff dff_B_kISjt9Nd0_2(.din(n19155), .dout(n19158));
    jdff dff_B_6d1qojQz1_1(.din(n4486), .dout(n19161));
    jdff dff_B_arPmkPW94_2(.din(n4132), .dout(n19164));
    jdff dff_B_eYb4nYSB6_2(.din(n19164), .dout(n19167));
    jdff dff_B_UA0qZu8p6_2(.din(n19167), .dout(n19170));
    jdff dff_B_ycShQNNf1_2(.din(n19170), .dout(n19173));
    jdff dff_B_vwywIjc38_2(.din(n19173), .dout(n19176));
    jdff dff_B_at1gFTkX8_2(.din(n19176), .dout(n19179));
    jdff dff_B_cmhlqIXG9_2(.din(n19179), .dout(n19182));
    jdff dff_B_pISZsA3N8_2(.din(n19182), .dout(n19185));
    jdff dff_B_mMikUdx37_2(.din(n19185), .dout(n19188));
    jdff dff_B_QLYrlFXX6_2(.din(n19188), .dout(n19191));
    jdff dff_B_jHcBvwUM4_2(.din(n19191), .dout(n19194));
    jdff dff_B_1QeLrvrj9_2(.din(n19194), .dout(n19197));
    jdff dff_B_y537y5px3_2(.din(n19197), .dout(n19200));
    jdff dff_B_7EOGJAyi0_2(.din(n19200), .dout(n19203));
    jdff dff_B_SRZiTzNW4_2(.din(n19203), .dout(n19206));
    jdff dff_B_BBsEUafp8_2(.din(n19206), .dout(n19209));
    jdff dff_B_SuLWa2X11_2(.din(n19209), .dout(n19212));
    jdff dff_B_N1fq99Ep3_2(.din(n19212), .dout(n19215));
    jdff dff_B_LbBO6qaN2_2(.din(n19215), .dout(n19218));
    jdff dff_B_TyOotS5b3_2(.din(n19218), .dout(n19221));
    jdff dff_B_sG5fA6rP3_2(.din(n19221), .dout(n19224));
    jdff dff_B_9Mr5x8V88_2(.din(n19224), .dout(n19227));
    jdff dff_B_5rC9Sz629_2(.din(n19227), .dout(n19230));
    jdff dff_B_2XOD3RCs5_2(.din(n19230), .dout(n19233));
    jdff dff_B_iUV9ddRP3_2(.din(n19233), .dout(n19236));
    jdff dff_B_lmhbLABn6_2(.din(n19236), .dout(n19239));
    jdff dff_B_gd9OMT3T3_2(.din(n19239), .dout(n19242));
    jdff dff_B_LDYzMncT7_2(.din(n19242), .dout(n19245));
    jdff dff_B_kP9rWVYB7_2(.din(n19245), .dout(n19248));
    jdff dff_B_0lC176QA7_2(.din(n19248), .dout(n19251));
    jdff dff_B_hQAH83qA2_2(.din(n19251), .dout(n19254));
    jdff dff_B_kq3TksPn3_2(.din(n19254), .dout(n19257));
    jdff dff_B_9RGTEren2_2(.din(n19257), .dout(n19260));
    jdff dff_B_eo8HzTsY9_2(.din(n19260), .dout(n19263));
    jdff dff_B_vCCULbSY1_2(.din(n19263), .dout(n19266));
    jdff dff_B_K4Sn2Y1Z6_2(.din(n19266), .dout(n19269));
    jdff dff_B_LiVhcqFl1_1(.din(n4136), .dout(n19272));
    jdff dff_B_5T1BUQmj0_2(.din(n3756), .dout(n19275));
    jdff dff_B_6hDLsMDT8_2(.din(n19275), .dout(n19278));
    jdff dff_B_sA8hbA520_2(.din(n19278), .dout(n19281));
    jdff dff_B_THETvd4u5_2(.din(n19281), .dout(n19284));
    jdff dff_B_VxDt8xz84_2(.din(n19284), .dout(n19287));
    jdff dff_B_xFbP1kHF3_2(.din(n19287), .dout(n19290));
    jdff dff_B_silobUlP7_2(.din(n19290), .dout(n19293));
    jdff dff_B_0jBhBDnc6_2(.din(n19293), .dout(n19296));
    jdff dff_B_04O1bZi03_2(.din(n19296), .dout(n19299));
    jdff dff_B_t02yxgQk1_2(.din(n19299), .dout(n19302));
    jdff dff_B_MewjG7D89_2(.din(n19302), .dout(n19305));
    jdff dff_B_dFCn7i5V6_2(.din(n19305), .dout(n19308));
    jdff dff_B_aVcUdzfJ1_2(.din(n19308), .dout(n19311));
    jdff dff_B_5CNxMRfU1_2(.din(n19311), .dout(n19314));
    jdff dff_B_cFdAtfq98_2(.din(n19314), .dout(n19317));
    jdff dff_B_CqDelUtY8_2(.din(n19317), .dout(n19320));
    jdff dff_B_HN26A4Ni0_2(.din(n19320), .dout(n19323));
    jdff dff_B_ESmp7wAC2_2(.din(n19323), .dout(n19326));
    jdff dff_B_6SQQFuWk0_2(.din(n19326), .dout(n19329));
    jdff dff_B_ZdHZhSpi1_2(.din(n19329), .dout(n19332));
    jdff dff_B_ydtLEszk5_2(.din(n19332), .dout(n19335));
    jdff dff_B_yJlNFCTq1_2(.din(n19335), .dout(n19338));
    jdff dff_B_T9STk5IL3_2(.din(n19338), .dout(n19341));
    jdff dff_B_jr5fRvJ45_2(.din(n19341), .dout(n19344));
    jdff dff_B_EdQo7zSe0_2(.din(n19344), .dout(n19347));
    jdff dff_B_GCfu9r2u5_2(.din(n19347), .dout(n19350));
    jdff dff_B_GbPeGblU3_2(.din(n19350), .dout(n19353));
    jdff dff_B_ETSuWgpd3_2(.din(n19353), .dout(n19356));
    jdff dff_B_BBvFPJw66_2(.din(n19356), .dout(n19359));
    jdff dff_B_ZkoKZYV51_2(.din(n19359), .dout(n19362));
    jdff dff_B_Tv3gA1nG5_2(.din(n19362), .dout(n19365));
    jdff dff_B_ExnYwyxT1_2(.din(n19365), .dout(n19368));
    jdff dff_B_bJ48C7vN1_2(.din(n19368), .dout(n19371));
    jdff dff_B_TOvxfCyx5_1(.din(n3760), .dout(n19374));
    jdff dff_B_OOBUTOR80_2(.din(n3376), .dout(n19377));
    jdff dff_B_D8hCKFkA6_2(.din(n19377), .dout(n19380));
    jdff dff_B_b1EnRnaB3_2(.din(n19380), .dout(n19383));
    jdff dff_B_BXIPDdgF9_2(.din(n19383), .dout(n19386));
    jdff dff_B_v2VkihFM1_2(.din(n19386), .dout(n19389));
    jdff dff_B_AVv2Zxrm7_2(.din(n19389), .dout(n19392));
    jdff dff_B_MH4fLmfQ2_2(.din(n19392), .dout(n19395));
    jdff dff_B_fPbrqTmk8_2(.din(n19395), .dout(n19398));
    jdff dff_B_jT1SUDCg2_2(.din(n19398), .dout(n19401));
    jdff dff_B_WKMyKDQw5_2(.din(n19401), .dout(n19404));
    jdff dff_B_mJQtkapL5_2(.din(n19404), .dout(n19407));
    jdff dff_B_1MfXvMZP2_2(.din(n19407), .dout(n19410));
    jdff dff_B_9DHT5X8f3_2(.din(n19410), .dout(n19413));
    jdff dff_B_351IfMQB1_2(.din(n19413), .dout(n19416));
    jdff dff_B_y4NHOxFn7_2(.din(n19416), .dout(n19419));
    jdff dff_B_YPCthopJ1_2(.din(n19419), .dout(n19422));
    jdff dff_B_4awknyCS9_2(.din(n19422), .dout(n19425));
    jdff dff_B_DWLC9RBZ3_2(.din(n19425), .dout(n19428));
    jdff dff_B_OqWSA1Nw7_2(.din(n19428), .dout(n19431));
    jdff dff_B_gCtn49xw4_2(.din(n19431), .dout(n19434));
    jdff dff_B_Pi0nXxgR0_2(.din(n19434), .dout(n19437));
    jdff dff_B_8AZnS9pP3_2(.din(n19437), .dout(n19440));
    jdff dff_B_Xxba8x8E1_2(.din(n19440), .dout(n19443));
    jdff dff_B_Ehs56RKh6_2(.din(n19443), .dout(n19446));
    jdff dff_B_HD4A2ZOK1_2(.din(n19446), .dout(n19449));
    jdff dff_B_tGNUhpZH2_2(.din(n19449), .dout(n19452));
    jdff dff_B_pfjyruZ24_2(.din(n19452), .dout(n19455));
    jdff dff_B_JbvP0yVV6_2(.din(n19455), .dout(n19458));
    jdff dff_B_Ob6Fd71d9_2(.din(n19458), .dout(n19461));
    jdff dff_B_pOWat9C22_2(.din(n19461), .dout(n19464));
    jdff dff_B_3pE5dkfD9_1(.din(n3380), .dout(n19467));
    jdff dff_B_Sdv33Ges1_2(.din(n2985), .dout(n19470));
    jdff dff_B_aGtrsy8H2_2(.din(n19470), .dout(n19473));
    jdff dff_B_gwpL6CsZ7_2(.din(n19473), .dout(n19476));
    jdff dff_B_JJvg7gsc7_2(.din(n19476), .dout(n19479));
    jdff dff_B_gFquDKE14_2(.din(n19479), .dout(n19482));
    jdff dff_B_IHxtHSjZ1_2(.din(n19482), .dout(n19485));
    jdff dff_B_SP6uV0Fr4_2(.din(n19485), .dout(n19488));
    jdff dff_B_EUc7JVss8_2(.din(n19488), .dout(n19491));
    jdff dff_B_Gq3OZvl68_2(.din(n19491), .dout(n19494));
    jdff dff_B_OlSijAxY2_2(.din(n19494), .dout(n19497));
    jdff dff_B_mvxnN1Jh5_2(.din(n19497), .dout(n19500));
    jdff dff_B_7WigKAb76_2(.din(n19500), .dout(n19503));
    jdff dff_B_mOah6vMx6_2(.din(n19503), .dout(n19506));
    jdff dff_B_bv47knXu4_2(.din(n19506), .dout(n19509));
    jdff dff_B_tujRlVA13_2(.din(n19509), .dout(n19512));
    jdff dff_B_ZTTkuLQJ6_2(.din(n19512), .dout(n19515));
    jdff dff_B_EJc5b1yF0_2(.din(n19515), .dout(n19518));
    jdff dff_B_ksKWp9c14_2(.din(n19518), .dout(n19521));
    jdff dff_B_SERcjpHn4_2(.din(n19521), .dout(n19524));
    jdff dff_B_tvqRN6p74_2(.din(n19524), .dout(n19527));
    jdff dff_B_QfL4rNG06_2(.din(n19527), .dout(n19530));
    jdff dff_B_CZvNo3Yr6_2(.din(n19530), .dout(n19533));
    jdff dff_B_ucpVJGBH3_2(.din(n19533), .dout(n19536));
    jdff dff_B_toF0Zfpz7_2(.din(n19536), .dout(n19539));
    jdff dff_B_28ZkR1Dl2_2(.din(n19539), .dout(n19542));
    jdff dff_B_nS4ZgaTO2_2(.din(n19542), .dout(n19545));
    jdff dff_B_oweQ0Jal5_2(.din(n19545), .dout(n19548));
    jdff dff_B_R0z19Jep3_1(.din(n2989), .dout(n19551));
    jdff dff_B_QXRnl56v5_2(.din(n2610), .dout(n19554));
    jdff dff_B_v8ZdHMr87_2(.din(n19554), .dout(n19557));
    jdff dff_B_V1zqU0I55_2(.din(n19557), .dout(n19560));
    jdff dff_B_CisTQMR80_2(.din(n19560), .dout(n19563));
    jdff dff_B_fe4cb1eZ6_2(.din(n19563), .dout(n19566));
    jdff dff_B_ijIuYNse6_2(.din(n19566), .dout(n19569));
    jdff dff_B_566cVKcr4_2(.din(n19569), .dout(n19572));
    jdff dff_B_WqcfleWR4_2(.din(n19572), .dout(n19575));
    jdff dff_B_S3eKu4XR9_2(.din(n19575), .dout(n19578));
    jdff dff_B_pQ4tXXlM0_2(.din(n19578), .dout(n19581));
    jdff dff_B_VWJBY6Ak9_2(.din(n19581), .dout(n19584));
    jdff dff_B_144ktcIl9_2(.din(n19584), .dout(n19587));
    jdff dff_B_rTcU2Qbc6_2(.din(n19587), .dout(n19590));
    jdff dff_B_5txrRGBZ7_2(.din(n19590), .dout(n19593));
    jdff dff_B_ceTNVhgU7_2(.din(n19593), .dout(n19596));
    jdff dff_B_oM1CwD9C8_2(.din(n19596), .dout(n19599));
    jdff dff_B_FCiStozC3_2(.din(n19599), .dout(n19602));
    jdff dff_B_uCabLax15_2(.din(n19602), .dout(n19605));
    jdff dff_B_MMFxZGqu2_2(.din(n19605), .dout(n19608));
    jdff dff_B_ptfX8f457_2(.din(n19608), .dout(n19611));
    jdff dff_B_Cnn5jTTL5_2(.din(n19611), .dout(n19614));
    jdff dff_B_2ydK2cuO5_2(.din(n19614), .dout(n19617));
    jdff dff_B_ZUEycug21_2(.din(n19617), .dout(n19620));
    jdff dff_B_QgQgfMTD9_2(.din(n19620), .dout(n19623));
    jdff dff_B_y8GhzqHs6_1(.din(n2614), .dout(n19626));
    jdff dff_B_wKUwr2961_2(.din(n2259), .dout(n19629));
    jdff dff_B_cAHx3hjm3_2(.din(n19629), .dout(n19632));
    jdff dff_B_hZNCI5Hf4_2(.din(n19632), .dout(n19635));
    jdff dff_B_sP1w03i44_2(.din(n19635), .dout(n19638));
    jdff dff_B_9iWZnr7B6_2(.din(n19638), .dout(n19641));
    jdff dff_B_knllvzOm7_2(.din(n19641), .dout(n19644));
    jdff dff_B_8Ck0rVff5_2(.din(n19644), .dout(n19647));
    jdff dff_B_9gBWMI4B5_2(.din(n19647), .dout(n19650));
    jdff dff_B_rgx9td3J4_2(.din(n19650), .dout(n19653));
    jdff dff_B_WQ171XwV0_2(.din(n19653), .dout(n19656));
    jdff dff_B_dwY2m9UF3_2(.din(n19656), .dout(n19659));
    jdff dff_B_JUxIufPX6_2(.din(n19659), .dout(n19662));
    jdff dff_B_PV8T9nrb8_2(.din(n19662), .dout(n19665));
    jdff dff_B_5h6mvSNl8_2(.din(n19665), .dout(n19668));
    jdff dff_B_Ojy9qFaM2_2(.din(n19668), .dout(n19671));
    jdff dff_B_dol2pIu93_2(.din(n19671), .dout(n19674));
    jdff dff_B_FRJtNm0V9_2(.din(n19674), .dout(n19677));
    jdff dff_B_YOq2of3r1_2(.din(n19677), .dout(n19680));
    jdff dff_B_IyBLy1eD9_2(.din(n19680), .dout(n19683));
    jdff dff_B_jQaiMMzj2_2(.din(n19683), .dout(n19686));
    jdff dff_B_N8U5UmxG3_2(.din(n19686), .dout(n19689));
    jdff dff_B_tzp9z56e2_1(.din(n2263), .dout(n19692));
    jdff dff_B_jPNCXNaj2_2(.din(n1935), .dout(n19695));
    jdff dff_B_Cpi0dReh1_2(.din(n19695), .dout(n19698));
    jdff dff_B_OWU55v149_2(.din(n19698), .dout(n19701));
    jdff dff_B_wvPkt51q9_2(.din(n19701), .dout(n19704));
    jdff dff_B_3juSFDU49_2(.din(n19704), .dout(n19707));
    jdff dff_B_Lrkf98dy0_2(.din(n19707), .dout(n19710));
    jdff dff_B_yl3iKIQG4_2(.din(n19710), .dout(n19713));
    jdff dff_B_yZdKaMai2_2(.din(n19713), .dout(n19716));
    jdff dff_B_DLeQDyfQ9_2(.din(n19716), .dout(n19719));
    jdff dff_B_2bPKmKWU6_2(.din(n19719), .dout(n19722));
    jdff dff_B_GcPNPhsu4_2(.din(n19722), .dout(n19725));
    jdff dff_B_rndqwl6u4_2(.din(n19725), .dout(n19728));
    jdff dff_B_DknIx0LD7_2(.din(n19728), .dout(n19731));
    jdff dff_B_t4DhqEG94_2(.din(n19731), .dout(n19734));
    jdff dff_B_Td7YVL914_2(.din(n19734), .dout(n19737));
    jdff dff_B_mlVKHcth2_2(.din(n19737), .dout(n19740));
    jdff dff_B_GZaXYlnM9_2(.din(n19740), .dout(n19743));
    jdff dff_B_ImxTX2uV5_2(.din(n19743), .dout(n19746));
    jdff dff_B_yLerp6T52_1(.din(n1939), .dout(n19749));
    jdff dff_B_xh23TJQr8_2(.din(n1638), .dout(n19752));
    jdff dff_B_09jGHuYQ8_2(.din(n19752), .dout(n19755));
    jdff dff_B_6ejMo3wB8_2(.din(n19755), .dout(n19758));
    jdff dff_B_c5X5DqdK8_2(.din(n19758), .dout(n19761));
    jdff dff_B_HGtgy4R34_2(.din(n19761), .dout(n19764));
    jdff dff_B_yCSnzhs16_2(.din(n19764), .dout(n19767));
    jdff dff_B_SFvSsLEM0_2(.din(n19767), .dout(n19770));
    jdff dff_B_1jqv8wRl7_2(.din(n19770), .dout(n19773));
    jdff dff_B_dBRo2nOc2_2(.din(n19773), .dout(n19776));
    jdff dff_B_ZzuDrKUA1_2(.din(n19776), .dout(n19779));
    jdff dff_B_fd8RLpn81_2(.din(n19779), .dout(n19782));
    jdff dff_B_HZl9l0B42_2(.din(n19782), .dout(n19785));
    jdff dff_B_TcTb2V1f6_2(.din(n19785), .dout(n19788));
    jdff dff_B_8kyQZQZ51_2(.din(n19788), .dout(n19791));
    jdff dff_B_JfRbc5xr0_2(.din(n19791), .dout(n19794));
    jdff dff_B_AwApN28D3_1(.din(n1642), .dout(n19797));
    jdff dff_B_ui3Vok8d8_2(.din(n1368), .dout(n19800));
    jdff dff_B_rycLXFoe9_2(.din(n19800), .dout(n19803));
    jdff dff_B_BAIFFObf8_2(.din(n19803), .dout(n19806));
    jdff dff_B_i6dKyt5G1_2(.din(n19806), .dout(n19809));
    jdff dff_B_zAncI7QG6_2(.din(n19809), .dout(n19812));
    jdff dff_B_duj50ZVH5_2(.din(n19812), .dout(n19815));
    jdff dff_B_5QHiVTBT2_2(.din(n19815), .dout(n19818));
    jdff dff_B_Eli7zVJp5_2(.din(n19818), .dout(n19821));
    jdff dff_B_HuYzGv3G8_2(.din(n19821), .dout(n19824));
    jdff dff_B_vM8hH5fA0_2(.din(n19824), .dout(n19827));
    jdff dff_B_2wEY9y9G1_2(.din(n19827), .dout(n19830));
    jdff dff_B_4Ews6Nh30_2(.din(n19830), .dout(n19833));
    jdff dff_B_NBaNDCuu2_1(.din(n1372), .dout(n19836));
    jdff dff_B_em16gT3f0_2(.din(n1128), .dout(n19839));
    jdff dff_B_UhREfVy77_2(.din(n19839), .dout(n19842));
    jdff dff_B_ZGV8XdVu4_2(.din(n19842), .dout(n19845));
    jdff dff_B_FiMxoM3v3_2(.din(n19845), .dout(n19848));
    jdff dff_B_NhkCPPxv1_2(.din(n19848), .dout(n19851));
    jdff dff_B_oWJ8I7fA0_2(.din(n19851), .dout(n19854));
    jdff dff_B_U5HSUCU58_2(.din(n19854), .dout(n19857));
    jdff dff_B_RIt4nk6Q7_2(.din(n19857), .dout(n19860));
    jdff dff_B_bhrnvtsu1_2(.din(n19860), .dout(n19863));
    jdff dff_B_AZjjbSdA3_2(.din(n1208), .dout(n19866));
    jdff dff_B_vTLeOGiF5_1(.din(n1132), .dout(n19869));
    jdff dff_B_96ZCAOpF3_2(.din(n915), .dout(n19872));
    jdff dff_B_yrshsnC17_2(.din(n19872), .dout(n19875));
    jdff dff_B_9AaqN74H3_2(.din(n19875), .dout(n19878));
    jdff dff_B_Tn8aBqFA4_2(.din(n19878), .dout(n19881));
    jdff dff_B_w4EXgv7l6_2(.din(n19881), .dout(n19884));
    jdff dff_B_uIrpoRSt3_2(.din(n19884), .dout(n19887));
    jdff dff_B_008ENNDH2_2(.din(n968), .dout(n19890));
    jdff dff_B_9mLinlEm2_2(.din(n732), .dout(n19893));
    jdff dff_B_lGbCP0C67_2(.din(n19893), .dout(n19896));
    jdff dff_B_lTV9VUfa5_2(.din(n19896), .dout(n19899));
    jdff dff_B_GV8eUhdT1_0(.din(n751), .dout(n19902));
    jdff dff_A_GLXUj7kV6_0(.din(n19907), .dout(n19904));
    jdff dff_A_PJAIXXDw9_0(.din(n562), .dout(n19907));
    jdff dff_A_yrorCRtU1_1(.din(n19913), .dout(n19910));
    jdff dff_A_q9M9gnBA4_1(.din(n562), .dout(n19913));
    jdff dff_B_w8ZEJdi97_2(.din(n5413), .dout(n19917));
    jdff dff_B_3QFD0j615_1(.din(n5405), .dout(n19920));
    jdff dff_B_k2wqKZQZ9_2(.din(n5126), .dout(n19923));
    jdff dff_B_SQ3Agozi2_2(.din(n19923), .dout(n19926));
    jdff dff_B_Ub5cjh3i8_2(.din(n19926), .dout(n19929));
    jdff dff_B_5c4vqkeX8_2(.din(n19929), .dout(n19932));
    jdff dff_B_3Nuek61q6_2(.din(n19932), .dout(n19935));
    jdff dff_B_sfNeiznr8_2(.din(n19935), .dout(n19938));
    jdff dff_B_Mp7ndH4q8_2(.din(n19938), .dout(n19941));
    jdff dff_B_ArSjtfMa1_2(.din(n19941), .dout(n19944));
    jdff dff_B_wnb6lGO95_2(.din(n19944), .dout(n19947));
    jdff dff_B_x3L7vdKr0_2(.din(n19947), .dout(n19950));
    jdff dff_B_3pbMwHA09_2(.din(n19950), .dout(n19953));
    jdff dff_B_CnP5aY734_2(.din(n19953), .dout(n19956));
    jdff dff_B_StkDG3hZ3_2(.din(n19956), .dout(n19959));
    jdff dff_B_eybkSGqS9_2(.din(n19959), .dout(n19962));
    jdff dff_B_AqZy4FWR8_2(.din(n19962), .dout(n19965));
    jdff dff_B_3fuGERfV3_2(.din(n19965), .dout(n19968));
    jdff dff_B_xO7fNMXW9_2(.din(n19968), .dout(n19971));
    jdff dff_B_MPmlsFHX5_2(.din(n19971), .dout(n19974));
    jdff dff_B_QflfAzRo9_2(.din(n19974), .dout(n19977));
    jdff dff_B_IPHjuRXg6_2(.din(n19977), .dout(n19980));
    jdff dff_B_iNBJO3Iw4_2(.din(n19980), .dout(n19983));
    jdff dff_B_p1UJ8gvY2_2(.din(n19983), .dout(n19986));
    jdff dff_B_A70XKMX65_2(.din(n19986), .dout(n19989));
    jdff dff_B_xVATjQpv2_2(.din(n19989), .dout(n19992));
    jdff dff_B_FfQGHvcz9_2(.din(n19992), .dout(n19995));
    jdff dff_B_tpDpCILF9_2(.din(n19995), .dout(n19998));
    jdff dff_B_y7UBxaVe9_2(.din(n19998), .dout(n20001));
    jdff dff_B_t3zvDPvW5_2(.din(n20001), .dout(n20004));
    jdff dff_B_sdIisz9O7_2(.din(n20004), .dout(n20007));
    jdff dff_B_j20DL4N69_2(.din(n20007), .dout(n20010));
    jdff dff_B_8ay992s14_2(.din(n20010), .dout(n20013));
    jdff dff_B_0a14F5911_2(.din(n20013), .dout(n20016));
    jdff dff_B_ljbBY7Lj5_2(.din(n20016), .dout(n20019));
    jdff dff_B_vAfuBllz1_2(.din(n20019), .dout(n20022));
    jdff dff_B_9R6hN7230_2(.din(n20022), .dout(n20025));
    jdff dff_B_6eoxZfhQ4_2(.din(n20025), .dout(n20028));
    jdff dff_B_6LRWDamo4_2(.din(n20028), .dout(n20031));
    jdff dff_B_8fNPFrdf1_2(.din(n20031), .dout(n20034));
    jdff dff_B_aapST4Cv0_2(.din(n20034), .dout(n20037));
    jdff dff_B_UJh4Cvpm5_2(.din(n20037), .dout(n20040));
    jdff dff_B_3Rj94cVZ0_2(.din(n20040), .dout(n20043));
    jdff dff_B_xrHz6jpY7_2(.din(n20043), .dout(n20046));
    jdff dff_B_UUKJBab72_2(.din(n20046), .dout(n20049));
    jdff dff_B_bWkcc7Z69_2(.din(n20049), .dout(n20052));
    jdff dff_B_Jayjf1Sp4_2(.din(n20052), .dout(n20055));
    jdff dff_B_okZPYfUy4_1(.din(n5130), .dout(n20058));
    jdff dff_B_2FHgVOBY5_2(.din(n4827), .dout(n20061));
    jdff dff_B_AiUKz9DE9_2(.din(n20061), .dout(n20064));
    jdff dff_B_GxH1MmvG7_2(.din(n20064), .dout(n20067));
    jdff dff_B_m4tnjpuY3_2(.din(n20067), .dout(n20070));
    jdff dff_B_cfai8G0e3_2(.din(n20070), .dout(n20073));
    jdff dff_B_KKUPwmjX8_2(.din(n20073), .dout(n20076));
    jdff dff_B_aDOm0Xx91_2(.din(n20076), .dout(n20079));
    jdff dff_B_Rj9sCT1D3_2(.din(n20079), .dout(n20082));
    jdff dff_B_CPqFrG2y8_2(.din(n20082), .dout(n20085));
    jdff dff_B_3tQuH77c7_2(.din(n20085), .dout(n20088));
    jdff dff_B_0e7vG31u5_2(.din(n20088), .dout(n20091));
    jdff dff_B_TdBal9S57_2(.din(n20091), .dout(n20094));
    jdff dff_B_ft8Dn88k7_2(.din(n20094), .dout(n20097));
    jdff dff_B_e01OjxXX3_2(.din(n20097), .dout(n20100));
    jdff dff_B_AW0MOot52_2(.din(n20100), .dout(n20103));
    jdff dff_B_jl81WEhp0_2(.din(n20103), .dout(n20106));
    jdff dff_B_rBITXdHJ1_2(.din(n20106), .dout(n20109));
    jdff dff_B_RMp93ep76_2(.din(n20109), .dout(n20112));
    jdff dff_B_Pq315Gmc5_2(.din(n20112), .dout(n20115));
    jdff dff_B_GjW8idSO6_2(.din(n20115), .dout(n20118));
    jdff dff_B_PcNx6c0N0_2(.din(n20118), .dout(n20121));
    jdff dff_B_7AyP6H7O7_2(.din(n20121), .dout(n20124));
    jdff dff_B_rY2At0qi5_2(.din(n20124), .dout(n20127));
    jdff dff_B_uQXcYRnD8_2(.din(n20127), .dout(n20130));
    jdff dff_B_3HOUjZ767_2(.din(n20130), .dout(n20133));
    jdff dff_B_Q8KQnlZG4_2(.din(n20133), .dout(n20136));
    jdff dff_B_BfZmWP7T6_2(.din(n20136), .dout(n20139));
    jdff dff_B_TsQO7Wvf1_2(.din(n20139), .dout(n20142));
    jdff dff_B_zzPrbLCm3_2(.din(n20142), .dout(n20145));
    jdff dff_B_Te1i66hV5_2(.din(n20145), .dout(n20148));
    jdff dff_B_htUOUhmr2_2(.din(n20148), .dout(n20151));
    jdff dff_B_SvxBL2CX5_2(.din(n20151), .dout(n20154));
    jdff dff_B_XFH8kGgb9_2(.din(n20154), .dout(n20157));
    jdff dff_B_Eat20wwF4_2(.din(n20157), .dout(n20160));
    jdff dff_B_p53BAToJ1_2(.din(n20160), .dout(n20163));
    jdff dff_B_1If2QCPg3_2(.din(n20163), .dout(n20166));
    jdff dff_B_QzXJUNAG0_2(.din(n20166), .dout(n20169));
    jdff dff_B_Yt2BTntV6_2(.din(n20169), .dout(n20172));
    jdff dff_B_5Tscc3mU5_2(.din(n20172), .dout(n20175));
    jdff dff_B_46wlq6IK4_2(.din(n20175), .dout(n20178));
    jdff dff_B_GkOsAjCA5_1(.din(n4831), .dout(n20181));
    jdff dff_B_qCfy96cX7_2(.din(n4501), .dout(n20184));
    jdff dff_B_qWFkwedW8_2(.din(n20184), .dout(n20187));
    jdff dff_B_ETqTeCqg5_2(.din(n20187), .dout(n20190));
    jdff dff_B_mrs8oaK01_2(.din(n20190), .dout(n20193));
    jdff dff_B_Ym8bGeRl2_2(.din(n20193), .dout(n20196));
    jdff dff_B_DsylCa3W7_2(.din(n20196), .dout(n20199));
    jdff dff_B_ij8RsBNT2_2(.din(n20199), .dout(n20202));
    jdff dff_B_s822BQXD2_2(.din(n20202), .dout(n20205));
    jdff dff_B_4LJR26Zz4_2(.din(n20205), .dout(n20208));
    jdff dff_B_I8FsOP383_2(.din(n20208), .dout(n20211));
    jdff dff_B_4TyCm9ea4_2(.din(n20211), .dout(n20214));
    jdff dff_B_jNm1oBz20_2(.din(n20214), .dout(n20217));
    jdff dff_B_yDvWNEvw1_2(.din(n20217), .dout(n20220));
    jdff dff_B_jQSi0nhl7_2(.din(n20220), .dout(n20223));
    jdff dff_B_zYfO4QD10_2(.din(n20223), .dout(n20226));
    jdff dff_B_npo0KMU07_2(.din(n20226), .dout(n20229));
    jdff dff_B_zNGsRY8g2_2(.din(n20229), .dout(n20232));
    jdff dff_B_rm5N9AZt7_2(.din(n20232), .dout(n20235));
    jdff dff_B_wgWjRY6A8_2(.din(n20235), .dout(n20238));
    jdff dff_B_BOFFIOU05_2(.din(n20238), .dout(n20241));
    jdff dff_B_Gxmvnb5R5_2(.din(n20241), .dout(n20244));
    jdff dff_B_XvF3he9e9_2(.din(n20244), .dout(n20247));
    jdff dff_B_3LlcdKAo3_2(.din(n20247), .dout(n20250));
    jdff dff_B_a6VJsaRx5_2(.din(n20250), .dout(n20253));
    jdff dff_B_fj0iVqtX8_2(.din(n20253), .dout(n20256));
    jdff dff_B_fhlgibW17_2(.din(n20256), .dout(n20259));
    jdff dff_B_Cp7XneBh6_2(.din(n20259), .dout(n20262));
    jdff dff_B_5IhKFno72_2(.din(n20262), .dout(n20265));
    jdff dff_B_SDTPaPew4_2(.din(n20265), .dout(n20268));
    jdff dff_B_LosGJHyD2_2(.din(n20268), .dout(n20271));
    jdff dff_B_olGrOOJb1_2(.din(n20271), .dout(n20274));
    jdff dff_B_2MIsppXc9_2(.din(n20274), .dout(n20277));
    jdff dff_B_t4jWqFVG6_2(.din(n20277), .dout(n20280));
    jdff dff_B_OZ6qpPTy4_2(.din(n20280), .dout(n20283));
    jdff dff_B_wnkFhy2N6_2(.din(n20283), .dout(n20286));
    jdff dff_B_XlSilwFu7_2(.din(n20286), .dout(n20289));
    jdff dff_B_yriLKFxM6_2(.din(n20289), .dout(n20292));
    jdff dff_B_eWRukfmw4_1(.din(n4505), .dout(n20295));
    jdff dff_B_ydnRlVpB3_2(.din(n4151), .dout(n20298));
    jdff dff_B_w7fsqj4P0_2(.din(n20298), .dout(n20301));
    jdff dff_B_ObquUWuS3_2(.din(n20301), .dout(n20304));
    jdff dff_B_HB8JQfSM1_2(.din(n20304), .dout(n20307));
    jdff dff_B_F02MSOvL3_2(.din(n20307), .dout(n20310));
    jdff dff_B_FGbvqy2Q7_2(.din(n20310), .dout(n20313));
    jdff dff_B_QQupTRmD1_2(.din(n20313), .dout(n20316));
    jdff dff_B_71fpE7MR4_2(.din(n20316), .dout(n20319));
    jdff dff_B_NauiZ4Fy0_2(.din(n20319), .dout(n20322));
    jdff dff_B_RX9WqM9h0_2(.din(n20322), .dout(n20325));
    jdff dff_B_XI0Fftw28_2(.din(n20325), .dout(n20328));
    jdff dff_B_JPYRxwGb9_2(.din(n20328), .dout(n20331));
    jdff dff_B_5PY4syl25_2(.din(n20331), .dout(n20334));
    jdff dff_B_rM1B12IR7_2(.din(n20334), .dout(n20337));
    jdff dff_B_kzbweZEn4_2(.din(n20337), .dout(n20340));
    jdff dff_B_hPe3EIBr9_2(.din(n20340), .dout(n20343));
    jdff dff_B_jlKiSpEy3_2(.din(n20343), .dout(n20346));
    jdff dff_B_SvRxmqY43_2(.din(n20346), .dout(n20349));
    jdff dff_B_sVpnHyj48_2(.din(n20349), .dout(n20352));
    jdff dff_B_ZtETKS3z6_2(.din(n20352), .dout(n20355));
    jdff dff_B_moEckjPF2_2(.din(n20355), .dout(n20358));
    jdff dff_B_go3ZHA9c7_2(.din(n20358), .dout(n20361));
    jdff dff_B_nbiclrTt7_2(.din(n20361), .dout(n20364));
    jdff dff_B_ZGsriYPt7_2(.din(n20364), .dout(n20367));
    jdff dff_B_H2jBMIvq9_2(.din(n20367), .dout(n20370));
    jdff dff_B_RGsD2Ahi9_2(.din(n20370), .dout(n20373));
    jdff dff_B_3h3hCPL00_2(.din(n20373), .dout(n20376));
    jdff dff_B_MAN844QY8_2(.din(n20376), .dout(n20379));
    jdff dff_B_iHtcMqOh4_2(.din(n20379), .dout(n20382));
    jdff dff_B_KCXcFZxf4_2(.din(n20382), .dout(n20385));
    jdff dff_B_Ba1c2bqR6_2(.din(n20385), .dout(n20388));
    jdff dff_B_nAh4pjQW7_2(.din(n20388), .dout(n20391));
    jdff dff_B_L0ho2uIT0_2(.din(n20391), .dout(n20394));
    jdff dff_B_2vJ0ECc04_2(.din(n20394), .dout(n20397));
    jdff dff_B_FmIUrn9u6_1(.din(n4155), .dout(n20400));
    jdff dff_B_YhOheFMg0_2(.din(n3775), .dout(n20403));
    jdff dff_B_5cIrRVT33_2(.din(n20403), .dout(n20406));
    jdff dff_B_kOYBXiHE9_2(.din(n20406), .dout(n20409));
    jdff dff_B_M6Wwa9E80_2(.din(n20409), .dout(n20412));
    jdff dff_B_IbJm1Q2G1_2(.din(n20412), .dout(n20415));
    jdff dff_B_o65yV4W44_2(.din(n20415), .dout(n20418));
    jdff dff_B_oq3h95fv5_2(.din(n20418), .dout(n20421));
    jdff dff_B_YPRjFFTg2_2(.din(n20421), .dout(n20424));
    jdff dff_B_9jWxiIwf0_2(.din(n20424), .dout(n20427));
    jdff dff_B_9oihohtO2_2(.din(n20427), .dout(n20430));
    jdff dff_B_3L40jCqf7_2(.din(n20430), .dout(n20433));
    jdff dff_B_zL8YWxPk1_2(.din(n20433), .dout(n20436));
    jdff dff_B_5xWILhr79_2(.din(n20436), .dout(n20439));
    jdff dff_B_gRWqRPTD8_2(.din(n20439), .dout(n20442));
    jdff dff_B_Xvrm9jtV6_2(.din(n20442), .dout(n20445));
    jdff dff_B_M2GUvrHP8_2(.din(n20445), .dout(n20448));
    jdff dff_B_ezwzdqy06_2(.din(n20448), .dout(n20451));
    jdff dff_B_UTwgntyC9_2(.din(n20451), .dout(n20454));
    jdff dff_B_SyqnNlG53_2(.din(n20454), .dout(n20457));
    jdff dff_B_dXG8MYI47_2(.din(n20457), .dout(n20460));
    jdff dff_B_bivUJdQg9_2(.din(n20460), .dout(n20463));
    jdff dff_B_0hyWc2yJ5_2(.din(n20463), .dout(n20466));
    jdff dff_B_YkUMhdsQ6_2(.din(n20466), .dout(n20469));
    jdff dff_B_ALrXiQfO9_2(.din(n20469), .dout(n20472));
    jdff dff_B_3o62TwvU7_2(.din(n20472), .dout(n20475));
    jdff dff_B_hv9kSpGt7_2(.din(n20475), .dout(n20478));
    jdff dff_B_Cl89ITno8_2(.din(n20478), .dout(n20481));
    jdff dff_B_bvYFSfcm1_2(.din(n20481), .dout(n20484));
    jdff dff_B_4xLBcRnD9_2(.din(n20484), .dout(n20487));
    jdff dff_B_pMWVECVB6_2(.din(n20487), .dout(n20490));
    jdff dff_B_UImGPrEg1_2(.din(n20490), .dout(n20493));
    jdff dff_B_X9x5eONG1_1(.din(n3779), .dout(n20496));
    jdff dff_B_lfBrzUrz6_2(.din(n3395), .dout(n20499));
    jdff dff_B_I4gDPI392_2(.din(n20499), .dout(n20502));
    jdff dff_B_BYaGUQBu7_2(.din(n20502), .dout(n20505));
    jdff dff_B_4SEIkHOT4_2(.din(n20505), .dout(n20508));
    jdff dff_B_FoWaM2DB1_2(.din(n20508), .dout(n20511));
    jdff dff_B_vtqDLHrl3_2(.din(n20511), .dout(n20514));
    jdff dff_B_qlO9WPcz7_2(.din(n20514), .dout(n20517));
    jdff dff_B_Gv3WRA0O5_2(.din(n20517), .dout(n20520));
    jdff dff_B_Hym1lT2v2_2(.din(n20520), .dout(n20523));
    jdff dff_B_QnELvtVC3_2(.din(n20523), .dout(n20526));
    jdff dff_B_z5fmOBeh4_2(.din(n20526), .dout(n20529));
    jdff dff_B_xfTH8nsm5_2(.din(n20529), .dout(n20532));
    jdff dff_B_PwRJ4YaM8_2(.din(n20532), .dout(n20535));
    jdff dff_B_VIYUXkdD6_2(.din(n20535), .dout(n20538));
    jdff dff_B_c2ygEIGp6_2(.din(n20538), .dout(n20541));
    jdff dff_B_8K4SJKp38_2(.din(n20541), .dout(n20544));
    jdff dff_B_8WTgtnfC7_2(.din(n20544), .dout(n20547));
    jdff dff_B_URCHDs8v9_2(.din(n20547), .dout(n20550));
    jdff dff_B_y35Sv2AP7_2(.din(n20550), .dout(n20553));
    jdff dff_B_Oyr3oh2T5_2(.din(n20553), .dout(n20556));
    jdff dff_B_kj4TQQJI6_2(.din(n20556), .dout(n20559));
    jdff dff_B_U5nNO81N0_2(.din(n20559), .dout(n20562));
    jdff dff_B_W06xmaZP0_2(.din(n20562), .dout(n20565));
    jdff dff_B_gq6YKjlZ3_2(.din(n20565), .dout(n20568));
    jdff dff_B_bm1ZlNgl4_2(.din(n20568), .dout(n20571));
    jdff dff_B_HD6R4fCa1_2(.din(n20571), .dout(n20574));
    jdff dff_B_GZNE8dma7_2(.din(n20574), .dout(n20577));
    jdff dff_B_VDExURbU0_2(.din(n20577), .dout(n20580));
    jdff dff_B_70voapNf1_1(.din(n3399), .dout(n20583));
    jdff dff_B_TnajQOjF5_2(.din(n3004), .dout(n20586));
    jdff dff_B_nX7Vn4xJ0_2(.din(n20586), .dout(n20589));
    jdff dff_B_T0Uzh5Y36_2(.din(n20589), .dout(n20592));
    jdff dff_B_x0u8nhnw7_2(.din(n20592), .dout(n20595));
    jdff dff_B_jaIlhc4N4_2(.din(n20595), .dout(n20598));
    jdff dff_B_e4TP2vWq7_2(.din(n20598), .dout(n20601));
    jdff dff_B_nxV8kibe6_2(.din(n20601), .dout(n20604));
    jdff dff_B_c0u3t53e8_2(.din(n20604), .dout(n20607));
    jdff dff_B_PIbZcqUT2_2(.din(n20607), .dout(n20610));
    jdff dff_B_91UUNVtU3_2(.din(n20610), .dout(n20613));
    jdff dff_B_wFMIMidM1_2(.din(n20613), .dout(n20616));
    jdff dff_B_8t7O4wBV8_2(.din(n20616), .dout(n20619));
    jdff dff_B_tRlUm20j6_2(.din(n20619), .dout(n20622));
    jdff dff_B_QyVkVUSp4_2(.din(n20622), .dout(n20625));
    jdff dff_B_YymKICMc9_2(.din(n20625), .dout(n20628));
    jdff dff_B_aCMHH9qC4_2(.din(n20628), .dout(n20631));
    jdff dff_B_hwY2v7cA7_2(.din(n20631), .dout(n20634));
    jdff dff_B_vVhDKRVx4_2(.din(n20634), .dout(n20637));
    jdff dff_B_6WwIKGxL4_2(.din(n20637), .dout(n20640));
    jdff dff_B_TRxvA4oM1_2(.din(n20640), .dout(n20643));
    jdff dff_B_QFo2R29W7_2(.din(n20643), .dout(n20646));
    jdff dff_B_lWDsRKFF7_2(.din(n20646), .dout(n20649));
    jdff dff_B_Wa67a40Z2_2(.din(n20649), .dout(n20652));
    jdff dff_B_2mA5JmjA2_2(.din(n20652), .dout(n20655));
    jdff dff_B_5ffPzOR82_2(.din(n20655), .dout(n20658));
    jdff dff_B_AojH413d8_1(.din(n3008), .dout(n20661));
    jdff dff_B_bojL8AXu1_2(.din(n2629), .dout(n20664));
    jdff dff_B_SFc7Rnd68_2(.din(n20664), .dout(n20667));
    jdff dff_B_UEQUFxnz8_2(.din(n20667), .dout(n20670));
    jdff dff_B_5pgdEYHc1_2(.din(n20670), .dout(n20673));
    jdff dff_B_Ek4SrkcL4_2(.din(n20673), .dout(n20676));
    jdff dff_B_Ykuj1MrY5_2(.din(n20676), .dout(n20679));
    jdff dff_B_Z8op9tpd0_2(.din(n20679), .dout(n20682));
    jdff dff_B_5E3MbnFt2_2(.din(n20682), .dout(n20685));
    jdff dff_B_WVyxDF8I4_2(.din(n20685), .dout(n20688));
    jdff dff_B_b1NwTAOJ4_2(.din(n20688), .dout(n20691));
    jdff dff_B_lNHeQRKb6_2(.din(n20691), .dout(n20694));
    jdff dff_B_VAyTxHL41_2(.din(n20694), .dout(n20697));
    jdff dff_B_fTBCHUgh1_2(.din(n20697), .dout(n20700));
    jdff dff_B_DQMvKJ7t2_2(.din(n20700), .dout(n20703));
    jdff dff_B_g8yulbvU8_2(.din(n20703), .dout(n20706));
    jdff dff_B_H6I1go5J2_2(.din(n20706), .dout(n20709));
    jdff dff_B_DWQ0Z7NF1_2(.din(n20709), .dout(n20712));
    jdff dff_B_3naLMSS43_2(.din(n20712), .dout(n20715));
    jdff dff_B_LKYOLMbw2_2(.din(n20715), .dout(n20718));
    jdff dff_B_Xe8hfpQ35_2(.din(n20718), .dout(n20721));
    jdff dff_B_djo0VUY31_2(.din(n20721), .dout(n20724));
    jdff dff_B_IUpPIGVx7_2(.din(n20724), .dout(n20727));
    jdff dff_B_fmHAL9ae8_1(.din(n2633), .dout(n20730));
    jdff dff_B_p0tE444d6_2(.din(n2278), .dout(n20733));
    jdff dff_B_K7UTe42L6_2(.din(n20733), .dout(n20736));
    jdff dff_B_usZ9fHwx7_2(.din(n20736), .dout(n20739));
    jdff dff_B_CbklaxfM4_2(.din(n20739), .dout(n20742));
    jdff dff_B_nYoSMv0S4_2(.din(n20742), .dout(n20745));
    jdff dff_B_Y01bI1t40_2(.din(n20745), .dout(n20748));
    jdff dff_B_lyYWGvSQ6_2(.din(n20748), .dout(n20751));
    jdff dff_B_SpMFarON3_2(.din(n20751), .dout(n20754));
    jdff dff_B_wHlfpW2R6_2(.din(n20754), .dout(n20757));
    jdff dff_B_2SCrIjwV1_2(.din(n20757), .dout(n20760));
    jdff dff_B_DAxOj5kw2_2(.din(n20760), .dout(n20763));
    jdff dff_B_F5LGktB03_2(.din(n20763), .dout(n20766));
    jdff dff_B_dL8pwDjZ5_2(.din(n20766), .dout(n20769));
    jdff dff_B_4125E9pF6_2(.din(n20769), .dout(n20772));
    jdff dff_B_ouX0EVPl2_2(.din(n20772), .dout(n20775));
    jdff dff_B_cMnm8UwX8_2(.din(n20775), .dout(n20778));
    jdff dff_B_YZicZTeH6_2(.din(n20778), .dout(n20781));
    jdff dff_B_JOVUyAjR9_2(.din(n20781), .dout(n20784));
    jdff dff_B_XIqTUG0R2_2(.din(n20784), .dout(n20787));
    jdff dff_B_C3gKgd3D9_1(.din(n2282), .dout(n20790));
    jdff dff_B_UIQ4Tq8K0_2(.din(n1954), .dout(n20793));
    jdff dff_B_xZKQC6Z66_2(.din(n20793), .dout(n20796));
    jdff dff_B_lNb5zbNw0_2(.din(n20796), .dout(n20799));
    jdff dff_B_ga64F56D5_2(.din(n20799), .dout(n20802));
    jdff dff_B_d7xdTB787_2(.din(n20802), .dout(n20805));
    jdff dff_B_2feWtac50_2(.din(n20805), .dout(n20808));
    jdff dff_B_WQK4Y9oX0_2(.din(n20808), .dout(n20811));
    jdff dff_B_Yk8M5kI21_2(.din(n20811), .dout(n20814));
    jdff dff_B_f4xQt3x57_2(.din(n20814), .dout(n20817));
    jdff dff_B_eYPa24kv9_2(.din(n20817), .dout(n20820));
    jdff dff_B_5xrQ4LJY0_2(.din(n20820), .dout(n20823));
    jdff dff_B_fErRU8Wa4_2(.din(n20823), .dout(n20826));
    jdff dff_B_Bd6Lq7wK7_2(.din(n20826), .dout(n20829));
    jdff dff_B_x36fGRs87_2(.din(n20829), .dout(n20832));
    jdff dff_B_D8eIa9Ef0_2(.din(n20832), .dout(n20835));
    jdff dff_B_uF078E1D9_2(.din(n20835), .dout(n20838));
    jdff dff_B_sw5cd2Qe4_1(.din(n1958), .dout(n20841));
    jdff dff_B_FGIlsyaX8_2(.din(n1657), .dout(n20844));
    jdff dff_B_n0mfdLxC7_2(.din(n20844), .dout(n20847));
    jdff dff_B_62jIwzj55_2(.din(n20847), .dout(n20850));
    jdff dff_B_XhVzmfEv7_2(.din(n20850), .dout(n20853));
    jdff dff_B_5eJCXF1s5_2(.din(n20853), .dout(n20856));
    jdff dff_B_NOQRRBaB4_2(.din(n20856), .dout(n20859));
    jdff dff_B_kHeG3J936_2(.din(n20859), .dout(n20862));
    jdff dff_B_YZ9xqlzj5_2(.din(n20862), .dout(n20865));
    jdff dff_B_iHiiKhso8_2(.din(n20865), .dout(n20868));
    jdff dff_B_1lthIbJN1_2(.din(n20868), .dout(n20871));
    jdff dff_B_ZEY1crJr7_2(.din(n20871), .dout(n20874));
    jdff dff_B_54IVPH8S9_2(.din(n20874), .dout(n20877));
    jdff dff_B_jEXVVydu5_2(.din(n20877), .dout(n20880));
    jdff dff_B_w72PYw6U1_1(.din(n1661), .dout(n20883));
    jdff dff_B_GVirOKkz8_2(.din(n1387), .dout(n20886));
    jdff dff_B_8VwgNTfV6_2(.din(n20886), .dout(n20889));
    jdff dff_B_LGWtgeBN4_2(.din(n20889), .dout(n20892));
    jdff dff_B_p1Qsan2p5_2(.din(n20892), .dout(n20895));
    jdff dff_B_KAxhzIm75_2(.din(n20895), .dout(n20898));
    jdff dff_B_FNNwejJq3_2(.din(n20898), .dout(n20901));
    jdff dff_B_BMlDPU3H2_2(.din(n20901), .dout(n20904));
    jdff dff_B_j38HnXvi8_2(.din(n20904), .dout(n20907));
    jdff dff_B_LmNVtie13_2(.din(n20907), .dout(n20910));
    jdff dff_B_LCG7Dk6n8_2(.din(n20910), .dout(n20913));
    jdff dff_B_JyHIx9uu1_2(.din(n1399), .dout(n20916));
    jdff dff_B_thuy0MMT4_1(.din(n1391), .dout(n20919));
    jdff dff_B_ljJHdLN36_2(.din(n1147), .dout(n20922));
    jdff dff_B_h6o6Ds5F7_2(.din(n20922), .dout(n20925));
    jdff dff_B_YtVsayaB5_2(.din(n20925), .dout(n20928));
    jdff dff_B_cjpEUtrF4_2(.din(n20928), .dout(n20931));
    jdff dff_B_5WzQe57n6_2(.din(n20931), .dout(n20934));
    jdff dff_B_sUOIGnBS8_2(.din(n20934), .dout(n20937));
    jdff dff_B_6texNomC5_2(.din(n1200), .dout(n20940));
    jdff dff_B_q5ZAGjY43_2(.din(n937), .dout(n20943));
    jdff dff_B_ZYfDr3Pu6_2(.din(n20943), .dout(n20946));
    jdff dff_B_rXwee7iy7_2(.din(n20946), .dout(n20949));
    jdff dff_B_z4cPPlU19_0(.din(n956), .dout(n20952));
    jdff dff_A_UHb6hdmf2_0(.din(n20957), .dout(n20954));
    jdff dff_A_OoN2Prmy8_0(.din(n740), .dout(n20957));
    jdff dff_A_xqfz72US4_1(.din(n20963), .dout(n20960));
    jdff dff_A_U7KNUsVf3_1(.din(n740), .dout(n20963));
    jdff dff_B_QvWK9LdJ4_1(.din(n5669), .dout(n20967));
    jdff dff_B_ppWMHWH82_2(.din(n5417), .dout(n20970));
    jdff dff_B_Du9yRvuv4_2(.din(n20970), .dout(n20973));
    jdff dff_B_rfOzPZWh0_2(.din(n20973), .dout(n20976));
    jdff dff_B_YRD4GLRA9_2(.din(n20976), .dout(n20979));
    jdff dff_B_qtVBLd7Y9_2(.din(n20979), .dout(n20982));
    jdff dff_B_xXxxeo2k8_2(.din(n20982), .dout(n20985));
    jdff dff_B_d8ZyoDXL4_2(.din(n20985), .dout(n20988));
    jdff dff_B_ZSyl96Lv8_2(.din(n20988), .dout(n20991));
    jdff dff_B_ty4Ue4Zf2_2(.din(n20991), .dout(n20994));
    jdff dff_B_QUKVixNC3_2(.din(n20994), .dout(n20997));
    jdff dff_B_EAF4somy5_2(.din(n20997), .dout(n21000));
    jdff dff_B_C9a3ZSxp0_2(.din(n21000), .dout(n21003));
    jdff dff_B_tNmU4ROw3_2(.din(n21003), .dout(n21006));
    jdff dff_B_8gGogAKO4_2(.din(n21006), .dout(n21009));
    jdff dff_B_iHw0yWVS2_2(.din(n21009), .dout(n21012));
    jdff dff_B_BfLDeT4F0_2(.din(n21012), .dout(n21015));
    jdff dff_B_HHnTZyAA9_2(.din(n21015), .dout(n21018));
    jdff dff_B_6myBpVsI6_2(.din(n21018), .dout(n21021));
    jdff dff_B_RKm6MBC72_2(.din(n21021), .dout(n21024));
    jdff dff_B_CYVv1W5i4_2(.din(n21024), .dout(n21027));
    jdff dff_B_l3al1kNK2_2(.din(n21027), .dout(n21030));
    jdff dff_B_6DiyvSLa4_2(.din(n21030), .dout(n21033));
    jdff dff_B_coAxeVZi2_2(.din(n21033), .dout(n21036));
    jdff dff_B_Bm9ZbwX94_2(.din(n21036), .dout(n21039));
    jdff dff_B_DSTJ5NN37_2(.din(n21039), .dout(n21042));
    jdff dff_B_bvZFtliG9_2(.din(n21042), .dout(n21045));
    jdff dff_B_U2I4LaUO3_2(.din(n21045), .dout(n21048));
    jdff dff_B_3EmoHhCN9_2(.din(n21048), .dout(n21051));
    jdff dff_B_vpWzQMEl9_2(.din(n21051), .dout(n21054));
    jdff dff_B_RaFgWQMW8_2(.din(n21054), .dout(n21057));
    jdff dff_B_85e4b9YS0_2(.din(n21057), .dout(n21060));
    jdff dff_B_TwqKLTjI6_2(.din(n21060), .dout(n21063));
    jdff dff_B_IJpz2FlE4_2(.din(n21063), .dout(n21066));
    jdff dff_B_RXGS2Cq57_2(.din(n21066), .dout(n21069));
    jdff dff_B_NqeVhiCF4_2(.din(n21069), .dout(n21072));
    jdff dff_B_KE23DJSF1_2(.din(n21072), .dout(n21075));
    jdff dff_B_27oEDSQy4_2(.din(n21075), .dout(n21078));
    jdff dff_B_WcwpsT4j7_2(.din(n21078), .dout(n21081));
    jdff dff_B_OhiqQqoW1_2(.din(n21081), .dout(n21084));
    jdff dff_B_e4TzaCi25_2(.din(n21084), .dout(n21087));
    jdff dff_B_zgaLzjm17_2(.din(n21087), .dout(n21090));
    jdff dff_B_ufmkUT7W0_2(.din(n21090), .dout(n21093));
    jdff dff_B_OfDykzgp6_2(.din(n21093), .dout(n21096));
    jdff dff_B_769FflUu8_2(.din(n21096), .dout(n21099));
    jdff dff_B_cWIKRbme5_2(.din(n21099), .dout(n21102));
    jdff dff_B_bG14cOkU1_2(.din(n21102), .dout(n21105));
    jdff dff_B_xTRmInr30_0(.din(n5665), .dout(n21108));
    jdff dff_A_Z1NK3AwW0_1(.din(n5622), .dout(n21110));
    jdff dff_B_JumOCHSu3_1(.din(n5421), .dout(n21114));
    jdff dff_B_djXDBNZ67_2(.din(n5145), .dout(n21117));
    jdff dff_B_rgShl3M96_2(.din(n21117), .dout(n21120));
    jdff dff_B_MbQSwguy8_2(.din(n21120), .dout(n21123));
    jdff dff_B_rTXAzY9u6_2(.din(n21123), .dout(n21126));
    jdff dff_B_TAxIsREk8_2(.din(n21126), .dout(n21129));
    jdff dff_B_SWI5FPZO2_2(.din(n21129), .dout(n21132));
    jdff dff_B_nES1lzeJ1_2(.din(n21132), .dout(n21135));
    jdff dff_B_6yVykT7u9_2(.din(n21135), .dout(n21138));
    jdff dff_B_X9DvH45u2_2(.din(n21138), .dout(n21141));
    jdff dff_B_TOFT54Yp0_2(.din(n21141), .dout(n21144));
    jdff dff_B_OdCsBtY38_2(.din(n21144), .dout(n21147));
    jdff dff_B_g10y2h3c7_2(.din(n21147), .dout(n21150));
    jdff dff_B_f3DeNnlr7_2(.din(n21150), .dout(n21153));
    jdff dff_B_SxCiQWFo4_2(.din(n21153), .dout(n21156));
    jdff dff_B_v9SIsnLb9_2(.din(n21156), .dout(n21159));
    jdff dff_B_ZNzTCBjo3_2(.din(n21159), .dout(n21162));
    jdff dff_B_egjYoBMq4_2(.din(n21162), .dout(n21165));
    jdff dff_B_k4CU2HWw1_2(.din(n21165), .dout(n21168));
    jdff dff_B_faOXZq9f7_2(.din(n21168), .dout(n21171));
    jdff dff_B_Ztrfcz5F5_2(.din(n21171), .dout(n21174));
    jdff dff_B_an9KytBv9_2(.din(n21174), .dout(n21177));
    jdff dff_B_LTd2AH0n9_2(.din(n21177), .dout(n21180));
    jdff dff_B_vd0NwYDS0_2(.din(n21180), .dout(n21183));
    jdff dff_B_jpAy5BiJ6_2(.din(n21183), .dout(n21186));
    jdff dff_B_Jx3w7Wv96_2(.din(n21186), .dout(n21189));
    jdff dff_B_mx0KoNRe1_2(.din(n21189), .dout(n21192));
    jdff dff_B_Lrim48jw3_2(.din(n21192), .dout(n21195));
    jdff dff_B_Gywrwyt91_2(.din(n21195), .dout(n21198));
    jdff dff_B_4stycAfw9_2(.din(n21198), .dout(n21201));
    jdff dff_B_5v1tJlmS4_2(.din(n21201), .dout(n21204));
    jdff dff_B_o9DQ50o20_2(.din(n21204), .dout(n21207));
    jdff dff_B_EMoVDda25_2(.din(n21207), .dout(n21210));
    jdff dff_B_480Yo4J14_2(.din(n21210), .dout(n21213));
    jdff dff_B_KftfVnJe9_2(.din(n21213), .dout(n21216));
    jdff dff_B_6Q6U5BxS6_2(.din(n21216), .dout(n21219));
    jdff dff_B_lgHEpE4d0_2(.din(n21219), .dout(n21222));
    jdff dff_B_KgXNBHXA8_2(.din(n21222), .dout(n21225));
    jdff dff_B_0qqmCVOu2_2(.din(n21225), .dout(n21228));
    jdff dff_B_cyDokG0S9_2(.din(n21228), .dout(n21231));
    jdff dff_B_GRujP2cX2_2(.din(n21231), .dout(n21234));
    jdff dff_B_sDfgSwXx5_2(.din(n21234), .dout(n21237));
    jdff dff_B_OeZSAjlN6_2(.din(n5350), .dout(n21240));
    jdff dff_B_48fLUiLC1_1(.din(n5149), .dout(n21243));
    jdff dff_B_Ze3kLx3K1_2(.din(n4846), .dout(n21246));
    jdff dff_B_D0RzeeaR9_2(.din(n21246), .dout(n21249));
    jdff dff_B_uvEPI7238_2(.din(n21249), .dout(n21252));
    jdff dff_B_1GtuQFdD7_2(.din(n21252), .dout(n21255));
    jdff dff_B_6I9bN3aj2_2(.din(n21255), .dout(n21258));
    jdff dff_B_pDkBuq3W4_2(.din(n21258), .dout(n21261));
    jdff dff_B_l6egQqTq1_2(.din(n21261), .dout(n21264));
    jdff dff_B_EeIx6lWu5_2(.din(n21264), .dout(n21267));
    jdff dff_B_ZKzze1G45_2(.din(n21267), .dout(n21270));
    jdff dff_B_5EIQBByw2_2(.din(n21270), .dout(n21273));
    jdff dff_B_WnUd9fAB9_2(.din(n21273), .dout(n21276));
    jdff dff_B_XJ7ye8VP4_2(.din(n21276), .dout(n21279));
    jdff dff_B_iATijlvg3_2(.din(n21279), .dout(n21282));
    jdff dff_B_WJsVMLVr2_2(.din(n21282), .dout(n21285));
    jdff dff_B_SoQN8u6O6_2(.din(n21285), .dout(n21288));
    jdff dff_B_WMpKEzfw9_2(.din(n21288), .dout(n21291));
    jdff dff_B_VyaUp4V64_2(.din(n21291), .dout(n21294));
    jdff dff_B_eOWDQZM86_2(.din(n21294), .dout(n21297));
    jdff dff_B_9fiXV1DK3_2(.din(n21297), .dout(n21300));
    jdff dff_B_cVKcOvl73_2(.din(n21300), .dout(n21303));
    jdff dff_B_2cCtsE6g0_2(.din(n21303), .dout(n21306));
    jdff dff_B_QFeoGzuf5_2(.din(n21306), .dout(n21309));
    jdff dff_B_MpVpW8QW2_2(.din(n21309), .dout(n21312));
    jdff dff_B_9I3MpTzM1_2(.din(n21312), .dout(n21315));
    jdff dff_B_FsC1pxoD0_2(.din(n21315), .dout(n21318));
    jdff dff_B_npHzAUx52_2(.din(n21318), .dout(n21321));
    jdff dff_B_lmkokJKy3_2(.din(n21321), .dout(n21324));
    jdff dff_B_Nla71nIv1_2(.din(n21324), .dout(n21327));
    jdff dff_B_rBTTfBLi3_2(.din(n21327), .dout(n21330));
    jdff dff_B_OsS6zM8y5_2(.din(n21330), .dout(n21333));
    jdff dff_B_j7TGoQOg7_2(.din(n21333), .dout(n21336));
    jdff dff_B_1xncBhks8_2(.din(n21336), .dout(n21339));
    jdff dff_B_aauT4CO23_2(.din(n21339), .dout(n21342));
    jdff dff_B_hK8ZzDrd1_2(.din(n21342), .dout(n21345));
    jdff dff_B_OzuIHOuw2_2(.din(n21345), .dout(n21348));
    jdff dff_B_SyOUUt9X8_2(.din(n21348), .dout(n21351));
    jdff dff_B_yX9rmHxl6_2(.din(n21351), .dout(n21354));
    jdff dff_B_tUH2K1Kj7_2(.din(n21354), .dout(n21357));
    jdff dff_B_lcTOel7j3_2(.din(n5051), .dout(n21360));
    jdff dff_B_uDtCWuTI2_1(.din(n4850), .dout(n21363));
    jdff dff_B_6Yaw6uqx5_2(.din(n4520), .dout(n21366));
    jdff dff_B_LKpBOd4S8_2(.din(n21366), .dout(n21369));
    jdff dff_B_yJLB6yw02_2(.din(n21369), .dout(n21372));
    jdff dff_B_GsbWfNwj8_2(.din(n21372), .dout(n21375));
    jdff dff_B_z9ITqEVW7_2(.din(n21375), .dout(n21378));
    jdff dff_B_p9IB5jVJ4_2(.din(n21378), .dout(n21381));
    jdff dff_B_EDkMg6i13_2(.din(n21381), .dout(n21384));
    jdff dff_B_lP6sjAII6_2(.din(n21384), .dout(n21387));
    jdff dff_B_8h7NaPld4_2(.din(n21387), .dout(n21390));
    jdff dff_B_J6f9wVXD2_2(.din(n21390), .dout(n21393));
    jdff dff_B_KD3qxIVs4_2(.din(n21393), .dout(n21396));
    jdff dff_B_txNDtw8o4_2(.din(n21396), .dout(n21399));
    jdff dff_B_GpM0pypo0_2(.din(n21399), .dout(n21402));
    jdff dff_B_iCeFsNNo9_2(.din(n21402), .dout(n21405));
    jdff dff_B_CUFHkhrZ5_2(.din(n21405), .dout(n21408));
    jdff dff_B_GIlZr1Dv9_2(.din(n21408), .dout(n21411));
    jdff dff_B_DEd7KeBy8_2(.din(n21411), .dout(n21414));
    jdff dff_B_NrOlrH518_2(.din(n21414), .dout(n21417));
    jdff dff_B_Lth8MXWF7_2(.din(n21417), .dout(n21420));
    jdff dff_B_GH5mXvln3_2(.din(n21420), .dout(n21423));
    jdff dff_B_nWFoS2jl6_2(.din(n21423), .dout(n21426));
    jdff dff_B_xiXCikwH9_2(.din(n21426), .dout(n21429));
    jdff dff_B_jQFxVyoR7_2(.din(n21429), .dout(n21432));
    jdff dff_B_i0DgvZ6z9_2(.din(n21432), .dout(n21435));
    jdff dff_B_psaKYNCg1_2(.din(n21435), .dout(n21438));
    jdff dff_B_zO67d4XR7_2(.din(n21438), .dout(n21441));
    jdff dff_B_PchzTo831_2(.din(n21441), .dout(n21444));
    jdff dff_B_FhYYglJE0_2(.din(n21444), .dout(n21447));
    jdff dff_B_0Z8dxuCq2_2(.din(n21447), .dout(n21450));
    jdff dff_B_raInsWt43_2(.din(n21450), .dout(n21453));
    jdff dff_B_xjhE7TFx1_2(.din(n21453), .dout(n21456));
    jdff dff_B_wtkhyI6N7_2(.din(n21456), .dout(n21459));
    jdff dff_B_MB2L94Ng8_2(.din(n21459), .dout(n21462));
    jdff dff_B_Jhi8veVz7_2(.din(n21462), .dout(n21465));
    jdff dff_B_1dOlMKis6_2(.din(n21465), .dout(n21468));
    jdff dff_B_Jne99qpP9_2(.din(n4725), .dout(n21471));
    jdff dff_B_wqdKiwbS9_1(.din(n4524), .dout(n21474));
    jdff dff_B_CHpjLhuk3_2(.din(n4170), .dout(n21477));
    jdff dff_B_LpyoHiG38_2(.din(n21477), .dout(n21480));
    jdff dff_B_oT9evhYB1_2(.din(n21480), .dout(n21483));
    jdff dff_B_YfPu9CoH1_2(.din(n21483), .dout(n21486));
    jdff dff_B_58QxJlSM5_2(.din(n21486), .dout(n21489));
    jdff dff_B_zteXz2tj4_2(.din(n21489), .dout(n21492));
    jdff dff_B_tzSbd6xs9_2(.din(n21492), .dout(n21495));
    jdff dff_B_QoKpxNwm7_2(.din(n21495), .dout(n21498));
    jdff dff_B_1HGe7cXS1_2(.din(n21498), .dout(n21501));
    jdff dff_B_btzooBeW8_2(.din(n21501), .dout(n21504));
    jdff dff_B_pWBrxOSL1_2(.din(n21504), .dout(n21507));
    jdff dff_B_DPu6pGJB2_2(.din(n21507), .dout(n21510));
    jdff dff_B_AzLLaukc4_2(.din(n21510), .dout(n21513));
    jdff dff_B_9VsHYNVU5_2(.din(n21513), .dout(n21516));
    jdff dff_B_R2wqIfy29_2(.din(n21516), .dout(n21519));
    jdff dff_B_61Mi9vDS6_2(.din(n21519), .dout(n21522));
    jdff dff_B_m9xDWTid6_2(.din(n21522), .dout(n21525));
    jdff dff_B_CcgNIaTM2_2(.din(n21525), .dout(n21528));
    jdff dff_B_h5OAkxsp3_2(.din(n21528), .dout(n21531));
    jdff dff_B_HEGYzhwY5_2(.din(n21531), .dout(n21534));
    jdff dff_B_kfbk9PY04_2(.din(n21534), .dout(n21537));
    jdff dff_B_jmaO7NWx0_2(.din(n21537), .dout(n21540));
    jdff dff_B_TShXzsna3_2(.din(n21540), .dout(n21543));
    jdff dff_B_pNS8rVN69_2(.din(n21543), .dout(n21546));
    jdff dff_B_hFPCJFyh2_2(.din(n21546), .dout(n21549));
    jdff dff_B_A0tafV0w9_2(.din(n21549), .dout(n21552));
    jdff dff_B_AEbfou5c6_2(.din(n21552), .dout(n21555));
    jdff dff_B_K75tx89b6_2(.din(n21555), .dout(n21558));
    jdff dff_B_wzPUwsfF3_2(.din(n21558), .dout(n21561));
    jdff dff_B_ZZcJZLBn4_2(.din(n21561), .dout(n21564));
    jdff dff_B_4VF6pijT7_2(.din(n21564), .dout(n21567));
    jdff dff_B_4HCmCGDr6_2(.din(n21567), .dout(n21570));
    jdff dff_B_xjUxkvVQ5_2(.din(n4375), .dout(n21573));
    jdff dff_B_Ks3Cgzof9_1(.din(n4174), .dout(n21576));
    jdff dff_B_LotTPgHT2_2(.din(n3794), .dout(n21579));
    jdff dff_B_eiVwXRlF0_2(.din(n21579), .dout(n21582));
    jdff dff_B_GApNkSkT3_2(.din(n21582), .dout(n21585));
    jdff dff_B_0UPiT9ic9_2(.din(n21585), .dout(n21588));
    jdff dff_B_Il2GKSpk7_2(.din(n21588), .dout(n21591));
    jdff dff_B_lUTGmdDb2_2(.din(n21591), .dout(n21594));
    jdff dff_B_xuW5NKz55_2(.din(n21594), .dout(n21597));
    jdff dff_B_w1R3Xp8i3_2(.din(n21597), .dout(n21600));
    jdff dff_B_DQw6JW6I5_2(.din(n21600), .dout(n21603));
    jdff dff_B_ThdgcyjF7_2(.din(n21603), .dout(n21606));
    jdff dff_B_Fm0jZ2AS0_2(.din(n21606), .dout(n21609));
    jdff dff_B_9hfurshI2_2(.din(n21609), .dout(n21612));
    jdff dff_B_fFRCeOFU6_2(.din(n21612), .dout(n21615));
    jdff dff_B_sL9yCUtx2_2(.din(n21615), .dout(n21618));
    jdff dff_B_zBNIm5ku7_2(.din(n21618), .dout(n21621));
    jdff dff_B_35zlfNO25_2(.din(n21621), .dout(n21624));
    jdff dff_B_ozIz7hsk9_2(.din(n21624), .dout(n21627));
    jdff dff_B_iBDx4kTa8_2(.din(n21627), .dout(n21630));
    jdff dff_B_FRqwOUtL0_2(.din(n21630), .dout(n21633));
    jdff dff_B_5SioB8bi0_2(.din(n21633), .dout(n21636));
    jdff dff_B_dRfhkIXO6_2(.din(n21636), .dout(n21639));
    jdff dff_B_meGfJ4Ml7_2(.din(n21639), .dout(n21642));
    jdff dff_B_THRXSfUE3_2(.din(n21642), .dout(n21645));
    jdff dff_B_djv53PIm9_2(.din(n21645), .dout(n21648));
    jdff dff_B_EQBEhJzu3_2(.din(n21648), .dout(n21651));
    jdff dff_B_SbD6dXDL5_2(.din(n21651), .dout(n21654));
    jdff dff_B_PZcz0VKj4_2(.din(n21654), .dout(n21657));
    jdff dff_B_Vv5vw15y6_2(.din(n21657), .dout(n21660));
    jdff dff_B_wqQfrI6j6_2(.din(n21660), .dout(n21663));
    jdff dff_B_xho3upNn0_2(.din(n3995), .dout(n21666));
    jdff dff_B_fiFeTNe63_1(.din(n3798), .dout(n21669));
    jdff dff_B_9HwILk8E8_2(.din(n3414), .dout(n21672));
    jdff dff_B_BmLP96EL6_2(.din(n21672), .dout(n21675));
    jdff dff_B_95OsEaqm3_2(.din(n21675), .dout(n21678));
    jdff dff_B_u1vD9SdR2_2(.din(n21678), .dout(n21681));
    jdff dff_B_iyhTj8nm2_2(.din(n21681), .dout(n21684));
    jdff dff_B_M4IeJZNd0_2(.din(n21684), .dout(n21687));
    jdff dff_B_ZEyAsnHN7_2(.din(n21687), .dout(n21690));
    jdff dff_B_4WlfT4Mr9_2(.din(n21690), .dout(n21693));
    jdff dff_B_tbs6DpMD0_2(.din(n21693), .dout(n21696));
    jdff dff_B_L8MrorfR3_2(.din(n21696), .dout(n21699));
    jdff dff_B_u8g5p00Q1_2(.din(n21699), .dout(n21702));
    jdff dff_B_5dMGJnKw8_2(.din(n21702), .dout(n21705));
    jdff dff_B_auTy16xV2_2(.din(n21705), .dout(n21708));
    jdff dff_B_jzl2WbeF3_2(.din(n21708), .dout(n21711));
    jdff dff_B_VAok8B1c7_2(.din(n21711), .dout(n21714));
    jdff dff_B_UYzEA5X27_2(.din(n21714), .dout(n21717));
    jdff dff_B_d2Gkv2e39_2(.din(n21717), .dout(n21720));
    jdff dff_B_0eXg0p0U9_2(.din(n21720), .dout(n21723));
    jdff dff_B_xiRj92M16_2(.din(n21723), .dout(n21726));
    jdff dff_B_u6oZYj6j5_2(.din(n21726), .dout(n21729));
    jdff dff_B_TnozkIyp2_2(.din(n21729), .dout(n21732));
    jdff dff_B_qnhEsylH2_2(.din(n21732), .dout(n21735));
    jdff dff_B_qkhO7al72_2(.din(n21735), .dout(n21738));
    jdff dff_B_y6kwC2sf6_2(.din(n21738), .dout(n21741));
    jdff dff_B_vV0bDt1L1_2(.din(n21741), .dout(n21744));
    jdff dff_B_lZ5Qjorr3_2(.din(n21744), .dout(n21747));
    jdff dff_B_bcP0E7Hi5_2(.din(n3612), .dout(n21750));
    jdff dff_B_PDENw4BN8_1(.din(n3418), .dout(n21753));
    jdff dff_B_hNgHePwe0_2(.din(n3023), .dout(n21756));
    jdff dff_B_LygJ5N0O7_2(.din(n21756), .dout(n21759));
    jdff dff_B_vLA6d5pQ6_2(.din(n21759), .dout(n21762));
    jdff dff_B_Cgfh33L38_2(.din(n21762), .dout(n21765));
    jdff dff_B_SlTnutle6_2(.din(n21765), .dout(n21768));
    jdff dff_B_piViiJcf3_2(.din(n21768), .dout(n21771));
    jdff dff_B_o90DMMD02_2(.din(n21771), .dout(n21774));
    jdff dff_B_4XRK2MfO1_2(.din(n21774), .dout(n21777));
    jdff dff_B_Umx2e0Ti1_2(.din(n21777), .dout(n21780));
    jdff dff_B_V9ZXbxxY2_2(.din(n21780), .dout(n21783));
    jdff dff_B_ptmoT6kf6_2(.din(n21783), .dout(n21786));
    jdff dff_B_uyGMp8xf6_2(.din(n21786), .dout(n21789));
    jdff dff_B_0aqzSceQ4_2(.din(n21789), .dout(n21792));
    jdff dff_B_WfaHkpyi8_2(.din(n21792), .dout(n21795));
    jdff dff_B_FQgo4IeQ5_2(.din(n21795), .dout(n21798));
    jdff dff_B_aHhwdnR76_2(.din(n21798), .dout(n21801));
    jdff dff_B_EZTUX7EG6_2(.din(n21801), .dout(n21804));
    jdff dff_B_11je3hXV5_2(.din(n21804), .dout(n21807));
    jdff dff_B_dNzfvh2j6_2(.din(n21807), .dout(n21810));
    jdff dff_B_ii4FWdKs3_2(.din(n21810), .dout(n21813));
    jdff dff_B_PMTWwnZD2_2(.din(n21813), .dout(n21816));
    jdff dff_B_2R7uQTqB7_2(.din(n21816), .dout(n21819));
    jdff dff_B_Jyz2QApv5_2(.din(n21819), .dout(n21822));
    jdff dff_B_JBIaOyn81_2(.din(n3207), .dout(n21825));
    jdff dff_B_yT5jobxk4_1(.din(n3027), .dout(n21828));
    jdff dff_B_7JAqNfso5_2(.din(n2648), .dout(n21831));
    jdff dff_B_retg5sal1_2(.din(n21831), .dout(n21834));
    jdff dff_B_A4vrtnSH3_2(.din(n21834), .dout(n21837));
    jdff dff_B_qlYry9lt8_2(.din(n21837), .dout(n21840));
    jdff dff_B_r1y2DTad6_2(.din(n21840), .dout(n21843));
    jdff dff_B_IpJS6Yjr3_2(.din(n21843), .dout(n21846));
    jdff dff_B_aSytTE3v5_2(.din(n21846), .dout(n21849));
    jdff dff_B_eA3eVsOS5_2(.din(n21849), .dout(n21852));
    jdff dff_B_NmyyoUbH7_2(.din(n21852), .dout(n21855));
    jdff dff_B_N30qgxtY5_2(.din(n21855), .dout(n21858));
    jdff dff_B_sBD5fOAS7_2(.din(n21858), .dout(n21861));
    jdff dff_B_ROiWYELl3_2(.din(n21861), .dout(n21864));
    jdff dff_B_JwGCPUiN1_2(.din(n21864), .dout(n21867));
    jdff dff_B_QP6oDmvm3_2(.din(n21867), .dout(n21870));
    jdff dff_B_IrJyoUG20_2(.din(n21870), .dout(n21873));
    jdff dff_B_Vh5xl8JH8_2(.din(n21873), .dout(n21876));
    jdff dff_B_uhyn0yt57_2(.din(n21876), .dout(n21879));
    jdff dff_B_8vJAl03n1_2(.din(n21879), .dout(n21882));
    jdff dff_B_3r6Rjrm44_2(.din(n21882), .dout(n21885));
    jdff dff_B_QJ1fA5oe5_2(.din(n21885), .dout(n21888));
    jdff dff_B_OBfPOlGw5_2(.din(n2812), .dout(n21891));
    jdff dff_B_Y00TVUep1_1(.din(n2652), .dout(n21894));
    jdff dff_B_GBVQ5kQi4_2(.din(n2297), .dout(n21897));
    jdff dff_B_emarn5hR8_2(.din(n21897), .dout(n21900));
    jdff dff_B_xo7lOydL0_2(.din(n21900), .dout(n21903));
    jdff dff_B_1y3bl1DT5_2(.din(n21903), .dout(n21906));
    jdff dff_B_S8pJRnZ08_2(.din(n21906), .dout(n21909));
    jdff dff_B_zyBgXcK69_2(.din(n21909), .dout(n21912));
    jdff dff_B_2l6JgLO20_2(.din(n21912), .dout(n21915));
    jdff dff_B_vvGstb3u6_2(.din(n21915), .dout(n21918));
    jdff dff_B_Ojxe2w5V1_2(.din(n21918), .dout(n21921));
    jdff dff_B_NJQC5RLN1_2(.din(n21921), .dout(n21924));
    jdff dff_B_xkyLc5QC5_2(.din(n21924), .dout(n21927));
    jdff dff_B_g4Xk05fy1_2(.din(n21927), .dout(n21930));
    jdff dff_B_LojWqOlZ3_2(.din(n21930), .dout(n21933));
    jdff dff_B_B9DS5n4x2_2(.din(n21933), .dout(n21936));
    jdff dff_B_UzAZefYP7_2(.din(n21936), .dout(n21939));
    jdff dff_B_zRtuluKM3_2(.din(n21939), .dout(n21942));
    jdff dff_B_uqRp0sXY8_2(.din(n21942), .dout(n21945));
    jdff dff_B_dnBmfhxP0_2(.din(n2434), .dout(n21948));
    jdff dff_B_3HGlLHHK0_1(.din(n2301), .dout(n21951));
    jdff dff_B_YfSYz0J25_2(.din(n1973), .dout(n21954));
    jdff dff_B_zRZmOvmZ9_2(.din(n21954), .dout(n21957));
    jdff dff_B_vHLmVdCp7_2(.din(n21957), .dout(n21960));
    jdff dff_B_WeDC8Aqf4_2(.din(n21960), .dout(n21963));
    jdff dff_B_pCDmsHui1_2(.din(n21963), .dout(n21966));
    jdff dff_B_A5EVWbOE0_2(.din(n21966), .dout(n21969));
    jdff dff_B_ygM08s7E1_2(.din(n21969), .dout(n21972));
    jdff dff_B_IIZZ6ubz3_2(.din(n21972), .dout(n21975));
    jdff dff_B_rCEn5z0B8_2(.din(n21975), .dout(n21978));
    jdff dff_B_Xo7uSpIc3_2(.din(n21978), .dout(n21981));
    jdff dff_B_AUIvz5kU7_2(.din(n21981), .dout(n21984));
    jdff dff_B_6J6Zapwv8_2(.din(n21984), .dout(n21987));
    jdff dff_B_Qds8q9tS3_2(.din(n21987), .dout(n21990));
    jdff dff_B_3uAKOUMy2_2(.din(n21990), .dout(n21993));
    jdff dff_B_aW03qvsr3_2(.din(n2083), .dout(n21996));
    jdff dff_B_5W1HNHhA0_1(.din(n1977), .dout(n21999));
    jdff dff_B_zeqJF3l42_2(.din(n1676), .dout(n22002));
    jdff dff_B_EX0KBTux0_2(.din(n22002), .dout(n22005));
    jdff dff_B_40DQ05gC1_2(.din(n22005), .dout(n22008));
    jdff dff_B_ispNmflQ4_2(.din(n22008), .dout(n22011));
    jdff dff_B_SUYk7Gpm9_2(.din(n22011), .dout(n22014));
    jdff dff_B_0wiadfvI9_2(.din(n22014), .dout(n22017));
    jdff dff_B_wCwrZ7sT0_2(.din(n22017), .dout(n22020));
    jdff dff_B_Ez6ZSNkI5_2(.din(n22020), .dout(n22023));
    jdff dff_B_9qG03qPU5_2(.din(n22023), .dout(n22026));
    jdff dff_B_lFuhzVqH5_2(.din(n22026), .dout(n22029));
    jdff dff_B_YFOUAA3M5_2(.din(n22029), .dout(n22032));
    jdff dff_B_H0YJAthz5_2(.din(n1759), .dout(n22035));
    jdff dff_B_TG7ggu479_1(.din(n1680), .dout(n22038));
    jdff dff_B_gICaoszp8_2(.din(n1406), .dout(n22041));
    jdff dff_B_AQ3BNbBd1_2(.din(n22041), .dout(n22044));
    jdff dff_B_LpODIpdX2_2(.din(n22044), .dout(n22047));
    jdff dff_B_qCK0mbns7_2(.din(n22047), .dout(n22050));
    jdff dff_B_yM5iZlxK9_2(.din(n22050), .dout(n22053));
    jdff dff_B_dE0RJCMY2_2(.din(n22053), .dout(n22056));
    jdff dff_B_BnSvBPJn0_2(.din(n22056), .dout(n22059));
    jdff dff_B_a5JaWE737_2(.din(n22059), .dout(n22062));
    jdff dff_B_StYRvpWz0_2(.din(n1462), .dout(n22065));
    jdff dff_B_xBcKVmxU9_2(.din(n22065), .dout(n22068));
    jdff dff_B_Baav93bQ4_2(.din(n22068), .dout(n22071));
    jdff dff_B_Cecb2C139_1(.din(n1410), .dout(n22074));
    jdff dff_B_LhXZKNt04_1(.din(n22074), .dout(n22077));
    jdff dff_B_GQQ7GrVa6_2(.din(n1169), .dout(n22080));
    jdff dff_B_tssskMr49_2(.din(n22080), .dout(n22083));
    jdff dff_B_XzIhFrPZ0_2(.din(n22083), .dout(n22086));
    jdff dff_B_wHOweIil2_0(.din(n1188), .dout(n22089));
    jdff dff_A_kPRBdduK3_0(.din(n22094), .dout(n22091));
    jdff dff_A_hmDCpiYY5_0(.din(n945), .dout(n22094));
    jdff dff_A_ONStMVIT2_1(.din(n22100), .dout(n22097));
    jdff dff_A_Cqil93OE8_1(.din(n945), .dout(n22100));
    jdff dff_B_tH64gZ2p2_1(.din(n5906), .dout(n22104));
    jdff dff_B_vsBkSVvQ9_2(.din(n5681), .dout(n22107));
    jdff dff_B_YDKIcx736_2(.din(n22107), .dout(n22110));
    jdff dff_B_wiQ12gCq0_2(.din(n22110), .dout(n22113));
    jdff dff_B_bc7mP5u12_2(.din(n22113), .dout(n22116));
    jdff dff_B_pJwiY3L16_2(.din(n22116), .dout(n22119));
    jdff dff_B_CfVTyzbr7_2(.din(n22119), .dout(n22122));
    jdff dff_B_3nC7AJco0_2(.din(n22122), .dout(n22125));
    jdff dff_B_z5Zy6f9Q3_2(.din(n22125), .dout(n22128));
    jdff dff_B_JiiRaLyT6_2(.din(n22128), .dout(n22131));
    jdff dff_B_dWWWBkCr0_2(.din(n22131), .dout(n22134));
    jdff dff_B_hVJNX2qw9_2(.din(n22134), .dout(n22137));
    jdff dff_B_8JGAj5iT2_2(.din(n22137), .dout(n22140));
    jdff dff_B_b6KKmoqP2_2(.din(n22140), .dout(n22143));
    jdff dff_B_p2xCU6m46_2(.din(n22143), .dout(n22146));
    jdff dff_B_uJrcZC8F0_2(.din(n22146), .dout(n22149));
    jdff dff_B_g1fcwlwt0_2(.din(n22149), .dout(n22152));
    jdff dff_B_gBggXZDR0_2(.din(n22152), .dout(n22155));
    jdff dff_B_qYAFNbPN4_2(.din(n22155), .dout(n22158));
    jdff dff_B_LXBC5JLy0_2(.din(n22158), .dout(n22161));
    jdff dff_B_BEpY2dra0_2(.din(n22161), .dout(n22164));
    jdff dff_B_oNRq0rgT5_2(.din(n22164), .dout(n22167));
    jdff dff_B_FUrM4H2e0_2(.din(n22167), .dout(n22170));
    jdff dff_B_hE4UHJNO5_2(.din(n22170), .dout(n22173));
    jdff dff_B_XpKPpW862_2(.din(n22173), .dout(n22176));
    jdff dff_B_Pukwssw95_2(.din(n22176), .dout(n22179));
    jdff dff_B_iDh9LQAv8_2(.din(n22179), .dout(n22182));
    jdff dff_B_zZ0kqyn91_2(.din(n22182), .dout(n22185));
    jdff dff_B_91ISSEBv4_2(.din(n22185), .dout(n22188));
    jdff dff_B_qPa29pS04_2(.din(n22188), .dout(n22191));
    jdff dff_B_kfwyd9nP9_2(.din(n22191), .dout(n22194));
    jdff dff_B_yrxVOoOE8_2(.din(n22194), .dout(n22197));
    jdff dff_B_AY7lYIUV9_2(.din(n22197), .dout(n22200));
    jdff dff_B_mrrtY6pt7_2(.din(n22200), .dout(n22203));
    jdff dff_B_LKQUuxjj8_2(.din(n22203), .dout(n22206));
    jdff dff_B_1kTDukAs5_2(.din(n22206), .dout(n22209));
    jdff dff_B_hUXzn7KH6_2(.din(n22209), .dout(n22212));
    jdff dff_B_njlmG7O59_2(.din(n22212), .dout(n22215));
    jdff dff_B_POyDQKv68_2(.din(n22215), .dout(n22218));
    jdff dff_B_4EvScwfw9_2(.din(n22218), .dout(n22221));
    jdff dff_B_Th3njhLC2_2(.din(n22221), .dout(n22224));
    jdff dff_B_w1gSjeAf4_2(.din(n22224), .dout(n22227));
    jdff dff_B_OsKlf9aE8_2(.din(n22227), .dout(n22230));
    jdff dff_B_2lysxwuL8_2(.din(n22230), .dout(n22233));
    jdff dff_B_NUZsT6f97_2(.din(n22233), .dout(n22236));
    jdff dff_B_ulbJp4165_2(.din(n22236), .dout(n22239));
    jdff dff_B_ERHUrecI3_2(.din(n22239), .dout(n22242));
    jdff dff_B_gnw9YzMm7_0(.din(n5902), .dout(n22245));
    jdff dff_A_0VYyg8st6_1(.din(n5859), .dout(n22247));
    jdff dff_B_mEub8Cht3_1(.din(n5685), .dout(n22251));
    jdff dff_B_04aaA9Pj2_2(.din(n5436), .dout(n22254));
    jdff dff_B_uGPEyDWy3_2(.din(n22254), .dout(n22257));
    jdff dff_B_Jw4gCK698_2(.din(n22257), .dout(n22260));
    jdff dff_B_4MHLehCB7_2(.din(n22260), .dout(n22263));
    jdff dff_B_mho9pv3N5_2(.din(n22263), .dout(n22266));
    jdff dff_B_9cKZPClz3_2(.din(n22266), .dout(n22269));
    jdff dff_B_aL7DujUi5_2(.din(n22269), .dout(n22272));
    jdff dff_B_WNed0ixx4_2(.din(n22272), .dout(n22275));
    jdff dff_B_RlHJfAZj3_2(.din(n22275), .dout(n22278));
    jdff dff_B_OXey3Q4g5_2(.din(n22278), .dout(n22281));
    jdff dff_B_Fb4TIpvM9_2(.din(n22281), .dout(n22284));
    jdff dff_B_hvDhxpSV8_2(.din(n22284), .dout(n22287));
    jdff dff_B_IlmlciXJ9_2(.din(n22287), .dout(n22290));
    jdff dff_B_NU3PDFub9_2(.din(n22290), .dout(n22293));
    jdff dff_B_kjDWGwKC5_2(.din(n22293), .dout(n22296));
    jdff dff_B_5EXv2p1d4_2(.din(n22296), .dout(n22299));
    jdff dff_B_f1JfoURg7_2(.din(n22299), .dout(n22302));
    jdff dff_B_VRDgX8f18_2(.din(n22302), .dout(n22305));
    jdff dff_B_GZkdl9En5_2(.din(n22305), .dout(n22308));
    jdff dff_B_I8KzF8wc2_2(.din(n22308), .dout(n22311));
    jdff dff_B_gaRqe6bL1_2(.din(n22311), .dout(n22314));
    jdff dff_B_kkHFDaT97_2(.din(n22314), .dout(n22317));
    jdff dff_B_SLCXx6yq3_2(.din(n22317), .dout(n22320));
    jdff dff_B_CIHttLD85_2(.din(n22320), .dout(n22323));
    jdff dff_B_LAMs7jrJ3_2(.din(n22323), .dout(n22326));
    jdff dff_B_Qp8Tv7Y91_2(.din(n22326), .dout(n22329));
    jdff dff_B_oeu70c2d3_2(.din(n22329), .dout(n22332));
    jdff dff_B_QyTblDHL5_2(.din(n22332), .dout(n22335));
    jdff dff_B_YqwMphmv2_2(.din(n22335), .dout(n22338));
    jdff dff_B_pC1cg0cG3_2(.din(n22338), .dout(n22341));
    jdff dff_B_D3KQpFdg0_2(.din(n22341), .dout(n22344));
    jdff dff_B_gDvfvCPO2_2(.din(n22344), .dout(n22347));
    jdff dff_B_zJAf4Cmw7_2(.din(n22347), .dout(n22350));
    jdff dff_B_IpZCzPRt6_2(.din(n22350), .dout(n22353));
    jdff dff_B_en0pEEKL1_2(.din(n22353), .dout(n22356));
    jdff dff_B_wsaxXHHs7_2(.din(n22356), .dout(n22359));
    jdff dff_B_IUhOhLE62_2(.din(n22359), .dout(n22362));
    jdff dff_B_jTOsY1Br4_2(.din(n22362), .dout(n22365));
    jdff dff_B_t6m14mr58_2(.din(n22365), .dout(n22368));
    jdff dff_B_7I4L68L81_2(.din(n22368), .dout(n22371));
    jdff dff_B_q3UgyzgI7_2(.din(n22371), .dout(n22374));
    jdff dff_B_LidCqk3d7_2(.din(n5614), .dout(n22377));
    jdff dff_B_0Um9Rg9s4_1(.din(n5440), .dout(n22380));
    jdff dff_B_FYeqss1r8_2(.din(n5164), .dout(n22383));
    jdff dff_B_0W5GxR8j8_2(.din(n22383), .dout(n22386));
    jdff dff_B_NEVodtvL7_2(.din(n22386), .dout(n22389));
    jdff dff_B_dS7nhfoN4_2(.din(n22389), .dout(n22392));
    jdff dff_B_DxMaCaeA6_2(.din(n22392), .dout(n22395));
    jdff dff_B_4DuoXHBK1_2(.din(n22395), .dout(n22398));
    jdff dff_B_xnHIWkkX9_2(.din(n22398), .dout(n22401));
    jdff dff_B_OguhmY5w5_2(.din(n22401), .dout(n22404));
    jdff dff_B_lrRq2WNd1_2(.din(n22404), .dout(n22407));
    jdff dff_B_LUS16xPf8_2(.din(n22407), .dout(n22410));
    jdff dff_B_0c9zDrv27_2(.din(n22410), .dout(n22413));
    jdff dff_B_2lR4bZBX6_2(.din(n22413), .dout(n22416));
    jdff dff_B_KgCCofJ52_2(.din(n22416), .dout(n22419));
    jdff dff_B_VJZliVqm8_2(.din(n22419), .dout(n22422));
    jdff dff_B_pbKSCjGs5_2(.din(n22422), .dout(n22425));
    jdff dff_B_XnRPovyT7_2(.din(n22425), .dout(n22428));
    jdff dff_B_u0kxdFDU7_2(.din(n22428), .dout(n22431));
    jdff dff_B_MNcbHyEE3_2(.din(n22431), .dout(n22434));
    jdff dff_B_Q4OwdjlL3_2(.din(n22434), .dout(n22437));
    jdff dff_B_o4bAO1UA8_2(.din(n22437), .dout(n22440));
    jdff dff_B_bBxnxwqF7_2(.din(n22440), .dout(n22443));
    jdff dff_B_nCngdcef7_2(.din(n22443), .dout(n22446));
    jdff dff_B_b1sbFnIp3_2(.din(n22446), .dout(n22449));
    jdff dff_B_Z51BpY3j1_2(.din(n22449), .dout(n22452));
    jdff dff_B_g0EJDHDJ5_2(.din(n22452), .dout(n22455));
    jdff dff_B_4gtwUJOe7_2(.din(n22455), .dout(n22458));
    jdff dff_B_XGXJ9S162_2(.din(n22458), .dout(n22461));
    jdff dff_B_lqSVTLqO9_2(.din(n22461), .dout(n22464));
    jdff dff_B_1ccNLfBt2_2(.din(n22464), .dout(n22467));
    jdff dff_B_ySeAm6lW3_2(.din(n22467), .dout(n22470));
    jdff dff_B_Tma7Mkyr4_2(.din(n22470), .dout(n22473));
    jdff dff_B_ry4mptlp7_2(.din(n22473), .dout(n22476));
    jdff dff_B_Y7zLzYTy3_2(.din(n22476), .dout(n22479));
    jdff dff_B_20eYAsih1_2(.din(n22479), .dout(n22482));
    jdff dff_B_WyUNR5Ew3_2(.din(n22482), .dout(n22485));
    jdff dff_B_P6uXQ72v4_2(.din(n22485), .dout(n22488));
    jdff dff_B_oSg6BDzv9_2(.din(n22488), .dout(n22491));
    jdff dff_B_i3Ve0M2d3_2(.din(n22491), .dout(n22494));
    jdff dff_B_389B8GSI6_2(.din(n5342), .dout(n22497));
    jdff dff_B_EEFDNy893_1(.din(n5168), .dout(n22500));
    jdff dff_B_9McnlYsm1_2(.din(n4865), .dout(n22503));
    jdff dff_B_pKf1HR1x4_2(.din(n22503), .dout(n22506));
    jdff dff_B_ZzQzMXrZ2_2(.din(n22506), .dout(n22509));
    jdff dff_B_rFb84YWB2_2(.din(n22509), .dout(n22512));
    jdff dff_B_7nHviEfH9_2(.din(n22512), .dout(n22515));
    jdff dff_B_81ooFWeb5_2(.din(n22515), .dout(n22518));
    jdff dff_B_YoHzIqbB8_2(.din(n22518), .dout(n22521));
    jdff dff_B_1ydIIUHn3_2(.din(n22521), .dout(n22524));
    jdff dff_B_s5ig4Y2j8_2(.din(n22524), .dout(n22527));
    jdff dff_B_rNt2kuqR7_2(.din(n22527), .dout(n22530));
    jdff dff_B_CgeR1ohU2_2(.din(n22530), .dout(n22533));
    jdff dff_B_0kXB4qhL2_2(.din(n22533), .dout(n22536));
    jdff dff_B_KB8LWmM05_2(.din(n22536), .dout(n22539));
    jdff dff_B_WiRQ99eB1_2(.din(n22539), .dout(n22542));
    jdff dff_B_suPLVpzt2_2(.din(n22542), .dout(n22545));
    jdff dff_B_XNBJe3SD3_2(.din(n22545), .dout(n22548));
    jdff dff_B_2Jcdb9cm1_2(.din(n22548), .dout(n22551));
    jdff dff_B_SxIBpEx52_2(.din(n22551), .dout(n22554));
    jdff dff_B_xp7BD0NP4_2(.din(n22554), .dout(n22557));
    jdff dff_B_fKc2By9A8_2(.din(n22557), .dout(n22560));
    jdff dff_B_x1gpd9tU7_2(.din(n22560), .dout(n22563));
    jdff dff_B_KWAnneZX5_2(.din(n22563), .dout(n22566));
    jdff dff_B_pK1bjzOe0_2(.din(n22566), .dout(n22569));
    jdff dff_B_qKvLM4Iq3_2(.din(n22569), .dout(n22572));
    jdff dff_B_nhlIYQLz9_2(.din(n22572), .dout(n22575));
    jdff dff_B_JB3bG6Ez7_2(.din(n22575), .dout(n22578));
    jdff dff_B_rE2btYBL6_2(.din(n22578), .dout(n22581));
    jdff dff_B_jamFC7LZ3_2(.din(n22581), .dout(n22584));
    jdff dff_B_4FG32wZ97_2(.din(n22584), .dout(n22587));
    jdff dff_B_sh2kcuiY3_2(.din(n22587), .dout(n22590));
    jdff dff_B_Cwv5OEyC3_2(.din(n22590), .dout(n22593));
    jdff dff_B_E6RTjQmc2_2(.din(n22593), .dout(n22596));
    jdff dff_B_b5uOftRa7_2(.din(n22596), .dout(n22599));
    jdff dff_B_m4B0bsaM0_2(.din(n22599), .dout(n22602));
    jdff dff_B_sJDrkbVR3_2(.din(n22602), .dout(n22605));
    jdff dff_B_IP2xz7gk6_2(.din(n5043), .dout(n22608));
    jdff dff_B_8fyuWS3C8_1(.din(n4869), .dout(n22611));
    jdff dff_B_CZ4lnBnU4_2(.din(n4539), .dout(n22614));
    jdff dff_B_uJTWmKKg9_2(.din(n22614), .dout(n22617));
    jdff dff_B_W8kdiqNn7_2(.din(n22617), .dout(n22620));
    jdff dff_B_DMpF30di2_2(.din(n22620), .dout(n22623));
    jdff dff_B_jObhIa4m8_2(.din(n22623), .dout(n22626));
    jdff dff_B_DkXtiUhh5_2(.din(n22626), .dout(n22629));
    jdff dff_B_3AZzWK5K9_2(.din(n22629), .dout(n22632));
    jdff dff_B_RB8EGyzc3_2(.din(n22632), .dout(n22635));
    jdff dff_B_2Rkc27738_2(.din(n22635), .dout(n22638));
    jdff dff_B_8bct5HR39_2(.din(n22638), .dout(n22641));
    jdff dff_B_TTeqG0FQ9_2(.din(n22641), .dout(n22644));
    jdff dff_B_blGsaODc0_2(.din(n22644), .dout(n22647));
    jdff dff_B_dC8F7YR52_2(.din(n22647), .dout(n22650));
    jdff dff_B_0CWn7SjJ2_2(.din(n22650), .dout(n22653));
    jdff dff_B_nwh0I2Wz3_2(.din(n22653), .dout(n22656));
    jdff dff_B_RUdayj0h1_2(.din(n22656), .dout(n22659));
    jdff dff_B_0taMoH0W1_2(.din(n22659), .dout(n22662));
    jdff dff_B_N06HOcfl0_2(.din(n22662), .dout(n22665));
    jdff dff_B_S6kSeQDQ7_2(.din(n22665), .dout(n22668));
    jdff dff_B_TnDkHids0_2(.din(n22668), .dout(n22671));
    jdff dff_B_QcMnnVQb5_2(.din(n22671), .dout(n22674));
    jdff dff_B_LZyd5xTg3_2(.din(n22674), .dout(n22677));
    jdff dff_B_jpyCYVHf7_2(.din(n22677), .dout(n22680));
    jdff dff_B_clxmQnR12_2(.din(n22680), .dout(n22683));
    jdff dff_B_tSSBfNa53_2(.din(n22683), .dout(n22686));
    jdff dff_B_EMA8cHjx2_2(.din(n22686), .dout(n22689));
    jdff dff_B_vPuxReyu7_2(.din(n22689), .dout(n22692));
    jdff dff_B_WpTXQUJm7_2(.din(n22692), .dout(n22695));
    jdff dff_B_ZwD6HCR57_2(.din(n22695), .dout(n22698));
    jdff dff_B_ywKQgdwa4_2(.din(n22698), .dout(n22701));
    jdff dff_B_j0Buq58s5_2(.din(n22701), .dout(n22704));
    jdff dff_B_yeqhcbgU8_2(.din(n22704), .dout(n22707));
    jdff dff_B_rRpQxRXk6_2(.din(n4717), .dout(n22710));
    jdff dff_B_CsyphyLd6_1(.din(n4543), .dout(n22713));
    jdff dff_B_hwIpHyGz5_2(.din(n4189), .dout(n22716));
    jdff dff_B_JaLNPF1R5_2(.din(n22716), .dout(n22719));
    jdff dff_B_Zoz5qMIX0_2(.din(n22719), .dout(n22722));
    jdff dff_B_3WYuB6Xe5_2(.din(n22722), .dout(n22725));
    jdff dff_B_O26byoBL3_2(.din(n22725), .dout(n22728));
    jdff dff_B_Wq22OHV66_2(.din(n22728), .dout(n22731));
    jdff dff_B_OMek1LYa7_2(.din(n22731), .dout(n22734));
    jdff dff_B_umbRiCSr6_2(.din(n22734), .dout(n22737));
    jdff dff_B_rLrmj8R86_2(.din(n22737), .dout(n22740));
    jdff dff_B_TGZvNaf38_2(.din(n22740), .dout(n22743));
    jdff dff_B_L6VddQaT1_2(.din(n22743), .dout(n22746));
    jdff dff_B_IeuTQqpa0_2(.din(n22746), .dout(n22749));
    jdff dff_B_bMmCb6Ng6_2(.din(n22749), .dout(n22752));
    jdff dff_B_3ObcaEG11_2(.din(n22752), .dout(n22755));
    jdff dff_B_1Nz5Iy0p0_2(.din(n22755), .dout(n22758));
    jdff dff_B_I8eRL6Ot3_2(.din(n22758), .dout(n22761));
    jdff dff_B_tlWbOF6S3_2(.din(n22761), .dout(n22764));
    jdff dff_B_JkJ5zbY76_2(.din(n22764), .dout(n22767));
    jdff dff_B_vJoA67bg3_2(.din(n22767), .dout(n22770));
    jdff dff_B_8zk7mE1u7_2(.din(n22770), .dout(n22773));
    jdff dff_B_4XKKqanO3_2(.din(n22773), .dout(n22776));
    jdff dff_B_4rGBuJul6_2(.din(n22776), .dout(n22779));
    jdff dff_B_bEemoxrx1_2(.din(n22779), .dout(n22782));
    jdff dff_B_xrQzQvAZ3_2(.din(n22782), .dout(n22785));
    jdff dff_B_gtHlNTOL7_2(.din(n22785), .dout(n22788));
    jdff dff_B_mwnWALYY4_2(.din(n22788), .dout(n22791));
    jdff dff_B_6rzBcZzE7_2(.din(n22791), .dout(n22794));
    jdff dff_B_eGjzVzzH4_2(.din(n22794), .dout(n22797));
    jdff dff_B_95Ba9HeD1_2(.din(n22797), .dout(n22800));
    jdff dff_B_Hv6YVCsr6_2(.din(n4367), .dout(n22803));
    jdff dff_B_LQq7XSgV1_1(.din(n4193), .dout(n22806));
    jdff dff_B_vcJIzG6e5_2(.din(n3813), .dout(n22809));
    jdff dff_B_KyAy0u7z2_2(.din(n22809), .dout(n22812));
    jdff dff_B_bwFVgsCd8_2(.din(n22812), .dout(n22815));
    jdff dff_B_ryv10emY7_2(.din(n22815), .dout(n22818));
    jdff dff_B_QLutS9cy4_2(.din(n22818), .dout(n22821));
    jdff dff_B_v9840jYK1_2(.din(n22821), .dout(n22824));
    jdff dff_B_BrCgUxQT1_2(.din(n22824), .dout(n22827));
    jdff dff_B_93aRqduI4_2(.din(n22827), .dout(n22830));
    jdff dff_B_PNnW47wB3_2(.din(n22830), .dout(n22833));
    jdff dff_B_rbEFlcNa3_2(.din(n22833), .dout(n22836));
    jdff dff_B_wvnIlnOQ6_2(.din(n22836), .dout(n22839));
    jdff dff_B_Dr87KwPU9_2(.din(n22839), .dout(n22842));
    jdff dff_B_iVVXmieo7_2(.din(n22842), .dout(n22845));
    jdff dff_B_XlvhNH716_2(.din(n22845), .dout(n22848));
    jdff dff_B_AgCiMPqe9_2(.din(n22848), .dout(n22851));
    jdff dff_B_7texvTvg8_2(.din(n22851), .dout(n22854));
    jdff dff_B_hYW46rO79_2(.din(n22854), .dout(n22857));
    jdff dff_B_tfZRLX5F1_2(.din(n22857), .dout(n22860));
    jdff dff_B_fdfRDlZi0_2(.din(n22860), .dout(n22863));
    jdff dff_B_KkekWbYD4_2(.din(n22863), .dout(n22866));
    jdff dff_B_DA453B0D7_2(.din(n22866), .dout(n22869));
    jdff dff_B_Tsr0aNow7_2(.din(n22869), .dout(n22872));
    jdff dff_B_bbOFfDPy5_2(.din(n22872), .dout(n22875));
    jdff dff_B_XGlQejHS2_2(.din(n22875), .dout(n22878));
    jdff dff_B_tpqpxOud6_2(.din(n22878), .dout(n22881));
    jdff dff_B_NgZUA2VO6_2(.din(n22881), .dout(n22884));
    jdff dff_B_a8DfgMyJ2_2(.din(n3987), .dout(n22887));
    jdff dff_B_VQ99M6Cp9_1(.din(n3817), .dout(n22890));
    jdff dff_B_fLOEm6OU5_2(.din(n3433), .dout(n22893));
    jdff dff_B_b7EgqpGf5_2(.din(n22893), .dout(n22896));
    jdff dff_B_IsKYsYA35_2(.din(n22896), .dout(n22899));
    jdff dff_B_mmaiWdOm9_2(.din(n22899), .dout(n22902));
    jdff dff_B_uifbmBo90_2(.din(n22902), .dout(n22905));
    jdff dff_B_VPp2sZDf3_2(.din(n22905), .dout(n22908));
    jdff dff_B_qSggmim50_2(.din(n22908), .dout(n22911));
    jdff dff_B_mvAoWqJI4_2(.din(n22911), .dout(n22914));
    jdff dff_B_QYgGxJNT9_2(.din(n22914), .dout(n22917));
    jdff dff_B_OjC2kcUA2_2(.din(n22917), .dout(n22920));
    jdff dff_B_ihnlVSrx3_2(.din(n22920), .dout(n22923));
    jdff dff_B_MMmXR79t3_2(.din(n22923), .dout(n22926));
    jdff dff_B_YZu4mbko4_2(.din(n22926), .dout(n22929));
    jdff dff_B_R2YHob0V1_2(.din(n22929), .dout(n22932));
    jdff dff_B_HGKn9FQW3_2(.din(n22932), .dout(n22935));
    jdff dff_B_KHbhU1An3_2(.din(n22935), .dout(n22938));
    jdff dff_B_dfrDS8QZ4_2(.din(n22938), .dout(n22941));
    jdff dff_B_VpsGrLNj7_2(.din(n22941), .dout(n22944));
    jdff dff_B_1iysCM1M1_2(.din(n22944), .dout(n22947));
    jdff dff_B_dbbJhbRE7_2(.din(n22947), .dout(n22950));
    jdff dff_B_m9jNYSza4_2(.din(n22950), .dout(n22953));
    jdff dff_B_fYo9iQxr0_2(.din(n22953), .dout(n22956));
    jdff dff_B_AJ278F735_2(.din(n22956), .dout(n22959));
    jdff dff_B_6UGA7hQZ1_2(.din(n3604), .dout(n22962));
    jdff dff_B_0oMYSq0L6_1(.din(n3437), .dout(n22965));
    jdff dff_B_loGNozgi9_2(.din(n3042), .dout(n22968));
    jdff dff_B_WwYCtl412_2(.din(n22968), .dout(n22971));
    jdff dff_B_0n1Jadz66_2(.din(n22971), .dout(n22974));
    jdff dff_B_PVehoIcG1_2(.din(n22974), .dout(n22977));
    jdff dff_B_vgegI7jV3_2(.din(n22977), .dout(n22980));
    jdff dff_B_1Pkxkatc6_2(.din(n22980), .dout(n22983));
    jdff dff_B_8YPRvzTG9_2(.din(n22983), .dout(n22986));
    jdff dff_B_5BL8usaY8_2(.din(n22986), .dout(n22989));
    jdff dff_B_5Wt5ibDr7_2(.din(n22989), .dout(n22992));
    jdff dff_B_HGp057y16_2(.din(n22992), .dout(n22995));
    jdff dff_B_N3HA4PbK2_2(.din(n22995), .dout(n22998));
    jdff dff_B_YP7WalGR7_2(.din(n22998), .dout(n23001));
    jdff dff_B_xXCczbKI4_2(.din(n23001), .dout(n23004));
    jdff dff_B_GG2LoV179_2(.din(n23004), .dout(n23007));
    jdff dff_B_7rTj1hxk0_2(.din(n23007), .dout(n23010));
    jdff dff_B_CU0GAnsS0_2(.din(n23010), .dout(n23013));
    jdff dff_B_lOPgQupd8_2(.din(n23013), .dout(n23016));
    jdff dff_B_r7yNn4561_2(.din(n23016), .dout(n23019));
    jdff dff_B_U5REUEV02_2(.din(n23019), .dout(n23022));
    jdff dff_B_nKiBMnI58_2(.din(n23022), .dout(n23025));
    jdff dff_B_OuUO3ksH5_2(.din(n3199), .dout(n23028));
    jdff dff_B_ze7CwRxD5_1(.din(n3046), .dout(n23031));
    jdff dff_B_t2qiqlq82_2(.din(n2667), .dout(n23034));
    jdff dff_B_hO8a1Kat6_2(.din(n23034), .dout(n23037));
    jdff dff_B_vIvEHoZA5_2(.din(n23037), .dout(n23040));
    jdff dff_B_M4VIBpVI8_2(.din(n23040), .dout(n23043));
    jdff dff_B_rie1OaCW6_2(.din(n23043), .dout(n23046));
    jdff dff_B_Q64ShAcO6_2(.din(n23046), .dout(n23049));
    jdff dff_B_0aDQFoDM4_2(.din(n23049), .dout(n23052));
    jdff dff_B_LU8Dum5u8_2(.din(n23052), .dout(n23055));
    jdff dff_B_cM3drlQI4_2(.din(n23055), .dout(n23058));
    jdff dff_B_Vl92Qsgo9_2(.din(n23058), .dout(n23061));
    jdff dff_B_uEBfFmQA5_2(.din(n23061), .dout(n23064));
    jdff dff_B_1JArMmMc1_2(.din(n23064), .dout(n23067));
    jdff dff_B_i5U1hvRO7_2(.din(n23067), .dout(n23070));
    jdff dff_B_SGnsI4oE7_2(.din(n23070), .dout(n23073));
    jdff dff_B_zEE62LWO5_2(.din(n23073), .dout(n23076));
    jdff dff_B_Y9rOaHPJ9_2(.din(n23076), .dout(n23079));
    jdff dff_B_XlNQGqbr8_2(.din(n23079), .dout(n23082));
    jdff dff_B_5kYk2Ixa5_2(.din(n2804), .dout(n23085));
    jdff dff_B_yZ1ZLZMX3_1(.din(n2671), .dout(n23088));
    jdff dff_B_9aoLueLy1_2(.din(n2316), .dout(n23091));
    jdff dff_B_NKCKydGn2_2(.din(n23091), .dout(n23094));
    jdff dff_B_EnS2MZHq4_2(.din(n23094), .dout(n23097));
    jdff dff_B_H4nkGOZq9_2(.din(n23097), .dout(n23100));
    jdff dff_B_I65d36uz4_2(.din(n23100), .dout(n23103));
    jdff dff_B_ODDEud1P6_2(.din(n23103), .dout(n23106));
    jdff dff_B_YOraFkZV4_2(.din(n23106), .dout(n23109));
    jdff dff_B_Do3QMKhj3_2(.din(n23109), .dout(n23112));
    jdff dff_B_5ngNZ9rE4_2(.din(n23112), .dout(n23115));
    jdff dff_B_MMv7rcA25_2(.din(n23115), .dout(n23118));
    jdff dff_B_PfO4DHBQ4_2(.din(n23118), .dout(n23121));
    jdff dff_B_LksThUh49_2(.din(n23121), .dout(n23124));
    jdff dff_B_o4GO084i3_2(.din(n23124), .dout(n23127));
    jdff dff_B_ZD8FogMh6_2(.din(n23127), .dout(n23130));
    jdff dff_B_YZpFnkvY4_2(.din(n2426), .dout(n23133));
    jdff dff_B_2TtZjgDR4_1(.din(n2320), .dout(n23136));
    jdff dff_B_Fjt8NB8M0_2(.din(n1992), .dout(n23139));
    jdff dff_B_u3Ye1c305_2(.din(n23139), .dout(n23142));
    jdff dff_B_gUTxaUXY9_2(.din(n23142), .dout(n23145));
    jdff dff_B_oevza0wB1_2(.din(n23145), .dout(n23148));
    jdff dff_B_a5k7dsn76_2(.din(n23148), .dout(n23151));
    jdff dff_B_jd9iXizh0_2(.din(n23151), .dout(n23154));
    jdff dff_B_Gg90a2hp3_2(.din(n23154), .dout(n23157));
    jdff dff_B_3CvsAI2d8_2(.din(n23157), .dout(n23160));
    jdff dff_B_yuFhykAK8_2(.din(n23160), .dout(n23163));
    jdff dff_B_7cHnDViy2_2(.din(n23163), .dout(n23166));
    jdff dff_B_hpCVcopu1_2(.din(n23166), .dout(n23169));
    jdff dff_B_N8xVdQVc1_2(.din(n2075), .dout(n23172));
    jdff dff_B_xDE2wZ4o5_1(.din(n1996), .dout(n23175));
    jdff dff_B_RVTKO89N5_2(.din(n1695), .dout(n23178));
    jdff dff_B_A9ghjFdp7_2(.din(n23178), .dout(n23181));
    jdff dff_B_WMQLPQZL3_2(.din(n23181), .dout(n23184));
    jdff dff_B_aFF7X2kQ6_2(.din(n23184), .dout(n23187));
    jdff dff_B_XU1FHgmb0_2(.din(n23187), .dout(n23190));
    jdff dff_B_DxLwwvlN7_2(.din(n23190), .dout(n23193));
    jdff dff_B_T9Gfyxhh1_2(.din(n23193), .dout(n23196));
    jdff dff_B_enx57Ify0_2(.din(n23196), .dout(n23199));
    jdff dff_B_NtmhkJ5H6_2(.din(n1751), .dout(n23202));
    jdff dff_B_s5WQ3C6t1_2(.din(n23202), .dout(n23205));
    jdff dff_B_HmdH1K3B2_2(.din(n23205), .dout(n23208));
    jdff dff_B_9yuZU2o59_1(.din(n1699), .dout(n23211));
    jdff dff_B_UTv53eIV5_1(.din(n23211), .dout(n23214));
    jdff dff_B_tWtgbXPF4_2(.din(n1431), .dout(n23217));
    jdff dff_B_ac57eWrJ6_2(.din(n23217), .dout(n23220));
    jdff dff_B_qT2GWI6i5_2(.din(n23220), .dout(n23223));
    jdff dff_B_tFhInTpS8_0(.din(n1450), .dout(n23226));
    jdff dff_A_Nr7FDlQy8_0(.din(n23231), .dout(n23228));
    jdff dff_A_ld5XHP2q6_0(.din(n1177), .dout(n23231));
    jdff dff_A_eYh6xHTD4_1(.din(n23237), .dout(n23234));
    jdff dff_A_iGOTVGdz2_1(.din(n1177), .dout(n23237));
    jdff dff_B_H4YrT5Qg7_2(.din(n6124), .dout(n23241));
    jdff dff_B_8u82OTEk1_1(.din(n6116), .dout(n23244));
    jdff dff_B_FGBf8jTf5_2(.din(n5918), .dout(n23247));
    jdff dff_B_U6B4oF6j0_2(.din(n23247), .dout(n23250));
    jdff dff_B_3fEIf1bE7_2(.din(n23250), .dout(n23253));
    jdff dff_B_yMlOjoPT8_2(.din(n23253), .dout(n23256));
    jdff dff_B_kCyg5rZc0_2(.din(n23256), .dout(n23259));
    jdff dff_B_ss9DrP9Y1_2(.din(n23259), .dout(n23262));
    jdff dff_B_dvk5yyze7_2(.din(n23262), .dout(n23265));
    jdff dff_B_4ywqs0yT2_2(.din(n23265), .dout(n23268));
    jdff dff_B_Gh7a08yD4_2(.din(n23268), .dout(n23271));
    jdff dff_B_JdaNaoCJ2_2(.din(n23271), .dout(n23274));
    jdff dff_B_pectrKqf5_2(.din(n23274), .dout(n23277));
    jdff dff_B_3R9HEZGO0_2(.din(n23277), .dout(n23280));
    jdff dff_B_9ygUsPbc1_2(.din(n23280), .dout(n23283));
    jdff dff_B_bOpPDq8M7_2(.din(n23283), .dout(n23286));
    jdff dff_B_Yj0muCWl6_2(.din(n23286), .dout(n23289));
    jdff dff_B_se3wxhWY6_2(.din(n23289), .dout(n23292));
    jdff dff_B_F3XBj8p07_2(.din(n23292), .dout(n23295));
    jdff dff_B_VVdkneR19_2(.din(n23295), .dout(n23298));
    jdff dff_B_LpBLNGRS6_2(.din(n23298), .dout(n23301));
    jdff dff_B_2VuZlde11_2(.din(n23301), .dout(n23304));
    jdff dff_B_nFCJ8jKP4_2(.din(n23304), .dout(n23307));
    jdff dff_B_KJT6IcWt6_2(.din(n23307), .dout(n23310));
    jdff dff_B_yRnuStW29_2(.din(n23310), .dout(n23313));
    jdff dff_B_f7ZKQCdD4_2(.din(n23313), .dout(n23316));
    jdff dff_B_cXNZhmIG1_2(.din(n23316), .dout(n23319));
    jdff dff_B_crvvGL4B9_2(.din(n23319), .dout(n23322));
    jdff dff_B_UhOpIEwD0_2(.din(n23322), .dout(n23325));
    jdff dff_B_ORNnKSAZ3_2(.din(n23325), .dout(n23328));
    jdff dff_B_O8kLOrDs2_2(.din(n23328), .dout(n23331));
    jdff dff_B_uDZeASMP8_2(.din(n23331), .dout(n23334));
    jdff dff_B_7PCcJPzQ8_2(.din(n23334), .dout(n23337));
    jdff dff_B_Wr61stAb9_2(.din(n23337), .dout(n23340));
    jdff dff_B_QiQR7aMu3_2(.din(n23340), .dout(n23343));
    jdff dff_B_i18PVtYj0_2(.din(n23343), .dout(n23346));
    jdff dff_B_CaZbuqti0_2(.din(n23346), .dout(n23349));
    jdff dff_B_KjIXxOAI4_2(.din(n23349), .dout(n23352));
    jdff dff_B_yNlJaCvY2_2(.din(n23352), .dout(n23355));
    jdff dff_B_0vT1vTWF3_2(.din(n23355), .dout(n23358));
    jdff dff_B_txootfBz2_2(.din(n23358), .dout(n23361));
    jdff dff_B_kNuXWdfu9_2(.din(n23361), .dout(n23364));
    jdff dff_B_detvEDeQ7_2(.din(n23364), .dout(n23367));
    jdff dff_B_sWByKdUo7_2(.din(n23367), .dout(n23370));
    jdff dff_B_2AclVfkZ8_2(.din(n23370), .dout(n23373));
    jdff dff_B_q3Jkis7o0_2(.din(n23373), .dout(n23376));
    jdff dff_B_Atz20Po82_2(.din(n23376), .dout(n23379));
    jdff dff_B_r2TRi9Mw7_2(.din(n23379), .dout(n23382));
    jdff dff_B_5fqpPpqw5_1(.din(n5922), .dout(n23385));
    jdff dff_B_QrfLMSFN7_2(.din(n5700), .dout(n23388));
    jdff dff_B_SwO2J2EG7_2(.din(n23388), .dout(n23391));
    jdff dff_B_Dhp19eWZ8_2(.din(n23391), .dout(n23394));
    jdff dff_B_oEFFDRTh8_2(.din(n23394), .dout(n23397));
    jdff dff_B_n4yAV2wC8_2(.din(n23397), .dout(n23400));
    jdff dff_B_3SGtO3pG8_2(.din(n23400), .dout(n23403));
    jdff dff_B_WPmYJb8g0_2(.din(n23403), .dout(n23406));
    jdff dff_B_vamdq46V0_2(.din(n23406), .dout(n23409));
    jdff dff_B_2c0lb1Bf7_2(.din(n23409), .dout(n23412));
    jdff dff_B_Sm94U7RC0_2(.din(n23412), .dout(n23415));
    jdff dff_B_tovPr3Gj6_2(.din(n23415), .dout(n23418));
    jdff dff_B_zPC9L6st9_2(.din(n23418), .dout(n23421));
    jdff dff_B_sTXdIzQA2_2(.din(n23421), .dout(n23424));
    jdff dff_B_x1NngZmO0_2(.din(n23424), .dout(n23427));
    jdff dff_B_azJUgKoO7_2(.din(n23427), .dout(n23430));
    jdff dff_B_u3P2LWv37_2(.din(n23430), .dout(n23433));
    jdff dff_B_cdPaMq575_2(.din(n23433), .dout(n23436));
    jdff dff_B_Zq5If9UR2_2(.din(n23436), .dout(n23439));
    jdff dff_B_w6kQEEtk9_2(.din(n23439), .dout(n23442));
    jdff dff_B_fbeGPNnm0_2(.din(n23442), .dout(n23445));
    jdff dff_B_BkEWtN9y7_2(.din(n23445), .dout(n23448));
    jdff dff_B_lvhUxNJ98_2(.din(n23448), .dout(n23451));
    jdff dff_B_ecqrKTUu2_2(.din(n23451), .dout(n23454));
    jdff dff_B_Y5dEumy19_2(.din(n23454), .dout(n23457));
    jdff dff_B_s2o6rmh26_2(.din(n23457), .dout(n23460));
    jdff dff_B_NMEG0RSD1_2(.din(n23460), .dout(n23463));
    jdff dff_B_JC3shGiu0_2(.din(n23463), .dout(n23466));
    jdff dff_B_pXr7CSBT4_2(.din(n23466), .dout(n23469));
    jdff dff_B_8w5qjcmb8_2(.din(n23469), .dout(n23472));
    jdff dff_B_z0CxYak16_2(.din(n23472), .dout(n23475));
    jdff dff_B_n8slCP0C6_2(.din(n23475), .dout(n23478));
    jdff dff_B_VT0uZWCC8_2(.din(n23478), .dout(n23481));
    jdff dff_B_bADfbBni1_2(.din(n23481), .dout(n23484));
    jdff dff_B_4BIGkTLY9_2(.din(n23484), .dout(n23487));
    jdff dff_B_4emyKrqa6_2(.din(n23487), .dout(n23490));
    jdff dff_B_m5RFnYi50_2(.din(n23490), .dout(n23493));
    jdff dff_B_HUgFLPur3_2(.din(n23493), .dout(n23496));
    jdff dff_B_a4usGJD99_2(.din(n23496), .dout(n23499));
    jdff dff_B_74qhYA3S4_2(.din(n23499), .dout(n23502));
    jdff dff_B_K35Yb9Sz9_2(.din(n23502), .dout(n23505));
    jdff dff_B_KK9cnNdY5_2(.din(n23505), .dout(n23508));
    jdff dff_B_qGDh7Zs29_2(.din(n5851), .dout(n23511));
    jdff dff_B_nhG2MuVO0_1(.din(n5704), .dout(n23514));
    jdff dff_B_a1J0J8zG7_2(.din(n5455), .dout(n23517));
    jdff dff_B_sLsiD19P3_2(.din(n23517), .dout(n23520));
    jdff dff_B_kZurIMWo1_2(.din(n23520), .dout(n23523));
    jdff dff_B_v1clK4ii3_2(.din(n23523), .dout(n23526));
    jdff dff_B_kbrYLWt37_2(.din(n23526), .dout(n23529));
    jdff dff_B_C1Pb4Yuh2_2(.din(n23529), .dout(n23532));
    jdff dff_B_Dut4g0gZ1_2(.din(n23532), .dout(n23535));
    jdff dff_B_MpKWRWAR2_2(.din(n23535), .dout(n23538));
    jdff dff_B_Fql4Qd7Y3_2(.din(n23538), .dout(n23541));
    jdff dff_B_HHxpagHl6_2(.din(n23541), .dout(n23544));
    jdff dff_B_PZ1KQNwm2_2(.din(n23544), .dout(n23547));
    jdff dff_B_nKl0y47p4_2(.din(n23547), .dout(n23550));
    jdff dff_B_OYBpVMMG4_2(.din(n23550), .dout(n23553));
    jdff dff_B_DhW66jAU8_2(.din(n23553), .dout(n23556));
    jdff dff_B_PKuxjvw20_2(.din(n23556), .dout(n23559));
    jdff dff_B_XO8h7PGg5_2(.din(n23559), .dout(n23562));
    jdff dff_B_6upL2GWj7_2(.din(n23562), .dout(n23565));
    jdff dff_B_GFhoQmhn0_2(.din(n23565), .dout(n23568));
    jdff dff_B_SY94yo6c3_2(.din(n23568), .dout(n23571));
    jdff dff_B_usDLdEv52_2(.din(n23571), .dout(n23574));
    jdff dff_B_sQZJRW9M8_2(.din(n23574), .dout(n23577));
    jdff dff_B_RS1zbws18_2(.din(n23577), .dout(n23580));
    jdff dff_B_oizmTqgH0_2(.din(n23580), .dout(n23583));
    jdff dff_B_7PiZW7l29_2(.din(n23583), .dout(n23586));
    jdff dff_B_A6TJtnUN1_2(.din(n23586), .dout(n23589));
    jdff dff_B_ohZEdczW6_2(.din(n23589), .dout(n23592));
    jdff dff_B_qy9MKSzC9_2(.din(n23592), .dout(n23595));
    jdff dff_B_iIQ3jMah6_2(.din(n23595), .dout(n23598));
    jdff dff_B_R38DuS625_2(.din(n23598), .dout(n23601));
    jdff dff_B_vIsaCBPL2_2(.din(n23601), .dout(n23604));
    jdff dff_B_cUbWS54X7_2(.din(n23604), .dout(n23607));
    jdff dff_B_eOyqHQmx1_2(.din(n23607), .dout(n23610));
    jdff dff_B_i0NGRoIy4_2(.din(n23610), .dout(n23613));
    jdff dff_B_QUAW3t0y8_2(.din(n23613), .dout(n23616));
    jdff dff_B_fLeIxoKr1_2(.din(n23616), .dout(n23619));
    jdff dff_B_hKsMYOUV6_2(.din(n23619), .dout(n23622));
    jdff dff_B_9uGbm21M2_2(.din(n23622), .dout(n23625));
    jdff dff_B_azQbmOOL5_2(.din(n23625), .dout(n23628));
    jdff dff_B_BHERS2qa9_2(.din(n5606), .dout(n23631));
    jdff dff_B_zf6t6t9G7_1(.din(n5459), .dout(n23634));
    jdff dff_B_dHAvEPUM8_2(.din(n5183), .dout(n23637));
    jdff dff_B_9vA585IV4_2(.din(n23637), .dout(n23640));
    jdff dff_B_5Ot79jrZ1_2(.din(n23640), .dout(n23643));
    jdff dff_B_bQt6pq1O5_2(.din(n23643), .dout(n23646));
    jdff dff_B_aCRvs3vO8_2(.din(n23646), .dout(n23649));
    jdff dff_B_OuMRJDx00_2(.din(n23649), .dout(n23652));
    jdff dff_B_7rnNunb37_2(.din(n23652), .dout(n23655));
    jdff dff_B_UNyA0LNQ6_2(.din(n23655), .dout(n23658));
    jdff dff_B_NkuPCib06_2(.din(n23658), .dout(n23661));
    jdff dff_B_HrWAqTVg2_2(.din(n23661), .dout(n23664));
    jdff dff_B_jr0H6M1h2_2(.din(n23664), .dout(n23667));
    jdff dff_B_SWrWulLa4_2(.din(n23667), .dout(n23670));
    jdff dff_B_Jct4dJkK5_2(.din(n23670), .dout(n23673));
    jdff dff_B_gvxPh2zu3_2(.din(n23673), .dout(n23676));
    jdff dff_B_irv6qS638_2(.din(n23676), .dout(n23679));
    jdff dff_B_77RqiY8q1_2(.din(n23679), .dout(n23682));
    jdff dff_B_4vLrbhgG4_2(.din(n23682), .dout(n23685));
    jdff dff_B_oshIgT4C9_2(.din(n23685), .dout(n23688));
    jdff dff_B_m3SBlrPt7_2(.din(n23688), .dout(n23691));
    jdff dff_B_tfumFg1C3_2(.din(n23691), .dout(n23694));
    jdff dff_B_wLCrObGZ6_2(.din(n23694), .dout(n23697));
    jdff dff_B_VVLKQ5Q39_2(.din(n23697), .dout(n23700));
    jdff dff_B_ezfXU9GF3_2(.din(n23700), .dout(n23703));
    jdff dff_B_cdb9Mvoj9_2(.din(n23703), .dout(n23706));
    jdff dff_B_lLLZcuUT7_2(.din(n23706), .dout(n23709));
    jdff dff_B_6O5EvuP08_2(.din(n23709), .dout(n23712));
    jdff dff_B_Ooj3M8kE1_2(.din(n23712), .dout(n23715));
    jdff dff_B_MKSnQWk41_2(.din(n23715), .dout(n23718));
    jdff dff_B_oLOudchR1_2(.din(n23718), .dout(n23721));
    jdff dff_B_zLTCYzRl5_2(.din(n23721), .dout(n23724));
    jdff dff_B_16exLBNQ7_2(.din(n23724), .dout(n23727));
    jdff dff_B_EdcHSJMl5_2(.din(n23727), .dout(n23730));
    jdff dff_B_shG9GEvp3_2(.din(n23730), .dout(n23733));
    jdff dff_B_27VPICdG5_2(.din(n23733), .dout(n23736));
    jdff dff_B_S6AkPJPj3_2(.din(n23736), .dout(n23739));
    jdff dff_B_YJTAuJ945_2(.din(n5334), .dout(n23742));
    jdff dff_B_vokYGC0b9_1(.din(n5187), .dout(n23745));
    jdff dff_B_Rs2hwzpB6_2(.din(n4884), .dout(n23748));
    jdff dff_B_aasmsvVd2_2(.din(n23748), .dout(n23751));
    jdff dff_B_4LFEAv2j1_2(.din(n23751), .dout(n23754));
    jdff dff_B_eaDDy6O16_2(.din(n23754), .dout(n23757));
    jdff dff_B_OcaGUfCW3_2(.din(n23757), .dout(n23760));
    jdff dff_B_PNv8s8b13_2(.din(n23760), .dout(n23763));
    jdff dff_B_vBZLomtJ0_2(.din(n23763), .dout(n23766));
    jdff dff_B_pFNvnAe62_2(.din(n23766), .dout(n23769));
    jdff dff_B_JH47gPyU9_2(.din(n23769), .dout(n23772));
    jdff dff_B_rV3xResR9_2(.din(n23772), .dout(n23775));
    jdff dff_B_63Ip9KMa2_2(.din(n23775), .dout(n23778));
    jdff dff_B_6M2EC8Sh4_2(.din(n23778), .dout(n23781));
    jdff dff_B_bcnpDTA37_2(.din(n23781), .dout(n23784));
    jdff dff_B_CZEdGSg04_2(.din(n23784), .dout(n23787));
    jdff dff_B_mm5R5TOt7_2(.din(n23787), .dout(n23790));
    jdff dff_B_60Pm7ex72_2(.din(n23790), .dout(n23793));
    jdff dff_B_PblsyD8d8_2(.din(n23793), .dout(n23796));
    jdff dff_B_RwT1Wr1B0_2(.din(n23796), .dout(n23799));
    jdff dff_B_vzNWISLk7_2(.din(n23799), .dout(n23802));
    jdff dff_B_3Kovejb60_2(.din(n23802), .dout(n23805));
    jdff dff_B_fYZ8xuDg6_2(.din(n23805), .dout(n23808));
    jdff dff_B_chM9taEi2_2(.din(n23808), .dout(n23811));
    jdff dff_B_74WmtdW34_2(.din(n23811), .dout(n23814));
    jdff dff_B_j07Wur1H8_2(.din(n23814), .dout(n23817));
    jdff dff_B_oqLzKfjo0_2(.din(n23817), .dout(n23820));
    jdff dff_B_AcLahKgS3_2(.din(n23820), .dout(n23823));
    jdff dff_B_t5uMJZv03_2(.din(n23823), .dout(n23826));
    jdff dff_B_3hXUBDKd9_2(.din(n23826), .dout(n23829));
    jdff dff_B_V6ganN2S2_2(.din(n23829), .dout(n23832));
    jdff dff_B_ZnWklMm30_2(.din(n23832), .dout(n23835));
    jdff dff_B_HPrd3aYp5_2(.din(n23835), .dout(n23838));
    jdff dff_B_FQxKZDL89_2(.din(n23838), .dout(n23841));
    jdff dff_B_Iax4cSnN7_2(.din(n5035), .dout(n23844));
    jdff dff_B_UmQpK0rO6_1(.din(n4888), .dout(n23847));
    jdff dff_B_FsbPAJqs4_2(.din(n4558), .dout(n23850));
    jdff dff_B_hr2bwteo6_2(.din(n23850), .dout(n23853));
    jdff dff_B_SPLLnP7V4_2(.din(n23853), .dout(n23856));
    jdff dff_B_ZQK7VYsx0_2(.din(n23856), .dout(n23859));
    jdff dff_B_eP6flCHu8_2(.din(n23859), .dout(n23862));
    jdff dff_B_brZIFypa5_2(.din(n23862), .dout(n23865));
    jdff dff_B_pqV4ZWSR7_2(.din(n23865), .dout(n23868));
    jdff dff_B_UYsBVN7x8_2(.din(n23868), .dout(n23871));
    jdff dff_B_tBOkJJb40_2(.din(n23871), .dout(n23874));
    jdff dff_B_nsVhCZI74_2(.din(n23874), .dout(n23877));
    jdff dff_B_cuijBt0D2_2(.din(n23877), .dout(n23880));
    jdff dff_B_9wj8SFYG0_2(.din(n23880), .dout(n23883));
    jdff dff_B_tsTS65vP0_2(.din(n23883), .dout(n23886));
    jdff dff_B_9Kcyb6XJ9_2(.din(n23886), .dout(n23889));
    jdff dff_B_9PupgfsD7_2(.din(n23889), .dout(n23892));
    jdff dff_B_6XqStstz9_2(.din(n23892), .dout(n23895));
    jdff dff_B_6eOq1zfV8_2(.din(n23895), .dout(n23898));
    jdff dff_B_ILwT88TU8_2(.din(n23898), .dout(n23901));
    jdff dff_B_BUWLskyo8_2(.din(n23901), .dout(n23904));
    jdff dff_B_N4sZZfxb6_2(.din(n23904), .dout(n23907));
    jdff dff_B_eqDd9iGy1_2(.din(n23907), .dout(n23910));
    jdff dff_B_wpPzMh8I8_2(.din(n23910), .dout(n23913));
    jdff dff_B_c7gFdwpw1_2(.din(n23913), .dout(n23916));
    jdff dff_B_cIlPVjOn5_2(.din(n23916), .dout(n23919));
    jdff dff_B_NqV9IsLF5_2(.din(n23919), .dout(n23922));
    jdff dff_B_Rb0pOu6w7_2(.din(n23922), .dout(n23925));
    jdff dff_B_662tQZJI7_2(.din(n23925), .dout(n23928));
    jdff dff_B_kSVCW75S1_2(.din(n23928), .dout(n23931));
    jdff dff_B_BJnENFj11_2(.din(n23931), .dout(n23934));
    jdff dff_B_iPNammup2_2(.din(n4709), .dout(n23937));
    jdff dff_B_kV5BDMjF1_1(.din(n4562), .dout(n23940));
    jdff dff_B_XhDtq3AJ2_2(.din(n4208), .dout(n23943));
    jdff dff_B_OtLSsN8s5_2(.din(n23943), .dout(n23946));
    jdff dff_B_bnGijKmp3_2(.din(n23946), .dout(n23949));
    jdff dff_B_hG63Xueq7_2(.din(n23949), .dout(n23952));
    jdff dff_B_n7O1Vi9l0_2(.din(n23952), .dout(n23955));
    jdff dff_B_EFcVe6XA3_2(.din(n23955), .dout(n23958));
    jdff dff_B_gUOyplqD7_2(.din(n23958), .dout(n23961));
    jdff dff_B_fOUSJ79E6_2(.din(n23961), .dout(n23964));
    jdff dff_B_C8o3RLos2_2(.din(n23964), .dout(n23967));
    jdff dff_B_pFQjw1tg7_2(.din(n23967), .dout(n23970));
    jdff dff_B_FI3zd4kB1_2(.din(n23970), .dout(n23973));
    jdff dff_B_2OInZIqZ2_2(.din(n23973), .dout(n23976));
    jdff dff_B_UZfuMZFs9_2(.din(n23976), .dout(n23979));
    jdff dff_B_7JcPBHQe5_2(.din(n23979), .dout(n23982));
    jdff dff_B_ndH0dVsQ9_2(.din(n23982), .dout(n23985));
    jdff dff_B_pkbBsHLO6_2(.din(n23985), .dout(n23988));
    jdff dff_B_NnntY5257_2(.din(n23988), .dout(n23991));
    jdff dff_B_iOERsrR15_2(.din(n23991), .dout(n23994));
    jdff dff_B_XxpYyPVq8_2(.din(n23994), .dout(n23997));
    jdff dff_B_Q5tekKKe3_2(.din(n23997), .dout(n24000));
    jdff dff_B_vLguwKsV5_2(.din(n24000), .dout(n24003));
    jdff dff_B_0dbO5Wv47_2(.din(n24003), .dout(n24006));
    jdff dff_B_OtmVuPkN3_2(.din(n24006), .dout(n24009));
    jdff dff_B_zByO5G0a4_2(.din(n24009), .dout(n24012));
    jdff dff_B_7Pig3tyK4_2(.din(n24012), .dout(n24015));
    jdff dff_B_JryGpri68_2(.din(n24015), .dout(n24018));
    jdff dff_B_Plxwei5y9_2(.din(n4359), .dout(n24021));
    jdff dff_B_OjcRlY2h2_1(.din(n4212), .dout(n24024));
    jdff dff_B_HPLnmYZ77_2(.din(n3832), .dout(n24027));
    jdff dff_B_LbOgLdUB8_2(.din(n24027), .dout(n24030));
    jdff dff_B_8NvYTmhn2_2(.din(n24030), .dout(n24033));
    jdff dff_B_MEBeBxjM5_2(.din(n24033), .dout(n24036));
    jdff dff_B_IGindAYx2_2(.din(n24036), .dout(n24039));
    jdff dff_B_ZQPs9dvB0_2(.din(n24039), .dout(n24042));
    jdff dff_B_ZCpSSidV1_2(.din(n24042), .dout(n24045));
    jdff dff_B_jXxu9ANi9_2(.din(n24045), .dout(n24048));
    jdff dff_B_tu67hxLv5_2(.din(n24048), .dout(n24051));
    jdff dff_B_0blAYzrs3_2(.din(n24051), .dout(n24054));
    jdff dff_B_TbBUV0R14_2(.din(n24054), .dout(n24057));
    jdff dff_B_JDREr97s5_2(.din(n24057), .dout(n24060));
    jdff dff_B_yb7PB9Q66_2(.din(n24060), .dout(n24063));
    jdff dff_B_nb3SKiOT1_2(.din(n24063), .dout(n24066));
    jdff dff_B_WWQgLknE4_2(.din(n24066), .dout(n24069));
    jdff dff_B_3O4752CT8_2(.din(n24069), .dout(n24072));
    jdff dff_B_vQ44mGwc6_2(.din(n24072), .dout(n24075));
    jdff dff_B_raAU1QSt2_2(.din(n24075), .dout(n24078));
    jdff dff_B_mvcsrnVc6_2(.din(n24078), .dout(n24081));
    jdff dff_B_TNAedXlp4_2(.din(n24081), .dout(n24084));
    jdff dff_B_UNstYPRl4_2(.din(n24084), .dout(n24087));
    jdff dff_B_86jlqXc21_2(.din(n24087), .dout(n24090));
    jdff dff_B_tSTxillR3_2(.din(n24090), .dout(n24093));
    jdff dff_B_hTlA5sbm7_2(.din(n3979), .dout(n24096));
    jdff dff_B_4uKjXcCu3_1(.din(n3836), .dout(n24099));
    jdff dff_B_fQlxMl3S2_2(.din(n3452), .dout(n24102));
    jdff dff_B_vOfmXFxe6_2(.din(n24102), .dout(n24105));
    jdff dff_B_Dnm3OYAp9_2(.din(n24105), .dout(n24108));
    jdff dff_B_6BoHQNdw7_2(.din(n24108), .dout(n24111));
    jdff dff_B_8skwEj4r5_2(.din(n24111), .dout(n24114));
    jdff dff_B_SDPVJy5z0_2(.din(n24114), .dout(n24117));
    jdff dff_B_1eEa4Tww7_2(.din(n24117), .dout(n24120));
    jdff dff_B_5oxYSuVg4_2(.din(n24120), .dout(n24123));
    jdff dff_B_qVWTOqfh8_2(.din(n24123), .dout(n24126));
    jdff dff_B_ebnHM4xV7_2(.din(n24126), .dout(n24129));
    jdff dff_B_NnQfzU9z1_2(.din(n24129), .dout(n24132));
    jdff dff_B_IozRSbbz6_2(.din(n24132), .dout(n24135));
    jdff dff_B_vM7YJ0Xz1_2(.din(n24135), .dout(n24138));
    jdff dff_B_qD9Fs3SU4_2(.din(n24138), .dout(n24141));
    jdff dff_B_xmQi2xox5_2(.din(n24141), .dout(n24144));
    jdff dff_B_jBhYpXq06_2(.din(n24144), .dout(n24147));
    jdff dff_B_CAA55B1Q4_2(.din(n24147), .dout(n24150));
    jdff dff_B_abYapm3v1_2(.din(n24150), .dout(n24153));
    jdff dff_B_x7NgL6XT6_2(.din(n24153), .dout(n24156));
    jdff dff_B_f5N2DkNH4_2(.din(n24156), .dout(n24159));
    jdff dff_B_D286X2Hh9_2(.din(n3596), .dout(n24162));
    jdff dff_B_UxsF3NTc2_1(.din(n3456), .dout(n24165));
    jdff dff_B_hX83ipm33_2(.din(n3061), .dout(n24168));
    jdff dff_B_zHvMk9Xz7_2(.din(n24168), .dout(n24171));
    jdff dff_B_HWcn8jjT1_2(.din(n24171), .dout(n24174));
    jdff dff_B_mGgKSy1w6_2(.din(n24174), .dout(n24177));
    jdff dff_B_LkwT9Bz25_2(.din(n24177), .dout(n24180));
    jdff dff_B_UygJsp3C1_2(.din(n24180), .dout(n24183));
    jdff dff_B_Fj9SQ95y6_2(.din(n24183), .dout(n24186));
    jdff dff_B_OOIce2499_2(.din(n24186), .dout(n24189));
    jdff dff_B_fCJYw80P6_2(.din(n24189), .dout(n24192));
    jdff dff_B_3bHjyah09_2(.din(n24192), .dout(n24195));
    jdff dff_B_Bz4Qlem84_2(.din(n24195), .dout(n24198));
    jdff dff_B_5G53VeFP1_2(.din(n24198), .dout(n24201));
    jdff dff_B_ydf0zOwQ6_2(.din(n24201), .dout(n24204));
    jdff dff_B_Mr9PeNBM7_2(.din(n24204), .dout(n24207));
    jdff dff_B_mijPNv5Q7_2(.din(n24207), .dout(n24210));
    jdff dff_B_EfAza7EV0_2(.din(n24210), .dout(n24213));
    jdff dff_B_QFBFxzKh3_2(.din(n24213), .dout(n24216));
    jdff dff_B_FYrpa1pl8_2(.din(n3191), .dout(n24219));
    jdff dff_B_0SQLVANx9_1(.din(n3065), .dout(n24222));
    jdff dff_B_JMyW1ypF9_2(.din(n2686), .dout(n24225));
    jdff dff_B_ZabHqtev9_2(.din(n24225), .dout(n24228));
    jdff dff_B_IgmttBZF3_2(.din(n24228), .dout(n24231));
    jdff dff_B_kxWji1ZO6_2(.din(n24231), .dout(n24234));
    jdff dff_B_d0AN3yjj9_2(.din(n24234), .dout(n24237));
    jdff dff_B_Yyo1N9A11_2(.din(n24237), .dout(n24240));
    jdff dff_B_vNMxwU1F8_2(.din(n24240), .dout(n24243));
    jdff dff_B_WhY8Jqys4_2(.din(n24243), .dout(n24246));
    jdff dff_B_E0b8Qx8l9_2(.din(n24246), .dout(n24249));
    jdff dff_B_FGUSWCTU2_2(.din(n24249), .dout(n24252));
    jdff dff_B_wZjoefnz4_2(.din(n24252), .dout(n24255));
    jdff dff_B_DLMpgKeL7_2(.din(n24255), .dout(n24258));
    jdff dff_B_KgWTyaJP3_2(.din(n24258), .dout(n24261));
    jdff dff_B_VRnjLZMF3_2(.din(n24261), .dout(n24264));
    jdff dff_B_1GKvZS0y0_2(.din(n2796), .dout(n24267));
    jdff dff_B_L9dAiNeY6_1(.din(n2690), .dout(n24270));
    jdff dff_B_2hQyrjfp5_2(.din(n2335), .dout(n24273));
    jdff dff_B_BOZk9Qht4_2(.din(n24273), .dout(n24276));
    jdff dff_B_r1xfYZN53_2(.din(n24276), .dout(n24279));
    jdff dff_B_EPQRGGMb7_2(.din(n24279), .dout(n24282));
    jdff dff_B_iIKiHArP0_2(.din(n24282), .dout(n24285));
    jdff dff_B_Eu9Ud1cb9_2(.din(n24285), .dout(n24288));
    jdff dff_B_kH1awpSJ2_2(.din(n24288), .dout(n24291));
    jdff dff_B_epbDVz3U0_2(.din(n24291), .dout(n24294));
    jdff dff_B_KZTDu68j0_2(.din(n24294), .dout(n24297));
    jdff dff_B_v20WeeIt3_2(.din(n24297), .dout(n24300));
    jdff dff_B_RmOrkIc96_2(.din(n24300), .dout(n24303));
    jdff dff_B_6vOacekQ0_2(.din(n2418), .dout(n24306));
    jdff dff_B_fhsB5pI32_1(.din(n2339), .dout(n24309));
    jdff dff_B_j6r1Pr0z6_2(.din(n2011), .dout(n24312));
    jdff dff_B_RyfUBfVm0_2(.din(n24312), .dout(n24315));
    jdff dff_B_ZW9y5cSy0_2(.din(n24315), .dout(n24318));
    jdff dff_B_zvjJeL4G4_2(.din(n24318), .dout(n24321));
    jdff dff_B_oPHvr82C4_2(.din(n24321), .dout(n24324));
    jdff dff_B_Gng1ttnp6_2(.din(n24324), .dout(n24327));
    jdff dff_B_IDqVQHuX0_2(.din(n24327), .dout(n24330));
    jdff dff_B_SF8nTlbT9_2(.din(n24330), .dout(n24333));
    jdff dff_B_1peuGQj02_2(.din(n2067), .dout(n24336));
    jdff dff_B_ioxh8fVC2_2(.din(n24336), .dout(n24339));
    jdff dff_B_7qNLUpmv4_2(.din(n24339), .dout(n24342));
    jdff dff_B_4LAuJUSU0_1(.din(n2015), .dout(n24345));
    jdff dff_B_Zdg8hQQA3_1(.din(n24345), .dout(n24348));
    jdff dff_B_ESJgNDMp1_2(.din(n1720), .dout(n24351));
    jdff dff_B_L6eWh6e09_2(.din(n24351), .dout(n24354));
    jdff dff_B_7ZZLxOsm6_2(.din(n24354), .dout(n24357));
    jdff dff_B_pZTOoJE89_0(.din(n1739), .dout(n24360));
    jdff dff_A_5Se624DU4_0(.din(n24365), .dout(n24362));
    jdff dff_A_tI7GeNyK3_0(.din(n1439), .dout(n24365));
    jdff dff_A_ZWzEZO8B7_1(.din(n24371), .dout(n24368));
    jdff dff_A_4MM8phz66_1(.din(n1439), .dout(n24371));
    jdff dff_B_GwYof2122_1(.din(n6424), .dout(n24375));
    jdff dff_A_SwQ6ri8m3_1(.din(n6301), .dout(n24377));
    jdff dff_B_2BO5H3Fh3_1(.din(n6293), .dout(n24381));
    jdff dff_B_RcXJoA6M0_2(.din(n6131), .dout(n24384));
    jdff dff_B_Y2oKoKr14_2(.din(n24384), .dout(n24387));
    jdff dff_B_AqPVFHW88_2(.din(n24387), .dout(n24390));
    jdff dff_B_LXSgQJGn9_2(.din(n24390), .dout(n24393));
    jdff dff_B_tnyuM3JP5_2(.din(n24393), .dout(n24396));
    jdff dff_B_EsATly1H6_2(.din(n24396), .dout(n24399));
    jdff dff_B_drNmJrFC1_2(.din(n24399), .dout(n24402));
    jdff dff_B_IZfbzlGw3_2(.din(n24402), .dout(n24405));
    jdff dff_B_kwFoYC738_2(.din(n24405), .dout(n24408));
    jdff dff_B_48rGiQOT0_2(.din(n24408), .dout(n24411));
    jdff dff_B_SJPeioDR3_2(.din(n24411), .dout(n24414));
    jdff dff_B_lFPka0Mg0_2(.din(n24414), .dout(n24417));
    jdff dff_B_q4jIGpo08_2(.din(n24417), .dout(n24420));
    jdff dff_B_6I0723fN9_2(.din(n24420), .dout(n24423));
    jdff dff_B_4Rmj2au51_2(.din(n24423), .dout(n24426));
    jdff dff_B_QsbgupvY5_2(.din(n24426), .dout(n24429));
    jdff dff_B_gR31hLuU8_2(.din(n24429), .dout(n24432));
    jdff dff_B_ayIruosr3_2(.din(n24432), .dout(n24435));
    jdff dff_B_FR4NXnEc2_2(.din(n24435), .dout(n24438));
    jdff dff_B_U8P0ZI8H6_2(.din(n24438), .dout(n24441));
    jdff dff_B_3uuSu37e9_2(.din(n24441), .dout(n24444));
    jdff dff_B_pJgnBA9L0_2(.din(n24444), .dout(n24447));
    jdff dff_B_oMVFEaJZ8_2(.din(n24447), .dout(n24450));
    jdff dff_B_SNcH6jEJ1_2(.din(n24450), .dout(n24453));
    jdff dff_B_Y9glgvmM9_2(.din(n24453), .dout(n24456));
    jdff dff_B_FSEjjpyd0_2(.din(n24456), .dout(n24459));
    jdff dff_B_1crG85sG9_2(.din(n24459), .dout(n24462));
    jdff dff_B_vTiA19Pk2_2(.din(n24462), .dout(n24465));
    jdff dff_B_Lyc5LJAo0_2(.din(n24465), .dout(n24468));
    jdff dff_B_bGXVEpuy0_2(.din(n24468), .dout(n24471));
    jdff dff_B_mSs1jPUu0_2(.din(n24471), .dout(n24474));
    jdff dff_B_Pku4wRHZ5_2(.din(n24474), .dout(n24477));
    jdff dff_B_B7nL4GdN8_2(.din(n24477), .dout(n24480));
    jdff dff_B_KGXfH1jC9_2(.din(n24480), .dout(n24483));
    jdff dff_B_J2KmmILp8_2(.din(n24483), .dout(n24486));
    jdff dff_B_OJ7Z7NdO4_2(.din(n24486), .dout(n24489));
    jdff dff_B_4gXtPzDy4_2(.din(n24489), .dout(n24492));
    jdff dff_B_JGdoBNXQ8_2(.din(n24492), .dout(n24495));
    jdff dff_B_VD9mQd8f7_2(.din(n24495), .dout(n24498));
    jdff dff_B_Ch4NS9AK4_2(.din(n24498), .dout(n24501));
    jdff dff_B_J1tycnE23_2(.din(n24501), .dout(n24504));
    jdff dff_B_aVyGAD361_2(.din(n24504), .dout(n24507));
    jdff dff_B_7v498nzy0_2(.din(n24507), .dout(n24510));
    jdff dff_B_JaHyIaEv7_2(.din(n24510), .dout(n24513));
    jdff dff_B_0Z2jdXNz8_2(.din(n24513), .dout(n24516));
    jdff dff_B_nBxfy3Zo3_2(.din(n24516), .dout(n24519));
    jdff dff_B_toABSUla3_2(.din(n6143), .dout(n24522));
    jdff dff_B_fL374ioq5_1(.din(n6135), .dout(n24525));
    jdff dff_B_srz84Pgv4_2(.din(n5937), .dout(n24528));
    jdff dff_B_sUGcgf2X2_2(.din(n24528), .dout(n24531));
    jdff dff_B_RUO0MwKQ6_2(.din(n24531), .dout(n24534));
    jdff dff_B_5CxXe5pG9_2(.din(n24534), .dout(n24537));
    jdff dff_B_50FqWL0Y6_2(.din(n24537), .dout(n24540));
    jdff dff_B_ArT0Qvck4_2(.din(n24540), .dout(n24543));
    jdff dff_B_QYaoqqG31_2(.din(n24543), .dout(n24546));
    jdff dff_B_bRblvbew7_2(.din(n24546), .dout(n24549));
    jdff dff_B_WLVMwxOw3_2(.din(n24549), .dout(n24552));
    jdff dff_B_vqFZ7Nlo6_2(.din(n24552), .dout(n24555));
    jdff dff_B_azEYAeet3_2(.din(n24555), .dout(n24558));
    jdff dff_B_6GDNLp3L0_2(.din(n24558), .dout(n24561));
    jdff dff_B_GR1mAU6h5_2(.din(n24561), .dout(n24564));
    jdff dff_B_iG84c0cQ4_2(.din(n24564), .dout(n24567));
    jdff dff_B_c0IoGkQP4_2(.din(n24567), .dout(n24570));
    jdff dff_B_gmBvsdYM9_2(.din(n24570), .dout(n24573));
    jdff dff_B_NrddrdD48_2(.din(n24573), .dout(n24576));
    jdff dff_B_qbGeRZxD1_2(.din(n24576), .dout(n24579));
    jdff dff_B_2ser7ZdF1_2(.din(n24579), .dout(n24582));
    jdff dff_B_47goirtf3_2(.din(n24582), .dout(n24585));
    jdff dff_B_D7XGDyVJ9_2(.din(n24585), .dout(n24588));
    jdff dff_B_sHbW1fKC7_2(.din(n24588), .dout(n24591));
    jdff dff_B_0Vhg79P96_2(.din(n24591), .dout(n24594));
    jdff dff_B_hvuTvXpA6_2(.din(n24594), .dout(n24597));
    jdff dff_B_5xX9sl2J5_2(.din(n24597), .dout(n24600));
    jdff dff_B_NQN0w1Pi1_2(.din(n24600), .dout(n24603));
    jdff dff_B_Ch0jz0Lk7_2(.din(n24603), .dout(n24606));
    jdff dff_B_6RVLTVQF5_2(.din(n24606), .dout(n24609));
    jdff dff_B_VKIDSFkq0_2(.din(n24609), .dout(n24612));
    jdff dff_B_6WOtqA6l9_2(.din(n24612), .dout(n24615));
    jdff dff_B_EUwzOq7b3_2(.din(n24615), .dout(n24618));
    jdff dff_B_YLDpHNXV0_2(.din(n24618), .dout(n24621));
    jdff dff_B_36NqWeYd2_2(.din(n24621), .dout(n24624));
    jdff dff_B_2brQbtMX9_2(.din(n24624), .dout(n24627));
    jdff dff_B_DqxQL4XO5_2(.din(n24627), .dout(n24630));
    jdff dff_B_NniZN1Ep7_2(.din(n24630), .dout(n24633));
    jdff dff_B_mgg01KfN9_2(.din(n24633), .dout(n24636));
    jdff dff_B_O9TiFwU31_2(.din(n24636), .dout(n24639));
    jdff dff_B_KzSalANb9_2(.din(n24639), .dout(n24642));
    jdff dff_B_Z8fkM5Ii2_2(.din(n24642), .dout(n24645));
    jdff dff_B_IPbenLDB9_2(.din(n24645), .dout(n24648));
    jdff dff_B_7sCSoUGO2_2(.din(n24648), .dout(n24651));
    jdff dff_B_JeVevLGF2_2(.din(n5949), .dout(n24654));
    jdff dff_B_72FCd2WI3_1(.din(n5941), .dout(n24657));
    jdff dff_B_0Vkd3RTi3_2(.din(n5719), .dout(n24660));
    jdff dff_B_viszoCbb1_2(.din(n24660), .dout(n24663));
    jdff dff_B_HKpayDrq0_2(.din(n24663), .dout(n24666));
    jdff dff_B_E9oVdWO76_2(.din(n24666), .dout(n24669));
    jdff dff_B_jhOmsjKU5_2(.din(n24669), .dout(n24672));
    jdff dff_B_xtnw1jPq3_2(.din(n24672), .dout(n24675));
    jdff dff_B_vMVUCDk53_2(.din(n24675), .dout(n24678));
    jdff dff_B_LLlFAXGO4_2(.din(n24678), .dout(n24681));
    jdff dff_B_WSTci83g3_2(.din(n24681), .dout(n24684));
    jdff dff_B_Sy19B0WV3_2(.din(n24684), .dout(n24687));
    jdff dff_B_hSeXNY4M3_2(.din(n24687), .dout(n24690));
    jdff dff_B_knrWhgjB0_2(.din(n24690), .dout(n24693));
    jdff dff_B_AlE2HCrZ7_2(.din(n24693), .dout(n24696));
    jdff dff_B_pUKBjtUL4_2(.din(n24696), .dout(n24699));
    jdff dff_B_x9Vc4eVj3_2(.din(n24699), .dout(n24702));
    jdff dff_B_YlLyWT2v8_2(.din(n24702), .dout(n24705));
    jdff dff_B_hE1A2bxz0_2(.din(n24705), .dout(n24708));
    jdff dff_B_RViGyZXN7_2(.din(n24708), .dout(n24711));
    jdff dff_B_js2biHo04_2(.din(n24711), .dout(n24714));
    jdff dff_B_WXYXMVMO7_2(.din(n24714), .dout(n24717));
    jdff dff_B_P71syNyq0_2(.din(n24717), .dout(n24720));
    jdff dff_B_3ubAaHD18_2(.din(n24720), .dout(n24723));
    jdff dff_B_ZKTx0qP55_2(.din(n24723), .dout(n24726));
    jdff dff_B_NRRn0mRd2_2(.din(n24726), .dout(n24729));
    jdff dff_B_qGaMJt2o9_2(.din(n24729), .dout(n24732));
    jdff dff_B_UOKfX48y1_2(.din(n24732), .dout(n24735));
    jdff dff_B_UAhTtrPE9_2(.din(n24735), .dout(n24738));
    jdff dff_B_qp6leGgL9_2(.din(n24738), .dout(n24741));
    jdff dff_B_Fun1EjNk6_2(.din(n24741), .dout(n24744));
    jdff dff_B_9F7rfMuK1_2(.din(n24744), .dout(n24747));
    jdff dff_B_N588Bo4B8_2(.din(n24747), .dout(n24750));
    jdff dff_B_jIJU7zvh7_2(.din(n24750), .dout(n24753));
    jdff dff_B_ywrMII1O9_2(.din(n24753), .dout(n24756));
    jdff dff_B_HHFWSoPB6_2(.din(n24756), .dout(n24759));
    jdff dff_B_FCpTu1Oa8_2(.din(n24759), .dout(n24762));
    jdff dff_B_Xjo0NHRN6_2(.din(n24762), .dout(n24765));
    jdff dff_B_6gaVyu1c2_2(.din(n24765), .dout(n24768));
    jdff dff_B_T9xSZq4u2_2(.din(n24768), .dout(n24771));
    jdff dff_B_rtoEWXzK4_1(.din(n5723), .dout(n24774));
    jdff dff_B_gnbereKi1_2(.din(n5474), .dout(n24777));
    jdff dff_B_4sCXKAMt1_2(.din(n24777), .dout(n24780));
    jdff dff_B_6isl9lQp4_2(.din(n24780), .dout(n24783));
    jdff dff_B_Hdl40UF99_2(.din(n24783), .dout(n24786));
    jdff dff_B_k3FqWsEE3_2(.din(n24786), .dout(n24789));
    jdff dff_B_iWKtQyWh8_2(.din(n24789), .dout(n24792));
    jdff dff_B_nvr54PpG3_2(.din(n24792), .dout(n24795));
    jdff dff_B_AK8tEOvm0_2(.din(n24795), .dout(n24798));
    jdff dff_B_1R9eaqrL3_2(.din(n24798), .dout(n24801));
    jdff dff_B_AtGAz6sJ3_2(.din(n24801), .dout(n24804));
    jdff dff_B_bxWflXCE9_2(.din(n24804), .dout(n24807));
    jdff dff_B_SIXSQ67O1_2(.din(n24807), .dout(n24810));
    jdff dff_B_7fkhM7wJ7_2(.din(n24810), .dout(n24813));
    jdff dff_B_zYeiN5JJ3_2(.din(n24813), .dout(n24816));
    jdff dff_B_JMkfEVJD1_2(.din(n24816), .dout(n24819));
    jdff dff_B_Tzx18ChG4_2(.din(n24819), .dout(n24822));
    jdff dff_B_yVYF2ret0_2(.din(n24822), .dout(n24825));
    jdff dff_B_VbsMSVfW1_2(.din(n24825), .dout(n24828));
    jdff dff_B_GRIBojrQ9_2(.din(n24828), .dout(n24831));
    jdff dff_B_ufNGh5Nz9_2(.din(n24831), .dout(n24834));
    jdff dff_B_DDVDSGGr2_2(.din(n24834), .dout(n24837));
    jdff dff_B_mNTMWGwj0_2(.din(n24837), .dout(n24840));
    jdff dff_B_VTye8jUV5_2(.din(n24840), .dout(n24843));
    jdff dff_B_UOQW4Sx61_2(.din(n24843), .dout(n24846));
    jdff dff_B_AXAewekX7_2(.din(n24846), .dout(n24849));
    jdff dff_B_I64BCFFe1_2(.din(n24849), .dout(n24852));
    jdff dff_B_GV3oyR2n5_2(.din(n24852), .dout(n24855));
    jdff dff_B_mjDJMCsb6_2(.din(n24855), .dout(n24858));
    jdff dff_B_8bAUqhY71_2(.din(n24858), .dout(n24861));
    jdff dff_B_WnYZ6jln3_2(.din(n24861), .dout(n24864));
    jdff dff_B_5mHy322U6_2(.din(n24864), .dout(n24867));
    jdff dff_B_w2IKrN7g5_2(.din(n24867), .dout(n24870));
    jdff dff_B_Qx7mxZdT6_2(.din(n24870), .dout(n24873));
    jdff dff_B_V8sIV8sd4_2(.din(n24873), .dout(n24876));
    jdff dff_B_YklFauZj3_2(.din(n24876), .dout(n24879));
    jdff dff_B_p7AWjSaB0_2(.din(n5598), .dout(n24882));
    jdff dff_B_ISJUd31I5_1(.din(n5478), .dout(n24885));
    jdff dff_B_ojx5wQ788_2(.din(n5202), .dout(n24888));
    jdff dff_B_QrGb6vKY1_2(.din(n24888), .dout(n24891));
    jdff dff_B_XmWNjiDD2_2(.din(n24891), .dout(n24894));
    jdff dff_B_U0fFuZLV2_2(.din(n24894), .dout(n24897));
    jdff dff_B_OcXYIF8E9_2(.din(n24897), .dout(n24900));
    jdff dff_B_gsfkJpD56_2(.din(n24900), .dout(n24903));
    jdff dff_B_lX7IsoW62_2(.din(n24903), .dout(n24906));
    jdff dff_B_R6nnz4UU4_2(.din(n24906), .dout(n24909));
    jdff dff_B_iseOWATe5_2(.din(n24909), .dout(n24912));
    jdff dff_B_ekQc6uMI0_2(.din(n24912), .dout(n24915));
    jdff dff_B_Tg2ton5F5_2(.din(n24915), .dout(n24918));
    jdff dff_B_NC6bMZWi2_2(.din(n24918), .dout(n24921));
    jdff dff_B_OV4Ev9ke2_2(.din(n24921), .dout(n24924));
    jdff dff_B_is4k58l98_2(.din(n24924), .dout(n24927));
    jdff dff_B_lyz9BWDG1_2(.din(n24927), .dout(n24930));
    jdff dff_B_guYPLWXn1_2(.din(n24930), .dout(n24933));
    jdff dff_B_mCemIItI9_2(.din(n24933), .dout(n24936));
    jdff dff_B_TqwFgypW8_2(.din(n24936), .dout(n24939));
    jdff dff_B_xYAQw4AV9_2(.din(n24939), .dout(n24942));
    jdff dff_B_EdqLmb3R3_2(.din(n24942), .dout(n24945));
    jdff dff_B_wCYtV0fA5_2(.din(n24945), .dout(n24948));
    jdff dff_B_C2u7cuHN4_2(.din(n24948), .dout(n24951));
    jdff dff_B_57zDsbaF2_2(.din(n24951), .dout(n24954));
    jdff dff_B_jHyEaw602_2(.din(n24954), .dout(n24957));
    jdff dff_B_EGWOWf9O9_2(.din(n24957), .dout(n24960));
    jdff dff_B_3Q829Jkz3_2(.din(n24960), .dout(n24963));
    jdff dff_B_sJTrjs2W8_2(.din(n24963), .dout(n24966));
    jdff dff_B_tCRWd8Nn7_2(.din(n24966), .dout(n24969));
    jdff dff_B_lgAIjsaz4_2(.din(n24969), .dout(n24972));
    jdff dff_B_gFPDvHSl5_2(.din(n24972), .dout(n24975));
    jdff dff_B_XWMtnGVA1_2(.din(n24975), .dout(n24978));
    jdff dff_B_b6jgOv2c9_2(.din(n24978), .dout(n24981));
    jdff dff_B_OMXvXjla2_2(.din(n5326), .dout(n24984));
    jdff dff_B_Np1v8xsj0_1(.din(n5206), .dout(n24987));
    jdff dff_B_r9gpkzOX2_2(.din(n4903), .dout(n24990));
    jdff dff_B_Q5FUyK8T8_2(.din(n24990), .dout(n24993));
    jdff dff_B_WR9kmS2X1_2(.din(n24993), .dout(n24996));
    jdff dff_B_1DoWVFXC1_2(.din(n24996), .dout(n24999));
    jdff dff_B_ZAbB7ElF1_2(.din(n24999), .dout(n25002));
    jdff dff_B_DPWgG65B2_2(.din(n25002), .dout(n25005));
    jdff dff_B_d4tDt8xY2_2(.din(n25005), .dout(n25008));
    jdff dff_B_SE9M4N407_2(.din(n25008), .dout(n25011));
    jdff dff_B_4KpCWajW6_2(.din(n25011), .dout(n25014));
    jdff dff_B_7rAnPWkD7_2(.din(n25014), .dout(n25017));
    jdff dff_B_OAgzgMeN7_2(.din(n25017), .dout(n25020));
    jdff dff_B_f3bO6ym16_2(.din(n25020), .dout(n25023));
    jdff dff_B_HesHG1wa0_2(.din(n25023), .dout(n25026));
    jdff dff_B_n536rLtD1_2(.din(n25026), .dout(n25029));
    jdff dff_B_6lxU23xG7_2(.din(n25029), .dout(n25032));
    jdff dff_B_oK34vapg7_2(.din(n25032), .dout(n25035));
    jdff dff_B_RIE4rCTD5_2(.din(n25035), .dout(n25038));
    jdff dff_B_tP5Jx9bR0_2(.din(n25038), .dout(n25041));
    jdff dff_B_jY14pEFG1_2(.din(n25041), .dout(n25044));
    jdff dff_B_MnnwXFB70_2(.din(n25044), .dout(n25047));
    jdff dff_B_3EnhQxlt8_2(.din(n25047), .dout(n25050));
    jdff dff_B_exRvzMEK2_2(.din(n25050), .dout(n25053));
    jdff dff_B_yAKnvj3u6_2(.din(n25053), .dout(n25056));
    jdff dff_B_j4vFqJ064_2(.din(n25056), .dout(n25059));
    jdff dff_B_yJX6VZx83_2(.din(n25059), .dout(n25062));
    jdff dff_B_GWUwXBzq6_2(.din(n25062), .dout(n25065));
    jdff dff_B_YFRCnf3a8_2(.din(n25065), .dout(n25068));
    jdff dff_B_8IqsvRsL8_2(.din(n25068), .dout(n25071));
    jdff dff_B_FIqkKil95_2(.din(n25071), .dout(n25074));
    jdff dff_B_QCqWFUuj5_2(.din(n5027), .dout(n25077));
    jdff dff_B_sVmjXq6O1_1(.din(n4907), .dout(n25080));
    jdff dff_B_EEabGscb2_2(.din(n4577), .dout(n25083));
    jdff dff_B_C5w2kazg8_2(.din(n25083), .dout(n25086));
    jdff dff_B_r9Sv5kHl7_2(.din(n25086), .dout(n25089));
    jdff dff_B_uGOE5r0T1_2(.din(n25089), .dout(n25092));
    jdff dff_B_9TwJOURK2_2(.din(n25092), .dout(n25095));
    jdff dff_B_TfOF2y5w2_2(.din(n25095), .dout(n25098));
    jdff dff_B_6IR98p932_2(.din(n25098), .dout(n25101));
    jdff dff_B_btSoseQP4_2(.din(n25101), .dout(n25104));
    jdff dff_B_fS0yraMI8_2(.din(n25104), .dout(n25107));
    jdff dff_B_scyRMOS63_2(.din(n25107), .dout(n25110));
    jdff dff_B_pVniVI5P7_2(.din(n25110), .dout(n25113));
    jdff dff_B_9uNclzfI9_2(.din(n25113), .dout(n25116));
    jdff dff_B_c3VBUoBz3_2(.din(n25116), .dout(n25119));
    jdff dff_B_4ifoD7h11_2(.din(n25119), .dout(n25122));
    jdff dff_B_hlolFbYN3_2(.din(n25122), .dout(n25125));
    jdff dff_B_GcVyUEG90_2(.din(n25125), .dout(n25128));
    jdff dff_B_IVrARRAJ7_2(.din(n25128), .dout(n25131));
    jdff dff_B_7JJpx3z64_2(.din(n25131), .dout(n25134));
    jdff dff_B_Jewm9tFG1_2(.din(n25134), .dout(n25137));
    jdff dff_B_p9A0L6m08_2(.din(n25137), .dout(n25140));
    jdff dff_B_lHK1nEr31_2(.din(n25140), .dout(n25143));
    jdff dff_B_xgDKfvmL6_2(.din(n25143), .dout(n25146));
    jdff dff_B_9SBAGRw60_2(.din(n25146), .dout(n25149));
    jdff dff_B_77LkU9Lp6_2(.din(n25149), .dout(n25152));
    jdff dff_B_oo3hJmBa6_2(.din(n25152), .dout(n25155));
    jdff dff_B_lI9bCXDS3_2(.din(n25155), .dout(n25158));
    jdff dff_B_vcCq38sD8_2(.din(n4701), .dout(n25161));
    jdff dff_B_D0MLO62s7_1(.din(n4581), .dout(n25164));
    jdff dff_B_lDD5EwiP7_2(.din(n4227), .dout(n25167));
    jdff dff_B_Hdwz1ovf6_2(.din(n25167), .dout(n25170));
    jdff dff_B_jqabLlTY0_2(.din(n25170), .dout(n25173));
    jdff dff_B_uKePzSI57_2(.din(n25173), .dout(n25176));
    jdff dff_B_gaOYESsH8_2(.din(n25176), .dout(n25179));
    jdff dff_B_CniT0wFX8_2(.din(n25179), .dout(n25182));
    jdff dff_B_dHg9dOE06_2(.din(n25182), .dout(n25185));
    jdff dff_B_NIVvBHeG0_2(.din(n25185), .dout(n25188));
    jdff dff_B_VzNCio8K6_2(.din(n25188), .dout(n25191));
    jdff dff_B_8w6j5v7y6_2(.din(n25191), .dout(n25194));
    jdff dff_B_pcyUuP953_2(.din(n25194), .dout(n25197));
    jdff dff_B_0Hiugs2T1_2(.din(n25197), .dout(n25200));
    jdff dff_B_BAdALqCA6_2(.din(n25200), .dout(n25203));
    jdff dff_B_mSwIxkXj7_2(.din(n25203), .dout(n25206));
    jdff dff_B_T0QRnaFX5_2(.din(n25206), .dout(n25209));
    jdff dff_B_GNuTaNYm0_2(.din(n25209), .dout(n25212));
    jdff dff_B_Dy29BoGg8_2(.din(n25212), .dout(n25215));
    jdff dff_B_tSwhzLp33_2(.din(n25215), .dout(n25218));
    jdff dff_B_gGSt85UG0_2(.din(n25218), .dout(n25221));
    jdff dff_B_YYxGgZYu9_2(.din(n25221), .dout(n25224));
    jdff dff_B_d5I3Ey5t8_2(.din(n25224), .dout(n25227));
    jdff dff_B_QuqzS3fK1_2(.din(n25227), .dout(n25230));
    jdff dff_B_mNza9tcW4_2(.din(n25230), .dout(n25233));
    jdff dff_B_WUYVu1hl2_2(.din(n4351), .dout(n25236));
    jdff dff_B_QMF8uRl06_1(.din(n4231), .dout(n25239));
    jdff dff_B_GWeOCnPO4_2(.din(n3851), .dout(n25242));
    jdff dff_B_dp9fFCs86_2(.din(n25242), .dout(n25245));
    jdff dff_B_VCj82tDn3_2(.din(n25245), .dout(n25248));
    jdff dff_B_vR181oxi7_2(.din(n25248), .dout(n25251));
    jdff dff_B_IxfaIcaT8_2(.din(n25251), .dout(n25254));
    jdff dff_B_IztkZPXG7_2(.din(n25254), .dout(n25257));
    jdff dff_B_hrt4Mc5x8_2(.din(n25257), .dout(n25260));
    jdff dff_B_8G0zxng01_2(.din(n25260), .dout(n25263));
    jdff dff_B_iSS9SgOM1_2(.din(n25263), .dout(n25266));
    jdff dff_B_61yb0ejX0_2(.din(n25266), .dout(n25269));
    jdff dff_B_DyhUzHgK1_2(.din(n25269), .dout(n25272));
    jdff dff_B_Q1Z70QoM6_2(.din(n25272), .dout(n25275));
    jdff dff_B_rKgbTX9Z3_2(.din(n25275), .dout(n25278));
    jdff dff_B_ZyRBvNaZ5_2(.din(n25278), .dout(n25281));
    jdff dff_B_JiEXtOrC9_2(.din(n25281), .dout(n25284));
    jdff dff_B_Ac5JdQf82_2(.din(n25284), .dout(n25287));
    jdff dff_B_QPIfgRm07_2(.din(n25287), .dout(n25290));
    jdff dff_B_dvVVJkmv8_2(.din(n25290), .dout(n25293));
    jdff dff_B_9c7T0okH9_2(.din(n25293), .dout(n25296));
    jdff dff_B_652yf0Nx1_2(.din(n25296), .dout(n25299));
    jdff dff_B_NeEOwLOI0_2(.din(n3971), .dout(n25302));
    jdff dff_B_Fipv8Gnp4_1(.din(n3855), .dout(n25305));
    jdff dff_B_D7jdRNo73_2(.din(n3471), .dout(n25308));
    jdff dff_B_BtA0HKAD4_2(.din(n25308), .dout(n25311));
    jdff dff_B_AhycjzWL7_2(.din(n25311), .dout(n25314));
    jdff dff_B_3xKiqqXz9_2(.din(n25314), .dout(n25317));
    jdff dff_B_T7FWyf9u6_2(.din(n25317), .dout(n25320));
    jdff dff_B_OU22KPS90_2(.din(n25320), .dout(n25323));
    jdff dff_B_RjM9ejhg4_2(.din(n25323), .dout(n25326));
    jdff dff_B_gab97HyR4_2(.din(n25326), .dout(n25329));
    jdff dff_B_rMKqRuTO1_2(.din(n25329), .dout(n25332));
    jdff dff_B_dSkZkfJE4_2(.din(n25332), .dout(n25335));
    jdff dff_B_sN3aDqCS2_2(.din(n25335), .dout(n25338));
    jdff dff_B_ncNNF4w89_2(.din(n25338), .dout(n25341));
    jdff dff_B_mNnMG2Nw2_2(.din(n25341), .dout(n25344));
    jdff dff_B_Nu24rtER5_2(.din(n25344), .dout(n25347));
    jdff dff_B_EH87Q9Ja2_2(.din(n25347), .dout(n25350));
    jdff dff_B_v7n9ZdN78_2(.din(n25350), .dout(n25353));
    jdff dff_B_vel3G9qh4_2(.din(n25353), .dout(n25356));
    jdff dff_B_BygthE7M4_2(.din(n3588), .dout(n25359));
    jdff dff_B_8eTRNjEg9_1(.din(n3475), .dout(n25362));
    jdff dff_B_dSdzBKzL6_2(.din(n3080), .dout(n25365));
    jdff dff_B_kRD1cGHm0_2(.din(n25365), .dout(n25368));
    jdff dff_B_XSB0ImkT2_2(.din(n25368), .dout(n25371));
    jdff dff_B_XFmF0o247_2(.din(n25371), .dout(n25374));
    jdff dff_B_PD1NDFcd8_2(.din(n25374), .dout(n25377));
    jdff dff_B_NB5zcMHp8_2(.din(n25377), .dout(n25380));
    jdff dff_B_LoTM9iGp8_2(.din(n25380), .dout(n25383));
    jdff dff_B_vh1z7EQf4_2(.din(n25383), .dout(n25386));
    jdff dff_B_zQxCkmZz4_2(.din(n25386), .dout(n25389));
    jdff dff_B_f8lY0Vet6_2(.din(n25389), .dout(n25392));
    jdff dff_B_dx4pguYu7_2(.din(n25392), .dout(n25395));
    jdff dff_B_QmuKa4eK6_2(.din(n25395), .dout(n25398));
    jdff dff_B_7X7O8SjT0_2(.din(n25398), .dout(n25401));
    jdff dff_B_y521lsx49_2(.din(n25401), .dout(n25404));
    jdff dff_B_nNHk4TPi9_2(.din(n3183), .dout(n25407));
    jdff dff_B_ls7eEVDF7_1(.din(n3084), .dout(n25410));
    jdff dff_B_zKkPmLf05_2(.din(n2705), .dout(n25413));
    jdff dff_B_TqMtYgbm1_2(.din(n25413), .dout(n25416));
    jdff dff_B_jE18dZpw0_2(.din(n25416), .dout(n25419));
    jdff dff_B_DJpvfd7x3_2(.din(n25419), .dout(n25422));
    jdff dff_B_RhTWUUQC2_2(.din(n25422), .dout(n25425));
    jdff dff_B_lUQaqNA31_2(.din(n25425), .dout(n25428));
    jdff dff_B_jhO1V4YD3_2(.din(n25428), .dout(n25431));
    jdff dff_B_OmTWrffi8_2(.din(n25431), .dout(n25434));
    jdff dff_B_6XF6CHzP5_2(.din(n25434), .dout(n25437));
    jdff dff_B_AZbtr5c57_2(.din(n25437), .dout(n25440));
    jdff dff_B_L4nzzlCr2_2(.din(n25440), .dout(n25443));
    jdff dff_B_t4bNrN1L3_2(.din(n2788), .dout(n25446));
    jdff dff_B_MeaEWRaU7_1(.din(n2709), .dout(n25449));
    jdff dff_B_BHp6WDKG1_2(.din(n2354), .dout(n25452));
    jdff dff_B_DSmInTRM0_2(.din(n25452), .dout(n25455));
    jdff dff_B_3QYMA24v9_2(.din(n25455), .dout(n25458));
    jdff dff_B_SFGCOXC16_2(.din(n25458), .dout(n25461));
    jdff dff_B_PjFtCOgg4_2(.din(n25461), .dout(n25464));
    jdff dff_B_gWzcO45F1_2(.din(n25464), .dout(n25467));
    jdff dff_B_e3dMIBCj6_2(.din(n25467), .dout(n25470));
    jdff dff_B_KiS2yLUk1_2(.din(n25470), .dout(n25473));
    jdff dff_B_5fbQ0Tdx8_2(.din(n2410), .dout(n25476));
    jdff dff_B_FXkMh77Y8_2(.din(n25476), .dout(n25479));
    jdff dff_B_BJLQn1AZ7_2(.din(n25479), .dout(n25482));
    jdff dff_B_HdovCmk45_1(.din(n2358), .dout(n25485));
    jdff dff_B_Q8Jhx20V3_1(.din(n25485), .dout(n25488));
    jdff dff_B_uImFXF9W3_2(.din(n2036), .dout(n25491));
    jdff dff_B_Mzhg2ssD0_2(.din(n25491), .dout(n25494));
    jdff dff_B_ts3WuSzZ2_2(.din(n25494), .dout(n25497));
    jdff dff_B_vPj7a03l5_0(.din(n2055), .dout(n25500));
    jdff dff_A_KX7Rd5572_0(.din(n25505), .dout(n25502));
    jdff dff_A_rWc83jMO0_0(.din(n1728), .dout(n25505));
    jdff dff_A_gy46G8l43_1(.din(n25511), .dout(n25508));
    jdff dff_A_mOLit72c0_1(.din(n1728), .dout(n25511));
    jdff dff_B_s9lPq6nu2_1(.din(n6550), .dout(n25515));
    jdff dff_A_xWpozIyr6_1(.din(n6454), .dout(n25517));
    jdff dff_B_iOR8SBie2_1(.din(n6446), .dout(n25521));
    jdff dff_B_xvidG6BS0_2(.din(n6308), .dout(n25524));
    jdff dff_B_H2JOajln6_2(.din(n25524), .dout(n25527));
    jdff dff_B_Ycn68z6x2_2(.din(n25527), .dout(n25530));
    jdff dff_B_Qkicp0Nj0_2(.din(n25530), .dout(n25533));
    jdff dff_B_zlxqnU5T9_2(.din(n25533), .dout(n25536));
    jdff dff_B_mSDuYZpA9_2(.din(n25536), .dout(n25539));
    jdff dff_B_vmDLUHHK1_2(.din(n25539), .dout(n25542));
    jdff dff_B_eHd2FTqC3_2(.din(n25542), .dout(n25545));
    jdff dff_B_uBOGlqrS6_2(.din(n25545), .dout(n25548));
    jdff dff_B_gyLmnItY4_2(.din(n25548), .dout(n25551));
    jdff dff_B_A0NbFXRA3_2(.din(n25551), .dout(n25554));
    jdff dff_B_KZ3Pl0a95_2(.din(n25554), .dout(n25557));
    jdff dff_B_68pFLTaF9_2(.din(n25557), .dout(n25560));
    jdff dff_B_Nblkd6oV4_2(.din(n25560), .dout(n25563));
    jdff dff_B_msA6pmMP5_2(.din(n25563), .dout(n25566));
    jdff dff_B_OTPIfpTj9_2(.din(n25566), .dout(n25569));
    jdff dff_B_ThheJh362_2(.din(n25569), .dout(n25572));
    jdff dff_B_78wLyOoW3_2(.din(n25572), .dout(n25575));
    jdff dff_B_K1WphjVx7_2(.din(n25575), .dout(n25578));
    jdff dff_B_y3jsG4hi1_2(.din(n25578), .dout(n25581));
    jdff dff_B_wBCu0QuX0_2(.din(n25581), .dout(n25584));
    jdff dff_B_k9OXH5N45_2(.din(n25584), .dout(n25587));
    jdff dff_B_mcAs9FME2_2(.din(n25587), .dout(n25590));
    jdff dff_B_xzlCFREP8_2(.din(n25590), .dout(n25593));
    jdff dff_B_EFUzlIud0_2(.din(n25593), .dout(n25596));
    jdff dff_B_0yo6G0Im4_2(.din(n25596), .dout(n25599));
    jdff dff_B_KIwlVoas2_2(.din(n25599), .dout(n25602));
    jdff dff_B_usAQ4Qhc7_2(.din(n25602), .dout(n25605));
    jdff dff_B_QKoOKo823_2(.din(n25605), .dout(n25608));
    jdff dff_B_D7HvH2q07_2(.din(n25608), .dout(n25611));
    jdff dff_B_iZ8Cg2jB2_2(.din(n25611), .dout(n25614));
    jdff dff_B_XrxrqQa70_2(.din(n25614), .dout(n25617));
    jdff dff_B_AimAZ4rY5_2(.din(n25617), .dout(n25620));
    jdff dff_B_0mGKjRwK7_2(.din(n25620), .dout(n25623));
    jdff dff_B_SLqgLeUz6_2(.din(n25623), .dout(n25626));
    jdff dff_B_0Notq8cF1_2(.din(n25626), .dout(n25629));
    jdff dff_B_cmmxr5wm9_2(.din(n25629), .dout(n25632));
    jdff dff_B_HsDwihJM1_2(.din(n25632), .dout(n25635));
    jdff dff_B_kU29M0Bi9_2(.din(n25635), .dout(n25638));
    jdff dff_B_OO6lC5Ma8_2(.din(n25638), .dout(n25641));
    jdff dff_B_u8os5wxt0_2(.din(n25641), .dout(n25644));
    jdff dff_B_9aw1YUF01_2(.din(n25644), .dout(n25647));
    jdff dff_B_H41Oumqr2_2(.din(n25647), .dout(n25650));
    jdff dff_B_MLozTtSE3_2(.din(n25650), .dout(n25653));
    jdff dff_B_u2iNC7Yd9_2(.din(n25653), .dout(n25656));
    jdff dff_B_lFhYoAov1_2(.din(n25656), .dout(n25659));
    jdff dff_B_FFxwMcAg2_2(.din(n25659), .dout(n25662));
    jdff dff_B_4Kjf9Xzu5_2(.din(n25662), .dout(n25665));
    jdff dff_B_AUJVVuZs7_2(.din(n6320), .dout(n25668));
    jdff dff_B_rhnCP9QY2_1(.din(n6312), .dout(n25671));
    jdff dff_B_C7LHpqBI3_2(.din(n6150), .dout(n25674));
    jdff dff_B_UeWfbcrz7_2(.din(n25674), .dout(n25677));
    jdff dff_B_n4tpqdkJ5_2(.din(n25677), .dout(n25680));
    jdff dff_B_G7YogIVE9_2(.din(n25680), .dout(n25683));
    jdff dff_B_J8LjVr9Z2_2(.din(n25683), .dout(n25686));
    jdff dff_B_Y0KJbX4N0_2(.din(n25686), .dout(n25689));
    jdff dff_B_4qNiEXOt8_2(.din(n25689), .dout(n25692));
    jdff dff_B_9kFeaxVf5_2(.din(n25692), .dout(n25695));
    jdff dff_B_HsptdJyG0_2(.din(n25695), .dout(n25698));
    jdff dff_B_TKzAi6Gl3_2(.din(n25698), .dout(n25701));
    jdff dff_B_6ynsMQ2l0_2(.din(n25701), .dout(n25704));
    jdff dff_B_bhnIZjwp3_2(.din(n25704), .dout(n25707));
    jdff dff_B_tXVk6FcT9_2(.din(n25707), .dout(n25710));
    jdff dff_B_58LdgK666_2(.din(n25710), .dout(n25713));
    jdff dff_B_gzIk7S020_2(.din(n25713), .dout(n25716));
    jdff dff_B_szxKorJG7_2(.din(n25716), .dout(n25719));
    jdff dff_B_f5OiTOd96_2(.din(n25719), .dout(n25722));
    jdff dff_B_e6WLPQm50_2(.din(n25722), .dout(n25725));
    jdff dff_B_2F000M8A6_2(.din(n25725), .dout(n25728));
    jdff dff_B_IFocsjVe8_2(.din(n25728), .dout(n25731));
    jdff dff_B_1Y0NbcHw4_2(.din(n25731), .dout(n25734));
    jdff dff_B_8w1rBpYa0_2(.din(n25734), .dout(n25737));
    jdff dff_B_eGCw48JR6_2(.din(n25737), .dout(n25740));
    jdff dff_B_Ym96BF5n5_2(.din(n25740), .dout(n25743));
    jdff dff_B_7GNR9CiQ1_2(.din(n25743), .dout(n25746));
    jdff dff_B_jydhBZkv3_2(.din(n25746), .dout(n25749));
    jdff dff_B_XwbwARax8_2(.din(n25749), .dout(n25752));
    jdff dff_B_XUXLl9PZ6_2(.din(n25752), .dout(n25755));
    jdff dff_B_9s5BgiKq1_2(.din(n25755), .dout(n25758));
    jdff dff_B_cbhmIanl0_2(.din(n25758), .dout(n25761));
    jdff dff_B_53C2nhS84_2(.din(n25761), .dout(n25764));
    jdff dff_B_UbLtddzG5_2(.din(n25764), .dout(n25767));
    jdff dff_B_KsXZ429F1_2(.din(n25767), .dout(n25770));
    jdff dff_B_rrGJcutx6_2(.din(n25770), .dout(n25773));
    jdff dff_B_mdjShcxc7_2(.din(n25773), .dout(n25776));
    jdff dff_B_6MPxDqRq9_2(.din(n25776), .dout(n25779));
    jdff dff_B_Uj77CKxn5_2(.din(n25779), .dout(n25782));
    jdff dff_B_VDZ8DIOG4_2(.din(n25782), .dout(n25785));
    jdff dff_B_lS3yPT7e4_2(.din(n25785), .dout(n25788));
    jdff dff_B_8uBAOWGH5_2(.din(n25788), .dout(n25791));
    jdff dff_B_26cPxGU03_2(.din(n25791), .dout(n25794));
    jdff dff_B_LrqcIO5M8_2(.din(n25794), .dout(n25797));
    jdff dff_B_aE2A8Mk01_2(.din(n25797), .dout(n25800));
    jdff dff_B_x0b2LiBp2_2(.din(n25800), .dout(n25803));
    jdff dff_B_oh5mULbq1_2(.din(n6162), .dout(n25806));
    jdff dff_B_eWtrvpIs8_1(.din(n6154), .dout(n25809));
    jdff dff_B_SEXWdAiT6_2(.din(n5956), .dout(n25812));
    jdff dff_B_mNob9bnb3_2(.din(n25812), .dout(n25815));
    jdff dff_B_Rq2NlqbI9_2(.din(n25815), .dout(n25818));
    jdff dff_B_Mx0VVGVZ5_2(.din(n25818), .dout(n25821));
    jdff dff_B_dViLjMkg3_2(.din(n25821), .dout(n25824));
    jdff dff_B_2ZNy9ijD6_2(.din(n25824), .dout(n25827));
    jdff dff_B_zYGaFDGy4_2(.din(n25827), .dout(n25830));
    jdff dff_B_tEeN3z9T5_2(.din(n25830), .dout(n25833));
    jdff dff_B_AxSFZzne9_2(.din(n25833), .dout(n25836));
    jdff dff_B_tWQnD0L75_2(.din(n25836), .dout(n25839));
    jdff dff_B_sDYprePW0_2(.din(n25839), .dout(n25842));
    jdff dff_B_WQqs7YsP8_2(.din(n25842), .dout(n25845));
    jdff dff_B_OG5ng1w95_2(.din(n25845), .dout(n25848));
    jdff dff_B_MiR8bfbQ0_2(.din(n25848), .dout(n25851));
    jdff dff_B_YZLiTGSk0_2(.din(n25851), .dout(n25854));
    jdff dff_B_EnkYOP629_2(.din(n25854), .dout(n25857));
    jdff dff_B_Mr0QJ2Rl2_2(.din(n25857), .dout(n25860));
    jdff dff_B_7Sbwzsal4_2(.din(n25860), .dout(n25863));
    jdff dff_B_ZBxEJg4i8_2(.din(n25863), .dout(n25866));
    jdff dff_B_D6LTuJuE5_2(.din(n25866), .dout(n25869));
    jdff dff_B_saW3zqss9_2(.din(n25869), .dout(n25872));
    jdff dff_B_KcjWQJfm3_2(.din(n25872), .dout(n25875));
    jdff dff_B_i9E5E1I67_2(.din(n25875), .dout(n25878));
    jdff dff_B_JW1bkQxN0_2(.din(n25878), .dout(n25881));
    jdff dff_B_e2OkxWGi5_2(.din(n25881), .dout(n25884));
    jdff dff_B_xJhJw2nF1_2(.din(n25884), .dout(n25887));
    jdff dff_B_wXwwq99M3_2(.din(n25887), .dout(n25890));
    jdff dff_B_GbvRjd4Z4_2(.din(n25890), .dout(n25893));
    jdff dff_B_wEKKARbf3_2(.din(n25893), .dout(n25896));
    jdff dff_B_Apw4MyEK7_2(.din(n25896), .dout(n25899));
    jdff dff_B_vVS5O0Tl3_2(.din(n25899), .dout(n25902));
    jdff dff_B_bhfZ3va88_2(.din(n25902), .dout(n25905));
    jdff dff_B_P4om3MHF6_2(.din(n25905), .dout(n25908));
    jdff dff_B_ulKX7iad3_2(.din(n25908), .dout(n25911));
    jdff dff_B_7qJFgdvK6_2(.din(n25911), .dout(n25914));
    jdff dff_B_1c96IQu83_2(.din(n25914), .dout(n25917));
    jdff dff_B_9Dh0EJpF6_2(.din(n25917), .dout(n25920));
    jdff dff_B_wYij6kNY8_2(.din(n25920), .dout(n25923));
    jdff dff_B_4GVMkThx5_2(.din(n25923), .dout(n25926));
    jdff dff_B_KFTi04Gr6_2(.din(n25926), .dout(n25929));
    jdff dff_B_lTDcgB0E7_2(.din(n5968), .dout(n25932));
    jdff dff_B_EBXg5wWk4_1(.din(n5960), .dout(n25935));
    jdff dff_B_CS0Eygq89_2(.din(n5738), .dout(n25938));
    jdff dff_B_tZDpSqCR3_2(.din(n25938), .dout(n25941));
    jdff dff_B_KbDKyaV90_2(.din(n25941), .dout(n25944));
    jdff dff_B_aNfeVkdx7_2(.din(n25944), .dout(n25947));
    jdff dff_B_HjDldspW8_2(.din(n25947), .dout(n25950));
    jdff dff_B_vsXKsXhd8_2(.din(n25950), .dout(n25953));
    jdff dff_B_mworufgv5_2(.din(n25953), .dout(n25956));
    jdff dff_B_EAgftY1d4_2(.din(n25956), .dout(n25959));
    jdff dff_B_5mH1526m9_2(.din(n25959), .dout(n25962));
    jdff dff_B_MGMWnnIC6_2(.din(n25962), .dout(n25965));
    jdff dff_B_gsLYPoQi5_2(.din(n25965), .dout(n25968));
    jdff dff_B_EznCGRIn1_2(.din(n25968), .dout(n25971));
    jdff dff_B_CHsZoZUY8_2(.din(n25971), .dout(n25974));
    jdff dff_B_JsWHldx16_2(.din(n25974), .dout(n25977));
    jdff dff_B_LYm6CVXr4_2(.din(n25977), .dout(n25980));
    jdff dff_B_jWypSJo20_2(.din(n25980), .dout(n25983));
    jdff dff_B_Sqw4sEgo6_2(.din(n25983), .dout(n25986));
    jdff dff_B_kVl59ngq4_2(.din(n25986), .dout(n25989));
    jdff dff_B_k48YUVn62_2(.din(n25989), .dout(n25992));
    jdff dff_B_JXehVPJs1_2(.din(n25992), .dout(n25995));
    jdff dff_B_d9IGH2WH9_2(.din(n25995), .dout(n25998));
    jdff dff_B_EFMcX0Bi4_2(.din(n25998), .dout(n26001));
    jdff dff_B_pBk6d6VG7_2(.din(n26001), .dout(n26004));
    jdff dff_B_B7dy0SCz9_2(.din(n26004), .dout(n26007));
    jdff dff_B_wV1OtUmf9_2(.din(n26007), .dout(n26010));
    jdff dff_B_0fkp3bTY3_2(.din(n26010), .dout(n26013));
    jdff dff_B_Jug4uxFi6_2(.din(n26013), .dout(n26016));
    jdff dff_B_dHAEEWK13_2(.din(n26016), .dout(n26019));
    jdff dff_B_fQPqUJfB7_2(.din(n26019), .dout(n26022));
    jdff dff_B_dsG3ScMA0_2(.din(n26022), .dout(n26025));
    jdff dff_B_xXtdYtIG7_2(.din(n26025), .dout(n26028));
    jdff dff_B_MJMUtV6s6_2(.din(n26028), .dout(n26031));
    jdff dff_B_JAChyVXO1_2(.din(n26031), .dout(n26034));
    jdff dff_B_cC53jNmb5_2(.din(n26034), .dout(n26037));
    jdff dff_B_Ypjycl5A1_2(.din(n26037), .dout(n26040));
    jdff dff_B_Qs83rpz59_2(.din(n26040), .dout(n26043));
    jdff dff_B_g95BrBah1_2(.din(n5750), .dout(n26046));
    jdff dff_B_kTo0wJwr9_1(.din(n5742), .dout(n26049));
    jdff dff_B_xXfvTIEd0_2(.din(n5493), .dout(n26052));
    jdff dff_B_ctNTb8Vz8_2(.din(n26052), .dout(n26055));
    jdff dff_B_OYTBoBDN5_2(.din(n26055), .dout(n26058));
    jdff dff_B_sxvJC70M6_2(.din(n26058), .dout(n26061));
    jdff dff_B_x7kPA3hh2_2(.din(n26061), .dout(n26064));
    jdff dff_B_A0qOBcfU0_2(.din(n26064), .dout(n26067));
    jdff dff_B_dNMv3fYf8_2(.din(n26067), .dout(n26070));
    jdff dff_B_MLygmdTh6_2(.din(n26070), .dout(n26073));
    jdff dff_B_qHf0FhW84_2(.din(n26073), .dout(n26076));
    jdff dff_B_hG1YzoXd2_2(.din(n26076), .dout(n26079));
    jdff dff_B_EyEr9Flw2_2(.din(n26079), .dout(n26082));
    jdff dff_B_Yq8VIdSQ8_2(.din(n26082), .dout(n26085));
    jdff dff_B_Gku1QtqH0_2(.din(n26085), .dout(n26088));
    jdff dff_B_RNxEJiZe6_2(.din(n26088), .dout(n26091));
    jdff dff_B_m2PhG3Yg5_2(.din(n26091), .dout(n26094));
    jdff dff_B_LxhWNwgI0_2(.din(n26094), .dout(n26097));
    jdff dff_B_l56bxpkC6_2(.din(n26097), .dout(n26100));
    jdff dff_B_YpCP5Imj6_2(.din(n26100), .dout(n26103));
    jdff dff_B_Bf7M6seD1_2(.din(n26103), .dout(n26106));
    jdff dff_B_MmXmCIyY0_2(.din(n26106), .dout(n26109));
    jdff dff_B_Spc6bhKa1_2(.din(n26109), .dout(n26112));
    jdff dff_B_r5cNsBke1_2(.din(n26112), .dout(n26115));
    jdff dff_B_nHrTzs1x6_2(.din(n26115), .dout(n26118));
    jdff dff_B_z8BuF0Ov7_2(.din(n26118), .dout(n26121));
    jdff dff_B_Qy6Ze7tF0_2(.din(n26121), .dout(n26124));
    jdff dff_B_g8XNXJmE1_2(.din(n26124), .dout(n26127));
    jdff dff_B_YcrhXcAJ0_2(.din(n26127), .dout(n26130));
    jdff dff_B_DyvprqCN1_2(.din(n26130), .dout(n26133));
    jdff dff_B_iVPqHczQ2_2(.din(n26133), .dout(n26136));
    jdff dff_B_Ui4cwZhr5_2(.din(n26136), .dout(n26139));
    jdff dff_B_ugUEf2eZ9_2(.din(n26139), .dout(n26142));
    jdff dff_B_6ZFVxRWY6_2(.din(n26142), .dout(n26145));
    jdff dff_B_IFTw00kJ0_1(.din(n5497), .dout(n26148));
    jdff dff_B_RdtKvNYk3_2(.din(n5221), .dout(n26151));
    jdff dff_B_PYP44jYz2_2(.din(n26151), .dout(n26154));
    jdff dff_B_VC9rdrPe5_2(.din(n26154), .dout(n26157));
    jdff dff_B_683VvSZM6_2(.din(n26157), .dout(n26160));
    jdff dff_B_HDIY0YNw2_2(.din(n26160), .dout(n26163));
    jdff dff_B_alUXG5IP2_2(.din(n26163), .dout(n26166));
    jdff dff_B_SH10VcSh0_2(.din(n26166), .dout(n26169));
    jdff dff_B_7aTyqGo02_2(.din(n26169), .dout(n26172));
    jdff dff_B_plSKXuKT6_2(.din(n26172), .dout(n26175));
    jdff dff_B_EPFTNTCF3_2(.din(n26175), .dout(n26178));
    jdff dff_B_Aqhfj5nR5_2(.din(n26178), .dout(n26181));
    jdff dff_B_YfFf0rx90_2(.din(n26181), .dout(n26184));
    jdff dff_B_59uJ2E770_2(.din(n26184), .dout(n26187));
    jdff dff_B_NU8mHIPF2_2(.din(n26187), .dout(n26190));
    jdff dff_B_Nh5cQURV0_2(.din(n26190), .dout(n26193));
    jdff dff_B_Qwg1tJgI4_2(.din(n26193), .dout(n26196));
    jdff dff_B_oBTCs1Ic9_2(.din(n26196), .dout(n26199));
    jdff dff_B_XklLRYk78_2(.din(n26199), .dout(n26202));
    jdff dff_B_GPxNX4dw3_2(.din(n26202), .dout(n26205));
    jdff dff_B_jDbtH2FR7_2(.din(n26205), .dout(n26208));
    jdff dff_B_7ezMDUGa6_2(.din(n26208), .dout(n26211));
    jdff dff_B_ieCxqmrM1_2(.din(n26211), .dout(n26214));
    jdff dff_B_58kcIXwr5_2(.din(n26214), .dout(n26217));
    jdff dff_B_jgVScGte7_2(.din(n26217), .dout(n26220));
    jdff dff_B_kVei2QwS4_2(.din(n26220), .dout(n26223));
    jdff dff_B_G6KMSaKk6_2(.din(n26223), .dout(n26226));
    jdff dff_B_0MYWOVCF2_2(.din(n26226), .dout(n26229));
    jdff dff_B_RqFGWpq18_2(.din(n26229), .dout(n26232));
    jdff dff_B_SaWBszGf8_2(.din(n26232), .dout(n26235));
    jdff dff_B_DMjZiILv3_2(.din(n5318), .dout(n26238));
    jdff dff_B_P7pV3xtN2_1(.din(n5225), .dout(n26241));
    jdff dff_B_cAv5JQXD4_2(.din(n4922), .dout(n26244));
    jdff dff_B_Ci97n3TX3_2(.din(n26244), .dout(n26247));
    jdff dff_B_QUZc3E899_2(.din(n26247), .dout(n26250));
    jdff dff_B_OXQttdKS8_2(.din(n26250), .dout(n26253));
    jdff dff_B_MrVLvbVi6_2(.din(n26253), .dout(n26256));
    jdff dff_B_2r5jHqnC5_2(.din(n26256), .dout(n26259));
    jdff dff_B_yNIcBTNp0_2(.din(n26259), .dout(n26262));
    jdff dff_B_uLGDsaIN0_2(.din(n26262), .dout(n26265));
    jdff dff_B_y1WSSNpM2_2(.din(n26265), .dout(n26268));
    jdff dff_B_YtGwdiAQ3_2(.din(n26268), .dout(n26271));
    jdff dff_B_qe8iiywU7_2(.din(n26271), .dout(n26274));
    jdff dff_B_6l0Wpm4N9_2(.din(n26274), .dout(n26277));
    jdff dff_B_VZVm6zFy0_2(.din(n26277), .dout(n26280));
    jdff dff_B_q2C1g8q56_2(.din(n26280), .dout(n26283));
    jdff dff_B_boap64Cn4_2(.din(n26283), .dout(n26286));
    jdff dff_B_oxSfq6k95_2(.din(n26286), .dout(n26289));
    jdff dff_B_WVnCnoJi5_2(.din(n26289), .dout(n26292));
    jdff dff_B_Q0dkQHni8_2(.din(n26292), .dout(n26295));
    jdff dff_B_xlSSTIkI9_2(.din(n26295), .dout(n26298));
    jdff dff_B_rUa4M8Eg4_2(.din(n26298), .dout(n26301));
    jdff dff_B_OTarkhj05_2(.din(n26301), .dout(n26304));
    jdff dff_B_Xh3xVpyD0_2(.din(n26304), .dout(n26307));
    jdff dff_B_7AhYg2xx1_2(.din(n26307), .dout(n26310));
    jdff dff_B_IDndbqFh3_2(.din(n26310), .dout(n26313));
    jdff dff_B_MbvSBqjA3_2(.din(n26313), .dout(n26316));
    jdff dff_B_59Rap77Z8_2(.din(n26316), .dout(n26319));
    jdff dff_B_8SaeRHr09_2(.din(n5019), .dout(n26322));
    jdff dff_B_fvBuavZm2_1(.din(n4926), .dout(n26325));
    jdff dff_B_rikRDUoQ1_2(.din(n4596), .dout(n26328));
    jdff dff_B_ODqYfBd60_2(.din(n26328), .dout(n26331));
    jdff dff_B_stjmCUix9_2(.din(n26331), .dout(n26334));
    jdff dff_B_W1CnToUL2_2(.din(n26334), .dout(n26337));
    jdff dff_B_nQibsh9b1_2(.din(n26337), .dout(n26340));
    jdff dff_B_kKp3HgM66_2(.din(n26340), .dout(n26343));
    jdff dff_B_umLtDdPn9_2(.din(n26343), .dout(n26346));
    jdff dff_B_BPR8izXS1_2(.din(n26346), .dout(n26349));
    jdff dff_B_qkOfTQAf0_2(.din(n26349), .dout(n26352));
    jdff dff_B_WLXmD37M5_2(.din(n26352), .dout(n26355));
    jdff dff_B_1jGcuY3J0_2(.din(n26355), .dout(n26358));
    jdff dff_B_MssQaZhz4_2(.din(n26358), .dout(n26361));
    jdff dff_B_4Y6TmLK67_2(.din(n26361), .dout(n26364));
    jdff dff_B_aI1Fc56f5_2(.din(n26364), .dout(n26367));
    jdff dff_B_3pmW3EdN4_2(.din(n26367), .dout(n26370));
    jdff dff_B_72SL8DNq3_2(.din(n26370), .dout(n26373));
    jdff dff_B_LGk9zbWS5_2(.din(n26373), .dout(n26376));
    jdff dff_B_O5NBdmpQ8_2(.din(n26376), .dout(n26379));
    jdff dff_B_2AiuQ0aa5_2(.din(n26379), .dout(n26382));
    jdff dff_B_R4gBO1sg1_2(.din(n26382), .dout(n26385));
    jdff dff_B_6S7DUVKu4_2(.din(n26385), .dout(n26388));
    jdff dff_B_s3V2nT0A2_2(.din(n26388), .dout(n26391));
    jdff dff_B_mIQobraJ3_2(.din(n26391), .dout(n26394));
    jdff dff_B_FU4KmCfZ3_2(.din(n4693), .dout(n26397));
    jdff dff_B_8eTcrcM07_1(.din(n4600), .dout(n26400));
    jdff dff_B_BpDJCnWy6_2(.din(n4246), .dout(n26403));
    jdff dff_B_c4Ac7gBD1_2(.din(n26403), .dout(n26406));
    jdff dff_B_q5sa0PWj0_2(.din(n26406), .dout(n26409));
    jdff dff_B_embPnHVU0_2(.din(n26409), .dout(n26412));
    jdff dff_B_VdXsQq5V5_2(.din(n26412), .dout(n26415));
    jdff dff_B_ClWm7J4h1_2(.din(n26415), .dout(n26418));
    jdff dff_B_96uQTumw9_2(.din(n26418), .dout(n26421));
    jdff dff_B_ZlA23hll0_2(.din(n26421), .dout(n26424));
    jdff dff_B_8DPtsfbq1_2(.din(n26424), .dout(n26427));
    jdff dff_B_1qKzQJJP8_2(.din(n26427), .dout(n26430));
    jdff dff_B_M0w7T2lc0_2(.din(n26430), .dout(n26433));
    jdff dff_B_mBifnvAS7_2(.din(n26433), .dout(n26436));
    jdff dff_B_8JcM7pM71_2(.din(n26436), .dout(n26439));
    jdff dff_B_EwOgen9I2_2(.din(n26439), .dout(n26442));
    jdff dff_B_Vcf7JBKS5_2(.din(n26442), .dout(n26445));
    jdff dff_B_e7VYbVbi1_2(.din(n26445), .dout(n26448));
    jdff dff_B_9pHvuOoV7_2(.din(n26448), .dout(n26451));
    jdff dff_B_83EA3s7T5_2(.din(n26451), .dout(n26454));
    jdff dff_B_V6q3kUu22_2(.din(n26454), .dout(n26457));
    jdff dff_B_sx23HeQZ2_2(.din(n26457), .dout(n26460));
    jdff dff_B_aZm2xLBW4_2(.din(n4343), .dout(n26463));
    jdff dff_B_S4B5uJt66_1(.din(n4250), .dout(n26466));
    jdff dff_B_WJNUuhNB8_2(.din(n3870), .dout(n26469));
    jdff dff_B_ErLCSPMA9_2(.din(n26469), .dout(n26472));
    jdff dff_B_3U4Xjlvm5_2(.din(n26472), .dout(n26475));
    jdff dff_B_7nm19qju8_2(.din(n26475), .dout(n26478));
    jdff dff_B_3fJvhWbh9_2(.din(n26478), .dout(n26481));
    jdff dff_B_oSfWurtQ4_2(.din(n26481), .dout(n26484));
    jdff dff_B_f4WRCaVE0_2(.din(n26484), .dout(n26487));
    jdff dff_B_2Mtrg2IV3_2(.din(n26487), .dout(n26490));
    jdff dff_B_1F4gxY6Q7_2(.din(n26490), .dout(n26493));
    jdff dff_B_NuWwU2qs6_2(.din(n26493), .dout(n26496));
    jdff dff_B_MIncjyIH1_2(.din(n26496), .dout(n26499));
    jdff dff_B_ZgAoVJIJ3_2(.din(n26499), .dout(n26502));
    jdff dff_B_efVkfXK28_2(.din(n26502), .dout(n26505));
    jdff dff_B_kFYl820U7_2(.din(n26505), .dout(n26508));
    jdff dff_B_M8n77AtN2_2(.din(n26508), .dout(n26511));
    jdff dff_B_qFN8LtCW0_2(.din(n26511), .dout(n26514));
    jdff dff_B_7weLBBiR8_2(.din(n26514), .dout(n26517));
    jdff dff_B_3TVnsZem2_2(.din(n3963), .dout(n26520));
    jdff dff_B_tEIsuwSY6_1(.din(n3874), .dout(n26523));
    jdff dff_B_7D12UUX70_2(.din(n3490), .dout(n26526));
    jdff dff_B_eHnnMSzG1_2(.din(n26526), .dout(n26529));
    jdff dff_B_S24SvMsw7_2(.din(n26529), .dout(n26532));
    jdff dff_B_345aMDvI1_2(.din(n26532), .dout(n26535));
    jdff dff_B_oLj4Ws795_2(.din(n26535), .dout(n26538));
    jdff dff_B_bq8Tivif7_2(.din(n26538), .dout(n26541));
    jdff dff_B_PKtjp3DY0_2(.din(n26541), .dout(n26544));
    jdff dff_B_D8Aa3MQq6_2(.din(n26544), .dout(n26547));
    jdff dff_B_kwYhMsJa9_2(.din(n26547), .dout(n26550));
    jdff dff_B_ShhZK4Dh8_2(.din(n26550), .dout(n26553));
    jdff dff_B_BrJCwibb1_2(.din(n26553), .dout(n26556));
    jdff dff_B_R3ndHCbo9_2(.din(n26556), .dout(n26559));
    jdff dff_B_YR6wcwMd9_2(.din(n26559), .dout(n26562));
    jdff dff_B_0qnDpiRu7_2(.din(n26562), .dout(n26565));
    jdff dff_B_8aMSco662_2(.din(n3580), .dout(n26568));
    jdff dff_B_dvYDu3121_1(.din(n3494), .dout(n26571));
    jdff dff_B_sGKYpW7A1_2(.din(n3099), .dout(n26574));
    jdff dff_B_bfIW92sH1_2(.din(n26574), .dout(n26577));
    jdff dff_B_Fsgw87Dp9_2(.din(n26577), .dout(n26580));
    jdff dff_B_9T1ypWOQ6_2(.din(n26580), .dout(n26583));
    jdff dff_B_OcvriUyv4_2(.din(n26583), .dout(n26586));
    jdff dff_B_1L2foCBo2_2(.din(n26586), .dout(n26589));
    jdff dff_B_dbicMcUa1_2(.din(n26589), .dout(n26592));
    jdff dff_B_2INhwtRo7_2(.din(n26592), .dout(n26595));
    jdff dff_B_WjTeDR5t1_2(.din(n26595), .dout(n26598));
    jdff dff_B_lhZez3Wi3_2(.din(n26598), .dout(n26601));
    jdff dff_B_lEt3Fjqo3_2(.din(n26601), .dout(n26604));
    jdff dff_B_Vd6fMmaD0_2(.din(n3175), .dout(n26607));
    jdff dff_B_rX2M1cWh8_1(.din(n3103), .dout(n26610));
    jdff dff_B_c50el4ku7_2(.din(n2724), .dout(n26613));
    jdff dff_B_c98Z24RB0_2(.din(n26613), .dout(n26616));
    jdff dff_B_h0AshvrR1_2(.din(n26616), .dout(n26619));
    jdff dff_B_Cl50itll5_2(.din(n26619), .dout(n26622));
    jdff dff_B_lq4ZSHCx9_2(.din(n26622), .dout(n26625));
    jdff dff_B_I93lvMkg4_2(.din(n26625), .dout(n26628));
    jdff dff_B_oe9DYwCn9_2(.din(n26628), .dout(n26631));
    jdff dff_B_GURg5o5w9_2(.din(n26631), .dout(n26634));
    jdff dff_B_VI1NDn6o2_2(.din(n2780), .dout(n26637));
    jdff dff_B_ifZxfT5A3_2(.din(n26637), .dout(n26640));
    jdff dff_B_9WGQxfkY6_2(.din(n26640), .dout(n26643));
    jdff dff_B_kuP3yNXd4_1(.din(n2728), .dout(n26646));
    jdff dff_B_6JvFeimc6_1(.din(n26646), .dout(n26649));
    jdff dff_B_j4e8ueRL0_2(.din(n2379), .dout(n26652));
    jdff dff_B_bJXOhhWn9_2(.din(n26652), .dout(n26655));
    jdff dff_B_3QPnI6HQ7_2(.din(n26655), .dout(n26658));
    jdff dff_B_P53qelmo0_0(.din(n2398), .dout(n26661));
    jdff dff_A_46UlZCZ00_0(.din(n26666), .dout(n26663));
    jdff dff_A_Y85roqRL0_0(.din(n2044), .dout(n26666));
    jdff dff_A_c6VNpxpW0_1(.din(n26672), .dout(n26669));
    jdff dff_A_as2XVWPH6_1(.din(n2044), .dout(n26672));
    jdff dff_B_IuxRMeHR7_1(.din(n6649), .dout(n26676));
    jdff dff_A_XICyd0S42_1(.din(n6580), .dout(n26678));
    jdff dff_B_cNIx8qef4_1(.din(n6572), .dout(n26682));
    jdff dff_B_5VH3S5KC4_2(.din(n6461), .dout(n26685));
    jdff dff_B_eonfFV8u8_2(.din(n26685), .dout(n26688));
    jdff dff_B_56vQnV2A8_2(.din(n26688), .dout(n26691));
    jdff dff_B_eO0lWiz65_2(.din(n26691), .dout(n26694));
    jdff dff_B_oC8nM5Yi5_2(.din(n26694), .dout(n26697));
    jdff dff_B_vwgx5DcS3_2(.din(n26697), .dout(n26700));
    jdff dff_B_fFVJZIG67_2(.din(n26700), .dout(n26703));
    jdff dff_B_d4FGOjfo9_2(.din(n26703), .dout(n26706));
    jdff dff_B_UILQIAy54_2(.din(n26706), .dout(n26709));
    jdff dff_B_KoF4gMht1_2(.din(n26709), .dout(n26712));
    jdff dff_B_Wn5ugI7L7_2(.din(n26712), .dout(n26715));
    jdff dff_B_rjqHnoJX9_2(.din(n26715), .dout(n26718));
    jdff dff_B_n6GBJcvL2_2(.din(n26718), .dout(n26721));
    jdff dff_B_Dt4sJqKx5_2(.din(n26721), .dout(n26724));
    jdff dff_B_BJI9yP0M9_2(.din(n26724), .dout(n26727));
    jdff dff_B_vrLlW9cl6_2(.din(n26727), .dout(n26730));
    jdff dff_B_3LRHKtQS9_2(.din(n26730), .dout(n26733));
    jdff dff_B_aCKGDVyq4_2(.din(n26733), .dout(n26736));
    jdff dff_B_ORugJqgg6_2(.din(n26736), .dout(n26739));
    jdff dff_B_5efZ3p6X7_2(.din(n26739), .dout(n26742));
    jdff dff_B_UwK4YVAB1_2(.din(n26742), .dout(n26745));
    jdff dff_B_euxLNvD36_2(.din(n26745), .dout(n26748));
    jdff dff_B_Dd2Sk7f24_2(.din(n26748), .dout(n26751));
    jdff dff_B_LVENd3dJ2_2(.din(n26751), .dout(n26754));
    jdff dff_B_73vxsRqY7_2(.din(n26754), .dout(n26757));
    jdff dff_B_lwlF5osT4_2(.din(n26757), .dout(n26760));
    jdff dff_B_E2oGo5wO3_2(.din(n26760), .dout(n26763));
    jdff dff_B_0ECbxJA31_2(.din(n26763), .dout(n26766));
    jdff dff_B_X4oyjOEb6_2(.din(n26766), .dout(n26769));
    jdff dff_B_mhVll2lE1_2(.din(n26769), .dout(n26772));
    jdff dff_B_f6oVvfJU1_2(.din(n26772), .dout(n26775));
    jdff dff_B_kyuORWib9_2(.din(n26775), .dout(n26778));
    jdff dff_B_xPcuBZK88_2(.din(n26778), .dout(n26781));
    jdff dff_B_5PC7VOl03_2(.din(n26781), .dout(n26784));
    jdff dff_B_u6CBGsXu3_2(.din(n26784), .dout(n26787));
    jdff dff_B_Jd60A3Jd8_2(.din(n26787), .dout(n26790));
    jdff dff_B_4ugWdidr7_2(.din(n26790), .dout(n26793));
    jdff dff_B_Wv25tivg8_2(.din(n26793), .dout(n26796));
    jdff dff_B_Fcmq35nS5_2(.din(n26796), .dout(n26799));
    jdff dff_B_6bRSeZ6Y0_2(.din(n26799), .dout(n26802));
    jdff dff_B_k9zFCfFa8_2(.din(n26802), .dout(n26805));
    jdff dff_B_UIxhGLUA5_2(.din(n26805), .dout(n26808));
    jdff dff_B_eTtUuq7z1_2(.din(n26808), .dout(n26811));
    jdff dff_B_eG0Dg59U6_2(.din(n26811), .dout(n26814));
    jdff dff_B_QtGIqCeq3_2(.din(n26814), .dout(n26817));
    jdff dff_B_Vd1YzWeS3_2(.din(n26817), .dout(n26820));
    jdff dff_B_Eq8KXynb3_2(.din(n26820), .dout(n26823));
    jdff dff_B_42Kb9K9Y3_2(.din(n26823), .dout(n26826));
    jdff dff_B_wOQWxcFM9_2(.din(n26826), .dout(n26829));
    jdff dff_B_kZfnxLQn1_2(.din(n26829), .dout(n26832));
    jdff dff_B_XI9aL1kA6_2(.din(n6473), .dout(n26835));
    jdff dff_B_YZ2J9A3L8_1(.din(n6465), .dout(n26838));
    jdff dff_B_qmakESc91_2(.din(n6327), .dout(n26841));
    jdff dff_B_eu2GnKC27_2(.din(n26841), .dout(n26844));
    jdff dff_B_PwLcmGNU4_2(.din(n26844), .dout(n26847));
    jdff dff_B_WAsqVksa8_2(.din(n26847), .dout(n26850));
    jdff dff_B_6WIRJcBQ2_2(.din(n26850), .dout(n26853));
    jdff dff_B_BhEidsID0_2(.din(n26853), .dout(n26856));
    jdff dff_B_GbCx0CF75_2(.din(n26856), .dout(n26859));
    jdff dff_B_PLhHUix31_2(.din(n26859), .dout(n26862));
    jdff dff_B_Gu0HUX2A1_2(.din(n26862), .dout(n26865));
    jdff dff_B_Sn5Vhz4B5_2(.din(n26865), .dout(n26868));
    jdff dff_B_FuwVTXdU6_2(.din(n26868), .dout(n26871));
    jdff dff_B_1rVF39iu2_2(.din(n26871), .dout(n26874));
    jdff dff_B_KsixzHA04_2(.din(n26874), .dout(n26877));
    jdff dff_B_fYltOazL9_2(.din(n26877), .dout(n26880));
    jdff dff_B_GK1aQCcu0_2(.din(n26880), .dout(n26883));
    jdff dff_B_eMqGJ8F13_2(.din(n26883), .dout(n26886));
    jdff dff_B_3zEYds2h1_2(.din(n26886), .dout(n26889));
    jdff dff_B_gcFnD3vg5_2(.din(n26889), .dout(n26892));
    jdff dff_B_rgjRzDTl7_2(.din(n26892), .dout(n26895));
    jdff dff_B_FGUL7rSd9_2(.din(n26895), .dout(n26898));
    jdff dff_B_AE4XgTMc7_2(.din(n26898), .dout(n26901));
    jdff dff_B_OpgnOYYm3_2(.din(n26901), .dout(n26904));
    jdff dff_B_GLwLq8Om5_2(.din(n26904), .dout(n26907));
    jdff dff_B_8IGFw4n75_2(.din(n26907), .dout(n26910));
    jdff dff_B_o3nhPfho0_2(.din(n26910), .dout(n26913));
    jdff dff_B_aBT5OuNh7_2(.din(n26913), .dout(n26916));
    jdff dff_B_NS0kfxfQ2_2(.din(n26916), .dout(n26919));
    jdff dff_B_emF6X8te7_2(.din(n26919), .dout(n26922));
    jdff dff_B_s1XKdGf11_2(.din(n26922), .dout(n26925));
    jdff dff_B_t5twnAwt4_2(.din(n26925), .dout(n26928));
    jdff dff_B_RWA8z1rd4_2(.din(n26928), .dout(n26931));
    jdff dff_B_tGQ1HdrO5_2(.din(n26931), .dout(n26934));
    jdff dff_B_cnVcqDy19_2(.din(n26934), .dout(n26937));
    jdff dff_B_YcoEt3Rc4_2(.din(n26937), .dout(n26940));
    jdff dff_B_Ke7e9Ui86_2(.din(n26940), .dout(n26943));
    jdff dff_B_8OtDWy1P2_2(.din(n26943), .dout(n26946));
    jdff dff_B_sG4f9neP9_2(.din(n26946), .dout(n26949));
    jdff dff_B_JRXAlELz5_2(.din(n26949), .dout(n26952));
    jdff dff_B_XoZAkpvS4_2(.din(n26952), .dout(n26955));
    jdff dff_B_LWMAvW8f8_2(.din(n26955), .dout(n26958));
    jdff dff_B_32XNziaG7_2(.din(n26958), .dout(n26961));
    jdff dff_B_zULAgVPI8_2(.din(n26961), .dout(n26964));
    jdff dff_B_Dc2eUq571_2(.din(n26964), .dout(n26967));
    jdff dff_B_9yEx8lTI4_2(.din(n26967), .dout(n26970));
    jdff dff_B_7wcgc0jE1_2(.din(n26970), .dout(n26973));
    jdff dff_B_R2b2iea10_2(.din(n26973), .dout(n26976));
    jdff dff_B_9JNkZehn3_2(.din(n6339), .dout(n26979));
    jdff dff_B_qIxe3vd75_1(.din(n6331), .dout(n26982));
    jdff dff_B_NVfbZG8w5_2(.din(n6169), .dout(n26985));
    jdff dff_B_q31nTGiS3_2(.din(n26985), .dout(n26988));
    jdff dff_B_yj1Oysll0_2(.din(n26988), .dout(n26991));
    jdff dff_B_NNh7bi0w6_2(.din(n26991), .dout(n26994));
    jdff dff_B_OMaqo4Ru2_2(.din(n26994), .dout(n26997));
    jdff dff_B_XHID7XCf1_2(.din(n26997), .dout(n27000));
    jdff dff_B_MOkMZ7Md9_2(.din(n27000), .dout(n27003));
    jdff dff_B_s9qYIOlf6_2(.din(n27003), .dout(n27006));
    jdff dff_B_9wN18sTM0_2(.din(n27006), .dout(n27009));
    jdff dff_B_nAWgq8vi1_2(.din(n27009), .dout(n27012));
    jdff dff_B_ZGYvdwqG6_2(.din(n27012), .dout(n27015));
    jdff dff_B_BwM7BUln4_2(.din(n27015), .dout(n27018));
    jdff dff_B_3DYt0mkP2_2(.din(n27018), .dout(n27021));
    jdff dff_B_TjitmiLP6_2(.din(n27021), .dout(n27024));
    jdff dff_B_B6KatWc69_2(.din(n27024), .dout(n27027));
    jdff dff_B_jJyY4cTE7_2(.din(n27027), .dout(n27030));
    jdff dff_B_ZDJN93Bu5_2(.din(n27030), .dout(n27033));
    jdff dff_B_4ybuubSP4_2(.din(n27033), .dout(n27036));
    jdff dff_B_qYAC7WbY1_2(.din(n27036), .dout(n27039));
    jdff dff_B_HYOiJHHU0_2(.din(n27039), .dout(n27042));
    jdff dff_B_slKoBVAO3_2(.din(n27042), .dout(n27045));
    jdff dff_B_v73g2qe33_2(.din(n27045), .dout(n27048));
    jdff dff_B_RRwZcDg88_2(.din(n27048), .dout(n27051));
    jdff dff_B_v7PMVfU24_2(.din(n27051), .dout(n27054));
    jdff dff_B_Ig3GQaC66_2(.din(n27054), .dout(n27057));
    jdff dff_B_UH5SJ1ty1_2(.din(n27057), .dout(n27060));
    jdff dff_B_gbY1j1Mp7_2(.din(n27060), .dout(n27063));
    jdff dff_B_Nan30Hjt2_2(.din(n27063), .dout(n27066));
    jdff dff_B_9PByZS5W8_2(.din(n27066), .dout(n27069));
    jdff dff_B_qwSj470X6_2(.din(n27069), .dout(n27072));
    jdff dff_B_9MKSPDSP3_2(.din(n27072), .dout(n27075));
    jdff dff_B_u8vTxEML2_2(.din(n27075), .dout(n27078));
    jdff dff_B_YXpqEmOj2_2(.din(n27078), .dout(n27081));
    jdff dff_B_9j7eYWqM0_2(.din(n27081), .dout(n27084));
    jdff dff_B_I7XImHNI4_2(.din(n27084), .dout(n27087));
    jdff dff_B_z9Rgkd8u4_2(.din(n27087), .dout(n27090));
    jdff dff_B_0pDl5VBX2_2(.din(n27090), .dout(n27093));
    jdff dff_B_ZkHN4mcn7_2(.din(n27093), .dout(n27096));
    jdff dff_B_JfmcWgGP3_2(.din(n27096), .dout(n27099));
    jdff dff_B_R82lrEbb0_2(.din(n27099), .dout(n27102));
    jdff dff_B_VDz2SiDw3_2(.din(n27102), .dout(n27105));
    jdff dff_B_QBDy5FYn6_2(.din(n27105), .dout(n27108));
    jdff dff_B_uQ6Ji3YS2_2(.din(n6181), .dout(n27111));
    jdff dff_B_2UH6Sju27_1(.din(n6173), .dout(n27114));
    jdff dff_B_KPqezL1z7_2(.din(n5975), .dout(n27117));
    jdff dff_B_LKVCHkt39_2(.din(n27117), .dout(n27120));
    jdff dff_B_Kub1RPoA5_2(.din(n27120), .dout(n27123));
    jdff dff_B_KxCVWRow4_2(.din(n27123), .dout(n27126));
    jdff dff_B_CCr9oJcR6_2(.din(n27126), .dout(n27129));
    jdff dff_B_BgfVez5E5_2(.din(n27129), .dout(n27132));
    jdff dff_B_JvFE5xG48_2(.din(n27132), .dout(n27135));
    jdff dff_B_wAeifTfD6_2(.din(n27135), .dout(n27138));
    jdff dff_B_r7SEr9GN3_2(.din(n27138), .dout(n27141));
    jdff dff_B_iWc8oDqp6_2(.din(n27141), .dout(n27144));
    jdff dff_B_PjOst9vO6_2(.din(n27144), .dout(n27147));
    jdff dff_B_KFSz1UYg8_2(.din(n27147), .dout(n27150));
    jdff dff_B_stk4p4U24_2(.din(n27150), .dout(n27153));
    jdff dff_B_LzvV4MbZ0_2(.din(n27153), .dout(n27156));
    jdff dff_B_SZIE7ewA0_2(.din(n27156), .dout(n27159));
    jdff dff_B_PSpzbNGq7_2(.din(n27159), .dout(n27162));
    jdff dff_B_6wEnHQ3O8_2(.din(n27162), .dout(n27165));
    jdff dff_B_9rBjxFsq1_2(.din(n27165), .dout(n27168));
    jdff dff_B_3QJIp8YZ9_2(.din(n27168), .dout(n27171));
    jdff dff_B_Yjt6tcos6_2(.din(n27171), .dout(n27174));
    jdff dff_B_nc5pdmiF8_2(.din(n27174), .dout(n27177));
    jdff dff_B_QDHaZHBr1_2(.din(n27177), .dout(n27180));
    jdff dff_B_g9QSn8kA9_2(.din(n27180), .dout(n27183));
    jdff dff_B_zzJ2wYow2_2(.din(n27183), .dout(n27186));
    jdff dff_B_xJW8AOW98_2(.din(n27186), .dout(n27189));
    jdff dff_B_YLOkRTk84_2(.din(n27189), .dout(n27192));
    jdff dff_B_c8afeDPF4_2(.din(n27192), .dout(n27195));
    jdff dff_B_6qhEYN629_2(.din(n27195), .dout(n27198));
    jdff dff_B_8L7B1R8z3_2(.din(n27198), .dout(n27201));
    jdff dff_B_MvYxJbrD3_2(.din(n27201), .dout(n27204));
    jdff dff_B_0hN6HVNw3_2(.din(n27204), .dout(n27207));
    jdff dff_B_MjmfVJrZ1_2(.din(n27207), .dout(n27210));
    jdff dff_B_ybvTQLDj6_2(.din(n27210), .dout(n27213));
    jdff dff_B_NBui3msE9_2(.din(n27213), .dout(n27216));
    jdff dff_B_b7o55a3V5_2(.din(n27216), .dout(n27219));
    jdff dff_B_bYHH4Yfc8_2(.din(n27219), .dout(n27222));
    jdff dff_B_N9AL9DrK6_2(.din(n27222), .dout(n27225));
    jdff dff_B_g4sqGszj0_2(.din(n27225), .dout(n27228));
    jdff dff_B_YuhbQnDV1_2(.din(n5987), .dout(n27231));
    jdff dff_B_QaZA6LOD3_1(.din(n5979), .dout(n27234));
    jdff dff_B_RzWB5iSg2_2(.din(n5757), .dout(n27237));
    jdff dff_B_NdfeGn7z7_2(.din(n27237), .dout(n27240));
    jdff dff_B_I4ubmTIl0_2(.din(n27240), .dout(n27243));
    jdff dff_B_iWz0g9oD4_2(.din(n27243), .dout(n27246));
    jdff dff_B_CjGinJYp1_2(.din(n27246), .dout(n27249));
    jdff dff_B_BLnkTZ9F0_2(.din(n27249), .dout(n27252));
    jdff dff_B_V1dW6LMn0_2(.din(n27252), .dout(n27255));
    jdff dff_B_UlYrC57j3_2(.din(n27255), .dout(n27258));
    jdff dff_B_oKIsmv7I1_2(.din(n27258), .dout(n27261));
    jdff dff_B_s0T3wLst3_2(.din(n27261), .dout(n27264));
    jdff dff_B_DsevGJRv5_2(.din(n27264), .dout(n27267));
    jdff dff_B_3HG2h4uj7_2(.din(n27267), .dout(n27270));
    jdff dff_B_bl2F6YaM6_2(.din(n27270), .dout(n27273));
    jdff dff_B_jW8y2dBd1_2(.din(n27273), .dout(n27276));
    jdff dff_B_XHAP7rNe0_2(.din(n27276), .dout(n27279));
    jdff dff_B_j5ZlGhP52_2(.din(n27279), .dout(n27282));
    jdff dff_B_7Nc3XTFA8_2(.din(n27282), .dout(n27285));
    jdff dff_B_5TvAHopH4_2(.din(n27285), .dout(n27288));
    jdff dff_B_uJ0AlV0R0_2(.din(n27288), .dout(n27291));
    jdff dff_B_c1mHGTGw3_2(.din(n27291), .dout(n27294));
    jdff dff_B_P2x1g1VB8_2(.din(n27294), .dout(n27297));
    jdff dff_B_T6aPQNht1_2(.din(n27297), .dout(n27300));
    jdff dff_B_70n6rwZV7_2(.din(n27300), .dout(n27303));
    jdff dff_B_YNZMNGWQ8_2(.din(n27303), .dout(n27306));
    jdff dff_B_dDnYqVIC0_2(.din(n27306), .dout(n27309));
    jdff dff_B_LCP5en5G1_2(.din(n27309), .dout(n27312));
    jdff dff_B_UDmQUMAb0_2(.din(n27312), .dout(n27315));
    jdff dff_B_1Rf4n2bq3_2(.din(n27315), .dout(n27318));
    jdff dff_B_KQuy6tPL7_2(.din(n27318), .dout(n27321));
    jdff dff_B_2SX8haRQ9_2(.din(n27321), .dout(n27324));
    jdff dff_B_kZx66CwO6_2(.din(n27324), .dout(n27327));
    jdff dff_B_5ix9SUyF4_2(.din(n27327), .dout(n27330));
    jdff dff_B_g8O4kjua5_2(.din(n27330), .dout(n27333));
    jdff dff_B_8XvW1uyN8_2(.din(n27333), .dout(n27336));
    jdff dff_B_mKfxyogV8_2(.din(n5769), .dout(n27339));
    jdff dff_B_iQ0mUJQH6_1(.din(n5761), .dout(n27342));
    jdff dff_B_dQdqVN723_2(.din(n5512), .dout(n27345));
    jdff dff_B_NTPd2rSh2_2(.din(n27345), .dout(n27348));
    jdff dff_B_zqV67sBM5_2(.din(n27348), .dout(n27351));
    jdff dff_B_n099u9Pv0_2(.din(n27351), .dout(n27354));
    jdff dff_B_6Sab7Gvb9_2(.din(n27354), .dout(n27357));
    jdff dff_B_gLeGkFh78_2(.din(n27357), .dout(n27360));
    jdff dff_B_ddkL6cTG5_2(.din(n27360), .dout(n27363));
    jdff dff_B_XCUWzEbc6_2(.din(n27363), .dout(n27366));
    jdff dff_B_UrPrCatm2_2(.din(n27366), .dout(n27369));
    jdff dff_B_eu3o8Ibq0_2(.din(n27369), .dout(n27372));
    jdff dff_B_hzY9z3lZ4_2(.din(n27372), .dout(n27375));
    jdff dff_B_n2NpeEVV3_2(.din(n27375), .dout(n27378));
    jdff dff_B_mNy4Cxjq4_2(.din(n27378), .dout(n27381));
    jdff dff_B_xZQFpAmx4_2(.din(n27381), .dout(n27384));
    jdff dff_B_HsqbjUEV3_2(.din(n27384), .dout(n27387));
    jdff dff_B_wCzqPmun3_2(.din(n27387), .dout(n27390));
    jdff dff_B_u0zIWOXM2_2(.din(n27390), .dout(n27393));
    jdff dff_B_UEzWtuxx1_2(.din(n27393), .dout(n27396));
    jdff dff_B_O71PxFAS5_2(.din(n27396), .dout(n27399));
    jdff dff_B_wIaZn0DU1_2(.din(n27399), .dout(n27402));
    jdff dff_B_s7c5mmix7_2(.din(n27402), .dout(n27405));
    jdff dff_B_G4522sUc5_2(.din(n27405), .dout(n27408));
    jdff dff_B_9Q1p4yba0_2(.din(n27408), .dout(n27411));
    jdff dff_B_jhCC9DdC0_2(.din(n27411), .dout(n27414));
    jdff dff_B_c6yzg8PN3_2(.din(n27414), .dout(n27417));
    jdff dff_B_LCNauuFj0_2(.din(n27417), .dout(n27420));
    jdff dff_B_xLJgt0sl3_2(.din(n27420), .dout(n27423));
    jdff dff_B_jx55aJCp5_2(.din(n27423), .dout(n27426));
    jdff dff_B_84X8Q3Iq5_2(.din(n27426), .dout(n27429));
    jdff dff_B_qrmTfwrb9_2(.din(n27429), .dout(n27432));
    jdff dff_B_KkbJhSEQ3_2(.din(n5524), .dout(n27435));
    jdff dff_B_ho8lWHFt5_1(.din(n5516), .dout(n27438));
    jdff dff_B_S58oYmMa0_2(.din(n5240), .dout(n27441));
    jdff dff_B_IKGTS3zP1_2(.din(n27441), .dout(n27444));
    jdff dff_B_DUCn5t4Q7_2(.din(n27444), .dout(n27447));
    jdff dff_B_1MiFA5151_2(.din(n27447), .dout(n27450));
    jdff dff_B_C6Zyxbbl3_2(.din(n27450), .dout(n27453));
    jdff dff_B_ZGPI2EY02_2(.din(n27453), .dout(n27456));
    jdff dff_B_DkH4Sp0K4_2(.din(n27456), .dout(n27459));
    jdff dff_B_BciaIpX67_2(.din(n27459), .dout(n27462));
    jdff dff_B_hPADyZlN8_2(.din(n27462), .dout(n27465));
    jdff dff_B_uN7n0fjF1_2(.din(n27465), .dout(n27468));
    jdff dff_B_LEEUnOa70_2(.din(n27468), .dout(n27471));
    jdff dff_B_KhVTjsAB2_2(.din(n27471), .dout(n27474));
    jdff dff_B_GcII21Rg3_2(.din(n27474), .dout(n27477));
    jdff dff_B_U71n6pbz7_2(.din(n27477), .dout(n27480));
    jdff dff_B_XulHHwSR3_2(.din(n27480), .dout(n27483));
    jdff dff_B_KpREJOeS1_2(.din(n27483), .dout(n27486));
    jdff dff_B_jTA3M3jC7_2(.din(n27486), .dout(n27489));
    jdff dff_B_vyF548bN1_2(.din(n27489), .dout(n27492));
    jdff dff_B_OMv3a6iv1_2(.din(n27492), .dout(n27495));
    jdff dff_B_Z8u58FAa3_2(.din(n27495), .dout(n27498));
    jdff dff_B_5p5T4rIz2_2(.din(n27498), .dout(n27501));
    jdff dff_B_vtpdGxVm4_2(.din(n27501), .dout(n27504));
    jdff dff_B_KMI7p34y5_2(.din(n27504), .dout(n27507));
    jdff dff_B_QH1yS4HV2_2(.din(n27507), .dout(n27510));
    jdff dff_B_AHxknJIR7_2(.din(n27510), .dout(n27513));
    jdff dff_B_1BL8Ahqj1_2(.din(n27513), .dout(n27516));
    jdff dff_B_XCPKuwD08_1(.din(n5244), .dout(n27519));
    jdff dff_B_8fWD4FDZ5_2(.din(n4941), .dout(n27522));
    jdff dff_B_0bmhFsBP2_2(.din(n27522), .dout(n27525));
    jdff dff_B_L8tmRKeS6_2(.din(n27525), .dout(n27528));
    jdff dff_B_Zq0PgvtI0_2(.din(n27528), .dout(n27531));
    jdff dff_B_bh9e0hKE9_2(.din(n27531), .dout(n27534));
    jdff dff_B_gvCo8ja90_2(.din(n27534), .dout(n27537));
    jdff dff_B_vPabyj2N4_2(.din(n27537), .dout(n27540));
    jdff dff_B_C4KObj3N2_2(.din(n27540), .dout(n27543));
    jdff dff_B_6tM6Bikm2_2(.din(n27543), .dout(n27546));
    jdff dff_B_Fxh8FrRE8_2(.din(n27546), .dout(n27549));
    jdff dff_B_1eMWfmE62_2(.din(n27549), .dout(n27552));
    jdff dff_B_iLlOrbvU8_2(.din(n27552), .dout(n27555));
    jdff dff_B_LoGDqp0X6_2(.din(n27555), .dout(n27558));
    jdff dff_B_24k2RjLd8_2(.din(n27558), .dout(n27561));
    jdff dff_B_2fR7Wl904_2(.din(n27561), .dout(n27564));
    jdff dff_B_k1RGTAP00_2(.din(n27564), .dout(n27567));
    jdff dff_B_ccpovmWP2_2(.din(n27567), .dout(n27570));
    jdff dff_B_fyHA7Bdf4_2(.din(n27570), .dout(n27573));
    jdff dff_B_fu7MWsCY7_2(.din(n27573), .dout(n27576));
    jdff dff_B_i43YjZIH4_2(.din(n27576), .dout(n27579));
    jdff dff_B_Wv5N0oYO3_2(.din(n27579), .dout(n27582));
    jdff dff_B_cb5H1mkX6_2(.din(n27582), .dout(n27585));
    jdff dff_B_QDSLTbY30_2(.din(n27585), .dout(n27588));
    jdff dff_B_HCQgwVJi0_2(.din(n5011), .dout(n27591));
    jdff dff_B_JqAWgDf77_1(.din(n4945), .dout(n27594));
    jdff dff_B_cjg5O9F09_2(.din(n4615), .dout(n27597));
    jdff dff_B_eD6PzqY11_2(.din(n27597), .dout(n27600));
    jdff dff_B_0mU4iFnm1_2(.din(n27600), .dout(n27603));
    jdff dff_B_sXGLcywk4_2(.din(n27603), .dout(n27606));
    jdff dff_B_83KL4U2s0_2(.din(n27606), .dout(n27609));
    jdff dff_B_qnPe1rC34_2(.din(n27609), .dout(n27612));
    jdff dff_B_FjH128Yc7_2(.din(n27612), .dout(n27615));
    jdff dff_B_3MVQSV9i7_2(.din(n27615), .dout(n27618));
    jdff dff_B_7RFmhv6M5_2(.din(n27618), .dout(n27621));
    jdff dff_B_9bqj45Az9_2(.din(n27621), .dout(n27624));
    jdff dff_B_jcI5yAf75_2(.din(n27624), .dout(n27627));
    jdff dff_B_e3mmbSYq6_2(.din(n27627), .dout(n27630));
    jdff dff_B_jtjhHmXu3_2(.din(n27630), .dout(n27633));
    jdff dff_B_BQSGshNK2_2(.din(n27633), .dout(n27636));
    jdff dff_B_hiE1BAur6_2(.din(n27636), .dout(n27639));
    jdff dff_B_PBJpxvx89_2(.din(n27639), .dout(n27642));
    jdff dff_B_2sugV3bU7_2(.din(n27642), .dout(n27645));
    jdff dff_B_xIxdlzct2_2(.din(n27645), .dout(n27648));
    jdff dff_B_swwuuHOT8_2(.din(n27648), .dout(n27651));
    jdff dff_B_f1fCDRhk4_2(.din(n27651), .dout(n27654));
    jdff dff_B_Xe6He2ej0_2(.din(n4685), .dout(n27657));
    jdff dff_B_bVIrtuqp5_1(.din(n4619), .dout(n27660));
    jdff dff_B_6m1xM35V8_2(.din(n4265), .dout(n27663));
    jdff dff_B_Cg7d4s2f6_2(.din(n27663), .dout(n27666));
    jdff dff_B_WXTTm8Gk6_2(.din(n27666), .dout(n27669));
    jdff dff_B_QmjzsAcW2_2(.din(n27669), .dout(n27672));
    jdff dff_B_LtJR30tu6_2(.din(n27672), .dout(n27675));
    jdff dff_B_Nsc63dWk3_2(.din(n27675), .dout(n27678));
    jdff dff_B_DompU1Mn5_2(.din(n27678), .dout(n27681));
    jdff dff_B_qNgr9wnv7_2(.din(n27681), .dout(n27684));
    jdff dff_B_7qLpwFRF7_2(.din(n27684), .dout(n27687));
    jdff dff_B_FMwohWg13_2(.din(n27687), .dout(n27690));
    jdff dff_B_sm3ZAiPd7_2(.din(n27690), .dout(n27693));
    jdff dff_B_PGvRhzpx8_2(.din(n27693), .dout(n27696));
    jdff dff_B_Ff6loTOH1_2(.din(n27696), .dout(n27699));
    jdff dff_B_JGntCBvc0_2(.din(n27699), .dout(n27702));
    jdff dff_B_tgJVvPhR1_2(.din(n27702), .dout(n27705));
    jdff dff_B_fYzdwXKl8_2(.din(n27705), .dout(n27708));
    jdff dff_B_n2dKzKE83_2(.din(n27708), .dout(n27711));
    jdff dff_B_I90VvDvk6_2(.din(n4335), .dout(n27714));
    jdff dff_B_RyEVqxOx9_1(.din(n4269), .dout(n27717));
    jdff dff_B_5y5m7if40_2(.din(n3889), .dout(n27720));
    jdff dff_B_C7NOqQmo0_2(.din(n27720), .dout(n27723));
    jdff dff_B_nOiyILY67_2(.din(n27723), .dout(n27726));
    jdff dff_B_Nr3nNIHK5_2(.din(n27726), .dout(n27729));
    jdff dff_B_Sldwm07Z4_2(.din(n27729), .dout(n27732));
    jdff dff_B_696ONaBT7_2(.din(n27732), .dout(n27735));
    jdff dff_B_5WJOaiIf6_2(.din(n27735), .dout(n27738));
    jdff dff_B_owGEMTNz7_2(.din(n27738), .dout(n27741));
    jdff dff_B_MTvfbLHM2_2(.din(n27741), .dout(n27744));
    jdff dff_B_QejiHL5P1_2(.din(n27744), .dout(n27747));
    jdff dff_B_blyeLdE39_2(.din(n27747), .dout(n27750));
    jdff dff_B_ftThUZDC8_2(.din(n27750), .dout(n27753));
    jdff dff_B_1OYb2m226_2(.din(n27753), .dout(n27756));
    jdff dff_B_Ci9wtgQJ5_2(.din(n27756), .dout(n27759));
    jdff dff_B_smVEtmv42_2(.din(n3955), .dout(n27762));
    jdff dff_B_zrwX1Wfj8_1(.din(n3893), .dout(n27765));
    jdff dff_B_Vyrvde2k7_2(.din(n3509), .dout(n27768));
    jdff dff_B_7dHNVaiX3_2(.din(n27768), .dout(n27771));
    jdff dff_B_Z07SO9pK4_2(.din(n27771), .dout(n27774));
    jdff dff_B_CU3VdFFs7_2(.din(n27774), .dout(n27777));
    jdff dff_B_1pRFknuG1_2(.din(n27777), .dout(n27780));
    jdff dff_B_pDyPHFbo8_2(.din(n27780), .dout(n27783));
    jdff dff_B_hW581FkD7_2(.din(n27783), .dout(n27786));
    jdff dff_B_ax2HaJUt4_2(.din(n27786), .dout(n27789));
    jdff dff_B_XyB4ET0e1_2(.din(n27789), .dout(n27792));
    jdff dff_B_7FkRkUes7_2(.din(n27792), .dout(n27795));
    jdff dff_B_imKGIIwC7_2(.din(n27795), .dout(n27798));
    jdff dff_B_NGWTcjpH5_2(.din(n3572), .dout(n27801));
    jdff dff_B_4oC1homs9_1(.din(n3513), .dout(n27804));
    jdff dff_B_aWKR5lhH0_2(.din(n3118), .dout(n27807));
    jdff dff_B_AciXEQ3X1_2(.din(n27807), .dout(n27810));
    jdff dff_B_RC2f9G3l3_2(.din(n27810), .dout(n27813));
    jdff dff_B_EuFkQLMU9_2(.din(n27813), .dout(n27816));
    jdff dff_B_d7qrxhmy8_2(.din(n27816), .dout(n27819));
    jdff dff_B_lKZInh7R6_2(.din(n27819), .dout(n27822));
    jdff dff_B_lvn5e4YR2_2(.din(n27822), .dout(n27825));
    jdff dff_B_wSpih1Qt8_2(.din(n27825), .dout(n27828));
    jdff dff_B_9x4o2KCf7_2(.din(n3167), .dout(n27831));
    jdff dff_B_OzCmzcbf7_2(.din(n27831), .dout(n27834));
    jdff dff_B_aL4m3DRC6_2(.din(n27834), .dout(n27837));
    jdff dff_B_9hdXcse39_1(.din(n3122), .dout(n27840));
    jdff dff_B_IPyqcC861_1(.din(n27840), .dout(n27843));
    jdff dff_B_U4bDjFzh5_2(.din(n2749), .dout(n27846));
    jdff dff_B_LYiWz5wH8_2(.din(n27846), .dout(n27849));
    jdff dff_B_BUBibZu93_2(.din(n27849), .dout(n27852));
    jdff dff_B_A0THsbh72_0(.din(n2768), .dout(n27855));
    jdff dff_A_sRUxz9k22_0(.din(n27860), .dout(n27857));
    jdff dff_A_sb8ifWuf6_0(.din(n2387), .dout(n27860));
    jdff dff_A_v5IQem1f2_1(.din(n27866), .dout(n27863));
    jdff dff_A_YptSCDAG8_1(.din(n2387), .dout(n27866));
    jdff dff_B_3khtPMZW2_1(.din(n6741), .dout(n27870));
    jdff dff_B_9DLV4WV10_1(.din(n6691), .dout(n27873));
    jdff dff_B_faZ3ZuPl5_1(.din(n27873), .dout(n27876));
    jdff dff_B_MfPpxzJJ9_2(.din(n6687), .dout(n27879));
    jdff dff_B_wqld1sS99_2(.din(n27879), .dout(n27882));
    jdff dff_B_TFMUueFe3_2(.din(n27882), .dout(n27885));
    jdff dff_B_meT1L5XU9_2(.din(n27885), .dout(n27888));
    jdff dff_B_eIGPAlFf5_2(.din(n27888), .dout(n27891));
    jdff dff_B_GYFatfmk0_2(.din(n27891), .dout(n27894));
    jdff dff_B_UFZSArsj2_2(.din(n27894), .dout(n27897));
    jdff dff_B_brlA7cSV0_2(.din(n27897), .dout(n27900));
    jdff dff_B_m91rymN61_2(.din(n27900), .dout(n27903));
    jdff dff_B_bZPLzYsL4_2(.din(n27903), .dout(n27906));
    jdff dff_B_g3fF2vhK7_2(.din(n27906), .dout(n27909));
    jdff dff_B_NSDCk7Dd7_2(.din(n27909), .dout(n27912));
    jdff dff_B_GX258PLG1_2(.din(n27912), .dout(n27915));
    jdff dff_B_GlgEY3dY5_2(.din(n27915), .dout(n27918));
    jdff dff_B_w9khd0Be5_2(.din(n27918), .dout(n27921));
    jdff dff_B_2lfrzC9f1_2(.din(n27921), .dout(n27924));
    jdff dff_B_9PLjGxQl9_2(.din(n27924), .dout(n27927));
    jdff dff_B_LiCwUIuV8_2(.din(n27927), .dout(n27930));
    jdff dff_B_hYnWIWjr6_2(.din(n27930), .dout(n27933));
    jdff dff_B_Xmzl4cMp4_2(.din(n27933), .dout(n27936));
    jdff dff_B_NoZ2XuEd6_2(.din(n27936), .dout(n27939));
    jdff dff_B_uHW3695z4_2(.din(n27939), .dout(n27942));
    jdff dff_B_YYFN2Zed4_2(.din(n27942), .dout(n27945));
    jdff dff_B_yYEalvjV5_2(.din(n27945), .dout(n27948));
    jdff dff_B_NvM6fDmN8_2(.din(n27948), .dout(n27951));
    jdff dff_B_BuhkKyiz1_2(.din(n27951), .dout(n27954));
    jdff dff_B_USWE1dzW0_2(.din(n27954), .dout(n27957));
    jdff dff_B_HpAjlrzA1_2(.din(n27957), .dout(n27960));
    jdff dff_B_vYBqpBVu4_2(.din(n27960), .dout(n27963));
    jdff dff_B_UJbJAONb9_2(.din(n27963), .dout(n27966));
    jdff dff_B_PHo3CXyP2_2(.din(n27966), .dout(n27969));
    jdff dff_B_mcM7JGJ51_2(.din(n27969), .dout(n27972));
    jdff dff_B_fdrUX4wB3_2(.din(n27972), .dout(n27975));
    jdff dff_B_s1gwsI996_2(.din(n27975), .dout(n27978));
    jdff dff_B_FQBwSGez0_2(.din(n27978), .dout(n27981));
    jdff dff_B_sHeUz6nC6_2(.din(n27981), .dout(n27984));
    jdff dff_B_cOsl4YVb1_2(.din(n27984), .dout(n27987));
    jdff dff_B_fTwFTflT5_2(.din(n27987), .dout(n27990));
    jdff dff_B_H5yL1yby8_2(.din(n27990), .dout(n27993));
    jdff dff_B_a8SEDwBz6_2(.din(n27993), .dout(n27996));
    jdff dff_B_TwxTjr6m7_2(.din(n27996), .dout(n27999));
    jdff dff_B_Yxnipmd05_2(.din(n27999), .dout(n28002));
    jdff dff_B_0gvTZBI68_2(.din(n28002), .dout(n28005));
    jdff dff_B_PB7KWXqT8_2(.din(n28005), .dout(n28008));
    jdff dff_B_Lko5MVvg3_2(.din(n28008), .dout(n28011));
    jdff dff_B_HSCpKC7y0_2(.din(n28011), .dout(n28014));
    jdff dff_B_OrMGwLI38_2(.din(n28014), .dout(n28017));
    jdff dff_B_uTO94k8z0_2(.din(n28017), .dout(n28020));
    jdff dff_B_Jj1COXCJ9_2(.din(n28020), .dout(n28023));
    jdff dff_B_Ar2B9dB93_2(.din(n28023), .dout(n28026));
    jdff dff_B_fkpKJ1nu2_2(.din(n28026), .dout(n28029));
    jdff dff_B_77zVpOrb5_2(.din(n28029), .dout(n28032));
    jdff dff_B_6aixUHpW2_2(.din(n28032), .dout(n28035));
    jdff dff_B_IGeMV9ib9_2(.din(n6683), .dout(n28038));
    jdff dff_B_1hXPoMWS8_2(.din(n28038), .dout(n28041));
    jdff dff_B_hTm9IOLP4_2(.din(n28041), .dout(n28044));
    jdff dff_B_lUSdTHp65_2(.din(n28044), .dout(n28047));
    jdff dff_B_nkhFoypa0_2(.din(n28047), .dout(n28050));
    jdff dff_B_hFKUTLDw7_2(.din(n28050), .dout(n28053));
    jdff dff_B_OlSnPDNG8_2(.din(n28053), .dout(n28056));
    jdff dff_B_MJVdG18b0_2(.din(n28056), .dout(n28059));
    jdff dff_B_uHrKPwcu2_2(.din(n28059), .dout(n28062));
    jdff dff_B_ARfFCk4c8_2(.din(n28062), .dout(n28065));
    jdff dff_B_0uOtnRUs4_2(.din(n28065), .dout(n28068));
    jdff dff_B_GgziSO107_2(.din(n28068), .dout(n28071));
    jdff dff_B_f2H1AQPX8_2(.din(n28071), .dout(n28074));
    jdff dff_B_Wbda1GtI8_2(.din(n28074), .dout(n28077));
    jdff dff_B_YzgAQTqb6_2(.din(n28077), .dout(n28080));
    jdff dff_B_5a1WIX7l3_2(.din(n28080), .dout(n28083));
    jdff dff_B_DGGBXSaQ6_2(.din(n28083), .dout(n28086));
    jdff dff_B_zKSRgERY3_2(.din(n28086), .dout(n28089));
    jdff dff_B_ZH41LcwF6_2(.din(n28089), .dout(n28092));
    jdff dff_B_JxGqPK4N2_2(.din(n28092), .dout(n28095));
    jdff dff_B_vdOInZ5o7_2(.din(n28095), .dout(n28098));
    jdff dff_B_wq5U4Wf54_2(.din(n28098), .dout(n28101));
    jdff dff_B_8DNgGRHO6_2(.din(n28101), .dout(n28104));
    jdff dff_B_hBdRicXW5_2(.din(n28104), .dout(n28107));
    jdff dff_B_y05gS8lc0_2(.din(n28107), .dout(n28110));
    jdff dff_B_CKs8n0Ga0_2(.din(n28110), .dout(n28113));
    jdff dff_B_QSqeWaxf5_2(.din(n28113), .dout(n28116));
    jdff dff_B_vkXyBreC2_2(.din(n28116), .dout(n28119));
    jdff dff_B_RH3bIGlB7_2(.din(n28119), .dout(n28122));
    jdff dff_B_nkG0x9KF5_2(.din(n28122), .dout(n28125));
    jdff dff_B_99JDZfRv1_2(.din(n28125), .dout(n28128));
    jdff dff_B_gC5WPp5f2_2(.din(n28128), .dout(n28131));
    jdff dff_B_9gwnppzM2_2(.din(n28131), .dout(n28134));
    jdff dff_B_UGPfeOys5_2(.din(n28134), .dout(n28137));
    jdff dff_B_1p3qAfnr3_2(.din(n28137), .dout(n28140));
    jdff dff_B_nzqDpM5g9_2(.din(n28140), .dout(n28143));
    jdff dff_B_j2gRuAmv6_2(.din(n28143), .dout(n28146));
    jdff dff_B_qjyyVmx96_2(.din(n28146), .dout(n28149));
    jdff dff_B_MOd2wavx1_2(.din(n28149), .dout(n28152));
    jdff dff_B_edEKACBM9_2(.din(n28152), .dout(n28155));
    jdff dff_B_iMCb9WWC1_2(.din(n28155), .dout(n28158));
    jdff dff_B_2EolgRcV6_2(.din(n28158), .dout(n28161));
    jdff dff_B_eQikfSyF9_2(.din(n28161), .dout(n28164));
    jdff dff_B_zZP6iBpU1_2(.din(n28164), .dout(n28167));
    jdff dff_B_sxPkbQoA5_2(.din(n28167), .dout(n28170));
    jdff dff_B_UVizJ9OA6_2(.din(n28170), .dout(n28173));
    jdff dff_B_Qmo4U34Y5_2(.din(n28173), .dout(n28176));
    jdff dff_B_PxKGak9c1_2(.din(n28176), .dout(n28179));
    jdff dff_B_bZvZbHM05_2(.din(n28179), .dout(n28182));
    jdff dff_B_BTIdkmGU8_2(.din(n28182), .dout(n28185));
    jdff dff_B_LjShF65B1_2(.din(n28185), .dout(n28188));
    jdff dff_B_Sx5j2Lhm8_2(.din(n28188), .dout(n28191));
    jdff dff_B_wGYfX4iD3_2(.din(n28191), .dout(n28194));
    jdff dff_B_77mgntCa2_2(.din(n28194), .dout(n28197));
    jdff dff_B_JTBAVYp00_2(.din(n28197), .dout(n28200));
    jdff dff_A_kIMEJZuV4_1(.din(n6679), .dout(n28202));
    jdff dff_B_kLCCYxg90_1(.din(n6671), .dout(n28206));
    jdff dff_B_6WvChU4n7_2(.din(n6587), .dout(n28209));
    jdff dff_B_VeE8k1Js9_2(.din(n28209), .dout(n28212));
    jdff dff_B_b0ffJJZ37_2(.din(n28212), .dout(n28215));
    jdff dff_B_qUAGjAFZ7_2(.din(n28215), .dout(n28218));
    jdff dff_B_HbUZ7giP6_2(.din(n28218), .dout(n28221));
    jdff dff_B_225T9Tfg2_2(.din(n28221), .dout(n28224));
    jdff dff_B_2Ebq5G2f8_2(.din(n28224), .dout(n28227));
    jdff dff_B_qLonYJt09_2(.din(n28227), .dout(n28230));
    jdff dff_B_rW4he9le3_2(.din(n28230), .dout(n28233));
    jdff dff_B_WltqSuis1_2(.din(n28233), .dout(n28236));
    jdff dff_B_WH1ZPVG68_2(.din(n28236), .dout(n28239));
    jdff dff_B_JxdmMQdi8_2(.din(n28239), .dout(n28242));
    jdff dff_B_YtQ5t4BL2_2(.din(n28242), .dout(n28245));
    jdff dff_B_9cMtjPah8_2(.din(n28245), .dout(n28248));
    jdff dff_B_T714fXWc2_2(.din(n28248), .dout(n28251));
    jdff dff_B_5ehTGXKN0_2(.din(n28251), .dout(n28254));
    jdff dff_B_U3HENvgj9_2(.din(n28254), .dout(n28257));
    jdff dff_B_sale1tLe9_2(.din(n28257), .dout(n28260));
    jdff dff_B_uG6YmGoK2_2(.din(n28260), .dout(n28263));
    jdff dff_B_ucI4AD7R8_2(.din(n28263), .dout(n28266));
    jdff dff_B_2AtVjVru3_2(.din(n28266), .dout(n28269));
    jdff dff_B_wi2x7uf67_2(.din(n28269), .dout(n28272));
    jdff dff_B_oWb3rbPn0_2(.din(n28272), .dout(n28275));
    jdff dff_B_GAs5Apbm0_2(.din(n28275), .dout(n28278));
    jdff dff_B_89P7xuT70_2(.din(n28278), .dout(n28281));
    jdff dff_B_UzxMRUuo1_2(.din(n28281), .dout(n28284));
    jdff dff_B_UtvfWYMs8_2(.din(n28284), .dout(n28287));
    jdff dff_B_vTVOUeVN0_2(.din(n28287), .dout(n28290));
    jdff dff_B_tnw1i2EO3_2(.din(n28290), .dout(n28293));
    jdff dff_B_utnlB5gF5_2(.din(n28293), .dout(n28296));
    jdff dff_B_0jtgF9Pa2_2(.din(n28296), .dout(n28299));
    jdff dff_B_ToWwYuCP9_2(.din(n28299), .dout(n28302));
    jdff dff_B_3ElCogYp8_2(.din(n28302), .dout(n28305));
    jdff dff_B_da2by9p20_2(.din(n28305), .dout(n28308));
    jdff dff_B_XiqeBoTE8_2(.din(n28308), .dout(n28311));
    jdff dff_B_7PW0mHnc6_2(.din(n28311), .dout(n28314));
    jdff dff_B_LvrPfIdk7_2(.din(n28314), .dout(n28317));
    jdff dff_B_DFZ8lVSh3_2(.din(n28317), .dout(n28320));
    jdff dff_B_pXOmb06k6_2(.din(n28320), .dout(n28323));
    jdff dff_B_FrGaBkqP7_2(.din(n28323), .dout(n28326));
    jdff dff_B_DRKSCwm95_2(.din(n28326), .dout(n28329));
    jdff dff_B_CfL2HHFE9_2(.din(n28329), .dout(n28332));
    jdff dff_B_R1wbpUy81_2(.din(n28332), .dout(n28335));
    jdff dff_B_u2A0zG2l8_2(.din(n28335), .dout(n28338));
    jdff dff_B_bGYF4gsT3_2(.din(n28338), .dout(n28341));
    jdff dff_B_5DYZp9407_2(.din(n28341), .dout(n28344));
    jdff dff_B_n49NGnNO7_2(.din(n28344), .dout(n28347));
    jdff dff_B_0p1ewIGR8_2(.din(n28347), .dout(n28350));
    jdff dff_B_pee5vlDs6_2(.din(n28350), .dout(n28353));
    jdff dff_B_Nu1GZGt17_2(.din(n28353), .dout(n28356));
    jdff dff_B_04UzHpm74_2(.din(n28356), .dout(n28359));
    jdff dff_B_vc5rPiNp8_2(.din(n28359), .dout(n28362));
    jdff dff_B_IIrK9S8e4_1(.din(n6611), .dout(n28365));
    jdff dff_B_KInWw2Ze8_1(.din(n28365), .dout(n28368));
    jdff dff_B_NvrZTT2W4_2(.din(n6607), .dout(n28371));
    jdff dff_B_De0raXHb8_2(.din(n28371), .dout(n28374));
    jdff dff_B_8ufEoUho1_2(.din(n28374), .dout(n28377));
    jdff dff_B_WfiKk9ED1_2(.din(n28377), .dout(n28380));
    jdff dff_B_RR8CyNt29_2(.din(n28380), .dout(n28383));
    jdff dff_B_fwbLCIO69_2(.din(n28383), .dout(n28386));
    jdff dff_B_bIZv65pX6_2(.din(n28386), .dout(n28389));
    jdff dff_B_WlTNzLHA3_2(.din(n28389), .dout(n28392));
    jdff dff_B_bZc4q3YB1_2(.din(n28392), .dout(n28395));
    jdff dff_B_IhhxcOd89_2(.din(n28395), .dout(n28398));
    jdff dff_B_bvdpctnm3_2(.din(n28398), .dout(n28401));
    jdff dff_B_GHdlnLmj6_2(.din(n28401), .dout(n28404));
    jdff dff_B_mtzGz4AY3_2(.din(n28404), .dout(n28407));
    jdff dff_B_QGx8HGMa5_2(.din(n28407), .dout(n28410));
    jdff dff_B_L91D3la25_2(.din(n28410), .dout(n28413));
    jdff dff_B_CZ8Y5NwY2_2(.din(n28413), .dout(n28416));
    jdff dff_B_tpEbFM308_2(.din(n28416), .dout(n28419));
    jdff dff_B_9NpQc4t86_2(.din(n28419), .dout(n28422));
    jdff dff_B_YCFMKMzF9_2(.din(n28422), .dout(n28425));
    jdff dff_B_B3EHuTda0_2(.din(n28425), .dout(n28428));
    jdff dff_B_JhLcc2yb1_2(.din(n28428), .dout(n28431));
    jdff dff_B_mquBrRvZ8_2(.din(n28431), .dout(n28434));
    jdff dff_B_QaQo3S3Q2_2(.din(n28434), .dout(n28437));
    jdff dff_B_3VG0ynRn9_2(.din(n28437), .dout(n28440));
    jdff dff_B_t2D9BH491_2(.din(n28440), .dout(n28443));
    jdff dff_B_wZwMO1n63_2(.din(n28443), .dout(n28446));
    jdff dff_B_CSEUDD1e1_2(.din(n28446), .dout(n28449));
    jdff dff_B_saawBkeW2_2(.din(n28449), .dout(n28452));
    jdff dff_B_UemBGa1j1_2(.din(n28452), .dout(n28455));
    jdff dff_B_98nErRHJ8_2(.din(n28455), .dout(n28458));
    jdff dff_B_11LC3EgX4_2(.din(n28458), .dout(n28461));
    jdff dff_B_MjhrhxhZ0_2(.din(n28461), .dout(n28464));
    jdff dff_B_EZjFtKMT9_2(.din(n28464), .dout(n28467));
    jdff dff_B_jdkNWGqi4_2(.din(n28467), .dout(n28470));
    jdff dff_B_BQuO9eMB8_2(.din(n28470), .dout(n28473));
    jdff dff_B_qwHNU55a6_2(.din(n28473), .dout(n28476));
    jdff dff_B_iciNOIY51_2(.din(n28476), .dout(n28479));
    jdff dff_B_S48muyIX0_2(.din(n28479), .dout(n28482));
    jdff dff_B_K7cPHnl28_2(.din(n28482), .dout(n28485));
    jdff dff_B_f6nEfctv1_2(.din(n28485), .dout(n28488));
    jdff dff_B_IDk7U9bE4_2(.din(n28488), .dout(n28491));
    jdff dff_B_e6LfYu1o8_2(.din(n28491), .dout(n28494));
    jdff dff_B_NxnBI4752_2(.din(n28494), .dout(n28497));
    jdff dff_B_ExZacyRm6_2(.din(n28497), .dout(n28500));
    jdff dff_B_x5WR6gah7_2(.din(n28500), .dout(n28503));
    jdff dff_B_PaHaOLhD0_2(.din(n28503), .dout(n28506));
    jdff dff_B_0IALB7UA1_2(.din(n28506), .dout(n28509));
    jdff dff_B_NBVbAG3x8_2(.din(n28509), .dout(n28512));
    jdff dff_B_PIWEmWL32_2(.din(n28512), .dout(n28515));
    jdff dff_B_iImEmESC3_2(.din(n6603), .dout(n28518));
    jdff dff_B_ioW0lsdf2_2(.din(n28518), .dout(n28521));
    jdff dff_B_b8avPETQ4_2(.din(n28521), .dout(n28524));
    jdff dff_B_Gl93NYTU5_2(.din(n28524), .dout(n28527));
    jdff dff_B_Bv4Iw56G1_2(.din(n28527), .dout(n28530));
    jdff dff_B_NFDbYbnJ8_2(.din(n28530), .dout(n28533));
    jdff dff_B_ZHjLGGQq6_2(.din(n28533), .dout(n28536));
    jdff dff_B_vHlc8EKC4_2(.din(n28536), .dout(n28539));
    jdff dff_B_aN7Pusvh5_2(.din(n28539), .dout(n28542));
    jdff dff_B_ZJeEpx7f1_2(.din(n28542), .dout(n28545));
    jdff dff_B_hNeWZUh13_2(.din(n28545), .dout(n28548));
    jdff dff_B_Wv0oDHv37_2(.din(n28548), .dout(n28551));
    jdff dff_B_DY2AlFEn3_2(.din(n28551), .dout(n28554));
    jdff dff_B_AxjmYavE4_2(.din(n28554), .dout(n28557));
    jdff dff_B_OFJpi7aV4_2(.din(n28557), .dout(n28560));
    jdff dff_B_viHaDg3n8_2(.din(n28560), .dout(n28563));
    jdff dff_B_6KAxKkF52_2(.din(n28563), .dout(n28566));
    jdff dff_B_WvUy9Xgj7_2(.din(n28566), .dout(n28569));
    jdff dff_B_yjPwEgj65_2(.din(n28569), .dout(n28572));
    jdff dff_B_ceBBZEjj7_2(.din(n28572), .dout(n28575));
    jdff dff_B_xn6GsXHo8_2(.din(n28575), .dout(n28578));
    jdff dff_B_cGsJNLJ77_2(.din(n28578), .dout(n28581));
    jdff dff_B_dibxXs7f9_2(.din(n28581), .dout(n28584));
    jdff dff_B_BVXcjW8O3_2(.din(n28584), .dout(n28587));
    jdff dff_B_WHKlnkAW0_2(.din(n28587), .dout(n28590));
    jdff dff_B_JS1aW1tV3_2(.din(n28590), .dout(n28593));
    jdff dff_B_TOrT2Hal9_2(.din(n28593), .dout(n28596));
    jdff dff_B_edlU4s8A5_2(.din(n28596), .dout(n28599));
    jdff dff_B_N2b6l1Lb9_2(.din(n28599), .dout(n28602));
    jdff dff_B_1Q8PyZCg0_2(.din(n28602), .dout(n28605));
    jdff dff_B_Ryb6VMY08_2(.din(n28605), .dout(n28608));
    jdff dff_B_mL8KOsxt8_2(.din(n28608), .dout(n28611));
    jdff dff_B_Lqpb9cmN6_2(.din(n28611), .dout(n28614));
    jdff dff_B_we1dICRd6_2(.din(n28614), .dout(n28617));
    jdff dff_B_hlQ9slZK8_2(.din(n28617), .dout(n28620));
    jdff dff_B_OTAyjO1U2_2(.din(n28620), .dout(n28623));
    jdff dff_B_0t2RPjdF7_2(.din(n28623), .dout(n28626));
    jdff dff_B_VNckG46C8_2(.din(n28626), .dout(n28629));
    jdff dff_B_5AnD0mq88_2(.din(n28629), .dout(n28632));
    jdff dff_B_64R7jRtM0_2(.din(n28632), .dout(n28635));
    jdff dff_B_yZFX5zYs1_2(.din(n28635), .dout(n28638));
    jdff dff_B_rat0vrnm5_2(.din(n28638), .dout(n28641));
    jdff dff_B_cjrXDAJm2_2(.din(n28641), .dout(n28644));
    jdff dff_B_SX2lUEYc6_2(.din(n28644), .dout(n28647));
    jdff dff_B_fP9B9w7o9_2(.din(n28647), .dout(n28650));
    jdff dff_B_YdQuE3et0_2(.din(n28650), .dout(n28653));
    jdff dff_B_mDd0gWwf2_2(.din(n28653), .dout(n28656));
    jdff dff_B_hEINZUw46_2(.din(n28656), .dout(n28659));
    jdff dff_B_4S6Z5FUH4_2(.din(n28659), .dout(n28662));
    jdff dff_B_GAvzG52H4_2(.din(n28662), .dout(n28665));
    jdff dff_B_Lam9kCm25_2(.din(n28665), .dout(n28668));
    jdff dff_B_962kAxAN4_2(.din(n6599), .dout(n28671));
    jdff dff_B_w3zmnl6r0_1(.din(n6591), .dout(n28674));
    jdff dff_B_doL0YCC16_2(.din(n6480), .dout(n28677));
    jdff dff_B_PO80Hljs3_2(.din(n28677), .dout(n28680));
    jdff dff_B_tAoJnxxI7_2(.din(n28680), .dout(n28683));
    jdff dff_B_I9tNYdXt6_2(.din(n28683), .dout(n28686));
    jdff dff_B_xVYa1lsO8_2(.din(n28686), .dout(n28689));
    jdff dff_B_eGZKkaC31_2(.din(n28689), .dout(n28692));
    jdff dff_B_ag97yKCq3_2(.din(n28692), .dout(n28695));
    jdff dff_B_r5LZPEN60_2(.din(n28695), .dout(n28698));
    jdff dff_B_8GMA7ssn8_2(.din(n28698), .dout(n28701));
    jdff dff_B_HZSYmuGw2_2(.din(n28701), .dout(n28704));
    jdff dff_B_zpNYHYiv5_2(.din(n28704), .dout(n28707));
    jdff dff_B_GK7qFWiW3_2(.din(n28707), .dout(n28710));
    jdff dff_B_Tv4ccQm50_2(.din(n28710), .dout(n28713));
    jdff dff_B_lx9X790e1_2(.din(n28713), .dout(n28716));
    jdff dff_B_69GtdHYW0_2(.din(n28716), .dout(n28719));
    jdff dff_B_H8BvjoBO4_2(.din(n28719), .dout(n28722));
    jdff dff_B_U0rRh0O24_2(.din(n28722), .dout(n28725));
    jdff dff_B_Yft8nIWx2_2(.din(n28725), .dout(n28728));
    jdff dff_B_TULcQlcD6_2(.din(n28728), .dout(n28731));
    jdff dff_B_I6nnn3an5_2(.din(n28731), .dout(n28734));
    jdff dff_B_4UavkAXR7_2(.din(n28734), .dout(n28737));
    jdff dff_B_meDrfdmn5_2(.din(n28737), .dout(n28740));
    jdff dff_B_mZmAkMTK6_2(.din(n28740), .dout(n28743));
    jdff dff_B_DWy7vFSZ3_2(.din(n28743), .dout(n28746));
    jdff dff_B_u9cOpx384_2(.din(n28746), .dout(n28749));
    jdff dff_B_PrUIrbZJ0_2(.din(n28749), .dout(n28752));
    jdff dff_B_d0RyFGEL1_2(.din(n28752), .dout(n28755));
    jdff dff_B_w4FEVQiI4_2(.din(n28755), .dout(n28758));
    jdff dff_B_2V7g2ufw7_2(.din(n28758), .dout(n28761));
    jdff dff_B_qmcX0Slb6_2(.din(n28761), .dout(n28764));
    jdff dff_B_bi3efb5G8_2(.din(n28764), .dout(n28767));
    jdff dff_B_GGyeunjO4_2(.din(n28767), .dout(n28770));
    jdff dff_B_YYY4kqJg7_2(.din(n28770), .dout(n28773));
    jdff dff_B_c2rmAP3l6_2(.din(n28773), .dout(n28776));
    jdff dff_B_usUNnHza6_2(.din(n28776), .dout(n28779));
    jdff dff_B_P4zJadhL9_2(.din(n28779), .dout(n28782));
    jdff dff_B_cc8eC8nn5_2(.din(n28782), .dout(n28785));
    jdff dff_B_A6n8MjoI5_2(.din(n28785), .dout(n28788));
    jdff dff_B_meZHDjPW6_2(.din(n28788), .dout(n28791));
    jdff dff_B_hYYQqhYG9_2(.din(n28791), .dout(n28794));
    jdff dff_B_h5C3FUQk0_2(.din(n28794), .dout(n28797));
    jdff dff_B_hgpcHUij2_2(.din(n28797), .dout(n28800));
    jdff dff_B_waOVNIE37_2(.din(n28800), .dout(n28803));
    jdff dff_B_xnqK7Byh6_2(.din(n28803), .dout(n28806));
    jdff dff_B_p7B7sbbP7_2(.din(n28806), .dout(n28809));
    jdff dff_B_DcLUZTiI2_2(.din(n28809), .dout(n28812));
    jdff dff_B_G20dCVcg1_2(.din(n28812), .dout(n28815));
    jdff dff_B_Gqhqk55Q6_2(.din(n28815), .dout(n28818));
    jdff dff_B_KSBx9hgd8_1(.din(n6504), .dout(n28821));
    jdff dff_B_HuYfgTST5_1(.din(n28821), .dout(n28824));
    jdff dff_B_NRarIm481_2(.din(n6500), .dout(n28827));
    jdff dff_B_bNkLPfhj3_2(.din(n28827), .dout(n28830));
    jdff dff_B_HsTrgkDH7_2(.din(n28830), .dout(n28833));
    jdff dff_B_WJ1K3ROM2_2(.din(n28833), .dout(n28836));
    jdff dff_B_Sy2gkp6g9_2(.din(n28836), .dout(n28839));
    jdff dff_B_vQw3N8xP1_2(.din(n28839), .dout(n28842));
    jdff dff_B_hu3d0up95_2(.din(n28842), .dout(n28845));
    jdff dff_B_bwTsxGle8_2(.din(n28845), .dout(n28848));
    jdff dff_B_ZVHMzRyU3_2(.din(n28848), .dout(n28851));
    jdff dff_B_Aa3Ruav88_2(.din(n28851), .dout(n28854));
    jdff dff_B_1hOm2KMg3_2(.din(n28854), .dout(n28857));
    jdff dff_B_PstwEAOL5_2(.din(n28857), .dout(n28860));
    jdff dff_B_SBC3Jut87_2(.din(n28860), .dout(n28863));
    jdff dff_B_1x4BOWQm9_2(.din(n28863), .dout(n28866));
    jdff dff_B_FPk5bM1R3_2(.din(n28866), .dout(n28869));
    jdff dff_B_AZNJ5v4x4_2(.din(n28869), .dout(n28872));
    jdff dff_B_TCdxf6yk6_2(.din(n28872), .dout(n28875));
    jdff dff_B_13eA2AlI8_2(.din(n28875), .dout(n28878));
    jdff dff_B_BneWj0V76_2(.din(n28878), .dout(n28881));
    jdff dff_B_4GUV5hjH8_2(.din(n28881), .dout(n28884));
    jdff dff_B_GytnC5GA3_2(.din(n28884), .dout(n28887));
    jdff dff_B_vgouNKQR2_2(.din(n28887), .dout(n28890));
    jdff dff_B_ARMT9Ao40_2(.din(n28890), .dout(n28893));
    jdff dff_B_KyBIYozU9_2(.din(n28893), .dout(n28896));
    jdff dff_B_EnifDq9L0_2(.din(n28896), .dout(n28899));
    jdff dff_B_6uVhiURb5_2(.din(n28899), .dout(n28902));
    jdff dff_B_doFOBq3C3_2(.din(n28902), .dout(n28905));
    jdff dff_B_PiALsGyr0_2(.din(n28905), .dout(n28908));
    jdff dff_B_edLLhkFo3_2(.din(n28908), .dout(n28911));
    jdff dff_B_SCokj42K4_2(.din(n28911), .dout(n28914));
    jdff dff_B_1UDNjSQa5_2(.din(n28914), .dout(n28917));
    jdff dff_B_RcZVIRtI1_2(.din(n28917), .dout(n28920));
    jdff dff_B_l14ZrkSU1_2(.din(n28920), .dout(n28923));
    jdff dff_B_nsUfkMOK9_2(.din(n28923), .dout(n28926));
    jdff dff_B_iYkn4oJr6_2(.din(n28926), .dout(n28929));
    jdff dff_B_qY0Midl32_2(.din(n28929), .dout(n28932));
    jdff dff_B_YrCBHve83_2(.din(n28932), .dout(n28935));
    jdff dff_B_RzP8ufSE6_2(.din(n28935), .dout(n28938));
    jdff dff_B_3OaYdXdL7_2(.din(n28938), .dout(n28941));
    jdff dff_B_sIdjzXAe4_2(.din(n28941), .dout(n28944));
    jdff dff_B_iNTIn2dh8_2(.din(n28944), .dout(n28947));
    jdff dff_B_eJivWHm39_2(.din(n28947), .dout(n28950));
    jdff dff_B_OsKF9fUF4_2(.din(n28950), .dout(n28953));
    jdff dff_B_7atpzyXC7_2(.din(n28953), .dout(n28956));
    jdff dff_B_f45WlC394_2(.din(n28956), .dout(n28959));
    jdff dff_B_hbLmOOlo1_2(.din(n6496), .dout(n28962));
    jdff dff_B_YjCazqQQ3_2(.din(n28962), .dout(n28965));
    jdff dff_B_t1xsbvDJ0_2(.din(n28965), .dout(n28968));
    jdff dff_B_ZgDqR1Pc8_2(.din(n28968), .dout(n28971));
    jdff dff_B_jC8a5Z0i6_2(.din(n28971), .dout(n28974));
    jdff dff_B_CtOC030R1_2(.din(n28974), .dout(n28977));
    jdff dff_B_KvAkGQWQ1_2(.din(n28977), .dout(n28980));
    jdff dff_B_GxhBTZam8_2(.din(n28980), .dout(n28983));
    jdff dff_B_hmvdfGcC1_2(.din(n28983), .dout(n28986));
    jdff dff_B_WofEt4Ay7_2(.din(n28986), .dout(n28989));
    jdff dff_B_Dq5naBde3_2(.din(n28989), .dout(n28992));
    jdff dff_B_tM7YFD2G3_2(.din(n28992), .dout(n28995));
    jdff dff_B_ES7BqhXo1_2(.din(n28995), .dout(n28998));
    jdff dff_B_04aS6UYb8_2(.din(n28998), .dout(n29001));
    jdff dff_B_bdSMKOBd5_2(.din(n29001), .dout(n29004));
    jdff dff_B_mF38fRtk7_2(.din(n29004), .dout(n29007));
    jdff dff_B_CutgmOio5_2(.din(n29007), .dout(n29010));
    jdff dff_B_SjFGFVOn6_2(.din(n29010), .dout(n29013));
    jdff dff_B_L0kR6tUv3_2(.din(n29013), .dout(n29016));
    jdff dff_B_KI5fYqMu0_2(.din(n29016), .dout(n29019));
    jdff dff_B_iX5CW8J70_2(.din(n29019), .dout(n29022));
    jdff dff_B_YDENOHEJ1_2(.din(n29022), .dout(n29025));
    jdff dff_B_0aMEzOUL1_2(.din(n29025), .dout(n29028));
    jdff dff_B_xbVwIZ758_2(.din(n29028), .dout(n29031));
    jdff dff_B_uCaqHB5Y1_2(.din(n29031), .dout(n29034));
    jdff dff_B_lnPNylQo6_2(.din(n29034), .dout(n29037));
    jdff dff_B_0edCn8cW7_2(.din(n29037), .dout(n29040));
    jdff dff_B_tlPVmLpa7_2(.din(n29040), .dout(n29043));
    jdff dff_B_CrNf6jlH1_2(.din(n29043), .dout(n29046));
    jdff dff_B_5uTOTLMr7_2(.din(n29046), .dout(n29049));
    jdff dff_B_ayMTJqjq5_2(.din(n29049), .dout(n29052));
    jdff dff_B_ZJSE5A6u8_2(.din(n29052), .dout(n29055));
    jdff dff_B_JOaVQVlj1_2(.din(n29055), .dout(n29058));
    jdff dff_B_87GpAEat4_2(.din(n29058), .dout(n29061));
    jdff dff_B_R4e1XHKk7_2(.din(n29061), .dout(n29064));
    jdff dff_B_acDlqHo75_2(.din(n29064), .dout(n29067));
    jdff dff_B_tzmShRyT4_2(.din(n29067), .dout(n29070));
    jdff dff_B_5gTMTT226_2(.din(n29070), .dout(n29073));
    jdff dff_B_qf7enKqJ3_2(.din(n29073), .dout(n29076));
    jdff dff_B_SjS9F0V23_2(.din(n29076), .dout(n29079));
    jdff dff_B_81SDYdzI1_2(.din(n29079), .dout(n29082));
    jdff dff_B_r6NlxRvS2_2(.din(n29082), .dout(n29085));
    jdff dff_B_honvnWC47_2(.din(n29085), .dout(n29088));
    jdff dff_B_Pm4lz2TE6_2(.din(n29088), .dout(n29091));
    jdff dff_B_qNm5DonE1_2(.din(n29091), .dout(n29094));
    jdff dff_B_SV2kvBoR0_2(.din(n29094), .dout(n29097));
    jdff dff_B_EBIpuuQR8_2(.din(n29097), .dout(n29100));
    jdff dff_B_WeM40RcL6_2(.din(n6492), .dout(n29103));
    jdff dff_B_ntpkS7Lg8_1(.din(n6484), .dout(n29106));
    jdff dff_B_lG7B0dfC4_2(.din(n6346), .dout(n29109));
    jdff dff_B_KJecEGLT1_2(.din(n29109), .dout(n29112));
    jdff dff_B_5mxEd2ES5_2(.din(n29112), .dout(n29115));
    jdff dff_B_p5mWZGv34_2(.din(n29115), .dout(n29118));
    jdff dff_B_ojpNVx150_2(.din(n29118), .dout(n29121));
    jdff dff_B_si9fCXoa2_2(.din(n29121), .dout(n29124));
    jdff dff_B_OCgk9N5P9_2(.din(n29124), .dout(n29127));
    jdff dff_B_WnmibGQH6_2(.din(n29127), .dout(n29130));
    jdff dff_B_ph9dCYgJ7_2(.din(n29130), .dout(n29133));
    jdff dff_B_5VGsv4e43_2(.din(n29133), .dout(n29136));
    jdff dff_B_XZbLP5Lf1_2(.din(n29136), .dout(n29139));
    jdff dff_B_MNC0GTuQ2_2(.din(n29139), .dout(n29142));
    jdff dff_B_JbaTNY7h6_2(.din(n29142), .dout(n29145));
    jdff dff_B_HQyyC0Ks2_2(.din(n29145), .dout(n29148));
    jdff dff_B_vY6PerlF7_2(.din(n29148), .dout(n29151));
    jdff dff_B_1hAp9e208_2(.din(n29151), .dout(n29154));
    jdff dff_B_XlhxLxdf4_2(.din(n29154), .dout(n29157));
    jdff dff_B_ya1aadhD8_2(.din(n29157), .dout(n29160));
    jdff dff_B_6b2jPVpP9_2(.din(n29160), .dout(n29163));
    jdff dff_B_ls1Z6PYf3_2(.din(n29163), .dout(n29166));
    jdff dff_B_Q32PWZgJ5_2(.din(n29166), .dout(n29169));
    jdff dff_B_nOu8jI8L3_2(.din(n29169), .dout(n29172));
    jdff dff_B_ThscDitp7_2(.din(n29172), .dout(n29175));
    jdff dff_B_RJkYcvaE6_2(.din(n29175), .dout(n29178));
    jdff dff_B_XxLkv4WB8_2(.din(n29178), .dout(n29181));
    jdff dff_B_4a0Znj3O4_2(.din(n29181), .dout(n29184));
    jdff dff_B_j9tULFLz3_2(.din(n29184), .dout(n29187));
    jdff dff_B_n8hs05Cd5_2(.din(n29187), .dout(n29190));
    jdff dff_B_LPoWhfUl3_2(.din(n29190), .dout(n29193));
    jdff dff_B_j1zwFrvm4_2(.din(n29193), .dout(n29196));
    jdff dff_B_xtrKM9KJ5_2(.din(n29196), .dout(n29199));
    jdff dff_B_gStlqySk1_2(.din(n29199), .dout(n29202));
    jdff dff_B_m1XEFau04_2(.din(n29202), .dout(n29205));
    jdff dff_B_rgFpqpQt5_2(.din(n29205), .dout(n29208));
    jdff dff_B_pJTzBIea4_2(.din(n29208), .dout(n29211));
    jdff dff_B_VmGD0QdK1_2(.din(n29211), .dout(n29214));
    jdff dff_B_tL8n37lo1_2(.din(n29214), .dout(n29217));
    jdff dff_B_1EEhgPRe6_2(.din(n29217), .dout(n29220));
    jdff dff_B_W2gLu4uP4_2(.din(n29220), .dout(n29223));
    jdff dff_B_zrvBGAS09_2(.din(n29223), .dout(n29226));
    jdff dff_B_k9bITiLT4_2(.din(n29226), .dout(n29229));
    jdff dff_B_BamoOFI32_2(.din(n29229), .dout(n29232));
    jdff dff_B_kY5qNx0X4_2(.din(n29232), .dout(n29235));
    jdff dff_B_hc8D6Meq7_2(.din(n29235), .dout(n29238));
    jdff dff_B_WENRyFSp3_1(.din(n6370), .dout(n29241));
    jdff dff_B_dofnAvnv2_1(.din(n29241), .dout(n29244));
    jdff dff_B_pSBUtnzf2_2(.din(n6366), .dout(n29247));
    jdff dff_B_O3wxnIq12_2(.din(n29247), .dout(n29250));
    jdff dff_B_14OyNwMz8_2(.din(n29250), .dout(n29253));
    jdff dff_B_R2UkBLZN6_2(.din(n29253), .dout(n29256));
    jdff dff_B_Ir5t8v328_2(.din(n29256), .dout(n29259));
    jdff dff_B_vvhWlZZ94_2(.din(n29259), .dout(n29262));
    jdff dff_B_p3wJfSXo4_2(.din(n29262), .dout(n29265));
    jdff dff_B_FI3lRxcy8_2(.din(n29265), .dout(n29268));
    jdff dff_B_hUfJYE093_2(.din(n29268), .dout(n29271));
    jdff dff_B_GnXh7Pqn2_2(.din(n29271), .dout(n29274));
    jdff dff_B_98zCHcyQ2_2(.din(n29274), .dout(n29277));
    jdff dff_B_e1qiWSwR7_2(.din(n29277), .dout(n29280));
    jdff dff_B_SOnsn3GE9_2(.din(n29280), .dout(n29283));
    jdff dff_B_S6xX9IMr5_2(.din(n29283), .dout(n29286));
    jdff dff_B_U2PTNmWC1_2(.din(n29286), .dout(n29289));
    jdff dff_B_HhKI1uqI6_2(.din(n29289), .dout(n29292));
    jdff dff_B_AuJP7aRH3_2(.din(n29292), .dout(n29295));
    jdff dff_B_E4oFzWpb5_2(.din(n29295), .dout(n29298));
    jdff dff_B_hR4v2NY77_2(.din(n29298), .dout(n29301));
    jdff dff_B_vFwUmgL80_2(.din(n29301), .dout(n29304));
    jdff dff_B_CUYVvrqS3_2(.din(n29304), .dout(n29307));
    jdff dff_B_C5fZiopT0_2(.din(n29307), .dout(n29310));
    jdff dff_B_QuAmi1I34_2(.din(n29310), .dout(n29313));
    jdff dff_B_vr3iXH2W2_2(.din(n29313), .dout(n29316));
    jdff dff_B_HotQv0NS4_2(.din(n29316), .dout(n29319));
    jdff dff_B_HCGhOKUu4_2(.din(n29319), .dout(n29322));
    jdff dff_B_1MuYgIjq2_2(.din(n29322), .dout(n29325));
    jdff dff_B_MB9s2mwy8_2(.din(n29325), .dout(n29328));
    jdff dff_B_g3DZWlK20_2(.din(n29328), .dout(n29331));
    jdff dff_B_Q1XIJ01N1_2(.din(n29331), .dout(n29334));
    jdff dff_B_pl1VKKq94_2(.din(n29334), .dout(n29337));
    jdff dff_B_6M08i3Rs0_2(.din(n29337), .dout(n29340));
    jdff dff_B_ueYOJYnk6_2(.din(n29340), .dout(n29343));
    jdff dff_B_RMmkhvFz7_2(.din(n29343), .dout(n29346));
    jdff dff_B_m1BpQfr49_2(.din(n29346), .dout(n29349));
    jdff dff_B_ScpP36Ta3_2(.din(n29349), .dout(n29352));
    jdff dff_B_y7uob3vh7_2(.din(n29352), .dout(n29355));
    jdff dff_B_cSZHN7Iz6_2(.din(n29355), .dout(n29358));
    jdff dff_B_T0aF33hJ2_2(.din(n29358), .dout(n29361));
    jdff dff_B_8V6d5mBP2_2(.din(n29361), .dout(n29364));
    jdff dff_B_qvorlkVc9_2(.din(n29364), .dout(n29367));
    jdff dff_B_ORVskRRL0_2(.din(n6362), .dout(n29370));
    jdff dff_B_uFLbA16n0_2(.din(n29370), .dout(n29373));
    jdff dff_B_hPPU42YS7_2(.din(n29373), .dout(n29376));
    jdff dff_B_zSHorKoy5_2(.din(n29376), .dout(n29379));
    jdff dff_B_Dsq5ntar3_2(.din(n29379), .dout(n29382));
    jdff dff_B_hkowsfGn2_2(.din(n29382), .dout(n29385));
    jdff dff_B_zzUlKvej9_2(.din(n29385), .dout(n29388));
    jdff dff_B_nlG2aPkr8_2(.din(n29388), .dout(n29391));
    jdff dff_B_hpD5bY4P9_2(.din(n29391), .dout(n29394));
    jdff dff_B_lwvS4Zqz8_2(.din(n29394), .dout(n29397));
    jdff dff_B_h47sk5SR6_2(.din(n29397), .dout(n29400));
    jdff dff_B_z07UA75T7_2(.din(n29400), .dout(n29403));
    jdff dff_B_hoiRqGj51_2(.din(n29403), .dout(n29406));
    jdff dff_B_BU8PtD0b4_2(.din(n29406), .dout(n29409));
    jdff dff_B_ruquY5fG5_2(.din(n29409), .dout(n29412));
    jdff dff_B_ZoTcBwNy0_2(.din(n29412), .dout(n29415));
    jdff dff_B_zHr4kXGj1_2(.din(n29415), .dout(n29418));
    jdff dff_B_ACzXzg0L4_2(.din(n29418), .dout(n29421));
    jdff dff_B_rP9G3l960_2(.din(n29421), .dout(n29424));
    jdff dff_B_Rp6DzqGG0_2(.din(n29424), .dout(n29427));
    jdff dff_B_GBP0cfjm9_2(.din(n29427), .dout(n29430));
    jdff dff_B_MVtfaO6K0_2(.din(n29430), .dout(n29433));
    jdff dff_B_QXqo12Wh5_2(.din(n29433), .dout(n29436));
    jdff dff_B_X11AiJN49_2(.din(n29436), .dout(n29439));
    jdff dff_B_rSkWizs21_2(.din(n29439), .dout(n29442));
    jdff dff_B_GbEMdghI6_2(.din(n29442), .dout(n29445));
    jdff dff_B_CghXusbL2_2(.din(n29445), .dout(n29448));
    jdff dff_B_AHRYWI4h6_2(.din(n29448), .dout(n29451));
    jdff dff_B_b10RUB805_2(.din(n29451), .dout(n29454));
    jdff dff_B_E0DuHRWX5_2(.din(n29454), .dout(n29457));
    jdff dff_B_DQki4TfN8_2(.din(n29457), .dout(n29460));
    jdff dff_B_BJxRN4Rq8_2(.din(n29460), .dout(n29463));
    jdff dff_B_gUA60vJn9_2(.din(n29463), .dout(n29466));
    jdff dff_B_NKbBbhAo5_2(.din(n29466), .dout(n29469));
    jdff dff_B_OY1yIeMD6_2(.din(n29469), .dout(n29472));
    jdff dff_B_1AsiLKXu0_2(.din(n29472), .dout(n29475));
    jdff dff_B_YOk2K5Xj7_2(.din(n29475), .dout(n29478));
    jdff dff_B_5QgVmLnI6_2(.din(n29478), .dout(n29481));
    jdff dff_B_6Qk5svwe4_2(.din(n29481), .dout(n29484));
    jdff dff_B_V6ItlT3I2_2(.din(n29484), .dout(n29487));
    jdff dff_B_82aBdxM65_2(.din(n29487), .dout(n29490));
    jdff dff_B_GZT2zF813_2(.din(n29490), .dout(n29493));
    jdff dff_B_Iwu0JBoY1_2(.din(n29493), .dout(n29496));
    jdff dff_B_fSAmthdF5_2(.din(n6358), .dout(n29499));
    jdff dff_B_so3bvXCA9_1(.din(n6350), .dout(n29502));
    jdff dff_B_vtEi4Kpz3_2(.din(n6188), .dout(n29505));
    jdff dff_B_rMh5kDWf4_2(.din(n29505), .dout(n29508));
    jdff dff_B_W3huiePw8_2(.din(n29508), .dout(n29511));
    jdff dff_B_GmeMhhA71_2(.din(n29511), .dout(n29514));
    jdff dff_B_C7QERlP91_2(.din(n29514), .dout(n29517));
    jdff dff_B_84s5c5Nz2_2(.din(n29517), .dout(n29520));
    jdff dff_B_7ZW0x3g02_2(.din(n29520), .dout(n29523));
    jdff dff_B_aPDhGeFP9_2(.din(n29523), .dout(n29526));
    jdff dff_B_KaUutlwy9_2(.din(n29526), .dout(n29529));
    jdff dff_B_bySvzJn36_2(.din(n29529), .dout(n29532));
    jdff dff_B_O66wpek53_2(.din(n29532), .dout(n29535));
    jdff dff_B_aizqsT1X0_2(.din(n29535), .dout(n29538));
    jdff dff_B_aiutfzTc1_2(.din(n29538), .dout(n29541));
    jdff dff_B_12oASWHn1_2(.din(n29541), .dout(n29544));
    jdff dff_B_alXqnom34_2(.din(n29544), .dout(n29547));
    jdff dff_B_ONerYRmf7_2(.din(n29547), .dout(n29550));
    jdff dff_B_Rrpl6yNC2_2(.din(n29550), .dout(n29553));
    jdff dff_B_ix0Gi1mB1_2(.din(n29553), .dout(n29556));
    jdff dff_B_zNqUTJr67_2(.din(n29556), .dout(n29559));
    jdff dff_B_EmUI2uyv6_2(.din(n29559), .dout(n29562));
    jdff dff_B_x5jrItde3_2(.din(n29562), .dout(n29565));
    jdff dff_B_PvovAB4y7_2(.din(n29565), .dout(n29568));
    jdff dff_B_Bh9Ch4t81_2(.din(n29568), .dout(n29571));
    jdff dff_B_i92uPmxT6_2(.din(n29571), .dout(n29574));
    jdff dff_B_raTTTJJC9_2(.din(n29574), .dout(n29577));
    jdff dff_B_niThLe7M3_2(.din(n29577), .dout(n29580));
    jdff dff_B_JuaK0qrj5_2(.din(n29580), .dout(n29583));
    jdff dff_B_NBcwkllt8_2(.din(n29583), .dout(n29586));
    jdff dff_B_aYlYT9TL0_2(.din(n29586), .dout(n29589));
    jdff dff_B_0rHLpv2Q3_2(.din(n29589), .dout(n29592));
    jdff dff_B_aspizn5w9_2(.din(n29592), .dout(n29595));
    jdff dff_B_Lh31jnUz8_2(.din(n29595), .dout(n29598));
    jdff dff_B_tQKoUhBA2_2(.din(n29598), .dout(n29601));
    jdff dff_B_BaVR6MCD1_2(.din(n29601), .dout(n29604));
    jdff dff_B_Eq2yXbdA5_2(.din(n29604), .dout(n29607));
    jdff dff_B_EW9AYF2q3_2(.din(n29607), .dout(n29610));
    jdff dff_B_rjDBiP412_2(.din(n29610), .dout(n29613));
    jdff dff_B_VlbZDsvX9_2(.din(n29613), .dout(n29616));
    jdff dff_B_EZofrVWs8_2(.din(n29616), .dout(n29619));
    jdff dff_B_YSlYmL2F6_2(.din(n29619), .dout(n29622));
    jdff dff_B_Jfqm8b2C2_1(.din(n6212), .dout(n29625));
    jdff dff_B_XGro1DDU8_1(.din(n29625), .dout(n29628));
    jdff dff_B_DCt7W3KY5_2(.din(n6208), .dout(n29631));
    jdff dff_B_Ze1Gbbtc4_2(.din(n29631), .dout(n29634));
    jdff dff_B_afN3qDdr6_2(.din(n29634), .dout(n29637));
    jdff dff_B_zNipOtPz0_2(.din(n29637), .dout(n29640));
    jdff dff_B_T48beAEl9_2(.din(n29640), .dout(n29643));
    jdff dff_B_zanLY2pj5_2(.din(n29643), .dout(n29646));
    jdff dff_B_o3WkWxfY1_2(.din(n29646), .dout(n29649));
    jdff dff_B_4ODzqni49_2(.din(n29649), .dout(n29652));
    jdff dff_B_Nd0ab4CN2_2(.din(n29652), .dout(n29655));
    jdff dff_B_ZQLpiDU95_2(.din(n29655), .dout(n29658));
    jdff dff_B_mGISbn4m9_2(.din(n29658), .dout(n29661));
    jdff dff_B_lSaa4y9E0_2(.din(n29661), .dout(n29664));
    jdff dff_B_bMaQ7bwB8_2(.din(n29664), .dout(n29667));
    jdff dff_B_V7dQB2OC2_2(.din(n29667), .dout(n29670));
    jdff dff_B_cyHswZPc6_2(.din(n29670), .dout(n29673));
    jdff dff_B_24iqTy5j5_2(.din(n29673), .dout(n29676));
    jdff dff_B_8xclsG7e0_2(.din(n29676), .dout(n29679));
    jdff dff_B_wOx0yO1d7_2(.din(n29679), .dout(n29682));
    jdff dff_B_HnLvbag86_2(.din(n29682), .dout(n29685));
    jdff dff_B_1dpNgc582_2(.din(n29685), .dout(n29688));
    jdff dff_B_inlD8xDw3_2(.din(n29688), .dout(n29691));
    jdff dff_B_rpjd2GH41_2(.din(n29691), .dout(n29694));
    jdff dff_B_DjxsCOey1_2(.din(n29694), .dout(n29697));
    jdff dff_B_EF4Ictk27_2(.din(n29697), .dout(n29700));
    jdff dff_B_Mbcn8u8I1_2(.din(n29700), .dout(n29703));
    jdff dff_B_KZy9Wzyl2_2(.din(n29703), .dout(n29706));
    jdff dff_B_oTyIkkL54_2(.din(n29706), .dout(n29709));
    jdff dff_B_2Eqq8dfa6_2(.din(n29709), .dout(n29712));
    jdff dff_B_RplELcYv5_2(.din(n29712), .dout(n29715));
    jdff dff_B_Mpd7KjoO9_2(.din(n29715), .dout(n29718));
    jdff dff_B_6ZIO1vSb3_2(.din(n29718), .dout(n29721));
    jdff dff_B_r1Iwv30N4_2(.din(n29721), .dout(n29724));
    jdff dff_B_7LBpGpU68_2(.din(n29724), .dout(n29727));
    jdff dff_B_jrTO1hzs4_2(.din(n29727), .dout(n29730));
    jdff dff_B_0dPZOt1m0_2(.din(n29730), .dout(n29733));
    jdff dff_B_Xqy7mTJH3_2(.din(n29733), .dout(n29736));
    jdff dff_B_nLDF5s0E1_2(.din(n29736), .dout(n29739));
    jdff dff_B_Gn5z5N8B7_2(.din(n6204), .dout(n29742));
    jdff dff_B_oxrMN8Kh5_2(.din(n29742), .dout(n29745));
    jdff dff_B_4Na5e2Ve2_2(.din(n29745), .dout(n29748));
    jdff dff_B_mqT7sGcI9_2(.din(n29748), .dout(n29751));
    jdff dff_B_I0wq4VfE7_2(.din(n29751), .dout(n29754));
    jdff dff_B_4p7ifI9w6_2(.din(n29754), .dout(n29757));
    jdff dff_B_8KitNCqB3_2(.din(n29757), .dout(n29760));
    jdff dff_B_E8h5qvUD1_2(.din(n29760), .dout(n29763));
    jdff dff_B_wDljcrXF6_2(.din(n29763), .dout(n29766));
    jdff dff_B_FGQZMneQ8_2(.din(n29766), .dout(n29769));
    jdff dff_B_S4IAZWVB1_2(.din(n29769), .dout(n29772));
    jdff dff_B_2Kh34KYl0_2(.din(n29772), .dout(n29775));
    jdff dff_B_ZPGuMP478_2(.din(n29775), .dout(n29778));
    jdff dff_B_xxvAtJO13_2(.din(n29778), .dout(n29781));
    jdff dff_B_w8vxuQ7V0_2(.din(n29781), .dout(n29784));
    jdff dff_B_IG7nORry1_2(.din(n29784), .dout(n29787));
    jdff dff_B_PSJ3wbRG5_2(.din(n29787), .dout(n29790));
    jdff dff_B_IwR4VEJz9_2(.din(n29790), .dout(n29793));
    jdff dff_B_0AN5FYnj7_2(.din(n29793), .dout(n29796));
    jdff dff_B_rUYiWd898_2(.din(n29796), .dout(n29799));
    jdff dff_B_YAml3ti30_2(.din(n29799), .dout(n29802));
    jdff dff_B_KXMdH0Dv1_2(.din(n29802), .dout(n29805));
    jdff dff_B_GoOFHact8_2(.din(n29805), .dout(n29808));
    jdff dff_B_y1NWIWDG0_2(.din(n29808), .dout(n29811));
    jdff dff_B_2PNBIXAu4_2(.din(n29811), .dout(n29814));
    jdff dff_B_rqmfBGFq8_2(.din(n29814), .dout(n29817));
    jdff dff_B_LlQ4oQ0Q5_2(.din(n29817), .dout(n29820));
    jdff dff_B_zXddmIFX4_2(.din(n29820), .dout(n29823));
    jdff dff_B_VMphltbY0_2(.din(n29823), .dout(n29826));
    jdff dff_B_mcgQLaqK0_2(.din(n29826), .dout(n29829));
    jdff dff_B_islzgUuV1_2(.din(n29829), .dout(n29832));
    jdff dff_B_HzXEvtSl7_2(.din(n29832), .dout(n29835));
    jdff dff_B_90Nz1PCK0_2(.din(n29835), .dout(n29838));
    jdff dff_B_QcZsuWx58_2(.din(n29838), .dout(n29841));
    jdff dff_B_qpxyykvy9_2(.din(n29841), .dout(n29844));
    jdff dff_B_tjsDtm5i5_2(.din(n29844), .dout(n29847));
    jdff dff_B_PwJXIweD9_2(.din(n29847), .dout(n29850));
    jdff dff_B_f2N7aWOk5_2(.din(n29850), .dout(n29853));
    jdff dff_B_SKoI0v3m4_2(.din(n29853), .dout(n29856));
    jdff dff_B_GhTEZuUV2_2(.din(n6200), .dout(n29859));
    jdff dff_B_egK88UFU6_1(.din(n6192), .dout(n29862));
    jdff dff_B_nuPRXyN19_2(.din(n5994), .dout(n29865));
    jdff dff_B_OV3k2TzR9_2(.din(n29865), .dout(n29868));
    jdff dff_B_AkPfrcEy4_2(.din(n29868), .dout(n29871));
    jdff dff_B_B9JU5BK58_2(.din(n29871), .dout(n29874));
    jdff dff_B_95thr4gk8_2(.din(n29874), .dout(n29877));
    jdff dff_B_3Qn4gqZ09_2(.din(n29877), .dout(n29880));
    jdff dff_B_5GvkDcz38_2(.din(n29880), .dout(n29883));
    jdff dff_B_EPcGO0WF1_2(.din(n29883), .dout(n29886));
    jdff dff_B_bnL5c9sb2_2(.din(n29886), .dout(n29889));
    jdff dff_B_T8XW9peQ7_2(.din(n29889), .dout(n29892));
    jdff dff_B_9Yad3EFy0_2(.din(n29892), .dout(n29895));
    jdff dff_B_zn8z2mBb6_2(.din(n29895), .dout(n29898));
    jdff dff_B_h4DXpltR5_2(.din(n29898), .dout(n29901));
    jdff dff_B_lKBVVANg4_2(.din(n29901), .dout(n29904));
    jdff dff_B_ENot0orb1_2(.din(n29904), .dout(n29907));
    jdff dff_B_D09HICv27_2(.din(n29907), .dout(n29910));
    jdff dff_B_OAfFfalN6_2(.din(n29910), .dout(n29913));
    jdff dff_B_nMq9dOsC3_2(.din(n29913), .dout(n29916));
    jdff dff_B_K0ZaFbJq8_2(.din(n29916), .dout(n29919));
    jdff dff_B_uvcL2WJG4_2(.din(n29919), .dout(n29922));
    jdff dff_B_CZZznmh27_2(.din(n29922), .dout(n29925));
    jdff dff_B_OhNPlfJw6_2(.din(n29925), .dout(n29928));
    jdff dff_B_kW2INgSM3_2(.din(n29928), .dout(n29931));
    jdff dff_B_9bj1JdwC4_2(.din(n29931), .dout(n29934));
    jdff dff_B_KpoYko7H8_2(.din(n29934), .dout(n29937));
    jdff dff_B_x6RjqWcj0_2(.din(n29937), .dout(n29940));
    jdff dff_B_HKZYHUZX9_2(.din(n29940), .dout(n29943));
    jdff dff_B_nGncQTUi1_2(.din(n29943), .dout(n29946));
    jdff dff_B_rwrnzylx8_2(.din(n29946), .dout(n29949));
    jdff dff_B_5rPQpd1L3_2(.din(n29949), .dout(n29952));
    jdff dff_B_bExroYum5_2(.din(n29952), .dout(n29955));
    jdff dff_B_yxQpWcGX6_2(.din(n29955), .dout(n29958));
    jdff dff_B_higTDy5o0_2(.din(n29958), .dout(n29961));
    jdff dff_B_lL1HJHi17_2(.din(n29961), .dout(n29964));
    jdff dff_B_uqQT0TR96_2(.din(n29964), .dout(n29967));
    jdff dff_B_MoL9CwpP0_2(.din(n29967), .dout(n29970));
    jdff dff_B_N4JfSr7n1_1(.din(n6018), .dout(n29973));
    jdff dff_B_5qq234Sr4_1(.din(n29973), .dout(n29976));
    jdff dff_B_K68rkaQn9_2(.din(n6014), .dout(n29979));
    jdff dff_B_CiM7q6Xq9_2(.din(n29979), .dout(n29982));
    jdff dff_B_dkzLxwFq0_2(.din(n29982), .dout(n29985));
    jdff dff_B_uDDFTSOm6_2(.din(n29985), .dout(n29988));
    jdff dff_B_mgJMzQa61_2(.din(n29988), .dout(n29991));
    jdff dff_B_VrpVDPnN9_2(.din(n29991), .dout(n29994));
    jdff dff_B_G4RSUY8j0_2(.din(n29994), .dout(n29997));
    jdff dff_B_4cME2GAL0_2(.din(n29997), .dout(n30000));
    jdff dff_B_ez5PiuDK8_2(.din(n30000), .dout(n30003));
    jdff dff_B_LLI0imW92_2(.din(n30003), .dout(n30006));
    jdff dff_B_QmHDANHS5_2(.din(n30006), .dout(n30009));
    jdff dff_B_kI9ytiqq9_2(.din(n30009), .dout(n30012));
    jdff dff_B_rjTU1pez0_2(.din(n30012), .dout(n30015));
    jdff dff_B_lpMXW1jg1_2(.din(n30015), .dout(n30018));
    jdff dff_B_hoUfVHa60_2(.din(n30018), .dout(n30021));
    jdff dff_B_j0iP1Hub7_2(.din(n30021), .dout(n30024));
    jdff dff_B_aLBmGYDK6_2(.din(n30024), .dout(n30027));
    jdff dff_B_fzDOd8fJ1_2(.din(n30027), .dout(n30030));
    jdff dff_B_TpOVAHZl7_2(.din(n30030), .dout(n30033));
    jdff dff_B_NKzhgmlF2_2(.din(n30033), .dout(n30036));
    jdff dff_B_bncAS4Pf5_2(.din(n30036), .dout(n30039));
    jdff dff_B_LlbdaGVx6_2(.din(n30039), .dout(n30042));
    jdff dff_B_u1oLIKQV6_2(.din(n30042), .dout(n30045));
    jdff dff_B_uq7RaOV39_2(.din(n30045), .dout(n30048));
    jdff dff_B_auCKxZI85_2(.din(n30048), .dout(n30051));
    jdff dff_B_X5V6IUaz7_2(.din(n30051), .dout(n30054));
    jdff dff_B_eiviAIJK3_2(.din(n30054), .dout(n30057));
    jdff dff_B_BGC8ItBU0_2(.din(n30057), .dout(n30060));
    jdff dff_B_K35cnsZx0_2(.din(n30060), .dout(n30063));
    jdff dff_B_WaZa6cDR7_2(.din(n30063), .dout(n30066));
    jdff dff_B_hvBdxNAh1_2(.din(n30066), .dout(n30069));
    jdff dff_B_1Bs6bCOl1_2(.din(n30069), .dout(n30072));
    jdff dff_B_3fu1YQq02_2(.din(n30072), .dout(n30075));
    jdff dff_B_R9BpI6KK7_2(.din(n6010), .dout(n30078));
    jdff dff_B_rgqCiTNK7_2(.din(n30078), .dout(n30081));
    jdff dff_B_pW0QKm1x8_2(.din(n30081), .dout(n30084));
    jdff dff_B_xg1axJwk5_2(.din(n30084), .dout(n30087));
    jdff dff_B_z8qdQBbT6_2(.din(n30087), .dout(n30090));
    jdff dff_B_xn1SH1mG0_2(.din(n30090), .dout(n30093));
    jdff dff_B_0A83RMKG1_2(.din(n30093), .dout(n30096));
    jdff dff_B_rb4pol9V8_2(.din(n30096), .dout(n30099));
    jdff dff_B_Ih7bEQca3_2(.din(n30099), .dout(n30102));
    jdff dff_B_CXOJ9m5j8_2(.din(n30102), .dout(n30105));
    jdff dff_B_AKdxi1Rf0_2(.din(n30105), .dout(n30108));
    jdff dff_B_dHN7jQjp8_2(.din(n30108), .dout(n30111));
    jdff dff_B_mcPNcui82_2(.din(n30111), .dout(n30114));
    jdff dff_B_rzKFESw93_2(.din(n30114), .dout(n30117));
    jdff dff_B_UhrocrFL1_2(.din(n30117), .dout(n30120));
    jdff dff_B_RU89xR409_2(.din(n30120), .dout(n30123));
    jdff dff_B_fHbRt2Nq6_2(.din(n30123), .dout(n30126));
    jdff dff_B_QJgFrR4p9_2(.din(n30126), .dout(n30129));
    jdff dff_B_Sxvk3fOd2_2(.din(n30129), .dout(n30132));
    jdff dff_B_pMUf683H6_2(.din(n30132), .dout(n30135));
    jdff dff_B_2pLBPppL5_2(.din(n30135), .dout(n30138));
    jdff dff_B_jsv79wMI0_2(.din(n30138), .dout(n30141));
    jdff dff_B_8vTgenk18_2(.din(n30141), .dout(n30144));
    jdff dff_B_V1SX7UNt0_2(.din(n30144), .dout(n30147));
    jdff dff_B_31X9wV946_2(.din(n30147), .dout(n30150));
    jdff dff_B_3NQYAGCw8_2(.din(n30150), .dout(n30153));
    jdff dff_B_zSEpyaj96_2(.din(n30153), .dout(n30156));
    jdff dff_B_HKUMPwgn9_2(.din(n30156), .dout(n30159));
    jdff dff_B_o7bljNKx1_2(.din(n30159), .dout(n30162));
    jdff dff_B_vBkPOOmw4_2(.din(n30162), .dout(n30165));
    jdff dff_B_QtazNloG8_2(.din(n30165), .dout(n30168));
    jdff dff_B_rRJOtmUo5_2(.din(n30168), .dout(n30171));
    jdff dff_B_tid6EDcB4_2(.din(n30171), .dout(n30174));
    jdff dff_B_ThuaIvl45_2(.din(n30174), .dout(n30177));
    jdff dff_B_UxFdy8pr2_2(.din(n30177), .dout(n30180));
    jdff dff_B_S9b9GWiV5_2(.din(n6006), .dout(n30183));
    jdff dff_B_HJZteJoN3_1(.din(n5998), .dout(n30186));
    jdff dff_B_OmvMAqTT0_2(.din(n5776), .dout(n30189));
    jdff dff_B_pvsZFsx15_2(.din(n30189), .dout(n30192));
    jdff dff_B_AXr4O4ty0_2(.din(n30192), .dout(n30195));
    jdff dff_B_862N7lLh1_2(.din(n30195), .dout(n30198));
    jdff dff_B_P7AhAO7I5_2(.din(n30198), .dout(n30201));
    jdff dff_B_x1kZzuYt4_2(.din(n30201), .dout(n30204));
    jdff dff_B_XKApxCph2_2(.din(n30204), .dout(n30207));
    jdff dff_B_JaHfiVvu5_2(.din(n30207), .dout(n30210));
    jdff dff_B_yvXraZ4b0_2(.din(n30210), .dout(n30213));
    jdff dff_B_osxJEzY77_2(.din(n30213), .dout(n30216));
    jdff dff_B_gtYJYOf66_2(.din(n30216), .dout(n30219));
    jdff dff_B_XqkQqxjt0_2(.din(n30219), .dout(n30222));
    jdff dff_B_Oh9Z1gqE0_2(.din(n30222), .dout(n30225));
    jdff dff_B_sJ956VoH2_2(.din(n30225), .dout(n30228));
    jdff dff_B_NFSfL3w03_2(.din(n30228), .dout(n30231));
    jdff dff_B_bhMsQ0N37_2(.din(n30231), .dout(n30234));
    jdff dff_B_dWoWhe207_2(.din(n30234), .dout(n30237));
    jdff dff_B_7FrM7QSE4_2(.din(n30237), .dout(n30240));
    jdff dff_B_jp38REXl8_2(.din(n30240), .dout(n30243));
    jdff dff_B_JVrL0fzG6_2(.din(n30243), .dout(n30246));
    jdff dff_B_rgx8hFa92_2(.din(n30246), .dout(n30249));
    jdff dff_B_mqpK7Xad6_2(.din(n30249), .dout(n30252));
    jdff dff_B_zeToHgRv0_2(.din(n30252), .dout(n30255));
    jdff dff_B_EbJNOq1D7_2(.din(n30255), .dout(n30258));
    jdff dff_B_ZIMh5qSI7_2(.din(n30258), .dout(n30261));
    jdff dff_B_Ln9EsESf0_2(.din(n30261), .dout(n30264));
    jdff dff_B_trsadETY7_2(.din(n30264), .dout(n30267));
    jdff dff_B_xqcF2OXE4_2(.din(n30267), .dout(n30270));
    jdff dff_B_LCJfPLE72_2(.din(n30270), .dout(n30273));
    jdff dff_B_snsH9h506_2(.din(n30273), .dout(n30276));
    jdff dff_B_If3bHUL46_2(.din(n30276), .dout(n30279));
    jdff dff_B_vCWHOO814_2(.din(n30279), .dout(n30282));
    jdff dff_B_lyZCPGs11_1(.din(n5800), .dout(n30285));
    jdff dff_B_R8uxWo708_1(.din(n30285), .dout(n30288));
    jdff dff_B_46WPqBBn2_2(.din(n5796), .dout(n30291));
    jdff dff_B_1XWtqaD66_2(.din(n30291), .dout(n30294));
    jdff dff_B_knW16qmU7_2(.din(n30294), .dout(n30297));
    jdff dff_B_4GCSMxTt4_2(.din(n30297), .dout(n30300));
    jdff dff_B_bcXDzk9i8_2(.din(n30300), .dout(n30303));
    jdff dff_B_ssevscCk1_2(.din(n30303), .dout(n30306));
    jdff dff_B_t9CUpARs6_2(.din(n30306), .dout(n30309));
    jdff dff_B_PKkvjSv16_2(.din(n30309), .dout(n30312));
    jdff dff_B_1tQLeOoh5_2(.din(n30312), .dout(n30315));
    jdff dff_B_iQ0u0b7B8_2(.din(n30315), .dout(n30318));
    jdff dff_B_2HVBPVYn0_2(.din(n30318), .dout(n30321));
    jdff dff_B_Tmz9uCix5_2(.din(n30321), .dout(n30324));
    jdff dff_B_1a7KvG528_2(.din(n30324), .dout(n30327));
    jdff dff_B_Y5s6eiW44_2(.din(n30327), .dout(n30330));
    jdff dff_B_kqvOaVKo7_2(.din(n30330), .dout(n30333));
    jdff dff_B_r9B0GuIM5_2(.din(n30333), .dout(n30336));
    jdff dff_B_ostB113k4_2(.din(n30336), .dout(n30339));
    jdff dff_B_ivdue0726_2(.din(n30339), .dout(n30342));
    jdff dff_B_SbTmByqZ9_2(.din(n30342), .dout(n30345));
    jdff dff_B_UpzIo9X63_2(.din(n30345), .dout(n30348));
    jdff dff_B_9M1mJqd92_2(.din(n30348), .dout(n30351));
    jdff dff_B_1jWpo7Xj0_2(.din(n30351), .dout(n30354));
    jdff dff_B_AGK4g5ti1_2(.din(n30354), .dout(n30357));
    jdff dff_B_vcJ09U567_2(.din(n30357), .dout(n30360));
    jdff dff_B_uhJs6o5p9_2(.din(n30360), .dout(n30363));
    jdff dff_B_ZgdaOcBh9_2(.din(n30363), .dout(n30366));
    jdff dff_B_N5MWngKd2_2(.din(n30366), .dout(n30369));
    jdff dff_B_BtMKTer00_2(.din(n30369), .dout(n30372));
    jdff dff_B_00H811zv5_2(.din(n30372), .dout(n30375));
    jdff dff_B_XI8wn8Uu3_2(.din(n5792), .dout(n30378));
    jdff dff_B_7BwIwi7Z2_2(.din(n30378), .dout(n30381));
    jdff dff_B_K3tdjOh04_2(.din(n30381), .dout(n30384));
    jdff dff_B_nluhx48n8_2(.din(n30384), .dout(n30387));
    jdff dff_B_NZIDjwhe7_2(.din(n30387), .dout(n30390));
    jdff dff_B_Zffxkm2s6_2(.din(n30390), .dout(n30393));
    jdff dff_B_1phQhY8Q9_2(.din(n30393), .dout(n30396));
    jdff dff_B_xKjVvZqP4_2(.din(n30396), .dout(n30399));
    jdff dff_B_l0ZUqaLf9_2(.din(n30399), .dout(n30402));
    jdff dff_B_MWaep3iz6_2(.din(n30402), .dout(n30405));
    jdff dff_B_hU9AkzUJ6_2(.din(n30405), .dout(n30408));
    jdff dff_B_AjQpZnQL2_2(.din(n30408), .dout(n30411));
    jdff dff_B_JC37OW3r9_2(.din(n30411), .dout(n30414));
    jdff dff_B_hXM82lQv5_2(.din(n30414), .dout(n30417));
    jdff dff_B_TVfRBuFz0_2(.din(n30417), .dout(n30420));
    jdff dff_B_4bp5GJi99_2(.din(n30420), .dout(n30423));
    jdff dff_B_a1Q1jioX6_2(.din(n30423), .dout(n30426));
    jdff dff_B_lUUGNdUr8_2(.din(n30426), .dout(n30429));
    jdff dff_B_fLdWDGxq5_2(.din(n30429), .dout(n30432));
    jdff dff_B_2m5bpYii5_2(.din(n30432), .dout(n30435));
    jdff dff_B_NTT9AYFE1_2(.din(n30435), .dout(n30438));
    jdff dff_B_g3vSHVBW2_2(.din(n30438), .dout(n30441));
    jdff dff_B_f1BJmZyr2_2(.din(n30441), .dout(n30444));
    jdff dff_B_ZJaPvM3o5_2(.din(n30444), .dout(n30447));
    jdff dff_B_KDPqWNWF0_2(.din(n30447), .dout(n30450));
    jdff dff_B_kTuf7nG95_2(.din(n30450), .dout(n30453));
    jdff dff_B_lCJyOdvc2_2(.din(n30453), .dout(n30456));
    jdff dff_B_IH3DPNQ59_2(.din(n30456), .dout(n30459));
    jdff dff_B_dymqQGsn2_2(.din(n30459), .dout(n30462));
    jdff dff_B_6ELLYYeu3_2(.din(n30462), .dout(n30465));
    jdff dff_B_VtqpH4MQ5_2(.din(n30465), .dout(n30468));
    jdff dff_B_ipKRWSpy6_2(.din(n5788), .dout(n30471));
    jdff dff_B_plcpmFsX2_1(.din(n5780), .dout(n30474));
    jdff dff_B_Av03ybjv7_2(.din(n5531), .dout(n30477));
    jdff dff_B_TOXOZ8v72_2(.din(n30477), .dout(n30480));
    jdff dff_B_8NNliQ6X1_2(.din(n30480), .dout(n30483));
    jdff dff_B_zKqFceEj0_2(.din(n30483), .dout(n30486));
    jdff dff_B_u8HlRG636_2(.din(n30486), .dout(n30489));
    jdff dff_B_1CTfZ9rO2_2(.din(n30489), .dout(n30492));
    jdff dff_B_NFOgvyNk0_2(.din(n30492), .dout(n30495));
    jdff dff_B_l4BH1Z9j0_2(.din(n30495), .dout(n30498));
    jdff dff_B_ps38PL8f9_2(.din(n30498), .dout(n30501));
    jdff dff_B_3yStKIJO4_2(.din(n30501), .dout(n30504));
    jdff dff_B_vekcYn1c4_2(.din(n30504), .dout(n30507));
    jdff dff_B_rUxGzJKf2_2(.din(n30507), .dout(n30510));
    jdff dff_B_0GKuh1zB5_2(.din(n30510), .dout(n30513));
    jdff dff_B_8JPsKB0k2_2(.din(n30513), .dout(n30516));
    jdff dff_B_dx6bcf6z5_2(.din(n30516), .dout(n30519));
    jdff dff_B_O1DiOXmJ6_2(.din(n30519), .dout(n30522));
    jdff dff_B_vkte66X21_2(.din(n30522), .dout(n30525));
    jdff dff_B_aDINbv7V1_2(.din(n30525), .dout(n30528));
    jdff dff_B_WzghUl385_2(.din(n30528), .dout(n30531));
    jdff dff_B_z03Ap8BX4_2(.din(n30531), .dout(n30534));
    jdff dff_B_WwKReFR89_2(.din(n30534), .dout(n30537));
    jdff dff_B_0huAPqU41_2(.din(n30537), .dout(n30540));
    jdff dff_B_ucANHPEB7_2(.din(n30540), .dout(n30543));
    jdff dff_B_ULZfgP8H2_2(.din(n30543), .dout(n30546));
    jdff dff_B_hsgHv1xE6_2(.din(n30546), .dout(n30549));
    jdff dff_B_aIIDjXAm4_2(.din(n30549), .dout(n30552));
    jdff dff_B_9CVhahh19_2(.din(n30552), .dout(n30555));
    jdff dff_B_B2JJaT8Y1_2(.din(n30555), .dout(n30558));
    jdff dff_B_YFMKMXf99_1(.din(n5555), .dout(n30561));
    jdff dff_B_zBIB7LIv3_1(.din(n30561), .dout(n30564));
    jdff dff_B_2lupi1eT7_2(.din(n5551), .dout(n30567));
    jdff dff_B_lDeJkaEL8_2(.din(n30567), .dout(n30570));
    jdff dff_B_m2ps2aC25_2(.din(n30570), .dout(n30573));
    jdff dff_B_QmTK3o6b0_2(.din(n30573), .dout(n30576));
    jdff dff_B_Z0VOmMi61_2(.din(n30576), .dout(n30579));
    jdff dff_B_XLWiyqa95_2(.din(n30579), .dout(n30582));
    jdff dff_B_EA0yKMqT5_2(.din(n30582), .dout(n30585));
    jdff dff_B_uYntsCLe6_2(.din(n30585), .dout(n30588));
    jdff dff_B_W7xGSPqc6_2(.din(n30588), .dout(n30591));
    jdff dff_B_8BqnZydY8_2(.din(n30591), .dout(n30594));
    jdff dff_B_KTe0YBW91_2(.din(n30594), .dout(n30597));
    jdff dff_B_TDNCuHUh6_2(.din(n30597), .dout(n30600));
    jdff dff_B_F7zplMgm0_2(.din(n30600), .dout(n30603));
    jdff dff_B_7ziRD5KS4_2(.din(n30603), .dout(n30606));
    jdff dff_B_Zhr77VUE0_2(.din(n30606), .dout(n30609));
    jdff dff_B_HvIRCMU08_2(.din(n30609), .dout(n30612));
    jdff dff_B_Pak5dTBC9_2(.din(n30612), .dout(n30615));
    jdff dff_B_s7w1pX6x4_2(.din(n30615), .dout(n30618));
    jdff dff_B_rlNnwseh7_2(.din(n30618), .dout(n30621));
    jdff dff_B_0GkVLFEq5_2(.din(n30621), .dout(n30624));
    jdff dff_B_I4XY41NH0_2(.din(n30624), .dout(n30627));
    jdff dff_B_8NyDsdmn2_2(.din(n30627), .dout(n30630));
    jdff dff_B_8Ql4FxcU6_2(.din(n30630), .dout(n30633));
    jdff dff_B_l6HYqmoc5_2(.din(n30633), .dout(n30636));
    jdff dff_B_7pxHhch97_2(.din(n30636), .dout(n30639));
    jdff dff_B_A2NDWBwO0_2(.din(n5547), .dout(n30642));
    jdff dff_B_YNYkrfAJ7_2(.din(n30642), .dout(n30645));
    jdff dff_B_bN5RRWSv1_2(.din(n30645), .dout(n30648));
    jdff dff_B_QlHe1He51_2(.din(n30648), .dout(n30651));
    jdff dff_B_g9NgCkTW4_2(.din(n30651), .dout(n30654));
    jdff dff_B_A4GuylTi0_2(.din(n30654), .dout(n30657));
    jdff dff_B_U0GPJpZ77_2(.din(n30657), .dout(n30660));
    jdff dff_B_fZoFfEII8_2(.din(n30660), .dout(n30663));
    jdff dff_B_HUKTMELg4_2(.din(n30663), .dout(n30666));
    jdff dff_B_jqEcdhi14_2(.din(n30666), .dout(n30669));
    jdff dff_B_z3aWz5gU4_2(.din(n30669), .dout(n30672));
    jdff dff_B_GoEvd0vC6_2(.din(n30672), .dout(n30675));
    jdff dff_B_AYPZjyLs3_2(.din(n30675), .dout(n30678));
    jdff dff_B_YE4EL8mj1_2(.din(n30678), .dout(n30681));
    jdff dff_B_WzOT6QaG6_2(.din(n30681), .dout(n30684));
    jdff dff_B_efoCT5ku6_2(.din(n30684), .dout(n30687));
    jdff dff_B_jD55L0qG7_2(.din(n30687), .dout(n30690));
    jdff dff_B_QFmHvdPf5_2(.din(n30690), .dout(n30693));
    jdff dff_B_VOFMawPP0_2(.din(n30693), .dout(n30696));
    jdff dff_B_iiUpzoe22_2(.din(n30696), .dout(n30699));
    jdff dff_B_Y30VZ7cH5_2(.din(n30699), .dout(n30702));
    jdff dff_B_wgDX7S5p8_2(.din(n30702), .dout(n30705));
    jdff dff_B_uOzOINEo1_2(.din(n30705), .dout(n30708));
    jdff dff_B_pmP1MQka3_2(.din(n30708), .dout(n30711));
    jdff dff_B_lCFVNw2c2_2(.din(n30711), .dout(n30714));
    jdff dff_B_Jm9w6RiA2_2(.din(n30714), .dout(n30717));
    jdff dff_B_2BeACS201_2(.din(n30717), .dout(n30720));
    jdff dff_B_8HqNMCiP7_2(.din(n5543), .dout(n30723));
    jdff dff_B_S026EZg56_1(.din(n5535), .dout(n30726));
    jdff dff_B_II4gFpzY7_2(.din(n5259), .dout(n30729));
    jdff dff_B_p6KibwD58_2(.din(n30729), .dout(n30732));
    jdff dff_B_0NSAln6R0_2(.din(n30732), .dout(n30735));
    jdff dff_B_6GJH66ZJ3_2(.din(n30735), .dout(n30738));
    jdff dff_B_arL3XSj35_2(.din(n30738), .dout(n30741));
    jdff dff_B_uXKY5agJ5_2(.din(n30741), .dout(n30744));
    jdff dff_B_C1ODHJfy8_2(.din(n30744), .dout(n30747));
    jdff dff_B_YPbSpx0w3_2(.din(n30747), .dout(n30750));
    jdff dff_B_GS2BtMHa6_2(.din(n30750), .dout(n30753));
    jdff dff_B_3S7Xee543_2(.din(n30753), .dout(n30756));
    jdff dff_B_YIlu3IVC2_2(.din(n30756), .dout(n30759));
    jdff dff_B_mJEY2d3L8_2(.din(n30759), .dout(n30762));
    jdff dff_B_BBMuspAo1_2(.din(n30762), .dout(n30765));
    jdff dff_B_FUoJSM8P2_2(.din(n30765), .dout(n30768));
    jdff dff_B_FarZG3x59_2(.din(n30768), .dout(n30771));
    jdff dff_B_D1blQciI4_2(.din(n30771), .dout(n30774));
    jdff dff_B_PSLsGNfR4_2(.din(n30774), .dout(n30777));
    jdff dff_B_GkV0GfZV3_2(.din(n30777), .dout(n30780));
    jdff dff_B_e2573Xix1_2(.din(n30780), .dout(n30783));
    jdff dff_B_S29BS6Mz3_2(.din(n30783), .dout(n30786));
    jdff dff_B_SLJeWLzc9_2(.din(n30786), .dout(n30789));
    jdff dff_B_6IidSZij5_2(.din(n30789), .dout(n30792));
    jdff dff_B_Yun8i6zT6_2(.din(n30792), .dout(n30795));
    jdff dff_B_uNJ5Rqbx3_2(.din(n30795), .dout(n30798));
    jdff dff_B_dfts3IKL9_1(.din(n5283), .dout(n30801));
    jdff dff_B_L7a03A1l4_1(.din(n30801), .dout(n30804));
    jdff dff_B_t5tatHDx5_2(.din(n5279), .dout(n30807));
    jdff dff_B_R4NCvGAC8_2(.din(n30807), .dout(n30810));
    jdff dff_B_iXGGVD222_2(.din(n30810), .dout(n30813));
    jdff dff_B_VcZm2RMr9_2(.din(n30813), .dout(n30816));
    jdff dff_B_7DCWxgRP0_2(.din(n30816), .dout(n30819));
    jdff dff_B_FfpEEnUS0_2(.din(n30819), .dout(n30822));
    jdff dff_B_bFwnEhbF0_2(.din(n30822), .dout(n30825));
    jdff dff_B_xAT24ykD2_2(.din(n30825), .dout(n30828));
    jdff dff_B_l9Ht3rWf6_2(.din(n30828), .dout(n30831));
    jdff dff_B_OhHNcRaJ6_2(.din(n30831), .dout(n30834));
    jdff dff_B_w8ltom5m9_2(.din(n30834), .dout(n30837));
    jdff dff_B_KRVmArpG9_2(.din(n30837), .dout(n30840));
    jdff dff_B_icWNlMFz9_2(.din(n30840), .dout(n30843));
    jdff dff_B_y7zRgHsx7_2(.din(n30843), .dout(n30846));
    jdff dff_B_292f23vW9_2(.din(n30846), .dout(n30849));
    jdff dff_B_lMtldrk21_2(.din(n30849), .dout(n30852));
    jdff dff_B_V0PjiF4E6_2(.din(n30852), .dout(n30855));
    jdff dff_B_JCtWA6Zp9_2(.din(n30855), .dout(n30858));
    jdff dff_B_6Kx7oBwQ2_2(.din(n30858), .dout(n30861));
    jdff dff_B_AjSzTbXd6_2(.din(n30861), .dout(n30864));
    jdff dff_B_KO8C55j57_2(.din(n30864), .dout(n30867));
    jdff dff_B_iHBpOj256_2(.din(n5275), .dout(n30870));
    jdff dff_B_aHWJISxO2_2(.din(n30870), .dout(n30873));
    jdff dff_B_figRRYyU9_2(.din(n30873), .dout(n30876));
    jdff dff_B_3ALz3QFj1_2(.din(n30876), .dout(n30879));
    jdff dff_B_ylZUh7nx1_2(.din(n30879), .dout(n30882));
    jdff dff_B_uJHYtz8k2_2(.din(n30882), .dout(n30885));
    jdff dff_B_RA6k6S0C9_2(.din(n30885), .dout(n30888));
    jdff dff_B_lllBzQUj4_2(.din(n30888), .dout(n30891));
    jdff dff_B_o1bQoWKX9_2(.din(n30891), .dout(n30894));
    jdff dff_B_qxNWYZJC9_2(.din(n30894), .dout(n30897));
    jdff dff_B_R9FC6olV1_2(.din(n30897), .dout(n30900));
    jdff dff_B_NUWo2WtU2_2(.din(n30900), .dout(n30903));
    jdff dff_B_IXZKlPZk1_2(.din(n30903), .dout(n30906));
    jdff dff_B_28AxlOWV2_2(.din(n30906), .dout(n30909));
    jdff dff_B_gvtEs4qI3_2(.din(n30909), .dout(n30912));
    jdff dff_B_n0tCGg293_2(.din(n30912), .dout(n30915));
    jdff dff_B_dfRpefxj8_2(.din(n30915), .dout(n30918));
    jdff dff_B_HKAXMSIQ3_2(.din(n30918), .dout(n30921));
    jdff dff_B_4lF1Wtn35_2(.din(n30921), .dout(n30924));
    jdff dff_B_Ywg0Cgk01_2(.din(n30924), .dout(n30927));
    jdff dff_B_qDAYAYTz6_2(.din(n30927), .dout(n30930));
    jdff dff_B_V6JVcxgo2_2(.din(n30930), .dout(n30933));
    jdff dff_B_oHPukJZ31_2(.din(n30933), .dout(n30936));
    jdff dff_B_q8jcn1tp2_2(.din(n5271), .dout(n30939));
    jdff dff_B_Ep9cpCXH0_1(.din(n5263), .dout(n30942));
    jdff dff_B_3ltbbv398_2(.din(n4960), .dout(n30945));
    jdff dff_B_bocfXfef2_2(.din(n30945), .dout(n30948));
    jdff dff_B_GaYdGWsG5_2(.din(n30948), .dout(n30951));
    jdff dff_B_q9gaTcDu3_2(.din(n30951), .dout(n30954));
    jdff dff_B_0QW5N3qY0_2(.din(n30954), .dout(n30957));
    jdff dff_B_Aowu6DMd5_2(.din(n30957), .dout(n30960));
    jdff dff_B_GvFDmbse0_2(.din(n30960), .dout(n30963));
    jdff dff_B_HdTcVjcR1_2(.din(n30963), .dout(n30966));
    jdff dff_B_0JOnG4MU9_2(.din(n30966), .dout(n30969));
    jdff dff_B_yVQYx5ct9_2(.din(n30969), .dout(n30972));
    jdff dff_B_pMrb1zjr9_2(.din(n30972), .dout(n30975));
    jdff dff_B_w9qkHa0X9_2(.din(n30975), .dout(n30978));
    jdff dff_B_0wIZXfFx6_2(.din(n30978), .dout(n30981));
    jdff dff_B_htGTtLG31_2(.din(n30981), .dout(n30984));
    jdff dff_B_SMleNtAW7_2(.din(n30984), .dout(n30987));
    jdff dff_B_E2neHheu8_2(.din(n30987), .dout(n30990));
    jdff dff_B_Rmk0nzYJ5_2(.din(n30990), .dout(n30993));
    jdff dff_B_4zsRuMEd9_2(.din(n30993), .dout(n30996));
    jdff dff_B_qy0GjkrA5_2(.din(n30996), .dout(n30999));
    jdff dff_B_9qLTKO0M8_2(.din(n30999), .dout(n31002));
    jdff dff_B_c8bSl9KV5_1(.din(n4984), .dout(n31005));
    jdff dff_B_niqKiDNW8_1(.din(n31005), .dout(n31008));
    jdff dff_B_p0P3BqH15_2(.din(n4980), .dout(n31011));
    jdff dff_B_I62c8JQI2_2(.din(n31011), .dout(n31014));
    jdff dff_B_28qhwm4P8_2(.din(n31014), .dout(n31017));
    jdff dff_B_D3dcFmjD0_2(.din(n31017), .dout(n31020));
    jdff dff_B_C1Fw9SYq6_2(.din(n31020), .dout(n31023));
    jdff dff_B_CEKibw6u6_2(.din(n31023), .dout(n31026));
    jdff dff_B_36SM1F5p9_2(.din(n31026), .dout(n31029));
    jdff dff_B_UVad4XiN1_2(.din(n31029), .dout(n31032));
    jdff dff_B_pX10OgSl7_2(.din(n31032), .dout(n31035));
    jdff dff_B_7Ffryffh8_2(.din(n31035), .dout(n31038));
    jdff dff_B_f6WdYUHc7_2(.din(n31038), .dout(n31041));
    jdff dff_B_P76XU3xn8_2(.din(n31041), .dout(n31044));
    jdff dff_B_WGSPOU760_2(.din(n31044), .dout(n31047));
    jdff dff_B_Nbcylzl11_2(.din(n31047), .dout(n31050));
    jdff dff_B_nI0JwNwB0_2(.din(n31050), .dout(n31053));
    jdff dff_B_NAIdpmZ68_2(.din(n31053), .dout(n31056));
    jdff dff_B_6BAj7eS14_2(.din(n31056), .dout(n31059));
    jdff dff_B_YNZ0gsHV9_2(.din(n4976), .dout(n31062));
    jdff dff_B_C5oaDWd87_2(.din(n31062), .dout(n31065));
    jdff dff_B_sTy8tjPG0_2(.din(n31065), .dout(n31068));
    jdff dff_B_oGCyOuvB8_2(.din(n31068), .dout(n31071));
    jdff dff_B_dWMT7Lpx4_2(.din(n31071), .dout(n31074));
    jdff dff_B_EfmG8clW0_2(.din(n31074), .dout(n31077));
    jdff dff_B_qAGUZoC20_2(.din(n31077), .dout(n31080));
    jdff dff_B_M8j8a8cD8_2(.din(n31080), .dout(n31083));
    jdff dff_B_6vxfeEe18_2(.din(n31083), .dout(n31086));
    jdff dff_B_HnYbGdPz3_2(.din(n31086), .dout(n31089));
    jdff dff_B_rMASGJuo7_2(.din(n31089), .dout(n31092));
    jdff dff_B_qFvWF0m06_2(.din(n31092), .dout(n31095));
    jdff dff_B_Y2SThVqk4_2(.din(n31095), .dout(n31098));
    jdff dff_B_xGwlfjck2_2(.din(n31098), .dout(n31101));
    jdff dff_B_QP6s4kkk8_2(.din(n31101), .dout(n31104));
    jdff dff_B_5g7jLAsm7_2(.din(n31104), .dout(n31107));
    jdff dff_B_djCIo45C6_2(.din(n31107), .dout(n31110));
    jdff dff_B_EiNPJyiw2_2(.din(n31110), .dout(n31113));
    jdff dff_B_5rhA6zGm7_2(.din(n31113), .dout(n31116));
    jdff dff_B_AqizxOau4_1(.din(n4964), .dout(n31119));
    jdff dff_B_nz9DrSU60_2(.din(n4634), .dout(n31122));
    jdff dff_B_ntXv2OJM3_2(.din(n31122), .dout(n31125));
    jdff dff_B_PG7YBjra7_2(.din(n31125), .dout(n31128));
    jdff dff_B_5aRFOs3S3_2(.din(n31128), .dout(n31131));
    jdff dff_B_VoPP6YrR0_2(.din(n31131), .dout(n31134));
    jdff dff_B_vEotDmyG3_2(.din(n31134), .dout(n31137));
    jdff dff_B_Yq6fbw8A8_2(.din(n31137), .dout(n31140));
    jdff dff_B_LZG5QkFe4_2(.din(n31140), .dout(n31143));
    jdff dff_B_YLNYEWHh0_2(.din(n31143), .dout(n31146));
    jdff dff_B_6ywo4OgW3_2(.din(n31146), .dout(n31149));
    jdff dff_B_wsuBI3Td1_2(.din(n31149), .dout(n31152));
    jdff dff_B_jt55LJ7J9_2(.din(n31152), .dout(n31155));
    jdff dff_B_1vZzD2DW9_2(.din(n31155), .dout(n31158));
    jdff dff_B_wxBL12NL9_2(.din(n31158), .dout(n31161));
    jdff dff_B_Hw4blZWM1_2(.din(n31161), .dout(n31164));
    jdff dff_B_dS6gl4Jj2_2(.din(n31164), .dout(n31167));
endmodule

