/*

c6288:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jdff: 1628
	jand: 664
	jor: 312

Summary:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jdff: 1628
	jand: 664
	jor: 312

The maximum logic level gap of any gate:
	c6288: 57
*/

module gf_c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G1gat_1;
	wire[2:0] w_G1gat_2;
	wire[2:0] w_G1gat_3;
	wire[2:0] w_G1gat_4;
	wire[2:0] w_G1gat_5;
	wire[2:0] w_G1gat_6;
	wire[1:0] w_G1gat_7;
	wire[2:0] w_G18gat_0;
	wire[2:0] w_G18gat_1;
	wire[2:0] w_G18gat_2;
	wire[2:0] w_G18gat_3;
	wire[2:0] w_G18gat_4;
	wire[2:0] w_G18gat_5;
	wire[2:0] w_G18gat_6;
	wire[1:0] w_G18gat_7;
	wire[2:0] w_G35gat_0;
	wire[2:0] w_G35gat_1;
	wire[2:0] w_G35gat_2;
	wire[2:0] w_G35gat_3;
	wire[2:0] w_G35gat_4;
	wire[2:0] w_G35gat_5;
	wire[2:0] w_G35gat_6;
	wire[2:0] w_G35gat_7;
	wire[2:0] w_G52gat_0;
	wire[2:0] w_G52gat_1;
	wire[2:0] w_G52gat_2;
	wire[2:0] w_G52gat_3;
	wire[2:0] w_G52gat_4;
	wire[2:0] w_G52gat_5;
	wire[2:0] w_G52gat_6;
	wire[2:0] w_G52gat_7;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G69gat_1;
	wire[2:0] w_G69gat_2;
	wire[2:0] w_G69gat_3;
	wire[2:0] w_G69gat_4;
	wire[2:0] w_G69gat_5;
	wire[2:0] w_G69gat_6;
	wire[1:0] w_G69gat_7;
	wire[2:0] w_G86gat_0;
	wire[2:0] w_G86gat_1;
	wire[2:0] w_G86gat_2;
	wire[2:0] w_G86gat_3;
	wire[2:0] w_G86gat_4;
	wire[2:0] w_G86gat_5;
	wire[2:0] w_G86gat_6;
	wire[1:0] w_G86gat_7;
	wire[2:0] w_G103gat_0;
	wire[2:0] w_G103gat_1;
	wire[2:0] w_G103gat_2;
	wire[2:0] w_G103gat_3;
	wire[2:0] w_G103gat_4;
	wire[2:0] w_G103gat_5;
	wire[2:0] w_G103gat_6;
	wire[1:0] w_G103gat_7;
	wire[2:0] w_G120gat_0;
	wire[2:0] w_G120gat_1;
	wire[2:0] w_G120gat_2;
	wire[2:0] w_G120gat_3;
	wire[2:0] w_G120gat_4;
	wire[2:0] w_G120gat_5;
	wire[2:0] w_G120gat_6;
	wire[1:0] w_G120gat_7;
	wire[2:0] w_G137gat_0;
	wire[2:0] w_G137gat_1;
	wire[2:0] w_G137gat_2;
	wire[2:0] w_G137gat_3;
	wire[2:0] w_G137gat_4;
	wire[2:0] w_G137gat_5;
	wire[2:0] w_G137gat_6;
	wire[1:0] w_G137gat_7;
	wire[2:0] w_G154gat_0;
	wire[2:0] w_G154gat_1;
	wire[2:0] w_G154gat_2;
	wire[2:0] w_G154gat_3;
	wire[2:0] w_G154gat_4;
	wire[2:0] w_G154gat_5;
	wire[2:0] w_G154gat_6;
	wire[1:0] w_G154gat_7;
	wire[2:0] w_G171gat_0;
	wire[2:0] w_G171gat_1;
	wire[2:0] w_G171gat_2;
	wire[2:0] w_G171gat_3;
	wire[2:0] w_G171gat_4;
	wire[2:0] w_G171gat_5;
	wire[2:0] w_G171gat_6;
	wire[1:0] w_G171gat_7;
	wire[2:0] w_G188gat_0;
	wire[2:0] w_G188gat_1;
	wire[2:0] w_G188gat_2;
	wire[2:0] w_G188gat_3;
	wire[2:0] w_G188gat_4;
	wire[2:0] w_G188gat_5;
	wire[2:0] w_G188gat_6;
	wire[1:0] w_G188gat_7;
	wire[2:0] w_G205gat_0;
	wire[2:0] w_G205gat_1;
	wire[2:0] w_G205gat_2;
	wire[2:0] w_G205gat_3;
	wire[2:0] w_G205gat_4;
	wire[2:0] w_G205gat_5;
	wire[2:0] w_G205gat_6;
	wire[1:0] w_G205gat_7;
	wire[2:0] w_G222gat_0;
	wire[2:0] w_G222gat_1;
	wire[2:0] w_G222gat_2;
	wire[2:0] w_G222gat_3;
	wire[2:0] w_G222gat_4;
	wire[2:0] w_G222gat_5;
	wire[2:0] w_G222gat_6;
	wire[1:0] w_G222gat_7;
	wire[2:0] w_G239gat_0;
	wire[2:0] w_G239gat_1;
	wire[2:0] w_G239gat_2;
	wire[2:0] w_G239gat_3;
	wire[2:0] w_G239gat_4;
	wire[2:0] w_G239gat_5;
	wire[2:0] w_G239gat_6;
	wire[1:0] w_G239gat_7;
	wire[2:0] w_G256gat_0;
	wire[2:0] w_G256gat_1;
	wire[2:0] w_G256gat_2;
	wire[2:0] w_G256gat_3;
	wire[2:0] w_G256gat_4;
	wire[2:0] w_G256gat_5;
	wire[2:0] w_G256gat_6;
	wire[1:0] w_G256gat_7;
	wire[2:0] w_G273gat_0;
	wire[2:0] w_G273gat_1;
	wire[2:0] w_G273gat_2;
	wire[2:0] w_G273gat_3;
	wire[2:0] w_G273gat_4;
	wire[2:0] w_G273gat_5;
	wire[2:0] w_G273gat_6;
	wire[1:0] w_G273gat_7;
	wire[2:0] w_G290gat_0;
	wire[2:0] w_G290gat_1;
	wire[2:0] w_G290gat_2;
	wire[2:0] w_G290gat_3;
	wire[2:0] w_G290gat_4;
	wire[2:0] w_G290gat_5;
	wire[2:0] w_G290gat_6;
	wire[2:0] w_G290gat_7;
	wire[2:0] w_G307gat_0;
	wire[2:0] w_G307gat_1;
	wire[2:0] w_G307gat_2;
	wire[2:0] w_G307gat_3;
	wire[2:0] w_G307gat_4;
	wire[2:0] w_G307gat_5;
	wire[2:0] w_G307gat_6;
	wire[1:0] w_G307gat_7;
	wire[2:0] w_G324gat_0;
	wire[2:0] w_G324gat_1;
	wire[2:0] w_G324gat_2;
	wire[2:0] w_G324gat_3;
	wire[2:0] w_G324gat_4;
	wire[2:0] w_G324gat_5;
	wire[2:0] w_G324gat_6;
	wire[1:0] w_G324gat_7;
	wire[2:0] w_G341gat_0;
	wire[2:0] w_G341gat_1;
	wire[2:0] w_G341gat_2;
	wire[2:0] w_G341gat_3;
	wire[2:0] w_G341gat_4;
	wire[2:0] w_G341gat_5;
	wire[2:0] w_G341gat_6;
	wire[1:0] w_G341gat_7;
	wire[2:0] w_G358gat_0;
	wire[2:0] w_G358gat_1;
	wire[2:0] w_G358gat_2;
	wire[2:0] w_G358gat_3;
	wire[2:0] w_G358gat_4;
	wire[2:0] w_G358gat_5;
	wire[2:0] w_G358gat_6;
	wire[1:0] w_G358gat_7;
	wire[2:0] w_G375gat_0;
	wire[2:0] w_G375gat_1;
	wire[2:0] w_G375gat_2;
	wire[2:0] w_G375gat_3;
	wire[2:0] w_G375gat_4;
	wire[2:0] w_G375gat_5;
	wire[2:0] w_G375gat_6;
	wire[1:0] w_G375gat_7;
	wire[2:0] w_G392gat_0;
	wire[2:0] w_G392gat_1;
	wire[2:0] w_G392gat_2;
	wire[2:0] w_G392gat_3;
	wire[2:0] w_G392gat_4;
	wire[2:0] w_G392gat_5;
	wire[2:0] w_G392gat_6;
	wire[1:0] w_G392gat_7;
	wire[2:0] w_G409gat_0;
	wire[2:0] w_G409gat_1;
	wire[2:0] w_G409gat_2;
	wire[2:0] w_G409gat_3;
	wire[2:0] w_G409gat_4;
	wire[2:0] w_G409gat_5;
	wire[2:0] w_G409gat_6;
	wire[1:0] w_G409gat_7;
	wire[2:0] w_G426gat_0;
	wire[2:0] w_G426gat_1;
	wire[2:0] w_G426gat_2;
	wire[2:0] w_G426gat_3;
	wire[2:0] w_G426gat_4;
	wire[2:0] w_G426gat_5;
	wire[2:0] w_G426gat_6;
	wire[1:0] w_G426gat_7;
	wire[2:0] w_G443gat_0;
	wire[2:0] w_G443gat_1;
	wire[2:0] w_G443gat_2;
	wire[2:0] w_G443gat_3;
	wire[2:0] w_G443gat_4;
	wire[2:0] w_G443gat_5;
	wire[2:0] w_G443gat_6;
	wire[1:0] w_G443gat_7;
	wire[2:0] w_G460gat_0;
	wire[2:0] w_G460gat_1;
	wire[2:0] w_G460gat_2;
	wire[2:0] w_G460gat_3;
	wire[2:0] w_G460gat_4;
	wire[2:0] w_G460gat_5;
	wire[2:0] w_G460gat_6;
	wire[1:0] w_G460gat_7;
	wire[2:0] w_G477gat_0;
	wire[2:0] w_G477gat_1;
	wire[2:0] w_G477gat_2;
	wire[2:0] w_G477gat_3;
	wire[2:0] w_G477gat_4;
	wire[2:0] w_G477gat_5;
	wire[2:0] w_G477gat_6;
	wire[1:0] w_G477gat_7;
	wire[2:0] w_G494gat_0;
	wire[2:0] w_G494gat_1;
	wire[2:0] w_G494gat_2;
	wire[2:0] w_G494gat_3;
	wire[2:0] w_G494gat_4;
	wire[2:0] w_G494gat_5;
	wire[2:0] w_G494gat_6;
	wire[1:0] w_G494gat_7;
	wire[2:0] w_G511gat_0;
	wire[2:0] w_G511gat_1;
	wire[2:0] w_G511gat_2;
	wire[2:0] w_G511gat_3;
	wire[2:0] w_G511gat_4;
	wire[2:0] w_G511gat_5;
	wire[2:0] w_G511gat_6;
	wire[1:0] w_G511gat_7;
	wire[2:0] w_G528gat_0;
	wire[2:0] w_G528gat_1;
	wire[2:0] w_G528gat_2;
	wire[2:0] w_G528gat_3;
	wire[2:0] w_G528gat_4;
	wire[2:0] w_G528gat_5;
	wire[2:0] w_G528gat_6;
	wire[1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire[1:0] w_n65_0;
	wire[1:0] w_n66_0;
	wire[1:0] w_n67_0;
	wire[1:0] w_n69_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n75_0;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[2:0] w_n80_0;
	wire[1:0] w_n83_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[1:0] w_n90_0;
	wire[1:0] w_n91_0;
	wire[1:0] w_n93_0;
	wire[1:0] w_n97_0;
	wire[1:0] w_n99_0;
	wire[2:0] w_n101_0;
	wire[1:0] w_n103_0;
	wire[1:0] w_n104_0;
	wire[1:0] w_n106_0;
	wire[1:0] w_n111_0;
	wire[1:0] w_n112_0;
	wire[2:0] w_n117_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[1:0] w_n121_0;
	wire[1:0] w_n122_0;
	wire[1:0] w_n123_0;
	wire[1:0] w_n125_0;
	wire[1:0] w_n127_0;
	wire[1:0] w_n128_0;
	wire[1:0] w_n129_0;
	wire[1:0] w_n130_0;
	wire[1:0] w_n132_0;
	wire[1:0] w_n133_0;
	wire[1:0] w_n135_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n141_0;
	wire[2:0] w_n146_0;
	wire[1:0] w_n148_0;
	wire[1:0] w_n152_0;
	wire[1:0] w_n154_0;
	wire[1:0] w_n155_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n157_0;
	wire[1:0] w_n158_0;
	wire[1:0] w_n160_0;
	wire[1:0] w_n161_0;
	wire[1:0] w_n162_0;
	wire[1:0] w_n163_0;
	wire[1:0] w_n164_0;
	wire[1:0] w_n165_0;
	wire[1:0] w_n167_0;
	wire[1:0] w_n168_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n175_0;
	wire[1:0] w_n176_0;
	wire[2:0] w_n181_0;
	wire[1:0] w_n183_0;
	wire[1:0] w_n186_0;
	wire[1:0] w_n188_0;
	wire[1:0] w_n192_0;
	wire[1:0] w_n194_0;
	wire[1:0] w_n195_0;
	wire[2:0] w_n196_0;
	wire[1:0] w_n198_0;
	wire[1:0] w_n200_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n202_0;
	wire[1:0] w_n203_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n205_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n207_0;
	wire[1:0] w_n209_0;
	wire[1:0] w_n210_0;
	wire[1:0] w_n212_0;
	wire[1:0] w_n217_0;
	wire[1:0] w_n218_0;
	wire[2:0] w_n223_0;
	wire[1:0] w_n225_0;
	wire[1:0] w_n228_0;
	wire[1:0] w_n230_0;
	wire[1:0] w_n233_0;
	wire[1:0] w_n235_0;
	wire[1:0] w_n239_0;
	wire[1:0] w_n241_0;
	wire[1:0] w_n242_0;
	wire[2:0] w_n243_0;
	wire[1:0] w_n245_0;
	wire[1:0] w_n247_0;
	wire[1:0] w_n248_0;
	wire[1:0] w_n249_0;
	wire[1:0] w_n250_0;
	wire[1:0] w_n251_0;
	wire[1:0] w_n252_0;
	wire[1:0] w_n253_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n255_0;
	wire[1:0] w_n256_0;
	wire[1:0] w_n258_0;
	wire[1:0] w_n259_0;
	wire[1:0] w_n261_0;
	wire[1:0] w_n266_0;
	wire[1:0] w_n267_0;
	wire[2:0] w_n272_0;
	wire[1:0] w_n274_0;
	wire[1:0] w_n277_0;
	wire[1:0] w_n279_0;
	wire[1:0] w_n282_0;
	wire[1:0] w_n284_0;
	wire[1:0] w_n287_0;
	wire[1:0] w_n289_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n295_0;
	wire[1:0] w_n296_0;
	wire[2:0] w_n297_0;
	wire[1:0] w_n299_0;
	wire[1:0] w_n301_0;
	wire[1:0] w_n302_0;
	wire[1:0] w_n303_0;
	wire[1:0] w_n304_0;
	wire[1:0] w_n305_0;
	wire[1:0] w_n306_0;
	wire[1:0] w_n307_0;
	wire[1:0] w_n308_0;
	wire[1:0] w_n309_0;
	wire[1:0] w_n310_0;
	wire[1:0] w_n311_0;
	wire[1:0] w_n312_0;
	wire[1:0] w_n314_0;
	wire[1:0] w_n315_0;
	wire[1:0] w_n317_0;
	wire[1:0] w_n322_0;
	wire[1:0] w_n323_0;
	wire[2:0] w_n328_0;
	wire[1:0] w_n330_0;
	wire[1:0] w_n333_0;
	wire[1:0] w_n335_0;
	wire[1:0] w_n338_0;
	wire[1:0] w_n340_0;
	wire[1:0] w_n343_0;
	wire[1:0] w_n345_0;
	wire[1:0] w_n348_0;
	wire[1:0] w_n350_0;
	wire[1:0] w_n354_0;
	wire[1:0] w_n356_0;
	wire[1:0] w_n357_0;
	wire[2:0] w_n358_0;
	wire[1:0] w_n360_0;
	wire[1:0] w_n362_0;
	wire[1:0] w_n363_0;
	wire[1:0] w_n364_0;
	wire[1:0] w_n365_0;
	wire[1:0] w_n366_0;
	wire[1:0] w_n367_0;
	wire[1:0] w_n368_0;
	wire[1:0] w_n369_0;
	wire[1:0] w_n370_0;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n373_0;
	wire[1:0] w_n374_0;
	wire[1:0] w_n375_0;
	wire[1:0] w_n377_0;
	wire[1:0] w_n378_0;
	wire[1:0] w_n380_0;
	wire[1:0] w_n385_0;
	wire[1:0] w_n386_0;
	wire[2:0] w_n391_0;
	wire[1:0] w_n393_0;
	wire[1:0] w_n396_0;
	wire[1:0] w_n398_0;
	wire[1:0] w_n401_0;
	wire[1:0] w_n403_0;
	wire[1:0] w_n406_0;
	wire[1:0] w_n408_0;
	wire[1:0] w_n411_0;
	wire[1:0] w_n413_0;
	wire[1:0] w_n416_0;
	wire[1:0] w_n418_0;
	wire[1:0] w_n423_0;
	wire[1:0] w_n425_0;
	wire[1:0] w_n426_0;
	wire[2:0] w_n427_0;
	wire[1:0] w_n429_0;
	wire[1:0] w_n431_0;
	wire[1:0] w_n432_0;
	wire[1:0] w_n433_0;
	wire[1:0] w_n434_0;
	wire[1:0] w_n435_0;
	wire[1:0] w_n436_0;
	wire[1:0] w_n437_0;
	wire[1:0] w_n438_0;
	wire[1:0] w_n439_0;
	wire[1:0] w_n440_0;
	wire[1:0] w_n441_0;
	wire[1:0] w_n442_0;
	wire[1:0] w_n443_0;
	wire[1:0] w_n444_0;
	wire[1:0] w_n445_0;
	wire[1:0] w_n446_0;
	wire[1:0] w_n448_0;
	wire[1:0] w_n449_0;
	wire[1:0] w_n451_0;
	wire[1:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[2:0] w_n462_0;
	wire[1:0] w_n464_0;
	wire[1:0] w_n467_0;
	wire[1:0] w_n469_0;
	wire[1:0] w_n472_0;
	wire[1:0] w_n474_0;
	wire[1:0] w_n477_0;
	wire[1:0] w_n479_0;
	wire[1:0] w_n482_0;
	wire[1:0] w_n484_0;
	wire[1:0] w_n487_0;
	wire[1:0] w_n489_0;
	wire[1:0] w_n492_0;
	wire[1:0] w_n494_0;
	wire[1:0] w_n499_0;
	wire[1:0] w_n501_0;
	wire[1:0] w_n502_0;
	wire[2:0] w_n503_0;
	wire[1:0] w_n505_0;
	wire[1:0] w_n507_0;
	wire[1:0] w_n508_0;
	wire[1:0] w_n509_0;
	wire[1:0] w_n510_0;
	wire[1:0] w_n511_0;
	wire[1:0] w_n512_0;
	wire[1:0] w_n513_0;
	wire[1:0] w_n514_0;
	wire[1:0] w_n515_0;
	wire[1:0] w_n516_0;
	wire[1:0] w_n517_0;
	wire[1:0] w_n518_0;
	wire[1:0] w_n519_0;
	wire[1:0] w_n520_0;
	wire[1:0] w_n521_0;
	wire[1:0] w_n522_0;
	wire[1:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n526_0;
	wire[1:0] w_n527_0;
	wire[1:0] w_n529_0;
	wire[1:0] w_n534_0;
	wire[1:0] w_n535_0;
	wire[2:0] w_n540_0;
	wire[1:0] w_n542_0;
	wire[1:0] w_n545_0;
	wire[1:0] w_n547_0;
	wire[1:0] w_n550_0;
	wire[1:0] w_n552_0;
	wire[1:0] w_n555_0;
	wire[1:0] w_n557_0;
	wire[1:0] w_n560_0;
	wire[1:0] w_n562_0;
	wire[1:0] w_n565_0;
	wire[1:0] w_n567_0;
	wire[1:0] w_n570_0;
	wire[1:0] w_n572_0;
	wire[1:0] w_n575_0;
	wire[1:0] w_n577_0;
	wire[1:0] w_n582_0;
	wire[1:0] w_n584_0;
	wire[1:0] w_n585_0;
	wire[2:0] w_n586_0;
	wire[1:0] w_n588_0;
	wire[1:0] w_n590_0;
	wire[1:0] w_n591_0;
	wire[1:0] w_n592_0;
	wire[1:0] w_n593_0;
	wire[1:0] w_n594_0;
	wire[1:0] w_n595_0;
	wire[1:0] w_n596_0;
	wire[1:0] w_n597_0;
	wire[1:0] w_n598_0;
	wire[1:0] w_n599_0;
	wire[1:0] w_n600_0;
	wire[1:0] w_n601_0;
	wire[1:0] w_n602_0;
	wire[1:0] w_n603_0;
	wire[1:0] w_n604_0;
	wire[1:0] w_n605_0;
	wire[1:0] w_n606_0;
	wire[1:0] w_n607_0;
	wire[1:0] w_n608_0;
	wire[1:0] w_n609_0;
	wire[1:0] w_n611_0;
	wire[1:0] w_n612_0;
	wire[1:0] w_n614_0;
	wire[1:0] w_n619_0;
	wire[1:0] w_n620_0;
	wire[2:0] w_n625_0;
	wire[1:0] w_n627_0;
	wire[1:0] w_n630_0;
	wire[1:0] w_n632_0;
	wire[1:0] w_n635_0;
	wire[1:0] w_n637_0;
	wire[1:0] w_n640_0;
	wire[1:0] w_n642_0;
	wire[1:0] w_n645_0;
	wire[1:0] w_n647_0;
	wire[1:0] w_n650_0;
	wire[1:0] w_n652_0;
	wire[1:0] w_n655_0;
	wire[1:0] w_n657_0;
	wire[1:0] w_n660_0;
	wire[1:0] w_n662_0;
	wire[1:0] w_n665_0;
	wire[1:0] w_n667_0;
	wire[1:0] w_n672_0;
	wire[1:0] w_n674_0;
	wire[1:0] w_n675_0;
	wire[2:0] w_n676_0;
	wire[1:0] w_n678_0;
	wire[1:0] w_n680_0;
	wire[1:0] w_n681_0;
	wire[1:0] w_n682_0;
	wire[1:0] w_n683_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n685_0;
	wire[1:0] w_n686_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n688_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n691_0;
	wire[1:0] w_n692_0;
	wire[1:0] w_n693_0;
	wire[1:0] w_n694_0;
	wire[1:0] w_n695_0;
	wire[1:0] w_n696_0;
	wire[1:0] w_n697_0;
	wire[1:0] w_n698_0;
	wire[1:0] w_n699_0;
	wire[1:0] w_n700_0;
	wire[1:0] w_n701_0;
	wire[1:0] w_n703_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n706_0;
	wire[1:0] w_n711_0;
	wire[1:0] w_n712_0;
	wire[2:0] w_n717_0;
	wire[1:0] w_n719_0;
	wire[1:0] w_n722_0;
	wire[1:0] w_n724_0;
	wire[1:0] w_n727_0;
	wire[1:0] w_n729_0;
	wire[1:0] w_n732_0;
	wire[1:0] w_n734_0;
	wire[1:0] w_n737_0;
	wire[1:0] w_n739_0;
	wire[1:0] w_n742_0;
	wire[1:0] w_n744_0;
	wire[1:0] w_n747_0;
	wire[1:0] w_n749_0;
	wire[1:0] w_n752_0;
	wire[1:0] w_n754_0;
	wire[1:0] w_n757_0;
	wire[1:0] w_n759_0;
	wire[1:0] w_n762_0;
	wire[1:0] w_n764_0;
	wire[1:0] w_n769_0;
	wire[1:0] w_n771_0;
	wire[1:0] w_n772_0;
	wire[1:0] w_n773_0;
	wire[1:0] w_n774_0;
	wire[1:0] w_n775_0;
	wire[1:0] w_n777_0;
	wire[1:0] w_n778_0;
	wire[1:0] w_n779_0;
	wire[1:0] w_n780_0;
	wire[1:0] w_n781_0;
	wire[1:0] w_n782_0;
	wire[1:0] w_n783_0;
	wire[1:0] w_n784_0;
	wire[1:0] w_n785_0;
	wire[1:0] w_n786_0;
	wire[1:0] w_n787_0;
	wire[1:0] w_n788_0;
	wire[1:0] w_n789_0;
	wire[1:0] w_n790_0;
	wire[1:0] w_n791_0;
	wire[1:0] w_n792_0;
	wire[1:0] w_n793_0;
	wire[1:0] w_n794_0;
	wire[1:0] w_n795_0;
	wire[1:0] w_n796_0;
	wire[1:0] w_n797_0;
	wire[1:0] w_n798_0;
	wire[1:0] w_n799_0;
	wire[1:0] w_n800_0;
	wire[1:0] w_n802_0;
	wire[1:0] w_n803_0;
	wire[1:0] w_n805_0;
	wire[1:0] w_n810_0;
	wire[1:0] w_n811_0;
	wire[1:0] w_n815_0;
	wire[1:0] w_n816_0;
	wire[2:0] w_n820_0;
	wire[1:0] w_n822_0;
	wire[1:0] w_n825_0;
	wire[1:0] w_n827_0;
	wire[1:0] w_n830_0;
	wire[1:0] w_n832_0;
	wire[1:0] w_n835_0;
	wire[1:0] w_n837_0;
	wire[1:0] w_n840_0;
	wire[1:0] w_n842_0;
	wire[1:0] w_n845_0;
	wire[1:0] w_n847_0;
	wire[1:0] w_n850_0;
	wire[1:0] w_n852_0;
	wire[1:0] w_n855_0;
	wire[1:0] w_n857_0;
	wire[1:0] w_n860_0;
	wire[1:0] w_n862_0;
	wire[1:0] w_n865_0;
	wire[1:0] w_n867_0;
	wire[1:0] w_n872_0;
	wire[1:0] w_n874_0;
	wire[1:0] w_n875_0;
	wire[1:0] w_n877_0;
	wire[1:0] w_n879_0;
	wire[1:0] w_n880_0;
	wire[1:0] w_n881_0;
	wire[1:0] w_n882_0;
	wire[1:0] w_n883_0;
	wire[1:0] w_n884_0;
	wire[1:0] w_n885_0;
	wire[1:0] w_n886_0;
	wire[1:0] w_n887_0;
	wire[1:0] w_n888_0;
	wire[1:0] w_n889_0;
	wire[1:0] w_n890_0;
	wire[1:0] w_n891_0;
	wire[1:0] w_n892_0;
	wire[1:0] w_n893_0;
	wire[1:0] w_n894_0;
	wire[1:0] w_n895_0;
	wire[1:0] w_n896_0;
	wire[1:0] w_n897_0;
	wire[1:0] w_n898_0;
	wire[1:0] w_n899_0;
	wire[2:0] w_n900_0;
	wire[1:0] w_n902_0;
	wire[1:0] w_n903_0;
	wire[1:0] w_n904_0;
	wire[1:0] w_n905_0;
	wire[1:0] w_n910_0;
	wire[1:0] w_n911_0;
	wire[2:0] w_n915_0;
	wire[1:0] w_n916_0;
	wire[1:0] w_n922_0;
	wire[1:0] w_n924_0;
	wire[1:0] w_n927_0;
	wire[1:0] w_n929_0;
	wire[1:0] w_n932_0;
	wire[1:0] w_n934_0;
	wire[1:0] w_n937_0;
	wire[1:0] w_n939_0;
	wire[1:0] w_n942_0;
	wire[1:0] w_n944_0;
	wire[1:0] w_n947_0;
	wire[1:0] w_n949_0;
	wire[1:0] w_n952_0;
	wire[1:0] w_n954_0;
	wire[1:0] w_n957_0;
	wire[1:0] w_n959_0;
	wire[1:0] w_n962_0;
	wire[1:0] w_n964_0;
	wire[1:0] w_n967_0;
	wire[1:0] w_n969_0;
	wire[1:0] w_n972_0;
	wire[1:0] w_n974_0;
	wire[1:0] w_n978_0;
	wire[1:0] w_n980_0;
	wire[1:0] w_n982_0;
	wire[1:0] w_n983_0;
	wire[1:0] w_n984_0;
	wire[1:0] w_n985_0;
	wire[1:0] w_n986_0;
	wire[1:0] w_n987_0;
	wire[1:0] w_n988_0;
	wire[1:0] w_n989_0;
	wire[1:0] w_n990_0;
	wire[1:0] w_n991_0;
	wire[1:0] w_n992_0;
	wire[1:0] w_n993_0;
	wire[1:0] w_n994_0;
	wire[1:0] w_n995_0;
	wire[1:0] w_n996_0;
	wire[1:0] w_n997_0;
	wire[1:0] w_n998_0;
	wire[1:0] w_n999_0;
	wire[1:0] w_n1000_0;
	wire[1:0] w_n1001_0;
	wire[1:0] w_n1002_0;
	wire[1:0] w_n1003_0;
	wire[1:0] w_n1004_0;
	wire[1:0] w_n1005_0;
	wire[1:0] w_n1006_0;
	wire[1:0] w_n1007_0;
	wire[1:0] w_n1008_0;
	wire[1:0] w_n1009_0;
	wire[1:0] w_n1011_0;
	wire[1:0] w_n1013_0;
	wire[1:0] w_n1017_0;
	wire[1:0] w_n1018_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1023_0;
	wire[1:0] w_n1026_0;
	wire[1:0] w_n1028_0;
	wire[1:0] w_n1031_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1036_0;
	wire[1:0] w_n1038_0;
	wire[1:0] w_n1041_0;
	wire[1:0] w_n1043_0;
	wire[1:0] w_n1046_0;
	wire[1:0] w_n1048_0;
	wire[1:0] w_n1051_0;
	wire[1:0] w_n1053_0;
	wire[1:0] w_n1056_0;
	wire[1:0] w_n1058_0;
	wire[1:0] w_n1061_0;
	wire[1:0] w_n1063_0;
	wire[1:0] w_n1066_0;
	wire[1:0] w_n1068_0;
	wire[1:0] w_n1071_0;
	wire[1:0] w_n1073_0;
	wire[1:0] w_n1076_0;
	wire[1:0] w_n1077_0;
	wire[1:0] w_n1078_0;
	wire[1:0] w_n1080_0;
	wire[1:0] w_n1082_0;
	wire[1:0] w_n1083_0;
	wire[1:0] w_n1084_0;
	wire[1:0] w_n1085_0;
	wire[1:0] w_n1086_0;
	wire[1:0] w_n1087_0;
	wire[1:0] w_n1088_0;
	wire[1:0] w_n1089_0;
	wire[1:0] w_n1090_0;
	wire[1:0] w_n1091_0;
	wire[1:0] w_n1092_0;
	wire[1:0] w_n1093_0;
	wire[1:0] w_n1094_0;
	wire[1:0] w_n1095_0;
	wire[1:0] w_n1096_0;
	wire[1:0] w_n1097_0;
	wire[1:0] w_n1098_0;
	wire[1:0] w_n1099_0;
	wire[1:0] w_n1100_0;
	wire[1:0] w_n1101_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1103_0;
	wire[1:0] w_n1105_0;
	wire[1:0] w_n1106_0;
	wire[1:0] w_n1107_0;
	wire[1:0] w_n1108_0;
	wire[1:0] w_n1109_0;
	wire[1:0] w_n1115_0;
	wire[1:0] w_n1119_0;
	wire[1:0] w_n1120_0;
	wire[1:0] w_n1124_0;
	wire[1:0] w_n1126_0;
	wire[1:0] w_n1129_0;
	wire[1:0] w_n1131_0;
	wire[1:0] w_n1134_0;
	wire[1:0] w_n1136_0;
	wire[1:0] w_n1139_0;
	wire[1:0] w_n1141_0;
	wire[1:0] w_n1144_0;
	wire[1:0] w_n1146_0;
	wire[1:0] w_n1149_0;
	wire[1:0] w_n1151_0;
	wire[1:0] w_n1154_0;
	wire[1:0] w_n1156_0;
	wire[1:0] w_n1159_0;
	wire[1:0] w_n1161_0;
	wire[1:0] w_n1164_0;
	wire[1:0] w_n1166_0;
	wire[1:0] w_n1169_0;
	wire[1:0] w_n1171_0;
	wire[1:0] w_n1174_0;
	wire[1:0] w_n1175_0;
	wire[1:0] w_n1176_0;
	wire[1:0] w_n1179_0;
	wire[1:0] w_n1181_0;
	wire[1:0] w_n1182_0;
	wire[1:0] w_n1183_0;
	wire[1:0] w_n1184_0;
	wire[1:0] w_n1185_0;
	wire[1:0] w_n1186_0;
	wire[1:0] w_n1187_0;
	wire[1:0] w_n1188_0;
	wire[1:0] w_n1189_0;
	wire[1:0] w_n1190_0;
	wire[1:0] w_n1191_0;
	wire[1:0] w_n1192_0;
	wire[1:0] w_n1193_0;
	wire[1:0] w_n1194_0;
	wire[1:0] w_n1195_0;
	wire[1:0] w_n1196_0;
	wire[1:0] w_n1197_0;
	wire[1:0] w_n1198_0;
	wire[1:0] w_n1199_0;
	wire[1:0] w_n1200_0;
	wire[1:0] w_n1201_0;
	wire[1:0] w_n1203_0;
	wire[1:0] w_n1205_0;
	wire[1:0] w_n1206_0;
	wire[1:0] w_n1207_0;
	wire[1:0] w_n1213_0;
	wire[1:0] w_n1216_0;
	wire[1:0] w_n1217_0;
	wire[1:0] w_n1220_0;
	wire[1:0] w_n1222_0;
	wire[1:0] w_n1225_0;
	wire[1:0] w_n1227_0;
	wire[1:0] w_n1230_0;
	wire[1:0] w_n1232_0;
	wire[1:0] w_n1235_0;
	wire[1:0] w_n1237_0;
	wire[1:0] w_n1240_0;
	wire[1:0] w_n1242_0;
	wire[1:0] w_n1245_0;
	wire[1:0] w_n1247_0;
	wire[1:0] w_n1250_0;
	wire[1:0] w_n1252_0;
	wire[1:0] w_n1255_0;
	wire[1:0] w_n1257_0;
	wire[1:0] w_n1260_0;
	wire[1:0] w_n1262_0;
	wire[1:0] w_n1265_0;
	wire[1:0] w_n1266_0;
	wire[1:0] w_n1267_0;
	wire[1:0] w_n1270_0;
	wire[1:0] w_n1272_0;
	wire[1:0] w_n1273_0;
	wire[1:0] w_n1274_0;
	wire[1:0] w_n1275_0;
	wire[1:0] w_n1276_0;
	wire[1:0] w_n1277_0;
	wire[1:0] w_n1278_0;
	wire[1:0] w_n1279_0;
	wire[1:0] w_n1280_0;
	wire[1:0] w_n1281_0;
	wire[1:0] w_n1282_0;
	wire[1:0] w_n1283_0;
	wire[1:0] w_n1284_0;
	wire[1:0] w_n1285_0;
	wire[1:0] w_n1286_0;
	wire[1:0] w_n1287_0;
	wire[1:0] w_n1288_0;
	wire[1:0] w_n1289_0;
	wire[1:0] w_n1290_0;
	wire[1:0] w_n1291_0;
	wire[1:0] w_n1293_0;
	wire[1:0] w_n1294_0;
	wire[1:0] w_n1295_0;
	wire[1:0] w_n1301_0;
	wire[1:0] w_n1306_0;
	wire[1:0] w_n1307_0;
	wire[1:0] w_n1310_0;
	wire[1:0] w_n1312_0;
	wire[1:0] w_n1315_0;
	wire[1:0] w_n1317_0;
	wire[1:0] w_n1320_0;
	wire[1:0] w_n1322_0;
	wire[1:0] w_n1325_0;
	wire[1:0] w_n1327_0;
	wire[1:0] w_n1330_0;
	wire[1:0] w_n1332_0;
	wire[1:0] w_n1335_0;
	wire[1:0] w_n1337_0;
	wire[1:0] w_n1340_0;
	wire[1:0] w_n1342_0;
	wire[1:0] w_n1345_0;
	wire[1:0] w_n1347_0;
	wire[1:0] w_n1350_0;
	wire[1:0] w_n1351_0;
	wire[1:0] w_n1352_0;
	wire[1:0] w_n1355_0;
	wire[1:0] w_n1357_0;
	wire[1:0] w_n1358_0;
	wire[1:0] w_n1359_0;
	wire[1:0] w_n1360_0;
	wire[1:0] w_n1361_0;
	wire[1:0] w_n1362_0;
	wire[1:0] w_n1363_0;
	wire[1:0] w_n1364_0;
	wire[1:0] w_n1365_0;
	wire[1:0] w_n1366_0;
	wire[1:0] w_n1367_0;
	wire[1:0] w_n1368_0;
	wire[1:0] w_n1369_0;
	wire[1:0] w_n1370_0;
	wire[1:0] w_n1371_0;
	wire[1:0] w_n1372_0;
	wire[1:0] w_n1373_0;
	wire[1:0] w_n1374_0;
	wire[1:0] w_n1376_0;
	wire[1:0] w_n1378_0;
	wire[1:0] w_n1379_0;
	wire[1:0] w_n1384_0;
	wire[1:0] w_n1389_0;
	wire[1:0] w_n1390_0;
	wire[1:0] w_n1393_0;
	wire[1:0] w_n1395_0;
	wire[1:0] w_n1398_0;
	wire[1:0] w_n1400_0;
	wire[1:0] w_n1403_0;
	wire[1:0] w_n1405_0;
	wire[1:0] w_n1408_0;
	wire[1:0] w_n1410_0;
	wire[1:0] w_n1413_0;
	wire[1:0] w_n1415_0;
	wire[1:0] w_n1418_0;
	wire[1:0] w_n1420_0;
	wire[1:0] w_n1423_0;
	wire[1:0] w_n1425_0;
	wire[1:0] w_n1428_0;
	wire[1:0] w_n1429_0;
	wire[1:0] w_n1430_0;
	wire[1:0] w_n1433_0;
	wire[1:0] w_n1435_0;
	wire[1:0] w_n1436_0;
	wire[1:0] w_n1437_0;
	wire[1:0] w_n1438_0;
	wire[1:0] w_n1439_0;
	wire[1:0] w_n1440_0;
	wire[1:0] w_n1441_0;
	wire[1:0] w_n1442_0;
	wire[1:0] w_n1443_0;
	wire[1:0] w_n1444_0;
	wire[1:0] w_n1445_0;
	wire[1:0] w_n1446_0;
	wire[1:0] w_n1447_0;
	wire[1:0] w_n1448_0;
	wire[1:0] w_n1449_0;
	wire[1:0] w_n1450_0;
	wire[1:0] w_n1452_0;
	wire[1:0] w_n1454_0;
	wire[1:0] w_n1455_0;
	wire[1:0] w_n1460_0;
	wire[1:0] w_n1465_0;
	wire[1:0] w_n1466_0;
	wire[1:0] w_n1469_0;
	wire[1:0] w_n1471_0;
	wire[1:0] w_n1474_0;
	wire[1:0] w_n1476_0;
	wire[1:0] w_n1479_0;
	wire[1:0] w_n1481_0;
	wire[1:0] w_n1484_0;
	wire[1:0] w_n1486_0;
	wire[1:0] w_n1489_0;
	wire[1:0] w_n1491_0;
	wire[1:0] w_n1494_0;
	wire[1:0] w_n1496_0;
	wire[1:0] w_n1499_0;
	wire[1:0] w_n1500_0;
	wire[1:0] w_n1501_0;
	wire[1:0] w_n1504_0;
	wire[1:0] w_n1506_0;
	wire[1:0] w_n1507_0;
	wire[1:0] w_n1508_0;
	wire[1:0] w_n1509_0;
	wire[1:0] w_n1510_0;
	wire[1:0] w_n1511_0;
	wire[1:0] w_n1512_0;
	wire[1:0] w_n1513_0;
	wire[1:0] w_n1514_0;
	wire[1:0] w_n1515_0;
	wire[1:0] w_n1516_0;
	wire[1:0] w_n1517_0;
	wire[1:0] w_n1518_0;
	wire[1:0] w_n1519_0;
	wire[1:0] w_n1521_0;
	wire[1:0] w_n1523_0;
	wire[1:0] w_n1524_0;
	wire[1:0] w_n1529_0;
	wire[1:0] w_n1534_0;
	wire[1:0] w_n1535_0;
	wire[1:0] w_n1538_0;
	wire[1:0] w_n1540_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1545_0;
	wire[1:0] w_n1548_0;
	wire[1:0] w_n1550_0;
	wire[1:0] w_n1553_0;
	wire[1:0] w_n1555_0;
	wire[1:0] w_n1558_0;
	wire[1:0] w_n1560_0;
	wire[1:0] w_n1563_0;
	wire[1:0] w_n1564_0;
	wire[1:0] w_n1565_0;
	wire[1:0] w_n1568_0;
	wire[1:0] w_n1570_0;
	wire[1:0] w_n1571_0;
	wire[1:0] w_n1572_0;
	wire[1:0] w_n1573_0;
	wire[1:0] w_n1574_0;
	wire[1:0] w_n1575_0;
	wire[1:0] w_n1576_0;
	wire[1:0] w_n1577_0;
	wire[1:0] w_n1578_0;
	wire[1:0] w_n1579_0;
	wire[1:0] w_n1580_0;
	wire[1:0] w_n1581_0;
	wire[1:0] w_n1583_0;
	wire[1:0] w_n1585_0;
	wire[1:0] w_n1586_0;
	wire[1:0] w_n1591_0;
	wire[1:0] w_n1596_0;
	wire[1:0] w_n1597_0;
	wire[1:0] w_n1600_0;
	wire[1:0] w_n1602_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1607_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1612_0;
	wire[1:0] w_n1615_0;
	wire[1:0] w_n1617_0;
	wire[1:0] w_n1620_0;
	wire[1:0] w_n1621_0;
	wire[1:0] w_n1622_0;
	wire[1:0] w_n1625_0;
	wire[1:0] w_n1627_0;
	wire[1:0] w_n1628_0;
	wire[1:0] w_n1629_0;
	wire[1:0] w_n1630_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1632_0;
	wire[1:0] w_n1633_0;
	wire[1:0] w_n1634_0;
	wire[1:0] w_n1635_0;
	wire[1:0] w_n1636_0;
	wire[1:0] w_n1638_0;
	wire[1:0] w_n1640_0;
	wire[1:0] w_n1641_0;
	wire[1:0] w_n1646_0;
	wire[1:0] w_n1651_0;
	wire[1:0] w_n1653_0;
	wire[1:0] w_n1656_0;
	wire[1:0] w_n1658_0;
	wire[1:0] w_n1661_0;
	wire[1:0] w_n1663_0;
	wire[1:0] w_n1666_0;
	wire[1:0] w_n1668_0;
	wire[1:0] w_n1671_0;
	wire[1:0] w_n1672_0;
	wire[1:0] w_n1673_0;
	wire[1:0] w_n1676_0;
	wire[1:0] w_n1678_0;
	wire[1:0] w_n1679_0;
	wire[1:0] w_n1680_0;
	wire[1:0] w_n1681_0;
	wire[1:0] w_n1682_0;
	wire[1:0] w_n1683_0;
	wire[1:0] w_n1684_0;
	wire[1:0] w_n1685_0;
	wire[1:0] w_n1686_0;
	wire[1:0] w_n1688_0;
	wire[1:0] w_n1689_0;
	wire[1:0] w_n1694_0;
	wire[1:0] w_n1697_0;
	wire[1:0] w_n1699_0;
	wire[1:0] w_n1702_0;
	wire[1:0] w_n1704_0;
	wire[1:0] w_n1707_0;
	wire[1:0] w_n1709_0;
	wire[1:0] w_n1712_0;
	wire[1:0] w_n1713_0;
	wire[1:0] w_n1714_0;
	wire[1:0] w_n1717_0;
	wire[1:0] w_n1719_0;
	wire[1:0] w_n1720_0;
	wire[1:0] w_n1721_0;
	wire[1:0] w_n1722_0;
	wire[1:0] w_n1723_0;
	wire[1:0] w_n1724_0;
	wire[1:0] w_n1725_0;
	wire[1:0] w_n1726_0;
	wire[1:0] w_n1727_0;
	wire[1:0] w_n1734_0;
	wire[1:0] w_n1737_0;
	wire[1:0] w_n1739_0;
	wire[1:0] w_n1742_0;
	wire[1:0] w_n1744_0;
	wire[1:0] w_n1747_0;
	wire[1:0] w_n1748_0;
	wire[1:0] w_n1749_0;
	wire[1:0] w_n1752_0;
	wire[1:0] w_n1754_0;
	wire[1:0] w_n1755_0;
	wire[1:0] w_n1756_0;
	wire[1:0] w_n1757_0;
	wire[1:0] w_n1758_0;
	wire[1:0] w_n1759_0;
	wire[1:0] w_n1760_0;
	wire[1:0] w_n1767_0;
	wire[1:0] w_n1770_0;
	wire[1:0] w_n1772_0;
	wire[1:0] w_n1775_0;
	wire[1:0] w_n1776_0;
	wire[1:0] w_n1777_0;
	wire[1:0] w_n1780_0;
	wire[1:0] w_n1782_0;
	wire[1:0] w_n1783_0;
	wire[1:0] w_n1784_0;
	wire[1:0] w_n1785_0;
	wire[1:0] w_n1786_0;
	wire[1:0] w_n1793_0;
	wire[1:0] w_n1796_0;
	wire[1:0] w_n1797_0;
	wire[1:0] w_n1798_0;
	wire[1:0] w_n1801_0;
	wire[1:0] w_n1803_0;
	wire[1:0] w_n1804_0;
	wire[1:0] w_n1805_0;
	wire[1:0] w_n1807_0;
	wire[1:0] w_n1810_0;
	wire[1:0] w_n1817_0;
	wire[1:0] w_n1818_0;
	wire w_dff_B_DmmoZnUj4_1;
	wire w_dff_B_O5UfwTMy7_1;
	wire w_dff_B_8vD6sN1d2_1;
	wire w_dff_B_Hiz3iM2k5_1;
	wire w_dff_B_m1Ii7war6_1;
	wire w_dff_B_hYO5RUoD3_1;
	wire w_dff_B_Hwgr4myO5_1;
	wire w_dff_B_qNxmAhNK9_1;
	wire w_dff_B_VEfEsqjZ4_1;
	wire w_dff_B_8KXu2Zag5_1;
	wire w_dff_B_uIY1MvCi2_1;
	wire w_dff_B_G16ejBdK8_1;
	wire w_dff_B_Njl0MimF5_1;
	wire w_dff_B_DdDQfMAb4_1;
	wire w_dff_B_08DDgJsb9_1;
	wire w_dff_B_6YBjp3va1_1;
	wire w_dff_B_pl8hv5cK9_1;
	wire w_dff_B_QGLP9ZNw7_1;
	wire w_dff_B_k6vZhay37_1;
	wire w_dff_B_PXqvL3oF9_1;
	wire w_dff_B_m525AQQ50_1;
	wire w_dff_B_nsx5O4Gl8_1;
	wire w_dff_B_Dw3YggC90_1;
	wire w_dff_B_oJoOm4SQ7_1;
	wire w_dff_B_LnvdU34o4_1;
	wire w_dff_B_6LbTY0Pz3_1;
	wire w_dff_B_uLNTgwOp2_1;
	wire w_dff_B_gwscHMSo7_1;
	wire w_dff_B_hMbcC3mw6_1;
	wire w_dff_B_zKlZiXNS1_1;
	wire w_dff_B_AnSItq1I2_1;
	wire w_dff_B_yjgmjPdQ9_1;
	wire w_dff_B_SdH9pkK08_1;
	wire w_dff_B_Ngrtt6ca2_1;
	wire w_dff_B_VMrmjhAN3_1;
	wire w_dff_B_gzsugydL4_1;
	wire w_dff_B_3T1e59ex9_1;
	wire w_dff_B_biLnVCNd4_1;
	wire w_dff_B_Z3eSmBT88_1;
	wire w_dff_B_hbLGiVVl0_1;
	wire w_dff_B_Oj9lc4aV7_1;
	wire w_dff_B_zo2drDBd7_1;
	wire w_dff_B_ouqWyAAx4_1;
	wire w_dff_B_v0WLDwnZ3_1;
	wire w_dff_B_GF8o5Vdy5_1;
	wire w_dff_B_iujrpnet2_1;
	wire w_dff_B_eJp8CXws4_1;
	wire w_dff_B_KgmnRMDg9_1;
	wire w_dff_B_4maCP0DT9_1;
	wire w_dff_B_fD0zaANk0_1;
	wire w_dff_B_frvYvEMt1_1;
	wire w_dff_B_C8DKEqdO0_1;
	wire w_dff_B_auOkeWc03_1;
	wire w_dff_B_ClUzhLj95_1;
	wire w_dff_B_pbZBQBQ81_1;
	wire w_dff_B_w5UJ3Hr82_1;
	wire w_dff_B_lzMtvHSY7_1;
	wire w_dff_B_3Uw4ZDel3_1;
	wire w_dff_B_IJvDkFa97_1;
	wire w_dff_B_GeJ4GHtm9_1;
	wire w_dff_B_n3OKOcXa8_1;
	wire w_dff_B_MHon3vc79_1;
	wire w_dff_B_789OLFB94_1;
	wire w_dff_B_b5QkdwGE9_1;
	wire w_dff_B_WAFfsglX3_1;
	wire w_dff_B_erwi466O1_1;
	wire w_dff_B_BWUk9T503_1;
	wire w_dff_B_riPkWCzu2_1;
	wire w_dff_B_TvYmVkVV7_1;
	wire w_dff_B_WSehINEJ4_1;
	wire w_dff_B_lKdWkEuU0_1;
	wire w_dff_B_YdG3jBos4_1;
	wire w_dff_B_iHggrrry0_1;
	wire w_dff_B_QQRsESRT6_1;
	wire w_dff_B_4nhTHUpg6_1;
	wire w_dff_B_jLRJMcJm6_1;
	wire w_dff_B_vF4XRc2B8_1;
	wire w_dff_B_2LLpG0Jk0_1;
	wire w_dff_B_xVKTvnKl8_1;
	wire w_dff_B_PtGgImiU4_1;
	wire w_dff_B_gXr6bPCJ7_1;
	wire w_dff_B_om5bBsvF4_1;
	wire w_dff_B_NsSxQTMb8_1;
	wire w_dff_B_fQ9WsX7z0_1;
	wire w_dff_B_01aOoW4c3_1;
	wire w_dff_B_IcpXjXpr1_1;
	wire w_dff_B_uZk2Emv61_1;
	wire w_dff_B_WoJNcMIQ1_1;
	wire w_dff_B_sgClU7AO7_1;
	wire w_dff_B_VPgk4d3B3_1;
	wire w_dff_B_l9WwO8Mz0_1;
	wire w_dff_B_oREOLxlD2_1;
	wire w_dff_B_Te1RunYj8_1;
	wire w_dff_B_MYxqiZYm4_1;
	wire w_dff_B_vBaHb8ij5_1;
	wire w_dff_B_HMSZy4Na2_1;
	wire w_dff_B_rwXOrWtG3_1;
	wire w_dff_B_T5SjFso25_1;
	wire w_dff_B_HdcJeoIO2_1;
	wire w_dff_B_VJtWhcZw1_1;
	wire w_dff_B_vzUVOpRP1_1;
	wire w_dff_B_PI3sUmll9_1;
	wire w_dff_B_P66p3rJ67_1;
	wire w_dff_B_MBRCpfmD5_1;
	wire w_dff_B_CiTjA84y9_1;
	wire w_dff_B_nun1b87I5_1;
	wire w_dff_B_SW6JTjmV5_1;
	wire w_dff_B_OHdJphC50_1;
	wire w_dff_B_E8fcmvup6_1;
	wire w_dff_B_E1nNgb8c2_1;
	wire w_dff_B_Bwgm8y2A6_1;
	wire w_dff_B_7S89rXFQ7_1;
	wire w_dff_B_iP6K61Sy2_1;
	wire w_dff_B_IF1kwRy05_1;
	wire w_dff_B_nG835zYk3_1;
	wire w_dff_B_YEgrd9ZL2_1;
	wire w_dff_B_fQSDUVuy2_1;
	wire w_dff_B_mmhX7XXn8_1;
	wire w_dff_B_S8LpbVQ87_1;
	wire w_dff_B_qnXRm3zS1_1;
	wire w_dff_B_QO6Z7H856_1;
	wire w_dff_B_8ZqH8pFz4_1;
	wire w_dff_B_jSivffm70_1;
	wire w_dff_B_yQQkW4Fa4_1;
	wire w_dff_B_JSeegWP58_1;
	wire w_dff_B_4yHvPCnb6_1;
	wire w_dff_B_RD7qAJwj2_1;
	wire w_dff_B_3TJDN0bk5_1;
	wire w_dff_B_0Qj6UhC57_1;
	wire w_dff_B_yGi0Wq9I4_1;
	wire w_dff_B_lOMoAspd9_1;
	wire w_dff_B_OySdTCav3_1;
	wire w_dff_B_g7bMOlFS4_1;
	wire w_dff_B_eL0bZyCn8_1;
	wire w_dff_B_1wTyjv7c3_1;
	wire w_dff_B_TfdwRd9M2_1;
	wire w_dff_B_1M7MlyqW0_1;
	wire w_dff_B_AwPOeHeQ5_1;
	wire w_dff_B_C2TYHHhe3_1;
	wire w_dff_B_Pj8V49Ek7_1;
	wire w_dff_B_3gJ76Ugx7_1;
	wire w_dff_B_Dbp9Iwf30_1;
	wire w_dff_B_tTTHKu3d4_1;
	wire w_dff_B_Itb1kBIT1_1;
	wire w_dff_B_g54LDIIB1_1;
	wire w_dff_B_Mzb6AKu96_1;
	wire w_dff_B_VcHvAqnl4_1;
	wire w_dff_B_NGjKnrUm7_1;
	wire w_dff_B_Tip0e28S9_1;
	wire w_dff_B_4ajDorjz4_1;
	wire w_dff_B_itTf6Q6w9_1;
	wire w_dff_B_Kx8XthuG6_1;
	wire w_dff_B_DrkKKcom5_1;
	wire w_dff_B_nzagnWGq2_1;
	wire w_dff_B_VXFgWWg23_1;
	wire w_dff_B_7vxnz7iE1_1;
	wire w_dff_B_GMLGlu8i1_1;
	wire w_dff_B_UFxdavHd9_1;
	wire w_dff_B_4QdrHxkM0_1;
	wire w_dff_B_d8Cvow7m9_1;
	wire w_dff_B_NgFZ1CPf8_1;
	wire w_dff_B_9G4RZfFC1_1;
	wire w_dff_B_SPh3Sak03_1;
	wire w_dff_B_Igyd8ruU9_1;
	wire w_dff_B_fjZoUprZ9_1;
	wire w_dff_B_Txky5zgy7_1;
	wire w_dff_B_k3FqqkVZ2_1;
	wire w_dff_B_J8ximAF64_1;
	wire w_dff_B_GpjNY5Oc5_1;
	wire w_dff_B_p4YATAlO1_1;
	wire w_dff_B_JiuUQjQD1_1;
	wire w_dff_B_zmFQ6Vpz1_1;
	wire w_dff_B_m5V3H9j18_1;
	wire w_dff_B_qWr93fEV4_1;
	wire w_dff_B_uHy60XbG0_1;
	wire w_dff_B_XUZEOL9G6_1;
	wire w_dff_B_8oyR6nEv8_1;
	wire w_dff_B_6PbOU3cd5_1;
	wire w_dff_B_uVd8zuOI9_1;
	wire w_dff_B_6bLfUHjx3_1;
	wire w_dff_B_kzudbABd2_1;
	wire w_dff_B_Q4jqvAR08_1;
	wire w_dff_B_W7TQf5g40_1;
	wire w_dff_B_Q72cJvuh4_1;
	wire w_dff_B_HbUHzykR5_1;
	wire w_dff_B_bdbcuCYw0_1;
	wire w_dff_B_watOFMiZ3_1;
	wire w_dff_B_wQVy7xhE5_1;
	wire w_dff_B_mF1QKGRy0_1;
	wire w_dff_B_1yUxJ1x12_1;
	wire w_dff_B_OFUJJxNn0_1;
	wire w_dff_B_6heiRbpb6_1;
	wire w_dff_B_BJJQTFvw0_1;
	wire w_dff_B_ZtoLuE4X5_1;
	wire w_dff_B_wYmjdvKH0_1;
	wire w_dff_B_U6UQxXkn3_1;
	wire w_dff_B_gr5e1xZr5_1;
	wire w_dff_B_r1iAy6MU3_1;
	wire w_dff_B_1QC1TQcj0_1;
	wire w_dff_B_2Md8l1sc6_1;
	wire w_dff_B_cKCw7bBK8_1;
	wire w_dff_B_GEJAlnEN5_1;
	wire w_dff_B_ek1jnSIg9_1;
	wire w_dff_B_YJIGeZAa9_1;
	wire w_dff_B_067TIfkz4_1;
	wire w_dff_B_48s9u1u96_1;
	wire w_dff_B_smNr4rDx2_1;
	wire w_dff_B_Em3nZ4jE4_1;
	wire w_dff_B_1I3uuWz87_1;
	wire w_dff_B_xt1bLtH50_1;
	wire w_dff_B_xdulWiE02_1;
	wire w_dff_B_QkcW4NYo0_1;
	wire w_dff_B_6lLVEvrx1_1;
	wire w_dff_B_xi943vMI6_1;
	wire w_dff_B_4iijnvTh3_1;
	wire w_dff_B_pfonSuJY5_1;
	wire w_dff_B_8BWcsDFe7_1;
	wire w_dff_B_mNNeMzGq2_1;
	wire w_dff_B_uZ9pkRDC2_1;
	wire w_dff_B_mbf7GveI3_1;
	wire w_dff_B_oScKx5Wf6_1;
	wire w_dff_B_4AsiEg0h4_1;
	wire w_dff_B_DVKnjaKG7_1;
	wire w_dff_B_aUekxOjk4_1;
	wire w_dff_B_jXgKvv612_1;
	wire w_dff_B_r6dfayWB3_1;
	wire w_dff_B_X2Jw8EXg6_1;
	wire w_dff_B_A46QaqN33_1;
	wire w_dff_B_Yx74BAga0_1;
	wire w_dff_B_P01OHjIW8_1;
	wire w_dff_B_4CgSfogD6_1;
	wire w_dff_B_WVCSxjUL1_1;
	wire w_dff_B_5qykt55W7_1;
	wire w_dff_B_Vb5ZFRw32_1;
	wire w_dff_B_k4jAsaKo7_1;
	wire w_dff_B_wpllafUx6_1;
	wire w_dff_B_EjYO7dmp8_1;
	wire w_dff_B_cxNaOFz90_1;
	wire w_dff_B_LYsPiCCA0_1;
	wire w_dff_B_xEiGVe7T2_1;
	wire w_dff_B_PmTPMPTs1_1;
	wire w_dff_B_gT3iJnmn0_1;
	wire w_dff_B_QpUILwRe9_1;
	wire w_dff_B_ehNSmuTL9_1;
	wire w_dff_B_9mU3c2q68_1;
	wire w_dff_B_zDrUJLFD3_1;
	wire w_dff_B_Uz5pXQIO1_1;
	wire w_dff_B_ZEtmJWfV7_1;
	wire w_dff_B_HmSXNsVh9_1;
	wire w_dff_B_mBI9FvqX1_1;
	wire w_dff_B_ojzThOHR2_1;
	wire w_dff_B_Q89DwB954_1;
	wire w_dff_B_Su6VguAg8_1;
	wire w_dff_B_0sUkPOSg7_1;
	wire w_dff_B_s0C5wQSf5_1;
	wire w_dff_B_sh8vrTxC4_1;
	wire w_dff_B_NFykJsdv1_1;
	wire w_dff_B_ms9B5Xkn0_1;
	wire w_dff_B_8LtNSkZM8_1;
	wire w_dff_B_Yp1W0ap52_1;
	wire w_dff_B_S0jgYNTv2_1;
	wire w_dff_B_IMlnEWuK7_1;
	wire w_dff_B_SafHHuqU4_1;
	wire w_dff_B_onCF08pC7_1;
	wire w_dff_B_tYhpkpMf6_1;
	wire w_dff_B_YSNgH7gA4_1;
	wire w_dff_B_0xOmQsRi1_1;
	wire w_dff_B_ZVn2BZEI0_1;
	wire w_dff_B_xKtPHTX48_1;
	wire w_dff_B_XZmhVAb25_1;
	wire w_dff_B_0Dv6C3xd8_1;
	wire w_dff_B_H12TUS8Q4_1;
	wire w_dff_B_khjF5Lua6_1;
	wire w_dff_B_OCgX8gW97_1;
	wire w_dff_B_G0f4VCiM3_1;
	wire w_dff_B_Ay1LnXh60_1;
	wire w_dff_B_eeV9nUrs1_1;
	wire w_dff_B_JQsVcHQJ0_1;
	wire w_dff_B_odtFOmT87_1;
	wire w_dff_B_eKMZstAZ6_1;
	wire w_dff_B_gqklguIX4_1;
	wire w_dff_B_pgUahyWQ2_1;
	wire w_dff_B_PIYxYIMU9_1;
	wire w_dff_B_MCDpiy712_1;
	wire w_dff_B_DbLOSDb16_1;
	wire w_dff_B_uQRAheUd0_1;
	wire w_dff_B_8VoKSApJ7_1;
	wire w_dff_B_s4ffzqGG3_1;
	wire w_dff_B_cSoUArzT0_1;
	wire w_dff_B_tnBYqjOd5_1;
	wire w_dff_B_IoUnQinS4_1;
	wire w_dff_B_2OxD9q6H5_1;
	wire w_dff_B_GaWogtCT2_1;
	wire w_dff_B_n5JMJ61k0_1;
	wire w_dff_B_Cs2OmUco5_1;
	wire w_dff_B_wdxefOFN0_1;
	wire w_dff_B_EFjaSjHT7_1;
	wire w_dff_B_2hZlOMVi8_1;
	wire w_dff_B_QRhjZZyp0_1;
	wire w_dff_B_lUE2hNpe3_1;
	wire w_dff_B_V2SsRoJB9_1;
	wire w_dff_B_0HyguaWJ1_1;
	wire w_dff_B_j7rUtNQ01_1;
	wire w_dff_B_UH7q5hBH3_1;
	wire w_dff_B_9PjiUSgH4_1;
	wire w_dff_B_sP81te7Z0_1;
	wire w_dff_B_Qm2w4L9n6_1;
	wire w_dff_B_NxbTxvB99_1;
	wire w_dff_B_p8VCotCh1_1;
	wire w_dff_B_pki0VitO5_1;
	wire w_dff_B_XxB3sXCL9_1;
	wire w_dff_B_OSzEtGV39_1;
	wire w_dff_B_VFotRj8h7_1;
	wire w_dff_B_6LtDBr7p7_1;
	wire w_dff_B_jf1zmcsS5_1;
	wire w_dff_B_A72U7TVO7_0;
	wire w_dff_B_2bXHW5pD2_1;
	wire w_dff_B_combaM0x6_1;
	wire w_dff_B_WJlDsVAg4_1;
	wire w_dff_B_6hfngCDd5_1;
	wire w_dff_B_Whl6dzRx7_1;
	wire w_dff_B_fowZhe165_1;
	wire w_dff_B_tn22G5N56_1;
	wire w_dff_B_5GRs5Cqd8_1;
	wire w_dff_B_Q9aBr6lV2_1;
	wire w_dff_B_PY7RO6Vt7_1;
	wire w_dff_B_Fo5D8mPH4_1;
	wire w_dff_B_amOp1eBC0_1;
	wire w_dff_B_uGmmzoV76_1;
	wire w_dff_B_8WpZYETE2_1;
	wire w_dff_B_I6ALDGFU2_1;
	wire w_dff_B_UODfp17m5_0;
	wire w_dff_B_C2fgywuC4_0;
	wire w_dff_B_iSNLeOj13_0;
	wire w_dff_B_ubllVIKr1_0;
	wire w_dff_B_sSHGz87U4_0;
	wire w_dff_B_WosEgbB53_0;
	wire w_dff_B_AA7GTO5r1_0;
	wire w_dff_B_F6O6CMhn6_0;
	wire w_dff_B_NDvo4c0r1_0;
	wire w_dff_B_28455s062_0;
	wire w_dff_B_rI9ZnYwA1_0;
	wire w_dff_B_hcUrSKa20_0;
	wire w_dff_B_7IAlXGz98_0;
	wire w_dff_B_vB92Z3wd0_1;
	wire w_dff_B_1z2SjFgn6_1;
	wire w_dff_B_s7f3VCWp9_1;
	wire w_dff_B_6f5bYo4b0_1;
	wire w_dff_B_sMYlibVf4_1;
	wire w_dff_B_y2bLOyBS9_1;
	wire w_dff_B_Ag21fRFK7_1;
	wire w_dff_B_NU2rreoE3_1;
	wire w_dff_B_20SpjbN58_1;
	wire w_dff_B_ni4MjmfM3_1;
	wire w_dff_B_U4FBYWht0_1;
	wire w_dff_B_6cBDMDFk1_1;
	wire w_dff_B_5v4CRyGD2_1;
	wire w_dff_B_C0lRgFtL6_0;
	wire w_dff_B_FaXRMAPW6_0;
	wire w_dff_B_bcklkbUS0_0;
	wire w_dff_B_OWWRXFVB1_0;
	wire w_dff_B_vFzvKk599_0;
	wire w_dff_B_wH2V0pic6_0;
	wire w_dff_B_KuaPtgtw3_0;
	wire w_dff_B_zcGSBZpn3_0;
	wire w_dff_B_yBE6hfya7_0;
	wire w_dff_B_QOyXFxXb1_0;
	wire w_dff_B_FTiyY0mW7_0;
	wire w_dff_B_MdmJGBM98_0;
	wire w_dff_B_l53WllE26_1;
	wire w_dff_B_vSbNmNzd5_1;
	wire w_dff_B_Mg9kBZZz1_1;
	wire w_dff_B_LiTXwJ6Q6_1;
	wire w_dff_B_PS8G7aWC1_1;
	wire w_dff_B_GZDCKJP06_1;
	wire w_dff_B_HNn22smk6_1;
	wire w_dff_B_pr6TljLb6_1;
	wire w_dff_B_5idRKmw72_1;
	wire w_dff_B_rc0gTyTh5_1;
	wire w_dff_B_tjpf42O52_1;
	wire w_dff_B_yk1vio3G0_1;
	wire w_dff_B_rfh8Azrx4_1;
	wire w_dff_B_DsiobYQn1_0;
	wire w_dff_B_YFdZIHOs6_0;
	wire w_dff_B_Zz9muBOd2_0;
	wire w_dff_B_4VYOsYnj6_0;
	wire w_dff_B_xaGkl7932_0;
	wire w_dff_B_ASUAg8o84_0;
	wire w_dff_B_HbqTf5TA5_0;
	wire w_dff_B_MnRayzoh5_0;
	wire w_dff_B_8EJkcAz10_0;
	wire w_dff_B_pWrvYSR92_0;
	wire w_dff_B_LaxHBH1F4_0;
	wire w_dff_B_zeHvFZoO8_0;
	wire w_dff_B_4rUrdJut2_1;
	wire w_dff_B_lSHDL41o8_1;
	wire w_dff_B_QVMOXoxm0_1;
	wire w_dff_B_wlaFYO1W2_1;
	wire w_dff_B_lLOn836r2_1;
	wire w_dff_B_i8CPTuLt7_1;
	wire w_dff_B_mNepDa3v0_1;
	wire w_dff_B_S3zaJXXc4_1;
	wire w_dff_B_Kv8ad9017_1;
	wire w_dff_B_u6KVBQwU1_1;
	wire w_dff_B_ikSOyS6r2_1;
	wire w_dff_B_Ywy5LDQw3_1;
	wire w_dff_B_cJe6CABx7_1;
	wire w_dff_B_uxFLB0it2_0;
	wire w_dff_B_j6bHU2QJ2_0;
	wire w_dff_B_RngWOTVA7_0;
	wire w_dff_B_CnngvG7H5_0;
	wire w_dff_B_CKE3EUF77_0;
	wire w_dff_B_55bo053C8_0;
	wire w_dff_B_AhNbvZ8F3_0;
	wire w_dff_B_l6tCg6yp8_0;
	wire w_dff_B_dFb3QVSD8_0;
	wire w_dff_B_uPqkqIb35_0;
	wire w_dff_B_q6KGRDOl4_0;
	wire w_dff_B_mlOdPv2S6_0;
	wire w_dff_B_xQCfkq6P2_1;
	wire w_dff_B_Gd4kUgaV9_1;
	wire w_dff_B_JjlNcBPv4_1;
	wire w_dff_B_bnx65bnW8_1;
	wire w_dff_B_wPSp4Poz7_1;
	wire w_dff_B_2l9hHGLC4_1;
	wire w_dff_B_k59GZeqv6_1;
	wire w_dff_B_6dnsRt8p2_1;
	wire w_dff_B_CXNy6fxz4_1;
	wire w_dff_B_ecas7eyI4_1;
	wire w_dff_B_PiU4xhR46_1;
	wire w_dff_B_SjMI8q2N3_1;
	wire w_dff_B_IZ4uEvw22_1;
	wire w_dff_B_yOdNxUpG8_0;
	wire w_dff_B_Ppaiyd0W7_0;
	wire w_dff_B_IIittGiD5_0;
	wire w_dff_B_RtQgXSsh1_0;
	wire w_dff_B_PciOO2LB1_0;
	wire w_dff_B_XsEugE3H9_0;
	wire w_dff_B_u1aeVSYb5_0;
	wire w_dff_B_Gz3MZsGO2_0;
	wire w_dff_B_GCobDsPT1_0;
	wire w_dff_B_jSkAOPfq3_0;
	wire w_dff_B_Am9jWcao0_0;
	wire w_dff_B_H4gx2No93_0;
	wire w_dff_B_XS0v6Yt94_1;
	wire w_dff_B_GzJukZws6_1;
	wire w_dff_B_SKcAnUJJ3_1;
	wire w_dff_B_nm6Woswp3_1;
	wire w_dff_B_IJgyw2lz5_1;
	wire w_dff_B_z14zVm0B2_1;
	wire w_dff_B_M8MFXSHL3_1;
	wire w_dff_B_SdVSy13N0_1;
	wire w_dff_B_AjupddhC6_1;
	wire w_dff_B_sCIEwXn17_1;
	wire w_dff_B_qadIgar63_1;
	wire w_dff_B_hrXwnM7u2_1;
	wire w_dff_B_FLzv5IFQ9_1;
	wire w_dff_B_AgH5C2HU5_0;
	wire w_dff_B_VSK6eRX65_0;
	wire w_dff_B_PqqA8cXq1_0;
	wire w_dff_B_SxAIVMtE8_0;
	wire w_dff_B_ZkV6EUFj9_0;
	wire w_dff_B_dAL4109h5_0;
	wire w_dff_B_emvDU7qz9_0;
	wire w_dff_B_Ci4zxg9i2_0;
	wire w_dff_B_NGl4n9je9_0;
	wire w_dff_B_49MfWjRv3_0;
	wire w_dff_B_XtoT0os52_0;
	wire w_dff_B_JYhckuGj9_1;
	wire w_dff_B_gNJ52H7k6_1;
	wire w_dff_B_QXGLSJiU0_1;
	wire w_dff_B_bmazQtKw7_1;
	wire w_dff_B_fvfPc0Y45_1;
	wire w_dff_B_rjErD65m3_1;
	wire w_dff_B_8C34pXR15_1;
	wire w_dff_B_60U9NIXZ2_1;
	wire w_dff_B_H8AGPWpd5_1;
	wire w_dff_B_IvcX5JtQ3_1;
	wire w_dff_B_ULhVCJZl1_1;
	wire w_dff_B_eDg4Wggn8_1;
	wire w_dff_B_i2yFD3pf6_0;
	wire w_dff_B_7bztS9jn8_0;
	wire w_dff_B_s0XxKT3p5_0;
	wire w_dff_B_Jx8nqwLq8_0;
	wire w_dff_B_mMJxiULn5_0;
	wire w_dff_B_XSrf3GsQ8_0;
	wire w_dff_B_LUQpthNW2_0;
	wire w_dff_B_fE3mV4bG3_0;
	wire w_dff_B_NyfWoSAF9_0;
	wire w_dff_B_17qFCh4f9_0;
	wire w_dff_B_ho1dLcXQ7_1;
	wire w_dff_B_MW0GOehu6_1;
	wire w_dff_B_d3imbFOs7_1;
	wire w_dff_B_DaYm668r7_1;
	wire w_dff_B_E99CDv9F1_1;
	wire w_dff_B_5YzPwp3N2_1;
	wire w_dff_B_UBvpm76y9_1;
	wire w_dff_B_OB4agIAn7_1;
	wire w_dff_B_lEQH5B4y9_1;
	wire w_dff_B_PekFeIzl8_1;
	wire w_dff_B_ROPNhEJH1_0;
	wire w_dff_B_v4FDHYhU7_0;
	wire w_dff_B_N9lZE66c9_0;
	wire w_dff_B_MlYzs8A12_0;
	wire w_dff_B_ot9XZPI12_0;
	wire w_dff_B_f32xVb5V9_0;
	wire w_dff_B_7d48Z0JU4_0;
	wire w_dff_B_BRq9R90W5_0;
	wire w_dff_B_0MOqRX8r1_1;
	wire w_dff_B_X3n6zlmJ0_1;
	wire w_dff_B_LHaoAXLB5_1;
	wire w_dff_B_Pi3L4iFl2_1;
	wire w_dff_B_u4MGejJa1_1;
	wire w_dff_B_EmbF5t6s7_1;
	wire w_dff_B_6zS7mczk2_1;
	wire w_dff_B_6XWUy8nb8_1;
	wire w_dff_B_4zhX4x6F4_0;
	wire w_dff_B_M4jVcfQi7_0;
	wire w_dff_B_PTz5t4lN2_0;
	wire w_dff_B_MS37GiVH4_0;
	wire w_dff_B_GptzSQq79_0;
	wire w_dff_B_tPp8Fugc9_0;
	wire w_dff_B_KllwmgZA0_1;
	wire w_dff_B_dw11LbjA5_1;
	wire w_dff_B_plwNbacf8_1;
	wire w_dff_B_onyABVuW4_1;
	wire w_dff_B_mmNgvumf7_1;
	wire w_dff_B_2zYF6yEk2_1;
	wire w_dff_B_S72RrKdf6_1;
	wire w_dff_B_bjDJvoz76_0;
	wire w_dff_B_1NnApfbK3_0;
	wire w_dff_B_Mz8I7oQ63_0;
	wire w_dff_B_kJ3TBsQJ6_0;
	wire w_dff_B_K8aNhHto4_0;
	wire w_dff_B_ZX58KJb36_1;
	wire w_dff_B_dmSDmjq87_1;
	wire w_dff_B_m4Ci5srJ3_1;
	wire w_dff_B_iyEaSrZ16_1;
	wire w_dff_B_DQMvCcBh2_1;
	wire w_dff_B_qh4TqmUH5_1;
	wire w_dff_B_s5EEVjOx9_0;
	wire w_dff_B_Lu1u8W6E1_0;
	wire w_dff_B_GwmRwY362_0;
	wire w_dff_B_d05Jrrm95_0;
	wire w_dff_B_i07KIMW05_1;
	wire w_dff_B_lDvUvXFE5_1;
	wire w_dff_B_vtqfyuMu0_1;
	wire w_dff_B_AmhI8UHA1_1;
	wire w_dff_B_nlpNDxfO7_1;
	wire w_dff_A_ldyRm5Sp4_1;
	wire w_dff_B_eoyEvq7x2_2;
	wire w_dff_B_tUJC509k0_1;
	wire w_dff_B_pDRcoDZO2_1;
	wire w_dff_B_LszaTL6P4_1;
	wire w_dff_B_sHrr4wRB8_1;
	wire w_dff_B_W13ktaNM2_1;
	wire w_dff_B_tzl0zDuC0_1;
	wire w_dff_B_8cIcvORO0_1;
	wire w_dff_B_x30379n46_1;
	wire w_dff_B_ZDi3jBiT2_1;
	wire w_dff_B_SFCaJsrj1_1;
	wire w_dff_B_WOBZxwkd3_1;
	wire w_dff_B_GrrYRaG21_1;
	wire w_dff_B_zyUCrIaE8_1;
	wire w_dff_B_hKWuVKxP1_1;
	wire w_dff_B_0KNpzkH01_2;
	wire w_dff_A_WP9bZbhQ6_0;
	wire w_dff_A_19rWTS8w4_0;
	wire w_dff_A_vQBAJatK4_1;
	wire w_dff_A_yDJmqpSx8_0;
	wire w_dff_A_lZwFM8ZI5_0;
	wire w_dff_A_pAecoUmY2_0;
	wire w_dff_A_uFXjBaex1_0;
	wire w_dff_A_PmFQJxZU4_0;
	wire w_dff_A_7516o1Wj1_0;
	wire w_dff_A_QR0VUwJA8_0;
	wire w_dff_A_GmH6zCB17_0;
	wire w_dff_A_U9nXheOp1_0;
	wire w_dff_A_B9BqP8PQ7_0;
	wire w_dff_A_lNLF2BjB4_0;
	wire w_dff_A_xR5oOP2r5_0;
	wire w_dff_A_EIvp8IWx3_0;
	wire w_dff_A_sL00PJx48_0;
	wire w_dff_A_sLW1frs88_0;
	wire w_dff_A_DGBD7lci8_0;
	wire w_dff_A_3hII8bb82_0;
	wire w_dff_A_lgYjaHiP5_0;
	wire w_dff_A_r3wG0ogX1_0;
	wire w_dff_A_2iu5bMul2_0;
	wire w_dff_A_xLU5Epjw5_0;
	wire w_dff_A_camGR4OS1_0;
	wire w_dff_A_8FjqrV9E6_0;
	wire w_dff_A_6xTW2Omh3_0;
	wire w_dff_A_JFAZPNSf9_0;
	wire w_dff_A_vJwNJk609_0;
	wire w_dff_A_f6xMlbQJ0_0;
	wire w_dff_A_rGMPTwGp0_0;
	wire w_dff_A_Yv3BvXIL8_0;
	wire w_dff_A_fyMvgymV0_0;
	wire w_dff_A_XuL0PMOG8_0;
	wire w_dff_A_DxWhPD141_0;
	wire w_dff_A_eEaul0dx2_0;
	wire w_dff_A_lsqm5opx1_0;
	wire w_dff_A_FiPshPat6_0;
	wire w_dff_A_B2Y1Nnml5_0;
	wire w_dff_A_ln96ecSa5_0;
	wire w_dff_A_K8Uc8uO82_0;
	wire w_dff_A_DnMtjMmI4_0;
	wire w_dff_A_tiJP9vMG7_0;
	wire w_dff_A_1EfO6lqI3_0;
	wire w_dff_A_sVOiuPDL6_0;
	wire w_dff_A_NkA4BtWt7_0;
	wire w_dff_A_hfstznWA8_0;
	wire w_dff_A_koaZlOGX7_0;
	wire w_dff_A_bpV6me7t3_0;
	wire w_dff_A_9cqNnkby4_0;
	wire w_dff_A_iMfraidZ2_0;
	wire w_dff_A_L6oQ0NhD3_0;
	wire w_dff_A_zvK8RSH07_0;
	wire w_dff_A_VnkAfI5P8_0;
	wire w_dff_A_uGrpNwGV6_0;
	wire w_dff_A_3ZRng7Ai9_0;
	wire w_dff_A_MCUPLppW4_0;
	wire w_dff_A_S61Jc8zR9_0;
	wire w_dff_A_v3rDdi969_0;
	wire w_dff_A_xv7cj5K92_0;
	wire w_dff_A_cwufwjbf6_0;
	wire w_dff_A_URs5L4D35_0;
	wire w_dff_A_EOt6XsKJ5_0;
	wire w_dff_A_ykR8CTuG2_0;
	wire w_dff_A_ubPgaL214_0;
	wire w_dff_A_axMy7jTL2_0;
	wire w_dff_A_H5xRXzh26_0;
	wire w_dff_A_PA8UFdlJ0_0;
	wire w_dff_A_UJNeqzmU5_0;
	wire w_dff_A_slxIVVxJ6_0;
	wire w_dff_A_Ghagossj9_0;
	wire w_dff_A_vEimH8TU6_0;
	wire w_dff_A_jufft8eE0_0;
	wire w_dff_A_1MWlUZeZ9_0;
	wire w_dff_A_y5q29IMO0_0;
	wire w_dff_A_w5aNIRF70_0;
	wire w_dff_A_HFwDfpPm3_2;
	wire w_dff_A_A4c8mjax2_0;
	wire w_dff_A_Njle6QaC8_0;
	wire w_dff_A_8GhHAcWv0_0;
	wire w_dff_A_FpePlT0U4_0;
	wire w_dff_A_K3ANNQyf9_0;
	wire w_dff_A_Qvg1yppC1_0;
	wire w_dff_A_3BucendH0_0;
	wire w_dff_A_7nMFY3eT0_0;
	wire w_dff_A_M8AfgK3h7_0;
	wire w_dff_A_Zu8ms7Rg8_0;
	wire w_dff_A_KvSSrMYO6_0;
	wire w_dff_A_ApJg33ru5_0;
	wire w_dff_A_hZFaVF6y3_0;
	wire w_dff_A_lOg3hT469_0;
	wire w_dff_A_nvTYsCxF4_0;
	wire w_dff_A_UOH1melP2_0;
	wire w_dff_A_hOSC90LA1_0;
	wire w_dff_A_zZgjbpdi2_0;
	wire w_dff_A_Uiwwkur33_0;
	wire w_dff_A_jolcGtlN3_0;
	wire w_dff_A_t8yUvLS06_0;
	wire w_dff_A_bprNHvkA9_0;
	wire w_dff_A_hqVSzu9O7_0;
	wire w_dff_A_BczsGttN5_0;
	wire w_dff_A_GWGiuHbv6_0;
	wire w_dff_A_sl5r2OFm7_0;
	wire w_dff_A_WKgYeipn3_0;
	wire w_dff_A_D25adAZR2_0;
	wire w_dff_A_KFf0f6sQ7_0;
	wire w_dff_A_kcDh5rxT7_0;
	wire w_dff_A_DrA9YxZp8_0;
	wire w_dff_A_WuUlyEvY4_0;
	wire w_dff_A_Mff4cG0V7_0;
	wire w_dff_A_c9hBSiem0_0;
	wire w_dff_A_FCgUzN3v7_0;
	wire w_dff_A_wOqsyxC38_0;
	wire w_dff_A_tqRN59FV1_0;
	wire w_dff_A_yIYHvv386_0;
	wire w_dff_A_LCTdrSdn8_0;
	wire w_dff_A_0cQgIh6a9_0;
	wire w_dff_A_Hmr0BAGN4_0;
	wire w_dff_A_Q3JbCeuL7_0;
	wire w_dff_A_2rE6LKwn7_0;
	wire w_dff_A_gOlzQcXr3_0;
	wire w_dff_A_zmuqQX1y4_0;
	wire w_dff_A_ey3pCS4B0_0;
	wire w_dff_A_Z7brXAli2_0;
	wire w_dff_A_TlzflgwK5_0;
	wire w_dff_A_7Rj678yq1_0;
	wire w_dff_A_AcnxaIQN5_0;
	wire w_dff_A_fJH9baaa4_0;
	wire w_dff_A_IIJctWqS5_0;
	wire w_dff_A_OrYl9Tm88_0;
	wire w_dff_A_P6h0nl4p4_0;
	wire w_dff_A_YxfdHJZr6_0;
	wire w_dff_A_6MOQtoeA0_0;
	wire w_dff_A_6RpKLiF12_0;
	wire w_dff_A_a2yxjw3a2_0;
	wire w_dff_A_qjzB4Z9t8_0;
	wire w_dff_A_jkkUfAJv6_0;
	wire w_dff_A_qKMfp8Dt5_0;
	wire w_dff_A_WoqI11ms6_0;
	wire w_dff_A_DlraXJsF2_0;
	wire w_dff_A_XR1bFcWX5_0;
	wire w_dff_A_seruZ6Fa5_0;
	wire w_dff_A_uECwVnlb2_0;
	wire w_dff_A_xTTaLZEK6_0;
	wire w_dff_A_VSXAMPib0_0;
	wire w_dff_A_gH9YZ6uC3_0;
	wire w_dff_A_RsDoFRkE0_2;
	wire w_dff_A_pBJQlEGq4_0;
	wire w_dff_A_RpRULNuW2_0;
	wire w_dff_A_e5HF90ds2_0;
	wire w_dff_A_xHzUFE0w9_0;
	wire w_dff_A_iOrBFzvF9_0;
	wire w_dff_A_uEMgeH9n2_0;
	wire w_dff_A_gor77tBY3_0;
	wire w_dff_A_lTGfop2H9_0;
	wire w_dff_A_5hbI78dF6_0;
	wire w_dff_A_ksLYVnJ73_0;
	wire w_dff_A_r89kxmHk7_0;
	wire w_dff_A_EdmRbVon5_0;
	wire w_dff_A_f8wQMqMZ5_0;
	wire w_dff_A_jB2IyY046_0;
	wire w_dff_A_FxiadecD1_0;
	wire w_dff_A_lVNUDG3p9_0;
	wire w_dff_A_xC5aIc0f4_0;
	wire w_dff_A_bSgQRPoh9_0;
	wire w_dff_A_KgaSOrHy6_0;
	wire w_dff_A_kOEpWpVj9_0;
	wire w_dff_A_y3FjiErL0_0;
	wire w_dff_A_NsKcCNXI8_0;
	wire w_dff_A_VJYGL9nz2_0;
	wire w_dff_A_fYR45Pcc6_0;
	wire w_dff_A_XQxi547z9_0;
	wire w_dff_A_aQkTh4fg4_0;
	wire w_dff_A_qCeRHAc97_0;
	wire w_dff_A_WbrauAlw8_0;
	wire w_dff_A_6R7MFucS8_0;
	wire w_dff_A_HVv8WAEd0_0;
	wire w_dff_A_yQOLCmJe4_0;
	wire w_dff_A_fChpvAtV5_0;
	wire w_dff_A_BVLGAnCp0_0;
	wire w_dff_A_LQGeLPW69_0;
	wire w_dff_A_oD6FFUYu2_0;
	wire w_dff_A_ZUlnMcF51_0;
	wire w_dff_A_M1tCmev92_0;
	wire w_dff_A_XjMUxa4I3_0;
	wire w_dff_A_ng7UeUqS7_0;
	wire w_dff_A_eZ3uWlS54_0;
	wire w_dff_A_CwRbadB94_0;
	wire w_dff_A_PfMru1ON8_0;
	wire w_dff_A_5eTsrVw56_0;
	wire w_dff_A_4RbthjPL5_0;
	wire w_dff_A_ivKjnPzW9_0;
	wire w_dff_A_i7bn42BC5_0;
	wire w_dff_A_P3QsJjAa4_0;
	wire w_dff_A_J7k8xNCL0_0;
	wire w_dff_A_YQ2HGsbt8_0;
	wire w_dff_A_NONL67SN7_0;
	wire w_dff_A_w6JVu9bk2_0;
	wire w_dff_A_qX4I8RST4_0;
	wire w_dff_A_oEw0h3W95_0;
	wire w_dff_A_I1mHrml95_0;
	wire w_dff_A_6kZC3iJ04_0;
	wire w_dff_A_9wRRePUh6_0;
	wire w_dff_A_jhNXnTh20_0;
	wire w_dff_A_fh7eCDxo5_0;
	wire w_dff_A_7AUygaGH5_0;
	wire w_dff_A_kaZy14qm6_0;
	wire w_dff_A_aYs1nTHT3_0;
	wire w_dff_A_8j8dHqgh7_0;
	wire w_dff_A_XAWMuwmi4_0;
	wire w_dff_A_H7UTNw2z5_0;
	wire w_dff_A_YznWS3Lm1_0;
	wire w_dff_A_RLSTf5Bj2_0;
	wire w_dff_A_MqlPqEgi9_0;
	wire w_dff_A_pjydccY89_0;
	wire w_dff_A_1xLXBDUh1_2;
	wire w_dff_A_xsu4rBt49_0;
	wire w_dff_A_k5BkWBtk7_0;
	wire w_dff_A_PQVsFRFi2_0;
	wire w_dff_A_uku0ZAZR9_0;
	wire w_dff_A_QfYY0DpD5_0;
	wire w_dff_A_jbDrEcJ23_0;
	wire w_dff_A_yROG9dB01_0;
	wire w_dff_A_CXPogtxx2_0;
	wire w_dff_A_PI1ULLSU5_0;
	wire w_dff_A_vkm5UZvG5_0;
	wire w_dff_A_yyMowZzA1_0;
	wire w_dff_A_LEaF1bsA9_0;
	wire w_dff_A_OEZJW24h5_0;
	wire w_dff_A_BBagiyHD6_0;
	wire w_dff_A_sdXcLymA1_0;
	wire w_dff_A_UCRcqDta2_0;
	wire w_dff_A_9jIW1bJN9_0;
	wire w_dff_A_FZ2ww8gG4_0;
	wire w_dff_A_7yokyOKu5_0;
	wire w_dff_A_ztLbhzp60_0;
	wire w_dff_A_0Cqhj6Rl1_0;
	wire w_dff_A_qahTg1QR1_0;
	wire w_dff_A_QfbEFPs25_0;
	wire w_dff_A_v8TmBlNa9_0;
	wire w_dff_A_GJoZHAUJ7_0;
	wire w_dff_A_nzm2KIE60_0;
	wire w_dff_A_PD83B6Xq1_0;
	wire w_dff_A_JjlHrhjj7_0;
	wire w_dff_A_YvhTfQmM9_0;
	wire w_dff_A_J01bPRDU4_0;
	wire w_dff_A_WI4akYC37_0;
	wire w_dff_A_Bcsxoab35_0;
	wire w_dff_A_sgOk7ufr0_0;
	wire w_dff_A_6NFXLFB45_0;
	wire w_dff_A_klwxy7Cy6_0;
	wire w_dff_A_G0fSCz8P5_0;
	wire w_dff_A_KInQa8R52_0;
	wire w_dff_A_IImVZS1d6_0;
	wire w_dff_A_SsgU5SUW7_0;
	wire w_dff_A_LW1yZJdS0_0;
	wire w_dff_A_XY7yEhb46_0;
	wire w_dff_A_YyDSFjD11_0;
	wire w_dff_A_NmETfZSo8_0;
	wire w_dff_A_ItpO6lpb2_0;
	wire w_dff_A_1qpEqiuq9_0;
	wire w_dff_A_tM64kL2f2_0;
	wire w_dff_A_ZtCEnyOQ6_0;
	wire w_dff_A_QHOWo0RC7_0;
	wire w_dff_A_o390FudG3_0;
	wire w_dff_A_OeteqeBr8_0;
	wire w_dff_A_nbB6fwHd1_0;
	wire w_dff_A_Xl6aWd1Q2_0;
	wire w_dff_A_pJ8IjpaS8_0;
	wire w_dff_A_yQiChqBE2_0;
	wire w_dff_A_Lps2nWTL1_0;
	wire w_dff_A_6D2gNe7X0_0;
	wire w_dff_A_aOa9I9ae0_0;
	wire w_dff_A_idDgyRDr6_0;
	wire w_dff_A_lWgC5v9h6_0;
	wire w_dff_A_HSrCP0S49_0;
	wire w_dff_A_PzcSGmdm1_0;
	wire w_dff_A_RTbgOhM20_0;
	wire w_dff_A_lWXAxUYh0_0;
	wire w_dff_A_F9LmMSId0_0;
	wire w_dff_A_CmXVFCyd7_0;
	wire w_dff_A_TeLedrld7_2;
	wire w_dff_A_bol0ejVz0_0;
	wire w_dff_A_t4LhVYjM3_0;
	wire w_dff_A_uacpOgHi5_0;
	wire w_dff_A_IU4O6lmQ3_0;
	wire w_dff_A_0VuVsBaC5_0;
	wire w_dff_A_wCLjnwhq7_0;
	wire w_dff_A_Ko6gxlib0_0;
	wire w_dff_A_3f08bY8f1_0;
	wire w_dff_A_8ijIKzc73_0;
	wire w_dff_A_n6T3EC4L6_0;
	wire w_dff_A_H1OWfJyx6_0;
	wire w_dff_A_oiTuYJ3v0_0;
	wire w_dff_A_eKp0PLuY3_0;
	wire w_dff_A_WUv6ZO6t9_0;
	wire w_dff_A_oT4gjTtw8_0;
	wire w_dff_A_EVMTMoUN5_0;
	wire w_dff_A_qMDPQIDd0_0;
	wire w_dff_A_t1zI0mwr3_0;
	wire w_dff_A_bs5lZ3yU2_0;
	wire w_dff_A_XnxGtaX32_0;
	wire w_dff_A_ZXXVlMKK2_0;
	wire w_dff_A_Vt9Hp3ou0_0;
	wire w_dff_A_yv2P0WMO0_0;
	wire w_dff_A_VKYp5l2u8_0;
	wire w_dff_A_9uwWeksb3_0;
	wire w_dff_A_7u72UeB25_0;
	wire w_dff_A_BJAw2yFA0_0;
	wire w_dff_A_JZWhghGf9_0;
	wire w_dff_A_X96sUsPH8_0;
	wire w_dff_A_v6cG4XWl5_0;
	wire w_dff_A_iEfdnanX3_0;
	wire w_dff_A_8dtyyjYc7_0;
	wire w_dff_A_dou3YUic3_0;
	wire w_dff_A_17qQnhVk4_0;
	wire w_dff_A_IqYsLYKj4_0;
	wire w_dff_A_BeU2OFCx0_0;
	wire w_dff_A_HnQaH6tW5_0;
	wire w_dff_A_drPL1Zui5_0;
	wire w_dff_A_LLT0fVxj1_0;
	wire w_dff_A_kDsHfPOj1_0;
	wire w_dff_A_5i3tz4Zv8_0;
	wire w_dff_A_qq3dITRB2_0;
	wire w_dff_A_ky4f0O2O2_0;
	wire w_dff_A_PvON90P24_0;
	wire w_dff_A_pF6tsaKP3_0;
	wire w_dff_A_atT6eD336_0;
	wire w_dff_A_Y3ohAWku0_0;
	wire w_dff_A_kLfdbApj6_0;
	wire w_dff_A_XqbapEyq8_0;
	wire w_dff_A_VjlNLbQz5_0;
	wire w_dff_A_DeEPtQdM3_0;
	wire w_dff_A_ZosguoP75_0;
	wire w_dff_A_cwWfmgn85_0;
	wire w_dff_A_bze71XGT3_0;
	wire w_dff_A_5mX8apPa9_0;
	wire w_dff_A_4YqBnL7B1_0;
	wire w_dff_A_cbasXw8a5_0;
	wire w_dff_A_zr21BW4f6_0;
	wire w_dff_A_cMAfwCVk0_0;
	wire w_dff_A_pJ33Hvnf2_0;
	wire w_dff_A_z7YRI3e49_0;
	wire w_dff_A_vT9YTuSq8_0;
	wire w_dff_A_TwM7lXbz1_2;
	wire w_dff_A_UAJW3X5l7_0;
	wire w_dff_A_j9B9Jvno8_0;
	wire w_dff_A_Q0c5kvtw1_0;
	wire w_dff_A_jIDC6kEQ7_0;
	wire w_dff_A_9JDPLOyP6_0;
	wire w_dff_A_sTrmOqhF6_0;
	wire w_dff_A_ZEdZut1c0_0;
	wire w_dff_A_4eYIvfCU3_0;
	wire w_dff_A_W9nowCdM3_0;
	wire w_dff_A_FCeCjAjz7_0;
	wire w_dff_A_RCFfnfy77_0;
	wire w_dff_A_PucO2c7U3_0;
	wire w_dff_A_Whz0sEPe6_0;
	wire w_dff_A_VeyoKap24_0;
	wire w_dff_A_jpfNtqAp9_0;
	wire w_dff_A_1miHCnrf2_0;
	wire w_dff_A_964Cxv4P3_0;
	wire w_dff_A_jDHBWnsD0_0;
	wire w_dff_A_0qfWCUNQ3_0;
	wire w_dff_A_YQudfU5M5_0;
	wire w_dff_A_CGmkKv4x4_0;
	wire w_dff_A_i8A7DZtS8_0;
	wire w_dff_A_WyQ2V4mb9_0;
	wire w_dff_A_8qSuFptH6_0;
	wire w_dff_A_qlC1par80_0;
	wire w_dff_A_6GLPw8WD8_0;
	wire w_dff_A_OxYs3xHo5_0;
	wire w_dff_A_VfmVkD5U5_0;
	wire w_dff_A_zXjrJcwF9_0;
	wire w_dff_A_6HQEtJCb3_0;
	wire w_dff_A_CqBS3ekW3_0;
	wire w_dff_A_39PURsZS2_0;
	wire w_dff_A_9BBI98LA7_0;
	wire w_dff_A_1AzSRlcb6_0;
	wire w_dff_A_SPKTtnlj1_0;
	wire w_dff_A_dknCnWo04_0;
	wire w_dff_A_g7BbC1sk9_0;
	wire w_dff_A_1pagNIXs4_0;
	wire w_dff_A_Rsnqd1pV2_0;
	wire w_dff_A_BdbkCvEe4_0;
	wire w_dff_A_aCSqIg5N2_0;
	wire w_dff_A_tHWsRnni2_0;
	wire w_dff_A_0Z0SbmFk8_0;
	wire w_dff_A_eL3TauJW9_0;
	wire w_dff_A_lu2ZM6HD0_0;
	wire w_dff_A_SNTgbLB45_0;
	wire w_dff_A_QK1XmSw77_0;
	wire w_dff_A_95mC63sH8_0;
	wire w_dff_A_Gis0XsyP0_0;
	wire w_dff_A_59nN0qvZ8_0;
	wire w_dff_A_xISAQfzA5_0;
	wire w_dff_A_D5gWjrEs7_0;
	wire w_dff_A_jYe5tZmU6_0;
	wire w_dff_A_xLRE8IRU5_0;
	wire w_dff_A_rmI08Fv90_0;
	wire w_dff_A_iyAoaOiS3_0;
	wire w_dff_A_f0ptJyQF8_0;
	wire w_dff_A_Axi3T5mV9_0;
	wire w_dff_A_Mslu13Cv9_0;
	wire w_dff_A_vUFKz7gI5_2;
	wire w_dff_A_1nGxUdwc0_0;
	wire w_dff_A_k2HBAkGy2_0;
	wire w_dff_A_zIuU1lhr8_0;
	wire w_dff_A_Iue0EIvQ9_0;
	wire w_dff_A_VmI0LVzu0_0;
	wire w_dff_A_r32ypvQj5_0;
	wire w_dff_A_9fQR6I3j3_0;
	wire w_dff_A_dms0CAFp0_0;
	wire w_dff_A_RRdA6QGb9_0;
	wire w_dff_A_2kgG5PXq3_0;
	wire w_dff_A_xDeq4DB57_0;
	wire w_dff_A_evdO9kTn3_0;
	wire w_dff_A_9P5ldShi1_0;
	wire w_dff_A_VMtbtwgH4_0;
	wire w_dff_A_5awSSqAp1_0;
	wire w_dff_A_yVS4wdMT3_0;
	wire w_dff_A_7wYmTe2D3_0;
	wire w_dff_A_ah3ui2GP6_0;
	wire w_dff_A_kNtpU5qE0_0;
	wire w_dff_A_P5BwMx4P8_0;
	wire w_dff_A_zbUnAbP68_0;
	wire w_dff_A_smQS5U6o0_0;
	wire w_dff_A_HkbiOc7H2_0;
	wire w_dff_A_98f1L4iL7_0;
	wire w_dff_A_p5ub0H2O5_0;
	wire w_dff_A_ALfQnhZL1_0;
	wire w_dff_A_0pAenHLj8_0;
	wire w_dff_A_E5Z5407s9_0;
	wire w_dff_A_PFF1U29P9_0;
	wire w_dff_A_ufi1obGv0_0;
	wire w_dff_A_4RIIh9zI9_0;
	wire w_dff_A_hFKqM5e91_0;
	wire w_dff_A_JOQPHkc96_0;
	wire w_dff_A_VLkM2l799_0;
	wire w_dff_A_RSeIIm0c1_0;
	wire w_dff_A_QOBVIXpe1_0;
	wire w_dff_A_T7LNFpVn4_0;
	wire w_dff_A_6GzhWNzm8_0;
	wire w_dff_A_PvxLyntL5_0;
	wire w_dff_A_6mtRfzYp9_0;
	wire w_dff_A_PBHcEw8k8_0;
	wire w_dff_A_zAHplGTV6_0;
	wire w_dff_A_wwhNBayJ5_0;
	wire w_dff_A_MM9i1v2l6_0;
	wire w_dff_A_hx3XmgLs4_0;
	wire w_dff_A_1tPG0c9q7_0;
	wire w_dff_A_5ymGjRTW1_0;
	wire w_dff_A_VQBN6s995_0;
	wire w_dff_A_RqPqsYCC1_0;
	wire w_dff_A_0ZYYcHJU3_0;
	wire w_dff_A_uT3NRADn6_0;
	wire w_dff_A_N1ZwoG8s4_0;
	wire w_dff_A_aiNHm7782_0;
	wire w_dff_A_zMA41CAZ9_0;
	wire w_dff_A_sEa4t8eO6_0;
	wire w_dff_A_NCFPQcXO1_0;
	wire w_dff_A_x5iNlZpF9_2;
	wire w_dff_A_lYD5SFbp2_0;
	wire w_dff_A_G7YWsEkZ1_0;
	wire w_dff_A_NBync2rf9_0;
	wire w_dff_A_EcTbDsa87_0;
	wire w_dff_A_t5VhvoHX0_0;
	wire w_dff_A_70OTFWmL8_0;
	wire w_dff_A_vO9UCCjL5_0;
	wire w_dff_A_MppMk7Nq5_0;
	wire w_dff_A_3rkWYmv03_0;
	wire w_dff_A_3wtYIhbw0_0;
	wire w_dff_A_lgQnK0hh6_0;
	wire w_dff_A_u2PABcCo6_0;
	wire w_dff_A_45FLl0c18_0;
	wire w_dff_A_jYK3K8x19_0;
	wire w_dff_A_wp7RYLUY5_0;
	wire w_dff_A_SLgo7Hm12_0;
	wire w_dff_A_VR4tcPvC9_0;
	wire w_dff_A_K3qZg2mx2_0;
	wire w_dff_A_WcyON9jG0_0;
	wire w_dff_A_fhbtDnig0_0;
	wire w_dff_A_SOMJbvNS3_0;
	wire w_dff_A_IbN7RXvn4_0;
	wire w_dff_A_sKbt3blr9_0;
	wire w_dff_A_rKPQto8e6_0;
	wire w_dff_A_iK1BqmU17_0;
	wire w_dff_A_JYff3aHV5_0;
	wire w_dff_A_6WG55EaU0_0;
	wire w_dff_A_z3kkVhEv8_0;
	wire w_dff_A_c3xRUcvx2_0;
	wire w_dff_A_kIM7Lkv92_0;
	wire w_dff_A_22NrmKdu1_0;
	wire w_dff_A_bAxytHLF9_0;
	wire w_dff_A_ueek6hZa8_0;
	wire w_dff_A_PfvWyb6E9_0;
	wire w_dff_A_V38DQqUm1_0;
	wire w_dff_A_YsJxLQ5t5_0;
	wire w_dff_A_8fpeffk00_0;
	wire w_dff_A_onlsQOkI3_0;
	wire w_dff_A_sT9b0ne13_0;
	wire w_dff_A_8QXdAe2M4_0;
	wire w_dff_A_5ULWgtiY9_0;
	wire w_dff_A_G0RJgVBj9_0;
	wire w_dff_A_d9T9VPEA3_0;
	wire w_dff_A_RNfkP6KG7_0;
	wire w_dff_A_zy7wlXDR1_0;
	wire w_dff_A_wA2la3kr3_0;
	wire w_dff_A_mcXzZJOI9_0;
	wire w_dff_A_itegJ70E7_0;
	wire w_dff_A_yaabpSOV7_0;
	wire w_dff_A_Ze7ewDjf8_0;
	wire w_dff_A_gnTNupHv5_0;
	wire w_dff_A_ib3Y8QpA0_0;
	wire w_dff_A_XkuYRI3a5_0;
	wire w_dff_A_tlP6TWHP5_2;
	wire w_dff_A_htKEXvld9_0;
	wire w_dff_A_eVa3qwvq5_0;
	wire w_dff_A_V91giNQZ4_0;
	wire w_dff_A_tiUeNl3k3_0;
	wire w_dff_A_8sAveCFd5_0;
	wire w_dff_A_zNw5rJOg1_0;
	wire w_dff_A_HGobqhKa8_0;
	wire w_dff_A_CPCuflJL8_0;
	wire w_dff_A_Y10nIyer7_0;
	wire w_dff_A_8N9H7D134_0;
	wire w_dff_A_hCwHbhsg6_0;
	wire w_dff_A_ygr39j160_0;
	wire w_dff_A_YuP7Jw1q2_0;
	wire w_dff_A_TVh0ArG66_0;
	wire w_dff_A_uyHRBDmb6_0;
	wire w_dff_A_564fWMVj5_0;
	wire w_dff_A_EgqQlhWB1_0;
	wire w_dff_A_3E5unMHL9_0;
	wire w_dff_A_ELdSFDX40_0;
	wire w_dff_A_QxzFyfou2_0;
	wire w_dff_A_KjZ2f8T25_0;
	wire w_dff_A_2o5DQ8Mt5_0;
	wire w_dff_A_IH5lNMX90_0;
	wire w_dff_A_mu0Z9Cv63_0;
	wire w_dff_A_hCjLP8dp6_0;
	wire w_dff_A_qDwBBmUR1_0;
	wire w_dff_A_ARlbxat40_0;
	wire w_dff_A_GOx0FYBK7_0;
	wire w_dff_A_I33b71Kd9_0;
	wire w_dff_A_XKtWoxgP6_0;
	wire w_dff_A_69iJw6Xi4_0;
	wire w_dff_A_QB7m5PNs8_0;
	wire w_dff_A_1FxkTZab5_0;
	wire w_dff_A_i5GSygaG3_0;
	wire w_dff_A_Bu3knTpj8_0;
	wire w_dff_A_P9d1Losl4_0;
	wire w_dff_A_v3ljCD6s3_0;
	wire w_dff_A_r8lg5iZI1_0;
	wire w_dff_A_AwGZmeen1_0;
	wire w_dff_A_xx6Hhrow5_0;
	wire w_dff_A_qomTXFr90_0;
	wire w_dff_A_DMEN1KHw8_0;
	wire w_dff_A_FbkpCx526_0;
	wire w_dff_A_yUyw4dIv6_0;
	wire w_dff_A_UxWic4sR2_0;
	wire w_dff_A_3uJZLNB75_0;
	wire w_dff_A_NtmaUURD2_0;
	wire w_dff_A_MFI1bAwp5_0;
	wire w_dff_A_6qzdKOMX1_0;
	wire w_dff_A_sXErAsAX8_0;
	wire w_dff_A_HcHGc8GI5_2;
	wire w_dff_A_qsoH4gB39_0;
	wire w_dff_A_nIP3F0dU4_0;
	wire w_dff_A_fvBVW7Tm8_0;
	wire w_dff_A_J8vI6M7I0_0;
	wire w_dff_A_sAcLa3sX6_0;
	wire w_dff_A_E95lJQPi8_0;
	wire w_dff_A_o93XOJ8P1_0;
	wire w_dff_A_40n6Vg5T0_0;
	wire w_dff_A_dKmeG3aR2_0;
	wire w_dff_A_AX1nK5VO6_0;
	wire w_dff_A_se1GDjip4_0;
	wire w_dff_A_Mmp8GNwa8_0;
	wire w_dff_A_AYvbEJrm8_0;
	wire w_dff_A_CJokU8Jk0_0;
	wire w_dff_A_nwawaXxH4_0;
	wire w_dff_A_hTsoAsnB1_0;
	wire w_dff_A_0ipCLz0L4_0;
	wire w_dff_A_UQQq3KWs9_0;
	wire w_dff_A_ibWbl1Nr1_0;
	wire w_dff_A_WV1P5eZ88_0;
	wire w_dff_A_nxvAh8NZ1_0;
	wire w_dff_A_QhpKQxvp0_0;
	wire w_dff_A_Rt0A6Q1L9_0;
	wire w_dff_A_XGf37ncy2_0;
	wire w_dff_A_i00ovWSt2_0;
	wire w_dff_A_pEuYcoju9_0;
	wire w_dff_A_Zn3mKGlE8_0;
	wire w_dff_A_mUCvp3GE2_0;
	wire w_dff_A_9kMotp116_0;
	wire w_dff_A_adUvZHCo2_0;
	wire w_dff_A_Pk1mll5I8_0;
	wire w_dff_A_0z0MehKw5_0;
	wire w_dff_A_UMdm7bR86_0;
	wire w_dff_A_WXZ0mLsa1_0;
	wire w_dff_A_Eh13WoxW3_0;
	wire w_dff_A_6SluiaN89_0;
	wire w_dff_A_lxDaDdos1_0;
	wire w_dff_A_6wMztMHk8_0;
	wire w_dff_A_44cAN4210_0;
	wire w_dff_A_UxijUgdI0_0;
	wire w_dff_A_ArdSPo6G5_0;
	wire w_dff_A_v5Xyjrb10_0;
	wire w_dff_A_h1Wl5xaf7_0;
	wire w_dff_A_JAvxWtIC6_0;
	wire w_dff_A_EZQkrqlz6_0;
	wire w_dff_A_LGB74pSN9_0;
	wire w_dff_A_F13iuZHC0_0;
	wire w_dff_A_Z99VGWH31_2;
	wire w_dff_A_0rPlNvCR0_0;
	wire w_dff_A_4At6yBK88_0;
	wire w_dff_A_E1mn4PEJ2_0;
	wire w_dff_A_HGjQL6Jk6_0;
	wire w_dff_A_yY0quIV29_0;
	wire w_dff_A_mQUd3zN64_0;
	wire w_dff_A_os0rrg7F4_0;
	wire w_dff_A_xei5nxWQ3_0;
	wire w_dff_A_ic61KOAc0_0;
	wire w_dff_A_ebianqhH1_0;
	wire w_dff_A_PLZnnfak3_0;
	wire w_dff_A_P5xy79OU0_0;
	wire w_dff_A_1YcfwdP87_0;
	wire w_dff_A_ra44eOUw8_0;
	wire w_dff_A_Fj8Eu6e52_0;
	wire w_dff_A_kIdF5RLh9_0;
	wire w_dff_A_6EO4qM4U7_0;
	wire w_dff_A_sWLnCkTn6_0;
	wire w_dff_A_kmsaJNrm5_0;
	wire w_dff_A_fwtl1zsk6_0;
	wire w_dff_A_qlvSIQUw9_0;
	wire w_dff_A_poZbm5i38_0;
	wire w_dff_A_CcAktltv3_0;
	wire w_dff_A_g9DfIthW7_0;
	wire w_dff_A_DItL0nNR3_0;
	wire w_dff_A_fWc5zKYH5_0;
	wire w_dff_A_rppv83j64_0;
	wire w_dff_A_iQGHrDZj3_0;
	wire w_dff_A_Mk6r4eNl7_0;
	wire w_dff_A_ZZ646FKw6_0;
	wire w_dff_A_ZBHma7Vm9_0;
	wire w_dff_A_XZgMTY9c5_0;
	wire w_dff_A_wAhbELF39_0;
	wire w_dff_A_YtxxQRmc1_0;
	wire w_dff_A_bABEPoPm6_0;
	wire w_dff_A_278nQgmT9_0;
	wire w_dff_A_mzMs0Jyu8_0;
	wire w_dff_A_cEKN8g9d7_0;
	wire w_dff_A_PPydyZsY3_0;
	wire w_dff_A_L6jSa4y59_0;
	wire w_dff_A_0ijJLyNe7_0;
	wire w_dff_A_zvxYt7Tv4_0;
	wire w_dff_A_LYTHLc343_0;
	wire w_dff_A_vilZNmuY8_0;
	wire w_dff_A_afeJhXAY4_2;
	wire w_dff_A_KLSSrEtu1_0;
	wire w_dff_A_gHp6ahtl2_0;
	wire w_dff_A_Mg8zQyCk3_0;
	wire w_dff_A_TlomVDoF6_0;
	wire w_dff_A_Alvdk1Bo6_0;
	wire w_dff_A_yoZXois07_0;
	wire w_dff_A_EAAkAPMg0_0;
	wire w_dff_A_fyOO9pcj6_0;
	wire w_dff_A_wcYj8kzg4_0;
	wire w_dff_A_jpQoDH987_0;
	wire w_dff_A_SMa2VANT8_0;
	wire w_dff_A_uOgRbNDV4_0;
	wire w_dff_A_wkrWorlu6_0;
	wire w_dff_A_05lb2NUr1_0;
	wire w_dff_A_0c39Pvsv8_0;
	wire w_dff_A_ZqlMTaoa4_0;
	wire w_dff_A_GCcWrlU12_0;
	wire w_dff_A_KqbgoRB20_0;
	wire w_dff_A_WHoVlYTy2_0;
	wire w_dff_A_rVpqoafh9_0;
	wire w_dff_A_bzX8rOTV5_0;
	wire w_dff_A_NzWoy8JQ3_0;
	wire w_dff_A_vWijRKai2_0;
	wire w_dff_A_1E1qQpmS1_0;
	wire w_dff_A_JJmaRRDd6_0;
	wire w_dff_A_T3WsZX3e0_0;
	wire w_dff_A_FN4zFvGm2_0;
	wire w_dff_A_Q9Wf0lyB1_0;
	wire w_dff_A_SRBgKef43_0;
	wire w_dff_A_7858yQTM7_0;
	wire w_dff_A_wCVTmF9v6_0;
	wire w_dff_A_wLUv0HrY8_0;
	wire w_dff_A_Ac974i1p7_0;
	wire w_dff_A_TNvEFM7X6_0;
	wire w_dff_A_vus6YOYj3_0;
	wire w_dff_A_RqfofxOU4_0;
	wire w_dff_A_DZQwGa1a9_0;
	wire w_dff_A_0fvfonUl5_0;
	wire w_dff_A_Lp5wsFC31_0;
	wire w_dff_A_JV1KtkJ67_0;
	wire w_dff_A_eRseWFyr5_0;
	wire w_dff_A_FoMYUxYC3_2;
	wire w_dff_A_gnvhzIGn4_0;
	wire w_dff_A_6izX916a9_0;
	wire w_dff_A_AcjGaaqB8_0;
	wire w_dff_A_qUUaUic41_0;
	wire w_dff_A_9HfdYidC8_0;
	wire w_dff_A_JdxyEs2o2_0;
	wire w_dff_A_g929yfn40_0;
	wire w_dff_A_jEPR9xl32_0;
	wire w_dff_A_q00CaeYe8_0;
	wire w_dff_A_KB3E3Z3z5_0;
	wire w_dff_A_bu7JjBvx2_0;
	wire w_dff_A_XAjSpPdI0_0;
	wire w_dff_A_2kz2U6hn6_0;
	wire w_dff_A_LLCGoYyS9_0;
	wire w_dff_A_WSdTx86Z0_0;
	wire w_dff_A_eOtDSeHO8_0;
	wire w_dff_A_lwQvF2y68_0;
	wire w_dff_A_ltxo5Jfm3_0;
	wire w_dff_A_jDGWNsFa2_0;
	wire w_dff_A_c6iRBxs45_0;
	wire w_dff_A_X5CZYujQ6_0;
	wire w_dff_A_rcVE5MdU7_0;
	wire w_dff_A_z0GMMdU54_0;
	wire w_dff_A_FTnuWQEh9_0;
	wire w_dff_A_fE3fl2JK8_0;
	wire w_dff_A_rRNZePuO7_0;
	wire w_dff_A_d9OqFF5V7_0;
	wire w_dff_A_etJLtNuo9_0;
	wire w_dff_A_lHIzLgsf4_0;
	wire w_dff_A_go9bXObM4_0;
	wire w_dff_A_0onAaVvQ7_0;
	wire w_dff_A_4TGbiVYl3_0;
	wire w_dff_A_GaMGoxSt0_0;
	wire w_dff_A_mYNbI0pB0_0;
	wire w_dff_A_PSrvcFwT1_0;
	wire w_dff_A_jEqiU7ii3_0;
	wire w_dff_A_T8rXtJu05_0;
	wire w_dff_A_8G1VuqpI6_0;
	wire w_dff_A_GmHJ0a9t0_2;
	wire w_dff_A_dSbbVZ3o7_0;
	wire w_dff_A_NZPOisht3_0;
	wire w_dff_A_SAjOOS886_0;
	wire w_dff_A_W8kKom7e5_0;
	wire w_dff_A_kWZP04ST6_0;
	wire w_dff_A_sbdJc6K36_0;
	wire w_dff_A_X4T6FdVr5_0;
	wire w_dff_A_RmsVUeVX5_0;
	wire w_dff_A_YkMKAMDb1_0;
	wire w_dff_A_MPxEYMBQ5_0;
	wire w_dff_A_Rs20P8xn1_0;
	wire w_dff_A_dPHorXnj0_0;
	wire w_dff_A_yzyNEFai1_0;
	wire w_dff_A_xwzNulXl4_0;
	wire w_dff_A_ZkaOgzgl6_0;
	wire w_dff_A_VKmschiw8_0;
	wire w_dff_A_HtKEXHjw5_0;
	wire w_dff_A_UhL7JSLh0_0;
	wire w_dff_A_tdiJykEE2_0;
	wire w_dff_A_cvEEGpoF9_0;
	wire w_dff_A_Q9JFcfxe0_0;
	wire w_dff_A_VvpZKsHW0_0;
	wire w_dff_A_R2k5lUdt0_0;
	wire w_dff_A_YbcYynJs9_0;
	wire w_dff_A_t3ukUg8n0_0;
	wire w_dff_A_hP5cGmAH5_0;
	wire w_dff_A_sW38N8fZ8_0;
	wire w_dff_A_nzYRjUJx3_0;
	wire w_dff_A_sD7fZ1M95_0;
	wire w_dff_A_QlQYNq4Y4_0;
	wire w_dff_A_qCfFwf2z5_0;
	wire w_dff_A_bXDfj5za1_0;
	wire w_dff_A_yu9252Xt7_0;
	wire w_dff_A_JBT4MzeO3_0;
	wire w_dff_A_XOBfWwGa2_0;
	wire w_dff_A_XaMEPoS81_2;
	wire w_dff_A_5QF3iZPZ9_0;
	wire w_dff_A_bQLsF19t0_0;
	wire w_dff_A_NBDITLYh6_0;
	wire w_dff_A_qiwKXeqI2_0;
	wire w_dff_A_OZcaRXYt3_0;
	wire w_dff_A_qjGaneWF7_0;
	wire w_dff_A_1YLz3UET5_0;
	wire w_dff_A_u7LQ7PlU6_0;
	wire w_dff_A_V20hFW2X6_0;
	wire w_dff_A_DPxxtKL94_0;
	wire w_dff_A_Wap2CB2h7_0;
	wire w_dff_A_UQaAL50u2_0;
	wire w_dff_A_S9snbeRI7_0;
	wire w_dff_A_7IQzRKXI5_0;
	wire w_dff_A_Utk6dRhz3_0;
	wire w_dff_A_RxYoKcRC1_0;
	wire w_dff_A_pPyncxk59_0;
	wire w_dff_A_KXhRlyXG2_0;
	wire w_dff_A_M1TIjveT3_0;
	wire w_dff_A_QcxhskVs4_0;
	wire w_dff_A_Cpsp4XmA0_0;
	wire w_dff_A_a3jxP59A5_0;
	wire w_dff_A_QOF6Jm5n6_0;
	wire w_dff_A_iiys9Ega1_0;
	wire w_dff_A_yl056mB47_0;
	wire w_dff_A_WY6T1iOP1_0;
	wire w_dff_A_Y6DoH7Lu0_0;
	wire w_dff_A_VjKk6thg6_0;
	wire w_dff_A_u6CIoNnq9_0;
	wire w_dff_A_RjEsBuRu8_0;
	wire w_dff_A_tTsaSnpf8_0;
	wire w_dff_A_8ZOo8LCE9_0;
	wire w_dff_A_r1aCngrq2_2;
	wire w_dff_A_XuFRjrVs3_0;
	wire w_dff_A_v9YqiqXu5_0;
	wire w_dff_A_9AXGyz639_0;
	wire w_dff_A_C35h2YZ36_0;
	wire w_dff_A_UHFQyyOC2_0;
	wire w_dff_A_VjVYa70F9_0;
	wire w_dff_A_AV07rs3B7_0;
	wire w_dff_A_OEBhgR793_0;
	wire w_dff_A_GVKpoXPD8_0;
	wire w_dff_A_3mwVx50J9_0;
	wire w_dff_A_OWo3gA2u8_0;
	wire w_dff_A_HjjsXZHh5_0;
	wire w_dff_A_BqowqEYv2_0;
	wire w_dff_A_Wd9GDAVx7_0;
	wire w_dff_A_yY3USx4c0_0;
	wire w_dff_A_vJDQ2GWV8_0;
	wire w_dff_A_9AdVyImf4_0;
	wire w_dff_A_u4N4Uje02_0;
	wire w_dff_A_9CxBwdcR8_0;
	wire w_dff_A_twn4eA197_0;
	wire w_dff_A_x361I8aL4_0;
	wire w_dff_A_fJuP8nTE4_0;
	wire w_dff_A_ehniVHbJ3_0;
	wire w_dff_A_uVQFxzYX4_0;
	wire w_dff_A_iXpVjrUq3_0;
	wire w_dff_A_clUjrJxA2_0;
	wire w_dff_A_pHNxuWoO9_0;
	wire w_dff_A_4nlKqnzp8_0;
	wire w_dff_A_i6PJMHws9_0;
	wire w_dff_A_Jo2F7egf8_2;
	wire w_dff_A_R1YbaEy04_0;
	wire w_dff_A_XG9gEGcT6_0;
	wire w_dff_A_ysQ9zyiw7_0;
	wire w_dff_A_ISRYGuJm7_0;
	wire w_dff_A_rjK2P2tH5_0;
	wire w_dff_A_IrYfBgBQ4_0;
	wire w_dff_A_5HGTNa9z9_0;
	wire w_dff_A_oCFTjAhD7_0;
	wire w_dff_A_eHkZvevr2_0;
	wire w_dff_A_NVe5xkYR6_0;
	wire w_dff_A_ei635nAD0_0;
	wire w_dff_A_Awg7C87t3_0;
	wire w_dff_A_9TWscmz96_0;
	wire w_dff_A_3WYPxpMa1_0;
	wire w_dff_A_qhsh2jpC2_0;
	wire w_dff_A_museoPD78_0;
	wire w_dff_A_bx0B8RLP8_0;
	wire w_dff_A_sDO8aYuP9_0;
	wire w_dff_A_mT9KQcqW7_0;
	wire w_dff_A_JKjdBYHm7_0;
	wire w_dff_A_ANsx75UK5_0;
	wire w_dff_A_WdxnNWbO0_0;
	wire w_dff_A_x5luIduw5_0;
	wire w_dff_A_DbbIKP4b6_0;
	wire w_dff_A_PtLRZelp4_0;
	wire w_dff_A_XbyGK9nu9_0;
	wire w_dff_A_sRgAlPUg1_0;
	wire w_dff_A_4izfRJkS6_2;
	wire w_dff_A_ppsMkLmp8_0;
	wire w_dff_A_zJoUeEbX8_0;
	wire w_dff_A_owbrdXYS4_0;
	wire w_dff_A_wP8pYvmu2_0;
	wire w_dff_A_Pj0roopd0_0;
	wire w_dff_A_bHuVC1ga7_0;
	wire w_dff_A_hqbjXSw79_0;
	wire w_dff_A_25DlQBwS8_0;
	wire w_dff_A_rBRUGHOt2_0;
	wire w_dff_A_1AatJLuc1_0;
	wire w_dff_A_zfOMHR2N7_0;
	wire w_dff_A_H6zG2bVS3_0;
	wire w_dff_A_ctlM9ASg1_0;
	wire w_dff_A_L6w3cSdp8_0;
	wire w_dff_A_KkFqToFD8_0;
	wire w_dff_A_vTI7170r4_0;
	wire w_dff_A_Ys7EmmBa4_0;
	wire w_dff_A_8xEIQZeC8_0;
	wire w_dff_A_wcm2MRYr4_0;
	wire w_dff_A_pvTt9bvg1_0;
	wire w_dff_A_0DoxGEUH1_0;
	wire w_dff_A_H0FKafym0_0;
	wire w_dff_A_6Z8AVGmP7_0;
	wire w_dff_A_dbUExD566_0;
	wire w_dff_A_L4JrPjBs8_0;
	wire w_dff_A_x9VZLpLG1_2;
	wire w_dff_A_hzCEB60T6_0;
	wire w_dff_A_VACDEFBw0_0;
	wire w_dff_A_j3WUboOe1_0;
	wire w_dff_A_7b85qm3S8_0;
	wire w_dff_A_W7pE5v2l1_0;
	wire w_dff_A_HQKdiD9s4_0;
	wire w_dff_A_F2xwVygP3_0;
	wire w_dff_A_PSnqNOKP1_0;
	wire w_dff_A_gA6GfLkW5_0;
	wire w_dff_A_57KLEFYh0_0;
	wire w_dff_A_TvW63X6d6_0;
	wire w_dff_A_o2MrrdRB9_0;
	wire w_dff_A_sKac6gYO8_0;
	wire w_dff_A_uDCZ8FDm6_0;
	wire w_dff_A_JNWJh7cx5_0;
	wire w_dff_A_hdd8L2608_0;
	wire w_dff_A_xLEkBZKi1_0;
	wire w_dff_A_8B1JFkR21_0;
	wire w_dff_A_XXhdQzVp9_0;
	wire w_dff_A_vpLYzyqZ6_0;
	wire w_dff_A_8B162l1j9_0;
	wire w_dff_A_fbjChCzp6_0;
	wire w_dff_A_d5G44bY50_0;
	wire w_dff_A_892Ip4n51_0;
	wire w_dff_A_4IuXdUMj6_2;
	wire w_dff_A_mD81bi5v7_0;
	wire w_dff_A_nMIKE5cS2_0;
	wire w_dff_A_UWiyTxOQ7_0;
	wire w_dff_A_2yv6LY7Y9_0;
	wire w_dff_A_2V2pQONp6_0;
	wire w_dff_A_iupM7qmo1_0;
	wire w_dff_A_M3lqxB9h1_0;
	wire w_dff_A_8ZtcXfmc8_0;
	wire w_dff_A_87cMEnYt4_0;
	wire w_dff_A_nh2SJF7z6_0;
	wire w_dff_A_UGjwBSOp4_0;
	wire w_dff_A_JkqT5Qtz2_0;
	wire w_dff_A_rAWPsB6q3_0;
	wire w_dff_A_TjZDc58h2_0;
	wire w_dff_A_ICaJKK2y7_0;
	wire w_dff_A_ybsYYklZ1_0;
	wire w_dff_A_DoG3Qxi32_0;
	wire w_dff_A_f5p4Rh8X5_0;
	wire w_dff_A_U33AsfOZ5_0;
	wire w_dff_A_wA95lBlI2_0;
	wire w_dff_A_pgP3a0OZ0_0;
	wire w_dff_A_FqZVic4Z9_0;
	wire w_dff_A_UJSpteTt5_2;
	wire w_dff_A_jkiZPCWk7_0;
	wire w_dff_A_AjsoM0Mb5_0;
	wire w_dff_A_oraR3IrY5_0;
	wire w_dff_A_WYhETyT44_0;
	wire w_dff_A_QsK3XZyc0_0;
	wire w_dff_A_1PeAAIgu1_0;
	wire w_dff_A_hF4jqLLM7_0;
	wire w_dff_A_5aH49PcP0_0;
	wire w_dff_A_tTJdCMNL7_0;
	wire w_dff_A_Fwjtbq3s0_0;
	wire w_dff_A_vYpDTAP79_0;
	wire w_dff_A_cUFFlbEi2_0;
	wire w_dff_A_ZFjfCiaE8_0;
	wire w_dff_A_NzUgoClu6_0;
	wire w_dff_A_2QzjacWM0_0;
	wire w_dff_A_41dcNXgg1_0;
	wire w_dff_A_mIbHVo4I9_0;
	wire w_dff_A_L1o6rsPk1_0;
	wire w_dff_A_Z4Azrdl98_0;
	wire w_dff_A_Vaodozu85_0;
	wire w_dff_A_X5zW4CkD5_2;
	wire w_dff_A_OMfjOz0S3_0;
	wire w_dff_A_TDJQUoIB6_0;
	wire w_dff_A_XebOGDqY7_0;
	wire w_dff_A_oCjiPegq0_0;
	wire w_dff_A_wn0Yqp8p2_0;
	wire w_dff_A_kD4AmjX62_0;
	wire w_dff_A_rIoUoEs72_0;
	wire w_dff_A_Hk1b5o689_0;
	wire w_dff_A_Y5soYLYw2_0;
	wire w_dff_A_OKWVZp9u2_0;
	wire w_dff_A_iLpN0RAr4_0;
	wire w_dff_A_olVfXW3u3_0;
	wire w_dff_A_RBXGyFvD1_0;
	wire w_dff_A_0AYV3bIS0_0;
	wire w_dff_A_uaBW9Ssy0_0;
	wire w_dff_A_fF9BKSPy9_0;
	wire w_dff_A_WbnvdjBE7_0;
	wire w_dff_A_2U9O2W6l1_0;
	wire w_dff_A_FtorKECO3_2;
	wire w_dff_A_U6FkGW781_0;
	wire w_dff_A_tB8FVRi90_0;
	wire w_dff_A_zvHMMnu73_0;
	wire w_dff_A_y1yEPVtH6_0;
	wire w_dff_A_pjl44f2L0_0;
	wire w_dff_A_XXla3sAj5_0;
	wire w_dff_A_ihL53V6l3_0;
	wire w_dff_A_YUYTSKZj1_0;
	wire w_dff_A_1qhbX22m1_0;
	wire w_dff_A_NXSUIUMR0_0;
	wire w_dff_A_T7wgGDDF9_0;
	wire w_dff_A_YKX4wmdg3_0;
	wire w_dff_A_yyGzkcoc7_0;
	wire w_dff_A_xX4xaIry1_0;
	wire w_dff_A_vq6Z7ur67_0;
	wire w_dff_A_sN8G1tc00_0;
	wire w_dff_A_EvWttnxa3_2;
	wire w_dff_A_zMc6k8E98_0;
	wire w_dff_A_lKKvZpJl4_0;
	wire w_dff_A_D9XZdQ9X8_0;
	wire w_dff_A_dtLH0Y6l3_0;
	wire w_dff_A_ltLPvjfK4_0;
	wire w_dff_A_kPu6HoWO2_0;
	wire w_dff_A_EPFWUV8h6_0;
	wire w_dff_A_ZMeag6LT5_0;
	wire w_dff_A_5w726Ijp3_0;
	wire w_dff_A_c8WMq0EH1_0;
	wire w_dff_A_X96knW085_0;
	wire w_dff_A_51tvmUTu7_0;
	wire w_dff_A_6ek4ZFL08_0;
	wire w_dff_A_phJnpuEk4_0;
	wire w_dff_A_TLmwHIhE1_2;
	wire w_dff_A_nXGdspfK3_0;
	wire w_dff_A_FIX0YiuS9_0;
	wire w_dff_A_5O5Qqwkd4_0;
	wire w_dff_A_29hlMrLC8_0;
	wire w_dff_A_so3Uc0T45_0;
	wire w_dff_A_HvjJnEIJ6_0;
	wire w_dff_A_K5Sk7pRt4_0;
	wire w_dff_A_Z9yG4cs03_0;
	wire w_dff_A_O7tpWd0y7_0;
	wire w_dff_A_L88DLSrW3_0;
	wire w_dff_A_9m8JFDcT3_0;
	wire w_dff_A_dixSqDUG8_0;
	wire w_dff_A_np4nDYGT0_2;
	wire w_dff_A_OQNzrkQT3_0;
	wire w_dff_A_yplJ0Ykl3_0;
	wire w_dff_A_fx1eFLLd6_0;
	wire w_dff_A_sxW095fL2_0;
	wire w_dff_A_7NrR5XjK2_0;
	wire w_dff_A_g8o6yiBn1_0;
	wire w_dff_A_VeNVzcJc0_0;
	wire w_dff_A_rvvPdYNb0_0;
	wire w_dff_A_fOgzutYn2_0;
	wire w_dff_A_40PEDUQR7_0;
	wire w_dff_A_MxA6KRqk3_2;
	wire w_dff_A_qty7FCa43_0;
	wire w_dff_A_rz1JjpZ09_0;
	wire w_dff_A_8YYLDw7X4_0;
	wire w_dff_A_gEc8NJbU0_0;
	wire w_dff_A_TkHTf4Y76_0;
	wire w_dff_A_hQAustIc1_0;
	wire w_dff_A_IGsU7fHb8_0;
	wire w_dff_A_LOpn4Y7Y4_0;
	wire w_dff_A_vaZ8kvun7_2;
	wire w_dff_A_fl4lL1AN3_0;
	wire w_dff_A_UiiR4dBg9_0;
	wire w_dff_A_4PeI1Z3o0_0;
	wire w_dff_A_bDg38os87_0;
	wire w_dff_A_AbQW1K2o9_0;
	wire w_dff_A_W4tUHAVz7_0;
	wire w_dff_A_QTxU36lP3_2;
	wire w_dff_A_SdRFDCEB9_0;
	wire w_dff_A_DUo9KVGb3_0;
	wire w_dff_A_gCpavY280_0;
	wire w_dff_A_nISZq5Dm2_0;
	wire w_dff_A_emw7PjXC7_2;
	wire w_dff_A_Ng3v1Jn62_0;
	wire w_dff_A_SZ5hnu3S8_0;
	wire w_dff_A_roQXFJyg9_2;
	jand g0000(.dina(w_G273gat_7[1]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G290gat_7[2]),.dinb(w_G18gat_7[1]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_n65_0[1]),.dinb(w_G545gat_0),.dout(n66),.clk(gclk));
	jnot g0003(.din(w_n66_0[1]),.dout(n67),.clk(gclk));
	jnot g0004(.din(w_G18gat_7[0]),.dout(n68),.clk(gclk));
	jnot g0005(.din(w_G273gat_7[0]),.dout(n69),.clk(gclk));
	jor g0006(.dina(w_n69_0[1]),.dinb(n68),.dout(n70),.clk(gclk));
	jnot g0007(.din(w_n70_0[1]),.dout(n71),.clk(gclk));
	jand g0008(.dina(w_G290gat_7[1]),.dinb(w_G1gat_7[0]),.dout(n72),.clk(gclk));
	jor g0009(.dina(n72),.dinb(n71),.dout(n73),.clk(gclk));
	jand g0010(.dina(n73),.dinb(w_n67_0[1]),.dout(w_dff_A_HFwDfpPm3_2),.clk(gclk));
	jand g0011(.dina(w_G307gat_7[1]),.dinb(w_G1gat_6[2]),.dout(n75),.clk(gclk));
	jnot g0012(.din(w_n75_0[1]),.dout(n76),.clk(gclk));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G290gat_7[0]),.dout(n78),.clk(gclk));
	jor g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79),.clk(gclk));
	jor g0016(.dina(n79),.dinb(w_n70_0[0]),.dout(n80),.clk(gclk));
	jand g0017(.dina(w_G273gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jor g0018(.dina(n81),.dinb(w_n65_0[0]),.dout(n82),.clk(gclk));
	jand g0019(.dina(n82),.dinb(w_n80_0[2]),.dout(n83),.clk(gclk));
	jxor g0020(.dina(w_n83_0[1]),.dinb(w_n67_0[0]),.dout(n84),.clk(gclk));
	jxor g0021(.dina(w_n84_0[1]),.dinb(w_dff_B_8vD6sN1d2_1),.dout(w_dff_A_RsDoFRkE0_2),.clk(gclk));
	jand g0022(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n86),.clk(gclk));
	jnot g0023(.din(w_n86_0[1]),.dout(n87),.clk(gclk));
	jor g0024(.dina(w_n83_0[0]),.dinb(w_n66_0[0]),.dout(n88),.clk(gclk));
	jor g0025(.dina(w_n84_0[0]),.dinb(w_n75_0[0]),.dout(n89),.clk(gclk));
	jand g0026(.dina(n89),.dinb(w_dff_B_hKWuVKxP1_1),.dout(n90),.clk(gclk));
	jand g0027(.dina(w_G307gat_7[0]),.dinb(w_G18gat_6[2]),.dout(n91),.clk(gclk));
	jnot g0028(.din(w_n91_0[1]),.dout(n92),.clk(gclk));
	jnot g0029(.din(w_n80_0[1]),.dout(n93),.clk(gclk));
	jor g0030(.dina(w_n69_0[0]),.dinb(w_n77_0[0]),.dout(n94),.clk(gclk));
	jnot g0031(.din(w_G52gat_7[2]),.dout(n95),.clk(gclk));
	jor g0032(.dina(w_n78_0[0]),.dinb(n95),.dout(n96),.clk(gclk));
	jor g0033(.dina(n96),.dinb(n94),.dout(n97),.clk(gclk));
	jand g0034(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G273gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jor g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100),.clk(gclk));
	jand g0037(.dina(n100),.dinb(w_n97_0[1]),.dout(n101),.clk(gclk));
	jxor g0038(.dina(w_n101_0[2]),.dinb(w_n93_0[1]),.dout(n102),.clk(gclk));
	jxor g0039(.dina(n102),.dinb(n92),.dout(n103),.clk(gclk));
	jxor g0040(.dina(w_n103_0[1]),.dinb(w_n90_0[1]),.dout(n104),.clk(gclk));
	jxor g0041(.dina(w_n104_0[1]),.dinb(w_dff_B_VEfEsqjZ4_1),.dout(w_dff_A_1xLXBDUh1_2),.clk(gclk));
	jand g0042(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n106),.clk(gclk));
	jnot g0043(.din(w_n106_0[1]),.dout(n107),.clk(gclk));
	jnot g0044(.din(w_n103_0[0]),.dout(n108),.clk(gclk));
	jor g0045(.dina(n108),.dinb(w_n90_0[0]),.dout(n109),.clk(gclk));
	jor g0046(.dina(w_n104_0[0]),.dinb(w_n86_0[0]),.dout(n110),.clk(gclk));
	jand g0047(.dina(n110),.dinb(w_dff_B_zyUCrIaE8_1),.dout(n111),.clk(gclk));
	jand g0048(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n112),.clk(gclk));
	jnot g0049(.din(w_n112_0[1]),.dout(n113),.clk(gclk));
	jor g0050(.dina(w_n101_0[1]),.dinb(w_n93_0[0]),.dout(n114),.clk(gclk));
	jxor g0051(.dina(w_n101_0[0]),.dinb(w_n80_0[0]),.dout(n115),.clk(gclk));
	jor g0052(.dina(n115),.dinb(w_n91_0[0]),.dout(n116),.clk(gclk));
	jand g0053(.dina(n116),.dinb(n114),.dout(n117),.clk(gclk));
	jand g0054(.dina(w_G307gat_6[2]),.dinb(w_G35gat_6[2]),.dout(n118),.clk(gclk));
	jnot g0055(.din(n118),.dout(n119),.clk(gclk));
	jnot g0056(.din(w_n97_0[0]),.dout(n120),.clk(gclk));
	jand g0057(.dina(w_G290gat_6[1]),.dinb(w_G69gat_7[1]),.dout(n121),.clk(gclk));
	jand g0058(.dina(w_n121_0[1]),.dinb(w_n99_0[0]),.dout(n122),.clk(gclk));
	jnot g0059(.din(w_n122_0[1]),.dout(n123),.clk(gclk));
	jand g0060(.dina(w_G290gat_6[0]),.dinb(w_G52gat_7[0]),.dout(n124),.clk(gclk));
	jand g0061(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n125),.clk(gclk));
	jor g0062(.dina(w_n125_0[1]),.dinb(n124),.dout(n126),.clk(gclk));
	jand g0063(.dina(n126),.dinb(w_n123_0[1]),.dout(n127),.clk(gclk));
	jxor g0064(.dina(w_n127_0[1]),.dinb(w_n120_0[1]),.dout(n128),.clk(gclk));
	jxor g0065(.dina(w_n128_0[1]),.dinb(w_n119_0[1]),.dout(n129),.clk(gclk));
	jnot g0066(.din(w_n129_0[1]),.dout(n130),.clk(gclk));
	jxor g0067(.dina(w_n130_0[1]),.dinb(w_n117_0[2]),.dout(n131),.clk(gclk));
	jxor g0068(.dina(n131),.dinb(n113),.dout(n132),.clk(gclk));
	jxor g0069(.dina(w_n132_0[1]),.dinb(w_n111_0[1]),.dout(n133),.clk(gclk));
	jxor g0070(.dina(w_n133_0[1]),.dinb(w_dff_B_QGLP9ZNw7_1),.dout(w_dff_A_TeLedrld7_2),.clk(gclk));
	jand g0071(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n135),.clk(gclk));
	jnot g0072(.din(w_n135_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(w_n132_0[0]),.dout(n137),.clk(gclk));
	jor g0074(.dina(n137),.dinb(w_n111_0[0]),.dout(n138),.clk(gclk));
	jor g0075(.dina(w_n133_0[0]),.dinb(w_n106_0[0]),.dout(n139),.clk(gclk));
	jand g0076(.dina(n139),.dinb(w_dff_B_GrrYRaG21_1),.dout(n140),.clk(gclk));
	jand g0077(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n141),.clk(gclk));
	jnot g0078(.din(w_n141_0[1]),.dout(n142),.clk(gclk));
	jor g0079(.dina(w_n130_0[0]),.dinb(w_n117_0[1]),.dout(n143),.clk(gclk));
	jxor g0080(.dina(w_n129_0[0]),.dinb(w_n117_0[0]),.dout(n144),.clk(gclk));
	jor g0081(.dina(n144),.dinb(w_n112_0[0]),.dout(n145),.clk(gclk));
	jand g0082(.dina(n145),.dinb(n143),.dout(n146),.clk(gclk));
	jand g0083(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n147),.clk(gclk));
	jnot g0084(.din(n147),.dout(n148),.clk(gclk));
	jor g0085(.dina(w_n127_0[0]),.dinb(w_n120_0[0]),.dout(n149),.clk(gclk));
	jnot g0086(.din(n149),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_n128_0[0]),.dinb(w_n119_0[0]),.dout(n151),.clk(gclk));
	jor g0088(.dina(n151),.dinb(n150),.dout(n152),.clk(gclk));
	jand g0089(.dina(w_G307gat_6[1]),.dinb(w_G52gat_6[2]),.dout(n153),.clk(gclk));
	jnot g0090(.din(n153),.dout(n154),.clk(gclk));
	jand g0091(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n155),.clk(gclk));
	jand g0092(.dina(w_n155_0[1]),.dinb(w_n125_0[0]),.dout(n156),.clk(gclk));
	jnot g0093(.din(w_n156_0[1]),.dout(n157),.clk(gclk));
	jand g0094(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n158),.clk(gclk));
	jor g0095(.dina(w_n158_0[1]),.dinb(w_n121_0[0]),.dout(n159),.clk(gclk));
	jand g0096(.dina(n159),.dinb(w_n157_0[1]),.dout(n160),.clk(gclk));
	jxor g0097(.dina(w_n160_0[1]),.dinb(w_n122_0[0]),.dout(n161),.clk(gclk));
	jxor g0098(.dina(w_n161_0[1]),.dinb(w_n154_0[1]),.dout(n162),.clk(gclk));
	jxor g0099(.dina(w_n162_0[1]),.dinb(w_n152_0[1]),.dout(n163),.clk(gclk));
	jxor g0100(.dina(w_n163_0[1]),.dinb(w_n148_0[1]),.dout(n164),.clk(gclk));
	jnot g0101(.din(w_n164_0[1]),.dout(n165),.clk(gclk));
	jxor g0102(.dina(w_n165_0[1]),.dinb(w_n146_0[2]),.dout(n166),.clk(gclk));
	jxor g0103(.dina(n166),.dinb(n142),.dout(n167),.clk(gclk));
	jxor g0104(.dina(w_n167_0[1]),.dinb(w_n140_0[1]),.dout(n168),.clk(gclk));
	jxor g0105(.dina(w_n168_0[1]),.dinb(w_dff_B_zKlZiXNS1_1),.dout(w_dff_A_TwM7lXbz1_2),.clk(gclk));
	jand g0106(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n170),.clk(gclk));
	jnot g0107(.din(w_n170_0[1]),.dout(n171),.clk(gclk));
	jnot g0108(.din(w_n167_0[0]),.dout(n172),.clk(gclk));
	jor g0109(.dina(n172),.dinb(w_n140_0[0]),.dout(n173),.clk(gclk));
	jor g0110(.dina(w_n168_0[0]),.dinb(w_n135_0[0]),.dout(n174),.clk(gclk));
	jand g0111(.dina(n174),.dinb(w_dff_B_WOBZxwkd3_1),.dout(n175),.clk(gclk));
	jand g0112(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n176),.clk(gclk));
	jnot g0113(.din(w_n176_0[1]),.dout(n177),.clk(gclk));
	jor g0114(.dina(w_n165_0[0]),.dinb(w_n146_0[1]),.dout(n178),.clk(gclk));
	jxor g0115(.dina(w_n164_0[0]),.dinb(w_n146_0[0]),.dout(n179),.clk(gclk));
	jor g0116(.dina(n179),.dinb(w_n141_0[0]),.dout(n180),.clk(gclk));
	jand g0117(.dina(n180),.dinb(n178),.dout(n181),.clk(gclk));
	jand g0118(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n182),.clk(gclk));
	jnot g0119(.din(n182),.dout(n183),.clk(gclk));
	jand g0120(.dina(w_n162_0[0]),.dinb(w_n152_0[0]),.dout(n184),.clk(gclk));
	jand g0121(.dina(w_n163_0[0]),.dinb(w_n148_0[0]),.dout(n185),.clk(gclk));
	jor g0122(.dina(n185),.dinb(n184),.dout(n186),.clk(gclk));
	jand g0123(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n187),.clk(gclk));
	jnot g0124(.din(n187),.dout(n188),.clk(gclk));
	jnot g0125(.din(w_n160_0[0]),.dout(n189),.clk(gclk));
	jand g0126(.dina(n189),.dinb(w_n123_0[0]),.dout(n190),.clk(gclk));
	jand g0127(.dina(w_n161_0[0]),.dinb(w_n154_0[0]),.dout(n191),.clk(gclk));
	jor g0128(.dina(n191),.dinb(n190),.dout(n192),.clk(gclk));
	jand g0129(.dina(w_G307gat_6[0]),.dinb(w_G69gat_6[2]),.dout(n193),.clk(gclk));
	jnot g0130(.din(n193),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n195),.clk(gclk));
	jand g0132(.dina(w_n195_0[1]),.dinb(w_n158_0[0]),.dout(n196),.clk(gclk));
	jnot g0133(.din(w_n196_0[2]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n198),.clk(gclk));
	jor g0135(.dina(w_n198_0[1]),.dinb(w_n155_0[0]),.dout(n199),.clk(gclk));
	jand g0136(.dina(n199),.dinb(n197),.dout(n200),.clk(gclk));
	jxor g0137(.dina(w_n200_0[1]),.dinb(w_n156_0[0]),.dout(n201),.clk(gclk));
	jxor g0138(.dina(w_n201_0[1]),.dinb(w_n194_0[1]),.dout(n202),.clk(gclk));
	jxor g0139(.dina(w_n202_0[1]),.dinb(w_n192_0[1]),.dout(n203),.clk(gclk));
	jxor g0140(.dina(w_n203_0[1]),.dinb(w_n188_0[1]),.dout(n204),.clk(gclk));
	jxor g0141(.dina(w_n204_0[1]),.dinb(w_n186_0[1]),.dout(n205),.clk(gclk));
	jxor g0142(.dina(w_n205_0[1]),.dinb(w_n183_0[1]),.dout(n206),.clk(gclk));
	jnot g0143(.din(w_n206_0[1]),.dout(n207),.clk(gclk));
	jxor g0144(.dina(w_n207_0[1]),.dinb(w_n181_0[2]),.dout(n208),.clk(gclk));
	jxor g0145(.dina(n208),.dinb(n177),.dout(n209),.clk(gclk));
	jxor g0146(.dina(w_n209_0[1]),.dinb(w_n175_0[1]),.dout(n210),.clk(gclk));
	jxor g0147(.dina(w_n210_0[1]),.dinb(w_dff_B_GF8o5Vdy5_1),.dout(w_dff_A_vUFKz7gI5_2),.clk(gclk));
	jand g0148(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n212),.clk(gclk));
	jnot g0149(.din(w_n212_0[1]),.dout(n213),.clk(gclk));
	jnot g0150(.din(w_n209_0[0]),.dout(n214),.clk(gclk));
	jor g0151(.dina(n214),.dinb(w_n175_0[0]),.dout(n215),.clk(gclk));
	jor g0152(.dina(w_n210_0[0]),.dinb(w_n170_0[0]),.dout(n216),.clk(gclk));
	jand g0153(.dina(n216),.dinb(w_dff_B_SFCaJsrj1_1),.dout(n217),.clk(gclk));
	jand g0154(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n218),.clk(gclk));
	jnot g0155(.din(w_n218_0[1]),.dout(n219),.clk(gclk));
	jor g0156(.dina(w_n207_0[0]),.dinb(w_n181_0[1]),.dout(n220),.clk(gclk));
	jxor g0157(.dina(w_n206_0[0]),.dinb(w_n181_0[0]),.dout(n221),.clk(gclk));
	jor g0158(.dina(n221),.dinb(w_n176_0[0]),.dout(n222),.clk(gclk));
	jand g0159(.dina(n222),.dinb(n220),.dout(n223),.clk(gclk));
	jand g0160(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n224),.clk(gclk));
	jnot g0161(.din(n224),.dout(n225),.clk(gclk));
	jand g0162(.dina(w_n204_0[0]),.dinb(w_n186_0[0]),.dout(n226),.clk(gclk));
	jand g0163(.dina(w_n205_0[0]),.dinb(w_n183_0[0]),.dout(n227),.clk(gclk));
	jor g0164(.dina(n227),.dinb(n226),.dout(n228),.clk(gclk));
	jand g0165(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n229),.clk(gclk));
	jnot g0166(.din(n229),.dout(n230),.clk(gclk));
	jand g0167(.dina(w_n202_0[0]),.dinb(w_n192_0[0]),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_n203_0[0]),.dinb(w_n188_0[0]),.dout(n232),.clk(gclk));
	jor g0169(.dina(n232),.dinb(n231),.dout(n233),.clk(gclk));
	jand g0170(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n234),.clk(gclk));
	jnot g0171(.din(n234),.dout(n235),.clk(gclk));
	jnot g0172(.din(w_n200_0[0]),.dout(n236),.clk(gclk));
	jand g0173(.dina(n236),.dinb(w_n157_0[0]),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_n201_0[0]),.dinb(w_n194_0[0]),.dout(n238),.clk(gclk));
	jor g0175(.dina(n238),.dinb(n237),.dout(n239),.clk(gclk));
	jand g0176(.dina(w_G307gat_5[2]),.dinb(w_G86gat_6[2]),.dout(n240),.clk(gclk));
	jnot g0177(.din(n240),.dout(n241),.clk(gclk));
	jand g0178(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n242),.clk(gclk));
	jand g0179(.dina(w_n242_0[1]),.dinb(w_n198_0[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(w_n243_0[2]),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n245),.clk(gclk));
	jor g0182(.dina(w_n245_0[1]),.dinb(w_n195_0[0]),.dout(n246),.clk(gclk));
	jand g0183(.dina(n246),.dinb(n244),.dout(n247),.clk(gclk));
	jxor g0184(.dina(w_n247_0[1]),.dinb(w_n196_0[1]),.dout(n248),.clk(gclk));
	jxor g0185(.dina(w_n248_0[1]),.dinb(w_n241_0[1]),.dout(n249),.clk(gclk));
	jxor g0186(.dina(w_n249_0[1]),.dinb(w_n239_0[1]),.dout(n250),.clk(gclk));
	jxor g0187(.dina(w_n250_0[1]),.dinb(w_n235_0[1]),.dout(n251),.clk(gclk));
	jxor g0188(.dina(w_n251_0[1]),.dinb(w_n233_0[1]),.dout(n252),.clk(gclk));
	jxor g0189(.dina(w_n252_0[1]),.dinb(w_n230_0[1]),.dout(n253),.clk(gclk));
	jxor g0190(.dina(w_n253_0[1]),.dinb(w_n228_0[1]),.dout(n254),.clk(gclk));
	jxor g0191(.dina(w_n254_0[1]),.dinb(w_n225_0[1]),.dout(n255),.clk(gclk));
	jnot g0192(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jxor g0193(.dina(w_n256_0[1]),.dinb(w_n223_0[2]),.dout(n257),.clk(gclk));
	jxor g0194(.dina(n257),.dinb(n219),.dout(n258),.clk(gclk));
	jxor g0195(.dina(w_n258_0[1]),.dinb(w_n217_0[1]),.dout(n259),.clk(gclk));
	jxor g0196(.dina(w_n259_0[1]),.dinb(w_dff_B_789OLFB94_1),.dout(w_dff_A_x5iNlZpF9_2),.clk(gclk));
	jand g0197(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n261),.clk(gclk));
	jnot g0198(.din(w_n261_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(w_n258_0[0]),.dout(n263),.clk(gclk));
	jor g0200(.dina(n263),.dinb(w_n217_0[0]),.dout(n264),.clk(gclk));
	jor g0201(.dina(w_n259_0[0]),.dinb(w_n212_0[0]),.dout(n265),.clk(gclk));
	jand g0202(.dina(n265),.dinb(w_dff_B_ZDi3jBiT2_1),.dout(n266),.clk(gclk));
	jand g0203(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n267),.clk(gclk));
	jnot g0204(.din(w_n267_0[1]),.dout(n268),.clk(gclk));
	jor g0205(.dina(w_n256_0[0]),.dinb(w_n223_0[1]),.dout(n269),.clk(gclk));
	jxor g0206(.dina(w_n255_0[0]),.dinb(w_n223_0[0]),.dout(n270),.clk(gclk));
	jor g0207(.dina(n270),.dinb(w_n218_0[0]),.dout(n271),.clk(gclk));
	jand g0208(.dina(n271),.dinb(n269),.dout(n272),.clk(gclk));
	jand g0209(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n273),.clk(gclk));
	jnot g0210(.din(n273),.dout(n274),.clk(gclk));
	jand g0211(.dina(w_n253_0[0]),.dinb(w_n228_0[0]),.dout(n275),.clk(gclk));
	jand g0212(.dina(w_n254_0[0]),.dinb(w_n225_0[0]),.dout(n276),.clk(gclk));
	jor g0213(.dina(n276),.dinb(n275),.dout(n277),.clk(gclk));
	jand g0214(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n278),.clk(gclk));
	jnot g0215(.din(n278),.dout(n279),.clk(gclk));
	jand g0216(.dina(w_n251_0[0]),.dinb(w_n233_0[0]),.dout(n280),.clk(gclk));
	jand g0217(.dina(w_n252_0[0]),.dinb(w_n230_0[0]),.dout(n281),.clk(gclk));
	jor g0218(.dina(n281),.dinb(n280),.dout(n282),.clk(gclk));
	jand g0219(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(n283),.dout(n284),.clk(gclk));
	jand g0221(.dina(w_n249_0[0]),.dinb(w_n239_0[0]),.dout(n285),.clk(gclk));
	jand g0222(.dina(w_n250_0[0]),.dinb(w_n235_0[0]),.dout(n286),.clk(gclk));
	jor g0223(.dina(n286),.dinb(n285),.dout(n287),.clk(gclk));
	jand g0224(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n288),.clk(gclk));
	jnot g0225(.din(n288),.dout(n289),.clk(gclk));
	jor g0226(.dina(w_n247_0[0]),.dinb(w_n196_0[0]),.dout(n290),.clk(gclk));
	jnot g0227(.din(n290),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n248_0[0]),.dinb(w_n241_0[0]),.dout(n292),.clk(gclk));
	jor g0229(.dina(n292),.dinb(n291),.dout(n293),.clk(gclk));
	jand g0230(.dina(w_G307gat_5[1]),.dinb(w_G103gat_6[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n296_0[1]),.dinb(w_n245_0[0]),.dout(n297),.clk(gclk));
	jnot g0234(.din(w_n297_0[2]),.dout(n298),.clk(gclk));
	jand g0235(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n299),.clk(gclk));
	jor g0236(.dina(w_n299_0[1]),.dinb(w_n242_0[0]),.dout(n300),.clk(gclk));
	jand g0237(.dina(n300),.dinb(n298),.dout(n301),.clk(gclk));
	jxor g0238(.dina(w_n301_0[1]),.dinb(w_n243_0[1]),.dout(n302),.clk(gclk));
	jxor g0239(.dina(w_n302_0[1]),.dinb(w_n295_0[1]),.dout(n303),.clk(gclk));
	jxor g0240(.dina(w_n303_0[1]),.dinb(w_n293_0[1]),.dout(n304),.clk(gclk));
	jxor g0241(.dina(w_n304_0[1]),.dinb(w_n289_0[1]),.dout(n305),.clk(gclk));
	jxor g0242(.dina(w_n305_0[1]),.dinb(w_n287_0[1]),.dout(n306),.clk(gclk));
	jxor g0243(.dina(w_n306_0[1]),.dinb(w_n284_0[1]),.dout(n307),.clk(gclk));
	jxor g0244(.dina(w_n307_0[1]),.dinb(w_n282_0[1]),.dout(n308),.clk(gclk));
	jxor g0245(.dina(w_n308_0[1]),.dinb(w_n279_0[1]),.dout(n309),.clk(gclk));
	jxor g0246(.dina(w_n309_0[1]),.dinb(w_n277_0[1]),.dout(n310),.clk(gclk));
	jxor g0247(.dina(w_n310_0[1]),.dinb(w_n274_0[1]),.dout(n311),.clk(gclk));
	jnot g0248(.din(w_n311_0[1]),.dout(n312),.clk(gclk));
	jxor g0249(.dina(w_n312_0[1]),.dinb(w_n272_0[2]),.dout(n313),.clk(gclk));
	jxor g0250(.dina(n313),.dinb(n268),.dout(n314),.clk(gclk));
	jxor g0251(.dina(w_n314_0[1]),.dinb(w_n266_0[1]),.dout(n315),.clk(gclk));
	jxor g0252(.dina(w_n315_0[1]),.dinb(w_dff_B_fQ9WsX7z0_1),.dout(w_dff_A_tlP6TWHP5_2),.clk(gclk));
	jand g0253(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n317),.clk(gclk));
	jnot g0254(.din(w_n317_0[1]),.dout(n318),.clk(gclk));
	jnot g0255(.din(w_n314_0[0]),.dout(n319),.clk(gclk));
	jor g0256(.dina(n319),.dinb(w_n266_0[0]),.dout(n320),.clk(gclk));
	jor g0257(.dina(w_n315_0[0]),.dinb(w_n261_0[0]),.dout(n321),.clk(gclk));
	jand g0258(.dina(n321),.dinb(w_dff_B_x30379n46_1),.dout(n322),.clk(gclk));
	jand g0259(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n323),.clk(gclk));
	jnot g0260(.din(w_n323_0[1]),.dout(n324),.clk(gclk));
	jor g0261(.dina(w_n312_0[0]),.dinb(w_n272_0[1]),.dout(n325),.clk(gclk));
	jxor g0262(.dina(w_n311_0[0]),.dinb(w_n272_0[0]),.dout(n326),.clk(gclk));
	jor g0263(.dina(n326),.dinb(w_n267_0[0]),.dout(n327),.clk(gclk));
	jand g0264(.dina(n327),.dinb(n325),.dout(n328),.clk(gclk));
	jand g0265(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n329),.clk(gclk));
	jnot g0266(.din(n329),.dout(n330),.clk(gclk));
	jand g0267(.dina(w_n309_0[0]),.dinb(w_n277_0[0]),.dout(n331),.clk(gclk));
	jand g0268(.dina(w_n310_0[0]),.dinb(w_n274_0[0]),.dout(n332),.clk(gclk));
	jor g0269(.dina(n332),.dinb(n331),.dout(n333),.clk(gclk));
	jand g0270(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n334),.clk(gclk));
	jnot g0271(.din(n334),.dout(n335),.clk(gclk));
	jand g0272(.dina(w_n307_0[0]),.dinb(w_n282_0[0]),.dout(n336),.clk(gclk));
	jand g0273(.dina(w_n308_0[0]),.dinb(w_n279_0[0]),.dout(n337),.clk(gclk));
	jor g0274(.dina(n337),.dinb(n336),.dout(n338),.clk(gclk));
	jand g0275(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n339),.clk(gclk));
	jnot g0276(.din(n339),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_n305_0[0]),.dinb(w_n287_0[0]),.dout(n341),.clk(gclk));
	jand g0278(.dina(w_n306_0[0]),.dinb(w_n284_0[0]),.dout(n342),.clk(gclk));
	jor g0279(.dina(n342),.dinb(n341),.dout(n343),.clk(gclk));
	jand g0280(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n344),.clk(gclk));
	jnot g0281(.din(n344),.dout(n345),.clk(gclk));
	jand g0282(.dina(w_n303_0[0]),.dinb(w_n293_0[0]),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_n304_0[0]),.dinb(w_n289_0[0]),.dout(n347),.clk(gclk));
	jor g0284(.dina(n347),.dinb(n346),.dout(n348),.clk(gclk));
	jand g0285(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n349),.clk(gclk));
	jnot g0286(.din(n349),.dout(n350),.clk(gclk));
	jor g0287(.dina(w_n301_0[0]),.dinb(w_n243_0[0]),.dout(n351),.clk(gclk));
	jnot g0288(.din(n351),.dout(n352),.clk(gclk));
	jand g0289(.dina(w_n302_0[0]),.dinb(w_n295_0[0]),.dout(n353),.clk(gclk));
	jor g0290(.dina(n353),.dinb(n352),.dout(n354),.clk(gclk));
	jand g0291(.dina(w_G307gat_5[0]),.dinb(w_G120gat_6[2]),.dout(n355),.clk(gclk));
	jnot g0292(.din(n355),.dout(n356),.clk(gclk));
	jand g0293(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n357),.clk(gclk));
	jand g0294(.dina(w_n357_0[1]),.dinb(w_n299_0[0]),.dout(n358),.clk(gclk));
	jnot g0295(.din(w_n358_0[2]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n360),.clk(gclk));
	jor g0297(.dina(w_n360_0[1]),.dinb(w_n296_0[0]),.dout(n361),.clk(gclk));
	jand g0298(.dina(n361),.dinb(n359),.dout(n362),.clk(gclk));
	jxor g0299(.dina(w_n362_0[1]),.dinb(w_n297_0[1]),.dout(n363),.clk(gclk));
	jxor g0300(.dina(w_n363_0[1]),.dinb(w_n356_0[1]),.dout(n364),.clk(gclk));
	jxor g0301(.dina(w_n364_0[1]),.dinb(w_n354_0[1]),.dout(n365),.clk(gclk));
	jxor g0302(.dina(w_n365_0[1]),.dinb(w_n350_0[1]),.dout(n366),.clk(gclk));
	jxor g0303(.dina(w_n366_0[1]),.dinb(w_n348_0[1]),.dout(n367),.clk(gclk));
	jxor g0304(.dina(w_n367_0[1]),.dinb(w_n345_0[1]),.dout(n368),.clk(gclk));
	jxor g0305(.dina(w_n368_0[1]),.dinb(w_n343_0[1]),.dout(n369),.clk(gclk));
	jxor g0306(.dina(w_n369_0[1]),.dinb(w_n340_0[1]),.dout(n370),.clk(gclk));
	jxor g0307(.dina(w_n370_0[1]),.dinb(w_n338_0[1]),.dout(n371),.clk(gclk));
	jxor g0308(.dina(w_n371_0[1]),.dinb(w_n335_0[1]),.dout(n372),.clk(gclk));
	jxor g0309(.dina(w_n372_0[1]),.dinb(w_n333_0[1]),.dout(n373),.clk(gclk));
	jxor g0310(.dina(w_n373_0[1]),.dinb(w_n330_0[1]),.dout(n374),.clk(gclk));
	jnot g0311(.din(w_n374_0[1]),.dout(n375),.clk(gclk));
	jxor g0312(.dina(w_n375_0[1]),.dinb(w_n328_0[2]),.dout(n376),.clk(gclk));
	jxor g0313(.dina(n376),.dinb(n324),.dout(n377),.clk(gclk));
	jxor g0314(.dina(w_n377_0[1]),.dinb(w_n322_0[1]),.dout(n378),.clk(gclk));
	jxor g0315(.dina(w_n378_0[1]),.dinb(w_dff_B_OHdJphC50_1),.dout(w_dff_A_HcHGc8GI5_2),.clk(gclk));
	jand g0316(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n380),.clk(gclk));
	jnot g0317(.din(w_n380_0[1]),.dout(n381),.clk(gclk));
	jnot g0318(.din(w_n377_0[0]),.dout(n382),.clk(gclk));
	jor g0319(.dina(n382),.dinb(w_n322_0[0]),.dout(n383),.clk(gclk));
	jor g0320(.dina(w_n378_0[0]),.dinb(w_n317_0[0]),.dout(n384),.clk(gclk));
	jand g0321(.dina(n384),.dinb(w_dff_B_8cIcvORO0_1),.dout(n385),.clk(gclk));
	jand g0322(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n386),.clk(gclk));
	jnot g0323(.din(w_n386_0[1]),.dout(n387),.clk(gclk));
	jor g0324(.dina(w_n375_0[0]),.dinb(w_n328_0[1]),.dout(n388),.clk(gclk));
	jxor g0325(.dina(w_n374_0[0]),.dinb(w_n328_0[0]),.dout(n389),.clk(gclk));
	jor g0326(.dina(n389),.dinb(w_n323_0[0]),.dout(n390),.clk(gclk));
	jand g0327(.dina(n390),.dinb(n388),.dout(n391),.clk(gclk));
	jand g0328(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n392),.clk(gclk));
	jnot g0329(.din(n392),.dout(n393),.clk(gclk));
	jand g0330(.dina(w_n372_0[0]),.dinb(w_n333_0[0]),.dout(n394),.clk(gclk));
	jand g0331(.dina(w_n373_0[0]),.dinb(w_n330_0[0]),.dout(n395),.clk(gclk));
	jor g0332(.dina(n395),.dinb(n394),.dout(n396),.clk(gclk));
	jand g0333(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n397),.clk(gclk));
	jnot g0334(.din(n397),.dout(n398),.clk(gclk));
	jand g0335(.dina(w_n370_0[0]),.dinb(w_n338_0[0]),.dout(n399),.clk(gclk));
	jand g0336(.dina(w_n371_0[0]),.dinb(w_n335_0[0]),.dout(n400),.clk(gclk));
	jor g0337(.dina(n400),.dinb(n399),.dout(n401),.clk(gclk));
	jand g0338(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n402),.clk(gclk));
	jnot g0339(.din(n402),.dout(n403),.clk(gclk));
	jand g0340(.dina(w_n368_0[0]),.dinb(w_n343_0[0]),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_n369_0[0]),.dinb(w_n340_0[0]),.dout(n405),.clk(gclk));
	jor g0342(.dina(n405),.dinb(n404),.dout(n406),.clk(gclk));
	jand g0343(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n407),.clk(gclk));
	jnot g0344(.din(n407),.dout(n408),.clk(gclk));
	jand g0345(.dina(w_n366_0[0]),.dinb(w_n348_0[0]),.dout(n409),.clk(gclk));
	jand g0346(.dina(w_n367_0[0]),.dinb(w_n345_0[0]),.dout(n410),.clk(gclk));
	jor g0347(.dina(n410),.dinb(n409),.dout(n411),.clk(gclk));
	jand g0348(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n412),.clk(gclk));
	jnot g0349(.din(n412),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n364_0[0]),.dinb(w_n354_0[0]),.dout(n414),.clk(gclk));
	jand g0351(.dina(w_n365_0[0]),.dinb(w_n350_0[0]),.dout(n415),.clk(gclk));
	jor g0352(.dina(n415),.dinb(n414),.dout(n416),.clk(gclk));
	jand g0353(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n417),.clk(gclk));
	jnot g0354(.din(n417),.dout(n418),.clk(gclk));
	jor g0355(.dina(w_n362_0[0]),.dinb(w_n297_0[0]),.dout(n419),.clk(gclk));
	jand g0356(.dina(w_n363_0[0]),.dinb(w_n356_0[0]),.dout(n420),.clk(gclk));
	jnot g0357(.din(n420),.dout(n421),.clk(gclk));
	jand g0358(.dina(n421),.dinb(n419),.dout(n422),.clk(gclk));
	jnot g0359(.din(n422),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_G307gat_4[2]),.dinb(w_G137gat_6[2]),.dout(n424),.clk(gclk));
	jnot g0361(.din(n424),.dout(n425),.clk(gclk));
	jand g0362(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n426),.clk(gclk));
	jand g0363(.dina(w_n426_0[1]),.dinb(w_n360_0[0]),.dout(n427),.clk(gclk));
	jnot g0364(.din(w_n427_0[2]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n429),.clk(gclk));
	jor g0366(.dina(w_n429_0[1]),.dinb(w_n357_0[0]),.dout(n430),.clk(gclk));
	jand g0367(.dina(n430),.dinb(n428),.dout(n431),.clk(gclk));
	jxor g0368(.dina(w_n431_0[1]),.dinb(w_n358_0[1]),.dout(n432),.clk(gclk));
	jxor g0369(.dina(w_n432_0[1]),.dinb(w_n425_0[1]),.dout(n433),.clk(gclk));
	jxor g0370(.dina(w_n433_0[1]),.dinb(w_n423_0[1]),.dout(n434),.clk(gclk));
	jxor g0371(.dina(w_n434_0[1]),.dinb(w_n418_0[1]),.dout(n435),.clk(gclk));
	jxor g0372(.dina(w_n435_0[1]),.dinb(w_n416_0[1]),.dout(n436),.clk(gclk));
	jxor g0373(.dina(w_n436_0[1]),.dinb(w_n413_0[1]),.dout(n437),.clk(gclk));
	jxor g0374(.dina(w_n437_0[1]),.dinb(w_n411_0[1]),.dout(n438),.clk(gclk));
	jxor g0375(.dina(w_n438_0[1]),.dinb(w_n408_0[1]),.dout(n439),.clk(gclk));
	jxor g0376(.dina(w_n439_0[1]),.dinb(w_n406_0[1]),.dout(n440),.clk(gclk));
	jxor g0377(.dina(w_n440_0[1]),.dinb(w_n403_0[1]),.dout(n441),.clk(gclk));
	jxor g0378(.dina(w_n441_0[1]),.dinb(w_n401_0[1]),.dout(n442),.clk(gclk));
	jxor g0379(.dina(w_n442_0[1]),.dinb(w_n398_0[1]),.dout(n443),.clk(gclk));
	jxor g0380(.dina(w_n443_0[1]),.dinb(w_n396_0[1]),.dout(n444),.clk(gclk));
	jxor g0381(.dina(w_n444_0[1]),.dinb(w_n393_0[1]),.dout(n445),.clk(gclk));
	jnot g0382(.din(w_n445_0[1]),.dout(n446),.clk(gclk));
	jxor g0383(.dina(w_n446_0[1]),.dinb(w_n391_0[2]),.dout(n447),.clk(gclk));
	jxor g0384(.dina(n447),.dinb(n387),.dout(n448),.clk(gclk));
	jxor g0385(.dina(w_n448_0[1]),.dinb(w_n385_0[1]),.dout(n449),.clk(gclk));
	jxor g0386(.dina(w_n449_0[1]),.dinb(w_dff_B_1wTyjv7c3_1),.dout(w_dff_A_Z99VGWH31_2),.clk(gclk));
	jand g0387(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n451),.clk(gclk));
	jnot g0388(.din(w_n451_0[1]),.dout(n452),.clk(gclk));
	jnot g0389(.din(w_n448_0[0]),.dout(n453),.clk(gclk));
	jor g0390(.dina(n453),.dinb(w_n385_0[0]),.dout(n454),.clk(gclk));
	jor g0391(.dina(w_n449_0[0]),.dinb(w_n380_0[0]),.dout(n455),.clk(gclk));
	jand g0392(.dina(n455),.dinb(w_dff_B_tzl0zDuC0_1),.dout(n456),.clk(gclk));
	jand g0393(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n457),.clk(gclk));
	jnot g0394(.din(w_n457_0[1]),.dout(n458),.clk(gclk));
	jor g0395(.dina(w_n446_0[0]),.dinb(w_n391_0[1]),.dout(n459),.clk(gclk));
	jxor g0396(.dina(w_n445_0[0]),.dinb(w_n391_0[0]),.dout(n460),.clk(gclk));
	jor g0397(.dina(n460),.dinb(w_n386_0[0]),.dout(n461),.clk(gclk));
	jand g0398(.dina(n461),.dinb(n459),.dout(n462),.clk(gclk));
	jand g0399(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n463),.clk(gclk));
	jnot g0400(.din(n463),.dout(n464),.clk(gclk));
	jand g0401(.dina(w_n443_0[0]),.dinb(w_n396_0[0]),.dout(n465),.clk(gclk));
	jand g0402(.dina(w_n444_0[0]),.dinb(w_n393_0[0]),.dout(n466),.clk(gclk));
	jor g0403(.dina(n466),.dinb(n465),.dout(n467),.clk(gclk));
	jand g0404(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n468),.clk(gclk));
	jnot g0405(.din(n468),.dout(n469),.clk(gclk));
	jand g0406(.dina(w_n441_0[0]),.dinb(w_n401_0[0]),.dout(n470),.clk(gclk));
	jand g0407(.dina(w_n442_0[0]),.dinb(w_n398_0[0]),.dout(n471),.clk(gclk));
	jor g0408(.dina(n471),.dinb(n470),.dout(n472),.clk(gclk));
	jand g0409(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n473),.clk(gclk));
	jnot g0410(.din(n473),.dout(n474),.clk(gclk));
	jand g0411(.dina(w_n439_0[0]),.dinb(w_n406_0[0]),.dout(n475),.clk(gclk));
	jand g0412(.dina(w_n440_0[0]),.dinb(w_n403_0[0]),.dout(n476),.clk(gclk));
	jor g0413(.dina(n476),.dinb(n475),.dout(n477),.clk(gclk));
	jand g0414(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n478),.clk(gclk));
	jnot g0415(.din(n478),.dout(n479),.clk(gclk));
	jand g0416(.dina(w_n437_0[0]),.dinb(w_n411_0[0]),.dout(n480),.clk(gclk));
	jand g0417(.dina(w_n438_0[0]),.dinb(w_n408_0[0]),.dout(n481),.clk(gclk));
	jor g0418(.dina(n481),.dinb(n480),.dout(n482),.clk(gclk));
	jand g0419(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n435_0[0]),.dinb(w_n416_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n436_0[0]),.dinb(w_n413_0[0]),.dout(n486),.clk(gclk));
	jor g0423(.dina(n486),.dinb(n485),.dout(n487),.clk(gclk));
	jand g0424(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n433_0[0]),.dinb(w_n423_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n434_0[0]),.dinb(w_n418_0[0]),.dout(n491),.clk(gclk));
	jor g0428(.dina(n491),.dinb(n490),.dout(n492),.clk(gclk));
	jand g0429(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jor g0431(.dina(w_n431_0[0]),.dinb(w_n358_0[0]),.dout(n495),.clk(gclk));
	jand g0432(.dina(w_n432_0[0]),.dinb(w_n425_0[0]),.dout(n496),.clk(gclk));
	jnot g0433(.din(n496),.dout(n497),.clk(gclk));
	jand g0434(.dina(n497),.dinb(n495),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_G307gat_4[1]),.dinb(w_G154gat_6[2]),.dout(n500),.clk(gclk));
	jnot g0437(.din(n500),.dout(n501),.clk(gclk));
	jand g0438(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n502),.clk(gclk));
	jand g0439(.dina(w_n502_0[1]),.dinb(w_n429_0[0]),.dout(n503),.clk(gclk));
	jnot g0440(.din(w_n503_0[2]),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n505),.clk(gclk));
	jor g0442(.dina(w_n505_0[1]),.dinb(w_n426_0[0]),.dout(n506),.clk(gclk));
	jand g0443(.dina(n506),.dinb(n504),.dout(n507),.clk(gclk));
	jxor g0444(.dina(w_n507_0[1]),.dinb(w_n427_0[1]),.dout(n508),.clk(gclk));
	jxor g0445(.dina(w_n508_0[1]),.dinb(w_n501_0[1]),.dout(n509),.clk(gclk));
	jxor g0446(.dina(w_n509_0[1]),.dinb(w_n499_0[1]),.dout(n510),.clk(gclk));
	jxor g0447(.dina(w_n510_0[1]),.dinb(w_n494_0[1]),.dout(n511),.clk(gclk));
	jxor g0448(.dina(w_n511_0[1]),.dinb(w_n492_0[1]),.dout(n512),.clk(gclk));
	jxor g0449(.dina(w_n512_0[1]),.dinb(w_n489_0[1]),.dout(n513),.clk(gclk));
	jxor g0450(.dina(w_n513_0[1]),.dinb(w_n487_0[1]),.dout(n514),.clk(gclk));
	jxor g0451(.dina(w_n514_0[1]),.dinb(w_n484_0[1]),.dout(n515),.clk(gclk));
	jxor g0452(.dina(w_n515_0[1]),.dinb(w_n482_0[1]),.dout(n516),.clk(gclk));
	jxor g0453(.dina(w_n516_0[1]),.dinb(w_n479_0[1]),.dout(n517),.clk(gclk));
	jxor g0454(.dina(w_n517_0[1]),.dinb(w_n477_0[1]),.dout(n518),.clk(gclk));
	jxor g0455(.dina(w_n518_0[1]),.dinb(w_n474_0[1]),.dout(n519),.clk(gclk));
	jxor g0456(.dina(w_n519_0[1]),.dinb(w_n472_0[1]),.dout(n520),.clk(gclk));
	jxor g0457(.dina(w_n520_0[1]),.dinb(w_n469_0[1]),.dout(n521),.clk(gclk));
	jxor g0458(.dina(w_n521_0[1]),.dinb(w_n467_0[1]),.dout(n522),.clk(gclk));
	jxor g0459(.dina(w_n522_0[1]),.dinb(w_n464_0[1]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[1]),.dout(n524),.clk(gclk));
	jxor g0461(.dina(w_n524_0[1]),.dinb(w_n462_0[2]),.dout(n525),.clk(gclk));
	jxor g0462(.dina(n525),.dinb(n458),.dout(n526),.clk(gclk));
	jxor g0463(.dina(w_n526_0[1]),.dinb(w_n456_0[1]),.dout(n527),.clk(gclk));
	jxor g0464(.dina(w_n527_0[1]),.dinb(w_dff_B_fjZoUprZ9_1),.dout(w_dff_A_afeJhXAY4_2),.clk(gclk));
	jand g0465(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n529),.clk(gclk));
	jnot g0466(.din(w_n529_0[1]),.dout(n530),.clk(gclk));
	jnot g0467(.din(w_n526_0[0]),.dout(n531),.clk(gclk));
	jor g0468(.dina(n531),.dinb(w_n456_0[0]),.dout(n532),.clk(gclk));
	jor g0469(.dina(w_n527_0[0]),.dinb(w_n451_0[0]),.dout(n533),.clk(gclk));
	jand g0470(.dina(n533),.dinb(w_dff_B_W13ktaNM2_1),.dout(n534),.clk(gclk));
	jand g0471(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n535),.clk(gclk));
	jnot g0472(.din(w_n535_0[1]),.dout(n536),.clk(gclk));
	jor g0473(.dina(w_n524_0[0]),.dinb(w_n462_0[1]),.dout(n537),.clk(gclk));
	jxor g0474(.dina(w_n523_0[0]),.dinb(w_n462_0[0]),.dout(n538),.clk(gclk));
	jor g0475(.dina(n538),.dinb(w_n457_0[0]),.dout(n539),.clk(gclk));
	jand g0476(.dina(n539),.dinb(n537),.dout(n540),.clk(gclk));
	jand g0477(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n541),.clk(gclk));
	jnot g0478(.din(n541),.dout(n542),.clk(gclk));
	jand g0479(.dina(w_n521_0[0]),.dinb(w_n467_0[0]),.dout(n543),.clk(gclk));
	jand g0480(.dina(w_n522_0[0]),.dinb(w_n464_0[0]),.dout(n544),.clk(gclk));
	jor g0481(.dina(n544),.dinb(n543),.dout(n545),.clk(gclk));
	jand g0482(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n546),.clk(gclk));
	jnot g0483(.din(n546),.dout(n547),.clk(gclk));
	jand g0484(.dina(w_n519_0[0]),.dinb(w_n472_0[0]),.dout(n548),.clk(gclk));
	jand g0485(.dina(w_n520_0[0]),.dinb(w_n469_0[0]),.dout(n549),.clk(gclk));
	jor g0486(.dina(n549),.dinb(n548),.dout(n550),.clk(gclk));
	jand g0487(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n551),.clk(gclk));
	jnot g0488(.din(n551),.dout(n552),.clk(gclk));
	jand g0489(.dina(w_n517_0[0]),.dinb(w_n477_0[0]),.dout(n553),.clk(gclk));
	jand g0490(.dina(w_n518_0[0]),.dinb(w_n474_0[0]),.dout(n554),.clk(gclk));
	jor g0491(.dina(n554),.dinb(n553),.dout(n555),.clk(gclk));
	jand g0492(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n556),.clk(gclk));
	jnot g0493(.din(n556),.dout(n557),.clk(gclk));
	jand g0494(.dina(w_n515_0[0]),.dinb(w_n482_0[0]),.dout(n558),.clk(gclk));
	jand g0495(.dina(w_n516_0[0]),.dinb(w_n479_0[0]),.dout(n559),.clk(gclk));
	jor g0496(.dina(n559),.dinb(n558),.dout(n560),.clk(gclk));
	jand g0497(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n561),.clk(gclk));
	jnot g0498(.din(n561),.dout(n562),.clk(gclk));
	jand g0499(.dina(w_n513_0[0]),.dinb(w_n487_0[0]),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n514_0[0]),.dinb(w_n484_0[0]),.dout(n564),.clk(gclk));
	jor g0501(.dina(n564),.dinb(n563),.dout(n565),.clk(gclk));
	jand g0502(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n566),.clk(gclk));
	jnot g0503(.din(n566),.dout(n567),.clk(gclk));
	jand g0504(.dina(w_n511_0[0]),.dinb(w_n492_0[0]),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n512_0[0]),.dinb(w_n489_0[0]),.dout(n569),.clk(gclk));
	jor g0506(.dina(n569),.dinb(n568),.dout(n570),.clk(gclk));
	jand g0507(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n571),.clk(gclk));
	jnot g0508(.din(n571),.dout(n572),.clk(gclk));
	jand g0509(.dina(w_n509_0[0]),.dinb(w_n499_0[0]),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n510_0[0]),.dinb(w_n494_0[0]),.dout(n574),.clk(gclk));
	jor g0511(.dina(n574),.dinb(n573),.dout(n575),.clk(gclk));
	jand g0512(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n576),.clk(gclk));
	jnot g0513(.din(n576),.dout(n577),.clk(gclk));
	jor g0514(.dina(w_n507_0[0]),.dinb(w_n427_0[0]),.dout(n578),.clk(gclk));
	jand g0515(.dina(w_n508_0[0]),.dinb(w_n501_0[0]),.dout(n579),.clk(gclk));
	jnot g0516(.din(n579),.dout(n580),.clk(gclk));
	jand g0517(.dina(n580),.dinb(n578),.dout(n581),.clk(gclk));
	jnot g0518(.din(n581),.dout(n582),.clk(gclk));
	jand g0519(.dina(w_G307gat_4[0]),.dinb(w_G171gat_6[2]),.dout(n583),.clk(gclk));
	jnot g0520(.din(n583),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n585),.clk(gclk));
	jand g0522(.dina(w_n585_0[1]),.dinb(w_n505_0[0]),.dout(n586),.clk(gclk));
	jnot g0523(.din(w_n586_0[2]),.dout(n587),.clk(gclk));
	jand g0524(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n588),.clk(gclk));
	jor g0525(.dina(w_n588_0[1]),.dinb(w_n502_0[0]),.dout(n589),.clk(gclk));
	jand g0526(.dina(n589),.dinb(n587),.dout(n590),.clk(gclk));
	jxor g0527(.dina(w_n590_0[1]),.dinb(w_n503_0[1]),.dout(n591),.clk(gclk));
	jxor g0528(.dina(w_n591_0[1]),.dinb(w_n584_0[1]),.dout(n592),.clk(gclk));
	jxor g0529(.dina(w_n592_0[1]),.dinb(w_n582_0[1]),.dout(n593),.clk(gclk));
	jxor g0530(.dina(w_n593_0[1]),.dinb(w_n577_0[1]),.dout(n594),.clk(gclk));
	jxor g0531(.dina(w_n594_0[1]),.dinb(w_n575_0[1]),.dout(n595),.clk(gclk));
	jxor g0532(.dina(w_n595_0[1]),.dinb(w_n572_0[1]),.dout(n596),.clk(gclk));
	jxor g0533(.dina(w_n596_0[1]),.dinb(w_n570_0[1]),.dout(n597),.clk(gclk));
	jxor g0534(.dina(w_n597_0[1]),.dinb(w_n567_0[1]),.dout(n598),.clk(gclk));
	jxor g0535(.dina(w_n598_0[1]),.dinb(w_n565_0[1]),.dout(n599),.clk(gclk));
	jxor g0536(.dina(w_n599_0[1]),.dinb(w_n562_0[1]),.dout(n600),.clk(gclk));
	jxor g0537(.dina(w_n600_0[1]),.dinb(w_n560_0[1]),.dout(n601),.clk(gclk));
	jxor g0538(.dina(w_n601_0[1]),.dinb(w_n557_0[1]),.dout(n602),.clk(gclk));
	jxor g0539(.dina(w_n602_0[1]),.dinb(w_n555_0[1]),.dout(n603),.clk(gclk));
	jxor g0540(.dina(w_n603_0[1]),.dinb(w_n552_0[1]),.dout(n604),.clk(gclk));
	jxor g0541(.dina(w_n604_0[1]),.dinb(w_n550_0[1]),.dout(n605),.clk(gclk));
	jxor g0542(.dina(w_n605_0[1]),.dinb(w_n547_0[1]),.dout(n606),.clk(gclk));
	jxor g0543(.dina(w_n606_0[1]),.dinb(w_n545_0[1]),.dout(n607),.clk(gclk));
	jxor g0544(.dina(w_n607_0[1]),.dinb(w_n542_0[1]),.dout(n608),.clk(gclk));
	jnot g0545(.din(w_n608_0[1]),.dout(n609),.clk(gclk));
	jxor g0546(.dina(w_n609_0[1]),.dinb(w_n540_0[2]),.dout(n610),.clk(gclk));
	jxor g0547(.dina(n610),.dinb(n536),.dout(n611),.clk(gclk));
	jxor g0548(.dina(w_n611_0[1]),.dinb(w_n534_0[1]),.dout(n612),.clk(gclk));
	jxor g0549(.dina(w_n612_0[1]),.dinb(w_dff_B_r1iAy6MU3_1),.dout(w_dff_A_FoMYUxYC3_2),.clk(gclk));
	jand g0550(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n614),.clk(gclk));
	jnot g0551(.din(w_n614_0[1]),.dout(n615),.clk(gclk));
	jnot g0552(.din(w_n611_0[0]),.dout(n616),.clk(gclk));
	jor g0553(.dina(n616),.dinb(w_n534_0[0]),.dout(n617),.clk(gclk));
	jor g0554(.dina(w_n612_0[0]),.dinb(w_n529_0[0]),.dout(n618),.clk(gclk));
	jand g0555(.dina(n618),.dinb(w_dff_B_sHrr4wRB8_1),.dout(n619),.clk(gclk));
	jand g0556(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n620),.clk(gclk));
	jnot g0557(.din(w_n620_0[1]),.dout(n621),.clk(gclk));
	jor g0558(.dina(w_n609_0[0]),.dinb(w_n540_0[1]),.dout(n622),.clk(gclk));
	jxor g0559(.dina(w_n608_0[0]),.dinb(w_n540_0[0]),.dout(n623),.clk(gclk));
	jor g0560(.dina(n623),.dinb(w_n535_0[0]),.dout(n624),.clk(gclk));
	jand g0561(.dina(n624),.dinb(n622),.dout(n625),.clk(gclk));
	jand g0562(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n626),.clk(gclk));
	jnot g0563(.din(n626),.dout(n627),.clk(gclk));
	jand g0564(.dina(w_n606_0[0]),.dinb(w_n545_0[0]),.dout(n628),.clk(gclk));
	jand g0565(.dina(w_n607_0[0]),.dinb(w_n542_0[0]),.dout(n629),.clk(gclk));
	jor g0566(.dina(n629),.dinb(n628),.dout(n630),.clk(gclk));
	jand g0567(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n631),.clk(gclk));
	jnot g0568(.din(n631),.dout(n632),.clk(gclk));
	jand g0569(.dina(w_n604_0[0]),.dinb(w_n550_0[0]),.dout(n633),.clk(gclk));
	jand g0570(.dina(w_n605_0[0]),.dinb(w_n547_0[0]),.dout(n634),.clk(gclk));
	jor g0571(.dina(n634),.dinb(n633),.dout(n635),.clk(gclk));
	jand g0572(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n636),.clk(gclk));
	jnot g0573(.din(n636),.dout(n637),.clk(gclk));
	jand g0574(.dina(w_n602_0[0]),.dinb(w_n555_0[0]),.dout(n638),.clk(gclk));
	jand g0575(.dina(w_n603_0[0]),.dinb(w_n552_0[0]),.dout(n639),.clk(gclk));
	jor g0576(.dina(n639),.dinb(n638),.dout(n640),.clk(gclk));
	jand g0577(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n641),.clk(gclk));
	jnot g0578(.din(n641),.dout(n642),.clk(gclk));
	jand g0579(.dina(w_n600_0[0]),.dinb(w_n560_0[0]),.dout(n643),.clk(gclk));
	jand g0580(.dina(w_n601_0[0]),.dinb(w_n557_0[0]),.dout(n644),.clk(gclk));
	jor g0581(.dina(n644),.dinb(n643),.dout(n645),.clk(gclk));
	jand g0582(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n646),.clk(gclk));
	jnot g0583(.din(n646),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_n598_0[0]),.dinb(w_n565_0[0]),.dout(n648),.clk(gclk));
	jand g0585(.dina(w_n599_0[0]),.dinb(w_n562_0[0]),.dout(n649),.clk(gclk));
	jor g0586(.dina(n649),.dinb(n648),.dout(n650),.clk(gclk));
	jand g0587(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n651),.clk(gclk));
	jnot g0588(.din(n651),.dout(n652),.clk(gclk));
	jand g0589(.dina(w_n596_0[0]),.dinb(w_n570_0[0]),.dout(n653),.clk(gclk));
	jand g0590(.dina(w_n597_0[0]),.dinb(w_n567_0[0]),.dout(n654),.clk(gclk));
	jor g0591(.dina(n654),.dinb(n653),.dout(n655),.clk(gclk));
	jand g0592(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n656),.clk(gclk));
	jnot g0593(.din(n656),.dout(n657),.clk(gclk));
	jand g0594(.dina(w_n594_0[0]),.dinb(w_n575_0[0]),.dout(n658),.clk(gclk));
	jand g0595(.dina(w_n595_0[0]),.dinb(w_n572_0[0]),.dout(n659),.clk(gclk));
	jor g0596(.dina(n659),.dinb(n658),.dout(n660),.clk(gclk));
	jand g0597(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n661),.clk(gclk));
	jnot g0598(.din(n661),.dout(n662),.clk(gclk));
	jand g0599(.dina(w_n592_0[0]),.dinb(w_n582_0[0]),.dout(n663),.clk(gclk));
	jand g0600(.dina(w_n593_0[0]),.dinb(w_n577_0[0]),.dout(n664),.clk(gclk));
	jor g0601(.dina(n664),.dinb(n663),.dout(n665),.clk(gclk));
	jand g0602(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n666),.clk(gclk));
	jnot g0603(.din(n666),.dout(n667),.clk(gclk));
	jor g0604(.dina(w_n590_0[0]),.dinb(w_n503_0[0]),.dout(n668),.clk(gclk));
	jand g0605(.dina(w_n591_0[0]),.dinb(w_n584_0[0]),.dout(n669),.clk(gclk));
	jnot g0606(.din(n669),.dout(n670),.clk(gclk));
	jand g0607(.dina(n670),.dinb(n668),.dout(n671),.clk(gclk));
	jnot g0608(.din(n671),.dout(n672),.clk(gclk));
	jand g0609(.dina(w_G307gat_3[2]),.dinb(w_G188gat_6[2]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n675_0[1]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jnot g0613(.din(w_n676_0[2]),.dout(n677),.clk(gclk));
	jand g0614(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n678),.clk(gclk));
	jor g0615(.dina(w_n678_0[1]),.dinb(w_n585_0[0]),.dout(n679),.clk(gclk));
	jand g0616(.dina(n679),.dinb(n677),.dout(n680),.clk(gclk));
	jxor g0617(.dina(w_n680_0[1]),.dinb(w_n586_0[1]),.dout(n681),.clk(gclk));
	jxor g0618(.dina(w_n681_0[1]),.dinb(w_n674_0[1]),.dout(n682),.clk(gclk));
	jxor g0619(.dina(w_n682_0[1]),.dinb(w_n672_0[1]),.dout(n683),.clk(gclk));
	jxor g0620(.dina(w_n683_0[1]),.dinb(w_n667_0[1]),.dout(n684),.clk(gclk));
	jxor g0621(.dina(w_n684_0[1]),.dinb(w_n665_0[1]),.dout(n685),.clk(gclk));
	jxor g0622(.dina(w_n685_0[1]),.dinb(w_n662_0[1]),.dout(n686),.clk(gclk));
	jxor g0623(.dina(w_n686_0[1]),.dinb(w_n660_0[1]),.dout(n687),.clk(gclk));
	jxor g0624(.dina(w_n687_0[1]),.dinb(w_n657_0[1]),.dout(n688),.clk(gclk));
	jxor g0625(.dina(w_n688_0[1]),.dinb(w_n655_0[1]),.dout(n689),.clk(gclk));
	jxor g0626(.dina(w_n689_0[1]),.dinb(w_n652_0[1]),.dout(n690),.clk(gclk));
	jxor g0627(.dina(w_n690_0[1]),.dinb(w_n650_0[1]),.dout(n691),.clk(gclk));
	jxor g0628(.dina(w_n691_0[1]),.dinb(w_n647_0[1]),.dout(n692),.clk(gclk));
	jxor g0629(.dina(w_n692_0[1]),.dinb(w_n645_0[1]),.dout(n693),.clk(gclk));
	jxor g0630(.dina(w_n693_0[1]),.dinb(w_n642_0[1]),.dout(n694),.clk(gclk));
	jxor g0631(.dina(w_n694_0[1]),.dinb(w_n640_0[1]),.dout(n695),.clk(gclk));
	jxor g0632(.dina(w_n695_0[1]),.dinb(w_n637_0[1]),.dout(n696),.clk(gclk));
	jxor g0633(.dina(w_n696_0[1]),.dinb(w_n635_0[1]),.dout(n697),.clk(gclk));
	jxor g0634(.dina(w_n697_0[1]),.dinb(w_n632_0[1]),.dout(n698),.clk(gclk));
	jxor g0635(.dina(w_n698_0[1]),.dinb(w_n630_0[1]),.dout(n699),.clk(gclk));
	jxor g0636(.dina(w_n699_0[1]),.dinb(w_n627_0[1]),.dout(n700),.clk(gclk));
	jnot g0637(.din(w_n700_0[1]),.dout(n701),.clk(gclk));
	jxor g0638(.dina(w_n701_0[1]),.dinb(w_n625_0[2]),.dout(n702),.clk(gclk));
	jxor g0639(.dina(n702),.dinb(n621),.dout(n703),.clk(gclk));
	jxor g0640(.dina(w_n703_0[1]),.dinb(w_n619_0[1]),.dout(n704),.clk(gclk));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_dff_B_Vb5ZFRw32_1),.dout(w_dff_A_GmHJ0a9t0_2),.clk(gclk));
	jand g0642(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n706),.clk(gclk));
	jnot g0643(.din(w_n706_0[1]),.dout(n707),.clk(gclk));
	jnot g0644(.din(w_n703_0[0]),.dout(n708),.clk(gclk));
	jor g0645(.dina(n708),.dinb(w_n619_0[0]),.dout(n709),.clk(gclk));
	jor g0646(.dina(w_n704_0[0]),.dinb(w_n614_0[0]),.dout(n710),.clk(gclk));
	jand g0647(.dina(n710),.dinb(w_dff_B_LszaTL6P4_1),.dout(n711),.clk(gclk));
	jand g0648(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n712),.clk(gclk));
	jnot g0649(.din(w_n712_0[1]),.dout(n713),.clk(gclk));
	jor g0650(.dina(w_n701_0[0]),.dinb(w_n625_0[1]),.dout(n714),.clk(gclk));
	jxor g0651(.dina(w_n700_0[0]),.dinb(w_n625_0[0]),.dout(n715),.clk(gclk));
	jor g0652(.dina(n715),.dinb(w_n620_0[0]),.dout(n716),.clk(gclk));
	jand g0653(.dina(n716),.dinb(n714),.dout(n717),.clk(gclk));
	jand g0654(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n718),.clk(gclk));
	jnot g0655(.din(n718),.dout(n719),.clk(gclk));
	jand g0656(.dina(w_n698_0[0]),.dinb(w_n630_0[0]),.dout(n720),.clk(gclk));
	jand g0657(.dina(w_n699_0[0]),.dinb(w_n627_0[0]),.dout(n721),.clk(gclk));
	jor g0658(.dina(n721),.dinb(n720),.dout(n722),.clk(gclk));
	jand g0659(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n723),.clk(gclk));
	jnot g0660(.din(n723),.dout(n724),.clk(gclk));
	jand g0661(.dina(w_n696_0[0]),.dinb(w_n635_0[0]),.dout(n725),.clk(gclk));
	jand g0662(.dina(w_n697_0[0]),.dinb(w_n632_0[0]),.dout(n726),.clk(gclk));
	jor g0663(.dina(n726),.dinb(n725),.dout(n727),.clk(gclk));
	jand g0664(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n728),.clk(gclk));
	jnot g0665(.din(n728),.dout(n729),.clk(gclk));
	jand g0666(.dina(w_n694_0[0]),.dinb(w_n640_0[0]),.dout(n730),.clk(gclk));
	jand g0667(.dina(w_n695_0[0]),.dinb(w_n637_0[0]),.dout(n731),.clk(gclk));
	jor g0668(.dina(n731),.dinb(n730),.dout(n732),.clk(gclk));
	jand g0669(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n733),.clk(gclk));
	jnot g0670(.din(n733),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_n692_0[0]),.dinb(w_n645_0[0]),.dout(n735),.clk(gclk));
	jand g0672(.dina(w_n693_0[0]),.dinb(w_n642_0[0]),.dout(n736),.clk(gclk));
	jor g0673(.dina(n736),.dinb(n735),.dout(n737),.clk(gclk));
	jand g0674(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n738),.clk(gclk));
	jnot g0675(.din(n738),.dout(n739),.clk(gclk));
	jand g0676(.dina(w_n690_0[0]),.dinb(w_n650_0[0]),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_n691_0[0]),.dinb(w_n647_0[0]),.dout(n741),.clk(gclk));
	jor g0678(.dina(n741),.dinb(n740),.dout(n742),.clk(gclk));
	jand g0679(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n743),.clk(gclk));
	jnot g0680(.din(n743),.dout(n744),.clk(gclk));
	jand g0681(.dina(w_n688_0[0]),.dinb(w_n655_0[0]),.dout(n745),.clk(gclk));
	jand g0682(.dina(w_n689_0[0]),.dinb(w_n652_0[0]),.dout(n746),.clk(gclk));
	jor g0683(.dina(n746),.dinb(n745),.dout(n747),.clk(gclk));
	jand g0684(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n748),.clk(gclk));
	jnot g0685(.din(n748),.dout(n749),.clk(gclk));
	jand g0686(.dina(w_n686_0[0]),.dinb(w_n660_0[0]),.dout(n750),.clk(gclk));
	jand g0687(.dina(w_n687_0[0]),.dinb(w_n657_0[0]),.dout(n751),.clk(gclk));
	jor g0688(.dina(n751),.dinb(n750),.dout(n752),.clk(gclk));
	jand g0689(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n753),.clk(gclk));
	jnot g0690(.din(n753),.dout(n754),.clk(gclk));
	jand g0691(.dina(w_n684_0[0]),.dinb(w_n665_0[0]),.dout(n755),.clk(gclk));
	jand g0692(.dina(w_n685_0[0]),.dinb(w_n662_0[0]),.dout(n756),.clk(gclk));
	jor g0693(.dina(n756),.dinb(n755),.dout(n757),.clk(gclk));
	jand g0694(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n758),.clk(gclk));
	jnot g0695(.din(n758),.dout(n759),.clk(gclk));
	jand g0696(.dina(w_n682_0[0]),.dinb(w_n672_0[0]),.dout(n760),.clk(gclk));
	jand g0697(.dina(w_n683_0[0]),.dinb(w_n667_0[0]),.dout(n761),.clk(gclk));
	jor g0698(.dina(n761),.dinb(n760),.dout(n762),.clk(gclk));
	jand g0699(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n763),.clk(gclk));
	jnot g0700(.din(n763),.dout(n764),.clk(gclk));
	jor g0701(.dina(w_n680_0[0]),.dinb(w_n586_0[0]),.dout(n765),.clk(gclk));
	jand g0702(.dina(w_n681_0[0]),.dinb(w_n674_0[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(n767),.dinb(n765),.dout(n768),.clk(gclk));
	jnot g0705(.din(n768),.dout(n769),.clk(gclk));
	jand g0706(.dina(w_G307gat_3[1]),.dinb(w_G205gat_6[2]),.dout(n770),.clk(gclk));
	jnot g0707(.din(n770),.dout(n771),.clk(gclk));
	jand g0708(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n772_0[1]),.dinb(w_n678_0[0]),.dout(n773),.clk(gclk));
	jnot g0710(.din(w_n773_0[1]),.dout(n774),.clk(gclk));
	jand g0711(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n775),.clk(gclk));
	jor g0712(.dina(w_n775_0[1]),.dinb(w_n675_0[0]),.dout(n776),.clk(gclk));
	jand g0713(.dina(n776),.dinb(w_n774_0[1]),.dout(n777),.clk(gclk));
	jxor g0714(.dina(w_n777_0[1]),.dinb(w_n676_0[1]),.dout(n778),.clk(gclk));
	jxor g0715(.dina(w_n778_0[1]),.dinb(w_n771_0[1]),.dout(n779),.clk(gclk));
	jxor g0716(.dina(w_n779_0[1]),.dinb(w_n769_0[1]),.dout(n780),.clk(gclk));
	jxor g0717(.dina(w_n780_0[1]),.dinb(w_n764_0[1]),.dout(n781),.clk(gclk));
	jxor g0718(.dina(w_n781_0[1]),.dinb(w_n762_0[1]),.dout(n782),.clk(gclk));
	jxor g0719(.dina(w_n782_0[1]),.dinb(w_n759_0[1]),.dout(n783),.clk(gclk));
	jxor g0720(.dina(w_n783_0[1]),.dinb(w_n757_0[1]),.dout(n784),.clk(gclk));
	jxor g0721(.dina(w_n784_0[1]),.dinb(w_n754_0[1]),.dout(n785),.clk(gclk));
	jxor g0722(.dina(w_n785_0[1]),.dinb(w_n752_0[1]),.dout(n786),.clk(gclk));
	jxor g0723(.dina(w_n786_0[1]),.dinb(w_n749_0[1]),.dout(n787),.clk(gclk));
	jxor g0724(.dina(w_n787_0[1]),.dinb(w_n747_0[1]),.dout(n788),.clk(gclk));
	jxor g0725(.dina(w_n788_0[1]),.dinb(w_n744_0[1]),.dout(n789),.clk(gclk));
	jxor g0726(.dina(w_n789_0[1]),.dinb(w_n742_0[1]),.dout(n790),.clk(gclk));
	jxor g0727(.dina(w_n790_0[1]),.dinb(w_n739_0[1]),.dout(n791),.clk(gclk));
	jxor g0728(.dina(w_n791_0[1]),.dinb(w_n737_0[1]),.dout(n792),.clk(gclk));
	jxor g0729(.dina(w_n792_0[1]),.dinb(w_n734_0[1]),.dout(n793),.clk(gclk));
	jxor g0730(.dina(w_n793_0[1]),.dinb(w_n732_0[1]),.dout(n794),.clk(gclk));
	jxor g0731(.dina(w_n794_0[1]),.dinb(w_n729_0[1]),.dout(n795),.clk(gclk));
	jxor g0732(.dina(w_n795_0[1]),.dinb(w_n727_0[1]),.dout(n796),.clk(gclk));
	jxor g0733(.dina(w_n796_0[1]),.dinb(w_n724_0[1]),.dout(n797),.clk(gclk));
	jxor g0734(.dina(w_n797_0[1]),.dinb(w_n722_0[1]),.dout(n798),.clk(gclk));
	jxor g0735(.dina(w_n798_0[1]),.dinb(w_n719_0[1]),.dout(n799),.clk(gclk));
	jnot g0736(.din(w_n799_0[1]),.dout(n800),.clk(gclk));
	jxor g0737(.dina(w_n800_0[1]),.dinb(w_n717_0[2]),.dout(n801),.clk(gclk));
	jxor g0738(.dina(n801),.dinb(n713),.dout(n802),.clk(gclk));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n711_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_dff_B_khjF5Lua6_1),.dout(w_dff_A_XaMEPoS81_2),.clk(gclk));
	jand g0741(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n805),.clk(gclk));
	jnot g0742(.din(w_n805_0[1]),.dout(n806),.clk(gclk));
	jnot g0743(.din(w_n802_0[0]),.dout(n807),.clk(gclk));
	jor g0744(.dina(n807),.dinb(w_n711_0[0]),.dout(n808),.clk(gclk));
	jor g0745(.dina(w_n803_0[0]),.dinb(w_n706_0[0]),.dout(n809),.clk(gclk));
	jand g0746(.dina(n809),.dinb(w_dff_B_pDRcoDZO2_1),.dout(n810),.clk(gclk));
	jand g0747(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n811),.clk(gclk));
	jor g0748(.dina(w_n800_0[0]),.dinb(w_n717_0[1]),.dout(n812),.clk(gclk));
	jxor g0749(.dina(w_n799_0[0]),.dinb(w_n717_0[0]),.dout(n813),.clk(gclk));
	jor g0750(.dina(n813),.dinb(w_n712_0[0]),.dout(n814),.clk(gclk));
	jand g0751(.dina(n814),.dinb(n812),.dout(n815),.clk(gclk));
	jand g0752(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n816),.clk(gclk));
	jnot g0753(.din(w_n816_0[1]),.dout(n817),.clk(gclk));
	jand g0754(.dina(w_n797_0[0]),.dinb(w_n722_0[0]),.dout(n818),.clk(gclk));
	jand g0755(.dina(w_n798_0[0]),.dinb(w_n719_0[0]),.dout(n819),.clk(gclk));
	jor g0756(.dina(n819),.dinb(n818),.dout(n820),.clk(gclk));
	jand g0757(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n821),.clk(gclk));
	jnot g0758(.din(n821),.dout(n822),.clk(gclk));
	jand g0759(.dina(w_n795_0[0]),.dinb(w_n727_0[0]),.dout(n823),.clk(gclk));
	jand g0760(.dina(w_n796_0[0]),.dinb(w_n724_0[0]),.dout(n824),.clk(gclk));
	jor g0761(.dina(n824),.dinb(n823),.dout(n825),.clk(gclk));
	jand g0762(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n826),.clk(gclk));
	jnot g0763(.din(n826),.dout(n827),.clk(gclk));
	jand g0764(.dina(w_n793_0[0]),.dinb(w_n732_0[0]),.dout(n828),.clk(gclk));
	jand g0765(.dina(w_n794_0[0]),.dinb(w_n729_0[0]),.dout(n829),.clk(gclk));
	jor g0766(.dina(n829),.dinb(n828),.dout(n830),.clk(gclk));
	jand g0767(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n831),.clk(gclk));
	jnot g0768(.din(n831),.dout(n832),.clk(gclk));
	jand g0769(.dina(w_n791_0[0]),.dinb(w_n737_0[0]),.dout(n833),.clk(gclk));
	jand g0770(.dina(w_n792_0[0]),.dinb(w_n734_0[0]),.dout(n834),.clk(gclk));
	jor g0771(.dina(n834),.dinb(n833),.dout(n835),.clk(gclk));
	jand g0772(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n836),.clk(gclk));
	jnot g0773(.din(n836),.dout(n837),.clk(gclk));
	jand g0774(.dina(w_n789_0[0]),.dinb(w_n742_0[0]),.dout(n838),.clk(gclk));
	jand g0775(.dina(w_n790_0[0]),.dinb(w_n739_0[0]),.dout(n839),.clk(gclk));
	jor g0776(.dina(n839),.dinb(n838),.dout(n840),.clk(gclk));
	jand g0777(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n841),.clk(gclk));
	jnot g0778(.din(n841),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n787_0[0]),.dinb(w_n747_0[0]),.dout(n843),.clk(gclk));
	jand g0780(.dina(w_n788_0[0]),.dinb(w_n744_0[0]),.dout(n844),.clk(gclk));
	jor g0781(.dina(n844),.dinb(n843),.dout(n845),.clk(gclk));
	jand g0782(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n846),.clk(gclk));
	jnot g0783(.din(n846),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n785_0[0]),.dinb(w_n752_0[0]),.dout(n848),.clk(gclk));
	jand g0785(.dina(w_n786_0[0]),.dinb(w_n749_0[0]),.dout(n849),.clk(gclk));
	jor g0786(.dina(n849),.dinb(n848),.dout(n850),.clk(gclk));
	jand g0787(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n851),.clk(gclk));
	jnot g0788(.din(n851),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n783_0[0]),.dinb(w_n757_0[0]),.dout(n853),.clk(gclk));
	jand g0790(.dina(w_n784_0[0]),.dinb(w_n754_0[0]),.dout(n854),.clk(gclk));
	jor g0791(.dina(n854),.dinb(n853),.dout(n855),.clk(gclk));
	jand g0792(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n856),.clk(gclk));
	jnot g0793(.din(n856),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n781_0[0]),.dinb(w_n762_0[0]),.dout(n858),.clk(gclk));
	jand g0795(.dina(w_n782_0[0]),.dinb(w_n759_0[0]),.dout(n859),.clk(gclk));
	jor g0796(.dina(n859),.dinb(n858),.dout(n860),.clk(gclk));
	jand g0797(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n861),.clk(gclk));
	jnot g0798(.din(n861),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n779_0[0]),.dinb(w_n769_0[0]),.dout(n863),.clk(gclk));
	jand g0800(.dina(w_n780_0[0]),.dinb(w_n764_0[0]),.dout(n864),.clk(gclk));
	jor g0801(.dina(n864),.dinb(n863),.dout(n865),.clk(gclk));
	jand g0802(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n866),.clk(gclk));
	jnot g0803(.din(n866),.dout(n867),.clk(gclk));
	jor g0804(.dina(w_n777_0[0]),.dinb(w_n676_0[0]),.dout(n868),.clk(gclk));
	jand g0805(.dina(w_n778_0[0]),.dinb(w_n771_0[0]),.dout(n869),.clk(gclk));
	jnot g0806(.din(n869),.dout(n870),.clk(gclk));
	jand g0807(.dina(n870),.dinb(n868),.dout(n871),.clk(gclk));
	jnot g0808(.din(n871),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_G307gat_3[0]),.dinb(w_G222gat_6[2]),.dout(n873),.clk(gclk));
	jnot g0810(.din(n873),.dout(n874),.clk(gclk));
	jand g0811(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n875),.clk(gclk));
	jxor g0812(.dina(w_n875_0[1]),.dinb(w_n772_0[0]),.dout(n876),.clk(gclk));
	jor g0813(.dina(n876),.dinb(w_n773_0[0]),.dout(n877),.clk(gclk));
	jor g0814(.dina(w_n875_0[0]),.dinb(w_n774_0[0]),.dout(n878),.clk(gclk));
	jand g0815(.dina(n878),.dinb(w_n877_0[1]),.dout(n879),.clk(gclk));
	jxor g0816(.dina(w_n879_0[1]),.dinb(w_n874_0[1]),.dout(n880),.clk(gclk));
	jxor g0817(.dina(w_n880_0[1]),.dinb(w_n872_0[1]),.dout(n881),.clk(gclk));
	jxor g0818(.dina(w_n881_0[1]),.dinb(w_n867_0[1]),.dout(n882),.clk(gclk));
	jxor g0819(.dina(w_n882_0[1]),.dinb(w_n865_0[1]),.dout(n883),.clk(gclk));
	jxor g0820(.dina(w_n883_0[1]),.dinb(w_n862_0[1]),.dout(n884),.clk(gclk));
	jxor g0821(.dina(w_n884_0[1]),.dinb(w_n860_0[1]),.dout(n885),.clk(gclk));
	jxor g0822(.dina(w_n885_0[1]),.dinb(w_n857_0[1]),.dout(n886),.clk(gclk));
	jxor g0823(.dina(w_n886_0[1]),.dinb(w_n855_0[1]),.dout(n887),.clk(gclk));
	jxor g0824(.dina(w_n887_0[1]),.dinb(w_n852_0[1]),.dout(n888),.clk(gclk));
	jxor g0825(.dina(w_n888_0[1]),.dinb(w_n850_0[1]),.dout(n889),.clk(gclk));
	jxor g0826(.dina(w_n889_0[1]),.dinb(w_n847_0[1]),.dout(n890),.clk(gclk));
	jxor g0827(.dina(w_n890_0[1]),.dinb(w_n845_0[1]),.dout(n891),.clk(gclk));
	jxor g0828(.dina(w_n891_0[1]),.dinb(w_n842_0[1]),.dout(n892),.clk(gclk));
	jxor g0829(.dina(w_n892_0[1]),.dinb(w_n840_0[1]),.dout(n893),.clk(gclk));
	jxor g0830(.dina(w_n893_0[1]),.dinb(w_n837_0[1]),.dout(n894),.clk(gclk));
	jxor g0831(.dina(w_n894_0[1]),.dinb(w_n835_0[1]),.dout(n895),.clk(gclk));
	jxor g0832(.dina(w_n895_0[1]),.dinb(w_n832_0[1]),.dout(n896),.clk(gclk));
	jxor g0833(.dina(w_n896_0[1]),.dinb(w_n830_0[1]),.dout(n897),.clk(gclk));
	jxor g0834(.dina(w_n897_0[1]),.dinb(w_n827_0[1]),.dout(n898),.clk(gclk));
	jxor g0835(.dina(w_n898_0[1]),.dinb(w_n825_0[1]),.dout(n899),.clk(gclk));
	jxor g0836(.dina(w_n899_0[1]),.dinb(w_n822_0[1]),.dout(n900),.clk(gclk));
	jxor g0837(.dina(w_n900_0[2]),.dinb(w_n820_0[2]),.dout(n901),.clk(gclk));
	jxor g0838(.dina(n901),.dinb(n817),.dout(n902),.clk(gclk));
	jxor g0839(.dina(w_n902_0[1]),.dinb(w_n815_0[1]),.dout(n903),.clk(gclk));
	jxor g0840(.dina(w_n903_0[1]),.dinb(w_n811_0[1]),.dout(n904),.clk(gclk));
	jxor g0841(.dina(w_n904_0[1]),.dinb(w_n810_0[1]),.dout(n905),.clk(gclk));
	jxor g0842(.dina(w_n905_0[1]),.dinb(w_dff_B_jf1zmcsS5_1),.dout(w_dff_A_r1aCngrq2_2),.clk(gclk));
	jnot g0843(.din(w_n904_0[0]),.dout(n907),.clk(gclk));
	jor g0844(.dina(n907),.dinb(w_n810_0[0]),.dout(n908),.clk(gclk));
	jor g0845(.dina(w_n905_0[0]),.dinb(w_n805_0[0]),.dout(n909),.clk(gclk));
	jand g0846(.dina(n909),.dinb(w_dff_B_tUJC509k0_1),.dout(n910),.clk(gclk));
	jand g0847(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n911),.clk(gclk));
	jnot g0848(.din(w_n902_0[0]),.dout(n912),.clk(gclk));
	jor g0849(.dina(n912),.dinb(w_n815_0[0]),.dout(n913),.clk(gclk));
	jor g0850(.dina(w_n903_0[0]),.dinb(w_n811_0[0]),.dout(n914),.clk(gclk));
	jand g0851(.dina(n914),.dinb(n913),.dout(n915),.clk(gclk));
	jand g0852(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n916),.clk(gclk));
	jand g0853(.dina(w_n900_0[1]),.dinb(w_n820_0[1]),.dout(n917),.clk(gclk));
	jnot g0854(.din(n917),.dout(n918),.clk(gclk));
	jnot g0855(.din(w_n900_0[0]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(n919),.dinb(w_n820_0[0]),.dout(n920),.clk(gclk));
	jor g0857(.dina(n920),.dinb(w_n816_0[0]),.dout(n921),.clk(gclk));
	jand g0858(.dina(n921),.dinb(n918),.dout(n922),.clk(gclk));
	jand g0859(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n923),.clk(gclk));
	jnot g0860(.din(n923),.dout(n924),.clk(gclk));
	jand g0861(.dina(w_n898_0[0]),.dinb(w_n825_0[0]),.dout(n925),.clk(gclk));
	jand g0862(.dina(w_n899_0[0]),.dinb(w_n822_0[0]),.dout(n926),.clk(gclk));
	jor g0863(.dina(n926),.dinb(n925),.dout(n927),.clk(gclk));
	jand g0864(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n928),.clk(gclk));
	jnot g0865(.din(n928),.dout(n929),.clk(gclk));
	jand g0866(.dina(w_n896_0[0]),.dinb(w_n830_0[0]),.dout(n930),.clk(gclk));
	jand g0867(.dina(w_n897_0[0]),.dinb(w_n827_0[0]),.dout(n931),.clk(gclk));
	jor g0868(.dina(n931),.dinb(n930),.dout(n932),.clk(gclk));
	jand g0869(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n933),.clk(gclk));
	jnot g0870(.din(n933),.dout(n934),.clk(gclk));
	jand g0871(.dina(w_n894_0[0]),.dinb(w_n835_0[0]),.dout(n935),.clk(gclk));
	jand g0872(.dina(w_n895_0[0]),.dinb(w_n832_0[0]),.dout(n936),.clk(gclk));
	jor g0873(.dina(n936),.dinb(n935),.dout(n937),.clk(gclk));
	jand g0874(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n938),.clk(gclk));
	jnot g0875(.din(n938),.dout(n939),.clk(gclk));
	jand g0876(.dina(w_n892_0[0]),.dinb(w_n840_0[0]),.dout(n940),.clk(gclk));
	jand g0877(.dina(w_n893_0[0]),.dinb(w_n837_0[0]),.dout(n941),.clk(gclk));
	jor g0878(.dina(n941),.dinb(n940),.dout(n942),.clk(gclk));
	jand g0879(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n943),.clk(gclk));
	jnot g0880(.din(n943),.dout(n944),.clk(gclk));
	jand g0881(.dina(w_n890_0[0]),.dinb(w_n845_0[0]),.dout(n945),.clk(gclk));
	jand g0882(.dina(w_n891_0[0]),.dinb(w_n842_0[0]),.dout(n946),.clk(gclk));
	jor g0883(.dina(n946),.dinb(n945),.dout(n947),.clk(gclk));
	jand g0884(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n948),.clk(gclk));
	jnot g0885(.din(n948),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_n888_0[0]),.dinb(w_n850_0[0]),.dout(n950),.clk(gclk));
	jand g0887(.dina(w_n889_0[0]),.dinb(w_n847_0[0]),.dout(n951),.clk(gclk));
	jor g0888(.dina(n951),.dinb(n950),.dout(n952),.clk(gclk));
	jand g0889(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n953),.clk(gclk));
	jnot g0890(.din(n953),.dout(n954),.clk(gclk));
	jand g0891(.dina(w_n886_0[0]),.dinb(w_n855_0[0]),.dout(n955),.clk(gclk));
	jand g0892(.dina(w_n887_0[0]),.dinb(w_n852_0[0]),.dout(n956),.clk(gclk));
	jor g0893(.dina(n956),.dinb(n955),.dout(n957),.clk(gclk));
	jand g0894(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n958),.clk(gclk));
	jnot g0895(.din(n958),.dout(n959),.clk(gclk));
	jand g0896(.dina(w_n884_0[0]),.dinb(w_n860_0[0]),.dout(n960),.clk(gclk));
	jand g0897(.dina(w_n885_0[0]),.dinb(w_n857_0[0]),.dout(n961),.clk(gclk));
	jor g0898(.dina(n961),.dinb(n960),.dout(n962),.clk(gclk));
	jand g0899(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n963),.clk(gclk));
	jnot g0900(.din(n963),.dout(n964),.clk(gclk));
	jand g0901(.dina(w_n882_0[0]),.dinb(w_n865_0[0]),.dout(n965),.clk(gclk));
	jand g0902(.dina(w_n883_0[0]),.dinb(w_n862_0[0]),.dout(n966),.clk(gclk));
	jor g0903(.dina(n966),.dinb(n965),.dout(n967),.clk(gclk));
	jand g0904(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n968),.clk(gclk));
	jnot g0905(.din(n968),.dout(n969),.clk(gclk));
	jand g0906(.dina(w_n880_0[0]),.dinb(w_n872_0[0]),.dout(n970),.clk(gclk));
	jand g0907(.dina(w_n881_0[0]),.dinb(w_n867_0[0]),.dout(n971),.clk(gclk));
	jor g0908(.dina(n971),.dinb(n970),.dout(n972),.clk(gclk));
	jand g0909(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n973),.clk(gclk));
	jnot g0910(.din(n973),.dout(n974),.clk(gclk));
	jand g0911(.dina(w_n879_0[0]),.dinb(w_n874_0[0]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(n976),.dinb(w_n877_0[0]),.dout(n977),.clk(gclk));
	jnot g0914(.din(n977),.dout(n978),.clk(gclk));
	jnot g0915(.din(w_n775_0[0]),.dout(n979),.clk(gclk));
	jand g0916(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n980),.clk(gclk));
	jand g0917(.dina(w_n980_0[1]),.dinb(n979),.dout(n981),.clk(gclk));
	jnot g0918(.din(n981),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_G307gat_2[2]),.dinb(w_G239gat_6[2]),.dout(n983),.clk(gclk));
	jxor g0920(.dina(w_n983_0[1]),.dinb(w_n982_0[1]),.dout(n984),.clk(gclk));
	jxor g0921(.dina(w_n984_0[1]),.dinb(w_n978_0[1]),.dout(n985),.clk(gclk));
	jxor g0922(.dina(w_n985_0[1]),.dinb(w_n974_0[1]),.dout(n986),.clk(gclk));
	jxor g0923(.dina(w_n986_0[1]),.dinb(w_n972_0[1]),.dout(n987),.clk(gclk));
	jxor g0924(.dina(w_n987_0[1]),.dinb(w_n969_0[1]),.dout(n988),.clk(gclk));
	jxor g0925(.dina(w_n988_0[1]),.dinb(w_n967_0[1]),.dout(n989),.clk(gclk));
	jxor g0926(.dina(w_n989_0[1]),.dinb(w_n964_0[1]),.dout(n990),.clk(gclk));
	jxor g0927(.dina(w_n990_0[1]),.dinb(w_n962_0[1]),.dout(n991),.clk(gclk));
	jxor g0928(.dina(w_n991_0[1]),.dinb(w_n959_0[1]),.dout(n992),.clk(gclk));
	jxor g0929(.dina(w_n992_0[1]),.dinb(w_n957_0[1]),.dout(n993),.clk(gclk));
	jxor g0930(.dina(w_n993_0[1]),.dinb(w_n954_0[1]),.dout(n994),.clk(gclk));
	jxor g0931(.dina(w_n994_0[1]),.dinb(w_n952_0[1]),.dout(n995),.clk(gclk));
	jxor g0932(.dina(w_n995_0[1]),.dinb(w_n949_0[1]),.dout(n996),.clk(gclk));
	jxor g0933(.dina(w_n996_0[1]),.dinb(w_n947_0[1]),.dout(n997),.clk(gclk));
	jxor g0934(.dina(w_n997_0[1]),.dinb(w_n944_0[1]),.dout(n998),.clk(gclk));
	jxor g0935(.dina(w_n998_0[1]),.dinb(w_n942_0[1]),.dout(n999),.clk(gclk));
	jxor g0936(.dina(w_n999_0[1]),.dinb(w_n939_0[1]),.dout(n1000),.clk(gclk));
	jxor g0937(.dina(w_n1000_0[1]),.dinb(w_n937_0[1]),.dout(n1001),.clk(gclk));
	jxor g0938(.dina(w_n1001_0[1]),.dinb(w_n934_0[1]),.dout(n1002),.clk(gclk));
	jxor g0939(.dina(w_n1002_0[1]),.dinb(w_n932_0[1]),.dout(n1003),.clk(gclk));
	jxor g0940(.dina(w_n1003_0[1]),.dinb(w_n929_0[1]),.dout(n1004),.clk(gclk));
	jxor g0941(.dina(w_n1004_0[1]),.dinb(w_n927_0[1]),.dout(n1005),.clk(gclk));
	jxor g0942(.dina(w_n1005_0[1]),.dinb(w_n924_0[1]),.dout(n1006),.clk(gclk));
	jxor g0943(.dina(w_n1006_0[1]),.dinb(w_n922_0[1]),.dout(n1007),.clk(gclk));
	jxor g0944(.dina(w_n1007_0[1]),.dinb(w_n916_0[1]),.dout(n1008),.clk(gclk));
	jnot g0945(.din(w_n1008_0[1]),.dout(n1009),.clk(gclk));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n915_0[2]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(n1010),.dinb(w_n911_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n910_0[1]),.dout(w_dff_A_Jo2F7egf8_2),.clk(gclk));
	jand g0949(.dina(w_n1011_0[0]),.dinb(w_n910_0[0]),.dout(n1013),.clk(gclk));
	jor g0950(.dina(w_n1009_0[0]),.dinb(w_n915_0[1]),.dout(n1014),.clk(gclk));
	jxor g0951(.dina(w_n1008_0[0]),.dinb(w_n915_0[0]),.dout(n1015),.clk(gclk));
	jor g0952(.dina(n1015),.dinb(w_n911_0[0]),.dout(n1016),.clk(gclk));
	jand g0953(.dina(n1016),.dinb(n1014),.dout(n1017),.clk(gclk));
	jand g0954(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1018),.clk(gclk));
	jnot g0955(.din(w_n1006_0[0]),.dout(n1019),.clk(gclk));
	jor g0956(.dina(n1019),.dinb(w_n922_0[0]),.dout(n1020),.clk(gclk));
	jor g0957(.dina(w_n1007_0[0]),.dinb(w_n916_0[0]),.dout(n1021),.clk(gclk));
	jand g0958(.dina(n1021),.dinb(n1020),.dout(n1022),.clk(gclk));
	jand g0959(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1023),.clk(gclk));
	jand g0960(.dina(w_n1004_0[0]),.dinb(w_n927_0[0]),.dout(n1024),.clk(gclk));
	jand g0961(.dina(w_n1005_0[0]),.dinb(w_n924_0[0]),.dout(n1025),.clk(gclk));
	jor g0962(.dina(n1025),.dinb(n1024),.dout(n1026),.clk(gclk));
	jand g0963(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1027),.clk(gclk));
	jnot g0964(.din(n1027),.dout(n1028),.clk(gclk));
	jand g0965(.dina(w_n1002_0[0]),.dinb(w_n932_0[0]),.dout(n1029),.clk(gclk));
	jand g0966(.dina(w_n1003_0[0]),.dinb(w_n929_0[0]),.dout(n1030),.clk(gclk));
	jor g0967(.dina(n1030),.dinb(n1029),.dout(n1031),.clk(gclk));
	jand g0968(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1032),.clk(gclk));
	jnot g0969(.din(n1032),.dout(n1033),.clk(gclk));
	jand g0970(.dina(w_n1000_0[0]),.dinb(w_n937_0[0]),.dout(n1034),.clk(gclk));
	jand g0971(.dina(w_n1001_0[0]),.dinb(w_n934_0[0]),.dout(n1035),.clk(gclk));
	jor g0972(.dina(n1035),.dinb(n1034),.dout(n1036),.clk(gclk));
	jand g0973(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1037),.clk(gclk));
	jnot g0974(.din(n1037),.dout(n1038),.clk(gclk));
	jand g0975(.dina(w_n998_0[0]),.dinb(w_n942_0[0]),.dout(n1039),.clk(gclk));
	jand g0976(.dina(w_n999_0[0]),.dinb(w_n939_0[0]),.dout(n1040),.clk(gclk));
	jor g0977(.dina(n1040),.dinb(n1039),.dout(n1041),.clk(gclk));
	jand g0978(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1042),.clk(gclk));
	jnot g0979(.din(n1042),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_n996_0[0]),.dinb(w_n947_0[0]),.dout(n1044),.clk(gclk));
	jand g0981(.dina(w_n997_0[0]),.dinb(w_n944_0[0]),.dout(n1045),.clk(gclk));
	jor g0982(.dina(n1045),.dinb(n1044),.dout(n1046),.clk(gclk));
	jand g0983(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1047),.clk(gclk));
	jnot g0984(.din(n1047),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_n994_0[0]),.dinb(w_n952_0[0]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n995_0[0]),.dinb(w_n949_0[0]),.dout(n1050),.clk(gclk));
	jor g0987(.dina(n1050),.dinb(n1049),.dout(n1051),.clk(gclk));
	jand g0988(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1052),.clk(gclk));
	jnot g0989(.din(n1052),.dout(n1053),.clk(gclk));
	jand g0990(.dina(w_n992_0[0]),.dinb(w_n957_0[0]),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n993_0[0]),.dinb(w_n954_0[0]),.dout(n1055),.clk(gclk));
	jor g0992(.dina(n1055),.dinb(n1054),.dout(n1056),.clk(gclk));
	jand g0993(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1057),.clk(gclk));
	jnot g0994(.din(n1057),.dout(n1058),.clk(gclk));
	jand g0995(.dina(w_n990_0[0]),.dinb(w_n962_0[0]),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n991_0[0]),.dinb(w_n959_0[0]),.dout(n1060),.clk(gclk));
	jor g0997(.dina(n1060),.dinb(n1059),.dout(n1061),.clk(gclk));
	jand g0998(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1062),.clk(gclk));
	jnot g0999(.din(n1062),.dout(n1063),.clk(gclk));
	jand g1000(.dina(w_n988_0[0]),.dinb(w_n967_0[0]),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n989_0[0]),.dinb(w_n964_0[0]),.dout(n1065),.clk(gclk));
	jor g1002(.dina(n1065),.dinb(n1064),.dout(n1066),.clk(gclk));
	jand g1003(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1067),.clk(gclk));
	jnot g1004(.din(n1067),.dout(n1068),.clk(gclk));
	jand g1005(.dina(w_n986_0[0]),.dinb(w_n972_0[0]),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n987_0[0]),.dinb(w_n969_0[0]),.dout(n1070),.clk(gclk));
	jor g1007(.dina(n1070),.dinb(n1069),.dout(n1071),.clk(gclk));
	jand g1008(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1072),.clk(gclk));
	jnot g1009(.din(n1072),.dout(n1073),.clk(gclk));
	jand g1010(.dina(w_n984_0[0]),.dinb(w_n978_0[0]),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n985_0[0]),.dinb(w_n974_0[0]),.dout(n1075),.clk(gclk));
	jor g1012(.dina(n1075),.dinb(n1074),.dout(n1076),.clk(gclk));
	jand g1013(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1077),.clk(gclk));
	jand g1014(.dina(w_G307gat_2[1]),.dinb(w_G256gat_6[2]),.dout(n1078),.clk(gclk));
	jor g1015(.dina(w_n983_0[0]),.dinb(w_n982_0[0]),.dout(n1079),.clk(gclk));
	jand g1016(.dina(n1079),.dinb(w_n980_0[0]),.dout(n1080),.clk(gclk));
	jxor g1017(.dina(w_n1080_0[1]),.dinb(w_n1078_0[1]),.dout(n1081),.clk(gclk));
	jnot g1018(.din(n1081),.dout(n1082),.clk(gclk));
	jxor g1019(.dina(w_n1082_0[1]),.dinb(w_n1077_0[1]),.dout(n1083),.clk(gclk));
	jxor g1020(.dina(w_n1083_0[1]),.dinb(w_n1076_0[1]),.dout(n1084),.clk(gclk));
	jxor g1021(.dina(w_n1084_0[1]),.dinb(w_n1073_0[1]),.dout(n1085),.clk(gclk));
	jxor g1022(.dina(w_n1085_0[1]),.dinb(w_n1071_0[1]),.dout(n1086),.clk(gclk));
	jxor g1023(.dina(w_n1086_0[1]),.dinb(w_n1068_0[1]),.dout(n1087),.clk(gclk));
	jxor g1024(.dina(w_n1087_0[1]),.dinb(w_n1066_0[1]),.dout(n1088),.clk(gclk));
	jxor g1025(.dina(w_n1088_0[1]),.dinb(w_n1063_0[1]),.dout(n1089),.clk(gclk));
	jxor g1026(.dina(w_n1089_0[1]),.dinb(w_n1061_0[1]),.dout(n1090),.clk(gclk));
	jxor g1027(.dina(w_n1090_0[1]),.dinb(w_n1058_0[1]),.dout(n1091),.clk(gclk));
	jxor g1028(.dina(w_n1091_0[1]),.dinb(w_n1056_0[1]),.dout(n1092),.clk(gclk));
	jxor g1029(.dina(w_n1092_0[1]),.dinb(w_n1053_0[1]),.dout(n1093),.clk(gclk));
	jxor g1030(.dina(w_n1093_0[1]),.dinb(w_n1051_0[1]),.dout(n1094),.clk(gclk));
	jxor g1031(.dina(w_n1094_0[1]),.dinb(w_n1048_0[1]),.dout(n1095),.clk(gclk));
	jxor g1032(.dina(w_n1095_0[1]),.dinb(w_n1046_0[1]),.dout(n1096),.clk(gclk));
	jxor g1033(.dina(w_n1096_0[1]),.dinb(w_n1043_0[1]),.dout(n1097),.clk(gclk));
	jxor g1034(.dina(w_n1097_0[1]),.dinb(w_n1041_0[1]),.dout(n1098),.clk(gclk));
	jxor g1035(.dina(w_n1098_0[1]),.dinb(w_n1038_0[1]),.dout(n1099),.clk(gclk));
	jxor g1036(.dina(w_n1099_0[1]),.dinb(w_n1036_0[1]),.dout(n1100),.clk(gclk));
	jxor g1037(.dina(w_n1100_0[1]),.dinb(w_n1033_0[1]),.dout(n1101),.clk(gclk));
	jxor g1038(.dina(w_n1101_0[1]),.dinb(w_n1031_0[1]),.dout(n1102),.clk(gclk));
	jxor g1039(.dina(w_n1102_0[1]),.dinb(w_n1028_0[1]),.dout(n1103),.clk(gclk));
	jxor g1040(.dina(w_n1103_0[1]),.dinb(w_n1026_0[1]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(n1104),.dout(n1105),.clk(gclk));
	jxor g1042(.dina(w_n1105_0[1]),.dinb(w_n1023_0[1]),.dout(n1106),.clk(gclk));
	jxor g1043(.dina(w_n1106_0[1]),.dinb(w_n1022_0[1]),.dout(n1107),.clk(gclk));
	jxor g1044(.dina(w_n1107_0[1]),.dinb(w_n1018_0[1]),.dout(n1108),.clk(gclk));
	jxor g1045(.dina(w_n1108_0[1]),.dinb(w_n1017_0[1]),.dout(n1109),.clk(gclk));
	jnot g1046(.din(w_n1109_0[1]),.dout(n1110),.clk(gclk));
	jxor g1047(.dina(n1110),.dinb(w_n1013_0[1]),.dout(w_dff_A_4izfRJkS6_2),.clk(gclk));
	jnot g1048(.din(w_n1108_0[0]),.dout(n1112),.clk(gclk));
	jor g1049(.dina(n1112),.dinb(w_n1017_0[0]),.dout(n1113),.clk(gclk));
	jor g1050(.dina(w_n1109_0[0]),.dinb(w_n1013_0[0]),.dout(n1114),.clk(gclk));
	jand g1051(.dina(n1114),.dinb(w_dff_B_nlpNDxfO7_1),.dout(n1115),.clk(gclk));
	jnot g1052(.din(w_n1106_0[0]),.dout(n1116),.clk(gclk));
	jor g1053(.dina(n1116),.dinb(w_n1022_0[0]),.dout(n1117),.clk(gclk));
	jor g1054(.dina(w_n1107_0[0]),.dinb(w_n1018_0[0]),.dout(n1118),.clk(gclk));
	jand g1055(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jand g1056(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1120),.clk(gclk));
	jand g1057(.dina(w_n1103_0[0]),.dinb(w_n1026_0[0]),.dout(n1121),.clk(gclk));
	jnot g1058(.din(n1121),.dout(n1122),.clk(gclk));
	jor g1059(.dina(w_n1105_0[0]),.dinb(w_n1023_0[0]),.dout(n1123),.clk(gclk));
	jand g1060(.dina(n1123),.dinb(n1122),.dout(n1124),.clk(gclk));
	jand g1061(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1125),.clk(gclk));
	jnot g1062(.din(n1125),.dout(n1126),.clk(gclk));
	jand g1063(.dina(w_n1101_0[0]),.dinb(w_n1031_0[0]),.dout(n1127),.clk(gclk));
	jand g1064(.dina(w_n1102_0[0]),.dinb(w_n1028_0[0]),.dout(n1128),.clk(gclk));
	jor g1065(.dina(n1128),.dinb(n1127),.dout(n1129),.clk(gclk));
	jand g1066(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1130),.clk(gclk));
	jnot g1067(.din(n1130),.dout(n1131),.clk(gclk));
	jand g1068(.dina(w_n1099_0[0]),.dinb(w_n1036_0[0]),.dout(n1132),.clk(gclk));
	jand g1069(.dina(w_n1100_0[0]),.dinb(w_n1033_0[0]),.dout(n1133),.clk(gclk));
	jor g1070(.dina(n1133),.dinb(n1132),.dout(n1134),.clk(gclk));
	jand g1071(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1135),.clk(gclk));
	jnot g1072(.din(n1135),.dout(n1136),.clk(gclk));
	jand g1073(.dina(w_n1097_0[0]),.dinb(w_n1041_0[0]),.dout(n1137),.clk(gclk));
	jand g1074(.dina(w_n1098_0[0]),.dinb(w_n1038_0[0]),.dout(n1138),.clk(gclk));
	jor g1075(.dina(n1138),.dinb(n1137),.dout(n1139),.clk(gclk));
	jand g1076(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1140),.clk(gclk));
	jnot g1077(.din(n1140),.dout(n1141),.clk(gclk));
	jand g1078(.dina(w_n1095_0[0]),.dinb(w_n1046_0[0]),.dout(n1142),.clk(gclk));
	jand g1079(.dina(w_n1096_0[0]),.dinb(w_n1043_0[0]),.dout(n1143),.clk(gclk));
	jor g1080(.dina(n1143),.dinb(n1142),.dout(n1144),.clk(gclk));
	jand g1081(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1145),.clk(gclk));
	jnot g1082(.din(n1145),.dout(n1146),.clk(gclk));
	jand g1083(.dina(w_n1093_0[0]),.dinb(w_n1051_0[0]),.dout(n1147),.clk(gclk));
	jand g1084(.dina(w_n1094_0[0]),.dinb(w_n1048_0[0]),.dout(n1148),.clk(gclk));
	jor g1085(.dina(n1148),.dinb(n1147),.dout(n1149),.clk(gclk));
	jand g1086(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1150),.clk(gclk));
	jnot g1087(.din(n1150),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_n1091_0[0]),.dinb(w_n1056_0[0]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1092_0[0]),.dinb(w_n1053_0[0]),.dout(n1153),.clk(gclk));
	jor g1090(.dina(n1153),.dinb(n1152),.dout(n1154),.clk(gclk));
	jand g1091(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1155),.clk(gclk));
	jnot g1092(.din(n1155),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_n1089_0[0]),.dinb(w_n1061_0[0]),.dout(n1157),.clk(gclk));
	jand g1094(.dina(w_n1090_0[0]),.dinb(w_n1058_0[0]),.dout(n1158),.clk(gclk));
	jor g1095(.dina(n1158),.dinb(n1157),.dout(n1159),.clk(gclk));
	jand g1096(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1160),.clk(gclk));
	jnot g1097(.din(n1160),.dout(n1161),.clk(gclk));
	jand g1098(.dina(w_n1087_0[0]),.dinb(w_n1066_0[0]),.dout(n1162),.clk(gclk));
	jand g1099(.dina(w_n1088_0[0]),.dinb(w_n1063_0[0]),.dout(n1163),.clk(gclk));
	jor g1100(.dina(n1163),.dinb(n1162),.dout(n1164),.clk(gclk));
	jand g1101(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1165),.clk(gclk));
	jnot g1102(.din(n1165),.dout(n1166),.clk(gclk));
	jand g1103(.dina(w_n1085_0[0]),.dinb(w_n1071_0[0]),.dout(n1167),.clk(gclk));
	jand g1104(.dina(w_n1086_0[0]),.dinb(w_n1068_0[0]),.dout(n1168),.clk(gclk));
	jor g1105(.dina(n1168),.dinb(n1167),.dout(n1169),.clk(gclk));
	jand g1106(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1170),.clk(gclk));
	jnot g1107(.din(n1170),.dout(n1171),.clk(gclk));
	jand g1108(.dina(w_n1083_0[0]),.dinb(w_n1076_0[0]),.dout(n1172),.clk(gclk));
	jand g1109(.dina(w_n1084_0[0]),.dinb(w_n1073_0[0]),.dout(n1173),.clk(gclk));
	jor g1110(.dina(n1173),.dinb(n1172),.dout(n1174),.clk(gclk));
	jand g1111(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1175),.clk(gclk));
	jand g1112(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1176),.clk(gclk));
	jor g1113(.dina(w_n1080_0[0]),.dinb(w_n1078_0[0]),.dout(n1177),.clk(gclk));
	jor g1114(.dina(w_n1082_0[0]),.dinb(w_n1077_0[0]),.dout(n1178),.clk(gclk));
	jand g1115(.dina(n1178),.dinb(n1177),.dout(n1179),.clk(gclk));
	jxor g1116(.dina(w_n1179_0[1]),.dinb(w_n1176_0[1]),.dout(n1180),.clk(gclk));
	jnot g1117(.din(n1180),.dout(n1181),.clk(gclk));
	jxor g1118(.dina(w_n1181_0[1]),.dinb(w_n1175_0[1]),.dout(n1182),.clk(gclk));
	jxor g1119(.dina(w_n1182_0[1]),.dinb(w_n1174_0[1]),.dout(n1183),.clk(gclk));
	jxor g1120(.dina(w_n1183_0[1]),.dinb(w_n1171_0[1]),.dout(n1184),.clk(gclk));
	jxor g1121(.dina(w_n1184_0[1]),.dinb(w_n1169_0[1]),.dout(n1185),.clk(gclk));
	jxor g1122(.dina(w_n1185_0[1]),.dinb(w_n1166_0[1]),.dout(n1186),.clk(gclk));
	jxor g1123(.dina(w_n1186_0[1]),.dinb(w_n1164_0[1]),.dout(n1187),.clk(gclk));
	jxor g1124(.dina(w_n1187_0[1]),.dinb(w_n1161_0[1]),.dout(n1188),.clk(gclk));
	jxor g1125(.dina(w_n1188_0[1]),.dinb(w_n1159_0[1]),.dout(n1189),.clk(gclk));
	jxor g1126(.dina(w_n1189_0[1]),.dinb(w_n1156_0[1]),.dout(n1190),.clk(gclk));
	jxor g1127(.dina(w_n1190_0[1]),.dinb(w_n1154_0[1]),.dout(n1191),.clk(gclk));
	jxor g1128(.dina(w_n1191_0[1]),.dinb(w_n1151_0[1]),.dout(n1192),.clk(gclk));
	jxor g1129(.dina(w_n1192_0[1]),.dinb(w_n1149_0[1]),.dout(n1193),.clk(gclk));
	jxor g1130(.dina(w_n1193_0[1]),.dinb(w_n1146_0[1]),.dout(n1194),.clk(gclk));
	jxor g1131(.dina(w_n1194_0[1]),.dinb(w_n1144_0[1]),.dout(n1195),.clk(gclk));
	jxor g1132(.dina(w_n1195_0[1]),.dinb(w_n1141_0[1]),.dout(n1196),.clk(gclk));
	jxor g1133(.dina(w_n1196_0[1]),.dinb(w_n1139_0[1]),.dout(n1197),.clk(gclk));
	jxor g1134(.dina(w_n1197_0[1]),.dinb(w_n1136_0[1]),.dout(n1198),.clk(gclk));
	jxor g1135(.dina(w_n1198_0[1]),.dinb(w_n1134_0[1]),.dout(n1199),.clk(gclk));
	jxor g1136(.dina(w_n1199_0[1]),.dinb(w_n1131_0[1]),.dout(n1200),.clk(gclk));
	jxor g1137(.dina(w_n1200_0[1]),.dinb(w_n1129_0[1]),.dout(n1201),.clk(gclk));
	jxor g1138(.dina(w_n1201_0[1]),.dinb(w_n1126_0[1]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jxor g1140(.dina(w_n1203_0[1]),.dinb(w_n1124_0[1]),.dout(n1204),.clk(gclk));
	jnot g1141(.din(n1204),.dout(n1205),.clk(gclk));
	jxor g1142(.dina(w_n1205_0[1]),.dinb(w_n1120_0[1]),.dout(n1206),.clk(gclk));
	jxor g1143(.dina(w_n1206_0[1]),.dinb(w_n1119_0[1]),.dout(n1207),.clk(gclk));
	jnot g1144(.din(w_n1207_0[1]),.dout(n1208),.clk(gclk));
	jxor g1145(.dina(n1208),.dinb(w_n1115_0[1]),.dout(w_dff_A_x9VZLpLG1_2),.clk(gclk));
	jnot g1146(.din(w_n1206_0[0]),.dout(n1210),.clk(gclk));
	jor g1147(.dina(n1210),.dinb(w_n1119_0[0]),.dout(n1211),.clk(gclk));
	jor g1148(.dina(w_n1207_0[0]),.dinb(w_n1115_0[0]),.dout(n1212),.clk(gclk));
	jand g1149(.dina(n1212),.dinb(w_dff_B_AmhI8UHA1_1),.dout(n1213),.clk(gclk));
	jor g1150(.dina(w_n1203_0[0]),.dinb(w_n1124_0[0]),.dout(n1214),.clk(gclk));
	jor g1151(.dina(w_n1205_0[0]),.dinb(w_n1120_0[0]),.dout(n1215),.clk(gclk));
	jand g1152(.dina(n1215),.dinb(n1214),.dout(n1216),.clk(gclk));
	jand g1153(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1217),.clk(gclk));
	jand g1154(.dina(w_n1200_0[0]),.dinb(w_n1129_0[0]),.dout(n1218),.clk(gclk));
	jand g1155(.dina(w_n1201_0[0]),.dinb(w_n1126_0[0]),.dout(n1219),.clk(gclk));
	jor g1156(.dina(n1219),.dinb(n1218),.dout(n1220),.clk(gclk));
	jand g1157(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1221),.clk(gclk));
	jnot g1158(.din(n1221),.dout(n1222),.clk(gclk));
	jand g1159(.dina(w_n1198_0[0]),.dinb(w_n1134_0[0]),.dout(n1223),.clk(gclk));
	jand g1160(.dina(w_n1199_0[0]),.dinb(w_n1131_0[0]),.dout(n1224),.clk(gclk));
	jor g1161(.dina(n1224),.dinb(n1223),.dout(n1225),.clk(gclk));
	jand g1162(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1226),.clk(gclk));
	jnot g1163(.din(n1226),.dout(n1227),.clk(gclk));
	jand g1164(.dina(w_n1196_0[0]),.dinb(w_n1139_0[0]),.dout(n1228),.clk(gclk));
	jand g1165(.dina(w_n1197_0[0]),.dinb(w_n1136_0[0]),.dout(n1229),.clk(gclk));
	jor g1166(.dina(n1229),.dinb(n1228),.dout(n1230),.clk(gclk));
	jand g1167(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1231),.clk(gclk));
	jnot g1168(.din(n1231),.dout(n1232),.clk(gclk));
	jand g1169(.dina(w_n1194_0[0]),.dinb(w_n1144_0[0]),.dout(n1233),.clk(gclk));
	jand g1170(.dina(w_n1195_0[0]),.dinb(w_n1141_0[0]),.dout(n1234),.clk(gclk));
	jor g1171(.dina(n1234),.dinb(n1233),.dout(n1235),.clk(gclk));
	jand g1172(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1236),.clk(gclk));
	jnot g1173(.din(n1236),.dout(n1237),.clk(gclk));
	jand g1174(.dina(w_n1192_0[0]),.dinb(w_n1149_0[0]),.dout(n1238),.clk(gclk));
	jand g1175(.dina(w_n1193_0[0]),.dinb(w_n1146_0[0]),.dout(n1239),.clk(gclk));
	jor g1176(.dina(n1239),.dinb(n1238),.dout(n1240),.clk(gclk));
	jand g1177(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1241),.clk(gclk));
	jnot g1178(.din(n1241),.dout(n1242),.clk(gclk));
	jand g1179(.dina(w_n1190_0[0]),.dinb(w_n1154_0[0]),.dout(n1243),.clk(gclk));
	jand g1180(.dina(w_n1191_0[0]),.dinb(w_n1151_0[0]),.dout(n1244),.clk(gclk));
	jor g1181(.dina(n1244),.dinb(n1243),.dout(n1245),.clk(gclk));
	jand g1182(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1246),.clk(gclk));
	jnot g1183(.din(n1246),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_n1188_0[0]),.dinb(w_n1159_0[0]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1189_0[0]),.dinb(w_n1156_0[0]),.dout(n1249),.clk(gclk));
	jor g1186(.dina(n1249),.dinb(n1248),.dout(n1250),.clk(gclk));
	jand g1187(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1251),.clk(gclk));
	jnot g1188(.din(n1251),.dout(n1252),.clk(gclk));
	jand g1189(.dina(w_n1186_0[0]),.dinb(w_n1164_0[0]),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1187_0[0]),.dinb(w_n1161_0[0]),.dout(n1254),.clk(gclk));
	jor g1191(.dina(n1254),.dinb(n1253),.dout(n1255),.clk(gclk));
	jand g1192(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1256),.clk(gclk));
	jnot g1193(.din(n1256),.dout(n1257),.clk(gclk));
	jand g1194(.dina(w_n1184_0[0]),.dinb(w_n1169_0[0]),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1185_0[0]),.dinb(w_n1166_0[0]),.dout(n1259),.clk(gclk));
	jor g1196(.dina(n1259),.dinb(n1258),.dout(n1260),.clk(gclk));
	jand g1197(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1261),.clk(gclk));
	jnot g1198(.din(n1261),.dout(n1262),.clk(gclk));
	jand g1199(.dina(w_n1182_0[0]),.dinb(w_n1174_0[0]),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1183_0[0]),.dinb(w_n1171_0[0]),.dout(n1264),.clk(gclk));
	jor g1201(.dina(n1264),.dinb(n1263),.dout(n1265),.clk(gclk));
	jand g1202(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1266),.clk(gclk));
	jand g1203(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1267),.clk(gclk));
	jor g1204(.dina(w_n1179_0[0]),.dinb(w_n1176_0[0]),.dout(n1268),.clk(gclk));
	jor g1205(.dina(w_n1181_0[0]),.dinb(w_n1175_0[0]),.dout(n1269),.clk(gclk));
	jand g1206(.dina(n1269),.dinb(n1268),.dout(n1270),.clk(gclk));
	jxor g1207(.dina(w_n1270_0[1]),.dinb(w_n1267_0[1]),.dout(n1271),.clk(gclk));
	jnot g1208(.din(n1271),.dout(n1272),.clk(gclk));
	jxor g1209(.dina(w_n1272_0[1]),.dinb(w_n1266_0[1]),.dout(n1273),.clk(gclk));
	jxor g1210(.dina(w_n1273_0[1]),.dinb(w_n1265_0[1]),.dout(n1274),.clk(gclk));
	jxor g1211(.dina(w_n1274_0[1]),.dinb(w_n1262_0[1]),.dout(n1275),.clk(gclk));
	jxor g1212(.dina(w_n1275_0[1]),.dinb(w_n1260_0[1]),.dout(n1276),.clk(gclk));
	jxor g1213(.dina(w_n1276_0[1]),.dinb(w_n1257_0[1]),.dout(n1277),.clk(gclk));
	jxor g1214(.dina(w_n1277_0[1]),.dinb(w_n1255_0[1]),.dout(n1278),.clk(gclk));
	jxor g1215(.dina(w_n1278_0[1]),.dinb(w_n1252_0[1]),.dout(n1279),.clk(gclk));
	jxor g1216(.dina(w_n1279_0[1]),.dinb(w_n1250_0[1]),.dout(n1280),.clk(gclk));
	jxor g1217(.dina(w_n1280_0[1]),.dinb(w_n1247_0[1]),.dout(n1281),.clk(gclk));
	jxor g1218(.dina(w_n1281_0[1]),.dinb(w_n1245_0[1]),.dout(n1282),.clk(gclk));
	jxor g1219(.dina(w_n1282_0[1]),.dinb(w_n1242_0[1]),.dout(n1283),.clk(gclk));
	jxor g1220(.dina(w_n1283_0[1]),.dinb(w_n1240_0[1]),.dout(n1284),.clk(gclk));
	jxor g1221(.dina(w_n1284_0[1]),.dinb(w_n1237_0[1]),.dout(n1285),.clk(gclk));
	jxor g1222(.dina(w_n1285_0[1]),.dinb(w_n1235_0[1]),.dout(n1286),.clk(gclk));
	jxor g1223(.dina(w_n1286_0[1]),.dinb(w_n1232_0[1]),.dout(n1287),.clk(gclk));
	jxor g1224(.dina(w_n1287_0[1]),.dinb(w_n1230_0[1]),.dout(n1288),.clk(gclk));
	jxor g1225(.dina(w_n1288_0[1]),.dinb(w_n1227_0[1]),.dout(n1289),.clk(gclk));
	jxor g1226(.dina(w_n1289_0[1]),.dinb(w_n1225_0[1]),.dout(n1290),.clk(gclk));
	jxor g1227(.dina(w_n1290_0[1]),.dinb(w_n1222_0[1]),.dout(n1291),.clk(gclk));
	jxor g1228(.dina(w_n1291_0[1]),.dinb(w_n1220_0[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jxor g1230(.dina(w_n1293_0[1]),.dinb(w_n1217_0[1]),.dout(n1294),.clk(gclk));
	jxor g1231(.dina(w_n1294_0[1]),.dinb(w_n1216_0[1]),.dout(n1295),.clk(gclk));
	jnot g1232(.din(w_n1295_0[1]),.dout(n1296),.clk(gclk));
	jxor g1233(.dina(w_dff_B_A72U7TVO7_0),.dinb(w_n1213_0[1]),.dout(w_dff_A_4IuXdUMj6_2),.clk(gclk));
	jnot g1234(.din(w_n1294_0[0]),.dout(n1298),.clk(gclk));
	jor g1235(.dina(n1298),.dinb(w_n1216_0[0]),.dout(n1299),.clk(gclk));
	jor g1236(.dina(w_n1295_0[0]),.dinb(w_n1213_0[0]),.dout(n1300),.clk(gclk));
	jand g1237(.dina(n1300),.dinb(w_dff_B_vtqfyuMu0_1),.dout(n1301),.clk(gclk));
	jnot g1238(.din(w_n1220_0[0]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(w_n1291_0[0]),.dout(n1303),.clk(gclk));
	jor g1240(.dina(n1303),.dinb(n1302),.dout(n1304),.clk(gclk));
	jor g1241(.dina(w_n1293_0[0]),.dinb(w_n1217_0[0]),.dout(n1305),.clk(gclk));
	jand g1242(.dina(n1305),.dinb(n1304),.dout(n1306),.clk(gclk));
	jand g1243(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1307),.clk(gclk));
	jand g1244(.dina(w_n1289_0[0]),.dinb(w_n1225_0[0]),.dout(n1308),.clk(gclk));
	jand g1245(.dina(w_n1290_0[0]),.dinb(w_n1222_0[0]),.dout(n1309),.clk(gclk));
	jor g1246(.dina(n1309),.dinb(n1308),.dout(n1310),.clk(gclk));
	jand g1247(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1311),.clk(gclk));
	jnot g1248(.din(n1311),.dout(n1312),.clk(gclk));
	jand g1249(.dina(w_n1287_0[0]),.dinb(w_n1230_0[0]),.dout(n1313),.clk(gclk));
	jand g1250(.dina(w_n1288_0[0]),.dinb(w_n1227_0[0]),.dout(n1314),.clk(gclk));
	jor g1251(.dina(n1314),.dinb(n1313),.dout(n1315),.clk(gclk));
	jand g1252(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1316),.clk(gclk));
	jnot g1253(.din(n1316),.dout(n1317),.clk(gclk));
	jand g1254(.dina(w_n1285_0[0]),.dinb(w_n1235_0[0]),.dout(n1318),.clk(gclk));
	jand g1255(.dina(w_n1286_0[0]),.dinb(w_n1232_0[0]),.dout(n1319),.clk(gclk));
	jor g1256(.dina(n1319),.dinb(n1318),.dout(n1320),.clk(gclk));
	jand g1257(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1321),.clk(gclk));
	jnot g1258(.din(n1321),.dout(n1322),.clk(gclk));
	jand g1259(.dina(w_n1283_0[0]),.dinb(w_n1240_0[0]),.dout(n1323),.clk(gclk));
	jand g1260(.dina(w_n1284_0[0]),.dinb(w_n1237_0[0]),.dout(n1324),.clk(gclk));
	jor g1261(.dina(n1324),.dinb(n1323),.dout(n1325),.clk(gclk));
	jand g1262(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(n1326),.dout(n1327),.clk(gclk));
	jand g1264(.dina(w_n1281_0[0]),.dinb(w_n1245_0[0]),.dout(n1328),.clk(gclk));
	jand g1265(.dina(w_n1282_0[0]),.dinb(w_n1242_0[0]),.dout(n1329),.clk(gclk));
	jor g1266(.dina(n1329),.dinb(n1328),.dout(n1330),.clk(gclk));
	jand g1267(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1331),.clk(gclk));
	jnot g1268(.din(n1331),.dout(n1332),.clk(gclk));
	jand g1269(.dina(w_n1279_0[0]),.dinb(w_n1250_0[0]),.dout(n1333),.clk(gclk));
	jand g1270(.dina(w_n1280_0[0]),.dinb(w_n1247_0[0]),.dout(n1334),.clk(gclk));
	jor g1271(.dina(n1334),.dinb(n1333),.dout(n1335),.clk(gclk));
	jand g1272(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1336),.clk(gclk));
	jnot g1273(.din(n1336),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_n1277_0[0]),.dinb(w_n1255_0[0]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1278_0[0]),.dinb(w_n1252_0[0]),.dout(n1339),.clk(gclk));
	jor g1276(.dina(n1339),.dinb(n1338),.dout(n1340),.clk(gclk));
	jand g1277(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1341),.clk(gclk));
	jnot g1278(.din(n1341),.dout(n1342),.clk(gclk));
	jand g1279(.dina(w_n1275_0[0]),.dinb(w_n1260_0[0]),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1276_0[0]),.dinb(w_n1257_0[0]),.dout(n1344),.clk(gclk));
	jor g1281(.dina(n1344),.dinb(n1343),.dout(n1345),.clk(gclk));
	jand g1282(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1346),.clk(gclk));
	jnot g1283(.din(n1346),.dout(n1347),.clk(gclk));
	jand g1284(.dina(w_n1273_0[0]),.dinb(w_n1265_0[0]),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1274_0[0]),.dinb(w_n1262_0[0]),.dout(n1349),.clk(gclk));
	jor g1286(.dina(n1349),.dinb(n1348),.dout(n1350),.clk(gclk));
	jand g1287(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1351),.clk(gclk));
	jand g1288(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1352),.clk(gclk));
	jor g1289(.dina(w_n1270_0[0]),.dinb(w_n1267_0[0]),.dout(n1353),.clk(gclk));
	jor g1290(.dina(w_n1272_0[0]),.dinb(w_n1266_0[0]),.dout(n1354),.clk(gclk));
	jand g1291(.dina(n1354),.dinb(n1353),.dout(n1355),.clk(gclk));
	jxor g1292(.dina(w_n1355_0[1]),.dinb(w_n1352_0[1]),.dout(n1356),.clk(gclk));
	jnot g1293(.din(n1356),.dout(n1357),.clk(gclk));
	jxor g1294(.dina(w_n1357_0[1]),.dinb(w_n1351_0[1]),.dout(n1358),.clk(gclk));
	jxor g1295(.dina(w_n1358_0[1]),.dinb(w_n1350_0[1]),.dout(n1359),.clk(gclk));
	jxor g1296(.dina(w_n1359_0[1]),.dinb(w_n1347_0[1]),.dout(n1360),.clk(gclk));
	jxor g1297(.dina(w_n1360_0[1]),.dinb(w_n1345_0[1]),.dout(n1361),.clk(gclk));
	jxor g1298(.dina(w_n1361_0[1]),.dinb(w_n1342_0[1]),.dout(n1362),.clk(gclk));
	jxor g1299(.dina(w_n1362_0[1]),.dinb(w_n1340_0[1]),.dout(n1363),.clk(gclk));
	jxor g1300(.dina(w_n1363_0[1]),.dinb(w_n1337_0[1]),.dout(n1364),.clk(gclk));
	jxor g1301(.dina(w_n1364_0[1]),.dinb(w_n1335_0[1]),.dout(n1365),.clk(gclk));
	jxor g1302(.dina(w_n1365_0[1]),.dinb(w_n1332_0[1]),.dout(n1366),.clk(gclk));
	jxor g1303(.dina(w_n1366_0[1]),.dinb(w_n1330_0[1]),.dout(n1367),.clk(gclk));
	jxor g1304(.dina(w_n1367_0[1]),.dinb(w_n1327_0[1]),.dout(n1368),.clk(gclk));
	jxor g1305(.dina(w_n1368_0[1]),.dinb(w_n1325_0[1]),.dout(n1369),.clk(gclk));
	jxor g1306(.dina(w_n1369_0[1]),.dinb(w_n1322_0[1]),.dout(n1370),.clk(gclk));
	jxor g1307(.dina(w_n1370_0[1]),.dinb(w_n1320_0[1]),.dout(n1371),.clk(gclk));
	jxor g1308(.dina(w_n1371_0[1]),.dinb(w_n1317_0[1]),.dout(n1372),.clk(gclk));
	jxor g1309(.dina(w_n1372_0[1]),.dinb(w_n1315_0[1]),.dout(n1373),.clk(gclk));
	jxor g1310(.dina(w_n1373_0[1]),.dinb(w_n1312_0[1]),.dout(n1374),.clk(gclk));
	jxor g1311(.dina(w_n1374_0[1]),.dinb(w_n1310_0[1]),.dout(n1375),.clk(gclk));
	jnot g1312(.din(n1375),.dout(n1376),.clk(gclk));
	jxor g1313(.dina(w_n1376_0[1]),.dinb(w_n1307_0[1]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jxor g1315(.dina(w_n1378_0[1]),.dinb(w_n1306_0[1]),.dout(n1379),.clk(gclk));
	jxor g1316(.dina(w_n1379_0[1]),.dinb(w_n1301_0[1]),.dout(w_dff_A_UJSpteTt5_2),.clk(gclk));
	jor g1317(.dina(w_n1378_0[0]),.dinb(w_n1306_0[0]),.dout(n1381),.clk(gclk));
	jnot g1318(.din(w_n1379_0[0]),.dout(n1382),.clk(gclk));
	jor g1319(.dina(w_dff_B_d05Jrrm95_0),.dinb(w_n1301_0[0]),.dout(n1383),.clk(gclk));
	jand g1320(.dina(n1383),.dinb(w_dff_B_qh4TqmUH5_1),.dout(n1384),.clk(gclk));
	jnot g1321(.din(w_n1310_0[0]),.dout(n1385),.clk(gclk));
	jnot g1322(.din(w_n1374_0[0]),.dout(n1386),.clk(gclk));
	jor g1323(.dina(n1386),.dinb(n1385),.dout(n1387),.clk(gclk));
	jor g1324(.dina(w_n1376_0[0]),.dinb(w_n1307_0[0]),.dout(n1388),.clk(gclk));
	jand g1325(.dina(n1388),.dinb(n1387),.dout(n1389),.clk(gclk));
	jand g1326(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1390),.clk(gclk));
	jand g1327(.dina(w_n1372_0[0]),.dinb(w_n1315_0[0]),.dout(n1391),.clk(gclk));
	jand g1328(.dina(w_n1373_0[0]),.dinb(w_n1312_0[0]),.dout(n1392),.clk(gclk));
	jor g1329(.dina(n1392),.dinb(n1391),.dout(n1393),.clk(gclk));
	jand g1330(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1394),.clk(gclk));
	jnot g1331(.din(n1394),.dout(n1395),.clk(gclk));
	jand g1332(.dina(w_n1370_0[0]),.dinb(w_n1320_0[0]),.dout(n1396),.clk(gclk));
	jand g1333(.dina(w_n1371_0[0]),.dinb(w_n1317_0[0]),.dout(n1397),.clk(gclk));
	jor g1334(.dina(n1397),.dinb(n1396),.dout(n1398),.clk(gclk));
	jand g1335(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1399),.clk(gclk));
	jnot g1336(.din(n1399),.dout(n1400),.clk(gclk));
	jand g1337(.dina(w_n1368_0[0]),.dinb(w_n1325_0[0]),.dout(n1401),.clk(gclk));
	jand g1338(.dina(w_n1369_0[0]),.dinb(w_n1322_0[0]),.dout(n1402),.clk(gclk));
	jor g1339(.dina(n1402),.dinb(n1401),.dout(n1403),.clk(gclk));
	jand g1340(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1404),.clk(gclk));
	jnot g1341(.din(n1404),.dout(n1405),.clk(gclk));
	jand g1342(.dina(w_n1366_0[0]),.dinb(w_n1330_0[0]),.dout(n1406),.clk(gclk));
	jand g1343(.dina(w_n1367_0[0]),.dinb(w_n1327_0[0]),.dout(n1407),.clk(gclk));
	jor g1344(.dina(n1407),.dinb(n1406),.dout(n1408),.clk(gclk));
	jand g1345(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1409),.clk(gclk));
	jnot g1346(.din(n1409),.dout(n1410),.clk(gclk));
	jand g1347(.dina(w_n1364_0[0]),.dinb(w_n1335_0[0]),.dout(n1411),.clk(gclk));
	jand g1348(.dina(w_n1365_0[0]),.dinb(w_n1332_0[0]),.dout(n1412),.clk(gclk));
	jor g1349(.dina(n1412),.dinb(n1411),.dout(n1413),.clk(gclk));
	jand g1350(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1414),.clk(gclk));
	jnot g1351(.din(n1414),.dout(n1415),.clk(gclk));
	jand g1352(.dina(w_n1362_0[0]),.dinb(w_n1340_0[0]),.dout(n1416),.clk(gclk));
	jand g1353(.dina(w_n1363_0[0]),.dinb(w_n1337_0[0]),.dout(n1417),.clk(gclk));
	jor g1354(.dina(n1417),.dinb(n1416),.dout(n1418),.clk(gclk));
	jand g1355(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1419),.clk(gclk));
	jnot g1356(.din(n1419),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_n1360_0[0]),.dinb(w_n1345_0[0]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1361_0[0]),.dinb(w_n1342_0[0]),.dout(n1422),.clk(gclk));
	jor g1359(.dina(n1422),.dinb(n1421),.dout(n1423),.clk(gclk));
	jand g1360(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1424),.clk(gclk));
	jnot g1361(.din(n1424),.dout(n1425),.clk(gclk));
	jand g1362(.dina(w_n1358_0[0]),.dinb(w_n1350_0[0]),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1359_0[0]),.dinb(w_n1347_0[0]),.dout(n1427),.clk(gclk));
	jor g1364(.dina(n1427),.dinb(n1426),.dout(n1428),.clk(gclk));
	jand g1365(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1429),.clk(gclk));
	jand g1366(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1430),.clk(gclk));
	jor g1367(.dina(w_n1355_0[0]),.dinb(w_n1352_0[0]),.dout(n1431),.clk(gclk));
	jor g1368(.dina(w_n1357_0[0]),.dinb(w_n1351_0[0]),.dout(n1432),.clk(gclk));
	jand g1369(.dina(n1432),.dinb(n1431),.dout(n1433),.clk(gclk));
	jxor g1370(.dina(w_n1433_0[1]),.dinb(w_n1430_0[1]),.dout(n1434),.clk(gclk));
	jnot g1371(.din(n1434),.dout(n1435),.clk(gclk));
	jxor g1372(.dina(w_n1435_0[1]),.dinb(w_n1429_0[1]),.dout(n1436),.clk(gclk));
	jxor g1373(.dina(w_n1436_0[1]),.dinb(w_n1428_0[1]),.dout(n1437),.clk(gclk));
	jxor g1374(.dina(w_n1437_0[1]),.dinb(w_n1425_0[1]),.dout(n1438),.clk(gclk));
	jxor g1375(.dina(w_n1438_0[1]),.dinb(w_n1423_0[1]),.dout(n1439),.clk(gclk));
	jxor g1376(.dina(w_n1439_0[1]),.dinb(w_n1420_0[1]),.dout(n1440),.clk(gclk));
	jxor g1377(.dina(w_n1440_0[1]),.dinb(w_n1418_0[1]),.dout(n1441),.clk(gclk));
	jxor g1378(.dina(w_n1441_0[1]),.dinb(w_n1415_0[1]),.dout(n1442),.clk(gclk));
	jxor g1379(.dina(w_n1442_0[1]),.dinb(w_n1413_0[1]),.dout(n1443),.clk(gclk));
	jxor g1380(.dina(w_n1443_0[1]),.dinb(w_n1410_0[1]),.dout(n1444),.clk(gclk));
	jxor g1381(.dina(w_n1444_0[1]),.dinb(w_n1408_0[1]),.dout(n1445),.clk(gclk));
	jxor g1382(.dina(w_n1445_0[1]),.dinb(w_n1405_0[1]),.dout(n1446),.clk(gclk));
	jxor g1383(.dina(w_n1446_0[1]),.dinb(w_n1403_0[1]),.dout(n1447),.clk(gclk));
	jxor g1384(.dina(w_n1447_0[1]),.dinb(w_n1400_0[1]),.dout(n1448),.clk(gclk));
	jxor g1385(.dina(w_n1448_0[1]),.dinb(w_n1398_0[1]),.dout(n1449),.clk(gclk));
	jxor g1386(.dina(w_n1449_0[1]),.dinb(w_n1395_0[1]),.dout(n1450),.clk(gclk));
	jxor g1387(.dina(w_n1450_0[1]),.dinb(w_n1393_0[1]),.dout(n1451),.clk(gclk));
	jnot g1388(.din(n1451),.dout(n1452),.clk(gclk));
	jxor g1389(.dina(w_n1452_0[1]),.dinb(w_n1390_0[1]),.dout(n1453),.clk(gclk));
	jnot g1390(.din(n1453),.dout(n1454),.clk(gclk));
	jxor g1391(.dina(w_n1454_0[1]),.dinb(w_n1389_0[1]),.dout(n1455),.clk(gclk));
	jxor g1392(.dina(w_n1455_0[1]),.dinb(w_n1384_0[1]),.dout(w_dff_A_X5zW4CkD5_2),.clk(gclk));
	jor g1393(.dina(w_n1454_0[0]),.dinb(w_n1389_0[0]),.dout(n1457),.clk(gclk));
	jnot g1394(.din(w_n1455_0[0]),.dout(n1458),.clk(gclk));
	jor g1395(.dina(w_dff_B_K8aNhHto4_0),.dinb(w_n1384_0[0]),.dout(n1459),.clk(gclk));
	jand g1396(.dina(n1459),.dinb(w_dff_B_S72RrKdf6_1),.dout(n1460),.clk(gclk));
	jnot g1397(.din(w_n1393_0[0]),.dout(n1461),.clk(gclk));
	jnot g1398(.din(w_n1450_0[0]),.dout(n1462),.clk(gclk));
	jor g1399(.dina(n1462),.dinb(n1461),.dout(n1463),.clk(gclk));
	jor g1400(.dina(w_n1452_0[0]),.dinb(w_n1390_0[0]),.dout(n1464),.clk(gclk));
	jand g1401(.dina(n1464),.dinb(n1463),.dout(n1465),.clk(gclk));
	jand g1402(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1466),.clk(gclk));
	jand g1403(.dina(w_n1448_0[0]),.dinb(w_n1398_0[0]),.dout(n1467),.clk(gclk));
	jand g1404(.dina(w_n1449_0[0]),.dinb(w_n1395_0[0]),.dout(n1468),.clk(gclk));
	jor g1405(.dina(n1468),.dinb(n1467),.dout(n1469),.clk(gclk));
	jand g1406(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1470),.clk(gclk));
	jnot g1407(.din(n1470),.dout(n1471),.clk(gclk));
	jand g1408(.dina(w_n1446_0[0]),.dinb(w_n1403_0[0]),.dout(n1472),.clk(gclk));
	jand g1409(.dina(w_n1447_0[0]),.dinb(w_n1400_0[0]),.dout(n1473),.clk(gclk));
	jor g1410(.dina(n1473),.dinb(n1472),.dout(n1474),.clk(gclk));
	jand g1411(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1475),.clk(gclk));
	jnot g1412(.din(n1475),.dout(n1476),.clk(gclk));
	jand g1413(.dina(w_n1444_0[0]),.dinb(w_n1408_0[0]),.dout(n1477),.clk(gclk));
	jand g1414(.dina(w_n1445_0[0]),.dinb(w_n1405_0[0]),.dout(n1478),.clk(gclk));
	jor g1415(.dina(n1478),.dinb(n1477),.dout(n1479),.clk(gclk));
	jand g1416(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1480),.clk(gclk));
	jnot g1417(.din(n1480),.dout(n1481),.clk(gclk));
	jand g1418(.dina(w_n1442_0[0]),.dinb(w_n1413_0[0]),.dout(n1482),.clk(gclk));
	jand g1419(.dina(w_n1443_0[0]),.dinb(w_n1410_0[0]),.dout(n1483),.clk(gclk));
	jor g1420(.dina(n1483),.dinb(n1482),.dout(n1484),.clk(gclk));
	jand g1421(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1485),.clk(gclk));
	jnot g1422(.din(n1485),.dout(n1486),.clk(gclk));
	jand g1423(.dina(w_n1440_0[0]),.dinb(w_n1418_0[0]),.dout(n1487),.clk(gclk));
	jand g1424(.dina(w_n1441_0[0]),.dinb(w_n1415_0[0]),.dout(n1488),.clk(gclk));
	jor g1425(.dina(n1488),.dinb(n1487),.dout(n1489),.clk(gclk));
	jand g1426(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1490),.clk(gclk));
	jnot g1427(.din(n1490),.dout(n1491),.clk(gclk));
	jand g1428(.dina(w_n1438_0[0]),.dinb(w_n1423_0[0]),.dout(n1492),.clk(gclk));
	jand g1429(.dina(w_n1439_0[0]),.dinb(w_n1420_0[0]),.dout(n1493),.clk(gclk));
	jor g1430(.dina(n1493),.dinb(n1492),.dout(n1494),.clk(gclk));
	jand g1431(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1495),.clk(gclk));
	jnot g1432(.din(n1495),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_n1436_0[0]),.dinb(w_n1428_0[0]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1437_0[0]),.dinb(w_n1425_0[0]),.dout(n1498),.clk(gclk));
	jor g1435(.dina(n1498),.dinb(n1497),.dout(n1499),.clk(gclk));
	jand g1436(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1500),.clk(gclk));
	jand g1437(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1501),.clk(gclk));
	jor g1438(.dina(w_n1433_0[0]),.dinb(w_n1430_0[0]),.dout(n1502),.clk(gclk));
	jor g1439(.dina(w_n1435_0[0]),.dinb(w_n1429_0[0]),.dout(n1503),.clk(gclk));
	jand g1440(.dina(n1503),.dinb(n1502),.dout(n1504),.clk(gclk));
	jxor g1441(.dina(w_n1504_0[1]),.dinb(w_n1501_0[1]),.dout(n1505),.clk(gclk));
	jnot g1442(.din(n1505),.dout(n1506),.clk(gclk));
	jxor g1443(.dina(w_n1506_0[1]),.dinb(w_n1500_0[1]),.dout(n1507),.clk(gclk));
	jxor g1444(.dina(w_n1507_0[1]),.dinb(w_n1499_0[1]),.dout(n1508),.clk(gclk));
	jxor g1445(.dina(w_n1508_0[1]),.dinb(w_n1496_0[1]),.dout(n1509),.clk(gclk));
	jxor g1446(.dina(w_n1509_0[1]),.dinb(w_n1494_0[1]),.dout(n1510),.clk(gclk));
	jxor g1447(.dina(w_n1510_0[1]),.dinb(w_n1491_0[1]),.dout(n1511),.clk(gclk));
	jxor g1448(.dina(w_n1511_0[1]),.dinb(w_n1489_0[1]),.dout(n1512),.clk(gclk));
	jxor g1449(.dina(w_n1512_0[1]),.dinb(w_n1486_0[1]),.dout(n1513),.clk(gclk));
	jxor g1450(.dina(w_n1513_0[1]),.dinb(w_n1484_0[1]),.dout(n1514),.clk(gclk));
	jxor g1451(.dina(w_n1514_0[1]),.dinb(w_n1481_0[1]),.dout(n1515),.clk(gclk));
	jxor g1452(.dina(w_n1515_0[1]),.dinb(w_n1479_0[1]),.dout(n1516),.clk(gclk));
	jxor g1453(.dina(w_n1516_0[1]),.dinb(w_n1476_0[1]),.dout(n1517),.clk(gclk));
	jxor g1454(.dina(w_n1517_0[1]),.dinb(w_n1474_0[1]),.dout(n1518),.clk(gclk));
	jxor g1455(.dina(w_n1518_0[1]),.dinb(w_n1471_0[1]),.dout(n1519),.clk(gclk));
	jxor g1456(.dina(w_n1519_0[1]),.dinb(w_n1469_0[1]),.dout(n1520),.clk(gclk));
	jnot g1457(.din(n1520),.dout(n1521),.clk(gclk));
	jxor g1458(.dina(w_n1521_0[1]),.dinb(w_n1466_0[1]),.dout(n1522),.clk(gclk));
	jnot g1459(.din(n1522),.dout(n1523),.clk(gclk));
	jxor g1460(.dina(w_n1523_0[1]),.dinb(w_n1465_0[1]),.dout(n1524),.clk(gclk));
	jxor g1461(.dina(w_n1524_0[1]),.dinb(w_n1460_0[1]),.dout(w_dff_A_FtorKECO3_2),.clk(gclk));
	jor g1462(.dina(w_n1523_0[0]),.dinb(w_n1465_0[0]),.dout(n1526),.clk(gclk));
	jnot g1463(.din(w_n1524_0[0]),.dout(n1527),.clk(gclk));
	jor g1464(.dina(w_dff_B_tPp8Fugc9_0),.dinb(w_n1460_0[0]),.dout(n1528),.clk(gclk));
	jand g1465(.dina(n1528),.dinb(w_dff_B_6XWUy8nb8_1),.dout(n1529),.clk(gclk));
	jnot g1466(.din(w_n1469_0[0]),.dout(n1530),.clk(gclk));
	jnot g1467(.din(w_n1519_0[0]),.dout(n1531),.clk(gclk));
	jor g1468(.dina(n1531),.dinb(n1530),.dout(n1532),.clk(gclk));
	jor g1469(.dina(w_n1521_0[0]),.dinb(w_n1466_0[0]),.dout(n1533),.clk(gclk));
	jand g1470(.dina(n1533),.dinb(n1532),.dout(n1534),.clk(gclk));
	jand g1471(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1535),.clk(gclk));
	jand g1472(.dina(w_n1517_0[0]),.dinb(w_n1474_0[0]),.dout(n1536),.clk(gclk));
	jand g1473(.dina(w_n1518_0[0]),.dinb(w_n1471_0[0]),.dout(n1537),.clk(gclk));
	jor g1474(.dina(n1537),.dinb(n1536),.dout(n1538),.clk(gclk));
	jand g1475(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1539),.clk(gclk));
	jnot g1476(.din(n1539),.dout(n1540),.clk(gclk));
	jand g1477(.dina(w_n1515_0[0]),.dinb(w_n1479_0[0]),.dout(n1541),.clk(gclk));
	jand g1478(.dina(w_n1516_0[0]),.dinb(w_n1476_0[0]),.dout(n1542),.clk(gclk));
	jor g1479(.dina(n1542),.dinb(n1541),.dout(n1543),.clk(gclk));
	jand g1480(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1544),.clk(gclk));
	jnot g1481(.din(n1544),.dout(n1545),.clk(gclk));
	jand g1482(.dina(w_n1513_0[0]),.dinb(w_n1484_0[0]),.dout(n1546),.clk(gclk));
	jand g1483(.dina(w_n1514_0[0]),.dinb(w_n1481_0[0]),.dout(n1547),.clk(gclk));
	jor g1484(.dina(n1547),.dinb(n1546),.dout(n1548),.clk(gclk));
	jand g1485(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1549),.clk(gclk));
	jnot g1486(.din(n1549),.dout(n1550),.clk(gclk));
	jand g1487(.dina(w_n1511_0[0]),.dinb(w_n1489_0[0]),.dout(n1551),.clk(gclk));
	jand g1488(.dina(w_n1512_0[0]),.dinb(w_n1486_0[0]),.dout(n1552),.clk(gclk));
	jor g1489(.dina(n1552),.dinb(n1551),.dout(n1553),.clk(gclk));
	jand g1490(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1554),.clk(gclk));
	jnot g1491(.din(n1554),.dout(n1555),.clk(gclk));
	jand g1492(.dina(w_n1509_0[0]),.dinb(w_n1494_0[0]),.dout(n1556),.clk(gclk));
	jand g1493(.dina(w_n1510_0[0]),.dinb(w_n1491_0[0]),.dout(n1557),.clk(gclk));
	jor g1494(.dina(n1557),.dinb(n1556),.dout(n1558),.clk(gclk));
	jand g1495(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1559),.clk(gclk));
	jnot g1496(.din(n1559),.dout(n1560),.clk(gclk));
	jand g1497(.dina(w_n1507_0[0]),.dinb(w_n1499_0[0]),.dout(n1561),.clk(gclk));
	jand g1498(.dina(w_n1508_0[0]),.dinb(w_n1496_0[0]),.dout(n1562),.clk(gclk));
	jor g1499(.dina(n1562),.dinb(n1561),.dout(n1563),.clk(gclk));
	jand g1500(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1564),.clk(gclk));
	jand g1501(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1565),.clk(gclk));
	jor g1502(.dina(w_n1504_0[0]),.dinb(w_n1501_0[0]),.dout(n1566),.clk(gclk));
	jor g1503(.dina(w_n1506_0[0]),.dinb(w_n1500_0[0]),.dout(n1567),.clk(gclk));
	jand g1504(.dina(n1567),.dinb(n1566),.dout(n1568),.clk(gclk));
	jxor g1505(.dina(w_n1568_0[1]),.dinb(w_n1565_0[1]),.dout(n1569),.clk(gclk));
	jnot g1506(.din(n1569),.dout(n1570),.clk(gclk));
	jxor g1507(.dina(w_n1570_0[1]),.dinb(w_n1564_0[1]),.dout(n1571),.clk(gclk));
	jxor g1508(.dina(w_n1571_0[1]),.dinb(w_n1563_0[1]),.dout(n1572),.clk(gclk));
	jxor g1509(.dina(w_n1572_0[1]),.dinb(w_n1560_0[1]),.dout(n1573),.clk(gclk));
	jxor g1510(.dina(w_n1573_0[1]),.dinb(w_n1558_0[1]),.dout(n1574),.clk(gclk));
	jxor g1511(.dina(w_n1574_0[1]),.dinb(w_n1555_0[1]),.dout(n1575),.clk(gclk));
	jxor g1512(.dina(w_n1575_0[1]),.dinb(w_n1553_0[1]),.dout(n1576),.clk(gclk));
	jxor g1513(.dina(w_n1576_0[1]),.dinb(w_n1550_0[1]),.dout(n1577),.clk(gclk));
	jxor g1514(.dina(w_n1577_0[1]),.dinb(w_n1548_0[1]),.dout(n1578),.clk(gclk));
	jxor g1515(.dina(w_n1578_0[1]),.dinb(w_n1545_0[1]),.dout(n1579),.clk(gclk));
	jxor g1516(.dina(w_n1579_0[1]),.dinb(w_n1543_0[1]),.dout(n1580),.clk(gclk));
	jxor g1517(.dina(w_n1580_0[1]),.dinb(w_n1540_0[1]),.dout(n1581),.clk(gclk));
	jxor g1518(.dina(w_n1581_0[1]),.dinb(w_n1538_0[1]),.dout(n1582),.clk(gclk));
	jnot g1519(.din(n1582),.dout(n1583),.clk(gclk));
	jxor g1520(.dina(w_n1583_0[1]),.dinb(w_n1535_0[1]),.dout(n1584),.clk(gclk));
	jnot g1521(.din(n1584),.dout(n1585),.clk(gclk));
	jxor g1522(.dina(w_n1585_0[1]),.dinb(w_n1534_0[1]),.dout(n1586),.clk(gclk));
	jxor g1523(.dina(w_n1586_0[1]),.dinb(w_n1529_0[1]),.dout(w_dff_A_EvWttnxa3_2),.clk(gclk));
	jor g1524(.dina(w_n1585_0[0]),.dinb(w_n1534_0[0]),.dout(n1588),.clk(gclk));
	jnot g1525(.din(w_n1586_0[0]),.dout(n1589),.clk(gclk));
	jor g1526(.dina(w_dff_B_BRq9R90W5_0),.dinb(w_n1529_0[0]),.dout(n1590),.clk(gclk));
	jand g1527(.dina(n1590),.dinb(w_dff_B_PekFeIzl8_1),.dout(n1591),.clk(gclk));
	jnot g1528(.din(w_n1538_0[0]),.dout(n1592),.clk(gclk));
	jnot g1529(.din(w_n1581_0[0]),.dout(n1593),.clk(gclk));
	jor g1530(.dina(n1593),.dinb(n1592),.dout(n1594),.clk(gclk));
	jor g1531(.dina(w_n1583_0[0]),.dinb(w_n1535_0[0]),.dout(n1595),.clk(gclk));
	jand g1532(.dina(n1595),.dinb(n1594),.dout(n1596),.clk(gclk));
	jand g1533(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1597),.clk(gclk));
	jand g1534(.dina(w_n1579_0[0]),.dinb(w_n1543_0[0]),.dout(n1598),.clk(gclk));
	jand g1535(.dina(w_n1580_0[0]),.dinb(w_n1540_0[0]),.dout(n1599),.clk(gclk));
	jor g1536(.dina(n1599),.dinb(n1598),.dout(n1600),.clk(gclk));
	jand g1537(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1601),.clk(gclk));
	jnot g1538(.din(n1601),.dout(n1602),.clk(gclk));
	jand g1539(.dina(w_n1577_0[0]),.dinb(w_n1548_0[0]),.dout(n1603),.clk(gclk));
	jand g1540(.dina(w_n1578_0[0]),.dinb(w_n1545_0[0]),.dout(n1604),.clk(gclk));
	jor g1541(.dina(n1604),.dinb(n1603),.dout(n1605),.clk(gclk));
	jand g1542(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1606),.clk(gclk));
	jnot g1543(.din(n1606),.dout(n1607),.clk(gclk));
	jand g1544(.dina(w_n1575_0[0]),.dinb(w_n1553_0[0]),.dout(n1608),.clk(gclk));
	jand g1545(.dina(w_n1576_0[0]),.dinb(w_n1550_0[0]),.dout(n1609),.clk(gclk));
	jor g1546(.dina(n1609),.dinb(n1608),.dout(n1610),.clk(gclk));
	jand g1547(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1611),.clk(gclk));
	jnot g1548(.din(n1611),.dout(n1612),.clk(gclk));
	jand g1549(.dina(w_n1573_0[0]),.dinb(w_n1558_0[0]),.dout(n1613),.clk(gclk));
	jand g1550(.dina(w_n1574_0[0]),.dinb(w_n1555_0[0]),.dout(n1614),.clk(gclk));
	jor g1551(.dina(n1614),.dinb(n1613),.dout(n1615),.clk(gclk));
	jand g1552(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1616),.clk(gclk));
	jnot g1553(.din(n1616),.dout(n1617),.clk(gclk));
	jand g1554(.dina(w_n1571_0[0]),.dinb(w_n1563_0[0]),.dout(n1618),.clk(gclk));
	jand g1555(.dina(w_n1572_0[0]),.dinb(w_n1560_0[0]),.dout(n1619),.clk(gclk));
	jor g1556(.dina(n1619),.dinb(n1618),.dout(n1620),.clk(gclk));
	jand g1557(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1621),.clk(gclk));
	jand g1558(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1622),.clk(gclk));
	jor g1559(.dina(w_n1568_0[0]),.dinb(w_n1565_0[0]),.dout(n1623),.clk(gclk));
	jor g1560(.dina(w_n1570_0[0]),.dinb(w_n1564_0[0]),.dout(n1624),.clk(gclk));
	jand g1561(.dina(n1624),.dinb(n1623),.dout(n1625),.clk(gclk));
	jxor g1562(.dina(w_n1625_0[1]),.dinb(w_n1622_0[1]),.dout(n1626),.clk(gclk));
	jnot g1563(.din(n1626),.dout(n1627),.clk(gclk));
	jxor g1564(.dina(w_n1627_0[1]),.dinb(w_n1621_0[1]),.dout(n1628),.clk(gclk));
	jxor g1565(.dina(w_n1628_0[1]),.dinb(w_n1620_0[1]),.dout(n1629),.clk(gclk));
	jxor g1566(.dina(w_n1629_0[1]),.dinb(w_n1617_0[1]),.dout(n1630),.clk(gclk));
	jxor g1567(.dina(w_n1630_0[1]),.dinb(w_n1615_0[1]),.dout(n1631),.clk(gclk));
	jxor g1568(.dina(w_n1631_0[1]),.dinb(w_n1612_0[1]),.dout(n1632),.clk(gclk));
	jxor g1569(.dina(w_n1632_0[1]),.dinb(w_n1610_0[1]),.dout(n1633),.clk(gclk));
	jxor g1570(.dina(w_n1633_0[1]),.dinb(w_n1607_0[1]),.dout(n1634),.clk(gclk));
	jxor g1571(.dina(w_n1634_0[1]),.dinb(w_n1605_0[1]),.dout(n1635),.clk(gclk));
	jxor g1572(.dina(w_n1635_0[1]),.dinb(w_n1602_0[1]),.dout(n1636),.clk(gclk));
	jxor g1573(.dina(w_n1636_0[1]),.dinb(w_n1600_0[1]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jxor g1575(.dina(w_n1638_0[1]),.dinb(w_n1597_0[1]),.dout(n1639),.clk(gclk));
	jnot g1576(.din(n1639),.dout(n1640),.clk(gclk));
	jxor g1577(.dina(w_n1640_0[1]),.dinb(w_n1596_0[1]),.dout(n1641),.clk(gclk));
	jxor g1578(.dina(w_n1641_0[1]),.dinb(w_n1591_0[1]),.dout(w_dff_A_TLmwHIhE1_2),.clk(gclk));
	jor g1579(.dina(w_n1640_0[0]),.dinb(w_n1596_0[0]),.dout(n1643),.clk(gclk));
	jnot g1580(.din(w_n1641_0[0]),.dout(n1644),.clk(gclk));
	jor g1581(.dina(w_dff_B_17qFCh4f9_0),.dinb(w_n1591_0[0]),.dout(n1645),.clk(gclk));
	jand g1582(.dina(n1645),.dinb(w_dff_B_eDg4Wggn8_1),.dout(n1646),.clk(gclk));
	jnot g1583(.din(w_n1600_0[0]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(w_n1636_0[0]),.dout(n1648),.clk(gclk));
	jor g1585(.dina(n1648),.dinb(n1647),.dout(n1649),.clk(gclk));
	jor g1586(.dina(w_n1638_0[0]),.dinb(w_n1597_0[0]),.dout(n1650),.clk(gclk));
	jand g1587(.dina(n1650),.dinb(n1649),.dout(n1651),.clk(gclk));
	jand g1588(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1652),.clk(gclk));
	jnot g1589(.din(n1652),.dout(n1653),.clk(gclk));
	jand g1590(.dina(w_n1634_0[0]),.dinb(w_n1605_0[0]),.dout(n1654),.clk(gclk));
	jand g1591(.dina(w_n1635_0[0]),.dinb(w_n1602_0[0]),.dout(n1655),.clk(gclk));
	jor g1592(.dina(n1655),.dinb(n1654),.dout(n1656),.clk(gclk));
	jand g1593(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jand g1595(.dina(w_n1632_0[0]),.dinb(w_n1610_0[0]),.dout(n1659),.clk(gclk));
	jand g1596(.dina(w_n1633_0[0]),.dinb(w_n1607_0[0]),.dout(n1660),.clk(gclk));
	jor g1597(.dina(n1660),.dinb(n1659),.dout(n1661),.clk(gclk));
	jand g1598(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1662),.clk(gclk));
	jnot g1599(.din(n1662),.dout(n1663),.clk(gclk));
	jand g1600(.dina(w_n1630_0[0]),.dinb(w_n1615_0[0]),.dout(n1664),.clk(gclk));
	jand g1601(.dina(w_n1631_0[0]),.dinb(w_n1612_0[0]),.dout(n1665),.clk(gclk));
	jor g1602(.dina(n1665),.dinb(n1664),.dout(n1666),.clk(gclk));
	jand g1603(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1667),.clk(gclk));
	jnot g1604(.din(n1667),.dout(n1668),.clk(gclk));
	jand g1605(.dina(w_n1628_0[0]),.dinb(w_n1620_0[0]),.dout(n1669),.clk(gclk));
	jand g1606(.dina(w_n1629_0[0]),.dinb(w_n1617_0[0]),.dout(n1670),.clk(gclk));
	jor g1607(.dina(n1670),.dinb(n1669),.dout(n1671),.clk(gclk));
	jand g1608(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1672),.clk(gclk));
	jand g1609(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1673),.clk(gclk));
	jor g1610(.dina(w_n1625_0[0]),.dinb(w_n1622_0[0]),.dout(n1674),.clk(gclk));
	jor g1611(.dina(w_n1627_0[0]),.dinb(w_n1621_0[0]),.dout(n1675),.clk(gclk));
	jand g1612(.dina(n1675),.dinb(n1674),.dout(n1676),.clk(gclk));
	jxor g1613(.dina(w_n1676_0[1]),.dinb(w_n1673_0[1]),.dout(n1677),.clk(gclk));
	jnot g1614(.din(n1677),.dout(n1678),.clk(gclk));
	jxor g1615(.dina(w_n1678_0[1]),.dinb(w_n1672_0[1]),.dout(n1679),.clk(gclk));
	jxor g1616(.dina(w_n1679_0[1]),.dinb(w_n1671_0[1]),.dout(n1680),.clk(gclk));
	jxor g1617(.dina(w_n1680_0[1]),.dinb(w_n1668_0[1]),.dout(n1681),.clk(gclk));
	jxor g1618(.dina(w_n1681_0[1]),.dinb(w_n1666_0[1]),.dout(n1682),.clk(gclk));
	jxor g1619(.dina(w_n1682_0[1]),.dinb(w_n1663_0[1]),.dout(n1683),.clk(gclk));
	jxor g1620(.dina(w_n1683_0[1]),.dinb(w_n1661_0[1]),.dout(n1684),.clk(gclk));
	jxor g1621(.dina(w_n1684_0[1]),.dinb(w_n1658_0[1]),.dout(n1685),.clk(gclk));
	jxor g1622(.dina(w_n1685_0[1]),.dinb(w_n1656_0[1]),.dout(n1686),.clk(gclk));
	jxor g1623(.dina(w_n1686_0[1]),.dinb(w_n1653_0[1]),.dout(n1687),.clk(gclk));
	jnot g1624(.din(n1687),.dout(n1688),.clk(gclk));
	jxor g1625(.dina(w_n1688_0[1]),.dinb(w_n1651_0[1]),.dout(n1689),.clk(gclk));
	jxor g1626(.dina(w_n1689_0[1]),.dinb(w_n1646_0[1]),.dout(w_dff_A_np4nDYGT0_2),.clk(gclk));
	jor g1627(.dina(w_n1688_0[0]),.dinb(w_n1651_0[0]),.dout(n1691),.clk(gclk));
	jnot g1628(.din(w_n1689_0[0]),.dout(n1692),.clk(gclk));
	jor g1629(.dina(w_dff_B_XtoT0os52_0),.dinb(w_n1646_0[0]),.dout(n1693),.clk(gclk));
	jand g1630(.dina(n1693),.dinb(w_dff_B_FLzv5IFQ9_1),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1685_0[0]),.dinb(w_n1656_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1686_0[0]),.dinb(w_n1653_0[0]),.dout(n1696),.clk(gclk));
	jor g1633(.dina(n1696),.dinb(n1695),.dout(n1697),.clk(gclk));
	jand g1634(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1683_0[0]),.dinb(w_n1661_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1684_0[0]),.dinb(w_n1658_0[0]),.dout(n1701),.clk(gclk));
	jor g1638(.dina(n1701),.dinb(n1700),.dout(n1702),.clk(gclk));
	jand g1639(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1703),.clk(gclk));
	jnot g1640(.din(n1703),.dout(n1704),.clk(gclk));
	jand g1641(.dina(w_n1681_0[0]),.dinb(w_n1666_0[0]),.dout(n1705),.clk(gclk));
	jand g1642(.dina(w_n1682_0[0]),.dinb(w_n1663_0[0]),.dout(n1706),.clk(gclk));
	jor g1643(.dina(n1706),.dinb(n1705),.dout(n1707),.clk(gclk));
	jand g1644(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jand g1646(.dina(w_n1679_0[0]),.dinb(w_n1671_0[0]),.dout(n1710),.clk(gclk));
	jand g1647(.dina(w_n1680_0[0]),.dinb(w_n1668_0[0]),.dout(n1711),.clk(gclk));
	jor g1648(.dina(n1711),.dinb(n1710),.dout(n1712),.clk(gclk));
	jand g1649(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1713),.clk(gclk));
	jand g1650(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1714),.clk(gclk));
	jor g1651(.dina(w_n1676_0[0]),.dinb(w_n1673_0[0]),.dout(n1715),.clk(gclk));
	jor g1652(.dina(w_n1678_0[0]),.dinb(w_n1672_0[0]),.dout(n1716),.clk(gclk));
	jand g1653(.dina(n1716),.dinb(n1715),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1714_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1713_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1712_0[1]),.dout(n1721),.clk(gclk));
	jxor g1658(.dina(w_n1721_0[1]),.dinb(w_n1709_0[1]),.dout(n1722),.clk(gclk));
	jxor g1659(.dina(w_n1722_0[1]),.dinb(w_n1707_0[1]),.dout(n1723),.clk(gclk));
	jxor g1660(.dina(w_n1723_0[1]),.dinb(w_n1704_0[1]),.dout(n1724),.clk(gclk));
	jxor g1661(.dina(w_n1724_0[1]),.dinb(w_n1702_0[1]),.dout(n1725),.clk(gclk));
	jxor g1662(.dina(w_n1725_0[1]),.dinb(w_n1699_0[1]),.dout(n1726),.clk(gclk));
	jxor g1663(.dina(w_n1726_0[1]),.dinb(w_n1697_0[1]),.dout(n1727),.clk(gclk));
	jxor g1664(.dina(w_n1727_0[1]),.dinb(w_n1694_0[1]),.dout(w_dff_A_MxA6KRqk3_2),.clk(gclk));
	jnot g1665(.din(w_n1697_0[0]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(w_n1726_0[0]),.dout(n1730),.clk(gclk));
	jor g1667(.dina(n1730),.dinb(n1729),.dout(n1731),.clk(gclk));
	jnot g1668(.din(w_n1727_0[0]),.dout(n1732),.clk(gclk));
	jor g1669(.dina(w_dff_B_H4gx2No93_0),.dinb(w_n1694_0[0]),.dout(n1733),.clk(gclk));
	jand g1670(.dina(n1733),.dinb(w_dff_B_IZ4uEvw22_1),.dout(n1734),.clk(gclk));
	jand g1671(.dina(w_n1724_0[0]),.dinb(w_n1702_0[0]),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1725_0[0]),.dinb(w_n1699_0[0]),.dout(n1736),.clk(gclk));
	jor g1673(.dina(n1736),.dinb(n1735),.dout(n1737),.clk(gclk));
	jand g1674(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1738),.clk(gclk));
	jnot g1675(.din(n1738),.dout(n1739),.clk(gclk));
	jand g1676(.dina(w_n1722_0[0]),.dinb(w_n1707_0[0]),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1723_0[0]),.dinb(w_n1704_0[0]),.dout(n1741),.clk(gclk));
	jor g1678(.dina(n1741),.dinb(n1740),.dout(n1742),.clk(gclk));
	jand g1679(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1743),.clk(gclk));
	jnot g1680(.din(n1743),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_n1720_0[0]),.dinb(w_n1712_0[0]),.dout(n1745),.clk(gclk));
	jand g1682(.dina(w_n1721_0[0]),.dinb(w_n1709_0[0]),.dout(n1746),.clk(gclk));
	jor g1683(.dina(n1746),.dinb(n1745),.dout(n1747),.clk(gclk));
	jand g1684(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1748),.clk(gclk));
	jand g1685(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1749),.clk(gclk));
	jor g1686(.dina(w_n1717_0[0]),.dinb(w_n1714_0[0]),.dout(n1750),.clk(gclk));
	jor g1687(.dina(w_n1719_0[0]),.dinb(w_n1713_0[0]),.dout(n1751),.clk(gclk));
	jand g1688(.dina(n1751),.dinb(n1750),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1749_0[1]),.dout(n1753),.clk(gclk));
	jnot g1690(.din(n1753),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1748_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1747_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1744_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1742_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1739_0[1]),.dout(n1759),.clk(gclk));
	jxor g1696(.dina(w_n1759_0[1]),.dinb(w_n1737_0[1]),.dout(n1760),.clk(gclk));
	jxor g1697(.dina(w_n1760_0[1]),.dinb(w_n1734_0[1]),.dout(w_dff_A_vaZ8kvun7_2),.clk(gclk));
	jnot g1698(.din(w_n1737_0[0]),.dout(n1762),.clk(gclk));
	jnot g1699(.din(w_n1759_0[0]),.dout(n1763),.clk(gclk));
	jor g1700(.dina(n1763),.dinb(n1762),.dout(n1764),.clk(gclk));
	jnot g1701(.din(w_n1760_0[0]),.dout(n1765),.clk(gclk));
	jor g1702(.dina(w_dff_B_mlOdPv2S6_0),.dinb(w_n1734_0[0]),.dout(n1766),.clk(gclk));
	jand g1703(.dina(n1766),.dinb(w_dff_B_cJe6CABx7_1),.dout(n1767),.clk(gclk));
	jand g1704(.dina(w_n1757_0[0]),.dinb(w_n1742_0[0]),.dout(n1768),.clk(gclk));
	jand g1705(.dina(w_n1758_0[0]),.dinb(w_n1739_0[0]),.dout(n1769),.clk(gclk));
	jor g1706(.dina(n1769),.dinb(n1768),.dout(n1770),.clk(gclk));
	jand g1707(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1771),.clk(gclk));
	jnot g1708(.din(n1771),.dout(n1772),.clk(gclk));
	jand g1709(.dina(w_n1755_0[0]),.dinb(w_n1747_0[0]),.dout(n1773),.clk(gclk));
	jand g1710(.dina(w_n1756_0[0]),.dinb(w_n1744_0[0]),.dout(n1774),.clk(gclk));
	jor g1711(.dina(n1774),.dinb(n1773),.dout(n1775),.clk(gclk));
	jand g1712(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1777),.clk(gclk));
	jor g1714(.dina(w_n1752_0[0]),.dinb(w_n1749_0[0]),.dout(n1778),.clk(gclk));
	jor g1715(.dina(w_n1754_0[0]),.dinb(w_n1748_0[0]),.dout(n1779),.clk(gclk));
	jand g1716(.dina(n1779),.dinb(n1778),.dout(n1780),.clk(gclk));
	jxor g1717(.dina(w_n1780_0[1]),.dinb(w_n1777_0[1]),.dout(n1781),.clk(gclk));
	jnot g1718(.din(n1781),.dout(n1782),.clk(gclk));
	jxor g1719(.dina(w_n1782_0[1]),.dinb(w_n1776_0[1]),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1775_0[1]),.dout(n1784),.clk(gclk));
	jxor g1721(.dina(w_n1784_0[1]),.dinb(w_n1772_0[1]),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1770_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1767_0[1]),.dout(w_dff_A_QTxU36lP3_2),.clk(gclk));
	jnot g1724(.din(w_n1770_0[0]),.dout(n1788),.clk(gclk));
	jnot g1725(.din(w_n1785_0[0]),.dout(n1789),.clk(gclk));
	jor g1726(.dina(n1789),.dinb(n1788),.dout(n1790),.clk(gclk));
	jnot g1727(.din(w_n1786_0[0]),.dout(n1791),.clk(gclk));
	jor g1728(.dina(w_dff_B_zeHvFZoO8_0),.dinb(w_n1767_0[0]),.dout(n1792),.clk(gclk));
	jand g1729(.dina(n1792),.dinb(w_dff_B_rfh8Azrx4_1),.dout(n1793),.clk(gclk));
	jand g1730(.dina(w_n1783_0[0]),.dinb(w_n1775_0[0]),.dout(n1794),.clk(gclk));
	jand g1731(.dina(w_n1784_0[0]),.dinb(w_n1772_0[0]),.dout(n1795),.clk(gclk));
	jor g1732(.dina(n1795),.dinb(n1794),.dout(n1796),.clk(gclk));
	jand g1733(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1797),.clk(gclk));
	jand g1734(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1798),.clk(gclk));
	jor g1735(.dina(w_n1780_0[0]),.dinb(w_n1777_0[0]),.dout(n1799),.clk(gclk));
	jor g1736(.dina(w_n1782_0[0]),.dinb(w_n1776_0[0]),.dout(n1800),.clk(gclk));
	jand g1737(.dina(n1800),.dinb(n1799),.dout(n1801),.clk(gclk));
	jxor g1738(.dina(w_n1801_0[1]),.dinb(w_n1798_0[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jxor g1740(.dina(w_n1803_0[1]),.dinb(w_n1797_0[1]),.dout(n1804),.clk(gclk));
	jxor g1741(.dina(w_n1804_0[1]),.dinb(w_n1796_0[1]),.dout(n1805),.clk(gclk));
	jxor g1742(.dina(w_n1805_0[1]),.dinb(w_n1793_0[1]),.dout(w_dff_A_emw7PjXC7_2),.clk(gclk));
	jand g1743(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1807),.clk(gclk));
	jor g1744(.dina(w_n1801_0[0]),.dinb(w_n1798_0[0]),.dout(n1808),.clk(gclk));
	jor g1745(.dina(w_n1803_0[0]),.dinb(w_n1797_0[0]),.dout(n1809),.clk(gclk));
	jand g1746(.dina(n1809),.dinb(n1808),.dout(n1810),.clk(gclk));
	jor g1747(.dina(w_n1810_0[1]),.dinb(w_n1807_0[1]),.dout(n1811),.clk(gclk));
	jnot g1748(.din(w_n1796_0[0]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(w_n1804_0[0]),.dout(n1813),.clk(gclk));
	jor g1750(.dina(n1813),.dinb(n1812),.dout(n1814),.clk(gclk));
	jnot g1751(.din(w_n1805_0[0]),.dout(n1815),.clk(gclk));
	jor g1752(.dina(w_dff_B_MdmJGBM98_0),.dinb(w_n1793_0[0]),.dout(n1816),.clk(gclk));
	jand g1753(.dina(n1816),.dinb(w_dff_B_5v4CRyGD2_1),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1810_0[0]),.dinb(w_n1807_0[0]),.dout(n1818),.clk(gclk));
	jnot g1755(.din(w_n1818_0[1]),.dout(n1819),.clk(gclk));
	jor g1756(.dina(w_dff_B_7IAlXGz98_0),.dinb(w_n1817_0[1]),.dout(n1820),.clk(gclk));
	jand g1757(.dina(n1820),.dinb(w_dff_B_I6ALDGFU2_1),.dout(G6287gat),.clk(gclk));
	jxor g1758(.dina(w_n1818_0[0]),.dinb(w_n1817_0[0]),.dout(w_dff_A_roQXFJyg9_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl jspl_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl jspl_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_G307gat_2[1]),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl jspl_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(w_dff_A_vQBAJatK4_1),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n66_0(.douta(w_dff_A_19rWTS8w4_0),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(w_dff_B_0KNpzkH01_2));
	jspl jspl_w_n69_0(.douta(w_n69_0[0]),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.doutc(w_n80_0[2]),.din(n80));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.din(n91));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.din(n103));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n106_0(.douta(w_n106_0[0]),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl jspl_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.din(n122));
	jspl jspl_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n129_0(.douta(w_n129_0[0]),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.din(n130));
	jspl jspl_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.din(n132));
	jspl jspl_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.din(n133));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.din(n135));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.doutc(w_n146_0[2]),.din(n146));
	jspl jspl_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.din(n148));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(n154));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(n158));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl jspl_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(n165));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl jspl_w_n183_0(.douta(w_n183_0[0]),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.din(n192));
	jspl jspl_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.din(n194));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.doutc(w_n196_0[2]),.din(n196));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(n203));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.din(n209));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.doutc(w_n223_0[2]),.din(n223));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(n225));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.din(n230));
	jspl jspl_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.din(n233));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_n235_0[1]),.din(n235));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(n239));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(n241));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n248_0(.douta(w_n248_0[0]),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.din(n251));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.din(n253));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n256_0(.douta(w_n256_0[0]),.doutb(w_n256_0[1]),.din(n256));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(n267));
	jspl3 jspl3_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.doutc(w_n272_0[2]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(n279));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n284_0(.douta(w_n284_0[0]),.doutb(w_n284_0[1]),.din(n284));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl jspl_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.din(n289));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(n295));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl3 jspl3_w_n297_0(.douta(w_n297_0[0]),.doutb(w_n297_0[1]),.doutc(w_n297_0[2]),.din(n297));
	jspl jspl_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.din(n299));
	jspl jspl_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.din(n301));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_n302_0[1]),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.din(n304));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(n305));
	jspl jspl_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.din(n306));
	jspl jspl_w_n307_0(.douta(w_n307_0[0]),.doutb(w_n307_0[1]),.din(n307));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(n309));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(n310));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.din(n312));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.din(n317));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(n323));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(n330));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.din(n335));
	jspl jspl_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.din(n338));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl jspl_w_n343_0(.douta(w_n343_0[0]),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(n345));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.din(n354));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(n356));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl3 jspl3_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.doutc(w_n358_0[2]),.din(n358));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(n363));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(n366));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(n368));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(n370));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.din(n374));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.din(n377));
	jspl jspl_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.din(n378));
	jspl jspl_w_n380_0(.douta(w_n380_0[0]),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.doutc(w_n391_0[2]),.din(n391));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.din(n396));
	jspl jspl_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.din(n398));
	jspl jspl_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.din(n401));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl jspl_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.din(n406));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl jspl_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.din(n411));
	jspl jspl_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.din(n413));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(n416));
	jspl jspl_w_n418_0(.douta(w_n418_0[0]),.doutb(w_n418_0[1]),.din(n418));
	jspl jspl_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.din(n423));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl3 jspl3_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.doutc(w_n427_0[2]),.din(n427));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl jspl_w_n431_0(.douta(w_n431_0[0]),.doutb(w_n431_0[1]),.din(n431));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(n432));
	jspl jspl_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.din(n433));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl jspl_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.din(n436));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl jspl_w_n438_0(.douta(w_n438_0[0]),.doutb(w_n438_0[1]),.din(n438));
	jspl jspl_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.din(n439));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_n442_0[1]),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n444_0(.douta(w_n444_0[0]),.doutb(w_n444_0[1]),.din(n444));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.din(n448));
	jspl jspl_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.din(n449));
	jspl jspl_w_n451_0(.douta(w_n451_0[0]),.doutb(w_n451_0[1]),.din(n451));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(n464));
	jspl jspl_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.din(n467));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(n469));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(n474));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(n479));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(n489));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(n499));
	jspl jspl_w_n501_0(.douta(w_n501_0[0]),.doutb(w_n501_0[1]),.din(n501));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl3 jspl3_w_n503_0(.douta(w_n503_0[0]),.doutb(w_n503_0[1]),.doutc(w_n503_0[2]),.din(n503));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(n509));
	jspl jspl_w_n510_0(.douta(w_n510_0[0]),.doutb(w_n510_0[1]),.din(n510));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.din(n513));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n515_0(.douta(w_n515_0[0]),.doutb(w_n515_0[1]),.din(n515));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(n519));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n521_0(.douta(w_n521_0[0]),.doutb(w_n521_0[1]),.din(n521));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl jspl_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n526_0(.douta(w_n526_0[0]),.doutb(w_n526_0[1]),.din(n526));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_n529_0[0]),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.din(n535));
	jspl3 jspl3_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.doutc(w_n540_0[2]),.din(n540));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(n547));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(n552));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(n567));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl jspl_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.din(n572));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(n577));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(n588));
	jspl jspl_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.din(n590));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(n592));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl jspl_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.din(n594));
	jspl jspl_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.din(n595));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(n596));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl jspl_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.din(n599));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(n600));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(n606));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.din(n609));
	jspl jspl_w_n611_0(.douta(w_n611_0[0]),.doutb(w_n611_0[1]),.din(n611));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl jspl_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.din(n614));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.din(n620));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl jspl_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.din(n635));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(n637));
	jspl jspl_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.din(n640));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(n647));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.din(n660));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(n662));
	jspl jspl_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.din(n665));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(n667));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(n674));
	jspl jspl_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.din(n675));
	jspl3 jspl3_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.doutc(w_n676_0[2]),.din(n676));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl jspl_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.din(n681));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n688_0(.douta(w_n688_0[0]),.doutb(w_n688_0[1]),.din(n688));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.din(n691));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.din(n692));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.din(n694));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.din(n696));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(n698));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_n700_0[1]),.din(n700));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.din(n712));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.doutc(w_n717_0[2]),.din(n717));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(n719));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(n724));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.din(n729));
	jspl jspl_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.din(n732));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(n734));
	jspl jspl_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.din(n737));
	jspl jspl_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.din(n739));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl jspl_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.din(n744));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(n747));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(n749));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(n762));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(n764));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.din(n774));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.din(n779));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.din(n781));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.din(n783));
	jspl jspl_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.din(n784));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(n787));
	jspl jspl_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.din(n788));
	jspl jspl_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.din(n789));
	jspl jspl_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.din(n790));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl jspl_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.din(n793));
	jspl jspl_w_n794_0(.douta(w_n794_0[0]),.doutb(w_n794_0[1]),.din(n794));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl jspl_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.din(n797));
	jspl jspl_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.din(n798));
	jspl jspl_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.din(n799));
	jspl jspl_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(n803));
	jspl jspl_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(n811));
	jspl jspl_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl3 jspl3_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.doutc(w_n820_0[2]),.din(n820));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(n822));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n830_0(.douta(w_n830_0[0]),.doutb(w_n830_0[1]),.din(n830));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl jspl_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.din(n837));
	jspl jspl_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.din(n840));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(n842));
	jspl jspl_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.din(n845));
	jspl jspl_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.din(n847));
	jspl jspl_w_n850_0(.douta(w_n850_0[0]),.doutb(w_n850_0[1]),.din(n850));
	jspl jspl_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.din(n852));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(n857));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(n862));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n872_0(.douta(w_n872_0[0]),.doutb(w_n872_0[1]),.din(n872));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(n874));
	jspl jspl_w_n875_0(.douta(w_n875_0[0]),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.din(n877));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.din(n880));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n882_0(.douta(w_n882_0[0]),.doutb(w_n882_0[1]),.din(n882));
	jspl jspl_w_n883_0(.douta(w_n883_0[0]),.doutb(w_n883_0[1]),.din(n883));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(n886));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.din(n887));
	jspl jspl_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.din(n888));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(n890));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(n891));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n893_0(.douta(w_n893_0[0]),.doutb(w_n893_0[1]),.din(n893));
	jspl jspl_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(n896));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(n898));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.din(n899));
	jspl3 jspl3_w_n900_0(.douta(w_n900_0[0]),.doutb(w_n900_0[1]),.doutc(w_n900_0[2]),.din(n900));
	jspl jspl_w_n902_0(.douta(w_n902_0[0]),.doutb(w_n902_0[1]),.din(n902));
	jspl jspl_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n904_0(.douta(w_n904_0[0]),.doutb(w_n904_0[1]),.din(n904));
	jspl jspl_w_n905_0(.douta(w_n905_0[0]),.doutb(w_n905_0[1]),.din(n905));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(n910));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(n911));
	jspl3 jspl3_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.doutc(w_n915_0[2]),.din(n915));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(n916));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(n924));
	jspl jspl_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(n929));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n934_0(.douta(w_n934_0[0]),.doutb(w_n934_0[1]),.din(n934));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n939_0(.douta(w_n939_0[0]),.doutb(w_n939_0[1]),.din(n939));
	jspl jspl_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.din(n942));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(n944));
	jspl jspl_w_n947_0(.douta(w_n947_0[0]),.doutb(w_n947_0[1]),.din(n947));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(n949));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(n959));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n967_0(.douta(w_n967_0[0]),.doutb(w_n967_0[1]),.din(n967));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n978_0(.douta(w_n978_0[0]),.doutb(w_n978_0[1]),.din(n978));
	jspl jspl_w_n980_0(.douta(w_n980_0[0]),.doutb(w_n980_0[1]),.din(n980));
	jspl jspl_w_n982_0(.douta(w_n982_0[0]),.doutb(w_n982_0[1]),.din(n982));
	jspl jspl_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.din(n983));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl jspl_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.din(n988));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.din(n990));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl jspl_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.din(n995));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(n996));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl jspl_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.din(n1002));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.din(n1004));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.din(n1006));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(w_dff_B_eoyEvq7x2_2));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_dff_A_ldyRm5Sp4_1),.din(n1013));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(n1018));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(n1023));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(n1028));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1036_0(.douta(w_n1036_0[0]),.doutb(w_n1036_0[1]),.din(n1036));
	jspl jspl_w_n1038_0(.douta(w_n1038_0[0]),.doutb(w_n1038_0[1]),.din(n1038));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(n1043));
	jspl jspl_w_n1046_0(.douta(w_n1046_0[0]),.doutb(w_n1046_0[1]),.din(n1046));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(n1048));
	jspl jspl_w_n1051_0(.douta(w_n1051_0[0]),.doutb(w_n1051_0[1]),.din(n1051));
	jspl jspl_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.din(n1053));
	jspl jspl_w_n1056_0(.douta(w_n1056_0[0]),.doutb(w_n1056_0[1]),.din(n1056));
	jspl jspl_w_n1058_0(.douta(w_n1058_0[0]),.doutb(w_n1058_0[1]),.din(n1058));
	jspl jspl_w_n1061_0(.douta(w_n1061_0[0]),.doutb(w_n1061_0[1]),.din(n1061));
	jspl jspl_w_n1063_0(.douta(w_n1063_0[0]),.doutb(w_n1063_0[1]),.din(n1063));
	jspl jspl_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.din(n1066));
	jspl jspl_w_n1068_0(.douta(w_n1068_0[0]),.doutb(w_n1068_0[1]),.din(n1068));
	jspl jspl_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.din(n1071));
	jspl jspl_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.din(n1073));
	jspl jspl_w_n1076_0(.douta(w_n1076_0[0]),.doutb(w_n1076_0[1]),.din(n1076));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(n1077));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(n1078));
	jspl jspl_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.din(n1080));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl jspl_w_n1083_0(.douta(w_n1083_0[0]),.doutb(w_n1083_0[1]),.din(n1083));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(n1084));
	jspl jspl_w_n1085_0(.douta(w_n1085_0[0]),.doutb(w_n1085_0[1]),.din(n1085));
	jspl jspl_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.din(n1086));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(n1087));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(n1089));
	jspl jspl_w_n1090_0(.douta(w_n1090_0[0]),.doutb(w_n1090_0[1]),.din(n1090));
	jspl jspl_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.din(n1091));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1093_0(.douta(w_n1093_0[0]),.doutb(w_n1093_0[1]),.din(n1093));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(n1094));
	jspl jspl_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.din(n1095));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1098_0(.douta(w_n1098_0[0]),.doutb(w_n1098_0[1]),.din(n1098));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1100_0(.douta(w_n1100_0[0]),.doutb(w_n1100_0[1]),.din(n1100));
	jspl jspl_w_n1101_0(.douta(w_n1101_0[0]),.doutb(w_n1101_0[1]),.din(n1101));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(n1103));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.din(n1105));
	jspl jspl_w_n1106_0(.douta(w_n1106_0[0]),.doutb(w_n1106_0[1]),.din(n1106));
	jspl jspl_w_n1107_0(.douta(w_n1107_0[0]),.doutb(w_n1107_0[1]),.din(n1107));
	jspl jspl_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_n1108_0[1]),.din(n1108));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(n1119));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(n1126));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(n1131));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1136_0(.douta(w_n1136_0[0]),.doutb(w_n1136_0[1]),.din(n1136));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(n1141));
	jspl jspl_w_n1144_0(.douta(w_n1144_0[0]),.doutb(w_n1144_0[1]),.din(n1144));
	jspl jspl_w_n1146_0(.douta(w_n1146_0[0]),.doutb(w_n1146_0[1]),.din(n1146));
	jspl jspl_w_n1149_0(.douta(w_n1149_0[0]),.doutb(w_n1149_0[1]),.din(n1149));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(n1151));
	jspl jspl_w_n1154_0(.douta(w_n1154_0[0]),.doutb(w_n1154_0[1]),.din(n1154));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(n1156));
	jspl jspl_w_n1159_0(.douta(w_n1159_0[0]),.doutb(w_n1159_0[1]),.din(n1159));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(n1161));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(n1164));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl jspl_w_n1169_0(.douta(w_n1169_0[0]),.doutb(w_n1169_0[1]),.din(n1169));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(n1171));
	jspl jspl_w_n1174_0(.douta(w_n1174_0[0]),.doutb(w_n1174_0[1]),.din(n1174));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_n1175_0[1]),.din(n1175));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(n1176));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1182_0(.douta(w_n1182_0[0]),.doutb(w_n1182_0[1]),.din(n1182));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.din(n1184));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(n1186));
	jspl jspl_w_n1187_0(.douta(w_n1187_0[0]),.doutb(w_n1187_0[1]),.din(n1187));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(n1188));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1190_0(.douta(w_n1190_0[0]),.doutb(w_n1190_0[1]),.din(n1190));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(n1191));
	jspl jspl_w_n1192_0(.douta(w_n1192_0[0]),.doutb(w_n1192_0[1]),.din(n1192));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(n1193));
	jspl jspl_w_n1194_0(.douta(w_n1194_0[0]),.doutb(w_n1194_0[1]),.din(n1194));
	jspl jspl_w_n1195_0(.douta(w_n1195_0[0]),.doutb(w_n1195_0[1]),.din(n1195));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.din(n1197));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(n1198));
	jspl jspl_w_n1199_0(.douta(w_n1199_0[0]),.doutb(w_n1199_0[1]),.din(n1199));
	jspl jspl_w_n1200_0(.douta(w_n1200_0[0]),.doutb(w_n1200_0[1]),.din(n1200));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(n1203));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(n1206));
	jspl jspl_w_n1207_0(.douta(w_n1207_0[0]),.doutb(w_n1207_0[1]),.din(n1207));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(n1217));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(n1222));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(n1225));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(n1227));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(n1232));
	jspl jspl_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.din(n1235));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(n1237));
	jspl jspl_w_n1240_0(.douta(w_n1240_0[0]),.doutb(w_n1240_0[1]),.din(n1240));
	jspl jspl_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.din(n1242));
	jspl jspl_w_n1245_0(.douta(w_n1245_0[0]),.doutb(w_n1245_0[1]),.din(n1245));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(n1247));
	jspl jspl_w_n1250_0(.douta(w_n1250_0[0]),.doutb(w_n1250_0[1]),.din(n1250));
	jspl jspl_w_n1252_0(.douta(w_n1252_0[0]),.doutb(w_n1252_0[1]),.din(n1252));
	jspl jspl_w_n1255_0(.douta(w_n1255_0[0]),.doutb(w_n1255_0[1]),.din(n1255));
	jspl jspl_w_n1257_0(.douta(w_n1257_0[0]),.doutb(w_n1257_0[1]),.din(n1257));
	jspl jspl_w_n1260_0(.douta(w_n1260_0[0]),.doutb(w_n1260_0[1]),.din(n1260));
	jspl jspl_w_n1262_0(.douta(w_n1262_0[0]),.doutb(w_n1262_0[1]),.din(n1262));
	jspl jspl_w_n1265_0(.douta(w_n1265_0[0]),.doutb(w_n1265_0[1]),.din(n1265));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(n1266));
	jspl jspl_w_n1267_0(.douta(w_n1267_0[0]),.doutb(w_n1267_0[1]),.din(n1267));
	jspl jspl_w_n1270_0(.douta(w_n1270_0[0]),.doutb(w_n1270_0[1]),.din(n1270));
	jspl jspl_w_n1272_0(.douta(w_n1272_0[0]),.doutb(w_n1272_0[1]),.din(n1272));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(n1273));
	jspl jspl_w_n1274_0(.douta(w_n1274_0[0]),.doutb(w_n1274_0[1]),.din(n1274));
	jspl jspl_w_n1275_0(.douta(w_n1275_0[0]),.doutb(w_n1275_0[1]),.din(n1275));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(n1276));
	jspl jspl_w_n1277_0(.douta(w_n1277_0[0]),.doutb(w_n1277_0[1]),.din(n1277));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(n1278));
	jspl jspl_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.din(n1279));
	jspl jspl_w_n1280_0(.douta(w_n1280_0[0]),.doutb(w_n1280_0[1]),.din(n1280));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(n1281));
	jspl jspl_w_n1282_0(.douta(w_n1282_0[0]),.doutb(w_n1282_0[1]),.din(n1282));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(n1283));
	jspl jspl_w_n1284_0(.douta(w_n1284_0[0]),.doutb(w_n1284_0[1]),.din(n1284));
	jspl jspl_w_n1285_0(.douta(w_n1285_0[0]),.doutb(w_n1285_0[1]),.din(n1285));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(n1286));
	jspl jspl_w_n1287_0(.douta(w_n1287_0[0]),.doutb(w_n1287_0[1]),.din(n1287));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(n1288));
	jspl jspl_w_n1289_0(.douta(w_n1289_0[0]),.doutb(w_n1289_0[1]),.din(n1289));
	jspl jspl_w_n1290_0(.douta(w_n1290_0[0]),.doutb(w_n1290_0[1]),.din(n1290));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_n1291_0[1]),.din(n1291));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(n1293));
	jspl jspl_w_n1294_0(.douta(w_n1294_0[0]),.doutb(w_n1294_0[1]),.din(n1294));
	jspl jspl_w_n1295_0(.douta(w_n1295_0[0]),.doutb(w_n1295_0[1]),.din(n1295));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(n1307));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(n1312));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.din(n1322));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl jspl_w_n1327_0(.douta(w_n1327_0[0]),.doutb(w_n1327_0[1]),.din(n1327));
	jspl jspl_w_n1330_0(.douta(w_n1330_0[0]),.doutb(w_n1330_0[1]),.din(n1330));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(n1332));
	jspl jspl_w_n1335_0(.douta(w_n1335_0[0]),.doutb(w_n1335_0[1]),.din(n1335));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(n1337));
	jspl jspl_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_n1340_0[1]),.din(n1340));
	jspl jspl_w_n1342_0(.douta(w_n1342_0[0]),.doutb(w_n1342_0[1]),.din(n1342));
	jspl jspl_w_n1345_0(.douta(w_n1345_0[0]),.doutb(w_n1345_0[1]),.din(n1345));
	jspl jspl_w_n1347_0(.douta(w_n1347_0[0]),.doutb(w_n1347_0[1]),.din(n1347));
	jspl jspl_w_n1350_0(.douta(w_n1350_0[0]),.doutb(w_n1350_0[1]),.din(n1350));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(n1351));
	jspl jspl_w_n1352_0(.douta(w_n1352_0[0]),.doutb(w_n1352_0[1]),.din(n1352));
	jspl jspl_w_n1355_0(.douta(w_n1355_0[0]),.doutb(w_n1355_0[1]),.din(n1355));
	jspl jspl_w_n1357_0(.douta(w_n1357_0[0]),.doutb(w_n1357_0[1]),.din(n1357));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.din(n1359));
	jspl jspl_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.din(n1360));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1362_0(.douta(w_n1362_0[0]),.doutb(w_n1362_0[1]),.din(n1362));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(n1363));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_n1364_0[1]),.din(n1364));
	jspl jspl_w_n1365_0(.douta(w_n1365_0[0]),.doutb(w_n1365_0[1]),.din(n1365));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(n1366));
	jspl jspl_w_n1367_0(.douta(w_n1367_0[0]),.doutb(w_n1367_0[1]),.din(n1367));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(n1368));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(n1369));
	jspl jspl_w_n1370_0(.douta(w_n1370_0[0]),.doutb(w_n1370_0[1]),.din(n1370));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(n1373));
	jspl jspl_w_n1374_0(.douta(w_n1374_0[0]),.doutb(w_n1374_0[1]),.din(n1374));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(n1376));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(n1378));
	jspl jspl_w_n1379_0(.douta(w_n1379_0[0]),.doutb(w_n1379_0[1]),.din(n1379));
	jspl jspl_w_n1384_0(.douta(w_n1384_0[0]),.doutb(w_n1384_0[1]),.din(n1384));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(n1389));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(n1390));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(n1395));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(n1400));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl jspl_w_n1408_0(.douta(w_n1408_0[0]),.doutb(w_n1408_0[1]),.din(n1408));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(n1410));
	jspl jspl_w_n1413_0(.douta(w_n1413_0[0]),.doutb(w_n1413_0[1]),.din(n1413));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(n1415));
	jspl jspl_w_n1418_0(.douta(w_n1418_0[0]),.doutb(w_n1418_0[1]),.din(n1418));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(n1420));
	jspl jspl_w_n1423_0(.douta(w_n1423_0[0]),.doutb(w_n1423_0[1]),.din(n1423));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(n1428));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1430_0(.douta(w_n1430_0[0]),.doutb(w_n1430_0[1]),.din(n1430));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1435_0(.douta(w_n1435_0[0]),.doutb(w_n1435_0[1]),.din(n1435));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(n1436));
	jspl jspl_w_n1437_0(.douta(w_n1437_0[0]),.doutb(w_n1437_0[1]),.din(n1437));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_n1438_0[1]),.din(n1438));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.din(n1440));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl jspl_w_n1442_0(.douta(w_n1442_0[0]),.doutb(w_n1442_0[1]),.din(n1442));
	jspl jspl_w_n1443_0(.douta(w_n1443_0[0]),.doutb(w_n1443_0[1]),.din(n1443));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(n1444));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1448_0(.douta(w_n1448_0[0]),.doutb(w_n1448_0[1]),.din(n1448));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(n1449));
	jspl jspl_w_n1450_0(.douta(w_n1450_0[0]),.doutb(w_n1450_0[1]),.din(n1450));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(n1454));
	jspl jspl_w_n1455_0(.douta(w_n1455_0[0]),.doutb(w_n1455_0[1]),.din(n1455));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(n1460));
	jspl jspl_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.din(n1465));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(n1466));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(n1471));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(n1474));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(n1476));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(n1479));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(n1481));
	jspl jspl_w_n1484_0(.douta(w_n1484_0[0]),.doutb(w_n1484_0[1]),.din(n1484));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(n1486));
	jspl jspl_w_n1489_0(.douta(w_n1489_0[0]),.doutb(w_n1489_0[1]),.din(n1489));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(n1491));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(n1494));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(n1496));
	jspl jspl_w_n1499_0(.douta(w_n1499_0[0]),.doutb(w_n1499_0[1]),.din(n1499));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(n1500));
	jspl jspl_w_n1501_0(.douta(w_n1501_0[0]),.doutb(w_n1501_0[1]),.din(n1501));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.din(n1506));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(n1507));
	jspl jspl_w_n1508_0(.douta(w_n1508_0[0]),.doutb(w_n1508_0[1]),.din(n1508));
	jspl jspl_w_n1509_0(.douta(w_n1509_0[0]),.doutb(w_n1509_0[1]),.din(n1509));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1511_0(.douta(w_n1511_0[0]),.doutb(w_n1511_0[1]),.din(n1511));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(n1512));
	jspl jspl_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.din(n1513));
	jspl jspl_w_n1514_0(.douta(w_n1514_0[0]),.doutb(w_n1514_0[1]),.din(n1514));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(n1515));
	jspl jspl_w_n1516_0(.douta(w_n1516_0[0]),.doutb(w_n1516_0[1]),.din(n1516));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(n1517));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1519_0(.douta(w_n1519_0[0]),.doutb(w_n1519_0[1]),.din(n1519));
	jspl jspl_w_n1521_0(.douta(w_n1521_0[0]),.doutb(w_n1521_0[1]),.din(n1521));
	jspl jspl_w_n1523_0(.douta(w_n1523_0[0]),.doutb(w_n1523_0[1]),.din(n1523));
	jspl jspl_w_n1524_0(.douta(w_n1524_0[0]),.doutb(w_n1524_0[1]),.din(n1524));
	jspl jspl_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.din(n1529));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(n1534));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(n1535));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(n1540));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(n1548));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_n1550_0[1]),.din(n1550));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(n1553));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(n1555));
	jspl jspl_w_n1558_0(.douta(w_n1558_0[0]),.doutb(w_n1558_0[1]),.din(n1558));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1563_0(.douta(w_n1563_0[0]),.doutb(w_n1563_0[1]),.din(n1563));
	jspl jspl_w_n1564_0(.douta(w_n1564_0[0]),.doutb(w_n1564_0[1]),.din(n1564));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(n1565));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_n1568_0[1]),.din(n1568));
	jspl jspl_w_n1570_0(.douta(w_n1570_0[0]),.doutb(w_n1570_0[1]),.din(n1570));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(n1571));
	jspl jspl_w_n1572_0(.douta(w_n1572_0[0]),.doutb(w_n1572_0[1]),.din(n1572));
	jspl jspl_w_n1573_0(.douta(w_n1573_0[0]),.doutb(w_n1573_0[1]),.din(n1573));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(n1574));
	jspl jspl_w_n1575_0(.douta(w_n1575_0[0]),.doutb(w_n1575_0[1]),.din(n1575));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(n1576));
	jspl jspl_w_n1577_0(.douta(w_n1577_0[0]),.doutb(w_n1577_0[1]),.din(n1577));
	jspl jspl_w_n1578_0(.douta(w_n1578_0[0]),.doutb(w_n1578_0[1]),.din(n1578));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(n1579));
	jspl jspl_w_n1580_0(.douta(w_n1580_0[0]),.doutb(w_n1580_0[1]),.din(n1580));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_n1581_0[1]),.din(n1581));
	jspl jspl_w_n1583_0(.douta(w_n1583_0[0]),.doutb(w_n1583_0[1]),.din(n1583));
	jspl jspl_w_n1585_0(.douta(w_n1585_0[0]),.doutb(w_n1585_0[1]),.din(n1585));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.din(n1586));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(n1597));
	jspl jspl_w_n1600_0(.douta(w_n1600_0[0]),.doutb(w_n1600_0[1]),.din(n1600));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(n1612));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(n1615));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_n1617_0[1]),.din(n1617));
	jspl jspl_w_n1620_0(.douta(w_n1620_0[0]),.doutb(w_n1620_0[1]),.din(n1620));
	jspl jspl_w_n1621_0(.douta(w_n1621_0[0]),.doutb(w_n1621_0[1]),.din(n1621));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(n1622));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(n1628));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1630_0(.douta(w_n1630_0[0]),.doutb(w_n1630_0[1]),.din(n1630));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(n1631));
	jspl jspl_w_n1632_0(.douta(w_n1632_0[0]),.doutb(w_n1632_0[1]),.din(n1632));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(n1633));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(n1634));
	jspl jspl_w_n1635_0(.douta(w_n1635_0[0]),.doutb(w_n1635_0[1]),.din(n1635));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(n1636));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(n1638));
	jspl jspl_w_n1640_0(.douta(w_n1640_0[0]),.doutb(w_n1640_0[1]),.din(n1640));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_n1641_0[1]),.din(n1641));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(n1646));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(n1651));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(n1653));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(n1656));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(n1658));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(n1661));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(n1663));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(n1666));
	jspl jspl_w_n1668_0(.douta(w_n1668_0[0]),.doutb(w_n1668_0[1]),.din(n1668));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(n1671));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(n1672));
	jspl jspl_w_n1673_0(.douta(w_n1673_0[0]),.doutb(w_n1673_0[1]),.din(n1673));
	jspl jspl_w_n1676_0(.douta(w_n1676_0[0]),.doutb(w_n1676_0[1]),.din(n1676));
	jspl jspl_w_n1678_0(.douta(w_n1678_0[0]),.doutb(w_n1678_0[1]),.din(n1678));
	jspl jspl_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1681_0(.douta(w_n1681_0[0]),.doutb(w_n1681_0[1]),.din(n1681));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(n1682));
	jspl jspl_w_n1683_0(.douta(w_n1683_0[0]),.doutb(w_n1683_0[1]),.din(n1683));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(n1684));
	jspl jspl_w_n1685_0(.douta(w_n1685_0[0]),.doutb(w_n1685_0[1]),.din(n1685));
	jspl jspl_w_n1686_0(.douta(w_n1686_0[0]),.doutb(w_n1686_0[1]),.din(n1686));
	jspl jspl_w_n1688_0(.douta(w_n1688_0[0]),.doutb(w_n1688_0[1]),.din(n1688));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(n1689));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(n1694));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_n1697_0[1]),.din(n1697));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(n1699));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(n1702));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(n1704));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(n1707));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(n1709));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(n1712));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(n1713));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(n1714));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_n1720_0[1]),.din(n1720));
	jspl jspl_w_n1721_0(.douta(w_n1721_0[0]),.doutb(w_n1721_0[1]),.din(n1721));
	jspl jspl_w_n1722_0(.douta(w_n1722_0[0]),.doutb(w_n1722_0[1]),.din(n1722));
	jspl jspl_w_n1723_0(.douta(w_n1723_0[0]),.doutb(w_n1723_0[1]),.din(n1723));
	jspl jspl_w_n1724_0(.douta(w_n1724_0[0]),.doutb(w_n1724_0[1]),.din(n1724));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1726_0(.douta(w_n1726_0[0]),.doutb(w_n1726_0[1]),.din(n1726));
	jspl jspl_w_n1727_0(.douta(w_n1727_0[0]),.doutb(w_n1727_0[1]),.din(n1727));
	jspl jspl_w_n1734_0(.douta(w_n1734_0[0]),.doutb(w_n1734_0[1]),.din(n1734));
	jspl jspl_w_n1737_0(.douta(w_n1737_0[0]),.doutb(w_n1737_0[1]),.din(n1737));
	jspl jspl_w_n1739_0(.douta(w_n1739_0[0]),.doutb(w_n1739_0[1]),.din(n1739));
	jspl jspl_w_n1742_0(.douta(w_n1742_0[0]),.doutb(w_n1742_0[1]),.din(n1742));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(n1744));
	jspl jspl_w_n1747_0(.douta(w_n1747_0[0]),.doutb(w_n1747_0[1]),.din(n1747));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(n1748));
	jspl jspl_w_n1749_0(.douta(w_n1749_0[0]),.doutb(w_n1749_0[1]),.din(n1749));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_n1758_0[1]),.din(n1758));
	jspl jspl_w_n1759_0(.douta(w_n1759_0[0]),.doutb(w_n1759_0[1]),.din(n1759));
	jspl jspl_w_n1760_0(.douta(w_n1760_0[0]),.doutb(w_n1760_0[1]),.din(n1760));
	jspl jspl_w_n1767_0(.douta(w_n1767_0[0]),.doutb(w_n1767_0[1]),.din(n1767));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(n1770));
	jspl jspl_w_n1772_0(.douta(w_n1772_0[0]),.doutb(w_n1772_0[1]),.din(n1772));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(n1775));
	jspl jspl_w_n1776_0(.douta(w_n1776_0[0]),.doutb(w_n1776_0[1]),.din(n1776));
	jspl jspl_w_n1777_0(.douta(w_n1777_0[0]),.doutb(w_n1777_0[1]),.din(n1777));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(n1780));
	jspl jspl_w_n1782_0(.douta(w_n1782_0[0]),.doutb(w_n1782_0[1]),.din(n1782));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1784_0(.douta(w_n1784_0[0]),.doutb(w_n1784_0[1]),.din(n1784));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_n1786_0[1]),.din(n1786));
	jspl jspl_w_n1793_0(.douta(w_n1793_0[0]),.doutb(w_n1793_0[1]),.din(n1793));
	jspl jspl_w_n1796_0(.douta(w_n1796_0[0]),.doutb(w_n1796_0[1]),.din(n1796));
	jspl jspl_w_n1797_0(.douta(w_n1797_0[0]),.doutb(w_n1797_0[1]),.din(n1797));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(n1798));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_n1801_0[1]),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(n1803));
	jspl jspl_w_n1804_0(.douta(w_n1804_0[0]),.doutb(w_n1804_0[1]),.din(n1804));
	jspl jspl_w_n1805_0(.douta(w_n1805_0[0]),.doutb(w_n1805_0[1]),.din(n1805));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(n1807));
	jspl jspl_w_n1810_0(.douta(w_n1810_0[0]),.doutb(w_n1810_0[1]),.din(n1810));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_n1817_0[1]),.din(n1817));
	jspl jspl_w_n1818_0(.douta(w_n1818_0[0]),.doutb(w_n1818_0[1]),.din(n1818));
	jdff dff_B_DmmoZnUj4_1(.din(n76),.dout(w_dff_B_DmmoZnUj4_1),.clk(gclk));
	jdff dff_B_O5UfwTMy7_1(.din(w_dff_B_DmmoZnUj4_1),.dout(w_dff_B_O5UfwTMy7_1),.clk(gclk));
	jdff dff_B_8vD6sN1d2_1(.din(w_dff_B_O5UfwTMy7_1),.dout(w_dff_B_8vD6sN1d2_1),.clk(gclk));
	jdff dff_B_Hiz3iM2k5_1(.din(n87),.dout(w_dff_B_Hiz3iM2k5_1),.clk(gclk));
	jdff dff_B_m1Ii7war6_1(.din(w_dff_B_Hiz3iM2k5_1),.dout(w_dff_B_m1Ii7war6_1),.clk(gclk));
	jdff dff_B_hYO5RUoD3_1(.din(w_dff_B_m1Ii7war6_1),.dout(w_dff_B_hYO5RUoD3_1),.clk(gclk));
	jdff dff_B_Hwgr4myO5_1(.din(w_dff_B_hYO5RUoD3_1),.dout(w_dff_B_Hwgr4myO5_1),.clk(gclk));
	jdff dff_B_qNxmAhNK9_1(.din(w_dff_B_Hwgr4myO5_1),.dout(w_dff_B_qNxmAhNK9_1),.clk(gclk));
	jdff dff_B_VEfEsqjZ4_1(.din(w_dff_B_qNxmAhNK9_1),.dout(w_dff_B_VEfEsqjZ4_1),.clk(gclk));
	jdff dff_B_8KXu2Zag5_1(.din(n107),.dout(w_dff_B_8KXu2Zag5_1),.clk(gclk));
	jdff dff_B_uIY1MvCi2_1(.din(w_dff_B_8KXu2Zag5_1),.dout(w_dff_B_uIY1MvCi2_1),.clk(gclk));
	jdff dff_B_G16ejBdK8_1(.din(w_dff_B_uIY1MvCi2_1),.dout(w_dff_B_G16ejBdK8_1),.clk(gclk));
	jdff dff_B_Njl0MimF5_1(.din(w_dff_B_G16ejBdK8_1),.dout(w_dff_B_Njl0MimF5_1),.clk(gclk));
	jdff dff_B_DdDQfMAb4_1(.din(w_dff_B_Njl0MimF5_1),.dout(w_dff_B_DdDQfMAb4_1),.clk(gclk));
	jdff dff_B_08DDgJsb9_1(.din(w_dff_B_DdDQfMAb4_1),.dout(w_dff_B_08DDgJsb9_1),.clk(gclk));
	jdff dff_B_6YBjp3va1_1(.din(w_dff_B_08DDgJsb9_1),.dout(w_dff_B_6YBjp3va1_1),.clk(gclk));
	jdff dff_B_pl8hv5cK9_1(.din(w_dff_B_6YBjp3va1_1),.dout(w_dff_B_pl8hv5cK9_1),.clk(gclk));
	jdff dff_B_QGLP9ZNw7_1(.din(w_dff_B_pl8hv5cK9_1),.dout(w_dff_B_QGLP9ZNw7_1),.clk(gclk));
	jdff dff_B_k6vZhay37_1(.din(n136),.dout(w_dff_B_k6vZhay37_1),.clk(gclk));
	jdff dff_B_PXqvL3oF9_1(.din(w_dff_B_k6vZhay37_1),.dout(w_dff_B_PXqvL3oF9_1),.clk(gclk));
	jdff dff_B_m525AQQ50_1(.din(w_dff_B_PXqvL3oF9_1),.dout(w_dff_B_m525AQQ50_1),.clk(gclk));
	jdff dff_B_nsx5O4Gl8_1(.din(w_dff_B_m525AQQ50_1),.dout(w_dff_B_nsx5O4Gl8_1),.clk(gclk));
	jdff dff_B_Dw3YggC90_1(.din(w_dff_B_nsx5O4Gl8_1),.dout(w_dff_B_Dw3YggC90_1),.clk(gclk));
	jdff dff_B_oJoOm4SQ7_1(.din(w_dff_B_Dw3YggC90_1),.dout(w_dff_B_oJoOm4SQ7_1),.clk(gclk));
	jdff dff_B_LnvdU34o4_1(.din(w_dff_B_oJoOm4SQ7_1),.dout(w_dff_B_LnvdU34o4_1),.clk(gclk));
	jdff dff_B_6LbTY0Pz3_1(.din(w_dff_B_LnvdU34o4_1),.dout(w_dff_B_6LbTY0Pz3_1),.clk(gclk));
	jdff dff_B_uLNTgwOp2_1(.din(w_dff_B_6LbTY0Pz3_1),.dout(w_dff_B_uLNTgwOp2_1),.clk(gclk));
	jdff dff_B_gwscHMSo7_1(.din(w_dff_B_uLNTgwOp2_1),.dout(w_dff_B_gwscHMSo7_1),.clk(gclk));
	jdff dff_B_hMbcC3mw6_1(.din(w_dff_B_gwscHMSo7_1),.dout(w_dff_B_hMbcC3mw6_1),.clk(gclk));
	jdff dff_B_zKlZiXNS1_1(.din(w_dff_B_hMbcC3mw6_1),.dout(w_dff_B_zKlZiXNS1_1),.clk(gclk));
	jdff dff_B_AnSItq1I2_1(.din(n171),.dout(w_dff_B_AnSItq1I2_1),.clk(gclk));
	jdff dff_B_yjgmjPdQ9_1(.din(w_dff_B_AnSItq1I2_1),.dout(w_dff_B_yjgmjPdQ9_1),.clk(gclk));
	jdff dff_B_SdH9pkK08_1(.din(w_dff_B_yjgmjPdQ9_1),.dout(w_dff_B_SdH9pkK08_1),.clk(gclk));
	jdff dff_B_Ngrtt6ca2_1(.din(w_dff_B_SdH9pkK08_1),.dout(w_dff_B_Ngrtt6ca2_1),.clk(gclk));
	jdff dff_B_VMrmjhAN3_1(.din(w_dff_B_Ngrtt6ca2_1),.dout(w_dff_B_VMrmjhAN3_1),.clk(gclk));
	jdff dff_B_gzsugydL4_1(.din(w_dff_B_VMrmjhAN3_1),.dout(w_dff_B_gzsugydL4_1),.clk(gclk));
	jdff dff_B_3T1e59ex9_1(.din(w_dff_B_gzsugydL4_1),.dout(w_dff_B_3T1e59ex9_1),.clk(gclk));
	jdff dff_B_biLnVCNd4_1(.din(w_dff_B_3T1e59ex9_1),.dout(w_dff_B_biLnVCNd4_1),.clk(gclk));
	jdff dff_B_Z3eSmBT88_1(.din(w_dff_B_biLnVCNd4_1),.dout(w_dff_B_Z3eSmBT88_1),.clk(gclk));
	jdff dff_B_hbLGiVVl0_1(.din(w_dff_B_Z3eSmBT88_1),.dout(w_dff_B_hbLGiVVl0_1),.clk(gclk));
	jdff dff_B_Oj9lc4aV7_1(.din(w_dff_B_hbLGiVVl0_1),.dout(w_dff_B_Oj9lc4aV7_1),.clk(gclk));
	jdff dff_B_zo2drDBd7_1(.din(w_dff_B_Oj9lc4aV7_1),.dout(w_dff_B_zo2drDBd7_1),.clk(gclk));
	jdff dff_B_ouqWyAAx4_1(.din(w_dff_B_zo2drDBd7_1),.dout(w_dff_B_ouqWyAAx4_1),.clk(gclk));
	jdff dff_B_v0WLDwnZ3_1(.din(w_dff_B_ouqWyAAx4_1),.dout(w_dff_B_v0WLDwnZ3_1),.clk(gclk));
	jdff dff_B_GF8o5Vdy5_1(.din(w_dff_B_v0WLDwnZ3_1),.dout(w_dff_B_GF8o5Vdy5_1),.clk(gclk));
	jdff dff_B_iujrpnet2_1(.din(n213),.dout(w_dff_B_iujrpnet2_1),.clk(gclk));
	jdff dff_B_eJp8CXws4_1(.din(w_dff_B_iujrpnet2_1),.dout(w_dff_B_eJp8CXws4_1),.clk(gclk));
	jdff dff_B_KgmnRMDg9_1(.din(w_dff_B_eJp8CXws4_1),.dout(w_dff_B_KgmnRMDg9_1),.clk(gclk));
	jdff dff_B_4maCP0DT9_1(.din(w_dff_B_KgmnRMDg9_1),.dout(w_dff_B_4maCP0DT9_1),.clk(gclk));
	jdff dff_B_fD0zaANk0_1(.din(w_dff_B_4maCP0DT9_1),.dout(w_dff_B_fD0zaANk0_1),.clk(gclk));
	jdff dff_B_frvYvEMt1_1(.din(w_dff_B_fD0zaANk0_1),.dout(w_dff_B_frvYvEMt1_1),.clk(gclk));
	jdff dff_B_C8DKEqdO0_1(.din(w_dff_B_frvYvEMt1_1),.dout(w_dff_B_C8DKEqdO0_1),.clk(gclk));
	jdff dff_B_auOkeWc03_1(.din(w_dff_B_C8DKEqdO0_1),.dout(w_dff_B_auOkeWc03_1),.clk(gclk));
	jdff dff_B_ClUzhLj95_1(.din(w_dff_B_auOkeWc03_1),.dout(w_dff_B_ClUzhLj95_1),.clk(gclk));
	jdff dff_B_pbZBQBQ81_1(.din(w_dff_B_ClUzhLj95_1),.dout(w_dff_B_pbZBQBQ81_1),.clk(gclk));
	jdff dff_B_w5UJ3Hr82_1(.din(w_dff_B_pbZBQBQ81_1),.dout(w_dff_B_w5UJ3Hr82_1),.clk(gclk));
	jdff dff_B_lzMtvHSY7_1(.din(w_dff_B_w5UJ3Hr82_1),.dout(w_dff_B_lzMtvHSY7_1),.clk(gclk));
	jdff dff_B_3Uw4ZDel3_1(.din(w_dff_B_lzMtvHSY7_1),.dout(w_dff_B_3Uw4ZDel3_1),.clk(gclk));
	jdff dff_B_IJvDkFa97_1(.din(w_dff_B_3Uw4ZDel3_1),.dout(w_dff_B_IJvDkFa97_1),.clk(gclk));
	jdff dff_B_GeJ4GHtm9_1(.din(w_dff_B_IJvDkFa97_1),.dout(w_dff_B_GeJ4GHtm9_1),.clk(gclk));
	jdff dff_B_n3OKOcXa8_1(.din(w_dff_B_GeJ4GHtm9_1),.dout(w_dff_B_n3OKOcXa8_1),.clk(gclk));
	jdff dff_B_MHon3vc79_1(.din(w_dff_B_n3OKOcXa8_1),.dout(w_dff_B_MHon3vc79_1),.clk(gclk));
	jdff dff_B_789OLFB94_1(.din(w_dff_B_MHon3vc79_1),.dout(w_dff_B_789OLFB94_1),.clk(gclk));
	jdff dff_B_b5QkdwGE9_1(.din(n262),.dout(w_dff_B_b5QkdwGE9_1),.clk(gclk));
	jdff dff_B_WAFfsglX3_1(.din(w_dff_B_b5QkdwGE9_1),.dout(w_dff_B_WAFfsglX3_1),.clk(gclk));
	jdff dff_B_erwi466O1_1(.din(w_dff_B_WAFfsglX3_1),.dout(w_dff_B_erwi466O1_1),.clk(gclk));
	jdff dff_B_BWUk9T503_1(.din(w_dff_B_erwi466O1_1),.dout(w_dff_B_BWUk9T503_1),.clk(gclk));
	jdff dff_B_riPkWCzu2_1(.din(w_dff_B_BWUk9T503_1),.dout(w_dff_B_riPkWCzu2_1),.clk(gclk));
	jdff dff_B_TvYmVkVV7_1(.din(w_dff_B_riPkWCzu2_1),.dout(w_dff_B_TvYmVkVV7_1),.clk(gclk));
	jdff dff_B_WSehINEJ4_1(.din(w_dff_B_TvYmVkVV7_1),.dout(w_dff_B_WSehINEJ4_1),.clk(gclk));
	jdff dff_B_lKdWkEuU0_1(.din(w_dff_B_WSehINEJ4_1),.dout(w_dff_B_lKdWkEuU0_1),.clk(gclk));
	jdff dff_B_YdG3jBos4_1(.din(w_dff_B_lKdWkEuU0_1),.dout(w_dff_B_YdG3jBos4_1),.clk(gclk));
	jdff dff_B_iHggrrry0_1(.din(w_dff_B_YdG3jBos4_1),.dout(w_dff_B_iHggrrry0_1),.clk(gclk));
	jdff dff_B_QQRsESRT6_1(.din(w_dff_B_iHggrrry0_1),.dout(w_dff_B_QQRsESRT6_1),.clk(gclk));
	jdff dff_B_4nhTHUpg6_1(.din(w_dff_B_QQRsESRT6_1),.dout(w_dff_B_4nhTHUpg6_1),.clk(gclk));
	jdff dff_B_jLRJMcJm6_1(.din(w_dff_B_4nhTHUpg6_1),.dout(w_dff_B_jLRJMcJm6_1),.clk(gclk));
	jdff dff_B_vF4XRc2B8_1(.din(w_dff_B_jLRJMcJm6_1),.dout(w_dff_B_vF4XRc2B8_1),.clk(gclk));
	jdff dff_B_2LLpG0Jk0_1(.din(w_dff_B_vF4XRc2B8_1),.dout(w_dff_B_2LLpG0Jk0_1),.clk(gclk));
	jdff dff_B_xVKTvnKl8_1(.din(w_dff_B_2LLpG0Jk0_1),.dout(w_dff_B_xVKTvnKl8_1),.clk(gclk));
	jdff dff_B_PtGgImiU4_1(.din(w_dff_B_xVKTvnKl8_1),.dout(w_dff_B_PtGgImiU4_1),.clk(gclk));
	jdff dff_B_gXr6bPCJ7_1(.din(w_dff_B_PtGgImiU4_1),.dout(w_dff_B_gXr6bPCJ7_1),.clk(gclk));
	jdff dff_B_om5bBsvF4_1(.din(w_dff_B_gXr6bPCJ7_1),.dout(w_dff_B_om5bBsvF4_1),.clk(gclk));
	jdff dff_B_NsSxQTMb8_1(.din(w_dff_B_om5bBsvF4_1),.dout(w_dff_B_NsSxQTMb8_1),.clk(gclk));
	jdff dff_B_fQ9WsX7z0_1(.din(w_dff_B_NsSxQTMb8_1),.dout(w_dff_B_fQ9WsX7z0_1),.clk(gclk));
	jdff dff_B_01aOoW4c3_1(.din(n318),.dout(w_dff_B_01aOoW4c3_1),.clk(gclk));
	jdff dff_B_IcpXjXpr1_1(.din(w_dff_B_01aOoW4c3_1),.dout(w_dff_B_IcpXjXpr1_1),.clk(gclk));
	jdff dff_B_uZk2Emv61_1(.din(w_dff_B_IcpXjXpr1_1),.dout(w_dff_B_uZk2Emv61_1),.clk(gclk));
	jdff dff_B_WoJNcMIQ1_1(.din(w_dff_B_uZk2Emv61_1),.dout(w_dff_B_WoJNcMIQ1_1),.clk(gclk));
	jdff dff_B_sgClU7AO7_1(.din(w_dff_B_WoJNcMIQ1_1),.dout(w_dff_B_sgClU7AO7_1),.clk(gclk));
	jdff dff_B_VPgk4d3B3_1(.din(w_dff_B_sgClU7AO7_1),.dout(w_dff_B_VPgk4d3B3_1),.clk(gclk));
	jdff dff_B_l9WwO8Mz0_1(.din(w_dff_B_VPgk4d3B3_1),.dout(w_dff_B_l9WwO8Mz0_1),.clk(gclk));
	jdff dff_B_oREOLxlD2_1(.din(w_dff_B_l9WwO8Mz0_1),.dout(w_dff_B_oREOLxlD2_1),.clk(gclk));
	jdff dff_B_Te1RunYj8_1(.din(w_dff_B_oREOLxlD2_1),.dout(w_dff_B_Te1RunYj8_1),.clk(gclk));
	jdff dff_B_MYxqiZYm4_1(.din(w_dff_B_Te1RunYj8_1),.dout(w_dff_B_MYxqiZYm4_1),.clk(gclk));
	jdff dff_B_vBaHb8ij5_1(.din(w_dff_B_MYxqiZYm4_1),.dout(w_dff_B_vBaHb8ij5_1),.clk(gclk));
	jdff dff_B_HMSZy4Na2_1(.din(w_dff_B_vBaHb8ij5_1),.dout(w_dff_B_HMSZy4Na2_1),.clk(gclk));
	jdff dff_B_rwXOrWtG3_1(.din(w_dff_B_HMSZy4Na2_1),.dout(w_dff_B_rwXOrWtG3_1),.clk(gclk));
	jdff dff_B_T5SjFso25_1(.din(w_dff_B_rwXOrWtG3_1),.dout(w_dff_B_T5SjFso25_1),.clk(gclk));
	jdff dff_B_HdcJeoIO2_1(.din(w_dff_B_T5SjFso25_1),.dout(w_dff_B_HdcJeoIO2_1),.clk(gclk));
	jdff dff_B_VJtWhcZw1_1(.din(w_dff_B_HdcJeoIO2_1),.dout(w_dff_B_VJtWhcZw1_1),.clk(gclk));
	jdff dff_B_vzUVOpRP1_1(.din(w_dff_B_VJtWhcZw1_1),.dout(w_dff_B_vzUVOpRP1_1),.clk(gclk));
	jdff dff_B_PI3sUmll9_1(.din(w_dff_B_vzUVOpRP1_1),.dout(w_dff_B_PI3sUmll9_1),.clk(gclk));
	jdff dff_B_P66p3rJ67_1(.din(w_dff_B_PI3sUmll9_1),.dout(w_dff_B_P66p3rJ67_1),.clk(gclk));
	jdff dff_B_MBRCpfmD5_1(.din(w_dff_B_P66p3rJ67_1),.dout(w_dff_B_MBRCpfmD5_1),.clk(gclk));
	jdff dff_B_CiTjA84y9_1(.din(w_dff_B_MBRCpfmD5_1),.dout(w_dff_B_CiTjA84y9_1),.clk(gclk));
	jdff dff_B_nun1b87I5_1(.din(w_dff_B_CiTjA84y9_1),.dout(w_dff_B_nun1b87I5_1),.clk(gclk));
	jdff dff_B_SW6JTjmV5_1(.din(w_dff_B_nun1b87I5_1),.dout(w_dff_B_SW6JTjmV5_1),.clk(gclk));
	jdff dff_B_OHdJphC50_1(.din(w_dff_B_SW6JTjmV5_1),.dout(w_dff_B_OHdJphC50_1),.clk(gclk));
	jdff dff_B_E8fcmvup6_1(.din(n381),.dout(w_dff_B_E8fcmvup6_1),.clk(gclk));
	jdff dff_B_E1nNgb8c2_1(.din(w_dff_B_E8fcmvup6_1),.dout(w_dff_B_E1nNgb8c2_1),.clk(gclk));
	jdff dff_B_Bwgm8y2A6_1(.din(w_dff_B_E1nNgb8c2_1),.dout(w_dff_B_Bwgm8y2A6_1),.clk(gclk));
	jdff dff_B_7S89rXFQ7_1(.din(w_dff_B_Bwgm8y2A6_1),.dout(w_dff_B_7S89rXFQ7_1),.clk(gclk));
	jdff dff_B_iP6K61Sy2_1(.din(w_dff_B_7S89rXFQ7_1),.dout(w_dff_B_iP6K61Sy2_1),.clk(gclk));
	jdff dff_B_IF1kwRy05_1(.din(w_dff_B_iP6K61Sy2_1),.dout(w_dff_B_IF1kwRy05_1),.clk(gclk));
	jdff dff_B_nG835zYk3_1(.din(w_dff_B_IF1kwRy05_1),.dout(w_dff_B_nG835zYk3_1),.clk(gclk));
	jdff dff_B_YEgrd9ZL2_1(.din(w_dff_B_nG835zYk3_1),.dout(w_dff_B_YEgrd9ZL2_1),.clk(gclk));
	jdff dff_B_fQSDUVuy2_1(.din(w_dff_B_YEgrd9ZL2_1),.dout(w_dff_B_fQSDUVuy2_1),.clk(gclk));
	jdff dff_B_mmhX7XXn8_1(.din(w_dff_B_fQSDUVuy2_1),.dout(w_dff_B_mmhX7XXn8_1),.clk(gclk));
	jdff dff_B_S8LpbVQ87_1(.din(w_dff_B_mmhX7XXn8_1),.dout(w_dff_B_S8LpbVQ87_1),.clk(gclk));
	jdff dff_B_qnXRm3zS1_1(.din(w_dff_B_S8LpbVQ87_1),.dout(w_dff_B_qnXRm3zS1_1),.clk(gclk));
	jdff dff_B_QO6Z7H856_1(.din(w_dff_B_qnXRm3zS1_1),.dout(w_dff_B_QO6Z7H856_1),.clk(gclk));
	jdff dff_B_8ZqH8pFz4_1(.din(w_dff_B_QO6Z7H856_1),.dout(w_dff_B_8ZqH8pFz4_1),.clk(gclk));
	jdff dff_B_jSivffm70_1(.din(w_dff_B_8ZqH8pFz4_1),.dout(w_dff_B_jSivffm70_1),.clk(gclk));
	jdff dff_B_yQQkW4Fa4_1(.din(w_dff_B_jSivffm70_1),.dout(w_dff_B_yQQkW4Fa4_1),.clk(gclk));
	jdff dff_B_JSeegWP58_1(.din(w_dff_B_yQQkW4Fa4_1),.dout(w_dff_B_JSeegWP58_1),.clk(gclk));
	jdff dff_B_4yHvPCnb6_1(.din(w_dff_B_JSeegWP58_1),.dout(w_dff_B_4yHvPCnb6_1),.clk(gclk));
	jdff dff_B_RD7qAJwj2_1(.din(w_dff_B_4yHvPCnb6_1),.dout(w_dff_B_RD7qAJwj2_1),.clk(gclk));
	jdff dff_B_3TJDN0bk5_1(.din(w_dff_B_RD7qAJwj2_1),.dout(w_dff_B_3TJDN0bk5_1),.clk(gclk));
	jdff dff_B_0Qj6UhC57_1(.din(w_dff_B_3TJDN0bk5_1),.dout(w_dff_B_0Qj6UhC57_1),.clk(gclk));
	jdff dff_B_yGi0Wq9I4_1(.din(w_dff_B_0Qj6UhC57_1),.dout(w_dff_B_yGi0Wq9I4_1),.clk(gclk));
	jdff dff_B_lOMoAspd9_1(.din(w_dff_B_yGi0Wq9I4_1),.dout(w_dff_B_lOMoAspd9_1),.clk(gclk));
	jdff dff_B_OySdTCav3_1(.din(w_dff_B_lOMoAspd9_1),.dout(w_dff_B_OySdTCav3_1),.clk(gclk));
	jdff dff_B_g7bMOlFS4_1(.din(w_dff_B_OySdTCav3_1),.dout(w_dff_B_g7bMOlFS4_1),.clk(gclk));
	jdff dff_B_eL0bZyCn8_1(.din(w_dff_B_g7bMOlFS4_1),.dout(w_dff_B_eL0bZyCn8_1),.clk(gclk));
	jdff dff_B_1wTyjv7c3_1(.din(w_dff_B_eL0bZyCn8_1),.dout(w_dff_B_1wTyjv7c3_1),.clk(gclk));
	jdff dff_B_TfdwRd9M2_1(.din(n452),.dout(w_dff_B_TfdwRd9M2_1),.clk(gclk));
	jdff dff_B_1M7MlyqW0_1(.din(w_dff_B_TfdwRd9M2_1),.dout(w_dff_B_1M7MlyqW0_1),.clk(gclk));
	jdff dff_B_AwPOeHeQ5_1(.din(w_dff_B_1M7MlyqW0_1),.dout(w_dff_B_AwPOeHeQ5_1),.clk(gclk));
	jdff dff_B_C2TYHHhe3_1(.din(w_dff_B_AwPOeHeQ5_1),.dout(w_dff_B_C2TYHHhe3_1),.clk(gclk));
	jdff dff_B_Pj8V49Ek7_1(.din(w_dff_B_C2TYHHhe3_1),.dout(w_dff_B_Pj8V49Ek7_1),.clk(gclk));
	jdff dff_B_3gJ76Ugx7_1(.din(w_dff_B_Pj8V49Ek7_1),.dout(w_dff_B_3gJ76Ugx7_1),.clk(gclk));
	jdff dff_B_Dbp9Iwf30_1(.din(w_dff_B_3gJ76Ugx7_1),.dout(w_dff_B_Dbp9Iwf30_1),.clk(gclk));
	jdff dff_B_tTTHKu3d4_1(.din(w_dff_B_Dbp9Iwf30_1),.dout(w_dff_B_tTTHKu3d4_1),.clk(gclk));
	jdff dff_B_Itb1kBIT1_1(.din(w_dff_B_tTTHKu3d4_1),.dout(w_dff_B_Itb1kBIT1_1),.clk(gclk));
	jdff dff_B_g54LDIIB1_1(.din(w_dff_B_Itb1kBIT1_1),.dout(w_dff_B_g54LDIIB1_1),.clk(gclk));
	jdff dff_B_Mzb6AKu96_1(.din(w_dff_B_g54LDIIB1_1),.dout(w_dff_B_Mzb6AKu96_1),.clk(gclk));
	jdff dff_B_VcHvAqnl4_1(.din(w_dff_B_Mzb6AKu96_1),.dout(w_dff_B_VcHvAqnl4_1),.clk(gclk));
	jdff dff_B_NGjKnrUm7_1(.din(w_dff_B_VcHvAqnl4_1),.dout(w_dff_B_NGjKnrUm7_1),.clk(gclk));
	jdff dff_B_Tip0e28S9_1(.din(w_dff_B_NGjKnrUm7_1),.dout(w_dff_B_Tip0e28S9_1),.clk(gclk));
	jdff dff_B_4ajDorjz4_1(.din(w_dff_B_Tip0e28S9_1),.dout(w_dff_B_4ajDorjz4_1),.clk(gclk));
	jdff dff_B_itTf6Q6w9_1(.din(w_dff_B_4ajDorjz4_1),.dout(w_dff_B_itTf6Q6w9_1),.clk(gclk));
	jdff dff_B_Kx8XthuG6_1(.din(w_dff_B_itTf6Q6w9_1),.dout(w_dff_B_Kx8XthuG6_1),.clk(gclk));
	jdff dff_B_DrkKKcom5_1(.din(w_dff_B_Kx8XthuG6_1),.dout(w_dff_B_DrkKKcom5_1),.clk(gclk));
	jdff dff_B_nzagnWGq2_1(.din(w_dff_B_DrkKKcom5_1),.dout(w_dff_B_nzagnWGq2_1),.clk(gclk));
	jdff dff_B_VXFgWWg23_1(.din(w_dff_B_nzagnWGq2_1),.dout(w_dff_B_VXFgWWg23_1),.clk(gclk));
	jdff dff_B_7vxnz7iE1_1(.din(w_dff_B_VXFgWWg23_1),.dout(w_dff_B_7vxnz7iE1_1),.clk(gclk));
	jdff dff_B_GMLGlu8i1_1(.din(w_dff_B_7vxnz7iE1_1),.dout(w_dff_B_GMLGlu8i1_1),.clk(gclk));
	jdff dff_B_UFxdavHd9_1(.din(w_dff_B_GMLGlu8i1_1),.dout(w_dff_B_UFxdavHd9_1),.clk(gclk));
	jdff dff_B_4QdrHxkM0_1(.din(w_dff_B_UFxdavHd9_1),.dout(w_dff_B_4QdrHxkM0_1),.clk(gclk));
	jdff dff_B_d8Cvow7m9_1(.din(w_dff_B_4QdrHxkM0_1),.dout(w_dff_B_d8Cvow7m9_1),.clk(gclk));
	jdff dff_B_NgFZ1CPf8_1(.din(w_dff_B_d8Cvow7m9_1),.dout(w_dff_B_NgFZ1CPf8_1),.clk(gclk));
	jdff dff_B_9G4RZfFC1_1(.din(w_dff_B_NgFZ1CPf8_1),.dout(w_dff_B_9G4RZfFC1_1),.clk(gclk));
	jdff dff_B_SPh3Sak03_1(.din(w_dff_B_9G4RZfFC1_1),.dout(w_dff_B_SPh3Sak03_1),.clk(gclk));
	jdff dff_B_Igyd8ruU9_1(.din(w_dff_B_SPh3Sak03_1),.dout(w_dff_B_Igyd8ruU9_1),.clk(gclk));
	jdff dff_B_fjZoUprZ9_1(.din(w_dff_B_Igyd8ruU9_1),.dout(w_dff_B_fjZoUprZ9_1),.clk(gclk));
	jdff dff_B_Txky5zgy7_1(.din(n530),.dout(w_dff_B_Txky5zgy7_1),.clk(gclk));
	jdff dff_B_k3FqqkVZ2_1(.din(w_dff_B_Txky5zgy7_1),.dout(w_dff_B_k3FqqkVZ2_1),.clk(gclk));
	jdff dff_B_J8ximAF64_1(.din(w_dff_B_k3FqqkVZ2_1),.dout(w_dff_B_J8ximAF64_1),.clk(gclk));
	jdff dff_B_GpjNY5Oc5_1(.din(w_dff_B_J8ximAF64_1),.dout(w_dff_B_GpjNY5Oc5_1),.clk(gclk));
	jdff dff_B_p4YATAlO1_1(.din(w_dff_B_GpjNY5Oc5_1),.dout(w_dff_B_p4YATAlO1_1),.clk(gclk));
	jdff dff_B_JiuUQjQD1_1(.din(w_dff_B_p4YATAlO1_1),.dout(w_dff_B_JiuUQjQD1_1),.clk(gclk));
	jdff dff_B_zmFQ6Vpz1_1(.din(w_dff_B_JiuUQjQD1_1),.dout(w_dff_B_zmFQ6Vpz1_1),.clk(gclk));
	jdff dff_B_m5V3H9j18_1(.din(w_dff_B_zmFQ6Vpz1_1),.dout(w_dff_B_m5V3H9j18_1),.clk(gclk));
	jdff dff_B_qWr93fEV4_1(.din(w_dff_B_m5V3H9j18_1),.dout(w_dff_B_qWr93fEV4_1),.clk(gclk));
	jdff dff_B_uHy60XbG0_1(.din(w_dff_B_qWr93fEV4_1),.dout(w_dff_B_uHy60XbG0_1),.clk(gclk));
	jdff dff_B_XUZEOL9G6_1(.din(w_dff_B_uHy60XbG0_1),.dout(w_dff_B_XUZEOL9G6_1),.clk(gclk));
	jdff dff_B_8oyR6nEv8_1(.din(w_dff_B_XUZEOL9G6_1),.dout(w_dff_B_8oyR6nEv8_1),.clk(gclk));
	jdff dff_B_6PbOU3cd5_1(.din(w_dff_B_8oyR6nEv8_1),.dout(w_dff_B_6PbOU3cd5_1),.clk(gclk));
	jdff dff_B_uVd8zuOI9_1(.din(w_dff_B_6PbOU3cd5_1),.dout(w_dff_B_uVd8zuOI9_1),.clk(gclk));
	jdff dff_B_6bLfUHjx3_1(.din(w_dff_B_uVd8zuOI9_1),.dout(w_dff_B_6bLfUHjx3_1),.clk(gclk));
	jdff dff_B_kzudbABd2_1(.din(w_dff_B_6bLfUHjx3_1),.dout(w_dff_B_kzudbABd2_1),.clk(gclk));
	jdff dff_B_Q4jqvAR08_1(.din(w_dff_B_kzudbABd2_1),.dout(w_dff_B_Q4jqvAR08_1),.clk(gclk));
	jdff dff_B_W7TQf5g40_1(.din(w_dff_B_Q4jqvAR08_1),.dout(w_dff_B_W7TQf5g40_1),.clk(gclk));
	jdff dff_B_Q72cJvuh4_1(.din(w_dff_B_W7TQf5g40_1),.dout(w_dff_B_Q72cJvuh4_1),.clk(gclk));
	jdff dff_B_HbUHzykR5_1(.din(w_dff_B_Q72cJvuh4_1),.dout(w_dff_B_HbUHzykR5_1),.clk(gclk));
	jdff dff_B_bdbcuCYw0_1(.din(w_dff_B_HbUHzykR5_1),.dout(w_dff_B_bdbcuCYw0_1),.clk(gclk));
	jdff dff_B_watOFMiZ3_1(.din(w_dff_B_bdbcuCYw0_1),.dout(w_dff_B_watOFMiZ3_1),.clk(gclk));
	jdff dff_B_wQVy7xhE5_1(.din(w_dff_B_watOFMiZ3_1),.dout(w_dff_B_wQVy7xhE5_1),.clk(gclk));
	jdff dff_B_mF1QKGRy0_1(.din(w_dff_B_wQVy7xhE5_1),.dout(w_dff_B_mF1QKGRy0_1),.clk(gclk));
	jdff dff_B_1yUxJ1x12_1(.din(w_dff_B_mF1QKGRy0_1),.dout(w_dff_B_1yUxJ1x12_1),.clk(gclk));
	jdff dff_B_OFUJJxNn0_1(.din(w_dff_B_1yUxJ1x12_1),.dout(w_dff_B_OFUJJxNn0_1),.clk(gclk));
	jdff dff_B_6heiRbpb6_1(.din(w_dff_B_OFUJJxNn0_1),.dout(w_dff_B_6heiRbpb6_1),.clk(gclk));
	jdff dff_B_BJJQTFvw0_1(.din(w_dff_B_6heiRbpb6_1),.dout(w_dff_B_BJJQTFvw0_1),.clk(gclk));
	jdff dff_B_ZtoLuE4X5_1(.din(w_dff_B_BJJQTFvw0_1),.dout(w_dff_B_ZtoLuE4X5_1),.clk(gclk));
	jdff dff_B_wYmjdvKH0_1(.din(w_dff_B_ZtoLuE4X5_1),.dout(w_dff_B_wYmjdvKH0_1),.clk(gclk));
	jdff dff_B_U6UQxXkn3_1(.din(w_dff_B_wYmjdvKH0_1),.dout(w_dff_B_U6UQxXkn3_1),.clk(gclk));
	jdff dff_B_gr5e1xZr5_1(.din(w_dff_B_U6UQxXkn3_1),.dout(w_dff_B_gr5e1xZr5_1),.clk(gclk));
	jdff dff_B_r1iAy6MU3_1(.din(w_dff_B_gr5e1xZr5_1),.dout(w_dff_B_r1iAy6MU3_1),.clk(gclk));
	jdff dff_B_1QC1TQcj0_1(.din(n615),.dout(w_dff_B_1QC1TQcj0_1),.clk(gclk));
	jdff dff_B_2Md8l1sc6_1(.din(w_dff_B_1QC1TQcj0_1),.dout(w_dff_B_2Md8l1sc6_1),.clk(gclk));
	jdff dff_B_cKCw7bBK8_1(.din(w_dff_B_2Md8l1sc6_1),.dout(w_dff_B_cKCw7bBK8_1),.clk(gclk));
	jdff dff_B_GEJAlnEN5_1(.din(w_dff_B_cKCw7bBK8_1),.dout(w_dff_B_GEJAlnEN5_1),.clk(gclk));
	jdff dff_B_ek1jnSIg9_1(.din(w_dff_B_GEJAlnEN5_1),.dout(w_dff_B_ek1jnSIg9_1),.clk(gclk));
	jdff dff_B_YJIGeZAa9_1(.din(w_dff_B_ek1jnSIg9_1),.dout(w_dff_B_YJIGeZAa9_1),.clk(gclk));
	jdff dff_B_067TIfkz4_1(.din(w_dff_B_YJIGeZAa9_1),.dout(w_dff_B_067TIfkz4_1),.clk(gclk));
	jdff dff_B_48s9u1u96_1(.din(w_dff_B_067TIfkz4_1),.dout(w_dff_B_48s9u1u96_1),.clk(gclk));
	jdff dff_B_smNr4rDx2_1(.din(w_dff_B_48s9u1u96_1),.dout(w_dff_B_smNr4rDx2_1),.clk(gclk));
	jdff dff_B_Em3nZ4jE4_1(.din(w_dff_B_smNr4rDx2_1),.dout(w_dff_B_Em3nZ4jE4_1),.clk(gclk));
	jdff dff_B_1I3uuWz87_1(.din(w_dff_B_Em3nZ4jE4_1),.dout(w_dff_B_1I3uuWz87_1),.clk(gclk));
	jdff dff_B_xt1bLtH50_1(.din(w_dff_B_1I3uuWz87_1),.dout(w_dff_B_xt1bLtH50_1),.clk(gclk));
	jdff dff_B_xdulWiE02_1(.din(w_dff_B_xt1bLtH50_1),.dout(w_dff_B_xdulWiE02_1),.clk(gclk));
	jdff dff_B_QkcW4NYo0_1(.din(w_dff_B_xdulWiE02_1),.dout(w_dff_B_QkcW4NYo0_1),.clk(gclk));
	jdff dff_B_6lLVEvrx1_1(.din(w_dff_B_QkcW4NYo0_1),.dout(w_dff_B_6lLVEvrx1_1),.clk(gclk));
	jdff dff_B_xi943vMI6_1(.din(w_dff_B_6lLVEvrx1_1),.dout(w_dff_B_xi943vMI6_1),.clk(gclk));
	jdff dff_B_4iijnvTh3_1(.din(w_dff_B_xi943vMI6_1),.dout(w_dff_B_4iijnvTh3_1),.clk(gclk));
	jdff dff_B_pfonSuJY5_1(.din(w_dff_B_4iijnvTh3_1),.dout(w_dff_B_pfonSuJY5_1),.clk(gclk));
	jdff dff_B_8BWcsDFe7_1(.din(w_dff_B_pfonSuJY5_1),.dout(w_dff_B_8BWcsDFe7_1),.clk(gclk));
	jdff dff_B_mNNeMzGq2_1(.din(w_dff_B_8BWcsDFe7_1),.dout(w_dff_B_mNNeMzGq2_1),.clk(gclk));
	jdff dff_B_uZ9pkRDC2_1(.din(w_dff_B_mNNeMzGq2_1),.dout(w_dff_B_uZ9pkRDC2_1),.clk(gclk));
	jdff dff_B_mbf7GveI3_1(.din(w_dff_B_uZ9pkRDC2_1),.dout(w_dff_B_mbf7GveI3_1),.clk(gclk));
	jdff dff_B_oScKx5Wf6_1(.din(w_dff_B_mbf7GveI3_1),.dout(w_dff_B_oScKx5Wf6_1),.clk(gclk));
	jdff dff_B_4AsiEg0h4_1(.din(w_dff_B_oScKx5Wf6_1),.dout(w_dff_B_4AsiEg0h4_1),.clk(gclk));
	jdff dff_B_DVKnjaKG7_1(.din(w_dff_B_4AsiEg0h4_1),.dout(w_dff_B_DVKnjaKG7_1),.clk(gclk));
	jdff dff_B_aUekxOjk4_1(.din(w_dff_B_DVKnjaKG7_1),.dout(w_dff_B_aUekxOjk4_1),.clk(gclk));
	jdff dff_B_jXgKvv612_1(.din(w_dff_B_aUekxOjk4_1),.dout(w_dff_B_jXgKvv612_1),.clk(gclk));
	jdff dff_B_r6dfayWB3_1(.din(w_dff_B_jXgKvv612_1),.dout(w_dff_B_r6dfayWB3_1),.clk(gclk));
	jdff dff_B_X2Jw8EXg6_1(.din(w_dff_B_r6dfayWB3_1),.dout(w_dff_B_X2Jw8EXg6_1),.clk(gclk));
	jdff dff_B_A46QaqN33_1(.din(w_dff_B_X2Jw8EXg6_1),.dout(w_dff_B_A46QaqN33_1),.clk(gclk));
	jdff dff_B_Yx74BAga0_1(.din(w_dff_B_A46QaqN33_1),.dout(w_dff_B_Yx74BAga0_1),.clk(gclk));
	jdff dff_B_P01OHjIW8_1(.din(w_dff_B_Yx74BAga0_1),.dout(w_dff_B_P01OHjIW8_1),.clk(gclk));
	jdff dff_B_4CgSfogD6_1(.din(w_dff_B_P01OHjIW8_1),.dout(w_dff_B_4CgSfogD6_1),.clk(gclk));
	jdff dff_B_WVCSxjUL1_1(.din(w_dff_B_4CgSfogD6_1),.dout(w_dff_B_WVCSxjUL1_1),.clk(gclk));
	jdff dff_B_5qykt55W7_1(.din(w_dff_B_WVCSxjUL1_1),.dout(w_dff_B_5qykt55W7_1),.clk(gclk));
	jdff dff_B_Vb5ZFRw32_1(.din(w_dff_B_5qykt55W7_1),.dout(w_dff_B_Vb5ZFRw32_1),.clk(gclk));
	jdff dff_B_k4jAsaKo7_1(.din(n707),.dout(w_dff_B_k4jAsaKo7_1),.clk(gclk));
	jdff dff_B_wpllafUx6_1(.din(w_dff_B_k4jAsaKo7_1),.dout(w_dff_B_wpllafUx6_1),.clk(gclk));
	jdff dff_B_EjYO7dmp8_1(.din(w_dff_B_wpllafUx6_1),.dout(w_dff_B_EjYO7dmp8_1),.clk(gclk));
	jdff dff_B_cxNaOFz90_1(.din(w_dff_B_EjYO7dmp8_1),.dout(w_dff_B_cxNaOFz90_1),.clk(gclk));
	jdff dff_B_LYsPiCCA0_1(.din(w_dff_B_cxNaOFz90_1),.dout(w_dff_B_LYsPiCCA0_1),.clk(gclk));
	jdff dff_B_xEiGVe7T2_1(.din(w_dff_B_LYsPiCCA0_1),.dout(w_dff_B_xEiGVe7T2_1),.clk(gclk));
	jdff dff_B_PmTPMPTs1_1(.din(w_dff_B_xEiGVe7T2_1),.dout(w_dff_B_PmTPMPTs1_1),.clk(gclk));
	jdff dff_B_gT3iJnmn0_1(.din(w_dff_B_PmTPMPTs1_1),.dout(w_dff_B_gT3iJnmn0_1),.clk(gclk));
	jdff dff_B_QpUILwRe9_1(.din(w_dff_B_gT3iJnmn0_1),.dout(w_dff_B_QpUILwRe9_1),.clk(gclk));
	jdff dff_B_ehNSmuTL9_1(.din(w_dff_B_QpUILwRe9_1),.dout(w_dff_B_ehNSmuTL9_1),.clk(gclk));
	jdff dff_B_9mU3c2q68_1(.din(w_dff_B_ehNSmuTL9_1),.dout(w_dff_B_9mU3c2q68_1),.clk(gclk));
	jdff dff_B_zDrUJLFD3_1(.din(w_dff_B_9mU3c2q68_1),.dout(w_dff_B_zDrUJLFD3_1),.clk(gclk));
	jdff dff_B_Uz5pXQIO1_1(.din(w_dff_B_zDrUJLFD3_1),.dout(w_dff_B_Uz5pXQIO1_1),.clk(gclk));
	jdff dff_B_ZEtmJWfV7_1(.din(w_dff_B_Uz5pXQIO1_1),.dout(w_dff_B_ZEtmJWfV7_1),.clk(gclk));
	jdff dff_B_HmSXNsVh9_1(.din(w_dff_B_ZEtmJWfV7_1),.dout(w_dff_B_HmSXNsVh9_1),.clk(gclk));
	jdff dff_B_mBI9FvqX1_1(.din(w_dff_B_HmSXNsVh9_1),.dout(w_dff_B_mBI9FvqX1_1),.clk(gclk));
	jdff dff_B_ojzThOHR2_1(.din(w_dff_B_mBI9FvqX1_1),.dout(w_dff_B_ojzThOHR2_1),.clk(gclk));
	jdff dff_B_Q89DwB954_1(.din(w_dff_B_ojzThOHR2_1),.dout(w_dff_B_Q89DwB954_1),.clk(gclk));
	jdff dff_B_Su6VguAg8_1(.din(w_dff_B_Q89DwB954_1),.dout(w_dff_B_Su6VguAg8_1),.clk(gclk));
	jdff dff_B_0sUkPOSg7_1(.din(w_dff_B_Su6VguAg8_1),.dout(w_dff_B_0sUkPOSg7_1),.clk(gclk));
	jdff dff_B_s0C5wQSf5_1(.din(w_dff_B_0sUkPOSg7_1),.dout(w_dff_B_s0C5wQSf5_1),.clk(gclk));
	jdff dff_B_sh8vrTxC4_1(.din(w_dff_B_s0C5wQSf5_1),.dout(w_dff_B_sh8vrTxC4_1),.clk(gclk));
	jdff dff_B_NFykJsdv1_1(.din(w_dff_B_sh8vrTxC4_1),.dout(w_dff_B_NFykJsdv1_1),.clk(gclk));
	jdff dff_B_ms9B5Xkn0_1(.din(w_dff_B_NFykJsdv1_1),.dout(w_dff_B_ms9B5Xkn0_1),.clk(gclk));
	jdff dff_B_8LtNSkZM8_1(.din(w_dff_B_ms9B5Xkn0_1),.dout(w_dff_B_8LtNSkZM8_1),.clk(gclk));
	jdff dff_B_Yp1W0ap52_1(.din(w_dff_B_8LtNSkZM8_1),.dout(w_dff_B_Yp1W0ap52_1),.clk(gclk));
	jdff dff_B_S0jgYNTv2_1(.din(w_dff_B_Yp1W0ap52_1),.dout(w_dff_B_S0jgYNTv2_1),.clk(gclk));
	jdff dff_B_IMlnEWuK7_1(.din(w_dff_B_S0jgYNTv2_1),.dout(w_dff_B_IMlnEWuK7_1),.clk(gclk));
	jdff dff_B_SafHHuqU4_1(.din(w_dff_B_IMlnEWuK7_1),.dout(w_dff_B_SafHHuqU4_1),.clk(gclk));
	jdff dff_B_onCF08pC7_1(.din(w_dff_B_SafHHuqU4_1),.dout(w_dff_B_onCF08pC7_1),.clk(gclk));
	jdff dff_B_tYhpkpMf6_1(.din(w_dff_B_onCF08pC7_1),.dout(w_dff_B_tYhpkpMf6_1),.clk(gclk));
	jdff dff_B_YSNgH7gA4_1(.din(w_dff_B_tYhpkpMf6_1),.dout(w_dff_B_YSNgH7gA4_1),.clk(gclk));
	jdff dff_B_0xOmQsRi1_1(.din(w_dff_B_YSNgH7gA4_1),.dout(w_dff_B_0xOmQsRi1_1),.clk(gclk));
	jdff dff_B_ZVn2BZEI0_1(.din(w_dff_B_0xOmQsRi1_1),.dout(w_dff_B_ZVn2BZEI0_1),.clk(gclk));
	jdff dff_B_xKtPHTX48_1(.din(w_dff_B_ZVn2BZEI0_1),.dout(w_dff_B_xKtPHTX48_1),.clk(gclk));
	jdff dff_B_XZmhVAb25_1(.din(w_dff_B_xKtPHTX48_1),.dout(w_dff_B_XZmhVAb25_1),.clk(gclk));
	jdff dff_B_0Dv6C3xd8_1(.din(w_dff_B_XZmhVAb25_1),.dout(w_dff_B_0Dv6C3xd8_1),.clk(gclk));
	jdff dff_B_H12TUS8Q4_1(.din(w_dff_B_0Dv6C3xd8_1),.dout(w_dff_B_H12TUS8Q4_1),.clk(gclk));
	jdff dff_B_khjF5Lua6_1(.din(w_dff_B_H12TUS8Q4_1),.dout(w_dff_B_khjF5Lua6_1),.clk(gclk));
	jdff dff_B_OCgX8gW97_1(.din(n806),.dout(w_dff_B_OCgX8gW97_1),.clk(gclk));
	jdff dff_B_G0f4VCiM3_1(.din(w_dff_B_OCgX8gW97_1),.dout(w_dff_B_G0f4VCiM3_1),.clk(gclk));
	jdff dff_B_Ay1LnXh60_1(.din(w_dff_B_G0f4VCiM3_1),.dout(w_dff_B_Ay1LnXh60_1),.clk(gclk));
	jdff dff_B_eeV9nUrs1_1(.din(w_dff_B_Ay1LnXh60_1),.dout(w_dff_B_eeV9nUrs1_1),.clk(gclk));
	jdff dff_B_JQsVcHQJ0_1(.din(w_dff_B_eeV9nUrs1_1),.dout(w_dff_B_JQsVcHQJ0_1),.clk(gclk));
	jdff dff_B_odtFOmT87_1(.din(w_dff_B_JQsVcHQJ0_1),.dout(w_dff_B_odtFOmT87_1),.clk(gclk));
	jdff dff_B_eKMZstAZ6_1(.din(w_dff_B_odtFOmT87_1),.dout(w_dff_B_eKMZstAZ6_1),.clk(gclk));
	jdff dff_B_gqklguIX4_1(.din(w_dff_B_eKMZstAZ6_1),.dout(w_dff_B_gqklguIX4_1),.clk(gclk));
	jdff dff_B_pgUahyWQ2_1(.din(w_dff_B_gqklguIX4_1),.dout(w_dff_B_pgUahyWQ2_1),.clk(gclk));
	jdff dff_B_PIYxYIMU9_1(.din(w_dff_B_pgUahyWQ2_1),.dout(w_dff_B_PIYxYIMU9_1),.clk(gclk));
	jdff dff_B_MCDpiy712_1(.din(w_dff_B_PIYxYIMU9_1),.dout(w_dff_B_MCDpiy712_1),.clk(gclk));
	jdff dff_B_DbLOSDb16_1(.din(w_dff_B_MCDpiy712_1),.dout(w_dff_B_DbLOSDb16_1),.clk(gclk));
	jdff dff_B_uQRAheUd0_1(.din(w_dff_B_DbLOSDb16_1),.dout(w_dff_B_uQRAheUd0_1),.clk(gclk));
	jdff dff_B_8VoKSApJ7_1(.din(w_dff_B_uQRAheUd0_1),.dout(w_dff_B_8VoKSApJ7_1),.clk(gclk));
	jdff dff_B_s4ffzqGG3_1(.din(w_dff_B_8VoKSApJ7_1),.dout(w_dff_B_s4ffzqGG3_1),.clk(gclk));
	jdff dff_B_cSoUArzT0_1(.din(w_dff_B_s4ffzqGG3_1),.dout(w_dff_B_cSoUArzT0_1),.clk(gclk));
	jdff dff_B_tnBYqjOd5_1(.din(w_dff_B_cSoUArzT0_1),.dout(w_dff_B_tnBYqjOd5_1),.clk(gclk));
	jdff dff_B_IoUnQinS4_1(.din(w_dff_B_tnBYqjOd5_1),.dout(w_dff_B_IoUnQinS4_1),.clk(gclk));
	jdff dff_B_2OxD9q6H5_1(.din(w_dff_B_IoUnQinS4_1),.dout(w_dff_B_2OxD9q6H5_1),.clk(gclk));
	jdff dff_B_GaWogtCT2_1(.din(w_dff_B_2OxD9q6H5_1),.dout(w_dff_B_GaWogtCT2_1),.clk(gclk));
	jdff dff_B_n5JMJ61k0_1(.din(w_dff_B_GaWogtCT2_1),.dout(w_dff_B_n5JMJ61k0_1),.clk(gclk));
	jdff dff_B_Cs2OmUco5_1(.din(w_dff_B_n5JMJ61k0_1),.dout(w_dff_B_Cs2OmUco5_1),.clk(gclk));
	jdff dff_B_wdxefOFN0_1(.din(w_dff_B_Cs2OmUco5_1),.dout(w_dff_B_wdxefOFN0_1),.clk(gclk));
	jdff dff_B_EFjaSjHT7_1(.din(w_dff_B_wdxefOFN0_1),.dout(w_dff_B_EFjaSjHT7_1),.clk(gclk));
	jdff dff_B_2hZlOMVi8_1(.din(w_dff_B_EFjaSjHT7_1),.dout(w_dff_B_2hZlOMVi8_1),.clk(gclk));
	jdff dff_B_QRhjZZyp0_1(.din(w_dff_B_2hZlOMVi8_1),.dout(w_dff_B_QRhjZZyp0_1),.clk(gclk));
	jdff dff_B_lUE2hNpe3_1(.din(w_dff_B_QRhjZZyp0_1),.dout(w_dff_B_lUE2hNpe3_1),.clk(gclk));
	jdff dff_B_V2SsRoJB9_1(.din(w_dff_B_lUE2hNpe3_1),.dout(w_dff_B_V2SsRoJB9_1),.clk(gclk));
	jdff dff_B_0HyguaWJ1_1(.din(w_dff_B_V2SsRoJB9_1),.dout(w_dff_B_0HyguaWJ1_1),.clk(gclk));
	jdff dff_B_j7rUtNQ01_1(.din(w_dff_B_0HyguaWJ1_1),.dout(w_dff_B_j7rUtNQ01_1),.clk(gclk));
	jdff dff_B_UH7q5hBH3_1(.din(w_dff_B_j7rUtNQ01_1),.dout(w_dff_B_UH7q5hBH3_1),.clk(gclk));
	jdff dff_B_9PjiUSgH4_1(.din(w_dff_B_UH7q5hBH3_1),.dout(w_dff_B_9PjiUSgH4_1),.clk(gclk));
	jdff dff_B_sP81te7Z0_1(.din(w_dff_B_9PjiUSgH4_1),.dout(w_dff_B_sP81te7Z0_1),.clk(gclk));
	jdff dff_B_Qm2w4L9n6_1(.din(w_dff_B_sP81te7Z0_1),.dout(w_dff_B_Qm2w4L9n6_1),.clk(gclk));
	jdff dff_B_NxbTxvB99_1(.din(w_dff_B_Qm2w4L9n6_1),.dout(w_dff_B_NxbTxvB99_1),.clk(gclk));
	jdff dff_B_p8VCotCh1_1(.din(w_dff_B_NxbTxvB99_1),.dout(w_dff_B_p8VCotCh1_1),.clk(gclk));
	jdff dff_B_pki0VitO5_1(.din(w_dff_B_p8VCotCh1_1),.dout(w_dff_B_pki0VitO5_1),.clk(gclk));
	jdff dff_B_XxB3sXCL9_1(.din(w_dff_B_pki0VitO5_1),.dout(w_dff_B_XxB3sXCL9_1),.clk(gclk));
	jdff dff_B_OSzEtGV39_1(.din(w_dff_B_XxB3sXCL9_1),.dout(w_dff_B_OSzEtGV39_1),.clk(gclk));
	jdff dff_B_VFotRj8h7_1(.din(w_dff_B_OSzEtGV39_1),.dout(w_dff_B_VFotRj8h7_1),.clk(gclk));
	jdff dff_B_6LtDBr7p7_1(.din(w_dff_B_VFotRj8h7_1),.dout(w_dff_B_6LtDBr7p7_1),.clk(gclk));
	jdff dff_B_jf1zmcsS5_1(.din(w_dff_B_6LtDBr7p7_1),.dout(w_dff_B_jf1zmcsS5_1),.clk(gclk));
	jdff dff_B_A72U7TVO7_0(.din(n1296),.dout(w_dff_B_A72U7TVO7_0),.clk(gclk));
	jdff dff_B_2bXHW5pD2_1(.din(n1811),.dout(w_dff_B_2bXHW5pD2_1),.clk(gclk));
	jdff dff_B_combaM0x6_1(.din(w_dff_B_2bXHW5pD2_1),.dout(w_dff_B_combaM0x6_1),.clk(gclk));
	jdff dff_B_WJlDsVAg4_1(.din(w_dff_B_combaM0x6_1),.dout(w_dff_B_WJlDsVAg4_1),.clk(gclk));
	jdff dff_B_6hfngCDd5_1(.din(w_dff_B_WJlDsVAg4_1),.dout(w_dff_B_6hfngCDd5_1),.clk(gclk));
	jdff dff_B_Whl6dzRx7_1(.din(w_dff_B_6hfngCDd5_1),.dout(w_dff_B_Whl6dzRx7_1),.clk(gclk));
	jdff dff_B_fowZhe165_1(.din(w_dff_B_Whl6dzRx7_1),.dout(w_dff_B_fowZhe165_1),.clk(gclk));
	jdff dff_B_tn22G5N56_1(.din(w_dff_B_fowZhe165_1),.dout(w_dff_B_tn22G5N56_1),.clk(gclk));
	jdff dff_B_5GRs5Cqd8_1(.din(w_dff_B_tn22G5N56_1),.dout(w_dff_B_5GRs5Cqd8_1),.clk(gclk));
	jdff dff_B_Q9aBr6lV2_1(.din(w_dff_B_5GRs5Cqd8_1),.dout(w_dff_B_Q9aBr6lV2_1),.clk(gclk));
	jdff dff_B_PY7RO6Vt7_1(.din(w_dff_B_Q9aBr6lV2_1),.dout(w_dff_B_PY7RO6Vt7_1),.clk(gclk));
	jdff dff_B_Fo5D8mPH4_1(.din(w_dff_B_PY7RO6Vt7_1),.dout(w_dff_B_Fo5D8mPH4_1),.clk(gclk));
	jdff dff_B_amOp1eBC0_1(.din(w_dff_B_Fo5D8mPH4_1),.dout(w_dff_B_amOp1eBC0_1),.clk(gclk));
	jdff dff_B_uGmmzoV76_1(.din(w_dff_B_amOp1eBC0_1),.dout(w_dff_B_uGmmzoV76_1),.clk(gclk));
	jdff dff_B_8WpZYETE2_1(.din(w_dff_B_uGmmzoV76_1),.dout(w_dff_B_8WpZYETE2_1),.clk(gclk));
	jdff dff_B_I6ALDGFU2_1(.din(w_dff_B_8WpZYETE2_1),.dout(w_dff_B_I6ALDGFU2_1),.clk(gclk));
	jdff dff_B_UODfp17m5_0(.din(n1819),.dout(w_dff_B_UODfp17m5_0),.clk(gclk));
	jdff dff_B_C2fgywuC4_0(.din(w_dff_B_UODfp17m5_0),.dout(w_dff_B_C2fgywuC4_0),.clk(gclk));
	jdff dff_B_iSNLeOj13_0(.din(w_dff_B_C2fgywuC4_0),.dout(w_dff_B_iSNLeOj13_0),.clk(gclk));
	jdff dff_B_ubllVIKr1_0(.din(w_dff_B_iSNLeOj13_0),.dout(w_dff_B_ubllVIKr1_0),.clk(gclk));
	jdff dff_B_sSHGz87U4_0(.din(w_dff_B_ubllVIKr1_0),.dout(w_dff_B_sSHGz87U4_0),.clk(gclk));
	jdff dff_B_WosEgbB53_0(.din(w_dff_B_sSHGz87U4_0),.dout(w_dff_B_WosEgbB53_0),.clk(gclk));
	jdff dff_B_AA7GTO5r1_0(.din(w_dff_B_WosEgbB53_0),.dout(w_dff_B_AA7GTO5r1_0),.clk(gclk));
	jdff dff_B_F6O6CMhn6_0(.din(w_dff_B_AA7GTO5r1_0),.dout(w_dff_B_F6O6CMhn6_0),.clk(gclk));
	jdff dff_B_NDvo4c0r1_0(.din(w_dff_B_F6O6CMhn6_0),.dout(w_dff_B_NDvo4c0r1_0),.clk(gclk));
	jdff dff_B_28455s062_0(.din(w_dff_B_NDvo4c0r1_0),.dout(w_dff_B_28455s062_0),.clk(gclk));
	jdff dff_B_rI9ZnYwA1_0(.din(w_dff_B_28455s062_0),.dout(w_dff_B_rI9ZnYwA1_0),.clk(gclk));
	jdff dff_B_hcUrSKa20_0(.din(w_dff_B_rI9ZnYwA1_0),.dout(w_dff_B_hcUrSKa20_0),.clk(gclk));
	jdff dff_B_7IAlXGz98_0(.din(w_dff_B_hcUrSKa20_0),.dout(w_dff_B_7IAlXGz98_0),.clk(gclk));
	jdff dff_B_vB92Z3wd0_1(.din(n1814),.dout(w_dff_B_vB92Z3wd0_1),.clk(gclk));
	jdff dff_B_1z2SjFgn6_1(.din(w_dff_B_vB92Z3wd0_1),.dout(w_dff_B_1z2SjFgn6_1),.clk(gclk));
	jdff dff_B_s7f3VCWp9_1(.din(w_dff_B_1z2SjFgn6_1),.dout(w_dff_B_s7f3VCWp9_1),.clk(gclk));
	jdff dff_B_6f5bYo4b0_1(.din(w_dff_B_s7f3VCWp9_1),.dout(w_dff_B_6f5bYo4b0_1),.clk(gclk));
	jdff dff_B_sMYlibVf4_1(.din(w_dff_B_6f5bYo4b0_1),.dout(w_dff_B_sMYlibVf4_1),.clk(gclk));
	jdff dff_B_y2bLOyBS9_1(.din(w_dff_B_sMYlibVf4_1),.dout(w_dff_B_y2bLOyBS9_1),.clk(gclk));
	jdff dff_B_Ag21fRFK7_1(.din(w_dff_B_y2bLOyBS9_1),.dout(w_dff_B_Ag21fRFK7_1),.clk(gclk));
	jdff dff_B_NU2rreoE3_1(.din(w_dff_B_Ag21fRFK7_1),.dout(w_dff_B_NU2rreoE3_1),.clk(gclk));
	jdff dff_B_20SpjbN58_1(.din(w_dff_B_NU2rreoE3_1),.dout(w_dff_B_20SpjbN58_1),.clk(gclk));
	jdff dff_B_ni4MjmfM3_1(.din(w_dff_B_20SpjbN58_1),.dout(w_dff_B_ni4MjmfM3_1),.clk(gclk));
	jdff dff_B_U4FBYWht0_1(.din(w_dff_B_ni4MjmfM3_1),.dout(w_dff_B_U4FBYWht0_1),.clk(gclk));
	jdff dff_B_6cBDMDFk1_1(.din(w_dff_B_U4FBYWht0_1),.dout(w_dff_B_6cBDMDFk1_1),.clk(gclk));
	jdff dff_B_5v4CRyGD2_1(.din(w_dff_B_6cBDMDFk1_1),.dout(w_dff_B_5v4CRyGD2_1),.clk(gclk));
	jdff dff_B_C0lRgFtL6_0(.din(n1815),.dout(w_dff_B_C0lRgFtL6_0),.clk(gclk));
	jdff dff_B_FaXRMAPW6_0(.din(w_dff_B_C0lRgFtL6_0),.dout(w_dff_B_FaXRMAPW6_0),.clk(gclk));
	jdff dff_B_bcklkbUS0_0(.din(w_dff_B_FaXRMAPW6_0),.dout(w_dff_B_bcklkbUS0_0),.clk(gclk));
	jdff dff_B_OWWRXFVB1_0(.din(w_dff_B_bcklkbUS0_0),.dout(w_dff_B_OWWRXFVB1_0),.clk(gclk));
	jdff dff_B_vFzvKk599_0(.din(w_dff_B_OWWRXFVB1_0),.dout(w_dff_B_vFzvKk599_0),.clk(gclk));
	jdff dff_B_wH2V0pic6_0(.din(w_dff_B_vFzvKk599_0),.dout(w_dff_B_wH2V0pic6_0),.clk(gclk));
	jdff dff_B_KuaPtgtw3_0(.din(w_dff_B_wH2V0pic6_0),.dout(w_dff_B_KuaPtgtw3_0),.clk(gclk));
	jdff dff_B_zcGSBZpn3_0(.din(w_dff_B_KuaPtgtw3_0),.dout(w_dff_B_zcGSBZpn3_0),.clk(gclk));
	jdff dff_B_yBE6hfya7_0(.din(w_dff_B_zcGSBZpn3_0),.dout(w_dff_B_yBE6hfya7_0),.clk(gclk));
	jdff dff_B_QOyXFxXb1_0(.din(w_dff_B_yBE6hfya7_0),.dout(w_dff_B_QOyXFxXb1_0),.clk(gclk));
	jdff dff_B_FTiyY0mW7_0(.din(w_dff_B_QOyXFxXb1_0),.dout(w_dff_B_FTiyY0mW7_0),.clk(gclk));
	jdff dff_B_MdmJGBM98_0(.din(w_dff_B_FTiyY0mW7_0),.dout(w_dff_B_MdmJGBM98_0),.clk(gclk));
	jdff dff_B_l53WllE26_1(.din(n1790),.dout(w_dff_B_l53WllE26_1),.clk(gclk));
	jdff dff_B_vSbNmNzd5_1(.din(w_dff_B_l53WllE26_1),.dout(w_dff_B_vSbNmNzd5_1),.clk(gclk));
	jdff dff_B_Mg9kBZZz1_1(.din(w_dff_B_vSbNmNzd5_1),.dout(w_dff_B_Mg9kBZZz1_1),.clk(gclk));
	jdff dff_B_LiTXwJ6Q6_1(.din(w_dff_B_Mg9kBZZz1_1),.dout(w_dff_B_LiTXwJ6Q6_1),.clk(gclk));
	jdff dff_B_PS8G7aWC1_1(.din(w_dff_B_LiTXwJ6Q6_1),.dout(w_dff_B_PS8G7aWC1_1),.clk(gclk));
	jdff dff_B_GZDCKJP06_1(.din(w_dff_B_PS8G7aWC1_1),.dout(w_dff_B_GZDCKJP06_1),.clk(gclk));
	jdff dff_B_HNn22smk6_1(.din(w_dff_B_GZDCKJP06_1),.dout(w_dff_B_HNn22smk6_1),.clk(gclk));
	jdff dff_B_pr6TljLb6_1(.din(w_dff_B_HNn22smk6_1),.dout(w_dff_B_pr6TljLb6_1),.clk(gclk));
	jdff dff_B_5idRKmw72_1(.din(w_dff_B_pr6TljLb6_1),.dout(w_dff_B_5idRKmw72_1),.clk(gclk));
	jdff dff_B_rc0gTyTh5_1(.din(w_dff_B_5idRKmw72_1),.dout(w_dff_B_rc0gTyTh5_1),.clk(gclk));
	jdff dff_B_tjpf42O52_1(.din(w_dff_B_rc0gTyTh5_1),.dout(w_dff_B_tjpf42O52_1),.clk(gclk));
	jdff dff_B_yk1vio3G0_1(.din(w_dff_B_tjpf42O52_1),.dout(w_dff_B_yk1vio3G0_1),.clk(gclk));
	jdff dff_B_rfh8Azrx4_1(.din(w_dff_B_yk1vio3G0_1),.dout(w_dff_B_rfh8Azrx4_1),.clk(gclk));
	jdff dff_B_DsiobYQn1_0(.din(n1791),.dout(w_dff_B_DsiobYQn1_0),.clk(gclk));
	jdff dff_B_YFdZIHOs6_0(.din(w_dff_B_DsiobYQn1_0),.dout(w_dff_B_YFdZIHOs6_0),.clk(gclk));
	jdff dff_B_Zz9muBOd2_0(.din(w_dff_B_YFdZIHOs6_0),.dout(w_dff_B_Zz9muBOd2_0),.clk(gclk));
	jdff dff_B_4VYOsYnj6_0(.din(w_dff_B_Zz9muBOd2_0),.dout(w_dff_B_4VYOsYnj6_0),.clk(gclk));
	jdff dff_B_xaGkl7932_0(.din(w_dff_B_4VYOsYnj6_0),.dout(w_dff_B_xaGkl7932_0),.clk(gclk));
	jdff dff_B_ASUAg8o84_0(.din(w_dff_B_xaGkl7932_0),.dout(w_dff_B_ASUAg8o84_0),.clk(gclk));
	jdff dff_B_HbqTf5TA5_0(.din(w_dff_B_ASUAg8o84_0),.dout(w_dff_B_HbqTf5TA5_0),.clk(gclk));
	jdff dff_B_MnRayzoh5_0(.din(w_dff_B_HbqTf5TA5_0),.dout(w_dff_B_MnRayzoh5_0),.clk(gclk));
	jdff dff_B_8EJkcAz10_0(.din(w_dff_B_MnRayzoh5_0),.dout(w_dff_B_8EJkcAz10_0),.clk(gclk));
	jdff dff_B_pWrvYSR92_0(.din(w_dff_B_8EJkcAz10_0),.dout(w_dff_B_pWrvYSR92_0),.clk(gclk));
	jdff dff_B_LaxHBH1F4_0(.din(w_dff_B_pWrvYSR92_0),.dout(w_dff_B_LaxHBH1F4_0),.clk(gclk));
	jdff dff_B_zeHvFZoO8_0(.din(w_dff_B_LaxHBH1F4_0),.dout(w_dff_B_zeHvFZoO8_0),.clk(gclk));
	jdff dff_B_4rUrdJut2_1(.din(n1764),.dout(w_dff_B_4rUrdJut2_1),.clk(gclk));
	jdff dff_B_lSHDL41o8_1(.din(w_dff_B_4rUrdJut2_1),.dout(w_dff_B_lSHDL41o8_1),.clk(gclk));
	jdff dff_B_QVMOXoxm0_1(.din(w_dff_B_lSHDL41o8_1),.dout(w_dff_B_QVMOXoxm0_1),.clk(gclk));
	jdff dff_B_wlaFYO1W2_1(.din(w_dff_B_QVMOXoxm0_1),.dout(w_dff_B_wlaFYO1W2_1),.clk(gclk));
	jdff dff_B_lLOn836r2_1(.din(w_dff_B_wlaFYO1W2_1),.dout(w_dff_B_lLOn836r2_1),.clk(gclk));
	jdff dff_B_i8CPTuLt7_1(.din(w_dff_B_lLOn836r2_1),.dout(w_dff_B_i8CPTuLt7_1),.clk(gclk));
	jdff dff_B_mNepDa3v0_1(.din(w_dff_B_i8CPTuLt7_1),.dout(w_dff_B_mNepDa3v0_1),.clk(gclk));
	jdff dff_B_S3zaJXXc4_1(.din(w_dff_B_mNepDa3v0_1),.dout(w_dff_B_S3zaJXXc4_1),.clk(gclk));
	jdff dff_B_Kv8ad9017_1(.din(w_dff_B_S3zaJXXc4_1),.dout(w_dff_B_Kv8ad9017_1),.clk(gclk));
	jdff dff_B_u6KVBQwU1_1(.din(w_dff_B_Kv8ad9017_1),.dout(w_dff_B_u6KVBQwU1_1),.clk(gclk));
	jdff dff_B_ikSOyS6r2_1(.din(w_dff_B_u6KVBQwU1_1),.dout(w_dff_B_ikSOyS6r2_1),.clk(gclk));
	jdff dff_B_Ywy5LDQw3_1(.din(w_dff_B_ikSOyS6r2_1),.dout(w_dff_B_Ywy5LDQw3_1),.clk(gclk));
	jdff dff_B_cJe6CABx7_1(.din(w_dff_B_Ywy5LDQw3_1),.dout(w_dff_B_cJe6CABx7_1),.clk(gclk));
	jdff dff_B_uxFLB0it2_0(.din(n1765),.dout(w_dff_B_uxFLB0it2_0),.clk(gclk));
	jdff dff_B_j6bHU2QJ2_0(.din(w_dff_B_uxFLB0it2_0),.dout(w_dff_B_j6bHU2QJ2_0),.clk(gclk));
	jdff dff_B_RngWOTVA7_0(.din(w_dff_B_j6bHU2QJ2_0),.dout(w_dff_B_RngWOTVA7_0),.clk(gclk));
	jdff dff_B_CnngvG7H5_0(.din(w_dff_B_RngWOTVA7_0),.dout(w_dff_B_CnngvG7H5_0),.clk(gclk));
	jdff dff_B_CKE3EUF77_0(.din(w_dff_B_CnngvG7H5_0),.dout(w_dff_B_CKE3EUF77_0),.clk(gclk));
	jdff dff_B_55bo053C8_0(.din(w_dff_B_CKE3EUF77_0),.dout(w_dff_B_55bo053C8_0),.clk(gclk));
	jdff dff_B_AhNbvZ8F3_0(.din(w_dff_B_55bo053C8_0),.dout(w_dff_B_AhNbvZ8F3_0),.clk(gclk));
	jdff dff_B_l6tCg6yp8_0(.din(w_dff_B_AhNbvZ8F3_0),.dout(w_dff_B_l6tCg6yp8_0),.clk(gclk));
	jdff dff_B_dFb3QVSD8_0(.din(w_dff_B_l6tCg6yp8_0),.dout(w_dff_B_dFb3QVSD8_0),.clk(gclk));
	jdff dff_B_uPqkqIb35_0(.din(w_dff_B_dFb3QVSD8_0),.dout(w_dff_B_uPqkqIb35_0),.clk(gclk));
	jdff dff_B_q6KGRDOl4_0(.din(w_dff_B_uPqkqIb35_0),.dout(w_dff_B_q6KGRDOl4_0),.clk(gclk));
	jdff dff_B_mlOdPv2S6_0(.din(w_dff_B_q6KGRDOl4_0),.dout(w_dff_B_mlOdPv2S6_0),.clk(gclk));
	jdff dff_B_xQCfkq6P2_1(.din(n1731),.dout(w_dff_B_xQCfkq6P2_1),.clk(gclk));
	jdff dff_B_Gd4kUgaV9_1(.din(w_dff_B_xQCfkq6P2_1),.dout(w_dff_B_Gd4kUgaV9_1),.clk(gclk));
	jdff dff_B_JjlNcBPv4_1(.din(w_dff_B_Gd4kUgaV9_1),.dout(w_dff_B_JjlNcBPv4_1),.clk(gclk));
	jdff dff_B_bnx65bnW8_1(.din(w_dff_B_JjlNcBPv4_1),.dout(w_dff_B_bnx65bnW8_1),.clk(gclk));
	jdff dff_B_wPSp4Poz7_1(.din(w_dff_B_bnx65bnW8_1),.dout(w_dff_B_wPSp4Poz7_1),.clk(gclk));
	jdff dff_B_2l9hHGLC4_1(.din(w_dff_B_wPSp4Poz7_1),.dout(w_dff_B_2l9hHGLC4_1),.clk(gclk));
	jdff dff_B_k59GZeqv6_1(.din(w_dff_B_2l9hHGLC4_1),.dout(w_dff_B_k59GZeqv6_1),.clk(gclk));
	jdff dff_B_6dnsRt8p2_1(.din(w_dff_B_k59GZeqv6_1),.dout(w_dff_B_6dnsRt8p2_1),.clk(gclk));
	jdff dff_B_CXNy6fxz4_1(.din(w_dff_B_6dnsRt8p2_1),.dout(w_dff_B_CXNy6fxz4_1),.clk(gclk));
	jdff dff_B_ecas7eyI4_1(.din(w_dff_B_CXNy6fxz4_1),.dout(w_dff_B_ecas7eyI4_1),.clk(gclk));
	jdff dff_B_PiU4xhR46_1(.din(w_dff_B_ecas7eyI4_1),.dout(w_dff_B_PiU4xhR46_1),.clk(gclk));
	jdff dff_B_SjMI8q2N3_1(.din(w_dff_B_PiU4xhR46_1),.dout(w_dff_B_SjMI8q2N3_1),.clk(gclk));
	jdff dff_B_IZ4uEvw22_1(.din(w_dff_B_SjMI8q2N3_1),.dout(w_dff_B_IZ4uEvw22_1),.clk(gclk));
	jdff dff_B_yOdNxUpG8_0(.din(n1732),.dout(w_dff_B_yOdNxUpG8_0),.clk(gclk));
	jdff dff_B_Ppaiyd0W7_0(.din(w_dff_B_yOdNxUpG8_0),.dout(w_dff_B_Ppaiyd0W7_0),.clk(gclk));
	jdff dff_B_IIittGiD5_0(.din(w_dff_B_Ppaiyd0W7_0),.dout(w_dff_B_IIittGiD5_0),.clk(gclk));
	jdff dff_B_RtQgXSsh1_0(.din(w_dff_B_IIittGiD5_0),.dout(w_dff_B_RtQgXSsh1_0),.clk(gclk));
	jdff dff_B_PciOO2LB1_0(.din(w_dff_B_RtQgXSsh1_0),.dout(w_dff_B_PciOO2LB1_0),.clk(gclk));
	jdff dff_B_XsEugE3H9_0(.din(w_dff_B_PciOO2LB1_0),.dout(w_dff_B_XsEugE3H9_0),.clk(gclk));
	jdff dff_B_u1aeVSYb5_0(.din(w_dff_B_XsEugE3H9_0),.dout(w_dff_B_u1aeVSYb5_0),.clk(gclk));
	jdff dff_B_Gz3MZsGO2_0(.din(w_dff_B_u1aeVSYb5_0),.dout(w_dff_B_Gz3MZsGO2_0),.clk(gclk));
	jdff dff_B_GCobDsPT1_0(.din(w_dff_B_Gz3MZsGO2_0),.dout(w_dff_B_GCobDsPT1_0),.clk(gclk));
	jdff dff_B_jSkAOPfq3_0(.din(w_dff_B_GCobDsPT1_0),.dout(w_dff_B_jSkAOPfq3_0),.clk(gclk));
	jdff dff_B_Am9jWcao0_0(.din(w_dff_B_jSkAOPfq3_0),.dout(w_dff_B_Am9jWcao0_0),.clk(gclk));
	jdff dff_B_H4gx2No93_0(.din(w_dff_B_Am9jWcao0_0),.dout(w_dff_B_H4gx2No93_0),.clk(gclk));
	jdff dff_B_XS0v6Yt94_1(.din(n1691),.dout(w_dff_B_XS0v6Yt94_1),.clk(gclk));
	jdff dff_B_GzJukZws6_1(.din(w_dff_B_XS0v6Yt94_1),.dout(w_dff_B_GzJukZws6_1),.clk(gclk));
	jdff dff_B_SKcAnUJJ3_1(.din(w_dff_B_GzJukZws6_1),.dout(w_dff_B_SKcAnUJJ3_1),.clk(gclk));
	jdff dff_B_nm6Woswp3_1(.din(w_dff_B_SKcAnUJJ3_1),.dout(w_dff_B_nm6Woswp3_1),.clk(gclk));
	jdff dff_B_IJgyw2lz5_1(.din(w_dff_B_nm6Woswp3_1),.dout(w_dff_B_IJgyw2lz5_1),.clk(gclk));
	jdff dff_B_z14zVm0B2_1(.din(w_dff_B_IJgyw2lz5_1),.dout(w_dff_B_z14zVm0B2_1),.clk(gclk));
	jdff dff_B_M8MFXSHL3_1(.din(w_dff_B_z14zVm0B2_1),.dout(w_dff_B_M8MFXSHL3_1),.clk(gclk));
	jdff dff_B_SdVSy13N0_1(.din(w_dff_B_M8MFXSHL3_1),.dout(w_dff_B_SdVSy13N0_1),.clk(gclk));
	jdff dff_B_AjupddhC6_1(.din(w_dff_B_SdVSy13N0_1),.dout(w_dff_B_AjupddhC6_1),.clk(gclk));
	jdff dff_B_sCIEwXn17_1(.din(w_dff_B_AjupddhC6_1),.dout(w_dff_B_sCIEwXn17_1),.clk(gclk));
	jdff dff_B_qadIgar63_1(.din(w_dff_B_sCIEwXn17_1),.dout(w_dff_B_qadIgar63_1),.clk(gclk));
	jdff dff_B_hrXwnM7u2_1(.din(w_dff_B_qadIgar63_1),.dout(w_dff_B_hrXwnM7u2_1),.clk(gclk));
	jdff dff_B_FLzv5IFQ9_1(.din(w_dff_B_hrXwnM7u2_1),.dout(w_dff_B_FLzv5IFQ9_1),.clk(gclk));
	jdff dff_B_AgH5C2HU5_0(.din(n1692),.dout(w_dff_B_AgH5C2HU5_0),.clk(gclk));
	jdff dff_B_VSK6eRX65_0(.din(w_dff_B_AgH5C2HU5_0),.dout(w_dff_B_VSK6eRX65_0),.clk(gclk));
	jdff dff_B_PqqA8cXq1_0(.din(w_dff_B_VSK6eRX65_0),.dout(w_dff_B_PqqA8cXq1_0),.clk(gclk));
	jdff dff_B_SxAIVMtE8_0(.din(w_dff_B_PqqA8cXq1_0),.dout(w_dff_B_SxAIVMtE8_0),.clk(gclk));
	jdff dff_B_ZkV6EUFj9_0(.din(w_dff_B_SxAIVMtE8_0),.dout(w_dff_B_ZkV6EUFj9_0),.clk(gclk));
	jdff dff_B_dAL4109h5_0(.din(w_dff_B_ZkV6EUFj9_0),.dout(w_dff_B_dAL4109h5_0),.clk(gclk));
	jdff dff_B_emvDU7qz9_0(.din(w_dff_B_dAL4109h5_0),.dout(w_dff_B_emvDU7qz9_0),.clk(gclk));
	jdff dff_B_Ci4zxg9i2_0(.din(w_dff_B_emvDU7qz9_0),.dout(w_dff_B_Ci4zxg9i2_0),.clk(gclk));
	jdff dff_B_NGl4n9je9_0(.din(w_dff_B_Ci4zxg9i2_0),.dout(w_dff_B_NGl4n9je9_0),.clk(gclk));
	jdff dff_B_49MfWjRv3_0(.din(w_dff_B_NGl4n9je9_0),.dout(w_dff_B_49MfWjRv3_0),.clk(gclk));
	jdff dff_B_XtoT0os52_0(.din(w_dff_B_49MfWjRv3_0),.dout(w_dff_B_XtoT0os52_0),.clk(gclk));
	jdff dff_B_JYhckuGj9_1(.din(n1643),.dout(w_dff_B_JYhckuGj9_1),.clk(gclk));
	jdff dff_B_gNJ52H7k6_1(.din(w_dff_B_JYhckuGj9_1),.dout(w_dff_B_gNJ52H7k6_1),.clk(gclk));
	jdff dff_B_QXGLSJiU0_1(.din(w_dff_B_gNJ52H7k6_1),.dout(w_dff_B_QXGLSJiU0_1),.clk(gclk));
	jdff dff_B_bmazQtKw7_1(.din(w_dff_B_QXGLSJiU0_1),.dout(w_dff_B_bmazQtKw7_1),.clk(gclk));
	jdff dff_B_fvfPc0Y45_1(.din(w_dff_B_bmazQtKw7_1),.dout(w_dff_B_fvfPc0Y45_1),.clk(gclk));
	jdff dff_B_rjErD65m3_1(.din(w_dff_B_fvfPc0Y45_1),.dout(w_dff_B_rjErD65m3_1),.clk(gclk));
	jdff dff_B_8C34pXR15_1(.din(w_dff_B_rjErD65m3_1),.dout(w_dff_B_8C34pXR15_1),.clk(gclk));
	jdff dff_B_60U9NIXZ2_1(.din(w_dff_B_8C34pXR15_1),.dout(w_dff_B_60U9NIXZ2_1),.clk(gclk));
	jdff dff_B_H8AGPWpd5_1(.din(w_dff_B_60U9NIXZ2_1),.dout(w_dff_B_H8AGPWpd5_1),.clk(gclk));
	jdff dff_B_IvcX5JtQ3_1(.din(w_dff_B_H8AGPWpd5_1),.dout(w_dff_B_IvcX5JtQ3_1),.clk(gclk));
	jdff dff_B_ULhVCJZl1_1(.din(w_dff_B_IvcX5JtQ3_1),.dout(w_dff_B_ULhVCJZl1_1),.clk(gclk));
	jdff dff_B_eDg4Wggn8_1(.din(w_dff_B_ULhVCJZl1_1),.dout(w_dff_B_eDg4Wggn8_1),.clk(gclk));
	jdff dff_B_i2yFD3pf6_0(.din(n1644),.dout(w_dff_B_i2yFD3pf6_0),.clk(gclk));
	jdff dff_B_7bztS9jn8_0(.din(w_dff_B_i2yFD3pf6_0),.dout(w_dff_B_7bztS9jn8_0),.clk(gclk));
	jdff dff_B_s0XxKT3p5_0(.din(w_dff_B_7bztS9jn8_0),.dout(w_dff_B_s0XxKT3p5_0),.clk(gclk));
	jdff dff_B_Jx8nqwLq8_0(.din(w_dff_B_s0XxKT3p5_0),.dout(w_dff_B_Jx8nqwLq8_0),.clk(gclk));
	jdff dff_B_mMJxiULn5_0(.din(w_dff_B_Jx8nqwLq8_0),.dout(w_dff_B_mMJxiULn5_0),.clk(gclk));
	jdff dff_B_XSrf3GsQ8_0(.din(w_dff_B_mMJxiULn5_0),.dout(w_dff_B_XSrf3GsQ8_0),.clk(gclk));
	jdff dff_B_LUQpthNW2_0(.din(w_dff_B_XSrf3GsQ8_0),.dout(w_dff_B_LUQpthNW2_0),.clk(gclk));
	jdff dff_B_fE3mV4bG3_0(.din(w_dff_B_LUQpthNW2_0),.dout(w_dff_B_fE3mV4bG3_0),.clk(gclk));
	jdff dff_B_NyfWoSAF9_0(.din(w_dff_B_fE3mV4bG3_0),.dout(w_dff_B_NyfWoSAF9_0),.clk(gclk));
	jdff dff_B_17qFCh4f9_0(.din(w_dff_B_NyfWoSAF9_0),.dout(w_dff_B_17qFCh4f9_0),.clk(gclk));
	jdff dff_B_ho1dLcXQ7_1(.din(n1588),.dout(w_dff_B_ho1dLcXQ7_1),.clk(gclk));
	jdff dff_B_MW0GOehu6_1(.din(w_dff_B_ho1dLcXQ7_1),.dout(w_dff_B_MW0GOehu6_1),.clk(gclk));
	jdff dff_B_d3imbFOs7_1(.din(w_dff_B_MW0GOehu6_1),.dout(w_dff_B_d3imbFOs7_1),.clk(gclk));
	jdff dff_B_DaYm668r7_1(.din(w_dff_B_d3imbFOs7_1),.dout(w_dff_B_DaYm668r7_1),.clk(gclk));
	jdff dff_B_E99CDv9F1_1(.din(w_dff_B_DaYm668r7_1),.dout(w_dff_B_E99CDv9F1_1),.clk(gclk));
	jdff dff_B_5YzPwp3N2_1(.din(w_dff_B_E99CDv9F1_1),.dout(w_dff_B_5YzPwp3N2_1),.clk(gclk));
	jdff dff_B_UBvpm76y9_1(.din(w_dff_B_5YzPwp3N2_1),.dout(w_dff_B_UBvpm76y9_1),.clk(gclk));
	jdff dff_B_OB4agIAn7_1(.din(w_dff_B_UBvpm76y9_1),.dout(w_dff_B_OB4agIAn7_1),.clk(gclk));
	jdff dff_B_lEQH5B4y9_1(.din(w_dff_B_OB4agIAn7_1),.dout(w_dff_B_lEQH5B4y9_1),.clk(gclk));
	jdff dff_B_PekFeIzl8_1(.din(w_dff_B_lEQH5B4y9_1),.dout(w_dff_B_PekFeIzl8_1),.clk(gclk));
	jdff dff_B_ROPNhEJH1_0(.din(n1589),.dout(w_dff_B_ROPNhEJH1_0),.clk(gclk));
	jdff dff_B_v4FDHYhU7_0(.din(w_dff_B_ROPNhEJH1_0),.dout(w_dff_B_v4FDHYhU7_0),.clk(gclk));
	jdff dff_B_N9lZE66c9_0(.din(w_dff_B_v4FDHYhU7_0),.dout(w_dff_B_N9lZE66c9_0),.clk(gclk));
	jdff dff_B_MlYzs8A12_0(.din(w_dff_B_N9lZE66c9_0),.dout(w_dff_B_MlYzs8A12_0),.clk(gclk));
	jdff dff_B_ot9XZPI12_0(.din(w_dff_B_MlYzs8A12_0),.dout(w_dff_B_ot9XZPI12_0),.clk(gclk));
	jdff dff_B_f32xVb5V9_0(.din(w_dff_B_ot9XZPI12_0),.dout(w_dff_B_f32xVb5V9_0),.clk(gclk));
	jdff dff_B_7d48Z0JU4_0(.din(w_dff_B_f32xVb5V9_0),.dout(w_dff_B_7d48Z0JU4_0),.clk(gclk));
	jdff dff_B_BRq9R90W5_0(.din(w_dff_B_7d48Z0JU4_0),.dout(w_dff_B_BRq9R90W5_0),.clk(gclk));
	jdff dff_B_0MOqRX8r1_1(.din(n1526),.dout(w_dff_B_0MOqRX8r1_1),.clk(gclk));
	jdff dff_B_X3n6zlmJ0_1(.din(w_dff_B_0MOqRX8r1_1),.dout(w_dff_B_X3n6zlmJ0_1),.clk(gclk));
	jdff dff_B_LHaoAXLB5_1(.din(w_dff_B_X3n6zlmJ0_1),.dout(w_dff_B_LHaoAXLB5_1),.clk(gclk));
	jdff dff_B_Pi3L4iFl2_1(.din(w_dff_B_LHaoAXLB5_1),.dout(w_dff_B_Pi3L4iFl2_1),.clk(gclk));
	jdff dff_B_u4MGejJa1_1(.din(w_dff_B_Pi3L4iFl2_1),.dout(w_dff_B_u4MGejJa1_1),.clk(gclk));
	jdff dff_B_EmbF5t6s7_1(.din(w_dff_B_u4MGejJa1_1),.dout(w_dff_B_EmbF5t6s7_1),.clk(gclk));
	jdff dff_B_6zS7mczk2_1(.din(w_dff_B_EmbF5t6s7_1),.dout(w_dff_B_6zS7mczk2_1),.clk(gclk));
	jdff dff_B_6XWUy8nb8_1(.din(w_dff_B_6zS7mczk2_1),.dout(w_dff_B_6XWUy8nb8_1),.clk(gclk));
	jdff dff_B_4zhX4x6F4_0(.din(n1527),.dout(w_dff_B_4zhX4x6F4_0),.clk(gclk));
	jdff dff_B_M4jVcfQi7_0(.din(w_dff_B_4zhX4x6F4_0),.dout(w_dff_B_M4jVcfQi7_0),.clk(gclk));
	jdff dff_B_PTz5t4lN2_0(.din(w_dff_B_M4jVcfQi7_0),.dout(w_dff_B_PTz5t4lN2_0),.clk(gclk));
	jdff dff_B_MS37GiVH4_0(.din(w_dff_B_PTz5t4lN2_0),.dout(w_dff_B_MS37GiVH4_0),.clk(gclk));
	jdff dff_B_GptzSQq79_0(.din(w_dff_B_MS37GiVH4_0),.dout(w_dff_B_GptzSQq79_0),.clk(gclk));
	jdff dff_B_tPp8Fugc9_0(.din(w_dff_B_GptzSQq79_0),.dout(w_dff_B_tPp8Fugc9_0),.clk(gclk));
	jdff dff_B_KllwmgZA0_1(.din(n1457),.dout(w_dff_B_KllwmgZA0_1),.clk(gclk));
	jdff dff_B_dw11LbjA5_1(.din(w_dff_B_KllwmgZA0_1),.dout(w_dff_B_dw11LbjA5_1),.clk(gclk));
	jdff dff_B_plwNbacf8_1(.din(w_dff_B_dw11LbjA5_1),.dout(w_dff_B_plwNbacf8_1),.clk(gclk));
	jdff dff_B_onyABVuW4_1(.din(w_dff_B_plwNbacf8_1),.dout(w_dff_B_onyABVuW4_1),.clk(gclk));
	jdff dff_B_mmNgvumf7_1(.din(w_dff_B_onyABVuW4_1),.dout(w_dff_B_mmNgvumf7_1),.clk(gclk));
	jdff dff_B_2zYF6yEk2_1(.din(w_dff_B_mmNgvumf7_1),.dout(w_dff_B_2zYF6yEk2_1),.clk(gclk));
	jdff dff_B_S72RrKdf6_1(.din(w_dff_B_2zYF6yEk2_1),.dout(w_dff_B_S72RrKdf6_1),.clk(gclk));
	jdff dff_B_bjDJvoz76_0(.din(n1458),.dout(w_dff_B_bjDJvoz76_0),.clk(gclk));
	jdff dff_B_1NnApfbK3_0(.din(w_dff_B_bjDJvoz76_0),.dout(w_dff_B_1NnApfbK3_0),.clk(gclk));
	jdff dff_B_Mz8I7oQ63_0(.din(w_dff_B_1NnApfbK3_0),.dout(w_dff_B_Mz8I7oQ63_0),.clk(gclk));
	jdff dff_B_kJ3TBsQJ6_0(.din(w_dff_B_Mz8I7oQ63_0),.dout(w_dff_B_kJ3TBsQJ6_0),.clk(gclk));
	jdff dff_B_K8aNhHto4_0(.din(w_dff_B_kJ3TBsQJ6_0),.dout(w_dff_B_K8aNhHto4_0),.clk(gclk));
	jdff dff_B_ZX58KJb36_1(.din(n1381),.dout(w_dff_B_ZX58KJb36_1),.clk(gclk));
	jdff dff_B_dmSDmjq87_1(.din(w_dff_B_ZX58KJb36_1),.dout(w_dff_B_dmSDmjq87_1),.clk(gclk));
	jdff dff_B_m4Ci5srJ3_1(.din(w_dff_B_dmSDmjq87_1),.dout(w_dff_B_m4Ci5srJ3_1),.clk(gclk));
	jdff dff_B_iyEaSrZ16_1(.din(w_dff_B_m4Ci5srJ3_1),.dout(w_dff_B_iyEaSrZ16_1),.clk(gclk));
	jdff dff_B_DQMvCcBh2_1(.din(w_dff_B_iyEaSrZ16_1),.dout(w_dff_B_DQMvCcBh2_1),.clk(gclk));
	jdff dff_B_qh4TqmUH5_1(.din(w_dff_B_DQMvCcBh2_1),.dout(w_dff_B_qh4TqmUH5_1),.clk(gclk));
	jdff dff_B_s5EEVjOx9_0(.din(n1382),.dout(w_dff_B_s5EEVjOx9_0),.clk(gclk));
	jdff dff_B_Lu1u8W6E1_0(.din(w_dff_B_s5EEVjOx9_0),.dout(w_dff_B_Lu1u8W6E1_0),.clk(gclk));
	jdff dff_B_GwmRwY362_0(.din(w_dff_B_Lu1u8W6E1_0),.dout(w_dff_B_GwmRwY362_0),.clk(gclk));
	jdff dff_B_d05Jrrm95_0(.din(w_dff_B_GwmRwY362_0),.dout(w_dff_B_d05Jrrm95_0),.clk(gclk));
	jdff dff_B_i07KIMW05_1(.din(n1299),.dout(w_dff_B_i07KIMW05_1),.clk(gclk));
	jdff dff_B_lDvUvXFE5_1(.din(w_dff_B_i07KIMW05_1),.dout(w_dff_B_lDvUvXFE5_1),.clk(gclk));
	jdff dff_B_vtqfyuMu0_1(.din(w_dff_B_lDvUvXFE5_1),.dout(w_dff_B_vtqfyuMu0_1),.clk(gclk));
	jdff dff_B_AmhI8UHA1_1(.din(n1211),.dout(w_dff_B_AmhI8UHA1_1),.clk(gclk));
	jdff dff_B_nlpNDxfO7_1(.din(n1113),.dout(w_dff_B_nlpNDxfO7_1),.clk(gclk));
	jdff dff_A_ldyRm5Sp4_1(.dout(w_n1013_0[1]),.din(w_dff_A_ldyRm5Sp4_1),.clk(gclk));
	jdff dff_B_eoyEvq7x2_2(.din(n1011),.dout(w_dff_B_eoyEvq7x2_2),.clk(gclk));
	jdff dff_B_tUJC509k0_1(.din(n908),.dout(w_dff_B_tUJC509k0_1),.clk(gclk));
	jdff dff_B_pDRcoDZO2_1(.din(n808),.dout(w_dff_B_pDRcoDZO2_1),.clk(gclk));
	jdff dff_B_LszaTL6P4_1(.din(n709),.dout(w_dff_B_LszaTL6P4_1),.clk(gclk));
	jdff dff_B_sHrr4wRB8_1(.din(n617),.dout(w_dff_B_sHrr4wRB8_1),.clk(gclk));
	jdff dff_B_W13ktaNM2_1(.din(n532),.dout(w_dff_B_W13ktaNM2_1),.clk(gclk));
	jdff dff_B_tzl0zDuC0_1(.din(n454),.dout(w_dff_B_tzl0zDuC0_1),.clk(gclk));
	jdff dff_B_8cIcvORO0_1(.din(n383),.dout(w_dff_B_8cIcvORO0_1),.clk(gclk));
	jdff dff_B_x30379n46_1(.din(n320),.dout(w_dff_B_x30379n46_1),.clk(gclk));
	jdff dff_B_ZDi3jBiT2_1(.din(n264),.dout(w_dff_B_ZDi3jBiT2_1),.clk(gclk));
	jdff dff_B_SFCaJsrj1_1(.din(n215),.dout(w_dff_B_SFCaJsrj1_1),.clk(gclk));
	jdff dff_B_WOBZxwkd3_1(.din(n173),.dout(w_dff_B_WOBZxwkd3_1),.clk(gclk));
	jdff dff_B_GrrYRaG21_1(.din(n138),.dout(w_dff_B_GrrYRaG21_1),.clk(gclk));
	jdff dff_B_zyUCrIaE8_1(.din(n109),.dout(w_dff_B_zyUCrIaE8_1),.clk(gclk));
	jdff dff_B_hKWuVKxP1_1(.din(n88),.dout(w_dff_B_hKWuVKxP1_1),.clk(gclk));
	jdff dff_B_0KNpzkH01_2(.din(n67),.dout(w_dff_B_0KNpzkH01_2),.clk(gclk));
	jdff dff_A_WP9bZbhQ6_0(.dout(w_n66_0[0]),.din(w_dff_A_WP9bZbhQ6_0),.clk(gclk));
	jdff dff_A_19rWTS8w4_0(.dout(w_dff_A_WP9bZbhQ6_0),.din(w_dff_A_19rWTS8w4_0),.clk(gclk));
	jdff dff_A_vQBAJatK4_1(.dout(w_dff_A_yDJmqpSx8_0),.din(w_dff_A_vQBAJatK4_1),.clk(gclk));
	jdff dff_A_yDJmqpSx8_0(.dout(w_dff_A_lZwFM8ZI5_0),.din(w_dff_A_yDJmqpSx8_0),.clk(gclk));
	jdff dff_A_lZwFM8ZI5_0(.dout(w_dff_A_pAecoUmY2_0),.din(w_dff_A_lZwFM8ZI5_0),.clk(gclk));
	jdff dff_A_pAecoUmY2_0(.dout(w_dff_A_uFXjBaex1_0),.din(w_dff_A_pAecoUmY2_0),.clk(gclk));
	jdff dff_A_uFXjBaex1_0(.dout(w_dff_A_PmFQJxZU4_0),.din(w_dff_A_uFXjBaex1_0),.clk(gclk));
	jdff dff_A_PmFQJxZU4_0(.dout(w_dff_A_7516o1Wj1_0),.din(w_dff_A_PmFQJxZU4_0),.clk(gclk));
	jdff dff_A_7516o1Wj1_0(.dout(w_dff_A_QR0VUwJA8_0),.din(w_dff_A_7516o1Wj1_0),.clk(gclk));
	jdff dff_A_QR0VUwJA8_0(.dout(w_dff_A_GmH6zCB17_0),.din(w_dff_A_QR0VUwJA8_0),.clk(gclk));
	jdff dff_A_GmH6zCB17_0(.dout(w_dff_A_U9nXheOp1_0),.din(w_dff_A_GmH6zCB17_0),.clk(gclk));
	jdff dff_A_U9nXheOp1_0(.dout(w_dff_A_B9BqP8PQ7_0),.din(w_dff_A_U9nXheOp1_0),.clk(gclk));
	jdff dff_A_B9BqP8PQ7_0(.dout(w_dff_A_lNLF2BjB4_0),.din(w_dff_A_B9BqP8PQ7_0),.clk(gclk));
	jdff dff_A_lNLF2BjB4_0(.dout(w_dff_A_xR5oOP2r5_0),.din(w_dff_A_lNLF2BjB4_0),.clk(gclk));
	jdff dff_A_xR5oOP2r5_0(.dout(w_dff_A_EIvp8IWx3_0),.din(w_dff_A_xR5oOP2r5_0),.clk(gclk));
	jdff dff_A_EIvp8IWx3_0(.dout(w_dff_A_sL00PJx48_0),.din(w_dff_A_EIvp8IWx3_0),.clk(gclk));
	jdff dff_A_sL00PJx48_0(.dout(w_dff_A_sLW1frs88_0),.din(w_dff_A_sL00PJx48_0),.clk(gclk));
	jdff dff_A_sLW1frs88_0(.dout(w_dff_A_DGBD7lci8_0),.din(w_dff_A_sLW1frs88_0),.clk(gclk));
	jdff dff_A_DGBD7lci8_0(.dout(w_dff_A_3hII8bb82_0),.din(w_dff_A_DGBD7lci8_0),.clk(gclk));
	jdff dff_A_3hII8bb82_0(.dout(w_dff_A_lgYjaHiP5_0),.din(w_dff_A_3hII8bb82_0),.clk(gclk));
	jdff dff_A_lgYjaHiP5_0(.dout(w_dff_A_r3wG0ogX1_0),.din(w_dff_A_lgYjaHiP5_0),.clk(gclk));
	jdff dff_A_r3wG0ogX1_0(.dout(w_dff_A_2iu5bMul2_0),.din(w_dff_A_r3wG0ogX1_0),.clk(gclk));
	jdff dff_A_2iu5bMul2_0(.dout(w_dff_A_xLU5Epjw5_0),.din(w_dff_A_2iu5bMul2_0),.clk(gclk));
	jdff dff_A_xLU5Epjw5_0(.dout(w_dff_A_camGR4OS1_0),.din(w_dff_A_xLU5Epjw5_0),.clk(gclk));
	jdff dff_A_camGR4OS1_0(.dout(w_dff_A_8FjqrV9E6_0),.din(w_dff_A_camGR4OS1_0),.clk(gclk));
	jdff dff_A_8FjqrV9E6_0(.dout(w_dff_A_6xTW2Omh3_0),.din(w_dff_A_8FjqrV9E6_0),.clk(gclk));
	jdff dff_A_6xTW2Omh3_0(.dout(w_dff_A_JFAZPNSf9_0),.din(w_dff_A_6xTW2Omh3_0),.clk(gclk));
	jdff dff_A_JFAZPNSf9_0(.dout(w_dff_A_vJwNJk609_0),.din(w_dff_A_JFAZPNSf9_0),.clk(gclk));
	jdff dff_A_vJwNJk609_0(.dout(w_dff_A_f6xMlbQJ0_0),.din(w_dff_A_vJwNJk609_0),.clk(gclk));
	jdff dff_A_f6xMlbQJ0_0(.dout(w_dff_A_rGMPTwGp0_0),.din(w_dff_A_f6xMlbQJ0_0),.clk(gclk));
	jdff dff_A_rGMPTwGp0_0(.dout(w_dff_A_Yv3BvXIL8_0),.din(w_dff_A_rGMPTwGp0_0),.clk(gclk));
	jdff dff_A_Yv3BvXIL8_0(.dout(w_dff_A_fyMvgymV0_0),.din(w_dff_A_Yv3BvXIL8_0),.clk(gclk));
	jdff dff_A_fyMvgymV0_0(.dout(w_dff_A_XuL0PMOG8_0),.din(w_dff_A_fyMvgymV0_0),.clk(gclk));
	jdff dff_A_XuL0PMOG8_0(.dout(w_dff_A_DxWhPD141_0),.din(w_dff_A_XuL0PMOG8_0),.clk(gclk));
	jdff dff_A_DxWhPD141_0(.dout(w_dff_A_eEaul0dx2_0),.din(w_dff_A_DxWhPD141_0),.clk(gclk));
	jdff dff_A_eEaul0dx2_0(.dout(w_dff_A_lsqm5opx1_0),.din(w_dff_A_eEaul0dx2_0),.clk(gclk));
	jdff dff_A_lsqm5opx1_0(.dout(w_dff_A_FiPshPat6_0),.din(w_dff_A_lsqm5opx1_0),.clk(gclk));
	jdff dff_A_FiPshPat6_0(.dout(w_dff_A_B2Y1Nnml5_0),.din(w_dff_A_FiPshPat6_0),.clk(gclk));
	jdff dff_A_B2Y1Nnml5_0(.dout(w_dff_A_ln96ecSa5_0),.din(w_dff_A_B2Y1Nnml5_0),.clk(gclk));
	jdff dff_A_ln96ecSa5_0(.dout(w_dff_A_K8Uc8uO82_0),.din(w_dff_A_ln96ecSa5_0),.clk(gclk));
	jdff dff_A_K8Uc8uO82_0(.dout(w_dff_A_DnMtjMmI4_0),.din(w_dff_A_K8Uc8uO82_0),.clk(gclk));
	jdff dff_A_DnMtjMmI4_0(.dout(w_dff_A_tiJP9vMG7_0),.din(w_dff_A_DnMtjMmI4_0),.clk(gclk));
	jdff dff_A_tiJP9vMG7_0(.dout(w_dff_A_1EfO6lqI3_0),.din(w_dff_A_tiJP9vMG7_0),.clk(gclk));
	jdff dff_A_1EfO6lqI3_0(.dout(w_dff_A_sVOiuPDL6_0),.din(w_dff_A_1EfO6lqI3_0),.clk(gclk));
	jdff dff_A_sVOiuPDL6_0(.dout(w_dff_A_NkA4BtWt7_0),.din(w_dff_A_sVOiuPDL6_0),.clk(gclk));
	jdff dff_A_NkA4BtWt7_0(.dout(w_dff_A_hfstznWA8_0),.din(w_dff_A_NkA4BtWt7_0),.clk(gclk));
	jdff dff_A_hfstznWA8_0(.dout(w_dff_A_koaZlOGX7_0),.din(w_dff_A_hfstznWA8_0),.clk(gclk));
	jdff dff_A_koaZlOGX7_0(.dout(w_dff_A_bpV6me7t3_0),.din(w_dff_A_koaZlOGX7_0),.clk(gclk));
	jdff dff_A_bpV6me7t3_0(.dout(w_dff_A_9cqNnkby4_0),.din(w_dff_A_bpV6me7t3_0),.clk(gclk));
	jdff dff_A_9cqNnkby4_0(.dout(w_dff_A_iMfraidZ2_0),.din(w_dff_A_9cqNnkby4_0),.clk(gclk));
	jdff dff_A_iMfraidZ2_0(.dout(w_dff_A_L6oQ0NhD3_0),.din(w_dff_A_iMfraidZ2_0),.clk(gclk));
	jdff dff_A_L6oQ0NhD3_0(.dout(w_dff_A_zvK8RSH07_0),.din(w_dff_A_L6oQ0NhD3_0),.clk(gclk));
	jdff dff_A_zvK8RSH07_0(.dout(w_dff_A_VnkAfI5P8_0),.din(w_dff_A_zvK8RSH07_0),.clk(gclk));
	jdff dff_A_VnkAfI5P8_0(.dout(w_dff_A_uGrpNwGV6_0),.din(w_dff_A_VnkAfI5P8_0),.clk(gclk));
	jdff dff_A_uGrpNwGV6_0(.dout(w_dff_A_3ZRng7Ai9_0),.din(w_dff_A_uGrpNwGV6_0),.clk(gclk));
	jdff dff_A_3ZRng7Ai9_0(.dout(w_dff_A_MCUPLppW4_0),.din(w_dff_A_3ZRng7Ai9_0),.clk(gclk));
	jdff dff_A_MCUPLppW4_0(.dout(w_dff_A_S61Jc8zR9_0),.din(w_dff_A_MCUPLppW4_0),.clk(gclk));
	jdff dff_A_S61Jc8zR9_0(.dout(w_dff_A_v3rDdi969_0),.din(w_dff_A_S61Jc8zR9_0),.clk(gclk));
	jdff dff_A_v3rDdi969_0(.dout(w_dff_A_xv7cj5K92_0),.din(w_dff_A_v3rDdi969_0),.clk(gclk));
	jdff dff_A_xv7cj5K92_0(.dout(w_dff_A_cwufwjbf6_0),.din(w_dff_A_xv7cj5K92_0),.clk(gclk));
	jdff dff_A_cwufwjbf6_0(.dout(w_dff_A_URs5L4D35_0),.din(w_dff_A_cwufwjbf6_0),.clk(gclk));
	jdff dff_A_URs5L4D35_0(.dout(w_dff_A_EOt6XsKJ5_0),.din(w_dff_A_URs5L4D35_0),.clk(gclk));
	jdff dff_A_EOt6XsKJ5_0(.dout(w_dff_A_ykR8CTuG2_0),.din(w_dff_A_EOt6XsKJ5_0),.clk(gclk));
	jdff dff_A_ykR8CTuG2_0(.dout(w_dff_A_ubPgaL214_0),.din(w_dff_A_ykR8CTuG2_0),.clk(gclk));
	jdff dff_A_ubPgaL214_0(.dout(w_dff_A_axMy7jTL2_0),.din(w_dff_A_ubPgaL214_0),.clk(gclk));
	jdff dff_A_axMy7jTL2_0(.dout(w_dff_A_H5xRXzh26_0),.din(w_dff_A_axMy7jTL2_0),.clk(gclk));
	jdff dff_A_H5xRXzh26_0(.dout(w_dff_A_PA8UFdlJ0_0),.din(w_dff_A_H5xRXzh26_0),.clk(gclk));
	jdff dff_A_PA8UFdlJ0_0(.dout(w_dff_A_UJNeqzmU5_0),.din(w_dff_A_PA8UFdlJ0_0),.clk(gclk));
	jdff dff_A_UJNeqzmU5_0(.dout(w_dff_A_slxIVVxJ6_0),.din(w_dff_A_UJNeqzmU5_0),.clk(gclk));
	jdff dff_A_slxIVVxJ6_0(.dout(w_dff_A_Ghagossj9_0),.din(w_dff_A_slxIVVxJ6_0),.clk(gclk));
	jdff dff_A_Ghagossj9_0(.dout(w_dff_A_vEimH8TU6_0),.din(w_dff_A_Ghagossj9_0),.clk(gclk));
	jdff dff_A_vEimH8TU6_0(.dout(w_dff_A_jufft8eE0_0),.din(w_dff_A_vEimH8TU6_0),.clk(gclk));
	jdff dff_A_jufft8eE0_0(.dout(w_dff_A_1MWlUZeZ9_0),.din(w_dff_A_jufft8eE0_0),.clk(gclk));
	jdff dff_A_1MWlUZeZ9_0(.dout(w_dff_A_y5q29IMO0_0),.din(w_dff_A_1MWlUZeZ9_0),.clk(gclk));
	jdff dff_A_y5q29IMO0_0(.dout(w_dff_A_w5aNIRF70_0),.din(w_dff_A_y5q29IMO0_0),.clk(gclk));
	jdff dff_A_w5aNIRF70_0(.dout(G545gat),.din(w_dff_A_w5aNIRF70_0),.clk(gclk));
	jdff dff_A_HFwDfpPm3_2(.dout(w_dff_A_A4c8mjax2_0),.din(w_dff_A_HFwDfpPm3_2),.clk(gclk));
	jdff dff_A_A4c8mjax2_0(.dout(w_dff_A_Njle6QaC8_0),.din(w_dff_A_A4c8mjax2_0),.clk(gclk));
	jdff dff_A_Njle6QaC8_0(.dout(w_dff_A_8GhHAcWv0_0),.din(w_dff_A_Njle6QaC8_0),.clk(gclk));
	jdff dff_A_8GhHAcWv0_0(.dout(w_dff_A_FpePlT0U4_0),.din(w_dff_A_8GhHAcWv0_0),.clk(gclk));
	jdff dff_A_FpePlT0U4_0(.dout(w_dff_A_K3ANNQyf9_0),.din(w_dff_A_FpePlT0U4_0),.clk(gclk));
	jdff dff_A_K3ANNQyf9_0(.dout(w_dff_A_Qvg1yppC1_0),.din(w_dff_A_K3ANNQyf9_0),.clk(gclk));
	jdff dff_A_Qvg1yppC1_0(.dout(w_dff_A_3BucendH0_0),.din(w_dff_A_Qvg1yppC1_0),.clk(gclk));
	jdff dff_A_3BucendH0_0(.dout(w_dff_A_7nMFY3eT0_0),.din(w_dff_A_3BucendH0_0),.clk(gclk));
	jdff dff_A_7nMFY3eT0_0(.dout(w_dff_A_M8AfgK3h7_0),.din(w_dff_A_7nMFY3eT0_0),.clk(gclk));
	jdff dff_A_M8AfgK3h7_0(.dout(w_dff_A_Zu8ms7Rg8_0),.din(w_dff_A_M8AfgK3h7_0),.clk(gclk));
	jdff dff_A_Zu8ms7Rg8_0(.dout(w_dff_A_KvSSrMYO6_0),.din(w_dff_A_Zu8ms7Rg8_0),.clk(gclk));
	jdff dff_A_KvSSrMYO6_0(.dout(w_dff_A_ApJg33ru5_0),.din(w_dff_A_KvSSrMYO6_0),.clk(gclk));
	jdff dff_A_ApJg33ru5_0(.dout(w_dff_A_hZFaVF6y3_0),.din(w_dff_A_ApJg33ru5_0),.clk(gclk));
	jdff dff_A_hZFaVF6y3_0(.dout(w_dff_A_lOg3hT469_0),.din(w_dff_A_hZFaVF6y3_0),.clk(gclk));
	jdff dff_A_lOg3hT469_0(.dout(w_dff_A_nvTYsCxF4_0),.din(w_dff_A_lOg3hT469_0),.clk(gclk));
	jdff dff_A_nvTYsCxF4_0(.dout(w_dff_A_UOH1melP2_0),.din(w_dff_A_nvTYsCxF4_0),.clk(gclk));
	jdff dff_A_UOH1melP2_0(.dout(w_dff_A_hOSC90LA1_0),.din(w_dff_A_UOH1melP2_0),.clk(gclk));
	jdff dff_A_hOSC90LA1_0(.dout(w_dff_A_zZgjbpdi2_0),.din(w_dff_A_hOSC90LA1_0),.clk(gclk));
	jdff dff_A_zZgjbpdi2_0(.dout(w_dff_A_Uiwwkur33_0),.din(w_dff_A_zZgjbpdi2_0),.clk(gclk));
	jdff dff_A_Uiwwkur33_0(.dout(w_dff_A_jolcGtlN3_0),.din(w_dff_A_Uiwwkur33_0),.clk(gclk));
	jdff dff_A_jolcGtlN3_0(.dout(w_dff_A_t8yUvLS06_0),.din(w_dff_A_jolcGtlN3_0),.clk(gclk));
	jdff dff_A_t8yUvLS06_0(.dout(w_dff_A_bprNHvkA9_0),.din(w_dff_A_t8yUvLS06_0),.clk(gclk));
	jdff dff_A_bprNHvkA9_0(.dout(w_dff_A_hqVSzu9O7_0),.din(w_dff_A_bprNHvkA9_0),.clk(gclk));
	jdff dff_A_hqVSzu9O7_0(.dout(w_dff_A_BczsGttN5_0),.din(w_dff_A_hqVSzu9O7_0),.clk(gclk));
	jdff dff_A_BczsGttN5_0(.dout(w_dff_A_GWGiuHbv6_0),.din(w_dff_A_BczsGttN5_0),.clk(gclk));
	jdff dff_A_GWGiuHbv6_0(.dout(w_dff_A_sl5r2OFm7_0),.din(w_dff_A_GWGiuHbv6_0),.clk(gclk));
	jdff dff_A_sl5r2OFm7_0(.dout(w_dff_A_WKgYeipn3_0),.din(w_dff_A_sl5r2OFm7_0),.clk(gclk));
	jdff dff_A_WKgYeipn3_0(.dout(w_dff_A_D25adAZR2_0),.din(w_dff_A_WKgYeipn3_0),.clk(gclk));
	jdff dff_A_D25adAZR2_0(.dout(w_dff_A_KFf0f6sQ7_0),.din(w_dff_A_D25adAZR2_0),.clk(gclk));
	jdff dff_A_KFf0f6sQ7_0(.dout(w_dff_A_kcDh5rxT7_0),.din(w_dff_A_KFf0f6sQ7_0),.clk(gclk));
	jdff dff_A_kcDh5rxT7_0(.dout(w_dff_A_DrA9YxZp8_0),.din(w_dff_A_kcDh5rxT7_0),.clk(gclk));
	jdff dff_A_DrA9YxZp8_0(.dout(w_dff_A_WuUlyEvY4_0),.din(w_dff_A_DrA9YxZp8_0),.clk(gclk));
	jdff dff_A_WuUlyEvY4_0(.dout(w_dff_A_Mff4cG0V7_0),.din(w_dff_A_WuUlyEvY4_0),.clk(gclk));
	jdff dff_A_Mff4cG0V7_0(.dout(w_dff_A_c9hBSiem0_0),.din(w_dff_A_Mff4cG0V7_0),.clk(gclk));
	jdff dff_A_c9hBSiem0_0(.dout(w_dff_A_FCgUzN3v7_0),.din(w_dff_A_c9hBSiem0_0),.clk(gclk));
	jdff dff_A_FCgUzN3v7_0(.dout(w_dff_A_wOqsyxC38_0),.din(w_dff_A_FCgUzN3v7_0),.clk(gclk));
	jdff dff_A_wOqsyxC38_0(.dout(w_dff_A_tqRN59FV1_0),.din(w_dff_A_wOqsyxC38_0),.clk(gclk));
	jdff dff_A_tqRN59FV1_0(.dout(w_dff_A_yIYHvv386_0),.din(w_dff_A_tqRN59FV1_0),.clk(gclk));
	jdff dff_A_yIYHvv386_0(.dout(w_dff_A_LCTdrSdn8_0),.din(w_dff_A_yIYHvv386_0),.clk(gclk));
	jdff dff_A_LCTdrSdn8_0(.dout(w_dff_A_0cQgIh6a9_0),.din(w_dff_A_LCTdrSdn8_0),.clk(gclk));
	jdff dff_A_0cQgIh6a9_0(.dout(w_dff_A_Hmr0BAGN4_0),.din(w_dff_A_0cQgIh6a9_0),.clk(gclk));
	jdff dff_A_Hmr0BAGN4_0(.dout(w_dff_A_Q3JbCeuL7_0),.din(w_dff_A_Hmr0BAGN4_0),.clk(gclk));
	jdff dff_A_Q3JbCeuL7_0(.dout(w_dff_A_2rE6LKwn7_0),.din(w_dff_A_Q3JbCeuL7_0),.clk(gclk));
	jdff dff_A_2rE6LKwn7_0(.dout(w_dff_A_gOlzQcXr3_0),.din(w_dff_A_2rE6LKwn7_0),.clk(gclk));
	jdff dff_A_gOlzQcXr3_0(.dout(w_dff_A_zmuqQX1y4_0),.din(w_dff_A_gOlzQcXr3_0),.clk(gclk));
	jdff dff_A_zmuqQX1y4_0(.dout(w_dff_A_ey3pCS4B0_0),.din(w_dff_A_zmuqQX1y4_0),.clk(gclk));
	jdff dff_A_ey3pCS4B0_0(.dout(w_dff_A_Z7brXAli2_0),.din(w_dff_A_ey3pCS4B0_0),.clk(gclk));
	jdff dff_A_Z7brXAli2_0(.dout(w_dff_A_TlzflgwK5_0),.din(w_dff_A_Z7brXAli2_0),.clk(gclk));
	jdff dff_A_TlzflgwK5_0(.dout(w_dff_A_7Rj678yq1_0),.din(w_dff_A_TlzflgwK5_0),.clk(gclk));
	jdff dff_A_7Rj678yq1_0(.dout(w_dff_A_AcnxaIQN5_0),.din(w_dff_A_7Rj678yq1_0),.clk(gclk));
	jdff dff_A_AcnxaIQN5_0(.dout(w_dff_A_fJH9baaa4_0),.din(w_dff_A_AcnxaIQN5_0),.clk(gclk));
	jdff dff_A_fJH9baaa4_0(.dout(w_dff_A_IIJctWqS5_0),.din(w_dff_A_fJH9baaa4_0),.clk(gclk));
	jdff dff_A_IIJctWqS5_0(.dout(w_dff_A_OrYl9Tm88_0),.din(w_dff_A_IIJctWqS5_0),.clk(gclk));
	jdff dff_A_OrYl9Tm88_0(.dout(w_dff_A_P6h0nl4p4_0),.din(w_dff_A_OrYl9Tm88_0),.clk(gclk));
	jdff dff_A_P6h0nl4p4_0(.dout(w_dff_A_YxfdHJZr6_0),.din(w_dff_A_P6h0nl4p4_0),.clk(gclk));
	jdff dff_A_YxfdHJZr6_0(.dout(w_dff_A_6MOQtoeA0_0),.din(w_dff_A_YxfdHJZr6_0),.clk(gclk));
	jdff dff_A_6MOQtoeA0_0(.dout(w_dff_A_6RpKLiF12_0),.din(w_dff_A_6MOQtoeA0_0),.clk(gclk));
	jdff dff_A_6RpKLiF12_0(.dout(w_dff_A_a2yxjw3a2_0),.din(w_dff_A_6RpKLiF12_0),.clk(gclk));
	jdff dff_A_a2yxjw3a2_0(.dout(w_dff_A_qjzB4Z9t8_0),.din(w_dff_A_a2yxjw3a2_0),.clk(gclk));
	jdff dff_A_qjzB4Z9t8_0(.dout(w_dff_A_jkkUfAJv6_0),.din(w_dff_A_qjzB4Z9t8_0),.clk(gclk));
	jdff dff_A_jkkUfAJv6_0(.dout(w_dff_A_qKMfp8Dt5_0),.din(w_dff_A_jkkUfAJv6_0),.clk(gclk));
	jdff dff_A_qKMfp8Dt5_0(.dout(w_dff_A_WoqI11ms6_0),.din(w_dff_A_qKMfp8Dt5_0),.clk(gclk));
	jdff dff_A_WoqI11ms6_0(.dout(w_dff_A_DlraXJsF2_0),.din(w_dff_A_WoqI11ms6_0),.clk(gclk));
	jdff dff_A_DlraXJsF2_0(.dout(w_dff_A_XR1bFcWX5_0),.din(w_dff_A_DlraXJsF2_0),.clk(gclk));
	jdff dff_A_XR1bFcWX5_0(.dout(w_dff_A_seruZ6Fa5_0),.din(w_dff_A_XR1bFcWX5_0),.clk(gclk));
	jdff dff_A_seruZ6Fa5_0(.dout(w_dff_A_uECwVnlb2_0),.din(w_dff_A_seruZ6Fa5_0),.clk(gclk));
	jdff dff_A_uECwVnlb2_0(.dout(w_dff_A_xTTaLZEK6_0),.din(w_dff_A_uECwVnlb2_0),.clk(gclk));
	jdff dff_A_xTTaLZEK6_0(.dout(w_dff_A_VSXAMPib0_0),.din(w_dff_A_xTTaLZEK6_0),.clk(gclk));
	jdff dff_A_VSXAMPib0_0(.dout(w_dff_A_gH9YZ6uC3_0),.din(w_dff_A_VSXAMPib0_0),.clk(gclk));
	jdff dff_A_gH9YZ6uC3_0(.dout(G1581gat),.din(w_dff_A_gH9YZ6uC3_0),.clk(gclk));
	jdff dff_A_RsDoFRkE0_2(.dout(w_dff_A_pBJQlEGq4_0),.din(w_dff_A_RsDoFRkE0_2),.clk(gclk));
	jdff dff_A_pBJQlEGq4_0(.dout(w_dff_A_RpRULNuW2_0),.din(w_dff_A_pBJQlEGq4_0),.clk(gclk));
	jdff dff_A_RpRULNuW2_0(.dout(w_dff_A_e5HF90ds2_0),.din(w_dff_A_RpRULNuW2_0),.clk(gclk));
	jdff dff_A_e5HF90ds2_0(.dout(w_dff_A_xHzUFE0w9_0),.din(w_dff_A_e5HF90ds2_0),.clk(gclk));
	jdff dff_A_xHzUFE0w9_0(.dout(w_dff_A_iOrBFzvF9_0),.din(w_dff_A_xHzUFE0w9_0),.clk(gclk));
	jdff dff_A_iOrBFzvF9_0(.dout(w_dff_A_uEMgeH9n2_0),.din(w_dff_A_iOrBFzvF9_0),.clk(gclk));
	jdff dff_A_uEMgeH9n2_0(.dout(w_dff_A_gor77tBY3_0),.din(w_dff_A_uEMgeH9n2_0),.clk(gclk));
	jdff dff_A_gor77tBY3_0(.dout(w_dff_A_lTGfop2H9_0),.din(w_dff_A_gor77tBY3_0),.clk(gclk));
	jdff dff_A_lTGfop2H9_0(.dout(w_dff_A_5hbI78dF6_0),.din(w_dff_A_lTGfop2H9_0),.clk(gclk));
	jdff dff_A_5hbI78dF6_0(.dout(w_dff_A_ksLYVnJ73_0),.din(w_dff_A_5hbI78dF6_0),.clk(gclk));
	jdff dff_A_ksLYVnJ73_0(.dout(w_dff_A_r89kxmHk7_0),.din(w_dff_A_ksLYVnJ73_0),.clk(gclk));
	jdff dff_A_r89kxmHk7_0(.dout(w_dff_A_EdmRbVon5_0),.din(w_dff_A_r89kxmHk7_0),.clk(gclk));
	jdff dff_A_EdmRbVon5_0(.dout(w_dff_A_f8wQMqMZ5_0),.din(w_dff_A_EdmRbVon5_0),.clk(gclk));
	jdff dff_A_f8wQMqMZ5_0(.dout(w_dff_A_jB2IyY046_0),.din(w_dff_A_f8wQMqMZ5_0),.clk(gclk));
	jdff dff_A_jB2IyY046_0(.dout(w_dff_A_FxiadecD1_0),.din(w_dff_A_jB2IyY046_0),.clk(gclk));
	jdff dff_A_FxiadecD1_0(.dout(w_dff_A_lVNUDG3p9_0),.din(w_dff_A_FxiadecD1_0),.clk(gclk));
	jdff dff_A_lVNUDG3p9_0(.dout(w_dff_A_xC5aIc0f4_0),.din(w_dff_A_lVNUDG3p9_0),.clk(gclk));
	jdff dff_A_xC5aIc0f4_0(.dout(w_dff_A_bSgQRPoh9_0),.din(w_dff_A_xC5aIc0f4_0),.clk(gclk));
	jdff dff_A_bSgQRPoh9_0(.dout(w_dff_A_KgaSOrHy6_0),.din(w_dff_A_bSgQRPoh9_0),.clk(gclk));
	jdff dff_A_KgaSOrHy6_0(.dout(w_dff_A_kOEpWpVj9_0),.din(w_dff_A_KgaSOrHy6_0),.clk(gclk));
	jdff dff_A_kOEpWpVj9_0(.dout(w_dff_A_y3FjiErL0_0),.din(w_dff_A_kOEpWpVj9_0),.clk(gclk));
	jdff dff_A_y3FjiErL0_0(.dout(w_dff_A_NsKcCNXI8_0),.din(w_dff_A_y3FjiErL0_0),.clk(gclk));
	jdff dff_A_NsKcCNXI8_0(.dout(w_dff_A_VJYGL9nz2_0),.din(w_dff_A_NsKcCNXI8_0),.clk(gclk));
	jdff dff_A_VJYGL9nz2_0(.dout(w_dff_A_fYR45Pcc6_0),.din(w_dff_A_VJYGL9nz2_0),.clk(gclk));
	jdff dff_A_fYR45Pcc6_0(.dout(w_dff_A_XQxi547z9_0),.din(w_dff_A_fYR45Pcc6_0),.clk(gclk));
	jdff dff_A_XQxi547z9_0(.dout(w_dff_A_aQkTh4fg4_0),.din(w_dff_A_XQxi547z9_0),.clk(gclk));
	jdff dff_A_aQkTh4fg4_0(.dout(w_dff_A_qCeRHAc97_0),.din(w_dff_A_aQkTh4fg4_0),.clk(gclk));
	jdff dff_A_qCeRHAc97_0(.dout(w_dff_A_WbrauAlw8_0),.din(w_dff_A_qCeRHAc97_0),.clk(gclk));
	jdff dff_A_WbrauAlw8_0(.dout(w_dff_A_6R7MFucS8_0),.din(w_dff_A_WbrauAlw8_0),.clk(gclk));
	jdff dff_A_6R7MFucS8_0(.dout(w_dff_A_HVv8WAEd0_0),.din(w_dff_A_6R7MFucS8_0),.clk(gclk));
	jdff dff_A_HVv8WAEd0_0(.dout(w_dff_A_yQOLCmJe4_0),.din(w_dff_A_HVv8WAEd0_0),.clk(gclk));
	jdff dff_A_yQOLCmJe4_0(.dout(w_dff_A_fChpvAtV5_0),.din(w_dff_A_yQOLCmJe4_0),.clk(gclk));
	jdff dff_A_fChpvAtV5_0(.dout(w_dff_A_BVLGAnCp0_0),.din(w_dff_A_fChpvAtV5_0),.clk(gclk));
	jdff dff_A_BVLGAnCp0_0(.dout(w_dff_A_LQGeLPW69_0),.din(w_dff_A_BVLGAnCp0_0),.clk(gclk));
	jdff dff_A_LQGeLPW69_0(.dout(w_dff_A_oD6FFUYu2_0),.din(w_dff_A_LQGeLPW69_0),.clk(gclk));
	jdff dff_A_oD6FFUYu2_0(.dout(w_dff_A_ZUlnMcF51_0),.din(w_dff_A_oD6FFUYu2_0),.clk(gclk));
	jdff dff_A_ZUlnMcF51_0(.dout(w_dff_A_M1tCmev92_0),.din(w_dff_A_ZUlnMcF51_0),.clk(gclk));
	jdff dff_A_M1tCmev92_0(.dout(w_dff_A_XjMUxa4I3_0),.din(w_dff_A_M1tCmev92_0),.clk(gclk));
	jdff dff_A_XjMUxa4I3_0(.dout(w_dff_A_ng7UeUqS7_0),.din(w_dff_A_XjMUxa4I3_0),.clk(gclk));
	jdff dff_A_ng7UeUqS7_0(.dout(w_dff_A_eZ3uWlS54_0),.din(w_dff_A_ng7UeUqS7_0),.clk(gclk));
	jdff dff_A_eZ3uWlS54_0(.dout(w_dff_A_CwRbadB94_0),.din(w_dff_A_eZ3uWlS54_0),.clk(gclk));
	jdff dff_A_CwRbadB94_0(.dout(w_dff_A_PfMru1ON8_0),.din(w_dff_A_CwRbadB94_0),.clk(gclk));
	jdff dff_A_PfMru1ON8_0(.dout(w_dff_A_5eTsrVw56_0),.din(w_dff_A_PfMru1ON8_0),.clk(gclk));
	jdff dff_A_5eTsrVw56_0(.dout(w_dff_A_4RbthjPL5_0),.din(w_dff_A_5eTsrVw56_0),.clk(gclk));
	jdff dff_A_4RbthjPL5_0(.dout(w_dff_A_ivKjnPzW9_0),.din(w_dff_A_4RbthjPL5_0),.clk(gclk));
	jdff dff_A_ivKjnPzW9_0(.dout(w_dff_A_i7bn42BC5_0),.din(w_dff_A_ivKjnPzW9_0),.clk(gclk));
	jdff dff_A_i7bn42BC5_0(.dout(w_dff_A_P3QsJjAa4_0),.din(w_dff_A_i7bn42BC5_0),.clk(gclk));
	jdff dff_A_P3QsJjAa4_0(.dout(w_dff_A_J7k8xNCL0_0),.din(w_dff_A_P3QsJjAa4_0),.clk(gclk));
	jdff dff_A_J7k8xNCL0_0(.dout(w_dff_A_YQ2HGsbt8_0),.din(w_dff_A_J7k8xNCL0_0),.clk(gclk));
	jdff dff_A_YQ2HGsbt8_0(.dout(w_dff_A_NONL67SN7_0),.din(w_dff_A_YQ2HGsbt8_0),.clk(gclk));
	jdff dff_A_NONL67SN7_0(.dout(w_dff_A_w6JVu9bk2_0),.din(w_dff_A_NONL67SN7_0),.clk(gclk));
	jdff dff_A_w6JVu9bk2_0(.dout(w_dff_A_qX4I8RST4_0),.din(w_dff_A_w6JVu9bk2_0),.clk(gclk));
	jdff dff_A_qX4I8RST4_0(.dout(w_dff_A_oEw0h3W95_0),.din(w_dff_A_qX4I8RST4_0),.clk(gclk));
	jdff dff_A_oEw0h3W95_0(.dout(w_dff_A_I1mHrml95_0),.din(w_dff_A_oEw0h3W95_0),.clk(gclk));
	jdff dff_A_I1mHrml95_0(.dout(w_dff_A_6kZC3iJ04_0),.din(w_dff_A_I1mHrml95_0),.clk(gclk));
	jdff dff_A_6kZC3iJ04_0(.dout(w_dff_A_9wRRePUh6_0),.din(w_dff_A_6kZC3iJ04_0),.clk(gclk));
	jdff dff_A_9wRRePUh6_0(.dout(w_dff_A_jhNXnTh20_0),.din(w_dff_A_9wRRePUh6_0),.clk(gclk));
	jdff dff_A_jhNXnTh20_0(.dout(w_dff_A_fh7eCDxo5_0),.din(w_dff_A_jhNXnTh20_0),.clk(gclk));
	jdff dff_A_fh7eCDxo5_0(.dout(w_dff_A_7AUygaGH5_0),.din(w_dff_A_fh7eCDxo5_0),.clk(gclk));
	jdff dff_A_7AUygaGH5_0(.dout(w_dff_A_kaZy14qm6_0),.din(w_dff_A_7AUygaGH5_0),.clk(gclk));
	jdff dff_A_kaZy14qm6_0(.dout(w_dff_A_aYs1nTHT3_0),.din(w_dff_A_kaZy14qm6_0),.clk(gclk));
	jdff dff_A_aYs1nTHT3_0(.dout(w_dff_A_8j8dHqgh7_0),.din(w_dff_A_aYs1nTHT3_0),.clk(gclk));
	jdff dff_A_8j8dHqgh7_0(.dout(w_dff_A_XAWMuwmi4_0),.din(w_dff_A_8j8dHqgh7_0),.clk(gclk));
	jdff dff_A_XAWMuwmi4_0(.dout(w_dff_A_H7UTNw2z5_0),.din(w_dff_A_XAWMuwmi4_0),.clk(gclk));
	jdff dff_A_H7UTNw2z5_0(.dout(w_dff_A_YznWS3Lm1_0),.din(w_dff_A_H7UTNw2z5_0),.clk(gclk));
	jdff dff_A_YznWS3Lm1_0(.dout(w_dff_A_RLSTf5Bj2_0),.din(w_dff_A_YznWS3Lm1_0),.clk(gclk));
	jdff dff_A_RLSTf5Bj2_0(.dout(w_dff_A_MqlPqEgi9_0),.din(w_dff_A_RLSTf5Bj2_0),.clk(gclk));
	jdff dff_A_MqlPqEgi9_0(.dout(w_dff_A_pjydccY89_0),.din(w_dff_A_MqlPqEgi9_0),.clk(gclk));
	jdff dff_A_pjydccY89_0(.dout(G1901gat),.din(w_dff_A_pjydccY89_0),.clk(gclk));
	jdff dff_A_1xLXBDUh1_2(.dout(w_dff_A_xsu4rBt49_0),.din(w_dff_A_1xLXBDUh1_2),.clk(gclk));
	jdff dff_A_xsu4rBt49_0(.dout(w_dff_A_k5BkWBtk7_0),.din(w_dff_A_xsu4rBt49_0),.clk(gclk));
	jdff dff_A_k5BkWBtk7_0(.dout(w_dff_A_PQVsFRFi2_0),.din(w_dff_A_k5BkWBtk7_0),.clk(gclk));
	jdff dff_A_PQVsFRFi2_0(.dout(w_dff_A_uku0ZAZR9_0),.din(w_dff_A_PQVsFRFi2_0),.clk(gclk));
	jdff dff_A_uku0ZAZR9_0(.dout(w_dff_A_QfYY0DpD5_0),.din(w_dff_A_uku0ZAZR9_0),.clk(gclk));
	jdff dff_A_QfYY0DpD5_0(.dout(w_dff_A_jbDrEcJ23_0),.din(w_dff_A_QfYY0DpD5_0),.clk(gclk));
	jdff dff_A_jbDrEcJ23_0(.dout(w_dff_A_yROG9dB01_0),.din(w_dff_A_jbDrEcJ23_0),.clk(gclk));
	jdff dff_A_yROG9dB01_0(.dout(w_dff_A_CXPogtxx2_0),.din(w_dff_A_yROG9dB01_0),.clk(gclk));
	jdff dff_A_CXPogtxx2_0(.dout(w_dff_A_PI1ULLSU5_0),.din(w_dff_A_CXPogtxx2_0),.clk(gclk));
	jdff dff_A_PI1ULLSU5_0(.dout(w_dff_A_vkm5UZvG5_0),.din(w_dff_A_PI1ULLSU5_0),.clk(gclk));
	jdff dff_A_vkm5UZvG5_0(.dout(w_dff_A_yyMowZzA1_0),.din(w_dff_A_vkm5UZvG5_0),.clk(gclk));
	jdff dff_A_yyMowZzA1_0(.dout(w_dff_A_LEaF1bsA9_0),.din(w_dff_A_yyMowZzA1_0),.clk(gclk));
	jdff dff_A_LEaF1bsA9_0(.dout(w_dff_A_OEZJW24h5_0),.din(w_dff_A_LEaF1bsA9_0),.clk(gclk));
	jdff dff_A_OEZJW24h5_0(.dout(w_dff_A_BBagiyHD6_0),.din(w_dff_A_OEZJW24h5_0),.clk(gclk));
	jdff dff_A_BBagiyHD6_0(.dout(w_dff_A_sdXcLymA1_0),.din(w_dff_A_BBagiyHD6_0),.clk(gclk));
	jdff dff_A_sdXcLymA1_0(.dout(w_dff_A_UCRcqDta2_0),.din(w_dff_A_sdXcLymA1_0),.clk(gclk));
	jdff dff_A_UCRcqDta2_0(.dout(w_dff_A_9jIW1bJN9_0),.din(w_dff_A_UCRcqDta2_0),.clk(gclk));
	jdff dff_A_9jIW1bJN9_0(.dout(w_dff_A_FZ2ww8gG4_0),.din(w_dff_A_9jIW1bJN9_0),.clk(gclk));
	jdff dff_A_FZ2ww8gG4_0(.dout(w_dff_A_7yokyOKu5_0),.din(w_dff_A_FZ2ww8gG4_0),.clk(gclk));
	jdff dff_A_7yokyOKu5_0(.dout(w_dff_A_ztLbhzp60_0),.din(w_dff_A_7yokyOKu5_0),.clk(gclk));
	jdff dff_A_ztLbhzp60_0(.dout(w_dff_A_0Cqhj6Rl1_0),.din(w_dff_A_ztLbhzp60_0),.clk(gclk));
	jdff dff_A_0Cqhj6Rl1_0(.dout(w_dff_A_qahTg1QR1_0),.din(w_dff_A_0Cqhj6Rl1_0),.clk(gclk));
	jdff dff_A_qahTg1QR1_0(.dout(w_dff_A_QfbEFPs25_0),.din(w_dff_A_qahTg1QR1_0),.clk(gclk));
	jdff dff_A_QfbEFPs25_0(.dout(w_dff_A_v8TmBlNa9_0),.din(w_dff_A_QfbEFPs25_0),.clk(gclk));
	jdff dff_A_v8TmBlNa9_0(.dout(w_dff_A_GJoZHAUJ7_0),.din(w_dff_A_v8TmBlNa9_0),.clk(gclk));
	jdff dff_A_GJoZHAUJ7_0(.dout(w_dff_A_nzm2KIE60_0),.din(w_dff_A_GJoZHAUJ7_0),.clk(gclk));
	jdff dff_A_nzm2KIE60_0(.dout(w_dff_A_PD83B6Xq1_0),.din(w_dff_A_nzm2KIE60_0),.clk(gclk));
	jdff dff_A_PD83B6Xq1_0(.dout(w_dff_A_JjlHrhjj7_0),.din(w_dff_A_PD83B6Xq1_0),.clk(gclk));
	jdff dff_A_JjlHrhjj7_0(.dout(w_dff_A_YvhTfQmM9_0),.din(w_dff_A_JjlHrhjj7_0),.clk(gclk));
	jdff dff_A_YvhTfQmM9_0(.dout(w_dff_A_J01bPRDU4_0),.din(w_dff_A_YvhTfQmM9_0),.clk(gclk));
	jdff dff_A_J01bPRDU4_0(.dout(w_dff_A_WI4akYC37_0),.din(w_dff_A_J01bPRDU4_0),.clk(gclk));
	jdff dff_A_WI4akYC37_0(.dout(w_dff_A_Bcsxoab35_0),.din(w_dff_A_WI4akYC37_0),.clk(gclk));
	jdff dff_A_Bcsxoab35_0(.dout(w_dff_A_sgOk7ufr0_0),.din(w_dff_A_Bcsxoab35_0),.clk(gclk));
	jdff dff_A_sgOk7ufr0_0(.dout(w_dff_A_6NFXLFB45_0),.din(w_dff_A_sgOk7ufr0_0),.clk(gclk));
	jdff dff_A_6NFXLFB45_0(.dout(w_dff_A_klwxy7Cy6_0),.din(w_dff_A_6NFXLFB45_0),.clk(gclk));
	jdff dff_A_klwxy7Cy6_0(.dout(w_dff_A_G0fSCz8P5_0),.din(w_dff_A_klwxy7Cy6_0),.clk(gclk));
	jdff dff_A_G0fSCz8P5_0(.dout(w_dff_A_KInQa8R52_0),.din(w_dff_A_G0fSCz8P5_0),.clk(gclk));
	jdff dff_A_KInQa8R52_0(.dout(w_dff_A_IImVZS1d6_0),.din(w_dff_A_KInQa8R52_0),.clk(gclk));
	jdff dff_A_IImVZS1d6_0(.dout(w_dff_A_SsgU5SUW7_0),.din(w_dff_A_IImVZS1d6_0),.clk(gclk));
	jdff dff_A_SsgU5SUW7_0(.dout(w_dff_A_LW1yZJdS0_0),.din(w_dff_A_SsgU5SUW7_0),.clk(gclk));
	jdff dff_A_LW1yZJdS0_0(.dout(w_dff_A_XY7yEhb46_0),.din(w_dff_A_LW1yZJdS0_0),.clk(gclk));
	jdff dff_A_XY7yEhb46_0(.dout(w_dff_A_YyDSFjD11_0),.din(w_dff_A_XY7yEhb46_0),.clk(gclk));
	jdff dff_A_YyDSFjD11_0(.dout(w_dff_A_NmETfZSo8_0),.din(w_dff_A_YyDSFjD11_0),.clk(gclk));
	jdff dff_A_NmETfZSo8_0(.dout(w_dff_A_ItpO6lpb2_0),.din(w_dff_A_NmETfZSo8_0),.clk(gclk));
	jdff dff_A_ItpO6lpb2_0(.dout(w_dff_A_1qpEqiuq9_0),.din(w_dff_A_ItpO6lpb2_0),.clk(gclk));
	jdff dff_A_1qpEqiuq9_0(.dout(w_dff_A_tM64kL2f2_0),.din(w_dff_A_1qpEqiuq9_0),.clk(gclk));
	jdff dff_A_tM64kL2f2_0(.dout(w_dff_A_ZtCEnyOQ6_0),.din(w_dff_A_tM64kL2f2_0),.clk(gclk));
	jdff dff_A_ZtCEnyOQ6_0(.dout(w_dff_A_QHOWo0RC7_0),.din(w_dff_A_ZtCEnyOQ6_0),.clk(gclk));
	jdff dff_A_QHOWo0RC7_0(.dout(w_dff_A_o390FudG3_0),.din(w_dff_A_QHOWo0RC7_0),.clk(gclk));
	jdff dff_A_o390FudG3_0(.dout(w_dff_A_OeteqeBr8_0),.din(w_dff_A_o390FudG3_0),.clk(gclk));
	jdff dff_A_OeteqeBr8_0(.dout(w_dff_A_nbB6fwHd1_0),.din(w_dff_A_OeteqeBr8_0),.clk(gclk));
	jdff dff_A_nbB6fwHd1_0(.dout(w_dff_A_Xl6aWd1Q2_0),.din(w_dff_A_nbB6fwHd1_0),.clk(gclk));
	jdff dff_A_Xl6aWd1Q2_0(.dout(w_dff_A_pJ8IjpaS8_0),.din(w_dff_A_Xl6aWd1Q2_0),.clk(gclk));
	jdff dff_A_pJ8IjpaS8_0(.dout(w_dff_A_yQiChqBE2_0),.din(w_dff_A_pJ8IjpaS8_0),.clk(gclk));
	jdff dff_A_yQiChqBE2_0(.dout(w_dff_A_Lps2nWTL1_0),.din(w_dff_A_yQiChqBE2_0),.clk(gclk));
	jdff dff_A_Lps2nWTL1_0(.dout(w_dff_A_6D2gNe7X0_0),.din(w_dff_A_Lps2nWTL1_0),.clk(gclk));
	jdff dff_A_6D2gNe7X0_0(.dout(w_dff_A_aOa9I9ae0_0),.din(w_dff_A_6D2gNe7X0_0),.clk(gclk));
	jdff dff_A_aOa9I9ae0_0(.dout(w_dff_A_idDgyRDr6_0),.din(w_dff_A_aOa9I9ae0_0),.clk(gclk));
	jdff dff_A_idDgyRDr6_0(.dout(w_dff_A_lWgC5v9h6_0),.din(w_dff_A_idDgyRDr6_0),.clk(gclk));
	jdff dff_A_lWgC5v9h6_0(.dout(w_dff_A_HSrCP0S49_0),.din(w_dff_A_lWgC5v9h6_0),.clk(gclk));
	jdff dff_A_HSrCP0S49_0(.dout(w_dff_A_PzcSGmdm1_0),.din(w_dff_A_HSrCP0S49_0),.clk(gclk));
	jdff dff_A_PzcSGmdm1_0(.dout(w_dff_A_RTbgOhM20_0),.din(w_dff_A_PzcSGmdm1_0),.clk(gclk));
	jdff dff_A_RTbgOhM20_0(.dout(w_dff_A_lWXAxUYh0_0),.din(w_dff_A_RTbgOhM20_0),.clk(gclk));
	jdff dff_A_lWXAxUYh0_0(.dout(w_dff_A_F9LmMSId0_0),.din(w_dff_A_lWXAxUYh0_0),.clk(gclk));
	jdff dff_A_F9LmMSId0_0(.dout(w_dff_A_CmXVFCyd7_0),.din(w_dff_A_F9LmMSId0_0),.clk(gclk));
	jdff dff_A_CmXVFCyd7_0(.dout(G2223gat),.din(w_dff_A_CmXVFCyd7_0),.clk(gclk));
	jdff dff_A_TeLedrld7_2(.dout(w_dff_A_bol0ejVz0_0),.din(w_dff_A_TeLedrld7_2),.clk(gclk));
	jdff dff_A_bol0ejVz0_0(.dout(w_dff_A_t4LhVYjM3_0),.din(w_dff_A_bol0ejVz0_0),.clk(gclk));
	jdff dff_A_t4LhVYjM3_0(.dout(w_dff_A_uacpOgHi5_0),.din(w_dff_A_t4LhVYjM3_0),.clk(gclk));
	jdff dff_A_uacpOgHi5_0(.dout(w_dff_A_IU4O6lmQ3_0),.din(w_dff_A_uacpOgHi5_0),.clk(gclk));
	jdff dff_A_IU4O6lmQ3_0(.dout(w_dff_A_0VuVsBaC5_0),.din(w_dff_A_IU4O6lmQ3_0),.clk(gclk));
	jdff dff_A_0VuVsBaC5_0(.dout(w_dff_A_wCLjnwhq7_0),.din(w_dff_A_0VuVsBaC5_0),.clk(gclk));
	jdff dff_A_wCLjnwhq7_0(.dout(w_dff_A_Ko6gxlib0_0),.din(w_dff_A_wCLjnwhq7_0),.clk(gclk));
	jdff dff_A_Ko6gxlib0_0(.dout(w_dff_A_3f08bY8f1_0),.din(w_dff_A_Ko6gxlib0_0),.clk(gclk));
	jdff dff_A_3f08bY8f1_0(.dout(w_dff_A_8ijIKzc73_0),.din(w_dff_A_3f08bY8f1_0),.clk(gclk));
	jdff dff_A_8ijIKzc73_0(.dout(w_dff_A_n6T3EC4L6_0),.din(w_dff_A_8ijIKzc73_0),.clk(gclk));
	jdff dff_A_n6T3EC4L6_0(.dout(w_dff_A_H1OWfJyx6_0),.din(w_dff_A_n6T3EC4L6_0),.clk(gclk));
	jdff dff_A_H1OWfJyx6_0(.dout(w_dff_A_oiTuYJ3v0_0),.din(w_dff_A_H1OWfJyx6_0),.clk(gclk));
	jdff dff_A_oiTuYJ3v0_0(.dout(w_dff_A_eKp0PLuY3_0),.din(w_dff_A_oiTuYJ3v0_0),.clk(gclk));
	jdff dff_A_eKp0PLuY3_0(.dout(w_dff_A_WUv6ZO6t9_0),.din(w_dff_A_eKp0PLuY3_0),.clk(gclk));
	jdff dff_A_WUv6ZO6t9_0(.dout(w_dff_A_oT4gjTtw8_0),.din(w_dff_A_WUv6ZO6t9_0),.clk(gclk));
	jdff dff_A_oT4gjTtw8_0(.dout(w_dff_A_EVMTMoUN5_0),.din(w_dff_A_oT4gjTtw8_0),.clk(gclk));
	jdff dff_A_EVMTMoUN5_0(.dout(w_dff_A_qMDPQIDd0_0),.din(w_dff_A_EVMTMoUN5_0),.clk(gclk));
	jdff dff_A_qMDPQIDd0_0(.dout(w_dff_A_t1zI0mwr3_0),.din(w_dff_A_qMDPQIDd0_0),.clk(gclk));
	jdff dff_A_t1zI0mwr3_0(.dout(w_dff_A_bs5lZ3yU2_0),.din(w_dff_A_t1zI0mwr3_0),.clk(gclk));
	jdff dff_A_bs5lZ3yU2_0(.dout(w_dff_A_XnxGtaX32_0),.din(w_dff_A_bs5lZ3yU2_0),.clk(gclk));
	jdff dff_A_XnxGtaX32_0(.dout(w_dff_A_ZXXVlMKK2_0),.din(w_dff_A_XnxGtaX32_0),.clk(gclk));
	jdff dff_A_ZXXVlMKK2_0(.dout(w_dff_A_Vt9Hp3ou0_0),.din(w_dff_A_ZXXVlMKK2_0),.clk(gclk));
	jdff dff_A_Vt9Hp3ou0_0(.dout(w_dff_A_yv2P0WMO0_0),.din(w_dff_A_Vt9Hp3ou0_0),.clk(gclk));
	jdff dff_A_yv2P0WMO0_0(.dout(w_dff_A_VKYp5l2u8_0),.din(w_dff_A_yv2P0WMO0_0),.clk(gclk));
	jdff dff_A_VKYp5l2u8_0(.dout(w_dff_A_9uwWeksb3_0),.din(w_dff_A_VKYp5l2u8_0),.clk(gclk));
	jdff dff_A_9uwWeksb3_0(.dout(w_dff_A_7u72UeB25_0),.din(w_dff_A_9uwWeksb3_0),.clk(gclk));
	jdff dff_A_7u72UeB25_0(.dout(w_dff_A_BJAw2yFA0_0),.din(w_dff_A_7u72UeB25_0),.clk(gclk));
	jdff dff_A_BJAw2yFA0_0(.dout(w_dff_A_JZWhghGf9_0),.din(w_dff_A_BJAw2yFA0_0),.clk(gclk));
	jdff dff_A_JZWhghGf9_0(.dout(w_dff_A_X96sUsPH8_0),.din(w_dff_A_JZWhghGf9_0),.clk(gclk));
	jdff dff_A_X96sUsPH8_0(.dout(w_dff_A_v6cG4XWl5_0),.din(w_dff_A_X96sUsPH8_0),.clk(gclk));
	jdff dff_A_v6cG4XWl5_0(.dout(w_dff_A_iEfdnanX3_0),.din(w_dff_A_v6cG4XWl5_0),.clk(gclk));
	jdff dff_A_iEfdnanX3_0(.dout(w_dff_A_8dtyyjYc7_0),.din(w_dff_A_iEfdnanX3_0),.clk(gclk));
	jdff dff_A_8dtyyjYc7_0(.dout(w_dff_A_dou3YUic3_0),.din(w_dff_A_8dtyyjYc7_0),.clk(gclk));
	jdff dff_A_dou3YUic3_0(.dout(w_dff_A_17qQnhVk4_0),.din(w_dff_A_dou3YUic3_0),.clk(gclk));
	jdff dff_A_17qQnhVk4_0(.dout(w_dff_A_IqYsLYKj4_0),.din(w_dff_A_17qQnhVk4_0),.clk(gclk));
	jdff dff_A_IqYsLYKj4_0(.dout(w_dff_A_BeU2OFCx0_0),.din(w_dff_A_IqYsLYKj4_0),.clk(gclk));
	jdff dff_A_BeU2OFCx0_0(.dout(w_dff_A_HnQaH6tW5_0),.din(w_dff_A_BeU2OFCx0_0),.clk(gclk));
	jdff dff_A_HnQaH6tW5_0(.dout(w_dff_A_drPL1Zui5_0),.din(w_dff_A_HnQaH6tW5_0),.clk(gclk));
	jdff dff_A_drPL1Zui5_0(.dout(w_dff_A_LLT0fVxj1_0),.din(w_dff_A_drPL1Zui5_0),.clk(gclk));
	jdff dff_A_LLT0fVxj1_0(.dout(w_dff_A_kDsHfPOj1_0),.din(w_dff_A_LLT0fVxj1_0),.clk(gclk));
	jdff dff_A_kDsHfPOj1_0(.dout(w_dff_A_5i3tz4Zv8_0),.din(w_dff_A_kDsHfPOj1_0),.clk(gclk));
	jdff dff_A_5i3tz4Zv8_0(.dout(w_dff_A_qq3dITRB2_0),.din(w_dff_A_5i3tz4Zv8_0),.clk(gclk));
	jdff dff_A_qq3dITRB2_0(.dout(w_dff_A_ky4f0O2O2_0),.din(w_dff_A_qq3dITRB2_0),.clk(gclk));
	jdff dff_A_ky4f0O2O2_0(.dout(w_dff_A_PvON90P24_0),.din(w_dff_A_ky4f0O2O2_0),.clk(gclk));
	jdff dff_A_PvON90P24_0(.dout(w_dff_A_pF6tsaKP3_0),.din(w_dff_A_PvON90P24_0),.clk(gclk));
	jdff dff_A_pF6tsaKP3_0(.dout(w_dff_A_atT6eD336_0),.din(w_dff_A_pF6tsaKP3_0),.clk(gclk));
	jdff dff_A_atT6eD336_0(.dout(w_dff_A_Y3ohAWku0_0),.din(w_dff_A_atT6eD336_0),.clk(gclk));
	jdff dff_A_Y3ohAWku0_0(.dout(w_dff_A_kLfdbApj6_0),.din(w_dff_A_Y3ohAWku0_0),.clk(gclk));
	jdff dff_A_kLfdbApj6_0(.dout(w_dff_A_XqbapEyq8_0),.din(w_dff_A_kLfdbApj6_0),.clk(gclk));
	jdff dff_A_XqbapEyq8_0(.dout(w_dff_A_VjlNLbQz5_0),.din(w_dff_A_XqbapEyq8_0),.clk(gclk));
	jdff dff_A_VjlNLbQz5_0(.dout(w_dff_A_DeEPtQdM3_0),.din(w_dff_A_VjlNLbQz5_0),.clk(gclk));
	jdff dff_A_DeEPtQdM3_0(.dout(w_dff_A_ZosguoP75_0),.din(w_dff_A_DeEPtQdM3_0),.clk(gclk));
	jdff dff_A_ZosguoP75_0(.dout(w_dff_A_cwWfmgn85_0),.din(w_dff_A_ZosguoP75_0),.clk(gclk));
	jdff dff_A_cwWfmgn85_0(.dout(w_dff_A_bze71XGT3_0),.din(w_dff_A_cwWfmgn85_0),.clk(gclk));
	jdff dff_A_bze71XGT3_0(.dout(w_dff_A_5mX8apPa9_0),.din(w_dff_A_bze71XGT3_0),.clk(gclk));
	jdff dff_A_5mX8apPa9_0(.dout(w_dff_A_4YqBnL7B1_0),.din(w_dff_A_5mX8apPa9_0),.clk(gclk));
	jdff dff_A_4YqBnL7B1_0(.dout(w_dff_A_cbasXw8a5_0),.din(w_dff_A_4YqBnL7B1_0),.clk(gclk));
	jdff dff_A_cbasXw8a5_0(.dout(w_dff_A_zr21BW4f6_0),.din(w_dff_A_cbasXw8a5_0),.clk(gclk));
	jdff dff_A_zr21BW4f6_0(.dout(w_dff_A_cMAfwCVk0_0),.din(w_dff_A_zr21BW4f6_0),.clk(gclk));
	jdff dff_A_cMAfwCVk0_0(.dout(w_dff_A_pJ33Hvnf2_0),.din(w_dff_A_cMAfwCVk0_0),.clk(gclk));
	jdff dff_A_pJ33Hvnf2_0(.dout(w_dff_A_z7YRI3e49_0),.din(w_dff_A_pJ33Hvnf2_0),.clk(gclk));
	jdff dff_A_z7YRI3e49_0(.dout(w_dff_A_vT9YTuSq8_0),.din(w_dff_A_z7YRI3e49_0),.clk(gclk));
	jdff dff_A_vT9YTuSq8_0(.dout(G2548gat),.din(w_dff_A_vT9YTuSq8_0),.clk(gclk));
	jdff dff_A_TwM7lXbz1_2(.dout(w_dff_A_UAJW3X5l7_0),.din(w_dff_A_TwM7lXbz1_2),.clk(gclk));
	jdff dff_A_UAJW3X5l7_0(.dout(w_dff_A_j9B9Jvno8_0),.din(w_dff_A_UAJW3X5l7_0),.clk(gclk));
	jdff dff_A_j9B9Jvno8_0(.dout(w_dff_A_Q0c5kvtw1_0),.din(w_dff_A_j9B9Jvno8_0),.clk(gclk));
	jdff dff_A_Q0c5kvtw1_0(.dout(w_dff_A_jIDC6kEQ7_0),.din(w_dff_A_Q0c5kvtw1_0),.clk(gclk));
	jdff dff_A_jIDC6kEQ7_0(.dout(w_dff_A_9JDPLOyP6_0),.din(w_dff_A_jIDC6kEQ7_0),.clk(gclk));
	jdff dff_A_9JDPLOyP6_0(.dout(w_dff_A_sTrmOqhF6_0),.din(w_dff_A_9JDPLOyP6_0),.clk(gclk));
	jdff dff_A_sTrmOqhF6_0(.dout(w_dff_A_ZEdZut1c0_0),.din(w_dff_A_sTrmOqhF6_0),.clk(gclk));
	jdff dff_A_ZEdZut1c0_0(.dout(w_dff_A_4eYIvfCU3_0),.din(w_dff_A_ZEdZut1c0_0),.clk(gclk));
	jdff dff_A_4eYIvfCU3_0(.dout(w_dff_A_W9nowCdM3_0),.din(w_dff_A_4eYIvfCU3_0),.clk(gclk));
	jdff dff_A_W9nowCdM3_0(.dout(w_dff_A_FCeCjAjz7_0),.din(w_dff_A_W9nowCdM3_0),.clk(gclk));
	jdff dff_A_FCeCjAjz7_0(.dout(w_dff_A_RCFfnfy77_0),.din(w_dff_A_FCeCjAjz7_0),.clk(gclk));
	jdff dff_A_RCFfnfy77_0(.dout(w_dff_A_PucO2c7U3_0),.din(w_dff_A_RCFfnfy77_0),.clk(gclk));
	jdff dff_A_PucO2c7U3_0(.dout(w_dff_A_Whz0sEPe6_0),.din(w_dff_A_PucO2c7U3_0),.clk(gclk));
	jdff dff_A_Whz0sEPe6_0(.dout(w_dff_A_VeyoKap24_0),.din(w_dff_A_Whz0sEPe6_0),.clk(gclk));
	jdff dff_A_VeyoKap24_0(.dout(w_dff_A_jpfNtqAp9_0),.din(w_dff_A_VeyoKap24_0),.clk(gclk));
	jdff dff_A_jpfNtqAp9_0(.dout(w_dff_A_1miHCnrf2_0),.din(w_dff_A_jpfNtqAp9_0),.clk(gclk));
	jdff dff_A_1miHCnrf2_0(.dout(w_dff_A_964Cxv4P3_0),.din(w_dff_A_1miHCnrf2_0),.clk(gclk));
	jdff dff_A_964Cxv4P3_0(.dout(w_dff_A_jDHBWnsD0_0),.din(w_dff_A_964Cxv4P3_0),.clk(gclk));
	jdff dff_A_jDHBWnsD0_0(.dout(w_dff_A_0qfWCUNQ3_0),.din(w_dff_A_jDHBWnsD0_0),.clk(gclk));
	jdff dff_A_0qfWCUNQ3_0(.dout(w_dff_A_YQudfU5M5_0),.din(w_dff_A_0qfWCUNQ3_0),.clk(gclk));
	jdff dff_A_YQudfU5M5_0(.dout(w_dff_A_CGmkKv4x4_0),.din(w_dff_A_YQudfU5M5_0),.clk(gclk));
	jdff dff_A_CGmkKv4x4_0(.dout(w_dff_A_i8A7DZtS8_0),.din(w_dff_A_CGmkKv4x4_0),.clk(gclk));
	jdff dff_A_i8A7DZtS8_0(.dout(w_dff_A_WyQ2V4mb9_0),.din(w_dff_A_i8A7DZtS8_0),.clk(gclk));
	jdff dff_A_WyQ2V4mb9_0(.dout(w_dff_A_8qSuFptH6_0),.din(w_dff_A_WyQ2V4mb9_0),.clk(gclk));
	jdff dff_A_8qSuFptH6_0(.dout(w_dff_A_qlC1par80_0),.din(w_dff_A_8qSuFptH6_0),.clk(gclk));
	jdff dff_A_qlC1par80_0(.dout(w_dff_A_6GLPw8WD8_0),.din(w_dff_A_qlC1par80_0),.clk(gclk));
	jdff dff_A_6GLPw8WD8_0(.dout(w_dff_A_OxYs3xHo5_0),.din(w_dff_A_6GLPw8WD8_0),.clk(gclk));
	jdff dff_A_OxYs3xHo5_0(.dout(w_dff_A_VfmVkD5U5_0),.din(w_dff_A_OxYs3xHo5_0),.clk(gclk));
	jdff dff_A_VfmVkD5U5_0(.dout(w_dff_A_zXjrJcwF9_0),.din(w_dff_A_VfmVkD5U5_0),.clk(gclk));
	jdff dff_A_zXjrJcwF9_0(.dout(w_dff_A_6HQEtJCb3_0),.din(w_dff_A_zXjrJcwF9_0),.clk(gclk));
	jdff dff_A_6HQEtJCb3_0(.dout(w_dff_A_CqBS3ekW3_0),.din(w_dff_A_6HQEtJCb3_0),.clk(gclk));
	jdff dff_A_CqBS3ekW3_0(.dout(w_dff_A_39PURsZS2_0),.din(w_dff_A_CqBS3ekW3_0),.clk(gclk));
	jdff dff_A_39PURsZS2_0(.dout(w_dff_A_9BBI98LA7_0),.din(w_dff_A_39PURsZS2_0),.clk(gclk));
	jdff dff_A_9BBI98LA7_0(.dout(w_dff_A_1AzSRlcb6_0),.din(w_dff_A_9BBI98LA7_0),.clk(gclk));
	jdff dff_A_1AzSRlcb6_0(.dout(w_dff_A_SPKTtnlj1_0),.din(w_dff_A_1AzSRlcb6_0),.clk(gclk));
	jdff dff_A_SPKTtnlj1_0(.dout(w_dff_A_dknCnWo04_0),.din(w_dff_A_SPKTtnlj1_0),.clk(gclk));
	jdff dff_A_dknCnWo04_0(.dout(w_dff_A_g7BbC1sk9_0),.din(w_dff_A_dknCnWo04_0),.clk(gclk));
	jdff dff_A_g7BbC1sk9_0(.dout(w_dff_A_1pagNIXs4_0),.din(w_dff_A_g7BbC1sk9_0),.clk(gclk));
	jdff dff_A_1pagNIXs4_0(.dout(w_dff_A_Rsnqd1pV2_0),.din(w_dff_A_1pagNIXs4_0),.clk(gclk));
	jdff dff_A_Rsnqd1pV2_0(.dout(w_dff_A_BdbkCvEe4_0),.din(w_dff_A_Rsnqd1pV2_0),.clk(gclk));
	jdff dff_A_BdbkCvEe4_0(.dout(w_dff_A_aCSqIg5N2_0),.din(w_dff_A_BdbkCvEe4_0),.clk(gclk));
	jdff dff_A_aCSqIg5N2_0(.dout(w_dff_A_tHWsRnni2_0),.din(w_dff_A_aCSqIg5N2_0),.clk(gclk));
	jdff dff_A_tHWsRnni2_0(.dout(w_dff_A_0Z0SbmFk8_0),.din(w_dff_A_tHWsRnni2_0),.clk(gclk));
	jdff dff_A_0Z0SbmFk8_0(.dout(w_dff_A_eL3TauJW9_0),.din(w_dff_A_0Z0SbmFk8_0),.clk(gclk));
	jdff dff_A_eL3TauJW9_0(.dout(w_dff_A_lu2ZM6HD0_0),.din(w_dff_A_eL3TauJW9_0),.clk(gclk));
	jdff dff_A_lu2ZM6HD0_0(.dout(w_dff_A_SNTgbLB45_0),.din(w_dff_A_lu2ZM6HD0_0),.clk(gclk));
	jdff dff_A_SNTgbLB45_0(.dout(w_dff_A_QK1XmSw77_0),.din(w_dff_A_SNTgbLB45_0),.clk(gclk));
	jdff dff_A_QK1XmSw77_0(.dout(w_dff_A_95mC63sH8_0),.din(w_dff_A_QK1XmSw77_0),.clk(gclk));
	jdff dff_A_95mC63sH8_0(.dout(w_dff_A_Gis0XsyP0_0),.din(w_dff_A_95mC63sH8_0),.clk(gclk));
	jdff dff_A_Gis0XsyP0_0(.dout(w_dff_A_59nN0qvZ8_0),.din(w_dff_A_Gis0XsyP0_0),.clk(gclk));
	jdff dff_A_59nN0qvZ8_0(.dout(w_dff_A_xISAQfzA5_0),.din(w_dff_A_59nN0qvZ8_0),.clk(gclk));
	jdff dff_A_xISAQfzA5_0(.dout(w_dff_A_D5gWjrEs7_0),.din(w_dff_A_xISAQfzA5_0),.clk(gclk));
	jdff dff_A_D5gWjrEs7_0(.dout(w_dff_A_jYe5tZmU6_0),.din(w_dff_A_D5gWjrEs7_0),.clk(gclk));
	jdff dff_A_jYe5tZmU6_0(.dout(w_dff_A_xLRE8IRU5_0),.din(w_dff_A_jYe5tZmU6_0),.clk(gclk));
	jdff dff_A_xLRE8IRU5_0(.dout(w_dff_A_rmI08Fv90_0),.din(w_dff_A_xLRE8IRU5_0),.clk(gclk));
	jdff dff_A_rmI08Fv90_0(.dout(w_dff_A_iyAoaOiS3_0),.din(w_dff_A_rmI08Fv90_0),.clk(gclk));
	jdff dff_A_iyAoaOiS3_0(.dout(w_dff_A_f0ptJyQF8_0),.din(w_dff_A_iyAoaOiS3_0),.clk(gclk));
	jdff dff_A_f0ptJyQF8_0(.dout(w_dff_A_Axi3T5mV9_0),.din(w_dff_A_f0ptJyQF8_0),.clk(gclk));
	jdff dff_A_Axi3T5mV9_0(.dout(w_dff_A_Mslu13Cv9_0),.din(w_dff_A_Axi3T5mV9_0),.clk(gclk));
	jdff dff_A_Mslu13Cv9_0(.dout(G2877gat),.din(w_dff_A_Mslu13Cv9_0),.clk(gclk));
	jdff dff_A_vUFKz7gI5_2(.dout(w_dff_A_1nGxUdwc0_0),.din(w_dff_A_vUFKz7gI5_2),.clk(gclk));
	jdff dff_A_1nGxUdwc0_0(.dout(w_dff_A_k2HBAkGy2_0),.din(w_dff_A_1nGxUdwc0_0),.clk(gclk));
	jdff dff_A_k2HBAkGy2_0(.dout(w_dff_A_zIuU1lhr8_0),.din(w_dff_A_k2HBAkGy2_0),.clk(gclk));
	jdff dff_A_zIuU1lhr8_0(.dout(w_dff_A_Iue0EIvQ9_0),.din(w_dff_A_zIuU1lhr8_0),.clk(gclk));
	jdff dff_A_Iue0EIvQ9_0(.dout(w_dff_A_VmI0LVzu0_0),.din(w_dff_A_Iue0EIvQ9_0),.clk(gclk));
	jdff dff_A_VmI0LVzu0_0(.dout(w_dff_A_r32ypvQj5_0),.din(w_dff_A_VmI0LVzu0_0),.clk(gclk));
	jdff dff_A_r32ypvQj5_0(.dout(w_dff_A_9fQR6I3j3_0),.din(w_dff_A_r32ypvQj5_0),.clk(gclk));
	jdff dff_A_9fQR6I3j3_0(.dout(w_dff_A_dms0CAFp0_0),.din(w_dff_A_9fQR6I3j3_0),.clk(gclk));
	jdff dff_A_dms0CAFp0_0(.dout(w_dff_A_RRdA6QGb9_0),.din(w_dff_A_dms0CAFp0_0),.clk(gclk));
	jdff dff_A_RRdA6QGb9_0(.dout(w_dff_A_2kgG5PXq3_0),.din(w_dff_A_RRdA6QGb9_0),.clk(gclk));
	jdff dff_A_2kgG5PXq3_0(.dout(w_dff_A_xDeq4DB57_0),.din(w_dff_A_2kgG5PXq3_0),.clk(gclk));
	jdff dff_A_xDeq4DB57_0(.dout(w_dff_A_evdO9kTn3_0),.din(w_dff_A_xDeq4DB57_0),.clk(gclk));
	jdff dff_A_evdO9kTn3_0(.dout(w_dff_A_9P5ldShi1_0),.din(w_dff_A_evdO9kTn3_0),.clk(gclk));
	jdff dff_A_9P5ldShi1_0(.dout(w_dff_A_VMtbtwgH4_0),.din(w_dff_A_9P5ldShi1_0),.clk(gclk));
	jdff dff_A_VMtbtwgH4_0(.dout(w_dff_A_5awSSqAp1_0),.din(w_dff_A_VMtbtwgH4_0),.clk(gclk));
	jdff dff_A_5awSSqAp1_0(.dout(w_dff_A_yVS4wdMT3_0),.din(w_dff_A_5awSSqAp1_0),.clk(gclk));
	jdff dff_A_yVS4wdMT3_0(.dout(w_dff_A_7wYmTe2D3_0),.din(w_dff_A_yVS4wdMT3_0),.clk(gclk));
	jdff dff_A_7wYmTe2D3_0(.dout(w_dff_A_ah3ui2GP6_0),.din(w_dff_A_7wYmTe2D3_0),.clk(gclk));
	jdff dff_A_ah3ui2GP6_0(.dout(w_dff_A_kNtpU5qE0_0),.din(w_dff_A_ah3ui2GP6_0),.clk(gclk));
	jdff dff_A_kNtpU5qE0_0(.dout(w_dff_A_P5BwMx4P8_0),.din(w_dff_A_kNtpU5qE0_0),.clk(gclk));
	jdff dff_A_P5BwMx4P8_0(.dout(w_dff_A_zbUnAbP68_0),.din(w_dff_A_P5BwMx4P8_0),.clk(gclk));
	jdff dff_A_zbUnAbP68_0(.dout(w_dff_A_smQS5U6o0_0),.din(w_dff_A_zbUnAbP68_0),.clk(gclk));
	jdff dff_A_smQS5U6o0_0(.dout(w_dff_A_HkbiOc7H2_0),.din(w_dff_A_smQS5U6o0_0),.clk(gclk));
	jdff dff_A_HkbiOc7H2_0(.dout(w_dff_A_98f1L4iL7_0),.din(w_dff_A_HkbiOc7H2_0),.clk(gclk));
	jdff dff_A_98f1L4iL7_0(.dout(w_dff_A_p5ub0H2O5_0),.din(w_dff_A_98f1L4iL7_0),.clk(gclk));
	jdff dff_A_p5ub0H2O5_0(.dout(w_dff_A_ALfQnhZL1_0),.din(w_dff_A_p5ub0H2O5_0),.clk(gclk));
	jdff dff_A_ALfQnhZL1_0(.dout(w_dff_A_0pAenHLj8_0),.din(w_dff_A_ALfQnhZL1_0),.clk(gclk));
	jdff dff_A_0pAenHLj8_0(.dout(w_dff_A_E5Z5407s9_0),.din(w_dff_A_0pAenHLj8_0),.clk(gclk));
	jdff dff_A_E5Z5407s9_0(.dout(w_dff_A_PFF1U29P9_0),.din(w_dff_A_E5Z5407s9_0),.clk(gclk));
	jdff dff_A_PFF1U29P9_0(.dout(w_dff_A_ufi1obGv0_0),.din(w_dff_A_PFF1U29P9_0),.clk(gclk));
	jdff dff_A_ufi1obGv0_0(.dout(w_dff_A_4RIIh9zI9_0),.din(w_dff_A_ufi1obGv0_0),.clk(gclk));
	jdff dff_A_4RIIh9zI9_0(.dout(w_dff_A_hFKqM5e91_0),.din(w_dff_A_4RIIh9zI9_0),.clk(gclk));
	jdff dff_A_hFKqM5e91_0(.dout(w_dff_A_JOQPHkc96_0),.din(w_dff_A_hFKqM5e91_0),.clk(gclk));
	jdff dff_A_JOQPHkc96_0(.dout(w_dff_A_VLkM2l799_0),.din(w_dff_A_JOQPHkc96_0),.clk(gclk));
	jdff dff_A_VLkM2l799_0(.dout(w_dff_A_RSeIIm0c1_0),.din(w_dff_A_VLkM2l799_0),.clk(gclk));
	jdff dff_A_RSeIIm0c1_0(.dout(w_dff_A_QOBVIXpe1_0),.din(w_dff_A_RSeIIm0c1_0),.clk(gclk));
	jdff dff_A_QOBVIXpe1_0(.dout(w_dff_A_T7LNFpVn4_0),.din(w_dff_A_QOBVIXpe1_0),.clk(gclk));
	jdff dff_A_T7LNFpVn4_0(.dout(w_dff_A_6GzhWNzm8_0),.din(w_dff_A_T7LNFpVn4_0),.clk(gclk));
	jdff dff_A_6GzhWNzm8_0(.dout(w_dff_A_PvxLyntL5_0),.din(w_dff_A_6GzhWNzm8_0),.clk(gclk));
	jdff dff_A_PvxLyntL5_0(.dout(w_dff_A_6mtRfzYp9_0),.din(w_dff_A_PvxLyntL5_0),.clk(gclk));
	jdff dff_A_6mtRfzYp9_0(.dout(w_dff_A_PBHcEw8k8_0),.din(w_dff_A_6mtRfzYp9_0),.clk(gclk));
	jdff dff_A_PBHcEw8k8_0(.dout(w_dff_A_zAHplGTV6_0),.din(w_dff_A_PBHcEw8k8_0),.clk(gclk));
	jdff dff_A_zAHplGTV6_0(.dout(w_dff_A_wwhNBayJ5_0),.din(w_dff_A_zAHplGTV6_0),.clk(gclk));
	jdff dff_A_wwhNBayJ5_0(.dout(w_dff_A_MM9i1v2l6_0),.din(w_dff_A_wwhNBayJ5_0),.clk(gclk));
	jdff dff_A_MM9i1v2l6_0(.dout(w_dff_A_hx3XmgLs4_0),.din(w_dff_A_MM9i1v2l6_0),.clk(gclk));
	jdff dff_A_hx3XmgLs4_0(.dout(w_dff_A_1tPG0c9q7_0),.din(w_dff_A_hx3XmgLs4_0),.clk(gclk));
	jdff dff_A_1tPG0c9q7_0(.dout(w_dff_A_5ymGjRTW1_0),.din(w_dff_A_1tPG0c9q7_0),.clk(gclk));
	jdff dff_A_5ymGjRTW1_0(.dout(w_dff_A_VQBN6s995_0),.din(w_dff_A_5ymGjRTW1_0),.clk(gclk));
	jdff dff_A_VQBN6s995_0(.dout(w_dff_A_RqPqsYCC1_0),.din(w_dff_A_VQBN6s995_0),.clk(gclk));
	jdff dff_A_RqPqsYCC1_0(.dout(w_dff_A_0ZYYcHJU3_0),.din(w_dff_A_RqPqsYCC1_0),.clk(gclk));
	jdff dff_A_0ZYYcHJU3_0(.dout(w_dff_A_uT3NRADn6_0),.din(w_dff_A_0ZYYcHJU3_0),.clk(gclk));
	jdff dff_A_uT3NRADn6_0(.dout(w_dff_A_N1ZwoG8s4_0),.din(w_dff_A_uT3NRADn6_0),.clk(gclk));
	jdff dff_A_N1ZwoG8s4_0(.dout(w_dff_A_aiNHm7782_0),.din(w_dff_A_N1ZwoG8s4_0),.clk(gclk));
	jdff dff_A_aiNHm7782_0(.dout(w_dff_A_zMA41CAZ9_0),.din(w_dff_A_aiNHm7782_0),.clk(gclk));
	jdff dff_A_zMA41CAZ9_0(.dout(w_dff_A_sEa4t8eO6_0),.din(w_dff_A_zMA41CAZ9_0),.clk(gclk));
	jdff dff_A_sEa4t8eO6_0(.dout(w_dff_A_NCFPQcXO1_0),.din(w_dff_A_sEa4t8eO6_0),.clk(gclk));
	jdff dff_A_NCFPQcXO1_0(.dout(G3211gat),.din(w_dff_A_NCFPQcXO1_0),.clk(gclk));
	jdff dff_A_x5iNlZpF9_2(.dout(w_dff_A_lYD5SFbp2_0),.din(w_dff_A_x5iNlZpF9_2),.clk(gclk));
	jdff dff_A_lYD5SFbp2_0(.dout(w_dff_A_G7YWsEkZ1_0),.din(w_dff_A_lYD5SFbp2_0),.clk(gclk));
	jdff dff_A_G7YWsEkZ1_0(.dout(w_dff_A_NBync2rf9_0),.din(w_dff_A_G7YWsEkZ1_0),.clk(gclk));
	jdff dff_A_NBync2rf9_0(.dout(w_dff_A_EcTbDsa87_0),.din(w_dff_A_NBync2rf9_0),.clk(gclk));
	jdff dff_A_EcTbDsa87_0(.dout(w_dff_A_t5VhvoHX0_0),.din(w_dff_A_EcTbDsa87_0),.clk(gclk));
	jdff dff_A_t5VhvoHX0_0(.dout(w_dff_A_70OTFWmL8_0),.din(w_dff_A_t5VhvoHX0_0),.clk(gclk));
	jdff dff_A_70OTFWmL8_0(.dout(w_dff_A_vO9UCCjL5_0),.din(w_dff_A_70OTFWmL8_0),.clk(gclk));
	jdff dff_A_vO9UCCjL5_0(.dout(w_dff_A_MppMk7Nq5_0),.din(w_dff_A_vO9UCCjL5_0),.clk(gclk));
	jdff dff_A_MppMk7Nq5_0(.dout(w_dff_A_3rkWYmv03_0),.din(w_dff_A_MppMk7Nq5_0),.clk(gclk));
	jdff dff_A_3rkWYmv03_0(.dout(w_dff_A_3wtYIhbw0_0),.din(w_dff_A_3rkWYmv03_0),.clk(gclk));
	jdff dff_A_3wtYIhbw0_0(.dout(w_dff_A_lgQnK0hh6_0),.din(w_dff_A_3wtYIhbw0_0),.clk(gclk));
	jdff dff_A_lgQnK0hh6_0(.dout(w_dff_A_u2PABcCo6_0),.din(w_dff_A_lgQnK0hh6_0),.clk(gclk));
	jdff dff_A_u2PABcCo6_0(.dout(w_dff_A_45FLl0c18_0),.din(w_dff_A_u2PABcCo6_0),.clk(gclk));
	jdff dff_A_45FLl0c18_0(.dout(w_dff_A_jYK3K8x19_0),.din(w_dff_A_45FLl0c18_0),.clk(gclk));
	jdff dff_A_jYK3K8x19_0(.dout(w_dff_A_wp7RYLUY5_0),.din(w_dff_A_jYK3K8x19_0),.clk(gclk));
	jdff dff_A_wp7RYLUY5_0(.dout(w_dff_A_SLgo7Hm12_0),.din(w_dff_A_wp7RYLUY5_0),.clk(gclk));
	jdff dff_A_SLgo7Hm12_0(.dout(w_dff_A_VR4tcPvC9_0),.din(w_dff_A_SLgo7Hm12_0),.clk(gclk));
	jdff dff_A_VR4tcPvC9_0(.dout(w_dff_A_K3qZg2mx2_0),.din(w_dff_A_VR4tcPvC9_0),.clk(gclk));
	jdff dff_A_K3qZg2mx2_0(.dout(w_dff_A_WcyON9jG0_0),.din(w_dff_A_K3qZg2mx2_0),.clk(gclk));
	jdff dff_A_WcyON9jG0_0(.dout(w_dff_A_fhbtDnig0_0),.din(w_dff_A_WcyON9jG0_0),.clk(gclk));
	jdff dff_A_fhbtDnig0_0(.dout(w_dff_A_SOMJbvNS3_0),.din(w_dff_A_fhbtDnig0_0),.clk(gclk));
	jdff dff_A_SOMJbvNS3_0(.dout(w_dff_A_IbN7RXvn4_0),.din(w_dff_A_SOMJbvNS3_0),.clk(gclk));
	jdff dff_A_IbN7RXvn4_0(.dout(w_dff_A_sKbt3blr9_0),.din(w_dff_A_IbN7RXvn4_0),.clk(gclk));
	jdff dff_A_sKbt3blr9_0(.dout(w_dff_A_rKPQto8e6_0),.din(w_dff_A_sKbt3blr9_0),.clk(gclk));
	jdff dff_A_rKPQto8e6_0(.dout(w_dff_A_iK1BqmU17_0),.din(w_dff_A_rKPQto8e6_0),.clk(gclk));
	jdff dff_A_iK1BqmU17_0(.dout(w_dff_A_JYff3aHV5_0),.din(w_dff_A_iK1BqmU17_0),.clk(gclk));
	jdff dff_A_JYff3aHV5_0(.dout(w_dff_A_6WG55EaU0_0),.din(w_dff_A_JYff3aHV5_0),.clk(gclk));
	jdff dff_A_6WG55EaU0_0(.dout(w_dff_A_z3kkVhEv8_0),.din(w_dff_A_6WG55EaU0_0),.clk(gclk));
	jdff dff_A_z3kkVhEv8_0(.dout(w_dff_A_c3xRUcvx2_0),.din(w_dff_A_z3kkVhEv8_0),.clk(gclk));
	jdff dff_A_c3xRUcvx2_0(.dout(w_dff_A_kIM7Lkv92_0),.din(w_dff_A_c3xRUcvx2_0),.clk(gclk));
	jdff dff_A_kIM7Lkv92_0(.dout(w_dff_A_22NrmKdu1_0),.din(w_dff_A_kIM7Lkv92_0),.clk(gclk));
	jdff dff_A_22NrmKdu1_0(.dout(w_dff_A_bAxytHLF9_0),.din(w_dff_A_22NrmKdu1_0),.clk(gclk));
	jdff dff_A_bAxytHLF9_0(.dout(w_dff_A_ueek6hZa8_0),.din(w_dff_A_bAxytHLF9_0),.clk(gclk));
	jdff dff_A_ueek6hZa8_0(.dout(w_dff_A_PfvWyb6E9_0),.din(w_dff_A_ueek6hZa8_0),.clk(gclk));
	jdff dff_A_PfvWyb6E9_0(.dout(w_dff_A_V38DQqUm1_0),.din(w_dff_A_PfvWyb6E9_0),.clk(gclk));
	jdff dff_A_V38DQqUm1_0(.dout(w_dff_A_YsJxLQ5t5_0),.din(w_dff_A_V38DQqUm1_0),.clk(gclk));
	jdff dff_A_YsJxLQ5t5_0(.dout(w_dff_A_8fpeffk00_0),.din(w_dff_A_YsJxLQ5t5_0),.clk(gclk));
	jdff dff_A_8fpeffk00_0(.dout(w_dff_A_onlsQOkI3_0),.din(w_dff_A_8fpeffk00_0),.clk(gclk));
	jdff dff_A_onlsQOkI3_0(.dout(w_dff_A_sT9b0ne13_0),.din(w_dff_A_onlsQOkI3_0),.clk(gclk));
	jdff dff_A_sT9b0ne13_0(.dout(w_dff_A_8QXdAe2M4_0),.din(w_dff_A_sT9b0ne13_0),.clk(gclk));
	jdff dff_A_8QXdAe2M4_0(.dout(w_dff_A_5ULWgtiY9_0),.din(w_dff_A_8QXdAe2M4_0),.clk(gclk));
	jdff dff_A_5ULWgtiY9_0(.dout(w_dff_A_G0RJgVBj9_0),.din(w_dff_A_5ULWgtiY9_0),.clk(gclk));
	jdff dff_A_G0RJgVBj9_0(.dout(w_dff_A_d9T9VPEA3_0),.din(w_dff_A_G0RJgVBj9_0),.clk(gclk));
	jdff dff_A_d9T9VPEA3_0(.dout(w_dff_A_RNfkP6KG7_0),.din(w_dff_A_d9T9VPEA3_0),.clk(gclk));
	jdff dff_A_RNfkP6KG7_0(.dout(w_dff_A_zy7wlXDR1_0),.din(w_dff_A_RNfkP6KG7_0),.clk(gclk));
	jdff dff_A_zy7wlXDR1_0(.dout(w_dff_A_wA2la3kr3_0),.din(w_dff_A_zy7wlXDR1_0),.clk(gclk));
	jdff dff_A_wA2la3kr3_0(.dout(w_dff_A_mcXzZJOI9_0),.din(w_dff_A_wA2la3kr3_0),.clk(gclk));
	jdff dff_A_mcXzZJOI9_0(.dout(w_dff_A_itegJ70E7_0),.din(w_dff_A_mcXzZJOI9_0),.clk(gclk));
	jdff dff_A_itegJ70E7_0(.dout(w_dff_A_yaabpSOV7_0),.din(w_dff_A_itegJ70E7_0),.clk(gclk));
	jdff dff_A_yaabpSOV7_0(.dout(w_dff_A_Ze7ewDjf8_0),.din(w_dff_A_yaabpSOV7_0),.clk(gclk));
	jdff dff_A_Ze7ewDjf8_0(.dout(w_dff_A_gnTNupHv5_0),.din(w_dff_A_Ze7ewDjf8_0),.clk(gclk));
	jdff dff_A_gnTNupHv5_0(.dout(w_dff_A_ib3Y8QpA0_0),.din(w_dff_A_gnTNupHv5_0),.clk(gclk));
	jdff dff_A_ib3Y8QpA0_0(.dout(w_dff_A_XkuYRI3a5_0),.din(w_dff_A_ib3Y8QpA0_0),.clk(gclk));
	jdff dff_A_XkuYRI3a5_0(.dout(G3552gat),.din(w_dff_A_XkuYRI3a5_0),.clk(gclk));
	jdff dff_A_tlP6TWHP5_2(.dout(w_dff_A_htKEXvld9_0),.din(w_dff_A_tlP6TWHP5_2),.clk(gclk));
	jdff dff_A_htKEXvld9_0(.dout(w_dff_A_eVa3qwvq5_0),.din(w_dff_A_htKEXvld9_0),.clk(gclk));
	jdff dff_A_eVa3qwvq5_0(.dout(w_dff_A_V91giNQZ4_0),.din(w_dff_A_eVa3qwvq5_0),.clk(gclk));
	jdff dff_A_V91giNQZ4_0(.dout(w_dff_A_tiUeNl3k3_0),.din(w_dff_A_V91giNQZ4_0),.clk(gclk));
	jdff dff_A_tiUeNl3k3_0(.dout(w_dff_A_8sAveCFd5_0),.din(w_dff_A_tiUeNl3k3_0),.clk(gclk));
	jdff dff_A_8sAveCFd5_0(.dout(w_dff_A_zNw5rJOg1_0),.din(w_dff_A_8sAveCFd5_0),.clk(gclk));
	jdff dff_A_zNw5rJOg1_0(.dout(w_dff_A_HGobqhKa8_0),.din(w_dff_A_zNw5rJOg1_0),.clk(gclk));
	jdff dff_A_HGobqhKa8_0(.dout(w_dff_A_CPCuflJL8_0),.din(w_dff_A_HGobqhKa8_0),.clk(gclk));
	jdff dff_A_CPCuflJL8_0(.dout(w_dff_A_Y10nIyer7_0),.din(w_dff_A_CPCuflJL8_0),.clk(gclk));
	jdff dff_A_Y10nIyer7_0(.dout(w_dff_A_8N9H7D134_0),.din(w_dff_A_Y10nIyer7_0),.clk(gclk));
	jdff dff_A_8N9H7D134_0(.dout(w_dff_A_hCwHbhsg6_0),.din(w_dff_A_8N9H7D134_0),.clk(gclk));
	jdff dff_A_hCwHbhsg6_0(.dout(w_dff_A_ygr39j160_0),.din(w_dff_A_hCwHbhsg6_0),.clk(gclk));
	jdff dff_A_ygr39j160_0(.dout(w_dff_A_YuP7Jw1q2_0),.din(w_dff_A_ygr39j160_0),.clk(gclk));
	jdff dff_A_YuP7Jw1q2_0(.dout(w_dff_A_TVh0ArG66_0),.din(w_dff_A_YuP7Jw1q2_0),.clk(gclk));
	jdff dff_A_TVh0ArG66_0(.dout(w_dff_A_uyHRBDmb6_0),.din(w_dff_A_TVh0ArG66_0),.clk(gclk));
	jdff dff_A_uyHRBDmb6_0(.dout(w_dff_A_564fWMVj5_0),.din(w_dff_A_uyHRBDmb6_0),.clk(gclk));
	jdff dff_A_564fWMVj5_0(.dout(w_dff_A_EgqQlhWB1_0),.din(w_dff_A_564fWMVj5_0),.clk(gclk));
	jdff dff_A_EgqQlhWB1_0(.dout(w_dff_A_3E5unMHL9_0),.din(w_dff_A_EgqQlhWB1_0),.clk(gclk));
	jdff dff_A_3E5unMHL9_0(.dout(w_dff_A_ELdSFDX40_0),.din(w_dff_A_3E5unMHL9_0),.clk(gclk));
	jdff dff_A_ELdSFDX40_0(.dout(w_dff_A_QxzFyfou2_0),.din(w_dff_A_ELdSFDX40_0),.clk(gclk));
	jdff dff_A_QxzFyfou2_0(.dout(w_dff_A_KjZ2f8T25_0),.din(w_dff_A_QxzFyfou2_0),.clk(gclk));
	jdff dff_A_KjZ2f8T25_0(.dout(w_dff_A_2o5DQ8Mt5_0),.din(w_dff_A_KjZ2f8T25_0),.clk(gclk));
	jdff dff_A_2o5DQ8Mt5_0(.dout(w_dff_A_IH5lNMX90_0),.din(w_dff_A_2o5DQ8Mt5_0),.clk(gclk));
	jdff dff_A_IH5lNMX90_0(.dout(w_dff_A_mu0Z9Cv63_0),.din(w_dff_A_IH5lNMX90_0),.clk(gclk));
	jdff dff_A_mu0Z9Cv63_0(.dout(w_dff_A_hCjLP8dp6_0),.din(w_dff_A_mu0Z9Cv63_0),.clk(gclk));
	jdff dff_A_hCjLP8dp6_0(.dout(w_dff_A_qDwBBmUR1_0),.din(w_dff_A_hCjLP8dp6_0),.clk(gclk));
	jdff dff_A_qDwBBmUR1_0(.dout(w_dff_A_ARlbxat40_0),.din(w_dff_A_qDwBBmUR1_0),.clk(gclk));
	jdff dff_A_ARlbxat40_0(.dout(w_dff_A_GOx0FYBK7_0),.din(w_dff_A_ARlbxat40_0),.clk(gclk));
	jdff dff_A_GOx0FYBK7_0(.dout(w_dff_A_I33b71Kd9_0),.din(w_dff_A_GOx0FYBK7_0),.clk(gclk));
	jdff dff_A_I33b71Kd9_0(.dout(w_dff_A_XKtWoxgP6_0),.din(w_dff_A_I33b71Kd9_0),.clk(gclk));
	jdff dff_A_XKtWoxgP6_0(.dout(w_dff_A_69iJw6Xi4_0),.din(w_dff_A_XKtWoxgP6_0),.clk(gclk));
	jdff dff_A_69iJw6Xi4_0(.dout(w_dff_A_QB7m5PNs8_0),.din(w_dff_A_69iJw6Xi4_0),.clk(gclk));
	jdff dff_A_QB7m5PNs8_0(.dout(w_dff_A_1FxkTZab5_0),.din(w_dff_A_QB7m5PNs8_0),.clk(gclk));
	jdff dff_A_1FxkTZab5_0(.dout(w_dff_A_i5GSygaG3_0),.din(w_dff_A_1FxkTZab5_0),.clk(gclk));
	jdff dff_A_i5GSygaG3_0(.dout(w_dff_A_Bu3knTpj8_0),.din(w_dff_A_i5GSygaG3_0),.clk(gclk));
	jdff dff_A_Bu3knTpj8_0(.dout(w_dff_A_P9d1Losl4_0),.din(w_dff_A_Bu3knTpj8_0),.clk(gclk));
	jdff dff_A_P9d1Losl4_0(.dout(w_dff_A_v3ljCD6s3_0),.din(w_dff_A_P9d1Losl4_0),.clk(gclk));
	jdff dff_A_v3ljCD6s3_0(.dout(w_dff_A_r8lg5iZI1_0),.din(w_dff_A_v3ljCD6s3_0),.clk(gclk));
	jdff dff_A_r8lg5iZI1_0(.dout(w_dff_A_AwGZmeen1_0),.din(w_dff_A_r8lg5iZI1_0),.clk(gclk));
	jdff dff_A_AwGZmeen1_0(.dout(w_dff_A_xx6Hhrow5_0),.din(w_dff_A_AwGZmeen1_0),.clk(gclk));
	jdff dff_A_xx6Hhrow5_0(.dout(w_dff_A_qomTXFr90_0),.din(w_dff_A_xx6Hhrow5_0),.clk(gclk));
	jdff dff_A_qomTXFr90_0(.dout(w_dff_A_DMEN1KHw8_0),.din(w_dff_A_qomTXFr90_0),.clk(gclk));
	jdff dff_A_DMEN1KHw8_0(.dout(w_dff_A_FbkpCx526_0),.din(w_dff_A_DMEN1KHw8_0),.clk(gclk));
	jdff dff_A_FbkpCx526_0(.dout(w_dff_A_yUyw4dIv6_0),.din(w_dff_A_FbkpCx526_0),.clk(gclk));
	jdff dff_A_yUyw4dIv6_0(.dout(w_dff_A_UxWic4sR2_0),.din(w_dff_A_yUyw4dIv6_0),.clk(gclk));
	jdff dff_A_UxWic4sR2_0(.dout(w_dff_A_3uJZLNB75_0),.din(w_dff_A_UxWic4sR2_0),.clk(gclk));
	jdff dff_A_3uJZLNB75_0(.dout(w_dff_A_NtmaUURD2_0),.din(w_dff_A_3uJZLNB75_0),.clk(gclk));
	jdff dff_A_NtmaUURD2_0(.dout(w_dff_A_MFI1bAwp5_0),.din(w_dff_A_NtmaUURD2_0),.clk(gclk));
	jdff dff_A_MFI1bAwp5_0(.dout(w_dff_A_6qzdKOMX1_0),.din(w_dff_A_MFI1bAwp5_0),.clk(gclk));
	jdff dff_A_6qzdKOMX1_0(.dout(w_dff_A_sXErAsAX8_0),.din(w_dff_A_6qzdKOMX1_0),.clk(gclk));
	jdff dff_A_sXErAsAX8_0(.dout(G3895gat),.din(w_dff_A_sXErAsAX8_0),.clk(gclk));
	jdff dff_A_HcHGc8GI5_2(.dout(w_dff_A_qsoH4gB39_0),.din(w_dff_A_HcHGc8GI5_2),.clk(gclk));
	jdff dff_A_qsoH4gB39_0(.dout(w_dff_A_nIP3F0dU4_0),.din(w_dff_A_qsoH4gB39_0),.clk(gclk));
	jdff dff_A_nIP3F0dU4_0(.dout(w_dff_A_fvBVW7Tm8_0),.din(w_dff_A_nIP3F0dU4_0),.clk(gclk));
	jdff dff_A_fvBVW7Tm8_0(.dout(w_dff_A_J8vI6M7I0_0),.din(w_dff_A_fvBVW7Tm8_0),.clk(gclk));
	jdff dff_A_J8vI6M7I0_0(.dout(w_dff_A_sAcLa3sX6_0),.din(w_dff_A_J8vI6M7I0_0),.clk(gclk));
	jdff dff_A_sAcLa3sX6_0(.dout(w_dff_A_E95lJQPi8_0),.din(w_dff_A_sAcLa3sX6_0),.clk(gclk));
	jdff dff_A_E95lJQPi8_0(.dout(w_dff_A_o93XOJ8P1_0),.din(w_dff_A_E95lJQPi8_0),.clk(gclk));
	jdff dff_A_o93XOJ8P1_0(.dout(w_dff_A_40n6Vg5T0_0),.din(w_dff_A_o93XOJ8P1_0),.clk(gclk));
	jdff dff_A_40n6Vg5T0_0(.dout(w_dff_A_dKmeG3aR2_0),.din(w_dff_A_40n6Vg5T0_0),.clk(gclk));
	jdff dff_A_dKmeG3aR2_0(.dout(w_dff_A_AX1nK5VO6_0),.din(w_dff_A_dKmeG3aR2_0),.clk(gclk));
	jdff dff_A_AX1nK5VO6_0(.dout(w_dff_A_se1GDjip4_0),.din(w_dff_A_AX1nK5VO6_0),.clk(gclk));
	jdff dff_A_se1GDjip4_0(.dout(w_dff_A_Mmp8GNwa8_0),.din(w_dff_A_se1GDjip4_0),.clk(gclk));
	jdff dff_A_Mmp8GNwa8_0(.dout(w_dff_A_AYvbEJrm8_0),.din(w_dff_A_Mmp8GNwa8_0),.clk(gclk));
	jdff dff_A_AYvbEJrm8_0(.dout(w_dff_A_CJokU8Jk0_0),.din(w_dff_A_AYvbEJrm8_0),.clk(gclk));
	jdff dff_A_CJokU8Jk0_0(.dout(w_dff_A_nwawaXxH4_0),.din(w_dff_A_CJokU8Jk0_0),.clk(gclk));
	jdff dff_A_nwawaXxH4_0(.dout(w_dff_A_hTsoAsnB1_0),.din(w_dff_A_nwawaXxH4_0),.clk(gclk));
	jdff dff_A_hTsoAsnB1_0(.dout(w_dff_A_0ipCLz0L4_0),.din(w_dff_A_hTsoAsnB1_0),.clk(gclk));
	jdff dff_A_0ipCLz0L4_0(.dout(w_dff_A_UQQq3KWs9_0),.din(w_dff_A_0ipCLz0L4_0),.clk(gclk));
	jdff dff_A_UQQq3KWs9_0(.dout(w_dff_A_ibWbl1Nr1_0),.din(w_dff_A_UQQq3KWs9_0),.clk(gclk));
	jdff dff_A_ibWbl1Nr1_0(.dout(w_dff_A_WV1P5eZ88_0),.din(w_dff_A_ibWbl1Nr1_0),.clk(gclk));
	jdff dff_A_WV1P5eZ88_0(.dout(w_dff_A_nxvAh8NZ1_0),.din(w_dff_A_WV1P5eZ88_0),.clk(gclk));
	jdff dff_A_nxvAh8NZ1_0(.dout(w_dff_A_QhpKQxvp0_0),.din(w_dff_A_nxvAh8NZ1_0),.clk(gclk));
	jdff dff_A_QhpKQxvp0_0(.dout(w_dff_A_Rt0A6Q1L9_0),.din(w_dff_A_QhpKQxvp0_0),.clk(gclk));
	jdff dff_A_Rt0A6Q1L9_0(.dout(w_dff_A_XGf37ncy2_0),.din(w_dff_A_Rt0A6Q1L9_0),.clk(gclk));
	jdff dff_A_XGf37ncy2_0(.dout(w_dff_A_i00ovWSt2_0),.din(w_dff_A_XGf37ncy2_0),.clk(gclk));
	jdff dff_A_i00ovWSt2_0(.dout(w_dff_A_pEuYcoju9_0),.din(w_dff_A_i00ovWSt2_0),.clk(gclk));
	jdff dff_A_pEuYcoju9_0(.dout(w_dff_A_Zn3mKGlE8_0),.din(w_dff_A_pEuYcoju9_0),.clk(gclk));
	jdff dff_A_Zn3mKGlE8_0(.dout(w_dff_A_mUCvp3GE2_0),.din(w_dff_A_Zn3mKGlE8_0),.clk(gclk));
	jdff dff_A_mUCvp3GE2_0(.dout(w_dff_A_9kMotp116_0),.din(w_dff_A_mUCvp3GE2_0),.clk(gclk));
	jdff dff_A_9kMotp116_0(.dout(w_dff_A_adUvZHCo2_0),.din(w_dff_A_9kMotp116_0),.clk(gclk));
	jdff dff_A_adUvZHCo2_0(.dout(w_dff_A_Pk1mll5I8_0),.din(w_dff_A_adUvZHCo2_0),.clk(gclk));
	jdff dff_A_Pk1mll5I8_0(.dout(w_dff_A_0z0MehKw5_0),.din(w_dff_A_Pk1mll5I8_0),.clk(gclk));
	jdff dff_A_0z0MehKw5_0(.dout(w_dff_A_UMdm7bR86_0),.din(w_dff_A_0z0MehKw5_0),.clk(gclk));
	jdff dff_A_UMdm7bR86_0(.dout(w_dff_A_WXZ0mLsa1_0),.din(w_dff_A_UMdm7bR86_0),.clk(gclk));
	jdff dff_A_WXZ0mLsa1_0(.dout(w_dff_A_Eh13WoxW3_0),.din(w_dff_A_WXZ0mLsa1_0),.clk(gclk));
	jdff dff_A_Eh13WoxW3_0(.dout(w_dff_A_6SluiaN89_0),.din(w_dff_A_Eh13WoxW3_0),.clk(gclk));
	jdff dff_A_6SluiaN89_0(.dout(w_dff_A_lxDaDdos1_0),.din(w_dff_A_6SluiaN89_0),.clk(gclk));
	jdff dff_A_lxDaDdos1_0(.dout(w_dff_A_6wMztMHk8_0),.din(w_dff_A_lxDaDdos1_0),.clk(gclk));
	jdff dff_A_6wMztMHk8_0(.dout(w_dff_A_44cAN4210_0),.din(w_dff_A_6wMztMHk8_0),.clk(gclk));
	jdff dff_A_44cAN4210_0(.dout(w_dff_A_UxijUgdI0_0),.din(w_dff_A_44cAN4210_0),.clk(gclk));
	jdff dff_A_UxijUgdI0_0(.dout(w_dff_A_ArdSPo6G5_0),.din(w_dff_A_UxijUgdI0_0),.clk(gclk));
	jdff dff_A_ArdSPo6G5_0(.dout(w_dff_A_v5Xyjrb10_0),.din(w_dff_A_ArdSPo6G5_0),.clk(gclk));
	jdff dff_A_v5Xyjrb10_0(.dout(w_dff_A_h1Wl5xaf7_0),.din(w_dff_A_v5Xyjrb10_0),.clk(gclk));
	jdff dff_A_h1Wl5xaf7_0(.dout(w_dff_A_JAvxWtIC6_0),.din(w_dff_A_h1Wl5xaf7_0),.clk(gclk));
	jdff dff_A_JAvxWtIC6_0(.dout(w_dff_A_EZQkrqlz6_0),.din(w_dff_A_JAvxWtIC6_0),.clk(gclk));
	jdff dff_A_EZQkrqlz6_0(.dout(w_dff_A_LGB74pSN9_0),.din(w_dff_A_EZQkrqlz6_0),.clk(gclk));
	jdff dff_A_LGB74pSN9_0(.dout(w_dff_A_F13iuZHC0_0),.din(w_dff_A_LGB74pSN9_0),.clk(gclk));
	jdff dff_A_F13iuZHC0_0(.dout(G4241gat),.din(w_dff_A_F13iuZHC0_0),.clk(gclk));
	jdff dff_A_Z99VGWH31_2(.dout(w_dff_A_0rPlNvCR0_0),.din(w_dff_A_Z99VGWH31_2),.clk(gclk));
	jdff dff_A_0rPlNvCR0_0(.dout(w_dff_A_4At6yBK88_0),.din(w_dff_A_0rPlNvCR0_0),.clk(gclk));
	jdff dff_A_4At6yBK88_0(.dout(w_dff_A_E1mn4PEJ2_0),.din(w_dff_A_4At6yBK88_0),.clk(gclk));
	jdff dff_A_E1mn4PEJ2_0(.dout(w_dff_A_HGjQL6Jk6_0),.din(w_dff_A_E1mn4PEJ2_0),.clk(gclk));
	jdff dff_A_HGjQL6Jk6_0(.dout(w_dff_A_yY0quIV29_0),.din(w_dff_A_HGjQL6Jk6_0),.clk(gclk));
	jdff dff_A_yY0quIV29_0(.dout(w_dff_A_mQUd3zN64_0),.din(w_dff_A_yY0quIV29_0),.clk(gclk));
	jdff dff_A_mQUd3zN64_0(.dout(w_dff_A_os0rrg7F4_0),.din(w_dff_A_mQUd3zN64_0),.clk(gclk));
	jdff dff_A_os0rrg7F4_0(.dout(w_dff_A_xei5nxWQ3_0),.din(w_dff_A_os0rrg7F4_0),.clk(gclk));
	jdff dff_A_xei5nxWQ3_0(.dout(w_dff_A_ic61KOAc0_0),.din(w_dff_A_xei5nxWQ3_0),.clk(gclk));
	jdff dff_A_ic61KOAc0_0(.dout(w_dff_A_ebianqhH1_0),.din(w_dff_A_ic61KOAc0_0),.clk(gclk));
	jdff dff_A_ebianqhH1_0(.dout(w_dff_A_PLZnnfak3_0),.din(w_dff_A_ebianqhH1_0),.clk(gclk));
	jdff dff_A_PLZnnfak3_0(.dout(w_dff_A_P5xy79OU0_0),.din(w_dff_A_PLZnnfak3_0),.clk(gclk));
	jdff dff_A_P5xy79OU0_0(.dout(w_dff_A_1YcfwdP87_0),.din(w_dff_A_P5xy79OU0_0),.clk(gclk));
	jdff dff_A_1YcfwdP87_0(.dout(w_dff_A_ra44eOUw8_0),.din(w_dff_A_1YcfwdP87_0),.clk(gclk));
	jdff dff_A_ra44eOUw8_0(.dout(w_dff_A_Fj8Eu6e52_0),.din(w_dff_A_ra44eOUw8_0),.clk(gclk));
	jdff dff_A_Fj8Eu6e52_0(.dout(w_dff_A_kIdF5RLh9_0),.din(w_dff_A_Fj8Eu6e52_0),.clk(gclk));
	jdff dff_A_kIdF5RLh9_0(.dout(w_dff_A_6EO4qM4U7_0),.din(w_dff_A_kIdF5RLh9_0),.clk(gclk));
	jdff dff_A_6EO4qM4U7_0(.dout(w_dff_A_sWLnCkTn6_0),.din(w_dff_A_6EO4qM4U7_0),.clk(gclk));
	jdff dff_A_sWLnCkTn6_0(.dout(w_dff_A_kmsaJNrm5_0),.din(w_dff_A_sWLnCkTn6_0),.clk(gclk));
	jdff dff_A_kmsaJNrm5_0(.dout(w_dff_A_fwtl1zsk6_0),.din(w_dff_A_kmsaJNrm5_0),.clk(gclk));
	jdff dff_A_fwtl1zsk6_0(.dout(w_dff_A_qlvSIQUw9_0),.din(w_dff_A_fwtl1zsk6_0),.clk(gclk));
	jdff dff_A_qlvSIQUw9_0(.dout(w_dff_A_poZbm5i38_0),.din(w_dff_A_qlvSIQUw9_0),.clk(gclk));
	jdff dff_A_poZbm5i38_0(.dout(w_dff_A_CcAktltv3_0),.din(w_dff_A_poZbm5i38_0),.clk(gclk));
	jdff dff_A_CcAktltv3_0(.dout(w_dff_A_g9DfIthW7_0),.din(w_dff_A_CcAktltv3_0),.clk(gclk));
	jdff dff_A_g9DfIthW7_0(.dout(w_dff_A_DItL0nNR3_0),.din(w_dff_A_g9DfIthW7_0),.clk(gclk));
	jdff dff_A_DItL0nNR3_0(.dout(w_dff_A_fWc5zKYH5_0),.din(w_dff_A_DItL0nNR3_0),.clk(gclk));
	jdff dff_A_fWc5zKYH5_0(.dout(w_dff_A_rppv83j64_0),.din(w_dff_A_fWc5zKYH5_0),.clk(gclk));
	jdff dff_A_rppv83j64_0(.dout(w_dff_A_iQGHrDZj3_0),.din(w_dff_A_rppv83j64_0),.clk(gclk));
	jdff dff_A_iQGHrDZj3_0(.dout(w_dff_A_Mk6r4eNl7_0),.din(w_dff_A_iQGHrDZj3_0),.clk(gclk));
	jdff dff_A_Mk6r4eNl7_0(.dout(w_dff_A_ZZ646FKw6_0),.din(w_dff_A_Mk6r4eNl7_0),.clk(gclk));
	jdff dff_A_ZZ646FKw6_0(.dout(w_dff_A_ZBHma7Vm9_0),.din(w_dff_A_ZZ646FKw6_0),.clk(gclk));
	jdff dff_A_ZBHma7Vm9_0(.dout(w_dff_A_XZgMTY9c5_0),.din(w_dff_A_ZBHma7Vm9_0),.clk(gclk));
	jdff dff_A_XZgMTY9c5_0(.dout(w_dff_A_wAhbELF39_0),.din(w_dff_A_XZgMTY9c5_0),.clk(gclk));
	jdff dff_A_wAhbELF39_0(.dout(w_dff_A_YtxxQRmc1_0),.din(w_dff_A_wAhbELF39_0),.clk(gclk));
	jdff dff_A_YtxxQRmc1_0(.dout(w_dff_A_bABEPoPm6_0),.din(w_dff_A_YtxxQRmc1_0),.clk(gclk));
	jdff dff_A_bABEPoPm6_0(.dout(w_dff_A_278nQgmT9_0),.din(w_dff_A_bABEPoPm6_0),.clk(gclk));
	jdff dff_A_278nQgmT9_0(.dout(w_dff_A_mzMs0Jyu8_0),.din(w_dff_A_278nQgmT9_0),.clk(gclk));
	jdff dff_A_mzMs0Jyu8_0(.dout(w_dff_A_cEKN8g9d7_0),.din(w_dff_A_mzMs0Jyu8_0),.clk(gclk));
	jdff dff_A_cEKN8g9d7_0(.dout(w_dff_A_PPydyZsY3_0),.din(w_dff_A_cEKN8g9d7_0),.clk(gclk));
	jdff dff_A_PPydyZsY3_0(.dout(w_dff_A_L6jSa4y59_0),.din(w_dff_A_PPydyZsY3_0),.clk(gclk));
	jdff dff_A_L6jSa4y59_0(.dout(w_dff_A_0ijJLyNe7_0),.din(w_dff_A_L6jSa4y59_0),.clk(gclk));
	jdff dff_A_0ijJLyNe7_0(.dout(w_dff_A_zvxYt7Tv4_0),.din(w_dff_A_0ijJLyNe7_0),.clk(gclk));
	jdff dff_A_zvxYt7Tv4_0(.dout(w_dff_A_LYTHLc343_0),.din(w_dff_A_zvxYt7Tv4_0),.clk(gclk));
	jdff dff_A_LYTHLc343_0(.dout(w_dff_A_vilZNmuY8_0),.din(w_dff_A_LYTHLc343_0),.clk(gclk));
	jdff dff_A_vilZNmuY8_0(.dout(G4591gat),.din(w_dff_A_vilZNmuY8_0),.clk(gclk));
	jdff dff_A_afeJhXAY4_2(.dout(w_dff_A_KLSSrEtu1_0),.din(w_dff_A_afeJhXAY4_2),.clk(gclk));
	jdff dff_A_KLSSrEtu1_0(.dout(w_dff_A_gHp6ahtl2_0),.din(w_dff_A_KLSSrEtu1_0),.clk(gclk));
	jdff dff_A_gHp6ahtl2_0(.dout(w_dff_A_Mg8zQyCk3_0),.din(w_dff_A_gHp6ahtl2_0),.clk(gclk));
	jdff dff_A_Mg8zQyCk3_0(.dout(w_dff_A_TlomVDoF6_0),.din(w_dff_A_Mg8zQyCk3_0),.clk(gclk));
	jdff dff_A_TlomVDoF6_0(.dout(w_dff_A_Alvdk1Bo6_0),.din(w_dff_A_TlomVDoF6_0),.clk(gclk));
	jdff dff_A_Alvdk1Bo6_0(.dout(w_dff_A_yoZXois07_0),.din(w_dff_A_Alvdk1Bo6_0),.clk(gclk));
	jdff dff_A_yoZXois07_0(.dout(w_dff_A_EAAkAPMg0_0),.din(w_dff_A_yoZXois07_0),.clk(gclk));
	jdff dff_A_EAAkAPMg0_0(.dout(w_dff_A_fyOO9pcj6_0),.din(w_dff_A_EAAkAPMg0_0),.clk(gclk));
	jdff dff_A_fyOO9pcj6_0(.dout(w_dff_A_wcYj8kzg4_0),.din(w_dff_A_fyOO9pcj6_0),.clk(gclk));
	jdff dff_A_wcYj8kzg4_0(.dout(w_dff_A_jpQoDH987_0),.din(w_dff_A_wcYj8kzg4_0),.clk(gclk));
	jdff dff_A_jpQoDH987_0(.dout(w_dff_A_SMa2VANT8_0),.din(w_dff_A_jpQoDH987_0),.clk(gclk));
	jdff dff_A_SMa2VANT8_0(.dout(w_dff_A_uOgRbNDV4_0),.din(w_dff_A_SMa2VANT8_0),.clk(gclk));
	jdff dff_A_uOgRbNDV4_0(.dout(w_dff_A_wkrWorlu6_0),.din(w_dff_A_uOgRbNDV4_0),.clk(gclk));
	jdff dff_A_wkrWorlu6_0(.dout(w_dff_A_05lb2NUr1_0),.din(w_dff_A_wkrWorlu6_0),.clk(gclk));
	jdff dff_A_05lb2NUr1_0(.dout(w_dff_A_0c39Pvsv8_0),.din(w_dff_A_05lb2NUr1_0),.clk(gclk));
	jdff dff_A_0c39Pvsv8_0(.dout(w_dff_A_ZqlMTaoa4_0),.din(w_dff_A_0c39Pvsv8_0),.clk(gclk));
	jdff dff_A_ZqlMTaoa4_0(.dout(w_dff_A_GCcWrlU12_0),.din(w_dff_A_ZqlMTaoa4_0),.clk(gclk));
	jdff dff_A_GCcWrlU12_0(.dout(w_dff_A_KqbgoRB20_0),.din(w_dff_A_GCcWrlU12_0),.clk(gclk));
	jdff dff_A_KqbgoRB20_0(.dout(w_dff_A_WHoVlYTy2_0),.din(w_dff_A_KqbgoRB20_0),.clk(gclk));
	jdff dff_A_WHoVlYTy2_0(.dout(w_dff_A_rVpqoafh9_0),.din(w_dff_A_WHoVlYTy2_0),.clk(gclk));
	jdff dff_A_rVpqoafh9_0(.dout(w_dff_A_bzX8rOTV5_0),.din(w_dff_A_rVpqoafh9_0),.clk(gclk));
	jdff dff_A_bzX8rOTV5_0(.dout(w_dff_A_NzWoy8JQ3_0),.din(w_dff_A_bzX8rOTV5_0),.clk(gclk));
	jdff dff_A_NzWoy8JQ3_0(.dout(w_dff_A_vWijRKai2_0),.din(w_dff_A_NzWoy8JQ3_0),.clk(gclk));
	jdff dff_A_vWijRKai2_0(.dout(w_dff_A_1E1qQpmS1_0),.din(w_dff_A_vWijRKai2_0),.clk(gclk));
	jdff dff_A_1E1qQpmS1_0(.dout(w_dff_A_JJmaRRDd6_0),.din(w_dff_A_1E1qQpmS1_0),.clk(gclk));
	jdff dff_A_JJmaRRDd6_0(.dout(w_dff_A_T3WsZX3e0_0),.din(w_dff_A_JJmaRRDd6_0),.clk(gclk));
	jdff dff_A_T3WsZX3e0_0(.dout(w_dff_A_FN4zFvGm2_0),.din(w_dff_A_T3WsZX3e0_0),.clk(gclk));
	jdff dff_A_FN4zFvGm2_0(.dout(w_dff_A_Q9Wf0lyB1_0),.din(w_dff_A_FN4zFvGm2_0),.clk(gclk));
	jdff dff_A_Q9Wf0lyB1_0(.dout(w_dff_A_SRBgKef43_0),.din(w_dff_A_Q9Wf0lyB1_0),.clk(gclk));
	jdff dff_A_SRBgKef43_0(.dout(w_dff_A_7858yQTM7_0),.din(w_dff_A_SRBgKef43_0),.clk(gclk));
	jdff dff_A_7858yQTM7_0(.dout(w_dff_A_wCVTmF9v6_0),.din(w_dff_A_7858yQTM7_0),.clk(gclk));
	jdff dff_A_wCVTmF9v6_0(.dout(w_dff_A_wLUv0HrY8_0),.din(w_dff_A_wCVTmF9v6_0),.clk(gclk));
	jdff dff_A_wLUv0HrY8_0(.dout(w_dff_A_Ac974i1p7_0),.din(w_dff_A_wLUv0HrY8_0),.clk(gclk));
	jdff dff_A_Ac974i1p7_0(.dout(w_dff_A_TNvEFM7X6_0),.din(w_dff_A_Ac974i1p7_0),.clk(gclk));
	jdff dff_A_TNvEFM7X6_0(.dout(w_dff_A_vus6YOYj3_0),.din(w_dff_A_TNvEFM7X6_0),.clk(gclk));
	jdff dff_A_vus6YOYj3_0(.dout(w_dff_A_RqfofxOU4_0),.din(w_dff_A_vus6YOYj3_0),.clk(gclk));
	jdff dff_A_RqfofxOU4_0(.dout(w_dff_A_DZQwGa1a9_0),.din(w_dff_A_RqfofxOU4_0),.clk(gclk));
	jdff dff_A_DZQwGa1a9_0(.dout(w_dff_A_0fvfonUl5_0),.din(w_dff_A_DZQwGa1a9_0),.clk(gclk));
	jdff dff_A_0fvfonUl5_0(.dout(w_dff_A_Lp5wsFC31_0),.din(w_dff_A_0fvfonUl5_0),.clk(gclk));
	jdff dff_A_Lp5wsFC31_0(.dout(w_dff_A_JV1KtkJ67_0),.din(w_dff_A_Lp5wsFC31_0),.clk(gclk));
	jdff dff_A_JV1KtkJ67_0(.dout(w_dff_A_eRseWFyr5_0),.din(w_dff_A_JV1KtkJ67_0),.clk(gclk));
	jdff dff_A_eRseWFyr5_0(.dout(G4946gat),.din(w_dff_A_eRseWFyr5_0),.clk(gclk));
	jdff dff_A_FoMYUxYC3_2(.dout(w_dff_A_gnvhzIGn4_0),.din(w_dff_A_FoMYUxYC3_2),.clk(gclk));
	jdff dff_A_gnvhzIGn4_0(.dout(w_dff_A_6izX916a9_0),.din(w_dff_A_gnvhzIGn4_0),.clk(gclk));
	jdff dff_A_6izX916a9_0(.dout(w_dff_A_AcjGaaqB8_0),.din(w_dff_A_6izX916a9_0),.clk(gclk));
	jdff dff_A_AcjGaaqB8_0(.dout(w_dff_A_qUUaUic41_0),.din(w_dff_A_AcjGaaqB8_0),.clk(gclk));
	jdff dff_A_qUUaUic41_0(.dout(w_dff_A_9HfdYidC8_0),.din(w_dff_A_qUUaUic41_0),.clk(gclk));
	jdff dff_A_9HfdYidC8_0(.dout(w_dff_A_JdxyEs2o2_0),.din(w_dff_A_9HfdYidC8_0),.clk(gclk));
	jdff dff_A_JdxyEs2o2_0(.dout(w_dff_A_g929yfn40_0),.din(w_dff_A_JdxyEs2o2_0),.clk(gclk));
	jdff dff_A_g929yfn40_0(.dout(w_dff_A_jEPR9xl32_0),.din(w_dff_A_g929yfn40_0),.clk(gclk));
	jdff dff_A_jEPR9xl32_0(.dout(w_dff_A_q00CaeYe8_0),.din(w_dff_A_jEPR9xl32_0),.clk(gclk));
	jdff dff_A_q00CaeYe8_0(.dout(w_dff_A_KB3E3Z3z5_0),.din(w_dff_A_q00CaeYe8_0),.clk(gclk));
	jdff dff_A_KB3E3Z3z5_0(.dout(w_dff_A_bu7JjBvx2_0),.din(w_dff_A_KB3E3Z3z5_0),.clk(gclk));
	jdff dff_A_bu7JjBvx2_0(.dout(w_dff_A_XAjSpPdI0_0),.din(w_dff_A_bu7JjBvx2_0),.clk(gclk));
	jdff dff_A_XAjSpPdI0_0(.dout(w_dff_A_2kz2U6hn6_0),.din(w_dff_A_XAjSpPdI0_0),.clk(gclk));
	jdff dff_A_2kz2U6hn6_0(.dout(w_dff_A_LLCGoYyS9_0),.din(w_dff_A_2kz2U6hn6_0),.clk(gclk));
	jdff dff_A_LLCGoYyS9_0(.dout(w_dff_A_WSdTx86Z0_0),.din(w_dff_A_LLCGoYyS9_0),.clk(gclk));
	jdff dff_A_WSdTx86Z0_0(.dout(w_dff_A_eOtDSeHO8_0),.din(w_dff_A_WSdTx86Z0_0),.clk(gclk));
	jdff dff_A_eOtDSeHO8_0(.dout(w_dff_A_lwQvF2y68_0),.din(w_dff_A_eOtDSeHO8_0),.clk(gclk));
	jdff dff_A_lwQvF2y68_0(.dout(w_dff_A_ltxo5Jfm3_0),.din(w_dff_A_lwQvF2y68_0),.clk(gclk));
	jdff dff_A_ltxo5Jfm3_0(.dout(w_dff_A_jDGWNsFa2_0),.din(w_dff_A_ltxo5Jfm3_0),.clk(gclk));
	jdff dff_A_jDGWNsFa2_0(.dout(w_dff_A_c6iRBxs45_0),.din(w_dff_A_jDGWNsFa2_0),.clk(gclk));
	jdff dff_A_c6iRBxs45_0(.dout(w_dff_A_X5CZYujQ6_0),.din(w_dff_A_c6iRBxs45_0),.clk(gclk));
	jdff dff_A_X5CZYujQ6_0(.dout(w_dff_A_rcVE5MdU7_0),.din(w_dff_A_X5CZYujQ6_0),.clk(gclk));
	jdff dff_A_rcVE5MdU7_0(.dout(w_dff_A_z0GMMdU54_0),.din(w_dff_A_rcVE5MdU7_0),.clk(gclk));
	jdff dff_A_z0GMMdU54_0(.dout(w_dff_A_FTnuWQEh9_0),.din(w_dff_A_z0GMMdU54_0),.clk(gclk));
	jdff dff_A_FTnuWQEh9_0(.dout(w_dff_A_fE3fl2JK8_0),.din(w_dff_A_FTnuWQEh9_0),.clk(gclk));
	jdff dff_A_fE3fl2JK8_0(.dout(w_dff_A_rRNZePuO7_0),.din(w_dff_A_fE3fl2JK8_0),.clk(gclk));
	jdff dff_A_rRNZePuO7_0(.dout(w_dff_A_d9OqFF5V7_0),.din(w_dff_A_rRNZePuO7_0),.clk(gclk));
	jdff dff_A_d9OqFF5V7_0(.dout(w_dff_A_etJLtNuo9_0),.din(w_dff_A_d9OqFF5V7_0),.clk(gclk));
	jdff dff_A_etJLtNuo9_0(.dout(w_dff_A_lHIzLgsf4_0),.din(w_dff_A_etJLtNuo9_0),.clk(gclk));
	jdff dff_A_lHIzLgsf4_0(.dout(w_dff_A_go9bXObM4_0),.din(w_dff_A_lHIzLgsf4_0),.clk(gclk));
	jdff dff_A_go9bXObM4_0(.dout(w_dff_A_0onAaVvQ7_0),.din(w_dff_A_go9bXObM4_0),.clk(gclk));
	jdff dff_A_0onAaVvQ7_0(.dout(w_dff_A_4TGbiVYl3_0),.din(w_dff_A_0onAaVvQ7_0),.clk(gclk));
	jdff dff_A_4TGbiVYl3_0(.dout(w_dff_A_GaMGoxSt0_0),.din(w_dff_A_4TGbiVYl3_0),.clk(gclk));
	jdff dff_A_GaMGoxSt0_0(.dout(w_dff_A_mYNbI0pB0_0),.din(w_dff_A_GaMGoxSt0_0),.clk(gclk));
	jdff dff_A_mYNbI0pB0_0(.dout(w_dff_A_PSrvcFwT1_0),.din(w_dff_A_mYNbI0pB0_0),.clk(gclk));
	jdff dff_A_PSrvcFwT1_0(.dout(w_dff_A_jEqiU7ii3_0),.din(w_dff_A_PSrvcFwT1_0),.clk(gclk));
	jdff dff_A_jEqiU7ii3_0(.dout(w_dff_A_T8rXtJu05_0),.din(w_dff_A_jEqiU7ii3_0),.clk(gclk));
	jdff dff_A_T8rXtJu05_0(.dout(w_dff_A_8G1VuqpI6_0),.din(w_dff_A_T8rXtJu05_0),.clk(gclk));
	jdff dff_A_8G1VuqpI6_0(.dout(G5308gat),.din(w_dff_A_8G1VuqpI6_0),.clk(gclk));
	jdff dff_A_GmHJ0a9t0_2(.dout(w_dff_A_dSbbVZ3o7_0),.din(w_dff_A_GmHJ0a9t0_2),.clk(gclk));
	jdff dff_A_dSbbVZ3o7_0(.dout(w_dff_A_NZPOisht3_0),.din(w_dff_A_dSbbVZ3o7_0),.clk(gclk));
	jdff dff_A_NZPOisht3_0(.dout(w_dff_A_SAjOOS886_0),.din(w_dff_A_NZPOisht3_0),.clk(gclk));
	jdff dff_A_SAjOOS886_0(.dout(w_dff_A_W8kKom7e5_0),.din(w_dff_A_SAjOOS886_0),.clk(gclk));
	jdff dff_A_W8kKom7e5_0(.dout(w_dff_A_kWZP04ST6_0),.din(w_dff_A_W8kKom7e5_0),.clk(gclk));
	jdff dff_A_kWZP04ST6_0(.dout(w_dff_A_sbdJc6K36_0),.din(w_dff_A_kWZP04ST6_0),.clk(gclk));
	jdff dff_A_sbdJc6K36_0(.dout(w_dff_A_X4T6FdVr5_0),.din(w_dff_A_sbdJc6K36_0),.clk(gclk));
	jdff dff_A_X4T6FdVr5_0(.dout(w_dff_A_RmsVUeVX5_0),.din(w_dff_A_X4T6FdVr5_0),.clk(gclk));
	jdff dff_A_RmsVUeVX5_0(.dout(w_dff_A_YkMKAMDb1_0),.din(w_dff_A_RmsVUeVX5_0),.clk(gclk));
	jdff dff_A_YkMKAMDb1_0(.dout(w_dff_A_MPxEYMBQ5_0),.din(w_dff_A_YkMKAMDb1_0),.clk(gclk));
	jdff dff_A_MPxEYMBQ5_0(.dout(w_dff_A_Rs20P8xn1_0),.din(w_dff_A_MPxEYMBQ5_0),.clk(gclk));
	jdff dff_A_Rs20P8xn1_0(.dout(w_dff_A_dPHorXnj0_0),.din(w_dff_A_Rs20P8xn1_0),.clk(gclk));
	jdff dff_A_dPHorXnj0_0(.dout(w_dff_A_yzyNEFai1_0),.din(w_dff_A_dPHorXnj0_0),.clk(gclk));
	jdff dff_A_yzyNEFai1_0(.dout(w_dff_A_xwzNulXl4_0),.din(w_dff_A_yzyNEFai1_0),.clk(gclk));
	jdff dff_A_xwzNulXl4_0(.dout(w_dff_A_ZkaOgzgl6_0),.din(w_dff_A_xwzNulXl4_0),.clk(gclk));
	jdff dff_A_ZkaOgzgl6_0(.dout(w_dff_A_VKmschiw8_0),.din(w_dff_A_ZkaOgzgl6_0),.clk(gclk));
	jdff dff_A_VKmschiw8_0(.dout(w_dff_A_HtKEXHjw5_0),.din(w_dff_A_VKmschiw8_0),.clk(gclk));
	jdff dff_A_HtKEXHjw5_0(.dout(w_dff_A_UhL7JSLh0_0),.din(w_dff_A_HtKEXHjw5_0),.clk(gclk));
	jdff dff_A_UhL7JSLh0_0(.dout(w_dff_A_tdiJykEE2_0),.din(w_dff_A_UhL7JSLh0_0),.clk(gclk));
	jdff dff_A_tdiJykEE2_0(.dout(w_dff_A_cvEEGpoF9_0),.din(w_dff_A_tdiJykEE2_0),.clk(gclk));
	jdff dff_A_cvEEGpoF9_0(.dout(w_dff_A_Q9JFcfxe0_0),.din(w_dff_A_cvEEGpoF9_0),.clk(gclk));
	jdff dff_A_Q9JFcfxe0_0(.dout(w_dff_A_VvpZKsHW0_0),.din(w_dff_A_Q9JFcfxe0_0),.clk(gclk));
	jdff dff_A_VvpZKsHW0_0(.dout(w_dff_A_R2k5lUdt0_0),.din(w_dff_A_VvpZKsHW0_0),.clk(gclk));
	jdff dff_A_R2k5lUdt0_0(.dout(w_dff_A_YbcYynJs9_0),.din(w_dff_A_R2k5lUdt0_0),.clk(gclk));
	jdff dff_A_YbcYynJs9_0(.dout(w_dff_A_t3ukUg8n0_0),.din(w_dff_A_YbcYynJs9_0),.clk(gclk));
	jdff dff_A_t3ukUg8n0_0(.dout(w_dff_A_hP5cGmAH5_0),.din(w_dff_A_t3ukUg8n0_0),.clk(gclk));
	jdff dff_A_hP5cGmAH5_0(.dout(w_dff_A_sW38N8fZ8_0),.din(w_dff_A_hP5cGmAH5_0),.clk(gclk));
	jdff dff_A_sW38N8fZ8_0(.dout(w_dff_A_nzYRjUJx3_0),.din(w_dff_A_sW38N8fZ8_0),.clk(gclk));
	jdff dff_A_nzYRjUJx3_0(.dout(w_dff_A_sD7fZ1M95_0),.din(w_dff_A_nzYRjUJx3_0),.clk(gclk));
	jdff dff_A_sD7fZ1M95_0(.dout(w_dff_A_QlQYNq4Y4_0),.din(w_dff_A_sD7fZ1M95_0),.clk(gclk));
	jdff dff_A_QlQYNq4Y4_0(.dout(w_dff_A_qCfFwf2z5_0),.din(w_dff_A_QlQYNq4Y4_0),.clk(gclk));
	jdff dff_A_qCfFwf2z5_0(.dout(w_dff_A_bXDfj5za1_0),.din(w_dff_A_qCfFwf2z5_0),.clk(gclk));
	jdff dff_A_bXDfj5za1_0(.dout(w_dff_A_yu9252Xt7_0),.din(w_dff_A_bXDfj5za1_0),.clk(gclk));
	jdff dff_A_yu9252Xt7_0(.dout(w_dff_A_JBT4MzeO3_0),.din(w_dff_A_yu9252Xt7_0),.clk(gclk));
	jdff dff_A_JBT4MzeO3_0(.dout(w_dff_A_XOBfWwGa2_0),.din(w_dff_A_JBT4MzeO3_0),.clk(gclk));
	jdff dff_A_XOBfWwGa2_0(.dout(G5672gat),.din(w_dff_A_XOBfWwGa2_0),.clk(gclk));
	jdff dff_A_XaMEPoS81_2(.dout(w_dff_A_5QF3iZPZ9_0),.din(w_dff_A_XaMEPoS81_2),.clk(gclk));
	jdff dff_A_5QF3iZPZ9_0(.dout(w_dff_A_bQLsF19t0_0),.din(w_dff_A_5QF3iZPZ9_0),.clk(gclk));
	jdff dff_A_bQLsF19t0_0(.dout(w_dff_A_NBDITLYh6_0),.din(w_dff_A_bQLsF19t0_0),.clk(gclk));
	jdff dff_A_NBDITLYh6_0(.dout(w_dff_A_qiwKXeqI2_0),.din(w_dff_A_NBDITLYh6_0),.clk(gclk));
	jdff dff_A_qiwKXeqI2_0(.dout(w_dff_A_OZcaRXYt3_0),.din(w_dff_A_qiwKXeqI2_0),.clk(gclk));
	jdff dff_A_OZcaRXYt3_0(.dout(w_dff_A_qjGaneWF7_0),.din(w_dff_A_OZcaRXYt3_0),.clk(gclk));
	jdff dff_A_qjGaneWF7_0(.dout(w_dff_A_1YLz3UET5_0),.din(w_dff_A_qjGaneWF7_0),.clk(gclk));
	jdff dff_A_1YLz3UET5_0(.dout(w_dff_A_u7LQ7PlU6_0),.din(w_dff_A_1YLz3UET5_0),.clk(gclk));
	jdff dff_A_u7LQ7PlU6_0(.dout(w_dff_A_V20hFW2X6_0),.din(w_dff_A_u7LQ7PlU6_0),.clk(gclk));
	jdff dff_A_V20hFW2X6_0(.dout(w_dff_A_DPxxtKL94_0),.din(w_dff_A_V20hFW2X6_0),.clk(gclk));
	jdff dff_A_DPxxtKL94_0(.dout(w_dff_A_Wap2CB2h7_0),.din(w_dff_A_DPxxtKL94_0),.clk(gclk));
	jdff dff_A_Wap2CB2h7_0(.dout(w_dff_A_UQaAL50u2_0),.din(w_dff_A_Wap2CB2h7_0),.clk(gclk));
	jdff dff_A_UQaAL50u2_0(.dout(w_dff_A_S9snbeRI7_0),.din(w_dff_A_UQaAL50u2_0),.clk(gclk));
	jdff dff_A_S9snbeRI7_0(.dout(w_dff_A_7IQzRKXI5_0),.din(w_dff_A_S9snbeRI7_0),.clk(gclk));
	jdff dff_A_7IQzRKXI5_0(.dout(w_dff_A_Utk6dRhz3_0),.din(w_dff_A_7IQzRKXI5_0),.clk(gclk));
	jdff dff_A_Utk6dRhz3_0(.dout(w_dff_A_RxYoKcRC1_0),.din(w_dff_A_Utk6dRhz3_0),.clk(gclk));
	jdff dff_A_RxYoKcRC1_0(.dout(w_dff_A_pPyncxk59_0),.din(w_dff_A_RxYoKcRC1_0),.clk(gclk));
	jdff dff_A_pPyncxk59_0(.dout(w_dff_A_KXhRlyXG2_0),.din(w_dff_A_pPyncxk59_0),.clk(gclk));
	jdff dff_A_KXhRlyXG2_0(.dout(w_dff_A_M1TIjveT3_0),.din(w_dff_A_KXhRlyXG2_0),.clk(gclk));
	jdff dff_A_M1TIjveT3_0(.dout(w_dff_A_QcxhskVs4_0),.din(w_dff_A_M1TIjveT3_0),.clk(gclk));
	jdff dff_A_QcxhskVs4_0(.dout(w_dff_A_Cpsp4XmA0_0),.din(w_dff_A_QcxhskVs4_0),.clk(gclk));
	jdff dff_A_Cpsp4XmA0_0(.dout(w_dff_A_a3jxP59A5_0),.din(w_dff_A_Cpsp4XmA0_0),.clk(gclk));
	jdff dff_A_a3jxP59A5_0(.dout(w_dff_A_QOF6Jm5n6_0),.din(w_dff_A_a3jxP59A5_0),.clk(gclk));
	jdff dff_A_QOF6Jm5n6_0(.dout(w_dff_A_iiys9Ega1_0),.din(w_dff_A_QOF6Jm5n6_0),.clk(gclk));
	jdff dff_A_iiys9Ega1_0(.dout(w_dff_A_yl056mB47_0),.din(w_dff_A_iiys9Ega1_0),.clk(gclk));
	jdff dff_A_yl056mB47_0(.dout(w_dff_A_WY6T1iOP1_0),.din(w_dff_A_yl056mB47_0),.clk(gclk));
	jdff dff_A_WY6T1iOP1_0(.dout(w_dff_A_Y6DoH7Lu0_0),.din(w_dff_A_WY6T1iOP1_0),.clk(gclk));
	jdff dff_A_Y6DoH7Lu0_0(.dout(w_dff_A_VjKk6thg6_0),.din(w_dff_A_Y6DoH7Lu0_0),.clk(gclk));
	jdff dff_A_VjKk6thg6_0(.dout(w_dff_A_u6CIoNnq9_0),.din(w_dff_A_VjKk6thg6_0),.clk(gclk));
	jdff dff_A_u6CIoNnq9_0(.dout(w_dff_A_RjEsBuRu8_0),.din(w_dff_A_u6CIoNnq9_0),.clk(gclk));
	jdff dff_A_RjEsBuRu8_0(.dout(w_dff_A_tTsaSnpf8_0),.din(w_dff_A_RjEsBuRu8_0),.clk(gclk));
	jdff dff_A_tTsaSnpf8_0(.dout(w_dff_A_8ZOo8LCE9_0),.din(w_dff_A_tTsaSnpf8_0),.clk(gclk));
	jdff dff_A_8ZOo8LCE9_0(.dout(G5971gat),.din(w_dff_A_8ZOo8LCE9_0),.clk(gclk));
	jdff dff_A_r1aCngrq2_2(.dout(w_dff_A_XuFRjrVs3_0),.din(w_dff_A_r1aCngrq2_2),.clk(gclk));
	jdff dff_A_XuFRjrVs3_0(.dout(w_dff_A_v9YqiqXu5_0),.din(w_dff_A_XuFRjrVs3_0),.clk(gclk));
	jdff dff_A_v9YqiqXu5_0(.dout(w_dff_A_9AXGyz639_0),.din(w_dff_A_v9YqiqXu5_0),.clk(gclk));
	jdff dff_A_9AXGyz639_0(.dout(w_dff_A_C35h2YZ36_0),.din(w_dff_A_9AXGyz639_0),.clk(gclk));
	jdff dff_A_C35h2YZ36_0(.dout(w_dff_A_UHFQyyOC2_0),.din(w_dff_A_C35h2YZ36_0),.clk(gclk));
	jdff dff_A_UHFQyyOC2_0(.dout(w_dff_A_VjVYa70F9_0),.din(w_dff_A_UHFQyyOC2_0),.clk(gclk));
	jdff dff_A_VjVYa70F9_0(.dout(w_dff_A_AV07rs3B7_0),.din(w_dff_A_VjVYa70F9_0),.clk(gclk));
	jdff dff_A_AV07rs3B7_0(.dout(w_dff_A_OEBhgR793_0),.din(w_dff_A_AV07rs3B7_0),.clk(gclk));
	jdff dff_A_OEBhgR793_0(.dout(w_dff_A_GVKpoXPD8_0),.din(w_dff_A_OEBhgR793_0),.clk(gclk));
	jdff dff_A_GVKpoXPD8_0(.dout(w_dff_A_3mwVx50J9_0),.din(w_dff_A_GVKpoXPD8_0),.clk(gclk));
	jdff dff_A_3mwVx50J9_0(.dout(w_dff_A_OWo3gA2u8_0),.din(w_dff_A_3mwVx50J9_0),.clk(gclk));
	jdff dff_A_OWo3gA2u8_0(.dout(w_dff_A_HjjsXZHh5_0),.din(w_dff_A_OWo3gA2u8_0),.clk(gclk));
	jdff dff_A_HjjsXZHh5_0(.dout(w_dff_A_BqowqEYv2_0),.din(w_dff_A_HjjsXZHh5_0),.clk(gclk));
	jdff dff_A_BqowqEYv2_0(.dout(w_dff_A_Wd9GDAVx7_0),.din(w_dff_A_BqowqEYv2_0),.clk(gclk));
	jdff dff_A_Wd9GDAVx7_0(.dout(w_dff_A_yY3USx4c0_0),.din(w_dff_A_Wd9GDAVx7_0),.clk(gclk));
	jdff dff_A_yY3USx4c0_0(.dout(w_dff_A_vJDQ2GWV8_0),.din(w_dff_A_yY3USx4c0_0),.clk(gclk));
	jdff dff_A_vJDQ2GWV8_0(.dout(w_dff_A_9AdVyImf4_0),.din(w_dff_A_vJDQ2GWV8_0),.clk(gclk));
	jdff dff_A_9AdVyImf4_0(.dout(w_dff_A_u4N4Uje02_0),.din(w_dff_A_9AdVyImf4_0),.clk(gclk));
	jdff dff_A_u4N4Uje02_0(.dout(w_dff_A_9CxBwdcR8_0),.din(w_dff_A_u4N4Uje02_0),.clk(gclk));
	jdff dff_A_9CxBwdcR8_0(.dout(w_dff_A_twn4eA197_0),.din(w_dff_A_9CxBwdcR8_0),.clk(gclk));
	jdff dff_A_twn4eA197_0(.dout(w_dff_A_x361I8aL4_0),.din(w_dff_A_twn4eA197_0),.clk(gclk));
	jdff dff_A_x361I8aL4_0(.dout(w_dff_A_fJuP8nTE4_0),.din(w_dff_A_x361I8aL4_0),.clk(gclk));
	jdff dff_A_fJuP8nTE4_0(.dout(w_dff_A_ehniVHbJ3_0),.din(w_dff_A_fJuP8nTE4_0),.clk(gclk));
	jdff dff_A_ehniVHbJ3_0(.dout(w_dff_A_uVQFxzYX4_0),.din(w_dff_A_ehniVHbJ3_0),.clk(gclk));
	jdff dff_A_uVQFxzYX4_0(.dout(w_dff_A_iXpVjrUq3_0),.din(w_dff_A_uVQFxzYX4_0),.clk(gclk));
	jdff dff_A_iXpVjrUq3_0(.dout(w_dff_A_clUjrJxA2_0),.din(w_dff_A_iXpVjrUq3_0),.clk(gclk));
	jdff dff_A_clUjrJxA2_0(.dout(w_dff_A_pHNxuWoO9_0),.din(w_dff_A_clUjrJxA2_0),.clk(gclk));
	jdff dff_A_pHNxuWoO9_0(.dout(w_dff_A_4nlKqnzp8_0),.din(w_dff_A_pHNxuWoO9_0),.clk(gclk));
	jdff dff_A_4nlKqnzp8_0(.dout(w_dff_A_i6PJMHws9_0),.din(w_dff_A_4nlKqnzp8_0),.clk(gclk));
	jdff dff_A_i6PJMHws9_0(.dout(G6123gat),.din(w_dff_A_i6PJMHws9_0),.clk(gclk));
	jdff dff_A_Jo2F7egf8_2(.dout(w_dff_A_R1YbaEy04_0),.din(w_dff_A_Jo2F7egf8_2),.clk(gclk));
	jdff dff_A_R1YbaEy04_0(.dout(w_dff_A_XG9gEGcT6_0),.din(w_dff_A_R1YbaEy04_0),.clk(gclk));
	jdff dff_A_XG9gEGcT6_0(.dout(w_dff_A_ysQ9zyiw7_0),.din(w_dff_A_XG9gEGcT6_0),.clk(gclk));
	jdff dff_A_ysQ9zyiw7_0(.dout(w_dff_A_ISRYGuJm7_0),.din(w_dff_A_ysQ9zyiw7_0),.clk(gclk));
	jdff dff_A_ISRYGuJm7_0(.dout(w_dff_A_rjK2P2tH5_0),.din(w_dff_A_ISRYGuJm7_0),.clk(gclk));
	jdff dff_A_rjK2P2tH5_0(.dout(w_dff_A_IrYfBgBQ4_0),.din(w_dff_A_rjK2P2tH5_0),.clk(gclk));
	jdff dff_A_IrYfBgBQ4_0(.dout(w_dff_A_5HGTNa9z9_0),.din(w_dff_A_IrYfBgBQ4_0),.clk(gclk));
	jdff dff_A_5HGTNa9z9_0(.dout(w_dff_A_oCFTjAhD7_0),.din(w_dff_A_5HGTNa9z9_0),.clk(gclk));
	jdff dff_A_oCFTjAhD7_0(.dout(w_dff_A_eHkZvevr2_0),.din(w_dff_A_oCFTjAhD7_0),.clk(gclk));
	jdff dff_A_eHkZvevr2_0(.dout(w_dff_A_NVe5xkYR6_0),.din(w_dff_A_eHkZvevr2_0),.clk(gclk));
	jdff dff_A_NVe5xkYR6_0(.dout(w_dff_A_ei635nAD0_0),.din(w_dff_A_NVe5xkYR6_0),.clk(gclk));
	jdff dff_A_ei635nAD0_0(.dout(w_dff_A_Awg7C87t3_0),.din(w_dff_A_ei635nAD0_0),.clk(gclk));
	jdff dff_A_Awg7C87t3_0(.dout(w_dff_A_9TWscmz96_0),.din(w_dff_A_Awg7C87t3_0),.clk(gclk));
	jdff dff_A_9TWscmz96_0(.dout(w_dff_A_3WYPxpMa1_0),.din(w_dff_A_9TWscmz96_0),.clk(gclk));
	jdff dff_A_3WYPxpMa1_0(.dout(w_dff_A_qhsh2jpC2_0),.din(w_dff_A_3WYPxpMa1_0),.clk(gclk));
	jdff dff_A_qhsh2jpC2_0(.dout(w_dff_A_museoPD78_0),.din(w_dff_A_qhsh2jpC2_0),.clk(gclk));
	jdff dff_A_museoPD78_0(.dout(w_dff_A_bx0B8RLP8_0),.din(w_dff_A_museoPD78_0),.clk(gclk));
	jdff dff_A_bx0B8RLP8_0(.dout(w_dff_A_sDO8aYuP9_0),.din(w_dff_A_bx0B8RLP8_0),.clk(gclk));
	jdff dff_A_sDO8aYuP9_0(.dout(w_dff_A_mT9KQcqW7_0),.din(w_dff_A_sDO8aYuP9_0),.clk(gclk));
	jdff dff_A_mT9KQcqW7_0(.dout(w_dff_A_JKjdBYHm7_0),.din(w_dff_A_mT9KQcqW7_0),.clk(gclk));
	jdff dff_A_JKjdBYHm7_0(.dout(w_dff_A_ANsx75UK5_0),.din(w_dff_A_JKjdBYHm7_0),.clk(gclk));
	jdff dff_A_ANsx75UK5_0(.dout(w_dff_A_WdxnNWbO0_0),.din(w_dff_A_ANsx75UK5_0),.clk(gclk));
	jdff dff_A_WdxnNWbO0_0(.dout(w_dff_A_x5luIduw5_0),.din(w_dff_A_WdxnNWbO0_0),.clk(gclk));
	jdff dff_A_x5luIduw5_0(.dout(w_dff_A_DbbIKP4b6_0),.din(w_dff_A_x5luIduw5_0),.clk(gclk));
	jdff dff_A_DbbIKP4b6_0(.dout(w_dff_A_PtLRZelp4_0),.din(w_dff_A_DbbIKP4b6_0),.clk(gclk));
	jdff dff_A_PtLRZelp4_0(.dout(w_dff_A_XbyGK9nu9_0),.din(w_dff_A_PtLRZelp4_0),.clk(gclk));
	jdff dff_A_XbyGK9nu9_0(.dout(w_dff_A_sRgAlPUg1_0),.din(w_dff_A_XbyGK9nu9_0),.clk(gclk));
	jdff dff_A_sRgAlPUg1_0(.dout(G6150gat),.din(w_dff_A_sRgAlPUg1_0),.clk(gclk));
	jdff dff_A_4izfRJkS6_2(.dout(w_dff_A_ppsMkLmp8_0),.din(w_dff_A_4izfRJkS6_2),.clk(gclk));
	jdff dff_A_ppsMkLmp8_0(.dout(w_dff_A_zJoUeEbX8_0),.din(w_dff_A_ppsMkLmp8_0),.clk(gclk));
	jdff dff_A_zJoUeEbX8_0(.dout(w_dff_A_owbrdXYS4_0),.din(w_dff_A_zJoUeEbX8_0),.clk(gclk));
	jdff dff_A_owbrdXYS4_0(.dout(w_dff_A_wP8pYvmu2_0),.din(w_dff_A_owbrdXYS4_0),.clk(gclk));
	jdff dff_A_wP8pYvmu2_0(.dout(w_dff_A_Pj0roopd0_0),.din(w_dff_A_wP8pYvmu2_0),.clk(gclk));
	jdff dff_A_Pj0roopd0_0(.dout(w_dff_A_bHuVC1ga7_0),.din(w_dff_A_Pj0roopd0_0),.clk(gclk));
	jdff dff_A_bHuVC1ga7_0(.dout(w_dff_A_hqbjXSw79_0),.din(w_dff_A_bHuVC1ga7_0),.clk(gclk));
	jdff dff_A_hqbjXSw79_0(.dout(w_dff_A_25DlQBwS8_0),.din(w_dff_A_hqbjXSw79_0),.clk(gclk));
	jdff dff_A_25DlQBwS8_0(.dout(w_dff_A_rBRUGHOt2_0),.din(w_dff_A_25DlQBwS8_0),.clk(gclk));
	jdff dff_A_rBRUGHOt2_0(.dout(w_dff_A_1AatJLuc1_0),.din(w_dff_A_rBRUGHOt2_0),.clk(gclk));
	jdff dff_A_1AatJLuc1_0(.dout(w_dff_A_zfOMHR2N7_0),.din(w_dff_A_1AatJLuc1_0),.clk(gclk));
	jdff dff_A_zfOMHR2N7_0(.dout(w_dff_A_H6zG2bVS3_0),.din(w_dff_A_zfOMHR2N7_0),.clk(gclk));
	jdff dff_A_H6zG2bVS3_0(.dout(w_dff_A_ctlM9ASg1_0),.din(w_dff_A_H6zG2bVS3_0),.clk(gclk));
	jdff dff_A_ctlM9ASg1_0(.dout(w_dff_A_L6w3cSdp8_0),.din(w_dff_A_ctlM9ASg1_0),.clk(gclk));
	jdff dff_A_L6w3cSdp8_0(.dout(w_dff_A_KkFqToFD8_0),.din(w_dff_A_L6w3cSdp8_0),.clk(gclk));
	jdff dff_A_KkFqToFD8_0(.dout(w_dff_A_vTI7170r4_0),.din(w_dff_A_KkFqToFD8_0),.clk(gclk));
	jdff dff_A_vTI7170r4_0(.dout(w_dff_A_Ys7EmmBa4_0),.din(w_dff_A_vTI7170r4_0),.clk(gclk));
	jdff dff_A_Ys7EmmBa4_0(.dout(w_dff_A_8xEIQZeC8_0),.din(w_dff_A_Ys7EmmBa4_0),.clk(gclk));
	jdff dff_A_8xEIQZeC8_0(.dout(w_dff_A_wcm2MRYr4_0),.din(w_dff_A_8xEIQZeC8_0),.clk(gclk));
	jdff dff_A_wcm2MRYr4_0(.dout(w_dff_A_pvTt9bvg1_0),.din(w_dff_A_wcm2MRYr4_0),.clk(gclk));
	jdff dff_A_pvTt9bvg1_0(.dout(w_dff_A_0DoxGEUH1_0),.din(w_dff_A_pvTt9bvg1_0),.clk(gclk));
	jdff dff_A_0DoxGEUH1_0(.dout(w_dff_A_H0FKafym0_0),.din(w_dff_A_0DoxGEUH1_0),.clk(gclk));
	jdff dff_A_H0FKafym0_0(.dout(w_dff_A_6Z8AVGmP7_0),.din(w_dff_A_H0FKafym0_0),.clk(gclk));
	jdff dff_A_6Z8AVGmP7_0(.dout(w_dff_A_dbUExD566_0),.din(w_dff_A_6Z8AVGmP7_0),.clk(gclk));
	jdff dff_A_dbUExD566_0(.dout(w_dff_A_L4JrPjBs8_0),.din(w_dff_A_dbUExD566_0),.clk(gclk));
	jdff dff_A_L4JrPjBs8_0(.dout(G6160gat),.din(w_dff_A_L4JrPjBs8_0),.clk(gclk));
	jdff dff_A_x9VZLpLG1_2(.dout(w_dff_A_hzCEB60T6_0),.din(w_dff_A_x9VZLpLG1_2),.clk(gclk));
	jdff dff_A_hzCEB60T6_0(.dout(w_dff_A_VACDEFBw0_0),.din(w_dff_A_hzCEB60T6_0),.clk(gclk));
	jdff dff_A_VACDEFBw0_0(.dout(w_dff_A_j3WUboOe1_0),.din(w_dff_A_VACDEFBw0_0),.clk(gclk));
	jdff dff_A_j3WUboOe1_0(.dout(w_dff_A_7b85qm3S8_0),.din(w_dff_A_j3WUboOe1_0),.clk(gclk));
	jdff dff_A_7b85qm3S8_0(.dout(w_dff_A_W7pE5v2l1_0),.din(w_dff_A_7b85qm3S8_0),.clk(gclk));
	jdff dff_A_W7pE5v2l1_0(.dout(w_dff_A_HQKdiD9s4_0),.din(w_dff_A_W7pE5v2l1_0),.clk(gclk));
	jdff dff_A_HQKdiD9s4_0(.dout(w_dff_A_F2xwVygP3_0),.din(w_dff_A_HQKdiD9s4_0),.clk(gclk));
	jdff dff_A_F2xwVygP3_0(.dout(w_dff_A_PSnqNOKP1_0),.din(w_dff_A_F2xwVygP3_0),.clk(gclk));
	jdff dff_A_PSnqNOKP1_0(.dout(w_dff_A_gA6GfLkW5_0),.din(w_dff_A_PSnqNOKP1_0),.clk(gclk));
	jdff dff_A_gA6GfLkW5_0(.dout(w_dff_A_57KLEFYh0_0),.din(w_dff_A_gA6GfLkW5_0),.clk(gclk));
	jdff dff_A_57KLEFYh0_0(.dout(w_dff_A_TvW63X6d6_0),.din(w_dff_A_57KLEFYh0_0),.clk(gclk));
	jdff dff_A_TvW63X6d6_0(.dout(w_dff_A_o2MrrdRB9_0),.din(w_dff_A_TvW63X6d6_0),.clk(gclk));
	jdff dff_A_o2MrrdRB9_0(.dout(w_dff_A_sKac6gYO8_0),.din(w_dff_A_o2MrrdRB9_0),.clk(gclk));
	jdff dff_A_sKac6gYO8_0(.dout(w_dff_A_uDCZ8FDm6_0),.din(w_dff_A_sKac6gYO8_0),.clk(gclk));
	jdff dff_A_uDCZ8FDm6_0(.dout(w_dff_A_JNWJh7cx5_0),.din(w_dff_A_uDCZ8FDm6_0),.clk(gclk));
	jdff dff_A_JNWJh7cx5_0(.dout(w_dff_A_hdd8L2608_0),.din(w_dff_A_JNWJh7cx5_0),.clk(gclk));
	jdff dff_A_hdd8L2608_0(.dout(w_dff_A_xLEkBZKi1_0),.din(w_dff_A_hdd8L2608_0),.clk(gclk));
	jdff dff_A_xLEkBZKi1_0(.dout(w_dff_A_8B1JFkR21_0),.din(w_dff_A_xLEkBZKi1_0),.clk(gclk));
	jdff dff_A_8B1JFkR21_0(.dout(w_dff_A_XXhdQzVp9_0),.din(w_dff_A_8B1JFkR21_0),.clk(gclk));
	jdff dff_A_XXhdQzVp9_0(.dout(w_dff_A_vpLYzyqZ6_0),.din(w_dff_A_XXhdQzVp9_0),.clk(gclk));
	jdff dff_A_vpLYzyqZ6_0(.dout(w_dff_A_8B162l1j9_0),.din(w_dff_A_vpLYzyqZ6_0),.clk(gclk));
	jdff dff_A_8B162l1j9_0(.dout(w_dff_A_fbjChCzp6_0),.din(w_dff_A_8B162l1j9_0),.clk(gclk));
	jdff dff_A_fbjChCzp6_0(.dout(w_dff_A_d5G44bY50_0),.din(w_dff_A_fbjChCzp6_0),.clk(gclk));
	jdff dff_A_d5G44bY50_0(.dout(w_dff_A_892Ip4n51_0),.din(w_dff_A_d5G44bY50_0),.clk(gclk));
	jdff dff_A_892Ip4n51_0(.dout(G6170gat),.din(w_dff_A_892Ip4n51_0),.clk(gclk));
	jdff dff_A_4IuXdUMj6_2(.dout(w_dff_A_mD81bi5v7_0),.din(w_dff_A_4IuXdUMj6_2),.clk(gclk));
	jdff dff_A_mD81bi5v7_0(.dout(w_dff_A_nMIKE5cS2_0),.din(w_dff_A_mD81bi5v7_0),.clk(gclk));
	jdff dff_A_nMIKE5cS2_0(.dout(w_dff_A_UWiyTxOQ7_0),.din(w_dff_A_nMIKE5cS2_0),.clk(gclk));
	jdff dff_A_UWiyTxOQ7_0(.dout(w_dff_A_2yv6LY7Y9_0),.din(w_dff_A_UWiyTxOQ7_0),.clk(gclk));
	jdff dff_A_2yv6LY7Y9_0(.dout(w_dff_A_2V2pQONp6_0),.din(w_dff_A_2yv6LY7Y9_0),.clk(gclk));
	jdff dff_A_2V2pQONp6_0(.dout(w_dff_A_iupM7qmo1_0),.din(w_dff_A_2V2pQONp6_0),.clk(gclk));
	jdff dff_A_iupM7qmo1_0(.dout(w_dff_A_M3lqxB9h1_0),.din(w_dff_A_iupM7qmo1_0),.clk(gclk));
	jdff dff_A_M3lqxB9h1_0(.dout(w_dff_A_8ZtcXfmc8_0),.din(w_dff_A_M3lqxB9h1_0),.clk(gclk));
	jdff dff_A_8ZtcXfmc8_0(.dout(w_dff_A_87cMEnYt4_0),.din(w_dff_A_8ZtcXfmc8_0),.clk(gclk));
	jdff dff_A_87cMEnYt4_0(.dout(w_dff_A_nh2SJF7z6_0),.din(w_dff_A_87cMEnYt4_0),.clk(gclk));
	jdff dff_A_nh2SJF7z6_0(.dout(w_dff_A_UGjwBSOp4_0),.din(w_dff_A_nh2SJF7z6_0),.clk(gclk));
	jdff dff_A_UGjwBSOp4_0(.dout(w_dff_A_JkqT5Qtz2_0),.din(w_dff_A_UGjwBSOp4_0),.clk(gclk));
	jdff dff_A_JkqT5Qtz2_0(.dout(w_dff_A_rAWPsB6q3_0),.din(w_dff_A_JkqT5Qtz2_0),.clk(gclk));
	jdff dff_A_rAWPsB6q3_0(.dout(w_dff_A_TjZDc58h2_0),.din(w_dff_A_rAWPsB6q3_0),.clk(gclk));
	jdff dff_A_TjZDc58h2_0(.dout(w_dff_A_ICaJKK2y7_0),.din(w_dff_A_TjZDc58h2_0),.clk(gclk));
	jdff dff_A_ICaJKK2y7_0(.dout(w_dff_A_ybsYYklZ1_0),.din(w_dff_A_ICaJKK2y7_0),.clk(gclk));
	jdff dff_A_ybsYYklZ1_0(.dout(w_dff_A_DoG3Qxi32_0),.din(w_dff_A_ybsYYklZ1_0),.clk(gclk));
	jdff dff_A_DoG3Qxi32_0(.dout(w_dff_A_f5p4Rh8X5_0),.din(w_dff_A_DoG3Qxi32_0),.clk(gclk));
	jdff dff_A_f5p4Rh8X5_0(.dout(w_dff_A_U33AsfOZ5_0),.din(w_dff_A_f5p4Rh8X5_0),.clk(gclk));
	jdff dff_A_U33AsfOZ5_0(.dout(w_dff_A_wA95lBlI2_0),.din(w_dff_A_U33AsfOZ5_0),.clk(gclk));
	jdff dff_A_wA95lBlI2_0(.dout(w_dff_A_pgP3a0OZ0_0),.din(w_dff_A_wA95lBlI2_0),.clk(gclk));
	jdff dff_A_pgP3a0OZ0_0(.dout(w_dff_A_FqZVic4Z9_0),.din(w_dff_A_pgP3a0OZ0_0),.clk(gclk));
	jdff dff_A_FqZVic4Z9_0(.dout(G6180gat),.din(w_dff_A_FqZVic4Z9_0),.clk(gclk));
	jdff dff_A_UJSpteTt5_2(.dout(w_dff_A_jkiZPCWk7_0),.din(w_dff_A_UJSpteTt5_2),.clk(gclk));
	jdff dff_A_jkiZPCWk7_0(.dout(w_dff_A_AjsoM0Mb5_0),.din(w_dff_A_jkiZPCWk7_0),.clk(gclk));
	jdff dff_A_AjsoM0Mb5_0(.dout(w_dff_A_oraR3IrY5_0),.din(w_dff_A_AjsoM0Mb5_0),.clk(gclk));
	jdff dff_A_oraR3IrY5_0(.dout(w_dff_A_WYhETyT44_0),.din(w_dff_A_oraR3IrY5_0),.clk(gclk));
	jdff dff_A_WYhETyT44_0(.dout(w_dff_A_QsK3XZyc0_0),.din(w_dff_A_WYhETyT44_0),.clk(gclk));
	jdff dff_A_QsK3XZyc0_0(.dout(w_dff_A_1PeAAIgu1_0),.din(w_dff_A_QsK3XZyc0_0),.clk(gclk));
	jdff dff_A_1PeAAIgu1_0(.dout(w_dff_A_hF4jqLLM7_0),.din(w_dff_A_1PeAAIgu1_0),.clk(gclk));
	jdff dff_A_hF4jqLLM7_0(.dout(w_dff_A_5aH49PcP0_0),.din(w_dff_A_hF4jqLLM7_0),.clk(gclk));
	jdff dff_A_5aH49PcP0_0(.dout(w_dff_A_tTJdCMNL7_0),.din(w_dff_A_5aH49PcP0_0),.clk(gclk));
	jdff dff_A_tTJdCMNL7_0(.dout(w_dff_A_Fwjtbq3s0_0),.din(w_dff_A_tTJdCMNL7_0),.clk(gclk));
	jdff dff_A_Fwjtbq3s0_0(.dout(w_dff_A_vYpDTAP79_0),.din(w_dff_A_Fwjtbq3s0_0),.clk(gclk));
	jdff dff_A_vYpDTAP79_0(.dout(w_dff_A_cUFFlbEi2_0),.din(w_dff_A_vYpDTAP79_0),.clk(gclk));
	jdff dff_A_cUFFlbEi2_0(.dout(w_dff_A_ZFjfCiaE8_0),.din(w_dff_A_cUFFlbEi2_0),.clk(gclk));
	jdff dff_A_ZFjfCiaE8_0(.dout(w_dff_A_NzUgoClu6_0),.din(w_dff_A_ZFjfCiaE8_0),.clk(gclk));
	jdff dff_A_NzUgoClu6_0(.dout(w_dff_A_2QzjacWM0_0),.din(w_dff_A_NzUgoClu6_0),.clk(gclk));
	jdff dff_A_2QzjacWM0_0(.dout(w_dff_A_41dcNXgg1_0),.din(w_dff_A_2QzjacWM0_0),.clk(gclk));
	jdff dff_A_41dcNXgg1_0(.dout(w_dff_A_mIbHVo4I9_0),.din(w_dff_A_41dcNXgg1_0),.clk(gclk));
	jdff dff_A_mIbHVo4I9_0(.dout(w_dff_A_L1o6rsPk1_0),.din(w_dff_A_mIbHVo4I9_0),.clk(gclk));
	jdff dff_A_L1o6rsPk1_0(.dout(w_dff_A_Z4Azrdl98_0),.din(w_dff_A_L1o6rsPk1_0),.clk(gclk));
	jdff dff_A_Z4Azrdl98_0(.dout(w_dff_A_Vaodozu85_0),.din(w_dff_A_Z4Azrdl98_0),.clk(gclk));
	jdff dff_A_Vaodozu85_0(.dout(G6190gat),.din(w_dff_A_Vaodozu85_0),.clk(gclk));
	jdff dff_A_X5zW4CkD5_2(.dout(w_dff_A_OMfjOz0S3_0),.din(w_dff_A_X5zW4CkD5_2),.clk(gclk));
	jdff dff_A_OMfjOz0S3_0(.dout(w_dff_A_TDJQUoIB6_0),.din(w_dff_A_OMfjOz0S3_0),.clk(gclk));
	jdff dff_A_TDJQUoIB6_0(.dout(w_dff_A_XebOGDqY7_0),.din(w_dff_A_TDJQUoIB6_0),.clk(gclk));
	jdff dff_A_XebOGDqY7_0(.dout(w_dff_A_oCjiPegq0_0),.din(w_dff_A_XebOGDqY7_0),.clk(gclk));
	jdff dff_A_oCjiPegq0_0(.dout(w_dff_A_wn0Yqp8p2_0),.din(w_dff_A_oCjiPegq0_0),.clk(gclk));
	jdff dff_A_wn0Yqp8p2_0(.dout(w_dff_A_kD4AmjX62_0),.din(w_dff_A_wn0Yqp8p2_0),.clk(gclk));
	jdff dff_A_kD4AmjX62_0(.dout(w_dff_A_rIoUoEs72_0),.din(w_dff_A_kD4AmjX62_0),.clk(gclk));
	jdff dff_A_rIoUoEs72_0(.dout(w_dff_A_Hk1b5o689_0),.din(w_dff_A_rIoUoEs72_0),.clk(gclk));
	jdff dff_A_Hk1b5o689_0(.dout(w_dff_A_Y5soYLYw2_0),.din(w_dff_A_Hk1b5o689_0),.clk(gclk));
	jdff dff_A_Y5soYLYw2_0(.dout(w_dff_A_OKWVZp9u2_0),.din(w_dff_A_Y5soYLYw2_0),.clk(gclk));
	jdff dff_A_OKWVZp9u2_0(.dout(w_dff_A_iLpN0RAr4_0),.din(w_dff_A_OKWVZp9u2_0),.clk(gclk));
	jdff dff_A_iLpN0RAr4_0(.dout(w_dff_A_olVfXW3u3_0),.din(w_dff_A_iLpN0RAr4_0),.clk(gclk));
	jdff dff_A_olVfXW3u3_0(.dout(w_dff_A_RBXGyFvD1_0),.din(w_dff_A_olVfXW3u3_0),.clk(gclk));
	jdff dff_A_RBXGyFvD1_0(.dout(w_dff_A_0AYV3bIS0_0),.din(w_dff_A_RBXGyFvD1_0),.clk(gclk));
	jdff dff_A_0AYV3bIS0_0(.dout(w_dff_A_uaBW9Ssy0_0),.din(w_dff_A_0AYV3bIS0_0),.clk(gclk));
	jdff dff_A_uaBW9Ssy0_0(.dout(w_dff_A_fF9BKSPy9_0),.din(w_dff_A_uaBW9Ssy0_0),.clk(gclk));
	jdff dff_A_fF9BKSPy9_0(.dout(w_dff_A_WbnvdjBE7_0),.din(w_dff_A_fF9BKSPy9_0),.clk(gclk));
	jdff dff_A_WbnvdjBE7_0(.dout(w_dff_A_2U9O2W6l1_0),.din(w_dff_A_WbnvdjBE7_0),.clk(gclk));
	jdff dff_A_2U9O2W6l1_0(.dout(G6200gat),.din(w_dff_A_2U9O2W6l1_0),.clk(gclk));
	jdff dff_A_FtorKECO3_2(.dout(w_dff_A_U6FkGW781_0),.din(w_dff_A_FtorKECO3_2),.clk(gclk));
	jdff dff_A_U6FkGW781_0(.dout(w_dff_A_tB8FVRi90_0),.din(w_dff_A_U6FkGW781_0),.clk(gclk));
	jdff dff_A_tB8FVRi90_0(.dout(w_dff_A_zvHMMnu73_0),.din(w_dff_A_tB8FVRi90_0),.clk(gclk));
	jdff dff_A_zvHMMnu73_0(.dout(w_dff_A_y1yEPVtH6_0),.din(w_dff_A_zvHMMnu73_0),.clk(gclk));
	jdff dff_A_y1yEPVtH6_0(.dout(w_dff_A_pjl44f2L0_0),.din(w_dff_A_y1yEPVtH6_0),.clk(gclk));
	jdff dff_A_pjl44f2L0_0(.dout(w_dff_A_XXla3sAj5_0),.din(w_dff_A_pjl44f2L0_0),.clk(gclk));
	jdff dff_A_XXla3sAj5_0(.dout(w_dff_A_ihL53V6l3_0),.din(w_dff_A_XXla3sAj5_0),.clk(gclk));
	jdff dff_A_ihL53V6l3_0(.dout(w_dff_A_YUYTSKZj1_0),.din(w_dff_A_ihL53V6l3_0),.clk(gclk));
	jdff dff_A_YUYTSKZj1_0(.dout(w_dff_A_1qhbX22m1_0),.din(w_dff_A_YUYTSKZj1_0),.clk(gclk));
	jdff dff_A_1qhbX22m1_0(.dout(w_dff_A_NXSUIUMR0_0),.din(w_dff_A_1qhbX22m1_0),.clk(gclk));
	jdff dff_A_NXSUIUMR0_0(.dout(w_dff_A_T7wgGDDF9_0),.din(w_dff_A_NXSUIUMR0_0),.clk(gclk));
	jdff dff_A_T7wgGDDF9_0(.dout(w_dff_A_YKX4wmdg3_0),.din(w_dff_A_T7wgGDDF9_0),.clk(gclk));
	jdff dff_A_YKX4wmdg3_0(.dout(w_dff_A_yyGzkcoc7_0),.din(w_dff_A_YKX4wmdg3_0),.clk(gclk));
	jdff dff_A_yyGzkcoc7_0(.dout(w_dff_A_xX4xaIry1_0),.din(w_dff_A_yyGzkcoc7_0),.clk(gclk));
	jdff dff_A_xX4xaIry1_0(.dout(w_dff_A_vq6Z7ur67_0),.din(w_dff_A_xX4xaIry1_0),.clk(gclk));
	jdff dff_A_vq6Z7ur67_0(.dout(w_dff_A_sN8G1tc00_0),.din(w_dff_A_vq6Z7ur67_0),.clk(gclk));
	jdff dff_A_sN8G1tc00_0(.dout(G6210gat),.din(w_dff_A_sN8G1tc00_0),.clk(gclk));
	jdff dff_A_EvWttnxa3_2(.dout(w_dff_A_zMc6k8E98_0),.din(w_dff_A_EvWttnxa3_2),.clk(gclk));
	jdff dff_A_zMc6k8E98_0(.dout(w_dff_A_lKKvZpJl4_0),.din(w_dff_A_zMc6k8E98_0),.clk(gclk));
	jdff dff_A_lKKvZpJl4_0(.dout(w_dff_A_D9XZdQ9X8_0),.din(w_dff_A_lKKvZpJl4_0),.clk(gclk));
	jdff dff_A_D9XZdQ9X8_0(.dout(w_dff_A_dtLH0Y6l3_0),.din(w_dff_A_D9XZdQ9X8_0),.clk(gclk));
	jdff dff_A_dtLH0Y6l3_0(.dout(w_dff_A_ltLPvjfK4_0),.din(w_dff_A_dtLH0Y6l3_0),.clk(gclk));
	jdff dff_A_ltLPvjfK4_0(.dout(w_dff_A_kPu6HoWO2_0),.din(w_dff_A_ltLPvjfK4_0),.clk(gclk));
	jdff dff_A_kPu6HoWO2_0(.dout(w_dff_A_EPFWUV8h6_0),.din(w_dff_A_kPu6HoWO2_0),.clk(gclk));
	jdff dff_A_EPFWUV8h6_0(.dout(w_dff_A_ZMeag6LT5_0),.din(w_dff_A_EPFWUV8h6_0),.clk(gclk));
	jdff dff_A_ZMeag6LT5_0(.dout(w_dff_A_5w726Ijp3_0),.din(w_dff_A_ZMeag6LT5_0),.clk(gclk));
	jdff dff_A_5w726Ijp3_0(.dout(w_dff_A_c8WMq0EH1_0),.din(w_dff_A_5w726Ijp3_0),.clk(gclk));
	jdff dff_A_c8WMq0EH1_0(.dout(w_dff_A_X96knW085_0),.din(w_dff_A_c8WMq0EH1_0),.clk(gclk));
	jdff dff_A_X96knW085_0(.dout(w_dff_A_51tvmUTu7_0),.din(w_dff_A_X96knW085_0),.clk(gclk));
	jdff dff_A_51tvmUTu7_0(.dout(w_dff_A_6ek4ZFL08_0),.din(w_dff_A_51tvmUTu7_0),.clk(gclk));
	jdff dff_A_6ek4ZFL08_0(.dout(w_dff_A_phJnpuEk4_0),.din(w_dff_A_6ek4ZFL08_0),.clk(gclk));
	jdff dff_A_phJnpuEk4_0(.dout(G6220gat),.din(w_dff_A_phJnpuEk4_0),.clk(gclk));
	jdff dff_A_TLmwHIhE1_2(.dout(w_dff_A_nXGdspfK3_0),.din(w_dff_A_TLmwHIhE1_2),.clk(gclk));
	jdff dff_A_nXGdspfK3_0(.dout(w_dff_A_FIX0YiuS9_0),.din(w_dff_A_nXGdspfK3_0),.clk(gclk));
	jdff dff_A_FIX0YiuS9_0(.dout(w_dff_A_5O5Qqwkd4_0),.din(w_dff_A_FIX0YiuS9_0),.clk(gclk));
	jdff dff_A_5O5Qqwkd4_0(.dout(w_dff_A_29hlMrLC8_0),.din(w_dff_A_5O5Qqwkd4_0),.clk(gclk));
	jdff dff_A_29hlMrLC8_0(.dout(w_dff_A_so3Uc0T45_0),.din(w_dff_A_29hlMrLC8_0),.clk(gclk));
	jdff dff_A_so3Uc0T45_0(.dout(w_dff_A_HvjJnEIJ6_0),.din(w_dff_A_so3Uc0T45_0),.clk(gclk));
	jdff dff_A_HvjJnEIJ6_0(.dout(w_dff_A_K5Sk7pRt4_0),.din(w_dff_A_HvjJnEIJ6_0),.clk(gclk));
	jdff dff_A_K5Sk7pRt4_0(.dout(w_dff_A_Z9yG4cs03_0),.din(w_dff_A_K5Sk7pRt4_0),.clk(gclk));
	jdff dff_A_Z9yG4cs03_0(.dout(w_dff_A_O7tpWd0y7_0),.din(w_dff_A_Z9yG4cs03_0),.clk(gclk));
	jdff dff_A_O7tpWd0y7_0(.dout(w_dff_A_L88DLSrW3_0),.din(w_dff_A_O7tpWd0y7_0),.clk(gclk));
	jdff dff_A_L88DLSrW3_0(.dout(w_dff_A_9m8JFDcT3_0),.din(w_dff_A_L88DLSrW3_0),.clk(gclk));
	jdff dff_A_9m8JFDcT3_0(.dout(w_dff_A_dixSqDUG8_0),.din(w_dff_A_9m8JFDcT3_0),.clk(gclk));
	jdff dff_A_dixSqDUG8_0(.dout(G6230gat),.din(w_dff_A_dixSqDUG8_0),.clk(gclk));
	jdff dff_A_np4nDYGT0_2(.dout(w_dff_A_OQNzrkQT3_0),.din(w_dff_A_np4nDYGT0_2),.clk(gclk));
	jdff dff_A_OQNzrkQT3_0(.dout(w_dff_A_yplJ0Ykl3_0),.din(w_dff_A_OQNzrkQT3_0),.clk(gclk));
	jdff dff_A_yplJ0Ykl3_0(.dout(w_dff_A_fx1eFLLd6_0),.din(w_dff_A_yplJ0Ykl3_0),.clk(gclk));
	jdff dff_A_fx1eFLLd6_0(.dout(w_dff_A_sxW095fL2_0),.din(w_dff_A_fx1eFLLd6_0),.clk(gclk));
	jdff dff_A_sxW095fL2_0(.dout(w_dff_A_7NrR5XjK2_0),.din(w_dff_A_sxW095fL2_0),.clk(gclk));
	jdff dff_A_7NrR5XjK2_0(.dout(w_dff_A_g8o6yiBn1_0),.din(w_dff_A_7NrR5XjK2_0),.clk(gclk));
	jdff dff_A_g8o6yiBn1_0(.dout(w_dff_A_VeNVzcJc0_0),.din(w_dff_A_g8o6yiBn1_0),.clk(gclk));
	jdff dff_A_VeNVzcJc0_0(.dout(w_dff_A_rvvPdYNb0_0),.din(w_dff_A_VeNVzcJc0_0),.clk(gclk));
	jdff dff_A_rvvPdYNb0_0(.dout(w_dff_A_fOgzutYn2_0),.din(w_dff_A_rvvPdYNb0_0),.clk(gclk));
	jdff dff_A_fOgzutYn2_0(.dout(w_dff_A_40PEDUQR7_0),.din(w_dff_A_fOgzutYn2_0),.clk(gclk));
	jdff dff_A_40PEDUQR7_0(.dout(G6240gat),.din(w_dff_A_40PEDUQR7_0),.clk(gclk));
	jdff dff_A_MxA6KRqk3_2(.dout(w_dff_A_qty7FCa43_0),.din(w_dff_A_MxA6KRqk3_2),.clk(gclk));
	jdff dff_A_qty7FCa43_0(.dout(w_dff_A_rz1JjpZ09_0),.din(w_dff_A_qty7FCa43_0),.clk(gclk));
	jdff dff_A_rz1JjpZ09_0(.dout(w_dff_A_8YYLDw7X4_0),.din(w_dff_A_rz1JjpZ09_0),.clk(gclk));
	jdff dff_A_8YYLDw7X4_0(.dout(w_dff_A_gEc8NJbU0_0),.din(w_dff_A_8YYLDw7X4_0),.clk(gclk));
	jdff dff_A_gEc8NJbU0_0(.dout(w_dff_A_TkHTf4Y76_0),.din(w_dff_A_gEc8NJbU0_0),.clk(gclk));
	jdff dff_A_TkHTf4Y76_0(.dout(w_dff_A_hQAustIc1_0),.din(w_dff_A_TkHTf4Y76_0),.clk(gclk));
	jdff dff_A_hQAustIc1_0(.dout(w_dff_A_IGsU7fHb8_0),.din(w_dff_A_hQAustIc1_0),.clk(gclk));
	jdff dff_A_IGsU7fHb8_0(.dout(w_dff_A_LOpn4Y7Y4_0),.din(w_dff_A_IGsU7fHb8_0),.clk(gclk));
	jdff dff_A_LOpn4Y7Y4_0(.dout(G6250gat),.din(w_dff_A_LOpn4Y7Y4_0),.clk(gclk));
	jdff dff_A_vaZ8kvun7_2(.dout(w_dff_A_fl4lL1AN3_0),.din(w_dff_A_vaZ8kvun7_2),.clk(gclk));
	jdff dff_A_fl4lL1AN3_0(.dout(w_dff_A_UiiR4dBg9_0),.din(w_dff_A_fl4lL1AN3_0),.clk(gclk));
	jdff dff_A_UiiR4dBg9_0(.dout(w_dff_A_4PeI1Z3o0_0),.din(w_dff_A_UiiR4dBg9_0),.clk(gclk));
	jdff dff_A_4PeI1Z3o0_0(.dout(w_dff_A_bDg38os87_0),.din(w_dff_A_4PeI1Z3o0_0),.clk(gclk));
	jdff dff_A_bDg38os87_0(.dout(w_dff_A_AbQW1K2o9_0),.din(w_dff_A_bDg38os87_0),.clk(gclk));
	jdff dff_A_AbQW1K2o9_0(.dout(w_dff_A_W4tUHAVz7_0),.din(w_dff_A_AbQW1K2o9_0),.clk(gclk));
	jdff dff_A_W4tUHAVz7_0(.dout(G6260gat),.din(w_dff_A_W4tUHAVz7_0),.clk(gclk));
	jdff dff_A_QTxU36lP3_2(.dout(w_dff_A_SdRFDCEB9_0),.din(w_dff_A_QTxU36lP3_2),.clk(gclk));
	jdff dff_A_SdRFDCEB9_0(.dout(w_dff_A_DUo9KVGb3_0),.din(w_dff_A_SdRFDCEB9_0),.clk(gclk));
	jdff dff_A_DUo9KVGb3_0(.dout(w_dff_A_gCpavY280_0),.din(w_dff_A_DUo9KVGb3_0),.clk(gclk));
	jdff dff_A_gCpavY280_0(.dout(w_dff_A_nISZq5Dm2_0),.din(w_dff_A_gCpavY280_0),.clk(gclk));
	jdff dff_A_nISZq5Dm2_0(.dout(G6270gat),.din(w_dff_A_nISZq5Dm2_0),.clk(gclk));
	jdff dff_A_emw7PjXC7_2(.dout(w_dff_A_Ng3v1Jn62_0),.din(w_dff_A_emw7PjXC7_2),.clk(gclk));
	jdff dff_A_Ng3v1Jn62_0(.dout(w_dff_A_SZ5hnu3S8_0),.din(w_dff_A_Ng3v1Jn62_0),.clk(gclk));
	jdff dff_A_SZ5hnu3S8_0(.dout(G6280gat),.din(w_dff_A_SZ5hnu3S8_0),.clk(gclk));
	jdff dff_A_roQXFJyg9_2(.dout(G6288gat),.din(w_dff_A_roQXFJyg9_2),.clk(gclk));
endmodule

