module rf_c1908(G902, G900, G116, G143, G125, G227, G134, G952, G122, G221, G119, G898, G224, G107, G101, G140, G472, G110, G478, G104, G128, G131, G234, G137, G146, G210, G217, G953, G113, G237, G214, G469, G475, G57, G66, G69, G63, G54, G51, G72, G42, G39, G36, G3, G45, G6, G9, G27, G12, G30, G48, G15, G18, G21, G24, G60, G75, G33);
    input G902, G900, G116, G143, G125, G227, G134, G952, G122, G221, G119, G898, G224, G107, G101, G140, G472, G110, G478, G104, G128, G131, G234, G137, G146, G210, G217, G953, G113, G237, G214, G469, G475;
    output G57, G66, G69, G63, G54, G51, G72, G42, G39, G36, G3, G45, G6, G9, G27, G12, G30, G48, G15, G18, G21, G24, G60, G75, G33;
    wire n60;
    wire n64;
    wire n68;
    wire n71;
    wire n75;
    wire n79;
    wire n83;
    wire n87;
    wire n91;
    wire n95;
    wire n99;
    wire n103;
    wire n106;
    wire n110;
    wire n113;
    wire n117;
    wire n121;
    wire n124;
    wire n128;
    wire n131;
    wire n135;
    wire n139;
    wire n143;
    wire n147;
    wire n150;
    wire n154;
    wire n158;
    wire n161;
    wire n165;
    wire n169;
    wire n173;
    wire n177;
    wire n181;
    wire n185;
    wire n189;
    wire n193;
    wire n197;
    wire n201;
    wire n204;
    wire n208;
    wire n211;
    wire n215;
    wire n219;
    wire n223;
    wire n227;
    wire n231;
    wire n235;
    wire n239;
    wire n243;
    wire n247;
    wire n251;
    wire n255;
    wire n259;
    wire n262;
    wire n266;
    wire n270;
    wire n274;
    wire n278;
    wire n282;
    wire n286;
    wire n290;
    wire n294;
    wire n298;
    wire n302;
    wire n306;
    wire n309;
    wire n313;
    wire n317;
    wire n321;
    wire n325;
    wire n329;
    wire n333;
    wire n337;
    wire n341;
    wire n345;
    wire n348;
    wire n352;
    wire n356;
    wire n360;
    wire n363;
    wire n367;
    wire n371;
    wire n375;
    wire n379;
    wire n383;
    wire n387;
    wire n391;
    wire n395;
    wire n399;
    wire n403;
    wire n407;
    wire n410;
    wire n414;
    wire n418;
    wire n421;
    wire n425;
    wire n428;
    wire n432;
    wire n436;
    wire n440;
    wire n443;
    wire n447;
    wire n451;
    wire n455;
    wire n459;
    wire n463;
    wire n467;
    wire n471;
    wire n475;
    wire n479;
    wire n483;
    wire n487;
    wire n491;
    wire n494;
    wire n498;
    wire n502;
    wire n506;
    wire n510;
    wire n514;
    wire n518;
    wire n522;
    wire n526;
    wire n530;
    wire n534;
    wire n538;
    wire n542;
    wire n545;
    wire n549;
    wire n553;
    wire n557;
    wire n561;
    wire n565;
    wire n569;
    wire n573;
    wire n577;
    wire n581;
    wire n585;
    wire n588;
    wire n592;
    wire n596;
    wire n600;
    wire n604;
    wire n608;
    wire n612;
    wire n616;
    wire n620;
    wire n624;
    wire n628;
    wire n632;
    wire n636;
    wire n640;
    wire n644;
    wire n648;
    wire n652;
    wire n656;
    wire n660;
    wire n664;
    wire n667;
    wire n671;
    wire n675;
    wire n679;
    wire n683;
    wire n687;
    wire n691;
    wire n695;
    wire n699;
    wire n703;
    wire n707;
    wire n711;
    wire n715;
    wire n719;
    wire n723;
    wire n727;
    wire n731;
    wire n735;
    wire n739;
    wire n743;
    wire n747;
    wire n751;
    wire n755;
    wire n759;
    wire n763;
    wire n767;
    wire n771;
    wire n775;
    wire n779;
    wire n783;
    wire n787;
    wire n791;
    wire n795;
    wire n799;
    wire n803;
    wire n807;
    wire n811;
    wire n815;
    wire n819;
    wire n823;
    wire n827;
    wire n831;
    wire n835;
    wire n839;
    wire n843;
    wire n847;
    wire n851;
    wire n855;
    wire n859;
    wire n863;
    wire n867;
    wire n871;
    wire n875;
    wire n879;
    wire n883;
    wire n887;
    wire n891;
    wire n894;
    wire n898;
    wire n901;
    wire n905;
    wire n909;
    wire n913;
    wire n916;
    wire n920;
    wire n924;
    wire n928;
    wire n932;
    wire n936;
    wire n940;
    wire n944;
    wire n947;
    wire n951;
    wire n955;
    wire n959;
    wire n963;
    wire n967;
    wire n971;
    wire n975;
    wire n979;
    wire n983;
    wire n987;
    wire n991;
    wire n995;
    wire n999;
    wire n1003;
    wire n1007;
    wire n1010;
    wire n1014;
    wire n1018;
    wire n1022;
    wire n1026;
    wire n1030;
    wire n1034;
    wire n1038;
    wire n1042;
    wire n1046;
    wire n1050;
    wire n1054;
    wire n1058;
    wire n1062;
    wire n1066;
    wire n1070;
    wire n1073;
    wire n1077;
    wire n1081;
    wire n1085;
    wire n1089;
    wire n1092;
    wire n1096;
    wire n1100;
    wire n1104;
    wire n1108;
    wire n1112;
    wire n1116;
    wire n1120;
    wire n1124;
    wire n1128;
    wire n1132;
    wire n1136;
    wire n1140;
    wire n1144;
    wire n1147;
    wire n1151;
    wire n1155;
    wire n1159;
    wire n1163;
    wire n1167;
    wire n1171;
    wire n1178;
    wire n1182;
    wire n1185;
    wire n1189;
    wire n1193;
    wire n1197;
    wire n1201;
    wire n1205;
    wire n1212;
    wire n1216;
    wire n1219;
    wire n1223;
    wire n1227;
    wire n1231;
    wire n1235;
    wire n1239;
    wire n1246;
    wire n1250;
    wire n1253;
    wire n1257;
    wire n1261;
    wire n1265;
    wire n1269;
    wire n1273;
    wire n1281;
    wire n1285;
    wire n1289;
    wire n1292;
    wire n1296;
    wire n1300;
    wire n1304;
    wire n1311;
    wire n1315;
    wire n1319;
    wire n1323;
    wire n1327;
    wire n1331;
    wire n1335;
    wire n1339;
    wire n1343;
    wire n1347;
    wire n1350;
    wire n1354;
    wire n1358;
    wire n1362;
    wire n1365;
    wire n1369;
    wire n1372;
    wire n1376;
    wire n1380;
    wire n1384;
    wire n1388;
    wire n1392;
    wire n2097;
    wire n2100;
    wire n2103;
    wire n2106;
    wire n2109;
    wire n2112;
    wire n2115;
    wire n2118;
    wire n2121;
    wire n2124;
    wire n2127;
    wire n2130;
    wire n2132;
    wire n2136;
    wire n2139;
    wire n2142;
    wire n2145;
    wire n2148;
    wire n2151;
    wire n2154;
    wire n2157;
    wire n2160;
    wire n2163;
    wire n2166;
    wire n2169;
    wire n2172;
    wire n2175;
    wire n2178;
    wire n2181;
    wire n2184;
    wire n2187;
    wire n2190;
    wire n2193;
    wire n2196;
    wire n2199;
    wire n2202;
    wire n2205;
    wire n2208;
    wire n2211;
    wire n2214;
    wire n2217;
    wire n2220;
    wire n2223;
    wire n2225;
    wire n2228;
    wire n2231;
    wire n2234;
    wire n2237;
    wire n2240;
    wire n2243;
    wire n2246;
    wire n2249;
    wire n2252;
    wire n2255;
    wire n2258;
    wire n2261;
    wire n2264;
    wire n2267;
    wire n2271;
    wire n2274;
    wire n2277;
    wire n2280;
    wire n2283;
    wire n2286;
    wire n2289;
    wire n2292;
    wire n2295;
    wire n2298;
    wire n2301;
    wire n2304;
    wire n2307;
    wire n2310;
    wire n2313;
    wire n2316;
    wire n2319;
    wire n2322;
    wire n2325;
    wire n2328;
    wire n2331;
    wire n2334;
    wire n2337;
    wire n2340;
    wire n2343;
    wire n2346;
    wire n2348;
    wire n2351;
    wire n2354;
    wire n2357;
    wire n2360;
    wire n2363;
    wire n2366;
    wire n2369;
    wire n2372;
    wire n2375;
    wire n2378;
    wire n2381;
    wire n2384;
    wire n2387;
    wire n2390;
    wire n2394;
    wire n2397;
    wire n2400;
    wire n2403;
    wire n2406;
    wire n2409;
    wire n2412;
    wire n2415;
    wire n2418;
    wire n2421;
    wire n2424;
    wire n2427;
    wire n2430;
    wire n2433;
    wire n2436;
    wire n2439;
    wire n2442;
    wire n2445;
    wire n2448;
    wire n2451;
    wire n2454;
    wire n2457;
    wire n2460;
    wire n2463;
    wire n2466;
    wire n2469;
    wire n2471;
    wire n2474;
    wire n2477;
    wire n2480;
    wire n2483;
    wire n2486;
    wire n2489;
    wire n2492;
    wire n2495;
    wire n2498;
    wire n2501;
    wire n2504;
    wire n2507;
    wire n2510;
    wire n2513;
    wire n2517;
    wire n2520;
    wire n2523;
    wire n2526;
    wire n2529;
    wire n2532;
    wire n2535;
    wire n2538;
    wire n2541;
    wire n2544;
    wire n2547;
    wire n2550;
    wire n2553;
    wire n2556;
    wire n2559;
    wire n2562;
    wire n2565;
    wire n2568;
    wire n2571;
    wire n2574;
    wire n2577;
    wire n2580;
    wire n2583;
    wire n2586;
    wire n2589;
    wire n2592;
    wire n2594;
    wire n2597;
    wire n2600;
    wire n2603;
    wire n2606;
    wire n2609;
    wire n2612;
    wire n2615;
    wire n2618;
    wire n2621;
    wire n2624;
    wire n2627;
    wire n2630;
    wire n2633;
    wire n2636;
    wire n2640;
    wire n2643;
    wire n2646;
    wire n2649;
    wire n2652;
    wire n2655;
    wire n2658;
    wire n2661;
    wire n2664;
    wire n2667;
    wire n2670;
    wire n2673;
    wire n2676;
    wire n2679;
    wire n2682;
    wire n2684;
    wire n2687;
    wire n2690;
    wire n2693;
    wire n2696;
    wire n2699;
    wire n2702;
    wire n2705;
    wire n2708;
    wire n2711;
    wire n2714;
    wire n2717;
    wire n2720;
    wire n2723;
    wire n2726;
    wire n2730;
    wire n2733;
    wire n2736;
    wire n2739;
    wire n2742;
    wire n2745;
    wire n2748;
    wire n2751;
    wire n2754;
    wire n2757;
    wire n2760;
    wire n2763;
    wire n2766;
    wire n2769;
    wire n2772;
    wire n2775;
    wire n2778;
    wire n2781;
    wire n2784;
    wire n2787;
    wire n2790;
    wire n2793;
    wire n2796;
    wire n2799;
    wire n2802;
    wire n2805;
    wire n2808;
    wire n2811;
    wire n2814;
    wire n2817;
    wire n2820;
    wire n2823;
    wire n2826;
    wire n2829;
    wire n2832;
    wire n2835;
    wire n2838;
    wire n2841;
    wire n2844;
    wire n2847;
    wire n2850;
    wire n2853;
    wire n2856;
    wire n2859;
    wire n2862;
    wire n2865;
    wire n2868;
    wire n2871;
    wire n2874;
    wire n2877;
    wire n2880;
    wire n2883;
    wire n2886;
    wire n2889;
    wire n2892;
    wire n2895;
    wire n2898;
    wire n2900;
    wire n2903;
    wire n2906;
    wire n2909;
    wire n2912;
    wire n2915;
    wire n2919;
    wire n2922;
    wire n2924;
    wire n2927;
    wire n2930;
    wire n2933;
    wire n2936;
    wire n2939;
    wire n2942;
    wire n2945;
    wire n2948;
    wire n2952;
    wire n2954;
    wire n2957;
    wire n2960;
    wire n2963;
    wire n2966;
    wire n2969;
    wire n2972;
    wire n2976;
    wire n2978;
    wire n2981;
    wire n2984;
    wire n2987;
    wire n2990;
    wire n2993;
    wire n2996;
    wire n2999;
    wire n3003;
    wire n3006;
    wire n3009;
    wire n3012;
    wire n3015;
    wire n3018;
    wire n3021;
    wire n3024;
    wire n3027;
    wire n3030;
    wire n3033;
    wire n3036;
    wire n3039;
    wire n3042;
    wire n3045;
    wire n3048;
    wire n3051;
    wire n3054;
    wire n3057;
    wire n3060;
    wire n3063;
    wire n3066;
    wire n3069;
    wire n3072;
    wire n3075;
    wire n3078;
    wire n3081;
    wire n3084;
    wire n3087;
    wire n3090;
    wire n3093;
    wire n3096;
    wire n3099;
    wire n3102;
    wire n3105;
    wire n3108;
    wire n3111;
    wire n3114;
    wire n3117;
    wire n3120;
    wire n3123;
    wire n3125;
    wire n3128;
    wire n3131;
    wire n3134;
    wire n3137;
    wire n3140;
    wire n3143;
    wire n3146;
    wire n3149;
    wire n3152;
    wire n3155;
    wire n3158;
    wire n3161;
    wire n3164;
    wire n3167;
    wire n3171;
    wire n3174;
    wire n3176;
    wire n3179;
    wire n3183;
    wire n3185;
    wire n3188;
    wire n3191;
    wire n3194;
    wire n3198;
    wire n3201;
    wire n3203;
    wire n3206;
    wire n3210;
    wire n3212;
    wire n3215;
    wire n3219;
    wire n3221;
    wire n3224;
    wire n3227;
    wire n3230;
    wire n3233;
    wire n3236;
    wire n3240;
    wire n3243;
    wire n3246;
    wire n3248;
    wire n3251;
    wire n3255;
    wire n3257;
    wire n3260;
    wire n3264;
    wire n3266;
    wire n3269;
    wire n3272;
    wire n3275;
    wire n3279;
    wire n3281;
    wire n3284;
    wire n3287;
    wire n3290;
    wire n3294;
    wire n3297;
    wire n3300;
    wire n3303;
    wire n3306;
    wire n3308;
    wire n3311;
    wire n3314;
    wire n3317;
    wire n3320;
    wire n3323;
    wire n3326;
    wire n3329;
    wire n3332;
    wire n3335;
    wire n3338;
    wire n3341;
    wire n3345;
    wire n3348;
    wire n3350;
    wire n3353;
    wire n3356;
    wire n3359;
    wire n3363;
    wire n3366;
    wire n3369;
    wire n3372;
    wire n3375;
    wire n3377;
    wire n3380;
    wire n3383;
    wire n3386;
    wire n3389;
    wire n3392;
    wire n3395;
    wire n3398;
    wire n3401;
    wire n3404;
    wire n3407;
    wire n3410;
    wire n3414;
    wire n3417;
    wire n3419;
    wire n3422;
    wire n3425;
    wire n3428;
    wire n3431;
    wire n3434;
    wire n3437;
    wire n3440;
    wire n3443;
    wire n3446;
    wire n3449;
    wire n3452;
    wire n3455;
    wire n3458;
    wire n3461;
    wire n3464;
    wire n3467;
    wire n3470;
    wire n3474;
    wire n3477;
    wire n3480;
    wire n3483;
    wire n3485;
    wire n3488;
    wire n3491;
    wire n3494;
    wire n3497;
    wire n3500;
    wire n3504;
    wire n3507;
    wire n3509;
    wire n3512;
    wire n3515;
    wire n3518;
    wire n3521;
    wire n3524;
    wire n3528;
    wire n3530;
    wire n3533;
    wire n3536;
    wire n3539;
    wire n3542;
    wire n3545;
    wire n3548;
    wire n3551;
    wire n3554;
    wire n3557;
    wire n3560;
    wire n3563;
    wire n3566;
    wire n3569;
    wire n3572;
    wire n3575;
    wire n3578;
    wire n3581;
    wire n3584;
    wire n3587;
    wire n3590;
    wire n3593;
    wire n3596;
    wire n3599;
    wire n3602;
    wire n3605;
    wire n3608;
    wire n3611;
    wire n3615;
    wire n3618;
    wire n3620;
    wire n3623;
    wire n3626;
    wire n3629;
    wire n3632;
    wire n3635;
    wire n3638;
    wire n3641;
    wire n3644;
    wire n3647;
    wire n3650;
    wire n3654;
    wire n3657;
    wire n3660;
    wire n3663;
    wire n3665;
    wire n3668;
    wire n3671;
    wire n3674;
    wire n3677;
    wire n3680;
    wire n3683;
    wire n3686;
    wire n3689;
    wire n3692;
    wire n3695;
    wire n3698;
    wire n3701;
    wire n3704;
    wire n3707;
    wire n3711;
    wire n3714;
    wire n3717;
    wire n3720;
    wire n3723;
    wire n3726;
    wire n3728;
    wire n3731;
    wire n3734;
    wire n3737;
    wire n3740;
    wire n3743;
    wire n3746;
    wire n3749;
    wire n3752;
    wire n3755;
    wire n3758;
    wire n3761;
    wire n3764;
    wire n3767;
    wire n3770;
    wire n3773;
    wire n3776;
    wire n3779;
    wire n3783;
    wire n3786;
    wire n3789;
    wire n3792;
    wire n3795;
    wire n3798;
    wire n3800;
    wire n3803;
    wire n3806;
    wire n3809;
    wire n3812;
    wire n3815;
    wire n3818;
    wire n3821;
    wire n3824;
    wire n3827;
    wire n3830;
    wire n3833;
    wire n3837;
    wire n3840;
    wire n3843;
    wire n3845;
    wire n3848;
    wire n3851;
    wire n3854;
    wire n3857;
    wire n3860;
    wire n3863;
    wire n3866;
    wire n3869;
    wire n3872;
    wire n3875;
    wire n3878;
    wire n3881;
    wire n3884;
    wire n3887;
    wire n3890;
    wire n3893;
    wire n3896;
    wire n3900;
    wire n3903;
    wire n3906;
    wire n3908;
    wire n3911;
    wire n3914;
    wire n3917;
    wire n3921;
    wire n3923;
    wire n3926;
    wire n3929;
    wire n3932;
    wire n3935;
    wire n3938;
    wire n3941;
    wire n3944;
    wire n3947;
    wire n3951;
    wire n3954;
    wire n3957;
    wire n3959;
    wire n3962;
    wire n3965;
    wire n3968;
    wire n3971;
    wire n3974;
    wire n3977;
    wire n3980;
    wire n3983;
    wire n3986;
    wire n3989;
    wire n3992;
    wire n3996;
    wire n3998;
    wire n4001;
    wire n4004;
    wire n4007;
    wire n4010;
    wire n4013;
    wire n4016;
    wire n4019;
    wire n4022;
    wire n4025;
    wire n4028;
    wire n4031;
    wire n4034;
    wire n4037;
    wire n4041;
    wire n4043;
    wire n4046;
    wire n4049;
    wire n4052;
    wire n4055;
    wire n4058;
    wire n4061;
    wire n4064;
    wire n4067;
    wire n4070;
    wire n4073;
    wire n4076;
    wire n4079;
    wire n4083;
    wire n4085;
    wire n4088;
    wire n4091;
    wire n4094;
    wire n4097;
    wire n4100;
    wire n4103;
    wire n4106;
    wire n4109;
    wire n4112;
    wire n4115;
    wire n4118;
    wire n4121;
    wire n4124;
    wire n4127;
    wire n4130;
    wire n4133;
    wire n4136;
    wire n4139;
    wire n4142;
    wire n4145;
    wire n4148;
    wire n4151;
    wire n4154;
    wire n4157;
    wire n4160;
    wire n4163;
    wire n4166;
    wire n4169;
    wire n4172;
    wire n4175;
    wire n4178;
    wire n4181;
    wire n4184;
    wire n4187;
    wire n4190;
    wire n4193;
    wire n4196;
    wire n4199;
    wire n4202;
    wire n4205;
    wire n4208;
    wire n4211;
    wire n4214;
    wire n4217;
    wire n4220;
    wire n4223;
    wire n4226;
    wire n4229;
    wire n4232;
    wire n4235;
    wire n4238;
    wire n4241;
    wire n4244;
    wire n4247;
    wire n4250;
    wire n4253;
    wire n4256;
    wire n4259;
    wire n4262;
    wire n4265;
    wire n4268;
    wire n4271;
    wire n4274;
    wire n4277;
    wire n4280;
    wire n4283;
    wire n4286;
    wire n4289;
    wire n4292;
    wire n4295;
    wire n4298;
    wire n4301;
    wire n4304;
    wire n4307;
    wire n4310;
    wire n4313;
    wire n4316;
    wire n4319;
    wire n4322;
    wire n4325;
    wire n4328;
    wire n4331;
    wire n4334;
    wire n4337;
    wire n4340;
    wire n4343;
    wire n4346;
    wire n4349;
    wire n4352;
    wire n4355;
    wire n4358;
    wire n4361;
    wire n4364;
    wire n4367;
    wire n4370;
    wire n4373;
    wire n4376;
    wire n4379;
    wire n4382;
    wire n4385;
    wire n4388;
    wire n4391;
    wire n4394;
    wire n4397;
    wire n4400;
    wire n4403;
    wire n4406;
    wire n4409;
    wire n4412;
    wire n4415;
    wire n4418;
    wire n4421;
    wire n4424;
    wire n4427;
    wire n4430;
    wire n4433;
    wire n4436;
    wire n4439;
    wire n4442;
    wire n4445;
    wire n4448;
    wire n4451;
    wire n4454;
    wire n4457;
    wire n4460;
    wire n4463;
    wire n4466;
    wire n4469;
    wire n4472;
    wire n4475;
    wire n4478;
    wire n4481;
    wire n4484;
    wire n4487;
    wire n4490;
    wire n4493;
    wire n4496;
    wire n4499;
    wire n4502;
    wire n4505;
    wire n4508;
    wire n4511;
    wire n4514;
    wire n4517;
    wire n4520;
    wire n4523;
    wire n4526;
    wire n4529;
    wire n4532;
    wire n4536;
    wire n4538;
    wire n4541;
    wire n4544;
    wire n4547;
    wire n4550;
    wire n4553;
    wire n4556;
    wire n4559;
    wire n4562;
    wire n4565;
    wire n4568;
    wire n4571;
    wire n4574;
    wire n4577;
    wire n4580;
    wire n4583;
    wire n4586;
    wire n4589;
    wire n4592;
    wire n4595;
    wire n4598;
    wire n4601;
    wire n4604;
    wire n4607;
    wire n4610;
    wire n4613;
    wire n4616;
    wire n4619;
    wire n4622;
    wire n4625;
    wire n4628;
    wire n4631;
    wire n4634;
    wire n4637;
    wire n4640;
    wire n4643;
    wire n4646;
    wire n4650;
    wire n4652;
    wire n4655;
    wire n4658;
    wire n4661;
    wire n4664;
    wire n4667;
    wire n4670;
    wire n4673;
    wire n4676;
    wire n4679;
    wire n4682;
    wire n4685;
    wire n4688;
    wire n4691;
    wire n4694;
    wire n4697;
    wire n4700;
    wire n4703;
    wire n4706;
    wire n4709;
    wire n4712;
    wire n4715;
    wire n4718;
    wire n4721;
    wire n4724;
    wire n4727;
    wire n4730;
    wire n4733;
    wire n4736;
    wire n4739;
    wire n4742;
    wire n4745;
    wire n4748;
    wire n4751;
    wire n4754;
    wire n4757;
    wire n4760;
    wire n4763;
    wire n4766;
    wire n4769;
    wire n4772;
    wire n4775;
    wire n4778;
    wire n4781;
    wire n4784;
    wire n4787;
    wire n4790;
    wire n4793;
    wire n4796;
    wire n4799;
    wire n4802;
    wire n4805;
    wire n4808;
    wire n4811;
    wire n4814;
    wire n4817;
    wire n4820;
    wire n4823;
    wire n4826;
    wire n4829;
    wire n4832;
    wire n4835;
    wire n4838;
    wire n4841;
    wire n4845;
    wire n4847;
    wire n4850;
    wire n4853;
    wire n4856;
    wire n4859;
    wire n4862;
    wire n4865;
    wire n4868;
    wire n4871;
    wire n4874;
    wire n4877;
    wire n4880;
    wire n4883;
    wire n4886;
    wire n4889;
    wire n4892;
    wire n4895;
    wire n4898;
    wire n4904;
    wire n4907;
    wire n4910;
    wire n4913;
    wire n4916;
    wire n4919;
    wire n4925;
    wire n4928;
    wire n4931;
    wire n4934;
    wire n4937;
    wire n4940;
    wire n4946;
    wire n4949;
    wire n4952;
    wire n4955;
    wire n4958;
    wire n4961;
    wire n4967;
    wire n4970;
    wire n4973;
    wire n4976;
    wire n4979;
    wire n4982;
    wire n4988;
    wire n4991;
    wire n4994;
    wire n4997;
    wire n5000;
    wire n5003;
    wire n5009;
    wire n5012;
    wire n5015;
    wire n5018;
    wire n5021;
    wire n5024;
    wire n5030;
    wire n5033;
    wire n5036;
    wire n5039;
    wire n5042;
    wire n5045;
    wire n5051;
    wire n5054;
    wire n5057;
    wire n5060;
    wire n5063;
    wire n5066;
    wire n5072;
    wire n5075;
    wire n5078;
    wire n5081;
    wire n5084;
    wire n5087;
    wire n5093;
    wire n5096;
    wire n5099;
    wire n5102;
    wire n5105;
    wire n5108;
    wire n5114;
    wire n5117;
    wire n5120;
    wire n5123;
    wire n5126;
    wire n5129;
    wire n5135;
    wire n5138;
    wire n5141;
    wire n5144;
    wire n5147;
    wire n5150;
    wire n5156;
    wire n5159;
    wire n5162;
    wire n5165;
    wire n5168;
    wire n5171;
    wire n5177;
    wire n5180;
    wire n5183;
    wire n5186;
    wire n5189;
    wire n5192;
    wire n5198;
    wire n5201;
    wire n5204;
    wire n5207;
    wire n5210;
    wire n5213;
    wire n5225;
    jnot g000(.din(G146), .dout(n60));
    jxor g001(.dinb(G125), .dina(G140), .dout(n64));
    jxor g002(.dinb(n60), .dina(n64), .dout(n68));
    jdff g003(.din(G953), .dout(n71));
    jand g004(.dinb(n3938), .dina(n71), .dout(n75));
    jand g005(.dinb(n3941), .dina(n75), .dout(n79));
    jxor g006(.dinb(n4838), .dina(n79), .dout(n83));
    jxor g007(.dinb(G119), .dina(G128), .dout(n87));
    jor g008(.dinb(n83), .dina(n3726), .dout(n91));
    jxor g009(.dinb(n4205), .dina(n91), .dout(n95));
    jxor g010(.dinb(n3728), .dina(n95), .dout(n99));
    jor g011(.dinb(n4310), .dina(n99), .dout(n103));
    jnot g012(.din(G902), .dout(n106));
    jand g013(.dinb(n3935), .dina(n106), .dout(n110));
    jnot g014(.din(n110), .dout(n113));
    jand g015(.dinb(n3671), .dina(n113), .dout(n117));
    jxor g016(.dinb(n103), .dina(n3663), .dout(n121));
    jnot g017(.din(G134), .dout(n124));
    jxor g018(.dinb(n124), .dina(n4845), .dout(n128));
    jnot g019(.din(G131), .dout(n131));
    jxor g020(.dinb(G143), .dina(G146), .dout(n135));
    jxor g021(.dinb(n4727), .dina(n135), .dout(n139));
    jxor g022(.dinb(n4766), .dina(n139), .dout(n143));
    jxor g023(.dinb(n4650), .dina(n143), .dout(n147));
    jnot g024(.din(G113), .dout(n150));
    jxor g025(.dinb(G116), .dina(G119), .dout(n154));
    jxor g026(.dinb(n150), .dina(n154), .dout(n158));
    jnot g027(.din(G210), .dout(n161));
    jor g028(.dinb(G237), .dina(G953), .dout(n165));
    jor g029(.dinb(n161), .dina(n165), .dout(n169));
    jxor g030(.dinb(n4532), .dina(n169), .dout(n173));
    jxor g031(.dinb(n4538), .dina(n173), .dout(n177));
    jxor g032(.dinb(n147), .dina(n177), .dout(n181));
    jand g033(.dinb(n3923), .dina(n181), .dout(n185));
    jxor g034(.dinb(n3635), .dina(n185), .dout(n189));
    jand g035(.dinb(n121), .dina(n3272), .dout(n193));
    jor g036(.dinb(G237), .dina(G902), .dout(n197));
    jand g037(.dinb(n4331), .dina(n197), .dout(n201));
    jnot g038(.din(n201), .dout(n204));
    jand g039(.dinb(n4496), .dina(n197), .dout(n208));
    jnot g040(.din(G110), .dout(n211));
    jxor g041(.dinb(n211), .dina(n4163), .dout(n215));
    jxor g042(.dinb(G104), .dina(G107), .dout(n219));
    jxor g043(.dinb(n4536), .dina(n219), .dout(n223));
    jxor g044(.dinb(n158), .dina(n223), .dout(n227));
    jxor g045(.dinb(n4083), .dina(n227), .dout(n231));
    jand g046(.dinb(n4041), .dina(n71), .dout(n235));
    jxor g047(.dinb(n4034), .dina(n139), .dout(n239));
    jxor g048(.dinb(n3996), .dina(n239), .dout(n243));
    jxor g049(.dinb(n231), .dina(n243), .dout(n247));
    jand g050(.dinb(n4256), .dina(n247), .dout(n251));
    jxor g051(.dinb(n4268), .dina(n251), .dout(n255));
    jand g052(.dinb(n2990), .dina(n255), .dout(n259));
    jnot g053(.din(G221), .dout(n262));
    jor g054(.dinb(n3921), .dina(n110), .dout(n266));
    jxor g055(.dinb(G110), .dina(G140), .dout(n270));
    jand g056(.dinb(n3843), .dina(n71), .dout(n274));
    jxor g057(.dinb(n223), .dina(n274), .dout(n278));
    jxor g058(.dinb(n3840), .dina(n278), .dout(n282));
    jxor g059(.dinb(n147), .dina(n282), .dout(n286));
    jand g060(.dinb(n4256), .dina(n286), .dout(n290));
    jxor g061(.dinb(n3881), .dina(n290), .dout(n294));
    jand g062(.dinb(n3908), .dina(n294), .dout(n298));
    jand g063(.dinb(n259), .dina(n298), .dout(n302));
    jand g064(.dinb(n193), .dina(n2976), .dout(n306));
    jnot g065(.din(G478), .dout(n309));
    jxor g066(.dinb(G128), .dina(G143), .dout(n313));
    jand g067(.dinb(n3665), .dina(n75), .dout(n317));
    jxor g068(.dinb(G116), .dina(G122), .dout(n321));
    jxor g069(.dinb(G107), .dina(G134), .dout(n325));
    jxor g070(.dinb(n321), .dina(n325), .dout(n329));
    jxor g071(.dinb(n317), .dina(n3483), .dout(n333));
    jxor g072(.dinb(n3480), .dina(n333), .dout(n337));
    jand g073(.dinb(n4256), .dina(n337), .dout(n341));
    jxor g074(.dinb(n3306), .dina(n341), .dout(n345));
    jnot g075(.din(G475), .dout(n348));
    jxor g076(.dinb(n131), .dina(n4724), .dout(n352));
    jxor g077(.dinb(n150), .dina(n4202), .dout(n356));
    jxor g078(.dinb(n4157), .dina(n356), .dout(n360));
    jnot g079(.din(G214), .dout(n363));
    jor g080(.dinb(n363), .dina(n165), .dout(n367));
    jxor g081(.dinb(n68), .dina(n367), .dout(n371));
    jxor g082(.dinb(n360), .dina(n371), .dout(n375));
    jxor g083(.dinb(n3417), .dina(n375), .dout(n379));
    jand g084(.dinb(n3767), .dina(n379), .dout(n383));
    jxor g085(.dinb(n3375), .dina(n383), .dout(n387));
    jand g086(.dinb(n345), .dina(n387), .dout(n391));
    jor g087(.dinb(n3618), .dina(n71), .dout(n395));
    jand g088(.dinb(G234), .dina(G237), .dout(n399));
    jor g089(.dinb(n106), .dina(n399), .dout(n403));
    jor g090(.dinb(n395), .dina(n403), .dout(n407));
    jnot g091(.din(n399), .dout(n410));
    jand g092(.dinb(n3615), .dina(n71), .dout(n414));
    jand g093(.dinb(n410), .dina(n414), .dout(n418));
    jnot g094(.din(n418), .dout(n421));
    jand g095(.dinb(n3528), .dina(n421), .dout(n425));
    jnot g096(.din(n425), .dout(n428));
    jand g097(.dinb(n391), .dina(n3507), .dout(n432));
    jand g098(.dinb(n306), .dina(n2948), .dout(n436));
    jxor g099(.dinb(n4499), .dina(n436), .dout(n440));
    jnot g100(.din(n189), .dout(n443));
    jand g101(.dinb(n121), .dina(n3264), .dout(n447));
    jand g102(.dinb(n2976), .dina(n447), .dout(n451));
    jxor g103(.dinb(n3419), .dina(n383), .dout(n455));
    jand g104(.dinb(n345), .dina(n455), .dout(n459));
    jand g105(.dinb(n3507), .dina(n459), .dout(n463));
    jand g106(.dinb(n451), .dina(n3287), .dout(n467));
    jxor g107(.dinb(n4121), .dina(n467), .dout(n471));
    jxor g108(.dinb(n3485), .dina(n341), .dout(n475));
    jand g109(.dinb(n475), .dina(n387), .dout(n479));
    jand g110(.dinb(n3507), .dina(n479), .dout(n483));
    jand g111(.dinb(n451), .dina(n3356), .dout(n487));
    jxor g112(.dinb(n4085), .dina(n487), .dout(n491));
    jnot g113(.din(n68), .dout(n494));
    jxor g114(.dinb(n3717), .dina(n95), .dout(n498));
    jand g115(.dinb(n3749), .dina(n498), .dout(n502));
    jxor g116(.dinb(n502), .dina(n3663), .dout(n506));
    jand g117(.dinb(n506), .dina(n3264), .dout(n510));
    jand g118(.dinb(n2952), .dina(n510), .dout(n514));
    jand g119(.dinb(n2972), .dina(n514), .dout(n518));
    jxor g120(.dinb(n4220), .dina(n518), .dout(n522));
    jand g121(.dinb(n506), .dina(n3266), .dout(n526));
    jand g122(.dinb(n2976), .dina(n526), .dout(n530));
    jor g123(.dinb(n3243), .dina(n71), .dout(n534));
    jor g124(.dinb(n403), .dina(n534), .dout(n538));
    jand g125(.dinb(n421), .dina(n3240), .dout(n542));
    jnot g126(.din(n542), .dout(n545));
    jand g127(.dinb(n479), .dina(n3201), .dout(n549));
    jand g128(.dinb(n530), .dina(n3191), .dout(n553));
    jxor g129(.dinb(n4730), .dina(n553), .dout(n557));
    jand g130(.dinb(n475), .dina(n455), .dout(n561));
    jand g131(.dinb(n3201), .dina(n561), .dout(n565));
    jand g132(.dinb(n306), .dina(n3176), .dout(n569));
    jxor g133(.dinb(n4688), .dina(n569), .dout(n573));
    jand g134(.dinb(n459), .dina(n3201), .dout(n577));
    jand g135(.dinb(n530), .dina(n2915), .dout(n581));
    jxor g136(.dinb(n4652), .dina(n581), .dout(n585));
    jnot g137(.din(G469), .dout(n588));
    jxor g138(.dinb(n3798), .dina(n290), .dout(n592));
    jand g139(.dinb(n3908), .dina(n592), .dout(n596));
    jand g140(.dinb(n259), .dina(n596), .dout(n600));
    jand g141(.dinb(n193), .dina(n2924), .dout(n604));
    jand g142(.dinb(n3281), .dina(n604), .dout(n608));
    jxor g143(.dinb(n4613), .dina(n608), .dout(n612));
    jand g144(.dinb(n3350), .dina(n604), .dout(n616));
    jxor g145(.dinb(n4577), .dina(n616), .dout(n620));
    jand g146(.dinb(n526), .dina(n2924), .dout(n624));
    jand g147(.dinb(n2945), .dina(n624), .dout(n628));
    jxor g148(.dinb(n4541), .dina(n628), .dout(n632));
    jand g149(.dinb(n447), .dina(n2933), .dout(n636));
    jand g150(.dinb(n259), .dina(n3507), .dout(n640));
    jand g151(.dinb(n3248), .dina(n640), .dout(n644));
    jand g152(.dinb(n636), .dina(n2922), .dout(n648));
    jxor g153(.dinb(n4166), .dina(n648), .dout(n652));
    jand g154(.dinb(n510), .dina(n2919), .dout(n656));
    jand g155(.dinb(n2927), .dina(n656), .dout(n660));
    jxor g156(.dinb(n3998), .dina(n660), .dout(n664));
    jnot g157(.din(n208), .dout(n667));
    jxor g158(.dinb(n3957), .dina(n251), .dout(n671));
    jand g159(.dinb(n2978), .dina(n671), .dout(n675));
    jand g160(.dinb(n298), .dina(n675), .dout(n679));
    jand g161(.dinb(n193), .dina(n2903), .dout(n683));
    jand g162(.dinb(n2912), .dina(n683), .dout(n687));
    jxor g163(.dinb(n4769), .dina(n687), .dout(n691));
    jand g164(.dinb(n3185), .dina(n683), .dout(n695));
    jxor g165(.dinb(n4847), .dina(n695), .dout(n699));
    jand g166(.dinb(n391), .dina(n3201), .dout(n703));
    jand g167(.dinb(n526), .dina(n2898), .dout(n707));
    jand g168(.dinb(n2900), .dina(n707), .dout(n711));
    jxor g169(.dinb(n4805), .dina(n711), .dout(n715));
    jand g170(.dinb(n656), .dina(n2906), .dout(n719));
    jxor g171(.dinb(n3845), .dina(n719), .dout(n723));
    jor g172(.dinb(n487), .dina(n518), .dout(n727));
    jor g173(.dinb(n467), .dina(n616), .dout(n731));
    jor g174(.dinb(n727), .dina(n731), .dout(n735));
    jor g175(.dinb(n436), .dina(n628), .dout(n739));
    jor g176(.dinb(n608), .dina(n648), .dout(n743));
    jor g177(.dinb(n739), .dina(n743), .dout(n747));
    jor g178(.dinb(n735), .dina(n747), .dout(n751));
    jor g179(.dinb(n581), .dina(n687), .dout(n755));
    jor g180(.dinb(n553), .dina(n695), .dout(n759));
    jor g181(.dinb(n755), .dina(n759), .dout(n763));
    jor g182(.dinb(n569), .dina(n719), .dout(n767));
    jor g183(.dinb(n660), .dina(n711), .dout(n771));
    jor g184(.dinb(n767), .dina(n771), .dout(n775));
    jor g185(.dinb(n763), .dina(n775), .dout(n779));
    jor g186(.dinb(n751), .dina(n779), .dout(n783));
    jor g187(.dinb(n600), .dina(n679), .dout(n787));
    jand g188(.dinb(n2954), .dina(n787), .dout(n791));
    jand g189(.dinb(n596), .dina(n675), .dout(n795));
    jxor g190(.dinb(n345), .dina(n387), .dout(n799));
    jand g191(.dinb(n795), .dina(n2145), .dout(n803));
    jor g192(.dinb(n791), .dina(n2142), .dout(n807));
    jand g193(.dinb(n2966), .dina(n807), .dout(n811));
    jand g194(.dinb(n391), .dina(n675), .dout(n815));
    jor g195(.dinb(n506), .dina(n3629), .dout(n819));
    jor g196(.dinb(n121), .dina(n3264), .dout(n823));
    jand g197(.dinb(n823), .dina(n2939), .dout(n827));
    jand g198(.dinb(n3620), .dina(n827), .dout(n831));
    jand g199(.dinb(n2132), .dina(n831), .dout(n835));
    jor g200(.dinb(n811), .dina(n835), .dout(n839));
    jand g201(.dinb(n3533), .dina(n839), .dout(n843));
    jxor g202(.dinb(n204), .dina(n266), .dout(n847));
    jand g203(.dinb(n3530), .dina(n847), .dout(n851));
    jand g204(.dinb(n592), .dina(n2130), .dout(n855));
    jand g205(.dinb(n3947), .dina(n855), .dout(n859));
    jand g206(.dinb(n2960), .dina(n447), .dout(n863));
    jand g207(.dinb(n2124), .dina(n863), .dout(n867));
    jor g208(.dinb(n843), .dina(n2118), .dout(n871));
    jor g209(.dinb(n783), .dina(n871), .dout(n875));
    jand g210(.dinb(n3566), .dina(n875), .dout(n879));
    jand g211(.dinb(n636), .dina(n2139), .dout(n883));
    jor g212(.dinb(n4370), .dina(n883), .dout(n887));
    jor g213(.dinb(n879), .dina(n2109), .dout(n891));
    jnot g214(.din(n247), .dout(n894));
    jor g215(.dinb(n4295), .dina(n671), .dout(n898));
    jnot g216(.din(n266), .dout(n901));
    jor g217(.dinb(n3906), .dina(n592), .dout(n905));
    jor g218(.dinb(n898), .dina(n905), .dout(n909));
    jor g219(.dinb(n3783), .dina(n819), .dout(n913));
    jnot g220(.din(n483), .dout(n916));
    jor g221(.dinb(n913), .dina(n3348), .dout(n920));
    jor g222(.dinb(n475), .dina(n455), .dout(n924));
    jor g223(.dinb(n924), .dina(n3518), .dout(n928));
    jor g224(.dinb(n121), .dina(n3623), .dout(n932));
    jor g225(.dinb(n3345), .dina(n932), .dout(n936));
    jor g226(.dinb(n3779), .dina(n936), .dout(n940));
    jand g227(.dinb(n920), .dina(n940), .dout(n944));
    jnot g228(.din(n463), .dout(n947));
    jor g229(.dinb(n913), .dina(n3279), .dout(n951));
    jor g230(.dinb(n506), .dina(n3264), .dout(n955));
    jor g231(.dinb(n3906), .dina(n294), .dout(n959));
    jor g232(.dinb(n898), .dina(n959), .dout(n963));
    jor g233(.dinb(n955), .dina(n3255), .dout(n967));
    jor g234(.dinb(n3348), .dina(n967), .dout(n971));
    jand g235(.dinb(n951), .dina(n971), .dout(n975));
    jand g236(.dinb(n944), .dina(n975), .dout(n979));
    jor g237(.dinb(n955), .dina(n3783), .dout(n983));
    jor g238(.dinb(n983), .dina(n3341), .dout(n987));
    jor g239(.dinb(n823), .dina(n3255), .dout(n991));
    jor g240(.dinb(n3338), .dina(n991), .dout(n995));
    jand g241(.dinb(n987), .dina(n995), .dout(n999));
    jor g242(.dinb(n3279), .dina(n967), .dout(n1003));
    jor g243(.dinb(n819), .dina(n3257), .dout(n1007));
    jnot g244(.din(n561), .dout(n1010));
    jor g245(.dinb(n898), .dina(n3509), .dout(n1014));
    jor g246(.dinb(n1010), .dina(n1014), .dout(n1018));
    jor g247(.dinb(n1007), .dina(n3246), .dout(n1022));
    jand g248(.dinb(n1003), .dina(n1022), .dout(n1026));
    jand g249(.dinb(n999), .dina(n1026), .dout(n1030));
    jand g250(.dinb(n979), .dina(n1030), .dout(n1034));
    jor g251(.dinb(n3783), .dina(n823), .dout(n1038));
    jor g252(.dinb(n475), .dina(n387), .dout(n1042));
    jor g253(.dinb(n1042), .dina(n3230), .dout(n1046));
    jor g254(.dinb(n1038), .dina(n3215), .dout(n1050));
    jor g255(.dinb(n4280), .dina(n255), .dout(n1054));
    jor g256(.dinb(n905), .dina(n1054), .dout(n1058));
    jor g257(.dinb(n955), .dina(n3210), .dout(n1062));
    jor g258(.dinb(n3212), .dina(n1062), .dout(n1066));
    jand g259(.dinb(n1050), .dina(n1066), .dout(n1070));
    jnot g260(.din(n549), .dout(n1073));
    jor g261(.dinb(n1038), .dina(n3183), .dout(n1077));
    jor g262(.dinb(n3183), .dina(n1062), .dout(n1081));
    jand g263(.dinb(n1077), .dina(n1081), .dout(n1085));
    jand g264(.dinb(n1070), .dina(n1085), .dout(n1089));
    jnot g265(.din(n565), .dout(n1092));
    jor g266(.dinb(n983), .dina(n3174), .dout(n1096));
    jor g267(.dinb(n932), .dina(n3219), .dout(n1100));
    jor g268(.dinb(n1100), .dina(n3206), .dout(n1104));
    jand g269(.dinb(n1096), .dina(n1104), .dout(n1108));
    jor g270(.dinb(n3251), .dina(n1100), .dout(n1112));
    jor g271(.dinb(n924), .dina(n3221), .dout(n1116));
    jor g272(.dinb(n823), .dina(n3171), .dout(n1120));
    jor g273(.dinb(n3203), .dina(n1120), .dout(n1124));
    jand g274(.dinb(n1112), .dina(n1124), .dout(n1128));
    jand g275(.dinb(n1108), .dina(n1128), .dout(n1132));
    jand g276(.dinb(n1089), .dina(n1132), .dout(n1136));
    jand g277(.dinb(n1034), .dina(n1136), .dout(n1140));
    jand g278(.dinb(G210), .dina(G902), .dout(n1144));
    jnot g279(.din(n1144), .dout(n1147));
    jor g280(.dinb(n1140), .dina(n2223), .dout(n1151));
    jor g281(.dinb(n2181), .dina(n1151), .dout(n1155));
    jor g282(.dinb(n3615), .dina(n71), .dout(n1159));
    jand g283(.dinb(n783), .dina(n2225), .dout(n1163));
    jor g284(.dinb(n3959), .dina(n1163), .dout(n1167));
    jand g285(.dinb(n3048), .dina(n1167), .dout(n1171));
    jand g286(.dinb(n2148), .dina(n1171), .dout(G51));
    jnot g287(.din(n286), .dout(n1178));
    jand g288(.dinb(G469), .dina(G902), .dout(n1182));
    jnot g289(.din(n1182), .dout(n1185));
    jor g290(.dinb(n1140), .dina(n2346), .dout(n1189));
    jor g291(.dinb(n2304), .dina(n1189), .dout(n1193));
    jand g292(.dinb(n783), .dina(n2348), .dout(n1197));
    jor g293(.dinb(n3800), .dina(n1197), .dout(n1201));
    jand g294(.dinb(n3048), .dina(n1201), .dout(n1205));
    jand g295(.dinb(n2271), .dina(n1205), .dout(G54));
    jnot g296(.din(n379), .dout(n1212));
    jand g297(.dinb(G475), .dina(G902), .dout(n1216));
    jnot g298(.din(n1216), .dout(n1219));
    jor g299(.dinb(n1140), .dina(n2469), .dout(n1223));
    jor g300(.dinb(n2427), .dina(n1223), .dout(n1227));
    jand g301(.dinb(n783), .dina(n2471), .dout(n1231));
    jor g302(.dinb(n3377), .dina(n1231), .dout(n1235));
    jand g303(.dinb(n3048), .dina(n1235), .dout(n1239));
    jand g304(.dinb(n2394), .dina(n1239), .dout(G60));
    jnot g305(.din(n337), .dout(n1246));
    jand g306(.dinb(G478), .dina(G902), .dout(n1250));
    jnot g307(.din(n1250), .dout(n1253));
    jor g308(.dinb(n1140), .dina(n2592), .dout(n1257));
    jor g309(.dinb(n2550), .dina(n1257), .dout(n1261));
    jand g310(.dinb(n783), .dina(n2594), .dout(n1265));
    jor g311(.dinb(n3437), .dina(n1265), .dout(n1269));
    jand g312(.dinb(n3048), .dina(n1269), .dout(n1273));
    jand g313(.dinb(n2517), .dina(n1273), .dout(G63));
    jand g314(.dinb(G217), .dina(G902), .dout(n1281));
    jand g315(.dinb(n783), .dina(n2684), .dout(n1285));
    jor g316(.dinb(n3680), .dina(n1285), .dout(n1289));
    jnot g317(.din(n1281), .dout(n1292));
    jor g318(.dinb(n1140), .dina(n2682), .dout(n1296));
    jor g319(.dinb(n3308), .dina(n1296), .dout(n1300));
    jand g320(.dinb(n3048), .dina(n1300), .dout(n1304));
    jand g321(.dinb(n2640), .dina(n1304), .dout(G66));
    jnot g322(.din(n395), .dout(n1311));
    jor g323(.dinb(n4451), .dina(n1034), .dout(n1315));
    jor g324(.dinb(n4041), .dina(n71), .dout(n1319));
    jand g325(.dinb(n1315), .dina(n2814), .dout(n1323));
    jxor g326(.dinb(n4043), .dina(n1323), .dout(n1327));
    jor g327(.dinb(n2772), .dina(n1327), .dout(n1331));
    jor g328(.dinb(n4406), .dina(n1136), .dout(n1335));
    jor g329(.dinb(n3843), .dina(n71), .dout(n1339));
    jand g330(.dinb(n534), .dina(n1339), .dout(n1343));
    jand g331(.dinb(n1335), .dina(n2892), .dout(n1347));
    jnot g332(.din(n534), .dout(n1350));
    jxor g333(.dinb(n3740), .dina(n147), .dout(n1354));
    jor g334(.dinb(n2853), .dina(n1354), .dout(n1358));
    jxor g335(.dinb(n1347), .dina(n2847), .dout(n1362));
    jnot g336(.din(n181), .dout(n1365));
    jand g337(.dinb(G472), .dina(G902), .dout(n1369));
    jnot g338(.din(n1369), .dout(n1372));
    jor g339(.dinb(n1140), .dina(n3123), .dout(n1376));
    jor g340(.dinb(n3081), .dina(n1376), .dout(n1380));
    jand g341(.dinb(n783), .dina(n3125), .dout(n1384));
    jor g342(.dinb(n4334), .dina(n1384), .dout(n1388));
    jand g343(.dinb(n3048), .dina(n1388), .dout(n1392));
    jand g344(.dinb(n2895), .dina(n1392), .dout(G57));
    jdff dff_A_PknvDO025_0(.din(n5225), .dout(G72));
    jdff dff_A_BblxUM767_2(.din(n1362), .dout(n5225));
    jdff dff_A_STzXy76t1_2(.din(n1331), .dout(G69));
    jdff dff_A_76IhHjB45_2(.din(n891), .dout(G75));
    jdff dff_A_Y2dIFbtx4_0(.din(n5213), .dout(G42));
    jdff dff_A_8OmdQrkT4_0(.din(n5210), .dout(n5213));
    jdff dff_A_7f5mwdfI9_0(.din(n5207), .dout(n5210));
    jdff dff_A_axJWYsxJ5_0(.din(n5204), .dout(n5207));
    jdff dff_A_EzXgRwKQ9_0(.din(n5201), .dout(n5204));
    jdff dff_A_M4OfibrF1_0(.din(n5198), .dout(n5201));
    jdff dff_A_5MAg6puK2_2(.din(n723), .dout(n5198));
    jdff dff_A_teud1nbE4_0(.din(n5192), .dout(G39));
    jdff dff_A_hm112p493_0(.din(n5189), .dout(n5192));
    jdff dff_A_vT75EyGY5_0(.din(n5186), .dout(n5189));
    jdff dff_A_DHl6Y7IQ9_0(.din(n5183), .dout(n5186));
    jdff dff_A_0hRpRr789_0(.din(n5180), .dout(n5183));
    jdff dff_A_BQvTciW99_0(.din(n5177), .dout(n5180));
    jdff dff_A_5ZGcPxwR6_2(.din(n715), .dout(n5177));
    jdff dff_A_sZZkANDc0_0(.din(n5171), .dout(G36));
    jdff dff_A_jp2Wqpe77_0(.din(n5168), .dout(n5171));
    jdff dff_A_1NG3OYxR8_0(.din(n5165), .dout(n5168));
    jdff dff_A_pI5WLpcv6_0(.din(n5162), .dout(n5165));
    jdff dff_A_Bz7H5Wjt7_0(.din(n5159), .dout(n5162));
    jdff dff_A_ilTLLlxC8_0(.din(n5156), .dout(n5159));
    jdff dff_A_wxTTumbh8_2(.din(n699), .dout(n5156));
    jdff dff_A_o6BgCzU64_0(.din(n5150), .dout(G33));
    jdff dff_A_Li6WKKvL4_0(.din(n5147), .dout(n5150));
    jdff dff_A_TMpfrc1Q8_0(.din(n5144), .dout(n5147));
    jdff dff_A_5gkAEx7I0_0(.din(n5141), .dout(n5144));
    jdff dff_A_xBgBFEHM7_0(.din(n5138), .dout(n5141));
    jdff dff_A_fy9LOIPT8_0(.din(n5135), .dout(n5138));
    jdff dff_A_XeL5ESXH3_2(.din(n691), .dout(n5135));
    jdff dff_A_mCHTSb2L3_0(.din(n5129), .dout(G27));
    jdff dff_A_xqSZaXoR3_0(.din(n5126), .dout(n5129));
    jdff dff_A_IhFQEkMO9_0(.din(n5123), .dout(n5126));
    jdff dff_A_cpS9pvUm5_0(.din(n5120), .dout(n5123));
    jdff dff_A_pVO7JxRf3_0(.din(n5117), .dout(n5120));
    jdff dff_A_muRMUgys2_0(.din(n5114), .dout(n5117));
    jdff dff_A_PCaNejM41_2(.din(n664), .dout(n5114));
    jdff dff_A_edZ4euLr7_0(.din(n5108), .dout(G24));
    jdff dff_A_lHlNJP5b7_0(.din(n5105), .dout(n5108));
    jdff dff_A_Aaedy9gb5_0(.din(n5102), .dout(n5105));
    jdff dff_A_4j4wXiaz0_0(.din(n5099), .dout(n5102));
    jdff dff_A_qJrzVuab9_0(.din(n5096), .dout(n5099));
    jdff dff_A_UI9HFpeL2_0(.din(n5093), .dout(n5096));
    jdff dff_A_VxBgzGut5_2(.din(n652), .dout(n5093));
    jdff dff_A_W8bPgPiJ6_0(.din(n5087), .dout(G21));
    jdff dff_A_xxeOSZzt9_0(.din(n5084), .dout(n5087));
    jdff dff_A_Q1qrKJZf1_0(.din(n5081), .dout(n5084));
    jdff dff_A_CAVjaFLi4_0(.din(n5078), .dout(n5081));
    jdff dff_A_fFYUbEWo4_0(.din(n5075), .dout(n5078));
    jdff dff_A_2jZUzQMO3_0(.din(n5072), .dout(n5075));
    jdff dff_A_Fko9CuZr6_2(.din(n632), .dout(n5072));
    jdff dff_A_JJWlIZNC0_0(.din(n5066), .dout(G18));
    jdff dff_A_8joY4mYZ5_0(.din(n5063), .dout(n5066));
    jdff dff_A_Tu2aKiaE8_0(.din(n5060), .dout(n5063));
    jdff dff_A_TrxtfwNt8_0(.din(n5057), .dout(n5060));
    jdff dff_A_d0NGJUAT7_0(.din(n5054), .dout(n5057));
    jdff dff_A_x7HgaYxP9_0(.din(n5051), .dout(n5054));
    jdff dff_A_OvTispEG5_2(.din(n620), .dout(n5051));
    jdff dff_A_h4SaEFY61_0(.din(n5045), .dout(G15));
    jdff dff_A_68iq09Iz0_0(.din(n5042), .dout(n5045));
    jdff dff_A_hi7LkfJQ5_0(.din(n5039), .dout(n5042));
    jdff dff_A_Ly8Z3pCD4_0(.din(n5036), .dout(n5039));
    jdff dff_A_sFpjpHVR7_0(.din(n5033), .dout(n5036));
    jdff dff_A_IExpIc7W2_0(.din(n5030), .dout(n5033));
    jdff dff_A_iA9pP22X1_2(.din(n612), .dout(n5030));
    jdff dff_A_pHmFZTGV1_0(.din(n5024), .dout(G48));
    jdff dff_A_WlEz4kmI8_0(.din(n5021), .dout(n5024));
    jdff dff_A_vt6MVxkA5_0(.din(n5018), .dout(n5021));
    jdff dff_A_BfppoD9q8_0(.din(n5015), .dout(n5018));
    jdff dff_A_D67fBNeB0_0(.din(n5012), .dout(n5015));
    jdff dff_A_lByYvY8H8_0(.din(n5009), .dout(n5012));
    jdff dff_A_CxV5R3S41_2(.din(n585), .dout(n5009));
    jdff dff_A_AYMvHAtF2_0(.din(n5003), .dout(G45));
    jdff dff_A_u7j7UB2c4_0(.din(n5000), .dout(n5003));
    jdff dff_A_ukcVafbV1_0(.din(n4997), .dout(n5000));
    jdff dff_A_CkySIeNS0_0(.din(n4994), .dout(n4997));
    jdff dff_A_QLAX8zKf4_0(.din(n4991), .dout(n4994));
    jdff dff_A_IaTZkgip1_0(.din(n4988), .dout(n4991));
    jdff dff_A_ehYWmLY91_2(.din(n573), .dout(n4988));
    jdff dff_A_ijmCbDwn1_0(.din(n4982), .dout(G30));
    jdff dff_A_ASjJGAdI0_0(.din(n4979), .dout(n4982));
    jdff dff_A_AY5bFrSp1_0(.din(n4976), .dout(n4979));
    jdff dff_A_U4KfyalL5_0(.din(n4973), .dout(n4976));
    jdff dff_A_9cQjYvRQ1_0(.din(n4970), .dout(n4973));
    jdff dff_A_QjzFVJyZ8_0(.din(n4967), .dout(n4970));
    jdff dff_A_3yefOgGp2_2(.din(n557), .dout(n4967));
    jdff dff_A_ZfoTHkX01_0(.din(n4961), .dout(G12));
    jdff dff_A_SOBVLc7F8_0(.din(n4958), .dout(n4961));
    jdff dff_A_scRGQsfY4_0(.din(n4955), .dout(n4958));
    jdff dff_A_pLYsoq2Q2_0(.din(n4952), .dout(n4955));
    jdff dff_A_FcBOieOs8_0(.din(n4949), .dout(n4952));
    jdff dff_A_R4yd7DBk4_0(.din(n4946), .dout(n4949));
    jdff dff_A_0f7i80Nd1_2(.din(n522), .dout(n4946));
    jdff dff_A_y16Uu0qQ7_0(.din(n4940), .dout(G9));
    jdff dff_A_5zyebfVW4_0(.din(n4937), .dout(n4940));
    jdff dff_A_STmyObGg3_0(.din(n4934), .dout(n4937));
    jdff dff_A_3aZ33zEw3_0(.din(n4931), .dout(n4934));
    jdff dff_A_AOZGbwPt8_0(.din(n4928), .dout(n4931));
    jdff dff_A_yM9yP70s3_0(.din(n4925), .dout(n4928));
    jdff dff_A_B8eR28a40_2(.din(n491), .dout(n4925));
    jdff dff_A_NWx4ToN48_0(.din(n4919), .dout(G6));
    jdff dff_A_PpPLHoD77_0(.din(n4916), .dout(n4919));
    jdff dff_A_3MEcD3C63_0(.din(n4913), .dout(n4916));
    jdff dff_A_fcLWlC2l7_0(.din(n4910), .dout(n4913));
    jdff dff_A_FLxDXH7i7_0(.din(n4907), .dout(n4910));
    jdff dff_A_h6B22lMB2_0(.din(n4904), .dout(n4907));
    jdff dff_A_1jvHz01S6_2(.din(n471), .dout(n4904));
    jdff dff_A_irGhth8U4_0(.din(n4898), .dout(G3));
    jdff dff_A_9CGrs0b87_0(.din(n4895), .dout(n4898));
    jdff dff_A_1yTGniJ24_0(.din(n4892), .dout(n4895));
    jdff dff_A_Oo8xOv4Z2_0(.din(n4889), .dout(n4892));
    jdff dff_A_lQQ7OrNU9_0(.din(n4886), .dout(n4889));
    jdff dff_A_Jo05WalF4_0(.din(n4883), .dout(n4886));
    jdff dff_A_tgsGGwUG3_2(.din(n440), .dout(n4883));
    jdff dff_A_etucNoNa4_0(.din(G134), .dout(n4880));
    jdff dff_A_AwtVxnWA7_0(.din(n4880), .dout(n4877));
    jdff dff_A_Pr4o3CpU3_0(.din(n4877), .dout(n4874));
    jdff dff_A_j27VBrhb1_0(.din(n4874), .dout(n4871));
    jdff dff_A_1bPf2LbR7_0(.din(n4871), .dout(n4868));
    jdff dff_A_Ji5K9ZSn0_0(.din(n4868), .dout(n4865));
    jdff dff_A_sSivf5sT5_0(.din(n4865), .dout(n4862));
    jdff dff_A_4qiJJOE21_0(.din(n4862), .dout(n4859));
    jdff dff_A_CrhC5AA46_0(.din(n4859), .dout(n4856));
    jdff dff_A_b5eJjfJ28_0(.din(n4856), .dout(n4853));
    jdff dff_A_BmZUYzin4_0(.din(n4853), .dout(n4850));
    jdff dff_A_Hk3nXfqo8_0(.din(n4850), .dout(n4847));
    jdff dff_B_TYwom6MH1_3(.din(G137), .dout(n4845));
    jdff dff_A_0jUAIR0N0_2(.din(n4845), .dout(n4841));
    jdff dff_A_gwoGQgPo3_2(.din(n4841), .dout(n4838));
    jdff dff_A_kaFOH6IU9_0(.din(n4845), .dout(n4835));
    jdff dff_A_VkgiVfXZ7_0(.din(n4835), .dout(n4832));
    jdff dff_A_WZ3AznBH3_0(.din(n4832), .dout(n4829));
    jdff dff_A_9nhakWyN2_0(.din(n4829), .dout(n4826));
    jdff dff_A_hvHGuKJ83_0(.din(n4826), .dout(n4823));
    jdff dff_A_A7GFZBeo0_0(.din(n4823), .dout(n4820));
    jdff dff_A_rEzsa2tP4_0(.din(n4820), .dout(n4817));
    jdff dff_A_p1WLYOiw3_0(.din(n4817), .dout(n4814));
    jdff dff_A_6wgcFCk43_0(.din(n4814), .dout(n4811));
    jdff dff_A_GtPlbU3g8_0(.din(n4811), .dout(n4808));
    jdff dff_A_TKgBSNOc3_0(.din(n4808), .dout(n4805));
    jdff dff_A_3crr4E687_0(.din(G131), .dout(n4802));
    jdff dff_A_hApYUv2t3_0(.din(n4802), .dout(n4799));
    jdff dff_A_UsCn5THH1_0(.din(n4799), .dout(n4796));
    jdff dff_A_1MXo40gh8_0(.din(n4796), .dout(n4793));
    jdff dff_A_9EuIiA1r1_0(.din(n4793), .dout(n4790));
    jdff dff_A_VxZaGK1w3_0(.din(n4790), .dout(n4787));
    jdff dff_A_oQ8MpKlk1_0(.din(n4787), .dout(n4784));
    jdff dff_A_MatWtpgi3_0(.din(n4784), .dout(n4781));
    jdff dff_A_OiKv6x1P3_0(.din(n4781), .dout(n4778));
    jdff dff_A_HiXB6ErV1_0(.din(n4778), .dout(n4775));
    jdff dff_A_zXIWKv336_0(.din(n4775), .dout(n4772));
    jdff dff_A_mQkGIWB23_0(.din(n4772), .dout(n4769));
    jdff dff_A_wOV34ZYg8_1(.din(n131), .dout(n4766));
    jdff dff_A_TOF1ISug0_1(.din(G128), .dout(n4763));
    jdff dff_A_j6eTlFGV7_1(.din(n4763), .dout(n4760));
    jdff dff_A_AaxeuSG62_1(.din(n4760), .dout(n4757));
    jdff dff_A_f9Epro6U8_1(.din(n4757), .dout(n4754));
    jdff dff_A_ZbpgyP838_1(.din(n4754), .dout(n4751));
    jdff dff_A_HJTlownT6_1(.din(n4751), .dout(n4748));
    jdff dff_A_pasSz2kO4_1(.din(n4748), .dout(n4745));
    jdff dff_A_ML9fB5ek4_1(.din(n4745), .dout(n4742));
    jdff dff_A_4a5ZjSeF2_1(.din(n4742), .dout(n4739));
    jdff dff_A_bAvRgBrY7_1(.din(n4739), .dout(n4736));
    jdff dff_A_SKEkCR5y1_1(.din(n4736), .dout(n4733));
    jdff dff_A_8dGNuAjS6_1(.din(n4733), .dout(n4730));
    jdff dff_A_uPQtcYLi3_0(.din(G128), .dout(n4727));
    jdff dff_A_tAIPdC814_2(.din(G143), .dout(n4724));
    jdff dff_A_KvChh7Xe5_1(.din(G143), .dout(n4721));
    jdff dff_A_PtVCZn1s7_1(.din(n4721), .dout(n4718));
    jdff dff_A_iOJCDytV9_1(.din(n4718), .dout(n4715));
    jdff dff_A_RiPSRki43_1(.din(n4715), .dout(n4712));
    jdff dff_A_0FBt5On70_1(.din(n4712), .dout(n4709));
    jdff dff_A_gjJLpUjO2_1(.din(n4709), .dout(n4706));
    jdff dff_A_xjC3xC1f3_1(.din(n4706), .dout(n4703));
    jdff dff_A_qtqbA7TE2_1(.din(n4703), .dout(n4700));
    jdff dff_A_CZgREzlJ7_1(.din(n4700), .dout(n4697));
    jdff dff_A_4NJCaWES2_1(.din(n4697), .dout(n4694));
    jdff dff_A_V2GnYsRI4_1(.din(n4694), .dout(n4691));
    jdff dff_A_iwuOnkwX7_1(.din(n4691), .dout(n4688));
    jdff dff_A_Ooj9orFX9_0(.din(G146), .dout(n4685));
    jdff dff_A_nil8ntDj1_0(.din(n4685), .dout(n4682));
    jdff dff_A_C0Oae3SM7_0(.din(n4682), .dout(n4679));
    jdff dff_A_7pcJFWUh4_0(.din(n4679), .dout(n4676));
    jdff dff_A_ch50iC326_0(.din(n4676), .dout(n4673));
    jdff dff_A_bcKuHTcd4_0(.din(n4673), .dout(n4670));
    jdff dff_A_np2tc0dK7_0(.din(n4670), .dout(n4667));
    jdff dff_A_kP1S94qw3_0(.din(n4667), .dout(n4664));
    jdff dff_A_qyhQuvCh2_0(.din(n4664), .dout(n4661));
    jdff dff_A_3GdzA8GT8_0(.din(n4661), .dout(n4658));
    jdff dff_A_XUxXPWpj3_0(.din(n4658), .dout(n4655));
    jdff dff_A_QFbJyn4L1_0(.din(n4655), .dout(n4652));
    jdff dff_B_rrIwJGG22_1(.din(n128), .dout(n4650));
    jdff dff_A_uGUkLdGk8_0(.din(G113), .dout(n4646));
    jdff dff_A_wW6jRfOH3_0(.din(n4646), .dout(n4643));
    jdff dff_A_YZHVwf6Q8_0(.din(n4643), .dout(n4640));
    jdff dff_A_tNRargS47_0(.din(n4640), .dout(n4637));
    jdff dff_A_MGD9JNrL1_0(.din(n4637), .dout(n4634));
    jdff dff_A_ge88EaDK2_0(.din(n4634), .dout(n4631));
    jdff dff_A_Z7vQxSIJ0_0(.din(n4631), .dout(n4628));
    jdff dff_B_LWkzKn8m7_0(.din(n887), .dout(n2097));
    jdff dff_B_Be0JuueW8_0(.din(n2097), .dout(n2100));
    jdff dff_B_feKD8TAg8_0(.din(n2100), .dout(n2103));
    jdff dff_B_lkPmwJSH6_0(.din(n2103), .dout(n2106));
    jdff dff_B_Dus5asfn5_0(.din(n2106), .dout(n2109));
    jdff dff_B_Mh6gqh832_0(.din(n867), .dout(n2112));
    jdff dff_B_Iqg5cNID3_0(.din(n2112), .dout(n2115));
    jdff dff_B_WhPzckqG5_0(.din(n2115), .dout(n2118));
    jdff dff_B_Y1HlTLS96_1(.din(n859), .dout(n2121));
    jdff dff_B_k74NkQxL3_1(.din(n2121), .dout(n2124));
    jdff dff_B_3oUgQuJh8_0(.din(n851), .dout(n2127));
    jdff dff_B_cnGFPP2K6_0(.din(n2127), .dout(n2130));
    jdff dff_A_3ue1GCAa6_1(.din(n2139), .dout(n2132));
    jdff dff_B_pbGQtWSj8_2(.din(n815), .dout(n2136));
    jdff dff_B_fXGOIhMh3_2(.din(n2136), .dout(n2139));
    jdff dff_B_1z3qikvk4_0(.din(n803), .dout(n2142));
    jdff dff_B_OjrxPkoz1_0(.din(n799), .dout(n2145));
    jdff dff_B_0NusGIpQ1_1(.din(n1155), .dout(n2148));
    jdff dff_B_hdCoarWM4_1(.din(n894), .dout(n2151));
    jdff dff_B_DsJPWdlA2_1(.din(n2151), .dout(n2154));
    jdff dff_B_u0O1DsPH2_1(.din(n2154), .dout(n2157));
    jdff dff_B_JakKkpps1_1(.din(n2157), .dout(n2160));
    jdff dff_B_E6lrRoBW0_1(.din(n2160), .dout(n2163));
    jdff dff_B_VuZcRjQM4_1(.din(n2163), .dout(n2166));
    jdff dff_B_q5HVwXmD5_1(.din(n2166), .dout(n2169));
    jdff dff_B_13uuITfG2_1(.din(n2169), .dout(n2172));
    jdff dff_B_QL5mamIM6_1(.din(n2172), .dout(n2175));
    jdff dff_B_LnVkTcjl3_1(.din(n2175), .dout(n2178));
    jdff dff_B_8v4Z0UIu6_1(.din(n2178), .dout(n2181));
    jdff dff_B_7u0DeLhZ9_0(.din(n1147), .dout(n2184));
    jdff dff_B_lYykZK1E7_0(.din(n2184), .dout(n2187));
    jdff dff_B_fKrfXaD88_0(.din(n2187), .dout(n2190));
    jdff dff_B_wKbd32w60_0(.din(n2190), .dout(n2193));
    jdff dff_B_FuQIJ1E44_0(.din(n2193), .dout(n2196));
    jdff dff_B_H9cCylnh8_0(.din(n2196), .dout(n2199));
    jdff dff_B_uuXwp87y5_0(.din(n2199), .dout(n2202));
    jdff dff_B_WQ0cvmw84_0(.din(n2202), .dout(n2205));
    jdff dff_B_i2Ue4JlN0_0(.din(n2205), .dout(n2208));
    jdff dff_B_OXR17nlL7_0(.din(n2208), .dout(n2211));
    jdff dff_B_thlH4yks4_0(.din(n2211), .dout(n2214));
    jdff dff_B_mimsbmED9_0(.din(n2214), .dout(n2217));
    jdff dff_B_DzktRynN5_0(.din(n2217), .dout(n2220));
    jdff dff_B_dr0BwsTl6_0(.din(n2220), .dout(n2223));
    jdff dff_A_PWhc653A2_0(.din(n2228), .dout(n2225));
    jdff dff_A_T55N1r1Y9_0(.din(n2231), .dout(n2228));
    jdff dff_A_KFFnJt7d9_0(.din(n2234), .dout(n2231));
    jdff dff_A_s8VJWkIA8_0(.din(n2237), .dout(n2234));
    jdff dff_A_GwVN9RiE3_0(.din(n2240), .dout(n2237));
    jdff dff_A_jRpf3phO1_0(.din(n2243), .dout(n2240));
    jdff dff_A_E9kIB8ML0_0(.din(n2246), .dout(n2243));
    jdff dff_A_6So5Xe162_0(.din(n2249), .dout(n2246));
    jdff dff_A_vj5pcntQ1_0(.din(n2252), .dout(n2249));
    jdff dff_A_58eoaMGF4_0(.din(n2255), .dout(n2252));
    jdff dff_A_z9WPkE0c8_0(.din(n2258), .dout(n2255));
    jdff dff_A_Tns3PYmN2_0(.din(n2261), .dout(n2258));
    jdff dff_A_Xs4reAsg9_0(.din(n2264), .dout(n2261));
    jdff dff_A_yE2KYfAC7_0(.din(n2267), .dout(n2264));
    jdff dff_A_wK8xo0ih4_0(.din(n1144), .dout(n2267));
    jdff dff_B_ANQgRK140_1(.din(n1193), .dout(n2271));
    jdff dff_B_4EnfuEyv7_1(.din(n1178), .dout(n2274));
    jdff dff_B_Oro06xku4_1(.din(n2274), .dout(n2277));
    jdff dff_B_XzmnYfwm7_1(.din(n2277), .dout(n2280));
    jdff dff_B_o5wRrX1u5_1(.din(n2280), .dout(n2283));
    jdff dff_B_DOqRJtRL1_1(.din(n2283), .dout(n2286));
    jdff dff_B_RB58VdCH1_1(.din(n2286), .dout(n2289));
    jdff dff_B_CRDkqrFk2_1(.din(n2289), .dout(n2292));
    jdff dff_B_8GAmCsxX6_1(.din(n2292), .dout(n2295));
    jdff dff_B_Rd0PAMwQ7_1(.din(n2295), .dout(n2298));
    jdff dff_B_jV8dr14K4_1(.din(n2298), .dout(n2301));
    jdff dff_B_fuB4YbjP6_1(.din(n2301), .dout(n2304));
    jdff dff_B_74JaBsIo5_0(.din(n1185), .dout(n2307));
    jdff dff_B_euM955On1_0(.din(n2307), .dout(n2310));
    jdff dff_B_cQbWAykn8_0(.din(n2310), .dout(n2313));
    jdff dff_B_luXDGkTp1_0(.din(n2313), .dout(n2316));
    jdff dff_B_05lhf9A88_0(.din(n2316), .dout(n2319));
    jdff dff_B_sZFyscMk1_0(.din(n2319), .dout(n2322));
    jdff dff_B_1vOjhKA85_0(.din(n2322), .dout(n2325));
    jdff dff_B_E0OyvjAW3_0(.din(n2325), .dout(n2328));
    jdff dff_B_hPzftarw4_0(.din(n2328), .dout(n2331));
    jdff dff_B_9TK02zqz0_0(.din(n2331), .dout(n2334));
    jdff dff_B_zCSJrkjM3_0(.din(n2334), .dout(n2337));
    jdff dff_B_0eEjCKXP5_0(.din(n2337), .dout(n2340));
    jdff dff_B_b6LaWH4c2_0(.din(n2340), .dout(n2343));
    jdff dff_B_Hz6UxcGC4_0(.din(n2343), .dout(n2346));
    jdff dff_A_WHafdpbG5_0(.din(n2351), .dout(n2348));
    jdff dff_A_M81hBMB46_0(.din(n2354), .dout(n2351));
    jdff dff_A_mFIrA8nf3_0(.din(n2357), .dout(n2354));
    jdff dff_A_SKUTIPTp3_0(.din(n2360), .dout(n2357));
    jdff dff_A_ZUbskobr6_0(.din(n2363), .dout(n2360));
    jdff dff_A_FIT1i4QH2_0(.din(n2366), .dout(n2363));
    jdff dff_A_xWOzoEwx6_0(.din(n2369), .dout(n2366));
    jdff dff_A_SVMe4flY6_0(.din(n2372), .dout(n2369));
    jdff dff_A_J79ltrwf6_0(.din(n2375), .dout(n2372));
    jdff dff_A_mCJiZiea9_0(.din(n2378), .dout(n2375));
    jdff dff_A_2w90mkWU1_0(.din(n2381), .dout(n2378));
    jdff dff_A_4SjneQ7j3_0(.din(n2384), .dout(n2381));
    jdff dff_A_3VrIdUWG7_0(.din(n2387), .dout(n2384));
    jdff dff_A_TKIxaGy19_0(.din(n2390), .dout(n2387));
    jdff dff_A_8J7Opxhj7_0(.din(n1182), .dout(n2390));
    jdff dff_B_SQh2gQdA3_1(.din(n1227), .dout(n2394));
    jdff dff_B_BJ6Rooop7_1(.din(n1212), .dout(n2397));
    jdff dff_B_748Igfu64_1(.din(n2397), .dout(n2400));
    jdff dff_B_DcC6rqkx2_1(.din(n2400), .dout(n2403));
    jdff dff_B_JVUOG1LR0_1(.din(n2403), .dout(n2406));
    jdff dff_B_xKDCvSCA8_1(.din(n2406), .dout(n2409));
    jdff dff_B_6kyTUGvp2_1(.din(n2409), .dout(n2412));
    jdff dff_B_OAGK93mI9_1(.din(n2412), .dout(n2415));
    jdff dff_B_hypuAYjm0_1(.din(n2415), .dout(n2418));
    jdff dff_B_6pDOdZjL4_1(.din(n2418), .dout(n2421));
    jdff dff_B_7hEdY94K4_1(.din(n2421), .dout(n2424));
    jdff dff_B_Slxm1lx63_1(.din(n2424), .dout(n2427));
    jdff dff_B_BBvIKtNP1_0(.din(n1219), .dout(n2430));
    jdff dff_B_xciTNEE36_0(.din(n2430), .dout(n2433));
    jdff dff_B_Ro86NhZw8_0(.din(n2433), .dout(n2436));
    jdff dff_B_jwgBJArJ6_0(.din(n2436), .dout(n2439));
    jdff dff_B_jGNFm7hT8_0(.din(n2439), .dout(n2442));
    jdff dff_B_dd85IcJm3_0(.din(n2442), .dout(n2445));
    jdff dff_B_udz6a51B2_0(.din(n2445), .dout(n2448));
    jdff dff_B_8R9AMw6g2_0(.din(n2448), .dout(n2451));
    jdff dff_B_BuFks82O4_0(.din(n2451), .dout(n2454));
    jdff dff_B_Imz9GHSJ2_0(.din(n2454), .dout(n2457));
    jdff dff_B_xxDbMDP82_0(.din(n2457), .dout(n2460));
    jdff dff_B_D7WhIya89_0(.din(n2460), .dout(n2463));
    jdff dff_B_zyeN6HZ17_0(.din(n2463), .dout(n2466));
    jdff dff_B_uPAk3PsE8_0(.din(n2466), .dout(n2469));
    jdff dff_A_dXEIWgDr5_0(.din(n2474), .dout(n2471));
    jdff dff_A_UblRcr5H7_0(.din(n2477), .dout(n2474));
    jdff dff_A_GbX3sqRV6_0(.din(n2480), .dout(n2477));
    jdff dff_A_jNwtQAJy2_0(.din(n2483), .dout(n2480));
    jdff dff_A_SBVTTQf23_0(.din(n2486), .dout(n2483));
    jdff dff_A_txZ7Byz38_0(.din(n2489), .dout(n2486));
    jdff dff_A_8uVVB5dg1_0(.din(n2492), .dout(n2489));
    jdff dff_A_3CkFEYoY8_0(.din(n2495), .dout(n2492));
    jdff dff_A_EYRVDabA5_0(.din(n2498), .dout(n2495));
    jdff dff_A_PsEwy2V65_0(.din(n2501), .dout(n2498));
    jdff dff_A_3G1Q4sZu6_0(.din(n2504), .dout(n2501));
    jdff dff_A_fZa86WO57_0(.din(n2507), .dout(n2504));
    jdff dff_A_DBUrhVvv0_0(.din(n2510), .dout(n2507));
    jdff dff_A_amj7g5Eo1_0(.din(n2513), .dout(n2510));
    jdff dff_A_TB6WP7ZL0_0(.din(n1216), .dout(n2513));
    jdff dff_B_kP0FXXRz4_1(.din(n1261), .dout(n2517));
    jdff dff_B_v6jcs1Tw1_1(.din(n1246), .dout(n2520));
    jdff dff_B_7SdlZiU25_1(.din(n2520), .dout(n2523));
    jdff dff_B_IcRwO1FJ6_1(.din(n2523), .dout(n2526));
    jdff dff_B_gQBk2m2P4_1(.din(n2526), .dout(n2529));
    jdff dff_B_iVlEzbxa0_1(.din(n2529), .dout(n2532));
    jdff dff_B_p0rppZQ87_1(.din(n2532), .dout(n2535));
    jdff dff_B_2nxCeAFo6_1(.din(n2535), .dout(n2538));
    jdff dff_B_bzqeEy5W3_1(.din(n2538), .dout(n2541));
    jdff dff_B_ic9vLmhp3_1(.din(n2541), .dout(n2544));
    jdff dff_B_233cQcXb5_1(.din(n2544), .dout(n2547));
    jdff dff_B_LUDNu2k16_1(.din(n2547), .dout(n2550));
    jdff dff_B_3laqQ3w85_0(.din(n1253), .dout(n2553));
    jdff dff_B_MRvqB5mu9_0(.din(n2553), .dout(n2556));
    jdff dff_B_SzAMrhsn1_0(.din(n2556), .dout(n2559));
    jdff dff_B_tsYHOX1q3_0(.din(n2559), .dout(n2562));
    jdff dff_B_u7wycnjS7_0(.din(n2562), .dout(n2565));
    jdff dff_B_rwp3hnEd4_0(.din(n2565), .dout(n2568));
    jdff dff_B_GKklkikf7_0(.din(n2568), .dout(n2571));
    jdff dff_B_V3T70aNx7_0(.din(n2571), .dout(n2574));
    jdff dff_B_Ujlr2ZEg2_0(.din(n2574), .dout(n2577));
    jdff dff_B_fzpbSU6a7_0(.din(n2577), .dout(n2580));
    jdff dff_B_rK25yWXp3_0(.din(n2580), .dout(n2583));
    jdff dff_B_wBy5jWGb1_0(.din(n2583), .dout(n2586));
    jdff dff_B_VmD68pLY4_0(.din(n2586), .dout(n2589));
    jdff dff_B_0pIk17TD5_0(.din(n2589), .dout(n2592));
    jdff dff_A_hJW82m2V4_0(.din(n2597), .dout(n2594));
    jdff dff_A_qcHMD30S9_0(.din(n2600), .dout(n2597));
    jdff dff_A_N7O9EOkX8_0(.din(n2603), .dout(n2600));
    jdff dff_A_j6zj1VIC0_0(.din(n2606), .dout(n2603));
    jdff dff_A_nhDcfOLW9_0(.din(n2609), .dout(n2606));
    jdff dff_A_Ckdu4Zry7_0(.din(n2612), .dout(n2609));
    jdff dff_A_PLKzdo2s9_0(.din(n2615), .dout(n2612));
    jdff dff_A_25FElTfP6_0(.din(n2618), .dout(n2615));
    jdff dff_A_tnZHCPXS6_0(.din(n2621), .dout(n2618));
    jdff dff_A_9I41b1se1_0(.din(n2624), .dout(n2621));
    jdff dff_A_4Ete7m1f1_0(.din(n2627), .dout(n2624));
    jdff dff_A_528SSXMD5_0(.din(n2630), .dout(n2627));
    jdff dff_A_2rWGtBLo2_0(.din(n2633), .dout(n2630));
    jdff dff_A_5o1TCmD08_0(.din(n2636), .dout(n2633));
    jdff dff_A_CcABDC6X3_0(.din(n1250), .dout(n2636));
    jdff dff_B_hhH2xC3T0_1(.din(n1289), .dout(n2640));
    jdff dff_B_c0dvw7ia2_0(.din(n1292), .dout(n2643));
    jdff dff_B_DoWwuulz7_0(.din(n2643), .dout(n2646));
    jdff dff_B_8o2Hng001_0(.din(n2646), .dout(n2649));
    jdff dff_B_zfNmRqNX3_0(.din(n2649), .dout(n2652));
    jdff dff_B_boihjMx19_0(.din(n2652), .dout(n2655));
    jdff dff_B_c1jH6Jpe8_0(.din(n2655), .dout(n2658));
    jdff dff_B_nhcB0gVo4_0(.din(n2658), .dout(n2661));
    jdff dff_B_8taZhUz01_0(.din(n2661), .dout(n2664));
    jdff dff_B_PoYWSBeP3_0(.din(n2664), .dout(n2667));
    jdff dff_B_rpsa5okZ2_0(.din(n2667), .dout(n2670));
    jdff dff_B_v1dQ2yPZ9_0(.din(n2670), .dout(n2673));
    jdff dff_B_NEupvcRc5_0(.din(n2673), .dout(n2676));
    jdff dff_B_LsTfgIb25_0(.din(n2676), .dout(n2679));
    jdff dff_B_6ZN0m6354_0(.din(n2679), .dout(n2682));
    jdff dff_A_mBkQ8FAy0_1(.din(n2687), .dout(n2684));
    jdff dff_A_YN62kmNa5_1(.din(n2690), .dout(n2687));
    jdff dff_A_aNi0VYs67_1(.din(n2693), .dout(n2690));
    jdff dff_A_f5GXX9C38_1(.din(n2696), .dout(n2693));
    jdff dff_A_DD2Q51WV7_1(.din(n2699), .dout(n2696));
    jdff dff_A_76QmUyYJ1_1(.din(n2702), .dout(n2699));
    jdff dff_A_hXQ8m05g6_1(.din(n2705), .dout(n2702));
    jdff dff_A_zYPqyOQZ3_1(.din(n2708), .dout(n2705));
    jdff dff_A_iKRB8Wsv9_1(.din(n2711), .dout(n2708));
    jdff dff_A_MT0lSSNP4_1(.din(n2714), .dout(n2711));
    jdff dff_A_MfaGeG4A4_1(.din(n2717), .dout(n2714));
    jdff dff_A_s8bj5XiD9_1(.din(n2720), .dout(n2717));
    jdff dff_A_7sHtpric0_1(.din(n2723), .dout(n2720));
    jdff dff_A_XhwenyFf1_1(.din(n2726), .dout(n2723));
    jdff dff_A_6mnfjbqs5_1(.din(n1281), .dout(n2726));
    jdff dff_B_6Mcs3N3a4_1(.din(n1311), .dout(n2730));
    jdff dff_B_IquWU2O29_1(.din(n2730), .dout(n2733));
    jdff dff_B_TyHydjQp0_1(.din(n2733), .dout(n2736));
    jdff dff_B_mD54nwjh4_1(.din(n2736), .dout(n2739));
    jdff dff_B_z8h3506y6_1(.din(n2739), .dout(n2742));
    jdff dff_B_2GaigCDV5_1(.din(n2742), .dout(n2745));
    jdff dff_B_lQkRj6Iz3_1(.din(n2745), .dout(n2748));
    jdff dff_B_LudLZ19a0_1(.din(n2748), .dout(n2751));
    jdff dff_B_VsWPvjX49_1(.din(n2751), .dout(n2754));
    jdff dff_B_qbYWJHA10_1(.din(n2754), .dout(n2757));
    jdff dff_B_O9sw4Yu05_1(.din(n2757), .dout(n2760));
    jdff dff_B_sSDWAtkI3_1(.din(n2760), .dout(n2763));
    jdff dff_B_Le9lD93B3_1(.din(n2763), .dout(n2766));
    jdff dff_B_GnHCDVG52_1(.din(n2766), .dout(n2769));
    jdff dff_B_PUcHH9zB0_1(.din(n2769), .dout(n2772));
    jdff dff_B_H800PHkW1_0(.din(n1319), .dout(n2775));
    jdff dff_B_XO80HZbQ7_0(.din(n2775), .dout(n2778));
    jdff dff_B_HyClYrg89_0(.din(n2778), .dout(n2781));
    jdff dff_B_PkibqWmq9_0(.din(n2781), .dout(n2784));
    jdff dff_B_Hqj4vDCg5_0(.din(n2784), .dout(n2787));
    jdff dff_B_Hgqy3dFk0_0(.din(n2787), .dout(n2790));
    jdff dff_B_v8gxKJNi0_0(.din(n2790), .dout(n2793));
    jdff dff_B_1tux3dAl5_0(.din(n2793), .dout(n2796));
    jdff dff_B_z6c6gTAI4_0(.din(n2796), .dout(n2799));
    jdff dff_B_9P16P36S9_0(.din(n2799), .dout(n2802));
    jdff dff_B_kzZdAeqh0_0(.din(n2802), .dout(n2805));
    jdff dff_B_nEajhgS89_0(.din(n2805), .dout(n2808));
    jdff dff_B_vUCbUvtk0_0(.din(n2808), .dout(n2811));
    jdff dff_B_vItphulR1_0(.din(n2811), .dout(n2814));
    jdff dff_B_HCeY6Xsg9_0(.din(n1358), .dout(n2817));
    jdff dff_B_wMfhvqXj8_0(.din(n2817), .dout(n2820));
    jdff dff_B_V7RppE9K3_0(.din(n2820), .dout(n2823));
    jdff dff_B_hNunlZQT5_0(.din(n2823), .dout(n2826));
    jdff dff_B_FabcnBuR2_0(.din(n2826), .dout(n2829));
    jdff dff_B_EEEa5WqG6_0(.din(n2829), .dout(n2832));
    jdff dff_B_CBw6WWyj2_0(.din(n2832), .dout(n2835));
    jdff dff_B_vE20W2EV6_0(.din(n2835), .dout(n2838));
    jdff dff_B_wJ4gMpo62_0(.din(n2838), .dout(n2841));
    jdff dff_B_21naDq6z9_0(.din(n2841), .dout(n2844));
    jdff dff_B_03H9PegJ1_0(.din(n2844), .dout(n2847));
    jdff dff_B_utAAeGFS6_1(.din(n1350), .dout(n2850));
    jdff dff_B_vd9YvGa17_1(.din(n2850), .dout(n2853));
    jdff dff_B_ooi95S6u9_0(.din(n1343), .dout(n2856));
    jdff dff_B_i5PDVMKi8_0(.din(n2856), .dout(n2859));
    jdff dff_B_FMRsiVLd6_0(.din(n2859), .dout(n2862));
    jdff dff_B_6EiM8kwb2_0(.din(n2862), .dout(n2865));
    jdff dff_B_cyxcypYz0_0(.din(n2865), .dout(n2868));
    jdff dff_B_N3mjGSh68_0(.din(n2868), .dout(n2871));
    jdff dff_B_CTe91qRz2_0(.din(n2871), .dout(n2874));
    jdff dff_B_IgAnoSEi5_0(.din(n2874), .dout(n2877));
    jdff dff_B_w8VI9R5M8_0(.din(n2877), .dout(n2880));
    jdff dff_B_fdQnRn6U8_0(.din(n2880), .dout(n2883));
    jdff dff_B_KCOZqQJA1_0(.din(n2883), .dout(n2886));
    jdff dff_B_6twX056v2_0(.din(n2886), .dout(n2889));
    jdff dff_B_oKxb8BLI3_0(.din(n2889), .dout(n2892));
    jdff dff_B_bNBiZI2c2_1(.din(n1380), .dout(n2895));
    jdff dff_B_0kZ2z18R8_0(.din(n703), .dout(n2898));
    jdff dff_A_A0xHajm72_0(.din(n2903), .dout(n2900));
    jdff dff_A_2Qa4mDst8_0(.din(n679), .dout(n2903));
    jdff dff_A_qkEZTYbq6_2(.din(n2909), .dout(n2906));
    jdff dff_A_Q9G6vVgF3_2(.din(n679), .dout(n2909));
    jdff dff_A_jsAhbsnF8_0(.din(n2919), .dout(n2912));
    jdff dff_A_AqRVZuO56_2(.din(n2919), .dout(n2915));
    jdff dff_B_xAj10c8M8_3(.din(n577), .dout(n2919));
    jdff dff_B_VWqHtd9m4_0(.din(n644), .dout(n2922));
    jdff dff_A_l0EIxeY21_0(.din(n600), .dout(n2924));
    jdff dff_A_KXlByAQf7_2(.din(n2930), .dout(n2927));
    jdff dff_A_jQgXWgqB0_2(.din(n600), .dout(n2930));
    jdff dff_A_2MC35eKk5_0(.din(n2936), .dout(n2933));
    jdff dff_A_bIOKmwFE6_0(.din(n596), .dout(n2936));
    jdff dff_A_7hU9kEf18_1(.din(n2942), .dout(n2939));
    jdff dff_A_HHgnVmET5_1(.din(n596), .dout(n2942));
    jdff dff_A_L8M4JS3W9_0(.din(n2952), .dout(n2945));
    jdff dff_A_e0hOEbT09_2(.din(n2952), .dout(n2948));
    jdff dff_B_XXYDJJC69_3(.din(n432), .dout(n2952));
    jdff dff_A_uOwPDkx45_0(.din(n2957), .dout(n2954));
    jdff dff_A_ALtmhgTc6_0(.din(n391), .dout(n2957));
    jdff dff_A_8RuVw5tC8_1(.din(n2963), .dout(n2960));
    jdff dff_A_EGYRcwBO5_1(.din(n391), .dout(n2963));
    jdff dff_A_9SSMtdeU1_2(.din(n2969), .dout(n2966));
    jdff dff_A_gtbJ1B1o4_2(.din(n447), .dout(n2969));
    jdff dff_A_fOwRUP1N3_2(.din(n2976), .dout(n2972));
    jdff dff_B_W1OUvgBT0_3(.din(n302), .dout(n2976));
    jdff dff_A_Shzbzd048_1(.din(n2981), .dout(n2978));
    jdff dff_A_W6SoiKOo9_1(.din(n2984), .dout(n2981));
    jdff dff_A_VFOZdRBQ2_1(.din(n2987), .dout(n2984));
    jdff dff_A_FvrCfnJD3_1(.din(n204), .dout(n2987));
    jdff dff_A_I348fSb59_2(.din(n2993), .dout(n2990));
    jdff dff_A_Mogc7lRq2_2(.din(n2996), .dout(n2993));
    jdff dff_A_y4d6FUuI4_2(.din(n2999), .dout(n2996));
    jdff dff_A_hDLlR9aU9_2(.din(n204), .dout(n2999));
    jdff dff_B_fmX5IGTT2_3(.din(n1159), .dout(n3003));
    jdff dff_B_VihuQQtv3_3(.din(n3003), .dout(n3006));
    jdff dff_B_iqoVMd6k3_3(.din(n3006), .dout(n3009));
    jdff dff_B_ylKjk9M09_3(.din(n3009), .dout(n3012));
    jdff dff_B_ugbwOPxA9_3(.din(n3012), .dout(n3015));
    jdff dff_B_91GUwpgB9_3(.din(n3015), .dout(n3018));
    jdff dff_B_PtF5RnJI4_3(.din(n3018), .dout(n3021));
    jdff dff_B_ews6HzcO6_3(.din(n3021), .dout(n3024));
    jdff dff_B_x22F5vcs9_3(.din(n3024), .dout(n3027));
    jdff dff_B_OwRWhq653_3(.din(n3027), .dout(n3030));
    jdff dff_B_iRIJRMt13_3(.din(n3030), .dout(n3033));
    jdff dff_B_8eHgVTOX8_3(.din(n3033), .dout(n3036));
    jdff dff_B_aqMOPiYk9_3(.din(n3036), .dout(n3039));
    jdff dff_B_AiVg1xue0_3(.din(n3039), .dout(n3042));
    jdff dff_B_LKvHw9nw2_3(.din(n3042), .dout(n3045));
    jdff dff_B_XEK9xg8v1_3(.din(n3045), .dout(n3048));
    jdff dff_B_qrCXNbTi1_1(.din(n1365), .dout(n3051));
    jdff dff_B_kmet4QdL0_1(.din(n3051), .dout(n3054));
    jdff dff_B_UIP3Bl9K0_1(.din(n3054), .dout(n3057));
    jdff dff_B_fC369nER5_1(.din(n3057), .dout(n3060));
    jdff dff_B_fFhIUMYH7_1(.din(n3060), .dout(n3063));
    jdff dff_B_MSky3R4C5_1(.din(n3063), .dout(n3066));
    jdff dff_B_8etoQi9d5_1(.din(n3066), .dout(n3069));
    jdff dff_B_Z35LIqLt5_1(.din(n3069), .dout(n3072));
    jdff dff_B_CxMlmehe3_1(.din(n3072), .dout(n3075));
    jdff dff_B_rM6vO3xV6_1(.din(n3075), .dout(n3078));
    jdff dff_B_rg16n2yA1_1(.din(n3078), .dout(n3081));
    jdff dff_B_dn0deQQx3_0(.din(n1372), .dout(n3084));
    jdff dff_B_rHLRHm304_0(.din(n3084), .dout(n3087));
    jdff dff_B_dBUl07bo3_0(.din(n3087), .dout(n3090));
    jdff dff_B_nFgPMPZJ8_0(.din(n3090), .dout(n3093));
    jdff dff_B_e6POofZE0_0(.din(n3093), .dout(n3096));
    jdff dff_B_k9as2cgn9_0(.din(n3096), .dout(n3099));
    jdff dff_B_iJ1Sgwnx8_0(.din(n3099), .dout(n3102));
    jdff dff_B_MHYNxXFv3_0(.din(n3102), .dout(n3105));
    jdff dff_B_xh2IlJkJ3_0(.din(n3105), .dout(n3108));
    jdff dff_B_TpthdZRQ8_0(.din(n3108), .dout(n3111));
    jdff dff_B_ZItEWuXN2_0(.din(n3111), .dout(n3114));
    jdff dff_B_VNNNKHBf2_0(.din(n3114), .dout(n3117));
    jdff dff_B_YYTIRybh0_0(.din(n3117), .dout(n3120));
    jdff dff_B_dl0Rx4Pp3_0(.din(n3120), .dout(n3123));
    jdff dff_A_1fyWL2jF4_0(.din(n3128), .dout(n3125));
    jdff dff_A_73TrNSFc1_0(.din(n3131), .dout(n3128));
    jdff dff_A_hmd0lHZm7_0(.din(n3134), .dout(n3131));
    jdff dff_A_oxJmmROU8_0(.din(n3137), .dout(n3134));
    jdff dff_A_T0lDex9y5_0(.din(n3140), .dout(n3137));
    jdff dff_A_F0V9QpbM3_0(.din(n3143), .dout(n3140));
    jdff dff_A_UBbUylUN6_0(.din(n3146), .dout(n3143));
    jdff dff_A_PVzqeHDp0_0(.din(n3149), .dout(n3146));
    jdff dff_A_hGkt8E1k4_0(.din(n3152), .dout(n3149));
    jdff dff_A_mSLNJsGa4_0(.din(n3155), .dout(n3152));
    jdff dff_A_pMrlqy470_0(.din(n3158), .dout(n3155));
    jdff dff_A_m6Qx9DAJ2_0(.din(n3161), .dout(n3158));
    jdff dff_A_LhM1B9Pt1_0(.din(n3164), .dout(n3161));
    jdff dff_A_fd4PZKEL4_0(.din(n3167), .dout(n3164));
    jdff dff_A_U46uTslA6_0(.din(n1369), .dout(n3167));
    jdff dff_B_qRJjuky49_0(.din(n1116), .dout(n3171));
    jdff dff_B_P1oev6OL7_0(.din(n1092), .dout(n3174));
    jdff dff_A_O4s2vHtd0_1(.din(n3179), .dout(n3176));
    jdff dff_A_eRcrnQaJ8_1(.din(n565), .dout(n3179));
    jdff dff_B_0F73FT6u8_2(.din(n1073), .dout(n3183));
    jdff dff_A_CtB0uMGN2_1(.din(n3188), .dout(n3185));
    jdff dff_A_NtqSXtuH4_1(.din(n549), .dout(n3188));
    jdff dff_A_hBG93Yhh6_2(.din(n3194), .dout(n3191));
    jdff dff_A_7XvFw0v89_2(.din(n549), .dout(n3194));
    jdff dff_B_6TFqzJ3w3_3(.din(n545), .dout(n3198));
    jdff dff_B_IEPWR7JI3_3(.din(n3198), .dout(n3201));
    jdff dff_A_DjGGIK7h6_0(.din(n3210), .dout(n3203));
    jdff dff_A_FKtcFAdn1_1(.din(n3210), .dout(n3206));
    jdff dff_B_IwweuLLc4_3(.din(n1058), .dout(n3210));
    jdff dff_A_n1nyfuVj7_1(.din(n3219), .dout(n3212));
    jdff dff_A_OZ8KK12W0_2(.din(n3219), .dout(n3215));
    jdff dff_B_xgSN3V3V7_3(.din(n1046), .dout(n3219));
    jdff dff_A_pbPmsnQ15_0(.din(n3224), .dout(n3221));
    jdff dff_A_aL9ZvaMz2_0(.din(n3227), .dout(n3224));
    jdff dff_A_EWqnEigz3_0(.din(n542), .dout(n3227));
    jdff dff_A_WrjgMOFJ0_1(.din(n3233), .dout(n3230));
    jdff dff_A_E73AQ5V10_1(.din(n3236), .dout(n3233));
    jdff dff_A_CpOdx5Gu0_1(.din(n542), .dout(n3236));
    jdff dff_B_wOFWd6LP3_0(.din(n538), .dout(n3240));
    jdff dff_B_GAw23NGM7_1(.din(G900), .dout(n3243));
    jdff dff_B_nCvU86gK5_0(.din(n1018), .dout(n3246));
    jdff dff_A_REGWZ8k48_1(.din(n561), .dout(n3248));
    jdff dff_A_n2Tcoh2U6_0(.din(n3255), .dout(n3251));
    jdff dff_B_vBdGNBbj5_3(.din(n963), .dout(n3255));
    jdff dff_A_VrzoVLr50_0(.din(n3260), .dout(n3257));
    jdff dff_A_lnNYhLRA3_0(.din(n959), .dout(n3260));
    jdff dff_B_sJq7yOVI7_3(.din(n443), .dout(n3264));
    jdff dff_A_IANGZgsD2_0(.din(n3269), .dout(n3266));
    jdff dff_A_OK5if8aX3_0(.din(n189), .dout(n3269));
    jdff dff_A_tmxZjWrt0_2(.din(n3275), .dout(n3272));
    jdff dff_A_XI8h2cgr0_2(.din(n189), .dout(n3275));
    jdff dff_B_E2Ozntam6_2(.din(n947), .dout(n3279));
    jdff dff_A_X1itAvbh4_1(.din(n3284), .dout(n3281));
    jdff dff_A_L4GXIG7G1_1(.din(n463), .dout(n3284));
    jdff dff_A_T3WBiKFQ5_2(.din(n3290), .dout(n3287));
    jdff dff_A_19nn0ZKO9_2(.din(n463), .dout(n3290));
    jdff dff_B_RlcOllUj0_1(.din(n309), .dout(n3294));
    jdff dff_B_BttTsZuX8_1(.din(n3294), .dout(n3297));
    jdff dff_B_2NvLaf0d2_1(.din(n3297), .dout(n3300));
    jdff dff_B_E6KpvIQS1_1(.din(n3300), .dout(n3303));
    jdff dff_B_tgqTKjST6_1(.din(n3303), .dout(n3306));
    jdff dff_A_3uMTGr290_0(.din(n3311), .dout(n3308));
    jdff dff_A_enOvBShm0_0(.din(n3314), .dout(n3311));
    jdff dff_A_ENUTJ48H9_0(.din(n3317), .dout(n3314));
    jdff dff_A_8LcSwH8V3_0(.din(n3320), .dout(n3317));
    jdff dff_A_1W7IgUaM5_0(.din(n3323), .dout(n3320));
    jdff dff_A_58imru5c5_0(.din(n3326), .dout(n3323));
    jdff dff_A_TsBU1uMv0_0(.din(n3329), .dout(n3326));
    jdff dff_A_sPGb23ld7_0(.din(n3332), .dout(n3329));
    jdff dff_A_k3v7wEYI1_0(.din(n3335), .dout(n3332));
    jdff dff_A_6AJDCdFE1_0(.din(n99), .dout(n3335));
    jdff dff_A_XLhE6Odj0_0(.din(n3345), .dout(n3338));
    jdff dff_A_sTQzwxcp3_1(.din(n3345), .dout(n3341));
    jdff dff_B_RiIbFyzW2_3(.din(n928), .dout(n3345));
    jdff dff_B_GQ5WKW4Z3_2(.din(n916), .dout(n3348));
    jdff dff_A_LPKtXx3w1_1(.din(n3353), .dout(n3350));
    jdff dff_A_375026EZ7_1(.din(n483), .dout(n3353));
    jdff dff_A_4M3NhlzX8_2(.din(n3359), .dout(n3356));
    jdff dff_A_MM0cDStJ0_2(.din(n483), .dout(n3359));
    jdff dff_B_RYP7aEv24_1(.din(n348), .dout(n3363));
    jdff dff_B_iB72dv0Z8_1(.din(n3363), .dout(n3366));
    jdff dff_B_al3r44FB2_1(.din(n3366), .dout(n3369));
    jdff dff_B_A7iquh0X4_1(.din(n3369), .dout(n3372));
    jdff dff_B_gkBWQhNm3_1(.din(n3372), .dout(n3375));
    jdff dff_A_gg5hEwhF8_0(.din(n3380), .dout(n3377));
    jdff dff_A_WenNg6Ky8_0(.din(n3383), .dout(n3380));
    jdff dff_A_MwJvXmnu9_0(.din(n3386), .dout(n3383));
    jdff dff_A_pDQ020eG4_0(.din(n3389), .dout(n3386));
    jdff dff_A_Q68tyZJT3_0(.din(n3392), .dout(n3389));
    jdff dff_A_LC3rQaQt4_0(.din(n3395), .dout(n3392));
    jdff dff_A_ZmC3SGWn1_0(.din(n3398), .dout(n3395));
    jdff dff_A_Ljyw1Tfj2_0(.din(n3401), .dout(n3398));
    jdff dff_A_0ya4Ojth2_0(.din(n3404), .dout(n3401));
    jdff dff_A_gRXzx6lV4_0(.din(n3407), .dout(n3404));
    jdff dff_A_ehwNMh3i9_0(.din(n3410), .dout(n3407));
    jdff dff_A_gV3TYRGf2_0(.din(n379), .dout(n3410));
    jdff dff_B_wGKmiluw8_1(.din(n352), .dout(n3414));
    jdff dff_B_32cs7bWc2_1(.din(n3414), .dout(n3417));
    jdff dff_A_iMghNJmt4_1(.din(n3422), .dout(n3419));
    jdff dff_A_r5EtnzcC9_1(.din(n3425), .dout(n3422));
    jdff dff_A_hAaYs4WB6_1(.din(n3428), .dout(n3425));
    jdff dff_A_Teu1UDtW7_1(.din(n3431), .dout(n3428));
    jdff dff_A_Yd45RafL0_1(.din(n3434), .dout(n3431));
    jdff dff_A_CEab87fn1_1(.din(G475), .dout(n3434));
    jdff dff_A_PEcKYvTo2_0(.din(n3440), .dout(n3437));
    jdff dff_A_09Ithtd01_0(.din(n3443), .dout(n3440));
    jdff dff_A_0AGzoZu19_0(.din(n3446), .dout(n3443));
    jdff dff_A_YDij4JRz9_0(.din(n3449), .dout(n3446));
    jdff dff_A_NYwfiaWO3_0(.din(n3452), .dout(n3449));
    jdff dff_A_XnX1efKo4_0(.din(n3455), .dout(n3452));
    jdff dff_A_PYpkFaEB2_0(.din(n3458), .dout(n3455));
    jdff dff_A_FIvoixvh8_0(.din(n3461), .dout(n3458));
    jdff dff_A_ULOqf1aM8_0(.din(n3464), .dout(n3461));
    jdff dff_A_HFst59VX1_0(.din(n3467), .dout(n3464));
    jdff dff_A_VSiWk4ZR0_0(.din(n3470), .dout(n3467));
    jdff dff_A_BIDb6lWi9_0(.din(n337), .dout(n3470));
    jdff dff_B_Po8Zbi7a6_1(.din(n313), .dout(n3474));
    jdff dff_B_Q3GIcbza0_1(.din(n3474), .dout(n3477));
    jdff dff_B_KYf5x2SV2_1(.din(n3477), .dout(n3480));
    jdff dff_B_vWcuUjsK6_0(.din(n329), .dout(n3483));
    jdff dff_A_uWZcgsMi2_1(.din(n3488), .dout(n3485));
    jdff dff_A_ScB36H0X3_1(.din(n3491), .dout(n3488));
    jdff dff_A_4c38AGAK5_1(.din(n3494), .dout(n3491));
    jdff dff_A_azIz4Y8S7_1(.din(n3497), .dout(n3494));
    jdff dff_A_xzz8La4D7_1(.din(n3500), .dout(n3497));
    jdff dff_A_WWtRK1vQ1_1(.din(G478), .dout(n3500));
    jdff dff_B_Ecqpcddf1_3(.din(n428), .dout(n3504));
    jdff dff_B_3tMQlBob3_3(.din(n3504), .dout(n3507));
    jdff dff_A_tw9iMYm32_0(.din(n3512), .dout(n3509));
    jdff dff_A_7f6FhRxn3_0(.din(n3515), .dout(n3512));
    jdff dff_A_qAr5oImy2_0(.din(n425), .dout(n3515));
    jdff dff_A_y39Ir1fy5_1(.din(n3521), .dout(n3518));
    jdff dff_A_ZNGFzyY63_1(.din(n3524), .dout(n3521));
    jdff dff_A_SAYeAZFS1_1(.din(n425), .dout(n3524));
    jdff dff_B_jF5kPCUT9_1(.din(n407), .dout(n3528));
    jdff dff_A_AizOC6QN4_0(.din(n418), .dout(n3530));
    jdff dff_A_IZaReYdH1_1(.din(n3536), .dout(n3533));
    jdff dff_A_GEijYecu8_1(.din(n3539), .dout(n3536));
    jdff dff_A_5Qhka2Bg4_1(.din(n3542), .dout(n3539));
    jdff dff_A_E7JR0M4V6_1(.din(n3545), .dout(n3542));
    jdff dff_A_wSuxgyHR1_1(.din(n3548), .dout(n3545));
    jdff dff_A_edH96Hus4_1(.din(n3551), .dout(n3548));
    jdff dff_A_A1IDbqi44_1(.din(n3554), .dout(n3551));
    jdff dff_A_SI7If7WT8_1(.din(n3557), .dout(n3554));
    jdff dff_A_m2SUxvgv9_1(.din(n3560), .dout(n3557));
    jdff dff_A_Wp07xHDd0_1(.din(n3563), .dout(n3560));
    jdff dff_A_CJMSy18s4_1(.din(n418), .dout(n3563));
    jdff dff_A_E0bkq6j93_1(.din(n3569), .dout(n3566));
    jdff dff_A_o6mUYrvZ4_1(.din(n3572), .dout(n3569));
    jdff dff_A_6XTcObx51_1(.din(n3575), .dout(n3572));
    jdff dff_A_nbxBiWfY8_1(.din(n3578), .dout(n3575));
    jdff dff_A_anU5sl0X7_1(.din(n3581), .dout(n3578));
    jdff dff_A_AlhORJZi8_1(.din(n3584), .dout(n3581));
    jdff dff_A_Ji7TlELM7_1(.din(n3587), .dout(n3584));
    jdff dff_A_zVcPylW94_1(.din(n3590), .dout(n3587));
    jdff dff_A_FY0A5AWO0_1(.din(n3593), .dout(n3590));
    jdff dff_A_oQtaNTI90_1(.din(n3596), .dout(n3593));
    jdff dff_A_7BQyAf1X2_1(.din(n3599), .dout(n3596));
    jdff dff_A_aCpNVqY13_1(.din(n3602), .dout(n3599));
    jdff dff_A_LqDRUReX2_1(.din(n3605), .dout(n3602));
    jdff dff_A_iI3HD5Bp2_1(.din(n3608), .dout(n3605));
    jdff dff_A_BYruvW6t9_1(.din(n3611), .dout(n3608));
    jdff dff_A_BsR5A8Rq5_1(.din(n3615), .dout(n3611));
    jdff dff_B_MxIFyWbc9_3(.din(G952), .dout(n3615));
    jdff dff_B_R6cGR84L7_1(.din(G898), .dout(n3618));
    jdff dff_A_VuuFiaHe4_2(.din(n819), .dout(n3620));
    jdff dff_A_4n5YnmTu4_1(.din(n3626), .dout(n3623));
    jdff dff_A_IIDNdxzU7_1(.din(n189), .dout(n3626));
    jdff dff_A_UNtvUHGa2_2(.din(n3632), .dout(n3629));
    jdff dff_A_1kIMQEqV3_2(.din(n189), .dout(n3632));
    jdff dff_A_yKYSx1j20_1(.din(n3638), .dout(n3635));
    jdff dff_A_pnq9SN502_1(.din(n3641), .dout(n3638));
    jdff dff_A_i5PFSqNZ8_1(.din(n3644), .dout(n3641));
    jdff dff_A_J05vdRn43_1(.din(n3647), .dout(n3644));
    jdff dff_A_BA8qXEPg4_1(.din(n3650), .dout(n3647));
    jdff dff_A_J4ywwvin4_1(.din(G472), .dout(n3650));
    jdff dff_B_DyUFSELa6_2(.din(n117), .dout(n3654));
    jdff dff_B_LVp1aPXk1_2(.din(n3654), .dout(n3657));
    jdff dff_B_AE97KynP0_2(.din(n3657), .dout(n3660));
    jdff dff_B_d1Qt6Vw90_2(.din(n3660), .dout(n3663));
    jdff dff_A_90bTC5ic7_1(.din(n3668), .dout(n3665));
    jdff dff_A_UVej9Q6S7_1(.din(G217), .dout(n3668));
    jdff dff_A_749vA3zO2_2(.din(n3674), .dout(n3671));
    jdff dff_A_mEDlAG3r4_2(.din(n3677), .dout(n3674));
    jdff dff_A_cIAEdAzU8_2(.din(G217), .dout(n3677));
    jdff dff_A_tPK35H4x3_0(.din(n3683), .dout(n3680));
    jdff dff_A_UQwIdcxJ2_0(.din(n3686), .dout(n3683));
    jdff dff_A_xCadTaOD3_0(.din(n3689), .dout(n3686));
    jdff dff_A_Co9J3NuT7_0(.din(n3692), .dout(n3689));
    jdff dff_A_dmJ8NtAT6_0(.din(n3695), .dout(n3692));
    jdff dff_A_5OU4Hzhe9_0(.din(n3698), .dout(n3695));
    jdff dff_A_ZrJcMgV21_0(.din(n3701), .dout(n3698));
    jdff dff_A_XOWBeYFi1_0(.din(n3704), .dout(n3701));
    jdff dff_A_4vKkhNU22_0(.din(n3707), .dout(n3704));
    jdff dff_A_4opZYrHl7_0(.din(n498), .dout(n3707));
    jdff dff_B_aY3Muk5q7_1(.din(n494), .dout(n3711));
    jdff dff_B_hdLbOZDB0_1(.din(n3711), .dout(n3714));
    jdff dff_B_pKaR8eaA2_1(.din(n3714), .dout(n3717));
    jdff dff_B_Z3x4UZAt1_0(.din(n87), .dout(n3720));
    jdff dff_B_qBlcKSpa6_0(.din(n3720), .dout(n3723));
    jdff dff_B_HZXyvK1o2_0(.din(n3723), .dout(n3726));
    jdff dff_A_lWle4vzx4_2(.din(n3731), .dout(n3728));
    jdff dff_A_ND1zml4C2_2(.din(n3734), .dout(n3731));
    jdff dff_A_zGKtC6DJ0_2(.din(n3737), .dout(n3734));
    jdff dff_A_qbrnQueL8_2(.din(n68), .dout(n3737));
    jdff dff_A_DE4xhmAQ3_0(.din(n3743), .dout(n3740));
    jdff dff_A_wrXkq0xj6_0(.din(n3746), .dout(n3743));
    jdff dff_A_F0OlzLAD1_0(.din(n64), .dout(n3746));
    jdff dff_A_NYHFwaqr6_0(.din(n3752), .dout(n3749));
    jdff dff_A_LY3FGZA26_0(.din(n3755), .dout(n3752));
    jdff dff_A_09DJ5dNl8_0(.din(n3758), .dout(n3755));
    jdff dff_A_ZsGqYRqj6_0(.din(n3761), .dout(n3758));
    jdff dff_A_TJWDZQVb4_0(.din(n3764), .dout(n3761));
    jdff dff_A_dkTleeez0_0(.din(n106), .dout(n3764));
    jdff dff_A_KgoQ2qci2_2(.din(n3770), .dout(n3767));
    jdff dff_A_5C5HgrQm5_2(.din(n3773), .dout(n3770));
    jdff dff_A_g1cQAKUA6_2(.din(n3776), .dout(n3773));
    jdff dff_A_iVMlshMV6_2(.din(n106), .dout(n3776));
    jdff dff_A_yQejMPDK3_0(.din(n3783), .dout(n3779));
    jdff dff_B_UXWqgLLL9_3(.din(n909), .dout(n3783));
    jdff dff_B_7FRH8gBm4_1(.din(n588), .dout(n3786));
    jdff dff_B_wYNYSM4x6_1(.din(n3786), .dout(n3789));
    jdff dff_B_fMGbrcGh6_1(.din(n3789), .dout(n3792));
    jdff dff_B_gK9l3Sqx9_1(.din(n3792), .dout(n3795));
    jdff dff_B_Jx9tTa653_1(.din(n3795), .dout(n3798));
    jdff dff_A_ID1k2XuY2_0(.din(n3803), .dout(n3800));
    jdff dff_A_d7FDJCNO2_0(.din(n3806), .dout(n3803));
    jdff dff_A_XvdFCzrw3_0(.din(n3809), .dout(n3806));
    jdff dff_A_plQxmdKp7_0(.din(n3812), .dout(n3809));
    jdff dff_A_vUaupqrr8_0(.din(n3815), .dout(n3812));
    jdff dff_A_gB9U7PJY9_0(.din(n3818), .dout(n3815));
    jdff dff_A_cMugvh9q4_0(.din(n3821), .dout(n3818));
    jdff dff_A_TDbpR4YG0_0(.din(n3824), .dout(n3821));
    jdff dff_A_2UAMgQJC5_0(.din(n3827), .dout(n3824));
    jdff dff_A_0FoaCd5f8_0(.din(n3830), .dout(n3827));
    jdff dff_A_c18q2Jzj9_0(.din(n3833), .dout(n3830));
    jdff dff_A_O0ethJcU8_0(.din(n286), .dout(n3833));
    jdff dff_B_EMzFG6GW9_1(.din(n270), .dout(n3837));
    jdff dff_B_2VYMP6Op9_1(.din(n3837), .dout(n3840));
    jdff dff_B_skuoW42i7_2(.din(G227), .dout(n3843));
    jdff dff_A_6D5aWB4x7_0(.din(n3848), .dout(n3845));
    jdff dff_A_O3vkfvPD5_0(.din(n3851), .dout(n3848));
    jdff dff_A_xNFSjN763_0(.din(n3854), .dout(n3851));
    jdff dff_A_euZgJ5on4_0(.din(n3857), .dout(n3854));
    jdff dff_A_ZlbdMtWu2_0(.din(n3860), .dout(n3857));
    jdff dff_A_QbEWsmZH7_0(.din(n3863), .dout(n3860));
    jdff dff_A_TdzEgtCD0_0(.din(n3866), .dout(n3863));
    jdff dff_A_y8dDQ0a08_0(.din(n3869), .dout(n3866));
    jdff dff_A_5zEdiTvk8_0(.din(n3872), .dout(n3869));
    jdff dff_A_RJ5QVG8f1_0(.din(n3875), .dout(n3872));
    jdff dff_A_wKRISSfC8_0(.din(n3878), .dout(n3875));
    jdff dff_A_ErJwq7to0_0(.din(G140), .dout(n3878));
    jdff dff_A_e3lVX8gh2_2(.din(n3884), .dout(n3881));
    jdff dff_A_gIN7R3uf1_2(.din(n3887), .dout(n3884));
    jdff dff_A_mERP0ZkL1_2(.din(n3890), .dout(n3887));
    jdff dff_A_c70Dbpyw4_2(.din(n3893), .dout(n3890));
    jdff dff_A_7ZWMuhfi8_2(.din(n3896), .dout(n3893));
    jdff dff_A_TyI5Y8M08_2(.din(G469), .dout(n3896));
    jdff dff_B_WcRU6Qft7_2(.din(n901), .dout(n3900));
    jdff dff_B_7quUQe1I0_2(.din(n3900), .dout(n3903));
    jdff dff_B_pJ0ykcTy3_2(.din(n3903), .dout(n3906));
    jdff dff_A_aO2f3qcc7_0(.din(n3911), .dout(n3908));
    jdff dff_A_XNfeC4qt2_0(.din(n3914), .dout(n3911));
    jdff dff_A_VthqGAlY9_0(.din(n3917), .dout(n3914));
    jdff dff_A_tqhHZpRV0_0(.din(n266), .dout(n3917));
    jdff dff_B_7iPPSUpd2_1(.din(n262), .dout(n3921));
    jdff dff_A_5VXt3w777_0(.din(n3926), .dout(n3923));
    jdff dff_A_7Jpnt4JB2_0(.din(n3929), .dout(n3926));
    jdff dff_A_PqzGkrR80_0(.din(n3932), .dout(n3929));
    jdff dff_A_HEbrDUYk4_0(.din(n106), .dout(n3932));
    jdff dff_A_xGppPr3k5_1(.din(G234), .dout(n3935));
    jdff dff_A_3T0Mu2XP9_2(.din(G234), .dout(n3938));
    jdff dff_A_0asksFzo1_1(.din(n3944), .dout(n3941));
    jdff dff_A_WhLdinJl8_1(.din(G221), .dout(n3944));
    jdff dff_A_L7rbIXSV3_1(.din(n671), .dout(n3947));
    jdff dff_B_f02cB3R30_1(.din(n667), .dout(n3951));
    jdff dff_B_JeWlBlYS1_1(.din(n3951), .dout(n3954));
    jdff dff_B_hXeRC8QT0_1(.din(n3954), .dout(n3957));
    jdff dff_A_x1lg016P1_0(.din(n3962), .dout(n3959));
    jdff dff_A_j272sTqQ3_0(.din(n3965), .dout(n3962));
    jdff dff_A_gLpiljix5_0(.din(n3968), .dout(n3965));
    jdff dff_A_9Vav6S578_0(.din(n3971), .dout(n3968));
    jdff dff_A_vhbPjJiy3_0(.din(n3974), .dout(n3971));
    jdff dff_A_H88aFHDB1_0(.din(n3977), .dout(n3974));
    jdff dff_A_DHK4VAkF2_0(.din(n3980), .dout(n3977));
    jdff dff_A_ft3kdH7l3_0(.din(n3983), .dout(n3980));
    jdff dff_A_OI8DS2hM9_0(.din(n3986), .dout(n3983));
    jdff dff_A_oNSKDJch6_0(.din(n3989), .dout(n3986));
    jdff dff_A_EBXwMR433_0(.din(n3992), .dout(n3989));
    jdff dff_A_ZhXSyGLz0_0(.din(n247), .dout(n3992));
    jdff dff_B_jhzHQqfo5_1(.din(n235), .dout(n3996));
    jdff dff_A_hGaPrqic9_0(.din(n4001), .dout(n3998));
    jdff dff_A_BUEBrPCd2_0(.din(n4004), .dout(n4001));
    jdff dff_A_hKYDeIqG7_0(.din(n4007), .dout(n4004));
    jdff dff_A_LK2anFOc8_0(.din(n4010), .dout(n4007));
    jdff dff_A_GoHPD5xI5_0(.din(n4013), .dout(n4010));
    jdff dff_A_MP3BtIz50_0(.din(n4016), .dout(n4013));
    jdff dff_A_2EprVAK18_0(.din(n4019), .dout(n4016));
    jdff dff_A_e5FFRQJK9_0(.din(n4022), .dout(n4019));
    jdff dff_A_71AJuITo6_0(.din(n4025), .dout(n4022));
    jdff dff_A_ABJqDcHw9_0(.din(n4028), .dout(n4025));
    jdff dff_A_WCLJcx8e0_0(.din(n4031), .dout(n4028));
    jdff dff_A_wEwstavb2_0(.din(G125), .dout(n4031));
    jdff dff_A_guNlDc5m9_1(.din(n4037), .dout(n4034));
    jdff dff_A_oICwdoW57_1(.din(G125), .dout(n4037));
    jdff dff_B_8hXZiefv1_2(.din(G224), .dout(n4041));
    jdff dff_A_rfpRIPBm1_0(.din(n4046), .dout(n4043));
    jdff dff_A_w8A4JYm67_0(.din(n4049), .dout(n4046));
    jdff dff_A_ADPXycaA9_0(.din(n4052), .dout(n4049));
    jdff dff_A_FdJbRLZR0_0(.din(n4055), .dout(n4052));
    jdff dff_A_JAW0FIg22_0(.din(n4058), .dout(n4055));
    jdff dff_A_LW17otL16_0(.din(n4061), .dout(n4058));
    jdff dff_A_eFpoyJQ54_0(.din(n4064), .dout(n4061));
    jdff dff_A_0ztDfp9y9_0(.din(n4067), .dout(n4064));
    jdff dff_A_7MthCdBr7_0(.din(n4070), .dout(n4067));
    jdff dff_A_TzaH7j9q2_0(.din(n4073), .dout(n4070));
    jdff dff_A_yMA7LU7d8_0(.din(n4076), .dout(n4073));
    jdff dff_A_9wStfIcu0_0(.din(n4079), .dout(n4076));
    jdff dff_A_Mjp2c5pP9_0(.din(n231), .dout(n4079));
    jdff dff_B_FXE00Kze7_1(.din(n215), .dout(n4083));
    jdff dff_A_SZ1Nm9Cs6_0(.din(n4088), .dout(n4085));
    jdff dff_A_b8kOHhoQ6_0(.din(n4091), .dout(n4088));
    jdff dff_A_3BvIEyqz4_0(.din(n4094), .dout(n4091));
    jdff dff_A_fl5DajHF6_0(.din(n4097), .dout(n4094));
    jdff dff_A_f9VF20vk0_0(.din(n4100), .dout(n4097));
    jdff dff_A_N8KbK16P5_0(.din(n4103), .dout(n4100));
    jdff dff_A_ZrfOKXBg8_0(.din(n4106), .dout(n4103));
    jdff dff_A_XTL9CeRp9_0(.din(n4109), .dout(n4106));
    jdff dff_A_TeErh5ES0_0(.din(n4112), .dout(n4109));
    jdff dff_A_w9oDyhL51_0(.din(n4115), .dout(n4112));
    jdff dff_A_DYKoNI6Y5_0(.din(n4118), .dout(n4115));
    jdff dff_A_w6XTsMsq8_0(.din(G107), .dout(n4118));
    jdff dff_A_97FbSwfK4_0(.din(n4124), .dout(n4121));
    jdff dff_A_GoqsyYIm8_0(.din(n4127), .dout(n4124));
    jdff dff_A_T4Eaq92Z3_0(.din(n4130), .dout(n4127));
    jdff dff_A_zElM6zFu1_0(.din(n4133), .dout(n4130));
    jdff dff_A_DRxUm7kI2_0(.din(n4136), .dout(n4133));
    jdff dff_A_3yPtjfDy8_0(.din(n4139), .dout(n4136));
    jdff dff_A_e8loeeor5_0(.din(n4142), .dout(n4139));
    jdff dff_A_05FENPcz7_0(.din(n4145), .dout(n4142));
    jdff dff_A_ec6pBWD25_0(.din(n4148), .dout(n4145));
    jdff dff_A_9IfFmerl9_0(.din(n4151), .dout(n4148));
    jdff dff_A_W4DPFxFO0_0(.din(n4154), .dout(n4151));
    jdff dff_A_PB4RuL8e9_0(.din(G104), .dout(n4154));
    jdff dff_A_WtxmHIdG9_1(.din(n4160), .dout(n4157));
    jdff dff_A_ADaMUmKc6_1(.din(G104), .dout(n4160));
    jdff dff_A_Xk15ibSQ5_1(.din(G122), .dout(n4163));
    jdff dff_A_kOA2vvfP0_1(.din(n4169), .dout(n4166));
    jdff dff_A_GoWajBuW7_1(.din(n4172), .dout(n4169));
    jdff dff_A_UdgX3NmM7_1(.din(n4175), .dout(n4172));
    jdff dff_A_huAXcbKv0_1(.din(n4178), .dout(n4175));
    jdff dff_A_Jqqv8qbg7_1(.din(n4181), .dout(n4178));
    jdff dff_A_vATM0Lp49_1(.din(n4184), .dout(n4181));
    jdff dff_A_RV81MCiQ5_1(.din(n4187), .dout(n4184));
    jdff dff_A_f7OK7zOE3_1(.din(n4190), .dout(n4187));
    jdff dff_A_YsiZRDlq9_1(.din(n4193), .dout(n4190));
    jdff dff_A_lJjo43g72_1(.din(n4196), .dout(n4193));
    jdff dff_A_d0Eel5RY2_1(.din(n4199), .dout(n4196));
    jdff dff_A_EyY3UJfQ7_1(.din(G122), .dout(n4199));
    jdff dff_A_EeE4pWsK2_2(.din(G122), .dout(n4202));
    jdff dff_A_tyLlt4Ug9_1(.din(n4208), .dout(n4205));
    jdff dff_A_etytuETZ9_1(.din(n4211), .dout(n4208));
    jdff dff_A_11apbKMy5_1(.din(n4214), .dout(n4211));
    jdff dff_A_GI9ubTPs6_1(.din(n4217), .dout(n4214));
    jdff dff_A_1FZCsts23_1(.din(G110), .dout(n4217));
    jdff dff_A_S7LbMjC51_1(.din(n4223), .dout(n4220));
    jdff dff_A_ObpxlGIK4_1(.din(n4226), .dout(n4223));
    jdff dff_A_0NJh9BDP9_1(.din(n4229), .dout(n4226));
    jdff dff_A_xzrtJekW4_1(.din(n4232), .dout(n4229));
    jdff dff_A_wNZ0DuLF0_1(.din(n4235), .dout(n4232));
    jdff dff_A_95ahYNiN7_1(.din(n4238), .dout(n4235));
    jdff dff_A_6vbxWAv54_1(.din(n4241), .dout(n4238));
    jdff dff_A_O4L5RZ7b7_1(.din(n4244), .dout(n4241));
    jdff dff_A_9G3HKwwo0_1(.din(n4247), .dout(n4244));
    jdff dff_A_qFoE6ANk9_1(.din(n4250), .dout(n4247));
    jdff dff_A_fxY1ZImU6_1(.din(n4253), .dout(n4250));
    jdff dff_A_6FnxbwUU6_1(.din(G110), .dout(n4253));
    jdff dff_A_wCCgcxh21_1(.din(n4259), .dout(n4256));
    jdff dff_A_hjgtmlav3_1(.din(n4262), .dout(n4259));
    jdff dff_A_ntsyURLv6_1(.din(n4265), .dout(n4262));
    jdff dff_A_sq6nP6G67_1(.din(n106), .dout(n4265));
    jdff dff_A_dSjSA72F1_1(.din(n4271), .dout(n4268));
    jdff dff_A_hwV4ctbQ9_1(.din(n4274), .dout(n4271));
    jdff dff_A_RT5C6dx18_1(.din(n4277), .dout(n4274));
    jdff dff_A_5QxyESWo5_1(.din(n208), .dout(n4277));
    jdff dff_A_3twR1F1A9_0(.din(n4283), .dout(n4280));
    jdff dff_A_lly5St5y0_0(.din(n4286), .dout(n4283));
    jdff dff_A_E0hdVmTV6_0(.din(n4289), .dout(n4286));
    jdff dff_A_izuiToZY1_0(.din(n4292), .dout(n4289));
    jdff dff_A_ASA7AT1X9_0(.din(n201), .dout(n4292));
    jdff dff_A_GezeG4B26_1(.din(n4298), .dout(n4295));
    jdff dff_A_94DAfcxq4_1(.din(n4301), .dout(n4298));
    jdff dff_A_2Qz32MAY7_1(.din(n4304), .dout(n4301));
    jdff dff_A_3vajMS4s9_1(.din(n4307), .dout(n4304));
    jdff dff_A_xnFTH5ZX1_1(.din(n201), .dout(n4307));
    jdff dff_A_9v5QviIV3_2(.din(n4313), .dout(n4310));
    jdff dff_A_tUC0hJ4s2_2(.din(n4316), .dout(n4313));
    jdff dff_A_uj7b49bG5_2(.din(n4319), .dout(n4316));
    jdff dff_A_71sARR4R6_2(.din(n4322), .dout(n4319));
    jdff dff_A_dFpJWWmH4_2(.din(n4325), .dout(n4322));
    jdff dff_A_eXeabmUB1_2(.din(n4328), .dout(n4325));
    jdff dff_A_WylMPeS41_2(.din(G902), .dout(n4328));
    jdff dff_A_C8ITO4682_1(.din(G214), .dout(n4331));
    jdff dff_A_omvqrot23_0(.din(n4337), .dout(n4334));
    jdff dff_A_z1FKsQwb4_0(.din(n4340), .dout(n4337));
    jdff dff_A_LVNl98VB2_0(.din(n4343), .dout(n4340));
    jdff dff_A_YdIrpSVj6_0(.din(n4346), .dout(n4343));
    jdff dff_A_LJ8Gi4uF8_0(.din(n4349), .dout(n4346));
    jdff dff_A_DZEGczG83_0(.din(n4352), .dout(n4349));
    jdff dff_A_KMClJIRV1_0(.din(n4355), .dout(n4352));
    jdff dff_A_M1oAQNKf2_0(.din(n4358), .dout(n4355));
    jdff dff_A_cNNtsd1I4_0(.din(n4361), .dout(n4358));
    jdff dff_A_qtYt3qJj9_0(.din(n4364), .dout(n4361));
    jdff dff_A_QEH7dcRk1_0(.din(n4367), .dout(n4364));
    jdff dff_A_wSqvZeYI9_0(.din(n181), .dout(n4367));
    jdff dff_A_UaBnAubx0_0(.din(n4373), .dout(n4370));
    jdff dff_A_c6EKCiTg3_0(.din(n4376), .dout(n4373));
    jdff dff_A_dAvRHgeN0_0(.din(n4379), .dout(n4376));
    jdff dff_A_hkaXSMhD4_0(.din(n4382), .dout(n4379));
    jdff dff_A_ceF5DLAr8_0(.din(n4385), .dout(n4382));
    jdff dff_A_v9tLWDIF1_0(.din(n4388), .dout(n4385));
    jdff dff_A_xgo6MV9X2_0(.din(n4391), .dout(n4388));
    jdff dff_A_CBh5iyhF0_0(.din(n4394), .dout(n4391));
    jdff dff_A_VLo057qZ4_0(.din(n4397), .dout(n4394));
    jdff dff_A_TyYdHk1b8_0(.din(n4400), .dout(n4397));
    jdff dff_A_OnKm0gGs9_0(.din(n4403), .dout(n4400));
    jdff dff_A_kfRW8fpl9_0(.din(G953), .dout(n4403));
    jdff dff_A_1DgrQCxR4_1(.din(n4409), .dout(n4406));
    jdff dff_A_QPs4KyXP2_1(.din(n4412), .dout(n4409));
    jdff dff_A_ItqCFU3O9_1(.din(n4415), .dout(n4412));
    jdff dff_A_uLPdK8m11_1(.din(n4418), .dout(n4415));
    jdff dff_A_sj9vVAaV6_1(.din(n4421), .dout(n4418));
    jdff dff_A_c9chWVhq5_1(.din(n4424), .dout(n4421));
    jdff dff_A_eWvczxoQ7_1(.din(n4427), .dout(n4424));
    jdff dff_A_NzHc1JiS4_1(.din(n4430), .dout(n4427));
    jdff dff_A_5CQyyH1w0_1(.din(n4433), .dout(n4430));
    jdff dff_A_t9EyqNw49_1(.din(n4436), .dout(n4433));
    jdff dff_A_HKSalTAP3_1(.din(n4439), .dout(n4436));
    jdff dff_A_CpSt5fEB7_1(.din(n4442), .dout(n4439));
    jdff dff_A_17b44fcI5_1(.din(n4445), .dout(n4442));
    jdff dff_A_8BXKGvxZ3_1(.din(n4448), .dout(n4445));
    jdff dff_A_NfEoZtfz9_1(.din(G953), .dout(n4448));
    jdff dff_A_aJrrWy2t9_2(.din(n4454), .dout(n4451));
    jdff dff_A_aypXjXkt3_2(.din(n4457), .dout(n4454));
    jdff dff_A_PNIcb18Q8_2(.din(n4460), .dout(n4457));
    jdff dff_A_OHQTwM1G8_2(.din(n4463), .dout(n4460));
    jdff dff_A_KHcooSNk5_2(.din(n4466), .dout(n4463));
    jdff dff_A_4ckL2wm82_2(.din(n4469), .dout(n4466));
    jdff dff_A_sgmh0wWz7_2(.din(n4472), .dout(n4469));
    jdff dff_A_NwLwOxON9_2(.din(n4475), .dout(n4472));
    jdff dff_A_1IFijKqr5_2(.din(n4478), .dout(n4475));
    jdff dff_A_Dr0R36Qq2_2(.din(n4481), .dout(n4478));
    jdff dff_A_FAXEgT0e3_2(.din(n4484), .dout(n4481));
    jdff dff_A_3VXP8UtH9_2(.din(n4487), .dout(n4484));
    jdff dff_A_PqbbI6gb8_2(.din(n4490), .dout(n4487));
    jdff dff_A_BnXwzpHc0_2(.din(n4493), .dout(n4490));
    jdff dff_A_MewQL7980_2(.din(G953), .dout(n4493));
    jdff dff_A_jtdazSx98_1(.din(G210), .dout(n4496));
    jdff dff_A_32dO2mgZ8_0(.din(n4502), .dout(n4499));
    jdff dff_A_y6vKYzLK4_0(.din(n4505), .dout(n4502));
    jdff dff_A_nSLHMqQ46_0(.din(n4508), .dout(n4505));
    jdff dff_A_q1UogLyh4_0(.din(n4511), .dout(n4508));
    jdff dff_A_z87XFPGG2_0(.din(n4514), .dout(n4511));
    jdff dff_A_I9lUJXPJ2_0(.din(n4517), .dout(n4514));
    jdff dff_A_tkXz10Lf5_0(.din(n4520), .dout(n4517));
    jdff dff_A_eVRXWvqv9_0(.din(n4523), .dout(n4520));
    jdff dff_A_YqIhGlMJ0_0(.din(n4526), .dout(n4523));
    jdff dff_A_7FVeCVei6_0(.din(n4529), .dout(n4526));
    jdff dff_A_fjjRkyM94_0(.din(n4536), .dout(n4529));
    jdff dff_A_xokxmThT8_2(.din(n4536), .dout(n4532));
    jdff dff_B_nhW2gutN0_3(.din(G101), .dout(n4536));
    jdff dff_A_zw6Yoo2x9_1(.din(n158), .dout(n4538));
    jdff dff_A_QYrbG5kf3_0(.din(n4544), .dout(n4541));
    jdff dff_A_g1ggyjHE6_0(.din(n4547), .dout(n4544));
    jdff dff_A_qlAwMW466_0(.din(n4550), .dout(n4547));
    jdff dff_A_uoLsdpJJ8_0(.din(n4553), .dout(n4550));
    jdff dff_A_TLRcHvBK0_0(.din(n4556), .dout(n4553));
    jdff dff_A_G3SHcqRu0_0(.din(n4559), .dout(n4556));
    jdff dff_A_F5vqeNN54_0(.din(n4562), .dout(n4559));
    jdff dff_A_4QrWqADd8_0(.din(n4565), .dout(n4562));
    jdff dff_A_HqrT7uBB3_0(.din(n4568), .dout(n4565));
    jdff dff_A_uqjWhDGs4_0(.din(n4571), .dout(n4568));
    jdff dff_A_rEvntC530_0(.din(n4574), .dout(n4571));
    jdff dff_A_kWji1Z9g6_0(.din(G119), .dout(n4574));
    jdff dff_A_ixzV3uN88_0(.din(n4580), .dout(n4577));
    jdff dff_A_7QMqde7C1_0(.din(n4583), .dout(n4580));
    jdff dff_A_fTN0M8Nl9_0(.din(n4586), .dout(n4583));
    jdff dff_A_Xvs9Klv14_0(.din(n4589), .dout(n4586));
    jdff dff_A_kYAyEiQQ5_0(.din(n4592), .dout(n4589));
    jdff dff_A_E4mlpWHo2_0(.din(n4595), .dout(n4592));
    jdff dff_A_hlClqw9d9_0(.din(n4598), .dout(n4595));
    jdff dff_A_NKLr0QsT4_0(.din(n4601), .dout(n4598));
    jdff dff_A_9lrOEVyf1_0(.din(n4604), .dout(n4601));
    jdff dff_A_1jlZLf9J6_0(.din(n4607), .dout(n4604));
    jdff dff_A_UbfACKGM5_0(.din(n4610), .dout(n4607));
    jdff dff_A_AQxkgjvZ4_0(.din(G116), .dout(n4610));
    jdff dff_A_vFPHv5Kn6_0(.din(n4616), .dout(n4613));
    jdff dff_A_5uLjVev71_0(.din(n4619), .dout(n4616));
    jdff dff_A_mhvx7r855_0(.din(n4622), .dout(n4619));
    jdff dff_A_RNYdsNw95_0(.din(n4625), .dout(n4622));
    jdff dff_A_LqK2UbH56_0(.din(n4628), .dout(n4625));
endmodule

