/*

c3540:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jdff: 1943
	jand: 535
	jor: 374

Summary:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jdff: 1943
	jand: 535
	jor: 374
*/

module c3540(gclk, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402);
	input gclk;
	input G1;
	input G13;
	input G20;
	input G33;
	input G41;
	input G45;
	input G50;
	input G58;
	input G68;
	input G77;
	input G87;
	input G97;
	input G107;
	input G116;
	input G124;
	input G125;
	input G128;
	input G132;
	input G137;
	input G143;
	input G150;
	input G159;
	input G169;
	input G179;
	input G190;
	input G200;
	input G213;
	input G222;
	input G223;
	input G226;
	input G232;
	input G238;
	input G244;
	input G250;
	input G257;
	input G264;
	input G270;
	input G274;
	input G283;
	input G294;
	input G303;
	input G311;
	input G317;
	input G322;
	input G326;
	input G329;
	input G330;
	input G343;
	input G1698;
	input G2897;
	output G353;
	output G355;
	output G361;
	output G358;
	output G351;
	output G372;
	output G369;
	output G399;
	output G364;
	output G396;
	output G384;
	output G367;
	output G387;
	output G393;
	output G390;
	output G378;
	output G375;
	output G381;
	output G407;
	output G409;
	output G405;
	output G402;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[2:0] w_G1_2;
	wire[1:0] w_G1_3;
	wire[2:0] w_G13_0;
	wire[1:0] w_G13_1;
	wire[2:0] w_G20_0;
	wire[2:0] w_G20_1;
	wire[2:0] w_G20_2;
	wire[2:0] w_G20_3;
	wire[2:0] w_G20_4;
	wire[2:0] w_G20_5;
	wire[2:0] w_G20_6;
	wire[1:0] w_G20_7;
	wire[2:0] w_G33_0;
	wire[2:0] w_G33_1;
	wire[2:0] w_G33_2;
	wire[2:0] w_G33_3;
	wire[2:0] w_G33_4;
	wire[2:0] w_G33_5;
	wire[2:0] w_G33_6;
	wire[2:0] w_G33_7;
	wire[2:0] w_G33_8;
	wire[2:0] w_G33_9;
	wire[2:0] w_G33_10;
	wire[2:0] w_G33_11;
	wire[2:0] w_G41_0;
	wire[1:0] w_G41_1;
	wire[2:0] w_G45_0;
	wire[2:0] w_G45_1;
	wire[2:0] w_G50_0;
	wire[2:0] w_G50_1;
	wire[2:0] w_G50_2;
	wire[2:0] w_G50_3;
	wire[2:0] w_G50_4;
	wire[2:0] w_G50_5;
	wire[2:0] w_G58_0;
	wire[2:0] w_G58_1;
	wire[2:0] w_G58_2;
	wire[2:0] w_G58_3;
	wire[2:0] w_G58_4;
	wire[1:0] w_G58_5;
	wire[2:0] w_G68_0;
	wire[2:0] w_G68_1;
	wire[2:0] w_G68_2;
	wire[2:0] w_G68_3;
	wire[2:0] w_G68_4;
	wire[1:0] w_G68_5;
	wire[2:0] w_G77_0;
	wire[2:0] w_G77_1;
	wire[2:0] w_G77_2;
	wire[2:0] w_G77_3;
	wire[2:0] w_G77_4;
	wire[1:0] w_G77_5;
	wire[2:0] w_G87_0;
	wire[2:0] w_G87_1;
	wire[2:0] w_G87_2;
	wire[2:0] w_G87_3;
	wire[2:0] w_G97_0;
	wire[2:0] w_G97_1;
	wire[2:0] w_G97_2;
	wire[2:0] w_G97_3;
	wire[2:0] w_G97_4;
	wire[1:0] w_G97_5;
	wire[2:0] w_G107_0;
	wire[2:0] w_G107_1;
	wire[2:0] w_G107_2;
	wire[2:0] w_G107_3;
	wire[2:0] w_G107_4;
	wire[1:0] w_G107_5;
	wire[2:0] w_G116_0;
	wire[2:0] w_G116_1;
	wire[2:0] w_G116_2;
	wire[2:0] w_G116_3;
	wire[2:0] w_G116_4;
	wire[1:0] w_G125_0;
	wire[2:0] w_G128_0;
	wire[2:0] w_G132_0;
	wire[1:0] w_G132_1;
	wire[2:0] w_G137_0;
	wire[2:0] w_G137_1;
	wire[2:0] w_G143_0;
	wire[2:0] w_G143_1;
	wire[1:0] w_G143_2;
	wire[2:0] w_G150_0;
	wire[2:0] w_G150_1;
	wire[2:0] w_G150_2;
	wire[1:0] w_G150_3;
	wire[2:0] w_G159_0;
	wire[2:0] w_G159_1;
	wire[2:0] w_G159_2;
	wire[2:0] w_G159_3;
	wire[2:0] w_G169_0;
	wire[1:0] w_G169_1;
	wire[2:0] w_G179_0;
	wire[2:0] w_G179_1;
	wire[2:0] w_G179_2;
	wire[2:0] w_G190_0;
	wire[2:0] w_G190_1;
	wire[2:0] w_G190_2;
	wire[2:0] w_G190_3;
	wire[1:0] w_G190_4;
	wire[2:0] w_G200_0;
	wire[2:0] w_G200_1;
	wire[2:0] w_G200_2;
	wire[2:0] w_G200_3;
	wire[2:0] w_G200_4;
	wire[2:0] w_G213_0;
	wire[1:0] w_G223_0;
	wire[2:0] w_G226_0;
	wire[1:0] w_G226_1;
	wire[2:0] w_G232_0;
	wire[2:0] w_G232_1;
	wire[2:0] w_G238_0;
	wire[2:0] w_G238_1;
	wire[2:0] w_G244_0;
	wire[2:0] w_G244_1;
	wire[2:0] w_G250_0;
	wire[2:0] w_G257_0;
	wire[2:0] w_G257_1;
	wire[2:0] w_G264_0;
	wire[1:0] w_G264_1;
	wire[2:0] w_G270_0;
	wire[2:0] w_G274_0;
	wire[2:0] w_G283_0;
	wire[2:0] w_G283_1;
	wire[2:0] w_G283_2;
	wire[2:0] w_G283_3;
	wire[2:0] w_G294_0;
	wire[2:0] w_G294_1;
	wire[2:0] w_G294_2;
	wire[1:0] w_G294_3;
	wire[2:0] w_G303_0;
	wire[2:0] w_G303_1;
	wire[2:0] w_G303_2;
	wire[2:0] w_G311_0;
	wire[2:0] w_G311_1;
	wire[2:0] w_G317_0;
	wire[1:0] w_G317_1;
	wire[2:0] w_G322_0;
	wire[1:0] w_G326_0;
	wire[1:0] w_G330_0;
	wire[1:0] w_G343_0;
	wire[2:0] w_G1698_0;
	wire w_G355_0;
	wire G355_fa_;
	wire[1:0] w_G396_0;
	wire G396_fa_;
	wire w_G384_0;
	wire G384_fa_;
	wire[1:0] w_G387_0;
	wire G387_fa_;
	wire[2:0] w_n72_0;
	wire[1:0] w_n72_1;
	wire[2:0] w_n73_0;
	wire[2:0] w_n73_1;
	wire[2:0] w_n73_2;
	wire[2:0] w_n74_0;
	wire[1:0] w_n74_1;
	wire[2:0] w_n75_0;
	wire[1:0] w_n75_1;
	wire[1:0] w_n76_0;
	wire[1:0] w_n77_0;
	wire[2:0] w_n79_0;
	wire[2:0] w_n80_0;
	wire[1:0] w_n80_1;
	wire[2:0] w_n81_0;
	wire[2:0] w_n85_0;
	wire[1:0] w_n86_0;
	wire[2:0] w_n88_0;
	wire[1:0] w_n88_1;
	wire[2:0] w_n91_0;
	wire[2:0] w_n91_1;
	wire[1:0] w_n93_0;
	wire[2:0] w_n97_0;
	wire[2:0] w_n97_1;
	wire[1:0] w_n97_2;
	wire[2:0] w_n98_0;
	wire[2:0] w_n98_1;
	wire[1:0] w_n98_2;
	wire[2:0] w_n103_0;
	wire[2:0] w_n105_0;
	wire[2:0] w_n105_1;
	wire[1:0] w_n105_2;
	wire[1:0] w_n106_0;
	wire[2:0] w_n112_0;
	wire[2:0] w_n112_1;
	wire[2:0] w_n112_2;
	wire[2:0] w_n112_3;
	wire[2:0] w_n112_4;
	wire[2:0] w_n112_5;
	wire[2:0] w_n113_0;
	wire[2:0] w_n113_1;
	wire[2:0] w_n113_2;
	wire[1:0] w_n113_3;
	wire[2:0] w_n114_0;
	wire[2:0] w_n114_1;
	wire[2:0] w_n115_0;
	wire[1:0] w_n115_1;
	wire[1:0] w_n116_0;
	wire[2:0] w_n118_0;
	wire[2:0] w_n121_0;
	wire[2:0] w_n122_0;
	wire[1:0] w_n122_1;
	wire[2:0] w_n123_0;
	wire[2:0] w_n123_1;
	wire[1:0] w_n131_0;
	wire[1:0] w_n135_0;
	wire[2:0] w_n137_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n144_0;
	wire[2:0] w_n146_0;
	wire[2:0] w_n146_1;
	wire[2:0] w_n146_2;
	wire[2:0] w_n146_3;
	wire[2:0] w_n147_0;
	wire[2:0] w_n148_0;
	wire[2:0] w_n148_1;
	wire[2:0] w_n148_2;
	wire[2:0] w_n148_3;
	wire[2:0] w_n148_4;
	wire[2:0] w_n148_5;
	wire[2:0] w_n148_6;
	wire[2:0] w_n148_7;
	wire[2:0] w_n148_8;
	wire[2:0] w_n148_9;
	wire[2:0] w_n149_0;
	wire[2:0] w_n149_1;
	wire[1:0] w_n149_2;
	wire[2:0] w_n151_0;
	wire[2:0] w_n151_1;
	wire[2:0] w_n151_2;
	wire[2:0] w_n151_3;
	wire[2:0] w_n151_4;
	wire[2:0] w_n152_0;
	wire[2:0] w_n152_1;
	wire[2:0] w_n152_2;
	wire[1:0] w_n152_3;
	wire[1:0] w_n154_0;
	wire[2:0] w_n155_0;
	wire[2:0] w_n155_1;
	wire[2:0] w_n155_2;
	wire[1:0] w_n155_3;
	wire[2:0] w_n157_0;
	wire[2:0] w_n161_0;
	wire[1:0] w_n161_1;
	wire[2:0] w_n162_0;
	wire[1:0] w_n163_0;
	wire[2:0] w_n166_0;
	wire[2:0] w_n166_1;
	wire[2:0] w_n166_2;
	wire[1:0] w_n166_3;
	wire[2:0] w_n170_0;
	wire[1:0] w_n172_0;
	wire[2:0] w_n179_0;
	wire[2:0] w_n179_1;
	wire[1:0] w_n180_0;
	wire[2:0] w_n185_0;
	wire[2:0] w_n185_1;
	wire[2:0] w_n185_2;
	wire[2:0] w_n185_3;
	wire[2:0] w_n189_0;
	wire[2:0] w_n189_1;
	wire[1:0] w_n189_2;
	wire[2:0] w_n190_0;
	wire[2:0] w_n190_1;
	wire[2:0] w_n191_0;
	wire[1:0] w_n195_0;
	wire[2:0] w_n196_0;
	wire[2:0] w_n196_1;
	wire[2:0] w_n196_2;
	wire[2:0] w_n197_0;
	wire[1:0] w_n197_1;
	wire[2:0] w_n199_0;
	wire[1:0] w_n199_1;
	wire[1:0] w_n201_0;
	wire[1:0] w_n205_0;
	wire[1:0] w_n206_0;
	wire[2:0] w_n210_0;
	wire[1:0] w_n213_0;
	wire[1:0] w_n214_0;
	wire[1:0] w_n218_0;
	wire[1:0] w_n219_0;
	wire[2:0] w_n221_0;
	wire[1:0] w_n228_0;
	wire[2:0] w_n229_0;
	wire[1:0] w_n230_0;
	wire[2:0] w_n231_0;
	wire[2:0] w_n234_0;
	wire[1:0] w_n241_0;
	wire[2:0] w_n242_0;
	wire[2:0] w_n243_0;
	wire[2:0] w_n246_0;
	wire[1:0] w_n246_1;
	wire[1:0] w_n249_0;
	wire[1:0] w_n255_0;
	wire[1:0] w_n257_0;
	wire[1:0] w_n259_0;
	wire[1:0] w_n261_0;
	wire[1:0] w_n262_0;
	wire[2:0] w_n269_0;
	wire[2:0] w_n269_1;
	wire[1:0] w_n270_0;
	wire[2:0] w_n271_0;
	wire[2:0] w_n271_1;
	wire[2:0] w_n274_0;
	wire[1:0] w_n278_0;
	wire[1:0] w_n279_0;
	wire[1:0] w_n281_0;
	wire[2:0] w_n288_0;
	wire[1:0] w_n288_1;
	wire[1:0] w_n296_0;
	wire[1:0] w_n298_0;
	wire[1:0] w_n300_0;
	wire[1:0] w_n303_0;
	wire[2:0] w_n312_0;
	wire[1:0] w_n312_1;
	wire[1:0] w_n315_0;
	wire[1:0] w_n320_0;
	wire[1:0] w_n324_0;
	wire[1:0] w_n328_0;
	wire[1:0] w_n334_0;
	wire[1:0] w_n339_0;
	wire[2:0] w_n346_0;
	wire[1:0] w_n346_1;
	wire[2:0] w_n355_0;
	wire[1:0] w_n355_1;
	wire[1:0] w_n362_0;
	wire[2:0] w_n367_0;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n374_0;
	wire[1:0] w_n381_0;
	wire[2:0] w_n382_0;
	wire[1:0] w_n382_1;
	wire[2:0] w_n385_0;
	wire[1:0] w_n385_1;
	wire[2:0] w_n387_0;
	wire[1:0] w_n387_1;
	wire[1:0] w_n390_0;
	wire[2:0] w_n401_0;
	wire[2:0] w_n404_0;
	wire[1:0] w_n405_0;
	wire[2:0] w_n407_0;
	wire[2:0] w_n407_1;
	wire[1:0] w_n407_2;
	wire[1:0] w_n412_0;
	wire[2:0] w_n420_0;
	wire[1:0] w_n420_1;
	wire[2:0] w_n425_0;
	wire[2:0] w_n425_1;
	wire[1:0] w_n426_0;
	wire[1:0] w_n430_0;
	wire[2:0] w_n436_0;
	wire[2:0] w_n439_0;
	wire[1:0] w_n439_1;
	wire[1:0] w_n445_0;
	wire[1:0] w_n446_0;
	wire[2:0] w_n455_0;
	wire[2:0] w_n462_0;
	wire[1:0] w_n465_0;
	wire[1:0] w_n474_0;
	wire[1:0] w_n475_0;
	wire[1:0] w_n478_0;
	wire[1:0] w_n479_0;
	wire[1:0] w_n483_0;
	wire[1:0] w_n484_0;
	wire[2:0] w_n492_0;
	wire[1:0] w_n507_0;
	wire[1:0] w_n508_0;
	wire[1:0] w_n511_0;
	wire[1:0] w_n512_0;
	wire[1:0] w_n516_0;
	wire[1:0] w_n517_0;
	wire[2:0] w_n519_0;
	wire[2:0] w_n519_1;
	wire[1:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n528_0;
	wire[1:0] w_n532_0;
	wire[1:0] w_n534_0;
	wire[2:0] w_n536_0;
	wire[1:0] w_n539_0;
	wire[1:0] w_n541_0;
	wire[2:0] w_n542_0;
	wire[1:0] w_n543_0;
	wire[2:0] w_n548_0;
	wire[1:0] w_n550_0;
	wire[2:0] w_n552_0;
	wire[1:0] w_n552_1;
	wire[2:0] w_n553_0;
	wire[2:0] w_n553_1;
	wire[2:0] w_n553_2;
	wire[2:0] w_n554_0;
	wire[2:0] w_n554_1;
	wire[2:0] w_n554_2;
	wire[2:0] w_n554_3;
	wire[1:0] w_n556_0;
	wire[1:0] w_n557_0;
	wire[2:0] w_n561_0;
	wire[2:0] w_n563_0;
	wire[1:0] w_n564_0;
	wire[1:0] w_n565_0;
	wire[1:0] w_n567_0;
	wire[2:0] w_n571_0;
	wire[2:0] w_n572_0;
	wire[2:0] w_n573_0;
	wire[2:0] w_n576_0;
	wire[1:0] w_n576_1;
	wire[2:0] w_n588_0;
	wire[1:0] w_n588_1;
	wire[2:0] w_n589_0;
	wire[2:0] w_n589_1;
	wire[2:0] w_n591_0;
	wire[1:0] w_n591_1;
	wire[2:0] w_n592_0;
	wire[2:0] w_n592_1;
	wire[1:0] w_n592_2;
	wire[2:0] w_n593_0;
	wire[1:0] w_n602_0;
	wire[2:0] w_n603_0;
	wire[2:0] w_n603_1;
	wire[1:0] w_n603_2;
	wire[2:0] w_n604_0;
	wire[2:0] w_n604_1;
	wire[1:0] w_n604_2;
	wire[2:0] w_n605_0;
	wire[2:0] w_n605_1;
	wire[2:0] w_n608_0;
	wire[2:0] w_n608_1;
	wire[2:0] w_n612_0;
	wire[2:0] w_n612_1;
	wire[2:0] w_n612_2;
	wire[2:0] w_n612_3;
	wire[1:0] w_n612_4;
	wire[2:0] w_n613_0;
	wire[1:0] w_n613_1;
	wire[1:0] w_n615_0;
	wire[1:0] w_n616_0;
	wire[2:0] w_n617_0;
	wire[2:0] w_n617_1;
	wire[2:0] w_n617_2;
	wire[2:0] w_n617_3;
	wire[2:0] w_n617_4;
	wire[2:0] w_n617_5;
	wire[1:0] w_n617_6;
	wire[1:0] w_n619_0;
	wire[1:0] w_n622_0;
	wire[2:0] w_n623_0;
	wire[2:0] w_n623_1;
	wire[2:0] w_n623_2;
	wire[2:0] w_n623_3;
	wire[2:0] w_n623_4;
	wire[1:0] w_n623_5;
	wire[1:0] w_n626_0;
	wire[2:0] w_n627_0;
	wire[2:0] w_n627_1;
	wire[2:0] w_n627_2;
	wire[2:0] w_n627_3;
	wire[2:0] w_n627_4;
	wire[2:0] w_n627_5;
	wire[2:0] w_n627_6;
	wire[1:0] w_n627_7;
	wire[2:0] w_n631_0;
	wire[2:0] w_n631_1;
	wire[2:0] w_n631_2;
	wire[2:0] w_n631_3;
	wire[2:0] w_n631_4;
	wire[2:0] w_n631_5;
	wire[2:0] w_n631_6;
	wire[1:0] w_n631_7;
	wire[2:0] w_n634_0;
	wire[2:0] w_n634_1;
	wire[2:0] w_n634_2;
	wire[2:0] w_n634_3;
	wire[1:0] w_n634_4;
	wire[2:0] w_n636_0;
	wire[2:0] w_n636_1;
	wire[2:0] w_n636_2;
	wire[2:0] w_n636_3;
	wire[2:0] w_n636_4;
	wire[2:0] w_n636_5;
	wire[2:0] w_n636_6;
	wire[1:0] w_n636_7;
	wire[1:0] w_n639_0;
	wire[2:0] w_n640_0;
	wire[2:0] w_n640_1;
	wire[2:0] w_n640_2;
	wire[2:0] w_n640_3;
	wire[2:0] w_n640_4;
	wire[2:0] w_n640_5;
	wire[2:0] w_n640_6;
	wire[1:0] w_n640_7;
	wire[2:0] w_n642_0;
	wire[2:0] w_n642_1;
	wire[2:0] w_n642_2;
	wire[2:0] w_n642_3;
	wire[2:0] w_n642_4;
	wire[2:0] w_n642_5;
	wire[2:0] w_n642_6;
	wire[1:0] w_n642_7;
	wire[1:0] w_n654_0;
	wire[1:0] w_n657_0;
	wire[1:0] w_n661_0;
	wire[2:0] w_n672_0;
	wire[1:0] w_n672_1;
	wire[2:0] w_n675_0;
	wire[1:0] w_n676_0;
	wire[1:0] w_n680_0;
	wire[1:0] w_n692_0;
	wire[2:0] w_n696_0;
	wire[2:0] w_n696_1;
	wire[1:0] w_n717_0;
	wire[1:0] w_n728_0;
	wire[2:0] w_n743_0;
	wire[1:0] w_n743_1;
	wire[1:0] w_n750_0;
	wire[1:0] w_n754_0;
	wire[2:0] w_n758_0;
	wire[1:0] w_n758_1;
	wire[1:0] w_n759_0;
	wire[1:0] w_n760_0;
	wire[2:0] w_n764_0;
	wire[2:0] w_n764_1;
	wire[1:0] w_n769_0;
	wire[2:0] w_n771_0;
	wire[1:0] w_n779_0;
	wire[1:0] w_n797_0;
	wire[1:0] w_n801_0;
	wire[1:0] w_n816_0;
	wire[1:0] w_n823_0;
	wire[1:0] w_n825_0;
	wire[2:0] w_n853_0;
	wire[2:0] w_n855_0;
	wire[2:0] w_n861_0;
	wire[1:0] w_n861_1;
	wire[1:0] w_n863_0;
	wire[1:0] w_n864_0;
	wire[1:0] w_n899_0;
	wire[1:0] w_n909_0;
	wire[2:0] w_n937_0;
	wire[1:0] w_n940_0;
	wire[1:0] w_n962_0;
	wire[2:0] w_n988_0;
	wire[1:0] w_n990_0;
	wire[2:0] w_n991_0;
	wire[1:0] w_n992_0;
	wire[2:0] w_n994_0;
	wire[2:0] w_n996_0;
	wire[1:0] w_n999_0;
	wire[2:0] w_n1001_0;
	wire[2:0] w_n1002_0;
	wire[1:0] w_n1003_0;
	wire[2:0] w_n1049_0;
	wire[1:0] w_n1052_0;
	wire[1:0] w_n1057_0;
	wire[1:0] w_n1059_0;
	wire[1:0] w_n1088_0;
	wire[2:0] w_n1114_0;
	wire[2:0] w_n1162_0;
	wire[1:0] w_n1164_0;
	wire[1:0] w_n1172_0;
	wire[1:0] w_n1175_0;
	wire[1:0] w_n1183_0;
	wire[1:0] w_n1184_0;
	wire[1:0] w_n1187_0;
	wire w_dff_B_8aZMsUSg1_1;
	wire w_dff_B_nTRQHFet8_0;
	wire w_dff_B_FHdOARZ04_0;
	wire w_dff_A_MDs6Vcnr7_1;
	wire w_dff_A_Cy55RF5Q7_1;
	wire w_dff_A_Fnp8WRIn0_0;
	wire w_dff_B_ldRFVe202_1;
	wire w_dff_B_j6waDMC76_0;
	wire w_dff_B_3gI0awUS0_0;
	wire w_dff_B_njzexcSK1_0;
	wire w_dff_B_t4i66qn88_0;
	wire w_dff_B_kVySOI6Y1_0;
	wire w_dff_B_rDlpP4Tm2_0;
	wire w_dff_B_7lYQBcTU9_0;
	wire w_dff_B_k6hK0ZL41_0;
	wire w_dff_B_MJ4Ko4900_0;
	wire w_dff_B_FFN7T7lW1_0;
	wire w_dff_B_Meiy2dWM6_0;
	wire w_dff_B_jmc7yEn00_0;
	wire w_dff_B_FBAA0OiE4_0;
	wire w_dff_B_qg1WDuVP3_0;
	wire w_dff_B_ll4EBX4T5_0;
	wire w_dff_B_rOe93E8Z0_0;
	wire w_dff_B_MIeghigj1_0;
	wire w_dff_B_toQfQAC32_0;
	wire w_dff_B_ZElfSDKJ4_0;
	wire w_dff_B_gfFi0Bru6_0;
	wire w_dff_B_rWmrLOuI8_0;
	wire w_dff_B_xcToyw074_0;
	wire w_dff_B_oXeKlS7g6_0;
	wire w_dff_B_SVhmJNuT3_0;
	wire w_dff_B_UazcTnMj9_0;
	wire w_dff_B_fMbyyNtm4_0;
	wire w_dff_B_9HLj2MZf8_0;
	wire w_dff_B_a03BJKRD2_0;
	wire w_dff_B_h20AqAp38_1;
	wire w_dff_B_KGWBjATJ3_0;
	wire w_dff_B_8dhPwf6t8_0;
	wire w_dff_B_A73Inxk12_0;
	wire w_dff_B_iUQfLqnQ3_0;
	wire w_dff_B_qUNMdAgl3_0;
	wire w_dff_B_5xQQZF0D0_0;
	wire w_dff_B_GKzjQE1R3_0;
	wire w_dff_B_WJA4ZsAw5_0;
	wire w_dff_B_sYnYWvBN0_0;
	wire w_dff_B_BIXpI8E30_0;
	wire w_dff_B_az5NFJ6w8_0;
	wire w_dff_B_xrkJsPzh4_0;
	wire w_dff_B_VBqfAsvq8_0;
	wire w_dff_B_GgxeHxsu5_0;
	wire w_dff_B_01o3erlq4_0;
	wire w_dff_B_kWKl3YgX2_0;
	wire w_dff_B_uToLvsbu0_0;
	wire w_dff_B_DrwagBmw7_0;
	wire w_dff_B_08UZhAAQ1_0;
	wire w_dff_A_kWsQxzyD4_1;
	wire w_dff_A_XPpM07ww0_1;
	wire w_dff_B_1ebv9Ywc6_0;
	wire w_dff_A_JrPOuNJj8_0;
	wire w_dff_B_C6myuNG13_1;
	wire w_dff_A_l8FyxM895_0;
	wire w_dff_B_YxMyLRdw2_1;
	wire w_dff_B_IhQIpIaA0_1;
	wire w_dff_B_B6DW9lbj3_1;
	wire w_dff_B_gtIhX11Z3_1;
	wire w_dff_B_96h1m6QL5_1;
	wire w_dff_B_G272gM9Z8_1;
	wire w_dff_B_ykvTJ1bc3_1;
	wire w_dff_B_mM3jbKiG4_1;
	wire w_dff_B_RO0M0pTf6_1;
	wire w_dff_B_TEkBKpVL7_1;
	wire w_dff_B_XpZeYqJT5_1;
	wire w_dff_B_yP207U600_1;
	wire w_dff_B_x4m8ajeN6_1;
	wire w_dff_B_5bux0arX6_1;
	wire w_dff_B_1mEcKKrc8_1;
	wire w_dff_B_k3KVRscA8_1;
	wire w_dff_B_Bq0kVR0O9_1;
	wire w_dff_B_aYZVBZi78_1;
	wire w_dff_B_ZqXARUce0_1;
	wire w_dff_B_xILg8HgC6_1;
	wire w_dff_B_aLbDCmTi0_1;
	wire w_dff_B_wXcETJsI9_1;
	wire w_dff_B_TJxq1Y5N5_1;
	wire w_dff_B_OvWgd3B04_1;
	wire w_dff_B_Ifi2zEUX1_1;
	wire w_dff_B_70Lh1d4I4_1;
	wire w_dff_A_RuAtsRXB7_0;
	wire w_dff_B_BIcvvNtC5_1;
	wire w_dff_B_0z1zdyUY5_1;
	wire w_dff_B_pDDrbT6h3_1;
	wire w_dff_B_Nua3Uscy5_1;
	wire w_dff_B_8ucCZc955_1;
	wire w_dff_B_vOUZ7sJR2_1;
	wire w_dff_B_OryVXVYG8_1;
	wire w_dff_B_L4z9TSUs1_1;
	wire w_dff_B_v3N1Brr01_1;
	wire w_dff_B_U8Syk4L07_1;
	wire w_dff_B_qiEjx3fb9_1;
	wire w_dff_B_ugKgAaRj7_1;
	wire w_dff_B_bsYBlFQC6_1;
	wire w_dff_B_r0Zni9ip3_1;
	wire w_dff_B_PHIVRap49_1;
	wire w_dff_B_3BXgcVFQ4_1;
	wire w_dff_B_8kFOkYio2_1;
	wire w_dff_B_HbyLvWG12_1;
	wire w_dff_B_9xpwargc1_1;
	wire w_dff_B_zEbeDmnE8_1;
	wire w_dff_B_AbOrrKBs0_1;
	wire w_dff_B_3gnqDvH62_1;
	wire w_dff_B_1Frq4AFi1_1;
	wire w_dff_B_r6us2hmd6_1;
	wire w_dff_B_kXptMM8s9_1;
	wire w_dff_B_ymAn6tCn5_1;
	wire w_dff_B_sJSKpJ2F1_1;
	wire w_dff_B_QHOGV6Yf9_1;
	wire w_dff_A_mHZxPKWf3_0;
	wire w_dff_A_VH2U8Oq64_0;
	wire w_dff_A_XBIBSthK4_0;
	wire w_dff_A_poTCiQoY4_0;
	wire w_dff_A_wAbsF8o51_0;
	wire w_dff_A_geEesXKv6_0;
	wire w_dff_A_Tmwd6mbF1_0;
	wire w_dff_A_vwSIPiSD5_0;
	wire w_dff_A_wVgi0O2n8_0;
	wire w_dff_A_UUiwvjWN7_0;
	wire w_dff_A_0ep7acPz3_0;
	wire w_dff_A_TBpBjb3h4_0;
	wire w_dff_A_Zko62mKg4_0;
	wire w_dff_A_5rFFZyZ71_0;
	wire w_dff_A_6oNImClC8_0;
	wire w_dff_A_NXl4ivyk3_0;
	wire w_dff_A_YobG7PX29_0;
	wire w_dff_A_7i5c9rVa5_0;
	wire w_dff_A_yHeClDfL7_0;
	wire w_dff_A_o4Y9rtJm4_0;
	wire w_dff_A_YCjAZHWK0_0;
	wire w_dff_A_LdsCSEZI6_0;
	wire w_dff_A_ChRngGDO9_0;
	wire w_dff_A_TiAQk5Re1_0;
	wire w_dff_A_zj7SLwyd6_1;
	wire w_dff_A_MlWFf3bL3_1;
	wire w_dff_A_GDrDJWA68_1;
	wire w_dff_A_X7uxLpvT9_1;
	wire w_dff_A_ZdNri9a43_1;
	wire w_dff_A_H3PqiOfo1_1;
	wire w_dff_A_Jie2WfFc5_1;
	wire w_dff_A_kUwnmmrZ7_1;
	wire w_dff_A_FETIMacw5_1;
	wire w_dff_A_WQ1bN8qa7_1;
	wire w_dff_A_otMMfgfO8_1;
	wire w_dff_A_3EpVKPhz5_1;
	wire w_dff_A_cMoJ2o695_1;
	wire w_dff_A_AzeBjmfW0_1;
	wire w_dff_A_0USWjrUG2_1;
	wire w_dff_A_oZZG3HHc4_1;
	wire w_dff_A_WWeEPOPW1_1;
	wire w_dff_A_3uhekAjo8_1;
	wire w_dff_A_0tZXxpk23_1;
	wire w_dff_A_tugRnaRv1_1;
	wire w_dff_A_oPtuWTSr1_1;
	wire w_dff_A_VRBojeX93_1;
	wire w_dff_A_B6w6EnVH3_1;
	wire w_dff_A_yM4DEeYD2_1;
	wire w_dff_A_2l8Hn0jK5_1;
	wire w_dff_A_r9l106aC1_0;
	wire w_dff_B_HbZ2tRBn8_1;
	wire w_dff_B_GJyJzrYg5_0;
	wire w_dff_B_m6mt5lgo3_0;
	wire w_dff_B_FnDaVBy43_0;
	wire w_dff_B_nWFepMSS1_0;
	wire w_dff_B_ApGIYt5O2_0;
	wire w_dff_B_M5crVnnZ1_0;
	wire w_dff_B_2ZzevI7Z5_0;
	wire w_dff_B_6RlGO1el5_0;
	wire w_dff_B_g6NpZbtg4_0;
	wire w_dff_B_9LYSI1eH6_0;
	wire w_dff_B_zfiVbqXR4_0;
	wire w_dff_B_jkxPcBk06_0;
	wire w_dff_B_R0XxsxpC1_0;
	wire w_dff_B_VX0yxNuR9_0;
	wire w_dff_B_eWTdcCEz0_0;
	wire w_dff_B_8XoYZ3G05_1;
	wire w_dff_B_Z3t2a2eE8_1;
	wire w_dff_B_6Zgzeqpj6_1;
	wire w_dff_B_GjLlNvMz7_1;
	wire w_dff_B_h1ZxgAE56_1;
	wire w_dff_B_1i38jL5G9_1;
	wire w_dff_B_pEMQrzCV0_1;
	wire w_dff_B_Dc1teHUy7_1;
	wire w_dff_B_ms8W2Lke6_1;
	wire w_dff_B_IOZhVMyW2_0;
	wire w_dff_B_MVmd3Uho4_0;
	wire w_dff_B_9w95WRaS0_0;
	wire w_dff_B_mxzQYyCT8_0;
	wire w_dff_B_cqhd36od9_0;
	wire w_dff_B_y6Vqf3g16_0;
	wire w_dff_B_jTIuBr0a9_0;
	wire w_dff_B_Ie3G75Ik7_0;
	wire w_dff_B_yfineotg2_1;
	wire w_dff_B_o3f2Divt9_1;
	wire w_dff_B_ZsBPbCzM7_1;
	wire w_dff_B_EHAmpLNC1_0;
	wire w_dff_B_NNe1iWJ31_0;
	wire w_dff_B_8nbF8iv83_0;
	wire w_dff_B_0VEg4nU59_0;
	wire w_dff_B_401L7AbP2_1;
	wire w_dff_B_Of5oisTA5_1;
	wire w_dff_B_DyzEanKZ7_0;
	wire w_dff_B_llo0HSNX3_1;
	wire w_dff_B_UbgWf2mq6_1;
	wire w_dff_B_SYxa1nNY0_1;
	wire w_dff_B_4Ks4C6Wa7_1;
	wire w_dff_B_rOBnvl9s1_1;
	wire w_dff_B_zOJ8wkxH1_1;
	wire w_dff_B_erZgD98O7_1;
	wire w_dff_B_BPeRjwXy5_1;
	wire w_dff_B_nl3pMGxk3_0;
	wire w_dff_B_xmWiSD9n9_0;
	wire w_dff_B_VUrcezlU8_0;
	wire w_dff_B_poS95E5R3_0;
	wire w_dff_B_cgxjWMuI9_1;
	wire w_dff_B_ES2YB4tC6_1;
	wire w_dff_B_BcRE7Wck8_1;
	wire w_dff_B_ZPHCc3s71_1;
	wire w_dff_B_0Wh4mUwg8_1;
	wire w_dff_A_t7KsM1fg9_1;
	wire w_dff_A_iyAYWHzH5_1;
	wire w_dff_A_jGO7FZbT7_1;
	wire w_dff_A_SlwfD1su5_1;
	wire w_dff_A_gu9V6RPw5_1;
	wire w_dff_A_0jptbRSB0_0;
	wire w_dff_B_FalOaTVm9_1;
	wire w_dff_B_LmEkCVDf8_1;
	wire w_dff_B_MIstKFXz0_1;
	wire w_dff_B_PpII1eyy4_1;
	wire w_dff_B_P9jroFVj2_1;
	wire w_dff_B_JsDsytI55_1;
	wire w_dff_A_SJmOnuzi0_1;
	wire w_dff_A_8L0DwhXT3_1;
	wire w_dff_A_hXcPV68U0_1;
	wire w_dff_B_9BqoDOAJ9_0;
	wire w_dff_B_0MIFE1Bw3_0;
	wire w_dff_B_nlp9xfky9_0;
	wire w_dff_B_s2xF01Tw8_0;
	wire w_dff_B_x53bLicH9_0;
	wire w_dff_B_7K6smtvZ2_0;
	wire w_dff_B_hlrUaGM92_0;
	wire w_dff_B_A1m94hoT3_0;
	wire w_dff_A_eiLXe4z73_0;
	wire w_dff_A_VyKc0K8E5_0;
	wire w_dff_A_ErRjlPQp7_1;
	wire w_dff_A_d0PiL9Ll8_1;
	wire w_dff_B_zF4bDGEv2_0;
	wire w_dff_B_yo14BoqS2_0;
	wire w_dff_B_9n6A3Gqv3_0;
	wire w_dff_B_752wZbhv8_0;
	wire w_dff_B_tlh8MtPP5_0;
	wire w_dff_B_81nv7xqY1_0;
	wire w_dff_B_fHRJB02K1_0;
	wire w_dff_B_ZHxKTDeG8_0;
	wire w_dff_B_y7op2Qz88_0;
	wire w_dff_B_tXmdT7kn9_0;
	wire w_dff_B_tM3qn2Od9_0;
	wire w_dff_B_k4bCUjyl2_1;
	wire w_dff_B_kvLmbFC01_1;
	wire w_dff_B_KHdMP5A09_1;
	wire w_dff_B_v6lCpZNv0_1;
	wire w_dff_B_sHvM5Zr10_1;
	wire w_dff_B_ksxvGuGo3_0;
	wire w_dff_B_p51TAtIC9_1;
	wire w_dff_B_W72VKEnG4_1;
	wire w_dff_B_cJrdyOfY6_1;
	wire w_dff_B_AGdyaDFT8_1;
	wire w_dff_B_t1VZo9LU6_1;
	wire w_dff_B_deyEznqR1_0;
	wire w_dff_A_zYWUnwFe9_1;
	wire w_dff_B_z6jI8JOq8_2;
	wire w_dff_B_xzqu5O5B4_2;
	wire w_dff_B_KScad4zf5_2;
	wire w_dff_A_cVaFdaMv6_1;
	wire w_dff_A_5CpDEeKf6_1;
	wire w_dff_A_eiKxvlwp6_0;
	wire w_dff_A_GonUom6y9_1;
	wire w_dff_A_4S7ROmRl3_1;
	wire w_dff_A_FYu6yqkl2_1;
	wire w_dff_A_um81YCu52_0;
	wire w_dff_B_6DSs9HIL1_0;
	wire w_dff_B_EcZ0iLGm0_0;
	wire w_dff_B_SMxFCpd09_0;
	wire w_dff_B_hlRPCz2F6_0;
	wire w_dff_A_WKicSeMw9_2;
	wire w_dff_A_S7H7Geem3_2;
	wire w_dff_A_DxjuNRJs4_1;
	wire w_dff_B_CR3BjyFH6_1;
	wire w_dff_B_ZOIj791h4_1;
	wire w_dff_B_PLRJ6Etj9_1;
	wire w_dff_B_lEZiYtB29_1;
	wire w_dff_B_oBSGK8As4_1;
	wire w_dff_A_CngO7eVm1_0;
	wire w_dff_A_qKqgdtiq5_0;
	wire w_dff_A_Z6o3NE1T2_1;
	wire w_dff_B_eB3cxISy9_0;
	wire w_dff_B_oI9jQJTi4_0;
	wire w_dff_B_tikuyAyg4_0;
	wire w_dff_B_5nXq0wmB1_0;
	wire w_dff_B_33rMplyV5_0;
	wire w_dff_B_iMrcfwYr1_0;
	wire w_dff_B_6sQkVDE55_0;
	wire w_dff_B_Qr37CMcf9_0;
	wire w_dff_B_yRhTEGI11_1;
	wire w_dff_B_K02sLONx8_1;
	wire w_dff_B_s7OrRFQo7_0;
	wire w_dff_A_nM5IVhfx6_2;
	wire w_dff_B_Bm1gAG0j2_2;
	wire w_dff_B_R0hu89kZ0_1;
	wire w_dff_B_Ir9qfCf96_1;
	wire w_dff_B_gXHOsSIl6_1;
	wire w_dff_B_X01pjMDj1_1;
	wire w_dff_B_GlulZvDF5_0;
	wire w_dff_A_fBl11jYt5_0;
	wire w_dff_A_7O4GBKmN5_2;
	wire w_dff_A_zHTm3kUb4_1;
	wire w_dff_A_4DfnUYM06_1;
	wire w_dff_A_BQrbGPB64_1;
	wire w_dff_A_b9LAaO2V4_1;
	wire w_dff_A_1ReQ3rI60_2;
	wire w_dff_A_sRJo8vKp0_2;
	wire w_dff_A_c6IZV7De9_2;
	wire w_dff_A_o4VBRHSQ5_2;
	wire w_dff_B_p93FT1pd2_0;
	wire w_dff_A_ESKtCnJ84_1;
	wire w_dff_B_DvXIxyGf4_1;
	wire w_dff_B_0qytQobt8_1;
	wire w_dff_B_Sa8S6l657_1;
	wire w_dff_B_LXJkArUv7_0;
	wire w_dff_B_3BYFU6wk9_1;
	wire w_dff_B_5wy3jEUG6_0;
	wire w_dff_A_tkWQIFCO0_0;
	wire w_dff_A_KXPvJ4ay2_0;
	wire w_dff_A_dYboeQ0R9_0;
	wire w_dff_B_3E3bFULf8_1;
	wire w_dff_B_mkW20p8i4_1;
	wire w_dff_B_hyFfmExd2_1;
	wire w_dff_B_O7F5IWIJ2_1;
	wire w_dff_B_9yN6e0JT4_1;
	wire w_dff_B_enNp6FUD9_1;
	wire w_dff_B_wBvIRgVB2_0;
	wire w_dff_B_i61UwHm20_0;
	wire w_dff_B_XYbubFso9_1;
	wire w_dff_B_lULTa84t5_1;
	wire w_dff_B_xGC1GvKU7_1;
	wire w_dff_B_21piD6Tr0_1;
	wire w_dff_B_RDsmvoLr7_1;
	wire w_dff_B_cj0UxHTU6_1;
	wire w_dff_A_oKGk8L4T6_1;
	wire w_dff_A_yC7bLEO03_1;
	wire w_dff_A_dDvpsJed7_2;
	wire w_dff_A_eTrHz4jv8_2;
	wire w_dff_B_2BHfzlba9_0;
	wire w_dff_B_0fop6hgz9_0;
	wire w_dff_B_R8jO07tz9_0;
	wire w_dff_B_oPHEf5Ne0_0;
	wire w_dff_A_gSZHdEuL1_1;
	wire w_dff_A_5IFVUyto1_1;
	wire w_dff_A_uXJjowcO9_2;
	wire w_dff_A_6Uj6uu5l7_2;
	wire w_dff_B_7uHF89Yi2_1;
	wire w_dff_B_OGNkaMNl4_1;
	wire w_dff_B_wzSXzrlF4_1;
	wire w_dff_B_pAxHbsCu2_0;
	wire w_dff_B_Aj2D0Oer9_0;
	wire w_dff_B_8eWT5FLm1_0;
	wire w_dff_B_UMGtMZK97_0;
	wire w_dff_B_dCLelrxZ8_0;
	wire w_dff_B_qBCX1vVK1_0;
	wire w_dff_B_WX1OM9gd9_1;
	wire w_dff_B_xoQRnqys4_1;
	wire w_dff_B_kFkvmHd54_0;
	wire w_dff_A_R8JEbloF5_0;
	wire w_dff_B_kUtKdGEd3_1;
	wire w_dff_B_8Mwsvgde1_1;
	wire w_dff_B_fgFE3RpO0_1;
	wire w_dff_B_L0ZsuJQK0_1;
	wire w_dff_B_9AAzravt8_1;
	wire w_dff_B_1vTMB9525_1;
	wire w_dff_B_gaXse5MV6_1;
	wire w_dff_B_PnW7Xyv40_1;
	wire w_dff_B_Ndnd0jB51_1;
	wire w_dff_B_yM0ra25v9_1;
	wire w_dff_B_AHrNX2v01_1;
	wire w_dff_B_KHWzBYxD2_1;
	wire w_dff_B_oPSouTSc8_1;
	wire w_dff_B_GKEavJx33_1;
	wire w_dff_B_AFA9y1HW5_0;
	wire w_dff_A_8nC7ayYu1_2;
	wire w_dff_A_pZGfTmqq0_0;
	wire w_dff_A_GPNj94e26_0;
	wire w_dff_A_Wsg0HdUG1_0;
	wire w_dff_A_ETicKf2s9_0;
	wire w_dff_B_GTkGHyzu7_0;
	wire w_dff_B_t8wk4rsF8_0;
	wire w_dff_A_i3FCZTXW0_0;
	wire w_dff_B_YUHFmixx5_0;
	wire w_dff_B_U9NVKsvB8_0;
	wire w_dff_B_Lcvoh0Hp3_0;
	wire w_dff_B_v8COqiHe8_0;
	wire w_dff_B_GFBcvfg54_0;
	wire w_dff_B_GmrysAj40_1;
	wire w_dff_B_MUofsgPe6_1;
	wire w_dff_B_BDtRMv4D3_1;
	wire w_dff_B_c9gsHbY27_1;
	wire w_dff_B_9szqQOzh1_1;
	wire w_dff_A_zyINY7Mr6_1;
	wire w_dff_A_pt9RtHEF4_1;
	wire w_dff_B_tZwGx5NQ2_1;
	wire w_dff_B_snBJIKE72_1;
	wire w_dff_B_T0JGSakf5_1;
	wire w_dff_B_m1toFi2Z4_1;
	wire w_dff_B_w8ZFtNkY0_1;
	wire w_dff_A_h0HBtqJs8_0;
	wire w_dff_A_1Rn6NAIO0_1;
	wire w_dff_A_zKbeWLTF1_1;
	wire w_dff_A_6c3adLdN9_1;
	wire w_dff_A_UxMnkg5s0_2;
	wire w_dff_A_hQjLbY4h4_2;
	wire w_dff_A_enpvF3rt7_2;
	wire w_dff_A_JUOYulXY2_2;
	wire w_dff_A_iF5cVrWG1_1;
	wire w_dff_B_qmhAqa5p4_0;
	wire w_dff_A_3nb9wQt70_0;
	wire w_dff_A_SLHqwUK49_0;
	wire w_dff_A_tqFOGh5y3_2;
	wire w_dff_A_gfeH5r0M2_2;
	wire w_dff_B_7xFu4Mi80_1;
	wire w_dff_B_1ecaiyHG9_1;
	wire w_dff_B_rwqpw1ea0_0;
	wire w_dff_B_eC3jd1QQ4_0;
	wire w_dff_A_Mokb2Ozp2_1;
	wire w_dff_A_wPCjnRXx0_2;
	wire w_dff_B_dxEGLWIz7_1;
	wire w_dff_B_xN7FYkZb6_0;
	wire w_dff_A_5d8bTIn96_0;
	wire w_dff_A_WFItt2iM5_1;
	wire w_dff_A_xeZgGkv54_1;
	wire w_dff_B_YfXokUhJ7_1;
	wire w_dff_B_J8ntFLjC9_1;
	wire w_dff_A_bJUmiIhN1_0;
	wire w_dff_A_DJibnqLW6_0;
	wire w_dff_A_vSvLhwb24_0;
	wire w_dff_A_DKsOg8qe2_0;
	wire w_dff_A_hhZyU8L87_0;
	wire w_dff_A_jQ3tBIKF0_1;
	wire w_dff_B_nXU4JbEZ0_0;
	wire w_dff_B_Po7JYX890_0;
	wire w_dff_B_PYgns8GG8_2;
	wire w_dff_B_ce4VxpCZ8_2;
	wire w_dff_A_YBcPvg7h7_0;
	wire w_dff_A_yv4guX720_0;
	wire w_dff_A_lE3ItQU19_0;
	wire w_dff_B_OPDiObkS2_0;
	wire w_dff_B_B7tUwYuz5_0;
	wire w_dff_B_1XT9siGY6_0;
	wire w_dff_B_9ylm8g6g4_0;
	wire w_dff_B_7n2j4Y9q1_1;
	wire w_dff_B_ni6NVzVi8_1;
	wire w_dff_B_WhCIUObC5_2;
	wire w_dff_B_ydfoAbKT5_1;
	wire w_dff_B_LvqtFccj9_1;
	wire w_dff_B_0eotRJax5_0;
	wire w_dff_A_H2vgC6kq4_1;
	wire w_dff_A_rukccQz65_1;
	wire w_dff_A_z8l9MxUk1_1;
	wire w_dff_A_kcV6abiy0_2;
	wire w_dff_A_q1KqtH6B0_2;
	wire w_dff_A_7ujfS0FO3_2;
	wire w_dff_B_hhfAUHHD0_1;
	wire w_dff_B_zPnQWszI8_1;
	wire w_dff_B_KVHLBWXp4_1;
	wire w_dff_B_vOi2AvAE7_1;
	wire w_dff_B_x8aIJJoV5_1;
	wire w_dff_B_KEhFo1TO7_1;
	wire w_dff_B_3b1YSCjC9_0;
	wire w_dff_B_28z0T09I2_1;
	wire w_dff_B_grn3rGDj5_1;
	wire w_dff_B_R2fQozyq6_0;
	wire w_dff_A_ph7TJQJV6_0;
	wire w_dff_B_3ps9KR4y8_3;
	wire w_dff_B_CKqL7Gir9_3;
	wire w_dff_B_CDR6Suz05_3;
	wire w_dff_A_yyHutWcL6_0;
	wire w_dff_B_ndqBDG7m5_2;
	wire w_dff_B_wb4jpeK49_2;
	wire w_dff_B_P0A9yaRt5_2;
	wire w_dff_B_ueObpH249_0;
	wire w_dff_B_jKyiDPet0_1;
	wire w_dff_B_mCyouFB74_1;
	wire w_dff_B_ogfKhUUA1_1;
	wire w_dff_B_X6hvEvIb3_1;
	wire w_dff_A_85JoKlax6_1;
	wire w_dff_A_Dv6O1XCu5_1;
	wire w_dff_A_tblrHz7F0_1;
	wire w_dff_A_9hkqwx6q6_2;
	wire w_dff_A_kXzz8afe8_2;
	wire w_dff_B_P6h9LSyK6_1;
	wire w_dff_B_iv6e9eD24_0;
	wire w_dff_A_vhYSnYkN0_0;
	wire w_dff_B_u7mi6eWz7_3;
	wire w_dff_B_2nFbqOQB2_3;
	wire w_dff_B_Y4As0ua57_3;
	wire w_dff_A_MvBFLSK72_1;
	wire w_dff_A_h7TBsyZ56_1;
	wire w_dff_A_ShlU2W4v1_1;
	wire w_dff_A_cHxiyPDX9_1;
	wire w_dff_A_liyqeJHw8_1;
	wire w_dff_A_4sp08cSE4_1;
	wire w_dff_A_tgRMtliv9_1;
	wire w_dff_A_Jnrfl8BP3_1;
	wire w_dff_A_ljCR1h082_0;
	wire w_dff_A_cX0ulFsR7_0;
	wire w_dff_A_9W79FXkf7_0;
	wire w_dff_A_dMNaZEgX4_0;
	wire w_dff_A_PuiCmZd40_0;
	wire w_dff_A_v1azH6f15_0;
	wire w_dff_A_SYZxXsO99_0;
	wire w_dff_A_rLgAvqL93_0;
	wire w_dff_A_vrwR2ugt4_0;
	wire w_dff_A_oZzRsgcd3_0;
	wire w_dff_A_UK7zN0hx1_0;
	wire w_dff_A_xEbno4Bc2_2;
	wire w_dff_A_cKNOEeHX5_2;
	wire w_dff_A_tOdF6zHU2_2;
	wire w_dff_A_8DEhp2Yc7_2;
	wire w_dff_A_RaGEzzcA5_2;
	wire w_dff_A_6oFbUtcT3_2;
	wire w_dff_A_I8RgdFMX2_2;
	wire w_dff_A_sRVzXlW13_2;
	wire w_dff_A_bkxMkfld2_2;
	wire w_dff_A_HqH1KDj88_2;
	wire w_dff_A_JRZ2oKPU4_2;
	wire w_dff_A_z5QvvfQZ2_1;
	wire w_dff_A_KQa0EXTd1_1;
	wire w_dff_A_05YmZwlX5_1;
	wire w_dff_A_S88yINAh8_1;
	wire w_dff_A_1ametKsg4_1;
	wire w_dff_A_ceTfrecR8_1;
	wire w_dff_A_VzSK2nFp8_1;
	wire w_dff_A_UMGNIApm0_1;
	wire w_dff_A_3k9j5T8S9_1;
	wire w_dff_A_n0HXTEJQ5_1;
	wire w_dff_A_mquicPis4_1;
	wire w_dff_A_iu21Zqse8_2;
	wire w_dff_A_bNb2Uc5A9_2;
	wire w_dff_A_Mho3DNf74_2;
	wire w_dff_A_CWuBi4A70_2;
	wire w_dff_A_fYj21vvD2_2;
	wire w_dff_A_2Yj3U0Ip8_2;
	wire w_dff_A_fETiwb8L9_2;
	wire w_dff_A_424xl1M53_2;
	wire w_dff_A_Axf6eWiB8_2;
	wire w_dff_A_e4gAfepL0_2;
	wire w_dff_A_cVKG9rir9_2;
	wire w_dff_B_pfinCzPT2_0;
	wire w_dff_B_6MOx5bXI0_0;
	wire w_dff_B_GlnTseJ03_0;
	wire w_dff_B_ub5IZ7f08_0;
	wire w_dff_B_hlze2NKO0_0;
	wire w_dff_A_5C6bK9Er7_0;
	wire w_dff_A_Mr9KwjKC5_0;
	wire w_dff_A_qLDdam202_1;
	wire w_dff_A_Q4wI0UC29_1;
	wire w_dff_A_VCWSou9t2_1;
	wire w_dff_A_W2tZn6oo0_2;
	wire w_dff_A_vZavnI3J3_2;
	wire w_dff_A_21XGM9dY5_2;
	wire w_dff_B_DVg5wLGo7_2;
	wire w_dff_B_od8OPG3C2_2;
	wire w_dff_B_XuZ320K68_2;
	wire w_dff_B_qi5F0OtT9_2;
	wire w_dff_B_E8dVdOKK3_2;
	wire w_dff_B_GUthqoH39_2;
	wire w_dff_B_kv6xiJAF2_2;
	wire w_dff_B_4b2PzjOD8_2;
	wire w_dff_B_MXXFSrIR7_2;
	wire w_dff_B_awJynNY93_2;
	wire w_dff_B_lKGVZogW8_2;
	wire w_dff_B_prryET5Y2_2;
	wire w_dff_B_ixLNvbGt5_2;
	wire w_dff_A_h6FWygUN2_1;
	wire w_dff_B_db7XWevs2_0;
	wire w_dff_B_S5C3hmwv6_0;
	wire w_dff_B_9KNlN64E5_0;
	wire w_dff_B_grSwZci18_0;
	wire w_dff_B_YFXLITn83_0;
	wire w_dff_B_c0lgAy7I6_0;
	wire w_dff_B_OnyCKrrI0_0;
	wire w_dff_B_Vmqt1nVN1_0;
	wire w_dff_B_emuLrLSO1_0;
	wire w_dff_B_G2gKboAY4_0;
	wire w_dff_B_ZCKLYel97_0;
	wire w_dff_B_T7YRSEFI8_1;
	wire w_dff_B_nFwzypT18_1;
	wire w_dff_B_OlxLIZKe6_1;
	wire w_dff_B_yCLnCPdg4_1;
	wire w_dff_A_HHcohrtA2_1;
	wire w_dff_A_PhMWxTnj9_1;
	wire w_dff_A_0IN0JfWw8_2;
	wire w_dff_A_kFX52wfa6_1;
	wire w_dff_A_qOiP1xr63_1;
	wire w_dff_A_NlxxDMZS6_1;
	wire w_dff_A_2qfylIWC6_1;
	wire w_dff_A_FaEIrqfd4_2;
	wire w_dff_A_RZ9Ybcvo7_2;
	wire w_dff_A_ai5X3qVU2_2;
	wire w_dff_A_k3RzfDcU5_2;
	wire w_dff_A_aX2enYOS0_1;
	wire w_dff_A_bMRvYAOp3_0;
	wire w_dff_A_VOzgwAf71_0;
	wire w_dff_A_f5eZqiSk3_0;
	wire w_dff_A_7dahFntp7_0;
	wire w_dff_A_hCdCIPgc2_2;
	wire w_dff_A_4mN2gque2_2;
	wire w_dff_A_dzJCSBPn5_2;
	wire w_dff_A_FGQPDyVV7_1;
	wire w_dff_B_QIWtjCoA8_1;
	wire w_dff_B_NeUMlFJp7_1;
	wire w_dff_B_3i5y8pxZ4_1;
	wire w_dff_B_Pd0enkjG3_0;
	wire w_dff_A_hNX5uZgb5_1;
	wire w_dff_A_57GtZJ4n5_2;
	wire w_dff_A_rM240p1f9_0;
	wire w_dff_B_LpsyiCaf0_3;
	wire w_dff_B_MfiL7xzF9_3;
	wire w_dff_B_0VZex3Hm5_3;
	wire w_dff_B_HEvNRcaN0_1;
	wire w_dff_B_7KXg4KOM0_0;
	wire w_dff_A_oB6lzMDA6_0;
	wire w_dff_A_j4Uv2WQa9_1;
	wire w_dff_A_hepERO6O0_1;
	wire w_dff_A_EQNe65gU1_1;
	wire w_dff_A_6nr5mi6s0_1;
	wire w_dff_A_An8P9YTY1_1;
	wire w_dff_A_FMuJZgSB0_1;
	wire w_dff_A_AJINMCdz2_1;
	wire w_dff_A_O8ofyVi79_1;
	wire w_dff_A_lNLgv9sO2_2;
	wire w_dff_A_znYIGwJu5_2;
	wire w_dff_B_dfYfCtd01_0;
	wire w_dff_B_HDbb506a3_0;
	wire w_dff_B_JEGIYvPq9_0;
	wire w_dff_B_2SXwo92r8_0;
	wire w_dff_A_fk5jWGnA9_0;
	wire w_dff_B_q0aTz60I1_0;
	wire w_dff_B_dOt1Tn671_0;
	wire w_dff_B_aX6P7Wmo8_0;
	wire w_dff_B_Rk8nBEIU8_0;
	wire w_dff_B_LnzMSa2X5_0;
	wire w_dff_A_SAJ9ZYRz3_2;
	wire w_dff_A_sX2QTqjo1_1;
	wire w_dff_A_08DYid1T7_1;
	wire w_dff_A_rUG6UDsZ7_2;
	wire w_dff_A_54pKiNtS3_2;
	wire w_dff_A_tzrtAI7m3_0;
	wire w_dff_A_K7dgk8tN8_1;
	wire w_dff_A_VGFuQtq12_1;
	wire w_dff_A_iLZMufHi7_1;
	wire w_dff_A_jdrnQAet0_1;
	wire w_dff_B_RWpjDFmZ9_1;
	wire w_dff_B_zINCodE96_1;
	wire w_dff_A_Omws4HRf0_1;
	wire w_dff_B_ofPosrps6_1;
	wire w_dff_B_GJ14VP5H9_0;
	wire w_dff_B_zFyNKBy09_0;
	wire w_dff_B_aqhacGvo0_0;
	wire w_dff_B_gnYSGXxX9_1;
	wire w_dff_A_QYJ1XEN48_0;
	wire w_dff_A_xhqleR399_0;
	wire w_dff_B_Z9DRwtjf7_1;
	wire w_dff_B_29U80Tha0_1;
	wire w_dff_A_Svx1ceIm9_0;
	wire w_dff_A_mDKt5XaW3_0;
	wire w_dff_B_ynRXNWFL6_0;
	wire w_dff_B_x12Dlwfq6_1;
	wire w_dff_B_kOs3fhSF4_1;
	wire w_dff_B_slMstrte5_1;
	wire w_dff_B_cshKiaOQ2_1;
	wire w_dff_B_zxbaoMfp4_0;
	wire w_dff_B_yOxgi82s2_0;
	wire w_dff_B_VmG7eHiP2_1;
	wire w_dff_B_EPNAo89L3_1;
	wire w_dff_B_B7COo6eY8_1;
	wire w_dff_A_ungVqv2X1_1;
	wire w_dff_A_C0LML8KC2_1;
	wire w_dff_B_d35W7zc98_1;
	wire w_dff_B_zWcwDe4Y2_1;
	wire w_dff_A_lWlnWEgN4_0;
	wire w_dff_A_Dqkbk04K2_0;
	wire w_dff_A_8FXxH05R3_0;
	wire w_dff_A_umKsocQE8_0;
	wire w_dff_B_npcdkGxv1_0;
	wire w_dff_A_eQgjJxiJ5_1;
	wire w_dff_A_DGM43qRJ8_1;
	wire w_dff_A_kTJVhsh78_2;
	wire w_dff_A_Mec99Jkt8_2;
	wire w_dff_A_KhBqDzzW3_2;
	wire w_dff_A_fJlaCSEw5_2;
	wire w_dff_B_0Azvf9Fl7_1;
	wire w_dff_B_ITbc963N6_1;
	wire w_dff_B_PRok0oYL4_1;
	wire w_dff_A_cpviNkYV1_0;
	wire w_dff_B_Qrej3fvK6_2;
	wire w_dff_A_DYWWZoxZ8_1;
	wire w_dff_A_PqId0mA34_1;
	wire w_dff_A_hIXBk1Sm1_1;
	wire w_dff_B_jhsR9Bgj6_2;
	wire w_dff_B_fru2YtIE1_2;
	wire w_dff_B_yiDorP7l7_1;
	wire w_dff_B_OSnglj877_1;
	wire w_dff_B_Mpdsynv86_1;
	wire w_dff_B_Ar0CnoHU5_0;
	wire w_dff_B_F9tTvFqz1_0;
	wire w_dff_A_bHunUFF88_2;
	wire w_dff_B_pHiKbyQ42_1;
	wire w_dff_B_dCHAiDYb7_1;
	wire w_dff_B_E8v5SAeS1_1;
	wire w_dff_A_PgdpENDr5_1;
	wire w_dff_A_9nFqy9n97_1;
	wire w_dff_A_H77SgCYr7_1;
	wire w_dff_A_64sbxD039_2;
	wire w_dff_A_FqNKuP124_2;
	wire w_dff_A_6WVgIdG06_2;
	wire w_dff_A_OvbUSvio9_2;
	wire w_dff_A_kxpL3vxm7_1;
	wire w_dff_A_4KT7QmGz5_1;
	wire w_dff_A_3idra0BX3_1;
	wire w_dff_A_CuR1NTLR6_2;
	wire w_dff_A_cHL9pHTy1_2;
	wire w_dff_A_IS82ssZ56_0;
	wire w_dff_A_vmV6BBVp7_0;
	wire w_dff_A_w6X8EAcp6_2;
	wire w_dff_A_6x8J0fqr0_2;
	wire w_dff_A_kUor1Urz2_2;
	wire w_dff_A_3meGaPFs8_2;
	wire w_dff_A_IMqtcTZr3_1;
	wire w_dff_A_kNeAsqV88_1;
	wire w_dff_A_RNGblkSf3_1;
	wire w_dff_A_LlrkQsaX4_0;
	wire w_dff_A_fRSggduI5_0;
	wire w_dff_A_uDnNAuvx7_1;
	wire w_dff_A_cO4jwKc07_0;
	wire w_dff_A_bX5NXgyS0_2;
	wire w_dff_A_uVQZlh898_2;
	wire w_dff_A_Np93gKq95_2;
	wire w_dff_A_k3YJBcmu3_2;
	wire w_dff_A_IMewhTWL3_0;
	wire w_dff_A_4vDcmayi0_0;
	wire w_dff_A_4WlSrDkw0_0;
	wire w_dff_A_nU0xe2hO8_0;
	wire w_dff_B_nz0k8Dpq6_0;
	wire w_dff_B_8OUHYnjW1_0;
	wire w_dff_B_zcaO3fTP5_0;
	wire w_dff_B_Jm8RHGg78_0;
	wire w_dff_B_pEm7TDq81_0;
	wire w_dff_B_dbbEQrdT0_0;
	wire w_dff_B_RMjq1yaJ2_0;
	wire w_dff_B_Df4TBVsa6_0;
	wire w_dff_B_zCZBW35C3_0;
	wire w_dff_A_UnD3muEz2_2;
	wire w_dff_A_7DsqpNYG0_2;
	wire w_dff_A_IwS5gG914_2;
	wire w_dff_A_GF8jmkDA1_2;
	wire w_dff_A_3EaRjSST1_2;
	wire w_dff_A_V97YHEA45_2;
	wire w_dff_A_0ufxqKr63_2;
	wire w_dff_A_H2OdbD9J3_2;
	wire w_dff_A_Aahst3tl4_0;
	wire w_dff_A_Lz1zNJb54_0;
	wire w_dff_A_kwqkkcbr4_0;
	wire w_dff_A_id0GhgZb4_0;
	wire w_dff_B_NU8ATwn54_1;
	wire w_dff_B_C5aySXOr5_1;
	wire w_dff_B_yxqJN0WG9_1;
	wire w_dff_B_lcR5Qci74_1;
	wire w_dff_B_cWpeFl2z9_1;
	wire w_dff_B_NRsKYzsN1_0;
	wire w_dff_A_PhvWA9S78_0;
	wire w_dff_A_QSc45vXT9_0;
	wire w_dff_A_epaqPPby9_0;
	wire w_dff_A_ryAzrpiQ6_0;
	wire w_dff_A_1OmPXXXf3_2;
	wire w_dff_A_fd8aelqm7_2;
	wire w_dff_A_cjnYpDZZ3_0;
	wire w_dff_A_hOC88yrv1_2;
	wire w_dff_A_S7K7j6zJ5_2;
	wire w_dff_B_F3OXA4Xb4_1;
	wire w_dff_B_OhJl4kWT7_0;
	wire w_dff_A_XbIQ92Om5_1;
	wire w_dff_B_rwito7iL8_3;
	wire w_dff_B_1HeEAX3R0_3;
	wire w_dff_B_dHAKO5Ky6_3;
	wire w_dff_B_xjOizQFs3_1;
	wire w_dff_B_uc1cmXy18_1;
	wire w_dff_B_JdtGa10D5_1;
	wire w_dff_B_OWwWer5e5_1;
	wire w_dff_A_j6sSd1G47_1;
	wire w_dff_A_rPzBLQIM3_1;
	wire w_dff_A_3ljWBAJk4_1;
	wire w_dff_A_KzTG18MI1_2;
	wire w_dff_A_YLSKHkFy7_2;
	wire w_dff_A_qfTcccIv9_1;
	wire w_dff_B_QUDIr1v97_3;
	wire w_dff_B_KNh74oeF5_3;
	wire w_dff_B_Q4pTqb6Z2_3;
	wire w_dff_B_0Ak9n4Gf5_3;
	wire w_dff_B_ZT2Fy5OR0_3;
	wire w_dff_B_UfJBKIYt5_3;
	wire w_dff_A_D7VmnP0H6_0;
	wire w_dff_A_VyqhLvL34_1;
	wire w_dff_A_ag9PAe2Q7_1;
	wire w_dff_A_2ISeGub15_0;
	wire w_dff_A_pFsDiY7u2_0;
	wire w_dff_A_YFMzVTqr9_1;
	wire w_dff_B_wpdkgUXj5_3;
	wire w_dff_B_qEsBJxUD4_3;
	wire w_dff_A_5QsPzIWS9_1;
	wire w_dff_A_tbwDyGZi6_1;
	wire w_dff_A_I7En2C3i0_1;
	wire w_dff_A_RkLGsPvh1_1;
	wire w_dff_A_BzFwJUiJ7_1;
	wire w_dff_A_zBquLsHA5_2;
	wire w_dff_A_l9kBWW3d9_2;
	wire w_dff_A_G0SkIRPB5_2;
	wire w_dff_A_Nru9sjMX0_2;
	wire w_dff_A_O8MIMKtL8_2;
	wire w_dff_A_l2StL5735_0;
	wire w_dff_A_STYJgthL2_0;
	wire w_dff_A_ViKm35nZ0_0;
	wire w_dff_A_6xd4p2ig0_2;
	wire w_dff_A_YnW30gqB9_2;
	wire w_dff_A_VTa9wZt32_2;
	wire w_dff_A_O3QSvosB8_2;
	wire w_dff_A_E4shbBiG7_1;
	wire w_dff_A_Ul7sozB86_1;
	wire w_dff_A_ceiHMDiR8_1;
	wire w_dff_A_awF8wFPy0_0;
	wire w_dff_A_x1TuvTHU1_0;
	wire w_dff_A_Vskg1MDg6_0;
	wire w_dff_A_vodn5zpv1_0;
	wire w_dff_A_WTvG5u597_1;
	wire w_dff_A_J9nVbyfr6_1;
	wire w_dff_A_MDmMMSEI6_1;
	wire w_dff_A_nX47WIO03_1;
	wire w_dff_A_jyy5vK6a4_1;
	wire w_dff_B_qnbmHtnG0_1;
	wire w_dff_B_NxTT5afB0_0;
	wire w_dff_A_SJzdCyfz2_0;
	wire w_dff_A_Hf6WpMvU3_0;
	wire w_dff_A_NYg96YUV4_0;
	wire w_dff_A_2jGD6EWq2_0;
	wire w_dff_A_hsQkJUjs5_0;
	wire w_dff_A_99Lyr7EB8_0;
	wire w_dff_A_I1ysKMfU3_1;
	wire w_dff_A_WuVLOwsN2_1;
	wire w_dff_A_KeaK6sWc8_1;
	wire w_dff_A_0J2BOCin4_0;
	wire w_dff_A_NfVWJxMP8_1;
	wire w_dff_A_OFz0DY0G5_1;
	wire w_dff_A_IygjiqAm7_1;
	wire w_dff_A_DjwTDdgY0_1;
	wire w_dff_A_WbsNak8x0_1;
	wire w_dff_A_Sr2PvNhv5_1;
	wire w_dff_A_zfneC0I78_1;
	wire w_dff_A_nM2dE7mB2_1;
	wire w_dff_A_DgfAJj4N8_1;
	wire w_dff_A_wXWYsxiw2_2;
	wire w_dff_A_haOV4gqD4_2;
	wire w_dff_A_rWBDxUmw4_2;
	wire w_dff_A_EvvZ3X4i9_2;
	wire w_dff_A_rabhZ6A95_2;
	wire w_dff_A_GNYgQhL69_2;
	wire w_dff_A_9GwzyXxU8_2;
	wire w_dff_A_5A63NY9a2_0;
	wire w_dff_A_QYNBuYWH1_0;
	wire w_dff_A_uw12bGCa6_1;
	wire w_dff_A_aqXJWKtH7_1;
	wire w_dff_A_hzAYjnOD2_1;
	wire w_dff_B_qAclKrdA2_3;
	wire w_dff_B_w3b5geSx4_3;
	wire w_dff_B_Fqzti0kV8_3;
	wire w_dff_A_lntjXngU7_0;
	wire w_dff_A_yPEQ2pZA0_0;
	wire w_dff_A_HBZAUb3Z2_0;
	wire w_dff_A_0KOZ3ZLX5_0;
	wire w_dff_A_0I2AnvN35_0;
	wire w_dff_A_oY6PDkZN7_0;
	wire w_dff_A_fMPXNQTL7_0;
	wire w_dff_A_vMAkBAe16_0;
	wire w_dff_A_TD28eZi25_0;
	wire w_dff_A_nejF3chI5_2;
	wire w_dff_A_eG28GnkY8_2;
	wire w_dff_A_Ys3imqdp0_2;
	wire w_dff_A_m4UV112b5_2;
	wire w_dff_A_rXrpx5k01_2;
	wire w_dff_A_96vV0G517_2;
	wire w_dff_A_nQN5faLv3_2;
	wire w_dff_A_dnxCFmOJ2_2;
	wire w_dff_A_TJa5PZqy0_2;
	wire w_dff_A_tTKLcRNg1_1;
	wire w_dff_A_VX52WHcy1_1;
	wire w_dff_A_YxEwIlRF2_1;
	wire w_dff_A_hZhPsBRS8_1;
	wire w_dff_A_WyR0C5My1_1;
	wire w_dff_A_SKjdGmfI2_1;
	wire w_dff_A_xYUjHr2C0_1;
	wire w_dff_A_hgHfYdiD1_1;
	wire w_dff_A_uXbz31cQ1_1;
	wire w_dff_A_blrUEFU90_1;
	wire w_dff_A_jJGCuiG54_1;
	wire w_dff_A_rk3LxFqX6_1;
	wire w_dff_A_xTp5TZ9O0_1;
	wire w_dff_A_XzxTgkJR1_2;
	wire w_dff_A_maUJpcYL6_2;
	wire w_dff_A_Y2tVyCbG7_2;
	wire w_dff_A_p7w6alMI1_2;
	wire w_dff_A_6pStX4yu2_2;
	wire w_dff_A_fzJDj07o3_2;
	wire w_dff_A_CwmetvLJ4_0;
	wire w_dff_A_KMhfDZJK4_0;
	wire w_dff_A_xZOQaMZ18_0;
	wire w_dff_A_HIIdMCc72_0;
	wire w_dff_A_DmgrzdGC2_0;
	wire w_dff_A_4qaDxOO28_0;
	wire w_dff_A_NYjhC4kM6_0;
	wire w_dff_A_cMZDIVR50_0;
	wire w_dff_A_yhKvvx4i3_0;
	wire w_dff_A_aaG5i23a4_0;
	wire w_dff_A_OU3GV55K4_0;
	wire w_dff_A_f05HXOnv4_0;
	wire w_dff_A_2tBscZ9S4_0;
	wire w_dff_A_wY2BFypZ0_1;
	wire w_dff_A_dpp6i8I67_1;
	wire w_dff_A_IVvQ347e1_1;
	wire w_dff_A_cnVrDyCU7_1;
	wire w_dff_A_8IVjR0xI3_1;
	wire w_dff_A_3Jxab8y11_1;
	wire w_dff_A_uN7FRiqQ5_1;
	wire w_dff_A_gJrVJFWp4_1;
	wire w_dff_A_2YLmKrwW2_1;
	wire w_dff_A_woculaxd1_1;
	wire w_dff_A_BIxKP5jb2_1;
	wire w_dff_A_gmUxuLte6_1;
	wire w_dff_A_IVH6G14y3_1;
	wire w_dff_A_zULqCA694_1;
	wire w_dff_A_mOQ1Rf9X4_1;
	wire w_dff_A_wMf7uVbY8_1;
	wire w_dff_A_X5uEQ9JW1_1;
	wire w_dff_A_brqX0PSN0_1;
	wire w_dff_A_hzkHJ7Cn2_1;
	wire w_dff_A_zwsVJ1Jd6_1;
	wire w_dff_A_QUlRRTAD9_1;
	wire w_dff_A_5r2OHNgV7_1;
	wire w_dff_A_cOX1wknL5_1;
	wire w_dff_A_UBMxUog21_1;
	wire w_dff_A_SBlFO4oN4_1;
	wire w_dff_A_Nog6MXY70_1;
	wire w_dff_A_selQeCpb8_2;
	wire w_dff_A_ZGjm3VWB7_2;
	wire w_dff_A_wt1jgVp02_2;
	wire w_dff_A_dE4yIXIU6_2;
	wire w_dff_A_aSLQIEMQ7_2;
	wire w_dff_A_f8ZhtnEk9_2;
	wire w_dff_A_pZMcA2zf2_2;
	wire w_dff_A_hcHaolDj0_2;
	wire w_dff_A_3UsKYpRU8_2;
	wire w_dff_A_auz1LV600_2;
	wire w_dff_A_K8NbMXzY1_2;
	wire w_dff_A_4oGrtiqL7_2;
	wire w_dff_A_n6eLtSK16_2;
	wire w_dff_A_9Ris1djT8_0;
	wire w_dff_A_vAB9WeN85_0;
	wire w_dff_A_8oI67hMM8_0;
	wire w_dff_A_cRzoOTxt2_0;
	wire w_dff_A_3FWaDXEN4_1;
	wire w_dff_A_ch7PBlMN5_1;
	wire w_dff_B_nKnuInHT5_0;
	wire w_dff_A_HFB9aPQp9_0;
	wire w_dff_A_SYDBoXsz1_0;
	wire w_dff_A_Bg85DPP36_2;
	wire w_dff_A_qpTm1GQJ9_2;
	wire w_dff_A_SOoMbCl00_2;
	wire w_dff_A_jgbfN1vM5_2;
	wire w_dff_A_EP4rSHyd8_2;
	wire w_dff_A_Ismp3crw7_2;
	wire w_dff_A_ZNyGVDGL9_2;
	wire w_dff_A_nKyYHsfW0_2;
	wire w_dff_A_FtLvesBI1_0;
	wire w_dff_A_ZrQMDoap6_0;
	wire w_dff_A_bfes5KM11_2;
	wire w_dff_A_GCtHfPh14_2;
	wire w_dff_A_F4JM2YFm9_0;
	wire w_dff_A_K84degn92_0;
	wire w_dff_A_nKuWQFIl5_0;
	wire w_dff_A_OIHgNgxR0_0;
	wire w_dff_A_Y2A7gShM2_0;
	wire w_dff_A_b50Re8nB5_0;
	wire w_dff_A_e2VBHxhv5_0;
	wire w_dff_A_0KIsQ1mU5_0;
	wire w_dff_A_7oO9CIoC1_0;
	wire w_dff_A_RSzZWXVj4_0;
	wire w_dff_A_rWmU1MjV1_0;
	wire w_dff_A_k1NkJp7b0_0;
	wire w_dff_A_xtv4nyuw3_0;
	wire w_dff_A_YC8evA8F3_0;
	wire w_dff_A_Ok1a3AvL2_0;
	wire w_dff_A_R18cgiXf1_0;
	wire w_dff_A_4LeNu4Fx5_0;
	wire w_dff_A_goZeSfFy0_0;
	wire w_dff_A_7ufrZGyP7_0;
	wire w_dff_A_9zjWDTx27_0;
	wire w_dff_A_A3zbijFr1_0;
	wire w_dff_A_Rvoneyhf2_0;
	wire w_dff_A_sefXaNOh3_0;
	wire w_dff_A_7GWS8WTE9_0;
	wire w_dff_A_5a96gD1R9_0;
	wire w_dff_A_E57cqyLp5_2;
	wire w_dff_A_3djHRfyX3_2;
	wire w_dff_A_anl4YDs76_2;
	wire w_dff_A_Mfi644JQ0_2;
	wire w_dff_A_BKiHM41L6_2;
	wire w_dff_A_jwf3RqY31_2;
	wire w_dff_A_s0qAwI177_2;
	wire w_dff_A_shISe07W1_2;
	wire w_dff_A_timhTuNW9_2;
	wire w_dff_A_XgT1hNsl5_2;
	wire w_dff_A_6FBUvdrw1_2;
	wire w_dff_A_s6e0nStv1_2;
	wire w_dff_A_G1RDL8658_2;
	wire w_dff_A_XXvBEiAi5_0;
	wire w_dff_A_RDrg7y4S0_0;
	wire w_dff_A_f9Cpt51i1_0;
	wire w_dff_A_cPKpNQWS6_0;
	wire w_dff_A_7hcUo6Fw6_0;
	wire w_dff_A_4l2dCGDJ4_0;
	wire w_dff_A_DwmwnVAX6_0;
	wire w_dff_A_YoxkjmP48_0;
	wire w_dff_A_EOKouaho4_0;
	wire w_dff_A_PBhybKyN1_0;
	wire w_dff_A_ZvsNFf2l9_0;
	wire w_dff_A_5O6qQtgB8_0;
	wire w_dff_A_7cPgEucv5_0;
	wire w_dff_A_ixKVzI3j3_0;
	wire w_dff_A_6h4ZecNt6_0;
	wire w_dff_A_w0tPuwmj0_0;
	wire w_dff_A_8ZO8nfsg0_0;
	wire w_dff_A_5NHNfACy9_0;
	wire w_dff_A_G18Mxl004_0;
	wire w_dff_A_usf1N4f43_0;
	wire w_dff_A_KNfKET0q1_0;
	wire w_dff_A_kz1yxDR71_0;
	wire w_dff_A_LHxeaux42_0;
	wire w_dff_A_5sTCyrqc9_0;
	wire w_dff_A_FX7F36bV1_0;
	wire w_dff_A_aCotgp3k1_0;
	wire w_dff_A_hkReL28n0_0;
	wire w_dff_A_d30irgnH5_0;
	wire w_dff_A_rzjd6yL58_0;
	wire w_dff_A_XVsKrCdE7_0;
	wire w_dff_A_eFeoRqT64_2;
	wire w_dff_A_n66LXlKa5_2;
	wire w_dff_A_4tE8wuxC2_2;
	wire w_dff_A_7K543ZXj6_2;
	wire w_dff_A_ucrzRESH3_2;
	wire w_dff_A_7HADqwTF6_2;
	wire w_dff_A_8EGHPGrd4_2;
	wire w_dff_A_U3Hu6lUw8_2;
	wire w_dff_A_rkloMUJm8_2;
	wire w_dff_A_DxSbFAvt0_2;
	wire w_dff_A_ss6FeutD6_2;
	wire w_dff_A_dZdSFfP14_2;
	wire w_dff_A_VLQxYgqR3_2;
	wire w_dff_A_S7M87JQ34_2;
	wire w_dff_A_9bEojj280_2;
	wire w_dff_A_8uzhtFKJ3_2;
	wire w_dff_A_CpoKBqtE8_1;
	wire w_dff_A_p1EYyQHN3_1;
	wire w_dff_A_JLk0Odgx0_1;
	wire w_dff_A_YCOGnO5v7_1;
	wire w_dff_A_HFqTF5Yr7_1;
	wire w_dff_A_ZIn8C9WS7_1;
	wire w_dff_A_oisPxduo3_1;
	wire w_dff_A_VZRWOjUT8_1;
	wire w_dff_A_cMAy5yxu0_1;
	wire w_dff_A_f3400uJP9_1;
	wire w_dff_A_URtKe4Ir6_1;
	wire w_dff_A_SNlLy2Sr3_1;
	wire w_dff_A_Zj24YKqJ9_1;
	wire w_dff_A_mLacGsv77_1;
	wire w_dff_A_JNRB8m2A6_1;
	wire w_dff_A_yvJ5Qhd01_2;
	wire w_dff_A_eHn2MEGk4_2;
	wire w_dff_A_EYMn6Bug8_2;
	wire w_dff_A_MyUmvZKc4_2;
	wire w_dff_A_wsQ58IRP9_2;
	wire w_dff_A_LMtJko6c3_2;
	wire w_dff_A_FCIy9CXr2_2;
	wire w_dff_A_CyvMBjUf4_2;
	wire w_dff_A_sSQQ3S9O4_2;
	wire w_dff_A_kXLpwcdx6_2;
	wire w_dff_A_vjqMPCmp1_2;
	wire w_dff_A_Kziu9Gxh6_2;
	wire w_dff_A_u9j690ft2_2;
	wire w_dff_A_dXO5iyXF3_2;
	wire w_dff_A_eK5Mpd8I8_2;
	wire w_dff_A_2rQ3bUW76_2;
	wire w_dff_A_ccXMLJM11_0;
	wire w_dff_B_RGswLtgJ5_1;
	wire w_dff_A_TGkm35os1_0;
	wire w_dff_A_Z5GVPtXq1_2;
	wire w_dff_A_aeOguVQ19_1;
	wire w_dff_A_bc0Bi0ZA8_1;
	wire w_dff_B_X3IijG2u6_2;
	wire w_dff_B_SfXOQchI0_1;
	wire w_dff_B_NL5dvISo6_1;
	wire w_dff_A_pQUuYADs3_1;
	wire w_dff_A_sTeDeewm0_1;
	wire w_dff_A_vPBdSlVK8_1;
	wire w_dff_A_93WQQBLH2_1;
	wire w_dff_A_abu25aDs1_1;
	wire w_dff_A_RstvUsjn8_1;
	wire w_dff_A_OUBqBLoT3_2;
	wire w_dff_A_ZIQFC32R1_1;
	wire w_dff_B_63h7EG696_1;
	wire w_dff_B_StYp0G5t7_1;
	wire w_dff_B_Z9Mxv1hA2_1;
	wire w_dff_B_HvNdSAf63_1;
	wire w_dff_B_oNpQ3xAu0_0;
	wire w_dff_B_3kuTcEeI7_0;
	wire w_dff_A_Fwg64vac3_1;
	wire w_dff_A_aNrypkVs1_1;
	wire w_dff_A_EUoXFZbj8_1;
	wire w_dff_A_isgYk3tV9_2;
	wire w_dff_A_OFAGcWOO5_2;
	wire w_dff_B_2tWgEd0F4_0;
	wire w_dff_A_cPFeS07j5_0;
	wire w_dff_A_xeprSQiT4_0;
	wire w_dff_A_vW5kdLoO4_1;
	wire w_dff_A_fGpFw67W2_1;
	wire w_dff_A_3WNCWLUH0_0;
	wire w_dff_A_8kvExLf64_1;
	wire w_dff_A_QTvtvopw5_0;
	wire w_dff_A_SxZL3EJ99_2;
	wire w_dff_A_KxezhIql8_2;
	wire w_dff_A_V113hr1Z0_2;
	wire w_dff_A_dVMNW22K3_2;
	wire w_dff_A_QXcKkVHt5_1;
	wire w_dff_A_1P7dtv694_2;
	wire w_dff_A_U8GyUu3t4_2;
	wire w_dff_A_XwAUHr957_2;
	wire w_dff_A_lo75t7xT1_1;
	wire w_dff_A_Z8t0bqlT9_2;
	wire w_dff_A_cuKsTYLP9_2;
	wire w_dff_B_lpv1eGNU2_2;
	wire w_dff_B_q5J8ugWw8_2;
	wire w_dff_A_8Yt8kIRK5_0;
	wire w_dff_A_fyUY5LK18_0;
	wire w_dff_A_VwQATvQA5_0;
	wire w_dff_A_USAElrpB3_0;
	wire w_dff_A_KdVX5pSY1_1;
	wire w_dff_A_KXXiqvSB0_1;
	wire w_dff_A_bGh2cSlv5_1;
	wire w_dff_A_wKnIhUQ70_1;
	wire w_dff_A_6TU1WaPJ5_1;
	wire w_dff_A_s0awC98P6_1;
	wire w_dff_B_PTmXAk1V4_1;
	wire w_dff_A_mI2UI2xn8_0;
	wire w_dff_A_dzTU3Vk73_0;
	wire w_dff_A_2feKBVo45_1;
	wire w_dff_A_ZD5WqsF17_1;
	wire w_dff_A_4h9kr1yV2_1;
	wire w_dff_A_rwkKLZMV3_1;
	wire w_dff_A_3ESCjbCr0_1;
	wire w_dff_A_8P9ooGNz3_2;
	wire w_dff_A_TFUnVYZP2_2;
	wire w_dff_B_Se6rDN258_0;
	wire w_dff_A_QuFQc92y8_1;
	wire w_dff_B_MbbpWLVQ2_1;
	wire w_dff_A_5FWxVWEW6_1;
	wire w_dff_A_hGqcwpXw6_0;
	wire w_dff_A_j22ZuSF67_2;
	wire w_dff_A_jNGD2hGt5_2;
	wire w_dff_B_Rk1Okfz02_0;
	wire w_dff_B_rmTxIiOP8_1;
	wire w_dff_B_lWHQMiHx3_1;
	wire w_dff_A_tcJ3l1fM8_1;
	wire w_dff_A_XfCasgZQ5_2;
	wire w_dff_A_URbIeJxJ0_2;
	wire w_dff_A_D5qewFWh0_2;
	wire w_dff_A_NC2qA0Je7_2;
	wire w_dff_A_EgEJlBtd7_2;
	wire w_dff_A_v7eCRbFV2_0;
	wire w_dff_A_oFnLsIPX9_0;
	wire w_dff_A_wpfbVsDK0_0;
	wire w_dff_A_flNQp3ij0_1;
	wire w_dff_A_vR3aIkMQ4_1;
	wire w_dff_B_OjW9Vqor4_3;
	wire w_dff_B_3sFmpLJj0_3;
	wire w_dff_A_QCZ4uVcY2_0;
	wire w_dff_A_pu7qAetM1_0;
	wire w_dff_A_zBRlUt1m9_0;
	wire w_dff_A_yHfWBgP21_0;
	wire w_dff_A_vMdL48KJ7_0;
	wire w_dff_A_WitXuKAx9_0;
	wire w_dff_A_LnxMytRQ4_0;
	wire w_dff_A_AsFGWGqn1_0;
	wire w_dff_A_w7hLjyjp5_0;
	wire w_dff_A_AuvwHplx0_0;
	wire w_dff_A_Hp6CzNv34_0;
	wire w_dff_A_Yw1MRRPk8_0;
	wire w_dff_A_ivacLBdj2_0;
	wire w_dff_A_ONiH80fW8_0;
	wire w_dff_A_Qga8kDwT0_0;
	wire w_dff_A_hIiMCyqd5_0;
	wire w_dff_A_9LQ1UWGS1_0;
	wire w_dff_A_wGWEvXks2_0;
	wire w_dff_A_PPgkTpKD3_0;
	wire w_dff_A_TIhhQQDF5_0;
	wire w_dff_A_pbBn6JLd6_0;
	wire w_dff_A_LuFLmaxL6_0;
	wire w_dff_A_c6Fd7P0W7_1;
	wire w_dff_A_IsVMXQcS6_1;
	wire w_dff_A_6naygO3F7_1;
	wire w_dff_A_DKq2xQ6u8_1;
	wire w_dff_A_NKo3CyIm1_1;
	wire w_dff_A_yR7tohNl7_0;
	wire w_dff_A_tCDrSdfO1_0;
	wire w_dff_A_wfnlm8TV8_0;
	wire w_dff_A_9d4p2KhZ4_0;
	wire w_dff_A_sLxuViSS4_2;
	wire w_dff_A_TSxV9rCA7_2;
	wire w_dff_A_qzHAvkSR4_2;
	wire w_dff_A_2ev2g0lR9_2;
	wire w_dff_A_9qtZupMq0_2;
	wire w_dff_A_hDnjk1EL9_2;
	wire w_dff_A_NnQ7vhNI6_1;
	wire w_dff_A_F8I1H2sb2_1;
	wire w_dff_A_UV4VtZOZ0_1;
	wire w_dff_A_yNMjwTIC6_1;
	wire w_dff_A_TMobsgdo7_1;
	wire w_dff_A_y4GBWH5w5_1;
	wire w_dff_A_DLDWHXGW0_1;
	wire w_dff_A_gmu7h94X8_2;
	wire w_dff_A_xh99m26B7_2;
	wire w_dff_A_EEcE2K3w7_2;
	wire w_dff_A_7J9ktyR82_2;
	wire w_dff_A_pY5Wevk57_2;
	wire w_dff_A_XitxJwXg7_2;
	wire w_dff_A_bbdjmFzC1_2;
	wire w_dff_A_i7KpoBFg0_0;
	wire w_dff_A_OZZpiNyz2_2;
	wire w_dff_A_xOFY8sRx8_0;
	wire w_dff_A_31dEtmIx9_0;
	wire w_dff_A_uTS2VDkH1_1;
	wire w_dff_A_xhApSxfL6_1;
	wire w_dff_A_QSjvWHOz2_1;
	wire w_dff_A_L8MHFwn28_1;
	wire w_dff_A_HDnpnNPw1_1;
	wire w_dff_A_eA1RIcGE2_1;
	wire w_dff_A_475euyrk0_1;
	wire w_dff_A_Ak4a31pQ8_1;
	wire w_dff_A_zbv5gQFc3_1;
	wire w_dff_A_APQK90eA1_1;
	wire w_dff_A_sSlKkMgd4_1;
	wire w_dff_A_d5cGi8cl6_1;
	wire w_dff_A_97odbeVd7_1;
	wire w_dff_A_JjQpRUKt4_1;
	wire w_dff_A_oaT70Ert9_1;
	wire w_dff_A_KMEJokLl8_1;
	wire w_dff_A_yxanHp4w4_1;
	wire w_dff_A_hdHP6RrK9_1;
	wire w_dff_A_uYaC6xKx9_1;
	wire w_dff_B_qaOjpxk54_0;
	wire w_dff_B_lBI3HOGf2_1;
	wire w_dff_B_Ob1JtJHk1_1;
	wire w_dff_A_8MqtPDd34_0;
	wire w_dff_A_scipC3JV3_0;
	wire w_dff_A_hlJK438k8_0;
	wire w_dff_A_lBD9smrQ6_0;
	wire w_dff_A_xMGadafd5_0;
	wire w_dff_A_Z0FLKKmW4_0;
	wire w_dff_A_fMy63A7W0_0;
	wire w_dff_A_FzlvnR3r4_0;
	wire w_dff_A_UoXAoSkh7_0;
	wire w_dff_A_OtJncsHi2_1;
	wire w_dff_A_HwBBcvxQ0_1;
	wire w_dff_A_zA8cSDbK4_1;
	wire w_dff_A_ofqVPrrA0_0;
	wire w_dff_A_5oFpw9a35_1;
	wire w_dff_B_0ZqnHgth1_0;
	wire w_dff_A_5dVkZH5j0_0;
	wire w_dff_A_UaLXOGn53_0;
	wire w_dff_B_rBOlzuRi6_0;
	wire w_dff_A_HgI6wU3w3_0;
	wire w_dff_A_vTk5FaV18_1;
	wire w_dff_B_CckvPW0B8_0;
	wire w_dff_B_FItYXkBg8_1;
	wire w_dff_A_LnP6kG3p1_1;
	wire w_dff_A_vWUGqqlo7_1;
	wire w_dff_A_I3zk9c6d7_1;
	wire w_dff_A_YVQlmWJZ8_1;
	wire w_dff_A_qwKoobid7_1;
	wire w_dff_A_d09YCIYx6_1;
	wire w_dff_A_8Y5cjDrJ2_1;
	wire w_dff_A_nQrwdI367_2;
	wire w_dff_A_NMLBWp9v4_2;
	wire w_dff_A_lZhEDrAO9_2;
	wire w_dff_A_AVRwB63d9_2;
	wire w_dff_A_2EK5RY1d5_2;
	wire w_dff_A_CAEEaN0d5_2;
	wire w_dff_A_pX9m3u7g3_2;
	wire w_dff_B_YUhf0cSD3_0;
	wire w_dff_B_2Ups4ZUZ1_1;
	wire w_dff_A_r9xSnZwN3_1;
	wire w_dff_B_ESiqQjT38_1;
	wire w_dff_A_Z1wBMHEA7_0;
	wire w_dff_A_IQoxZCL04_0;
	wire w_dff_A_k0B8T4cV2_0;
	wire w_dff_A_X3OGsQtv9_1;
	wire w_dff_A_kryDyheK3_1;
	wire w_dff_A_JLnUbvKH6_1;
	wire w_dff_A_8vJy3UYI7_2;
	wire w_dff_A_HO9wEOsL3_1;
	wire w_dff_A_y18LBZqP9_2;
	wire w_dff_A_JyxRLC5D6_1;
	wire w_dff_A_4V7aPM779_1;
	wire w_dff_A_FPAyaDou3_0;
	wire w_dff_A_BjWdFFvn0_0;
	wire w_dff_A_IkzaHFq56_1;
	wire w_dff_A_ExKRS7R52_1;
	wire w_dff_A_DgwHk2E26_0;
	wire w_dff_A_yvlK8xgo9_2;
	wire w_dff_A_2nabn6W25_0;
	wire w_dff_A_KluREwqb8_0;
	wire w_dff_A_bOauCHnq3_0;
	wire w_dff_A_XGRbaAcM7_2;
	wire w_dff_A_qMub9GaM3_2;
	wire w_dff_A_olsPP0wh9_2;
	wire w_dff_A_w57tCPB92_0;
	wire w_dff_A_Doideh6u1_1;
	wire w_dff_A_UDaGBK512_1;
	wire w_dff_A_dCzj3Zxc8_1;
	wire w_dff_A_iypLFhgt0_1;
	wire w_dff_A_3U20ts2s3_1;
	wire w_dff_A_voGAwgge3_0;
	wire w_dff_A_2m34iBkZ9_0;
	wire w_dff_A_Gn9pDYYA7_0;
	wire w_dff_A_z5vr8YyK9_1;
	wire w_dff_A_mdV8smXh6_1;
	wire w_dff_A_rSAM8eBC8_1;
	wire w_dff_A_DYzNfhCS8_0;
	wire w_dff_A_87s3fh111_0;
	wire w_dff_A_HKylwl923_0;
	wire w_dff_A_cQ54mkdH5_0;
	wire w_dff_B_KP5W2ISa8_1;
	wire w_dff_A_82NHEE7b0_1;
	wire w_dff_A_aWCZ3PV36_1;
	wire w_dff_A_6i5ky61a5_0;
	wire w_dff_A_kIdF8Lbd6_0;
	wire w_dff_A_dRIFEpXE2_0;
	wire w_dff_A_hRLX5UKi5_1;
	wire w_dff_A_e2w0AW7a7_1;
	wire w_dff_A_ntHYKpwE3_1;
	wire w_dff_A_zHbiGjTa4_1;
	wire w_dff_A_2rZxIfci9_0;
	wire w_dff_A_wySlA28l1_0;
	wire w_dff_A_rs9LaVd82_0;
	wire w_dff_A_NgDrAnaq0_2;
	wire w_dff_A_3JGXcpoo3_2;
	wire w_dff_A_oCBzW6XC8_2;
	wire w_dff_A_r4fvZwfG5_2;
	wire w_dff_A_xM3lupbG2_1;
	wire w_dff_A_UCe6xSXk1_1;
	wire w_dff_A_FVoRFnKk5_1;
	wire w_dff_A_JKOTdtIu3_1;
	wire w_dff_A_sz6Xv0Vz2_2;
	wire w_dff_A_DpVal63g7_2;
	wire w_dff_B_g8zLtGBf1_1;
	wire w_dff_A_CvAUyHMO4_1;
	wire w_dff_A_SAu8rnnx7_0;
	wire w_dff_B_JTvsNzW86_2;
	wire w_dff_A_2QHmvWhb3_0;
	wire w_dff_A_5e450z2C9_0;
	wire w_dff_A_kV7y1LTJ4_0;
	wire w_dff_A_Scn0bNSL3_0;
	wire w_dff_A_3MA49UyW2_1;
	wire w_dff_A_5Ud1X3uD6_0;
	wire w_dff_A_5ICkNZKZ6_0;
	wire w_dff_A_8JtEjNTX7_0;
	wire w_dff_A_6SIYP9g29_1;
	wire w_dff_B_eeystC7o7_0;
	wire w_dff_B_cumdVIoI3_1;
	wire w_dff_A_Zr3jYwrt4_0;
	wire w_dff_A_K44SgIkp8_0;
	wire w_dff_A_2284LzIR3_0;
	wire w_dff_A_JmzGA6ll1_0;
	wire w_dff_A_IQNMlTkt4_1;
	wire w_dff_A_3qbxSaiM9_0;
	wire w_dff_A_yO1GxoUW4_0;
	wire w_dff_A_S3RsoBOp6_2;
	wire w_dff_A_wpN8eSkS4_2;
	wire w_dff_A_qlA9x71M5_2;
	wire w_dff_A_tDndV5yl1_2;
	wire w_dff_B_jOlQVX3f4_2;
	wire w_dff_B_XWyL3vEe4_2;
	wire w_dff_A_D9ebEIyT2_0;
	wire w_dff_A_5wqENpGk3_0;
	wire w_dff_A_MGIj5Kmt6_0;
	wire w_dff_A_MLMpndjC3_0;
	wire w_dff_A_Ww2dKrqe4_0;
	wire w_dff_A_eoP6Xd8S5_0;
	wire w_dff_A_KXzl8J1t1_0;
	wire w_dff_B_AdmWGaOe4_1;
	wire w_dff_B_97RKkF8C6_1;
	wire w_dff_A_bf5y3ZLr2_0;
	wire w_dff_A_7m6aJFYP6_0;
	wire w_dff_A_iUfZNA4n8_0;
	wire w_dff_A_dRMR1wIA9_1;
	wire w_dff_A_LdnhFLWB7_1;
	wire w_dff_A_cpfsNo8c5_0;
	wire w_dff_A_S7CcMjSb9_0;
	wire w_dff_A_dnvwvo7A0_0;
	wire w_dff_A_vrlGWjLz1_1;
	wire w_dff_A_7ehDI4M01_0;
	wire w_dff_A_iW93BtpF8_0;
	wire w_dff_A_VQhbRkxc1_0;
	wire w_dff_A_PVlXVh3K7_0;
	wire w_dff_A_R8TMyVsb5_1;
	wire w_dff_A_vWbAlTR88_1;
	wire w_dff_A_ltqoHmBF3_1;
	wire w_dff_A_xWL67o6i4_2;
	wire w_dff_A_U2PfyQfO1_2;
	wire w_dff_A_amvJWUy39_1;
	wire w_dff_A_LSUBSLPz7_0;
	wire w_dff_A_wRipiJfK3_0;
	wire w_dff_A_IDwFqbWc2_1;
	wire w_dff_A_wmPnpOg62_1;
	wire w_dff_A_70MqtVLv0_0;
	wire w_dff_A_CMYqqWq50_0;
	wire w_dff_A_qJosGXVx0_0;
	wire w_dff_A_yggG9FsL8_1;
	wire w_dff_A_nbD8OjSx0_1;
	wire w_dff_A_sfpgrEtx3_1;
	wire w_dff_A_qEGcM8sZ4_1;
	wire w_dff_A_xWkutRy76_0;
	wire w_dff_A_o2zAMAZe0_0;
	wire w_dff_A_HFEcO3OZ4_0;
	wire w_dff_A_ZXAphjHl9_1;
	wire w_dff_A_kQ9ZolWv4_1;
	wire w_dff_A_FRy2ruUc6_1;
	wire w_dff_A_Lrq5l9tN6_2;
	wire w_dff_B_WGGkR6IG8_1;
	wire w_dff_A_TFuT86eL8_0;
	wire w_dff_A_D1ne4K4h6_0;
	wire w_dff_A_sOPCTEl24_0;
	wire w_dff_A_mXjksGXB1_0;
	wire w_dff_A_DQBLRFxv6_0;
	wire w_dff_A_NMUsM9wm2_0;
	wire w_dff_A_YqcSp3Kl9_0;
	wire w_dff_A_nM2frNaL4_1;
	wire w_dff_A_DmpEb5RY1_2;
	wire w_dff_A_CCTZdFk07_2;
	wire w_dff_A_PC7hCPp52_2;
	wire w_dff_A_lrrUXja13_2;
	wire w_dff_A_KadsinUX2_2;
	wire w_dff_A_TkAhIzsv6_2;
	wire w_dff_A_qRkE6gDE0_2;
	wire w_dff_A_6bRW6Qnl2_0;
	wire w_dff_A_TcCrMEl05_0;
	wire w_dff_A_2ypiILTb6_0;
	wire w_dff_A_6NH8agMt2_0;
	wire w_dff_A_nw8f0R964_0;
	wire w_dff_A_hrPLdJey5_0;
	wire w_dff_A_e5MdD5iH7_0;
	wire w_dff_A_iEO4TAKl5_1;
	wire w_dff_A_od4RnqI36_1;
	wire w_dff_A_J7ajIevY0_1;
	wire w_dff_A_Qdhww1xq6_1;
	wire w_dff_A_n7LAqGNU5_1;
	wire w_dff_A_nBJU71419_0;
	wire w_dff_A_xlZw4z332_0;
	wire w_dff_B_VCunKxQB3_2;
	wire w_dff_A_yBIm5AGK6_0;
	wire w_dff_A_RJ3ehxuJ6_2;
	wire w_dff_A_dXo3rnxy2_1;
	wire w_dff_A_Yu58xckM0_0;
	wire w_dff_A_5DkLtjcb4_1;
	wire w_dff_A_jXJ1oX4K0_0;
	wire w_dff_A_vV1USWCc7_2;
	wire w_dff_B_8fRgtUxn3_3;
	wire w_dff_B_t0pyKXGU0_3;
	wire w_dff_B_aViKNqFt3_3;
	wire w_dff_B_jUizMbAi8_3;
	wire w_dff_B_gHcHtbaM1_3;
	wire w_dff_A_KMlib6jm0_0;
	wire w_dff_A_B2p8k5Fz8_0;
	wire w_dff_A_sCVs6zPD6_0;
	wire w_dff_A_brn168q66_0;
	wire w_dff_A_3JfNc2cQ6_0;
	wire w_dff_A_b5dhTsKc6_0;
	wire w_dff_A_J9O08y4f3_0;
	wire w_dff_A_Ogmw8Xod0_1;
	wire w_dff_A_S8rupHTl9_1;
	wire w_dff_A_Wd21yO0Q4_1;
	wire w_dff_A_OlEhyq3b3_1;
	wire w_dff_A_oLA0qMKS8_1;
	wire w_dff_A_EmEmE86E6_1;
	wire w_dff_A_Xfg6H6d67_1;
	wire w_dff_A_YJh1HPjB0_0;
	wire w_dff_A_tU4FM3tT9_0;
	wire w_dff_A_ccDNE53y1_0;
	wire w_dff_A_lpebNB3R4_0;
	wire w_dff_A_WHln3AV55_0;
	wire w_dff_A_XOhSyQFY7_0;
	wire w_dff_A_g2I0R6IE3_0;
	wire w_dff_B_wLkV8Msg4_0;
	wire w_dff_A_oUx6ewKo9_1;
	wire w_dff_A_nNOwGfR79_0;
	wire w_dff_A_0ImIa9oz1_0;
	wire w_dff_A_es4OKvcI0_2;
	wire w_dff_A_4rBuxrm07_0;
	wire w_dff_A_o5EKPjlR2_0;
	wire w_dff_A_9VJYIO237_2;
	wire w_dff_A_S0f0OtKf4_2;
	wire w_dff_A_5kn7p0kp0_2;
	wire w_dff_A_6naw0bNr9_2;
	wire w_dff_A_ln2asg344_0;
	wire w_dff_A_FGDdilbX4_1;
	wire w_dff_A_JWPKIpRZ9_1;
	wire w_dff_A_vnfRPm0D1_1;
	wire w_dff_A_6XzsJmGb0_1;
	wire w_dff_A_IVFQEA879_2;
	wire w_dff_A_f9Vx7bTT7_2;
	wire w_dff_A_C8ItDbhr4_2;
	wire w_dff_A_JzOAiOhW1_2;
	wire w_dff_A_j1CPUTnK0_2;
	wire w_dff_A_QN1UTpGE1_2;
	wire w_dff_A_IWIbbCRv4_2;
	wire w_dff_A_KLhsMzL80_2;
	wire w_dff_A_o2dkQw2X6_1;
	wire w_dff_A_Q72I1szT1_1;
	wire w_dff_A_t00ToI546_1;
	wire w_dff_A_hzSNvali3_2;
	wire w_dff_A_UQjn3JcF8_2;
	wire w_dff_A_5RDm4RVr9_2;
	wire w_dff_A_S8uciYKb7_0;
	wire w_dff_A_BmhYXBOh6_0;
	wire w_dff_A_fbC376HG6_0;
	wire w_dff_A_602sP49u2_1;
	wire w_dff_A_NBWhMjeI7_0;
	wire w_dff_A_aExwiZ3Z6_0;
	wire w_dff_A_LbDMwrdX5_2;
	wire w_dff_A_JtiMkx3W9_2;
	wire w_dff_A_s2DAGwOv7_2;
	wire w_dff_A_GWoSYVQn1_0;
	wire w_dff_A_W6NPhmPO4_0;
	wire w_dff_A_Ngq5RurS5_0;
	wire w_dff_A_v1DIj67w8_1;
	wire w_dff_A_aLKewj3f7_1;
	wire w_dff_A_81DlHO2N5_2;
	wire w_dff_A_ldhGD3Gr7_2;
	wire w_dff_A_oio6ptqe1_2;
	wire w_dff_A_Xs3u2aA27_1;
	wire w_dff_A_sVih4rfd4_0;
	wire w_dff_A_BiYpS19j7_1;
	wire w_dff_A_EXr1nqMF9_0;
	wire w_dff_A_ybmlZtvC9_2;
	wire w_dff_A_VQfRxLjO4_2;
	wire w_dff_A_wdiVNzGw5_2;
	wire w_dff_A_O2WVEmuP0_2;
	wire w_dff_A_nJpYmbT09_2;
	wire w_dff_A_7iLGToeL6_1;
	wire w_dff_A_N9Azsqpu1_0;
	wire w_dff_A_gKX85fBz5_2;
	wire w_dff_A_U7WxENXP3_0;
	wire w_dff_B_hMBDDOzB3_2;
	wire w_dff_B_Mf2fnBMK2_2;
	wire w_dff_A_Q9teBhin7_0;
	wire w_dff_A_Rwdh5tfI4_0;
	wire w_dff_A_mP813Pcd7_0;
	wire w_dff_A_cCjyevy15_2;
	wire w_dff_A_NGRSvjyA2_2;
	wire w_dff_A_hupm6H9s3_2;
	wire w_dff_A_qFESAoza9_2;
	wire w_dff_A_bh8X36zm6_1;
	wire w_dff_A_rAs9fs752_1;
	wire w_dff_A_zFlKy9Tf6_1;
	wire w_dff_A_37h6aHQw9_2;
	wire w_dff_A_RIYLDndJ8_0;
	wire w_dff_A_Hdd3lQoJ9_1;
	wire w_dff_A_OEIpwxEF5_0;
	wire w_dff_B_c3EoQMcj3_0;
	wire w_dff_A_F9yCgSqd8_0;
	wire w_dff_A_vFfXoTgA4_0;
	wire w_dff_A_LfpceVR85_0;
	wire w_dff_A_Z8i083sN4_2;
	wire w_dff_A_wNbrbeh79_2;
	wire w_dff_A_JZDmjjWv3_0;
	wire w_dff_B_sfNk1m3n4_0;
	wire w_dff_A_sflOr6SE6_2;
	wire w_dff_A_FHTOnRU44_0;
	wire w_dff_A_ruaDa1ua8_1;
	wire w_dff_A_plqwpa2X5_0;
	wire w_dff_A_MIU4X5zD8_2;
	wire w_dff_A_O4SyOYIf4_2;
	wire w_dff_A_AkNA0WSt5_2;
	wire w_dff_A_GjEuVDQb9_0;
	wire w_dff_A_Gg30chY37_0;
	wire w_dff_A_zAnPpuHg8_1;
	wire w_dff_A_YAkzqEdY8_1;
	wire w_dff_A_hz0rqOpc4_1;
	wire w_dff_A_O7RBQmC53_1;
	wire w_dff_A_ZqoXkDEg9_2;
	wire w_dff_A_MWBJbelM4_2;
	wire w_dff_A_mlsnI8yO0_2;
	wire w_dff_A_wnamHytM4_0;
	wire w_dff_A_Nhy7Pxuv0_1;
	wire w_dff_A_y1kiTWae9_0;
	wire w_dff_A_WgYvqrS63_0;
	wire w_dff_A_vVsBMaPY2_1;
	wire w_dff_A_72UFADII8_1;
	wire w_dff_B_CvdKY4r86_1;
	wire w_dff_A_Lqeye15K4_0;
	wire w_dff_A_IC5fUeBa9_0;
	wire w_dff_A_Jqq4jghV2_2;
	wire w_dff_A_mjO8ion64_2;
	wire w_dff_A_N71CIgGb6_1;
	wire w_dff_A_x1gD1Ai78_1;
	wire w_dff_A_wubsV4sU3_1;
	wire w_dff_A_bxeGtGKh1_2;
	wire w_dff_A_kCRtpCFN6_2;
	wire w_dff_A_0FigtYqf8_2;
	wire w_dff_A_7N9VqluI2_1;
	wire w_dff_A_lPXlGRsb0_1;
	wire w_dff_A_QBQC4kG27_1;
	wire w_dff_A_8pOBQB5E3_2;
	wire w_dff_A_Uj6RaHaN7_0;
	wire w_dff_A_SKieoeJM9_0;
	wire w_dff_A_jcx56kjk5_1;
	wire w_dff_A_Rb6IF7670_1;
	wire w_dff_A_tI7E6PyX4_1;
	wire w_dff_A_M9xudvUV9_1;
	wire w_dff_A_2x8NneIi5_2;
	wire w_dff_A_zG3jJkC47_2;
	wire w_dff_A_eZH5iZ0n7_2;
	wire w_dff_A_eXpKzxeD8_0;
	wire w_dff_A_XaWl6EhB4_0;
	wire w_dff_A_X4sKCKie2_1;
	wire w_dff_A_Bbp2fDwr8_1;
	wire w_dff_A_pBzLVghr5_1;
	wire w_dff_A_FjTqQqIS7_1;
	wire w_dff_A_NQqXkoGO5_2;
	wire w_dff_A_RKxoHzft5_2;
	wire w_dff_A_Zu2QdsRX7_2;
	wire w_dff_A_MvEArPr95_2;
	wire w_dff_A_lhwi2Cs43_1;
	wire w_dff_A_qojIAw5P2_1;
	wire w_dff_A_lMIT5JCa7_2;
	wire w_dff_A_LQBuzSCm1_2;
	wire w_dff_A_guEi5ejR3_1;
	wire w_dff_A_TQ9Ulg3a7_1;
	wire w_dff_A_SOrcP7xY6_0;
	wire w_dff_A_imXvUDCW9_1;
	wire w_dff_A_eAWEYyPb0_2;
	wire w_dff_A_bIepQwPZ9_2;
	wire w_dff_A_ztKs9EU99_2;
	wire w_dff_A_emGDu4J31_2;
	wire w_dff_A_HBy6B4246_2;
	wire w_dff_A_qDRWEKsA1_2;
	wire w_dff_A_YKI0fE2C8_2;
	wire w_dff_A_L884xvOs1_0;
	wire w_dff_A_Zcca7dj56_1;
	wire w_dff_A_gOULqPpa3_2;
	wire w_dff_A_ojIQhcSW4_1;
	wire w_dff_A_U5T40sHc3_2;
	wire w_dff_A_zTZXqXCx5_2;
	wire w_dff_A_IexZa1a62_0;
	wire w_dff_A_NB7BrxW80_2;
	wire w_dff_A_M6s2GyiG1_0;
	wire w_dff_A_cSmSc4Xu5_1;
	wire w_dff_A_KHhMTtkU8_1;
	wire w_dff_A_yrPrpbg44_1;
	wire w_dff_A_UuUqAC6S6_1;
	wire w_dff_A_GvZz6AZU1_1;
	wire w_dff_A_aWjUpErp0_1;
	wire w_dff_A_j9RaDmuA2_2;
	wire w_dff_A_w5GE8PKU8_2;
	wire w_dff_A_wKI40e3k2_2;
	wire w_dff_A_gkHTHtTR2_2;
	wire w_dff_A_HzDq4ZSw5_2;
	wire w_dff_A_EF4gWOik0_2;
	wire w_dff_A_Z9Ua2TPN8_0;
	wire w_dff_A_mwPkPso39_0;
	wire w_dff_A_yOV1ySzR8_0;
	wire w_dff_A_F4uQ5KSq5_0;
	wire w_dff_A_uAtBLhjT8_0;
	wire w_dff_A_Q10g6KuD1_0;
	wire w_dff_A_0eQoAOf32_0;
	wire w_dff_A_soBXMpL87_1;
	wire w_dff_A_0Itur3Zy0_1;
	wire w_dff_A_WTVt3mkB8_1;
	wire w_dff_A_raZPFetv9_1;
	wire w_dff_A_jSs7c7wO4_1;
	wire w_dff_A_JtQve0o20_1;
	wire w_dff_A_tbnSXAeN5_1;
	wire w_dff_A_cXLjNAtl1_2;
	wire w_dff_A_cjRJxW1x0_2;
	wire w_dff_A_tGIt2dJ92_2;
	wire w_dff_A_9yVzYEyV9_2;
	wire w_dff_A_pnsng7Im4_2;
	wire w_dff_A_2DD56qok2_2;
	wire w_dff_A_gYcfZmMb5_2;
	wire w_dff_A_9UgON85M6_2;
	wire w_dff_A_UX4Td7kW7_0;
	wire w_dff_A_BftYGRw05_0;
	wire w_dff_A_jnQOSjw22_0;
	wire w_dff_A_zq8GjPoa7_0;
	wire w_dff_A_UkQKU8MN8_0;
	wire w_dff_A_iZ0swn2t3_0;
	wire w_dff_A_YmiDJlxs6_0;
	wire w_dff_A_twUMrmTp5_0;
	wire w_dff_A_QGh853AF7_0;
	wire w_dff_A_4vmu8yGq9_0;
	wire w_dff_A_lLTWS1Wl1_0;
	wire w_dff_A_mwubIDYI7_0;
	wire w_dff_A_5aDZiB8w5_0;
	wire w_dff_A_j6Y7nI6U2_0;
	wire w_dff_A_pGiHP5Wr6_0;
	wire w_dff_A_68XgBR0N1_0;
	wire w_dff_A_KOoupgFN8_0;
	wire w_dff_A_bwYMGR4O4_0;
	wire w_dff_A_JPlebdm77_0;
	wire w_dff_A_qX5tQoTy3_0;
	wire w_dff_A_IQsoLb6z3_0;
	wire w_dff_A_i8MqfCfC3_0;
	wire w_dff_A_tugXxbQl4_0;
	wire w_dff_A_7LtWy9ON6_0;
	wire w_dff_A_VGKJsJxE9_1;
	wire w_dff_A_ig4PozfA5_0;
	wire w_dff_A_uzwQkORy9_0;
	wire w_dff_A_3ALl68WS6_0;
	wire w_dff_A_V35gbC4i6_0;
	wire w_dff_A_tCxKm7xA9_0;
	wire w_dff_A_t6XBcfqj6_0;
	wire w_dff_A_xL0zm0Fl5_0;
	wire w_dff_A_nJAOgdCd9_0;
	wire w_dff_A_FrnaEkXg9_0;
	wire w_dff_A_6fqnp5KR3_0;
	wire w_dff_A_ce7h9YRo9_0;
	wire w_dff_A_zNDDkFbe2_0;
	wire w_dff_A_fVPSZAq72_0;
	wire w_dff_A_I5PU5NZb9_0;
	wire w_dff_A_jUbTQsvT2_0;
	wire w_dff_A_N3xBY6Le3_0;
	wire w_dff_A_pNbxZHaQ8_0;
	wire w_dff_A_xwMGWpNP1_0;
	wire w_dff_A_414Rv4rQ6_0;
	wire w_dff_A_uY7Sf3477_0;
	wire w_dff_A_b3LfsZFr3_0;
	wire w_dff_A_iTN280Lp2_0;
	wire w_dff_A_f35KXooB9_0;
	wire w_dff_A_OClhKNEQ1_2;
	wire w_dff_A_FTUjRZ7L7_0;
	wire w_dff_A_2cCv4Uq26_0;
	wire w_dff_A_uZeBWyBl2_0;
	wire w_dff_A_q8aNVWan7_0;
	wire w_dff_A_U5jYb0Me2_0;
	wire w_dff_A_ACAoiT623_0;
	wire w_dff_A_1bHwmezi1_0;
	wire w_dff_A_D2Rjg7pc7_0;
	wire w_dff_A_L3LjZnyL1_0;
	wire w_dff_A_aFU4Geun3_0;
	wire w_dff_A_WziQ7ikS4_0;
	wire w_dff_A_GBsQMOTJ8_0;
	wire w_dff_A_lmkQI2SK4_0;
	wire w_dff_A_RJnLx0Ps7_0;
	wire w_dff_A_x1g1cW3Z6_0;
	wire w_dff_A_Hrh5qpCW6_0;
	wire w_dff_A_OQeLCToq2_0;
	wire w_dff_A_VuyDDf5T1_0;
	wire w_dff_A_9Mt7Ovpk7_0;
	wire w_dff_A_bk5lb8nL8_0;
	wire w_dff_A_CBmIP1Be0_2;
	wire w_dff_A_Gpm2Gb564_0;
	wire w_dff_A_W9RtSmlw4_0;
	wire w_dff_A_V1MY2djm8_0;
	wire w_dff_A_aIeawZzs5_0;
	wire w_dff_A_ZT55nFUa8_0;
	wire w_dff_A_4QVdc3U34_0;
	wire w_dff_A_lgQSOq4c1_0;
	wire w_dff_A_J4Br3uUv6_0;
	wire w_dff_A_yLPWMbr66_0;
	wire w_dff_A_SvvJkNuU9_0;
	wire w_dff_A_pSz1K8PI5_0;
	wire w_dff_A_VIAjZZZN7_0;
	wire w_dff_A_btfzpc5T9_0;
	wire w_dff_A_VQItuOtk3_0;
	wire w_dff_A_auBXnjy44_0;
	wire w_dff_A_9TKneLFD7_0;
	wire w_dff_A_wgvgXfY93_0;
	wire w_dff_A_4hQXFrDq2_0;
	wire w_dff_A_pnfM9AFv1_0;
	wire w_dff_A_Je0TwSxO1_0;
	wire w_dff_A_yl28ZcZy7_0;
	wire w_dff_A_kuuk5Rv47_0;
	wire w_dff_A_hUGUhDUA2_0;
	wire w_dff_A_xhxNDiQP5_2;
	wire w_dff_A_G8sReFIO7_0;
	wire w_dff_A_GOlZdwVX1_0;
	wire w_dff_A_g7Usebxg6_0;
	wire w_dff_A_OsqYQmCQ7_0;
	wire w_dff_A_hBCpgmvG9_0;
	wire w_dff_A_euATcaSn0_0;
	wire w_dff_A_JA7TipuW1_0;
	wire w_dff_A_krocCZFq9_0;
	wire w_dff_A_z0qIjVrv3_0;
	wire w_dff_A_qBxhkwf92_0;
	wire w_dff_A_JKZTHmqS5_0;
	wire w_dff_A_QOuv3Btq8_0;
	wire w_dff_A_gEiVgxUV9_0;
	wire w_dff_A_9Hv7a4ML5_0;
	wire w_dff_A_Qv4XXsdJ1_0;
	wire w_dff_A_3a5I1Iz07_0;
	wire w_dff_A_4OCRONKN0_0;
	wire w_dff_A_eqFUR6LR2_0;
	wire w_dff_A_bZDZd1ym5_0;
	wire w_dff_A_Zk1YGLwI3_0;
	wire w_dff_A_ieGty0Vc3_0;
	wire w_dff_A_ldNqHtrp9_0;
	wire w_dff_A_xa8ZCa0C5_0;
	wire w_dff_A_U1r5udv24_2;
	wire w_dff_A_ansNdKhk9_0;
	wire w_dff_A_6BMiPlfg1_0;
	wire w_dff_A_jXO6Q5Gk2_0;
	wire w_dff_A_1GjBFRWh5_0;
	wire w_dff_A_4IT75zj88_0;
	wire w_dff_A_576dMHkL5_0;
	wire w_dff_A_k1MVbUaM9_0;
	wire w_dff_A_jRHX9TTv0_0;
	wire w_dff_A_qZalfgYi8_0;
	wire w_dff_A_lDMgdEmu1_0;
	wire w_dff_A_CI0WGJSA8_0;
	wire w_dff_A_5UYdZsCK3_0;
	wire w_dff_A_U6EaKE1v6_0;
	wire w_dff_A_Rrj7Q0eY0_2;
	wire w_dff_A_sMvGYYQz5_0;
	wire w_dff_A_9zs5oxww3_0;
	wire w_dff_A_9s9YW4Cz7_0;
	wire w_dff_A_OELFuOV88_0;
	wire w_dff_A_F1weehSI0_0;
	wire w_dff_A_DE6tKUmO5_0;
	wire w_dff_A_zXoUCZGe1_0;
	wire w_dff_A_vufGJQ6A9_0;
	wire w_dff_A_rrHNbRHj1_0;
	wire w_dff_A_RAFXNA2R7_0;
	wire w_dff_A_Pv2N3cy47_0;
	wire w_dff_A_ePxRogil5_2;
	wire w_dff_A_896ZXHP37_0;
	wire w_dff_A_29WEVTCJ7_0;
	wire w_dff_A_XGLceOqF2_0;
	wire w_dff_A_lIJF73m14_0;
	wire w_dff_A_31zOZi8z4_0;
	wire w_dff_A_ASPMRDqh1_0;
	wire w_dff_A_4InhCdb05_0;
	wire w_dff_A_QBdaBEbx3_0;
	wire w_dff_A_6cz7jF5L6_0;
	wire w_dff_A_F6Fwcihu2_0;
	wire w_dff_A_FcBxUslg3_2;
	wire w_dff_A_YfmPqORr1_0;
	wire w_dff_A_zMLiY6PE5_0;
	wire w_dff_A_obHbBVlV0_0;
	wire w_dff_A_5oymxLVk5_0;
	wire w_dff_A_1wo000Vw3_0;
	wire w_dff_A_LCowYuNM1_0;
	wire w_dff_A_kRkRToyy2_0;
	wire w_dff_A_601qsepq9_0;
	wire w_dff_A_h8q06yD68_0;
	wire w_dff_A_plNEmITS6_0;
	wire w_dff_A_xU860ofM7_2;
	wire w_dff_A_2aK7iVgO7_0;
	wire w_dff_A_c6vS7XhE7_0;
	wire w_dff_A_nEIZ7oaJ9_0;
	wire w_dff_A_RsJWmTEr0_0;
	wire w_dff_A_nxGsCySq0_0;
	wire w_dff_A_L4ElTozG3_0;
	wire w_dff_A_tOCJwP9o9_0;
	wire w_dff_A_Nmw7ct6Y4_0;
	wire w_dff_A_RGK8DXxp7_0;
	wire w_dff_A_e0tgGeMz8_0;
	wire w_dff_A_du0s43qn6_1;
	wire w_dff_A_zNIYIL1a4_0;
	wire w_dff_A_mLjXaajH3_0;
	wire w_dff_A_8EMbMuO37_0;
	wire w_dff_A_nl32DYBz4_0;
	wire w_dff_A_yIiR2RH77_0;
	wire w_dff_A_FSORTYGC7_0;
	wire w_dff_A_CfeXRRy36_0;
	wire w_dff_A_WtxJkxnW0_2;
	wire w_dff_A_kvZW2pNS3_0;
	wire w_dff_A_q8kxXbp53_0;
	wire w_dff_A_dMo2TFOl9_0;
	wire w_dff_A_2PnyNn0i6_0;
	wire w_dff_A_FnlWl4Ri9_2;
	wire w_dff_A_lCWnU55g8_0;
	wire w_dff_A_3G595ny84_0;
	wire w_dff_A_1xfDIt8f7_0;
	wire w_dff_A_KJ62ScuT9_0;
	wire w_dff_A_HbcdcMhN5_1;
	wire w_dff_A_56KqB1r02_0;
	wire w_dff_A_7N4LheIH7_0;
	wire w_dff_A_qekMxyrJ1_0;
	wire w_dff_A_qsCD0GK29_0;
	wire w_dff_A_ndSfgAv18_0;
	wire w_dff_A_9u21ON9p7_0;
	wire w_dff_A_Xq1tvspa5_1;
	wire w_dff_A_nnOmNew95_0;
	wire w_dff_A_KuCBcFFz1_0;
	wire w_dff_A_HGJsfUsS7_0;
	wire w_dff_A_g3M5ctib2_0;
	wire w_dff_A_CXI4NZcl3_0;
	wire w_dff_A_XeMRgOBq9_1;
	wire w_dff_A_tRgQlSEG7_0;
	wire w_dff_A_TugvvbVr3_0;
	wire w_dff_A_e7jcRQLs2_0;
	wire w_dff_A_3x8hGX1b5_0;
	wire w_dff_A_suoffQtL3_1;
	wire w_dff_A_WkLmf1A43_0;
	wire w_dff_A_TBa6wdVG1_0;
	wire w_dff_A_BWmK6cNT5_1;
	wire w_dff_A_Svc0U3fn9_0;
	wire w_dff_A_Wir5E6q46_0;
	wire w_dff_A_QW8FzAo49_0;
	wire w_dff_A_Tn1IrHG90_0;
	wire w_dff_A_cajdjt8l9_1;
	wire w_dff_A_AmqgxAwU4_2;
	jnot g0000(.din(w_G77_5[1]),.dout(n72),.clk(gclk));
	jnot g0001(.din(w_G50_5[2]),.dout(n73),.clk(gclk));
	jnot g0002(.din(w_G58_5[1]),.dout(n74),.clk(gclk));
	jnot g0003(.din(w_G68_5[1]),.dout(n75),.clk(gclk));
	jand g0004(.dina(w_n75_1[1]),.dinb(w_n74_1[1]),.dout(n76),.clk(gclk));
	jand g0005(.dina(w_n76_0[1]),.dinb(w_n73_2[2]),.dout(n77),.clk(gclk));
	jand g0006(.dina(w_n77_0[1]),.dinb(w_n72_1[1]),.dout(w_dff_A_9UgON85M6_2),.clk(gclk));
	jnot g0007(.din(w_G97_5[1]),.dout(n79),.clk(gclk));
	jnot g0008(.din(w_G107_5[1]),.dout(n80),.clk(gclk));
	jand g0009(.dina(w_n80_1[1]),.dinb(w_n79_0[2]),.dout(n81),.clk(gclk));
	jnot g0010(.din(w_n81_0[2]),.dout(n82),.clk(gclk));
	jand g0011(.dina(n82),.dinb(w_G87_3[2]),.dout(n83),.clk(gclk));
	jnot g0012(.din(n83),.dout(G355_fa_),.clk(gclk));
	jand g0013(.dina(w_G20_7[1]),.dinb(w_G1_3[1]),.dout(n85),.clk(gclk));
	jnot g0014(.din(w_G226_1[1]),.dout(n86),.clk(gclk));
	jor g0015(.dina(w_n86_0[1]),.dinb(w_n73_2[1]),.dout(n87),.clk(gclk));
	jnot g0016(.din(w_G264_1[1]),.dout(n88),.clk(gclk));
	jor g0017(.dina(w_n88_1[1]),.dinb(w_n80_1[0]),.dout(n89),.clk(gclk));
	jand g0018(.dina(n89),.dinb(n87),.dout(n90),.clk(gclk));
	jnot g0019(.din(w_G257_1[2]),.dout(n91),.clk(gclk));
	jor g0020(.dina(w_n91_1[2]),.dinb(w_n79_0[1]),.dout(n92),.clk(gclk));
	jnot g0021(.din(w_G238_1[2]),.dout(n93),.clk(gclk));
	jor g0022(.dina(w_n93_0[1]),.dinb(w_n75_1[0]),.dout(n94),.clk(gclk));
	jand g0023(.dina(n94),.dinb(n92),.dout(n95),.clk(gclk));
	jand g0024(.dina(n95),.dinb(n90),.dout(n96),.clk(gclk));
	jnot g0025(.din(w_G87_3[1]),.dout(n97),.clk(gclk));
	jnot g0026(.din(w_G250_0[2]),.dout(n98),.clk(gclk));
	jor g0027(.dina(w_n98_2[1]),.dinb(w_n97_2[1]),.dout(n99),.clk(gclk));
	jnot g0028(.din(w_G232_1[2]),.dout(n100),.clk(gclk));
	jor g0029(.dina(n100),.dinb(w_n74_1[0]),.dout(n101),.clk(gclk));
	jand g0030(.dina(n101),.dinb(n99),.dout(n102),.clk(gclk));
	jnot g0031(.din(w_G244_1[2]),.dout(n103),.clk(gclk));
	jor g0032(.dina(w_n103_0[2]),.dinb(w_n72_1[0]),.dout(n104),.clk(gclk));
	jnot g0033(.din(w_G116_4[2]),.dout(n105),.clk(gclk));
	jnot g0034(.din(w_G270_0[2]),.dout(n106),.clk(gclk));
	jor g0035(.dina(w_n106_0[1]),.dinb(w_n105_2[1]),.dout(n107),.clk(gclk));
	jand g0036(.dina(n107),.dinb(n104),.dout(n108),.clk(gclk));
	jand g0037(.dina(n108),.dinb(n102),.dout(n109),.clk(gclk));
	jand g0038(.dina(n109),.dinb(n96),.dout(n110),.clk(gclk));
	jor g0039(.dina(n110),.dinb(w_n85_0[2]),.dout(n111),.clk(gclk));
	jnot g0040(.din(w_G20_7[0]),.dout(n112),.clk(gclk));
	jnot g0041(.din(w_G1_3[0]),.dout(n113),.clk(gclk));
	jnot g0042(.din(w_G13_1[1]),.dout(n114),.clk(gclk));
	jor g0043(.dina(w_n114_1[2]),.dinb(w_n113_3[1]),.dout(n115),.clk(gclk));
	jor g0044(.dina(w_n115_1[1]),.dinb(w_n112_5[2]),.dout(n116),.clk(gclk));
	jnot g0045(.din(w_n76_0[0]),.dout(n117),.clk(gclk));
	jand g0046(.dina(n117),.dinb(w_G50_5[1]),.dout(n118),.clk(gclk));
	jnot g0047(.din(w_n118_0[2]),.dout(n119),.clk(gclk));
	jor g0048(.dina(n119),.dinb(w_n116_0[1]),.dout(n120),.clk(gclk));
	jand g0049(.dina(w_n114_1[1]),.dinb(w_G1_2[2]),.dout(n121),.clk(gclk));
	jand g0050(.dina(w_n121_0[2]),.dinb(w_G20_6[2]),.dout(n122),.clk(gclk));
	jnot g0051(.din(w_n122_1[1]),.dout(n123),.clk(gclk));
	jand g0052(.dina(w_n88_1[0]),.dinb(w_n91_1[1]),.dout(n124),.clk(gclk));
	jor g0053(.dina(n124),.dinb(w_n98_2[0]),.dout(n125),.clk(gclk));
	jor g0054(.dina(w_dff_B_FHdOARZ04_0),.dinb(w_n123_1[2]),.dout(n126),.clk(gclk));
	jand g0055(.dina(w_dff_B_nTRQHFet8_0),.dinb(n120),.dout(n127),.clk(gclk));
	jand g0056(.dina(n127),.dinb(w_dff_B_8aZMsUSg1_1),.dout(w_dff_A_OClhKNEQ1_2),.clk(gclk));
	jxor g0057(.dina(w_G270_0[1]),.dinb(w_G264_1[0]),.dout(n129),.clk(gclk));
	jxor g0058(.dina(w_G257_1[1]),.dinb(w_n98_1[2]),.dout(n130),.clk(gclk));
	jxor g0059(.dina(n130),.dinb(w_dff_B_kUtKdGEd3_1),.dout(n131),.clk(gclk));
	jnot g0060(.din(w_n131_0[1]),.dout(n132),.clk(gclk));
	jxor g0061(.dina(w_G244_1[1]),.dinb(w_G238_1[1]),.dout(n133),.clk(gclk));
	jxor g0062(.dina(w_G232_1[1]),.dinb(w_n86_0[0]),.dout(n134),.clk(gclk));
	jxor g0063(.dina(n134),.dinb(w_dff_B_tZwGx5NQ2_1),.dout(n135),.clk(gclk));
	jxor g0064(.dina(w_n135_0[1]),.dinb(n132),.dout(w_dff_A_CBmIP1Be0_2),.clk(gclk));
	jxor g0065(.dina(w_G68_5[0]),.dinb(w_G58_5[0]),.dout(n137),.clk(gclk));
	jnot g0066(.din(w_n137_0[2]),.dout(n138),.clk(gclk));
	jxor g0067(.dina(w_G77_5[0]),.dinb(w_G50_5[0]),.dout(n139),.clk(gclk));
	jxor g0068(.dina(w_dff_B_0eotRJax5_0),.dinb(n138),.dout(n140),.clk(gclk));
	jnot g0069(.din(w_n140_0[1]),.dout(n141),.clk(gclk));
	jxor g0070(.dina(w_G116_4[1]),.dinb(w_G107_5[0]),.dout(n142),.clk(gclk));
	jxor g0071(.dina(w_G97_5[0]),.dinb(w_n97_2[0]),.dout(n143),.clk(gclk));
	jxor g0072(.dina(n143),.dinb(w_dff_B_R0hu89kZ0_1),.dout(n144),.clk(gclk));
	jxor g0073(.dina(w_n144_0[1]),.dinb(n141),.dout(w_dff_A_xhxNDiQP5_2),.clk(gclk));
	jnot g0074(.din(w_G169_1[1]),.dout(n146),.clk(gclk));
	jand g0075(.dina(w_G13_1[0]),.dinb(w_G1_2[1]),.dout(n147),.clk(gclk));
	jnot g0076(.din(w_G33_11[2]),.dout(n148),.clk(gclk));
	jnot g0077(.din(w_G41_1[1]),.dout(n149),.clk(gclk));
	jor g0078(.dina(w_n149_2[1]),.dinb(w_n148_9[2]),.dout(n150),.clk(gclk));
	jand g0079(.dina(n150),.dinb(w_n147_0[2]),.dout(n151),.clk(gclk));
	jand g0080(.dina(w_G1698_0[2]),.dinb(w_n148_9[1]),.dout(n152),.clk(gclk));
	jand g0081(.dina(w_n152_3[1]),.dinb(w_G244_1[0]),.dout(n153),.clk(gclk));
	jnot g0082(.din(w_G1698_0[1]),.dout(n154),.clk(gclk));
	jand g0083(.dina(w_n154_0[1]),.dinb(w_n148_9[0]),.dout(n155),.clk(gclk));
	jand g0084(.dina(w_n155_3[1]),.dinb(w_G238_1[0]),.dout(n156),.clk(gclk));
	jand g0085(.dina(w_G116_4[0]),.dinb(w_G33_11[1]),.dout(n157),.clk(gclk));
	jor g0086(.dina(w_n157_0[2]),.dinb(n156),.dout(n158),.clk(gclk));
	jor g0087(.dina(n158),.dinb(w_dff_B_CvdKY4r86_1),.dout(n159),.clk(gclk));
	jand g0088(.dina(n159),.dinb(w_n151_4[2]),.dout(n160),.clk(gclk));
	jnot g0089(.din(w_G45_1[2]),.dout(n161),.clk(gclk));
	jor g0090(.dina(w_n161_1[1]),.dinb(w_G1_2[0]),.dout(n162),.clk(gclk));
	jand g0091(.dina(w_n162_0[2]),.dinb(w_n98_1[1]),.dout(n163),.clk(gclk));
	jnot g0092(.din(w_n163_0[1]),.dout(n164),.clk(gclk));
	jand g0093(.dina(w_G41_1[0]),.dinb(w_G33_11[0]),.dout(n165),.clk(gclk));
	jor g0094(.dina(w_dff_B_sfNk1m3n4_0),.dinb(w_n115_1[0]),.dout(n166),.clk(gclk));
	jor g0095(.dina(w_n162_0[1]),.dinb(w_G274_0[2]),.dout(n167),.clk(gclk));
	jand g0096(.dina(n167),.dinb(w_n166_3[1]),.dout(n168),.clk(gclk));
	jand g0097(.dina(n168),.dinb(n164),.dout(n169),.clk(gclk));
	jor g0098(.dina(w_dff_B_c3EoQMcj3_0),.dinb(n160),.dout(n170),.clk(gclk));
	jand g0099(.dina(w_n170_0[2]),.dinb(w_n146_3[2]),.dout(n171),.clk(gclk));
	jand g0100(.dina(w_G97_4[2]),.dinb(w_G33_10[2]),.dout(n172),.clk(gclk));
	jand g0101(.dina(w_G68_4[2]),.dinb(w_n148_8[2]),.dout(n173),.clk(gclk));
	jor g0102(.dina(n173),.dinb(w_G20_6[1]),.dout(n174),.clk(gclk));
	jor g0103(.dina(n174),.dinb(w_n172_0[1]),.dout(n175),.clk(gclk));
	jnot g0104(.din(n175),.dout(n176),.clk(gclk));
	jor g0105(.dina(w_n112_5[1]),.dinb(w_n113_3[0]),.dout(n177),.clk(gclk));
	jor g0106(.dina(n177),.dinb(w_n148_8[1]),.dout(n178),.clk(gclk));
	jand g0107(.dina(n178),.dinb(w_n115_0[2]),.dout(n179),.clk(gclk));
	jand g0108(.dina(w_n81_0[1]),.dinb(w_n97_1[2]),.dout(n180),.clk(gclk));
	jand g0109(.dina(w_n180_0[1]),.dinb(w_G20_6[0]),.dout(n181),.clk(gclk));
	jor g0110(.dina(n181),.dinb(w_n179_1[2]),.dout(n182),.clk(gclk));
	jor g0111(.dina(n182),.dinb(n176),.dout(n183),.clk(gclk));
	jand g0112(.dina(w_G20_5[2]),.dinb(w_n113_2[2]),.dout(n184),.clk(gclk));
	jand g0113(.dina(n184),.dinb(w_G13_0[2]),.dout(n185),.clk(gclk));
	jand g0114(.dina(w_n185_3[2]),.dinb(w_n97_1[1]),.dout(n186),.clk(gclk));
	jnot g0115(.din(n186),.dout(n187),.clk(gclk));
	jand g0116(.dina(w_n85_0[1]),.dinb(w_G33_10[1]),.dout(n188),.clk(gclk));
	jor g0117(.dina(n188),.dinb(w_n147_0[1]),.dout(n189),.clk(gclk));
	jor g0118(.dina(w_n185_3[1]),.dinb(w_n189_2[1]),.dout(n190),.clk(gclk));
	jand g0119(.dina(w_G33_10[0]),.dinb(w_n113_2[1]),.dout(n191),.clk(gclk));
	jor g0120(.dina(w_n191_0[2]),.dinb(w_n97_1[0]),.dout(n192),.clk(gclk));
	jor g0121(.dina(w_dff_B_wLkV8Msg4_0),.dinb(w_n190_1[2]),.dout(n193),.clk(gclk));
	jand g0122(.dina(n193),.dinb(n187),.dout(n194),.clk(gclk));
	jand g0123(.dina(n194),.dinb(n183),.dout(n195),.clk(gclk));
	jnot g0124(.din(w_G179_2[2]),.dout(n196),.clk(gclk));
	jor g0125(.dina(w_n154_0[0]),.dinb(w_G33_9[2]),.dout(n197),.clk(gclk));
	jor g0126(.dina(w_n197_1[1]),.dinb(w_n103_0[1]),.dout(n198),.clk(gclk));
	jor g0127(.dina(w_G1698_0[0]),.dinb(w_G33_9[1]),.dout(n199),.clk(gclk));
	jor g0128(.dina(w_n199_1[1]),.dinb(w_n93_0[0]),.dout(n200),.clk(gclk));
	jnot g0129(.din(w_n157_0[1]),.dout(n201),.clk(gclk));
	jand g0130(.dina(w_n201_0[1]),.dinb(n200),.dout(n202),.clk(gclk));
	jand g0131(.dina(n202),.dinb(n198),.dout(n203),.clk(gclk));
	jor g0132(.dina(n203),.dinb(w_n166_3[0]),.dout(n204),.clk(gclk));
	jnot g0133(.din(w_G274_0[1]),.dout(n205),.clk(gclk));
	jand g0134(.dina(w_G45_1[1]),.dinb(w_n113_2[0]),.dout(n206),.clk(gclk));
	jand g0135(.dina(w_n206_0[1]),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jor g0136(.dina(n207),.dinb(w_n151_4[1]),.dout(n208),.clk(gclk));
	jor g0137(.dina(n208),.dinb(w_n163_0[0]),.dout(n209),.clk(gclk));
	jand g0138(.dina(n209),.dinb(n204),.dout(n210),.clk(gclk));
	jand g0139(.dina(w_n210_0[2]),.dinb(w_n196_2[2]),.dout(n211),.clk(gclk));
	jor g0140(.dina(n211),.dinb(w_n195_0[1]),.dout(n212),.clk(gclk));
	jor g0141(.dina(n212),.dinb(n171),.dout(n213),.clk(gclk));
	jnot g0142(.din(w_n195_0[0]),.dout(n214),.clk(gclk));
	jand g0143(.dina(w_n210_0[1]),.dinb(w_G190_4[1]),.dout(n215),.clk(gclk));
	jand g0144(.dina(w_n170_0[1]),.dinb(w_G200_4[2]),.dout(n216),.clk(gclk));
	jor g0145(.dina(n216),.dinb(w_dff_B_WGGkR6IG8_1),.dout(n217),.clk(gclk));
	jor g0146(.dina(n217),.dinb(w_n214_0[1]),.dout(n218),.clk(gclk));
	jand g0147(.dina(w_n218_0[1]),.dinb(w_n213_0[1]),.dout(n219),.clk(gclk));
	jor g0148(.dina(w_n197_1[0]),.dinb(w_n98_1[0]),.dout(n220),.clk(gclk));
	jand g0149(.dina(w_G283_3[2]),.dinb(w_G33_9[0]),.dout(n221),.clk(gclk));
	jnot g0150(.din(w_n221_0[2]),.dout(n222),.clk(gclk));
	jor g0151(.dina(w_n199_1[0]),.dinb(w_n103_0[0]),.dout(n223),.clk(gclk));
	jand g0152(.dina(n223),.dinb(n222),.dout(n224),.clk(gclk));
	jand g0153(.dina(n224),.dinb(n220),.dout(n225),.clk(gclk));
	jor g0154(.dina(n225),.dinb(w_n166_2[2]),.dout(n226),.clk(gclk));
	jor g0155(.dina(w_n151_4[0]),.dinb(w_n205_0[0]),.dout(n227),.clk(gclk));
	jor g0156(.dina(w_n162_0[0]),.dinb(w_G41_0[2]),.dout(n228),.clk(gclk));
	jor g0157(.dina(w_n228_0[1]),.dinb(n227),.dout(n229),.clk(gclk));
	jand g0158(.dina(w_n206_0[0]),.dinb(w_n149_2[0]),.dout(n230),.clk(gclk));
	jor g0159(.dina(w_n230_0[1]),.dinb(w_n151_3[2]),.dout(n231),.clk(gclk));
	jor g0160(.dina(w_n231_0[2]),.dinb(w_n91_1[0]),.dout(n232),.clk(gclk));
	jand g0161(.dina(n232),.dinb(w_n229_0[2]),.dout(n233),.clk(gclk));
	jand g0162(.dina(n233),.dinb(w_dff_B_97RKkF8C6_1),.dout(n234),.clk(gclk));
	jor g0163(.dina(w_n234_0[2]),.dinb(w_n146_3[1]),.dout(n235),.clk(gclk));
	jand g0164(.dina(w_n152_3[0]),.dinb(w_G250_0[1]),.dout(n236),.clk(gclk));
	jand g0165(.dina(w_n155_3[0]),.dinb(w_G244_0[2]),.dout(n237),.clk(gclk));
	jor g0166(.dina(n237),.dinb(w_n221_0[1]),.dout(n238),.clk(gclk));
	jor g0167(.dina(n238),.dinb(w_dff_B_AdmWGaOe4_1),.dout(n239),.clk(gclk));
	jand g0168(.dina(n239),.dinb(w_n151_3[1]),.dout(n240),.clk(gclk));
	jand g0169(.dina(w_n166_2[1]),.dinb(w_G274_0[0]),.dout(n241),.clk(gclk));
	jand g0170(.dina(w_n230_0[0]),.dinb(w_n241_0[1]),.dout(n242),.clk(gclk));
	jand g0171(.dina(w_n228_0[0]),.dinb(w_n166_2[0]),.dout(n243),.clk(gclk));
	jand g0172(.dina(w_n243_0[2]),.dinb(w_G257_1[0]),.dout(n244),.clk(gclk));
	jor g0173(.dina(n244),.dinb(w_n242_0[2]),.dout(n245),.clk(gclk));
	jor g0174(.dina(n245),.dinb(n240),.dout(n246),.clk(gclk));
	jor g0175(.dina(w_n246_1[1]),.dinb(w_n196_2[1]),.dout(n247),.clk(gclk));
	jand g0176(.dina(n247),.dinb(n235),.dout(n248),.clk(gclk));
	jand g0177(.dina(w_G107_4[2]),.dinb(w_G33_8[2]),.dout(n249),.clk(gclk));
	jand g0178(.dina(w_G77_4[2]),.dinb(w_n148_8[0]),.dout(n250),.clk(gclk));
	jor g0179(.dina(n250),.dinb(w_G20_5[1]),.dout(n251),.clk(gclk));
	jor g0180(.dina(n251),.dinb(w_n249_0[1]),.dout(n252),.clk(gclk));
	jand g0181(.dina(w_G107_4[1]),.dinb(w_G97_4[1]),.dout(n253),.clk(gclk));
	jor g0182(.dina(n253),.dinb(w_n112_5[0]),.dout(n254),.clk(gclk));
	jor g0183(.dina(n254),.dinb(w_n81_0[0]),.dout(n255),.clk(gclk));
	jand g0184(.dina(w_n255_0[1]),.dinb(n252),.dout(n256),.clk(gclk));
	jand g0185(.dina(n256),.dinb(w_n189_2[0]),.dout(n257),.clk(gclk));
	jnot g0186(.din(w_n257_0[1]),.dout(n258),.clk(gclk));
	jand g0187(.dina(w_n185_3[0]),.dinb(w_n79_0[0]),.dout(n259),.clk(gclk));
	jnot g0188(.din(w_n259_0[1]),.dout(n260),.clk(gclk));
	jnot g0189(.din(w_n191_0[1]),.dout(n261),.clk(gclk));
	jand g0190(.dina(w_n261_0[1]),.dinb(w_G97_4[0]),.dout(n262),.clk(gclk));
	jnot g0191(.din(w_n262_0[1]),.dout(n263),.clk(gclk));
	jor g0192(.dina(n263),.dinb(w_n190_1[1]),.dout(n264),.clk(gclk));
	jand g0193(.dina(n264),.dinb(w_dff_B_cumdVIoI3_1),.dout(n265),.clk(gclk));
	jand g0194(.dina(n265),.dinb(n258),.dout(n266),.clk(gclk));
	jor g0195(.dina(w_dff_B_eeystC7o7_0),.dinb(n248),.dout(n267),.clk(gclk));
	jand g0196(.dina(w_n246_1[0]),.dinb(w_G200_4[1]),.dout(n268),.clk(gclk));
	jor g0197(.dina(w_n112_4[2]),.dinb(w_G1_1[2]),.dout(n269),.clk(gclk));
	jor g0198(.dina(w_n269_1[2]),.dinb(w_n114_1[0]),.dout(n270),.clk(gclk));
	jand g0199(.dina(w_n270_0[1]),.dinb(w_n179_1[1]),.dout(n271),.clk(gclk));
	jand g0200(.dina(w_n262_0[0]),.dinb(w_n271_1[2]),.dout(n272),.clk(gclk));
	jor g0201(.dina(n272),.dinb(w_n259_0[0]),.dout(n273),.clk(gclk));
	jor g0202(.dina(n273),.dinb(w_n257_0[0]),.dout(n274),.clk(gclk));
	jand g0203(.dina(w_n234_0[1]),.dinb(w_G190_4[0]),.dout(n275),.clk(gclk));
	jor g0204(.dina(n275),.dinb(w_n274_0[2]),.dout(n276),.clk(gclk));
	jor g0205(.dina(n276),.dinb(w_dff_B_g8zLtGBf1_1),.dout(n277),.clk(gclk));
	jand g0206(.dina(n277),.dinb(n267),.dout(n278),.clk(gclk));
	jand g0207(.dina(w_n278_0[1]),.dinb(w_n219_0[1]),.dout(n279),.clk(gclk));
	jand g0208(.dina(w_n152_2[2]),.dinb(w_G264_0[2]),.dout(n280),.clk(gclk));
	jand g0209(.dina(w_G303_2[2]),.dinb(w_G33_8[1]),.dout(n281),.clk(gclk));
	jand g0210(.dina(w_n155_2[2]),.dinb(w_G257_0[2]),.dout(n282),.clk(gclk));
	jor g0211(.dina(n282),.dinb(w_n281_0[1]),.dout(n283),.clk(gclk));
	jor g0212(.dina(n283),.dinb(w_dff_B_KP5W2ISa8_1),.dout(n284),.clk(gclk));
	jand g0213(.dina(n284),.dinb(w_n151_3[0]),.dout(n285),.clk(gclk));
	jand g0214(.dina(w_n243_0[1]),.dinb(w_G270_0[0]),.dout(n286),.clk(gclk));
	jor g0215(.dina(n286),.dinb(w_n242_0[1]),.dout(n287),.clk(gclk));
	jor g0216(.dina(n287),.dinb(n285),.dout(n288),.clk(gclk));
	jand g0217(.dina(w_n288_1[1]),.dinb(w_n146_3[0]),.dout(n289),.clk(gclk));
	jand g0218(.dina(w_G97_3[2]),.dinb(w_n148_7[2]),.dout(n290),.clk(gclk));
	jor g0219(.dina(n290),.dinb(w_G20_5[0]),.dout(n291),.clk(gclk));
	jor g0220(.dina(n291),.dinb(w_n221_0[0]),.dout(n292),.clk(gclk));
	jand g0221(.dina(w_n105_2[0]),.dinb(w_G20_4[2]),.dout(n293),.clk(gclk));
	jnot g0222(.din(n293),.dout(n294),.clk(gclk));
	jand g0223(.dina(n294),.dinb(w_n189_1[2]),.dout(n295),.clk(gclk));
	jand g0224(.dina(n295),.dinb(n292),.dout(n296),.clk(gclk));
	jnot g0225(.din(w_n296_0[1]),.dout(n297),.clk(gclk));
	jand g0226(.dina(w_n185_2[2]),.dinb(w_n105_1[2]),.dout(n298),.clk(gclk));
	jnot g0227(.din(w_n298_0[1]),.dout(n299),.clk(gclk));
	jor g0228(.dina(w_n191_0[0]),.dinb(w_n105_1[1]),.dout(n300),.clk(gclk));
	jor g0229(.dina(w_n300_0[1]),.dinb(w_n190_1[0]),.dout(n301),.clk(gclk));
	jand g0230(.dina(n301),.dinb(n299),.dout(n302),.clk(gclk));
	jand g0231(.dina(n302),.dinb(n297),.dout(n303),.clk(gclk));
	jor g0232(.dina(w_n197_0[2]),.dinb(w_n88_0[2]),.dout(n304),.clk(gclk));
	jnot g0233(.din(w_n281_0[0]),.dout(n305),.clk(gclk));
	jor g0234(.dina(w_n199_0[2]),.dinb(w_n91_0[2]),.dout(n306),.clk(gclk));
	jand g0235(.dina(n306),.dinb(n305),.dout(n307),.clk(gclk));
	jand g0236(.dina(n307),.dinb(n304),.dout(n308),.clk(gclk));
	jor g0237(.dina(n308),.dinb(w_n166_1[2]),.dout(n309),.clk(gclk));
	jor g0238(.dina(w_n231_0[1]),.dinb(w_n106_0[0]),.dout(n310),.clk(gclk));
	jand g0239(.dina(n310),.dinb(w_n229_0[1]),.dout(n311),.clk(gclk));
	jand g0240(.dina(n311),.dinb(w_dff_B_ESiqQjT38_1),.dout(n312),.clk(gclk));
	jand g0241(.dina(w_n312_1[1]),.dinb(w_n196_2[0]),.dout(n313),.clk(gclk));
	jor g0242(.dina(n313),.dinb(w_n303_0[1]),.dout(n314),.clk(gclk));
	jor g0243(.dina(n314),.dinb(w_dff_B_2Ups4ZUZ1_1),.dout(n315),.clk(gclk));
	jand g0244(.dina(w_n288_1[0]),.dinb(w_G200_4[0]),.dout(n316),.clk(gclk));
	jnot g0245(.din(w_n300_0[0]),.dout(n317),.clk(gclk));
	jand g0246(.dina(w_dff_B_YUhf0cSD3_0),.dinb(w_n271_1[1]),.dout(n318),.clk(gclk));
	jor g0247(.dina(n318),.dinb(w_n298_0[0]),.dout(n319),.clk(gclk));
	jor g0248(.dina(n319),.dinb(w_n296_0[0]),.dout(n320),.clk(gclk));
	jand g0249(.dina(w_n312_1[0]),.dinb(w_G190_3[2]),.dout(n321),.clk(gclk));
	jor g0250(.dina(n321),.dinb(w_n320_0[1]),.dout(n322),.clk(gclk));
	jor g0251(.dina(n322),.dinb(w_dff_B_FItYXkBg8_1),.dout(n323),.clk(gclk));
	jand g0252(.dina(n323),.dinb(w_n315_0[1]),.dout(n324),.clk(gclk));
	jor g0253(.dina(w_n97_0[2]),.dinb(w_G33_8[0]),.dout(n325),.clk(gclk));
	jand g0254(.dina(n325),.dinb(w_n112_4[1]),.dout(n326),.clk(gclk));
	jand g0255(.dina(n326),.dinb(w_n201_0[0]),.dout(n327),.clk(gclk));
	jor g0256(.dina(n327),.dinb(w_n179_1[0]),.dout(n328),.clk(gclk));
	jor g0257(.dina(w_n328_0[1]),.dinb(w_G20_4[1]),.dout(n329),.clk(gclk));
	jand g0258(.dina(n329),.dinb(w_G107_4[0]),.dout(n330),.clk(gclk));
	jand g0259(.dina(w_n328_0[0]),.dinb(w_n270_0[0]),.dout(n331),.clk(gclk));
	jor g0260(.dina(w_dff_B_CckvPW0B8_0),.dinb(n330),.dout(n332),.clk(gclk));
	jand g0261(.dina(w_n261_0[0]),.dinb(w_G107_3[2]),.dout(n333),.clk(gclk));
	jand g0262(.dina(w_dff_B_rBOlzuRi6_0),.dinb(w_n271_1[0]),.dout(n334),.clk(gclk));
	jnot g0263(.din(w_n334_0[1]),.dout(n335),.clk(gclk));
	jand g0264(.dina(w_dff_B_0ZqnHgth1_0),.dinb(n332),.dout(n336),.clk(gclk));
	jor g0265(.dina(w_n197_0[1]),.dinb(w_n91_0[1]),.dout(n337),.clk(gclk));
	jor g0266(.dina(w_n199_0[1]),.dinb(w_n98_0[2]),.dout(n338),.clk(gclk));
	jand g0267(.dina(w_G294_3[1]),.dinb(w_G33_7[2]),.dout(n339),.clk(gclk));
	jnot g0268(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jand g0269(.dina(n340),.dinb(n338),.dout(n341),.clk(gclk));
	jand g0270(.dina(n341),.dinb(n337),.dout(n342),.clk(gclk));
	jor g0271(.dina(n342),.dinb(w_n166_1[1]),.dout(n343),.clk(gclk));
	jor g0272(.dina(w_n231_0[0]),.dinb(w_n88_0[1]),.dout(n344),.clk(gclk));
	jand g0273(.dina(n344),.dinb(w_n229_0[0]),.dout(n345),.clk(gclk));
	jand g0274(.dina(n345),.dinb(w_dff_B_Ob1JtJHk1_1),.dout(n346),.clk(gclk));
	jand g0275(.dina(w_n346_1[1]),.dinb(w_n196_1[2]),.dout(n347),.clk(gclk));
	jand g0276(.dina(w_n152_2[1]),.dinb(w_G257_0[1]),.dout(n348),.clk(gclk));
	jand g0277(.dina(w_n155_2[1]),.dinb(w_G250_0[0]),.dout(n349),.clk(gclk));
	jor g0278(.dina(w_n339_0[0]),.dinb(n349),.dout(n350),.clk(gclk));
	jor g0279(.dina(n350),.dinb(w_dff_B_lBI3HOGf2_1),.dout(n351),.clk(gclk));
	jand g0280(.dina(n351),.dinb(w_n151_2[2]),.dout(n352),.clk(gclk));
	jand g0281(.dina(w_n243_0[0]),.dinb(w_G264_0[1]),.dout(n353),.clk(gclk));
	jor g0282(.dina(n353),.dinb(w_n242_0[0]),.dout(n354),.clk(gclk));
	jor g0283(.dina(n354),.dinb(n352),.dout(n355),.clk(gclk));
	jand g0284(.dina(w_n355_1[1]),.dinb(w_n146_2[2]),.dout(n356),.clk(gclk));
	jor g0285(.dina(n356),.dinb(n347),.dout(n357),.clk(gclk));
	jor g0286(.dina(n357),.dinb(n336),.dout(n358),.clk(gclk));
	jand g0287(.dina(w_G87_3[0]),.dinb(w_n148_7[1]),.dout(n359),.clk(gclk));
	jor g0288(.dina(n359),.dinb(w_G20_4[0]),.dout(n360),.clk(gclk));
	jor g0289(.dina(n360),.dinb(w_n157_0[0]),.dout(n361),.clk(gclk));
	jand g0290(.dina(n361),.dinb(w_n189_1[1]),.dout(n362),.clk(gclk));
	jand g0291(.dina(w_n362_0[1]),.dinb(w_n112_4[0]),.dout(n363),.clk(gclk));
	jor g0292(.dina(n363),.dinb(w_n80_0[2]),.dout(n364),.clk(gclk));
	jor g0293(.dina(w_n362_0[0]),.dinb(w_n185_2[1]),.dout(n365),.clk(gclk));
	jand g0294(.dina(w_dff_B_qaOjpxk54_0),.dinb(n364),.dout(n366),.clk(gclk));
	jor g0295(.dina(w_n334_0[0]),.dinb(n366),.dout(n367),.clk(gclk));
	jor g0296(.dina(w_n355_1[0]),.dinb(w_G190_3[1]),.dout(n368),.clk(gclk));
	jor g0297(.dina(w_n346_1[0]),.dinb(w_G200_3[2]),.dout(n369),.clk(gclk));
	jand g0298(.dina(n369),.dinb(n368),.dout(n370),.clk(gclk));
	jor g0299(.dina(n370),.dinb(w_n367_0[2]),.dout(n371),.clk(gclk));
	jand g0300(.dina(w_n371_0[1]),.dinb(n358),.dout(n372),.clk(gclk));
	jand g0301(.dina(w_n372_0[1]),.dinb(w_n324_0[1]),.dout(n373),.clk(gclk));
	jand g0302(.dina(n373),.dinb(w_n279_0[1]),.dout(n374),.clk(gclk));
	jand g0303(.dina(w_n155_2[0]),.dinb(w_G232_1[0]),.dout(n375),.clk(gclk));
	jand g0304(.dina(w_n152_2[0]),.dinb(w_G238_0[2]),.dout(n376),.clk(gclk));
	jor g0305(.dina(n376),.dinb(w_n249_0[0]),.dout(n377),.clk(gclk));
	jor g0306(.dina(n377),.dinb(w_dff_B_PTmXAk1V4_1),.dout(n378),.clk(gclk));
	jand g0307(.dina(n378),.dinb(w_n151_2[1]),.dout(n379),.clk(gclk));
	jand g0308(.dina(w_n161_1[0]),.dinb(w_n149_1[2]),.dout(n380),.clk(gclk));
	jor g0309(.dina(n380),.dinb(w_G1_1[1]),.dout(n381),.clk(gclk));
	jand g0310(.dina(w_n381_0[1]),.dinb(w_n166_1[0]),.dout(n382),.clk(gclk));
	jand g0311(.dina(w_n382_1[1]),.dinb(w_G244_0[1]),.dout(n383),.clk(gclk));
	jnot g0312(.din(w_n381_0[0]),.dout(n384),.clk(gclk));
	jand g0313(.dina(n384),.dinb(w_n241_0[0]),.dout(n385),.clk(gclk));
	jor g0314(.dina(w_n385_1[1]),.dinb(n383),.dout(n386),.clk(gclk));
	jor g0315(.dina(n386),.dinb(n379),.dout(n387),.clk(gclk));
	jand g0316(.dina(w_n387_1[1]),.dinb(w_n146_2[1]),.dout(n388),.clk(gclk));
	jnot g0317(.din(n388),.dout(n389),.clk(gclk));
	jand g0318(.dina(w_G87_2[2]),.dinb(w_G33_7[1]),.dout(n390),.clk(gclk));
	jand g0319(.dina(w_G58_4[2]),.dinb(w_n148_7[0]),.dout(n391),.clk(gclk));
	jor g0320(.dina(n391),.dinb(w_G20_3[2]),.dout(n392),.clk(gclk));
	jor g0321(.dina(n392),.dinb(w_n390_0[1]),.dout(n393),.clk(gclk));
	jor g0322(.dina(w_G77_4[1]),.dinb(w_n112_3[2]),.dout(n394),.clk(gclk));
	jand g0323(.dina(w_dff_B_2tWgEd0F4_0),.dinb(w_n189_1[0]),.dout(n395),.clk(gclk));
	jand g0324(.dina(n395),.dinb(n393),.dout(n396),.clk(gclk));
	jand g0325(.dina(w_n185_2[0]),.dinb(w_n72_0[2]),.dout(n397),.clk(gclk));
	jand g0326(.dina(w_n269_1[1]),.dinb(w_G77_4[0]),.dout(n398),.clk(gclk));
	jand g0327(.dina(w_dff_B_3kuTcEeI7_0),.dinb(w_n271_0[2]),.dout(n399),.clk(gclk));
	jor g0328(.dina(n399),.dinb(w_dff_B_HvNdSAf63_1),.dout(n400),.clk(gclk));
	jor g0329(.dina(n400),.dinb(w_dff_B_StYp0G5t7_1),.dout(n401),.clk(gclk));
	jor g0330(.dina(w_n387_1[0]),.dinb(w_G179_2[1]),.dout(n402),.clk(gclk));
	jand g0331(.dina(n402),.dinb(w_n401_0[2]),.dout(n403),.clk(gclk));
	jand g0332(.dina(n403),.dinb(n389),.dout(n404),.clk(gclk));
	jnot g0333(.din(w_n404_0[2]),.dout(n405),.clk(gclk));
	jand g0334(.dina(w_n387_0[2]),.dinb(w_G200_3[1]),.dout(n406),.clk(gclk));
	jnot g0335(.din(w_G190_3[0]),.dout(n407),.clk(gclk));
	jor g0336(.dina(w_n387_0[1]),.dinb(w_n407_2[1]),.dout(n408),.clk(gclk));
	jnot g0337(.din(n408),.dout(n409),.clk(gclk));
	jor g0338(.dina(n409),.dinb(w_n401_0[1]),.dout(n410),.clk(gclk));
	jor g0339(.dina(n410),.dinb(w_dff_B_NL5dvISo6_1),.dout(n411),.clk(gclk));
	jand g0340(.dina(n411),.dinb(w_n405_0[1]),.dout(n412),.clk(gclk));
	jand g0341(.dina(w_n155_1[2]),.dinb(w_G226_1[0]),.dout(n413),.clk(gclk));
	jand g0342(.dina(w_n152_1[2]),.dinb(w_G232_0[2]),.dout(n414),.clk(gclk));
	jor g0343(.dina(n414),.dinb(w_n172_0[0]),.dout(n415),.clk(gclk));
	jor g0344(.dina(n415),.dinb(w_dff_B_gnYSGXxX9_1),.dout(n416),.clk(gclk));
	jand g0345(.dina(n416),.dinb(w_n151_2[0]),.dout(n417),.clk(gclk));
	jand g0346(.dina(w_n382_1[0]),.dinb(w_G238_0[1]),.dout(n418),.clk(gclk));
	jor g0347(.dina(n418),.dinb(w_n385_1[0]),.dout(n419),.clk(gclk));
	jor g0348(.dina(n419),.dinb(n417),.dout(n420),.clk(gclk));
	jand g0349(.dina(w_n420_1[1]),.dinb(w_n146_2[0]),.dout(n421),.clk(gclk));
	jnot g0350(.din(n421),.dout(n422),.clk(gclk));
	jand g0351(.dina(w_n269_1[0]),.dinb(w_G68_4[1]),.dout(n423),.clk(gclk));
	jand g0352(.dina(w_dff_B_aqhacGvo0_0),.dinb(w_n271_0[1]),.dout(n424),.clk(gclk));
	jand g0353(.dina(w_n148_6[2]),.dinb(w_n114_0[2]),.dout(n425),.clk(gclk));
	jnot g0354(.din(w_n425_1[2]),.dout(n426),.clk(gclk));
	jand g0355(.dina(w_n426_0[1]),.dinb(w_n85_0[0]),.dout(n427),.clk(gclk));
	jor g0356(.dina(n427),.dinb(w_n185_1[2]),.dout(n428),.clk(gclk));
	jand g0357(.dina(n428),.dinb(w_n75_0[2]),.dout(n429),.clk(gclk));
	jand g0358(.dina(w_G77_3[2]),.dinb(w_G33_7[0]),.dout(n430),.clk(gclk));
	jand g0359(.dina(w_G50_4[2]),.dinb(w_n148_6[1]),.dout(n431),.clk(gclk));
	jor g0360(.dina(n431),.dinb(w_n430_0[1]),.dout(n432),.clk(gclk));
	jand g0361(.dina(n432),.dinb(w_n112_3[1]),.dout(n433),.clk(gclk));
	jand g0362(.dina(n433),.dinb(w_n189_0[2]),.dout(n434),.clk(gclk));
	jor g0363(.dina(w_dff_B_GJ14VP5H9_0),.dinb(n429),.dout(n435),.clk(gclk));
	jor g0364(.dina(n435),.dinb(w_dff_B_ofPosrps6_1),.dout(n436),.clk(gclk));
	jor g0365(.dina(w_n420_1[0]),.dinb(w_G179_2[0]),.dout(n437),.clk(gclk));
	jand g0366(.dina(n437),.dinb(w_n436_0[2]),.dout(n438),.clk(gclk));
	jand g0367(.dina(n438),.dinb(n422),.dout(n439),.clk(gclk));
	jnot g0368(.din(w_n439_1[1]),.dout(n440),.clk(gclk));
	jand g0369(.dina(w_n420_0[2]),.dinb(w_G200_3[0]),.dout(n441),.clk(gclk));
	jor g0370(.dina(w_n420_0[1]),.dinb(w_n407_2[0]),.dout(n442),.clk(gclk));
	jnot g0371(.din(n442),.dout(n443),.clk(gclk));
	jor g0372(.dina(n443),.dinb(w_n436_0[1]),.dout(n444),.clk(gclk));
	jor g0373(.dina(n444),.dinb(w_dff_B_zINCodE96_1),.dout(n445),.clk(gclk));
	jand g0374(.dina(w_n445_0[1]),.dinb(n440),.dout(n446),.clk(gclk));
	jand g0375(.dina(w_n446_0[1]),.dinb(w_n412_0[1]),.dout(n447),.clk(gclk));
	jand g0376(.dina(w_n152_1[1]),.dinb(w_G223_0[1]),.dout(n448),.clk(gclk));
	jand g0377(.dina(w_n155_1[1]),.dinb(w_dff_B_PRok0oYL4_1),.dout(n449),.clk(gclk));
	jor g0378(.dina(n449),.dinb(w_n430_0[0]),.dout(n450),.clk(gclk));
	jor g0379(.dina(n450),.dinb(w_dff_B_0Azvf9Fl7_1),.dout(n451),.clk(gclk));
	jand g0380(.dina(n451),.dinb(w_n151_1[2]),.dout(n452),.clk(gclk));
	jand g0381(.dina(w_n382_0[2]),.dinb(w_G226_0[2]),.dout(n453),.clk(gclk));
	jor g0382(.dina(n453),.dinb(w_n385_0[2]),.dout(n454),.clk(gclk));
	jor g0383(.dina(n454),.dinb(n452),.dout(n455),.clk(gclk));
	jand g0384(.dina(w_n455_0[2]),.dinb(w_n146_1[2]),.dout(n456),.clk(gclk));
	jand g0385(.dina(w_n269_0[2]),.dinb(w_G50_4[1]),.dout(n457),.clk(gclk));
	jnot g0386(.din(n457),.dout(n458),.clk(gclk));
	jor g0387(.dina(n458),.dinb(w_n190_0[2]),.dout(n459),.clk(gclk));
	jor g0388(.dina(w_n77_0[0]),.dinb(w_n112_3[0]),.dout(n460),.clk(gclk));
	jnot g0389(.din(w_G150_3[1]),.dout(n461),.clk(gclk));
	jand g0390(.dina(w_n148_6[0]),.dinb(w_n112_2[2]),.dout(n462),.clk(gclk));
	jnot g0391(.din(w_n462_0[2]),.dout(n463),.clk(gclk));
	jor g0392(.dina(n463),.dinb(w_dff_B_E8v5SAeS1_1),.dout(n464),.clk(gclk));
	jand g0393(.dina(w_G33_6[2]),.dinb(w_n112_2[1]),.dout(n465),.clk(gclk));
	jand g0394(.dina(w_n465_0[1]),.dinb(w_G58_4[1]),.dout(n466),.clk(gclk));
	jnot g0395(.din(n466),.dout(n467),.clk(gclk));
	jand g0396(.dina(n467),.dinb(n464),.dout(n468),.clk(gclk));
	jand g0397(.dina(n468),.dinb(w_dff_B_pHiKbyQ42_1),.dout(n469),.clk(gclk));
	jor g0398(.dina(n469),.dinb(w_n179_0[2]),.dout(n470),.clk(gclk));
	jand g0399(.dina(w_n185_1[1]),.dinb(w_n73_2[0]),.dout(n471),.clk(gclk));
	jnot g0400(.din(n471),.dout(n472),.clk(gclk));
	jand g0401(.dina(w_dff_B_F9tTvFqz1_0),.dinb(n470),.dout(n473),.clk(gclk));
	jand g0402(.dina(n473),.dinb(w_dff_B_Mpdsynv86_1),.dout(n474),.clk(gclk));
	jnot g0403(.din(w_n455_0[1]),.dout(n475),.clk(gclk));
	jand g0404(.dina(w_n475_0[1]),.dinb(w_n196_1[1]),.dout(n476),.clk(gclk));
	jor g0405(.dina(n476),.dinb(w_n474_0[1]),.dout(n477),.clk(gclk));
	jor g0406(.dina(n477),.dinb(w_dff_B_zWcwDe4Y2_1),.dout(n478),.clk(gclk));
	jnot g0407(.din(w_n474_0[0]),.dout(n479),.clk(gclk));
	jand g0408(.dina(w_n475_0[0]),.dinb(w_G190_2[2]),.dout(n480),.clk(gclk));
	jand g0409(.dina(w_n455_0[0]),.dinb(w_G200_2[2]),.dout(n481),.clk(gclk));
	jor g0410(.dina(w_dff_B_npcdkGxv1_0),.dinb(n480),.dout(n482),.clk(gclk));
	jor g0411(.dina(n482),.dinb(w_n479_0[1]),.dout(n483),.clk(gclk));
	jand g0412(.dina(w_n483_0[1]),.dinb(w_n478_0[1]),.dout(n484),.clk(gclk));
	jand g0413(.dina(w_n152_1[0]),.dinb(w_G226_0[1]),.dout(n485),.clk(gclk));
	jand g0414(.dina(w_n155_1[0]),.dinb(w_G223_0[0]),.dout(n486),.clk(gclk));
	jor g0415(.dina(n486),.dinb(w_n390_0[0]),.dout(n487),.clk(gclk));
	jor g0416(.dina(n487),.dinb(w_dff_B_x12Dlwfq6_1),.dout(n488),.clk(gclk));
	jand g0417(.dina(n488),.dinb(w_n151_1[1]),.dout(n489),.clk(gclk));
	jand g0418(.dina(w_n382_0[1]),.dinb(w_G232_0[1]),.dout(n490),.clk(gclk));
	jor g0419(.dina(n490),.dinb(w_n385_0[1]),.dout(n491),.clk(gclk));
	jor g0420(.dina(n491),.dinb(n489),.dout(n492),.clk(gclk));
	jand g0421(.dina(w_n492_0[2]),.dinb(w_n146_1[1]),.dout(n493),.clk(gclk));
	jand g0422(.dina(w_n269_0[1]),.dinb(w_G58_4[0]),.dout(n494),.clk(gclk));
	jnot g0423(.din(n494),.dout(n495),.clk(gclk));
	jor g0424(.dina(n495),.dinb(w_n190_0[1]),.dout(n496),.clk(gclk));
	jor g0425(.dina(w_n137_0[1]),.dinb(w_n112_2[0]),.dout(n497),.clk(gclk));
	jand g0426(.dina(w_n462_0[1]),.dinb(w_G159_3[2]),.dout(n498),.clk(gclk));
	jand g0427(.dina(w_n465_0[0]),.dinb(w_G68_4[0]),.dout(n499),.clk(gclk));
	jor g0428(.dina(n499),.dinb(n498),.dout(n500),.clk(gclk));
	jnot g0429(.din(n500),.dout(n501),.clk(gclk));
	jand g0430(.dina(n501),.dinb(w_dff_B_B7COo6eY8_1),.dout(n502),.clk(gclk));
	jor g0431(.dina(n502),.dinb(w_n179_0[1]),.dout(n503),.clk(gclk));
	jand g0432(.dina(w_n185_1[0]),.dinb(w_n74_0[2]),.dout(n504),.clk(gclk));
	jnot g0433(.din(n504),.dout(n505),.clk(gclk));
	jand g0434(.dina(w_dff_B_yOxgi82s2_0),.dinb(n503),.dout(n506),.clk(gclk));
	jand g0435(.dina(n506),.dinb(w_dff_B_cshKiaOQ2_1),.dout(n507),.clk(gclk));
	jnot g0436(.din(w_n492_0[1]),.dout(n508),.clk(gclk));
	jand g0437(.dina(w_n508_0[1]),.dinb(w_n196_1[0]),.dout(n509),.clk(gclk));
	jor g0438(.dina(n509),.dinb(w_n507_0[1]),.dout(n510),.clk(gclk));
	jor g0439(.dina(n510),.dinb(w_dff_B_29U80Tha0_1),.dout(n511),.clk(gclk));
	jnot g0440(.din(w_n507_0[0]),.dout(n512),.clk(gclk));
	jand g0441(.dina(w_n508_0[0]),.dinb(w_G190_2[1]),.dout(n513),.clk(gclk));
	jand g0442(.dina(w_n492_0[0]),.dinb(w_G200_2[1]),.dout(n514),.clk(gclk));
	jor g0443(.dina(w_dff_B_ynRXNWFL6_0),.dinb(n513),.dout(n515),.clk(gclk));
	jor g0444(.dina(n515),.dinb(w_n512_0[1]),.dout(n516),.clk(gclk));
	jand g0445(.dina(w_n516_0[1]),.dinb(w_n511_0[1]),.dout(n517),.clk(gclk));
	jand g0446(.dina(w_n517_0[1]),.dinb(w_n484_0[1]),.dout(n518),.clk(gclk));
	jand g0447(.dina(n518),.dinb(n447),.dout(n519),.clk(gclk));
	jand g0448(.dina(w_n519_1[2]),.dinb(w_n374_0[1]),.dout(w_dff_A_U1r5udv24_2),.clk(gclk));
	jor g0449(.dina(w_n355_0[2]),.dinb(w_G179_1[2]),.dout(n521),.clk(gclk));
	jor g0450(.dina(w_n346_0[2]),.dinb(w_G169_1[0]),.dout(n522),.clk(gclk));
	jand g0451(.dina(n522),.dinb(n521),.dout(n523),.clk(gclk));
	jand g0452(.dina(w_n523_0[1]),.dinb(w_n367_0[1]),.dout(n524),.clk(gclk));
	jor g0453(.dina(w_n312_0[2]),.dinb(w_G169_0[2]),.dout(n525),.clk(gclk));
	jor g0454(.dina(w_n288_0[2]),.dinb(w_G179_1[1]),.dout(n526),.clk(gclk));
	jand g0455(.dina(n526),.dinb(w_n320_0[0]),.dout(n527),.clk(gclk));
	jand g0456(.dina(n527),.dinb(w_dff_B_MbbpWLVQ2_1),.dout(n528),.clk(gclk));
	jand g0457(.dina(w_n371_0[0]),.dinb(w_n528_0[1]),.dout(n529),.clk(gclk));
	jor g0458(.dina(n529),.dinb(w_n524_0[1]),.dout(n530),.clk(gclk));
	jand g0459(.dina(n530),.dinb(w_n279_0[0]),.dout(n531),.clk(gclk));
	jnot g0460(.din(w_n213_0[0]),.dout(n532),.clk(gclk));
	jand g0461(.dina(w_n246_0[2]),.dinb(w_G169_0[1]),.dout(n533),.clk(gclk));
	jand g0462(.dina(w_n234_0[0]),.dinb(w_G179_1[0]),.dout(n534),.clk(gclk));
	jor g0463(.dina(w_n534_0[1]),.dinb(n533),.dout(n535),.clk(gclk));
	jand g0464(.dina(w_n274_0[1]),.dinb(n535),.dout(n536),.clk(gclk));
	jand g0465(.dina(w_n536_0[2]),.dinb(w_n218_0[0]),.dout(n537),.clk(gclk));
	jor g0466(.dina(n537),.dinb(w_n532_0[1]),.dout(n538),.clk(gclk));
	jor g0467(.dina(w_dff_B_Se6rDN258_0),.dinb(n531),.dout(n539),.clk(gclk));
	jand g0468(.dina(w_n539_0[1]),.dinb(w_n519_1[1]),.dout(n540),.clk(gclk));
	jnot g0469(.din(w_n478_0[0]),.dout(n541),.clk(gclk));
	jnot g0470(.din(w_n511_0[0]),.dout(n542),.clk(gclk));
	jor g0471(.dina(w_n439_1[0]),.dinb(w_n404_0[1]),.dout(n543),.clk(gclk));
	jand g0472(.dina(w_n543_0[1]),.dinb(w_n445_0[0]),.dout(n544),.clk(gclk));
	jor g0473(.dina(n544),.dinb(w_n542_0[2]),.dout(n545),.clk(gclk));
	jand g0474(.dina(n545),.dinb(w_n516_0[0]),.dout(n546),.clk(gclk));
	jor g0475(.dina(n546),.dinb(w_n541_0[1]),.dout(n547),.clk(gclk));
	jand g0476(.dina(n547),.dinb(w_n483_0[0]),.dout(n548),.clk(gclk));
	jor g0477(.dina(w_n548_0[2]),.dinb(w_dff_B_ldRFVe202_1),.dout(w_dff_A_Rrj7Q0eY0_2),.clk(gclk));
	jand g0478(.dina(w_n112_1[2]),.dinb(w_G13_0[1]),.dout(n550),.clk(gclk));
	jand g0479(.dina(w_G213_0[2]),.dinb(w_n113_1[2]),.dout(n551),.clk(gclk));
	jand g0480(.dina(n551),.dinb(w_n550_0[1]),.dout(n552),.clk(gclk));
	jand g0481(.dina(w_n552_1[1]),.dinb(w_G343_0[1]),.dout(n553),.clk(gclk));
	jnot g0482(.din(w_n553_2[2]),.dout(n554),.clk(gclk));
	jand g0483(.dina(w_n554_3[2]),.dinb(w_n524_0[0]),.dout(n555),.clk(gclk));
	jand g0484(.dina(w_n554_3[1]),.dinb(w_n528_0[0]),.dout(n556),.clk(gclk));
	jand g0485(.dina(w_n553_2[1]),.dinb(w_n367_0[0]),.dout(n557),.clk(gclk));
	jnot g0486(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jand g0487(.dina(n558),.dinb(w_n372_0[0]),.dout(n559),.clk(gclk));
	jand g0488(.dina(w_n557_0[0]),.dinb(w_n523_0[0]),.dout(n560),.clk(gclk));
	jor g0489(.dina(w_dff_B_Po7JYX890_0),.dinb(n559),.dout(n561),.clk(gclk));
	jand g0490(.dina(w_n561_0[2]),.dinb(w_n556_0[1]),.dout(n562),.clk(gclk));
	jor g0491(.dina(n562),.dinb(w_dff_B_wzSXzrlF4_1),.dout(n563),.clk(gclk));
	jnot g0492(.din(w_n561_0[1]),.dout(n564),.clk(gclk));
	jnot g0493(.din(w_G330_0[1]),.dout(n565),.clk(gclk));
	jnot g0494(.din(w_n324_0[0]),.dout(n566),.clk(gclk));
	jor g0495(.dina(w_n554_3[0]),.dinb(w_n303_0[0]),.dout(n567),.clk(gclk));
	jnot g0496(.din(w_n567_0[1]),.dout(n568),.clk(gclk));
	jor g0497(.dina(w_dff_B_hlze2NKO0_0),.dinb(n566),.dout(n569),.clk(gclk));
	jor g0498(.dina(w_n567_0[0]),.dinb(w_n315_0[0]),.dout(n570),.clk(gclk));
	jand g0499(.dina(w_dff_B_6MOx5bXI0_0),.dinb(n569),.dout(n571),.clk(gclk));
	jor g0500(.dina(w_n571_0[2]),.dinb(w_n565_0[1]),.dout(n572),.clk(gclk));
	jor g0501(.dina(w_n572_0[2]),.dinb(w_n564_0[1]),.dout(n573),.clk(gclk));
	jnot g0502(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jor g0503(.dina(n574),.dinb(w_n563_0[2]),.dout(w_dff_A_ePxRogil5_2),.clk(gclk));
	jand g0504(.dina(w_n554_2[2]),.dinb(w_n539_0[0]),.dout(n576),.clk(gclk));
	jor g0505(.dina(w_n553_2[0]),.dinb(w_n374_0[0]),.dout(n577),.clk(gclk));
	jand g0506(.dina(w_n346_0[1]),.dinb(w_n210_0[0]),.dout(n578),.clk(gclk));
	jand g0507(.dina(n578),.dinb(w_n312_0[1]),.dout(n579),.clk(gclk));
	jand g0508(.dina(n579),.dinb(w_n534_0[0]),.dout(n580),.clk(gclk));
	jand g0509(.dina(w_n288_0[1]),.dinb(w_n196_0[2]),.dout(n581),.clk(gclk));
	jand g0510(.dina(w_n355_0[1]),.dinb(w_n246_0[1]),.dout(n582),.clk(gclk));
	jand g0511(.dina(n582),.dinb(w_n170_0[0]),.dout(n583),.clk(gclk));
	jand g0512(.dina(n583),.dinb(w_dff_B_lWHQMiHx3_1),.dout(n584),.clk(gclk));
	jor g0513(.dina(n584),.dinb(w_n554_2[1]),.dout(n585),.clk(gclk));
	jor g0514(.dina(n585),.dinb(w_dff_B_rmTxIiOP8_1),.dout(n586),.clk(gclk));
	jand g0515(.dina(n586),.dinb(w_G330_0[0]),.dout(n587),.clk(gclk));
	jand g0516(.dina(w_dff_B_Rk1Okfz02_0),.dinb(n577),.dout(n588),.clk(gclk));
	jor g0517(.dina(w_n588_1[1]),.dinb(w_n576_1[1]),.dout(n589),.clk(gclk));
	jand g0518(.dina(w_n589_1[2]),.dinb(w_n113_1[1]),.dout(n590),.clk(gclk));
	jand g0519(.dina(w_n122_1[0]),.dinb(w_n149_1[1]),.dout(n591),.clk(gclk));
	jnot g0520(.din(w_n591_1[1]),.dout(n592),.clk(gclk));
	jand g0521(.dina(w_n180_0[0]),.dinb(w_n105_1[0]),.dout(n593),.clk(gclk));
	jand g0522(.dina(w_n593_0[2]),.dinb(w_G1_1[0]),.dout(n594),.clk(gclk));
	jand g0523(.dina(n594),.dinb(w_n592_2[1]),.dout(n595),.clk(gclk));
	jand g0524(.dina(w_n591_1[0]),.dinb(w_n118_0[1]),.dout(n596),.clk(gclk));
	jor g0525(.dina(w_dff_B_Meiy2dWM6_0),.dinb(n595),.dout(n597),.clk(gclk));
	jor g0526(.dina(w_dff_B_FFN7T7lW1_0),.dinb(n590),.dout(w_dff_A_FcBxUslg3_2),.clk(gclk));
	jand g0527(.dina(w_n571_0[1]),.dinb(w_n565_0[0]),.dout(n599),.clk(gclk));
	jnot g0528(.din(n599),.dout(n600),.clk(gclk));
	jand g0529(.dina(w_n550_0[0]),.dinb(w_G45_1[0]),.dout(n601),.clk(gclk));
	jor g0530(.dina(n601),.dinb(w_n113_1[0]),.dout(n602),.clk(gclk));
	jnot g0531(.din(w_n602_0[1]),.dout(n603),.clk(gclk));
	jand g0532(.dina(w_n603_2[1]),.dinb(w_n592_2[0]),.dout(n604),.clk(gclk));
	jnot g0533(.din(w_n604_2[1]),.dout(n605),.clk(gclk));
	jand g0534(.dina(w_n605_1[2]),.dinb(w_n572_0[1]),.dout(n606),.clk(gclk));
	jand g0535(.dina(n606),.dinb(n600),.dout(n607),.clk(gclk));
	jand g0536(.dina(w_n462_0[0]),.dinb(w_n114_0[1]),.dout(n608),.clk(gclk));
	jand g0537(.dina(w_n608_1[2]),.dinb(w_n571_0[0]),.dout(n609),.clk(gclk));
	jnot g0538(.din(n609),.dout(n610),.clk(gclk));
	jand g0539(.dina(w_n146_1[0]),.dinb(w_G20_3[1]),.dout(n611),.clk(gclk));
	jor g0540(.dina(n611),.dinb(w_n115_0[1]),.dout(n612),.clk(gclk));
	jand g0541(.dina(w_G179_0[2]),.dinb(w_G20_3[0]),.dout(n613),.clk(gclk));
	jnot g0542(.din(w_n613_1[1]),.dout(n614),.clk(gclk));
	jand g0543(.dina(w_G200_2[0]),.dinb(w_G20_2[2]),.dout(n615),.clk(gclk));
	jand g0544(.dina(w_n615_0[1]),.dinb(n614),.dout(n616),.clk(gclk));
	jand g0545(.dina(w_n616_0[1]),.dinb(w_G190_2[0]),.dout(n617),.clk(gclk));
	jand g0546(.dina(w_n617_6[1]),.dinb(w_G303_2[1]),.dout(n618),.clk(gclk));
	jand g0547(.dina(w_n407_1[2]),.dinb(w_G20_2[1]),.dout(n619),.clk(gclk));
	jnot g0548(.din(w_n619_0[1]),.dout(n620),.clk(gclk));
	jor g0549(.dina(w_n615_0[0]),.dinb(w_n613_1[0]),.dout(n621),.clk(gclk));
	jnot g0550(.din(n621),.dout(n622),.clk(gclk));
	jand g0551(.dina(w_n622_0[1]),.dinb(n620),.dout(n623),.clk(gclk));
	jand g0552(.dina(w_n623_5[1]),.dinb(w_G294_3[0]),.dout(n624),.clk(gclk));
	jnot g0553(.din(w_G200_1[2]),.dout(n625),.clk(gclk));
	jand g0554(.dina(w_n613_0[2]),.dinb(n625),.dout(n626),.clk(gclk));
	jand g0555(.dina(w_n626_0[1]),.dinb(w_G190_1[2]),.dout(n627),.clk(gclk));
	jand g0556(.dina(w_n627_7[1]),.dinb(w_G322_0[2]),.dout(n628),.clk(gclk));
	jor g0557(.dina(w_dff_B_iv6e9eD24_0),.dinb(n624),.dout(n629),.clk(gclk));
	jor g0558(.dina(n629),.dinb(w_dff_B_P6h9LSyK6_1),.dout(n630),.clk(gclk));
	jand g0559(.dina(w_n622_0[0]),.dinb(w_n619_0[0]),.dout(n631),.clk(gclk));
	jand g0560(.dina(w_n631_7[1]),.dinb(w_dff_B_X6hvEvIb3_1),.dout(n632),.clk(gclk));
	jor g0561(.dina(n632),.dinb(w_n148_5[2]),.dout(n633),.clk(gclk));
	jand g0562(.dina(w_n616_0[0]),.dinb(w_n407_1[1]),.dout(n634),.clk(gclk));
	jand g0563(.dina(w_n634_4[1]),.dinb(w_G283_3[1]),.dout(n635),.clk(gclk));
	jand g0564(.dina(w_n626_0[0]),.dinb(w_n407_1[0]),.dout(n636),.clk(gclk));
	jand g0565(.dina(w_n636_7[1]),.dinb(w_G311_1[2]),.dout(n637),.clk(gclk));
	jor g0566(.dina(w_dff_B_ueObpH249_0),.dinb(n635),.dout(n638),.clk(gclk));
	jand g0567(.dina(w_n613_0[1]),.dinb(w_G200_1[1]),.dout(n639),.clk(gclk));
	jand g0568(.dina(w_n639_0[1]),.dinb(w_G190_1[1]),.dout(n640),.clk(gclk));
	jand g0569(.dina(w_n640_7[1]),.dinb(w_G326_0[1]),.dout(n641),.clk(gclk));
	jand g0570(.dina(w_n639_0[0]),.dinb(w_n407_0[2]),.dout(n642),.clk(gclk));
	jand g0571(.dina(w_n642_7[1]),.dinb(w_G317_1[1]),.dout(n643),.clk(gclk));
	jor g0572(.dina(n643),.dinb(n641),.dout(n644),.clk(gclk));
	jor g0573(.dina(w_dff_B_R2fQozyq6_0),.dinb(n638),.dout(n645),.clk(gclk));
	jor g0574(.dina(n645),.dinb(w_dff_B_grn3rGDj5_1),.dout(n646),.clk(gclk));
	jor g0575(.dina(n646),.dinb(w_dff_B_28z0T09I2_1),.dout(n647),.clk(gclk));
	jand g0576(.dina(w_n631_7[0]),.dinb(w_G159_3[1]),.dout(n648),.clk(gclk));
	jand g0577(.dina(w_n640_7[0]),.dinb(w_G50_4[0]),.dout(n649),.clk(gclk));
	jand g0578(.dina(w_n642_7[0]),.dinb(w_G68_3[2]),.dout(n650),.clk(gclk));
	jor g0579(.dina(n650),.dinb(n649),.dout(n651),.clk(gclk));
	jor g0580(.dina(n651),.dinb(n648),.dout(n652),.clk(gclk));
	jnot g0581(.din(n652),.dout(n653),.clk(gclk));
	jand g0582(.dina(w_n617_6[0]),.dinb(w_G87_2[1]),.dout(n654),.clk(gclk));
	jnot g0583(.din(w_n654_0[1]),.dout(n655),.clk(gclk));
	jand g0584(.dina(n655),.dinb(w_n148_5[1]),.dout(n656),.clk(gclk));
	jand g0585(.dina(w_n634_4[0]),.dinb(w_G107_3[1]),.dout(n657),.clk(gclk));
	jand g0586(.dina(w_n636_7[0]),.dinb(w_G77_3[1]),.dout(n658),.clk(gclk));
	jor g0587(.dina(w_dff_B_3b1YSCjC9_0),.dinb(w_n657_0[1]),.dout(n659),.clk(gclk));
	jand g0588(.dina(w_n627_7[0]),.dinb(w_G58_3[2]),.dout(n660),.clk(gclk));
	jand g0589(.dina(w_n623_5[0]),.dinb(w_G97_3[1]),.dout(n661),.clk(gclk));
	jor g0590(.dina(w_n661_0[1]),.dinb(w_dff_B_KEhFo1TO7_1),.dout(n662),.clk(gclk));
	jor g0591(.dina(n662),.dinb(n659),.dout(n663),.clk(gclk));
	jnot g0592(.din(n663),.dout(n664),.clk(gclk));
	jand g0593(.dina(n664),.dinb(w_dff_B_x8aIJJoV5_1),.dout(n665),.clk(gclk));
	jand g0594(.dina(n665),.dinb(w_dff_B_vOi2AvAE7_1),.dout(n666),.clk(gclk));
	jnot g0595(.din(n666),.dout(n667),.clk(gclk));
	jand g0596(.dina(n667),.dinb(w_dff_B_zPnQWszI8_1),.dout(n668),.clk(gclk));
	jor g0597(.dina(n668),.dinb(w_n612_4[1]),.dout(n669),.clk(gclk));
	jnot g0598(.din(w_n608_1[1]),.dout(n670),.clk(gclk));
	jand g0599(.dina(w_n612_4[0]),.dinb(n670),.dout(n671),.clk(gclk));
	jnot g0600(.din(n671),.dout(n672),.clk(gclk));
	jand g0601(.dina(w_n140_0[0]),.dinb(w_G45_0[2]),.dout(n673),.clk(gclk));
	jand g0602(.dina(w_n118_0[0]),.dinb(w_n161_0[2]),.dout(n674),.clk(gclk));
	jand g0603(.dina(w_n122_0[2]),.dinb(w_G33_6[1]),.dout(n675),.clk(gclk));
	jnot g0604(.din(w_n675_0[2]),.dout(n676),.clk(gclk));
	jor g0605(.dina(w_n676_0[1]),.dinb(n674),.dout(n677),.clk(gclk));
	jor g0606(.dina(n677),.dinb(w_dff_B_LvqtFccj9_1),.dout(n678),.clk(gclk));
	jand g0607(.dina(w_n123_1[1]),.dinb(w_n105_0[2]),.dout(n679),.clk(gclk));
	jand g0608(.dina(w_n122_0[1]),.dinb(w_n148_5[0]),.dout(n680),.clk(gclk));
	jand g0609(.dina(w_n680_0[1]),.dinb(w_G355_0),.dout(n681),.clk(gclk));
	jor g0610(.dina(n681),.dinb(w_dff_B_ni6NVzVi8_1),.dout(n682),.clk(gclk));
	jnot g0611(.din(n682),.dout(n683),.clk(gclk));
	jand g0612(.dina(n683),.dinb(w_dff_B_7n2j4Y9q1_1),.dout(n684),.clk(gclk));
	jor g0613(.dina(n684),.dinb(w_n672_1[1]),.dout(n685),.clk(gclk));
	jand g0614(.dina(n685),.dinb(w_n604_2[0]),.dout(n686),.clk(gclk));
	jand g0615(.dina(w_dff_B_9ylm8g6g4_0),.dinb(n669),.dout(n687),.clk(gclk));
	jand g0616(.dina(w_dff_B_B7tUwYuz5_0),.dinb(n610),.dout(n688),.clk(gclk));
	jor g0617(.dina(n688),.dinb(n607),.dout(G396_fa_),.clk(gclk));
	jnot g0618(.din(w_n588_1[0]),.dout(n690),.clk(gclk));
	jnot g0619(.din(w_n401_0[0]),.dout(n691),.clk(gclk));
	jor g0620(.dina(w_n554_2[0]),.dinb(n691),.dout(n692),.clk(gclk));
	jand g0621(.dina(w_n692_0[1]),.dinb(w_n412_0[0]),.dout(n693),.clk(gclk));
	jor g0622(.dina(w_n692_0[0]),.dinb(w_n405_0[0]),.dout(n694),.clk(gclk));
	jnot g0623(.din(n694),.dout(n695),.clk(gclk));
	jor g0624(.dina(n695),.dinb(n693),.dout(n696),.clk(gclk));
	jxor g0625(.dina(w_n696_1[2]),.dinb(w_n576_1[0]),.dout(n697),.clk(gclk));
	jnot g0626(.din(n697),.dout(n698),.clk(gclk));
	jand g0627(.dina(n698),.dinb(w_dff_B_RGswLtgJ5_1),.dout(n699),.clk(gclk));
	jor g0628(.dina(w_n991_0[2]),.dinb(w_n604_1[2]),.dout(n701),.clk(gclk));
	jor g0629(.dina(w_dff_B_nKnuInHT5_0),.dinb(n699),.dout(n702),.clk(gclk));
	jnot g0630(.din(w_n696_1[1]),.dout(n703),.clk(gclk));
	jand g0631(.dina(n703),.dinb(w_n425_1[1]),.dout(n704),.clk(gclk));
	jnot g0632(.din(n704),.dout(n705),.clk(gclk));
	jand g0633(.dina(w_n631_6[2]),.dinb(w_G132_1[1]),.dout(n706),.clk(gclk));
	jand g0634(.dina(w_n623_4[2]),.dinb(w_G58_3[1]),.dout(n707),.clk(gclk));
	jand g0635(.dina(w_n642_6[2]),.dinb(w_G150_3[0]),.dout(n708),.clk(gclk));
	jor g0636(.dina(w_dff_B_NxTT5afB0_0),.dinb(n707),.dout(n709),.clk(gclk));
	jor g0637(.dina(n709),.dinb(w_dff_B_qnbmHtnG0_1),.dout(n710),.clk(gclk));
	jand g0638(.dina(w_n617_5[2]),.dinb(w_G50_3[2]),.dout(n711),.clk(gclk));
	jor g0639(.dina(n711),.dinb(w_G33_6[0]),.dout(n712),.clk(gclk));
	jand g0640(.dina(w_n636_6[2]),.dinb(w_G159_3[0]),.dout(n713),.clk(gclk));
	jand g0641(.dina(w_n627_6[2]),.dinb(w_G143_2[1]),.dout(n714),.clk(gclk));
	jor g0642(.dina(n714),.dinb(n713),.dout(n715),.clk(gclk));
	jand g0643(.dina(w_n640_6[2]),.dinb(w_G137_1[2]),.dout(n716),.clk(gclk));
	jand g0644(.dina(w_n634_3[2]),.dinb(w_G68_3[1]),.dout(n717),.clk(gclk));
	jor g0645(.dina(w_n717_0[1]),.dinb(w_dff_B_OWwWer5e5_1),.dout(n718),.clk(gclk));
	jor g0646(.dina(n718),.dinb(w_dff_B_JdtGa10D5_1),.dout(n719),.clk(gclk));
	jor g0647(.dina(n719),.dinb(w_dff_B_uc1cmXy18_1),.dout(n720),.clk(gclk));
	jor g0648(.dina(n720),.dinb(w_dff_B_xjOizQFs3_1),.dout(n721),.clk(gclk));
	jand g0649(.dina(w_n631_6[1]),.dinb(w_G311_1[1]),.dout(n722),.clk(gclk));
	jand g0650(.dina(w_n617_5[1]),.dinb(w_G107_3[0]),.dout(n723),.clk(gclk));
	jand g0651(.dina(w_n642_6[1]),.dinb(w_G283_3[0]),.dout(n724),.clk(gclk));
	jor g0652(.dina(w_dff_B_OhJl4kWT7_0),.dinb(n723),.dout(n725),.clk(gclk));
	jor g0653(.dina(n725),.dinb(w_dff_B_F3OXA4Xb4_1),.dout(n726),.clk(gclk));
	jnot g0654(.din(n726),.dout(n727),.clk(gclk));
	jand g0655(.dina(w_n634_3[1]),.dinb(w_G87_2[0]),.dout(n728),.clk(gclk));
	jnot g0656(.din(w_n728_0[1]),.dout(n729),.clk(gclk));
	jand g0657(.dina(n729),.dinb(w_G33_5[2]),.dout(n730),.clk(gclk));
	jand g0658(.dina(w_n636_6[1]),.dinb(w_G116_3[2]),.dout(n731),.clk(gclk));
	jand g0659(.dina(w_n627_6[1]),.dinb(w_G294_2[2]),.dout(n732),.clk(gclk));
	jor g0660(.dina(n732),.dinb(n731),.dout(n733),.clk(gclk));
	jand g0661(.dina(w_n640_6[1]),.dinb(w_G303_2[0]),.dout(n734),.clk(gclk));
	jor g0662(.dina(w_dff_B_NRsKYzsN1_0),.dinb(w_n661_0[0]),.dout(n735),.clk(gclk));
	jor g0663(.dina(n735),.dinb(w_dff_B_cWpeFl2z9_1),.dout(n736),.clk(gclk));
	jnot g0664(.din(n736),.dout(n737),.clk(gclk));
	jand g0665(.dina(n737),.dinb(w_dff_B_lcR5Qci74_1),.dout(n738),.clk(gclk));
	jand g0666(.dina(n738),.dinb(w_dff_B_yxqJN0WG9_1),.dout(n739),.clk(gclk));
	jnot g0667(.din(n739),.dout(n740),.clk(gclk));
	jand g0668(.dina(n740),.dinb(w_dff_B_C5aySXOr5_1),.dout(n741),.clk(gclk));
	jor g0669(.dina(n741),.dinb(w_n612_3[2]),.dout(n742),.clk(gclk));
	jand g0670(.dina(w_n612_3[1]),.dinb(w_n426_0[0]),.dout(n743),.clk(gclk));
	jand g0671(.dina(w_n743_1[1]),.dinb(w_n72_0[1]),.dout(n744),.clk(gclk));
	jor g0672(.dina(w_dff_B_zCZBW35C3_0),.dinb(w_n605_1[1]),.dout(n745),.clk(gclk));
	jnot g0673(.din(n745),.dout(n746),.clk(gclk));
	jand g0674(.dina(w_dff_B_RMjq1yaJ2_0),.dinb(n742),.dout(n747),.clk(gclk));
	jand g0675(.dina(w_dff_B_zcaO3fTP5_0),.dinb(n705),.dout(n748),.clk(gclk));
	jnot g0676(.din(n748),.dout(n749),.clk(gclk));
	jand g0677(.dina(n749),.dinb(n702),.dout(n750),.clk(gclk));
	jnot g0678(.din(w_n750_0[1]),.dout(G384_fa_),.clk(gclk));
	jnot g0679(.din(w_n552_1[0]),.dout(n752),.clk(gclk));
	jand g0680(.dina(w_dff_B_A1m94hoT3_0),.dinb(w_n542_0[1]),.dout(n753),.clk(gclk));
	jand g0681(.dina(w_n552_0[2]),.dinb(w_n512_0[0]),.dout(n754),.clk(gclk));
	jnot g0682(.din(w_n754_0[1]),.dout(n755),.clk(gclk));
	jand g0683(.dina(n755),.dinb(w_n517_0[0]),.dout(n756),.clk(gclk));
	jand g0684(.dina(w_n754_0[0]),.dinb(w_n542_0[0]),.dout(n757),.clk(gclk));
	jor g0685(.dina(n757),.dinb(n756),.dout(n758),.clk(gclk));
	jand g0686(.dina(w_n696_1[0]),.dinb(w_n576_0[2]),.dout(n759),.clk(gclk));
	jand g0687(.dina(w_n553_1[2]),.dinb(w_n436_0[0]),.dout(n760),.clk(gclk));
	jnot g0688(.din(w_n760_0[1]),.dout(n761),.clk(gclk));
	jand g0689(.dina(w_dff_B_2SXwo92r8_0),.dinb(w_n446_0[0]),.dout(n762),.clk(gclk));
	jand g0690(.dina(w_n760_0[0]),.dinb(w_n439_0[2]),.dout(n763),.clk(gclk));
	jor g0691(.dina(w_dff_B_HDbb506a3_0),.dinb(n762),.dout(n764),.clk(gclk));
	jand g0692(.dina(w_n764_1[2]),.dinb(w_n759_0[1]),.dout(n765),.clk(gclk));
	jor g0693(.dina(w_n764_1[1]),.dinb(w_n439_0[1]),.dout(n766),.clk(gclk));
	jand g0694(.dina(w_n554_1[2]),.dinb(w_n543_0[0]),.dout(n767),.clk(gclk));
	jand g0695(.dina(w_dff_B_hlRPCz2F6_0),.dinb(n766),.dout(n768),.clk(gclk));
	jor g0696(.dina(w_dff_B_6DSs9HIL1_0),.dinb(n765),.dout(n769),.clk(gclk));
	jand g0697(.dina(w_n769_0[1]),.dinb(w_n758_1[1]),.dout(n770),.clk(gclk));
	jor g0698(.dina(n770),.dinb(w_dff_B_JsDsytI55_1),.dout(n771),.clk(gclk));
	jnot g0699(.din(w_n771_0[2]),.dout(n772),.clk(gclk));
	jand g0700(.dina(w_n576_0[1]),.dinb(w_n519_1[0]),.dout(n773),.clk(gclk));
	jor g0701(.dina(n773),.dinb(w_n548_0[1]),.dout(n774),.clk(gclk));
	jand g0702(.dina(w_n764_1[0]),.dinb(w_n696_0[2]),.dout(n775),.clk(gclk));
	jand g0703(.dina(n775),.dinb(w_n758_1[0]),.dout(n776),.clk(gclk));
	jxor g0704(.dina(n776),.dinb(w_n519_0[2]),.dout(n777),.clk(gclk));
	jand g0705(.dina(n777),.dinb(w_n588_0[2]),.dout(n778),.clk(gclk));
	jxor g0706(.dina(n778),.dinb(w_dff_B_C6myuNG13_1),.dout(n779),.clk(gclk));
	jnot g0707(.din(w_n779_0[1]),.dout(n780),.clk(gclk));
	jor g0708(.dina(w_dff_B_1ebv9Ywc6_0),.dinb(n772),.dout(n781),.clk(gclk));
	jor g0709(.dina(w_n779_0[0]),.dinb(w_n771_0[1]),.dout(n782),.clk(gclk));
	jnot g0710(.din(w_n121_0[1]),.dout(n783),.clk(gclk));
	jand g0711(.dina(n783),.dinb(w_n116_0[0]),.dout(n784),.clk(gclk));
	jand g0712(.dina(w_dff_B_08UZhAAQ1_0),.dinb(n782),.dout(n785),.clk(gclk));
	jand g0713(.dina(n785),.dinb(n781),.dout(n786),.clk(gclk));
	jand g0714(.dina(w_G77_3[0]),.dinb(w_G50_3[1]),.dout(n787),.clk(gclk));
	jand g0715(.dina(n787),.dinb(w_n137_0[0]),.dout(n788),.clk(gclk));
	jand g0716(.dina(w_G68_3[0]),.dinb(w_n73_1[2]),.dout(n789),.clk(gclk));
	jor g0717(.dina(n789),.dinb(n788),.dout(n790),.clk(gclk));
	jand g0718(.dina(n790),.dinb(w_n121_0[0]),.dout(n791),.clk(gclk));
	jnot g0719(.din(w_n255_0[0]),.dout(n792),.clk(gclk));
	jand g0720(.dina(w_n147_0[0]),.dinb(w_G116_3[1]),.dout(n793),.clk(gclk));
	jand g0721(.dina(w_dff_B_8dhPwf6t8_0),.dinb(n792),.dout(n794),.clk(gclk));
	jor g0722(.dina(n794),.dinb(w_dff_B_h20AqAp38_1),.dout(n795),.clk(gclk));
	jor g0723(.dina(w_dff_B_a03BJKRD2_0),.dinb(n786),.dout(w_dff_A_WtxJkxnW0_2),.clk(gclk));
	jand g0724(.dina(w_n553_1[1]),.dinb(w_n214_0[0]),.dout(n797),.clk(gclk));
	jnot g0725(.din(w_n797_0[1]),.dout(n798),.clk(gclk));
	jand g0726(.dina(w_dff_B_t8wk4rsF8_0),.dinb(w_n219_0[0]),.dout(n799),.clk(gclk));
	jand g0727(.dina(w_n797_0[0]),.dinb(w_n532_0[0]),.dout(n800),.clk(gclk));
	jor g0728(.dina(w_dff_B_GTkGHyzu7_0),.dinb(n799),.dout(n801),.clk(gclk));
	jnot g0729(.din(w_n801_0[1]),.dout(n802),.clk(gclk));
	jand g0730(.dina(n802),.dinb(w_n608_1[0]),.dout(n803),.clk(gclk));
	jnot g0731(.din(n803),.dout(n804),.clk(gclk));
	jand g0732(.dina(w_n631_6[0]),.dinb(w_G317_1[0]),.dout(n805),.clk(gclk));
	jand g0733(.dina(w_n623_4[1]),.dinb(w_G107_2[2]),.dout(n806),.clk(gclk));
	jand g0734(.dina(w_n642_6[0]),.dinb(w_G294_2[1]),.dout(n807),.clk(gclk));
	jor g0735(.dina(w_dff_B_AFA9y1HW5_0),.dinb(n806),.dout(n808),.clk(gclk));
	jor g0736(.dina(n808),.dinb(w_dff_B_GKEavJx33_1),.dout(n809),.clk(gclk));
	jand g0737(.dina(w_n617_5[0]),.dinb(w_G116_3[0]),.dout(n810),.clk(gclk));
	jor g0738(.dina(n810),.dinb(w_n148_4[2]),.dout(n811),.clk(gclk));
	jand g0739(.dina(w_n636_6[0]),.dinb(w_G283_2[2]),.dout(n812),.clk(gclk));
	jand g0740(.dina(w_n627_6[0]),.dinb(w_G303_1[2]),.dout(n813),.clk(gclk));
	jor g0741(.dina(n813),.dinb(n812),.dout(n814),.clk(gclk));
	jand g0742(.dina(w_n640_6[0]),.dinb(w_G311_1[0]),.dout(n815),.clk(gclk));
	jand g0743(.dina(w_n634_3[0]),.dinb(w_G97_3[0]),.dout(n816),.clk(gclk));
	jor g0744(.dina(w_n816_0[1]),.dinb(w_dff_B_oPSouTSc8_1),.dout(n817),.clk(gclk));
	jor g0745(.dina(n817),.dinb(w_dff_B_KHWzBYxD2_1),.dout(n818),.clk(gclk));
	jor g0746(.dina(n818),.dinb(w_dff_B_AHrNX2v01_1),.dout(n819),.clk(gclk));
	jor g0747(.dina(n819),.dinb(w_dff_B_yM0ra25v9_1),.dout(n820),.clk(gclk));
	jand g0748(.dina(w_n631_5[2]),.dinb(w_G137_1[1]),.dout(n821),.clk(gclk));
	jnot g0749(.din(n821),.dout(n822),.clk(gclk));
	jand g0750(.dina(w_n623_4[0]),.dinb(w_G68_2[2]),.dout(n823),.clk(gclk));
	jnot g0751(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jand g0752(.dina(w_n634_2[2]),.dinb(w_G77_2[2]),.dout(n825),.clk(gclk));
	jnot g0753(.din(w_n825_0[1]),.dout(n826),.clk(gclk));
	jand g0754(.dina(n826),.dinb(n824),.dout(n827),.clk(gclk));
	jand g0755(.dina(n827),.dinb(w_dff_B_Ndnd0jB51_1),.dout(n828),.clk(gclk));
	jand g0756(.dina(w_n642_5[2]),.dinb(w_G159_2[2]),.dout(n829),.clk(gclk));
	jor g0757(.dina(n829),.dinb(w_G33_5[1]),.dout(n830),.clk(gclk));
	jand g0758(.dina(w_n640_5[2]),.dinb(w_G143_2[0]),.dout(n831),.clk(gclk));
	jand g0759(.dina(w_n627_5[2]),.dinb(w_G150_2[2]),.dout(n832),.clk(gclk));
	jor g0760(.dina(n832),.dinb(n831),.dout(n833),.clk(gclk));
	jand g0761(.dina(w_n636_5[2]),.dinb(w_G50_3[0]),.dout(n834),.clk(gclk));
	jand g0762(.dina(w_n617_4[2]),.dinb(w_G58_3[0]),.dout(n835),.clk(gclk));
	jor g0763(.dina(n835),.dinb(w_dff_B_PnW7Xyv40_1),.dout(n836),.clk(gclk));
	jor g0764(.dina(n836),.dinb(w_dff_B_gaXse5MV6_1),.dout(n837),.clk(gclk));
	jor g0765(.dina(n837),.dinb(w_dff_B_1vTMB9525_1),.dout(n838),.clk(gclk));
	jnot g0766(.din(n838),.dout(n839),.clk(gclk));
	jand g0767(.dina(n839),.dinb(w_dff_B_L0ZsuJQK0_1),.dout(n840),.clk(gclk));
	jnot g0768(.din(n840),.dout(n841),.clk(gclk));
	jand g0769(.dina(n841),.dinb(w_dff_B_fgFE3RpO0_1),.dout(n842),.clk(gclk));
	jor g0770(.dina(n842),.dinb(w_n612_3[0]),.dout(n843),.clk(gclk));
	jand g0771(.dina(w_n675_0[1]),.dinb(w_n131_0[0]),.dout(n844),.clk(gclk));
	jand g0772(.dina(w_n123_1[0]),.dinb(w_G87_1[2]),.dout(n845),.clk(gclk));
	jor g0773(.dina(w_dff_B_kFkvmHd54_0),.dinb(w_n672_1[0]),.dout(n846),.clk(gclk));
	jor g0774(.dina(n846),.dinb(w_dff_B_xoQRnqys4_1),.dout(n847),.clk(gclk));
	jand g0775(.dina(n847),.dinb(w_n604_1[1]),.dout(n848),.clk(gclk));
	jand g0776(.dina(w_dff_B_qBCX1vVK1_0),.dinb(n843),.dout(n849),.clk(gclk));
	jand g0777(.dina(w_dff_B_Aj2D0Oer9_0),.dinb(n804),.dout(n850),.clk(gclk));
	jnot g0778(.din(w_n589_1[1]),.dout(n851),.clk(gclk));
	jxor g0779(.dina(w_n561_0[0]),.dinb(w_n556_0[0]),.dout(n852),.clk(gclk));
	jxor g0780(.dina(w_dff_B_nXU4JbEZ0_0),.dinb(w_n572_0[0]),.dout(n853),.clk(gclk));
	jnot g0781(.din(w_n853_0[2]),.dout(n854),.clk(gclk));
	jand g0782(.dina(n854),.dinb(n851),.dout(n855),.clk(gclk));
	jnot g0783(.din(w_n278_0[0]),.dout(n856),.clk(gclk));
	jand g0784(.dina(w_n553_1[0]),.dinb(w_n274_0[0]),.dout(n857),.clk(gclk));
	jor g0785(.dina(w_dff_B_oPHEf5Ne0_0),.dinb(n856),.dout(n858),.clk(gclk));
	jand g0786(.dina(w_n553_0[2]),.dinb(w_n536_0[1]),.dout(n859),.clk(gclk));
	jnot g0787(.din(n859),.dout(n860),.clk(gclk));
	jand g0788(.dina(w_dff_B_2BHfzlba9_0),.dinb(n858),.dout(n861),.clk(gclk));
	jxor g0789(.dina(w_n861_1[1]),.dinb(w_n573_0[1]),.dout(n862),.clk(gclk));
	jxor g0790(.dina(n862),.dinb(w_n563_0[1]),.dout(n863),.clk(gclk));
	jand g0791(.dina(w_n863_0[1]),.dinb(w_n855_0[2]),.dout(n864),.clk(gclk));
	jor g0792(.dina(w_n864_0[1]),.dinb(w_n589_1[0]),.dout(n865),.clk(gclk));
	jand g0793(.dina(n865),.dinb(w_n591_0[2]),.dout(n866),.clk(gclk));
	jor g0794(.dina(n866),.dinb(w_n602_0[0]),.dout(n867),.clk(gclk));
	jand g0795(.dina(w_n554_1[1]),.dinb(w_n536_0[0]),.dout(n868),.clk(gclk));
	jnot g0796(.din(w_n861_1[0]),.dout(n869),.clk(gclk));
	jand g0797(.dina(n869),.dinb(w_n563_0[0]),.dout(n870),.clk(gclk));
	jor g0798(.dina(n870),.dinb(w_dff_B_cj0UxHTU6_1),.dout(n871),.clk(gclk));
	jor g0799(.dina(w_n861_0[2]),.dinb(w_n573_0[0]),.dout(n872),.clk(gclk));
	jxor g0800(.dina(n872),.dinb(w_n801_0[0]),.dout(n873),.clk(gclk));
	jxor g0801(.dina(n873),.dinb(w_dff_B_XYbubFso9_1),.dout(n874),.clk(gclk));
	jnot g0802(.din(n874),.dout(n875),.clk(gclk));
	jand g0803(.dina(w_dff_B_i61UwHm20_0),.dinb(n867),.dout(n876),.clk(gclk));
	jor g0804(.dina(n876),.dinb(w_dff_B_enNp6FUD9_1),.dout(G387_fa_),.clk(gclk));
	jand g0805(.dina(w_n853_0[1]),.dinb(w_n589_0[2]),.dout(n878),.clk(gclk));
	jor g0806(.dina(w_n855_0[1]),.dinb(w_n592_1[2]),.dout(n879),.clk(gclk));
	jor g0807(.dina(n879),.dinb(w_dff_B_J8ntFLjC9_1),.dout(n880),.clk(gclk));
	jor g0808(.dina(w_n853_0[0]),.dinb(w_n603_2[0]),.dout(n881),.clk(gclk));
	jand g0809(.dina(w_n608_0[2]),.dinb(w_n564_0[0]),.dout(n882),.clk(gclk));
	jand g0810(.dina(w_n631_5[1]),.dinb(w_G326_0[0]),.dout(n883),.clk(gclk));
	jand g0811(.dina(w_n623_3[2]),.dinb(w_G283_2[1]),.dout(n884),.clk(gclk));
	jand g0812(.dina(w_n627_5[1]),.dinb(w_G317_0[2]),.dout(n885),.clk(gclk));
	jor g0813(.dina(w_dff_B_xN7FYkZb6_0),.dinb(n884),.dout(n886),.clk(gclk));
	jor g0814(.dina(n886),.dinb(w_dff_B_dxEGLWIz7_1),.dout(n887),.clk(gclk));
	jand g0815(.dina(w_n617_4[1]),.dinb(w_G294_2[0]),.dout(n888),.clk(gclk));
	jor g0816(.dina(n888),.dinb(w_n148_4[1]),.dout(n889),.clk(gclk));
	jand g0817(.dina(w_n634_2[1]),.dinb(w_G116_2[2]),.dout(n890),.clk(gclk));
	jand g0818(.dina(w_n636_5[1]),.dinb(w_G303_1[1]),.dout(n891),.clk(gclk));
	jor g0819(.dina(w_dff_B_eC3jd1QQ4_0),.dinb(n890),.dout(n892),.clk(gclk));
	jand g0820(.dina(w_n640_5[1]),.dinb(w_G322_0[1]),.dout(n893),.clk(gclk));
	jand g0821(.dina(w_n642_5[1]),.dinb(w_G311_0[2]),.dout(n894),.clk(gclk));
	jor g0822(.dina(n894),.dinb(n893),.dout(n895),.clk(gclk));
	jor g0823(.dina(w_dff_B_rwqpw1ea0_0),.dinb(n892),.dout(n896),.clk(gclk));
	jor g0824(.dina(n896),.dinb(w_dff_B_1ecaiyHG9_1),.dout(n897),.clk(gclk));
	jor g0825(.dina(n897),.dinb(w_dff_B_7xFu4Mi80_1),.dout(n898),.clk(gclk));
	jand g0826(.dina(w_n623_3[1]),.dinb(w_G87_1[1]),.dout(n899),.clk(gclk));
	jand g0827(.dina(w_n642_5[0]),.dinb(w_G58_2[2]),.dout(n900),.clk(gclk));
	jor g0828(.dina(w_dff_B_qmhAqa5p4_0),.dinb(w_n816_0[0]),.dout(n901),.clk(gclk));
	jor g0829(.dina(n901),.dinb(w_n899_0[1]),.dout(n902),.clk(gclk));
	jand g0830(.dina(w_n631_5[0]),.dinb(w_G150_2[1]),.dout(n903),.clk(gclk));
	jor g0831(.dina(n903),.dinb(w_G33_5[0]),.dout(n904),.clk(gclk));
	jand g0832(.dina(w_n640_5[0]),.dinb(w_G159_2[1]),.dout(n905),.clk(gclk));
	jand g0833(.dina(w_n636_5[0]),.dinb(w_G68_2[1]),.dout(n906),.clk(gclk));
	jor g0834(.dina(n906),.dinb(n905),.dout(n907),.clk(gclk));
	jand g0835(.dina(w_n627_5[0]),.dinb(w_G50_2[2]),.dout(n908),.clk(gclk));
	jand g0836(.dina(w_n617_4[0]),.dinb(w_G77_2[1]),.dout(n909),.clk(gclk));
	jor g0837(.dina(w_n909_0[1]),.dinb(w_dff_B_w8ZFtNkY0_1),.dout(n910),.clk(gclk));
	jor g0838(.dina(n910),.dinb(w_dff_B_m1toFi2Z4_1),.dout(n911),.clk(gclk));
	jor g0839(.dina(n911),.dinb(w_dff_B_T0JGSakf5_1),.dout(n912),.clk(gclk));
	jor g0840(.dina(n912),.dinb(w_dff_B_snBJIKE72_1),.dout(n913),.clk(gclk));
	jand g0841(.dina(n913),.dinb(n898),.dout(n914),.clk(gclk));
	jor g0842(.dina(n914),.dinb(w_n612_2[2]),.dout(n915),.clk(gclk));
	jand g0843(.dina(w_n135_0[0]),.dinb(w_G45_0[1]),.dout(n916),.clk(gclk));
	jand g0844(.dina(w_G77_2[0]),.dinb(w_G68_2[0]),.dout(n917),.clk(gclk));
	jnot g0845(.din(n917),.dout(n918),.clk(gclk));
	jand g0846(.dina(w_G58_2[1]),.dinb(w_n161_0[1]),.dout(n919),.clk(gclk));
	jand g0847(.dina(n919),.dinb(w_n73_1[1]),.dout(n920),.clk(gclk));
	jand g0848(.dina(n920),.dinb(w_dff_B_9szqQOzh1_1),.dout(n921),.clk(gclk));
	jand g0849(.dina(n921),.dinb(w_n593_0[1]),.dout(n922),.clk(gclk));
	jor g0850(.dina(n922),.dinb(w_n676_0[0]),.dout(n923),.clk(gclk));
	jor g0851(.dina(n923),.dinb(w_dff_B_c9gsHbY27_1),.dout(n924),.clk(gclk));
	jand g0852(.dina(w_n123_0[2]),.dinb(w_n80_0[1]),.dout(n925),.clk(gclk));
	jnot g0853(.din(w_n593_0[0]),.dout(n926),.clk(gclk));
	jand g0854(.dina(w_n680_0[0]),.dinb(n926),.dout(n927),.clk(gclk));
	jor g0855(.dina(n927),.dinb(w_dff_B_MUofsgPe6_1),.dout(n928),.clk(gclk));
	jnot g0856(.din(n928),.dout(n929),.clk(gclk));
	jand g0857(.dina(n929),.dinb(w_dff_B_GmrysAj40_1),.dout(n930),.clk(gclk));
	jor g0858(.dina(n930),.dinb(w_n672_0[2]),.dout(n931),.clk(gclk));
	jand g0859(.dina(n931),.dinb(w_n604_1[0]),.dout(n932),.clk(gclk));
	jand g0860(.dina(n932),.dinb(n915),.dout(n933),.clk(gclk));
	jnot g0861(.din(n933),.dout(n934),.clk(gclk));
	jor g0862(.dina(w_dff_B_GFBcvfg54_0),.dinb(n882),.dout(n935),.clk(gclk));
	jand g0863(.dina(w_dff_B_Lcvoh0Hp3_0),.dinb(n881),.dout(n936),.clk(gclk));
	jand g0864(.dina(w_dff_B_U9NVKsvB8_0),.dinb(n880),.dout(n937),.clk(gclk));
	jnot g0865(.din(w_n937_0[2]),.dout(w_dff_A_HbcdcMhN5_1),.clk(gclk));
	jnot g0866(.din(w_n855_0[0]),.dout(n939),.clk(gclk));
	jnot g0867(.din(w_n863_0[0]),.dout(n940),.clk(gclk));
	jand g0868(.dina(w_n940_0[1]),.dinb(n939),.dout(n941),.clk(gclk));
	jor g0869(.dina(w_n864_0[0]),.dinb(w_n592_1[1]),.dout(n942),.clk(gclk));
	jor g0870(.dina(n942),.dinb(n941),.dout(n943),.clk(gclk));
	jor g0871(.dina(w_n940_0[0]),.dinb(w_n603_1[2]),.dout(n944),.clk(gclk));
	jand g0872(.dina(w_n861_0[1]),.dinb(w_n608_0[1]),.dout(n945),.clk(gclk));
	jnot g0873(.din(n945),.dout(n946),.clk(gclk));
	jand g0874(.dina(w_n623_3[0]),.dinb(w_G116_2[1]),.dout(n947),.clk(gclk));
	jand g0875(.dina(w_n617_3[2]),.dinb(w_G283_2[0]),.dout(n948),.clk(gclk));
	jand g0876(.dina(w_n642_4[2]),.dinb(w_G303_1[0]),.dout(n949),.clk(gclk));
	jor g0877(.dina(w_dff_B_5wy3jEUG6_0),.dinb(n948),.dout(n950),.clk(gclk));
	jor g0878(.dina(n950),.dinb(w_dff_B_3BYFU6wk9_1),.dout(n951),.clk(gclk));
	jand g0879(.dina(w_n631_4[2]),.dinb(w_G322_0[0]),.dout(n952),.clk(gclk));
	jor g0880(.dina(n952),.dinb(w_n148_4[0]),.dout(n953),.clk(gclk));
	jand g0881(.dina(w_n636_4[2]),.dinb(w_G294_1[2]),.dout(n954),.clk(gclk));
	jand g0882(.dina(w_n627_4[2]),.dinb(w_G311_0[1]),.dout(n955),.clk(gclk));
	jor g0883(.dina(n955),.dinb(n954),.dout(n956),.clk(gclk));
	jand g0884(.dina(w_n640_4[2]),.dinb(w_G317_0[1]),.dout(n957),.clk(gclk));
	jor g0885(.dina(w_dff_B_LXJkArUv7_0),.dinb(w_n657_0[0]),.dout(n958),.clk(gclk));
	jor g0886(.dina(n958),.dinb(w_dff_B_Sa8S6l657_1),.dout(n959),.clk(gclk));
	jor g0887(.dina(n959),.dinb(w_dff_B_0qytQobt8_1),.dout(n960),.clk(gclk));
	jor g0888(.dina(n960),.dinb(w_dff_B_DvXIxyGf4_1),.dout(n961),.clk(gclk));
	jand g0889(.dina(w_n623_2[2]),.dinb(w_G77_1[2]),.dout(n962),.clk(gclk));
	jand g0890(.dina(w_n617_3[1]),.dinb(w_G68_1[2]),.dout(n963),.clk(gclk));
	jand g0891(.dina(w_n642_4[1]),.dinb(w_G50_2[1]),.dout(n964),.clk(gclk));
	jor g0892(.dina(w_dff_B_p93FT1pd2_0),.dinb(n963),.dout(n965),.clk(gclk));
	jor g0893(.dina(n965),.dinb(w_n962_0[1]),.dout(n966),.clk(gclk));
	jand g0894(.dina(w_n631_4[1]),.dinb(w_G143_1[2]),.dout(n967),.clk(gclk));
	jor g0895(.dina(n967),.dinb(w_G33_4[2]),.dout(n968),.clk(gclk));
	jand g0896(.dina(w_n636_4[1]),.dinb(w_G58_2[0]),.dout(n969),.clk(gclk));
	jand g0897(.dina(w_n627_4[1]),.dinb(w_G159_2[0]),.dout(n970),.clk(gclk));
	jor g0898(.dina(n970),.dinb(n969),.dout(n971),.clk(gclk));
	jand g0899(.dina(w_n640_4[1]),.dinb(w_G150_2[0]),.dout(n972),.clk(gclk));
	jor g0900(.dina(w_dff_B_GlulZvDF5_0),.dinb(w_n728_0[0]),.dout(n973),.clk(gclk));
	jor g0901(.dina(n973),.dinb(w_dff_B_X01pjMDj1_1),.dout(n974),.clk(gclk));
	jor g0902(.dina(n974),.dinb(w_dff_B_gXHOsSIl6_1),.dout(n975),.clk(gclk));
	jor g0903(.dina(n975),.dinb(w_dff_B_Ir9qfCf96_1),.dout(n976),.clk(gclk));
	jand g0904(.dina(n976),.dinb(n961),.dout(n977),.clk(gclk));
	jor g0905(.dina(n977),.dinb(w_n612_2[1]),.dout(n978),.clk(gclk));
	jand g0906(.dina(w_n675_0[0]),.dinb(w_n144_0[0]),.dout(n979),.clk(gclk));
	jand g0907(.dina(w_n123_0[1]),.dinb(w_G97_2[2]),.dout(n980),.clk(gclk));
	jor g0908(.dina(w_dff_B_s7OrRFQo7_0),.dinb(w_n672_0[1]),.dout(n981),.clk(gclk));
	jor g0909(.dina(n981),.dinb(w_dff_B_K02sLONx8_1),.dout(n982),.clk(gclk));
	jand g0910(.dina(n982),.dinb(w_n604_0[2]),.dout(n983),.clk(gclk));
	jand g0911(.dina(w_dff_B_Qr37CMcf9_0),.dinb(n978),.dout(n984),.clk(gclk));
	jand g0912(.dina(w_dff_B_iMrcfwYr1_0),.dinb(n946),.dout(n985),.clk(gclk));
	jnot g0913(.din(n985),.dout(n986),.clk(gclk));
	jand g0914(.dina(w_dff_B_oI9jQJTi4_0),.dinb(n944),.dout(n987),.clk(gclk));
	jand g0915(.dina(n987),.dinb(n943),.dout(n988),.clk(gclk));
	jnot g0916(.din(w_n988_0[2]),.dout(w_dff_A_Xq1tvspa5_1),.clk(gclk));
	jnot g0917(.din(w_n758_0[2]),.dout(n990),.clk(gclk));
	jand g0918(.dina(w_n696_0[1]),.dinb(w_n588_0[1]),.dout(n991),.clk(gclk));
	jand g0919(.dina(w_n991_0[1]),.dinb(w_n764_0[2]),.dout(n992),.clk(gclk));
	jxor g0920(.dina(w_n992_0[1]),.dinb(w_n990_0[1]),.dout(n993),.clk(gclk));
	jxor g0921(.dina(n993),.dinb(w_n769_0[0]),.dout(n994),.clk(gclk));
	jand g0922(.dina(w_n589_0[1]),.dinb(w_n519_0[1]),.dout(n995),.clk(gclk));
	jor g0923(.dina(n995),.dinb(w_n548_0[0]),.dout(n996),.clk(gclk));
	jand g0924(.dina(w_n554_1[0]),.dinb(w_n404_0[0]),.dout(n997),.clk(gclk));
	jor g0925(.dina(w_dff_B_LnzMSa2X5_0),.dinb(w_n759_0[0]),.dout(n998),.clk(gclk));
	jnot g0926(.din(w_n764_0[1]),.dout(n999),.clk(gclk));
	jxor g0927(.dina(w_n991_0[0]),.dinb(w_n999_0[1]),.dout(n1000),.clk(gclk));
	jxor g0928(.dina(n1000),.dinb(n998),.dout(n1001),.clk(gclk));
	jor g0929(.dina(w_n1001_0[2]),.dinb(w_n996_0[2]),.dout(n1002),.clk(gclk));
	jor g0930(.dina(w_n1002_0[2]),.dinb(w_n994_0[2]),.dout(n1003),.clk(gclk));
	jnot g0931(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jand g0932(.dina(w_n1002_0[1]),.dinb(w_n994_0[1]),.dout(n1005),.clk(gclk));
	jor g0933(.dina(n1005),.dinb(w_n592_1[0]),.dout(n1006),.clk(gclk));
	jor g0934(.dina(n1006),.dinb(n1004),.dout(n1007),.clk(gclk));
	jor g0935(.dina(w_n994_0[0]),.dinb(w_n603_1[1]),.dout(n1008),.clk(gclk));
	jand g0936(.dina(w_n990_0[0]),.dinb(w_n425_1[0]),.dout(n1009),.clk(gclk));
	jnot g0937(.din(n1009),.dout(n1010),.clk(gclk));
	jand g0938(.dina(w_n631_4[0]),.dinb(w_G125_0[1]),.dout(n1011),.clk(gclk));
	jand g0939(.dina(w_n623_2[1]),.dinb(w_G159_1[2]),.dout(n1012),.clk(gclk));
	jand g0940(.dina(w_n642_4[0]),.dinb(w_G137_1[0]),.dout(n1013),.clk(gclk));
	jor g0941(.dina(w_dff_B_deyEznqR1_0),.dinb(n1012),.dout(n1014),.clk(gclk));
	jor g0942(.dina(n1014),.dinb(w_dff_B_t1VZo9LU6_1),.dout(n1015),.clk(gclk));
	jand g0943(.dina(w_n617_3[0]),.dinb(w_G150_1[2]),.dout(n1016),.clk(gclk));
	jor g0944(.dina(n1016),.dinb(w_G33_4[1]),.dout(n1017),.clk(gclk));
	jand g0945(.dina(w_n636_4[0]),.dinb(w_G143_1[1]),.dout(n1018),.clk(gclk));
	jand g0946(.dina(w_n627_4[0]),.dinb(w_G132_1[0]),.dout(n1019),.clk(gclk));
	jor g0947(.dina(n1019),.dinb(n1018),.dout(n1020),.clk(gclk));
	jand g0948(.dina(w_n640_4[0]),.dinb(w_G128_0[2]),.dout(n1021),.clk(gclk));
	jand g0949(.dina(w_n634_2[0]),.dinb(w_G50_2[0]),.dout(n1022),.clk(gclk));
	jor g0950(.dina(n1022),.dinb(w_dff_B_AGdyaDFT8_1),.dout(n1023),.clk(gclk));
	jor g0951(.dina(n1023),.dinb(w_dff_B_cJrdyOfY6_1),.dout(n1024),.clk(gclk));
	jor g0952(.dina(n1024),.dinb(w_dff_B_W72VKEnG4_1),.dout(n1025),.clk(gclk));
	jor g0953(.dina(n1025),.dinb(w_dff_B_p51TAtIC9_1),.dout(n1026),.clk(gclk));
	jand g0954(.dina(w_n631_3[2]),.dinb(w_G294_1[1]),.dout(n1027),.clk(gclk));
	jand g0955(.dina(w_n642_3[2]),.dinb(w_G107_2[1]),.dout(n1028),.clk(gclk));
	jor g0956(.dina(w_dff_B_ksxvGuGo3_0),.dinb(w_n962_0[0]),.dout(n1029),.clk(gclk));
	jor g0957(.dina(n1029),.dinb(w_dff_B_sHvM5Zr10_1),.dout(n1030),.clk(gclk));
	jand g0958(.dina(w_n640_3[2]),.dinb(w_G283_1[2]),.dout(n1031),.clk(gclk));
	jor g0959(.dina(n1031),.dinb(w_n148_3[2]),.dout(n1032),.clk(gclk));
	jand g0960(.dina(w_n636_3[2]),.dinb(w_G97_2[1]),.dout(n1033),.clk(gclk));
	jand g0961(.dina(w_n627_3[2]),.dinb(w_G116_2[0]),.dout(n1034),.clk(gclk));
	jor g0962(.dina(n1034),.dinb(n1033),.dout(n1035),.clk(gclk));
	jor g0963(.dina(w_n717_0[0]),.dinb(w_n654_0[0]),.dout(n1036),.clk(gclk));
	jor g0964(.dina(n1036),.dinb(w_dff_B_v6lCpZNv0_1),.dout(n1037),.clk(gclk));
	jor g0965(.dina(n1037),.dinb(w_dff_B_KHdMP5A09_1),.dout(n1038),.clk(gclk));
	jor g0966(.dina(n1038),.dinb(w_dff_B_k4bCUjyl2_1),.dout(n1039),.clk(gclk));
	jand g0967(.dina(n1039),.dinb(n1026),.dout(n1040),.clk(gclk));
	jor g0968(.dina(n1040),.dinb(w_n612_2[0]),.dout(n1041),.clk(gclk));
	jand g0969(.dina(w_n743_1[0]),.dinb(w_n74_0[1]),.dout(n1042),.clk(gclk));
	jor g0970(.dina(w_dff_B_tM3qn2Od9_0),.dinb(w_n605_1[0]),.dout(n1043),.clk(gclk));
	jnot g0971(.din(n1043),.dout(n1044),.clk(gclk));
	jand g0972(.dina(w_dff_B_y7op2Qz88_0),.dinb(n1041),.dout(n1045),.clk(gclk));
	jand g0973(.dina(w_dff_B_fHRJB02K1_0),.dinb(n1010),.dout(n1046),.clk(gclk));
	jnot g0974(.din(n1046),.dout(n1047),.clk(gclk));
	jand g0975(.dina(w_dff_B_yo14BoqS2_0),.dinb(n1008),.dout(n1048),.clk(gclk));
	jand g0976(.dina(w_dff_B_zF4bDGEv2_0),.dinb(n1007),.dout(n1049),.clk(gclk));
	jnot g0977(.din(w_n1049_0[2]),.dout(w_dff_A_XeMRgOBq9_1),.clk(gclk));
	jand g0978(.dina(w_n992_0[0]),.dinb(w_n758_0[1]),.dout(n1051),.clk(gclk));
	jand g0979(.dina(w_n552_0[1]),.dinb(w_n479_0[0]),.dout(n1052),.clk(gclk));
	jnot g0980(.din(w_n1052_0[1]),.dout(n1053),.clk(gclk));
	jand g0981(.dina(n1053),.dinb(w_n484_0[0]),.dout(n1054),.clk(gclk));
	jand g0982(.dina(w_n1052_0[0]),.dinb(w_n541_0[0]),.dout(n1055),.clk(gclk));
	jor g0983(.dina(n1055),.dinb(n1054),.dout(n1056),.clk(gclk));
	jnot g0984(.din(n1056),.dout(n1057),.clk(gclk));
	jxor g0985(.dina(w_n1057_0[1]),.dinb(w_n771_0[0]),.dout(n1058),.clk(gclk));
	jxor g0986(.dina(n1058),.dinb(w_dff_B_0Wh4mUwg8_1),.dout(n1059),.clk(gclk));
	jor g0987(.dina(w_n1059_0[1]),.dinb(w_n603_1[0]),.dout(n1060),.clk(gclk));
	jnot g0988(.din(w_n996_0[1]),.dout(n1061),.clk(gclk));
	jand g0989(.dina(w_n1003_0[0]),.dinb(w_dff_B_ES2YB4tC6_1),.dout(n1062),.clk(gclk));
	jor g0990(.dina(n1062),.dinb(w_n592_0[2]),.dout(n1063),.clk(gclk));
	jor g0991(.dina(n1063),.dinb(w_n1059_0[0]),.dout(n1064),.clk(gclk));
	jand g0992(.dina(w_n1057_0[0]),.dinb(w_n425_0[2]),.dout(n1065),.clk(gclk));
	jnot g0993(.din(w_n612_1[2]),.dout(n1066),.clk(gclk));
	jand g0994(.dina(w_n642_3[1]),.dinb(w_G132_0[2]),.dout(n1067),.clk(gclk));
	jand g0995(.dina(w_n627_3[1]),.dinb(w_G128_0[1]),.dout(n1068),.clk(gclk));
	jand g0996(.dina(w_n636_3[1]),.dinb(w_G137_0[2]),.dout(n1069),.clk(gclk));
	jor g0997(.dina(n1069),.dinb(n1068),.dout(n1070),.clk(gclk));
	jor g0998(.dina(n1070),.dinb(w_dff_B_cgxjWMuI9_1),.dout(n1071),.clk(gclk));
	jnot g0999(.din(n1071),.dout(n1072),.clk(gclk));
	jand g1000(.dina(w_n623_2[0]),.dinb(w_G150_1[1]),.dout(n1073),.clk(gclk));
	jnot g1001(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1002(.dina(w_n149_1[0]),.dinb(w_n148_3[1]),.dout(n1075),.clk(gclk));
	jand g1003(.dina(w_dff_B_poS95E5R3_0),.dinb(n1074),.dout(n1076),.clk(gclk));
	jand g1004(.dina(w_n640_3[1]),.dinb(w_G125_0[0]),.dout(n1077),.clk(gclk));
	jand g1005(.dina(w_n617_2[2]),.dinb(w_G143_1[0]),.dout(n1078),.clk(gclk));
	jor g1006(.dina(n1078),.dinb(w_dff_B_BPeRjwXy5_1),.dout(n1079),.clk(gclk));
	jand g1007(.dina(w_n631_3[1]),.dinb(w_dff_B_erZgD98O7_1),.dout(n1080),.clk(gclk));
	jand g1008(.dina(w_n634_1[2]),.dinb(w_G159_1[1]),.dout(n1081),.clk(gclk));
	jor g1009(.dina(n1081),.dinb(n1080),.dout(n1082),.clk(gclk));
	jor g1010(.dina(n1082),.dinb(n1079),.dout(n1083),.clk(gclk));
	jnot g1011(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1012(.dina(n1084),.dinb(w_dff_B_SYxa1nNY0_1),.dout(n1085),.clk(gclk));
	jand g1013(.dina(n1085),.dinb(w_dff_B_UbgWf2mq6_1),.dout(n1086),.clk(gclk));
	jand g1014(.dina(w_n627_3[0]),.dinb(w_G107_2[0]),.dout(n1087),.clk(gclk));
	jand g1015(.dina(w_n634_1[1]),.dinb(w_G58_1[2]),.dout(n1088),.clk(gclk));
	jand g1016(.dina(w_n636_3[0]),.dinb(w_G87_1[0]),.dout(n1089),.clk(gclk));
	jor g1017(.dina(w_dff_B_DyzEanKZ7_0),.dinb(w_n1088_0[1]),.dout(n1090),.clk(gclk));
	jor g1018(.dina(n1090),.dinb(w_dff_B_Of5oisTA5_1),.dout(n1091),.clk(gclk));
	jnot g1019(.din(n1091),.dout(n1092),.clk(gclk));
	jand g1020(.dina(w_n642_3[0]),.dinb(w_G97_2[0]),.dout(n1093),.clk(gclk));
	jnot g1021(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1022(.dina(w_n149_0[2]),.dinb(w_G33_4[0]),.dout(n1095),.clk(gclk));
	jand g1023(.dina(w_dff_B_0VEg4nU59_0),.dinb(n1094),.dout(n1096),.clk(gclk));
	jand g1024(.dina(w_n631_3[0]),.dinb(w_G283_1[1]),.dout(n1097),.clk(gclk));
	jor g1025(.dina(n1097),.dinb(w_n823_0[0]),.dout(n1098),.clk(gclk));
	jand g1026(.dina(w_n640_3[0]),.dinb(w_G116_1[2]),.dout(n1099),.clk(gclk));
	jor g1027(.dina(w_dff_B_EHAmpLNC1_0),.dinb(w_n909_0[0]),.dout(n1100),.clk(gclk));
	jor g1028(.dina(n1100),.dinb(n1098),.dout(n1101),.clk(gclk));
	jnot g1029(.din(n1101),.dout(n1102),.clk(gclk));
	jand g1030(.dina(n1102),.dinb(w_dff_B_ZsBPbCzM7_1),.dout(n1103),.clk(gclk));
	jand g1031(.dina(n1103),.dinb(w_dff_B_yfineotg2_1),.dout(n1104),.clk(gclk));
	jand g1032(.dina(w_n73_1[0]),.dinb(w_G41_0[1]),.dout(n1105),.clk(gclk));
	jor g1033(.dina(w_dff_B_Ie3G75Ik7_0),.dinb(n1104),.dout(n1106),.clk(gclk));
	jor g1034(.dina(n1106),.dinb(w_dff_B_ms8W2Lke6_1),.dout(n1107),.clk(gclk));
	jand g1035(.dina(n1107),.dinb(w_dff_B_Dc1teHUy7_1),.dout(n1108),.clk(gclk));
	jand g1036(.dina(w_n743_0[2]),.dinb(w_n73_0[2]),.dout(n1109),.clk(gclk));
	jor g1037(.dina(w_dff_B_eWTdcCEz0_0),.dinb(w_n605_0[2]),.dout(n1110),.clk(gclk));
	jor g1038(.dina(w_dff_B_R0XxsxpC1_0),.dinb(n1108),.dout(n1111),.clk(gclk));
	jor g1039(.dina(w_dff_B_6RlGO1el5_0),.dinb(n1065),.dout(n1112),.clk(gclk));
	jand g1040(.dina(w_dff_B_M5crVnnZ1_0),.dinb(n1064),.dout(n1113),.clk(gclk));
	jand g1041(.dina(n1113),.dinb(w_dff_B_HbZ2tRBn8_1),.dout(n1114),.clk(gclk));
	jnot g1042(.din(w_n1114_0[2]),.dout(w_dff_A_suoffQtL3_1),.clk(gclk));
	jand g1043(.dina(w_n1001_0[1]),.dinb(w_n996_0[0]),.dout(n1116),.clk(gclk));
	jnot g1044(.din(n1116),.dout(n1117),.clk(gclk));
	jand g1045(.dina(w_n1002_0[0]),.dinb(w_n591_0[1]),.dout(n1118),.clk(gclk));
	jand g1046(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jnot g1047(.din(n1119),.dout(n1120),.clk(gclk));
	jor g1048(.dina(w_n1001_0[0]),.dinb(w_n603_0[2]),.dout(n1121),.clk(gclk));
	jand g1049(.dina(w_n999_0[0]),.dinb(w_n425_0[1]),.dout(n1122),.clk(gclk));
	jnot g1050(.din(n1122),.dout(n1123),.clk(gclk));
	jand g1051(.dina(w_n623_1[2]),.dinb(w_G50_1[2]),.dout(n1124),.clk(gclk));
	jand g1052(.dina(w_n617_2[1]),.dinb(w_G159_1[0]),.dout(n1125),.clk(gclk));
	jand g1053(.dina(w_n642_2[2]),.dinb(w_G143_0[2]),.dout(n1126),.clk(gclk));
	jor g1054(.dina(w_dff_B_7KXg4KOM0_0),.dinb(n1125),.dout(n1127),.clk(gclk));
	jor g1055(.dina(n1127),.dinb(w_dff_B_HEvNRcaN0_1),.dout(n1128),.clk(gclk));
	jand g1056(.dina(w_n631_2[2]),.dinb(w_G128_0[0]),.dout(n1129),.clk(gclk));
	jor g1057(.dina(n1129),.dinb(w_G33_3[2]),.dout(n1130),.clk(gclk));
	jand g1058(.dina(w_n636_2[2]),.dinb(w_G150_1[0]),.dout(n1131),.clk(gclk));
	jand g1059(.dina(w_n627_2[2]),.dinb(w_G137_0[1]),.dout(n1132),.clk(gclk));
	jor g1060(.dina(n1132),.dinb(n1131),.dout(n1133),.clk(gclk));
	jand g1061(.dina(w_n640_2[2]),.dinb(w_G132_0[1]),.dout(n1134),.clk(gclk));
	jor g1062(.dina(w_dff_B_Pd0enkjG3_0),.dinb(w_n1088_0[0]),.dout(n1135),.clk(gclk));
	jor g1063(.dina(n1135),.dinb(w_dff_B_3i5y8pxZ4_1),.dout(n1136),.clk(gclk));
	jor g1064(.dina(n1136),.dinb(w_dff_B_NeUMlFJp7_1),.dout(n1137),.clk(gclk));
	jor g1065(.dina(n1137),.dinb(w_dff_B_QIWtjCoA8_1),.dout(n1138),.clk(gclk));
	jand g1066(.dina(w_n617_2[0]),.dinb(w_G97_1[2]),.dout(n1139),.clk(gclk));
	jand g1067(.dina(w_n640_2[1]),.dinb(w_G294_1[0]),.dout(n1140),.clk(gclk));
	jand g1068(.dina(w_n642_2[1]),.dinb(w_G116_1[1]),.dout(n1141),.clk(gclk));
	jor g1069(.dina(n1141),.dinb(n1140),.dout(n1142),.clk(gclk));
	jor g1070(.dina(n1142),.dinb(n1139),.dout(n1143),.clk(gclk));
	jand g1071(.dina(w_n631_2[1]),.dinb(w_G303_0[2]),.dout(n1144),.clk(gclk));
	jor g1072(.dina(n1144),.dinb(w_n148_3[0]),.dout(n1145),.clk(gclk));
	jand g1073(.dina(w_n636_2[1]),.dinb(w_G107_1[2]),.dout(n1146),.clk(gclk));
	jand g1074(.dina(w_n627_2[1]),.dinb(w_G283_1[0]),.dout(n1147),.clk(gclk));
	jor g1075(.dina(n1147),.dinb(n1146),.dout(n1148),.clk(gclk));
	jor g1076(.dina(w_n899_0[0]),.dinb(w_n825_0[0]),.dout(n1149),.clk(gclk));
	jor g1077(.dina(n1149),.dinb(w_dff_B_yCLnCPdg4_1),.dout(n1150),.clk(gclk));
	jor g1078(.dina(n1150),.dinb(w_dff_B_OlxLIZKe6_1),.dout(n1151),.clk(gclk));
	jor g1079(.dina(n1151),.dinb(w_dff_B_nFwzypT18_1),.dout(n1152),.clk(gclk));
	jand g1080(.dina(n1152),.dinb(n1138),.dout(n1153),.clk(gclk));
	jor g1081(.dina(n1153),.dinb(w_n612_1[1]),.dout(n1154),.clk(gclk));
	jand g1082(.dina(w_n743_0[1]),.dinb(w_n75_0[1]),.dout(n1155),.clk(gclk));
	jor g1083(.dina(w_dff_B_ZCKLYel97_0),.dinb(w_n605_0[1]),.dout(n1156),.clk(gclk));
	jnot g1084(.din(n1156),.dout(n1157),.clk(gclk));
	jand g1085(.dina(w_dff_B_emuLrLSO1_0),.dinb(n1154),.dout(n1158),.clk(gclk));
	jand g1086(.dina(w_dff_B_OnyCKrrI0_0),.dinb(n1123),.dout(n1159),.clk(gclk));
	jnot g1087(.din(n1159),.dout(n1160),.clk(gclk));
	jand g1088(.dina(n1160),.dinb(n1121),.dout(n1161),.clk(gclk));
	jand g1089(.dina(w_dff_B_S5C3hmwv6_0),.dinb(n1120),.dout(n1162),.clk(gclk));
	jnot g1090(.din(w_n1162_0[2]),.dout(w_dff_A_BWmK6cNT5_1),.clk(gclk));
	jand g1091(.dina(w_n1114_0[1]),.dinb(w_n1049_0[1]),.dout(n1164),.clk(gclk));
	jnot g1092(.din(w_G387_0[1]),.dout(n1165),.clk(gclk));
	jnot g1093(.din(w_G396_0[1]),.dout(n1166),.clk(gclk));
	jand g1094(.dina(w_n937_0[1]),.dinb(w_dff_B_0z1zdyUY5_1),.dout(n1167),.clk(gclk));
	jand g1095(.dina(n1167),.dinb(w_n750_0[0]),.dout(n1168),.clk(gclk));
	jand g1096(.dina(n1168),.dinb(w_n988_0[1]),.dout(n1169),.clk(gclk));
	jand g1097(.dina(n1169),.dinb(w_n1162_0[1]),.dout(n1170),.clk(gclk));
	jand g1098(.dina(n1170),.dinb(n1165),.dout(n1171),.clk(gclk));
	jand g1099(.dina(n1171),.dinb(w_n1164_0[1]),.dout(n1172),.clk(gclk));
	jnot g1100(.din(w_n1172_0[1]),.dout(w_dff_A_cajdjt8l9_1),.clk(gclk));
	jnot g1101(.din(w_G213_0[1]),.dout(n1174),.clk(gclk));
	jnot g1102(.din(w_G343_0[0]),.dout(n1175),.clk(gclk));
	jand g1103(.dina(w_n1164_0[0]),.dinb(w_n1175_0[1]),.dout(n1176),.clk(gclk));
	jor g1104(.dina(n1176),.dinb(w_dff_B_70Lh1d4I4_1),.dout(n1177),.clk(gclk));
	jor g1105(.dina(n1177),.dinb(w_n1172_0[0]),.dout(G409),.clk(gclk));
	jxor g1106(.dina(w_n1162_0[0]),.dinb(w_G384_0),.dout(n1179),.clk(gclk));
	jxor g1107(.dina(w_n937_0[0]),.dinb(w_G396_0[0]),.dout(n1180),.clk(gclk));
	jxor g1108(.dina(w_n988_0[0]),.dinb(w_G387_0[0]),.dout(n1181),.clk(gclk));
	jxor g1109(.dina(n1181),.dinb(w_dff_B_oBSGK8As4_1),.dout(n1182),.clk(gclk));
	jxor g1110(.dina(n1182),.dinb(w_dff_B_ZOIj791h4_1),.dout(n1183),.clk(gclk));
	jand g1111(.dina(w_n1175_0[0]),.dinb(w_G213_0[0]),.dout(n1184),.clk(gclk));
	jnot g1112(.din(w_n1184_0[1]),.dout(n1185),.clk(gclk));
	jor g1113(.dina(n1185),.dinb(w_dff_B_QHOGV6Yf9_1),.dout(n1186),.clk(gclk));
	jxor g1114(.dina(w_n1114_0[0]),.dinb(w_n1049_0[0]),.dout(n1187),.clk(gclk));
	jor g1115(.dina(w_n1187_0[1]),.dinb(w_n1184_0[0]),.dout(n1188),.clk(gclk));
	jand g1116(.dina(n1188),.dinb(w_dff_B_kXptMM8s9_1),.dout(n1189),.clk(gclk));
	jxor g1117(.dina(n1189),.dinb(w_n1183_0[1]),.dout(G405),.clk(gclk));
	jxor g1118(.dina(w_n1187_0[0]),.dinb(w_n1183_0[0]),.dout(w_dff_A_AmqgxAwU4_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_dff_A_M6s2GyiG1_0),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_dff_A_8JtEjNTX7_0),.doutb(w_dff_A_6SIYP9g29_1),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G1_2(.douta(w_dff_A_IexZa1a62_0),.doutb(w_G1_2[1]),.doutc(w_dff_A_NB7BrxW80_2),.din(w_G1_0[1]));
	jspl jspl_w_G1_3(.douta(w_G1_3[0]),.doutb(w_G1_3[1]),.din(w_G1_0[2]));
	jspl3 jspl3_w_G13_0(.douta(w_G13_0[0]),.doutb(w_dff_A_ojIQhcSW4_1),.doutc(w_dff_A_zTZXqXCx5_2),.din(G13));
	jspl jspl_w_G13_1(.douta(w_G13_1[0]),.doutb(w_G13_1[1]),.din(w_G13_0[0]));
	jspl3 jspl3_w_G20_0(.douta(w_dff_A_U7WxENXP3_0),.doutb(w_G20_0[1]),.doutc(w_G20_0[2]),.din(G20));
	jspl3 jspl3_w_G20_1(.douta(w_G20_1[0]),.doutb(w_G20_1[1]),.doutc(w_dff_A_gKX85fBz5_2),.din(w_G20_0[0]));
	jspl3 jspl3_w_G20_2(.douta(w_G20_2[0]),.doutb(w_dff_A_Xs3u2aA27_1),.doutc(w_G20_2[2]),.din(w_G20_0[1]));
	jspl3 jspl3_w_G20_3(.douta(w_G20_3[0]),.doutb(w_dff_A_lo75t7xT1_1),.doutc(w_dff_A_cuKsTYLP9_2),.din(w_G20_0[2]));
	jspl3 jspl3_w_G20_4(.douta(w_dff_A_w57tCPB92_0),.doutb(w_dff_A_iypLFhgt0_1),.doutc(w_G20_4[2]),.din(w_G20_1[0]));
	jspl3 jspl3_w_G20_5(.douta(w_dff_A_ln2asg344_0),.doutb(w_dff_A_FGDdilbX4_1),.doutc(w_G20_5[2]),.din(w_G20_1[1]));
	jspl3 jspl3_w_G20_6(.douta(w_dff_A_N9Azsqpu1_0),.doutb(w_G20_6[1]),.doutc(w_G20_6[2]),.din(w_G20_1[2]));
	jspl jspl_w_G20_7(.douta(w_G20_7[0]),.doutb(w_G20_7[1]),.din(w_G20_2[0]));
	jspl3 jspl3_w_G33_0(.douta(w_dff_A_L884xvOs1_0),.doutb(w_G33_0[1]),.doutc(w_G33_0[2]),.din(G33));
	jspl3 jspl3_w_G33_1(.douta(w_G33_1[0]),.doutb(w_dff_A_jyy5vK6a4_1),.doutc(w_G33_1[2]),.din(w_G33_0[0]));
	jspl3 jspl3_w_G33_2(.douta(w_G33_2[0]),.doutb(w_G33_2[1]),.doutc(w_G33_2[2]),.din(w_G33_0[1]));
	jspl3 jspl3_w_G33_3(.douta(w_G33_3[0]),.doutb(w_G33_3[1]),.doutc(w_dff_A_YKI0fE2C8_2),.din(w_G33_0[2]));
	jspl3 jspl3_w_G33_4(.douta(w_G33_4[0]),.doutb(w_dff_A_b9LAaO2V4_1),.doutc(w_dff_A_o4VBRHSQ5_2),.din(w_G33_1[0]));
	jspl3 jspl3_w_G33_5(.douta(w_dff_A_cjnYpDZZ3_0),.doutb(w_G33_5[1]),.doutc(w_dff_A_S7K7j6zJ5_2),.din(w_G33_1[1]));
	jspl3 jspl3_w_G33_6(.douta(w_dff_A_vodn5zpv1_0),.doutb(w_dff_A_J9nVbyfr6_1),.doutc(w_G33_6[2]),.din(w_G33_1[2]));
	jspl3 jspl3_w_G33_7(.douta(w_G33_7[0]),.doutb(w_G33_7[1]),.doutc(w_G33_7[2]),.din(w_G33_2[0]));
	jspl3 jspl3_w_G33_8(.douta(w_dff_A_KXzl8J1t1_0),.doutb(w_G33_8[1]),.doutc(w_G33_8[2]),.din(w_G33_2[1]));
	jspl3 jspl3_w_G33_9(.douta(w_G33_9[0]),.doutb(w_G33_9[1]),.doutc(w_dff_A_RJ3ehxuJ6_2),.din(w_G33_2[2]));
	jspl3 jspl3_w_G33_10(.douta(w_dff_A_RIYLDndJ8_0),.doutb(w_dff_A_Hdd3lQoJ9_1),.doutc(w_G33_10[2]),.din(w_G33_3[0]));
	jspl3 jspl3_w_G33_11(.douta(w_G33_11[0]),.doutb(w_G33_11[1]),.doutc(w_G33_11[2]),.din(w_G33_3[1]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_dff_A_imXvUDCW9_1),.doutc(w_dff_A_bIepQwPZ9_2),.din(G41));
	jspl jspl_w_G41_1(.douta(w_G41_1[0]),.doutb(w_G41_1[1]),.din(w_G41_0[0]));
	jspl3 jspl3_w_G45_0(.douta(w_G45_0[0]),.doutb(w_dff_A_O7RBQmC53_1),.doutc(w_dff_A_mlsnI8yO0_2),.din(G45));
	jspl3 jspl3_w_G45_1(.douta(w_dff_A_Gg30chY37_0),.doutb(w_dff_A_zAnPpuHg8_1),.doutc(w_G45_1[2]),.din(w_G45_0[0]));
	jspl3 jspl3_w_G50_0(.douta(w_G50_0[0]),.doutb(w_dff_A_ceiHMDiR8_1),.doutc(w_G50_0[2]),.din(G50));
	jspl3 jspl3_w_G50_1(.douta(w_dff_A_cO4jwKc07_0),.doutb(w_G50_1[1]),.doutc(w_dff_A_k3YJBcmu3_2),.din(w_G50_0[0]));
	jspl3 jspl3_w_G50_2(.douta(w_dff_A_h0HBtqJs8_0),.doutb(w_G50_2[1]),.doutc(w_G50_2[2]),.din(w_G50_0[1]));
	jspl3 jspl3_w_G50_3(.douta(w_dff_A_ViKm35nZ0_0),.doutb(w_G50_3[1]),.doutc(w_dff_A_O3QSvosB8_2),.din(w_G50_0[2]));
	jspl3 jspl3_w_G50_4(.douta(w_dff_A_fRSggduI5_0),.doutb(w_dff_A_uDnNAuvx7_1),.doutc(w_G50_4[2]),.din(w_G50_1[0]));
	jspl3 jspl3_w_G50_5(.douta(w_G50_5[0]),.doutb(w_dff_A_RNGblkSf3_1),.doutc(w_G50_5[2]),.din(w_G50_1[1]));
	jspl3 jspl3_w_G58_0(.douta(w_G58_0[0]),.doutb(w_dff_A_QXcKkVHt5_1),.doutc(w_dff_A_XwAUHr957_2),.din(G58));
	jspl3 jspl3_w_G58_1(.douta(w_dff_A_QTvtvopw5_0),.doutb(w_G58_1[1]),.doutc(w_dff_A_dVMNW22K3_2),.din(w_G58_0[0]));
	jspl3 jspl3_w_G58_2(.douta(w_dff_A_SLHqwUK49_0),.doutb(w_G58_2[1]),.doutc(w_dff_A_gfeH5r0M2_2),.din(w_G58_0[1]));
	jspl3 jspl3_w_G58_3(.douta(w_dff_A_0J2BOCin4_0),.doutb(w_dff_A_NfVWJxMP8_1),.doutc(w_G58_3[2]),.din(w_G58_0[2]));
	jspl3 jspl3_w_G58_4(.douta(w_dff_A_3WNCWLUH0_0),.doutb(w_dff_A_8kvExLf64_1),.doutc(w_G58_4[2]),.din(w_G58_1[0]));
	jspl jspl_w_G58_5(.douta(w_G58_5[0]),.doutb(w_G58_5[1]),.din(w_G58_1[1]));
	jspl3 jspl3_w_G68_0(.douta(w_G68_0[0]),.doutb(w_G68_0[1]),.doutc(w_dff_A_nJpYmbT09_2),.din(G68));
	jspl3 jspl3_w_G68_1(.douta(w_dff_A_EXr1nqMF9_0),.doutb(w_G68_1[1]),.doutc(w_dff_A_O2WVEmuP0_2),.din(w_G68_0[0]));
	jspl3 jspl3_w_G68_2(.douta(w_G68_2[0]),.doutb(w_dff_A_6c3adLdN9_1),.doutc(w_dff_A_JUOYulXY2_2),.din(w_G68_0[1]));
	jspl3 jspl3_w_G68_3(.douta(w_G68_3[0]),.doutb(w_dff_A_3ljWBAJk4_1),.doutc(w_dff_A_YLSKHkFy7_2),.din(w_G68_0[2]));
	jspl3 jspl3_w_G68_4(.douta(w_dff_A_sVih4rfd4_0),.doutb(w_dff_A_BiYpS19j7_1),.doutc(w_G68_4[2]),.din(w_G68_1[0]));
	jspl jspl_w_G68_5(.douta(w_G68_5[0]),.doutb(w_G68_5[1]),.din(w_G68_1[1]));
	jspl3 jspl3_w_G77_0(.douta(w_G77_0[0]),.doutb(w_G77_0[1]),.doutc(w_G77_0[2]),.din(G77));
	jspl3 jspl3_w_G77_1(.douta(w_dff_A_yO1GxoUW4_0),.doutb(w_G77_1[1]),.doutc(w_dff_A_tDndV5yl1_2),.din(w_G77_0[0]));
	jspl3 jspl3_w_G77_2(.douta(w_G77_2[0]),.doutb(w_dff_A_2qfylIWC6_1),.doutc(w_dff_A_k3RzfDcU5_2),.din(w_G77_0[1]));
	jspl3 jspl3_w_G77_3(.douta(w_G77_3[0]),.doutb(w_dff_A_hIXBk1Sm1_1),.doutc(w_G77_3[2]),.din(w_G77_0[2]));
	jspl3 jspl3_w_G77_4(.douta(w_dff_A_3qbxSaiM9_0),.doutb(w_G77_4[1]),.doutc(w_G77_4[2]),.din(w_G77_1[0]));
	jspl jspl_w_G77_5(.douta(w_G77_5[0]),.doutb(w_G77_5[1]),.din(w_G77_1[1]));
	jspl3 jspl3_w_G87_0(.douta(w_dff_A_Ngq5RurS5_0),.doutb(w_G87_0[1]),.doutc(w_G87_0[2]),.din(G87));
	jspl3 jspl3_w_G87_1(.douta(w_G87_1[0]),.doutb(w_dff_A_PhMWxTnj9_1),.doutc(w_dff_A_0IN0JfWw8_2),.din(w_G87_0[0]));
	jspl3 jspl3_w_G87_2(.douta(w_dff_A_USAElrpB3_0),.doutb(w_dff_A_wKnIhUQ70_1),.doutc(w_G87_2[2]),.din(w_G87_0[1]));
	jspl3 jspl3_w_G87_3(.douta(w_dff_A_aExwiZ3Z6_0),.doutb(w_G87_3[1]),.doutc(w_dff_A_s2DAGwOv7_2),.din(w_G87_0[2]));
	jspl3 jspl3_w_G97_0(.douta(w_G97_0[0]),.doutb(w_dff_A_zFlKy9Tf6_1),.doutc(w_dff_A_37h6aHQw9_2),.din(G97));
	jspl3 jspl3_w_G97_1(.douta(w_G97_1[0]),.doutb(w_G97_1[1]),.doutc(w_dff_A_qFESAoza9_2),.din(w_G97_0[0]));
	jspl3 jspl3_w_G97_2(.douta(w_G97_2[0]),.doutb(w_G97_2[1]),.doutc(w_dff_A_nM5IVhfx6_2),.din(w_G97_0[1]));
	jspl3 jspl3_w_G97_3(.douta(w_dff_A_Gn9pDYYA7_0),.doutb(w_dff_A_rSAM8eBC8_1),.doutc(w_G97_3[2]),.din(w_G97_0[2]));
	jspl3 jspl3_w_G97_4(.douta(w_dff_A_mP813Pcd7_0),.doutb(w_G97_4[1]),.doutc(w_G97_4[2]),.din(w_G97_1[0]));
	jspl jspl_w_G97_5(.douta(w_dff_A_fbC376HG6_0),.doutb(w_G97_5[1]),.din(w_G97_1[1]));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_dff_A_t00ToI546_1),.doutc(w_dff_A_5RDm4RVr9_2),.din(G107));
	jspl3 jspl3_w_G107_1(.douta(w_G107_1[0]),.doutb(w_G107_1[1]),.doutc(w_dff_A_KLhsMzL80_2),.din(w_G107_0[0]));
	jspl3 jspl3_w_G107_2(.douta(w_G107_2[0]),.doutb(w_G107_2[1]),.doutc(w_dff_A_8nC7ayYu1_2),.din(w_G107_0[1]));
	jspl3 jspl3_w_G107_3(.douta(w_dff_A_HgI6wU3w3_0),.doutb(w_dff_A_vTk5FaV18_1),.doutc(w_G107_3[2]),.din(w_G107_0[2]));
	jspl3 jspl3_w_G107_4(.douta(w_dff_A_eoP6Xd8S5_0),.doutb(w_G107_4[1]),.doutc(w_G107_4[2]),.din(w_G107_1[0]));
	jspl jspl_w_G107_5(.douta(w_G107_5[0]),.doutb(w_G107_5[1]),.din(w_G107_1[1]));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_dff_A_QBQC4kG27_1),.doutc(w_dff_A_8pOBQB5E3_2),.din(G116));
	jspl3 jspl3_w_G116_1(.douta(w_G116_1[0]),.doutb(w_dff_A_wubsV4sU3_1),.doutc(w_dff_A_0FigtYqf8_2),.din(w_G116_0[0]));
	jspl3 jspl3_w_G116_2(.douta(w_G116_2[0]),.doutb(w_dff_A_Mokb2Ozp2_1),.doutc(w_dff_A_wPCjnRXx0_2),.din(w_G116_0[1]));
	jspl3 jspl3_w_G116_3(.douta(w_dff_A_ryAzrpiQ6_0),.doutb(w_G116_3[1]),.doutc(w_dff_A_fd8aelqm7_2),.din(w_G116_0[2]));
	jspl3 jspl3_w_G116_4(.douta(w_G116_4[0]),.doutb(w_G116_4[1]),.doutc(w_G116_4[2]),.din(w_G116_1[0]));
	jspl jspl_w_G125_0(.douta(w_G125_0[0]),.doutb(w_dff_A_zYWUnwFe9_1),.din(w_dff_B_KScad4zf5_2));
	jspl3 jspl3_w_G128_0(.douta(w_dff_A_rM240p1f9_0),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(w_dff_B_0VZex3Hm5_3));
	jspl3 jspl3_w_G132_0(.douta(w_G132_0[0]),.doutb(w_G132_0[1]),.doutc(w_G132_0[2]),.din(w_dff_B_Fqzti0kV8_3));
	jspl jspl_w_G132_1(.douta(w_G132_1[0]),.doutb(w_dff_A_hzAYjnOD2_1),.din(w_G132_0[0]));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(w_dff_B_Q4pTqb6Z2_3));
	jspl3 jspl3_w_G137_1(.douta(w_G137_1[0]),.doutb(w_dff_A_qfTcccIv9_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(w_dff_B_UfJBKIYt5_3));
	jspl3 jspl3_w_G143_1(.douta(w_dff_A_fBl11jYt5_0),.doutb(w_G143_1[1]),.doutc(w_dff_A_7O4GBKmN5_2),.din(w_G143_0[0]));
	jspl jspl_w_G143_2(.douta(w_G143_2[0]),.doutb(w_G143_2[1]),.din(w_G143_0[1]));
	jspl3 jspl3_w_G150_0(.douta(w_dff_A_99Lyr7EB8_0),.doutb(w_dff_A_KeaK6sWc8_1),.doutc(w_G150_0[2]),.din(G150));
	jspl3 jspl3_w_G150_1(.douta(w_G150_1[0]),.doutb(w_dff_A_hNX5uZgb5_1),.doutc(w_dff_A_57GtZJ4n5_2),.din(w_G150_0[0]));
	jspl3 jspl3_w_G150_2(.douta(w_G150_2[0]),.doutb(w_dff_A_iF5cVrWG1_1),.doutc(w_G150_2[2]),.din(w_G150_0[1]));
	jspl jspl_w_G150_3(.douta(w_dff_A_NYg96YUV4_0),.doutb(w_G150_3[1]),.din(w_G150_0[2]));
	jspl3 jspl3_w_G159_0(.douta(w_dff_A_pFsDiY7u2_0),.doutb(w_dff_A_YFMzVTqr9_1),.doutc(w_G159_0[2]),.din(w_dff_B_qEsBJxUD4_3));
	jspl3 jspl3_w_G159_1(.douta(w_G159_1[0]),.doutb(w_G159_1[1]),.doutc(w_G159_1[2]),.din(w_G159_0[0]));
	jspl3 jspl3_w_G159_2(.douta(w_G159_2[0]),.doutb(w_G159_2[1]),.doutc(w_G159_2[2]),.din(w_G159_0[1]));
	jspl3 jspl3_w_G159_3(.douta(w_dff_A_D7VmnP0H6_0),.doutb(w_dff_A_ag9PAe2Q7_1),.doutc(w_G159_3[2]),.din(w_G159_0[2]));
	jspl3 jspl3_w_G169_0(.douta(w_G169_0[0]),.doutb(w_dff_A_tbnSXAeN5_1),.doutc(w_dff_A_gYcfZmMb5_2),.din(G169));
	jspl jspl_w_G169_1(.douta(w_dff_A_0eQoAOf32_0),.doutb(w_G169_1[1]),.din(w_G169_0[0]));
	jspl3 jspl3_w_G179_0(.douta(w_dff_A_g2I0R6IE3_0),.doutb(w_G179_0[1]),.doutc(w_G179_0[2]),.din(G179));
	jspl3 jspl3_w_G179_1(.douta(w_G179_1[0]),.doutb(w_G179_1[1]),.doutc(w_G179_1[2]),.din(w_G179_0[0]));
	jspl3 jspl3_w_G179_2(.douta(w_dff_A_J9O08y4f3_0),.doutb(w_dff_A_Xfg6H6d67_1),.doutc(w_G179_2[2]),.din(w_G179_0[1]));
	jspl3 jspl3_w_G190_0(.douta(w_dff_A_e5MdD5iH7_0),.doutb(w_dff_A_J7ajIevY0_1),.doutc(w_G190_0[2]),.din(G190));
	jspl3 jspl3_w_G190_1(.douta(w_dff_A_nw8f0R964_0),.doutb(w_G190_1[1]),.doutc(w_G190_1[2]),.din(w_G190_0[0]));
	jspl3 jspl3_w_G190_2(.douta(w_G190_2[0]),.doutb(w_dff_A_BzFwJUiJ7_1),.doutc(w_dff_A_O8MIMKtL8_2),.din(w_G190_0[1]));
	jspl3 jspl3_w_G190_3(.douta(w_G190_3[0]),.doutb(w_dff_A_8Y5cjDrJ2_1),.doutc(w_dff_A_pX9m3u7g3_2),.din(w_G190_0[2]));
	jspl jspl_w_G190_4(.douta(w_dff_A_6bRW6Qnl2_0),.doutb(w_G190_4[1]),.din(w_G190_1[0]));
	jspl3 jspl3_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.doutc(w_dff_A_qRkE6gDE0_2),.din(G200));
	jspl3 jspl3_w_G200_1(.douta(w_dff_A_YqcSp3Kl9_0),.doutb(w_dff_A_nM2frNaL4_1),.doutc(w_G200_1[2]),.din(w_G200_0[0]));
	jspl3 jspl3_w_G200_2(.douta(w_G200_2[0]),.doutb(w_dff_A_DgfAJj4N8_1),.doutc(w_dff_A_9GwzyXxU8_2),.din(w_G200_0[1]));
	jspl3 jspl3_w_G200_3(.douta(w_G200_3[0]),.doutb(w_G200_3[1]),.doutc(w_G200_3[2]),.din(w_G200_0[2]));
	jspl3 jspl3_w_G200_4(.douta(w_G200_4[0]),.doutb(w_G200_4[1]),.doutc(w_G200_4[2]),.din(w_G200_1[0]));
	jspl3 jspl3_w_G213_0(.douta(w_dff_A_i7KpoBFg0_0),.doutb(w_G213_0[1]),.doutc(w_dff_A_OZZpiNyz2_2),.din(G213));
	jspl jspl_w_G223_0(.douta(w_G223_0[0]),.doutb(w_G223_0[1]),.din(w_dff_B_fru2YtIE1_2));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_dff_A_DGM43qRJ8_1),.doutc(w_dff_A_fJlaCSEw5_2),.din(G226));
	jspl jspl_w_G226_1(.douta(w_dff_A_xhqleR399_0),.doutb(w_G226_1[1]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G232_0(.douta(w_G232_0[0]),.doutb(w_dff_A_3ESCjbCr0_1),.doutc(w_dff_A_TFUnVYZP2_2),.din(G232));
	jspl3 jspl3_w_G232_1(.douta(w_dff_A_dzTU3Vk73_0),.doutb(w_dff_A_2feKBVo45_1),.doutc(w_G232_1[2]),.din(w_G232_0[0]));
	jspl3 jspl3_w_G238_0(.douta(w_G238_0[0]),.doutb(w_dff_A_M9xudvUV9_1),.doutc(w_dff_A_zG3jJkC47_2),.din(G238));
	jspl3 jspl3_w_G238_1(.douta(w_dff_A_SKieoeJM9_0),.doutb(w_G238_1[1]),.doutc(w_G238_1[2]),.din(w_G238_0[0]));
	jspl3 jspl3_w_G244_0(.douta(w_G244_0[0]),.doutb(w_dff_A_FjTqQqIS7_1),.doutc(w_dff_A_RKxoHzft5_2),.din(G244));
	jspl3 jspl3_w_G244_1(.douta(w_dff_A_XaWl6EhB4_0),.doutb(w_G244_1[1]),.doutc(w_G244_1[2]),.din(w_G244_0[0]));
	jspl3 jspl3_w_G250_0(.douta(w_dff_A_WgYvqrS63_0),.doutb(w_dff_A_72UFADII8_1),.doutc(w_G250_0[2]),.din(G250));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_dff_A_ltqoHmBF3_1),.doutc(w_dff_A_U2PfyQfO1_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_PVlXVh3K7_0),.doutb(w_dff_A_R8TMyVsb5_1),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G264_0(.douta(w_G264_0[0]),.doutb(w_dff_A_JKOTdtIu3_1),.doutc(w_dff_A_DpVal63g7_2),.din(G264));
	jspl jspl_w_G264_1(.douta(w_G264_1[0]),.doutb(w_G264_1[1]),.din(w_G264_0[0]));
	jspl3 jspl3_w_G270_0(.douta(w_dff_A_cQ54mkdH5_0),.doutb(w_G270_0[1]),.doutc(w_G270_0[2]),.din(G270));
	jspl3 jspl3_w_G274_0(.douta(w_dff_A_LfpceVR85_0),.doutb(w_G274_0[1]),.doutc(w_dff_A_wNbrbeh79_2),.din(G274));
	jspl3 jspl3_w_G283_0(.douta(w_dff_A_HFEcO3OZ4_0),.doutb(w_dff_A_FRy2ruUc6_1),.doutc(w_G283_0[2]),.din(G283));
	jspl3 jspl3_w_G283_1(.douta(w_G283_1[0]),.doutb(w_dff_A_aX2enYOS0_1),.doutc(w_G283_1[2]),.din(w_G283_0[0]));
	jspl3 jspl3_w_G283_2(.douta(w_dff_A_5d8bTIn96_0),.doutb(w_dff_A_WFItt2iM5_1),.doutc(w_G283_2[2]),.din(w_G283_0[1]));
	jspl3 jspl3_w_G283_3(.douta(w_dff_A_qJosGXVx0_0),.doutb(w_dff_A_qEGcM8sZ4_1),.doutc(w_G283_3[2]),.din(w_G283_0[2]));
	jspl3 jspl3_w_G294_0(.douta(w_dff_A_UoXAoSkh7_0),.doutb(w_dff_A_zA8cSDbK4_1),.doutc(w_G294_0[2]),.din(G294));
	jspl3 jspl3_w_G294_1(.douta(w_G294_1[0]),.doutb(w_dff_A_FGQPDyVV7_1),.doutc(w_G294_1[2]),.din(w_G294_0[0]));
	jspl3 jspl3_w_G294_2(.douta(w_dff_A_PhvWA9S78_0),.doutb(w_G294_2[1]),.doutc(w_G294_2[2]),.din(w_G294_0[1]));
	jspl jspl_w_G294_3(.douta(w_dff_A_Z0FLKKmW4_0),.doutb(w_G294_3[1]),.din(w_G294_0[2]));
	jspl3 jspl3_w_G303_0(.douta(w_dff_A_rs9LaVd82_0),.doutb(w_G303_0[1]),.doutc(w_dff_A_r4fvZwfG5_2),.din(G303));
	jspl3 jspl3_w_G303_1(.douta(w_G303_1[0]),.doutb(w_G303_1[1]),.doutc(w_G303_1[2]),.din(w_G303_0[0]));
	jspl3 jspl3_w_G303_2(.douta(w_dff_A_dRIFEpXE2_0),.doutb(w_dff_A_zHbiGjTa4_1),.doutc(w_G303_2[2]),.din(w_G303_0[1]));
	jspl3 jspl3_w_G311_0(.douta(w_G311_0[0]),.doutb(w_G311_0[1]),.doutc(w_G311_0[2]),.din(w_dff_B_dHAKO5Ky6_3));
	jspl3 jspl3_w_G311_1(.douta(w_G311_1[0]),.doutb(w_dff_A_XbIQ92Om5_1),.doutc(w_G311_1[2]),.din(w_G311_0[0]));
	jspl3 jspl3_w_G317_0(.douta(w_G317_0[0]),.doutb(w_G317_0[1]),.doutc(w_G317_0[2]),.din(w_dff_B_CDR6Suz05_3));
	jspl jspl_w_G317_1(.douta(w_dff_A_ph7TJQJV6_0),.doutb(w_G317_1[1]),.din(w_G317_0[0]));
	jspl3 jspl3_w_G322_0(.douta(w_dff_A_vhYSnYkN0_0),.doutb(w_G322_0[1]),.doutc(w_G322_0[2]),.din(w_dff_B_Y4As0ua57_3));
	jspl jspl_w_G326_0(.douta(w_dff_A_yyHutWcL6_0),.doutb(w_G326_0[1]),.din(w_dff_B_P0A9yaRt5_2));
	jspl jspl_w_G330_0(.douta(w_dff_A_ivacLBdj2_0),.doutb(w_G330_0[1]),.din(G330));
	jspl jspl_w_G343_0(.douta(w_G343_0[0]),.doutb(w_dff_A_hdHP6RrK9_1),.din(G343));
	jspl3 jspl3_w_G1698_0(.douta(w_G1698_0[0]),.doutb(w_G1698_0[1]),.doutc(w_dff_A_eZH5iZ0n7_2),.din(G1698));
	jspl jspl_w_G355_0(.douta(w_G355_0),.doutb(w_dff_A_VGKJsJxE9_1),.din(G355_fa_));
	jspl3 jspl3_w_G396_0(.douta(w_dff_A_lE3ItQU19_0),.doutb(w_G396_0[1]),.doutc(w_dff_A_xU860ofM7_2),.din(G396_fa_));
	jspl jspl_w_G384_0(.douta(w_dff_A_4vDcmayi0_0),.doutb(w_dff_A_du0s43qn6_1),.din(G384_fa_));
	jspl3 jspl3_w_G387_0(.douta(w_G387_0[0]),.doutb(w_G387_0[1]),.doutc(w_dff_A_FnlWl4Ri9_2),.din(G387_fa_));
	jspl3 jspl3_w_n72_0(.douta(w_n72_0[0]),.doutb(w_dff_A_EUoXFZbj8_1),.doutc(w_dff_A_OFAGcWOO5_2),.din(n72));
	jspl jspl_w_n72_1(.douta(w_n72_1[0]),.doutb(w_dff_A_Cy55RF5Q7_1),.din(w_n72_0[0]));
	jspl3 jspl3_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.doutc(w_dff_A_3meGaPFs8_2),.din(n73));
	jspl3 jspl3_w_n73_1(.douta(w_n73_1[0]),.doutb(w_dff_A_zyINY7Mr6_1),.doutc(w_n73_1[2]),.din(w_n73_0[0]));
	jspl3 jspl3_w_n73_2(.douta(w_dff_A_vmV6BBVp7_0),.doutb(w_n73_2[1]),.doutc(w_dff_A_w6X8EAcp6_2),.din(w_n73_0[1]));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_dff_A_3idra0BX3_1),.doutc(w_dff_A_cHL9pHTy1_2),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_dff_A_H77SgCYr7_1),.doutc(w_dff_A_OvbUSvio9_2),.din(n75));
	jspl jspl_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.din(w_n75_0[0]));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.din(n76));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl3 jspl3_w_n79_0(.douta(w_dff_A_BmhYXBOh6_0),.doutb(w_n79_0[1]),.doutc(w_n79_0[2]),.din(n79));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_dff_A_6XzsJmGb0_1),.doutc(w_dff_A_j1CPUTnK0_2),.din(n80));
	jspl jspl_w_n80_1(.douta(w_n80_1[0]),.doutb(w_n80_1[1]),.din(w_n80_0[0]));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_o5EKPjlR2_0),.doutb(w_n85_0[1]),.doutc(w_dff_A_6naw0bNr9_2),.din(n85));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n88_0(.douta(w_n88_0[0]),.doutb(w_dff_A_JLnUbvKH6_1),.doutc(w_dff_A_8vJy3UYI7_2),.din(n88));
	jspl jspl_w_n88_1(.douta(w_n88_1[0]),.doutb(w_n88_1[1]),.din(w_n88_0[0]));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_dff_A_vrlGWjLz1_1),.doutc(w_n91_0[2]),.din(n91));
	jspl3 jspl3_w_n91_1(.douta(w_dff_A_dnvwvo7A0_0),.doutb(w_n91_1[1]),.doutc(w_n91_1[2]),.din(w_n91_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n97_0(.douta(w_dff_A_NBWhMjeI7_0),.doutb(w_n97_0[1]),.doutc(w_n97_0[2]),.din(n97));
	jspl3 jspl3_w_n97_1(.douta(w_n97_1[0]),.doutb(w_dff_A_602sP49u2_1),.doutc(w_n97_1[2]),.din(w_n97_0[0]));
	jspl jspl_w_n97_2(.douta(w_n97_2[0]),.doutb(w_n97_2[1]),.din(w_n97_0[1]));
	jspl3 jspl3_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.doutc(w_n98_0[2]),.din(n98));
	jspl3 jspl3_w_n98_1(.douta(w_dff_A_wnamHytM4_0),.doutb(w_dff_A_Nhy7Pxuv0_1),.doutc(w_n98_1[2]),.din(w_n98_0[0]));
	jspl jspl_w_n98_2(.douta(w_dff_A_Fnp8WRIn0_0),.doutb(w_n98_2[1]),.din(w_n98_0[1]));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_dXo3rnxy2_1),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n105_0(.douta(w_dff_A_bOauCHnq3_0),.doutb(w_n105_0[1]),.doutc(w_dff_A_olsPP0wh9_2),.din(n105));
	jspl3 jspl3_w_n105_1(.douta(w_dff_A_DgwHk2E26_0),.doutb(w_n105_1[1]),.doutc(w_dff_A_yvlK8xgo9_2),.din(w_n105_0[0]));
	jspl jspl_w_n105_2(.douta(w_n105_2[0]),.doutb(w_n105_2[1]),.din(w_n105_0[1]));
	jspl jspl_w_n106_0(.douta(w_dff_A_k0B8T4cV2_0),.doutb(w_n106_0[1]),.din(n106));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl3 jspl3_w_n112_3(.douta(w_dff_A_xeprSQiT4_0),.doutb(w_dff_A_fGpFw67W2_1),.doutc(w_n112_3[2]),.din(w_n112_0[2]));
	jspl3 jspl3_w_n112_4(.douta(w_dff_A_Scn0bNSL3_0),.doutb(w_dff_A_3MA49UyW2_1),.doutc(w_n112_4[2]),.din(w_n112_1[0]));
	jspl3 jspl3_w_n112_5(.douta(w_n112_5[0]),.doutb(w_n112_5[1]),.doutc(w_dff_A_oio6ptqe1_2),.din(w_n112_1[1]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.doutc(w_n113_0[2]),.din(n113));
	jspl3 jspl3_w_n113_1(.douta(w_dff_A_31dEtmIx9_0),.doutb(w_dff_A_oaT70Ert9_1),.doutc(w_n113_1[2]),.din(w_n113_0[0]));
	jspl3 jspl3_w_n113_2(.douta(w_n113_2[0]),.doutb(w_n113_2[1]),.doutc(w_n113_2[2]),.din(w_n113_0[1]));
	jspl jspl_w_n113_3(.douta(w_n113_3[0]),.doutb(w_n113_3[1]),.din(w_n113_0[2]));
	jspl3 jspl3_w_n114_0(.douta(w_n114_0[0]),.doutb(w_dff_A_ruaDa1ua8_1),.doutc(w_n114_0[2]),.din(n114));
	jspl3 jspl3_w_n114_1(.douta(w_dff_A_FHTOnRU44_0),.doutb(w_n114_1[1]),.doutc(w_n114_1[2]),.din(w_n114_0[0]));
	jspl3 jspl3_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.doutc(w_dff_A_sflOr6SE6_2),.din(n115));
	jspl jspl_w_n115_1(.douta(w_n115_1[0]),.doutb(w_n115_1[1]),.din(w_n115_0[0]));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_dff_A_XPpM07ww0_1),.din(n116));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl3 jspl3_w_n121_0(.douta(w_dff_A_ccXMLJM11_0),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.doutc(w_n122_0[2]),.din(n122));
	jspl jspl_w_n122_1(.douta(w_n122_1[0]),.doutb(w_n122_1[1]),.din(w_n122_0[0]));
	jspl3 jspl3_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.doutc(w_n123_0[2]),.din(n123));
	jspl3 jspl3_w_n123_1(.douta(w_n123_1[0]),.doutb(w_n123_1[1]),.doutc(w_n123_1[2]),.din(w_n123_0[0]));
	jspl jspl_w_n131_0(.douta(w_dff_A_R8JEbloF5_0),.doutb(w_n131_0[1]),.din(n131));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_dff_A_pt9RtHEF4_1),.din(n135));
	jspl3 jspl3_w_n137_0(.douta(w_n137_0[0]),.doutb(w_n137_0[1]),.doutc(w_n137_0[2]),.din(n137));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(w_dff_B_Bm1gAG0j2_2));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_aWjUpErp0_1),.doutc(w_dff_A_EF4gWOik0_2),.din(n146));
	jspl3 jspl3_w_n146_1(.douta(w_n146_1[0]),.doutb(w_dff_A_xTp5TZ9O0_1),.doutc(w_dff_A_fzJDj07o3_2),.din(w_n146_0[0]));
	jspl3 jspl3_w_n146_2(.douta(w_n146_2[0]),.doutb(w_n146_2[1]),.doutc(w_n146_2[2]),.din(w_n146_0[1]));
	jspl3 jspl3_w_n146_3(.douta(w_n146_3[0]),.doutb(w_n146_3[1]),.doutc(w_n146_3[2]),.din(w_n146_0[2]));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_dff_A_Zcca7dj56_1),.doutc(w_dff_A_gOULqPpa3_2),.din(n147));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_dff_A_cRzoOTxt2_0),.doutb(w_dff_A_ch7PBlMN5_1),.doutc(w_n148_1[2]),.din(w_n148_0[0]));
	jspl3 jspl3_w_n148_2(.douta(w_n148_2[0]),.doutb(w_n148_2[1]),.doutc(w_n148_2[2]),.din(w_n148_0[1]));
	jspl3 jspl3_w_n148_3(.douta(w_dff_A_7dahFntp7_0),.doutb(w_n148_3[1]),.doutc(w_dff_A_dzJCSBPn5_2),.din(w_n148_0[2]));
	jspl3 jspl3_w_n148_4(.douta(w_n148_4[0]),.doutb(w_n148_4[1]),.doutc(w_n148_4[2]),.din(w_n148_1[0]));
	jspl3 jspl3_w_n148_5(.douta(w_n148_5[0]),.doutb(w_dff_A_tblrHz7F0_1),.doutc(w_dff_A_kXzz8afe8_2),.din(w_n148_1[1]));
	jspl3 jspl3_w_n148_6(.douta(w_n148_6[0]),.doutb(w_n148_6[1]),.doutc(w_n148_6[2]),.din(w_n148_1[2]));
	jspl3 jspl3_w_n148_7(.douta(w_n148_7[0]),.doutb(w_n148_7[1]),.doutc(w_n148_7[2]),.din(w_n148_2[0]));
	jspl3 jspl3_w_n148_8(.douta(w_n148_8[0]),.doutb(w_dff_A_7iLGToeL6_1),.doutc(w_n148_8[2]),.din(w_n148_2[1]));
	jspl3 jspl3_w_n148_9(.douta(w_n148_9[0]),.doutb(w_n148_9[1]),.doutc(w_n148_9[2]),.din(w_n148_2[2]));
	jspl3 jspl3_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.doutc(w_n149_0[2]),.din(n149));
	jspl3 jspl3_w_n149_1(.douta(w_n149_1[0]),.doutb(w_dff_A_s0awC98P6_1),.doutc(w_n149_1[2]),.din(w_n149_0[0]));
	jspl jspl_w_n149_2(.douta(w_dff_A_SOrcP7xY6_0),.doutb(w_n149_2[1]),.din(w_n149_0[1]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_TQ9Ulg3a7_1),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_dff_A_qojIAw5P2_1),.doutc(w_dff_A_LQBuzSCm1_2),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_n151_2[0]),.doutb(w_n151_2[1]),.doutc(w_n151_2[2]),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_dff_A_iUfZNA4n8_0),.doutb(w_dff_A_LdnhFLWB7_1),.doutc(w_n151_3[2]),.din(w_n151_0[2]));
	jspl3 jspl3_w_n151_4(.douta(w_n151_4[0]),.doutb(w_n151_4[1]),.doutc(w_dff_A_MvEArPr95_2),.din(w_n151_1[0]));
	jspl3 jspl3_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.doutc(w_n152_0[2]),.din(n152));
	jspl3 jspl3_w_n152_1(.douta(w_n152_1[0]),.doutb(w_n152_1[1]),.doutc(w_n152_1[2]),.din(w_n152_0[0]));
	jspl3 jspl3_w_n152_2(.douta(w_n152_2[0]),.doutb(w_n152_2[1]),.doutc(w_n152_2[2]),.din(w_n152_0[1]));
	jspl jspl_w_n152_3(.douta(w_n152_3[0]),.doutb(w_n152_3[1]),.din(w_n152_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(n154));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl3 jspl3_w_n155_1(.douta(w_n155_1[0]),.doutb(w_n155_1[1]),.doutc(w_n155_1[2]),.din(w_n155_0[0]));
	jspl3 jspl3_w_n155_2(.douta(w_n155_2[0]),.doutb(w_n155_2[1]),.doutc(w_n155_2[2]),.din(w_n155_0[1]));
	jspl jspl_w_n155_3(.douta(w_n155_3[0]),.doutb(w_n155_3[1]),.din(w_n155_0[2]));
	jspl3 jspl3_w_n157_0(.douta(w_dff_A_IC5fUeBa9_0),.doutb(w_n157_0[1]),.doutc(w_dff_A_mjO8ion64_2),.din(n157));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_dff_A_AkNA0WSt5_2),.din(n161));
	jspl jspl_w_n161_1(.douta(w_n161_1[0]),.doutb(w_n161_1[1]),.din(w_n161_0[0]));
	jspl3 jspl3_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.doutc(w_n162_0[2]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_dff_A_plqwpa2X5_0),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_dff_A_HO9wEOsL3_1),.doutc(w_dff_A_y18LBZqP9_2),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_dff_A_Lrq5l9tN6_2),.din(w_n166_0[1]));
	jspl jspl_w_n166_3(.douta(w_dff_A_JZDmjjWv3_0),.doutb(w_n166_3[1]),.din(w_n166_0[2]));
	jspl3 jspl3_w_n170_0(.douta(w_dff_A_OEIpwxEF5_0),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(w_dff_B_Mf2fnBMK2_2));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_dff_A_aLKewj3f7_1),.doutc(w_dff_A_ldhGD3Gr7_2),.din(n179));
	jspl3 jspl3_w_n179_1(.douta(w_n179_1[0]),.doutb(w_n179_1[1]),.doutc(w_n179_1[2]),.din(w_n179_0[0]));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.doutc(w_n185_0[2]),.din(n185));
	jspl3 jspl3_w_n185_1(.douta(w_n185_1[0]),.doutb(w_n185_1[1]),.doutc(w_dff_A_bHunUFF88_2),.din(w_n185_0[0]));
	jspl3 jspl3_w_n185_2(.douta(w_n185_2[0]),.doutb(w_dff_A_ExKRS7R52_1),.doutc(w_n185_2[2]),.din(w_n185_0[1]));
	jspl3 jspl3_w_n185_3(.douta(w_n185_3[0]),.doutb(w_n185_3[1]),.doutc(w_n185_3[2]),.din(w_n185_0[2]));
	jspl3 jspl3_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.doutc(w_dff_A_es4OKvcI0_2),.din(n189));
	jspl3 jspl3_w_n189_1(.douta(w_n189_1[0]),.doutb(w_dff_A_3U20ts2s3_1),.doutc(w_n189_1[2]),.din(w_n189_0[0]));
	jspl jspl_w_n189_2(.douta(w_dff_A_0ImIa9oz1_0),.doutb(w_n189_2[1]),.din(w_n189_0[1]));
	jspl3 jspl3_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.doutc(w_n190_0[2]),.din(n190));
	jspl3 jspl3_w_n190_1(.douta(w_n190_1[0]),.doutb(w_dff_A_oUx6ewKo9_1),.doutc(w_n190_1[2]),.din(w_n190_0[0]));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_dff_A_jXJ1oX4K0_0),.doutb(w_n196_0[1]),.doutc(w_dff_A_vV1USWCc7_2),.din(w_dff_B_gHcHtbaM1_3));
	jspl3 jspl3_w_n196_1(.douta(w_dff_A_ofqVPrrA0_0),.doutb(w_dff_A_5oFpw9a35_1),.doutc(w_n196_1[2]),.din(w_n196_0[0]));
	jspl3 jspl3_w_n196_2(.douta(w_dff_A_Yu58xckM0_0),.doutb(w_dff_A_5DkLtjcb4_1),.doutc(w_n196_2[2]),.din(w_n196_0[1]));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_n197_1[0]),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n199_1(.douta(w_n199_1[0]),.doutb(w_n199_1[1]),.din(w_n199_0[0]));
	jspl jspl_w_n201_0(.douta(w_dff_A_yBIm5AGK6_0),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n205_0(.douta(w_dff_A_xlZw4z332_0),.doutb(w_n205_0[1]),.din(w_dff_B_VCunKxQB3_2));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl3 jspl3_w_n210_0(.douta(w_dff_A_nBJU71419_0),.doutb(w_n210_0[1]),.doutc(w_n210_0[2]),.din(n210));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_dff_A_n7LAqGNU5_1),.din(n213));
	jspl jspl_w_n214_0(.douta(w_n214_0[0]),.doutb(w_dff_A_Qdhww1xq6_1),.din(n214));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl3 jspl3_w_n221_0(.douta(w_dff_A_wRipiJfK3_0),.doutb(w_dff_A_wmPnpOg62_1),.doutc(w_n221_0[2]),.din(n221));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_dff_A_amvJWUy39_1),.din(n228));
	jspl3 jspl3_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.doutc(w_n229_0[2]),.din(n229));
	jspl jspl_w_n230_0(.douta(w_dff_A_bf5y3ZLr2_0),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.doutc(w_n231_0[2]),.din(n231));
	jspl3 jspl3_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.doutc(w_n234_0[2]),.din(n234));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(n241));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl jspl_w_n246_1(.douta(w_n246_1[0]),.doutb(w_n246_1[1]),.din(w_n246_0[0]));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_XWyL3vEe4_2));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_dff_A_IQNMlTkt4_1),.din(n255));
	jspl jspl_w_n257_0(.douta(w_dff_A_JmzGA6ll1_0),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n259_0(.douta(w_dff_A_2284LzIR3_0),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n262_0(.douta(w_dff_A_Zr3jYwrt4_0),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.doutc(w_n269_1[2]),.din(w_n269_0[0]));
	jspl jspl_w_n270_0(.douta(w_dff_A_SAu8rnnx7_0),.doutb(w_n270_0[1]),.din(w_dff_B_JTvsNzW86_2));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_n271_1[0]),.doutb(w_n271_1[1]),.doutc(w_n271_1[2]),.din(w_n271_0[0]));
	jspl3 jspl3_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_CvAUyHMO4_1),.doutc(w_n274_0[2]),.din(n274));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(n278));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(n279));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_dff_A_aWCZ3PV36_1),.din(n281));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n288_1(.douta(w_n288_1[0]),.doutb(w_n288_1[1]),.din(w_n288_0[0]));
	jspl jspl_w_n296_0(.douta(w_dff_A_KluREwqb8_0),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n298_0(.douta(w_dff_A_BjWdFFvn0_0),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_dff_A_4V7aPM779_1),.din(n300));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_JyxRLC5D6_1),.din(n303));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_dff_A_r9xSnZwN3_1),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n334_0(.douta(w_dff_A_UaLXOGn53_0),.doutb(w_n334_0[1]),.din(n334));
	jspl jspl_w_n339_0(.douta(w_dff_A_scipC3JV3_0),.doutb(w_n339_0[1]),.din(n339));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl jspl_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.din(w_n355_0[0]));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_dff_A_uYaC6xKx9_1),.din(n374));
	jspl jspl_w_n381_0(.douta(w_n381_0[0]),.doutb(w_n381_0[1]),.din(n381));
	jspl3 jspl3_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.doutc(w_n382_0[2]),.din(n382));
	jspl jspl_w_n382_1(.douta(w_n382_1[0]),.doutb(w_n382_1[1]),.din(w_n382_0[0]));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl jspl_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(w_dff_B_q5J8ugWw8_2));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_dff_A_ZIQFC32R1_1),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n407_0(.douta(w_n407_0[0]),.doutb(w_dff_A_RstvUsjn8_1),.doutc(w_dff_A_OUBqBLoT3_2),.din(n407));
	jspl3 jspl3_w_n407_1(.douta(w_dff_A_QYNBuYWH1_0),.doutb(w_dff_A_aqXJWKtH7_1),.doutc(w_n407_1[2]),.din(w_n407_0[0]));
	jspl jspl_w_n407_2(.douta(w_n407_2[0]),.doutb(w_n407_2[1]),.din(w_n407_0[1]));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(n412));
	jspl3 jspl3_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jspl jspl_w_n420_1(.douta(w_n420_1[0]),.doutb(w_n420_1[1]),.din(w_n420_0[0]));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_dff_A_Nog6MXY70_1),.doutc(w_dff_A_n6eLtSK16_2),.din(n425));
	jspl3 jspl3_w_n425_1(.douta(w_dff_A_2tBscZ9S4_0),.doutb(w_dff_A_IVH6G14y3_1),.doutc(w_n425_1[2]),.din(w_n425_0[0]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl jspl_w_n430_0(.douta(w_dff_A_cpviNkYV1_0),.doutb(w_n430_0[1]),.din(w_dff_B_Qrej3fvK6_2));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_dff_A_Omws4HRf0_1),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_dff_A_jdrnQAet0_1),.doutc(w_n439_0[2]),.din(n439));
	jspl jspl_w_n439_1(.douta(w_n439_1[0]),.doutb(w_n439_1[1]),.din(w_n439_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl3 jspl3_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.doutc(w_n455_0[2]),.din(n455));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(n474));
	jspl jspl_w_n475_0(.douta(w_n475_0[0]),.doutb(w_n475_0[1]),.din(n475));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(n479));
	jspl jspl_w_n483_0(.douta(w_dff_A_umKsocQE8_0),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl3 jspl3_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.doutc(w_n492_0[2]),.din(n492));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n516_0(.douta(w_dff_A_mDKt5XaW3_0),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n519_0(.douta(w_n519_0[0]),.doutb(w_dff_A_08DYid1T7_1),.doutc(w_dff_A_54pKiNtS3_2),.din(n519));
	jspl3 jspl3_w_n519_1(.douta(w_dff_A_l8FyxM895_0),.doutb(w_n519_1[1]),.doutc(w_n519_1[2]),.din(w_n519_0[0]));
	jspl jspl_w_n523_0(.douta(w_dff_A_hGqcwpXw6_0),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_dff_A_5FWxVWEW6_1),.din(n524));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_dff_A_QuFQc92y8_1),.din(n532));
	jspl jspl_w_n534_0(.douta(w_dff_A_QCZ4uVcY2_0),.doutb(w_n534_0[1]),.din(n534));
	jspl3 jspl3_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.doutc(w_n536_0[2]),.din(n536));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_dff_A_C0LML8KC2_1),.din(n541));
	jspl3 jspl3_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.doutc(w_n542_0[2]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n548_0(.douta(w_dff_A_tzrtAI7m3_0),.doutb(w_n548_0[1]),.doutc(w_n548_0[2]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl3 jspl3_w_n552_0(.douta(w_n552_0[0]),.doutb(w_dff_A_DLDWHXGW0_1),.doutc(w_dff_A_bbdjmFzC1_2),.din(n552));
	jspl jspl_w_n552_1(.douta(w_n552_1[0]),.doutb(w_n552_1[1]),.din(w_n552_0[0]));
	jspl3 jspl3_w_n553_0(.douta(w_dff_A_9d4p2KhZ4_0),.doutb(w_n553_0[1]),.doutc(w_dff_A_hDnjk1EL9_2),.din(n553));
	jspl3 jspl3_w_n553_1(.douta(w_n553_1[0]),.doutb(w_n553_1[1]),.doutc(w_n553_1[2]),.din(w_n553_0[0]));
	jspl3 jspl3_w_n553_2(.douta(w_dff_A_LuFLmaxL6_0),.doutb(w_dff_A_NKo3CyIm1_1),.doutc(w_n553_2[2]),.din(w_n553_0[1]));
	jspl3 jspl3_w_n554_0(.douta(w_dff_A_wpfbVsDK0_0),.doutb(w_dff_A_vR3aIkMQ4_1),.doutc(w_n554_0[2]),.din(w_dff_B_3sFmpLJj0_3));
	jspl3 jspl3_w_n554_1(.douta(w_n554_1[0]),.doutb(w_n554_1[1]),.doutc(w_dff_A_SAJ9ZYRz3_2),.din(w_n554_0[0]));
	jspl3 jspl3_w_n554_2(.douta(w_n554_2[0]),.doutb(w_dff_A_tcJ3l1fM8_1),.doutc(w_dff_A_EgEJlBtd7_2),.din(w_n554_0[1]));
	jspl3 jspl3_w_n554_3(.douta(w_n554_3[0]),.doutb(w_dff_A_VCWSou9t2_1),.doutc(w_dff_A_21XGM9dY5_2),.din(w_n554_0[2]));
	jspl jspl_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.din(w_dff_B_ce4VxpCZ8_2));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl3 jspl3_w_n563_0(.douta(w_n563_0[0]),.doutb(w_dff_A_5IFVUyto1_1),.doutc(w_dff_A_6Uj6uu5l7_2),.din(n563));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_xeZgGkv54_1),.din(n564));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(w_dff_B_ixLNvbGt5_2));
	jspl jspl_w_n567_0(.douta(w_dff_A_Mr9KwjKC5_0),.doutb(w_n567_0[1]),.din(n567));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_n571_0[2]),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n576_1(.douta(w_n576_1[0]),.doutb(w_n576_1[1]),.din(w_n576_0[0]));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_dff_A_jNGD2hGt5_2),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n589_0(.douta(w_n589_0[0]),.doutb(w_n589_0[1]),.doutc(w_n589_0[2]),.din(n589));
	jspl3 jspl3_w_n589_1(.douta(w_dff_A_vSvLhwb24_0),.doutb(w_n589_1[1]),.doutc(w_n589_1[2]),.din(w_n589_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_dff_A_JNRB8m2A6_1),.doutc(w_dff_A_2rQ3bUW76_2),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_dff_A_XVsKrCdE7_0),.doutb(w_n592_0[1]),.doutc(w_dff_A_8uzhtFKJ3_2),.din(n592));
	jspl3 jspl3_w_n592_1(.douta(w_dff_A_hhZyU8L87_0),.doutb(w_dff_A_jQ3tBIKF0_1),.doutc(w_n592_1[2]),.din(w_n592_0[0]));
	jspl jspl_w_n592_2(.douta(w_n592_2[0]),.doutb(w_n592_2[1]),.din(w_n592_0[1]));
	jspl3 jspl3_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.doutc(w_n593_0[2]),.din(n593));
	jspl jspl_w_n602_0(.douta(w_dff_A_8ZO8nfsg0_0),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n603_0(.douta(w_dff_A_5a96gD1R9_0),.doutb(w_n603_0[1]),.doutc(w_dff_A_G1RDL8658_2),.din(n603));
	jspl3 jspl3_w_n603_1(.douta(w_dff_A_dYboeQ0R9_0),.doutb(w_n603_1[1]),.doutc(w_n603_1[2]),.din(w_n603_0[0]));
	jspl jspl_w_n603_2(.douta(w_dff_A_rWmU1MjV1_0),.doutb(w_n603_2[1]),.din(w_n603_0[1]));
	jspl3 jspl3_w_n604_0(.douta(w_dff_A_ZrQMDoap6_0),.doutb(w_n604_0[1]),.doutc(w_dff_A_GCtHfPh14_2),.din(n604));
	jspl3 jspl3_w_n604_1(.douta(w_dff_A_SYDBoXsz1_0),.doutb(w_n604_1[1]),.doutc(w_dff_A_nKyYHsfW0_2),.din(w_n604_0[0]));
	jspl jspl_w_n604_2(.douta(w_dff_A_id0GhgZb4_0),.doutb(w_n604_2[1]),.din(w_n604_0[1]));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_dff_A_H2OdbD9J3_2),.din(w_n605_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_dff_A_mquicPis4_1),.doutc(w_dff_A_cVKG9rir9_2),.din(n608));
	jspl3 jspl3_w_n608_1(.douta(w_dff_A_UK7zN0hx1_0),.doutb(w_n608_1[1]),.doutc(w_dff_A_JRZ2oKPU4_2),.din(w_n608_0[0]));
	jspl3 jspl3_w_n612_0(.douta(w_n612_0[0]),.doutb(w_dff_A_xYUjHr2C0_1),.doutc(w_n612_0[2]),.din(n612));
	jspl3 jspl3_w_n612_1(.douta(w_dff_A_oB6lzMDA6_0),.doutb(w_dff_A_AJINMCdz2_1),.doutc(w_n612_1[2]),.din(w_n612_0[0]));
	jspl3 jspl3_w_n612_2(.douta(w_n612_2[0]),.doutb(w_n612_2[1]),.doutc(w_n612_2[2]),.din(w_n612_0[1]));
	jspl3 jspl3_w_n612_3(.douta(w_dff_A_TD28eZi25_0),.doutb(w_n612_3[1]),.doutc(w_dff_A_TJa5PZqy0_2),.din(w_n612_0[2]));
	jspl jspl_w_n612_4(.douta(w_n612_4[0]),.doutb(w_dff_A_Jnrfl8BP3_1),.din(w_n612_1[0]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl jspl_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.din(w_n613_0[0]));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_dff_A_OFz0DY0G5_1),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl3 jspl3_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.doutc(w_n617_1[2]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n617_2(.douta(w_n617_2[0]),.doutb(w_n617_2[1]),.doutc(w_n617_2[2]),.din(w_n617_0[1]));
	jspl3 jspl3_w_n617_3(.douta(w_n617_3[0]),.doutb(w_n617_3[1]),.doutc(w_n617_3[2]),.din(w_n617_0[2]));
	jspl3 jspl3_w_n617_4(.douta(w_n617_4[0]),.doutb(w_n617_4[1]),.doutc(w_n617_4[2]),.din(w_n617_1[0]));
	jspl3 jspl3_w_n617_5(.douta(w_n617_5[0]),.doutb(w_n617_5[1]),.doutc(w_n617_5[2]),.din(w_n617_1[1]));
	jspl jspl_w_n617_6(.douta(w_n617_6[0]),.doutb(w_n617_6[1]),.din(w_n617_1[2]));
	jspl jspl_w_n619_0(.douta(w_dff_A_5A63NY9a2_0),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl3 jspl3_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.doutc(w_n623_0[2]),.din(n623));
	jspl3 jspl3_w_n623_1(.douta(w_n623_1[0]),.doutb(w_n623_1[1]),.doutc(w_n623_1[2]),.din(w_n623_0[0]));
	jspl3 jspl3_w_n623_2(.douta(w_n623_2[0]),.doutb(w_n623_2[1]),.doutc(w_n623_2[2]),.din(w_n623_0[1]));
	jspl3 jspl3_w_n623_3(.douta(w_n623_3[0]),.doutb(w_n623_3[1]),.doutc(w_n623_3[2]),.din(w_n623_0[2]));
	jspl3 jspl3_w_n623_4(.douta(w_n623_4[0]),.doutb(w_n623_4[1]),.doutc(w_n623_4[2]),.din(w_n623_1[0]));
	jspl jspl_w_n623_5(.douta(w_n623_5[0]),.doutb(w_n623_5[1]),.din(w_n623_1[1]));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(n626));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl3 jspl3_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.doutc(w_n627_1[2]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n627_2(.douta(w_n627_2[0]),.doutb(w_n627_2[1]),.doutc(w_n627_2[2]),.din(w_n627_0[1]));
	jspl3 jspl3_w_n627_3(.douta(w_n627_3[0]),.doutb(w_n627_3[1]),.doutc(w_n627_3[2]),.din(w_n627_0[2]));
	jspl3 jspl3_w_n627_4(.douta(w_n627_4[0]),.doutb(w_n627_4[1]),.doutc(w_n627_4[2]),.din(w_n627_1[0]));
	jspl3 jspl3_w_n627_5(.douta(w_n627_5[0]),.doutb(w_n627_5[1]),.doutc(w_n627_5[2]),.din(w_n627_1[1]));
	jspl3 jspl3_w_n627_6(.douta(w_n627_6[0]),.doutb(w_n627_6[1]),.doutc(w_n627_6[2]),.din(w_n627_1[2]));
	jspl jspl_w_n627_7(.douta(w_n627_7[0]),.doutb(w_n627_7[1]),.din(w_n627_2[0]));
	jspl3 jspl3_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.doutc(w_n631_0[2]),.din(n631));
	jspl3 jspl3_w_n631_1(.douta(w_n631_1[0]),.doutb(w_n631_1[1]),.doutc(w_n631_1[2]),.din(w_n631_0[0]));
	jspl3 jspl3_w_n631_2(.douta(w_n631_2[0]),.doutb(w_n631_2[1]),.doutc(w_n631_2[2]),.din(w_n631_0[1]));
	jspl3 jspl3_w_n631_3(.douta(w_n631_3[0]),.doutb(w_n631_3[1]),.doutc(w_n631_3[2]),.din(w_n631_0[2]));
	jspl3 jspl3_w_n631_4(.douta(w_n631_4[0]),.doutb(w_n631_4[1]),.doutc(w_n631_4[2]),.din(w_n631_1[0]));
	jspl3 jspl3_w_n631_5(.douta(w_n631_5[0]),.doutb(w_n631_5[1]),.doutc(w_n631_5[2]),.din(w_n631_1[1]));
	jspl3 jspl3_w_n631_6(.douta(w_n631_6[0]),.doutb(w_n631_6[1]),.doutc(w_n631_6[2]),.din(w_n631_1[2]));
	jspl jspl_w_n631_7(.douta(w_n631_7[0]),.doutb(w_n631_7[1]),.din(w_n631_2[0]));
	jspl3 jspl3_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.doutc(w_n634_0[2]),.din(n634));
	jspl3 jspl3_w_n634_1(.douta(w_n634_1[0]),.doutb(w_n634_1[1]),.doutc(w_n634_1[2]),.din(w_n634_0[0]));
	jspl3 jspl3_w_n634_2(.douta(w_n634_2[0]),.doutb(w_n634_2[1]),.doutc(w_n634_2[2]),.din(w_n634_0[1]));
	jspl3 jspl3_w_n634_3(.douta(w_n634_3[0]),.doutb(w_n634_3[1]),.doutc(w_n634_3[2]),.din(w_n634_0[2]));
	jspl jspl_w_n634_4(.douta(w_n634_4[0]),.doutb(w_n634_4[1]),.din(w_n634_1[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n636_1(.douta(w_n636_1[0]),.doutb(w_n636_1[1]),.doutc(w_n636_1[2]),.din(w_n636_0[0]));
	jspl3 jspl3_w_n636_2(.douta(w_n636_2[0]),.doutb(w_n636_2[1]),.doutc(w_n636_2[2]),.din(w_n636_0[1]));
	jspl3 jspl3_w_n636_3(.douta(w_n636_3[0]),.doutb(w_n636_3[1]),.doutc(w_n636_3[2]),.din(w_n636_0[2]));
	jspl3 jspl3_w_n636_4(.douta(w_n636_4[0]),.doutb(w_n636_4[1]),.doutc(w_n636_4[2]),.din(w_n636_1[0]));
	jspl3 jspl3_w_n636_5(.douta(w_n636_5[0]),.doutb(w_n636_5[1]),.doutc(w_n636_5[2]),.din(w_n636_1[1]));
	jspl3 jspl3_w_n636_6(.douta(w_n636_6[0]),.doutb(w_n636_6[1]),.doutc(w_n636_6[2]),.din(w_n636_1[2]));
	jspl jspl_w_n636_7(.douta(w_n636_7[0]),.doutb(w_n636_7[1]),.din(w_n636_2[0]));
	jspl jspl_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.din(n639));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl3 jspl3_w_n640_2(.douta(w_n640_2[0]),.doutb(w_n640_2[1]),.doutc(w_n640_2[2]),.din(w_n640_0[1]));
	jspl3 jspl3_w_n640_3(.douta(w_n640_3[0]),.doutb(w_n640_3[1]),.doutc(w_n640_3[2]),.din(w_n640_0[2]));
	jspl3 jspl3_w_n640_4(.douta(w_n640_4[0]),.doutb(w_n640_4[1]),.doutc(w_n640_4[2]),.din(w_n640_1[0]));
	jspl3 jspl3_w_n640_5(.douta(w_n640_5[0]),.doutb(w_n640_5[1]),.doutc(w_n640_5[2]),.din(w_n640_1[1]));
	jspl3 jspl3_w_n640_6(.douta(w_n640_6[0]),.doutb(w_n640_6[1]),.doutc(w_n640_6[2]),.din(w_n640_1[2]));
	jspl jspl_w_n640_7(.douta(w_n640_7[0]),.doutb(w_n640_7[1]),.din(w_n640_2[0]));
	jspl3 jspl3_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.doutc(w_n642_0[2]),.din(n642));
	jspl3 jspl3_w_n642_1(.douta(w_n642_1[0]),.doutb(w_n642_1[1]),.doutc(w_n642_1[2]),.din(w_n642_0[0]));
	jspl3 jspl3_w_n642_2(.douta(w_n642_2[0]),.doutb(w_n642_2[1]),.doutc(w_n642_2[2]),.din(w_n642_0[1]));
	jspl3 jspl3_w_n642_3(.douta(w_n642_3[0]),.doutb(w_n642_3[1]),.doutc(w_n642_3[2]),.din(w_n642_0[2]));
	jspl3 jspl3_w_n642_4(.douta(w_n642_4[0]),.doutb(w_n642_4[1]),.doutc(w_n642_4[2]),.din(w_n642_1[0]));
	jspl3 jspl3_w_n642_5(.douta(w_n642_5[0]),.doutb(w_n642_5[1]),.doutc(w_n642_5[2]),.din(w_n642_1[1]));
	jspl3 jspl3_w_n642_6(.douta(w_n642_6[0]),.doutb(w_n642_6[1]),.doutc(w_n642_6[2]),.din(w_n642_1[2]));
	jspl jspl_w_n642_7(.douta(w_n642_7[0]),.doutb(w_n642_7[1]),.din(w_n642_2[0]));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(n654));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl3 jspl3_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.doutc(w_dff_A_7ujfS0FO3_2),.din(n672));
	jspl jspl_w_n672_1(.douta(w_n672_1[0]),.doutb(w_dff_A_z8l9MxUk1_1),.din(w_n672_0[0]));
	jspl3 jspl3_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.doutc(w_n675_0[2]),.din(n675));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(w_dff_B_WhCIUObC5_2));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_dff_A_bc0Bi0ZA8_1),.din(w_dff_B_X3IijG2u6_2));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_dff_A_aeOguVQ19_1),.doutc(w_n696_0[2]),.din(n696));
	jspl3 jspl3_w_n696_1(.douta(w_dff_A_TGkm35os1_0),.doutb(w_n696_1[1]),.doutc(w_dff_A_Z5GVPtXq1_2),.din(w_n696_0[0]));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.doutc(w_n743_0[2]),.din(n743));
	jspl jspl_w_n743_1(.douta(w_n743_1[0]),.doutb(w_n743_1[1]),.din(w_n743_0[0]));
	jspl jspl_w_n750_0(.douta(w_dff_A_nU0xe2hO8_0),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n754_0(.douta(w_dff_A_um81YCu52_0),.doutb(w_n754_0[1]),.din(n754));
	jspl3 jspl3_w_n758_0(.douta(w_dff_A_eiKxvlwp6_0),.doutb(w_dff_A_FYu6yqkl2_1),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n758_1(.douta(w_n758_1[0]),.doutb(w_dff_A_hXcPV68U0_1),.din(w_n758_0[0]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_dff_A_fk5jWGnA9_0),.doutb(w_n760_0[1]),.din(n760));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_dff_A_znYIGwJu5_2),.din(n764));
	jspl3 jspl3_w_n764_1(.douta(w_n764_1[0]),.doutb(w_n764_1[1]),.doutc(w_dff_A_S7H7Geem3_2),.din(w_n764_0[0]));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_n771_0[2]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_dff_A_JrPOuNJj8_0),.doutb(w_n779_0[1]),.din(n779));
	jspl jspl_w_n797_0(.douta(w_dff_A_i3FCZTXW0_0),.doutb(w_n797_0[1]),.din(n797));
	jspl jspl_w_n801_0(.douta(w_dff_A_ETicKf2s9_0),.doutb(w_n801_0[1]),.din(n801));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl3 jspl3_w_n853_0(.douta(w_n853_0[0]),.doutb(w_n853_0[1]),.doutc(w_n853_0[2]),.din(n853));
	jspl3 jspl3_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.doutc(w_n855_0[2]),.din(n855));
	jspl3 jspl3_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.doutc(w_dff_A_eTrHz4jv8_2),.din(n861));
	jspl jspl_w_n861_1(.douta(w_n861_1[0]),.doutb(w_dff_A_yC7bLEO03_1),.din(w_n861_0[0]));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.din(n863));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_dff_A_HHcohrtA2_1),.din(n899));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl3 jspl3_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.doutc(w_n937_0[2]),.din(n937));
	jspl jspl_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.din(n940));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_dff_A_ESKtCnJ84_1),.din(n962));
	jspl3 jspl3_w_n988_0(.douta(w_dff_A_qKqgdtiq5_0),.doutb(w_dff_A_Z6o3NE1T2_1),.doutc(w_n988_0[2]),.din(n988));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_dff_A_5CpDEeKf6_1),.din(n990));
	jspl3 jspl3_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.doutc(w_n991_0[2]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_dff_A_O8ofyVi79_1),.din(n999));
	jspl3 jspl3_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.doutc(w_n1001_0[2]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.doutc(w_n1002_0[2]),.din(n1002));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl3 jspl3_w_n1049_0(.douta(w_dff_A_VyKc0K8E5_0),.doutb(w_dff_A_d0PiL9Ll8_1),.doutc(w_n1049_0[2]),.din(n1049));
	jspl jspl_w_n1052_0(.douta(w_dff_A_0jptbRSB0_0),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_dff_A_gu9V6RPw5_1),.din(n1057));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(n1059));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl3 jspl3_w_n1162_0(.douta(w_n1162_0[0]),.doutb(w_dff_A_h6FWygUN2_1),.doutc(w_n1162_0[2]),.din(n1162));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(n1164));
	jspl jspl_w_n1172_0(.douta(w_dff_A_RuAtsRXB7_0),.doutb(w_n1172_0[1]),.din(n1172));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_dff_A_2l8Hn0jK5_1),.din(n1175));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_dff_A_DxjuNRJs4_1),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_dff_A_TiAQk5Re1_0),.doutb(w_n1184_0[1]),.din(n1184));
	jspl jspl_w_n1187_0(.douta(w_dff_A_r9l106aC1_0),.doutb(w_n1187_0[1]),.din(n1187));
	jdff dff_B_8aZMsUSg1_1(.din(n111),.dout(w_dff_B_8aZMsUSg1_1),.clk(gclk));
	jdff dff_B_nTRQHFet8_0(.din(n126),.dout(w_dff_B_nTRQHFet8_0),.clk(gclk));
	jdff dff_B_FHdOARZ04_0(.din(n125),.dout(w_dff_B_FHdOARZ04_0),.clk(gclk));
	jdff dff_A_MDs6Vcnr7_1(.dout(w_n72_1[1]),.din(w_dff_A_MDs6Vcnr7_1),.clk(gclk));
	jdff dff_A_Cy55RF5Q7_1(.dout(w_dff_A_MDs6Vcnr7_1),.din(w_dff_A_Cy55RF5Q7_1),.clk(gclk));
	jdff dff_A_Fnp8WRIn0_0(.dout(w_n98_2[0]),.din(w_dff_A_Fnp8WRIn0_0),.clk(gclk));
	jdff dff_B_ldRFVe202_1(.din(n540),.dout(w_dff_B_ldRFVe202_1),.clk(gclk));
	jdff dff_B_j6waDMC76_0(.din(n597),.dout(w_dff_B_j6waDMC76_0),.clk(gclk));
	jdff dff_B_3gI0awUS0_0(.din(w_dff_B_j6waDMC76_0),.dout(w_dff_B_3gI0awUS0_0),.clk(gclk));
	jdff dff_B_njzexcSK1_0(.din(w_dff_B_3gI0awUS0_0),.dout(w_dff_B_njzexcSK1_0),.clk(gclk));
	jdff dff_B_t4i66qn88_0(.din(w_dff_B_njzexcSK1_0),.dout(w_dff_B_t4i66qn88_0),.clk(gclk));
	jdff dff_B_kVySOI6Y1_0(.din(w_dff_B_t4i66qn88_0),.dout(w_dff_B_kVySOI6Y1_0),.clk(gclk));
	jdff dff_B_rDlpP4Tm2_0(.din(w_dff_B_kVySOI6Y1_0),.dout(w_dff_B_rDlpP4Tm2_0),.clk(gclk));
	jdff dff_B_7lYQBcTU9_0(.din(w_dff_B_rDlpP4Tm2_0),.dout(w_dff_B_7lYQBcTU9_0),.clk(gclk));
	jdff dff_B_k6hK0ZL41_0(.din(w_dff_B_7lYQBcTU9_0),.dout(w_dff_B_k6hK0ZL41_0),.clk(gclk));
	jdff dff_B_MJ4Ko4900_0(.din(w_dff_B_k6hK0ZL41_0),.dout(w_dff_B_MJ4Ko4900_0),.clk(gclk));
	jdff dff_B_FFN7T7lW1_0(.din(w_dff_B_MJ4Ko4900_0),.dout(w_dff_B_FFN7T7lW1_0),.clk(gclk));
	jdff dff_B_Meiy2dWM6_0(.din(n596),.dout(w_dff_B_Meiy2dWM6_0),.clk(gclk));
	jdff dff_B_jmc7yEn00_0(.din(n795),.dout(w_dff_B_jmc7yEn00_0),.clk(gclk));
	jdff dff_B_FBAA0OiE4_0(.din(w_dff_B_jmc7yEn00_0),.dout(w_dff_B_FBAA0OiE4_0),.clk(gclk));
	jdff dff_B_qg1WDuVP3_0(.din(w_dff_B_FBAA0OiE4_0),.dout(w_dff_B_qg1WDuVP3_0),.clk(gclk));
	jdff dff_B_ll4EBX4T5_0(.din(w_dff_B_qg1WDuVP3_0),.dout(w_dff_B_ll4EBX4T5_0),.clk(gclk));
	jdff dff_B_rOe93E8Z0_0(.din(w_dff_B_ll4EBX4T5_0),.dout(w_dff_B_rOe93E8Z0_0),.clk(gclk));
	jdff dff_B_MIeghigj1_0(.din(w_dff_B_rOe93E8Z0_0),.dout(w_dff_B_MIeghigj1_0),.clk(gclk));
	jdff dff_B_toQfQAC32_0(.din(w_dff_B_MIeghigj1_0),.dout(w_dff_B_toQfQAC32_0),.clk(gclk));
	jdff dff_B_ZElfSDKJ4_0(.din(w_dff_B_toQfQAC32_0),.dout(w_dff_B_ZElfSDKJ4_0),.clk(gclk));
	jdff dff_B_gfFi0Bru6_0(.din(w_dff_B_ZElfSDKJ4_0),.dout(w_dff_B_gfFi0Bru6_0),.clk(gclk));
	jdff dff_B_rWmrLOuI8_0(.din(w_dff_B_gfFi0Bru6_0),.dout(w_dff_B_rWmrLOuI8_0),.clk(gclk));
	jdff dff_B_xcToyw074_0(.din(w_dff_B_rWmrLOuI8_0),.dout(w_dff_B_xcToyw074_0),.clk(gclk));
	jdff dff_B_oXeKlS7g6_0(.din(w_dff_B_xcToyw074_0),.dout(w_dff_B_oXeKlS7g6_0),.clk(gclk));
	jdff dff_B_SVhmJNuT3_0(.din(w_dff_B_oXeKlS7g6_0),.dout(w_dff_B_SVhmJNuT3_0),.clk(gclk));
	jdff dff_B_UazcTnMj9_0(.din(w_dff_B_SVhmJNuT3_0),.dout(w_dff_B_UazcTnMj9_0),.clk(gclk));
	jdff dff_B_fMbyyNtm4_0(.din(w_dff_B_UazcTnMj9_0),.dout(w_dff_B_fMbyyNtm4_0),.clk(gclk));
	jdff dff_B_9HLj2MZf8_0(.din(w_dff_B_fMbyyNtm4_0),.dout(w_dff_B_9HLj2MZf8_0),.clk(gclk));
	jdff dff_B_a03BJKRD2_0(.din(w_dff_B_9HLj2MZf8_0),.dout(w_dff_B_a03BJKRD2_0),.clk(gclk));
	jdff dff_B_h20AqAp38_1(.din(n791),.dout(w_dff_B_h20AqAp38_1),.clk(gclk));
	jdff dff_B_KGWBjATJ3_0(.din(n793),.dout(w_dff_B_KGWBjATJ3_0),.clk(gclk));
	jdff dff_B_8dhPwf6t8_0(.din(w_dff_B_KGWBjATJ3_0),.dout(w_dff_B_8dhPwf6t8_0),.clk(gclk));
	jdff dff_B_A73Inxk12_0(.din(n784),.dout(w_dff_B_A73Inxk12_0),.clk(gclk));
	jdff dff_B_iUQfLqnQ3_0(.din(w_dff_B_A73Inxk12_0),.dout(w_dff_B_iUQfLqnQ3_0),.clk(gclk));
	jdff dff_B_qUNMdAgl3_0(.din(w_dff_B_iUQfLqnQ3_0),.dout(w_dff_B_qUNMdAgl3_0),.clk(gclk));
	jdff dff_B_5xQQZF0D0_0(.din(w_dff_B_qUNMdAgl3_0),.dout(w_dff_B_5xQQZF0D0_0),.clk(gclk));
	jdff dff_B_GKzjQE1R3_0(.din(w_dff_B_5xQQZF0D0_0),.dout(w_dff_B_GKzjQE1R3_0),.clk(gclk));
	jdff dff_B_WJA4ZsAw5_0(.din(w_dff_B_GKzjQE1R3_0),.dout(w_dff_B_WJA4ZsAw5_0),.clk(gclk));
	jdff dff_B_sYnYWvBN0_0(.din(w_dff_B_WJA4ZsAw5_0),.dout(w_dff_B_sYnYWvBN0_0),.clk(gclk));
	jdff dff_B_BIXpI8E30_0(.din(w_dff_B_sYnYWvBN0_0),.dout(w_dff_B_BIXpI8E30_0),.clk(gclk));
	jdff dff_B_az5NFJ6w8_0(.din(w_dff_B_BIXpI8E30_0),.dout(w_dff_B_az5NFJ6w8_0),.clk(gclk));
	jdff dff_B_xrkJsPzh4_0(.din(w_dff_B_az5NFJ6w8_0),.dout(w_dff_B_xrkJsPzh4_0),.clk(gclk));
	jdff dff_B_VBqfAsvq8_0(.din(w_dff_B_xrkJsPzh4_0),.dout(w_dff_B_VBqfAsvq8_0),.clk(gclk));
	jdff dff_B_GgxeHxsu5_0(.din(w_dff_B_VBqfAsvq8_0),.dout(w_dff_B_GgxeHxsu5_0),.clk(gclk));
	jdff dff_B_01o3erlq4_0(.din(w_dff_B_GgxeHxsu5_0),.dout(w_dff_B_01o3erlq4_0),.clk(gclk));
	jdff dff_B_kWKl3YgX2_0(.din(w_dff_B_01o3erlq4_0),.dout(w_dff_B_kWKl3YgX2_0),.clk(gclk));
	jdff dff_B_uToLvsbu0_0(.din(w_dff_B_kWKl3YgX2_0),.dout(w_dff_B_uToLvsbu0_0),.clk(gclk));
	jdff dff_B_DrwagBmw7_0(.din(w_dff_B_uToLvsbu0_0),.dout(w_dff_B_DrwagBmw7_0),.clk(gclk));
	jdff dff_B_08UZhAAQ1_0(.din(w_dff_B_DrwagBmw7_0),.dout(w_dff_B_08UZhAAQ1_0),.clk(gclk));
	jdff dff_A_kWsQxzyD4_1(.dout(w_n116_0[1]),.din(w_dff_A_kWsQxzyD4_1),.clk(gclk));
	jdff dff_A_XPpM07ww0_1(.dout(w_dff_A_kWsQxzyD4_1),.din(w_dff_A_XPpM07ww0_1),.clk(gclk));
	jdff dff_B_1ebv9Ywc6_0(.din(n780),.dout(w_dff_B_1ebv9Ywc6_0),.clk(gclk));
	jdff dff_A_JrPOuNJj8_0(.dout(w_n779_0[0]),.din(w_dff_A_JrPOuNJj8_0),.clk(gclk));
	jdff dff_B_C6myuNG13_1(.din(n774),.dout(w_dff_B_C6myuNG13_1),.clk(gclk));
	jdff dff_A_l8FyxM895_0(.dout(w_n519_1[0]),.din(w_dff_A_l8FyxM895_0),.clk(gclk));
	jdff dff_B_YxMyLRdw2_1(.din(n1174),.dout(w_dff_B_YxMyLRdw2_1),.clk(gclk));
	jdff dff_B_IhQIpIaA0_1(.din(w_dff_B_YxMyLRdw2_1),.dout(w_dff_B_IhQIpIaA0_1),.clk(gclk));
	jdff dff_B_B6DW9lbj3_1(.din(w_dff_B_IhQIpIaA0_1),.dout(w_dff_B_B6DW9lbj3_1),.clk(gclk));
	jdff dff_B_gtIhX11Z3_1(.din(w_dff_B_B6DW9lbj3_1),.dout(w_dff_B_gtIhX11Z3_1),.clk(gclk));
	jdff dff_B_96h1m6QL5_1(.din(w_dff_B_gtIhX11Z3_1),.dout(w_dff_B_96h1m6QL5_1),.clk(gclk));
	jdff dff_B_G272gM9Z8_1(.din(w_dff_B_96h1m6QL5_1),.dout(w_dff_B_G272gM9Z8_1),.clk(gclk));
	jdff dff_B_ykvTJ1bc3_1(.din(w_dff_B_G272gM9Z8_1),.dout(w_dff_B_ykvTJ1bc3_1),.clk(gclk));
	jdff dff_B_mM3jbKiG4_1(.din(w_dff_B_ykvTJ1bc3_1),.dout(w_dff_B_mM3jbKiG4_1),.clk(gclk));
	jdff dff_B_RO0M0pTf6_1(.din(w_dff_B_mM3jbKiG4_1),.dout(w_dff_B_RO0M0pTf6_1),.clk(gclk));
	jdff dff_B_TEkBKpVL7_1(.din(w_dff_B_RO0M0pTf6_1),.dout(w_dff_B_TEkBKpVL7_1),.clk(gclk));
	jdff dff_B_XpZeYqJT5_1(.din(w_dff_B_TEkBKpVL7_1),.dout(w_dff_B_XpZeYqJT5_1),.clk(gclk));
	jdff dff_B_yP207U600_1(.din(w_dff_B_XpZeYqJT5_1),.dout(w_dff_B_yP207U600_1),.clk(gclk));
	jdff dff_B_x4m8ajeN6_1(.din(w_dff_B_yP207U600_1),.dout(w_dff_B_x4m8ajeN6_1),.clk(gclk));
	jdff dff_B_5bux0arX6_1(.din(w_dff_B_x4m8ajeN6_1),.dout(w_dff_B_5bux0arX6_1),.clk(gclk));
	jdff dff_B_1mEcKKrc8_1(.din(w_dff_B_5bux0arX6_1),.dout(w_dff_B_1mEcKKrc8_1),.clk(gclk));
	jdff dff_B_k3KVRscA8_1(.din(w_dff_B_1mEcKKrc8_1),.dout(w_dff_B_k3KVRscA8_1),.clk(gclk));
	jdff dff_B_Bq0kVR0O9_1(.din(w_dff_B_k3KVRscA8_1),.dout(w_dff_B_Bq0kVR0O9_1),.clk(gclk));
	jdff dff_B_aYZVBZi78_1(.din(w_dff_B_Bq0kVR0O9_1),.dout(w_dff_B_aYZVBZi78_1),.clk(gclk));
	jdff dff_B_ZqXARUce0_1(.din(w_dff_B_aYZVBZi78_1),.dout(w_dff_B_ZqXARUce0_1),.clk(gclk));
	jdff dff_B_xILg8HgC6_1(.din(w_dff_B_ZqXARUce0_1),.dout(w_dff_B_xILg8HgC6_1),.clk(gclk));
	jdff dff_B_aLbDCmTi0_1(.din(w_dff_B_xILg8HgC6_1),.dout(w_dff_B_aLbDCmTi0_1),.clk(gclk));
	jdff dff_B_wXcETJsI9_1(.din(w_dff_B_aLbDCmTi0_1),.dout(w_dff_B_wXcETJsI9_1),.clk(gclk));
	jdff dff_B_TJxq1Y5N5_1(.din(w_dff_B_wXcETJsI9_1),.dout(w_dff_B_TJxq1Y5N5_1),.clk(gclk));
	jdff dff_B_OvWgd3B04_1(.din(w_dff_B_TJxq1Y5N5_1),.dout(w_dff_B_OvWgd3B04_1),.clk(gclk));
	jdff dff_B_Ifi2zEUX1_1(.din(w_dff_B_OvWgd3B04_1),.dout(w_dff_B_Ifi2zEUX1_1),.clk(gclk));
	jdff dff_B_70Lh1d4I4_1(.din(w_dff_B_Ifi2zEUX1_1),.dout(w_dff_B_70Lh1d4I4_1),.clk(gclk));
	jdff dff_A_RuAtsRXB7_0(.dout(w_n1172_0[0]),.din(w_dff_A_RuAtsRXB7_0),.clk(gclk));
	jdff dff_B_BIcvvNtC5_1(.din(n1166),.dout(w_dff_B_BIcvvNtC5_1),.clk(gclk));
	jdff dff_B_0z1zdyUY5_1(.din(w_dff_B_BIcvvNtC5_1),.dout(w_dff_B_0z1zdyUY5_1),.clk(gclk));
	jdff dff_B_pDDrbT6h3_1(.din(n1186),.dout(w_dff_B_pDDrbT6h3_1),.clk(gclk));
	jdff dff_B_Nua3Uscy5_1(.din(w_dff_B_pDDrbT6h3_1),.dout(w_dff_B_Nua3Uscy5_1),.clk(gclk));
	jdff dff_B_8ucCZc955_1(.din(w_dff_B_Nua3Uscy5_1),.dout(w_dff_B_8ucCZc955_1),.clk(gclk));
	jdff dff_B_vOUZ7sJR2_1(.din(w_dff_B_8ucCZc955_1),.dout(w_dff_B_vOUZ7sJR2_1),.clk(gclk));
	jdff dff_B_OryVXVYG8_1(.din(w_dff_B_vOUZ7sJR2_1),.dout(w_dff_B_OryVXVYG8_1),.clk(gclk));
	jdff dff_B_L4z9TSUs1_1(.din(w_dff_B_OryVXVYG8_1),.dout(w_dff_B_L4z9TSUs1_1),.clk(gclk));
	jdff dff_B_v3N1Brr01_1(.din(w_dff_B_L4z9TSUs1_1),.dout(w_dff_B_v3N1Brr01_1),.clk(gclk));
	jdff dff_B_U8Syk4L07_1(.din(w_dff_B_v3N1Brr01_1),.dout(w_dff_B_U8Syk4L07_1),.clk(gclk));
	jdff dff_B_qiEjx3fb9_1(.din(w_dff_B_U8Syk4L07_1),.dout(w_dff_B_qiEjx3fb9_1),.clk(gclk));
	jdff dff_B_ugKgAaRj7_1(.din(w_dff_B_qiEjx3fb9_1),.dout(w_dff_B_ugKgAaRj7_1),.clk(gclk));
	jdff dff_B_bsYBlFQC6_1(.din(w_dff_B_ugKgAaRj7_1),.dout(w_dff_B_bsYBlFQC6_1),.clk(gclk));
	jdff dff_B_r0Zni9ip3_1(.din(w_dff_B_bsYBlFQC6_1),.dout(w_dff_B_r0Zni9ip3_1),.clk(gclk));
	jdff dff_B_PHIVRap49_1(.din(w_dff_B_r0Zni9ip3_1),.dout(w_dff_B_PHIVRap49_1),.clk(gclk));
	jdff dff_B_3BXgcVFQ4_1(.din(w_dff_B_PHIVRap49_1),.dout(w_dff_B_3BXgcVFQ4_1),.clk(gclk));
	jdff dff_B_8kFOkYio2_1(.din(w_dff_B_3BXgcVFQ4_1),.dout(w_dff_B_8kFOkYio2_1),.clk(gclk));
	jdff dff_B_HbyLvWG12_1(.din(w_dff_B_8kFOkYio2_1),.dout(w_dff_B_HbyLvWG12_1),.clk(gclk));
	jdff dff_B_9xpwargc1_1(.din(w_dff_B_HbyLvWG12_1),.dout(w_dff_B_9xpwargc1_1),.clk(gclk));
	jdff dff_B_zEbeDmnE8_1(.din(w_dff_B_9xpwargc1_1),.dout(w_dff_B_zEbeDmnE8_1),.clk(gclk));
	jdff dff_B_AbOrrKBs0_1(.din(w_dff_B_zEbeDmnE8_1),.dout(w_dff_B_AbOrrKBs0_1),.clk(gclk));
	jdff dff_B_3gnqDvH62_1(.din(w_dff_B_AbOrrKBs0_1),.dout(w_dff_B_3gnqDvH62_1),.clk(gclk));
	jdff dff_B_1Frq4AFi1_1(.din(w_dff_B_3gnqDvH62_1),.dout(w_dff_B_1Frq4AFi1_1),.clk(gclk));
	jdff dff_B_r6us2hmd6_1(.din(w_dff_B_1Frq4AFi1_1),.dout(w_dff_B_r6us2hmd6_1),.clk(gclk));
	jdff dff_B_kXptMM8s9_1(.din(w_dff_B_r6us2hmd6_1),.dout(w_dff_B_kXptMM8s9_1),.clk(gclk));
	jdff dff_B_ymAn6tCn5_1(.din(G2897),.dout(w_dff_B_ymAn6tCn5_1),.clk(gclk));
	jdff dff_B_sJSKpJ2F1_1(.din(w_dff_B_ymAn6tCn5_1),.dout(w_dff_B_sJSKpJ2F1_1),.clk(gclk));
	jdff dff_B_QHOGV6Yf9_1(.din(w_dff_B_sJSKpJ2F1_1),.dout(w_dff_B_QHOGV6Yf9_1),.clk(gclk));
	jdff dff_A_mHZxPKWf3_0(.dout(w_n1184_0[0]),.din(w_dff_A_mHZxPKWf3_0),.clk(gclk));
	jdff dff_A_VH2U8Oq64_0(.dout(w_dff_A_mHZxPKWf3_0),.din(w_dff_A_VH2U8Oq64_0),.clk(gclk));
	jdff dff_A_XBIBSthK4_0(.dout(w_dff_A_VH2U8Oq64_0),.din(w_dff_A_XBIBSthK4_0),.clk(gclk));
	jdff dff_A_poTCiQoY4_0(.dout(w_dff_A_XBIBSthK4_0),.din(w_dff_A_poTCiQoY4_0),.clk(gclk));
	jdff dff_A_wAbsF8o51_0(.dout(w_dff_A_poTCiQoY4_0),.din(w_dff_A_wAbsF8o51_0),.clk(gclk));
	jdff dff_A_geEesXKv6_0(.dout(w_dff_A_wAbsF8o51_0),.din(w_dff_A_geEesXKv6_0),.clk(gclk));
	jdff dff_A_Tmwd6mbF1_0(.dout(w_dff_A_geEesXKv6_0),.din(w_dff_A_Tmwd6mbF1_0),.clk(gclk));
	jdff dff_A_vwSIPiSD5_0(.dout(w_dff_A_Tmwd6mbF1_0),.din(w_dff_A_vwSIPiSD5_0),.clk(gclk));
	jdff dff_A_wVgi0O2n8_0(.dout(w_dff_A_vwSIPiSD5_0),.din(w_dff_A_wVgi0O2n8_0),.clk(gclk));
	jdff dff_A_UUiwvjWN7_0(.dout(w_dff_A_wVgi0O2n8_0),.din(w_dff_A_UUiwvjWN7_0),.clk(gclk));
	jdff dff_A_0ep7acPz3_0(.dout(w_dff_A_UUiwvjWN7_0),.din(w_dff_A_0ep7acPz3_0),.clk(gclk));
	jdff dff_A_TBpBjb3h4_0(.dout(w_dff_A_0ep7acPz3_0),.din(w_dff_A_TBpBjb3h4_0),.clk(gclk));
	jdff dff_A_Zko62mKg4_0(.dout(w_dff_A_TBpBjb3h4_0),.din(w_dff_A_Zko62mKg4_0),.clk(gclk));
	jdff dff_A_5rFFZyZ71_0(.dout(w_dff_A_Zko62mKg4_0),.din(w_dff_A_5rFFZyZ71_0),.clk(gclk));
	jdff dff_A_6oNImClC8_0(.dout(w_dff_A_5rFFZyZ71_0),.din(w_dff_A_6oNImClC8_0),.clk(gclk));
	jdff dff_A_NXl4ivyk3_0(.dout(w_dff_A_6oNImClC8_0),.din(w_dff_A_NXl4ivyk3_0),.clk(gclk));
	jdff dff_A_YobG7PX29_0(.dout(w_dff_A_NXl4ivyk3_0),.din(w_dff_A_YobG7PX29_0),.clk(gclk));
	jdff dff_A_7i5c9rVa5_0(.dout(w_dff_A_YobG7PX29_0),.din(w_dff_A_7i5c9rVa5_0),.clk(gclk));
	jdff dff_A_yHeClDfL7_0(.dout(w_dff_A_7i5c9rVa5_0),.din(w_dff_A_yHeClDfL7_0),.clk(gclk));
	jdff dff_A_o4Y9rtJm4_0(.dout(w_dff_A_yHeClDfL7_0),.din(w_dff_A_o4Y9rtJm4_0),.clk(gclk));
	jdff dff_A_YCjAZHWK0_0(.dout(w_dff_A_o4Y9rtJm4_0),.din(w_dff_A_YCjAZHWK0_0),.clk(gclk));
	jdff dff_A_LdsCSEZI6_0(.dout(w_dff_A_YCjAZHWK0_0),.din(w_dff_A_LdsCSEZI6_0),.clk(gclk));
	jdff dff_A_ChRngGDO9_0(.dout(w_dff_A_LdsCSEZI6_0),.din(w_dff_A_ChRngGDO9_0),.clk(gclk));
	jdff dff_A_TiAQk5Re1_0(.dout(w_dff_A_ChRngGDO9_0),.din(w_dff_A_TiAQk5Re1_0),.clk(gclk));
	jdff dff_A_zj7SLwyd6_1(.dout(w_n1175_0[1]),.din(w_dff_A_zj7SLwyd6_1),.clk(gclk));
	jdff dff_A_MlWFf3bL3_1(.dout(w_dff_A_zj7SLwyd6_1),.din(w_dff_A_MlWFf3bL3_1),.clk(gclk));
	jdff dff_A_GDrDJWA68_1(.dout(w_dff_A_MlWFf3bL3_1),.din(w_dff_A_GDrDJWA68_1),.clk(gclk));
	jdff dff_A_X7uxLpvT9_1(.dout(w_dff_A_GDrDJWA68_1),.din(w_dff_A_X7uxLpvT9_1),.clk(gclk));
	jdff dff_A_ZdNri9a43_1(.dout(w_dff_A_X7uxLpvT9_1),.din(w_dff_A_ZdNri9a43_1),.clk(gclk));
	jdff dff_A_H3PqiOfo1_1(.dout(w_dff_A_ZdNri9a43_1),.din(w_dff_A_H3PqiOfo1_1),.clk(gclk));
	jdff dff_A_Jie2WfFc5_1(.dout(w_dff_A_H3PqiOfo1_1),.din(w_dff_A_Jie2WfFc5_1),.clk(gclk));
	jdff dff_A_kUwnmmrZ7_1(.dout(w_dff_A_Jie2WfFc5_1),.din(w_dff_A_kUwnmmrZ7_1),.clk(gclk));
	jdff dff_A_FETIMacw5_1(.dout(w_dff_A_kUwnmmrZ7_1),.din(w_dff_A_FETIMacw5_1),.clk(gclk));
	jdff dff_A_WQ1bN8qa7_1(.dout(w_dff_A_FETIMacw5_1),.din(w_dff_A_WQ1bN8qa7_1),.clk(gclk));
	jdff dff_A_otMMfgfO8_1(.dout(w_dff_A_WQ1bN8qa7_1),.din(w_dff_A_otMMfgfO8_1),.clk(gclk));
	jdff dff_A_3EpVKPhz5_1(.dout(w_dff_A_otMMfgfO8_1),.din(w_dff_A_3EpVKPhz5_1),.clk(gclk));
	jdff dff_A_cMoJ2o695_1(.dout(w_dff_A_3EpVKPhz5_1),.din(w_dff_A_cMoJ2o695_1),.clk(gclk));
	jdff dff_A_AzeBjmfW0_1(.dout(w_dff_A_cMoJ2o695_1),.din(w_dff_A_AzeBjmfW0_1),.clk(gclk));
	jdff dff_A_0USWjrUG2_1(.dout(w_dff_A_AzeBjmfW0_1),.din(w_dff_A_0USWjrUG2_1),.clk(gclk));
	jdff dff_A_oZZG3HHc4_1(.dout(w_dff_A_0USWjrUG2_1),.din(w_dff_A_oZZG3HHc4_1),.clk(gclk));
	jdff dff_A_WWeEPOPW1_1(.dout(w_dff_A_oZZG3HHc4_1),.din(w_dff_A_WWeEPOPW1_1),.clk(gclk));
	jdff dff_A_3uhekAjo8_1(.dout(w_dff_A_WWeEPOPW1_1),.din(w_dff_A_3uhekAjo8_1),.clk(gclk));
	jdff dff_A_0tZXxpk23_1(.dout(w_dff_A_3uhekAjo8_1),.din(w_dff_A_0tZXxpk23_1),.clk(gclk));
	jdff dff_A_tugRnaRv1_1(.dout(w_dff_A_0tZXxpk23_1),.din(w_dff_A_tugRnaRv1_1),.clk(gclk));
	jdff dff_A_oPtuWTSr1_1(.dout(w_dff_A_tugRnaRv1_1),.din(w_dff_A_oPtuWTSr1_1),.clk(gclk));
	jdff dff_A_VRBojeX93_1(.dout(w_dff_A_oPtuWTSr1_1),.din(w_dff_A_VRBojeX93_1),.clk(gclk));
	jdff dff_A_B6w6EnVH3_1(.dout(w_dff_A_VRBojeX93_1),.din(w_dff_A_B6w6EnVH3_1),.clk(gclk));
	jdff dff_A_yM4DEeYD2_1(.dout(w_dff_A_B6w6EnVH3_1),.din(w_dff_A_yM4DEeYD2_1),.clk(gclk));
	jdff dff_A_2l8Hn0jK5_1(.dout(w_dff_A_yM4DEeYD2_1),.din(w_dff_A_2l8Hn0jK5_1),.clk(gclk));
	jdff dff_A_r9l106aC1_0(.dout(w_n1187_0[0]),.din(w_dff_A_r9l106aC1_0),.clk(gclk));
	jdff dff_B_HbZ2tRBn8_1(.din(n1060),.dout(w_dff_B_HbZ2tRBn8_1),.clk(gclk));
	jdff dff_B_GJyJzrYg5_0(.din(n1112),.dout(w_dff_B_GJyJzrYg5_0),.clk(gclk));
	jdff dff_B_m6mt5lgo3_0(.din(w_dff_B_GJyJzrYg5_0),.dout(w_dff_B_m6mt5lgo3_0),.clk(gclk));
	jdff dff_B_FnDaVBy43_0(.din(w_dff_B_m6mt5lgo3_0),.dout(w_dff_B_FnDaVBy43_0),.clk(gclk));
	jdff dff_B_nWFepMSS1_0(.din(w_dff_B_FnDaVBy43_0),.dout(w_dff_B_nWFepMSS1_0),.clk(gclk));
	jdff dff_B_ApGIYt5O2_0(.din(w_dff_B_nWFepMSS1_0),.dout(w_dff_B_ApGIYt5O2_0),.clk(gclk));
	jdff dff_B_M5crVnnZ1_0(.din(w_dff_B_ApGIYt5O2_0),.dout(w_dff_B_M5crVnnZ1_0),.clk(gclk));
	jdff dff_B_2ZzevI7Z5_0(.din(n1111),.dout(w_dff_B_2ZzevI7Z5_0),.clk(gclk));
	jdff dff_B_6RlGO1el5_0(.din(w_dff_B_2ZzevI7Z5_0),.dout(w_dff_B_6RlGO1el5_0),.clk(gclk));
	jdff dff_B_g6NpZbtg4_0(.din(n1110),.dout(w_dff_B_g6NpZbtg4_0),.clk(gclk));
	jdff dff_B_9LYSI1eH6_0(.din(w_dff_B_g6NpZbtg4_0),.dout(w_dff_B_9LYSI1eH6_0),.clk(gclk));
	jdff dff_B_zfiVbqXR4_0(.din(w_dff_B_9LYSI1eH6_0),.dout(w_dff_B_zfiVbqXR4_0),.clk(gclk));
	jdff dff_B_jkxPcBk06_0(.din(w_dff_B_zfiVbqXR4_0),.dout(w_dff_B_jkxPcBk06_0),.clk(gclk));
	jdff dff_B_R0XxsxpC1_0(.din(w_dff_B_jkxPcBk06_0),.dout(w_dff_B_R0XxsxpC1_0),.clk(gclk));
	jdff dff_B_VX0yxNuR9_0(.din(n1109),.dout(w_dff_B_VX0yxNuR9_0),.clk(gclk));
	jdff dff_B_eWTdcCEz0_0(.din(w_dff_B_VX0yxNuR9_0),.dout(w_dff_B_eWTdcCEz0_0),.clk(gclk));
	jdff dff_B_8XoYZ3G05_1(.din(n1066),.dout(w_dff_B_8XoYZ3G05_1),.clk(gclk));
	jdff dff_B_Z3t2a2eE8_1(.din(w_dff_B_8XoYZ3G05_1),.dout(w_dff_B_Z3t2a2eE8_1),.clk(gclk));
	jdff dff_B_6Zgzeqpj6_1(.din(w_dff_B_Z3t2a2eE8_1),.dout(w_dff_B_6Zgzeqpj6_1),.clk(gclk));
	jdff dff_B_GjLlNvMz7_1(.din(w_dff_B_6Zgzeqpj6_1),.dout(w_dff_B_GjLlNvMz7_1),.clk(gclk));
	jdff dff_B_h1ZxgAE56_1(.din(w_dff_B_GjLlNvMz7_1),.dout(w_dff_B_h1ZxgAE56_1),.clk(gclk));
	jdff dff_B_1i38jL5G9_1(.din(w_dff_B_h1ZxgAE56_1),.dout(w_dff_B_1i38jL5G9_1),.clk(gclk));
	jdff dff_B_pEMQrzCV0_1(.din(w_dff_B_1i38jL5G9_1),.dout(w_dff_B_pEMQrzCV0_1),.clk(gclk));
	jdff dff_B_Dc1teHUy7_1(.din(w_dff_B_pEMQrzCV0_1),.dout(w_dff_B_Dc1teHUy7_1),.clk(gclk));
	jdff dff_B_ms8W2Lke6_1(.din(n1086),.dout(w_dff_B_ms8W2Lke6_1),.clk(gclk));
	jdff dff_B_IOZhVMyW2_0(.din(n1105),.dout(w_dff_B_IOZhVMyW2_0),.clk(gclk));
	jdff dff_B_MVmd3Uho4_0(.din(w_dff_B_IOZhVMyW2_0),.dout(w_dff_B_MVmd3Uho4_0),.clk(gclk));
	jdff dff_B_9w95WRaS0_0(.din(w_dff_B_MVmd3Uho4_0),.dout(w_dff_B_9w95WRaS0_0),.clk(gclk));
	jdff dff_B_mxzQYyCT8_0(.din(w_dff_B_9w95WRaS0_0),.dout(w_dff_B_mxzQYyCT8_0),.clk(gclk));
	jdff dff_B_cqhd36od9_0(.din(w_dff_B_mxzQYyCT8_0),.dout(w_dff_B_cqhd36od9_0),.clk(gclk));
	jdff dff_B_y6Vqf3g16_0(.din(w_dff_B_cqhd36od9_0),.dout(w_dff_B_y6Vqf3g16_0),.clk(gclk));
	jdff dff_B_jTIuBr0a9_0(.din(w_dff_B_y6Vqf3g16_0),.dout(w_dff_B_jTIuBr0a9_0),.clk(gclk));
	jdff dff_B_Ie3G75Ik7_0(.din(w_dff_B_jTIuBr0a9_0),.dout(w_dff_B_Ie3G75Ik7_0),.clk(gclk));
	jdff dff_B_yfineotg2_1(.din(n1092),.dout(w_dff_B_yfineotg2_1),.clk(gclk));
	jdff dff_B_o3f2Divt9_1(.din(n1096),.dout(w_dff_B_o3f2Divt9_1),.clk(gclk));
	jdff dff_B_ZsBPbCzM7_1(.din(w_dff_B_o3f2Divt9_1),.dout(w_dff_B_ZsBPbCzM7_1),.clk(gclk));
	jdff dff_B_EHAmpLNC1_0(.din(n1099),.dout(w_dff_B_EHAmpLNC1_0),.clk(gclk));
	jdff dff_B_NNe1iWJ31_0(.din(n1095),.dout(w_dff_B_NNe1iWJ31_0),.clk(gclk));
	jdff dff_B_8nbF8iv83_0(.din(w_dff_B_NNe1iWJ31_0),.dout(w_dff_B_8nbF8iv83_0),.clk(gclk));
	jdff dff_B_0VEg4nU59_0(.din(w_dff_B_8nbF8iv83_0),.dout(w_dff_B_0VEg4nU59_0),.clk(gclk));
	jdff dff_B_401L7AbP2_1(.din(n1087),.dout(w_dff_B_401L7AbP2_1),.clk(gclk));
	jdff dff_B_Of5oisTA5_1(.din(w_dff_B_401L7AbP2_1),.dout(w_dff_B_Of5oisTA5_1),.clk(gclk));
	jdff dff_B_DyzEanKZ7_0(.din(n1089),.dout(w_dff_B_DyzEanKZ7_0),.clk(gclk));
	jdff dff_B_llo0HSNX3_1(.din(n1072),.dout(w_dff_B_llo0HSNX3_1),.clk(gclk));
	jdff dff_B_UbgWf2mq6_1(.din(w_dff_B_llo0HSNX3_1),.dout(w_dff_B_UbgWf2mq6_1),.clk(gclk));
	jdff dff_B_SYxa1nNY0_1(.din(n1076),.dout(w_dff_B_SYxa1nNY0_1),.clk(gclk));
	jdff dff_B_4Ks4C6Wa7_1(.din(G124),.dout(w_dff_B_4Ks4C6Wa7_1),.clk(gclk));
	jdff dff_B_rOBnvl9s1_1(.din(w_dff_B_4Ks4C6Wa7_1),.dout(w_dff_B_rOBnvl9s1_1),.clk(gclk));
	jdff dff_B_zOJ8wkxH1_1(.din(w_dff_B_rOBnvl9s1_1),.dout(w_dff_B_zOJ8wkxH1_1),.clk(gclk));
	jdff dff_B_erZgD98O7_1(.din(w_dff_B_zOJ8wkxH1_1),.dout(w_dff_B_erZgD98O7_1),.clk(gclk));
	jdff dff_B_BPeRjwXy5_1(.din(n1077),.dout(w_dff_B_BPeRjwXy5_1),.clk(gclk));
	jdff dff_B_nl3pMGxk3_0(.din(n1075),.dout(w_dff_B_nl3pMGxk3_0),.clk(gclk));
	jdff dff_B_xmWiSD9n9_0(.din(w_dff_B_nl3pMGxk3_0),.dout(w_dff_B_xmWiSD9n9_0),.clk(gclk));
	jdff dff_B_VUrcezlU8_0(.din(w_dff_B_xmWiSD9n9_0),.dout(w_dff_B_VUrcezlU8_0),.clk(gclk));
	jdff dff_B_poS95E5R3_0(.din(w_dff_B_VUrcezlU8_0),.dout(w_dff_B_poS95E5R3_0),.clk(gclk));
	jdff dff_B_cgxjWMuI9_1(.din(n1067),.dout(w_dff_B_cgxjWMuI9_1),.clk(gclk));
	jdff dff_B_ES2YB4tC6_1(.din(n1061),.dout(w_dff_B_ES2YB4tC6_1),.clk(gclk));
	jdff dff_B_BcRE7Wck8_1(.din(n1051),.dout(w_dff_B_BcRE7Wck8_1),.clk(gclk));
	jdff dff_B_ZPHCc3s71_1(.din(w_dff_B_BcRE7Wck8_1),.dout(w_dff_B_ZPHCc3s71_1),.clk(gclk));
	jdff dff_B_0Wh4mUwg8_1(.din(w_dff_B_ZPHCc3s71_1),.dout(w_dff_B_0Wh4mUwg8_1),.clk(gclk));
	jdff dff_A_t7KsM1fg9_1(.dout(w_n1057_0[1]),.din(w_dff_A_t7KsM1fg9_1),.clk(gclk));
	jdff dff_A_iyAYWHzH5_1(.dout(w_dff_A_t7KsM1fg9_1),.din(w_dff_A_iyAYWHzH5_1),.clk(gclk));
	jdff dff_A_jGO7FZbT7_1(.dout(w_dff_A_iyAYWHzH5_1),.din(w_dff_A_jGO7FZbT7_1),.clk(gclk));
	jdff dff_A_SlwfD1su5_1(.dout(w_dff_A_jGO7FZbT7_1),.din(w_dff_A_SlwfD1su5_1),.clk(gclk));
	jdff dff_A_gu9V6RPw5_1(.dout(w_dff_A_SlwfD1su5_1),.din(w_dff_A_gu9V6RPw5_1),.clk(gclk));
	jdff dff_A_0jptbRSB0_0(.dout(w_n1052_0[0]),.din(w_dff_A_0jptbRSB0_0),.clk(gclk));
	jdff dff_B_FalOaTVm9_1(.din(n753),.dout(w_dff_B_FalOaTVm9_1),.clk(gclk));
	jdff dff_B_LmEkCVDf8_1(.din(w_dff_B_FalOaTVm9_1),.dout(w_dff_B_LmEkCVDf8_1),.clk(gclk));
	jdff dff_B_MIstKFXz0_1(.din(w_dff_B_LmEkCVDf8_1),.dout(w_dff_B_MIstKFXz0_1),.clk(gclk));
	jdff dff_B_PpII1eyy4_1(.din(w_dff_B_MIstKFXz0_1),.dout(w_dff_B_PpII1eyy4_1),.clk(gclk));
	jdff dff_B_P9jroFVj2_1(.din(w_dff_B_PpII1eyy4_1),.dout(w_dff_B_P9jroFVj2_1),.clk(gclk));
	jdff dff_B_JsDsytI55_1(.din(w_dff_B_P9jroFVj2_1),.dout(w_dff_B_JsDsytI55_1),.clk(gclk));
	jdff dff_A_SJmOnuzi0_1(.dout(w_n758_1[1]),.din(w_dff_A_SJmOnuzi0_1),.clk(gclk));
	jdff dff_A_8L0DwhXT3_1(.dout(w_dff_A_SJmOnuzi0_1),.din(w_dff_A_8L0DwhXT3_1),.clk(gclk));
	jdff dff_A_hXcPV68U0_1(.dout(w_dff_A_8L0DwhXT3_1),.din(w_dff_A_hXcPV68U0_1),.clk(gclk));
	jdff dff_B_9BqoDOAJ9_0(.din(n752),.dout(w_dff_B_9BqoDOAJ9_0),.clk(gclk));
	jdff dff_B_0MIFE1Bw3_0(.din(w_dff_B_9BqoDOAJ9_0),.dout(w_dff_B_0MIFE1Bw3_0),.clk(gclk));
	jdff dff_B_nlp9xfky9_0(.din(w_dff_B_0MIFE1Bw3_0),.dout(w_dff_B_nlp9xfky9_0),.clk(gclk));
	jdff dff_B_s2xF01Tw8_0(.din(w_dff_B_nlp9xfky9_0),.dout(w_dff_B_s2xF01Tw8_0),.clk(gclk));
	jdff dff_B_x53bLicH9_0(.din(w_dff_B_s2xF01Tw8_0),.dout(w_dff_B_x53bLicH9_0),.clk(gclk));
	jdff dff_B_7K6smtvZ2_0(.din(w_dff_B_x53bLicH9_0),.dout(w_dff_B_7K6smtvZ2_0),.clk(gclk));
	jdff dff_B_hlrUaGM92_0(.din(w_dff_B_7K6smtvZ2_0),.dout(w_dff_B_hlrUaGM92_0),.clk(gclk));
	jdff dff_B_A1m94hoT3_0(.din(w_dff_B_hlrUaGM92_0),.dout(w_dff_B_A1m94hoT3_0),.clk(gclk));
	jdff dff_A_eiLXe4z73_0(.dout(w_n1049_0[0]),.din(w_dff_A_eiLXe4z73_0),.clk(gclk));
	jdff dff_A_VyKc0K8E5_0(.dout(w_dff_A_eiLXe4z73_0),.din(w_dff_A_VyKc0K8E5_0),.clk(gclk));
	jdff dff_A_ErRjlPQp7_1(.dout(w_n1049_0[1]),.din(w_dff_A_ErRjlPQp7_1),.clk(gclk));
	jdff dff_A_d0PiL9Ll8_1(.dout(w_dff_A_ErRjlPQp7_1),.din(w_dff_A_d0PiL9Ll8_1),.clk(gclk));
	jdff dff_B_zF4bDGEv2_0(.din(n1048),.dout(w_dff_B_zF4bDGEv2_0),.clk(gclk));
	jdff dff_B_yo14BoqS2_0(.din(n1047),.dout(w_dff_B_yo14BoqS2_0),.clk(gclk));
	jdff dff_B_9n6A3Gqv3_0(.din(n1045),.dout(w_dff_B_9n6A3Gqv3_0),.clk(gclk));
	jdff dff_B_752wZbhv8_0(.din(w_dff_B_9n6A3Gqv3_0),.dout(w_dff_B_752wZbhv8_0),.clk(gclk));
	jdff dff_B_tlh8MtPP5_0(.din(w_dff_B_752wZbhv8_0),.dout(w_dff_B_tlh8MtPP5_0),.clk(gclk));
	jdff dff_B_81nv7xqY1_0(.din(w_dff_B_tlh8MtPP5_0),.dout(w_dff_B_81nv7xqY1_0),.clk(gclk));
	jdff dff_B_fHRJB02K1_0(.din(w_dff_B_81nv7xqY1_0),.dout(w_dff_B_fHRJB02K1_0),.clk(gclk));
	jdff dff_B_ZHxKTDeG8_0(.din(n1044),.dout(w_dff_B_ZHxKTDeG8_0),.clk(gclk));
	jdff dff_B_y7op2Qz88_0(.din(w_dff_B_ZHxKTDeG8_0),.dout(w_dff_B_y7op2Qz88_0),.clk(gclk));
	jdff dff_B_tXmdT7kn9_0(.din(n1042),.dout(w_dff_B_tXmdT7kn9_0),.clk(gclk));
	jdff dff_B_tM3qn2Od9_0(.din(w_dff_B_tXmdT7kn9_0),.dout(w_dff_B_tM3qn2Od9_0),.clk(gclk));
	jdff dff_B_k4bCUjyl2_1(.din(n1030),.dout(w_dff_B_k4bCUjyl2_1),.clk(gclk));
	jdff dff_B_kvLmbFC01_1(.din(n1032),.dout(w_dff_B_kvLmbFC01_1),.clk(gclk));
	jdff dff_B_KHdMP5A09_1(.din(w_dff_B_kvLmbFC01_1),.dout(w_dff_B_KHdMP5A09_1),.clk(gclk));
	jdff dff_B_v6lCpZNv0_1(.din(n1035),.dout(w_dff_B_v6lCpZNv0_1),.clk(gclk));
	jdff dff_B_sHvM5Zr10_1(.din(n1027),.dout(w_dff_B_sHvM5Zr10_1),.clk(gclk));
	jdff dff_B_ksxvGuGo3_0(.din(n1028),.dout(w_dff_B_ksxvGuGo3_0),.clk(gclk));
	jdff dff_B_p51TAtIC9_1(.din(n1015),.dout(w_dff_B_p51TAtIC9_1),.clk(gclk));
	jdff dff_B_W72VKEnG4_1(.din(n1017),.dout(w_dff_B_W72VKEnG4_1),.clk(gclk));
	jdff dff_B_cJrdyOfY6_1(.din(n1020),.dout(w_dff_B_cJrdyOfY6_1),.clk(gclk));
	jdff dff_B_AGdyaDFT8_1(.din(n1021),.dout(w_dff_B_AGdyaDFT8_1),.clk(gclk));
	jdff dff_B_t1VZo9LU6_1(.din(n1011),.dout(w_dff_B_t1VZo9LU6_1),.clk(gclk));
	jdff dff_B_deyEznqR1_0(.din(n1013),.dout(w_dff_B_deyEznqR1_0),.clk(gclk));
	jdff dff_A_zYWUnwFe9_1(.dout(w_G125_0[1]),.din(w_dff_A_zYWUnwFe9_1),.clk(gclk));
	jdff dff_B_z6jI8JOq8_2(.din(G125),.dout(w_dff_B_z6jI8JOq8_2),.clk(gclk));
	jdff dff_B_xzqu5O5B4_2(.din(w_dff_B_z6jI8JOq8_2),.dout(w_dff_B_xzqu5O5B4_2),.clk(gclk));
	jdff dff_B_KScad4zf5_2(.din(w_dff_B_xzqu5O5B4_2),.dout(w_dff_B_KScad4zf5_2),.clk(gclk));
	jdff dff_A_cVaFdaMv6_1(.dout(w_n990_0[1]),.din(w_dff_A_cVaFdaMv6_1),.clk(gclk));
	jdff dff_A_5CpDEeKf6_1(.dout(w_dff_A_cVaFdaMv6_1),.din(w_dff_A_5CpDEeKf6_1),.clk(gclk));
	jdff dff_A_eiKxvlwp6_0(.dout(w_n758_0[0]),.din(w_dff_A_eiKxvlwp6_0),.clk(gclk));
	jdff dff_A_GonUom6y9_1(.dout(w_n758_0[1]),.din(w_dff_A_GonUom6y9_1),.clk(gclk));
	jdff dff_A_4S7ROmRl3_1(.dout(w_dff_A_GonUom6y9_1),.din(w_dff_A_4S7ROmRl3_1),.clk(gclk));
	jdff dff_A_FYu6yqkl2_1(.dout(w_dff_A_4S7ROmRl3_1),.din(w_dff_A_FYu6yqkl2_1),.clk(gclk));
	jdff dff_A_um81YCu52_0(.dout(w_n754_0[0]),.din(w_dff_A_um81YCu52_0),.clk(gclk));
	jdff dff_B_6DSs9HIL1_0(.din(n768),.dout(w_dff_B_6DSs9HIL1_0),.clk(gclk));
	jdff dff_B_EcZ0iLGm0_0(.din(n767),.dout(w_dff_B_EcZ0iLGm0_0),.clk(gclk));
	jdff dff_B_SMxFCpd09_0(.din(w_dff_B_EcZ0iLGm0_0),.dout(w_dff_B_SMxFCpd09_0),.clk(gclk));
	jdff dff_B_hlRPCz2F6_0(.din(w_dff_B_SMxFCpd09_0),.dout(w_dff_B_hlRPCz2F6_0),.clk(gclk));
	jdff dff_A_WKicSeMw9_2(.dout(w_n764_1[2]),.din(w_dff_A_WKicSeMw9_2),.clk(gclk));
	jdff dff_A_S7H7Geem3_2(.dout(w_dff_A_WKicSeMw9_2),.din(w_dff_A_S7H7Geem3_2),.clk(gclk));
	jdff dff_A_DxjuNRJs4_1(.dout(w_n1183_0[1]),.din(w_dff_A_DxjuNRJs4_1),.clk(gclk));
	jdff dff_B_CR3BjyFH6_1(.din(n1179),.dout(w_dff_B_CR3BjyFH6_1),.clk(gclk));
	jdff dff_B_ZOIj791h4_1(.din(w_dff_B_CR3BjyFH6_1),.dout(w_dff_B_ZOIj791h4_1),.clk(gclk));
	jdff dff_B_PLRJ6Etj9_1(.din(n1180),.dout(w_dff_B_PLRJ6Etj9_1),.clk(gclk));
	jdff dff_B_lEZiYtB29_1(.din(w_dff_B_PLRJ6Etj9_1),.dout(w_dff_B_lEZiYtB29_1),.clk(gclk));
	jdff dff_B_oBSGK8As4_1(.din(w_dff_B_lEZiYtB29_1),.dout(w_dff_B_oBSGK8As4_1),.clk(gclk));
	jdff dff_A_CngO7eVm1_0(.dout(w_n988_0[0]),.din(w_dff_A_CngO7eVm1_0),.clk(gclk));
	jdff dff_A_qKqgdtiq5_0(.dout(w_dff_A_CngO7eVm1_0),.din(w_dff_A_qKqgdtiq5_0),.clk(gclk));
	jdff dff_A_Z6o3NE1T2_1(.dout(w_n988_0[1]),.din(w_dff_A_Z6o3NE1T2_1),.clk(gclk));
	jdff dff_B_eB3cxISy9_0(.din(n986),.dout(w_dff_B_eB3cxISy9_0),.clk(gclk));
	jdff dff_B_oI9jQJTi4_0(.din(w_dff_B_eB3cxISy9_0),.dout(w_dff_B_oI9jQJTi4_0),.clk(gclk));
	jdff dff_B_tikuyAyg4_0(.din(n984),.dout(w_dff_B_tikuyAyg4_0),.clk(gclk));
	jdff dff_B_5nXq0wmB1_0(.din(w_dff_B_tikuyAyg4_0),.dout(w_dff_B_5nXq0wmB1_0),.clk(gclk));
	jdff dff_B_33rMplyV5_0(.din(w_dff_B_5nXq0wmB1_0),.dout(w_dff_B_33rMplyV5_0),.clk(gclk));
	jdff dff_B_iMrcfwYr1_0(.din(w_dff_B_33rMplyV5_0),.dout(w_dff_B_iMrcfwYr1_0),.clk(gclk));
	jdff dff_B_6sQkVDE55_0(.din(n983),.dout(w_dff_B_6sQkVDE55_0),.clk(gclk));
	jdff dff_B_Qr37CMcf9_0(.din(w_dff_B_6sQkVDE55_0),.dout(w_dff_B_Qr37CMcf9_0),.clk(gclk));
	jdff dff_B_yRhTEGI11_1(.din(n979),.dout(w_dff_B_yRhTEGI11_1),.clk(gclk));
	jdff dff_B_K02sLONx8_1(.din(w_dff_B_yRhTEGI11_1),.dout(w_dff_B_K02sLONx8_1),.clk(gclk));
	jdff dff_B_s7OrRFQo7_0(.din(n980),.dout(w_dff_B_s7OrRFQo7_0),.clk(gclk));
	jdff dff_A_nM5IVhfx6_2(.dout(w_G97_2[2]),.din(w_dff_A_nM5IVhfx6_2),.clk(gclk));
	jdff dff_B_Bm1gAG0j2_2(.din(n144),.dout(w_dff_B_Bm1gAG0j2_2),.clk(gclk));
	jdff dff_B_R0hu89kZ0_1(.din(n142),.dout(w_dff_B_R0hu89kZ0_1),.clk(gclk));
	jdff dff_B_Ir9qfCf96_1(.din(n966),.dout(w_dff_B_Ir9qfCf96_1),.clk(gclk));
	jdff dff_B_gXHOsSIl6_1(.din(n968),.dout(w_dff_B_gXHOsSIl6_1),.clk(gclk));
	jdff dff_B_X01pjMDj1_1(.din(n971),.dout(w_dff_B_X01pjMDj1_1),.clk(gclk));
	jdff dff_B_GlulZvDF5_0(.din(n972),.dout(w_dff_B_GlulZvDF5_0),.clk(gclk));
	jdff dff_A_fBl11jYt5_0(.dout(w_G143_1[0]),.din(w_dff_A_fBl11jYt5_0),.clk(gclk));
	jdff dff_A_7O4GBKmN5_2(.dout(w_G143_1[2]),.din(w_dff_A_7O4GBKmN5_2),.clk(gclk));
	jdff dff_A_zHTm3kUb4_1(.dout(w_G33_4[1]),.din(w_dff_A_zHTm3kUb4_1),.clk(gclk));
	jdff dff_A_4DfnUYM06_1(.dout(w_dff_A_zHTm3kUb4_1),.din(w_dff_A_4DfnUYM06_1),.clk(gclk));
	jdff dff_A_BQrbGPB64_1(.dout(w_dff_A_4DfnUYM06_1),.din(w_dff_A_BQrbGPB64_1),.clk(gclk));
	jdff dff_A_b9LAaO2V4_1(.dout(w_dff_A_BQrbGPB64_1),.din(w_dff_A_b9LAaO2V4_1),.clk(gclk));
	jdff dff_A_1ReQ3rI60_2(.dout(w_G33_4[2]),.din(w_dff_A_1ReQ3rI60_2),.clk(gclk));
	jdff dff_A_sRJo8vKp0_2(.dout(w_dff_A_1ReQ3rI60_2),.din(w_dff_A_sRJo8vKp0_2),.clk(gclk));
	jdff dff_A_c6IZV7De9_2(.dout(w_dff_A_sRJo8vKp0_2),.din(w_dff_A_c6IZV7De9_2),.clk(gclk));
	jdff dff_A_o4VBRHSQ5_2(.dout(w_dff_A_c6IZV7De9_2),.din(w_dff_A_o4VBRHSQ5_2),.clk(gclk));
	jdff dff_B_p93FT1pd2_0(.din(n964),.dout(w_dff_B_p93FT1pd2_0),.clk(gclk));
	jdff dff_A_ESKtCnJ84_1(.dout(w_n962_0[1]),.din(w_dff_A_ESKtCnJ84_1),.clk(gclk));
	jdff dff_B_DvXIxyGf4_1(.din(n951),.dout(w_dff_B_DvXIxyGf4_1),.clk(gclk));
	jdff dff_B_0qytQobt8_1(.din(n953),.dout(w_dff_B_0qytQobt8_1),.clk(gclk));
	jdff dff_B_Sa8S6l657_1(.din(n956),.dout(w_dff_B_Sa8S6l657_1),.clk(gclk));
	jdff dff_B_LXJkArUv7_0(.din(n957),.dout(w_dff_B_LXJkArUv7_0),.clk(gclk));
	jdff dff_B_3BYFU6wk9_1(.din(n947),.dout(w_dff_B_3BYFU6wk9_1),.clk(gclk));
	jdff dff_B_5wy3jEUG6_0(.din(n949),.dout(w_dff_B_5wy3jEUG6_0),.clk(gclk));
	jdff dff_A_tkWQIFCO0_0(.dout(w_n603_1[0]),.din(w_dff_A_tkWQIFCO0_0),.clk(gclk));
	jdff dff_A_KXPvJ4ay2_0(.dout(w_dff_A_tkWQIFCO0_0),.din(w_dff_A_KXPvJ4ay2_0),.clk(gclk));
	jdff dff_A_dYboeQ0R9_0(.dout(w_dff_A_KXPvJ4ay2_0),.din(w_dff_A_dYboeQ0R9_0),.clk(gclk));
	jdff dff_B_3E3bFULf8_1(.din(n850),.dout(w_dff_B_3E3bFULf8_1),.clk(gclk));
	jdff dff_B_mkW20p8i4_1(.din(w_dff_B_3E3bFULf8_1),.dout(w_dff_B_mkW20p8i4_1),.clk(gclk));
	jdff dff_B_hyFfmExd2_1(.din(w_dff_B_mkW20p8i4_1),.dout(w_dff_B_hyFfmExd2_1),.clk(gclk));
	jdff dff_B_O7F5IWIJ2_1(.din(w_dff_B_hyFfmExd2_1),.dout(w_dff_B_O7F5IWIJ2_1),.clk(gclk));
	jdff dff_B_9yN6e0JT4_1(.din(w_dff_B_O7F5IWIJ2_1),.dout(w_dff_B_9yN6e0JT4_1),.clk(gclk));
	jdff dff_B_enNp6FUD9_1(.din(w_dff_B_9yN6e0JT4_1),.dout(w_dff_B_enNp6FUD9_1),.clk(gclk));
	jdff dff_B_wBvIRgVB2_0(.din(n875),.dout(w_dff_B_wBvIRgVB2_0),.clk(gclk));
	jdff dff_B_i61UwHm20_0(.din(w_dff_B_wBvIRgVB2_0),.dout(w_dff_B_i61UwHm20_0),.clk(gclk));
	jdff dff_B_XYbubFso9_1(.din(n871),.dout(w_dff_B_XYbubFso9_1),.clk(gclk));
	jdff dff_B_lULTa84t5_1(.din(n868),.dout(w_dff_B_lULTa84t5_1),.clk(gclk));
	jdff dff_B_xGC1GvKU7_1(.din(w_dff_B_lULTa84t5_1),.dout(w_dff_B_xGC1GvKU7_1),.clk(gclk));
	jdff dff_B_21piD6Tr0_1(.din(w_dff_B_xGC1GvKU7_1),.dout(w_dff_B_21piD6Tr0_1),.clk(gclk));
	jdff dff_B_RDsmvoLr7_1(.din(w_dff_B_21piD6Tr0_1),.dout(w_dff_B_RDsmvoLr7_1),.clk(gclk));
	jdff dff_B_cj0UxHTU6_1(.din(w_dff_B_RDsmvoLr7_1),.dout(w_dff_B_cj0UxHTU6_1),.clk(gclk));
	jdff dff_A_oKGk8L4T6_1(.dout(w_n861_1[1]),.din(w_dff_A_oKGk8L4T6_1),.clk(gclk));
	jdff dff_A_yC7bLEO03_1(.dout(w_dff_A_oKGk8L4T6_1),.din(w_dff_A_yC7bLEO03_1),.clk(gclk));
	jdff dff_A_dDvpsJed7_2(.dout(w_n861_0[2]),.din(w_dff_A_dDvpsJed7_2),.clk(gclk));
	jdff dff_A_eTrHz4jv8_2(.dout(w_dff_A_dDvpsJed7_2),.din(w_dff_A_eTrHz4jv8_2),.clk(gclk));
	jdff dff_B_2BHfzlba9_0(.din(n860),.dout(w_dff_B_2BHfzlba9_0),.clk(gclk));
	jdff dff_B_0fop6hgz9_0(.din(n857),.dout(w_dff_B_0fop6hgz9_0),.clk(gclk));
	jdff dff_B_R8jO07tz9_0(.din(w_dff_B_0fop6hgz9_0),.dout(w_dff_B_R8jO07tz9_0),.clk(gclk));
	jdff dff_B_oPHEf5Ne0_0(.din(w_dff_B_R8jO07tz9_0),.dout(w_dff_B_oPHEf5Ne0_0),.clk(gclk));
	jdff dff_A_gSZHdEuL1_1(.dout(w_n563_0[1]),.din(w_dff_A_gSZHdEuL1_1),.clk(gclk));
	jdff dff_A_5IFVUyto1_1(.dout(w_dff_A_gSZHdEuL1_1),.din(w_dff_A_5IFVUyto1_1),.clk(gclk));
	jdff dff_A_uXJjowcO9_2(.dout(w_n563_0[2]),.din(w_dff_A_uXJjowcO9_2),.clk(gclk));
	jdff dff_A_6Uj6uu5l7_2(.dout(w_dff_A_uXJjowcO9_2),.din(w_dff_A_6Uj6uu5l7_2),.clk(gclk));
	jdff dff_B_7uHF89Yi2_1(.din(n555),.dout(w_dff_B_7uHF89Yi2_1),.clk(gclk));
	jdff dff_B_OGNkaMNl4_1(.din(w_dff_B_7uHF89Yi2_1),.dout(w_dff_B_OGNkaMNl4_1),.clk(gclk));
	jdff dff_B_wzSXzrlF4_1(.din(w_dff_B_OGNkaMNl4_1),.dout(w_dff_B_wzSXzrlF4_1),.clk(gclk));
	jdff dff_B_pAxHbsCu2_0(.din(n849),.dout(w_dff_B_pAxHbsCu2_0),.clk(gclk));
	jdff dff_B_Aj2D0Oer9_0(.din(w_dff_B_pAxHbsCu2_0),.dout(w_dff_B_Aj2D0Oer9_0),.clk(gclk));
	jdff dff_B_8eWT5FLm1_0(.din(n848),.dout(w_dff_B_8eWT5FLm1_0),.clk(gclk));
	jdff dff_B_UMGtMZK97_0(.din(w_dff_B_8eWT5FLm1_0),.dout(w_dff_B_UMGtMZK97_0),.clk(gclk));
	jdff dff_B_dCLelrxZ8_0(.din(w_dff_B_UMGtMZK97_0),.dout(w_dff_B_dCLelrxZ8_0),.clk(gclk));
	jdff dff_B_qBCX1vVK1_0(.din(w_dff_B_dCLelrxZ8_0),.dout(w_dff_B_qBCX1vVK1_0),.clk(gclk));
	jdff dff_B_WX1OM9gd9_1(.din(n844),.dout(w_dff_B_WX1OM9gd9_1),.clk(gclk));
	jdff dff_B_xoQRnqys4_1(.din(w_dff_B_WX1OM9gd9_1),.dout(w_dff_B_xoQRnqys4_1),.clk(gclk));
	jdff dff_B_kFkvmHd54_0(.din(n845),.dout(w_dff_B_kFkvmHd54_0),.clk(gclk));
	jdff dff_A_R8JEbloF5_0(.dout(w_n131_0[0]),.din(w_dff_A_R8JEbloF5_0),.clk(gclk));
	jdff dff_B_kUtKdGEd3_1(.din(n129),.dout(w_dff_B_kUtKdGEd3_1),.clk(gclk));
	jdff dff_B_8Mwsvgde1_1(.din(n820),.dout(w_dff_B_8Mwsvgde1_1),.clk(gclk));
	jdff dff_B_fgFE3RpO0_1(.din(w_dff_B_8Mwsvgde1_1),.dout(w_dff_B_fgFE3RpO0_1),.clk(gclk));
	jdff dff_B_L0ZsuJQK0_1(.din(n828),.dout(w_dff_B_L0ZsuJQK0_1),.clk(gclk));
	jdff dff_B_9AAzravt8_1(.din(n830),.dout(w_dff_B_9AAzravt8_1),.clk(gclk));
	jdff dff_B_1vTMB9525_1(.din(w_dff_B_9AAzravt8_1),.dout(w_dff_B_1vTMB9525_1),.clk(gclk));
	jdff dff_B_gaXse5MV6_1(.din(n833),.dout(w_dff_B_gaXse5MV6_1),.clk(gclk));
	jdff dff_B_PnW7Xyv40_1(.din(n834),.dout(w_dff_B_PnW7Xyv40_1),.clk(gclk));
	jdff dff_B_Ndnd0jB51_1(.din(n822),.dout(w_dff_B_Ndnd0jB51_1),.clk(gclk));
	jdff dff_B_yM0ra25v9_1(.din(n809),.dout(w_dff_B_yM0ra25v9_1),.clk(gclk));
	jdff dff_B_AHrNX2v01_1(.din(n811),.dout(w_dff_B_AHrNX2v01_1),.clk(gclk));
	jdff dff_B_KHWzBYxD2_1(.din(n814),.dout(w_dff_B_KHWzBYxD2_1),.clk(gclk));
	jdff dff_B_oPSouTSc8_1(.din(n815),.dout(w_dff_B_oPSouTSc8_1),.clk(gclk));
	jdff dff_B_GKEavJx33_1(.din(n805),.dout(w_dff_B_GKEavJx33_1),.clk(gclk));
	jdff dff_B_AFA9y1HW5_0(.din(n807),.dout(w_dff_B_AFA9y1HW5_0),.clk(gclk));
	jdff dff_A_8nC7ayYu1_2(.dout(w_G107_2[2]),.din(w_dff_A_8nC7ayYu1_2),.clk(gclk));
	jdff dff_A_pZGfTmqq0_0(.dout(w_n801_0[0]),.din(w_dff_A_pZGfTmqq0_0),.clk(gclk));
	jdff dff_A_GPNj94e26_0(.dout(w_dff_A_pZGfTmqq0_0),.din(w_dff_A_GPNj94e26_0),.clk(gclk));
	jdff dff_A_Wsg0HdUG1_0(.dout(w_dff_A_GPNj94e26_0),.din(w_dff_A_Wsg0HdUG1_0),.clk(gclk));
	jdff dff_A_ETicKf2s9_0(.dout(w_dff_A_Wsg0HdUG1_0),.din(w_dff_A_ETicKf2s9_0),.clk(gclk));
	jdff dff_B_GTkGHyzu7_0(.din(n800),.dout(w_dff_B_GTkGHyzu7_0),.clk(gclk));
	jdff dff_B_t8wk4rsF8_0(.din(n798),.dout(w_dff_B_t8wk4rsF8_0),.clk(gclk));
	jdff dff_A_i3FCZTXW0_0(.dout(w_n797_0[0]),.din(w_dff_A_i3FCZTXW0_0),.clk(gclk));
	jdff dff_B_YUHFmixx5_0(.din(n936),.dout(w_dff_B_YUHFmixx5_0),.clk(gclk));
	jdff dff_B_U9NVKsvB8_0(.din(w_dff_B_YUHFmixx5_0),.dout(w_dff_B_U9NVKsvB8_0),.clk(gclk));
	jdff dff_B_Lcvoh0Hp3_0(.din(n935),.dout(w_dff_B_Lcvoh0Hp3_0),.clk(gclk));
	jdff dff_B_v8COqiHe8_0(.din(n934),.dout(w_dff_B_v8COqiHe8_0),.clk(gclk));
	jdff dff_B_GFBcvfg54_0(.din(w_dff_B_v8COqiHe8_0),.dout(w_dff_B_GFBcvfg54_0),.clk(gclk));
	jdff dff_B_GmrysAj40_1(.din(n924),.dout(w_dff_B_GmrysAj40_1),.clk(gclk));
	jdff dff_B_MUofsgPe6_1(.din(n925),.dout(w_dff_B_MUofsgPe6_1),.clk(gclk));
	jdff dff_B_BDtRMv4D3_1(.din(n916),.dout(w_dff_B_BDtRMv4D3_1),.clk(gclk));
	jdff dff_B_c9gsHbY27_1(.din(w_dff_B_BDtRMv4D3_1),.dout(w_dff_B_c9gsHbY27_1),.clk(gclk));
	jdff dff_B_9szqQOzh1_1(.din(n918),.dout(w_dff_B_9szqQOzh1_1),.clk(gclk));
	jdff dff_A_zyINY7Mr6_1(.dout(w_n73_1[1]),.din(w_dff_A_zyINY7Mr6_1),.clk(gclk));
	jdff dff_A_pt9RtHEF4_1(.dout(w_n135_0[1]),.din(w_dff_A_pt9RtHEF4_1),.clk(gclk));
	jdff dff_B_tZwGx5NQ2_1(.din(n133),.dout(w_dff_B_tZwGx5NQ2_1),.clk(gclk));
	jdff dff_B_snBJIKE72_1(.din(n902),.dout(w_dff_B_snBJIKE72_1),.clk(gclk));
	jdff dff_B_T0JGSakf5_1(.din(n904),.dout(w_dff_B_T0JGSakf5_1),.clk(gclk));
	jdff dff_B_m1toFi2Z4_1(.din(n907),.dout(w_dff_B_m1toFi2Z4_1),.clk(gclk));
	jdff dff_B_w8ZFtNkY0_1(.din(n908),.dout(w_dff_B_w8ZFtNkY0_1),.clk(gclk));
	jdff dff_A_h0HBtqJs8_0(.dout(w_G50_2[0]),.din(w_dff_A_h0HBtqJs8_0),.clk(gclk));
	jdff dff_A_1Rn6NAIO0_1(.dout(w_G68_2[1]),.din(w_dff_A_1Rn6NAIO0_1),.clk(gclk));
	jdff dff_A_zKbeWLTF1_1(.dout(w_dff_A_1Rn6NAIO0_1),.din(w_dff_A_zKbeWLTF1_1),.clk(gclk));
	jdff dff_A_6c3adLdN9_1(.dout(w_dff_A_zKbeWLTF1_1),.din(w_dff_A_6c3adLdN9_1),.clk(gclk));
	jdff dff_A_UxMnkg5s0_2(.dout(w_G68_2[2]),.din(w_dff_A_UxMnkg5s0_2),.clk(gclk));
	jdff dff_A_hQjLbY4h4_2(.dout(w_dff_A_UxMnkg5s0_2),.din(w_dff_A_hQjLbY4h4_2),.clk(gclk));
	jdff dff_A_enpvF3rt7_2(.dout(w_dff_A_hQjLbY4h4_2),.din(w_dff_A_enpvF3rt7_2),.clk(gclk));
	jdff dff_A_JUOYulXY2_2(.dout(w_dff_A_enpvF3rt7_2),.din(w_dff_A_JUOYulXY2_2),.clk(gclk));
	jdff dff_A_iF5cVrWG1_1(.dout(w_G150_2[1]),.din(w_dff_A_iF5cVrWG1_1),.clk(gclk));
	jdff dff_B_qmhAqa5p4_0(.din(n900),.dout(w_dff_B_qmhAqa5p4_0),.clk(gclk));
	jdff dff_A_3nb9wQt70_0(.dout(w_G58_2[0]),.din(w_dff_A_3nb9wQt70_0),.clk(gclk));
	jdff dff_A_SLHqwUK49_0(.dout(w_dff_A_3nb9wQt70_0),.din(w_dff_A_SLHqwUK49_0),.clk(gclk));
	jdff dff_A_tqFOGh5y3_2(.dout(w_G58_2[2]),.din(w_dff_A_tqFOGh5y3_2),.clk(gclk));
	jdff dff_A_gfeH5r0M2_2(.dout(w_dff_A_tqFOGh5y3_2),.din(w_dff_A_gfeH5r0M2_2),.clk(gclk));
	jdff dff_B_7xFu4Mi80_1(.din(n887),.dout(w_dff_B_7xFu4Mi80_1),.clk(gclk));
	jdff dff_B_1ecaiyHG9_1(.din(n889),.dout(w_dff_B_1ecaiyHG9_1),.clk(gclk));
	jdff dff_B_rwqpw1ea0_0(.din(n895),.dout(w_dff_B_rwqpw1ea0_0),.clk(gclk));
	jdff dff_B_eC3jd1QQ4_0(.din(n891),.dout(w_dff_B_eC3jd1QQ4_0),.clk(gclk));
	jdff dff_A_Mokb2Ozp2_1(.dout(w_G116_2[1]),.din(w_dff_A_Mokb2Ozp2_1),.clk(gclk));
	jdff dff_A_wPCjnRXx0_2(.dout(w_G116_2[2]),.din(w_dff_A_wPCjnRXx0_2),.clk(gclk));
	jdff dff_B_dxEGLWIz7_1(.din(n883),.dout(w_dff_B_dxEGLWIz7_1),.clk(gclk));
	jdff dff_B_xN7FYkZb6_0(.din(n885),.dout(w_dff_B_xN7FYkZb6_0),.clk(gclk));
	jdff dff_A_5d8bTIn96_0(.dout(w_G283_2[0]),.din(w_dff_A_5d8bTIn96_0),.clk(gclk));
	jdff dff_A_WFItt2iM5_1(.dout(w_G283_2[1]),.din(w_dff_A_WFItt2iM5_1),.clk(gclk));
	jdff dff_A_xeZgGkv54_1(.dout(w_n564_0[1]),.din(w_dff_A_xeZgGkv54_1),.clk(gclk));
	jdff dff_B_YfXokUhJ7_1(.din(n878),.dout(w_dff_B_YfXokUhJ7_1),.clk(gclk));
	jdff dff_B_J8ntFLjC9_1(.din(w_dff_B_YfXokUhJ7_1),.dout(w_dff_B_J8ntFLjC9_1),.clk(gclk));
	jdff dff_A_bJUmiIhN1_0(.dout(w_n589_1[0]),.din(w_dff_A_bJUmiIhN1_0),.clk(gclk));
	jdff dff_A_DJibnqLW6_0(.dout(w_dff_A_bJUmiIhN1_0),.din(w_dff_A_DJibnqLW6_0),.clk(gclk));
	jdff dff_A_vSvLhwb24_0(.dout(w_dff_A_DJibnqLW6_0),.din(w_dff_A_vSvLhwb24_0),.clk(gclk));
	jdff dff_A_DKsOg8qe2_0(.dout(w_n592_1[0]),.din(w_dff_A_DKsOg8qe2_0),.clk(gclk));
	jdff dff_A_hhZyU8L87_0(.dout(w_dff_A_DKsOg8qe2_0),.din(w_dff_A_hhZyU8L87_0),.clk(gclk));
	jdff dff_A_jQ3tBIKF0_1(.dout(w_n592_1[1]),.din(w_dff_A_jQ3tBIKF0_1),.clk(gclk));
	jdff dff_B_nXU4JbEZ0_0(.din(n852),.dout(w_dff_B_nXU4JbEZ0_0),.clk(gclk));
	jdff dff_B_Po7JYX890_0(.din(n560),.dout(w_dff_B_Po7JYX890_0),.clk(gclk));
	jdff dff_B_PYgns8GG8_2(.din(n556),.dout(w_dff_B_PYgns8GG8_2),.clk(gclk));
	jdff dff_B_ce4VxpCZ8_2(.din(w_dff_B_PYgns8GG8_2),.dout(w_dff_B_ce4VxpCZ8_2),.clk(gclk));
	jdff dff_A_YBcPvg7h7_0(.dout(w_G396_0[0]),.din(w_dff_A_YBcPvg7h7_0),.clk(gclk));
	jdff dff_A_yv4guX720_0(.dout(w_dff_A_YBcPvg7h7_0),.din(w_dff_A_yv4guX720_0),.clk(gclk));
	jdff dff_A_lE3ItQU19_0(.dout(w_dff_A_yv4guX720_0),.din(w_dff_A_lE3ItQU19_0),.clk(gclk));
	jdff dff_B_OPDiObkS2_0(.din(n687),.dout(w_dff_B_OPDiObkS2_0),.clk(gclk));
	jdff dff_B_B7tUwYuz5_0(.din(w_dff_B_OPDiObkS2_0),.dout(w_dff_B_B7tUwYuz5_0),.clk(gclk));
	jdff dff_B_1XT9siGY6_0(.din(n686),.dout(w_dff_B_1XT9siGY6_0),.clk(gclk));
	jdff dff_B_9ylm8g6g4_0(.din(w_dff_B_1XT9siGY6_0),.dout(w_dff_B_9ylm8g6g4_0),.clk(gclk));
	jdff dff_B_7n2j4Y9q1_1(.din(n678),.dout(w_dff_B_7n2j4Y9q1_1),.clk(gclk));
	jdff dff_B_ni6NVzVi8_1(.din(n679),.dout(w_dff_B_ni6NVzVi8_1),.clk(gclk));
	jdff dff_B_WhCIUObC5_2(.din(n680),.dout(w_dff_B_WhCIUObC5_2),.clk(gclk));
	jdff dff_B_ydfoAbKT5_1(.din(n673),.dout(w_dff_B_ydfoAbKT5_1),.clk(gclk));
	jdff dff_B_LvqtFccj9_1(.din(w_dff_B_ydfoAbKT5_1),.dout(w_dff_B_LvqtFccj9_1),.clk(gclk));
	jdff dff_B_0eotRJax5_0(.din(n139),.dout(w_dff_B_0eotRJax5_0),.clk(gclk));
	jdff dff_A_H2vgC6kq4_1(.dout(w_n672_1[1]),.din(w_dff_A_H2vgC6kq4_1),.clk(gclk));
	jdff dff_A_rukccQz65_1(.dout(w_dff_A_H2vgC6kq4_1),.din(w_dff_A_rukccQz65_1),.clk(gclk));
	jdff dff_A_z8l9MxUk1_1(.dout(w_dff_A_rukccQz65_1),.din(w_dff_A_z8l9MxUk1_1),.clk(gclk));
	jdff dff_A_kcV6abiy0_2(.dout(w_n672_0[2]),.din(w_dff_A_kcV6abiy0_2),.clk(gclk));
	jdff dff_A_q1KqtH6B0_2(.dout(w_dff_A_kcV6abiy0_2),.din(w_dff_A_q1KqtH6B0_2),.clk(gclk));
	jdff dff_A_7ujfS0FO3_2(.dout(w_dff_A_q1KqtH6B0_2),.din(w_dff_A_7ujfS0FO3_2),.clk(gclk));
	jdff dff_B_hhfAUHHD0_1(.din(n647),.dout(w_dff_B_hhfAUHHD0_1),.clk(gclk));
	jdff dff_B_zPnQWszI8_1(.din(w_dff_B_hhfAUHHD0_1),.dout(w_dff_B_zPnQWszI8_1),.clk(gclk));
	jdff dff_B_KVHLBWXp4_1(.din(n653),.dout(w_dff_B_KVHLBWXp4_1),.clk(gclk));
	jdff dff_B_vOi2AvAE7_1(.din(w_dff_B_KVHLBWXp4_1),.dout(w_dff_B_vOi2AvAE7_1),.clk(gclk));
	jdff dff_B_x8aIJJoV5_1(.din(n656),.dout(w_dff_B_x8aIJJoV5_1),.clk(gclk));
	jdff dff_B_KEhFo1TO7_1(.din(n660),.dout(w_dff_B_KEhFo1TO7_1),.clk(gclk));
	jdff dff_B_3b1YSCjC9_0(.din(n658),.dout(w_dff_B_3b1YSCjC9_0),.clk(gclk));
	jdff dff_B_28z0T09I2_1(.din(n630),.dout(w_dff_B_28z0T09I2_1),.clk(gclk));
	jdff dff_B_grn3rGDj5_1(.din(n633),.dout(w_dff_B_grn3rGDj5_1),.clk(gclk));
	jdff dff_B_R2fQozyq6_0(.din(n644),.dout(w_dff_B_R2fQozyq6_0),.clk(gclk));
	jdff dff_A_ph7TJQJV6_0(.dout(w_G317_1[0]),.din(w_dff_A_ph7TJQJV6_0),.clk(gclk));
	jdff dff_B_3ps9KR4y8_3(.din(G317),.dout(w_dff_B_3ps9KR4y8_3),.clk(gclk));
	jdff dff_B_CKqL7Gir9_3(.din(w_dff_B_3ps9KR4y8_3),.dout(w_dff_B_CKqL7Gir9_3),.clk(gclk));
	jdff dff_B_CDR6Suz05_3(.din(w_dff_B_CKqL7Gir9_3),.dout(w_dff_B_CDR6Suz05_3),.clk(gclk));
	jdff dff_A_yyHutWcL6_0(.dout(w_G326_0[0]),.din(w_dff_A_yyHutWcL6_0),.clk(gclk));
	jdff dff_B_ndqBDG7m5_2(.din(G326),.dout(w_dff_B_ndqBDG7m5_2),.clk(gclk));
	jdff dff_B_wb4jpeK49_2(.din(w_dff_B_ndqBDG7m5_2),.dout(w_dff_B_wb4jpeK49_2),.clk(gclk));
	jdff dff_B_P0A9yaRt5_2(.din(w_dff_B_wb4jpeK49_2),.dout(w_dff_B_P0A9yaRt5_2),.clk(gclk));
	jdff dff_B_ueObpH249_0(.din(n637),.dout(w_dff_B_ueObpH249_0),.clk(gclk));
	jdff dff_B_jKyiDPet0_1(.din(G329),.dout(w_dff_B_jKyiDPet0_1),.clk(gclk));
	jdff dff_B_mCyouFB74_1(.din(w_dff_B_jKyiDPet0_1),.dout(w_dff_B_mCyouFB74_1),.clk(gclk));
	jdff dff_B_ogfKhUUA1_1(.din(w_dff_B_mCyouFB74_1),.dout(w_dff_B_ogfKhUUA1_1),.clk(gclk));
	jdff dff_B_X6hvEvIb3_1(.din(w_dff_B_ogfKhUUA1_1),.dout(w_dff_B_X6hvEvIb3_1),.clk(gclk));
	jdff dff_A_85JoKlax6_1(.dout(w_n148_5[1]),.din(w_dff_A_85JoKlax6_1),.clk(gclk));
	jdff dff_A_Dv6O1XCu5_1(.dout(w_dff_A_85JoKlax6_1),.din(w_dff_A_Dv6O1XCu5_1),.clk(gclk));
	jdff dff_A_tblrHz7F0_1(.dout(w_dff_A_Dv6O1XCu5_1),.din(w_dff_A_tblrHz7F0_1),.clk(gclk));
	jdff dff_A_9hkqwx6q6_2(.dout(w_n148_5[2]),.din(w_dff_A_9hkqwx6q6_2),.clk(gclk));
	jdff dff_A_kXzz8afe8_2(.dout(w_dff_A_9hkqwx6q6_2),.din(w_dff_A_kXzz8afe8_2),.clk(gclk));
	jdff dff_B_P6h9LSyK6_1(.din(n618),.dout(w_dff_B_P6h9LSyK6_1),.clk(gclk));
	jdff dff_B_iv6e9eD24_0(.din(n628),.dout(w_dff_B_iv6e9eD24_0),.clk(gclk));
	jdff dff_A_vhYSnYkN0_0(.dout(w_G322_0[0]),.din(w_dff_A_vhYSnYkN0_0),.clk(gclk));
	jdff dff_B_u7mi6eWz7_3(.din(G322),.dout(w_dff_B_u7mi6eWz7_3),.clk(gclk));
	jdff dff_B_2nFbqOQB2_3(.din(w_dff_B_u7mi6eWz7_3),.dout(w_dff_B_2nFbqOQB2_3),.clk(gclk));
	jdff dff_B_Y4As0ua57_3(.din(w_dff_B_2nFbqOQB2_3),.dout(w_dff_B_Y4As0ua57_3),.clk(gclk));
	jdff dff_A_MvBFLSK72_1(.dout(w_n612_4[1]),.din(w_dff_A_MvBFLSK72_1),.clk(gclk));
	jdff dff_A_h7TBsyZ56_1(.dout(w_dff_A_MvBFLSK72_1),.din(w_dff_A_h7TBsyZ56_1),.clk(gclk));
	jdff dff_A_ShlU2W4v1_1(.dout(w_dff_A_h7TBsyZ56_1),.din(w_dff_A_ShlU2W4v1_1),.clk(gclk));
	jdff dff_A_cHxiyPDX9_1(.dout(w_dff_A_ShlU2W4v1_1),.din(w_dff_A_cHxiyPDX9_1),.clk(gclk));
	jdff dff_A_liyqeJHw8_1(.dout(w_dff_A_cHxiyPDX9_1),.din(w_dff_A_liyqeJHw8_1),.clk(gclk));
	jdff dff_A_4sp08cSE4_1(.dout(w_dff_A_liyqeJHw8_1),.din(w_dff_A_4sp08cSE4_1),.clk(gclk));
	jdff dff_A_tgRMtliv9_1(.dout(w_dff_A_4sp08cSE4_1),.din(w_dff_A_tgRMtliv9_1),.clk(gclk));
	jdff dff_A_Jnrfl8BP3_1(.dout(w_dff_A_tgRMtliv9_1),.din(w_dff_A_Jnrfl8BP3_1),.clk(gclk));
	jdff dff_A_ljCR1h082_0(.dout(w_n608_1[0]),.din(w_dff_A_ljCR1h082_0),.clk(gclk));
	jdff dff_A_cX0ulFsR7_0(.dout(w_dff_A_ljCR1h082_0),.din(w_dff_A_cX0ulFsR7_0),.clk(gclk));
	jdff dff_A_9W79FXkf7_0(.dout(w_dff_A_cX0ulFsR7_0),.din(w_dff_A_9W79FXkf7_0),.clk(gclk));
	jdff dff_A_dMNaZEgX4_0(.dout(w_dff_A_9W79FXkf7_0),.din(w_dff_A_dMNaZEgX4_0),.clk(gclk));
	jdff dff_A_PuiCmZd40_0(.dout(w_dff_A_dMNaZEgX4_0),.din(w_dff_A_PuiCmZd40_0),.clk(gclk));
	jdff dff_A_v1azH6f15_0(.dout(w_dff_A_PuiCmZd40_0),.din(w_dff_A_v1azH6f15_0),.clk(gclk));
	jdff dff_A_SYZxXsO99_0(.dout(w_dff_A_v1azH6f15_0),.din(w_dff_A_SYZxXsO99_0),.clk(gclk));
	jdff dff_A_rLgAvqL93_0(.dout(w_dff_A_SYZxXsO99_0),.din(w_dff_A_rLgAvqL93_0),.clk(gclk));
	jdff dff_A_vrwR2ugt4_0(.dout(w_dff_A_rLgAvqL93_0),.din(w_dff_A_vrwR2ugt4_0),.clk(gclk));
	jdff dff_A_oZzRsgcd3_0(.dout(w_dff_A_vrwR2ugt4_0),.din(w_dff_A_oZzRsgcd3_0),.clk(gclk));
	jdff dff_A_UK7zN0hx1_0(.dout(w_dff_A_oZzRsgcd3_0),.din(w_dff_A_UK7zN0hx1_0),.clk(gclk));
	jdff dff_A_xEbno4Bc2_2(.dout(w_n608_1[2]),.din(w_dff_A_xEbno4Bc2_2),.clk(gclk));
	jdff dff_A_cKNOEeHX5_2(.dout(w_dff_A_xEbno4Bc2_2),.din(w_dff_A_cKNOEeHX5_2),.clk(gclk));
	jdff dff_A_tOdF6zHU2_2(.dout(w_dff_A_cKNOEeHX5_2),.din(w_dff_A_tOdF6zHU2_2),.clk(gclk));
	jdff dff_A_8DEhp2Yc7_2(.dout(w_dff_A_tOdF6zHU2_2),.din(w_dff_A_8DEhp2Yc7_2),.clk(gclk));
	jdff dff_A_RaGEzzcA5_2(.dout(w_dff_A_8DEhp2Yc7_2),.din(w_dff_A_RaGEzzcA5_2),.clk(gclk));
	jdff dff_A_6oFbUtcT3_2(.dout(w_dff_A_RaGEzzcA5_2),.din(w_dff_A_6oFbUtcT3_2),.clk(gclk));
	jdff dff_A_I8RgdFMX2_2(.dout(w_dff_A_6oFbUtcT3_2),.din(w_dff_A_I8RgdFMX2_2),.clk(gclk));
	jdff dff_A_sRVzXlW13_2(.dout(w_dff_A_I8RgdFMX2_2),.din(w_dff_A_sRVzXlW13_2),.clk(gclk));
	jdff dff_A_bkxMkfld2_2(.dout(w_dff_A_sRVzXlW13_2),.din(w_dff_A_bkxMkfld2_2),.clk(gclk));
	jdff dff_A_HqH1KDj88_2(.dout(w_dff_A_bkxMkfld2_2),.din(w_dff_A_HqH1KDj88_2),.clk(gclk));
	jdff dff_A_JRZ2oKPU4_2(.dout(w_dff_A_HqH1KDj88_2),.din(w_dff_A_JRZ2oKPU4_2),.clk(gclk));
	jdff dff_A_z5QvvfQZ2_1(.dout(w_n608_0[1]),.din(w_dff_A_z5QvvfQZ2_1),.clk(gclk));
	jdff dff_A_KQa0EXTd1_1(.dout(w_dff_A_z5QvvfQZ2_1),.din(w_dff_A_KQa0EXTd1_1),.clk(gclk));
	jdff dff_A_05YmZwlX5_1(.dout(w_dff_A_KQa0EXTd1_1),.din(w_dff_A_05YmZwlX5_1),.clk(gclk));
	jdff dff_A_S88yINAh8_1(.dout(w_dff_A_05YmZwlX5_1),.din(w_dff_A_S88yINAh8_1),.clk(gclk));
	jdff dff_A_1ametKsg4_1(.dout(w_dff_A_S88yINAh8_1),.din(w_dff_A_1ametKsg4_1),.clk(gclk));
	jdff dff_A_ceTfrecR8_1(.dout(w_dff_A_1ametKsg4_1),.din(w_dff_A_ceTfrecR8_1),.clk(gclk));
	jdff dff_A_VzSK2nFp8_1(.dout(w_dff_A_ceTfrecR8_1),.din(w_dff_A_VzSK2nFp8_1),.clk(gclk));
	jdff dff_A_UMGNIApm0_1(.dout(w_dff_A_VzSK2nFp8_1),.din(w_dff_A_UMGNIApm0_1),.clk(gclk));
	jdff dff_A_3k9j5T8S9_1(.dout(w_dff_A_UMGNIApm0_1),.din(w_dff_A_3k9j5T8S9_1),.clk(gclk));
	jdff dff_A_n0HXTEJQ5_1(.dout(w_dff_A_3k9j5T8S9_1),.din(w_dff_A_n0HXTEJQ5_1),.clk(gclk));
	jdff dff_A_mquicPis4_1(.dout(w_dff_A_n0HXTEJQ5_1),.din(w_dff_A_mquicPis4_1),.clk(gclk));
	jdff dff_A_iu21Zqse8_2(.dout(w_n608_0[2]),.din(w_dff_A_iu21Zqse8_2),.clk(gclk));
	jdff dff_A_bNb2Uc5A9_2(.dout(w_dff_A_iu21Zqse8_2),.din(w_dff_A_bNb2Uc5A9_2),.clk(gclk));
	jdff dff_A_Mho3DNf74_2(.dout(w_dff_A_bNb2Uc5A9_2),.din(w_dff_A_Mho3DNf74_2),.clk(gclk));
	jdff dff_A_CWuBi4A70_2(.dout(w_dff_A_Mho3DNf74_2),.din(w_dff_A_CWuBi4A70_2),.clk(gclk));
	jdff dff_A_fYj21vvD2_2(.dout(w_dff_A_CWuBi4A70_2),.din(w_dff_A_fYj21vvD2_2),.clk(gclk));
	jdff dff_A_2Yj3U0Ip8_2(.dout(w_dff_A_fYj21vvD2_2),.din(w_dff_A_2Yj3U0Ip8_2),.clk(gclk));
	jdff dff_A_fETiwb8L9_2(.dout(w_dff_A_2Yj3U0Ip8_2),.din(w_dff_A_fETiwb8L9_2),.clk(gclk));
	jdff dff_A_424xl1M53_2(.dout(w_dff_A_fETiwb8L9_2),.din(w_dff_A_424xl1M53_2),.clk(gclk));
	jdff dff_A_Axf6eWiB8_2(.dout(w_dff_A_424xl1M53_2),.din(w_dff_A_Axf6eWiB8_2),.clk(gclk));
	jdff dff_A_e4gAfepL0_2(.dout(w_dff_A_Axf6eWiB8_2),.din(w_dff_A_e4gAfepL0_2),.clk(gclk));
	jdff dff_A_cVKG9rir9_2(.dout(w_dff_A_e4gAfepL0_2),.din(w_dff_A_cVKG9rir9_2),.clk(gclk));
	jdff dff_B_pfinCzPT2_0(.din(n570),.dout(w_dff_B_pfinCzPT2_0),.clk(gclk));
	jdff dff_B_6MOx5bXI0_0(.din(w_dff_B_pfinCzPT2_0),.dout(w_dff_B_6MOx5bXI0_0),.clk(gclk));
	jdff dff_B_GlnTseJ03_0(.din(n568),.dout(w_dff_B_GlnTseJ03_0),.clk(gclk));
	jdff dff_B_ub5IZ7f08_0(.din(w_dff_B_GlnTseJ03_0),.dout(w_dff_B_ub5IZ7f08_0),.clk(gclk));
	jdff dff_B_hlze2NKO0_0(.din(w_dff_B_ub5IZ7f08_0),.dout(w_dff_B_hlze2NKO0_0),.clk(gclk));
	jdff dff_A_5C6bK9Er7_0(.dout(w_n567_0[0]),.din(w_dff_A_5C6bK9Er7_0),.clk(gclk));
	jdff dff_A_Mr9KwjKC5_0(.dout(w_dff_A_5C6bK9Er7_0),.din(w_dff_A_Mr9KwjKC5_0),.clk(gclk));
	jdff dff_A_qLDdam202_1(.dout(w_n554_3[1]),.din(w_dff_A_qLDdam202_1),.clk(gclk));
	jdff dff_A_Q4wI0UC29_1(.dout(w_dff_A_qLDdam202_1),.din(w_dff_A_Q4wI0UC29_1),.clk(gclk));
	jdff dff_A_VCWSou9t2_1(.dout(w_dff_A_Q4wI0UC29_1),.din(w_dff_A_VCWSou9t2_1),.clk(gclk));
	jdff dff_A_W2tZn6oo0_2(.dout(w_n554_3[2]),.din(w_dff_A_W2tZn6oo0_2),.clk(gclk));
	jdff dff_A_vZavnI3J3_2(.dout(w_dff_A_W2tZn6oo0_2),.din(w_dff_A_vZavnI3J3_2),.clk(gclk));
	jdff dff_A_21XGM9dY5_2(.dout(w_dff_A_vZavnI3J3_2),.din(w_dff_A_21XGM9dY5_2),.clk(gclk));
	jdff dff_B_DVg5wLGo7_2(.din(n565),.dout(w_dff_B_DVg5wLGo7_2),.clk(gclk));
	jdff dff_B_od8OPG3C2_2(.din(w_dff_B_DVg5wLGo7_2),.dout(w_dff_B_od8OPG3C2_2),.clk(gclk));
	jdff dff_B_XuZ320K68_2(.din(w_dff_B_od8OPG3C2_2),.dout(w_dff_B_XuZ320K68_2),.clk(gclk));
	jdff dff_B_qi5F0OtT9_2(.din(w_dff_B_XuZ320K68_2),.dout(w_dff_B_qi5F0OtT9_2),.clk(gclk));
	jdff dff_B_E8dVdOKK3_2(.din(w_dff_B_qi5F0OtT9_2),.dout(w_dff_B_E8dVdOKK3_2),.clk(gclk));
	jdff dff_B_GUthqoH39_2(.din(w_dff_B_E8dVdOKK3_2),.dout(w_dff_B_GUthqoH39_2),.clk(gclk));
	jdff dff_B_kv6xiJAF2_2(.din(w_dff_B_GUthqoH39_2),.dout(w_dff_B_kv6xiJAF2_2),.clk(gclk));
	jdff dff_B_4b2PzjOD8_2(.din(w_dff_B_kv6xiJAF2_2),.dout(w_dff_B_4b2PzjOD8_2),.clk(gclk));
	jdff dff_B_MXXFSrIR7_2(.din(w_dff_B_4b2PzjOD8_2),.dout(w_dff_B_MXXFSrIR7_2),.clk(gclk));
	jdff dff_B_awJynNY93_2(.din(w_dff_B_MXXFSrIR7_2),.dout(w_dff_B_awJynNY93_2),.clk(gclk));
	jdff dff_B_lKGVZogW8_2(.din(w_dff_B_awJynNY93_2),.dout(w_dff_B_lKGVZogW8_2),.clk(gclk));
	jdff dff_B_prryET5Y2_2(.din(w_dff_B_lKGVZogW8_2),.dout(w_dff_B_prryET5Y2_2),.clk(gclk));
	jdff dff_B_ixLNvbGt5_2(.din(w_dff_B_prryET5Y2_2),.dout(w_dff_B_ixLNvbGt5_2),.clk(gclk));
	jdff dff_A_h6FWygUN2_1(.dout(w_n1162_0[1]),.din(w_dff_A_h6FWygUN2_1),.clk(gclk));
	jdff dff_B_db7XWevs2_0(.din(n1161),.dout(w_dff_B_db7XWevs2_0),.clk(gclk));
	jdff dff_B_S5C3hmwv6_0(.din(w_dff_B_db7XWevs2_0),.dout(w_dff_B_S5C3hmwv6_0),.clk(gclk));
	jdff dff_B_9KNlN64E5_0(.din(n1158),.dout(w_dff_B_9KNlN64E5_0),.clk(gclk));
	jdff dff_B_grSwZci18_0(.din(w_dff_B_9KNlN64E5_0),.dout(w_dff_B_grSwZci18_0),.clk(gclk));
	jdff dff_B_YFXLITn83_0(.din(w_dff_B_grSwZci18_0),.dout(w_dff_B_YFXLITn83_0),.clk(gclk));
	jdff dff_B_c0lgAy7I6_0(.din(w_dff_B_YFXLITn83_0),.dout(w_dff_B_c0lgAy7I6_0),.clk(gclk));
	jdff dff_B_OnyCKrrI0_0(.din(w_dff_B_c0lgAy7I6_0),.dout(w_dff_B_OnyCKrrI0_0),.clk(gclk));
	jdff dff_B_Vmqt1nVN1_0(.din(n1157),.dout(w_dff_B_Vmqt1nVN1_0),.clk(gclk));
	jdff dff_B_emuLrLSO1_0(.din(w_dff_B_Vmqt1nVN1_0),.dout(w_dff_B_emuLrLSO1_0),.clk(gclk));
	jdff dff_B_G2gKboAY4_0(.din(n1155),.dout(w_dff_B_G2gKboAY4_0),.clk(gclk));
	jdff dff_B_ZCKLYel97_0(.din(w_dff_B_G2gKboAY4_0),.dout(w_dff_B_ZCKLYel97_0),.clk(gclk));
	jdff dff_B_T7YRSEFI8_1(.din(n1143),.dout(w_dff_B_T7YRSEFI8_1),.clk(gclk));
	jdff dff_B_nFwzypT18_1(.din(w_dff_B_T7YRSEFI8_1),.dout(w_dff_B_nFwzypT18_1),.clk(gclk));
	jdff dff_B_OlxLIZKe6_1(.din(n1145),.dout(w_dff_B_OlxLIZKe6_1),.clk(gclk));
	jdff dff_B_yCLnCPdg4_1(.din(n1148),.dout(w_dff_B_yCLnCPdg4_1),.clk(gclk));
	jdff dff_A_HHcohrtA2_1(.dout(w_n899_0[1]),.din(w_dff_A_HHcohrtA2_1),.clk(gclk));
	jdff dff_A_PhMWxTnj9_1(.dout(w_G87_1[1]),.din(w_dff_A_PhMWxTnj9_1),.clk(gclk));
	jdff dff_A_0IN0JfWw8_2(.dout(w_G87_1[2]),.din(w_dff_A_0IN0JfWw8_2),.clk(gclk));
	jdff dff_A_kFX52wfa6_1(.dout(w_G77_2[1]),.din(w_dff_A_kFX52wfa6_1),.clk(gclk));
	jdff dff_A_qOiP1xr63_1(.dout(w_dff_A_kFX52wfa6_1),.din(w_dff_A_qOiP1xr63_1),.clk(gclk));
	jdff dff_A_NlxxDMZS6_1(.dout(w_dff_A_qOiP1xr63_1),.din(w_dff_A_NlxxDMZS6_1),.clk(gclk));
	jdff dff_A_2qfylIWC6_1(.dout(w_dff_A_NlxxDMZS6_1),.din(w_dff_A_2qfylIWC6_1),.clk(gclk));
	jdff dff_A_FaEIrqfd4_2(.dout(w_G77_2[2]),.din(w_dff_A_FaEIrqfd4_2),.clk(gclk));
	jdff dff_A_RZ9Ybcvo7_2(.dout(w_dff_A_FaEIrqfd4_2),.din(w_dff_A_RZ9Ybcvo7_2),.clk(gclk));
	jdff dff_A_ai5X3qVU2_2(.dout(w_dff_A_RZ9Ybcvo7_2),.din(w_dff_A_ai5X3qVU2_2),.clk(gclk));
	jdff dff_A_k3RzfDcU5_2(.dout(w_dff_A_ai5X3qVU2_2),.din(w_dff_A_k3RzfDcU5_2),.clk(gclk));
	jdff dff_A_aX2enYOS0_1(.dout(w_G283_1[1]),.din(w_dff_A_aX2enYOS0_1),.clk(gclk));
	jdff dff_A_bMRvYAOp3_0(.dout(w_n148_3[0]),.din(w_dff_A_bMRvYAOp3_0),.clk(gclk));
	jdff dff_A_VOzgwAf71_0(.dout(w_dff_A_bMRvYAOp3_0),.din(w_dff_A_VOzgwAf71_0),.clk(gclk));
	jdff dff_A_f5eZqiSk3_0(.dout(w_dff_A_VOzgwAf71_0),.din(w_dff_A_f5eZqiSk3_0),.clk(gclk));
	jdff dff_A_7dahFntp7_0(.dout(w_dff_A_f5eZqiSk3_0),.din(w_dff_A_7dahFntp7_0),.clk(gclk));
	jdff dff_A_hCdCIPgc2_2(.dout(w_n148_3[2]),.din(w_dff_A_hCdCIPgc2_2),.clk(gclk));
	jdff dff_A_4mN2gque2_2(.dout(w_dff_A_hCdCIPgc2_2),.din(w_dff_A_4mN2gque2_2),.clk(gclk));
	jdff dff_A_dzJCSBPn5_2(.dout(w_dff_A_4mN2gque2_2),.din(w_dff_A_dzJCSBPn5_2),.clk(gclk));
	jdff dff_A_FGQPDyVV7_1(.dout(w_G294_1[1]),.din(w_dff_A_FGQPDyVV7_1),.clk(gclk));
	jdff dff_B_QIWtjCoA8_1(.din(n1128),.dout(w_dff_B_QIWtjCoA8_1),.clk(gclk));
	jdff dff_B_NeUMlFJp7_1(.din(n1130),.dout(w_dff_B_NeUMlFJp7_1),.clk(gclk));
	jdff dff_B_3i5y8pxZ4_1(.din(n1133),.dout(w_dff_B_3i5y8pxZ4_1),.clk(gclk));
	jdff dff_B_Pd0enkjG3_0(.din(n1134),.dout(w_dff_B_Pd0enkjG3_0),.clk(gclk));
	jdff dff_A_hNX5uZgb5_1(.dout(w_G150_1[1]),.din(w_dff_A_hNX5uZgb5_1),.clk(gclk));
	jdff dff_A_57GtZJ4n5_2(.dout(w_G150_1[2]),.din(w_dff_A_57GtZJ4n5_2),.clk(gclk));
	jdff dff_A_rM240p1f9_0(.dout(w_G128_0[0]),.din(w_dff_A_rM240p1f9_0),.clk(gclk));
	jdff dff_B_LpsyiCaf0_3(.din(G128),.dout(w_dff_B_LpsyiCaf0_3),.clk(gclk));
	jdff dff_B_MfiL7xzF9_3(.din(w_dff_B_LpsyiCaf0_3),.dout(w_dff_B_MfiL7xzF9_3),.clk(gclk));
	jdff dff_B_0VZex3Hm5_3(.din(w_dff_B_MfiL7xzF9_3),.dout(w_dff_B_0VZex3Hm5_3),.clk(gclk));
	jdff dff_B_HEvNRcaN0_1(.din(n1124),.dout(w_dff_B_HEvNRcaN0_1),.clk(gclk));
	jdff dff_B_7KXg4KOM0_0(.din(n1126),.dout(w_dff_B_7KXg4KOM0_0),.clk(gclk));
	jdff dff_A_oB6lzMDA6_0(.dout(w_n612_1[0]),.din(w_dff_A_oB6lzMDA6_0),.clk(gclk));
	jdff dff_A_j4Uv2WQa9_1(.dout(w_n612_1[1]),.din(w_dff_A_j4Uv2WQa9_1),.clk(gclk));
	jdff dff_A_hepERO6O0_1(.dout(w_dff_A_j4Uv2WQa9_1),.din(w_dff_A_hepERO6O0_1),.clk(gclk));
	jdff dff_A_EQNe65gU1_1(.dout(w_dff_A_hepERO6O0_1),.din(w_dff_A_EQNe65gU1_1),.clk(gclk));
	jdff dff_A_6nr5mi6s0_1(.dout(w_dff_A_EQNe65gU1_1),.din(w_dff_A_6nr5mi6s0_1),.clk(gclk));
	jdff dff_A_An8P9YTY1_1(.dout(w_dff_A_6nr5mi6s0_1),.din(w_dff_A_An8P9YTY1_1),.clk(gclk));
	jdff dff_A_FMuJZgSB0_1(.dout(w_dff_A_An8P9YTY1_1),.din(w_dff_A_FMuJZgSB0_1),.clk(gclk));
	jdff dff_A_AJINMCdz2_1(.dout(w_dff_A_FMuJZgSB0_1),.din(w_dff_A_AJINMCdz2_1),.clk(gclk));
	jdff dff_A_O8ofyVi79_1(.dout(w_n999_0[1]),.din(w_dff_A_O8ofyVi79_1),.clk(gclk));
	jdff dff_A_lNLgv9sO2_2(.dout(w_n764_0[2]),.din(w_dff_A_lNLgv9sO2_2),.clk(gclk));
	jdff dff_A_znYIGwJu5_2(.dout(w_dff_A_lNLgv9sO2_2),.din(w_dff_A_znYIGwJu5_2),.clk(gclk));
	jdff dff_B_dfYfCtd01_0(.din(n763),.dout(w_dff_B_dfYfCtd01_0),.clk(gclk));
	jdff dff_B_HDbb506a3_0(.din(w_dff_B_dfYfCtd01_0),.dout(w_dff_B_HDbb506a3_0),.clk(gclk));
	jdff dff_B_JEGIYvPq9_0(.din(n761),.dout(w_dff_B_JEGIYvPq9_0),.clk(gclk));
	jdff dff_B_2SXwo92r8_0(.din(w_dff_B_JEGIYvPq9_0),.dout(w_dff_B_2SXwo92r8_0),.clk(gclk));
	jdff dff_A_fk5jWGnA9_0(.dout(w_n760_0[0]),.din(w_dff_A_fk5jWGnA9_0),.clk(gclk));
	jdff dff_B_q0aTz60I1_0(.din(n997),.dout(w_dff_B_q0aTz60I1_0),.clk(gclk));
	jdff dff_B_dOt1Tn671_0(.din(w_dff_B_q0aTz60I1_0),.dout(w_dff_B_dOt1Tn671_0),.clk(gclk));
	jdff dff_B_aX6P7Wmo8_0(.din(w_dff_B_dOt1Tn671_0),.dout(w_dff_B_aX6P7Wmo8_0),.clk(gclk));
	jdff dff_B_Rk8nBEIU8_0(.din(w_dff_B_aX6P7Wmo8_0),.dout(w_dff_B_Rk8nBEIU8_0),.clk(gclk));
	jdff dff_B_LnzMSa2X5_0(.din(w_dff_B_Rk8nBEIU8_0),.dout(w_dff_B_LnzMSa2X5_0),.clk(gclk));
	jdff dff_A_SAJ9ZYRz3_2(.dout(w_n554_1[2]),.din(w_dff_A_SAJ9ZYRz3_2),.clk(gclk));
	jdff dff_A_sX2QTqjo1_1(.dout(w_n519_0[1]),.din(w_dff_A_sX2QTqjo1_1),.clk(gclk));
	jdff dff_A_08DYid1T7_1(.dout(w_dff_A_sX2QTqjo1_1),.din(w_dff_A_08DYid1T7_1),.clk(gclk));
	jdff dff_A_rUG6UDsZ7_2(.dout(w_n519_0[2]),.din(w_dff_A_rUG6UDsZ7_2),.clk(gclk));
	jdff dff_A_54pKiNtS3_2(.dout(w_dff_A_rUG6UDsZ7_2),.din(w_dff_A_54pKiNtS3_2),.clk(gclk));
	jdff dff_A_tzrtAI7m3_0(.dout(w_n548_0[0]),.din(w_dff_A_tzrtAI7m3_0),.clk(gclk));
	jdff dff_A_K7dgk8tN8_1(.dout(w_n439_0[1]),.din(w_dff_A_K7dgk8tN8_1),.clk(gclk));
	jdff dff_A_VGFuQtq12_1(.dout(w_dff_A_K7dgk8tN8_1),.din(w_dff_A_VGFuQtq12_1),.clk(gclk));
	jdff dff_A_iLZMufHi7_1(.dout(w_dff_A_VGFuQtq12_1),.din(w_dff_A_iLZMufHi7_1),.clk(gclk));
	jdff dff_A_jdrnQAet0_1(.dout(w_dff_A_iLZMufHi7_1),.din(w_dff_A_jdrnQAet0_1),.clk(gclk));
	jdff dff_B_RWpjDFmZ9_1(.din(n441),.dout(w_dff_B_RWpjDFmZ9_1),.clk(gclk));
	jdff dff_B_zINCodE96_1(.din(w_dff_B_RWpjDFmZ9_1),.dout(w_dff_B_zINCodE96_1),.clk(gclk));
	jdff dff_A_Omws4HRf0_1(.dout(w_n436_0[1]),.din(w_dff_A_Omws4HRf0_1),.clk(gclk));
	jdff dff_B_ofPosrps6_1(.din(n424),.dout(w_dff_B_ofPosrps6_1),.clk(gclk));
	jdff dff_B_GJ14VP5H9_0(.din(n434),.dout(w_dff_B_GJ14VP5H9_0),.clk(gclk));
	jdff dff_B_zFyNKBy09_0(.din(n423),.dout(w_dff_B_zFyNKBy09_0),.clk(gclk));
	jdff dff_B_aqhacGvo0_0(.din(w_dff_B_zFyNKBy09_0),.dout(w_dff_B_aqhacGvo0_0),.clk(gclk));
	jdff dff_B_gnYSGXxX9_1(.din(n413),.dout(w_dff_B_gnYSGXxX9_1),.clk(gclk));
	jdff dff_A_QYJ1XEN48_0(.dout(w_G226_1[0]),.din(w_dff_A_QYJ1XEN48_0),.clk(gclk));
	jdff dff_A_xhqleR399_0(.dout(w_dff_A_QYJ1XEN48_0),.din(w_dff_A_xhqleR399_0),.clk(gclk));
	jdff dff_B_Z9DRwtjf7_1(.din(n493),.dout(w_dff_B_Z9DRwtjf7_1),.clk(gclk));
	jdff dff_B_29U80Tha0_1(.din(w_dff_B_Z9DRwtjf7_1),.dout(w_dff_B_29U80Tha0_1),.clk(gclk));
	jdff dff_A_Svx1ceIm9_0(.dout(w_n516_0[0]),.din(w_dff_A_Svx1ceIm9_0),.clk(gclk));
	jdff dff_A_mDKt5XaW3_0(.dout(w_dff_A_Svx1ceIm9_0),.din(w_dff_A_mDKt5XaW3_0),.clk(gclk));
	jdff dff_B_ynRXNWFL6_0(.din(n514),.dout(w_dff_B_ynRXNWFL6_0),.clk(gclk));
	jdff dff_B_x12Dlwfq6_1(.din(n485),.dout(w_dff_B_x12Dlwfq6_1),.clk(gclk));
	jdff dff_B_kOs3fhSF4_1(.din(n496),.dout(w_dff_B_kOs3fhSF4_1),.clk(gclk));
	jdff dff_B_slMstrte5_1(.din(w_dff_B_kOs3fhSF4_1),.dout(w_dff_B_slMstrte5_1),.clk(gclk));
	jdff dff_B_cshKiaOQ2_1(.din(w_dff_B_slMstrte5_1),.dout(w_dff_B_cshKiaOQ2_1),.clk(gclk));
	jdff dff_B_zxbaoMfp4_0(.din(n505),.dout(w_dff_B_zxbaoMfp4_0),.clk(gclk));
	jdff dff_B_yOxgi82s2_0(.din(w_dff_B_zxbaoMfp4_0),.dout(w_dff_B_yOxgi82s2_0),.clk(gclk));
	jdff dff_B_VmG7eHiP2_1(.din(n497),.dout(w_dff_B_VmG7eHiP2_1),.clk(gclk));
	jdff dff_B_EPNAo89L3_1(.din(w_dff_B_VmG7eHiP2_1),.dout(w_dff_B_EPNAo89L3_1),.clk(gclk));
	jdff dff_B_B7COo6eY8_1(.din(w_dff_B_EPNAo89L3_1),.dout(w_dff_B_B7COo6eY8_1),.clk(gclk));
	jdff dff_A_ungVqv2X1_1(.dout(w_n541_0[1]),.din(w_dff_A_ungVqv2X1_1),.clk(gclk));
	jdff dff_A_C0LML8KC2_1(.dout(w_dff_A_ungVqv2X1_1),.din(w_dff_A_C0LML8KC2_1),.clk(gclk));
	jdff dff_B_d35W7zc98_1(.din(n456),.dout(w_dff_B_d35W7zc98_1),.clk(gclk));
	jdff dff_B_zWcwDe4Y2_1(.din(w_dff_B_d35W7zc98_1),.dout(w_dff_B_zWcwDe4Y2_1),.clk(gclk));
	jdff dff_A_lWlnWEgN4_0(.dout(w_n483_0[0]),.din(w_dff_A_lWlnWEgN4_0),.clk(gclk));
	jdff dff_A_Dqkbk04K2_0(.dout(w_dff_A_lWlnWEgN4_0),.din(w_dff_A_Dqkbk04K2_0),.clk(gclk));
	jdff dff_A_8FXxH05R3_0(.dout(w_dff_A_Dqkbk04K2_0),.din(w_dff_A_8FXxH05R3_0),.clk(gclk));
	jdff dff_A_umKsocQE8_0(.dout(w_dff_A_8FXxH05R3_0),.din(w_dff_A_umKsocQE8_0),.clk(gclk));
	jdff dff_B_npcdkGxv1_0(.din(n481),.dout(w_dff_B_npcdkGxv1_0),.clk(gclk));
	jdff dff_A_eQgjJxiJ5_1(.dout(w_G226_0[1]),.din(w_dff_A_eQgjJxiJ5_1),.clk(gclk));
	jdff dff_A_DGM43qRJ8_1(.dout(w_dff_A_eQgjJxiJ5_1),.din(w_dff_A_DGM43qRJ8_1),.clk(gclk));
	jdff dff_A_kTJVhsh78_2(.dout(w_G226_0[2]),.din(w_dff_A_kTJVhsh78_2),.clk(gclk));
	jdff dff_A_Mec99Jkt8_2(.dout(w_dff_A_kTJVhsh78_2),.din(w_dff_A_Mec99Jkt8_2),.clk(gclk));
	jdff dff_A_KhBqDzzW3_2(.dout(w_dff_A_Mec99Jkt8_2),.din(w_dff_A_KhBqDzzW3_2),.clk(gclk));
	jdff dff_A_fJlaCSEw5_2(.dout(w_dff_A_KhBqDzzW3_2),.din(w_dff_A_fJlaCSEw5_2),.clk(gclk));
	jdff dff_B_0Azvf9Fl7_1(.din(n448),.dout(w_dff_B_0Azvf9Fl7_1),.clk(gclk));
	jdff dff_B_ITbc963N6_1(.din(G222),.dout(w_dff_B_ITbc963N6_1),.clk(gclk));
	jdff dff_B_PRok0oYL4_1(.din(w_dff_B_ITbc963N6_1),.dout(w_dff_B_PRok0oYL4_1),.clk(gclk));
	jdff dff_A_cpviNkYV1_0(.dout(w_n430_0[0]),.din(w_dff_A_cpviNkYV1_0),.clk(gclk));
	jdff dff_B_Qrej3fvK6_2(.din(n430),.dout(w_dff_B_Qrej3fvK6_2),.clk(gclk));
	jdff dff_A_DYWWZoxZ8_1(.dout(w_G77_3[1]),.din(w_dff_A_DYWWZoxZ8_1),.clk(gclk));
	jdff dff_A_PqId0mA34_1(.dout(w_dff_A_DYWWZoxZ8_1),.din(w_dff_A_PqId0mA34_1),.clk(gclk));
	jdff dff_A_hIXBk1Sm1_1(.dout(w_dff_A_PqId0mA34_1),.din(w_dff_A_hIXBk1Sm1_1),.clk(gclk));
	jdff dff_B_jhsR9Bgj6_2(.din(G223),.dout(w_dff_B_jhsR9Bgj6_2),.clk(gclk));
	jdff dff_B_fru2YtIE1_2(.din(w_dff_B_jhsR9Bgj6_2),.dout(w_dff_B_fru2YtIE1_2),.clk(gclk));
	jdff dff_B_yiDorP7l7_1(.din(n459),.dout(w_dff_B_yiDorP7l7_1),.clk(gclk));
	jdff dff_B_OSnglj877_1(.din(w_dff_B_yiDorP7l7_1),.dout(w_dff_B_OSnglj877_1),.clk(gclk));
	jdff dff_B_Mpdsynv86_1(.din(w_dff_B_OSnglj877_1),.dout(w_dff_B_Mpdsynv86_1),.clk(gclk));
	jdff dff_B_Ar0CnoHU5_0(.din(n472),.dout(w_dff_B_Ar0CnoHU5_0),.clk(gclk));
	jdff dff_B_F9tTvFqz1_0(.din(w_dff_B_Ar0CnoHU5_0),.dout(w_dff_B_F9tTvFqz1_0),.clk(gclk));
	jdff dff_A_bHunUFF88_2(.dout(w_n185_1[2]),.din(w_dff_A_bHunUFF88_2),.clk(gclk));
	jdff dff_B_pHiKbyQ42_1(.din(n460),.dout(w_dff_B_pHiKbyQ42_1),.clk(gclk));
	jdff dff_B_dCHAiDYb7_1(.din(n461),.dout(w_dff_B_dCHAiDYb7_1),.clk(gclk));
	jdff dff_B_E8v5SAeS1_1(.din(w_dff_B_dCHAiDYb7_1),.dout(w_dff_B_E8v5SAeS1_1),.clk(gclk));
	jdff dff_A_PgdpENDr5_1(.dout(w_n75_0[1]),.din(w_dff_A_PgdpENDr5_1),.clk(gclk));
	jdff dff_A_9nFqy9n97_1(.dout(w_dff_A_PgdpENDr5_1),.din(w_dff_A_9nFqy9n97_1),.clk(gclk));
	jdff dff_A_H77SgCYr7_1(.dout(w_dff_A_9nFqy9n97_1),.din(w_dff_A_H77SgCYr7_1),.clk(gclk));
	jdff dff_A_64sbxD039_2(.dout(w_n75_0[2]),.din(w_dff_A_64sbxD039_2),.clk(gclk));
	jdff dff_A_FqNKuP124_2(.dout(w_dff_A_64sbxD039_2),.din(w_dff_A_FqNKuP124_2),.clk(gclk));
	jdff dff_A_6WVgIdG06_2(.dout(w_dff_A_FqNKuP124_2),.din(w_dff_A_6WVgIdG06_2),.clk(gclk));
	jdff dff_A_OvbUSvio9_2(.dout(w_dff_A_6WVgIdG06_2),.din(w_dff_A_OvbUSvio9_2),.clk(gclk));
	jdff dff_A_kxpL3vxm7_1(.dout(w_n74_0[1]),.din(w_dff_A_kxpL3vxm7_1),.clk(gclk));
	jdff dff_A_4KT7QmGz5_1(.dout(w_dff_A_kxpL3vxm7_1),.din(w_dff_A_4KT7QmGz5_1),.clk(gclk));
	jdff dff_A_3idra0BX3_1(.dout(w_dff_A_4KT7QmGz5_1),.din(w_dff_A_3idra0BX3_1),.clk(gclk));
	jdff dff_A_CuR1NTLR6_2(.dout(w_n74_0[2]),.din(w_dff_A_CuR1NTLR6_2),.clk(gclk));
	jdff dff_A_cHL9pHTy1_2(.dout(w_dff_A_CuR1NTLR6_2),.din(w_dff_A_cHL9pHTy1_2),.clk(gclk));
	jdff dff_A_IS82ssZ56_0(.dout(w_n73_2[0]),.din(w_dff_A_IS82ssZ56_0),.clk(gclk));
	jdff dff_A_vmV6BBVp7_0(.dout(w_dff_A_IS82ssZ56_0),.din(w_dff_A_vmV6BBVp7_0),.clk(gclk));
	jdff dff_A_w6X8EAcp6_2(.dout(w_n73_2[2]),.din(w_dff_A_w6X8EAcp6_2),.clk(gclk));
	jdff dff_A_6x8J0fqr0_2(.dout(w_n73_0[2]),.din(w_dff_A_6x8J0fqr0_2),.clk(gclk));
	jdff dff_A_kUor1Urz2_2(.dout(w_dff_A_6x8J0fqr0_2),.din(w_dff_A_kUor1Urz2_2),.clk(gclk));
	jdff dff_A_3meGaPFs8_2(.dout(w_dff_A_kUor1Urz2_2),.din(w_dff_A_3meGaPFs8_2),.clk(gclk));
	jdff dff_A_IMqtcTZr3_1(.dout(w_G50_5[1]),.din(w_dff_A_IMqtcTZr3_1),.clk(gclk));
	jdff dff_A_kNeAsqV88_1(.dout(w_dff_A_IMqtcTZr3_1),.din(w_dff_A_kNeAsqV88_1),.clk(gclk));
	jdff dff_A_RNGblkSf3_1(.dout(w_dff_A_kNeAsqV88_1),.din(w_dff_A_RNGblkSf3_1),.clk(gclk));
	jdff dff_A_LlrkQsaX4_0(.dout(w_G50_4[0]),.din(w_dff_A_LlrkQsaX4_0),.clk(gclk));
	jdff dff_A_fRSggduI5_0(.dout(w_dff_A_LlrkQsaX4_0),.din(w_dff_A_fRSggduI5_0),.clk(gclk));
	jdff dff_A_uDnNAuvx7_1(.dout(w_G50_4[1]),.din(w_dff_A_uDnNAuvx7_1),.clk(gclk));
	jdff dff_A_cO4jwKc07_0(.dout(w_G50_1[0]),.din(w_dff_A_cO4jwKc07_0),.clk(gclk));
	jdff dff_A_bX5NXgyS0_2(.dout(w_G50_1[2]),.din(w_dff_A_bX5NXgyS0_2),.clk(gclk));
	jdff dff_A_uVQZlh898_2(.dout(w_dff_A_bX5NXgyS0_2),.din(w_dff_A_uVQZlh898_2),.clk(gclk));
	jdff dff_A_Np93gKq95_2(.dout(w_dff_A_uVQZlh898_2),.din(w_dff_A_Np93gKq95_2),.clk(gclk));
	jdff dff_A_k3YJBcmu3_2(.dout(w_dff_A_Np93gKq95_2),.din(w_dff_A_k3YJBcmu3_2),.clk(gclk));
	jdff dff_A_IMewhTWL3_0(.dout(w_G384_0),.din(w_dff_A_IMewhTWL3_0),.clk(gclk));
	jdff dff_A_4vDcmayi0_0(.dout(w_dff_A_IMewhTWL3_0),.din(w_dff_A_4vDcmayi0_0),.clk(gclk));
	jdff dff_A_4WlSrDkw0_0(.dout(w_n750_0[0]),.din(w_dff_A_4WlSrDkw0_0),.clk(gclk));
	jdff dff_A_nU0xe2hO8_0(.dout(w_dff_A_4WlSrDkw0_0),.din(w_dff_A_nU0xe2hO8_0),.clk(gclk));
	jdff dff_B_nz0k8Dpq6_0(.din(n747),.dout(w_dff_B_nz0k8Dpq6_0),.clk(gclk));
	jdff dff_B_8OUHYnjW1_0(.din(w_dff_B_nz0k8Dpq6_0),.dout(w_dff_B_8OUHYnjW1_0),.clk(gclk));
	jdff dff_B_zcaO3fTP5_0(.din(w_dff_B_8OUHYnjW1_0),.dout(w_dff_B_zcaO3fTP5_0),.clk(gclk));
	jdff dff_B_Jm8RHGg78_0(.din(n746),.dout(w_dff_B_Jm8RHGg78_0),.clk(gclk));
	jdff dff_B_pEm7TDq81_0(.din(w_dff_B_Jm8RHGg78_0),.dout(w_dff_B_pEm7TDq81_0),.clk(gclk));
	jdff dff_B_dbbEQrdT0_0(.din(w_dff_B_pEm7TDq81_0),.dout(w_dff_B_dbbEQrdT0_0),.clk(gclk));
	jdff dff_B_RMjq1yaJ2_0(.din(w_dff_B_dbbEQrdT0_0),.dout(w_dff_B_RMjq1yaJ2_0),.clk(gclk));
	jdff dff_B_Df4TBVsa6_0(.din(n744),.dout(w_dff_B_Df4TBVsa6_0),.clk(gclk));
	jdff dff_B_zCZBW35C3_0(.din(w_dff_B_Df4TBVsa6_0),.dout(w_dff_B_zCZBW35C3_0),.clk(gclk));
	jdff dff_A_UnD3muEz2_2(.dout(w_n605_1[2]),.din(w_dff_A_UnD3muEz2_2),.clk(gclk));
	jdff dff_A_7DsqpNYG0_2(.dout(w_dff_A_UnD3muEz2_2),.din(w_dff_A_7DsqpNYG0_2),.clk(gclk));
	jdff dff_A_IwS5gG914_2(.dout(w_dff_A_7DsqpNYG0_2),.din(w_dff_A_IwS5gG914_2),.clk(gclk));
	jdff dff_A_GF8jmkDA1_2(.dout(w_dff_A_IwS5gG914_2),.din(w_dff_A_GF8jmkDA1_2),.clk(gclk));
	jdff dff_A_3EaRjSST1_2(.dout(w_dff_A_GF8jmkDA1_2),.din(w_dff_A_3EaRjSST1_2),.clk(gclk));
	jdff dff_A_V97YHEA45_2(.dout(w_dff_A_3EaRjSST1_2),.din(w_dff_A_V97YHEA45_2),.clk(gclk));
	jdff dff_A_0ufxqKr63_2(.dout(w_dff_A_V97YHEA45_2),.din(w_dff_A_0ufxqKr63_2),.clk(gclk));
	jdff dff_A_H2OdbD9J3_2(.dout(w_dff_A_0ufxqKr63_2),.din(w_dff_A_H2OdbD9J3_2),.clk(gclk));
	jdff dff_A_Aahst3tl4_0(.dout(w_n604_2[0]),.din(w_dff_A_Aahst3tl4_0),.clk(gclk));
	jdff dff_A_Lz1zNJb54_0(.dout(w_dff_A_Aahst3tl4_0),.din(w_dff_A_Lz1zNJb54_0),.clk(gclk));
	jdff dff_A_kwqkkcbr4_0(.dout(w_dff_A_Lz1zNJb54_0),.din(w_dff_A_kwqkkcbr4_0),.clk(gclk));
	jdff dff_A_id0GhgZb4_0(.dout(w_dff_A_kwqkkcbr4_0),.din(w_dff_A_id0GhgZb4_0),.clk(gclk));
	jdff dff_B_NU8ATwn54_1(.din(n721),.dout(w_dff_B_NU8ATwn54_1),.clk(gclk));
	jdff dff_B_C5aySXOr5_1(.din(w_dff_B_NU8ATwn54_1),.dout(w_dff_B_C5aySXOr5_1),.clk(gclk));
	jdff dff_B_yxqJN0WG9_1(.din(n727),.dout(w_dff_B_yxqJN0WG9_1),.clk(gclk));
	jdff dff_B_lcR5Qci74_1(.din(n730),.dout(w_dff_B_lcR5Qci74_1),.clk(gclk));
	jdff dff_B_cWpeFl2z9_1(.din(n733),.dout(w_dff_B_cWpeFl2z9_1),.clk(gclk));
	jdff dff_B_NRsKYzsN1_0(.din(n734),.dout(w_dff_B_NRsKYzsN1_0),.clk(gclk));
	jdff dff_A_PhvWA9S78_0(.dout(w_G294_2[0]),.din(w_dff_A_PhvWA9S78_0),.clk(gclk));
	jdff dff_A_QSc45vXT9_0(.dout(w_G116_3[0]),.din(w_dff_A_QSc45vXT9_0),.clk(gclk));
	jdff dff_A_epaqPPby9_0(.dout(w_dff_A_QSc45vXT9_0),.din(w_dff_A_epaqPPby9_0),.clk(gclk));
	jdff dff_A_ryAzrpiQ6_0(.dout(w_dff_A_epaqPPby9_0),.din(w_dff_A_ryAzrpiQ6_0),.clk(gclk));
	jdff dff_A_1OmPXXXf3_2(.dout(w_G116_3[2]),.din(w_dff_A_1OmPXXXf3_2),.clk(gclk));
	jdff dff_A_fd8aelqm7_2(.dout(w_dff_A_1OmPXXXf3_2),.din(w_dff_A_fd8aelqm7_2),.clk(gclk));
	jdff dff_A_cjnYpDZZ3_0(.dout(w_G33_5[0]),.din(w_dff_A_cjnYpDZZ3_0),.clk(gclk));
	jdff dff_A_hOC88yrv1_2(.dout(w_G33_5[2]),.din(w_dff_A_hOC88yrv1_2),.clk(gclk));
	jdff dff_A_S7K7j6zJ5_2(.dout(w_dff_A_hOC88yrv1_2),.din(w_dff_A_S7K7j6zJ5_2),.clk(gclk));
	jdff dff_B_F3OXA4Xb4_1(.din(n722),.dout(w_dff_B_F3OXA4Xb4_1),.clk(gclk));
	jdff dff_B_OhJl4kWT7_0(.din(n724),.dout(w_dff_B_OhJl4kWT7_0),.clk(gclk));
	jdff dff_A_XbIQ92Om5_1(.dout(w_G311_1[1]),.din(w_dff_A_XbIQ92Om5_1),.clk(gclk));
	jdff dff_B_rwito7iL8_3(.din(G311),.dout(w_dff_B_rwito7iL8_3),.clk(gclk));
	jdff dff_B_1HeEAX3R0_3(.din(w_dff_B_rwito7iL8_3),.dout(w_dff_B_1HeEAX3R0_3),.clk(gclk));
	jdff dff_B_dHAKO5Ky6_3(.din(w_dff_B_1HeEAX3R0_3),.dout(w_dff_B_dHAKO5Ky6_3),.clk(gclk));
	jdff dff_B_xjOizQFs3_1(.din(n710),.dout(w_dff_B_xjOizQFs3_1),.clk(gclk));
	jdff dff_B_uc1cmXy18_1(.din(n712),.dout(w_dff_B_uc1cmXy18_1),.clk(gclk));
	jdff dff_B_JdtGa10D5_1(.din(n715),.dout(w_dff_B_JdtGa10D5_1),.clk(gclk));
	jdff dff_B_OWwWer5e5_1(.din(n716),.dout(w_dff_B_OWwWer5e5_1),.clk(gclk));
	jdff dff_A_j6sSd1G47_1(.dout(w_G68_3[1]),.din(w_dff_A_j6sSd1G47_1),.clk(gclk));
	jdff dff_A_rPzBLQIM3_1(.dout(w_dff_A_j6sSd1G47_1),.din(w_dff_A_rPzBLQIM3_1),.clk(gclk));
	jdff dff_A_3ljWBAJk4_1(.dout(w_dff_A_rPzBLQIM3_1),.din(w_dff_A_3ljWBAJk4_1),.clk(gclk));
	jdff dff_A_KzTG18MI1_2(.dout(w_G68_3[2]),.din(w_dff_A_KzTG18MI1_2),.clk(gclk));
	jdff dff_A_YLSKHkFy7_2(.dout(w_dff_A_KzTG18MI1_2),.din(w_dff_A_YLSKHkFy7_2),.clk(gclk));
	jdff dff_A_qfTcccIv9_1(.dout(w_G137_1[1]),.din(w_dff_A_qfTcccIv9_1),.clk(gclk));
	jdff dff_B_QUDIr1v97_3(.din(G137),.dout(w_dff_B_QUDIr1v97_3),.clk(gclk));
	jdff dff_B_KNh74oeF5_3(.din(w_dff_B_QUDIr1v97_3),.dout(w_dff_B_KNh74oeF5_3),.clk(gclk));
	jdff dff_B_Q4pTqb6Z2_3(.din(w_dff_B_KNh74oeF5_3),.dout(w_dff_B_Q4pTqb6Z2_3),.clk(gclk));
	jdff dff_B_0Ak9n4Gf5_3(.din(G143),.dout(w_dff_B_0Ak9n4Gf5_3),.clk(gclk));
	jdff dff_B_ZT2Fy5OR0_3(.din(w_dff_B_0Ak9n4Gf5_3),.dout(w_dff_B_ZT2Fy5OR0_3),.clk(gclk));
	jdff dff_B_UfJBKIYt5_3(.din(w_dff_B_ZT2Fy5OR0_3),.dout(w_dff_B_UfJBKIYt5_3),.clk(gclk));
	jdff dff_A_D7VmnP0H6_0(.dout(w_G159_3[0]),.din(w_dff_A_D7VmnP0H6_0),.clk(gclk));
	jdff dff_A_VyqhLvL34_1(.dout(w_G159_3[1]),.din(w_dff_A_VyqhLvL34_1),.clk(gclk));
	jdff dff_A_ag9PAe2Q7_1(.dout(w_dff_A_VyqhLvL34_1),.din(w_dff_A_ag9PAe2Q7_1),.clk(gclk));
	jdff dff_A_2ISeGub15_0(.dout(w_G159_0[0]),.din(w_dff_A_2ISeGub15_0),.clk(gclk));
	jdff dff_A_pFsDiY7u2_0(.dout(w_dff_A_2ISeGub15_0),.din(w_dff_A_pFsDiY7u2_0),.clk(gclk));
	jdff dff_A_YFMzVTqr9_1(.dout(w_G159_0[1]),.din(w_dff_A_YFMzVTqr9_1),.clk(gclk));
	jdff dff_B_wpdkgUXj5_3(.din(G159),.dout(w_dff_B_wpdkgUXj5_3),.clk(gclk));
	jdff dff_B_qEsBJxUD4_3(.din(w_dff_B_wpdkgUXj5_3),.dout(w_dff_B_qEsBJxUD4_3),.clk(gclk));
	jdff dff_A_5QsPzIWS9_1(.dout(w_G190_2[1]),.din(w_dff_A_5QsPzIWS9_1),.clk(gclk));
	jdff dff_A_tbwDyGZi6_1(.dout(w_dff_A_5QsPzIWS9_1),.din(w_dff_A_tbwDyGZi6_1),.clk(gclk));
	jdff dff_A_I7En2C3i0_1(.dout(w_dff_A_tbwDyGZi6_1),.din(w_dff_A_I7En2C3i0_1),.clk(gclk));
	jdff dff_A_RkLGsPvh1_1(.dout(w_dff_A_I7En2C3i0_1),.din(w_dff_A_RkLGsPvh1_1),.clk(gclk));
	jdff dff_A_BzFwJUiJ7_1(.dout(w_dff_A_RkLGsPvh1_1),.din(w_dff_A_BzFwJUiJ7_1),.clk(gclk));
	jdff dff_A_zBquLsHA5_2(.dout(w_G190_2[2]),.din(w_dff_A_zBquLsHA5_2),.clk(gclk));
	jdff dff_A_l9kBWW3d9_2(.dout(w_dff_A_zBquLsHA5_2),.din(w_dff_A_l9kBWW3d9_2),.clk(gclk));
	jdff dff_A_G0SkIRPB5_2(.dout(w_dff_A_l9kBWW3d9_2),.din(w_dff_A_G0SkIRPB5_2),.clk(gclk));
	jdff dff_A_Nru9sjMX0_2(.dout(w_dff_A_G0SkIRPB5_2),.din(w_dff_A_Nru9sjMX0_2),.clk(gclk));
	jdff dff_A_O8MIMKtL8_2(.dout(w_dff_A_Nru9sjMX0_2),.din(w_dff_A_O8MIMKtL8_2),.clk(gclk));
	jdff dff_A_l2StL5735_0(.dout(w_G50_3[0]),.din(w_dff_A_l2StL5735_0),.clk(gclk));
	jdff dff_A_STYJgthL2_0(.dout(w_dff_A_l2StL5735_0),.din(w_dff_A_STYJgthL2_0),.clk(gclk));
	jdff dff_A_ViKm35nZ0_0(.dout(w_dff_A_STYJgthL2_0),.din(w_dff_A_ViKm35nZ0_0),.clk(gclk));
	jdff dff_A_6xd4p2ig0_2(.dout(w_G50_3[2]),.din(w_dff_A_6xd4p2ig0_2),.clk(gclk));
	jdff dff_A_YnW30gqB9_2(.dout(w_dff_A_6xd4p2ig0_2),.din(w_dff_A_YnW30gqB9_2),.clk(gclk));
	jdff dff_A_VTa9wZt32_2(.dout(w_dff_A_YnW30gqB9_2),.din(w_dff_A_VTa9wZt32_2),.clk(gclk));
	jdff dff_A_O3QSvosB8_2(.dout(w_dff_A_VTa9wZt32_2),.din(w_dff_A_O3QSvosB8_2),.clk(gclk));
	jdff dff_A_E4shbBiG7_1(.dout(w_G50_0[1]),.din(w_dff_A_E4shbBiG7_1),.clk(gclk));
	jdff dff_A_Ul7sozB86_1(.dout(w_dff_A_E4shbBiG7_1),.din(w_dff_A_Ul7sozB86_1),.clk(gclk));
	jdff dff_A_ceiHMDiR8_1(.dout(w_dff_A_Ul7sozB86_1),.din(w_dff_A_ceiHMDiR8_1),.clk(gclk));
	jdff dff_A_awF8wFPy0_0(.dout(w_G33_6[0]),.din(w_dff_A_awF8wFPy0_0),.clk(gclk));
	jdff dff_A_x1TuvTHU1_0(.dout(w_dff_A_awF8wFPy0_0),.din(w_dff_A_x1TuvTHU1_0),.clk(gclk));
	jdff dff_A_Vskg1MDg6_0(.dout(w_dff_A_x1TuvTHU1_0),.din(w_dff_A_Vskg1MDg6_0),.clk(gclk));
	jdff dff_A_vodn5zpv1_0(.dout(w_dff_A_Vskg1MDg6_0),.din(w_dff_A_vodn5zpv1_0),.clk(gclk));
	jdff dff_A_WTvG5u597_1(.dout(w_G33_6[1]),.din(w_dff_A_WTvG5u597_1),.clk(gclk));
	jdff dff_A_J9nVbyfr6_1(.dout(w_dff_A_WTvG5u597_1),.din(w_dff_A_J9nVbyfr6_1),.clk(gclk));
	jdff dff_A_MDmMMSEI6_1(.dout(w_G33_1[1]),.din(w_dff_A_MDmMMSEI6_1),.clk(gclk));
	jdff dff_A_nX47WIO03_1(.dout(w_dff_A_MDmMMSEI6_1),.din(w_dff_A_nX47WIO03_1),.clk(gclk));
	jdff dff_A_jyy5vK6a4_1(.dout(w_dff_A_nX47WIO03_1),.din(w_dff_A_jyy5vK6a4_1),.clk(gclk));
	jdff dff_B_qnbmHtnG0_1(.din(n706),.dout(w_dff_B_qnbmHtnG0_1),.clk(gclk));
	jdff dff_B_NxTT5afB0_0(.din(n708),.dout(w_dff_B_NxTT5afB0_0),.clk(gclk));
	jdff dff_A_SJzdCyfz2_0(.dout(w_G150_3[0]),.din(w_dff_A_SJzdCyfz2_0),.clk(gclk));
	jdff dff_A_Hf6WpMvU3_0(.dout(w_dff_A_SJzdCyfz2_0),.din(w_dff_A_Hf6WpMvU3_0),.clk(gclk));
	jdff dff_A_NYg96YUV4_0(.dout(w_dff_A_Hf6WpMvU3_0),.din(w_dff_A_NYg96YUV4_0),.clk(gclk));
	jdff dff_A_2jGD6EWq2_0(.dout(w_G150_0[0]),.din(w_dff_A_2jGD6EWq2_0),.clk(gclk));
	jdff dff_A_hsQkJUjs5_0(.dout(w_dff_A_2jGD6EWq2_0),.din(w_dff_A_hsQkJUjs5_0),.clk(gclk));
	jdff dff_A_99Lyr7EB8_0(.dout(w_dff_A_hsQkJUjs5_0),.din(w_dff_A_99Lyr7EB8_0),.clk(gclk));
	jdff dff_A_I1ysKMfU3_1(.dout(w_G150_0[1]),.din(w_dff_A_I1ysKMfU3_1),.clk(gclk));
	jdff dff_A_WuVLOwsN2_1(.dout(w_dff_A_I1ysKMfU3_1),.din(w_dff_A_WuVLOwsN2_1),.clk(gclk));
	jdff dff_A_KeaK6sWc8_1(.dout(w_dff_A_WuVLOwsN2_1),.din(w_dff_A_KeaK6sWc8_1),.clk(gclk));
	jdff dff_A_0J2BOCin4_0(.dout(w_G58_3[0]),.din(w_dff_A_0J2BOCin4_0),.clk(gclk));
	jdff dff_A_NfVWJxMP8_1(.dout(w_G58_3[1]),.din(w_dff_A_NfVWJxMP8_1),.clk(gclk));
	jdff dff_A_OFz0DY0G5_1(.dout(w_n615_0[1]),.din(w_dff_A_OFz0DY0G5_1),.clk(gclk));
	jdff dff_A_IygjiqAm7_1(.dout(w_G200_2[1]),.din(w_dff_A_IygjiqAm7_1),.clk(gclk));
	jdff dff_A_DjwTDdgY0_1(.dout(w_dff_A_IygjiqAm7_1),.din(w_dff_A_DjwTDdgY0_1),.clk(gclk));
	jdff dff_A_WbsNak8x0_1(.dout(w_dff_A_DjwTDdgY0_1),.din(w_dff_A_WbsNak8x0_1),.clk(gclk));
	jdff dff_A_Sr2PvNhv5_1(.dout(w_dff_A_WbsNak8x0_1),.din(w_dff_A_Sr2PvNhv5_1),.clk(gclk));
	jdff dff_A_zfneC0I78_1(.dout(w_dff_A_Sr2PvNhv5_1),.din(w_dff_A_zfneC0I78_1),.clk(gclk));
	jdff dff_A_nM2dE7mB2_1(.dout(w_dff_A_zfneC0I78_1),.din(w_dff_A_nM2dE7mB2_1),.clk(gclk));
	jdff dff_A_DgfAJj4N8_1(.dout(w_dff_A_nM2dE7mB2_1),.din(w_dff_A_DgfAJj4N8_1),.clk(gclk));
	jdff dff_A_wXWYsxiw2_2(.dout(w_G200_2[2]),.din(w_dff_A_wXWYsxiw2_2),.clk(gclk));
	jdff dff_A_haOV4gqD4_2(.dout(w_dff_A_wXWYsxiw2_2),.din(w_dff_A_haOV4gqD4_2),.clk(gclk));
	jdff dff_A_rWBDxUmw4_2(.dout(w_dff_A_haOV4gqD4_2),.din(w_dff_A_rWBDxUmw4_2),.clk(gclk));
	jdff dff_A_EvvZ3X4i9_2(.dout(w_dff_A_rWBDxUmw4_2),.din(w_dff_A_EvvZ3X4i9_2),.clk(gclk));
	jdff dff_A_rabhZ6A95_2(.dout(w_dff_A_EvvZ3X4i9_2),.din(w_dff_A_rabhZ6A95_2),.clk(gclk));
	jdff dff_A_GNYgQhL69_2(.dout(w_dff_A_rabhZ6A95_2),.din(w_dff_A_GNYgQhL69_2),.clk(gclk));
	jdff dff_A_9GwzyXxU8_2(.dout(w_dff_A_GNYgQhL69_2),.din(w_dff_A_9GwzyXxU8_2),.clk(gclk));
	jdff dff_A_5A63NY9a2_0(.dout(w_n619_0[0]),.din(w_dff_A_5A63NY9a2_0),.clk(gclk));
	jdff dff_A_QYNBuYWH1_0(.dout(w_n407_1[0]),.din(w_dff_A_QYNBuYWH1_0),.clk(gclk));
	jdff dff_A_uw12bGCa6_1(.dout(w_n407_1[1]),.din(w_dff_A_uw12bGCa6_1),.clk(gclk));
	jdff dff_A_aqXJWKtH7_1(.dout(w_dff_A_uw12bGCa6_1),.din(w_dff_A_aqXJWKtH7_1),.clk(gclk));
	jdff dff_A_hzAYjnOD2_1(.dout(w_G132_1[1]),.din(w_dff_A_hzAYjnOD2_1),.clk(gclk));
	jdff dff_B_qAclKrdA2_3(.din(G132),.dout(w_dff_B_qAclKrdA2_3),.clk(gclk));
	jdff dff_B_w3b5geSx4_3(.din(w_dff_B_qAclKrdA2_3),.dout(w_dff_B_w3b5geSx4_3),.clk(gclk));
	jdff dff_B_Fqzti0kV8_3(.din(w_dff_B_w3b5geSx4_3),.dout(w_dff_B_Fqzti0kV8_3),.clk(gclk));
	jdff dff_A_lntjXngU7_0(.dout(w_n612_3[0]),.din(w_dff_A_lntjXngU7_0),.clk(gclk));
	jdff dff_A_yPEQ2pZA0_0(.dout(w_dff_A_lntjXngU7_0),.din(w_dff_A_yPEQ2pZA0_0),.clk(gclk));
	jdff dff_A_HBZAUb3Z2_0(.dout(w_dff_A_yPEQ2pZA0_0),.din(w_dff_A_HBZAUb3Z2_0),.clk(gclk));
	jdff dff_A_0KOZ3ZLX5_0(.dout(w_dff_A_HBZAUb3Z2_0),.din(w_dff_A_0KOZ3ZLX5_0),.clk(gclk));
	jdff dff_A_0I2AnvN35_0(.dout(w_dff_A_0KOZ3ZLX5_0),.din(w_dff_A_0I2AnvN35_0),.clk(gclk));
	jdff dff_A_oY6PDkZN7_0(.dout(w_dff_A_0I2AnvN35_0),.din(w_dff_A_oY6PDkZN7_0),.clk(gclk));
	jdff dff_A_fMPXNQTL7_0(.dout(w_dff_A_oY6PDkZN7_0),.din(w_dff_A_fMPXNQTL7_0),.clk(gclk));
	jdff dff_A_vMAkBAe16_0(.dout(w_dff_A_fMPXNQTL7_0),.din(w_dff_A_vMAkBAe16_0),.clk(gclk));
	jdff dff_A_TD28eZi25_0(.dout(w_dff_A_vMAkBAe16_0),.din(w_dff_A_TD28eZi25_0),.clk(gclk));
	jdff dff_A_nejF3chI5_2(.dout(w_n612_3[2]),.din(w_dff_A_nejF3chI5_2),.clk(gclk));
	jdff dff_A_eG28GnkY8_2(.dout(w_dff_A_nejF3chI5_2),.din(w_dff_A_eG28GnkY8_2),.clk(gclk));
	jdff dff_A_Ys3imqdp0_2(.dout(w_dff_A_eG28GnkY8_2),.din(w_dff_A_Ys3imqdp0_2),.clk(gclk));
	jdff dff_A_m4UV112b5_2(.dout(w_dff_A_Ys3imqdp0_2),.din(w_dff_A_m4UV112b5_2),.clk(gclk));
	jdff dff_A_rXrpx5k01_2(.dout(w_dff_A_m4UV112b5_2),.din(w_dff_A_rXrpx5k01_2),.clk(gclk));
	jdff dff_A_96vV0G517_2(.dout(w_dff_A_rXrpx5k01_2),.din(w_dff_A_96vV0G517_2),.clk(gclk));
	jdff dff_A_nQN5faLv3_2(.dout(w_dff_A_96vV0G517_2),.din(w_dff_A_nQN5faLv3_2),.clk(gclk));
	jdff dff_A_dnxCFmOJ2_2(.dout(w_dff_A_nQN5faLv3_2),.din(w_dff_A_dnxCFmOJ2_2),.clk(gclk));
	jdff dff_A_TJa5PZqy0_2(.dout(w_dff_A_dnxCFmOJ2_2),.din(w_dff_A_TJa5PZqy0_2),.clk(gclk));
	jdff dff_A_tTKLcRNg1_1(.dout(w_n612_0[1]),.din(w_dff_A_tTKLcRNg1_1),.clk(gclk));
	jdff dff_A_VX52WHcy1_1(.dout(w_dff_A_tTKLcRNg1_1),.din(w_dff_A_VX52WHcy1_1),.clk(gclk));
	jdff dff_A_YxEwIlRF2_1(.dout(w_dff_A_VX52WHcy1_1),.din(w_dff_A_YxEwIlRF2_1),.clk(gclk));
	jdff dff_A_hZhPsBRS8_1(.dout(w_dff_A_YxEwIlRF2_1),.din(w_dff_A_hZhPsBRS8_1),.clk(gclk));
	jdff dff_A_WyR0C5My1_1(.dout(w_dff_A_hZhPsBRS8_1),.din(w_dff_A_WyR0C5My1_1),.clk(gclk));
	jdff dff_A_SKjdGmfI2_1(.dout(w_dff_A_WyR0C5My1_1),.din(w_dff_A_SKjdGmfI2_1),.clk(gclk));
	jdff dff_A_xYUjHr2C0_1(.dout(w_dff_A_SKjdGmfI2_1),.din(w_dff_A_xYUjHr2C0_1),.clk(gclk));
	jdff dff_A_hgHfYdiD1_1(.dout(w_n146_1[1]),.din(w_dff_A_hgHfYdiD1_1),.clk(gclk));
	jdff dff_A_uXbz31cQ1_1(.dout(w_dff_A_hgHfYdiD1_1),.din(w_dff_A_uXbz31cQ1_1),.clk(gclk));
	jdff dff_A_blrUEFU90_1(.dout(w_dff_A_uXbz31cQ1_1),.din(w_dff_A_blrUEFU90_1),.clk(gclk));
	jdff dff_A_jJGCuiG54_1(.dout(w_dff_A_blrUEFU90_1),.din(w_dff_A_jJGCuiG54_1),.clk(gclk));
	jdff dff_A_rk3LxFqX6_1(.dout(w_dff_A_jJGCuiG54_1),.din(w_dff_A_rk3LxFqX6_1),.clk(gclk));
	jdff dff_A_xTp5TZ9O0_1(.dout(w_dff_A_rk3LxFqX6_1),.din(w_dff_A_xTp5TZ9O0_1),.clk(gclk));
	jdff dff_A_XzxTgkJR1_2(.dout(w_n146_1[2]),.din(w_dff_A_XzxTgkJR1_2),.clk(gclk));
	jdff dff_A_maUJpcYL6_2(.dout(w_dff_A_XzxTgkJR1_2),.din(w_dff_A_maUJpcYL6_2),.clk(gclk));
	jdff dff_A_Y2tVyCbG7_2(.dout(w_dff_A_maUJpcYL6_2),.din(w_dff_A_Y2tVyCbG7_2),.clk(gclk));
	jdff dff_A_p7w6alMI1_2(.dout(w_dff_A_Y2tVyCbG7_2),.din(w_dff_A_p7w6alMI1_2),.clk(gclk));
	jdff dff_A_6pStX4yu2_2(.dout(w_dff_A_p7w6alMI1_2),.din(w_dff_A_6pStX4yu2_2),.clk(gclk));
	jdff dff_A_fzJDj07o3_2(.dout(w_dff_A_6pStX4yu2_2),.din(w_dff_A_fzJDj07o3_2),.clk(gclk));
	jdff dff_A_CwmetvLJ4_0(.dout(w_n425_1[0]),.din(w_dff_A_CwmetvLJ4_0),.clk(gclk));
	jdff dff_A_KMhfDZJK4_0(.dout(w_dff_A_CwmetvLJ4_0),.din(w_dff_A_KMhfDZJK4_0),.clk(gclk));
	jdff dff_A_xZOQaMZ18_0(.dout(w_dff_A_KMhfDZJK4_0),.din(w_dff_A_xZOQaMZ18_0),.clk(gclk));
	jdff dff_A_HIIdMCc72_0(.dout(w_dff_A_xZOQaMZ18_0),.din(w_dff_A_HIIdMCc72_0),.clk(gclk));
	jdff dff_A_DmgrzdGC2_0(.dout(w_dff_A_HIIdMCc72_0),.din(w_dff_A_DmgrzdGC2_0),.clk(gclk));
	jdff dff_A_4qaDxOO28_0(.dout(w_dff_A_DmgrzdGC2_0),.din(w_dff_A_4qaDxOO28_0),.clk(gclk));
	jdff dff_A_NYjhC4kM6_0(.dout(w_dff_A_4qaDxOO28_0),.din(w_dff_A_NYjhC4kM6_0),.clk(gclk));
	jdff dff_A_cMZDIVR50_0(.dout(w_dff_A_NYjhC4kM6_0),.din(w_dff_A_cMZDIVR50_0),.clk(gclk));
	jdff dff_A_yhKvvx4i3_0(.dout(w_dff_A_cMZDIVR50_0),.din(w_dff_A_yhKvvx4i3_0),.clk(gclk));
	jdff dff_A_aaG5i23a4_0(.dout(w_dff_A_yhKvvx4i3_0),.din(w_dff_A_aaG5i23a4_0),.clk(gclk));
	jdff dff_A_OU3GV55K4_0(.dout(w_dff_A_aaG5i23a4_0),.din(w_dff_A_OU3GV55K4_0),.clk(gclk));
	jdff dff_A_f05HXOnv4_0(.dout(w_dff_A_OU3GV55K4_0),.din(w_dff_A_f05HXOnv4_0),.clk(gclk));
	jdff dff_A_2tBscZ9S4_0(.dout(w_dff_A_f05HXOnv4_0),.din(w_dff_A_2tBscZ9S4_0),.clk(gclk));
	jdff dff_A_wY2BFypZ0_1(.dout(w_n425_1[1]),.din(w_dff_A_wY2BFypZ0_1),.clk(gclk));
	jdff dff_A_dpp6i8I67_1(.dout(w_dff_A_wY2BFypZ0_1),.din(w_dff_A_dpp6i8I67_1),.clk(gclk));
	jdff dff_A_IVvQ347e1_1(.dout(w_dff_A_dpp6i8I67_1),.din(w_dff_A_IVvQ347e1_1),.clk(gclk));
	jdff dff_A_cnVrDyCU7_1(.dout(w_dff_A_IVvQ347e1_1),.din(w_dff_A_cnVrDyCU7_1),.clk(gclk));
	jdff dff_A_8IVjR0xI3_1(.dout(w_dff_A_cnVrDyCU7_1),.din(w_dff_A_8IVjR0xI3_1),.clk(gclk));
	jdff dff_A_3Jxab8y11_1(.dout(w_dff_A_8IVjR0xI3_1),.din(w_dff_A_3Jxab8y11_1),.clk(gclk));
	jdff dff_A_uN7FRiqQ5_1(.dout(w_dff_A_3Jxab8y11_1),.din(w_dff_A_uN7FRiqQ5_1),.clk(gclk));
	jdff dff_A_gJrVJFWp4_1(.dout(w_dff_A_uN7FRiqQ5_1),.din(w_dff_A_gJrVJFWp4_1),.clk(gclk));
	jdff dff_A_2YLmKrwW2_1(.dout(w_dff_A_gJrVJFWp4_1),.din(w_dff_A_2YLmKrwW2_1),.clk(gclk));
	jdff dff_A_woculaxd1_1(.dout(w_dff_A_2YLmKrwW2_1),.din(w_dff_A_woculaxd1_1),.clk(gclk));
	jdff dff_A_BIxKP5jb2_1(.dout(w_dff_A_woculaxd1_1),.din(w_dff_A_BIxKP5jb2_1),.clk(gclk));
	jdff dff_A_gmUxuLte6_1(.dout(w_dff_A_BIxKP5jb2_1),.din(w_dff_A_gmUxuLte6_1),.clk(gclk));
	jdff dff_A_IVH6G14y3_1(.dout(w_dff_A_gmUxuLte6_1),.din(w_dff_A_IVH6G14y3_1),.clk(gclk));
	jdff dff_A_zULqCA694_1(.dout(w_n425_0[1]),.din(w_dff_A_zULqCA694_1),.clk(gclk));
	jdff dff_A_mOQ1Rf9X4_1(.dout(w_dff_A_zULqCA694_1),.din(w_dff_A_mOQ1Rf9X4_1),.clk(gclk));
	jdff dff_A_wMf7uVbY8_1(.dout(w_dff_A_mOQ1Rf9X4_1),.din(w_dff_A_wMf7uVbY8_1),.clk(gclk));
	jdff dff_A_X5uEQ9JW1_1(.dout(w_dff_A_wMf7uVbY8_1),.din(w_dff_A_X5uEQ9JW1_1),.clk(gclk));
	jdff dff_A_brqX0PSN0_1(.dout(w_dff_A_X5uEQ9JW1_1),.din(w_dff_A_brqX0PSN0_1),.clk(gclk));
	jdff dff_A_hzkHJ7Cn2_1(.dout(w_dff_A_brqX0PSN0_1),.din(w_dff_A_hzkHJ7Cn2_1),.clk(gclk));
	jdff dff_A_zwsVJ1Jd6_1(.dout(w_dff_A_hzkHJ7Cn2_1),.din(w_dff_A_zwsVJ1Jd6_1),.clk(gclk));
	jdff dff_A_QUlRRTAD9_1(.dout(w_dff_A_zwsVJ1Jd6_1),.din(w_dff_A_QUlRRTAD9_1),.clk(gclk));
	jdff dff_A_5r2OHNgV7_1(.dout(w_dff_A_QUlRRTAD9_1),.din(w_dff_A_5r2OHNgV7_1),.clk(gclk));
	jdff dff_A_cOX1wknL5_1(.dout(w_dff_A_5r2OHNgV7_1),.din(w_dff_A_cOX1wknL5_1),.clk(gclk));
	jdff dff_A_UBMxUog21_1(.dout(w_dff_A_cOX1wknL5_1),.din(w_dff_A_UBMxUog21_1),.clk(gclk));
	jdff dff_A_SBlFO4oN4_1(.dout(w_dff_A_UBMxUog21_1),.din(w_dff_A_SBlFO4oN4_1),.clk(gclk));
	jdff dff_A_Nog6MXY70_1(.dout(w_dff_A_SBlFO4oN4_1),.din(w_dff_A_Nog6MXY70_1),.clk(gclk));
	jdff dff_A_selQeCpb8_2(.dout(w_n425_0[2]),.din(w_dff_A_selQeCpb8_2),.clk(gclk));
	jdff dff_A_ZGjm3VWB7_2(.dout(w_dff_A_selQeCpb8_2),.din(w_dff_A_ZGjm3VWB7_2),.clk(gclk));
	jdff dff_A_wt1jgVp02_2(.dout(w_dff_A_ZGjm3VWB7_2),.din(w_dff_A_wt1jgVp02_2),.clk(gclk));
	jdff dff_A_dE4yIXIU6_2(.dout(w_dff_A_wt1jgVp02_2),.din(w_dff_A_dE4yIXIU6_2),.clk(gclk));
	jdff dff_A_aSLQIEMQ7_2(.dout(w_dff_A_dE4yIXIU6_2),.din(w_dff_A_aSLQIEMQ7_2),.clk(gclk));
	jdff dff_A_f8ZhtnEk9_2(.dout(w_dff_A_aSLQIEMQ7_2),.din(w_dff_A_f8ZhtnEk9_2),.clk(gclk));
	jdff dff_A_pZMcA2zf2_2(.dout(w_dff_A_f8ZhtnEk9_2),.din(w_dff_A_pZMcA2zf2_2),.clk(gclk));
	jdff dff_A_hcHaolDj0_2(.dout(w_dff_A_pZMcA2zf2_2),.din(w_dff_A_hcHaolDj0_2),.clk(gclk));
	jdff dff_A_3UsKYpRU8_2(.dout(w_dff_A_hcHaolDj0_2),.din(w_dff_A_3UsKYpRU8_2),.clk(gclk));
	jdff dff_A_auz1LV600_2(.dout(w_dff_A_3UsKYpRU8_2),.din(w_dff_A_auz1LV600_2),.clk(gclk));
	jdff dff_A_K8NbMXzY1_2(.dout(w_dff_A_auz1LV600_2),.din(w_dff_A_K8NbMXzY1_2),.clk(gclk));
	jdff dff_A_4oGrtiqL7_2(.dout(w_dff_A_K8NbMXzY1_2),.din(w_dff_A_4oGrtiqL7_2),.clk(gclk));
	jdff dff_A_n6eLtSK16_2(.dout(w_dff_A_4oGrtiqL7_2),.din(w_dff_A_n6eLtSK16_2),.clk(gclk));
	jdff dff_A_9Ris1djT8_0(.dout(w_n148_1[0]),.din(w_dff_A_9Ris1djT8_0),.clk(gclk));
	jdff dff_A_vAB9WeN85_0(.dout(w_dff_A_9Ris1djT8_0),.din(w_dff_A_vAB9WeN85_0),.clk(gclk));
	jdff dff_A_8oI67hMM8_0(.dout(w_dff_A_vAB9WeN85_0),.din(w_dff_A_8oI67hMM8_0),.clk(gclk));
	jdff dff_A_cRzoOTxt2_0(.dout(w_dff_A_8oI67hMM8_0),.din(w_dff_A_cRzoOTxt2_0),.clk(gclk));
	jdff dff_A_3FWaDXEN4_1(.dout(w_n148_1[1]),.din(w_dff_A_3FWaDXEN4_1),.clk(gclk));
	jdff dff_A_ch7PBlMN5_1(.dout(w_dff_A_3FWaDXEN4_1),.din(w_dff_A_ch7PBlMN5_1),.clk(gclk));
	jdff dff_B_nKnuInHT5_0(.din(n701),.dout(w_dff_B_nKnuInHT5_0),.clk(gclk));
	jdff dff_A_HFB9aPQp9_0(.dout(w_n604_1[0]),.din(w_dff_A_HFB9aPQp9_0),.clk(gclk));
	jdff dff_A_SYDBoXsz1_0(.dout(w_dff_A_HFB9aPQp9_0),.din(w_dff_A_SYDBoXsz1_0),.clk(gclk));
	jdff dff_A_Bg85DPP36_2(.dout(w_n604_1[2]),.din(w_dff_A_Bg85DPP36_2),.clk(gclk));
	jdff dff_A_qpTm1GQJ9_2(.dout(w_dff_A_Bg85DPP36_2),.din(w_dff_A_qpTm1GQJ9_2),.clk(gclk));
	jdff dff_A_SOoMbCl00_2(.dout(w_dff_A_qpTm1GQJ9_2),.din(w_dff_A_SOoMbCl00_2),.clk(gclk));
	jdff dff_A_jgbfN1vM5_2(.dout(w_dff_A_SOoMbCl00_2),.din(w_dff_A_jgbfN1vM5_2),.clk(gclk));
	jdff dff_A_EP4rSHyd8_2(.dout(w_dff_A_jgbfN1vM5_2),.din(w_dff_A_EP4rSHyd8_2),.clk(gclk));
	jdff dff_A_Ismp3crw7_2(.dout(w_dff_A_EP4rSHyd8_2),.din(w_dff_A_Ismp3crw7_2),.clk(gclk));
	jdff dff_A_ZNyGVDGL9_2(.dout(w_dff_A_Ismp3crw7_2),.din(w_dff_A_ZNyGVDGL9_2),.clk(gclk));
	jdff dff_A_nKyYHsfW0_2(.dout(w_dff_A_ZNyGVDGL9_2),.din(w_dff_A_nKyYHsfW0_2),.clk(gclk));
	jdff dff_A_FtLvesBI1_0(.dout(w_n604_0[0]),.din(w_dff_A_FtLvesBI1_0),.clk(gclk));
	jdff dff_A_ZrQMDoap6_0(.dout(w_dff_A_FtLvesBI1_0),.din(w_dff_A_ZrQMDoap6_0),.clk(gclk));
	jdff dff_A_bfes5KM11_2(.dout(w_n604_0[2]),.din(w_dff_A_bfes5KM11_2),.clk(gclk));
	jdff dff_A_GCtHfPh14_2(.dout(w_dff_A_bfes5KM11_2),.din(w_dff_A_GCtHfPh14_2),.clk(gclk));
	jdff dff_A_F4JM2YFm9_0(.dout(w_n603_2[0]),.din(w_dff_A_F4JM2YFm9_0),.clk(gclk));
	jdff dff_A_K84degn92_0(.dout(w_dff_A_F4JM2YFm9_0),.din(w_dff_A_K84degn92_0),.clk(gclk));
	jdff dff_A_nKuWQFIl5_0(.dout(w_dff_A_K84degn92_0),.din(w_dff_A_nKuWQFIl5_0),.clk(gclk));
	jdff dff_A_OIHgNgxR0_0(.dout(w_dff_A_nKuWQFIl5_0),.din(w_dff_A_OIHgNgxR0_0),.clk(gclk));
	jdff dff_A_Y2A7gShM2_0(.dout(w_dff_A_OIHgNgxR0_0),.din(w_dff_A_Y2A7gShM2_0),.clk(gclk));
	jdff dff_A_b50Re8nB5_0(.dout(w_dff_A_Y2A7gShM2_0),.din(w_dff_A_b50Re8nB5_0),.clk(gclk));
	jdff dff_A_e2VBHxhv5_0(.dout(w_dff_A_b50Re8nB5_0),.din(w_dff_A_e2VBHxhv5_0),.clk(gclk));
	jdff dff_A_0KIsQ1mU5_0(.dout(w_dff_A_e2VBHxhv5_0),.din(w_dff_A_0KIsQ1mU5_0),.clk(gclk));
	jdff dff_A_7oO9CIoC1_0(.dout(w_dff_A_0KIsQ1mU5_0),.din(w_dff_A_7oO9CIoC1_0),.clk(gclk));
	jdff dff_A_RSzZWXVj4_0(.dout(w_dff_A_7oO9CIoC1_0),.din(w_dff_A_RSzZWXVj4_0),.clk(gclk));
	jdff dff_A_rWmU1MjV1_0(.dout(w_dff_A_RSzZWXVj4_0),.din(w_dff_A_rWmU1MjV1_0),.clk(gclk));
	jdff dff_A_k1NkJp7b0_0(.dout(w_n603_0[0]),.din(w_dff_A_k1NkJp7b0_0),.clk(gclk));
	jdff dff_A_xtv4nyuw3_0(.dout(w_dff_A_k1NkJp7b0_0),.din(w_dff_A_xtv4nyuw3_0),.clk(gclk));
	jdff dff_A_YC8evA8F3_0(.dout(w_dff_A_xtv4nyuw3_0),.din(w_dff_A_YC8evA8F3_0),.clk(gclk));
	jdff dff_A_Ok1a3AvL2_0(.dout(w_dff_A_YC8evA8F3_0),.din(w_dff_A_Ok1a3AvL2_0),.clk(gclk));
	jdff dff_A_R18cgiXf1_0(.dout(w_dff_A_Ok1a3AvL2_0),.din(w_dff_A_R18cgiXf1_0),.clk(gclk));
	jdff dff_A_4LeNu4Fx5_0(.dout(w_dff_A_R18cgiXf1_0),.din(w_dff_A_4LeNu4Fx5_0),.clk(gclk));
	jdff dff_A_goZeSfFy0_0(.dout(w_dff_A_4LeNu4Fx5_0),.din(w_dff_A_goZeSfFy0_0),.clk(gclk));
	jdff dff_A_7ufrZGyP7_0(.dout(w_dff_A_goZeSfFy0_0),.din(w_dff_A_7ufrZGyP7_0),.clk(gclk));
	jdff dff_A_9zjWDTx27_0(.dout(w_dff_A_7ufrZGyP7_0),.din(w_dff_A_9zjWDTx27_0),.clk(gclk));
	jdff dff_A_A3zbijFr1_0(.dout(w_dff_A_9zjWDTx27_0),.din(w_dff_A_A3zbijFr1_0),.clk(gclk));
	jdff dff_A_Rvoneyhf2_0(.dout(w_dff_A_A3zbijFr1_0),.din(w_dff_A_Rvoneyhf2_0),.clk(gclk));
	jdff dff_A_sefXaNOh3_0(.dout(w_dff_A_Rvoneyhf2_0),.din(w_dff_A_sefXaNOh3_0),.clk(gclk));
	jdff dff_A_7GWS8WTE9_0(.dout(w_dff_A_sefXaNOh3_0),.din(w_dff_A_7GWS8WTE9_0),.clk(gclk));
	jdff dff_A_5a96gD1R9_0(.dout(w_dff_A_7GWS8WTE9_0),.din(w_dff_A_5a96gD1R9_0),.clk(gclk));
	jdff dff_A_E57cqyLp5_2(.dout(w_n603_0[2]),.din(w_dff_A_E57cqyLp5_2),.clk(gclk));
	jdff dff_A_3djHRfyX3_2(.dout(w_dff_A_E57cqyLp5_2),.din(w_dff_A_3djHRfyX3_2),.clk(gclk));
	jdff dff_A_anl4YDs76_2(.dout(w_dff_A_3djHRfyX3_2),.din(w_dff_A_anl4YDs76_2),.clk(gclk));
	jdff dff_A_Mfi644JQ0_2(.dout(w_dff_A_anl4YDs76_2),.din(w_dff_A_Mfi644JQ0_2),.clk(gclk));
	jdff dff_A_BKiHM41L6_2(.dout(w_dff_A_Mfi644JQ0_2),.din(w_dff_A_BKiHM41L6_2),.clk(gclk));
	jdff dff_A_jwf3RqY31_2(.dout(w_dff_A_BKiHM41L6_2),.din(w_dff_A_jwf3RqY31_2),.clk(gclk));
	jdff dff_A_s0qAwI177_2(.dout(w_dff_A_jwf3RqY31_2),.din(w_dff_A_s0qAwI177_2),.clk(gclk));
	jdff dff_A_shISe07W1_2(.dout(w_dff_A_s0qAwI177_2),.din(w_dff_A_shISe07W1_2),.clk(gclk));
	jdff dff_A_timhTuNW9_2(.dout(w_dff_A_shISe07W1_2),.din(w_dff_A_timhTuNW9_2),.clk(gclk));
	jdff dff_A_XgT1hNsl5_2(.dout(w_dff_A_timhTuNW9_2),.din(w_dff_A_XgT1hNsl5_2),.clk(gclk));
	jdff dff_A_6FBUvdrw1_2(.dout(w_dff_A_XgT1hNsl5_2),.din(w_dff_A_6FBUvdrw1_2),.clk(gclk));
	jdff dff_A_s6e0nStv1_2(.dout(w_dff_A_6FBUvdrw1_2),.din(w_dff_A_s6e0nStv1_2),.clk(gclk));
	jdff dff_A_G1RDL8658_2(.dout(w_dff_A_s6e0nStv1_2),.din(w_dff_A_G1RDL8658_2),.clk(gclk));
	jdff dff_A_XXvBEiAi5_0(.dout(w_n602_0[0]),.din(w_dff_A_XXvBEiAi5_0),.clk(gclk));
	jdff dff_A_RDrg7y4S0_0(.dout(w_dff_A_XXvBEiAi5_0),.din(w_dff_A_RDrg7y4S0_0),.clk(gclk));
	jdff dff_A_f9Cpt51i1_0(.dout(w_dff_A_RDrg7y4S0_0),.din(w_dff_A_f9Cpt51i1_0),.clk(gclk));
	jdff dff_A_cPKpNQWS6_0(.dout(w_dff_A_f9Cpt51i1_0),.din(w_dff_A_cPKpNQWS6_0),.clk(gclk));
	jdff dff_A_7hcUo6Fw6_0(.dout(w_dff_A_cPKpNQWS6_0),.din(w_dff_A_7hcUo6Fw6_0),.clk(gclk));
	jdff dff_A_4l2dCGDJ4_0(.dout(w_dff_A_7hcUo6Fw6_0),.din(w_dff_A_4l2dCGDJ4_0),.clk(gclk));
	jdff dff_A_DwmwnVAX6_0(.dout(w_dff_A_4l2dCGDJ4_0),.din(w_dff_A_DwmwnVAX6_0),.clk(gclk));
	jdff dff_A_YoxkjmP48_0(.dout(w_dff_A_DwmwnVAX6_0),.din(w_dff_A_YoxkjmP48_0),.clk(gclk));
	jdff dff_A_EOKouaho4_0(.dout(w_dff_A_YoxkjmP48_0),.din(w_dff_A_EOKouaho4_0),.clk(gclk));
	jdff dff_A_PBhybKyN1_0(.dout(w_dff_A_EOKouaho4_0),.din(w_dff_A_PBhybKyN1_0),.clk(gclk));
	jdff dff_A_ZvsNFf2l9_0(.dout(w_dff_A_PBhybKyN1_0),.din(w_dff_A_ZvsNFf2l9_0),.clk(gclk));
	jdff dff_A_5O6qQtgB8_0(.dout(w_dff_A_ZvsNFf2l9_0),.din(w_dff_A_5O6qQtgB8_0),.clk(gclk));
	jdff dff_A_7cPgEucv5_0(.dout(w_dff_A_5O6qQtgB8_0),.din(w_dff_A_7cPgEucv5_0),.clk(gclk));
	jdff dff_A_ixKVzI3j3_0(.dout(w_dff_A_7cPgEucv5_0),.din(w_dff_A_ixKVzI3j3_0),.clk(gclk));
	jdff dff_A_6h4ZecNt6_0(.dout(w_dff_A_ixKVzI3j3_0),.din(w_dff_A_6h4ZecNt6_0),.clk(gclk));
	jdff dff_A_w0tPuwmj0_0(.dout(w_dff_A_6h4ZecNt6_0),.din(w_dff_A_w0tPuwmj0_0),.clk(gclk));
	jdff dff_A_8ZO8nfsg0_0(.dout(w_dff_A_w0tPuwmj0_0),.din(w_dff_A_8ZO8nfsg0_0),.clk(gclk));
	jdff dff_A_5NHNfACy9_0(.dout(w_n592_0[0]),.din(w_dff_A_5NHNfACy9_0),.clk(gclk));
	jdff dff_A_G18Mxl004_0(.dout(w_dff_A_5NHNfACy9_0),.din(w_dff_A_G18Mxl004_0),.clk(gclk));
	jdff dff_A_usf1N4f43_0(.dout(w_dff_A_G18Mxl004_0),.din(w_dff_A_usf1N4f43_0),.clk(gclk));
	jdff dff_A_KNfKET0q1_0(.dout(w_dff_A_usf1N4f43_0),.din(w_dff_A_KNfKET0q1_0),.clk(gclk));
	jdff dff_A_kz1yxDR71_0(.dout(w_dff_A_KNfKET0q1_0),.din(w_dff_A_kz1yxDR71_0),.clk(gclk));
	jdff dff_A_LHxeaux42_0(.dout(w_dff_A_kz1yxDR71_0),.din(w_dff_A_LHxeaux42_0),.clk(gclk));
	jdff dff_A_5sTCyrqc9_0(.dout(w_dff_A_LHxeaux42_0),.din(w_dff_A_5sTCyrqc9_0),.clk(gclk));
	jdff dff_A_FX7F36bV1_0(.dout(w_dff_A_5sTCyrqc9_0),.din(w_dff_A_FX7F36bV1_0),.clk(gclk));
	jdff dff_A_aCotgp3k1_0(.dout(w_dff_A_FX7F36bV1_0),.din(w_dff_A_aCotgp3k1_0),.clk(gclk));
	jdff dff_A_hkReL28n0_0(.dout(w_dff_A_aCotgp3k1_0),.din(w_dff_A_hkReL28n0_0),.clk(gclk));
	jdff dff_A_d30irgnH5_0(.dout(w_dff_A_hkReL28n0_0),.din(w_dff_A_d30irgnH5_0),.clk(gclk));
	jdff dff_A_rzjd6yL58_0(.dout(w_dff_A_d30irgnH5_0),.din(w_dff_A_rzjd6yL58_0),.clk(gclk));
	jdff dff_A_XVsKrCdE7_0(.dout(w_dff_A_rzjd6yL58_0),.din(w_dff_A_XVsKrCdE7_0),.clk(gclk));
	jdff dff_A_eFeoRqT64_2(.dout(w_n592_0[2]),.din(w_dff_A_eFeoRqT64_2),.clk(gclk));
	jdff dff_A_n66LXlKa5_2(.dout(w_dff_A_eFeoRqT64_2),.din(w_dff_A_n66LXlKa5_2),.clk(gclk));
	jdff dff_A_4tE8wuxC2_2(.dout(w_dff_A_n66LXlKa5_2),.din(w_dff_A_4tE8wuxC2_2),.clk(gclk));
	jdff dff_A_7K543ZXj6_2(.dout(w_dff_A_4tE8wuxC2_2),.din(w_dff_A_7K543ZXj6_2),.clk(gclk));
	jdff dff_A_ucrzRESH3_2(.dout(w_dff_A_7K543ZXj6_2),.din(w_dff_A_ucrzRESH3_2),.clk(gclk));
	jdff dff_A_7HADqwTF6_2(.dout(w_dff_A_ucrzRESH3_2),.din(w_dff_A_7HADqwTF6_2),.clk(gclk));
	jdff dff_A_8EGHPGrd4_2(.dout(w_dff_A_7HADqwTF6_2),.din(w_dff_A_8EGHPGrd4_2),.clk(gclk));
	jdff dff_A_U3Hu6lUw8_2(.dout(w_dff_A_8EGHPGrd4_2),.din(w_dff_A_U3Hu6lUw8_2),.clk(gclk));
	jdff dff_A_rkloMUJm8_2(.dout(w_dff_A_U3Hu6lUw8_2),.din(w_dff_A_rkloMUJm8_2),.clk(gclk));
	jdff dff_A_DxSbFAvt0_2(.dout(w_dff_A_rkloMUJm8_2),.din(w_dff_A_DxSbFAvt0_2),.clk(gclk));
	jdff dff_A_ss6FeutD6_2(.dout(w_dff_A_DxSbFAvt0_2),.din(w_dff_A_ss6FeutD6_2),.clk(gclk));
	jdff dff_A_dZdSFfP14_2(.dout(w_dff_A_ss6FeutD6_2),.din(w_dff_A_dZdSFfP14_2),.clk(gclk));
	jdff dff_A_VLQxYgqR3_2(.dout(w_dff_A_dZdSFfP14_2),.din(w_dff_A_VLQxYgqR3_2),.clk(gclk));
	jdff dff_A_S7M87JQ34_2(.dout(w_dff_A_VLQxYgqR3_2),.din(w_dff_A_S7M87JQ34_2),.clk(gclk));
	jdff dff_A_9bEojj280_2(.dout(w_dff_A_S7M87JQ34_2),.din(w_dff_A_9bEojj280_2),.clk(gclk));
	jdff dff_A_8uzhtFKJ3_2(.dout(w_dff_A_9bEojj280_2),.din(w_dff_A_8uzhtFKJ3_2),.clk(gclk));
	jdff dff_A_CpoKBqtE8_1(.dout(w_n591_0[1]),.din(w_dff_A_CpoKBqtE8_1),.clk(gclk));
	jdff dff_A_p1EYyQHN3_1(.dout(w_dff_A_CpoKBqtE8_1),.din(w_dff_A_p1EYyQHN3_1),.clk(gclk));
	jdff dff_A_JLk0Odgx0_1(.dout(w_dff_A_p1EYyQHN3_1),.din(w_dff_A_JLk0Odgx0_1),.clk(gclk));
	jdff dff_A_YCOGnO5v7_1(.dout(w_dff_A_JLk0Odgx0_1),.din(w_dff_A_YCOGnO5v7_1),.clk(gclk));
	jdff dff_A_HFqTF5Yr7_1(.dout(w_dff_A_YCOGnO5v7_1),.din(w_dff_A_HFqTF5Yr7_1),.clk(gclk));
	jdff dff_A_ZIn8C9WS7_1(.dout(w_dff_A_HFqTF5Yr7_1),.din(w_dff_A_ZIn8C9WS7_1),.clk(gclk));
	jdff dff_A_oisPxduo3_1(.dout(w_dff_A_ZIn8C9WS7_1),.din(w_dff_A_oisPxduo3_1),.clk(gclk));
	jdff dff_A_VZRWOjUT8_1(.dout(w_dff_A_oisPxduo3_1),.din(w_dff_A_VZRWOjUT8_1),.clk(gclk));
	jdff dff_A_cMAy5yxu0_1(.dout(w_dff_A_VZRWOjUT8_1),.din(w_dff_A_cMAy5yxu0_1),.clk(gclk));
	jdff dff_A_f3400uJP9_1(.dout(w_dff_A_cMAy5yxu0_1),.din(w_dff_A_f3400uJP9_1),.clk(gclk));
	jdff dff_A_URtKe4Ir6_1(.dout(w_dff_A_f3400uJP9_1),.din(w_dff_A_URtKe4Ir6_1),.clk(gclk));
	jdff dff_A_SNlLy2Sr3_1(.dout(w_dff_A_URtKe4Ir6_1),.din(w_dff_A_SNlLy2Sr3_1),.clk(gclk));
	jdff dff_A_Zj24YKqJ9_1(.dout(w_dff_A_SNlLy2Sr3_1),.din(w_dff_A_Zj24YKqJ9_1),.clk(gclk));
	jdff dff_A_mLacGsv77_1(.dout(w_dff_A_Zj24YKqJ9_1),.din(w_dff_A_mLacGsv77_1),.clk(gclk));
	jdff dff_A_JNRB8m2A6_1(.dout(w_dff_A_mLacGsv77_1),.din(w_dff_A_JNRB8m2A6_1),.clk(gclk));
	jdff dff_A_yvJ5Qhd01_2(.dout(w_n591_0[2]),.din(w_dff_A_yvJ5Qhd01_2),.clk(gclk));
	jdff dff_A_eHn2MEGk4_2(.dout(w_dff_A_yvJ5Qhd01_2),.din(w_dff_A_eHn2MEGk4_2),.clk(gclk));
	jdff dff_A_EYMn6Bug8_2(.dout(w_dff_A_eHn2MEGk4_2),.din(w_dff_A_EYMn6Bug8_2),.clk(gclk));
	jdff dff_A_MyUmvZKc4_2(.dout(w_dff_A_EYMn6Bug8_2),.din(w_dff_A_MyUmvZKc4_2),.clk(gclk));
	jdff dff_A_wsQ58IRP9_2(.dout(w_dff_A_MyUmvZKc4_2),.din(w_dff_A_wsQ58IRP9_2),.clk(gclk));
	jdff dff_A_LMtJko6c3_2(.dout(w_dff_A_wsQ58IRP9_2),.din(w_dff_A_LMtJko6c3_2),.clk(gclk));
	jdff dff_A_FCIy9CXr2_2(.dout(w_dff_A_LMtJko6c3_2),.din(w_dff_A_FCIy9CXr2_2),.clk(gclk));
	jdff dff_A_CyvMBjUf4_2(.dout(w_dff_A_FCIy9CXr2_2),.din(w_dff_A_CyvMBjUf4_2),.clk(gclk));
	jdff dff_A_sSQQ3S9O4_2(.dout(w_dff_A_CyvMBjUf4_2),.din(w_dff_A_sSQQ3S9O4_2),.clk(gclk));
	jdff dff_A_kXLpwcdx6_2(.dout(w_dff_A_sSQQ3S9O4_2),.din(w_dff_A_kXLpwcdx6_2),.clk(gclk));
	jdff dff_A_vjqMPCmp1_2(.dout(w_dff_A_kXLpwcdx6_2),.din(w_dff_A_vjqMPCmp1_2),.clk(gclk));
	jdff dff_A_Kziu9Gxh6_2(.dout(w_dff_A_vjqMPCmp1_2),.din(w_dff_A_Kziu9Gxh6_2),.clk(gclk));
	jdff dff_A_u9j690ft2_2(.dout(w_dff_A_Kziu9Gxh6_2),.din(w_dff_A_u9j690ft2_2),.clk(gclk));
	jdff dff_A_dXO5iyXF3_2(.dout(w_dff_A_u9j690ft2_2),.din(w_dff_A_dXO5iyXF3_2),.clk(gclk));
	jdff dff_A_eK5Mpd8I8_2(.dout(w_dff_A_dXO5iyXF3_2),.din(w_dff_A_eK5Mpd8I8_2),.clk(gclk));
	jdff dff_A_2rQ3bUW76_2(.dout(w_dff_A_eK5Mpd8I8_2),.din(w_dff_A_2rQ3bUW76_2),.clk(gclk));
	jdff dff_A_ccXMLJM11_0(.dout(w_n121_0[0]),.din(w_dff_A_ccXMLJM11_0),.clk(gclk));
	jdff dff_B_RGswLtgJ5_1(.din(n690),.dout(w_dff_B_RGswLtgJ5_1),.clk(gclk));
	jdff dff_A_TGkm35os1_0(.dout(w_n696_1[0]),.din(w_dff_A_TGkm35os1_0),.clk(gclk));
	jdff dff_A_Z5GVPtXq1_2(.dout(w_n696_1[2]),.din(w_dff_A_Z5GVPtXq1_2),.clk(gclk));
	jdff dff_A_aeOguVQ19_1(.dout(w_n696_0[1]),.din(w_dff_A_aeOguVQ19_1),.clk(gclk));
	jdff dff_A_bc0Bi0ZA8_1(.dout(w_n692_0[1]),.din(w_dff_A_bc0Bi0ZA8_1),.clk(gclk));
	jdff dff_B_X3IijG2u6_2(.din(n692),.dout(w_dff_B_X3IijG2u6_2),.clk(gclk));
	jdff dff_B_SfXOQchI0_1(.din(n406),.dout(w_dff_B_SfXOQchI0_1),.clk(gclk));
	jdff dff_B_NL5dvISo6_1(.din(w_dff_B_SfXOQchI0_1),.dout(w_dff_B_NL5dvISo6_1),.clk(gclk));
	jdff dff_A_pQUuYADs3_1(.dout(w_n407_0[1]),.din(w_dff_A_pQUuYADs3_1),.clk(gclk));
	jdff dff_A_sTeDeewm0_1(.dout(w_dff_A_pQUuYADs3_1),.din(w_dff_A_sTeDeewm0_1),.clk(gclk));
	jdff dff_A_vPBdSlVK8_1(.dout(w_dff_A_sTeDeewm0_1),.din(w_dff_A_vPBdSlVK8_1),.clk(gclk));
	jdff dff_A_93WQQBLH2_1(.dout(w_dff_A_vPBdSlVK8_1),.din(w_dff_A_93WQQBLH2_1),.clk(gclk));
	jdff dff_A_abu25aDs1_1(.dout(w_dff_A_93WQQBLH2_1),.din(w_dff_A_abu25aDs1_1),.clk(gclk));
	jdff dff_A_RstvUsjn8_1(.dout(w_dff_A_abu25aDs1_1),.din(w_dff_A_RstvUsjn8_1),.clk(gclk));
	jdff dff_A_OUBqBLoT3_2(.dout(w_n407_0[2]),.din(w_dff_A_OUBqBLoT3_2),.clk(gclk));
	jdff dff_A_ZIQFC32R1_1(.dout(w_n401_0[1]),.din(w_dff_A_ZIQFC32R1_1),.clk(gclk));
	jdff dff_B_63h7EG696_1(.din(n396),.dout(w_dff_B_63h7EG696_1),.clk(gclk));
	jdff dff_B_StYp0G5t7_1(.din(w_dff_B_63h7EG696_1),.dout(w_dff_B_StYp0G5t7_1),.clk(gclk));
	jdff dff_B_Z9Mxv1hA2_1(.din(n397),.dout(w_dff_B_Z9Mxv1hA2_1),.clk(gclk));
	jdff dff_B_HvNdSAf63_1(.din(w_dff_B_Z9Mxv1hA2_1),.dout(w_dff_B_HvNdSAf63_1),.clk(gclk));
	jdff dff_B_oNpQ3xAu0_0(.din(n398),.dout(w_dff_B_oNpQ3xAu0_0),.clk(gclk));
	jdff dff_B_3kuTcEeI7_0(.din(w_dff_B_oNpQ3xAu0_0),.dout(w_dff_B_3kuTcEeI7_0),.clk(gclk));
	jdff dff_A_Fwg64vac3_1(.dout(w_n72_0[1]),.din(w_dff_A_Fwg64vac3_1),.clk(gclk));
	jdff dff_A_aNrypkVs1_1(.dout(w_dff_A_Fwg64vac3_1),.din(w_dff_A_aNrypkVs1_1),.clk(gclk));
	jdff dff_A_EUoXFZbj8_1(.dout(w_dff_A_aNrypkVs1_1),.din(w_dff_A_EUoXFZbj8_1),.clk(gclk));
	jdff dff_A_isgYk3tV9_2(.dout(w_n72_0[2]),.din(w_dff_A_isgYk3tV9_2),.clk(gclk));
	jdff dff_A_OFAGcWOO5_2(.dout(w_dff_A_isgYk3tV9_2),.din(w_dff_A_OFAGcWOO5_2),.clk(gclk));
	jdff dff_B_2tWgEd0F4_0(.din(n394),.dout(w_dff_B_2tWgEd0F4_0),.clk(gclk));
	jdff dff_A_cPFeS07j5_0(.dout(w_n112_3[0]),.din(w_dff_A_cPFeS07j5_0),.clk(gclk));
	jdff dff_A_xeprSQiT4_0(.dout(w_dff_A_cPFeS07j5_0),.din(w_dff_A_xeprSQiT4_0),.clk(gclk));
	jdff dff_A_vW5kdLoO4_1(.dout(w_n112_3[1]),.din(w_dff_A_vW5kdLoO4_1),.clk(gclk));
	jdff dff_A_fGpFw67W2_1(.dout(w_dff_A_vW5kdLoO4_1),.din(w_dff_A_fGpFw67W2_1),.clk(gclk));
	jdff dff_A_3WNCWLUH0_0(.dout(w_G58_4[0]),.din(w_dff_A_3WNCWLUH0_0),.clk(gclk));
	jdff dff_A_8kvExLf64_1(.dout(w_G58_4[1]),.din(w_dff_A_8kvExLf64_1),.clk(gclk));
	jdff dff_A_QTvtvopw5_0(.dout(w_G58_1[0]),.din(w_dff_A_QTvtvopw5_0),.clk(gclk));
	jdff dff_A_SxZL3EJ99_2(.dout(w_G58_1[2]),.din(w_dff_A_SxZL3EJ99_2),.clk(gclk));
	jdff dff_A_KxezhIql8_2(.dout(w_dff_A_SxZL3EJ99_2),.din(w_dff_A_KxezhIql8_2),.clk(gclk));
	jdff dff_A_V113hr1Z0_2(.dout(w_dff_A_KxezhIql8_2),.din(w_dff_A_V113hr1Z0_2),.clk(gclk));
	jdff dff_A_dVMNW22K3_2(.dout(w_dff_A_V113hr1Z0_2),.din(w_dff_A_dVMNW22K3_2),.clk(gclk));
	jdff dff_A_QXcKkVHt5_1(.dout(w_G58_0[1]),.din(w_dff_A_QXcKkVHt5_1),.clk(gclk));
	jdff dff_A_1P7dtv694_2(.dout(w_G58_0[2]),.din(w_dff_A_1P7dtv694_2),.clk(gclk));
	jdff dff_A_U8GyUu3t4_2(.dout(w_dff_A_1P7dtv694_2),.din(w_dff_A_U8GyUu3t4_2),.clk(gclk));
	jdff dff_A_XwAUHr957_2(.dout(w_dff_A_U8GyUu3t4_2),.din(w_dff_A_XwAUHr957_2),.clk(gclk));
	jdff dff_A_lo75t7xT1_1(.dout(w_G20_3[1]),.din(w_dff_A_lo75t7xT1_1),.clk(gclk));
	jdff dff_A_Z8t0bqlT9_2(.dout(w_G20_3[2]),.din(w_dff_A_Z8t0bqlT9_2),.clk(gclk));
	jdff dff_A_cuKsTYLP9_2(.dout(w_dff_A_Z8t0bqlT9_2),.din(w_dff_A_cuKsTYLP9_2),.clk(gclk));
	jdff dff_B_lpv1eGNU2_2(.din(n390),.dout(w_dff_B_lpv1eGNU2_2),.clk(gclk));
	jdff dff_B_q5J8ugWw8_2(.din(w_dff_B_lpv1eGNU2_2),.dout(w_dff_B_q5J8ugWw8_2),.clk(gclk));
	jdff dff_A_8Yt8kIRK5_0(.dout(w_G87_2[0]),.din(w_dff_A_8Yt8kIRK5_0),.clk(gclk));
	jdff dff_A_fyUY5LK18_0(.dout(w_dff_A_8Yt8kIRK5_0),.din(w_dff_A_fyUY5LK18_0),.clk(gclk));
	jdff dff_A_VwQATvQA5_0(.dout(w_dff_A_fyUY5LK18_0),.din(w_dff_A_VwQATvQA5_0),.clk(gclk));
	jdff dff_A_USAElrpB3_0(.dout(w_dff_A_VwQATvQA5_0),.din(w_dff_A_USAElrpB3_0),.clk(gclk));
	jdff dff_A_KdVX5pSY1_1(.dout(w_G87_2[1]),.din(w_dff_A_KdVX5pSY1_1),.clk(gclk));
	jdff dff_A_KXXiqvSB0_1(.dout(w_dff_A_KdVX5pSY1_1),.din(w_dff_A_KXXiqvSB0_1),.clk(gclk));
	jdff dff_A_bGh2cSlv5_1(.dout(w_dff_A_KXXiqvSB0_1),.din(w_dff_A_bGh2cSlv5_1),.clk(gclk));
	jdff dff_A_wKnIhUQ70_1(.dout(w_dff_A_bGh2cSlv5_1),.din(w_dff_A_wKnIhUQ70_1),.clk(gclk));
	jdff dff_A_6TU1WaPJ5_1(.dout(w_n149_1[1]),.din(w_dff_A_6TU1WaPJ5_1),.clk(gclk));
	jdff dff_A_s0awC98P6_1(.dout(w_dff_A_6TU1WaPJ5_1),.din(w_dff_A_s0awC98P6_1),.clk(gclk));
	jdff dff_B_PTmXAk1V4_1(.din(n375),.dout(w_dff_B_PTmXAk1V4_1),.clk(gclk));
	jdff dff_A_mI2UI2xn8_0(.dout(w_G232_1[0]),.din(w_dff_A_mI2UI2xn8_0),.clk(gclk));
	jdff dff_A_dzTU3Vk73_0(.dout(w_dff_A_mI2UI2xn8_0),.din(w_dff_A_dzTU3Vk73_0),.clk(gclk));
	jdff dff_A_2feKBVo45_1(.dout(w_G232_1[1]),.din(w_dff_A_2feKBVo45_1),.clk(gclk));
	jdff dff_A_ZD5WqsF17_1(.dout(w_G232_0[1]),.din(w_dff_A_ZD5WqsF17_1),.clk(gclk));
	jdff dff_A_4h9kr1yV2_1(.dout(w_dff_A_ZD5WqsF17_1),.din(w_dff_A_4h9kr1yV2_1),.clk(gclk));
	jdff dff_A_rwkKLZMV3_1(.dout(w_dff_A_4h9kr1yV2_1),.din(w_dff_A_rwkKLZMV3_1),.clk(gclk));
	jdff dff_A_3ESCjbCr0_1(.dout(w_dff_A_rwkKLZMV3_1),.din(w_dff_A_3ESCjbCr0_1),.clk(gclk));
	jdff dff_A_8P9ooGNz3_2(.dout(w_G232_0[2]),.din(w_dff_A_8P9ooGNz3_2),.clk(gclk));
	jdff dff_A_TFUnVYZP2_2(.dout(w_dff_A_8P9ooGNz3_2),.din(w_dff_A_TFUnVYZP2_2),.clk(gclk));
	jdff dff_B_Se6rDN258_0(.din(n538),.dout(w_dff_B_Se6rDN258_0),.clk(gclk));
	jdff dff_A_QuFQc92y8_1(.dout(w_n532_0[1]),.din(w_dff_A_QuFQc92y8_1),.clk(gclk));
	jdff dff_B_MbbpWLVQ2_1(.din(n525),.dout(w_dff_B_MbbpWLVQ2_1),.clk(gclk));
	jdff dff_A_5FWxVWEW6_1(.dout(w_n524_0[1]),.din(w_dff_A_5FWxVWEW6_1),.clk(gclk));
	jdff dff_A_hGqcwpXw6_0(.dout(w_n523_0[0]),.din(w_dff_A_hGqcwpXw6_0),.clk(gclk));
	jdff dff_A_j22ZuSF67_2(.dout(w_n588_0[2]),.din(w_dff_A_j22ZuSF67_2),.clk(gclk));
	jdff dff_A_jNGD2hGt5_2(.dout(w_dff_A_j22ZuSF67_2),.din(w_dff_A_jNGD2hGt5_2),.clk(gclk));
	jdff dff_B_Rk1Okfz02_0(.din(n587),.dout(w_dff_B_Rk1Okfz02_0),.clk(gclk));
	jdff dff_B_rmTxIiOP8_1(.din(n580),.dout(w_dff_B_rmTxIiOP8_1),.clk(gclk));
	jdff dff_B_lWHQMiHx3_1(.din(n581),.dout(w_dff_B_lWHQMiHx3_1),.clk(gclk));
	jdff dff_A_tcJ3l1fM8_1(.dout(w_n554_2[1]),.din(w_dff_A_tcJ3l1fM8_1),.clk(gclk));
	jdff dff_A_XfCasgZQ5_2(.dout(w_n554_2[2]),.din(w_dff_A_XfCasgZQ5_2),.clk(gclk));
	jdff dff_A_URbIeJxJ0_2(.dout(w_dff_A_XfCasgZQ5_2),.din(w_dff_A_URbIeJxJ0_2),.clk(gclk));
	jdff dff_A_D5qewFWh0_2(.dout(w_dff_A_URbIeJxJ0_2),.din(w_dff_A_D5qewFWh0_2),.clk(gclk));
	jdff dff_A_NC2qA0Je7_2(.dout(w_dff_A_D5qewFWh0_2),.din(w_dff_A_NC2qA0Je7_2),.clk(gclk));
	jdff dff_A_EgEJlBtd7_2(.dout(w_dff_A_NC2qA0Je7_2),.din(w_dff_A_EgEJlBtd7_2),.clk(gclk));
	jdff dff_A_v7eCRbFV2_0(.dout(w_n554_0[0]),.din(w_dff_A_v7eCRbFV2_0),.clk(gclk));
	jdff dff_A_oFnLsIPX9_0(.dout(w_dff_A_v7eCRbFV2_0),.din(w_dff_A_oFnLsIPX9_0),.clk(gclk));
	jdff dff_A_wpfbVsDK0_0(.dout(w_dff_A_oFnLsIPX9_0),.din(w_dff_A_wpfbVsDK0_0),.clk(gclk));
	jdff dff_A_flNQp3ij0_1(.dout(w_n554_0[1]),.din(w_dff_A_flNQp3ij0_1),.clk(gclk));
	jdff dff_A_vR3aIkMQ4_1(.dout(w_dff_A_flNQp3ij0_1),.din(w_dff_A_vR3aIkMQ4_1),.clk(gclk));
	jdff dff_B_OjW9Vqor4_3(.din(n554),.dout(w_dff_B_OjW9Vqor4_3),.clk(gclk));
	jdff dff_B_3sFmpLJj0_3(.din(w_dff_B_OjW9Vqor4_3),.dout(w_dff_B_3sFmpLJj0_3),.clk(gclk));
	jdff dff_A_QCZ4uVcY2_0(.dout(w_n534_0[0]),.din(w_dff_A_QCZ4uVcY2_0),.clk(gclk));
	jdff dff_A_pu7qAetM1_0(.dout(w_G330_0[0]),.din(w_dff_A_pu7qAetM1_0),.clk(gclk));
	jdff dff_A_zBRlUt1m9_0(.dout(w_dff_A_pu7qAetM1_0),.din(w_dff_A_zBRlUt1m9_0),.clk(gclk));
	jdff dff_A_yHfWBgP21_0(.dout(w_dff_A_zBRlUt1m9_0),.din(w_dff_A_yHfWBgP21_0),.clk(gclk));
	jdff dff_A_vMdL48KJ7_0(.dout(w_dff_A_yHfWBgP21_0),.din(w_dff_A_vMdL48KJ7_0),.clk(gclk));
	jdff dff_A_WitXuKAx9_0(.dout(w_dff_A_vMdL48KJ7_0),.din(w_dff_A_WitXuKAx9_0),.clk(gclk));
	jdff dff_A_LnxMytRQ4_0(.dout(w_dff_A_WitXuKAx9_0),.din(w_dff_A_LnxMytRQ4_0),.clk(gclk));
	jdff dff_A_AsFGWGqn1_0(.dout(w_dff_A_LnxMytRQ4_0),.din(w_dff_A_AsFGWGqn1_0),.clk(gclk));
	jdff dff_A_w7hLjyjp5_0(.dout(w_dff_A_AsFGWGqn1_0),.din(w_dff_A_w7hLjyjp5_0),.clk(gclk));
	jdff dff_A_AuvwHplx0_0(.dout(w_dff_A_w7hLjyjp5_0),.din(w_dff_A_AuvwHplx0_0),.clk(gclk));
	jdff dff_A_Hp6CzNv34_0(.dout(w_dff_A_AuvwHplx0_0),.din(w_dff_A_Hp6CzNv34_0),.clk(gclk));
	jdff dff_A_Yw1MRRPk8_0(.dout(w_dff_A_Hp6CzNv34_0),.din(w_dff_A_Yw1MRRPk8_0),.clk(gclk));
	jdff dff_A_ivacLBdj2_0(.dout(w_dff_A_Yw1MRRPk8_0),.din(w_dff_A_ivacLBdj2_0),.clk(gclk));
	jdff dff_A_ONiH80fW8_0(.dout(w_n553_2[0]),.din(w_dff_A_ONiH80fW8_0),.clk(gclk));
	jdff dff_A_Qga8kDwT0_0(.dout(w_dff_A_ONiH80fW8_0),.din(w_dff_A_Qga8kDwT0_0),.clk(gclk));
	jdff dff_A_hIiMCyqd5_0(.dout(w_dff_A_Qga8kDwT0_0),.din(w_dff_A_hIiMCyqd5_0),.clk(gclk));
	jdff dff_A_9LQ1UWGS1_0(.dout(w_dff_A_hIiMCyqd5_0),.din(w_dff_A_9LQ1UWGS1_0),.clk(gclk));
	jdff dff_A_wGWEvXks2_0(.dout(w_dff_A_9LQ1UWGS1_0),.din(w_dff_A_wGWEvXks2_0),.clk(gclk));
	jdff dff_A_PPgkTpKD3_0(.dout(w_dff_A_wGWEvXks2_0),.din(w_dff_A_PPgkTpKD3_0),.clk(gclk));
	jdff dff_A_TIhhQQDF5_0(.dout(w_dff_A_PPgkTpKD3_0),.din(w_dff_A_TIhhQQDF5_0),.clk(gclk));
	jdff dff_A_pbBn6JLd6_0(.dout(w_dff_A_TIhhQQDF5_0),.din(w_dff_A_pbBn6JLd6_0),.clk(gclk));
	jdff dff_A_LuFLmaxL6_0(.dout(w_dff_A_pbBn6JLd6_0),.din(w_dff_A_LuFLmaxL6_0),.clk(gclk));
	jdff dff_A_c6Fd7P0W7_1(.dout(w_n553_2[1]),.din(w_dff_A_c6Fd7P0W7_1),.clk(gclk));
	jdff dff_A_IsVMXQcS6_1(.dout(w_dff_A_c6Fd7P0W7_1),.din(w_dff_A_IsVMXQcS6_1),.clk(gclk));
	jdff dff_A_6naygO3F7_1(.dout(w_dff_A_IsVMXQcS6_1),.din(w_dff_A_6naygO3F7_1),.clk(gclk));
	jdff dff_A_DKq2xQ6u8_1(.dout(w_dff_A_6naygO3F7_1),.din(w_dff_A_DKq2xQ6u8_1),.clk(gclk));
	jdff dff_A_NKo3CyIm1_1(.dout(w_dff_A_DKq2xQ6u8_1),.din(w_dff_A_NKo3CyIm1_1),.clk(gclk));
	jdff dff_A_yR7tohNl7_0(.dout(w_n553_0[0]),.din(w_dff_A_yR7tohNl7_0),.clk(gclk));
	jdff dff_A_tCDrSdfO1_0(.dout(w_dff_A_yR7tohNl7_0),.din(w_dff_A_tCDrSdfO1_0),.clk(gclk));
	jdff dff_A_wfnlm8TV8_0(.dout(w_dff_A_tCDrSdfO1_0),.din(w_dff_A_wfnlm8TV8_0),.clk(gclk));
	jdff dff_A_9d4p2KhZ4_0(.dout(w_dff_A_wfnlm8TV8_0),.din(w_dff_A_9d4p2KhZ4_0),.clk(gclk));
	jdff dff_A_sLxuViSS4_2(.dout(w_n553_0[2]),.din(w_dff_A_sLxuViSS4_2),.clk(gclk));
	jdff dff_A_TSxV9rCA7_2(.dout(w_dff_A_sLxuViSS4_2),.din(w_dff_A_TSxV9rCA7_2),.clk(gclk));
	jdff dff_A_qzHAvkSR4_2(.dout(w_dff_A_TSxV9rCA7_2),.din(w_dff_A_qzHAvkSR4_2),.clk(gclk));
	jdff dff_A_2ev2g0lR9_2(.dout(w_dff_A_qzHAvkSR4_2),.din(w_dff_A_2ev2g0lR9_2),.clk(gclk));
	jdff dff_A_9qtZupMq0_2(.dout(w_dff_A_2ev2g0lR9_2),.din(w_dff_A_9qtZupMq0_2),.clk(gclk));
	jdff dff_A_hDnjk1EL9_2(.dout(w_dff_A_9qtZupMq0_2),.din(w_dff_A_hDnjk1EL9_2),.clk(gclk));
	jdff dff_A_NnQ7vhNI6_1(.dout(w_n552_0[1]),.din(w_dff_A_NnQ7vhNI6_1),.clk(gclk));
	jdff dff_A_F8I1H2sb2_1(.dout(w_dff_A_NnQ7vhNI6_1),.din(w_dff_A_F8I1H2sb2_1),.clk(gclk));
	jdff dff_A_UV4VtZOZ0_1(.dout(w_dff_A_F8I1H2sb2_1),.din(w_dff_A_UV4VtZOZ0_1),.clk(gclk));
	jdff dff_A_yNMjwTIC6_1(.dout(w_dff_A_UV4VtZOZ0_1),.din(w_dff_A_yNMjwTIC6_1),.clk(gclk));
	jdff dff_A_TMobsgdo7_1(.dout(w_dff_A_yNMjwTIC6_1),.din(w_dff_A_TMobsgdo7_1),.clk(gclk));
	jdff dff_A_y4GBWH5w5_1(.dout(w_dff_A_TMobsgdo7_1),.din(w_dff_A_y4GBWH5w5_1),.clk(gclk));
	jdff dff_A_DLDWHXGW0_1(.dout(w_dff_A_y4GBWH5w5_1),.din(w_dff_A_DLDWHXGW0_1),.clk(gclk));
	jdff dff_A_gmu7h94X8_2(.dout(w_n552_0[2]),.din(w_dff_A_gmu7h94X8_2),.clk(gclk));
	jdff dff_A_xh99m26B7_2(.dout(w_dff_A_gmu7h94X8_2),.din(w_dff_A_xh99m26B7_2),.clk(gclk));
	jdff dff_A_EEcE2K3w7_2(.dout(w_dff_A_xh99m26B7_2),.din(w_dff_A_EEcE2K3w7_2),.clk(gclk));
	jdff dff_A_7J9ktyR82_2(.dout(w_dff_A_EEcE2K3w7_2),.din(w_dff_A_7J9ktyR82_2),.clk(gclk));
	jdff dff_A_pY5Wevk57_2(.dout(w_dff_A_7J9ktyR82_2),.din(w_dff_A_pY5Wevk57_2),.clk(gclk));
	jdff dff_A_XitxJwXg7_2(.dout(w_dff_A_pY5Wevk57_2),.din(w_dff_A_XitxJwXg7_2),.clk(gclk));
	jdff dff_A_bbdjmFzC1_2(.dout(w_dff_A_XitxJwXg7_2),.din(w_dff_A_bbdjmFzC1_2),.clk(gclk));
	jdff dff_A_i7KpoBFg0_0(.dout(w_G213_0[0]),.din(w_dff_A_i7KpoBFg0_0),.clk(gclk));
	jdff dff_A_OZZpiNyz2_2(.dout(w_G213_0[2]),.din(w_dff_A_OZZpiNyz2_2),.clk(gclk));
	jdff dff_A_xOFY8sRx8_0(.dout(w_n113_1[0]),.din(w_dff_A_xOFY8sRx8_0),.clk(gclk));
	jdff dff_A_31dEtmIx9_0(.dout(w_dff_A_xOFY8sRx8_0),.din(w_dff_A_31dEtmIx9_0),.clk(gclk));
	jdff dff_A_uTS2VDkH1_1(.dout(w_n113_1[1]),.din(w_dff_A_uTS2VDkH1_1),.clk(gclk));
	jdff dff_A_xhApSxfL6_1(.dout(w_dff_A_uTS2VDkH1_1),.din(w_dff_A_xhApSxfL6_1),.clk(gclk));
	jdff dff_A_QSjvWHOz2_1(.dout(w_dff_A_xhApSxfL6_1),.din(w_dff_A_QSjvWHOz2_1),.clk(gclk));
	jdff dff_A_L8MHFwn28_1(.dout(w_dff_A_QSjvWHOz2_1),.din(w_dff_A_L8MHFwn28_1),.clk(gclk));
	jdff dff_A_HDnpnNPw1_1(.dout(w_dff_A_L8MHFwn28_1),.din(w_dff_A_HDnpnNPw1_1),.clk(gclk));
	jdff dff_A_eA1RIcGE2_1(.dout(w_dff_A_HDnpnNPw1_1),.din(w_dff_A_eA1RIcGE2_1),.clk(gclk));
	jdff dff_A_475euyrk0_1(.dout(w_dff_A_eA1RIcGE2_1),.din(w_dff_A_475euyrk0_1),.clk(gclk));
	jdff dff_A_Ak4a31pQ8_1(.dout(w_dff_A_475euyrk0_1),.din(w_dff_A_Ak4a31pQ8_1),.clk(gclk));
	jdff dff_A_zbv5gQFc3_1(.dout(w_dff_A_Ak4a31pQ8_1),.din(w_dff_A_zbv5gQFc3_1),.clk(gclk));
	jdff dff_A_APQK90eA1_1(.dout(w_dff_A_zbv5gQFc3_1),.din(w_dff_A_APQK90eA1_1),.clk(gclk));
	jdff dff_A_sSlKkMgd4_1(.dout(w_dff_A_APQK90eA1_1),.din(w_dff_A_sSlKkMgd4_1),.clk(gclk));
	jdff dff_A_d5cGi8cl6_1(.dout(w_dff_A_sSlKkMgd4_1),.din(w_dff_A_d5cGi8cl6_1),.clk(gclk));
	jdff dff_A_97odbeVd7_1(.dout(w_dff_A_d5cGi8cl6_1),.din(w_dff_A_97odbeVd7_1),.clk(gclk));
	jdff dff_A_JjQpRUKt4_1(.dout(w_dff_A_97odbeVd7_1),.din(w_dff_A_JjQpRUKt4_1),.clk(gclk));
	jdff dff_A_oaT70Ert9_1(.dout(w_dff_A_JjQpRUKt4_1),.din(w_dff_A_oaT70Ert9_1),.clk(gclk));
	jdff dff_A_KMEJokLl8_1(.dout(w_G343_0[1]),.din(w_dff_A_KMEJokLl8_1),.clk(gclk));
	jdff dff_A_yxanHp4w4_1(.dout(w_dff_A_KMEJokLl8_1),.din(w_dff_A_yxanHp4w4_1),.clk(gclk));
	jdff dff_A_hdHP6RrK9_1(.dout(w_dff_A_yxanHp4w4_1),.din(w_dff_A_hdHP6RrK9_1),.clk(gclk));
	jdff dff_A_uYaC6xKx9_1(.dout(w_n374_0[1]),.din(w_dff_A_uYaC6xKx9_1),.clk(gclk));
	jdff dff_B_qaOjpxk54_0(.din(n365),.dout(w_dff_B_qaOjpxk54_0),.clk(gclk));
	jdff dff_B_lBI3HOGf2_1(.din(n348),.dout(w_dff_B_lBI3HOGf2_1),.clk(gclk));
	jdff dff_B_Ob1JtJHk1_1(.din(n343),.dout(w_dff_B_Ob1JtJHk1_1),.clk(gclk));
	jdff dff_A_8MqtPDd34_0(.dout(w_n339_0[0]),.din(w_dff_A_8MqtPDd34_0),.clk(gclk));
	jdff dff_A_scipC3JV3_0(.dout(w_dff_A_8MqtPDd34_0),.din(w_dff_A_scipC3JV3_0),.clk(gclk));
	jdff dff_A_hlJK438k8_0(.dout(w_G294_3[0]),.din(w_dff_A_hlJK438k8_0),.clk(gclk));
	jdff dff_A_lBD9smrQ6_0(.dout(w_dff_A_hlJK438k8_0),.din(w_dff_A_lBD9smrQ6_0),.clk(gclk));
	jdff dff_A_xMGadafd5_0(.dout(w_dff_A_lBD9smrQ6_0),.din(w_dff_A_xMGadafd5_0),.clk(gclk));
	jdff dff_A_Z0FLKKmW4_0(.dout(w_dff_A_xMGadafd5_0),.din(w_dff_A_Z0FLKKmW4_0),.clk(gclk));
	jdff dff_A_fMy63A7W0_0(.dout(w_G294_0[0]),.din(w_dff_A_fMy63A7W0_0),.clk(gclk));
	jdff dff_A_FzlvnR3r4_0(.dout(w_dff_A_fMy63A7W0_0),.din(w_dff_A_FzlvnR3r4_0),.clk(gclk));
	jdff dff_A_UoXAoSkh7_0(.dout(w_dff_A_FzlvnR3r4_0),.din(w_dff_A_UoXAoSkh7_0),.clk(gclk));
	jdff dff_A_OtJncsHi2_1(.dout(w_G294_0[1]),.din(w_dff_A_OtJncsHi2_1),.clk(gclk));
	jdff dff_A_HwBBcvxQ0_1(.dout(w_dff_A_OtJncsHi2_1),.din(w_dff_A_HwBBcvxQ0_1),.clk(gclk));
	jdff dff_A_zA8cSDbK4_1(.dout(w_dff_A_HwBBcvxQ0_1),.din(w_dff_A_zA8cSDbK4_1),.clk(gclk));
	jdff dff_A_ofqVPrrA0_0(.dout(w_n196_1[0]),.din(w_dff_A_ofqVPrrA0_0),.clk(gclk));
	jdff dff_A_5oFpw9a35_1(.dout(w_n196_1[1]),.din(w_dff_A_5oFpw9a35_1),.clk(gclk));
	jdff dff_B_0ZqnHgth1_0(.din(n335),.dout(w_dff_B_0ZqnHgth1_0),.clk(gclk));
	jdff dff_A_5dVkZH5j0_0(.dout(w_n334_0[0]),.din(w_dff_A_5dVkZH5j0_0),.clk(gclk));
	jdff dff_A_UaLXOGn53_0(.dout(w_dff_A_5dVkZH5j0_0),.din(w_dff_A_UaLXOGn53_0),.clk(gclk));
	jdff dff_B_rBOlzuRi6_0(.din(n333),.dout(w_dff_B_rBOlzuRi6_0),.clk(gclk));
	jdff dff_A_HgI6wU3w3_0(.dout(w_G107_3[0]),.din(w_dff_A_HgI6wU3w3_0),.clk(gclk));
	jdff dff_A_vTk5FaV18_1(.dout(w_G107_3[1]),.din(w_dff_A_vTk5FaV18_1),.clk(gclk));
	jdff dff_B_CckvPW0B8_0(.din(n331),.dout(w_dff_B_CckvPW0B8_0),.clk(gclk));
	jdff dff_B_FItYXkBg8_1(.din(n316),.dout(w_dff_B_FItYXkBg8_1),.clk(gclk));
	jdff dff_A_LnP6kG3p1_1(.dout(w_G190_3[1]),.din(w_dff_A_LnP6kG3p1_1),.clk(gclk));
	jdff dff_A_vWUGqqlo7_1(.dout(w_dff_A_LnP6kG3p1_1),.din(w_dff_A_vWUGqqlo7_1),.clk(gclk));
	jdff dff_A_I3zk9c6d7_1(.dout(w_dff_A_vWUGqqlo7_1),.din(w_dff_A_I3zk9c6d7_1),.clk(gclk));
	jdff dff_A_YVQlmWJZ8_1(.dout(w_dff_A_I3zk9c6d7_1),.din(w_dff_A_YVQlmWJZ8_1),.clk(gclk));
	jdff dff_A_qwKoobid7_1(.dout(w_dff_A_YVQlmWJZ8_1),.din(w_dff_A_qwKoobid7_1),.clk(gclk));
	jdff dff_A_d09YCIYx6_1(.dout(w_dff_A_qwKoobid7_1),.din(w_dff_A_d09YCIYx6_1),.clk(gclk));
	jdff dff_A_8Y5cjDrJ2_1(.dout(w_dff_A_d09YCIYx6_1),.din(w_dff_A_8Y5cjDrJ2_1),.clk(gclk));
	jdff dff_A_nQrwdI367_2(.dout(w_G190_3[2]),.din(w_dff_A_nQrwdI367_2),.clk(gclk));
	jdff dff_A_NMLBWp9v4_2(.dout(w_dff_A_nQrwdI367_2),.din(w_dff_A_NMLBWp9v4_2),.clk(gclk));
	jdff dff_A_lZhEDrAO9_2(.dout(w_dff_A_NMLBWp9v4_2),.din(w_dff_A_lZhEDrAO9_2),.clk(gclk));
	jdff dff_A_AVRwB63d9_2(.dout(w_dff_A_lZhEDrAO9_2),.din(w_dff_A_AVRwB63d9_2),.clk(gclk));
	jdff dff_A_2EK5RY1d5_2(.dout(w_dff_A_AVRwB63d9_2),.din(w_dff_A_2EK5RY1d5_2),.clk(gclk));
	jdff dff_A_CAEEaN0d5_2(.dout(w_dff_A_2EK5RY1d5_2),.din(w_dff_A_CAEEaN0d5_2),.clk(gclk));
	jdff dff_A_pX9m3u7g3_2(.dout(w_dff_A_CAEEaN0d5_2),.din(w_dff_A_pX9m3u7g3_2),.clk(gclk));
	jdff dff_B_YUhf0cSD3_0(.din(n317),.dout(w_dff_B_YUhf0cSD3_0),.clk(gclk));
	jdff dff_B_2Ups4ZUZ1_1(.din(n289),.dout(w_dff_B_2Ups4ZUZ1_1),.clk(gclk));
	jdff dff_A_r9xSnZwN3_1(.dout(w_n312_0[1]),.din(w_dff_A_r9xSnZwN3_1),.clk(gclk));
	jdff dff_B_ESiqQjT38_1(.din(n309),.dout(w_dff_B_ESiqQjT38_1),.clk(gclk));
	jdff dff_A_Z1wBMHEA7_0(.dout(w_n106_0[0]),.din(w_dff_A_Z1wBMHEA7_0),.clk(gclk));
	jdff dff_A_IQoxZCL04_0(.dout(w_dff_A_Z1wBMHEA7_0),.din(w_dff_A_IQoxZCL04_0),.clk(gclk));
	jdff dff_A_k0B8T4cV2_0(.dout(w_dff_A_IQoxZCL04_0),.din(w_dff_A_k0B8T4cV2_0),.clk(gclk));
	jdff dff_A_X3OGsQtv9_1(.dout(w_n88_0[1]),.din(w_dff_A_X3OGsQtv9_1),.clk(gclk));
	jdff dff_A_kryDyheK3_1(.dout(w_dff_A_X3OGsQtv9_1),.din(w_dff_A_kryDyheK3_1),.clk(gclk));
	jdff dff_A_JLnUbvKH6_1(.dout(w_dff_A_kryDyheK3_1),.din(w_dff_A_JLnUbvKH6_1),.clk(gclk));
	jdff dff_A_8vJy3UYI7_2(.dout(w_n88_0[2]),.din(w_dff_A_8vJy3UYI7_2),.clk(gclk));
	jdff dff_A_HO9wEOsL3_1(.dout(w_n166_1[1]),.din(w_dff_A_HO9wEOsL3_1),.clk(gclk));
	jdff dff_A_y18LBZqP9_2(.dout(w_n166_1[2]),.din(w_dff_A_y18LBZqP9_2),.clk(gclk));
	jdff dff_A_JyxRLC5D6_1(.dout(w_n303_0[1]),.din(w_dff_A_JyxRLC5D6_1),.clk(gclk));
	jdff dff_A_4V7aPM779_1(.dout(w_n300_0[1]),.din(w_dff_A_4V7aPM779_1),.clk(gclk));
	jdff dff_A_FPAyaDou3_0(.dout(w_n298_0[0]),.din(w_dff_A_FPAyaDou3_0),.clk(gclk));
	jdff dff_A_BjWdFFvn0_0(.dout(w_dff_A_FPAyaDou3_0),.din(w_dff_A_BjWdFFvn0_0),.clk(gclk));
	jdff dff_A_IkzaHFq56_1(.dout(w_n185_2[1]),.din(w_dff_A_IkzaHFq56_1),.clk(gclk));
	jdff dff_A_ExKRS7R52_1(.dout(w_dff_A_IkzaHFq56_1),.din(w_dff_A_ExKRS7R52_1),.clk(gclk));
	jdff dff_A_DgwHk2E26_0(.dout(w_n105_1[0]),.din(w_dff_A_DgwHk2E26_0),.clk(gclk));
	jdff dff_A_yvlK8xgo9_2(.dout(w_n105_1[2]),.din(w_dff_A_yvlK8xgo9_2),.clk(gclk));
	jdff dff_A_2nabn6W25_0(.dout(w_n296_0[0]),.din(w_dff_A_2nabn6W25_0),.clk(gclk));
	jdff dff_A_KluREwqb8_0(.dout(w_dff_A_2nabn6W25_0),.din(w_dff_A_KluREwqb8_0),.clk(gclk));
	jdff dff_A_bOauCHnq3_0(.dout(w_n105_0[0]),.din(w_dff_A_bOauCHnq3_0),.clk(gclk));
	jdff dff_A_XGRbaAcM7_2(.dout(w_n105_0[2]),.din(w_dff_A_XGRbaAcM7_2),.clk(gclk));
	jdff dff_A_qMub9GaM3_2(.dout(w_dff_A_XGRbaAcM7_2),.din(w_dff_A_qMub9GaM3_2),.clk(gclk));
	jdff dff_A_olsPP0wh9_2(.dout(w_dff_A_qMub9GaM3_2),.din(w_dff_A_olsPP0wh9_2),.clk(gclk));
	jdff dff_A_w57tCPB92_0(.dout(w_G20_4[0]),.din(w_dff_A_w57tCPB92_0),.clk(gclk));
	jdff dff_A_Doideh6u1_1(.dout(w_G20_4[1]),.din(w_dff_A_Doideh6u1_1),.clk(gclk));
	jdff dff_A_UDaGBK512_1(.dout(w_dff_A_Doideh6u1_1),.din(w_dff_A_UDaGBK512_1),.clk(gclk));
	jdff dff_A_dCzj3Zxc8_1(.dout(w_dff_A_UDaGBK512_1),.din(w_dff_A_dCzj3Zxc8_1),.clk(gclk));
	jdff dff_A_iypLFhgt0_1(.dout(w_dff_A_dCzj3Zxc8_1),.din(w_dff_A_iypLFhgt0_1),.clk(gclk));
	jdff dff_A_3U20ts2s3_1(.dout(w_n189_1[1]),.din(w_dff_A_3U20ts2s3_1),.clk(gclk));
	jdff dff_A_voGAwgge3_0(.dout(w_G97_3[0]),.din(w_dff_A_voGAwgge3_0),.clk(gclk));
	jdff dff_A_2m34iBkZ9_0(.dout(w_dff_A_voGAwgge3_0),.din(w_dff_A_2m34iBkZ9_0),.clk(gclk));
	jdff dff_A_Gn9pDYYA7_0(.dout(w_dff_A_2m34iBkZ9_0),.din(w_dff_A_Gn9pDYYA7_0),.clk(gclk));
	jdff dff_A_z5vr8YyK9_1(.dout(w_G97_3[1]),.din(w_dff_A_z5vr8YyK9_1),.clk(gclk));
	jdff dff_A_mdV8smXh6_1(.dout(w_dff_A_z5vr8YyK9_1),.din(w_dff_A_mdV8smXh6_1),.clk(gclk));
	jdff dff_A_rSAM8eBC8_1(.dout(w_dff_A_mdV8smXh6_1),.din(w_dff_A_rSAM8eBC8_1),.clk(gclk));
	jdff dff_A_DYzNfhCS8_0(.dout(w_G270_0[0]),.din(w_dff_A_DYzNfhCS8_0),.clk(gclk));
	jdff dff_A_87s3fh111_0(.dout(w_dff_A_DYzNfhCS8_0),.din(w_dff_A_87s3fh111_0),.clk(gclk));
	jdff dff_A_HKylwl923_0(.dout(w_dff_A_87s3fh111_0),.din(w_dff_A_HKylwl923_0),.clk(gclk));
	jdff dff_A_cQ54mkdH5_0(.dout(w_dff_A_HKylwl923_0),.din(w_dff_A_cQ54mkdH5_0),.clk(gclk));
	jdff dff_B_KP5W2ISa8_1(.din(n280),.dout(w_dff_B_KP5W2ISa8_1),.clk(gclk));
	jdff dff_A_82NHEE7b0_1(.dout(w_n281_0[1]),.din(w_dff_A_82NHEE7b0_1),.clk(gclk));
	jdff dff_A_aWCZ3PV36_1(.dout(w_dff_A_82NHEE7b0_1),.din(w_dff_A_aWCZ3PV36_1),.clk(gclk));
	jdff dff_A_6i5ky61a5_0(.dout(w_G303_2[0]),.din(w_dff_A_6i5ky61a5_0),.clk(gclk));
	jdff dff_A_kIdF8Lbd6_0(.dout(w_dff_A_6i5ky61a5_0),.din(w_dff_A_kIdF8Lbd6_0),.clk(gclk));
	jdff dff_A_dRIFEpXE2_0(.dout(w_dff_A_kIdF8Lbd6_0),.din(w_dff_A_dRIFEpXE2_0),.clk(gclk));
	jdff dff_A_hRLX5UKi5_1(.dout(w_G303_2[1]),.din(w_dff_A_hRLX5UKi5_1),.clk(gclk));
	jdff dff_A_e2w0AW7a7_1(.dout(w_dff_A_hRLX5UKi5_1),.din(w_dff_A_e2w0AW7a7_1),.clk(gclk));
	jdff dff_A_ntHYKpwE3_1(.dout(w_dff_A_e2w0AW7a7_1),.din(w_dff_A_ntHYKpwE3_1),.clk(gclk));
	jdff dff_A_zHbiGjTa4_1(.dout(w_dff_A_ntHYKpwE3_1),.din(w_dff_A_zHbiGjTa4_1),.clk(gclk));
	jdff dff_A_2rZxIfci9_0(.dout(w_G303_0[0]),.din(w_dff_A_2rZxIfci9_0),.clk(gclk));
	jdff dff_A_wySlA28l1_0(.dout(w_dff_A_2rZxIfci9_0),.din(w_dff_A_wySlA28l1_0),.clk(gclk));
	jdff dff_A_rs9LaVd82_0(.dout(w_dff_A_wySlA28l1_0),.din(w_dff_A_rs9LaVd82_0),.clk(gclk));
	jdff dff_A_NgDrAnaq0_2(.dout(w_G303_0[2]),.din(w_dff_A_NgDrAnaq0_2),.clk(gclk));
	jdff dff_A_3JGXcpoo3_2(.dout(w_dff_A_NgDrAnaq0_2),.din(w_dff_A_3JGXcpoo3_2),.clk(gclk));
	jdff dff_A_oCBzW6XC8_2(.dout(w_dff_A_3JGXcpoo3_2),.din(w_dff_A_oCBzW6XC8_2),.clk(gclk));
	jdff dff_A_r4fvZwfG5_2(.dout(w_dff_A_oCBzW6XC8_2),.din(w_dff_A_r4fvZwfG5_2),.clk(gclk));
	jdff dff_A_xM3lupbG2_1(.dout(w_G264_0[1]),.din(w_dff_A_xM3lupbG2_1),.clk(gclk));
	jdff dff_A_UCe6xSXk1_1(.dout(w_dff_A_xM3lupbG2_1),.din(w_dff_A_UCe6xSXk1_1),.clk(gclk));
	jdff dff_A_FVoRFnKk5_1(.dout(w_dff_A_UCe6xSXk1_1),.din(w_dff_A_FVoRFnKk5_1),.clk(gclk));
	jdff dff_A_JKOTdtIu3_1(.dout(w_dff_A_FVoRFnKk5_1),.din(w_dff_A_JKOTdtIu3_1),.clk(gclk));
	jdff dff_A_sz6Xv0Vz2_2(.dout(w_G264_0[2]),.din(w_dff_A_sz6Xv0Vz2_2),.clk(gclk));
	jdff dff_A_DpVal63g7_2(.dout(w_dff_A_sz6Xv0Vz2_2),.din(w_dff_A_DpVal63g7_2),.clk(gclk));
	jdff dff_B_g8zLtGBf1_1(.din(n268),.dout(w_dff_B_g8zLtGBf1_1),.clk(gclk));
	jdff dff_A_CvAUyHMO4_1(.dout(w_n274_0[1]),.din(w_dff_A_CvAUyHMO4_1),.clk(gclk));
	jdff dff_A_SAu8rnnx7_0(.dout(w_n270_0[0]),.din(w_dff_A_SAu8rnnx7_0),.clk(gclk));
	jdff dff_B_JTvsNzW86_2(.din(n270),.dout(w_dff_B_JTvsNzW86_2),.clk(gclk));
	jdff dff_A_2QHmvWhb3_0(.dout(w_n112_4[0]),.din(w_dff_A_2QHmvWhb3_0),.clk(gclk));
	jdff dff_A_5e450z2C9_0(.dout(w_dff_A_2QHmvWhb3_0),.din(w_dff_A_5e450z2C9_0),.clk(gclk));
	jdff dff_A_kV7y1LTJ4_0(.dout(w_dff_A_5e450z2C9_0),.din(w_dff_A_kV7y1LTJ4_0),.clk(gclk));
	jdff dff_A_Scn0bNSL3_0(.dout(w_dff_A_kV7y1LTJ4_0),.din(w_dff_A_Scn0bNSL3_0),.clk(gclk));
	jdff dff_A_3MA49UyW2_1(.dout(w_n112_4[1]),.din(w_dff_A_3MA49UyW2_1),.clk(gclk));
	jdff dff_A_5Ud1X3uD6_0(.dout(w_G1_1[0]),.din(w_dff_A_5Ud1X3uD6_0),.clk(gclk));
	jdff dff_A_5ICkNZKZ6_0(.dout(w_dff_A_5Ud1X3uD6_0),.din(w_dff_A_5ICkNZKZ6_0),.clk(gclk));
	jdff dff_A_8JtEjNTX7_0(.dout(w_dff_A_5ICkNZKZ6_0),.din(w_dff_A_8JtEjNTX7_0),.clk(gclk));
	jdff dff_A_6SIYP9g29_1(.dout(w_G1_1[1]),.din(w_dff_A_6SIYP9g29_1),.clk(gclk));
	jdff dff_B_eeystC7o7_0(.din(n266),.dout(w_dff_B_eeystC7o7_0),.clk(gclk));
	jdff dff_B_cumdVIoI3_1(.din(n260),.dout(w_dff_B_cumdVIoI3_1),.clk(gclk));
	jdff dff_A_Zr3jYwrt4_0(.dout(w_n262_0[0]),.din(w_dff_A_Zr3jYwrt4_0),.clk(gclk));
	jdff dff_A_K44SgIkp8_0(.dout(w_n259_0[0]),.din(w_dff_A_K44SgIkp8_0),.clk(gclk));
	jdff dff_A_2284LzIR3_0(.dout(w_dff_A_K44SgIkp8_0),.din(w_dff_A_2284LzIR3_0),.clk(gclk));
	jdff dff_A_JmzGA6ll1_0(.dout(w_n257_0[0]),.din(w_dff_A_JmzGA6ll1_0),.clk(gclk));
	jdff dff_A_IQNMlTkt4_1(.dout(w_n255_0[1]),.din(w_dff_A_IQNMlTkt4_1),.clk(gclk));
	jdff dff_A_3qbxSaiM9_0(.dout(w_G77_4[0]),.din(w_dff_A_3qbxSaiM9_0),.clk(gclk));
	jdff dff_A_yO1GxoUW4_0(.dout(w_G77_1[0]),.din(w_dff_A_yO1GxoUW4_0),.clk(gclk));
	jdff dff_A_S3RsoBOp6_2(.dout(w_G77_1[2]),.din(w_dff_A_S3RsoBOp6_2),.clk(gclk));
	jdff dff_A_wpN8eSkS4_2(.dout(w_dff_A_S3RsoBOp6_2),.din(w_dff_A_wpN8eSkS4_2),.clk(gclk));
	jdff dff_A_qlA9x71M5_2(.dout(w_dff_A_wpN8eSkS4_2),.din(w_dff_A_qlA9x71M5_2),.clk(gclk));
	jdff dff_A_tDndV5yl1_2(.dout(w_dff_A_qlA9x71M5_2),.din(w_dff_A_tDndV5yl1_2),.clk(gclk));
	jdff dff_B_jOlQVX3f4_2(.din(n249),.dout(w_dff_B_jOlQVX3f4_2),.clk(gclk));
	jdff dff_B_XWyL3vEe4_2(.din(w_dff_B_jOlQVX3f4_2),.dout(w_dff_B_XWyL3vEe4_2),.clk(gclk));
	jdff dff_A_D9ebEIyT2_0(.dout(w_G107_4[0]),.din(w_dff_A_D9ebEIyT2_0),.clk(gclk));
	jdff dff_A_5wqENpGk3_0(.dout(w_dff_A_D9ebEIyT2_0),.din(w_dff_A_5wqENpGk3_0),.clk(gclk));
	jdff dff_A_MGIj5Kmt6_0(.dout(w_dff_A_5wqENpGk3_0),.din(w_dff_A_MGIj5Kmt6_0),.clk(gclk));
	jdff dff_A_MLMpndjC3_0(.dout(w_dff_A_MGIj5Kmt6_0),.din(w_dff_A_MLMpndjC3_0),.clk(gclk));
	jdff dff_A_Ww2dKrqe4_0(.dout(w_dff_A_MLMpndjC3_0),.din(w_dff_A_Ww2dKrqe4_0),.clk(gclk));
	jdff dff_A_eoP6Xd8S5_0(.dout(w_dff_A_Ww2dKrqe4_0),.din(w_dff_A_eoP6Xd8S5_0),.clk(gclk));
	jdff dff_A_KXzl8J1t1_0(.dout(w_G33_8[0]),.din(w_dff_A_KXzl8J1t1_0),.clk(gclk));
	jdff dff_B_AdmWGaOe4_1(.din(n236),.dout(w_dff_B_AdmWGaOe4_1),.clk(gclk));
	jdff dff_B_97RKkF8C6_1(.din(n226),.dout(w_dff_B_97RKkF8C6_1),.clk(gclk));
	jdff dff_A_bf5y3ZLr2_0(.dout(w_n230_0[0]),.din(w_dff_A_bf5y3ZLr2_0),.clk(gclk));
	jdff dff_A_7m6aJFYP6_0(.dout(w_n151_3[0]),.din(w_dff_A_7m6aJFYP6_0),.clk(gclk));
	jdff dff_A_iUfZNA4n8_0(.dout(w_dff_A_7m6aJFYP6_0),.din(w_dff_A_iUfZNA4n8_0),.clk(gclk));
	jdff dff_A_dRMR1wIA9_1(.dout(w_n151_3[1]),.din(w_dff_A_dRMR1wIA9_1),.clk(gclk));
	jdff dff_A_LdnhFLWB7_1(.dout(w_dff_A_dRMR1wIA9_1),.din(w_dff_A_LdnhFLWB7_1),.clk(gclk));
	jdff dff_A_cpfsNo8c5_0(.dout(w_n91_1[0]),.din(w_dff_A_cpfsNo8c5_0),.clk(gclk));
	jdff dff_A_S7CcMjSb9_0(.dout(w_dff_A_cpfsNo8c5_0),.din(w_dff_A_S7CcMjSb9_0),.clk(gclk));
	jdff dff_A_dnvwvo7A0_0(.dout(w_dff_A_S7CcMjSb9_0),.din(w_dff_A_dnvwvo7A0_0),.clk(gclk));
	jdff dff_A_vrlGWjLz1_1(.dout(w_n91_0[1]),.din(w_dff_A_vrlGWjLz1_1),.clk(gclk));
	jdff dff_A_7ehDI4M01_0(.dout(w_G257_1[0]),.din(w_dff_A_7ehDI4M01_0),.clk(gclk));
	jdff dff_A_iW93BtpF8_0(.dout(w_dff_A_7ehDI4M01_0),.din(w_dff_A_iW93BtpF8_0),.clk(gclk));
	jdff dff_A_VQhbRkxc1_0(.dout(w_dff_A_iW93BtpF8_0),.din(w_dff_A_VQhbRkxc1_0),.clk(gclk));
	jdff dff_A_PVlXVh3K7_0(.dout(w_dff_A_VQhbRkxc1_0),.din(w_dff_A_PVlXVh3K7_0),.clk(gclk));
	jdff dff_A_R8TMyVsb5_1(.dout(w_G257_1[1]),.din(w_dff_A_R8TMyVsb5_1),.clk(gclk));
	jdff dff_A_vWbAlTR88_1(.dout(w_G257_0[1]),.din(w_dff_A_vWbAlTR88_1),.clk(gclk));
	jdff dff_A_ltqoHmBF3_1(.dout(w_dff_A_vWbAlTR88_1),.din(w_dff_A_ltqoHmBF3_1),.clk(gclk));
	jdff dff_A_xWL67o6i4_2(.dout(w_G257_0[2]),.din(w_dff_A_xWL67o6i4_2),.clk(gclk));
	jdff dff_A_U2PfyQfO1_2(.dout(w_dff_A_xWL67o6i4_2),.din(w_dff_A_U2PfyQfO1_2),.clk(gclk));
	jdff dff_A_amvJWUy39_1(.dout(w_n228_0[1]),.din(w_dff_A_amvJWUy39_1),.clk(gclk));
	jdff dff_A_LSUBSLPz7_0(.dout(w_n221_0[0]),.din(w_dff_A_LSUBSLPz7_0),.clk(gclk));
	jdff dff_A_wRipiJfK3_0(.dout(w_dff_A_LSUBSLPz7_0),.din(w_dff_A_wRipiJfK3_0),.clk(gclk));
	jdff dff_A_IDwFqbWc2_1(.dout(w_n221_0[1]),.din(w_dff_A_IDwFqbWc2_1),.clk(gclk));
	jdff dff_A_wmPnpOg62_1(.dout(w_dff_A_IDwFqbWc2_1),.din(w_dff_A_wmPnpOg62_1),.clk(gclk));
	jdff dff_A_70MqtVLv0_0(.dout(w_G283_3[0]),.din(w_dff_A_70MqtVLv0_0),.clk(gclk));
	jdff dff_A_CMYqqWq50_0(.dout(w_dff_A_70MqtVLv0_0),.din(w_dff_A_CMYqqWq50_0),.clk(gclk));
	jdff dff_A_qJosGXVx0_0(.dout(w_dff_A_CMYqqWq50_0),.din(w_dff_A_qJosGXVx0_0),.clk(gclk));
	jdff dff_A_yggG9FsL8_1(.dout(w_G283_3[1]),.din(w_dff_A_yggG9FsL8_1),.clk(gclk));
	jdff dff_A_nbD8OjSx0_1(.dout(w_dff_A_yggG9FsL8_1),.din(w_dff_A_nbD8OjSx0_1),.clk(gclk));
	jdff dff_A_sfpgrEtx3_1(.dout(w_dff_A_nbD8OjSx0_1),.din(w_dff_A_sfpgrEtx3_1),.clk(gclk));
	jdff dff_A_qEGcM8sZ4_1(.dout(w_dff_A_sfpgrEtx3_1),.din(w_dff_A_qEGcM8sZ4_1),.clk(gclk));
	jdff dff_A_xWkutRy76_0(.dout(w_G283_0[0]),.din(w_dff_A_xWkutRy76_0),.clk(gclk));
	jdff dff_A_o2zAMAZe0_0(.dout(w_dff_A_xWkutRy76_0),.din(w_dff_A_o2zAMAZe0_0),.clk(gclk));
	jdff dff_A_HFEcO3OZ4_0(.dout(w_dff_A_o2zAMAZe0_0),.din(w_dff_A_HFEcO3OZ4_0),.clk(gclk));
	jdff dff_A_ZXAphjHl9_1(.dout(w_G283_0[1]),.din(w_dff_A_ZXAphjHl9_1),.clk(gclk));
	jdff dff_A_kQ9ZolWv4_1(.dout(w_dff_A_ZXAphjHl9_1),.din(w_dff_A_kQ9ZolWv4_1),.clk(gclk));
	jdff dff_A_FRy2ruUc6_1(.dout(w_dff_A_kQ9ZolWv4_1),.din(w_dff_A_FRy2ruUc6_1),.clk(gclk));
	jdff dff_A_Lrq5l9tN6_2(.dout(w_n166_2[2]),.din(w_dff_A_Lrq5l9tN6_2),.clk(gclk));
	jdff dff_B_WGGkR6IG8_1(.din(n215),.dout(w_dff_B_WGGkR6IG8_1),.clk(gclk));
	jdff dff_A_TFuT86eL8_0(.dout(w_G200_1[0]),.din(w_dff_A_TFuT86eL8_0),.clk(gclk));
	jdff dff_A_D1ne4K4h6_0(.dout(w_dff_A_TFuT86eL8_0),.din(w_dff_A_D1ne4K4h6_0),.clk(gclk));
	jdff dff_A_sOPCTEl24_0(.dout(w_dff_A_D1ne4K4h6_0),.din(w_dff_A_sOPCTEl24_0),.clk(gclk));
	jdff dff_A_mXjksGXB1_0(.dout(w_dff_A_sOPCTEl24_0),.din(w_dff_A_mXjksGXB1_0),.clk(gclk));
	jdff dff_A_DQBLRFxv6_0(.dout(w_dff_A_mXjksGXB1_0),.din(w_dff_A_DQBLRFxv6_0),.clk(gclk));
	jdff dff_A_NMUsM9wm2_0(.dout(w_dff_A_DQBLRFxv6_0),.din(w_dff_A_NMUsM9wm2_0),.clk(gclk));
	jdff dff_A_YqcSp3Kl9_0(.dout(w_dff_A_NMUsM9wm2_0),.din(w_dff_A_YqcSp3Kl9_0),.clk(gclk));
	jdff dff_A_nM2frNaL4_1(.dout(w_G200_1[1]),.din(w_dff_A_nM2frNaL4_1),.clk(gclk));
	jdff dff_A_DmpEb5RY1_2(.dout(w_G200_0[2]),.din(w_dff_A_DmpEb5RY1_2),.clk(gclk));
	jdff dff_A_CCTZdFk07_2(.dout(w_dff_A_DmpEb5RY1_2),.din(w_dff_A_CCTZdFk07_2),.clk(gclk));
	jdff dff_A_PC7hCPp52_2(.dout(w_dff_A_CCTZdFk07_2),.din(w_dff_A_PC7hCPp52_2),.clk(gclk));
	jdff dff_A_lrrUXja13_2(.dout(w_dff_A_PC7hCPp52_2),.din(w_dff_A_lrrUXja13_2),.clk(gclk));
	jdff dff_A_KadsinUX2_2(.dout(w_dff_A_lrrUXja13_2),.din(w_dff_A_KadsinUX2_2),.clk(gclk));
	jdff dff_A_TkAhIzsv6_2(.dout(w_dff_A_KadsinUX2_2),.din(w_dff_A_TkAhIzsv6_2),.clk(gclk));
	jdff dff_A_qRkE6gDE0_2(.dout(w_dff_A_TkAhIzsv6_2),.din(w_dff_A_qRkE6gDE0_2),.clk(gclk));
	jdff dff_A_6bRW6Qnl2_0(.dout(w_G190_4[0]),.din(w_dff_A_6bRW6Qnl2_0),.clk(gclk));
	jdff dff_A_TcCrMEl05_0(.dout(w_G190_1[0]),.din(w_dff_A_TcCrMEl05_0),.clk(gclk));
	jdff dff_A_2ypiILTb6_0(.dout(w_dff_A_TcCrMEl05_0),.din(w_dff_A_2ypiILTb6_0),.clk(gclk));
	jdff dff_A_6NH8agMt2_0(.dout(w_dff_A_2ypiILTb6_0),.din(w_dff_A_6NH8agMt2_0),.clk(gclk));
	jdff dff_A_nw8f0R964_0(.dout(w_dff_A_6NH8agMt2_0),.din(w_dff_A_nw8f0R964_0),.clk(gclk));
	jdff dff_A_hrPLdJey5_0(.dout(w_G190_0[0]),.din(w_dff_A_hrPLdJey5_0),.clk(gclk));
	jdff dff_A_e5MdD5iH7_0(.dout(w_dff_A_hrPLdJey5_0),.din(w_dff_A_e5MdD5iH7_0),.clk(gclk));
	jdff dff_A_iEO4TAKl5_1(.dout(w_G190_0[1]),.din(w_dff_A_iEO4TAKl5_1),.clk(gclk));
	jdff dff_A_od4RnqI36_1(.dout(w_dff_A_iEO4TAKl5_1),.din(w_dff_A_od4RnqI36_1),.clk(gclk));
	jdff dff_A_J7ajIevY0_1(.dout(w_dff_A_od4RnqI36_1),.din(w_dff_A_J7ajIevY0_1),.clk(gclk));
	jdff dff_A_Qdhww1xq6_1(.dout(w_n214_0[1]),.din(w_dff_A_Qdhww1xq6_1),.clk(gclk));
	jdff dff_A_n7LAqGNU5_1(.dout(w_n213_0[1]),.din(w_dff_A_n7LAqGNU5_1),.clk(gclk));
	jdff dff_A_nBJU71419_0(.dout(w_n210_0[0]),.din(w_dff_A_nBJU71419_0),.clk(gclk));
	jdff dff_A_xlZw4z332_0(.dout(w_n205_0[0]),.din(w_dff_A_xlZw4z332_0),.clk(gclk));
	jdff dff_B_VCunKxQB3_2(.din(n205),.dout(w_dff_B_VCunKxQB3_2),.clk(gclk));
	jdff dff_A_yBIm5AGK6_0(.dout(w_n201_0[0]),.din(w_dff_A_yBIm5AGK6_0),.clk(gclk));
	jdff dff_A_RJ3ehxuJ6_2(.dout(w_G33_9[2]),.din(w_dff_A_RJ3ehxuJ6_2),.clk(gclk));
	jdff dff_A_dXo3rnxy2_1(.dout(w_n103_0[1]),.din(w_dff_A_dXo3rnxy2_1),.clk(gclk));
	jdff dff_A_Yu58xckM0_0(.dout(w_n196_2[0]),.din(w_dff_A_Yu58xckM0_0),.clk(gclk));
	jdff dff_A_5DkLtjcb4_1(.dout(w_n196_2[1]),.din(w_dff_A_5DkLtjcb4_1),.clk(gclk));
	jdff dff_A_jXJ1oX4K0_0(.dout(w_n196_0[0]),.din(w_dff_A_jXJ1oX4K0_0),.clk(gclk));
	jdff dff_A_vV1USWCc7_2(.dout(w_n196_0[2]),.din(w_dff_A_vV1USWCc7_2),.clk(gclk));
	jdff dff_B_8fRgtUxn3_3(.din(n196),.dout(w_dff_B_8fRgtUxn3_3),.clk(gclk));
	jdff dff_B_t0pyKXGU0_3(.din(w_dff_B_8fRgtUxn3_3),.dout(w_dff_B_t0pyKXGU0_3),.clk(gclk));
	jdff dff_B_aViKNqFt3_3(.din(w_dff_B_t0pyKXGU0_3),.dout(w_dff_B_aViKNqFt3_3),.clk(gclk));
	jdff dff_B_jUizMbAi8_3(.din(w_dff_B_aViKNqFt3_3),.dout(w_dff_B_jUizMbAi8_3),.clk(gclk));
	jdff dff_B_gHcHtbaM1_3(.din(w_dff_B_jUizMbAi8_3),.dout(w_dff_B_gHcHtbaM1_3),.clk(gclk));
	jdff dff_A_KMlib6jm0_0(.dout(w_G179_2[0]),.din(w_dff_A_KMlib6jm0_0),.clk(gclk));
	jdff dff_A_B2p8k5Fz8_0(.dout(w_dff_A_KMlib6jm0_0),.din(w_dff_A_B2p8k5Fz8_0),.clk(gclk));
	jdff dff_A_sCVs6zPD6_0(.dout(w_dff_A_B2p8k5Fz8_0),.din(w_dff_A_sCVs6zPD6_0),.clk(gclk));
	jdff dff_A_brn168q66_0(.dout(w_dff_A_sCVs6zPD6_0),.din(w_dff_A_brn168q66_0),.clk(gclk));
	jdff dff_A_3JfNc2cQ6_0(.dout(w_dff_A_brn168q66_0),.din(w_dff_A_3JfNc2cQ6_0),.clk(gclk));
	jdff dff_A_b5dhTsKc6_0(.dout(w_dff_A_3JfNc2cQ6_0),.din(w_dff_A_b5dhTsKc6_0),.clk(gclk));
	jdff dff_A_J9O08y4f3_0(.dout(w_dff_A_b5dhTsKc6_0),.din(w_dff_A_J9O08y4f3_0),.clk(gclk));
	jdff dff_A_Ogmw8Xod0_1(.dout(w_G179_2[1]),.din(w_dff_A_Ogmw8Xod0_1),.clk(gclk));
	jdff dff_A_S8rupHTl9_1(.dout(w_dff_A_Ogmw8Xod0_1),.din(w_dff_A_S8rupHTl9_1),.clk(gclk));
	jdff dff_A_Wd21yO0Q4_1(.dout(w_dff_A_S8rupHTl9_1),.din(w_dff_A_Wd21yO0Q4_1),.clk(gclk));
	jdff dff_A_OlEhyq3b3_1(.dout(w_dff_A_Wd21yO0Q4_1),.din(w_dff_A_OlEhyq3b3_1),.clk(gclk));
	jdff dff_A_oLA0qMKS8_1(.dout(w_dff_A_OlEhyq3b3_1),.din(w_dff_A_oLA0qMKS8_1),.clk(gclk));
	jdff dff_A_EmEmE86E6_1(.dout(w_dff_A_oLA0qMKS8_1),.din(w_dff_A_EmEmE86E6_1),.clk(gclk));
	jdff dff_A_Xfg6H6d67_1(.dout(w_dff_A_EmEmE86E6_1),.din(w_dff_A_Xfg6H6d67_1),.clk(gclk));
	jdff dff_A_YJh1HPjB0_0(.dout(w_G179_0[0]),.din(w_dff_A_YJh1HPjB0_0),.clk(gclk));
	jdff dff_A_tU4FM3tT9_0(.dout(w_dff_A_YJh1HPjB0_0),.din(w_dff_A_tU4FM3tT9_0),.clk(gclk));
	jdff dff_A_ccDNE53y1_0(.dout(w_dff_A_tU4FM3tT9_0),.din(w_dff_A_ccDNE53y1_0),.clk(gclk));
	jdff dff_A_lpebNB3R4_0(.dout(w_dff_A_ccDNE53y1_0),.din(w_dff_A_lpebNB3R4_0),.clk(gclk));
	jdff dff_A_WHln3AV55_0(.dout(w_dff_A_lpebNB3R4_0),.din(w_dff_A_WHln3AV55_0),.clk(gclk));
	jdff dff_A_XOhSyQFY7_0(.dout(w_dff_A_WHln3AV55_0),.din(w_dff_A_XOhSyQFY7_0),.clk(gclk));
	jdff dff_A_g2I0R6IE3_0(.dout(w_dff_A_XOhSyQFY7_0),.din(w_dff_A_g2I0R6IE3_0),.clk(gclk));
	jdff dff_B_wLkV8Msg4_0(.din(n192),.dout(w_dff_B_wLkV8Msg4_0),.clk(gclk));
	jdff dff_A_oUx6ewKo9_1(.dout(w_n190_1[1]),.din(w_dff_A_oUx6ewKo9_1),.clk(gclk));
	jdff dff_A_nNOwGfR79_0(.dout(w_n189_2[0]),.din(w_dff_A_nNOwGfR79_0),.clk(gclk));
	jdff dff_A_0ImIa9oz1_0(.dout(w_dff_A_nNOwGfR79_0),.din(w_dff_A_0ImIa9oz1_0),.clk(gclk));
	jdff dff_A_es4OKvcI0_2(.dout(w_n189_0[2]),.din(w_dff_A_es4OKvcI0_2),.clk(gclk));
	jdff dff_A_4rBuxrm07_0(.dout(w_n85_0[0]),.din(w_dff_A_4rBuxrm07_0),.clk(gclk));
	jdff dff_A_o5EKPjlR2_0(.dout(w_dff_A_4rBuxrm07_0),.din(w_dff_A_o5EKPjlR2_0),.clk(gclk));
	jdff dff_A_9VJYIO237_2(.dout(w_n85_0[2]),.din(w_dff_A_9VJYIO237_2),.clk(gclk));
	jdff dff_A_S0f0OtKf4_2(.dout(w_dff_A_9VJYIO237_2),.din(w_dff_A_S0f0OtKf4_2),.clk(gclk));
	jdff dff_A_5kn7p0kp0_2(.dout(w_dff_A_S0f0OtKf4_2),.din(w_dff_A_5kn7p0kp0_2),.clk(gclk));
	jdff dff_A_6naw0bNr9_2(.dout(w_dff_A_5kn7p0kp0_2),.din(w_dff_A_6naw0bNr9_2),.clk(gclk));
	jdff dff_A_ln2asg344_0(.dout(w_G20_5[0]),.din(w_dff_A_ln2asg344_0),.clk(gclk));
	jdff dff_A_FGDdilbX4_1(.dout(w_G20_5[1]),.din(w_dff_A_FGDdilbX4_1),.clk(gclk));
	jdff dff_A_JWPKIpRZ9_1(.dout(w_n80_0[1]),.din(w_dff_A_JWPKIpRZ9_1),.clk(gclk));
	jdff dff_A_vnfRPm0D1_1(.dout(w_dff_A_JWPKIpRZ9_1),.din(w_dff_A_vnfRPm0D1_1),.clk(gclk));
	jdff dff_A_6XzsJmGb0_1(.dout(w_dff_A_vnfRPm0D1_1),.din(w_dff_A_6XzsJmGb0_1),.clk(gclk));
	jdff dff_A_IVFQEA879_2(.dout(w_n80_0[2]),.din(w_dff_A_IVFQEA879_2),.clk(gclk));
	jdff dff_A_f9Vx7bTT7_2(.dout(w_dff_A_IVFQEA879_2),.din(w_dff_A_f9Vx7bTT7_2),.clk(gclk));
	jdff dff_A_C8ItDbhr4_2(.dout(w_dff_A_f9Vx7bTT7_2),.din(w_dff_A_C8ItDbhr4_2),.clk(gclk));
	jdff dff_A_JzOAiOhW1_2(.dout(w_dff_A_C8ItDbhr4_2),.din(w_dff_A_JzOAiOhW1_2),.clk(gclk));
	jdff dff_A_j1CPUTnK0_2(.dout(w_dff_A_JzOAiOhW1_2),.din(w_dff_A_j1CPUTnK0_2),.clk(gclk));
	jdff dff_A_QN1UTpGE1_2(.dout(w_G107_1[2]),.din(w_dff_A_QN1UTpGE1_2),.clk(gclk));
	jdff dff_A_IWIbbCRv4_2(.dout(w_dff_A_QN1UTpGE1_2),.din(w_dff_A_IWIbbCRv4_2),.clk(gclk));
	jdff dff_A_KLhsMzL80_2(.dout(w_dff_A_IWIbbCRv4_2),.din(w_dff_A_KLhsMzL80_2),.clk(gclk));
	jdff dff_A_o2dkQw2X6_1(.dout(w_G107_0[1]),.din(w_dff_A_o2dkQw2X6_1),.clk(gclk));
	jdff dff_A_Q72I1szT1_1(.dout(w_dff_A_o2dkQw2X6_1),.din(w_dff_A_Q72I1szT1_1),.clk(gclk));
	jdff dff_A_t00ToI546_1(.dout(w_dff_A_Q72I1szT1_1),.din(w_dff_A_t00ToI546_1),.clk(gclk));
	jdff dff_A_hzSNvali3_2(.dout(w_G107_0[2]),.din(w_dff_A_hzSNvali3_2),.clk(gclk));
	jdff dff_A_UQjn3JcF8_2(.dout(w_dff_A_hzSNvali3_2),.din(w_dff_A_UQjn3JcF8_2),.clk(gclk));
	jdff dff_A_5RDm4RVr9_2(.dout(w_dff_A_UQjn3JcF8_2),.din(w_dff_A_5RDm4RVr9_2),.clk(gclk));
	jdff dff_A_S8uciYKb7_0(.dout(w_n79_0[0]),.din(w_dff_A_S8uciYKb7_0),.clk(gclk));
	jdff dff_A_BmhYXBOh6_0(.dout(w_dff_A_S8uciYKb7_0),.din(w_dff_A_BmhYXBOh6_0),.clk(gclk));
	jdff dff_A_fbC376HG6_0(.dout(w_G97_5[0]),.din(w_dff_A_fbC376HG6_0),.clk(gclk));
	jdff dff_A_602sP49u2_1(.dout(w_n97_1[1]),.din(w_dff_A_602sP49u2_1),.clk(gclk));
	jdff dff_A_NBWhMjeI7_0(.dout(w_n97_0[0]),.din(w_dff_A_NBWhMjeI7_0),.clk(gclk));
	jdff dff_A_aExwiZ3Z6_0(.dout(w_G87_3[0]),.din(w_dff_A_aExwiZ3Z6_0),.clk(gclk));
	jdff dff_A_LbDMwrdX5_2(.dout(w_G87_3[2]),.din(w_dff_A_LbDMwrdX5_2),.clk(gclk));
	jdff dff_A_JtiMkx3W9_2(.dout(w_dff_A_LbDMwrdX5_2),.din(w_dff_A_JtiMkx3W9_2),.clk(gclk));
	jdff dff_A_s2DAGwOv7_2(.dout(w_dff_A_JtiMkx3W9_2),.din(w_dff_A_s2DAGwOv7_2),.clk(gclk));
	jdff dff_A_GWoSYVQn1_0(.dout(w_G87_0[0]),.din(w_dff_A_GWoSYVQn1_0),.clk(gclk));
	jdff dff_A_W6NPhmPO4_0(.dout(w_dff_A_GWoSYVQn1_0),.din(w_dff_A_W6NPhmPO4_0),.clk(gclk));
	jdff dff_A_Ngq5RurS5_0(.dout(w_dff_A_W6NPhmPO4_0),.din(w_dff_A_Ngq5RurS5_0),.clk(gclk));
	jdff dff_A_v1DIj67w8_1(.dout(w_n179_0[1]),.din(w_dff_A_v1DIj67w8_1),.clk(gclk));
	jdff dff_A_aLKewj3f7_1(.dout(w_dff_A_v1DIj67w8_1),.din(w_dff_A_aLKewj3f7_1),.clk(gclk));
	jdff dff_A_81DlHO2N5_2(.dout(w_n179_0[2]),.din(w_dff_A_81DlHO2N5_2),.clk(gclk));
	jdff dff_A_ldhGD3Gr7_2(.dout(w_dff_A_81DlHO2N5_2),.din(w_dff_A_ldhGD3Gr7_2),.clk(gclk));
	jdff dff_A_oio6ptqe1_2(.dout(w_n112_5[2]),.din(w_dff_A_oio6ptqe1_2),.clk(gclk));
	jdff dff_A_Xs3u2aA27_1(.dout(w_G20_2[1]),.din(w_dff_A_Xs3u2aA27_1),.clk(gclk));
	jdff dff_A_sVih4rfd4_0(.dout(w_G68_4[0]),.din(w_dff_A_sVih4rfd4_0),.clk(gclk));
	jdff dff_A_BiYpS19j7_1(.dout(w_G68_4[1]),.din(w_dff_A_BiYpS19j7_1),.clk(gclk));
	jdff dff_A_EXr1nqMF9_0(.dout(w_G68_1[0]),.din(w_dff_A_EXr1nqMF9_0),.clk(gclk));
	jdff dff_A_ybmlZtvC9_2(.dout(w_G68_1[2]),.din(w_dff_A_ybmlZtvC9_2),.clk(gclk));
	jdff dff_A_VQfRxLjO4_2(.dout(w_dff_A_ybmlZtvC9_2),.din(w_dff_A_VQfRxLjO4_2),.clk(gclk));
	jdff dff_A_wdiVNzGw5_2(.dout(w_dff_A_VQfRxLjO4_2),.din(w_dff_A_wdiVNzGw5_2),.clk(gclk));
	jdff dff_A_O2WVEmuP0_2(.dout(w_dff_A_wdiVNzGw5_2),.din(w_dff_A_O2WVEmuP0_2),.clk(gclk));
	jdff dff_A_nJpYmbT09_2(.dout(w_G68_0[2]),.din(w_dff_A_nJpYmbT09_2),.clk(gclk));
	jdff dff_A_7iLGToeL6_1(.dout(w_n148_8[1]),.din(w_dff_A_7iLGToeL6_1),.clk(gclk));
	jdff dff_A_N9Azsqpu1_0(.dout(w_G20_6[0]),.din(w_dff_A_N9Azsqpu1_0),.clk(gclk));
	jdff dff_A_gKX85fBz5_2(.dout(w_G20_1[2]),.din(w_dff_A_gKX85fBz5_2),.clk(gclk));
	jdff dff_A_U7WxENXP3_0(.dout(w_G20_0[0]),.din(w_dff_A_U7WxENXP3_0),.clk(gclk));
	jdff dff_B_hMBDDOzB3_2(.din(n172),.dout(w_dff_B_hMBDDOzB3_2),.clk(gclk));
	jdff dff_B_Mf2fnBMK2_2(.din(w_dff_B_hMBDDOzB3_2),.dout(w_dff_B_Mf2fnBMK2_2),.clk(gclk));
	jdff dff_A_Q9teBhin7_0(.dout(w_G97_4[0]),.din(w_dff_A_Q9teBhin7_0),.clk(gclk));
	jdff dff_A_Rwdh5tfI4_0(.dout(w_dff_A_Q9teBhin7_0),.din(w_dff_A_Rwdh5tfI4_0),.clk(gclk));
	jdff dff_A_mP813Pcd7_0(.dout(w_dff_A_Rwdh5tfI4_0),.din(w_dff_A_mP813Pcd7_0),.clk(gclk));
	jdff dff_A_cCjyevy15_2(.dout(w_G97_1[2]),.din(w_dff_A_cCjyevy15_2),.clk(gclk));
	jdff dff_A_NGRSvjyA2_2(.dout(w_dff_A_cCjyevy15_2),.din(w_dff_A_NGRSvjyA2_2),.clk(gclk));
	jdff dff_A_hupm6H9s3_2(.dout(w_dff_A_NGRSvjyA2_2),.din(w_dff_A_hupm6H9s3_2),.clk(gclk));
	jdff dff_A_qFESAoza9_2(.dout(w_dff_A_hupm6H9s3_2),.din(w_dff_A_qFESAoza9_2),.clk(gclk));
	jdff dff_A_bh8X36zm6_1(.dout(w_G97_0[1]),.din(w_dff_A_bh8X36zm6_1),.clk(gclk));
	jdff dff_A_rAs9fs752_1(.dout(w_dff_A_bh8X36zm6_1),.din(w_dff_A_rAs9fs752_1),.clk(gclk));
	jdff dff_A_zFlKy9Tf6_1(.dout(w_dff_A_rAs9fs752_1),.din(w_dff_A_zFlKy9Tf6_1),.clk(gclk));
	jdff dff_A_37h6aHQw9_2(.dout(w_G97_0[2]),.din(w_dff_A_37h6aHQw9_2),.clk(gclk));
	jdff dff_A_RIYLDndJ8_0(.dout(w_G33_10[0]),.din(w_dff_A_RIYLDndJ8_0),.clk(gclk));
	jdff dff_A_Hdd3lQoJ9_1(.dout(w_G33_10[1]),.din(w_dff_A_Hdd3lQoJ9_1),.clk(gclk));
	jdff dff_A_OEIpwxEF5_0(.dout(w_n170_0[0]),.din(w_dff_A_OEIpwxEF5_0),.clk(gclk));
	jdff dff_B_c3EoQMcj3_0(.din(n169),.dout(w_dff_B_c3EoQMcj3_0),.clk(gclk));
	jdff dff_A_F9yCgSqd8_0(.dout(w_G274_0[0]),.din(w_dff_A_F9yCgSqd8_0),.clk(gclk));
	jdff dff_A_vFfXoTgA4_0(.dout(w_dff_A_F9yCgSqd8_0),.din(w_dff_A_vFfXoTgA4_0),.clk(gclk));
	jdff dff_A_LfpceVR85_0(.dout(w_dff_A_vFfXoTgA4_0),.din(w_dff_A_LfpceVR85_0),.clk(gclk));
	jdff dff_A_Z8i083sN4_2(.dout(w_G274_0[2]),.din(w_dff_A_Z8i083sN4_2),.clk(gclk));
	jdff dff_A_wNbrbeh79_2(.dout(w_dff_A_Z8i083sN4_2),.din(w_dff_A_wNbrbeh79_2),.clk(gclk));
	jdff dff_A_JZDmjjWv3_0(.dout(w_n166_3[0]),.din(w_dff_A_JZDmjjWv3_0),.clk(gclk));
	jdff dff_B_sfNk1m3n4_0(.din(n165),.dout(w_dff_B_sfNk1m3n4_0),.clk(gclk));
	jdff dff_A_sflOr6SE6_2(.dout(w_n115_0[2]),.din(w_dff_A_sflOr6SE6_2),.clk(gclk));
	jdff dff_A_FHTOnRU44_0(.dout(w_n114_1[0]),.din(w_dff_A_FHTOnRU44_0),.clk(gclk));
	jdff dff_A_ruaDa1ua8_1(.dout(w_n114_0[1]),.din(w_dff_A_ruaDa1ua8_1),.clk(gclk));
	jdff dff_A_plqwpa2X5_0(.dout(w_n163_0[0]),.din(w_dff_A_plqwpa2X5_0),.clk(gclk));
	jdff dff_A_MIU4X5zD8_2(.dout(w_n161_0[2]),.din(w_dff_A_MIU4X5zD8_2),.clk(gclk));
	jdff dff_A_O4SyOYIf4_2(.dout(w_dff_A_MIU4X5zD8_2),.din(w_dff_A_O4SyOYIf4_2),.clk(gclk));
	jdff dff_A_AkNA0WSt5_2(.dout(w_dff_A_O4SyOYIf4_2),.din(w_dff_A_AkNA0WSt5_2),.clk(gclk));
	jdff dff_A_GjEuVDQb9_0(.dout(w_G45_1[0]),.din(w_dff_A_GjEuVDQb9_0),.clk(gclk));
	jdff dff_A_Gg30chY37_0(.dout(w_dff_A_GjEuVDQb9_0),.din(w_dff_A_Gg30chY37_0),.clk(gclk));
	jdff dff_A_zAnPpuHg8_1(.dout(w_G45_1[1]),.din(w_dff_A_zAnPpuHg8_1),.clk(gclk));
	jdff dff_A_YAkzqEdY8_1(.dout(w_G45_0[1]),.din(w_dff_A_YAkzqEdY8_1),.clk(gclk));
	jdff dff_A_hz0rqOpc4_1(.dout(w_dff_A_YAkzqEdY8_1),.din(w_dff_A_hz0rqOpc4_1),.clk(gclk));
	jdff dff_A_O7RBQmC53_1(.dout(w_dff_A_hz0rqOpc4_1),.din(w_dff_A_O7RBQmC53_1),.clk(gclk));
	jdff dff_A_ZqoXkDEg9_2(.dout(w_G45_0[2]),.din(w_dff_A_ZqoXkDEg9_2),.clk(gclk));
	jdff dff_A_MWBJbelM4_2(.dout(w_dff_A_ZqoXkDEg9_2),.din(w_dff_A_MWBJbelM4_2),.clk(gclk));
	jdff dff_A_mlsnI8yO0_2(.dout(w_dff_A_MWBJbelM4_2),.din(w_dff_A_mlsnI8yO0_2),.clk(gclk));
	jdff dff_A_wnamHytM4_0(.dout(w_n98_1[0]),.din(w_dff_A_wnamHytM4_0),.clk(gclk));
	jdff dff_A_Nhy7Pxuv0_1(.dout(w_n98_1[1]),.din(w_dff_A_Nhy7Pxuv0_1),.clk(gclk));
	jdff dff_A_y1kiTWae9_0(.dout(w_G250_0[0]),.din(w_dff_A_y1kiTWae9_0),.clk(gclk));
	jdff dff_A_WgYvqrS63_0(.dout(w_dff_A_y1kiTWae9_0),.din(w_dff_A_WgYvqrS63_0),.clk(gclk));
	jdff dff_A_vVsBMaPY2_1(.dout(w_G250_0[1]),.din(w_dff_A_vVsBMaPY2_1),.clk(gclk));
	jdff dff_A_72UFADII8_1(.dout(w_dff_A_vVsBMaPY2_1),.din(w_dff_A_72UFADII8_1),.clk(gclk));
	jdff dff_B_CvdKY4r86_1(.din(n153),.dout(w_dff_B_CvdKY4r86_1),.clk(gclk));
	jdff dff_A_Lqeye15K4_0(.dout(w_n157_0[0]),.din(w_dff_A_Lqeye15K4_0),.clk(gclk));
	jdff dff_A_IC5fUeBa9_0(.dout(w_dff_A_Lqeye15K4_0),.din(w_dff_A_IC5fUeBa9_0),.clk(gclk));
	jdff dff_A_Jqq4jghV2_2(.dout(w_n157_0[2]),.din(w_dff_A_Jqq4jghV2_2),.clk(gclk));
	jdff dff_A_mjO8ion64_2(.dout(w_dff_A_Jqq4jghV2_2),.din(w_dff_A_mjO8ion64_2),.clk(gclk));
	jdff dff_A_N71CIgGb6_1(.dout(w_G116_1[1]),.din(w_dff_A_N71CIgGb6_1),.clk(gclk));
	jdff dff_A_x1gD1Ai78_1(.dout(w_dff_A_N71CIgGb6_1),.din(w_dff_A_x1gD1Ai78_1),.clk(gclk));
	jdff dff_A_wubsV4sU3_1(.dout(w_dff_A_x1gD1Ai78_1),.din(w_dff_A_wubsV4sU3_1),.clk(gclk));
	jdff dff_A_bxeGtGKh1_2(.dout(w_G116_1[2]),.din(w_dff_A_bxeGtGKh1_2),.clk(gclk));
	jdff dff_A_kCRtpCFN6_2(.dout(w_dff_A_bxeGtGKh1_2),.din(w_dff_A_kCRtpCFN6_2),.clk(gclk));
	jdff dff_A_0FigtYqf8_2(.dout(w_dff_A_kCRtpCFN6_2),.din(w_dff_A_0FigtYqf8_2),.clk(gclk));
	jdff dff_A_7N9VqluI2_1(.dout(w_G116_0[1]),.din(w_dff_A_7N9VqluI2_1),.clk(gclk));
	jdff dff_A_lPXlGRsb0_1(.dout(w_dff_A_7N9VqluI2_1),.din(w_dff_A_lPXlGRsb0_1),.clk(gclk));
	jdff dff_A_QBQC4kG27_1(.dout(w_dff_A_lPXlGRsb0_1),.din(w_dff_A_QBQC4kG27_1),.clk(gclk));
	jdff dff_A_8pOBQB5E3_2(.dout(w_G116_0[2]),.din(w_dff_A_8pOBQB5E3_2),.clk(gclk));
	jdff dff_A_Uj6RaHaN7_0(.dout(w_G238_1[0]),.din(w_dff_A_Uj6RaHaN7_0),.clk(gclk));
	jdff dff_A_SKieoeJM9_0(.dout(w_dff_A_Uj6RaHaN7_0),.din(w_dff_A_SKieoeJM9_0),.clk(gclk));
	jdff dff_A_jcx56kjk5_1(.dout(w_G238_0[1]),.din(w_dff_A_jcx56kjk5_1),.clk(gclk));
	jdff dff_A_Rb6IF7670_1(.dout(w_dff_A_jcx56kjk5_1),.din(w_dff_A_Rb6IF7670_1),.clk(gclk));
	jdff dff_A_tI7E6PyX4_1(.dout(w_dff_A_Rb6IF7670_1),.din(w_dff_A_tI7E6PyX4_1),.clk(gclk));
	jdff dff_A_M9xudvUV9_1(.dout(w_dff_A_tI7E6PyX4_1),.din(w_dff_A_M9xudvUV9_1),.clk(gclk));
	jdff dff_A_2x8NneIi5_2(.dout(w_G238_0[2]),.din(w_dff_A_2x8NneIi5_2),.clk(gclk));
	jdff dff_A_zG3jJkC47_2(.dout(w_dff_A_2x8NneIi5_2),.din(w_dff_A_zG3jJkC47_2),.clk(gclk));
	jdff dff_A_eZH5iZ0n7_2(.dout(w_G1698_0[2]),.din(w_dff_A_eZH5iZ0n7_2),.clk(gclk));
	jdff dff_A_eXpKzxeD8_0(.dout(w_G244_1[0]),.din(w_dff_A_eXpKzxeD8_0),.clk(gclk));
	jdff dff_A_XaWl6EhB4_0(.dout(w_dff_A_eXpKzxeD8_0),.din(w_dff_A_XaWl6EhB4_0),.clk(gclk));
	jdff dff_A_X4sKCKie2_1(.dout(w_G244_0[1]),.din(w_dff_A_X4sKCKie2_1),.clk(gclk));
	jdff dff_A_Bbp2fDwr8_1(.dout(w_dff_A_X4sKCKie2_1),.din(w_dff_A_Bbp2fDwr8_1),.clk(gclk));
	jdff dff_A_pBzLVghr5_1(.dout(w_dff_A_Bbp2fDwr8_1),.din(w_dff_A_pBzLVghr5_1),.clk(gclk));
	jdff dff_A_FjTqQqIS7_1(.dout(w_dff_A_pBzLVghr5_1),.din(w_dff_A_FjTqQqIS7_1),.clk(gclk));
	jdff dff_A_NQqXkoGO5_2(.dout(w_G244_0[2]),.din(w_dff_A_NQqXkoGO5_2),.clk(gclk));
	jdff dff_A_RKxoHzft5_2(.dout(w_dff_A_NQqXkoGO5_2),.din(w_dff_A_RKxoHzft5_2),.clk(gclk));
	jdff dff_A_Zu2QdsRX7_2(.dout(w_n151_4[2]),.din(w_dff_A_Zu2QdsRX7_2),.clk(gclk));
	jdff dff_A_MvEArPr95_2(.dout(w_dff_A_Zu2QdsRX7_2),.din(w_dff_A_MvEArPr95_2),.clk(gclk));
	jdff dff_A_lhwi2Cs43_1(.dout(w_n151_1[1]),.din(w_dff_A_lhwi2Cs43_1),.clk(gclk));
	jdff dff_A_qojIAw5P2_1(.dout(w_dff_A_lhwi2Cs43_1),.din(w_dff_A_qojIAw5P2_1),.clk(gclk));
	jdff dff_A_lMIT5JCa7_2(.dout(w_n151_1[2]),.din(w_dff_A_lMIT5JCa7_2),.clk(gclk));
	jdff dff_A_LQBuzSCm1_2(.dout(w_dff_A_lMIT5JCa7_2),.din(w_dff_A_LQBuzSCm1_2),.clk(gclk));
	jdff dff_A_guEi5ejR3_1(.dout(w_n151_0[1]),.din(w_dff_A_guEi5ejR3_1),.clk(gclk));
	jdff dff_A_TQ9Ulg3a7_1(.dout(w_dff_A_guEi5ejR3_1),.din(w_dff_A_TQ9Ulg3a7_1),.clk(gclk));
	jdff dff_A_SOrcP7xY6_0(.dout(w_n149_2[0]),.din(w_dff_A_SOrcP7xY6_0),.clk(gclk));
	jdff dff_A_imXvUDCW9_1(.dout(w_G41_0[1]),.din(w_dff_A_imXvUDCW9_1),.clk(gclk));
	jdff dff_A_eAWEYyPb0_2(.dout(w_G41_0[2]),.din(w_dff_A_eAWEYyPb0_2),.clk(gclk));
	jdff dff_A_bIepQwPZ9_2(.dout(w_dff_A_eAWEYyPb0_2),.din(w_dff_A_bIepQwPZ9_2),.clk(gclk));
	jdff dff_A_ztKs9EU99_2(.dout(w_G33_3[2]),.din(w_dff_A_ztKs9EU99_2),.clk(gclk));
	jdff dff_A_emGDu4J31_2(.dout(w_dff_A_ztKs9EU99_2),.din(w_dff_A_emGDu4J31_2),.clk(gclk));
	jdff dff_A_HBy6B4246_2(.dout(w_dff_A_emGDu4J31_2),.din(w_dff_A_HBy6B4246_2),.clk(gclk));
	jdff dff_A_qDRWEKsA1_2(.dout(w_dff_A_HBy6B4246_2),.din(w_dff_A_qDRWEKsA1_2),.clk(gclk));
	jdff dff_A_YKI0fE2C8_2(.dout(w_dff_A_qDRWEKsA1_2),.din(w_dff_A_YKI0fE2C8_2),.clk(gclk));
	jdff dff_A_L884xvOs1_0(.dout(w_G33_0[0]),.din(w_dff_A_L884xvOs1_0),.clk(gclk));
	jdff dff_A_Zcca7dj56_1(.dout(w_n147_0[1]),.din(w_dff_A_Zcca7dj56_1),.clk(gclk));
	jdff dff_A_gOULqPpa3_2(.dout(w_n147_0[2]),.din(w_dff_A_gOULqPpa3_2),.clk(gclk));
	jdff dff_A_ojIQhcSW4_1(.dout(w_G13_0[1]),.din(w_dff_A_ojIQhcSW4_1),.clk(gclk));
	jdff dff_A_U5T40sHc3_2(.dout(w_G13_0[2]),.din(w_dff_A_U5T40sHc3_2),.clk(gclk));
	jdff dff_A_zTZXqXCx5_2(.dout(w_dff_A_U5T40sHc3_2),.din(w_dff_A_zTZXqXCx5_2),.clk(gclk));
	jdff dff_A_IexZa1a62_0(.dout(w_G1_2[0]),.din(w_dff_A_IexZa1a62_0),.clk(gclk));
	jdff dff_A_NB7BrxW80_2(.dout(w_G1_2[2]),.din(w_dff_A_NB7BrxW80_2),.clk(gclk));
	jdff dff_A_M6s2GyiG1_0(.dout(w_G1_0[0]),.din(w_dff_A_M6s2GyiG1_0),.clk(gclk));
	jdff dff_A_cSmSc4Xu5_1(.dout(w_n146_0[1]),.din(w_dff_A_cSmSc4Xu5_1),.clk(gclk));
	jdff dff_A_KHhMTtkU8_1(.dout(w_dff_A_cSmSc4Xu5_1),.din(w_dff_A_KHhMTtkU8_1),.clk(gclk));
	jdff dff_A_yrPrpbg44_1(.dout(w_dff_A_KHhMTtkU8_1),.din(w_dff_A_yrPrpbg44_1),.clk(gclk));
	jdff dff_A_UuUqAC6S6_1(.dout(w_dff_A_yrPrpbg44_1),.din(w_dff_A_UuUqAC6S6_1),.clk(gclk));
	jdff dff_A_GvZz6AZU1_1(.dout(w_dff_A_UuUqAC6S6_1),.din(w_dff_A_GvZz6AZU1_1),.clk(gclk));
	jdff dff_A_aWjUpErp0_1(.dout(w_dff_A_GvZz6AZU1_1),.din(w_dff_A_aWjUpErp0_1),.clk(gclk));
	jdff dff_A_j9RaDmuA2_2(.dout(w_n146_0[2]),.din(w_dff_A_j9RaDmuA2_2),.clk(gclk));
	jdff dff_A_w5GE8PKU8_2(.dout(w_dff_A_j9RaDmuA2_2),.din(w_dff_A_w5GE8PKU8_2),.clk(gclk));
	jdff dff_A_wKI40e3k2_2(.dout(w_dff_A_w5GE8PKU8_2),.din(w_dff_A_wKI40e3k2_2),.clk(gclk));
	jdff dff_A_gkHTHtTR2_2(.dout(w_dff_A_wKI40e3k2_2),.din(w_dff_A_gkHTHtTR2_2),.clk(gclk));
	jdff dff_A_HzDq4ZSw5_2(.dout(w_dff_A_gkHTHtTR2_2),.din(w_dff_A_HzDq4ZSw5_2),.clk(gclk));
	jdff dff_A_EF4gWOik0_2(.dout(w_dff_A_HzDq4ZSw5_2),.din(w_dff_A_EF4gWOik0_2),.clk(gclk));
	jdff dff_A_Z9Ua2TPN8_0(.dout(w_G169_1[0]),.din(w_dff_A_Z9Ua2TPN8_0),.clk(gclk));
	jdff dff_A_mwPkPso39_0(.dout(w_dff_A_Z9Ua2TPN8_0),.din(w_dff_A_mwPkPso39_0),.clk(gclk));
	jdff dff_A_yOV1ySzR8_0(.dout(w_dff_A_mwPkPso39_0),.din(w_dff_A_yOV1ySzR8_0),.clk(gclk));
	jdff dff_A_F4uQ5KSq5_0(.dout(w_dff_A_yOV1ySzR8_0),.din(w_dff_A_F4uQ5KSq5_0),.clk(gclk));
	jdff dff_A_uAtBLhjT8_0(.dout(w_dff_A_F4uQ5KSq5_0),.din(w_dff_A_uAtBLhjT8_0),.clk(gclk));
	jdff dff_A_Q10g6KuD1_0(.dout(w_dff_A_uAtBLhjT8_0),.din(w_dff_A_Q10g6KuD1_0),.clk(gclk));
	jdff dff_A_0eQoAOf32_0(.dout(w_dff_A_Q10g6KuD1_0),.din(w_dff_A_0eQoAOf32_0),.clk(gclk));
	jdff dff_A_soBXMpL87_1(.dout(w_G169_0[1]),.din(w_dff_A_soBXMpL87_1),.clk(gclk));
	jdff dff_A_0Itur3Zy0_1(.dout(w_dff_A_soBXMpL87_1),.din(w_dff_A_0Itur3Zy0_1),.clk(gclk));
	jdff dff_A_WTVt3mkB8_1(.dout(w_dff_A_0Itur3Zy0_1),.din(w_dff_A_WTVt3mkB8_1),.clk(gclk));
	jdff dff_A_raZPFetv9_1(.dout(w_dff_A_WTVt3mkB8_1),.din(w_dff_A_raZPFetv9_1),.clk(gclk));
	jdff dff_A_jSs7c7wO4_1(.dout(w_dff_A_raZPFetv9_1),.din(w_dff_A_jSs7c7wO4_1),.clk(gclk));
	jdff dff_A_JtQve0o20_1(.dout(w_dff_A_jSs7c7wO4_1),.din(w_dff_A_JtQve0o20_1),.clk(gclk));
	jdff dff_A_tbnSXAeN5_1(.dout(w_dff_A_JtQve0o20_1),.din(w_dff_A_tbnSXAeN5_1),.clk(gclk));
	jdff dff_A_cXLjNAtl1_2(.dout(w_G169_0[2]),.din(w_dff_A_cXLjNAtl1_2),.clk(gclk));
	jdff dff_A_cjRJxW1x0_2(.dout(w_dff_A_cXLjNAtl1_2),.din(w_dff_A_cjRJxW1x0_2),.clk(gclk));
	jdff dff_A_tGIt2dJ92_2(.dout(w_dff_A_cjRJxW1x0_2),.din(w_dff_A_tGIt2dJ92_2),.clk(gclk));
	jdff dff_A_9yVzYEyV9_2(.dout(w_dff_A_tGIt2dJ92_2),.din(w_dff_A_9yVzYEyV9_2),.clk(gclk));
	jdff dff_A_pnsng7Im4_2(.dout(w_dff_A_9yVzYEyV9_2),.din(w_dff_A_pnsng7Im4_2),.clk(gclk));
	jdff dff_A_2DD56qok2_2(.dout(w_dff_A_pnsng7Im4_2),.din(w_dff_A_2DD56qok2_2),.clk(gclk));
	jdff dff_A_gYcfZmMb5_2(.dout(w_dff_A_2DD56qok2_2),.din(w_dff_A_gYcfZmMb5_2),.clk(gclk));
	jdff dff_A_9UgON85M6_2(.dout(w_dff_A_UX4Td7kW7_0),.din(w_dff_A_9UgON85M6_2),.clk(gclk));
	jdff dff_A_UX4Td7kW7_0(.dout(w_dff_A_BftYGRw05_0),.din(w_dff_A_UX4Td7kW7_0),.clk(gclk));
	jdff dff_A_BftYGRw05_0(.dout(w_dff_A_jnQOSjw22_0),.din(w_dff_A_BftYGRw05_0),.clk(gclk));
	jdff dff_A_jnQOSjw22_0(.dout(w_dff_A_zq8GjPoa7_0),.din(w_dff_A_jnQOSjw22_0),.clk(gclk));
	jdff dff_A_zq8GjPoa7_0(.dout(w_dff_A_UkQKU8MN8_0),.din(w_dff_A_zq8GjPoa7_0),.clk(gclk));
	jdff dff_A_UkQKU8MN8_0(.dout(w_dff_A_iZ0swn2t3_0),.din(w_dff_A_UkQKU8MN8_0),.clk(gclk));
	jdff dff_A_iZ0swn2t3_0(.dout(w_dff_A_YmiDJlxs6_0),.din(w_dff_A_iZ0swn2t3_0),.clk(gclk));
	jdff dff_A_YmiDJlxs6_0(.dout(w_dff_A_twUMrmTp5_0),.din(w_dff_A_YmiDJlxs6_0),.clk(gclk));
	jdff dff_A_twUMrmTp5_0(.dout(w_dff_A_QGh853AF7_0),.din(w_dff_A_twUMrmTp5_0),.clk(gclk));
	jdff dff_A_QGh853AF7_0(.dout(w_dff_A_4vmu8yGq9_0),.din(w_dff_A_QGh853AF7_0),.clk(gclk));
	jdff dff_A_4vmu8yGq9_0(.dout(w_dff_A_lLTWS1Wl1_0),.din(w_dff_A_4vmu8yGq9_0),.clk(gclk));
	jdff dff_A_lLTWS1Wl1_0(.dout(w_dff_A_mwubIDYI7_0),.din(w_dff_A_lLTWS1Wl1_0),.clk(gclk));
	jdff dff_A_mwubIDYI7_0(.dout(w_dff_A_5aDZiB8w5_0),.din(w_dff_A_mwubIDYI7_0),.clk(gclk));
	jdff dff_A_5aDZiB8w5_0(.dout(w_dff_A_j6Y7nI6U2_0),.din(w_dff_A_5aDZiB8w5_0),.clk(gclk));
	jdff dff_A_j6Y7nI6U2_0(.dout(w_dff_A_pGiHP5Wr6_0),.din(w_dff_A_j6Y7nI6U2_0),.clk(gclk));
	jdff dff_A_pGiHP5Wr6_0(.dout(w_dff_A_68XgBR0N1_0),.din(w_dff_A_pGiHP5Wr6_0),.clk(gclk));
	jdff dff_A_68XgBR0N1_0(.dout(w_dff_A_KOoupgFN8_0),.din(w_dff_A_68XgBR0N1_0),.clk(gclk));
	jdff dff_A_KOoupgFN8_0(.dout(w_dff_A_bwYMGR4O4_0),.din(w_dff_A_KOoupgFN8_0),.clk(gclk));
	jdff dff_A_bwYMGR4O4_0(.dout(w_dff_A_JPlebdm77_0),.din(w_dff_A_bwYMGR4O4_0),.clk(gclk));
	jdff dff_A_JPlebdm77_0(.dout(w_dff_A_qX5tQoTy3_0),.din(w_dff_A_JPlebdm77_0),.clk(gclk));
	jdff dff_A_qX5tQoTy3_0(.dout(w_dff_A_IQsoLb6z3_0),.din(w_dff_A_qX5tQoTy3_0),.clk(gclk));
	jdff dff_A_IQsoLb6z3_0(.dout(w_dff_A_i8MqfCfC3_0),.din(w_dff_A_IQsoLb6z3_0),.clk(gclk));
	jdff dff_A_i8MqfCfC3_0(.dout(w_dff_A_tugXxbQl4_0),.din(w_dff_A_i8MqfCfC3_0),.clk(gclk));
	jdff dff_A_tugXxbQl4_0(.dout(w_dff_A_7LtWy9ON6_0),.din(w_dff_A_tugXxbQl4_0),.clk(gclk));
	jdff dff_A_7LtWy9ON6_0(.dout(G353),.din(w_dff_A_7LtWy9ON6_0),.clk(gclk));
	jdff dff_A_VGKJsJxE9_1(.dout(w_dff_A_ig4PozfA5_0),.din(w_dff_A_VGKJsJxE9_1),.clk(gclk));
	jdff dff_A_ig4PozfA5_0(.dout(w_dff_A_uzwQkORy9_0),.din(w_dff_A_ig4PozfA5_0),.clk(gclk));
	jdff dff_A_uzwQkORy9_0(.dout(w_dff_A_3ALl68WS6_0),.din(w_dff_A_uzwQkORy9_0),.clk(gclk));
	jdff dff_A_3ALl68WS6_0(.dout(w_dff_A_V35gbC4i6_0),.din(w_dff_A_3ALl68WS6_0),.clk(gclk));
	jdff dff_A_V35gbC4i6_0(.dout(w_dff_A_tCxKm7xA9_0),.din(w_dff_A_V35gbC4i6_0),.clk(gclk));
	jdff dff_A_tCxKm7xA9_0(.dout(w_dff_A_t6XBcfqj6_0),.din(w_dff_A_tCxKm7xA9_0),.clk(gclk));
	jdff dff_A_t6XBcfqj6_0(.dout(w_dff_A_xL0zm0Fl5_0),.din(w_dff_A_t6XBcfqj6_0),.clk(gclk));
	jdff dff_A_xL0zm0Fl5_0(.dout(w_dff_A_nJAOgdCd9_0),.din(w_dff_A_xL0zm0Fl5_0),.clk(gclk));
	jdff dff_A_nJAOgdCd9_0(.dout(w_dff_A_FrnaEkXg9_0),.din(w_dff_A_nJAOgdCd9_0),.clk(gclk));
	jdff dff_A_FrnaEkXg9_0(.dout(w_dff_A_6fqnp5KR3_0),.din(w_dff_A_FrnaEkXg9_0),.clk(gclk));
	jdff dff_A_6fqnp5KR3_0(.dout(w_dff_A_ce7h9YRo9_0),.din(w_dff_A_6fqnp5KR3_0),.clk(gclk));
	jdff dff_A_ce7h9YRo9_0(.dout(w_dff_A_zNDDkFbe2_0),.din(w_dff_A_ce7h9YRo9_0),.clk(gclk));
	jdff dff_A_zNDDkFbe2_0(.dout(w_dff_A_fVPSZAq72_0),.din(w_dff_A_zNDDkFbe2_0),.clk(gclk));
	jdff dff_A_fVPSZAq72_0(.dout(w_dff_A_I5PU5NZb9_0),.din(w_dff_A_fVPSZAq72_0),.clk(gclk));
	jdff dff_A_I5PU5NZb9_0(.dout(w_dff_A_jUbTQsvT2_0),.din(w_dff_A_I5PU5NZb9_0),.clk(gclk));
	jdff dff_A_jUbTQsvT2_0(.dout(w_dff_A_N3xBY6Le3_0),.din(w_dff_A_jUbTQsvT2_0),.clk(gclk));
	jdff dff_A_N3xBY6Le3_0(.dout(w_dff_A_pNbxZHaQ8_0),.din(w_dff_A_N3xBY6Le3_0),.clk(gclk));
	jdff dff_A_pNbxZHaQ8_0(.dout(w_dff_A_xwMGWpNP1_0),.din(w_dff_A_pNbxZHaQ8_0),.clk(gclk));
	jdff dff_A_xwMGWpNP1_0(.dout(w_dff_A_414Rv4rQ6_0),.din(w_dff_A_xwMGWpNP1_0),.clk(gclk));
	jdff dff_A_414Rv4rQ6_0(.dout(w_dff_A_uY7Sf3477_0),.din(w_dff_A_414Rv4rQ6_0),.clk(gclk));
	jdff dff_A_uY7Sf3477_0(.dout(w_dff_A_b3LfsZFr3_0),.din(w_dff_A_uY7Sf3477_0),.clk(gclk));
	jdff dff_A_b3LfsZFr3_0(.dout(w_dff_A_iTN280Lp2_0),.din(w_dff_A_b3LfsZFr3_0),.clk(gclk));
	jdff dff_A_iTN280Lp2_0(.dout(w_dff_A_f35KXooB9_0),.din(w_dff_A_iTN280Lp2_0),.clk(gclk));
	jdff dff_A_f35KXooB9_0(.dout(G355),.din(w_dff_A_f35KXooB9_0),.clk(gclk));
	jdff dff_A_OClhKNEQ1_2(.dout(w_dff_A_FTUjRZ7L7_0),.din(w_dff_A_OClhKNEQ1_2),.clk(gclk));
	jdff dff_A_FTUjRZ7L7_0(.dout(w_dff_A_2cCv4Uq26_0),.din(w_dff_A_FTUjRZ7L7_0),.clk(gclk));
	jdff dff_A_2cCv4Uq26_0(.dout(w_dff_A_uZeBWyBl2_0),.din(w_dff_A_2cCv4Uq26_0),.clk(gclk));
	jdff dff_A_uZeBWyBl2_0(.dout(w_dff_A_q8aNVWan7_0),.din(w_dff_A_uZeBWyBl2_0),.clk(gclk));
	jdff dff_A_q8aNVWan7_0(.dout(w_dff_A_U5jYb0Me2_0),.din(w_dff_A_q8aNVWan7_0),.clk(gclk));
	jdff dff_A_U5jYb0Me2_0(.dout(w_dff_A_ACAoiT623_0),.din(w_dff_A_U5jYb0Me2_0),.clk(gclk));
	jdff dff_A_ACAoiT623_0(.dout(w_dff_A_1bHwmezi1_0),.din(w_dff_A_ACAoiT623_0),.clk(gclk));
	jdff dff_A_1bHwmezi1_0(.dout(w_dff_A_D2Rjg7pc7_0),.din(w_dff_A_1bHwmezi1_0),.clk(gclk));
	jdff dff_A_D2Rjg7pc7_0(.dout(w_dff_A_L3LjZnyL1_0),.din(w_dff_A_D2Rjg7pc7_0),.clk(gclk));
	jdff dff_A_L3LjZnyL1_0(.dout(w_dff_A_aFU4Geun3_0),.din(w_dff_A_L3LjZnyL1_0),.clk(gclk));
	jdff dff_A_aFU4Geun3_0(.dout(w_dff_A_WziQ7ikS4_0),.din(w_dff_A_aFU4Geun3_0),.clk(gclk));
	jdff dff_A_WziQ7ikS4_0(.dout(w_dff_A_GBsQMOTJ8_0),.din(w_dff_A_WziQ7ikS4_0),.clk(gclk));
	jdff dff_A_GBsQMOTJ8_0(.dout(w_dff_A_lmkQI2SK4_0),.din(w_dff_A_GBsQMOTJ8_0),.clk(gclk));
	jdff dff_A_lmkQI2SK4_0(.dout(w_dff_A_RJnLx0Ps7_0),.din(w_dff_A_lmkQI2SK4_0),.clk(gclk));
	jdff dff_A_RJnLx0Ps7_0(.dout(w_dff_A_x1g1cW3Z6_0),.din(w_dff_A_RJnLx0Ps7_0),.clk(gclk));
	jdff dff_A_x1g1cW3Z6_0(.dout(w_dff_A_Hrh5qpCW6_0),.din(w_dff_A_x1g1cW3Z6_0),.clk(gclk));
	jdff dff_A_Hrh5qpCW6_0(.dout(w_dff_A_OQeLCToq2_0),.din(w_dff_A_Hrh5qpCW6_0),.clk(gclk));
	jdff dff_A_OQeLCToq2_0(.dout(w_dff_A_VuyDDf5T1_0),.din(w_dff_A_OQeLCToq2_0),.clk(gclk));
	jdff dff_A_VuyDDf5T1_0(.dout(w_dff_A_9Mt7Ovpk7_0),.din(w_dff_A_VuyDDf5T1_0),.clk(gclk));
	jdff dff_A_9Mt7Ovpk7_0(.dout(w_dff_A_bk5lb8nL8_0),.din(w_dff_A_9Mt7Ovpk7_0),.clk(gclk));
	jdff dff_A_bk5lb8nL8_0(.dout(G361),.din(w_dff_A_bk5lb8nL8_0),.clk(gclk));
	jdff dff_A_CBmIP1Be0_2(.dout(w_dff_A_Gpm2Gb564_0),.din(w_dff_A_CBmIP1Be0_2),.clk(gclk));
	jdff dff_A_Gpm2Gb564_0(.dout(w_dff_A_W9RtSmlw4_0),.din(w_dff_A_Gpm2Gb564_0),.clk(gclk));
	jdff dff_A_W9RtSmlw4_0(.dout(w_dff_A_V1MY2djm8_0),.din(w_dff_A_W9RtSmlw4_0),.clk(gclk));
	jdff dff_A_V1MY2djm8_0(.dout(w_dff_A_aIeawZzs5_0),.din(w_dff_A_V1MY2djm8_0),.clk(gclk));
	jdff dff_A_aIeawZzs5_0(.dout(w_dff_A_ZT55nFUa8_0),.din(w_dff_A_aIeawZzs5_0),.clk(gclk));
	jdff dff_A_ZT55nFUa8_0(.dout(w_dff_A_4QVdc3U34_0),.din(w_dff_A_ZT55nFUa8_0),.clk(gclk));
	jdff dff_A_4QVdc3U34_0(.dout(w_dff_A_lgQSOq4c1_0),.din(w_dff_A_4QVdc3U34_0),.clk(gclk));
	jdff dff_A_lgQSOq4c1_0(.dout(w_dff_A_J4Br3uUv6_0),.din(w_dff_A_lgQSOq4c1_0),.clk(gclk));
	jdff dff_A_J4Br3uUv6_0(.dout(w_dff_A_yLPWMbr66_0),.din(w_dff_A_J4Br3uUv6_0),.clk(gclk));
	jdff dff_A_yLPWMbr66_0(.dout(w_dff_A_SvvJkNuU9_0),.din(w_dff_A_yLPWMbr66_0),.clk(gclk));
	jdff dff_A_SvvJkNuU9_0(.dout(w_dff_A_pSz1K8PI5_0),.din(w_dff_A_SvvJkNuU9_0),.clk(gclk));
	jdff dff_A_pSz1K8PI5_0(.dout(w_dff_A_VIAjZZZN7_0),.din(w_dff_A_pSz1K8PI5_0),.clk(gclk));
	jdff dff_A_VIAjZZZN7_0(.dout(w_dff_A_btfzpc5T9_0),.din(w_dff_A_VIAjZZZN7_0),.clk(gclk));
	jdff dff_A_btfzpc5T9_0(.dout(w_dff_A_VQItuOtk3_0),.din(w_dff_A_btfzpc5T9_0),.clk(gclk));
	jdff dff_A_VQItuOtk3_0(.dout(w_dff_A_auBXnjy44_0),.din(w_dff_A_VQItuOtk3_0),.clk(gclk));
	jdff dff_A_auBXnjy44_0(.dout(w_dff_A_9TKneLFD7_0),.din(w_dff_A_auBXnjy44_0),.clk(gclk));
	jdff dff_A_9TKneLFD7_0(.dout(w_dff_A_wgvgXfY93_0),.din(w_dff_A_9TKneLFD7_0),.clk(gclk));
	jdff dff_A_wgvgXfY93_0(.dout(w_dff_A_4hQXFrDq2_0),.din(w_dff_A_wgvgXfY93_0),.clk(gclk));
	jdff dff_A_4hQXFrDq2_0(.dout(w_dff_A_pnfM9AFv1_0),.din(w_dff_A_4hQXFrDq2_0),.clk(gclk));
	jdff dff_A_pnfM9AFv1_0(.dout(w_dff_A_Je0TwSxO1_0),.din(w_dff_A_pnfM9AFv1_0),.clk(gclk));
	jdff dff_A_Je0TwSxO1_0(.dout(w_dff_A_yl28ZcZy7_0),.din(w_dff_A_Je0TwSxO1_0),.clk(gclk));
	jdff dff_A_yl28ZcZy7_0(.dout(w_dff_A_kuuk5Rv47_0),.din(w_dff_A_yl28ZcZy7_0),.clk(gclk));
	jdff dff_A_kuuk5Rv47_0(.dout(w_dff_A_hUGUhDUA2_0),.din(w_dff_A_kuuk5Rv47_0),.clk(gclk));
	jdff dff_A_hUGUhDUA2_0(.dout(G358),.din(w_dff_A_hUGUhDUA2_0),.clk(gclk));
	jdff dff_A_xhxNDiQP5_2(.dout(w_dff_A_G8sReFIO7_0),.din(w_dff_A_xhxNDiQP5_2),.clk(gclk));
	jdff dff_A_G8sReFIO7_0(.dout(w_dff_A_GOlZdwVX1_0),.din(w_dff_A_G8sReFIO7_0),.clk(gclk));
	jdff dff_A_GOlZdwVX1_0(.dout(w_dff_A_g7Usebxg6_0),.din(w_dff_A_GOlZdwVX1_0),.clk(gclk));
	jdff dff_A_g7Usebxg6_0(.dout(w_dff_A_OsqYQmCQ7_0),.din(w_dff_A_g7Usebxg6_0),.clk(gclk));
	jdff dff_A_OsqYQmCQ7_0(.dout(w_dff_A_hBCpgmvG9_0),.din(w_dff_A_OsqYQmCQ7_0),.clk(gclk));
	jdff dff_A_hBCpgmvG9_0(.dout(w_dff_A_euATcaSn0_0),.din(w_dff_A_hBCpgmvG9_0),.clk(gclk));
	jdff dff_A_euATcaSn0_0(.dout(w_dff_A_JA7TipuW1_0),.din(w_dff_A_euATcaSn0_0),.clk(gclk));
	jdff dff_A_JA7TipuW1_0(.dout(w_dff_A_krocCZFq9_0),.din(w_dff_A_JA7TipuW1_0),.clk(gclk));
	jdff dff_A_krocCZFq9_0(.dout(w_dff_A_z0qIjVrv3_0),.din(w_dff_A_krocCZFq9_0),.clk(gclk));
	jdff dff_A_z0qIjVrv3_0(.dout(w_dff_A_qBxhkwf92_0),.din(w_dff_A_z0qIjVrv3_0),.clk(gclk));
	jdff dff_A_qBxhkwf92_0(.dout(w_dff_A_JKZTHmqS5_0),.din(w_dff_A_qBxhkwf92_0),.clk(gclk));
	jdff dff_A_JKZTHmqS5_0(.dout(w_dff_A_QOuv3Btq8_0),.din(w_dff_A_JKZTHmqS5_0),.clk(gclk));
	jdff dff_A_QOuv3Btq8_0(.dout(w_dff_A_gEiVgxUV9_0),.din(w_dff_A_QOuv3Btq8_0),.clk(gclk));
	jdff dff_A_gEiVgxUV9_0(.dout(w_dff_A_9Hv7a4ML5_0),.din(w_dff_A_gEiVgxUV9_0),.clk(gclk));
	jdff dff_A_9Hv7a4ML5_0(.dout(w_dff_A_Qv4XXsdJ1_0),.din(w_dff_A_9Hv7a4ML5_0),.clk(gclk));
	jdff dff_A_Qv4XXsdJ1_0(.dout(w_dff_A_3a5I1Iz07_0),.din(w_dff_A_Qv4XXsdJ1_0),.clk(gclk));
	jdff dff_A_3a5I1Iz07_0(.dout(w_dff_A_4OCRONKN0_0),.din(w_dff_A_3a5I1Iz07_0),.clk(gclk));
	jdff dff_A_4OCRONKN0_0(.dout(w_dff_A_eqFUR6LR2_0),.din(w_dff_A_4OCRONKN0_0),.clk(gclk));
	jdff dff_A_eqFUR6LR2_0(.dout(w_dff_A_bZDZd1ym5_0),.din(w_dff_A_eqFUR6LR2_0),.clk(gclk));
	jdff dff_A_bZDZd1ym5_0(.dout(w_dff_A_Zk1YGLwI3_0),.din(w_dff_A_bZDZd1ym5_0),.clk(gclk));
	jdff dff_A_Zk1YGLwI3_0(.dout(w_dff_A_ieGty0Vc3_0),.din(w_dff_A_Zk1YGLwI3_0),.clk(gclk));
	jdff dff_A_ieGty0Vc3_0(.dout(w_dff_A_ldNqHtrp9_0),.din(w_dff_A_ieGty0Vc3_0),.clk(gclk));
	jdff dff_A_ldNqHtrp9_0(.dout(w_dff_A_xa8ZCa0C5_0),.din(w_dff_A_ldNqHtrp9_0),.clk(gclk));
	jdff dff_A_xa8ZCa0C5_0(.dout(G351),.din(w_dff_A_xa8ZCa0C5_0),.clk(gclk));
	jdff dff_A_U1r5udv24_2(.dout(w_dff_A_ansNdKhk9_0),.din(w_dff_A_U1r5udv24_2),.clk(gclk));
	jdff dff_A_ansNdKhk9_0(.dout(w_dff_A_6BMiPlfg1_0),.din(w_dff_A_ansNdKhk9_0),.clk(gclk));
	jdff dff_A_6BMiPlfg1_0(.dout(w_dff_A_jXO6Q5Gk2_0),.din(w_dff_A_6BMiPlfg1_0),.clk(gclk));
	jdff dff_A_jXO6Q5Gk2_0(.dout(w_dff_A_1GjBFRWh5_0),.din(w_dff_A_jXO6Q5Gk2_0),.clk(gclk));
	jdff dff_A_1GjBFRWh5_0(.dout(w_dff_A_4IT75zj88_0),.din(w_dff_A_1GjBFRWh5_0),.clk(gclk));
	jdff dff_A_4IT75zj88_0(.dout(w_dff_A_576dMHkL5_0),.din(w_dff_A_4IT75zj88_0),.clk(gclk));
	jdff dff_A_576dMHkL5_0(.dout(w_dff_A_k1MVbUaM9_0),.din(w_dff_A_576dMHkL5_0),.clk(gclk));
	jdff dff_A_k1MVbUaM9_0(.dout(w_dff_A_jRHX9TTv0_0),.din(w_dff_A_k1MVbUaM9_0),.clk(gclk));
	jdff dff_A_jRHX9TTv0_0(.dout(w_dff_A_qZalfgYi8_0),.din(w_dff_A_jRHX9TTv0_0),.clk(gclk));
	jdff dff_A_qZalfgYi8_0(.dout(w_dff_A_lDMgdEmu1_0),.din(w_dff_A_qZalfgYi8_0),.clk(gclk));
	jdff dff_A_lDMgdEmu1_0(.dout(w_dff_A_CI0WGJSA8_0),.din(w_dff_A_lDMgdEmu1_0),.clk(gclk));
	jdff dff_A_CI0WGJSA8_0(.dout(w_dff_A_5UYdZsCK3_0),.din(w_dff_A_CI0WGJSA8_0),.clk(gclk));
	jdff dff_A_5UYdZsCK3_0(.dout(w_dff_A_U6EaKE1v6_0),.din(w_dff_A_5UYdZsCK3_0),.clk(gclk));
	jdff dff_A_U6EaKE1v6_0(.dout(G372),.din(w_dff_A_U6EaKE1v6_0),.clk(gclk));
	jdff dff_A_Rrj7Q0eY0_2(.dout(w_dff_A_sMvGYYQz5_0),.din(w_dff_A_Rrj7Q0eY0_2),.clk(gclk));
	jdff dff_A_sMvGYYQz5_0(.dout(w_dff_A_9zs5oxww3_0),.din(w_dff_A_sMvGYYQz5_0),.clk(gclk));
	jdff dff_A_9zs5oxww3_0(.dout(w_dff_A_9s9YW4Cz7_0),.din(w_dff_A_9zs5oxww3_0),.clk(gclk));
	jdff dff_A_9s9YW4Cz7_0(.dout(w_dff_A_OELFuOV88_0),.din(w_dff_A_9s9YW4Cz7_0),.clk(gclk));
	jdff dff_A_OELFuOV88_0(.dout(w_dff_A_F1weehSI0_0),.din(w_dff_A_OELFuOV88_0),.clk(gclk));
	jdff dff_A_F1weehSI0_0(.dout(w_dff_A_DE6tKUmO5_0),.din(w_dff_A_F1weehSI0_0),.clk(gclk));
	jdff dff_A_DE6tKUmO5_0(.dout(w_dff_A_zXoUCZGe1_0),.din(w_dff_A_DE6tKUmO5_0),.clk(gclk));
	jdff dff_A_zXoUCZGe1_0(.dout(w_dff_A_vufGJQ6A9_0),.din(w_dff_A_zXoUCZGe1_0),.clk(gclk));
	jdff dff_A_vufGJQ6A9_0(.dout(w_dff_A_rrHNbRHj1_0),.din(w_dff_A_vufGJQ6A9_0),.clk(gclk));
	jdff dff_A_rrHNbRHj1_0(.dout(w_dff_A_RAFXNA2R7_0),.din(w_dff_A_rrHNbRHj1_0),.clk(gclk));
	jdff dff_A_RAFXNA2R7_0(.dout(w_dff_A_Pv2N3cy47_0),.din(w_dff_A_RAFXNA2R7_0),.clk(gclk));
	jdff dff_A_Pv2N3cy47_0(.dout(G369),.din(w_dff_A_Pv2N3cy47_0),.clk(gclk));
	jdff dff_A_ePxRogil5_2(.dout(w_dff_A_896ZXHP37_0),.din(w_dff_A_ePxRogil5_2),.clk(gclk));
	jdff dff_A_896ZXHP37_0(.dout(w_dff_A_29WEVTCJ7_0),.din(w_dff_A_896ZXHP37_0),.clk(gclk));
	jdff dff_A_29WEVTCJ7_0(.dout(w_dff_A_XGLceOqF2_0),.din(w_dff_A_29WEVTCJ7_0),.clk(gclk));
	jdff dff_A_XGLceOqF2_0(.dout(w_dff_A_lIJF73m14_0),.din(w_dff_A_XGLceOqF2_0),.clk(gclk));
	jdff dff_A_lIJF73m14_0(.dout(w_dff_A_31zOZi8z4_0),.din(w_dff_A_lIJF73m14_0),.clk(gclk));
	jdff dff_A_31zOZi8z4_0(.dout(w_dff_A_ASPMRDqh1_0),.din(w_dff_A_31zOZi8z4_0),.clk(gclk));
	jdff dff_A_ASPMRDqh1_0(.dout(w_dff_A_4InhCdb05_0),.din(w_dff_A_ASPMRDqh1_0),.clk(gclk));
	jdff dff_A_4InhCdb05_0(.dout(w_dff_A_QBdaBEbx3_0),.din(w_dff_A_4InhCdb05_0),.clk(gclk));
	jdff dff_A_QBdaBEbx3_0(.dout(w_dff_A_6cz7jF5L6_0),.din(w_dff_A_QBdaBEbx3_0),.clk(gclk));
	jdff dff_A_6cz7jF5L6_0(.dout(w_dff_A_F6Fwcihu2_0),.din(w_dff_A_6cz7jF5L6_0),.clk(gclk));
	jdff dff_A_F6Fwcihu2_0(.dout(G399),.din(w_dff_A_F6Fwcihu2_0),.clk(gclk));
	jdff dff_A_FcBxUslg3_2(.dout(w_dff_A_YfmPqORr1_0),.din(w_dff_A_FcBxUslg3_2),.clk(gclk));
	jdff dff_A_YfmPqORr1_0(.dout(w_dff_A_zMLiY6PE5_0),.din(w_dff_A_YfmPqORr1_0),.clk(gclk));
	jdff dff_A_zMLiY6PE5_0(.dout(w_dff_A_obHbBVlV0_0),.din(w_dff_A_zMLiY6PE5_0),.clk(gclk));
	jdff dff_A_obHbBVlV0_0(.dout(w_dff_A_5oymxLVk5_0),.din(w_dff_A_obHbBVlV0_0),.clk(gclk));
	jdff dff_A_5oymxLVk5_0(.dout(w_dff_A_1wo000Vw3_0),.din(w_dff_A_5oymxLVk5_0),.clk(gclk));
	jdff dff_A_1wo000Vw3_0(.dout(w_dff_A_LCowYuNM1_0),.din(w_dff_A_1wo000Vw3_0),.clk(gclk));
	jdff dff_A_LCowYuNM1_0(.dout(w_dff_A_kRkRToyy2_0),.din(w_dff_A_LCowYuNM1_0),.clk(gclk));
	jdff dff_A_kRkRToyy2_0(.dout(w_dff_A_601qsepq9_0),.din(w_dff_A_kRkRToyy2_0),.clk(gclk));
	jdff dff_A_601qsepq9_0(.dout(w_dff_A_h8q06yD68_0),.din(w_dff_A_601qsepq9_0),.clk(gclk));
	jdff dff_A_h8q06yD68_0(.dout(w_dff_A_plNEmITS6_0),.din(w_dff_A_h8q06yD68_0),.clk(gclk));
	jdff dff_A_plNEmITS6_0(.dout(G364),.din(w_dff_A_plNEmITS6_0),.clk(gclk));
	jdff dff_A_xU860ofM7_2(.dout(w_dff_A_2aK7iVgO7_0),.din(w_dff_A_xU860ofM7_2),.clk(gclk));
	jdff dff_A_2aK7iVgO7_0(.dout(w_dff_A_c6vS7XhE7_0),.din(w_dff_A_2aK7iVgO7_0),.clk(gclk));
	jdff dff_A_c6vS7XhE7_0(.dout(w_dff_A_nEIZ7oaJ9_0),.din(w_dff_A_c6vS7XhE7_0),.clk(gclk));
	jdff dff_A_nEIZ7oaJ9_0(.dout(w_dff_A_RsJWmTEr0_0),.din(w_dff_A_nEIZ7oaJ9_0),.clk(gclk));
	jdff dff_A_RsJWmTEr0_0(.dout(w_dff_A_nxGsCySq0_0),.din(w_dff_A_RsJWmTEr0_0),.clk(gclk));
	jdff dff_A_nxGsCySq0_0(.dout(w_dff_A_L4ElTozG3_0),.din(w_dff_A_nxGsCySq0_0),.clk(gclk));
	jdff dff_A_L4ElTozG3_0(.dout(w_dff_A_tOCJwP9o9_0),.din(w_dff_A_L4ElTozG3_0),.clk(gclk));
	jdff dff_A_tOCJwP9o9_0(.dout(w_dff_A_Nmw7ct6Y4_0),.din(w_dff_A_tOCJwP9o9_0),.clk(gclk));
	jdff dff_A_Nmw7ct6Y4_0(.dout(w_dff_A_RGK8DXxp7_0),.din(w_dff_A_Nmw7ct6Y4_0),.clk(gclk));
	jdff dff_A_RGK8DXxp7_0(.dout(w_dff_A_e0tgGeMz8_0),.din(w_dff_A_RGK8DXxp7_0),.clk(gclk));
	jdff dff_A_e0tgGeMz8_0(.dout(G396),.din(w_dff_A_e0tgGeMz8_0),.clk(gclk));
	jdff dff_A_du0s43qn6_1(.dout(w_dff_A_zNIYIL1a4_0),.din(w_dff_A_du0s43qn6_1),.clk(gclk));
	jdff dff_A_zNIYIL1a4_0(.dout(w_dff_A_mLjXaajH3_0),.din(w_dff_A_zNIYIL1a4_0),.clk(gclk));
	jdff dff_A_mLjXaajH3_0(.dout(w_dff_A_8EMbMuO37_0),.din(w_dff_A_mLjXaajH3_0),.clk(gclk));
	jdff dff_A_8EMbMuO37_0(.dout(w_dff_A_nl32DYBz4_0),.din(w_dff_A_8EMbMuO37_0),.clk(gclk));
	jdff dff_A_nl32DYBz4_0(.dout(w_dff_A_yIiR2RH77_0),.din(w_dff_A_nl32DYBz4_0),.clk(gclk));
	jdff dff_A_yIiR2RH77_0(.dout(w_dff_A_FSORTYGC7_0),.din(w_dff_A_yIiR2RH77_0),.clk(gclk));
	jdff dff_A_FSORTYGC7_0(.dout(w_dff_A_CfeXRRy36_0),.din(w_dff_A_FSORTYGC7_0),.clk(gclk));
	jdff dff_A_CfeXRRy36_0(.dout(G384),.din(w_dff_A_CfeXRRy36_0),.clk(gclk));
	jdff dff_A_WtxJkxnW0_2(.dout(w_dff_A_kvZW2pNS3_0),.din(w_dff_A_WtxJkxnW0_2),.clk(gclk));
	jdff dff_A_kvZW2pNS3_0(.dout(w_dff_A_q8kxXbp53_0),.din(w_dff_A_kvZW2pNS3_0),.clk(gclk));
	jdff dff_A_q8kxXbp53_0(.dout(w_dff_A_dMo2TFOl9_0),.din(w_dff_A_q8kxXbp53_0),.clk(gclk));
	jdff dff_A_dMo2TFOl9_0(.dout(w_dff_A_2PnyNn0i6_0),.din(w_dff_A_dMo2TFOl9_0),.clk(gclk));
	jdff dff_A_2PnyNn0i6_0(.dout(G367),.din(w_dff_A_2PnyNn0i6_0),.clk(gclk));
	jdff dff_A_FnlWl4Ri9_2(.dout(w_dff_A_lCWnU55g8_0),.din(w_dff_A_FnlWl4Ri9_2),.clk(gclk));
	jdff dff_A_lCWnU55g8_0(.dout(w_dff_A_3G595ny84_0),.din(w_dff_A_lCWnU55g8_0),.clk(gclk));
	jdff dff_A_3G595ny84_0(.dout(w_dff_A_1xfDIt8f7_0),.din(w_dff_A_3G595ny84_0),.clk(gclk));
	jdff dff_A_1xfDIt8f7_0(.dout(w_dff_A_KJ62ScuT9_0),.din(w_dff_A_1xfDIt8f7_0),.clk(gclk));
	jdff dff_A_KJ62ScuT9_0(.dout(G387),.din(w_dff_A_KJ62ScuT9_0),.clk(gclk));
	jdff dff_A_HbcdcMhN5_1(.dout(w_dff_A_56KqB1r02_0),.din(w_dff_A_HbcdcMhN5_1),.clk(gclk));
	jdff dff_A_56KqB1r02_0(.dout(w_dff_A_7N4LheIH7_0),.din(w_dff_A_56KqB1r02_0),.clk(gclk));
	jdff dff_A_7N4LheIH7_0(.dout(w_dff_A_qekMxyrJ1_0),.din(w_dff_A_7N4LheIH7_0),.clk(gclk));
	jdff dff_A_qekMxyrJ1_0(.dout(w_dff_A_qsCD0GK29_0),.din(w_dff_A_qekMxyrJ1_0),.clk(gclk));
	jdff dff_A_qsCD0GK29_0(.dout(w_dff_A_ndSfgAv18_0),.din(w_dff_A_qsCD0GK29_0),.clk(gclk));
	jdff dff_A_ndSfgAv18_0(.dout(w_dff_A_9u21ON9p7_0),.din(w_dff_A_ndSfgAv18_0),.clk(gclk));
	jdff dff_A_9u21ON9p7_0(.dout(G393),.din(w_dff_A_9u21ON9p7_0),.clk(gclk));
	jdff dff_A_Xq1tvspa5_1(.dout(w_dff_A_nnOmNew95_0),.din(w_dff_A_Xq1tvspa5_1),.clk(gclk));
	jdff dff_A_nnOmNew95_0(.dout(w_dff_A_KuCBcFFz1_0),.din(w_dff_A_nnOmNew95_0),.clk(gclk));
	jdff dff_A_KuCBcFFz1_0(.dout(w_dff_A_HGJsfUsS7_0),.din(w_dff_A_KuCBcFFz1_0),.clk(gclk));
	jdff dff_A_HGJsfUsS7_0(.dout(w_dff_A_g3M5ctib2_0),.din(w_dff_A_HGJsfUsS7_0),.clk(gclk));
	jdff dff_A_g3M5ctib2_0(.dout(w_dff_A_CXI4NZcl3_0),.din(w_dff_A_g3M5ctib2_0),.clk(gclk));
	jdff dff_A_CXI4NZcl3_0(.dout(G390),.din(w_dff_A_CXI4NZcl3_0),.clk(gclk));
	jdff dff_A_XeMRgOBq9_1(.dout(w_dff_A_tRgQlSEG7_0),.din(w_dff_A_XeMRgOBq9_1),.clk(gclk));
	jdff dff_A_tRgQlSEG7_0(.dout(w_dff_A_TugvvbVr3_0),.din(w_dff_A_tRgQlSEG7_0),.clk(gclk));
	jdff dff_A_TugvvbVr3_0(.dout(w_dff_A_e7jcRQLs2_0),.din(w_dff_A_TugvvbVr3_0),.clk(gclk));
	jdff dff_A_e7jcRQLs2_0(.dout(w_dff_A_3x8hGX1b5_0),.din(w_dff_A_e7jcRQLs2_0),.clk(gclk));
	jdff dff_A_3x8hGX1b5_0(.dout(G378),.din(w_dff_A_3x8hGX1b5_0),.clk(gclk));
	jdff dff_A_suoffQtL3_1(.dout(w_dff_A_WkLmf1A43_0),.din(w_dff_A_suoffQtL3_1),.clk(gclk));
	jdff dff_A_WkLmf1A43_0(.dout(w_dff_A_TBa6wdVG1_0),.din(w_dff_A_WkLmf1A43_0),.clk(gclk));
	jdff dff_A_TBa6wdVG1_0(.dout(G375),.din(w_dff_A_TBa6wdVG1_0),.clk(gclk));
	jdff dff_A_BWmK6cNT5_1(.dout(w_dff_A_Svc0U3fn9_0),.din(w_dff_A_BWmK6cNT5_1),.clk(gclk));
	jdff dff_A_Svc0U3fn9_0(.dout(w_dff_A_Wir5E6q46_0),.din(w_dff_A_Svc0U3fn9_0),.clk(gclk));
	jdff dff_A_Wir5E6q46_0(.dout(w_dff_A_QW8FzAo49_0),.din(w_dff_A_Wir5E6q46_0),.clk(gclk));
	jdff dff_A_QW8FzAo49_0(.dout(w_dff_A_Tn1IrHG90_0),.din(w_dff_A_QW8FzAo49_0),.clk(gclk));
	jdff dff_A_Tn1IrHG90_0(.dout(G381),.din(w_dff_A_Tn1IrHG90_0),.clk(gclk));
	jdff dff_A_cajdjt8l9_1(.dout(G407),.din(w_dff_A_cajdjt8l9_1),.clk(gclk));
	jdff dff_A_AmqgxAwU4_2(.dout(G402),.din(w_dff_A_AmqgxAwU4_2),.clk(gclk));
endmodule

