/*

c1355:
	jxor: 124
	jspl: 39
	jspl3: 79
	jnot: 9
	jdff: 400
	jand: 72
	jor: 10

Summary:
	jxor: 124
	jspl: 39
	jspl3: 79
	jnot: 9
	jdff: 400
	jand: 72
	jor: 10
*/

module c1355(gclk, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat, G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat, G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat, G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat, G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat, G1352gat, G1353gat, G1354gat, G1355gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G15gat;
	input G22gat;
	input G29gat;
	input G36gat;
	input G43gat;
	input G50gat;
	input G57gat;
	input G64gat;
	input G71gat;
	input G78gat;
	input G85gat;
	input G92gat;
	input G99gat;
	input G106gat;
	input G113gat;
	input G120gat;
	input G127gat;
	input G134gat;
	input G141gat;
	input G148gat;
	input G155gat;
	input G162gat;
	input G169gat;
	input G176gat;
	input G183gat;
	input G190gat;
	input G197gat;
	input G204gat;
	input G211gat;
	input G218gat;
	input G225gat;
	input G226gat;
	input G227gat;
	input G228gat;
	input G229gat;
	input G230gat;
	input G231gat;
	input G232gat;
	input G233gat;
	output G1324gat;
	output G1325gat;
	output G1326gat;
	output G1327gat;
	output G1328gat;
	output G1329gat;
	output G1330gat;
	output G1331gat;
	output G1332gat;
	output G1333gat;
	output G1334gat;
	output G1335gat;
	output G1336gat;
	output G1337gat;
	output G1338gat;
	output G1339gat;
	output G1340gat;
	output G1341gat;
	output G1342gat;
	output G1343gat;
	output G1344gat;
	output G1345gat;
	output G1346gat;
	output G1347gat;
	output G1348gat;
	output G1349gat;
	output G1350gat;
	output G1351gat;
	output G1352gat;
	output G1353gat;
	output G1354gat;
	output G1355gat;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n203;
	wire n205;
	wire n207;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n221;
	wire n223;
	wire n225;
	wire n227;
	wire n228;
	wire n229;
	wire n231;
	wire n233;
	wire n235;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n250;
	wire n252;
	wire n254;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n261;
	wire n263;
	wire n265;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n272;
	wire n274;
	wire n276;
	wire n278;
	wire n279;
	wire n280;
	wire n282;
	wire n284;
	wire n286;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G8gat_0;
	wire [2:0] w_G15gat_0;
	wire [2:0] w_G22gat_0;
	wire [2:0] w_G29gat_0;
	wire [2:0] w_G36gat_0;
	wire [2:0] w_G43gat_0;
	wire [2:0] w_G50gat_0;
	wire [2:0] w_G57gat_0;
	wire [2:0] w_G64gat_0;
	wire [2:0] w_G71gat_0;
	wire [2:0] w_G78gat_0;
	wire [2:0] w_G85gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G99gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G113gat_0;
	wire [2:0] w_G120gat_0;
	wire [2:0] w_G127gat_0;
	wire [2:0] w_G134gat_0;
	wire [2:0] w_G141gat_0;
	wire [2:0] w_G148gat_0;
	wire [2:0] w_G155gat_0;
	wire [2:0] w_G162gat_0;
	wire [2:0] w_G169gat_0;
	wire [2:0] w_G176gat_0;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G190gat_0;
	wire [2:0] w_G197gat_0;
	wire [2:0] w_G204gat_0;
	wire [2:0] w_G211gat_0;
	wire [2:0] w_G218gat_0;
	wire [1:0] w_G225gat_0;
	wire [1:0] w_G226gat_0;
	wire [1:0] w_G227gat_0;
	wire [1:0] w_G228gat_0;
	wire [1:0] w_G229gat_0;
	wire [1:0] w_G230gat_0;
	wire [1:0] w_G231gat_0;
	wire [1:0] w_G232gat_0;
	wire [2:0] w_G233gat_0;
	wire [2:0] w_G233gat_1;
	wire [2:0] w_G233gat_2;
	wire [2:0] w_G233gat_3;
	wire [2:0] w_n76_0;
	wire [1:0] w_n76_1;
	wire [2:0] w_n83_0;
	wire [1:0] w_n84_0;
	wire [2:0] w_n85_0;
	wire [2:0] w_n85_1;
	wire [2:0] w_n87_0;
	wire [2:0] w_n87_1;
	wire [2:0] w_n87_2;
	wire [1:0] w_n87_3;
	wire [2:0] w_n90_0;
	wire [2:0] w_n95_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n103_0;
	wire [2:0] w_n104_0;
	wire [1:0] w_n112_0;
	wire [2:0] w_n113_0;
	wire [1:0] w_n120_0;
	wire [2:0] w_n121_0;
	wire [2:0] w_n127_0;
	wire [1:0] w_n127_1;
	wire [2:0] w_n131_0;
	wire [1:0] w_n131_1;
	wire [2:0] w_n135_0;
	wire [1:0] w_n139_0;
	wire [2:0] w_n140_0;
	wire [2:0] w_n140_1;
	wire [2:0] w_n145_0;
	wire [1:0] w_n149_0;
	wire [1:0] w_n153_0;
	wire [2:0] w_n154_0;
	wire [1:0] w_n155_0;
	wire [1:0] w_n162_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n169_0;
	wire [2:0] w_n170_0;
	wire [2:0] w_n170_1;
	wire [1:0] w_n171_0;
	wire [2:0] w_n173_0;
	wire [1:0] w_n173_1;
	wire [2:0] w_n178_0;
	wire [2:0] w_n178_1;
	wire [2:0] w_n183_0;
	wire [2:0] w_n183_1;
	wire [2:0] w_n188_0;
	wire [2:0] w_n188_1;
	wire [2:0] w_n193_0;
	wire [2:0] w_n193_1;
	wire [2:0] w_n197_0;
	wire [1:0] w_n198_0;
	wire [2:0] w_n200_0;
	wire [1:0] w_n200_1;
	wire [2:0] w_n212_0;
	wire [2:0] w_n215_0;
	wire [2:0] w_n215_1;
	wire [1:0] w_n216_0;
	wire [2:0] w_n218_0;
	wire [1:0] w_n218_1;
	wire [2:0] w_n228_0;
	wire [1:0] w_n228_1;
	wire [2:0] w_n243_0;
	wire [1:0] w_n243_1;
	wire [1:0] w_n244_0;
	wire [1:0] w_n245_0;
	wire [2:0] w_n247_0;
	wire [1:0] w_n247_1;
	wire [1:0] w_n256_0;
	wire [2:0] w_n258_0;
	wire [1:0] w_n258_1;
	wire [1:0] w_n267_0;
	wire [2:0] w_n269_0;
	wire [1:0] w_n269_1;
	wire [2:0] w_n279_0;
	wire [1:0] w_n279_1;
	wire w_dff_B_JpMKVmZl9_0;
	wire w_dff_B_06NNXGq62_0;
	wire w_dff_B_btmg2ddw6_0;
	wire w_dff_B_pn2oIhGQ2_0;
	wire w_dff_B_2Km8CvHk0_0;
	wire w_dff_A_UEFCxbK25_0;
	wire w_dff_A_g1BfgCzT0_0;
	wire w_dff_A_v7xPrecR9_0;
	wire w_dff_A_af33HeQj4_0;
	wire w_dff_A_ZlG0OEia8_1;
	wire w_dff_A_cUtTnJo07_1;
	wire w_dff_A_PJl0B6a46_1;
	wire w_dff_A_HjKQHrjl4_1;
	wire w_dff_A_nlWAvpXB4_0;
	wire w_dff_A_xT1L5ZQw9_0;
	wire w_dff_A_rPUdUG9W3_0;
	wire w_dff_A_SReMXxCA6_0;
	wire w_dff_A_GYNK3MhN6_1;
	wire w_dff_A_1MgGcnkf2_1;
	wire w_dff_A_J2Qlhlvh1_1;
	wire w_dff_A_tX3pqyub1_1;
	wire w_dff_A_VUZMEUK57_0;
	wire w_dff_A_C2tTUdFW9_0;
	wire w_dff_A_hlETrfwt2_0;
	wire w_dff_A_RjilLUSm9_0;
	wire w_dff_A_zmb6Iz487_1;
	wire w_dff_A_RpJ5IAsl3_1;
	wire w_dff_A_vZXhAKHK9_1;
	wire w_dff_A_TP2le7tE4_1;
	wire w_dff_B_2INi8XQd3_0;
	wire w_dff_A_ITY20qju2_0;
	wire w_dff_A_XPZNI1cD3_0;
	wire w_dff_A_alsCGyvt9_0;
	wire w_dff_A_InqPmjAf2_0;
	wire w_dff_A_hjOrORjM4_2;
	wire w_dff_A_Zzioavus5_2;
	wire w_dff_A_05lu8w600_2;
	wire w_dff_A_jWD4RRAF2_2;
	wire w_dff_B_pdYoucrR6_1;
	wire w_dff_A_9yOWnLIP5_0;
	wire w_dff_A_4iPUKJBz0_0;
	wire w_dff_A_3BJoGveC8_0;
	wire w_dff_A_hmGuCVsx1_0;
	wire w_dff_A_jkZrImb09_1;
	wire w_dff_A_xpcBif0g1_1;
	wire w_dff_A_8qybLMO87_1;
	wire w_dff_A_Gmtn59Zy1_1;
	wire w_dff_B_1gFbPR9p4_0;
	wire w_dff_A_vDuh33W94_0;
	wire w_dff_A_CuHLstmq1_0;
	wire w_dff_A_iMxb8M8i4_0;
	wire w_dff_A_vjFuTVfN7_0;
	wire w_dff_A_Q3bxO8ma6_2;
	wire w_dff_A_gTpzAnOG5_2;
	wire w_dff_A_bpEI5ce25_2;
	wire w_dff_A_rEuNCYgm9_2;
	wire w_dff_B_qOd2XWaL1_0;
	wire w_dff_A_Kxc47GtV0_1;
	wire w_dff_A_iBZDce420_1;
	wire w_dff_A_jH4meBDb6_1;
	wire w_dff_A_gz6QLfLj0_1;
	wire w_dff_A_EovRSw7Z5_2;
	wire w_dff_A_l73MpFsM3_2;
	wire w_dff_A_5mg9CYSE6_2;
	wire w_dff_A_9jk7SHR34_2;
	wire w_dff_B_6HSWmL7A4_1;
	wire w_dff_A_6wht6jjS9_1;
	wire w_dff_A_CuUeb5F64_1;
	wire w_dff_A_4sK58bz96_1;
	wire w_dff_A_gtr1tQUw2_1;
	wire w_dff_A_QiFr9GKJ0_2;
	wire w_dff_A_L0zuODby1_2;
	wire w_dff_A_FOmorWB30_2;
	wire w_dff_A_mPztUbUJ7_2;
	wire w_dff_B_SoJaXzm66_1;
	wire w_dff_A_rszApFuE6_1;
	wire w_dff_A_CJhm6qde5_1;
	wire w_dff_A_QZ4juBak6_1;
	wire w_dff_A_wRehXAhG7_1;
	wire w_dff_A_bUlwPINx4_2;
	wire w_dff_A_QseusKqf2_2;
	wire w_dff_A_GzkFXzdh3_2;
	wire w_dff_A_zPPLunni8_2;
	wire w_dff_B_gH4FIO5Q8_0;
	wire w_dff_B_5ISMQj3O1_0;
	wire w_dff_A_Jh1Vr3280_0;
	wire w_dff_A_aAIfW8Qg4_0;
	wire w_dff_A_QlTneZLs8_0;
	wire w_dff_A_zFHeq7ah5_0;
	wire w_dff_A_J7XXJgdO6_2;
	wire w_dff_A_BC676bst6_2;
	wire w_dff_A_oGmJaPL98_2;
	wire w_dff_A_oSDLP5Yh7_2;
	wire w_dff_B_mkSFGFSU5_0;
	wire w_dff_A_rTPmh6yz8_0;
	wire w_dff_A_OUnsK4da7_0;
	wire w_dff_A_NuFlGr284_0;
	wire w_dff_A_agrTuzZR9_0;
	wire w_dff_A_NYSv60IV8_2;
	wire w_dff_A_9U3ZkJ0I8_2;
	wire w_dff_A_1WSdQZiH5_2;
	wire w_dff_A_3jjv8xX07_2;
	wire w_dff_B_6PMEPoOn5_1;
	wire w_dff_A_KbrTgli03_0;
	wire w_dff_A_Eet2dHw20_0;
	wire w_dff_A_x1mHxHrO7_0;
	wire w_dff_A_2ukqXYEG5_0;
	wire w_dff_A_EIvQluIV0_0;
	wire w_dff_A_QI1EBWci3_0;
	wire w_dff_A_BILdSeYm1_0;
	wire w_dff_A_H4KCkzPz9_0;
	wire w_dff_A_D6dAaGkh4_0;
	wire w_dff_A_v25iy4EA9_0;
	wire w_dff_A_6ws0EdZG4_0;
	wire w_dff_A_9npPaJRl3_0;
	wire w_dff_A_rKPIajl82_0;
	wire w_dff_A_fRmLfm376_0;
	wire w_dff_A_3apjY6hn4_0;
	wire w_dff_A_ANKXSSDB1_0;
	wire w_dff_A_3BNT17BE6_0;
	wire w_dff_A_OyAPfEGQ2_0;
	wire w_dff_A_rphy6nna1_0;
	wire w_dff_A_vhP9Nzv64_0;
	wire w_dff_A_XQXlRbjK0_0;
	wire w_dff_A_cM2lksrO9_0;
	wire w_dff_A_uQmCCl9M8_0;
	wire w_dff_A_lVWX8ZPp5_0;
	wire w_dff_A_fizDFYwF0_0;
	wire w_dff_A_rkxtQIjF0_0;
	wire w_dff_A_PxtJZ94Q4_0;
	wire w_dff_A_Q7Uv4kNI6_0;
	wire w_dff_A_PU5o12Yv5_0;
	wire w_dff_A_gK9Yriil2_0;
	wire w_dff_A_FRlZvOYt1_0;
	wire w_dff_A_ZotPLopL7_0;
	wire w_dff_A_yTmacIWl0_0;
	wire w_dff_A_JRw8BJae0_0;
	wire w_dff_A_O0GHoQSB5_0;
	wire w_dff_A_rk60w1u35_0;
	wire w_dff_A_GafMvStw1_0;
	wire w_dff_A_Ot2yuFw25_0;
	wire w_dff_A_4p02WoLu4_0;
	wire w_dff_A_izpkRR5Q9_0;
	wire w_dff_A_GFJ60qxS4_0;
	wire w_dff_A_LH3URp8V9_0;
	wire w_dff_A_9Q0hwyxl1_0;
	wire w_dff_A_eMLKePgr5_0;
	wire w_dff_A_MIJ29XG96_0;
	wire w_dff_A_JmQdnqEg1_0;
	wire w_dff_A_dV1zL4912_0;
	wire w_dff_A_CQGlUN0V0_0;
	wire w_dff_A_yHdzh8Fy5_0;
	wire w_dff_A_JsB1D3RH3_0;
	wire w_dff_A_NrcsKszJ3_0;
	wire w_dff_A_gF0cEuQl2_0;
	wire w_dff_A_CxkqJPHN1_0;
	wire w_dff_A_j9H4W8fS4_0;
	wire w_dff_A_vfGtvVCT7_0;
	wire w_dff_A_5iniG0Kh2_0;
	wire w_dff_A_tW67o2ko8_0;
	wire w_dff_A_YI8ihUHD9_0;
	wire w_dff_A_2f3bqegi4_0;
	wire w_dff_A_eBanHSkz1_0;
	wire w_dff_A_jc5aLY4O8_0;
	wire w_dff_A_2rokQqMN5_0;
	wire w_dff_A_Gw2FmiMh0_0;
	wire w_dff_A_3D0cCzIt9_0;
	wire w_dff_A_BhFxGBCj9_0;
	wire w_dff_A_HMn7Fy4c6_0;
	wire w_dff_A_slSttrwN2_0;
	wire w_dff_A_R1Hjm5YU9_0;
	wire w_dff_A_wUu2E1Tg6_0;
	wire w_dff_A_RbKkd4CZ7_0;
	wire w_dff_A_JGf72LPl7_0;
	wire w_dff_A_IWKs33zr3_0;
	wire w_dff_A_bHvBKiqW2_0;
	wire w_dff_A_vOk5WkIj4_0;
	wire w_dff_A_BQ855u9F3_0;
	wire w_dff_A_Nq4r9eQU4_0;
	wire w_dff_A_F8juxuHs6_0;
	wire w_dff_A_7CJVnmPL8_0;
	wire w_dff_A_LgLOrG210_0;
	wire w_dff_A_jQITJNMj2_0;
	wire w_dff_A_O0xEvHZB4_0;
	wire w_dff_A_YWECeiuH1_0;
	wire w_dff_A_K8ht5ClC1_0;
	wire w_dff_A_APuOohiE9_0;
	wire w_dff_A_qsbhR7XD2_0;
	wire w_dff_A_hJCevG5D6_0;
	wire w_dff_A_wfJVwl017_0;
	wire w_dff_A_CAd6zvoO0_0;
	wire w_dff_A_P3d78dXh2_0;
	wire w_dff_A_vUEa1tOP9_0;
	wire w_dff_A_JRmpj3vW1_0;
	wire w_dff_A_mIkq9KWc7_0;
	wire w_dff_A_kVgO0sV91_0;
	wire w_dff_A_ivwwygLT0_0;
	wire w_dff_A_tnoy1bpI3_0;
	wire w_dff_A_xl3vBmQY7_0;
	wire w_dff_A_lw9uu5et0_0;
	wire w_dff_A_ApUu8QX68_0;
	wire w_dff_A_SyaQvzUr9_0;
	wire w_dff_A_wqM4bRK39_0;
	wire w_dff_A_hmxSCtab0_0;
	wire w_dff_A_IiVfJ6Lt3_0;
	wire w_dff_A_dEnjAOzf4_0;
	wire w_dff_A_SMsC3kwI7_0;
	wire w_dff_A_JpiXpZXw7_0;
	wire w_dff_A_Q9tQXbC02_0;
	wire w_dff_A_MrFTOFe00_0;
	wire w_dff_A_bH14foRf7_0;
	wire w_dff_A_SS3Vkgin2_0;
	wire w_dff_A_lLV4X3S78_0;
	wire w_dff_A_ErAp9cSi4_0;
	wire w_dff_A_KDP32BWO9_0;
	wire w_dff_A_V7QMWGL00_0;
	wire w_dff_A_uNJqB8J02_0;
	wire w_dff_A_b8JYYJic6_0;
	wire w_dff_A_rmSHLCRY7_0;
	wire w_dff_A_i5rz0XZO0_0;
	wire w_dff_A_5xvVeZUQ1_0;
	wire w_dff_A_L926TgT70_0;
	wire w_dff_A_uGDL3LlH8_0;
	wire w_dff_A_LQnVihV25_0;
	wire w_dff_A_LARyHFiL2_0;
	wire w_dff_A_y93UQyjQ9_0;
	wire w_dff_A_mgdO3aCs5_0;
	wire w_dff_A_Cds15KqZ2_0;
	wire w_dff_A_RJtrtdK02_0;
	wire w_dff_A_8cZgt6PL3_0;
	wire w_dff_A_gyWsRh5u5_0;
	wire w_dff_A_cP7XeylB5_0;
	wire w_dff_A_WKBsu2kb7_0;
	wire w_dff_A_yk7MLahK2_0;
	wire w_dff_A_6IjGjCaJ9_0;
	wire w_dff_A_aBYOTLyX7_0;
	wire w_dff_A_xQl0VRP72_0;
	wire w_dff_A_DgsZDsXk0_0;
	wire w_dff_A_8tqHFnHw5_0;
	wire w_dff_A_gA4zrwt49_0;
	wire w_dff_A_0geqOlnf9_0;
	wire w_dff_A_OTtH03OS3_0;
	wire w_dff_A_7rsDzaEd8_0;
	wire w_dff_A_8msweTtN0_0;
	wire w_dff_A_P6twqtTa7_0;
	wire w_dff_A_HZ4p6TmS2_0;
	wire w_dff_A_fdC9aunC4_0;
	wire w_dff_A_qxa5TtMk0_0;
	wire w_dff_A_V76aXWiQ6_0;
	wire w_dff_A_WRnJI9Kl9_0;
	wire w_dff_A_kDVMhmEy5_0;
	wire w_dff_A_BvkTwHL13_0;
	wire w_dff_A_7I6nZD8M5_0;
	wire w_dff_A_jzEg5pm64_0;
	wire w_dff_A_nCG7rUg54_0;
	wire w_dff_A_gBnaavUD6_0;
	wire w_dff_A_d6pMsqyY1_0;
	wire w_dff_A_8XMPAys19_0;
	wire w_dff_A_YZJZwMlC4_0;
	wire w_dff_A_cMuuJ3HN3_0;
	wire w_dff_A_YsrSFMqX9_0;
	wire w_dff_A_aqUX2jBo3_0;
	wire w_dff_A_hQ7lpytX3_0;
	wire w_dff_A_3lu6ZQS50_0;
	wire w_dff_A_R1Kk3biT2_0;
	wire w_dff_A_z94p2JxK8_0;
	wire w_dff_A_6WvV3fa74_0;
	wire w_dff_A_eYngrMjt2_0;
	wire w_dff_A_7P5UDB3E3_0;
	wire w_dff_A_8uX3ycbG4_0;
	wire w_dff_A_EGVbRc0F9_0;
	wire w_dff_A_iDYW34Zv8_0;
	wire w_dff_A_FqZZi1YR1_0;
	wire w_dff_A_stWt3Lte9_0;
	wire w_dff_A_IqyTzLwR5_0;
	wire w_dff_A_845PcrZY6_0;
	wire w_dff_A_eWXkWq271_0;
	wire w_dff_A_KYjcePUD0_0;
	wire w_dff_A_izVBTHt02_0;
	wire w_dff_A_cKHFlPhF7_0;
	wire w_dff_A_Ppkqod837_0;
	wire w_dff_A_BrXcoD0H4_0;
	wire w_dff_A_1aKUPuaX8_0;
	wire w_dff_A_GWzDKBZD4_1;
	wire w_dff_A_btjalPWr6_1;
	wire w_dff_A_b8y4dfmI3_1;
	wire w_dff_A_mXsTGYGu8_1;
	wire w_dff_A_lNEaeZEi6_2;
	wire w_dff_A_xzS7HUuI9_2;
	wire w_dff_A_3yfnbr4L1_2;
	wire w_dff_A_zHWUR9p43_2;
	wire w_dff_A_ibsX1cxs4_0;
	wire w_dff_A_tCdREcKa2_0;
	wire w_dff_A_vFNQZEMZ1_0;
	wire w_dff_A_iUmeuBPm1_0;
	wire w_dff_A_PzxzdSoV4_0;
	wire w_dff_A_rjqeuLkK5_0;
	wire w_dff_A_jUz51r6j8_0;
	wire w_dff_A_Box9InxF9_0;
	wire w_dff_A_rAX5N1mb8_0;
	wire w_dff_A_3BfG94Lu2_0;
	wire w_dff_A_eHZZYIL78_0;
	wire w_dff_A_uBxlZuto1_0;
	wire w_dff_A_jAx6sNoT5_0;
	wire w_dff_A_rMxDDKKr1_0;
	wire w_dff_A_vUssrorw4_0;
	wire w_dff_A_sgcqp6yk5_0;
	wire w_dff_A_bh1PU6yV7_0;
	wire w_dff_A_R0VlCnVr4_0;
	wire w_dff_A_nh98z9qp3_0;
	wire w_dff_A_38qDdbeF7_0;
	wire w_dff_A_AVpyYFh75_0;
	wire w_dff_A_ODtt1Elw8_0;
	wire w_dff_A_ybj2aDPc2_0;
	wire w_dff_A_jKvWkiT39_0;
	wire w_dff_A_ui2ARFNK3_0;
	wire w_dff_A_pXC3GHm42_0;
	wire w_dff_A_4ix7yO1c6_0;
	wire w_dff_A_u4DOqvYj9_0;
	wire w_dff_A_mnUv4xHz2_0;
	wire w_dff_A_Zq7j6Wug3_0;
	wire w_dff_A_7kQCIwvX5_0;
	wire w_dff_A_cZZvKzC88_0;
	wire w_dff_A_xMa23chv2_0;
	wire w_dff_A_aLRmqX4y5_0;
	wire w_dff_A_0rgyHWSn3_0;
	wire w_dff_A_7bIcqB0f7_0;
	wire w_dff_A_HgIZFkTJ4_0;
	wire w_dff_A_S1zPxHxo4_0;
	wire w_dff_A_N5qQfwvz4_0;
	wire w_dff_A_SbXpIhpg1_0;
	wire w_dff_A_jARsJAHT1_0;
	wire w_dff_A_8bmxk5ct5_0;
	wire w_dff_A_YLBSHGtv6_0;
	wire w_dff_A_Wo2KMpZw1_0;
	wire w_dff_A_jq8KQ46T1_0;
	wire w_dff_A_dcTQargd2_0;
	wire w_dff_A_41sYUzFO3_0;
	wire w_dff_A_sJYDNqPR5_0;
	wire w_dff_A_pegcWvZv1_0;
	wire w_dff_A_iweDOZN63_0;
	wire w_dff_A_laIWXTMB6_0;
	wire w_dff_A_uiXBeY8o9_0;
	wire w_dff_A_oczNyP5o9_0;
	wire w_dff_A_VwcYzyRB8_0;
	wire w_dff_A_OzhPNIhy0_0;
	wire w_dff_A_2HuVFVWt7_0;
	wire w_dff_A_KoDAHiOe0_0;
	wire w_dff_A_JCRifkk40_0;
	wire w_dff_A_Uhqsz52h4_0;
	wire w_dff_A_cldGPkuk8_0;
	wire w_dff_A_N76rax1t8_0;
	wire w_dff_A_ik88G5GF9_0;
	wire w_dff_A_LGoqKOvX1_0;
	wire w_dff_A_hjYQRhIH2_0;
	wire w_dff_A_tNw4S6Df5_0;
	wire w_dff_A_FFLW49A00_0;
	wire w_dff_A_jsZlvTon1_0;
	wire w_dff_A_j6uKOymn5_0;
	wire w_dff_A_rAMLe7Y78_0;
	wire w_dff_A_eFPGJfq35_0;
	wire w_dff_A_1rgRVts25_0;
	wire w_dff_A_jpqv8m5G6_0;
	wire w_dff_B_lGXLKP903_0;
	wire w_dff_A_cHovN6V07_0;
	wire w_dff_A_bLhCn3Y76_0;
	wire w_dff_A_mBEEZ1aI1_0;
	wire w_dff_A_3jdHesJ14_0;
	wire w_dff_A_6PHoglSS2_0;
	wire w_dff_A_7DELWPFL7_0;
	wire w_dff_A_lP662Jqj8_0;
	wire w_dff_A_ZMWiXPVM8_0;
	wire w_dff_A_v7ED5tYc9_0;
	wire w_dff_A_VwB4v1RI5_0;
	wire w_dff_A_LaQyHxma8_0;
	wire w_dff_A_I3KZClPs6_0;
	wire w_dff_A_ht4nWXRa4_0;
	wire w_dff_A_FOQxKWTa0_0;
	wire w_dff_A_CbVdveOh1_0;
	wire w_dff_A_Kz7moYql1_0;
	wire w_dff_A_50J4jW6q2_0;
	wire w_dff_A_SDqRMGgO8_0;
	wire w_dff_A_x3xM2y5l7_0;
	wire w_dff_A_RGLLuGf07_0;
	wire w_dff_A_baFEwu9S7_0;
	wire w_dff_A_A8XbdSah2_0;
	wire w_dff_A_n2qcSHdG9_0;
	wire w_dff_A_apya2kGJ1_0;
	wire w_dff_A_qnaUJiEI2_0;
	wire w_dff_A_eD3q2sz12_0;
	wire w_dff_A_jrgtPD7H9_0;
	wire w_dff_A_3pmWagUy8_0;
	wire w_dff_A_v7PwXPi94_0;
	wire w_dff_A_cPhaBPVu6_0;
	wire w_dff_A_hxFmtyc21_0;
	wire w_dff_A_nc7ErHap5_0;
	wire w_dff_A_oKgMuC9Y5_0;
	wire w_dff_A_UBXeWElZ8_0;
	wire w_dff_A_7UIp3iqL5_0;
	wire w_dff_A_EHOuqmax2_0;
	jand g000(.dina(w_G233gat_3[2]),.dinb(w_G225gat_0[1]),.dout(n73),.clk(gclk));
	jxor g001(.dina(w_G134gat_0[2]),.dinb(w_G127gat_0[2]),.dout(n74),.clk(gclk));
	jxor g002(.dina(w_G120gat_0[2]),.dinb(w_G113gat_0[2]),.dout(n75),.clk(gclk));
	jxor g003(.dina(n75),.dinb(n74),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_n76_1[1]),.dinb(w_dff_B_pdYoucrR6_1),.dout(n77),.clk(gclk));
	jxor g005(.dina(w_G85gat_0[2]),.dinb(w_G57gat_0[2]),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_G29gat_0[2]),.dinb(w_G1gat_0[2]),.dout(n79),.clk(gclk));
	jxor g007(.dina(n79),.dinb(n78),.dout(n80),.clk(gclk));
	jxor g008(.dina(w_G162gat_0[2]),.dinb(w_G155gat_0[2]),.dout(n81),.clk(gclk));
	jxor g009(.dina(w_G148gat_0[2]),.dinb(w_G141gat_0[2]),.dout(n82),.clk(gclk));
	jxor g010(.dina(n82),.dinb(n81),.dout(n83),.clk(gclk));
	jxor g011(.dina(w_n83_0[2]),.dinb(n80),.dout(n84),.clk(gclk));
	jxor g012(.dina(w_n84_0[1]),.dinb(n77),.dout(n85),.clk(gclk));
	jnot g013(.din(w_G225gat_0[0]),.dout(n86),.clk(gclk));
	jnot g014(.din(w_G233gat_3[1]),.dout(n87),.clk(gclk));
	jor g015(.dina(w_n87_3[1]),.dinb(n86),.dout(n88),.clk(gclk));
	jxor g016(.dina(w_n76_1[0]),.dinb(n88),.dout(n89),.clk(gclk));
	jxor g017(.dina(w_n84_0[0]),.dinb(n89),.dout(n90),.clk(gclk));
	jnot g018(.din(w_G226gat_0[1]),.dout(n91),.clk(gclk));
	jor g019(.dina(w_n87_3[0]),.dinb(n91),.dout(n92),.clk(gclk));
	jxor g020(.dina(w_G218gat_0[2]),.dinb(w_G211gat_0[2]),.dout(n93),.clk(gclk));
	jxor g021(.dina(w_G204gat_0[2]),.dinb(w_G197gat_0[2]),.dout(n94),.clk(gclk));
	jxor g022(.dina(n94),.dinb(n93),.dout(n95),.clk(gclk));
	jxor g023(.dina(w_n95_0[2]),.dinb(n92),.dout(n96),.clk(gclk));
	jxor g024(.dina(w_G190gat_0[2]),.dinb(w_G183gat_0[2]),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_G176gat_0[2]),.dinb(w_G169gat_0[2]),.dout(n98),.clk(gclk));
	jxor g026(.dina(n98),.dinb(n97),.dout(n99),.clk(gclk));
	jxor g027(.dina(w_G92gat_0[2]),.dinb(w_G64gat_0[2]),.dout(n100),.clk(gclk));
	jxor g028(.dina(w_G36gat_0[2]),.dinb(w_G8gat_0[2]),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n100),.dout(n102),.clk(gclk));
	jxor g030(.dina(n102),.dinb(w_n99_0[1]),.dout(n103),.clk(gclk));
	jxor g031(.dina(w_n103_0[1]),.dinb(n96),.dout(n104),.clk(gclk));
	jxor g032(.dina(w_n104_0[2]),.dinb(w_n90_0[2]),.dout(n105),.clk(gclk));
	jnot g033(.din(w_G227gat_0[1]),.dout(n106),.clk(gclk));
	jor g034(.dina(w_n87_2[2]),.dinb(n106),.dout(n107),.clk(gclk));
	jxor g035(.dina(n107),.dinb(w_n76_0[2]),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_G99gat_0[2]),.dinb(w_G71gat_0[2]),.dout(n109),.clk(gclk));
	jxor g037(.dina(w_G43gat_0[2]),.dinb(w_G15gat_0[2]),.dout(n110),.clk(gclk));
	jxor g038(.dina(n110),.dinb(n109),.dout(n111),.clk(gclk));
	jxor g039(.dina(n111),.dinb(w_n99_0[0]),.dout(n112),.clk(gclk));
	jxor g040(.dina(w_n112_0[1]),.dinb(n108),.dout(n113),.clk(gclk));
	jnot g041(.din(w_G228gat_0[1]),.dout(n114),.clk(gclk));
	jor g042(.dina(w_n87_2[1]),.dinb(n114),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(w_n83_0[1]),.dout(n116),.clk(gclk));
	jxor g044(.dina(w_G106gat_0[2]),.dinb(w_G78gat_0[2]),.dout(n117),.clk(gclk));
	jxor g045(.dina(w_G50gat_0[2]),.dinb(w_G22gat_0[2]),.dout(n118),.clk(gclk));
	jxor g046(.dina(n118),.dinb(n117),.dout(n119),.clk(gclk));
	jxor g047(.dina(n119),.dinb(w_n95_0[1]),.dout(n120),.clk(gclk));
	jxor g048(.dina(w_n120_0[1]),.dinb(n116),.dout(n121),.clk(gclk));
	jand g049(.dina(w_n121_0[2]),.dinb(w_n113_0[2]),.dout(n122),.clk(gclk));
	jand g050(.dina(n122),.dinb(n105),.dout(n123),.clk(gclk));
	jxor g051(.dina(w_n121_0[1]),.dinb(w_n113_0[1]),.dout(n124),.clk(gclk));
	jand g052(.dina(w_n104_0[1]),.dinb(w_n90_0[1]),.dout(n125),.clk(gclk));
	jand g053(.dina(n125),.dinb(n124),.dout(n126),.clk(gclk));
	jor g054(.dina(n126),.dinb(n123),.dout(n127),.clk(gclk));
	jand g055(.dina(w_G233gat_3[0]),.dinb(w_G229gat_0[1]),.dout(n128),.clk(gclk));
	jxor g056(.dina(w_G50gat_0[1]),.dinb(w_G43gat_0[1]),.dout(n129),.clk(gclk));
	jxor g057(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n130),.clk(gclk));
	jxor g058(.dina(n130),.dinb(n129),.dout(n131),.clk(gclk));
	jxor g059(.dina(w_n131_1[1]),.dinb(w_dff_B_6HSWmL7A4_1),.dout(n132),.clk(gclk));
	jxor g060(.dina(w_G22gat_0[1]),.dinb(w_G15gat_0[1]),.dout(n133),.clk(gclk));
	jxor g061(.dina(w_G8gat_0[1]),.dinb(w_G1gat_0[1]),.dout(n134),.clk(gclk));
	jxor g062(.dina(n134),.dinb(n133),.dout(n135),.clk(gclk));
	jxor g063(.dina(w_G197gat_0[1]),.dinb(w_G169gat_0[1]),.dout(n136),.clk(gclk));
	jxor g064(.dina(w_G141gat_0[1]),.dinb(w_G113gat_0[1]),.dout(n137),.clk(gclk));
	jxor g065(.dina(n137),.dinb(n136),.dout(n138),.clk(gclk));
	jxor g066(.dina(n138),.dinb(w_n135_0[2]),.dout(n139),.clk(gclk));
	jxor g067(.dina(w_n139_0[1]),.dinb(n132),.dout(n140),.clk(gclk));
	jnot g068(.din(w_G230gat_0[1]),.dout(n141),.clk(gclk));
	jor g069(.dina(w_n87_2[0]),.dinb(n141),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_G106gat_0[1]),.dinb(w_G99gat_0[1]),.dout(n143),.clk(gclk));
	jxor g071(.dina(w_G92gat_0[1]),.dinb(w_G85gat_0[1]),.dout(n144),.clk(gclk));
	jxor g072(.dina(n144),.dinb(n143),.dout(n145),.clk(gclk));
	jxor g073(.dina(w_n145_0[2]),.dinb(n142),.dout(n146),.clk(gclk));
	jxor g074(.dina(w_G78gat_0[1]),.dinb(w_G71gat_0[1]),.dout(n147),.clk(gclk));
	jxor g075(.dina(w_G64gat_0[1]),.dinb(w_G57gat_0[1]),.dout(n148),.clk(gclk));
	jxor g076(.dina(n148),.dinb(n147),.dout(n149),.clk(gclk));
	jxor g077(.dina(w_G204gat_0[1]),.dinb(w_G176gat_0[1]),.dout(n150),.clk(gclk));
	jxor g078(.dina(w_G148gat_0[1]),.dinb(w_G120gat_0[1]),.dout(n151),.clk(gclk));
	jxor g079(.dina(n151),.dinb(n150),.dout(n152),.clk(gclk));
	jxor g080(.dina(n152),.dinb(w_n149_0[1]),.dout(n153),.clk(gclk));
	jxor g081(.dina(w_n153_0[1]),.dinb(n146),.dout(n154),.clk(gclk));
	jand g082(.dina(w_n154_0[2]),.dinb(w_n140_1[2]),.dout(n155),.clk(gclk));
	jnot g083(.din(w_G232gat_0[1]),.dout(n156),.clk(gclk));
	jor g084(.dina(w_n87_1[2]),.dinb(n156),.dout(n157),.clk(gclk));
	jxor g085(.dina(n157),.dinb(w_n131_1[0]),.dout(n158),.clk(gclk));
	jxor g086(.dina(w_G218gat_0[1]),.dinb(w_G190gat_0[1]),.dout(n159),.clk(gclk));
	jxor g087(.dina(w_G162gat_0[1]),.dinb(w_G134gat_0[1]),.dout(n160),.clk(gclk));
	jxor g088(.dina(n160),.dinb(n159),.dout(n161),.clk(gclk));
	jxor g089(.dina(n161),.dinb(w_n145_0[1]),.dout(n162),.clk(gclk));
	jxor g090(.dina(w_n162_0[1]),.dinb(n158),.dout(n163),.clk(gclk));
	jand g091(.dina(w_G233gat_2[2]),.dinb(w_G231gat_0[1]),.dout(n164),.clk(gclk));
	jxor g092(.dina(w_dff_B_gH4FIO5Q8_0),.dinb(w_n135_0[1]),.dout(n165),.clk(gclk));
	jxor g093(.dina(w_G211gat_0[1]),.dinb(w_G183gat_0[1]),.dout(n166),.clk(gclk));
	jxor g094(.dina(w_G155gat_0[1]),.dinb(w_G127gat_0[1]),.dout(n167),.clk(gclk));
	jxor g095(.dina(n167),.dinb(n166),.dout(n168),.clk(gclk));
	jxor g096(.dina(n168),.dinb(w_n149_0[0]),.dout(n169),.clk(gclk));
	jxor g097(.dina(w_n169_0[1]),.dinb(n165),.dout(n170),.clk(gclk));
	jand g098(.dina(w_n170_1[2]),.dinb(w_n163_0[2]),.dout(n171),.clk(gclk));
	jand g099(.dina(w_n171_0[1]),.dinb(w_n155_0[1]),.dout(n172),.clk(gclk));
	jand g100(.dina(w_dff_B_JpMKVmZl9_0),.dinb(w_n127_1[1]),.dout(n173),.clk(gclk));
	jand g101(.dina(w_n173_1[1]),.dinb(w_n85_1[2]),.dout(n174),.clk(gclk));
	jxor g102(.dina(n174),.dinb(w_G1gat_0[0]),.dout(G1324gat),.clk(gclk));
	jand g103(.dina(w_G233gat_2[1]),.dinb(w_G226gat_0[0]),.dout(n176),.clk(gclk));
	jxor g104(.dina(w_n95_0[0]),.dinb(w_dff_B_6PMEPoOn5_1),.dout(n177),.clk(gclk));
	jxor g105(.dina(w_n103_0[0]),.dinb(n177),.dout(n178),.clk(gclk));
	jand g106(.dina(w_n173_1[0]),.dinb(w_n178_1[2]),.dout(n179),.clk(gclk));
	jxor g107(.dina(n179),.dinb(w_G8gat_0[0]),.dout(G1325gat),.clk(gclk));
	jand g108(.dina(w_G233gat_2[0]),.dinb(w_G227gat_0[0]),.dout(n181),.clk(gclk));
	jxor g109(.dina(w_dff_B_qOd2XWaL1_0),.dinb(w_n76_0[1]),.dout(n182),.clk(gclk));
	jxor g110(.dina(w_n112_0[0]),.dinb(n182),.dout(n183),.clk(gclk));
	jand g111(.dina(w_n173_0[2]),.dinb(w_n183_1[2]),.dout(n184),.clk(gclk));
	jxor g112(.dina(n184),.dinb(w_G15gat_0[0]),.dout(G1326gat),.clk(gclk));
	jand g113(.dina(w_G233gat_1[2]),.dinb(w_G228gat_0[0]),.dout(n186),.clk(gclk));
	jxor g114(.dina(w_dff_B_mkSFGFSU5_0),.dinb(w_n83_0[0]),.dout(n187),.clk(gclk));
	jxor g115(.dina(w_n120_0[0]),.dinb(n187),.dout(n188),.clk(gclk));
	jand g116(.dina(w_n173_0[1]),.dinb(w_n188_1[2]),.dout(n189),.clk(gclk));
	jxor g117(.dina(n189),.dinb(w_G22gat_0[0]),.dout(G1327gat),.clk(gclk));
	jand g118(.dina(w_G233gat_1[1]),.dinb(w_G232gat_0[0]),.dout(n191),.clk(gclk));
	jxor g119(.dina(w_dff_B_lGXLKP903_0),.dinb(w_n131_0[2]),.dout(n192),.clk(gclk));
	jxor g120(.dina(w_n162_0[0]),.dinb(n192),.dout(n193),.clk(gclk));
	jnot g121(.din(w_G231gat_0[0]),.dout(n194),.clk(gclk));
	jor g122(.dina(w_n87_1[1]),.dinb(n194),.dout(n195),.clk(gclk));
	jxor g123(.dina(n195),.dinb(w_n135_0[0]),.dout(n196),.clk(gclk));
	jxor g124(.dina(w_n169_0[0]),.dinb(n196),.dout(n197),.clk(gclk));
	jand g125(.dina(w_n197_0[2]),.dinb(w_n193_1[2]),.dout(n198),.clk(gclk));
	jand g126(.dina(w_n198_0[1]),.dinb(w_n155_0[0]),.dout(n199),.clk(gclk));
	jand g127(.dina(w_dff_B_06NNXGq62_0),.dinb(w_n127_1[0]),.dout(n200),.clk(gclk));
	jand g128(.dina(w_n200_1[1]),.dinb(w_n85_1[1]),.dout(n201),.clk(gclk));
	jxor g129(.dina(n201),.dinb(w_G29gat_0[0]),.dout(G1328gat),.clk(gclk));
	jand g130(.dina(w_n200_1[0]),.dinb(w_n178_1[1]),.dout(n203),.clk(gclk));
	jxor g131(.dina(n203),.dinb(w_G36gat_0[0]),.dout(G1329gat),.clk(gclk));
	jand g132(.dina(w_n200_0[2]),.dinb(w_n183_1[1]),.dout(n205),.clk(gclk));
	jxor g133(.dina(n205),.dinb(w_G43gat_0[0]),.dout(G1330gat),.clk(gclk));
	jand g134(.dina(w_n200_0[1]),.dinb(w_n188_1[1]),.dout(n207),.clk(gclk));
	jxor g135(.dina(n207),.dinb(w_G50gat_0[0]),.dout(G1331gat),.clk(gclk));
	jnot g136(.din(w_G229gat_0[0]),.dout(n209),.clk(gclk));
	jor g137(.dina(w_n87_1[0]),.dinb(n209),.dout(n210),.clk(gclk));
	jxor g138(.dina(w_n131_0[1]),.dinb(n210),.dout(n211),.clk(gclk));
	jxor g139(.dina(w_n139_0[0]),.dinb(n211),.dout(n212),.clk(gclk));
	jand g140(.dina(w_G233gat_1[0]),.dinb(w_G230gat_0[0]),.dout(n213),.clk(gclk));
	jxor g141(.dina(w_n145_0[0]),.dinb(w_dff_B_SoJaXzm66_1),.dout(n214),.clk(gclk));
	jxor g142(.dina(w_n153_0[0]),.dinb(n214),.dout(n215),.clk(gclk));
	jand g143(.dina(w_n215_1[2]),.dinb(w_n212_0[2]),.dout(n216),.clk(gclk));
	jand g144(.dina(w_n216_0[1]),.dinb(w_n171_0[0]),.dout(n217),.clk(gclk));
	jand g145(.dina(w_dff_B_btmg2ddw6_0),.dinb(w_n127_0[2]),.dout(n218),.clk(gclk));
	jand g146(.dina(w_n218_1[1]),.dinb(w_n85_1[0]),.dout(n219),.clk(gclk));
	jxor g147(.dina(n219),.dinb(w_G57gat_0[0]),.dout(G1332gat),.clk(gclk));
	jand g148(.dina(w_n218_1[0]),.dinb(w_n178_1[0]),.dout(n221),.clk(gclk));
	jxor g149(.dina(n221),.dinb(w_G64gat_0[0]),.dout(G1333gat),.clk(gclk));
	jand g150(.dina(w_n218_0[2]),.dinb(w_n183_1[0]),.dout(n223),.clk(gclk));
	jxor g151(.dina(n223),.dinb(w_G71gat_0[0]),.dout(G1334gat),.clk(gclk));
	jand g152(.dina(w_n218_0[1]),.dinb(w_n188_1[0]),.dout(n225),.clk(gclk));
	jxor g153(.dina(n225),.dinb(w_G78gat_0[0]),.dout(G1335gat),.clk(gclk));
	jand g154(.dina(w_n216_0[0]),.dinb(w_n198_0[0]),.dout(n227),.clk(gclk));
	jand g155(.dina(w_dff_B_pn2oIhGQ2_0),.dinb(w_n127_0[1]),.dout(n228),.clk(gclk));
	jand g156(.dina(w_n228_1[1]),.dinb(w_n85_0[2]),.dout(n229),.clk(gclk));
	jxor g157(.dina(n229),.dinb(w_G85gat_0[0]),.dout(G1336gat),.clk(gclk));
	jand g158(.dina(w_n228_1[0]),.dinb(w_n178_0[2]),.dout(n231),.clk(gclk));
	jxor g159(.dina(n231),.dinb(w_G92gat_0[0]),.dout(G1337gat),.clk(gclk));
	jand g160(.dina(w_n228_0[2]),.dinb(w_n183_0[2]),.dout(n233),.clk(gclk));
	jxor g161(.dina(n233),.dinb(w_G99gat_0[0]),.dout(G1338gat),.clk(gclk));
	jand g162(.dina(w_n228_0[1]),.dinb(w_n188_0[2]),.dout(n235),.clk(gclk));
	jxor g163(.dina(n235),.dinb(w_G106gat_0[0]),.dout(G1339gat),.clk(gclk));
	jxor g164(.dina(w_n154_0[1]),.dinb(w_n212_0[1]),.dout(n237),.clk(gclk));
	jand g165(.dina(w_n197_0[1]),.dinb(w_n163_0[1]),.dout(n238),.clk(gclk));
	jand g166(.dina(n238),.dinb(n237),.dout(n239),.clk(gclk));
	jxor g167(.dina(w_n197_0[0]),.dinb(w_n163_0[0]),.dout(n240),.clk(gclk));
	jand g168(.dina(w_n154_0[0]),.dinb(w_n212_0[0]),.dout(n241),.clk(gclk));
	jand g169(.dina(n241),.dinb(n240),.dout(n242),.clk(gclk));
	jor g170(.dina(n242),.dinb(n239),.dout(n243),.clk(gclk));
	jand g171(.dina(w_n104_0[0]),.dinb(w_n85_0[1]),.dout(n244),.clk(gclk));
	jand g172(.dina(w_n121_0[0]),.dinb(w_n183_0[1]),.dout(n245),.clk(gclk));
	jand g173(.dina(w_n245_0[1]),.dinb(w_n244_0[1]),.dout(n246),.clk(gclk));
	jand g174(.dina(w_dff_B_2Km8CvHk0_0),.dinb(w_n243_1[1]),.dout(n247),.clk(gclk));
	jand g175(.dina(w_n247_1[1]),.dinb(w_n140_1[1]),.dout(n248),.clk(gclk));
	jxor g176(.dina(n248),.dinb(w_G113gat_0[0]),.dout(G1340gat),.clk(gclk));
	jand g177(.dina(w_n247_1[0]),.dinb(w_n215_1[1]),.dout(n250),.clk(gclk));
	jxor g178(.dina(n250),.dinb(w_G120gat_0[0]),.dout(G1341gat),.clk(gclk));
	jand g179(.dina(w_n247_0[2]),.dinb(w_n170_1[1]),.dout(n252),.clk(gclk));
	jxor g180(.dina(n252),.dinb(w_G127gat_0[0]),.dout(G1342gat),.clk(gclk));
	jand g181(.dina(w_n247_0[1]),.dinb(w_n193_1[1]),.dout(n254),.clk(gclk));
	jxor g182(.dina(n254),.dinb(w_G134gat_0[0]),.dout(G1343gat),.clk(gclk));
	jand g183(.dina(w_n188_0[1]),.dinb(w_n113_0[0]),.dout(n256),.clk(gclk));
	jand g184(.dina(w_n256_0[1]),.dinb(w_n244_0[0]),.dout(n257),.clk(gclk));
	jand g185(.dina(w_dff_B_2INi8XQd3_0),.dinb(w_n243_1[0]),.dout(n258),.clk(gclk));
	jand g186(.dina(w_n258_1[1]),.dinb(w_n140_1[0]),.dout(n259),.clk(gclk));
	jxor g187(.dina(n259),.dinb(w_G141gat_0[0]),.dout(G1344gat),.clk(gclk));
	jand g188(.dina(w_n258_1[0]),.dinb(w_n215_1[0]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_G148gat_0[0]),.dout(G1345gat),.clk(gclk));
	jand g190(.dina(w_n258_0[2]),.dinb(w_n170_1[0]),.dout(n263),.clk(gclk));
	jxor g191(.dina(n263),.dinb(w_G155gat_0[0]),.dout(G1346gat),.clk(gclk));
	jand g192(.dina(w_n258_0[1]),.dinb(w_n193_1[0]),.dout(n265),.clk(gclk));
	jxor g193(.dina(n265),.dinb(w_G162gat_0[0]),.dout(G1347gat),.clk(gclk));
	jand g194(.dina(w_n178_0[1]),.dinb(w_n90_0[0]),.dout(n267),.clk(gclk));
	jand g195(.dina(w_n245_0[0]),.dinb(w_n267_0[1]),.dout(n268),.clk(gclk));
	jand g196(.dina(w_dff_B_1gFbPR9p4_0),.dinb(w_n243_0[2]),.dout(n269),.clk(gclk));
	jand g197(.dina(w_n269_1[1]),.dinb(w_n140_0[2]),.dout(n270),.clk(gclk));
	jxor g198(.dina(n270),.dinb(w_G169gat_0[0]),.dout(G1348gat),.clk(gclk));
	jand g199(.dina(w_n269_1[0]),.dinb(w_n215_0[2]),.dout(n272),.clk(gclk));
	jxor g200(.dina(n272),.dinb(w_G176gat_0[0]),.dout(G1349gat),.clk(gclk));
	jand g201(.dina(w_n269_0[2]),.dinb(w_n170_0[2]),.dout(n274),.clk(gclk));
	jxor g202(.dina(n274),.dinb(w_G183gat_0[0]),.dout(G1350gat),.clk(gclk));
	jand g203(.dina(w_n269_0[1]),.dinb(w_n193_0[2]),.dout(n276),.clk(gclk));
	jxor g204(.dina(n276),.dinb(w_G190gat_0[0]),.dout(G1351gat),.clk(gclk));
	jand g205(.dina(w_n256_0[0]),.dinb(w_n267_0[0]),.dout(n278),.clk(gclk));
	jand g206(.dina(w_dff_B_5ISMQj3O1_0),.dinb(w_n243_0[1]),.dout(n279),.clk(gclk));
	jand g207(.dina(w_n279_1[1]),.dinb(w_n140_0[1]),.dout(n280),.clk(gclk));
	jxor g208(.dina(n280),.dinb(w_G197gat_0[0]),.dout(G1352gat),.clk(gclk));
	jand g209(.dina(w_n279_1[0]),.dinb(w_n215_0[1]),.dout(n282),.clk(gclk));
	jxor g210(.dina(n282),.dinb(w_G204gat_0[0]),.dout(G1353gat),.clk(gclk));
	jand g211(.dina(w_n279_0[2]),.dinb(w_n170_0[1]),.dout(n284),.clk(gclk));
	jxor g212(.dina(n284),.dinb(w_G211gat_0[0]),.dout(G1354gat),.clk(gclk));
	jand g213(.dina(w_n279_0[1]),.dinb(w_n193_0[1]),.dout(n286),.clk(gclk));
	jxor g214(.dina(n286),.dinb(w_G218gat_0[0]),.dout(G1355gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_R1Kk3biT2_0),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_gBnaavUD6_0),.doutb(w_G8gat_0[1]),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G15gat_0(.douta(w_dff_A_1aKUPuaX8_0),.doutb(w_G15gat_0[1]),.doutc(w_G15gat_0[2]),.din(G15gat));
	jspl3 jspl3_w_G22gat_0(.douta(w_dff_A_stWt3Lte9_0),.doutb(w_G22gat_0[1]),.doutc(w_G22gat_0[2]),.din(G22gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_dff_A_SDqRMGgO8_0),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl3 jspl3_w_G36gat_0(.douta(w_dff_A_v7ED5tYc9_0),.doutb(w_G36gat_0[1]),.doutc(w_G36gat_0[2]),.din(G36gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_dff_A_EHOuqmax2_0),.doutb(w_G43gat_0[1]),.doutc(w_G43gat_0[2]),.din(G43gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_dff_A_jrgtPD7H9_0),.doutb(w_G50gat_0[1]),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl3 jspl3_w_G57gat_0(.douta(w_dff_A_vUEa1tOP9_0),.doutb(w_G57gat_0[1]),.doutc(w_G57gat_0[2]),.din(G57gat));
	jspl3 jspl3_w_G64gat_0(.douta(w_dff_A_O0xEvHZB4_0),.doutb(w_G64gat_0[1]),.doutc(w_G64gat_0[2]),.din(G64gat));
	jspl3 jspl3_w_G71gat_0(.douta(w_dff_A_bH14foRf7_0),.doutb(w_G71gat_0[1]),.doutc(w_G71gat_0[2]),.din(G71gat));
	jspl3 jspl3_w_G78gat_0(.douta(w_dff_A_SyaQvzUr9_0),.doutb(w_G78gat_0[1]),.doutc(w_G78gat_0[2]),.din(G78gat));
	jspl3 jspl3_w_G85gat_0(.douta(w_dff_A_VwcYzyRB8_0),.doutb(w_G85gat_0[1]),.doutc(w_G85gat_0[2]),.din(G85gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_jq8KQ46T1_0),.doutb(w_G92gat_0[1]),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_jpqv8m5G6_0),.doutb(w_G99gat_0[1]),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_LGoqKOvX1_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G113gat_0(.douta(w_dff_A_RJtrtdK02_0),.doutb(w_G113gat_0[1]),.doutc(w_G113gat_0[2]),.din(G113gat));
	jspl3 jspl3_w_G120gat_0(.douta(w_dff_A_j9H4W8fS4_0),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G127gat_0(.douta(w_dff_A_OyAPfEGQ2_0),.doutb(w_G127gat_0[1]),.doutc(w_G127gat_0[2]),.din(G127gat));
	jspl3 jspl3_w_G134gat_0(.douta(w_dff_A_R0VlCnVr4_0),.doutb(w_G134gat_0[1]),.doutc(w_G134gat_0[2]),.din(G134gat));
	jspl3 jspl3_w_G141gat_0(.douta(w_dff_A_i5rz0XZO0_0),.doutb(w_G141gat_0[1]),.doutc(w_G141gat_0[2]),.din(G141gat));
	jspl3 jspl3_w_G148gat_0(.douta(w_dff_A_MIJ29XG96_0),.doutb(w_G148gat_0[1]),.doutc(w_G148gat_0[2]),.din(G148gat));
	jspl3 jspl3_w_G155gat_0(.douta(w_dff_A_D6dAaGkh4_0),.doutb(w_G155gat_0[1]),.doutc(w_G155gat_0[2]),.din(G155gat));
	jspl3 jspl3_w_G162gat_0(.douta(w_dff_A_rAX5N1mb8_0),.doutb(w_G162gat_0[1]),.doutc(w_G162gat_0[2]),.din(G162gat));
	jspl3 jspl3_w_G169gat_0(.douta(w_dff_A_fdC9aunC4_0),.doutb(w_G169gat_0[1]),.doutc(w_G169gat_0[2]),.din(G169gat));
	jspl3 jspl3_w_G176gat_0(.douta(w_dff_A_IWKs33zr3_0),.doutb(w_G176gat_0[1]),.doutc(w_G176gat_0[2]),.din(G176gat));
	jspl3 jspl3_w_G183gat_0(.douta(w_dff_A_rk60w1u35_0),.doutb(w_G183gat_0[1]),.doutc(w_G183gat_0[2]),.din(G183gat));
	jspl3 jspl3_w_G190gat_0(.douta(w_dff_A_7bIcqB0f7_0),.doutb(w_G190gat_0[1]),.doutc(w_G190gat_0[2]),.din(G190gat));
	jspl3 jspl3_w_G197gat_0(.douta(w_dff_A_DgsZDsXk0_0),.doutb(w_G197gat_0[1]),.doutc(w_G197gat_0[2]),.din(G197gat));
	jspl3 jspl3_w_G204gat_0(.douta(w_dff_A_Gw2FmiMh0_0),.doutb(w_G204gat_0[1]),.doutc(w_G204gat_0[2]),.din(G204gat));
	jspl3 jspl3_w_G211gat_0(.douta(w_dff_A_PxtJZ94Q4_0),.doutb(w_G211gat_0[1]),.doutc(w_G211gat_0[2]),.din(G211gat));
	jspl3 jspl3_w_G218gat_0(.douta(w_dff_A_4ix7yO1c6_0),.doutb(w_G218gat_0[1]),.doutc(w_G218gat_0[2]),.din(G218gat));
	jspl jspl_w_G225gat_0(.douta(w_G225gat_0[0]),.doutb(w_G225gat_0[1]),.din(G225gat));
	jspl jspl_w_G226gat_0(.douta(w_G226gat_0[0]),.doutb(w_G226gat_0[1]),.din(G226gat));
	jspl jspl_w_G227gat_0(.douta(w_G227gat_0[0]),.doutb(w_G227gat_0[1]),.din(G227gat));
	jspl jspl_w_G228gat_0(.douta(w_G228gat_0[0]),.doutb(w_G228gat_0[1]),.din(G228gat));
	jspl jspl_w_G229gat_0(.douta(w_G229gat_0[0]),.doutb(w_G229gat_0[1]),.din(G229gat));
	jspl jspl_w_G230gat_0(.douta(w_G230gat_0[0]),.doutb(w_G230gat_0[1]),.din(G230gat));
	jspl jspl_w_G231gat_0(.douta(w_G231gat_0[0]),.doutb(w_G231gat_0[1]),.din(G231gat));
	jspl jspl_w_G232gat_0(.douta(w_G232gat_0[0]),.doutb(w_G232gat_0[1]),.din(G232gat));
	jspl3 jspl3_w_G233gat_0(.douta(w_G233gat_0[0]),.doutb(w_G233gat_0[1]),.doutc(w_G233gat_0[2]),.din(G233gat));
	jspl3 jspl3_w_G233gat_1(.douta(w_G233gat_1[0]),.doutb(w_G233gat_1[1]),.doutc(w_G233gat_1[2]),.din(w_G233gat_0[0]));
	jspl3 jspl3_w_G233gat_2(.douta(w_G233gat_2[0]),.doutb(w_G233gat_2[1]),.doutc(w_G233gat_2[2]),.din(w_G233gat_0[1]));
	jspl3 jspl3_w_G233gat_3(.douta(w_G233gat_3[0]),.doutb(w_G233gat_3[1]),.doutc(w_G233gat_3[2]),.din(w_G233gat_0[2]));
	jspl3 jspl3_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.doutc(w_n76_0[2]),.din(n76));
	jspl jspl_w_n76_1(.douta(w_n76_1[0]),.doutb(w_n76_1[1]),.din(w_n76_0[0]));
	jspl3 jspl3_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.doutc(w_n83_0[2]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_InqPmjAf2_0),.doutb(w_n85_0[1]),.doutc(w_dff_A_jWD4RRAF2_2),.din(n85));
	jspl3 jspl3_w_n85_1(.douta(w_n85_1[0]),.doutb(w_n85_1[1]),.doutc(w_n85_1[2]),.din(w_n85_0[0]));
	jspl3 jspl3_w_n87_0(.douta(w_n87_0[0]),.doutb(w_n87_0[1]),.doutc(w_n87_0[2]),.din(n87));
	jspl3 jspl3_w_n87_1(.douta(w_n87_1[0]),.doutb(w_n87_1[1]),.doutc(w_n87_1[2]),.din(w_n87_0[0]));
	jspl3 jspl3_w_n87_2(.douta(w_n87_2[0]),.doutb(w_n87_2[1]),.doutc(w_n87_2[2]),.din(w_n87_0[1]));
	jspl jspl_w_n87_3(.douta(w_n87_3[0]),.doutb(w_n87_3[1]),.din(w_n87_0[2]));
	jspl3 jspl3_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n95_0(.douta(w_n95_0[0]),.doutb(w_n95_0[1]),.doutc(w_n95_0[2]),.din(n95));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.din(n103));
	jspl3 jspl3_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.doutc(w_n104_0[2]),.din(n104));
	jspl jspl_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.doutc(w_n113_0[2]),.din(n113));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.doutc(w_n127_0[2]),.din(n127));
	jspl jspl_w_n127_1(.douta(w_n127_1[0]),.doutb(w_n127_1[1]),.din(w_n127_0[0]));
	jspl3 jspl3_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.doutc(w_n131_0[2]),.din(n131));
	jspl jspl_w_n131_1(.douta(w_n131_1[0]),.doutb(w_n131_1[1]),.din(w_n131_0[0]));
	jspl3 jspl3_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.doutc(w_n135_0[2]),.din(n135));
	jspl jspl_w_n139_0(.douta(w_n139_0[0]),.doutb(w_n139_0[1]),.din(n139));
	jspl3 jspl3_w_n140_0(.douta(w_n140_0[0]),.doutb(w_dff_A_gz6QLfLj0_1),.doutc(w_dff_A_9jk7SHR34_2),.din(n140));
	jspl3 jspl3_w_n140_1(.douta(w_dff_A_af33HeQj4_0),.doutb(w_dff_A_HjKQHrjl4_1),.doutc(w_n140_1[2]),.din(w_n140_0[0]));
	jspl3 jspl3_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.doutc(w_n145_0[2]),.din(n145));
	jspl jspl_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.din(n149));
	jspl jspl_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.din(n153));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_n154_0[2]),.din(n154));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_n163_0[2]),.din(n163));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_dff_A_wRehXAhG7_1),.doutc(w_dff_A_zPPLunni8_2),.din(n170));
	jspl3 jspl3_w_n170_1(.douta(w_dff_A_RjilLUSm9_0),.doutb(w_dff_A_TP2le7tE4_1),.doutc(w_n170_1[2]),.din(w_n170_0[0]));
	jspl jspl_w_n171_0(.douta(w_n171_0[0]),.doutb(w_n171_0[1]),.din(n171));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl jspl_w_n173_1(.douta(w_n173_1[0]),.doutb(w_n173_1[1]),.din(w_n173_0[0]));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_agrTuzZR9_0),.doutb(w_n178_0[1]),.doutc(w_dff_A_3jjv8xX07_2),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_n178_1[1]),.doutc(w_n178_1[2]),.din(w_n178_0[0]));
	jspl3 jspl3_w_n183_0(.douta(w_dff_A_vjFuTVfN7_0),.doutb(w_n183_0[1]),.doutc(w_dff_A_rEuNCYgm9_2),.din(n183));
	jspl3 jspl3_w_n183_1(.douta(w_n183_1[0]),.doutb(w_n183_1[1]),.doutc(w_n183_1[2]),.din(w_n183_0[0]));
	jspl3 jspl3_w_n188_0(.douta(w_dff_A_zFHeq7ah5_0),.doutb(w_n188_0[1]),.doutc(w_dff_A_oSDLP5Yh7_2),.din(n188));
	jspl3 jspl3_w_n188_1(.douta(w_n188_1[0]),.doutb(w_n188_1[1]),.doutc(w_n188_1[2]),.din(w_n188_0[0]));
	jspl3 jspl3_w_n193_0(.douta(w_n193_0[0]),.doutb(w_dff_A_mXsTGYGu8_1),.doutc(w_dff_A_zHWUR9p43_2),.din(n193));
	jspl3 jspl3_w_n193_1(.douta(w_dff_A_hmGuCVsx1_0),.doutb(w_dff_A_Gmtn59Zy1_1),.doutc(w_n193_1[2]),.din(w_n193_0[0]));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl3 jspl3_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.doutc(w_n200_0[2]),.din(n200));
	jspl jspl_w_n200_1(.douta(w_n200_1[0]),.doutb(w_n200_1[1]),.din(w_n200_0[0]));
	jspl3 jspl3_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.doutc(w_n212_0[2]),.din(n212));
	jspl3 jspl3_w_n215_0(.douta(w_n215_0[0]),.doutb(w_dff_A_gtr1tQUw2_1),.doutc(w_dff_A_mPztUbUJ7_2),.din(n215));
	jspl3 jspl3_w_n215_1(.douta(w_dff_A_SReMXxCA6_0),.doutb(w_dff_A_tX3pqyub1_1),.doutc(w_n215_1[2]),.din(w_n215_0[0]));
	jspl jspl_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.din(n216));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_n218_0[2]),.din(n218));
	jspl jspl_w_n218_1(.douta(w_n218_1[0]),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl3 jspl3_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.doutc(w_n228_0[2]),.din(n228));
	jspl jspl_w_n228_1(.douta(w_n228_1[0]),.doutb(w_n228_1[1]),.din(w_n228_0[0]));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n243_1(.douta(w_n243_1[0]),.doutb(w_n243_1[1]),.din(w_n243_0[0]));
	jspl jspl_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.din(n244));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl3 jspl3_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.doutc(w_n247_0[2]),.din(n247));
	jspl jspl_w_n247_1(.douta(w_n247_1[0]),.doutb(w_n247_1[1]),.din(w_n247_0[0]));
	jspl jspl_w_n256_0(.douta(w_n256_0[0]),.doutb(w_n256_0[1]),.din(n256));
	jspl3 jspl3_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.doutc(w_n258_0[2]),.din(n258));
	jspl jspl_w_n258_1(.douta(w_n258_1[0]),.doutb(w_n258_1[1]),.din(w_n258_0[0]));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(n267));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl jspl_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.din(w_n269_0[0]));
	jspl3 jspl3_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.doutc(w_n279_0[2]),.din(n279));
	jspl jspl_w_n279_1(.douta(w_n279_1[0]),.doutb(w_n279_1[1]),.din(w_n279_0[0]));
	jdff dff_B_JpMKVmZl9_0(.din(n172),.dout(w_dff_B_JpMKVmZl9_0),.clk(gclk));
	jdff dff_B_06NNXGq62_0(.din(n199),.dout(w_dff_B_06NNXGq62_0),.clk(gclk));
	jdff dff_B_btmg2ddw6_0(.din(n217),.dout(w_dff_B_btmg2ddw6_0),.clk(gclk));
	jdff dff_B_pn2oIhGQ2_0(.din(n227),.dout(w_dff_B_pn2oIhGQ2_0),.clk(gclk));
	jdff dff_B_2Km8CvHk0_0(.din(n246),.dout(w_dff_B_2Km8CvHk0_0),.clk(gclk));
	jdff dff_A_UEFCxbK25_0(.dout(w_n140_1[0]),.din(w_dff_A_UEFCxbK25_0),.clk(gclk));
	jdff dff_A_g1BfgCzT0_0(.dout(w_dff_A_UEFCxbK25_0),.din(w_dff_A_g1BfgCzT0_0),.clk(gclk));
	jdff dff_A_v7xPrecR9_0(.dout(w_dff_A_g1BfgCzT0_0),.din(w_dff_A_v7xPrecR9_0),.clk(gclk));
	jdff dff_A_af33HeQj4_0(.dout(w_dff_A_v7xPrecR9_0),.din(w_dff_A_af33HeQj4_0),.clk(gclk));
	jdff dff_A_ZlG0OEia8_1(.dout(w_n140_1[1]),.din(w_dff_A_ZlG0OEia8_1),.clk(gclk));
	jdff dff_A_cUtTnJo07_1(.dout(w_dff_A_ZlG0OEia8_1),.din(w_dff_A_cUtTnJo07_1),.clk(gclk));
	jdff dff_A_PJl0B6a46_1(.dout(w_dff_A_cUtTnJo07_1),.din(w_dff_A_PJl0B6a46_1),.clk(gclk));
	jdff dff_A_HjKQHrjl4_1(.dout(w_dff_A_PJl0B6a46_1),.din(w_dff_A_HjKQHrjl4_1),.clk(gclk));
	jdff dff_A_nlWAvpXB4_0(.dout(w_n215_1[0]),.din(w_dff_A_nlWAvpXB4_0),.clk(gclk));
	jdff dff_A_xT1L5ZQw9_0(.dout(w_dff_A_nlWAvpXB4_0),.din(w_dff_A_xT1L5ZQw9_0),.clk(gclk));
	jdff dff_A_rPUdUG9W3_0(.dout(w_dff_A_xT1L5ZQw9_0),.din(w_dff_A_rPUdUG9W3_0),.clk(gclk));
	jdff dff_A_SReMXxCA6_0(.dout(w_dff_A_rPUdUG9W3_0),.din(w_dff_A_SReMXxCA6_0),.clk(gclk));
	jdff dff_A_GYNK3MhN6_1(.dout(w_n215_1[1]),.din(w_dff_A_GYNK3MhN6_1),.clk(gclk));
	jdff dff_A_1MgGcnkf2_1(.dout(w_dff_A_GYNK3MhN6_1),.din(w_dff_A_1MgGcnkf2_1),.clk(gclk));
	jdff dff_A_J2Qlhlvh1_1(.dout(w_dff_A_1MgGcnkf2_1),.din(w_dff_A_J2Qlhlvh1_1),.clk(gclk));
	jdff dff_A_tX3pqyub1_1(.dout(w_dff_A_J2Qlhlvh1_1),.din(w_dff_A_tX3pqyub1_1),.clk(gclk));
	jdff dff_A_VUZMEUK57_0(.dout(w_n170_1[0]),.din(w_dff_A_VUZMEUK57_0),.clk(gclk));
	jdff dff_A_C2tTUdFW9_0(.dout(w_dff_A_VUZMEUK57_0),.din(w_dff_A_C2tTUdFW9_0),.clk(gclk));
	jdff dff_A_hlETrfwt2_0(.dout(w_dff_A_C2tTUdFW9_0),.din(w_dff_A_hlETrfwt2_0),.clk(gclk));
	jdff dff_A_RjilLUSm9_0(.dout(w_dff_A_hlETrfwt2_0),.din(w_dff_A_RjilLUSm9_0),.clk(gclk));
	jdff dff_A_zmb6Iz487_1(.dout(w_n170_1[1]),.din(w_dff_A_zmb6Iz487_1),.clk(gclk));
	jdff dff_A_RpJ5IAsl3_1(.dout(w_dff_A_zmb6Iz487_1),.din(w_dff_A_RpJ5IAsl3_1),.clk(gclk));
	jdff dff_A_vZXhAKHK9_1(.dout(w_dff_A_RpJ5IAsl3_1),.din(w_dff_A_vZXhAKHK9_1),.clk(gclk));
	jdff dff_A_TP2le7tE4_1(.dout(w_dff_A_vZXhAKHK9_1),.din(w_dff_A_TP2le7tE4_1),.clk(gclk));
	jdff dff_B_2INi8XQd3_0(.din(n257),.dout(w_dff_B_2INi8XQd3_0),.clk(gclk));
	jdff dff_A_ITY20qju2_0(.dout(w_n85_0[0]),.din(w_dff_A_ITY20qju2_0),.clk(gclk));
	jdff dff_A_XPZNI1cD3_0(.dout(w_dff_A_ITY20qju2_0),.din(w_dff_A_XPZNI1cD3_0),.clk(gclk));
	jdff dff_A_alsCGyvt9_0(.dout(w_dff_A_XPZNI1cD3_0),.din(w_dff_A_alsCGyvt9_0),.clk(gclk));
	jdff dff_A_InqPmjAf2_0(.dout(w_dff_A_alsCGyvt9_0),.din(w_dff_A_InqPmjAf2_0),.clk(gclk));
	jdff dff_A_hjOrORjM4_2(.dout(w_n85_0[2]),.din(w_dff_A_hjOrORjM4_2),.clk(gclk));
	jdff dff_A_Zzioavus5_2(.dout(w_dff_A_hjOrORjM4_2),.din(w_dff_A_Zzioavus5_2),.clk(gclk));
	jdff dff_A_05lu8w600_2(.dout(w_dff_A_Zzioavus5_2),.din(w_dff_A_05lu8w600_2),.clk(gclk));
	jdff dff_A_jWD4RRAF2_2(.dout(w_dff_A_05lu8w600_2),.din(w_dff_A_jWD4RRAF2_2),.clk(gclk));
	jdff dff_B_pdYoucrR6_1(.din(n73),.dout(w_dff_B_pdYoucrR6_1),.clk(gclk));
	jdff dff_A_9yOWnLIP5_0(.dout(w_n193_1[0]),.din(w_dff_A_9yOWnLIP5_0),.clk(gclk));
	jdff dff_A_4iPUKJBz0_0(.dout(w_dff_A_9yOWnLIP5_0),.din(w_dff_A_4iPUKJBz0_0),.clk(gclk));
	jdff dff_A_3BJoGveC8_0(.dout(w_dff_A_4iPUKJBz0_0),.din(w_dff_A_3BJoGveC8_0),.clk(gclk));
	jdff dff_A_hmGuCVsx1_0(.dout(w_dff_A_3BJoGveC8_0),.din(w_dff_A_hmGuCVsx1_0),.clk(gclk));
	jdff dff_A_jkZrImb09_1(.dout(w_n193_1[1]),.din(w_dff_A_jkZrImb09_1),.clk(gclk));
	jdff dff_A_xpcBif0g1_1(.dout(w_dff_A_jkZrImb09_1),.din(w_dff_A_xpcBif0g1_1),.clk(gclk));
	jdff dff_A_8qybLMO87_1(.dout(w_dff_A_xpcBif0g1_1),.din(w_dff_A_8qybLMO87_1),.clk(gclk));
	jdff dff_A_Gmtn59Zy1_1(.dout(w_dff_A_8qybLMO87_1),.din(w_dff_A_Gmtn59Zy1_1),.clk(gclk));
	jdff dff_B_1gFbPR9p4_0(.din(n268),.dout(w_dff_B_1gFbPR9p4_0),.clk(gclk));
	jdff dff_A_vDuh33W94_0(.dout(w_n183_0[0]),.din(w_dff_A_vDuh33W94_0),.clk(gclk));
	jdff dff_A_CuHLstmq1_0(.dout(w_dff_A_vDuh33W94_0),.din(w_dff_A_CuHLstmq1_0),.clk(gclk));
	jdff dff_A_iMxb8M8i4_0(.dout(w_dff_A_CuHLstmq1_0),.din(w_dff_A_iMxb8M8i4_0),.clk(gclk));
	jdff dff_A_vjFuTVfN7_0(.dout(w_dff_A_iMxb8M8i4_0),.din(w_dff_A_vjFuTVfN7_0),.clk(gclk));
	jdff dff_A_Q3bxO8ma6_2(.dout(w_n183_0[2]),.din(w_dff_A_Q3bxO8ma6_2),.clk(gclk));
	jdff dff_A_gTpzAnOG5_2(.dout(w_dff_A_Q3bxO8ma6_2),.din(w_dff_A_gTpzAnOG5_2),.clk(gclk));
	jdff dff_A_bpEI5ce25_2(.dout(w_dff_A_gTpzAnOG5_2),.din(w_dff_A_bpEI5ce25_2),.clk(gclk));
	jdff dff_A_rEuNCYgm9_2(.dout(w_dff_A_bpEI5ce25_2),.din(w_dff_A_rEuNCYgm9_2),.clk(gclk));
	jdff dff_B_qOd2XWaL1_0(.din(n181),.dout(w_dff_B_qOd2XWaL1_0),.clk(gclk));
	jdff dff_A_Kxc47GtV0_1(.dout(w_n140_0[1]),.din(w_dff_A_Kxc47GtV0_1),.clk(gclk));
	jdff dff_A_iBZDce420_1(.dout(w_dff_A_Kxc47GtV0_1),.din(w_dff_A_iBZDce420_1),.clk(gclk));
	jdff dff_A_jH4meBDb6_1(.dout(w_dff_A_iBZDce420_1),.din(w_dff_A_jH4meBDb6_1),.clk(gclk));
	jdff dff_A_gz6QLfLj0_1(.dout(w_dff_A_jH4meBDb6_1),.din(w_dff_A_gz6QLfLj0_1),.clk(gclk));
	jdff dff_A_EovRSw7Z5_2(.dout(w_n140_0[2]),.din(w_dff_A_EovRSw7Z5_2),.clk(gclk));
	jdff dff_A_l73MpFsM3_2(.dout(w_dff_A_EovRSw7Z5_2),.din(w_dff_A_l73MpFsM3_2),.clk(gclk));
	jdff dff_A_5mg9CYSE6_2(.dout(w_dff_A_l73MpFsM3_2),.din(w_dff_A_5mg9CYSE6_2),.clk(gclk));
	jdff dff_A_9jk7SHR34_2(.dout(w_dff_A_5mg9CYSE6_2),.din(w_dff_A_9jk7SHR34_2),.clk(gclk));
	jdff dff_B_6HSWmL7A4_1(.din(n128),.dout(w_dff_B_6HSWmL7A4_1),.clk(gclk));
	jdff dff_A_6wht6jjS9_1(.dout(w_n215_0[1]),.din(w_dff_A_6wht6jjS9_1),.clk(gclk));
	jdff dff_A_CuUeb5F64_1(.dout(w_dff_A_6wht6jjS9_1),.din(w_dff_A_CuUeb5F64_1),.clk(gclk));
	jdff dff_A_4sK58bz96_1(.dout(w_dff_A_CuUeb5F64_1),.din(w_dff_A_4sK58bz96_1),.clk(gclk));
	jdff dff_A_gtr1tQUw2_1(.dout(w_dff_A_4sK58bz96_1),.din(w_dff_A_gtr1tQUw2_1),.clk(gclk));
	jdff dff_A_QiFr9GKJ0_2(.dout(w_n215_0[2]),.din(w_dff_A_QiFr9GKJ0_2),.clk(gclk));
	jdff dff_A_L0zuODby1_2(.dout(w_dff_A_QiFr9GKJ0_2),.din(w_dff_A_L0zuODby1_2),.clk(gclk));
	jdff dff_A_FOmorWB30_2(.dout(w_dff_A_L0zuODby1_2),.din(w_dff_A_FOmorWB30_2),.clk(gclk));
	jdff dff_A_mPztUbUJ7_2(.dout(w_dff_A_FOmorWB30_2),.din(w_dff_A_mPztUbUJ7_2),.clk(gclk));
	jdff dff_B_SoJaXzm66_1(.din(n213),.dout(w_dff_B_SoJaXzm66_1),.clk(gclk));
	jdff dff_A_rszApFuE6_1(.dout(w_n170_0[1]),.din(w_dff_A_rszApFuE6_1),.clk(gclk));
	jdff dff_A_CJhm6qde5_1(.dout(w_dff_A_rszApFuE6_1),.din(w_dff_A_CJhm6qde5_1),.clk(gclk));
	jdff dff_A_QZ4juBak6_1(.dout(w_dff_A_CJhm6qde5_1),.din(w_dff_A_QZ4juBak6_1),.clk(gclk));
	jdff dff_A_wRehXAhG7_1(.dout(w_dff_A_QZ4juBak6_1),.din(w_dff_A_wRehXAhG7_1),.clk(gclk));
	jdff dff_A_bUlwPINx4_2(.dout(w_n170_0[2]),.din(w_dff_A_bUlwPINx4_2),.clk(gclk));
	jdff dff_A_QseusKqf2_2(.dout(w_dff_A_bUlwPINx4_2),.din(w_dff_A_QseusKqf2_2),.clk(gclk));
	jdff dff_A_GzkFXzdh3_2(.dout(w_dff_A_QseusKqf2_2),.din(w_dff_A_GzkFXzdh3_2),.clk(gclk));
	jdff dff_A_zPPLunni8_2(.dout(w_dff_A_GzkFXzdh3_2),.din(w_dff_A_zPPLunni8_2),.clk(gclk));
	jdff dff_B_gH4FIO5Q8_0(.din(n164),.dout(w_dff_B_gH4FIO5Q8_0),.clk(gclk));
	jdff dff_B_5ISMQj3O1_0(.din(n278),.dout(w_dff_B_5ISMQj3O1_0),.clk(gclk));
	jdff dff_A_Jh1Vr3280_0(.dout(w_n188_0[0]),.din(w_dff_A_Jh1Vr3280_0),.clk(gclk));
	jdff dff_A_aAIfW8Qg4_0(.dout(w_dff_A_Jh1Vr3280_0),.din(w_dff_A_aAIfW8Qg4_0),.clk(gclk));
	jdff dff_A_QlTneZLs8_0(.dout(w_dff_A_aAIfW8Qg4_0),.din(w_dff_A_QlTneZLs8_0),.clk(gclk));
	jdff dff_A_zFHeq7ah5_0(.dout(w_dff_A_QlTneZLs8_0),.din(w_dff_A_zFHeq7ah5_0),.clk(gclk));
	jdff dff_A_J7XXJgdO6_2(.dout(w_n188_0[2]),.din(w_dff_A_J7XXJgdO6_2),.clk(gclk));
	jdff dff_A_BC676bst6_2(.dout(w_dff_A_J7XXJgdO6_2),.din(w_dff_A_BC676bst6_2),.clk(gclk));
	jdff dff_A_oGmJaPL98_2(.dout(w_dff_A_BC676bst6_2),.din(w_dff_A_oGmJaPL98_2),.clk(gclk));
	jdff dff_A_oSDLP5Yh7_2(.dout(w_dff_A_oGmJaPL98_2),.din(w_dff_A_oSDLP5Yh7_2),.clk(gclk));
	jdff dff_B_mkSFGFSU5_0(.din(n186),.dout(w_dff_B_mkSFGFSU5_0),.clk(gclk));
	jdff dff_A_rTPmh6yz8_0(.dout(w_n178_0[0]),.din(w_dff_A_rTPmh6yz8_0),.clk(gclk));
	jdff dff_A_OUnsK4da7_0(.dout(w_dff_A_rTPmh6yz8_0),.din(w_dff_A_OUnsK4da7_0),.clk(gclk));
	jdff dff_A_NuFlGr284_0(.dout(w_dff_A_OUnsK4da7_0),.din(w_dff_A_NuFlGr284_0),.clk(gclk));
	jdff dff_A_agrTuzZR9_0(.dout(w_dff_A_NuFlGr284_0),.din(w_dff_A_agrTuzZR9_0),.clk(gclk));
	jdff dff_A_NYSv60IV8_2(.dout(w_n178_0[2]),.din(w_dff_A_NYSv60IV8_2),.clk(gclk));
	jdff dff_A_9U3ZkJ0I8_2(.dout(w_dff_A_NYSv60IV8_2),.din(w_dff_A_9U3ZkJ0I8_2),.clk(gclk));
	jdff dff_A_1WSdQZiH5_2(.dout(w_dff_A_9U3ZkJ0I8_2),.din(w_dff_A_1WSdQZiH5_2),.clk(gclk));
	jdff dff_A_3jjv8xX07_2(.dout(w_dff_A_1WSdQZiH5_2),.din(w_dff_A_3jjv8xX07_2),.clk(gclk));
	jdff dff_B_6PMEPoOn5_1(.din(n176),.dout(w_dff_B_6PMEPoOn5_1),.clk(gclk));
	jdff dff_A_KbrTgli03_0(.dout(w_G155gat_0[0]),.din(w_dff_A_KbrTgli03_0),.clk(gclk));
	jdff dff_A_Eet2dHw20_0(.dout(w_dff_A_KbrTgli03_0),.din(w_dff_A_Eet2dHw20_0),.clk(gclk));
	jdff dff_A_x1mHxHrO7_0(.dout(w_dff_A_Eet2dHw20_0),.din(w_dff_A_x1mHxHrO7_0),.clk(gclk));
	jdff dff_A_2ukqXYEG5_0(.dout(w_dff_A_x1mHxHrO7_0),.din(w_dff_A_2ukqXYEG5_0),.clk(gclk));
	jdff dff_A_EIvQluIV0_0(.dout(w_dff_A_2ukqXYEG5_0),.din(w_dff_A_EIvQluIV0_0),.clk(gclk));
	jdff dff_A_QI1EBWci3_0(.dout(w_dff_A_EIvQluIV0_0),.din(w_dff_A_QI1EBWci3_0),.clk(gclk));
	jdff dff_A_BILdSeYm1_0(.dout(w_dff_A_QI1EBWci3_0),.din(w_dff_A_BILdSeYm1_0),.clk(gclk));
	jdff dff_A_H4KCkzPz9_0(.dout(w_dff_A_BILdSeYm1_0),.din(w_dff_A_H4KCkzPz9_0),.clk(gclk));
	jdff dff_A_D6dAaGkh4_0(.dout(w_dff_A_H4KCkzPz9_0),.din(w_dff_A_D6dAaGkh4_0),.clk(gclk));
	jdff dff_A_v25iy4EA9_0(.dout(w_G127gat_0[0]),.din(w_dff_A_v25iy4EA9_0),.clk(gclk));
	jdff dff_A_6ws0EdZG4_0(.dout(w_dff_A_v25iy4EA9_0),.din(w_dff_A_6ws0EdZG4_0),.clk(gclk));
	jdff dff_A_9npPaJRl3_0(.dout(w_dff_A_6ws0EdZG4_0),.din(w_dff_A_9npPaJRl3_0),.clk(gclk));
	jdff dff_A_rKPIajl82_0(.dout(w_dff_A_9npPaJRl3_0),.din(w_dff_A_rKPIajl82_0),.clk(gclk));
	jdff dff_A_fRmLfm376_0(.dout(w_dff_A_rKPIajl82_0),.din(w_dff_A_fRmLfm376_0),.clk(gclk));
	jdff dff_A_3apjY6hn4_0(.dout(w_dff_A_fRmLfm376_0),.din(w_dff_A_3apjY6hn4_0),.clk(gclk));
	jdff dff_A_ANKXSSDB1_0(.dout(w_dff_A_3apjY6hn4_0),.din(w_dff_A_ANKXSSDB1_0),.clk(gclk));
	jdff dff_A_3BNT17BE6_0(.dout(w_dff_A_ANKXSSDB1_0),.din(w_dff_A_3BNT17BE6_0),.clk(gclk));
	jdff dff_A_OyAPfEGQ2_0(.dout(w_dff_A_3BNT17BE6_0),.din(w_dff_A_OyAPfEGQ2_0),.clk(gclk));
	jdff dff_A_rphy6nna1_0(.dout(w_G211gat_0[0]),.din(w_dff_A_rphy6nna1_0),.clk(gclk));
	jdff dff_A_vhP9Nzv64_0(.dout(w_dff_A_rphy6nna1_0),.din(w_dff_A_vhP9Nzv64_0),.clk(gclk));
	jdff dff_A_XQXlRbjK0_0(.dout(w_dff_A_vhP9Nzv64_0),.din(w_dff_A_XQXlRbjK0_0),.clk(gclk));
	jdff dff_A_cM2lksrO9_0(.dout(w_dff_A_XQXlRbjK0_0),.din(w_dff_A_cM2lksrO9_0),.clk(gclk));
	jdff dff_A_uQmCCl9M8_0(.dout(w_dff_A_cM2lksrO9_0),.din(w_dff_A_uQmCCl9M8_0),.clk(gclk));
	jdff dff_A_lVWX8ZPp5_0(.dout(w_dff_A_uQmCCl9M8_0),.din(w_dff_A_lVWX8ZPp5_0),.clk(gclk));
	jdff dff_A_fizDFYwF0_0(.dout(w_dff_A_lVWX8ZPp5_0),.din(w_dff_A_fizDFYwF0_0),.clk(gclk));
	jdff dff_A_rkxtQIjF0_0(.dout(w_dff_A_fizDFYwF0_0),.din(w_dff_A_rkxtQIjF0_0),.clk(gclk));
	jdff dff_A_PxtJZ94Q4_0(.dout(w_dff_A_rkxtQIjF0_0),.din(w_dff_A_PxtJZ94Q4_0),.clk(gclk));
	jdff dff_A_Q7Uv4kNI6_0(.dout(w_G183gat_0[0]),.din(w_dff_A_Q7Uv4kNI6_0),.clk(gclk));
	jdff dff_A_PU5o12Yv5_0(.dout(w_dff_A_Q7Uv4kNI6_0),.din(w_dff_A_PU5o12Yv5_0),.clk(gclk));
	jdff dff_A_gK9Yriil2_0(.dout(w_dff_A_PU5o12Yv5_0),.din(w_dff_A_gK9Yriil2_0),.clk(gclk));
	jdff dff_A_FRlZvOYt1_0(.dout(w_dff_A_gK9Yriil2_0),.din(w_dff_A_FRlZvOYt1_0),.clk(gclk));
	jdff dff_A_ZotPLopL7_0(.dout(w_dff_A_FRlZvOYt1_0),.din(w_dff_A_ZotPLopL7_0),.clk(gclk));
	jdff dff_A_yTmacIWl0_0(.dout(w_dff_A_ZotPLopL7_0),.din(w_dff_A_yTmacIWl0_0),.clk(gclk));
	jdff dff_A_JRw8BJae0_0(.dout(w_dff_A_yTmacIWl0_0),.din(w_dff_A_JRw8BJae0_0),.clk(gclk));
	jdff dff_A_O0GHoQSB5_0(.dout(w_dff_A_JRw8BJae0_0),.din(w_dff_A_O0GHoQSB5_0),.clk(gclk));
	jdff dff_A_rk60w1u35_0(.dout(w_dff_A_O0GHoQSB5_0),.din(w_dff_A_rk60w1u35_0),.clk(gclk));
	jdff dff_A_GafMvStw1_0(.dout(w_G148gat_0[0]),.din(w_dff_A_GafMvStw1_0),.clk(gclk));
	jdff dff_A_Ot2yuFw25_0(.dout(w_dff_A_GafMvStw1_0),.din(w_dff_A_Ot2yuFw25_0),.clk(gclk));
	jdff dff_A_4p02WoLu4_0(.dout(w_dff_A_Ot2yuFw25_0),.din(w_dff_A_4p02WoLu4_0),.clk(gclk));
	jdff dff_A_izpkRR5Q9_0(.dout(w_dff_A_4p02WoLu4_0),.din(w_dff_A_izpkRR5Q9_0),.clk(gclk));
	jdff dff_A_GFJ60qxS4_0(.dout(w_dff_A_izpkRR5Q9_0),.din(w_dff_A_GFJ60qxS4_0),.clk(gclk));
	jdff dff_A_LH3URp8V9_0(.dout(w_dff_A_GFJ60qxS4_0),.din(w_dff_A_LH3URp8V9_0),.clk(gclk));
	jdff dff_A_9Q0hwyxl1_0(.dout(w_dff_A_LH3URp8V9_0),.din(w_dff_A_9Q0hwyxl1_0),.clk(gclk));
	jdff dff_A_eMLKePgr5_0(.dout(w_dff_A_9Q0hwyxl1_0),.din(w_dff_A_eMLKePgr5_0),.clk(gclk));
	jdff dff_A_MIJ29XG96_0(.dout(w_dff_A_eMLKePgr5_0),.din(w_dff_A_MIJ29XG96_0),.clk(gclk));
	jdff dff_A_JmQdnqEg1_0(.dout(w_G120gat_0[0]),.din(w_dff_A_JmQdnqEg1_0),.clk(gclk));
	jdff dff_A_dV1zL4912_0(.dout(w_dff_A_JmQdnqEg1_0),.din(w_dff_A_dV1zL4912_0),.clk(gclk));
	jdff dff_A_CQGlUN0V0_0(.dout(w_dff_A_dV1zL4912_0),.din(w_dff_A_CQGlUN0V0_0),.clk(gclk));
	jdff dff_A_yHdzh8Fy5_0(.dout(w_dff_A_CQGlUN0V0_0),.din(w_dff_A_yHdzh8Fy5_0),.clk(gclk));
	jdff dff_A_JsB1D3RH3_0(.dout(w_dff_A_yHdzh8Fy5_0),.din(w_dff_A_JsB1D3RH3_0),.clk(gclk));
	jdff dff_A_NrcsKszJ3_0(.dout(w_dff_A_JsB1D3RH3_0),.din(w_dff_A_NrcsKszJ3_0),.clk(gclk));
	jdff dff_A_gF0cEuQl2_0(.dout(w_dff_A_NrcsKszJ3_0),.din(w_dff_A_gF0cEuQl2_0),.clk(gclk));
	jdff dff_A_CxkqJPHN1_0(.dout(w_dff_A_gF0cEuQl2_0),.din(w_dff_A_CxkqJPHN1_0),.clk(gclk));
	jdff dff_A_j9H4W8fS4_0(.dout(w_dff_A_CxkqJPHN1_0),.din(w_dff_A_j9H4W8fS4_0),.clk(gclk));
	jdff dff_A_vfGtvVCT7_0(.dout(w_G204gat_0[0]),.din(w_dff_A_vfGtvVCT7_0),.clk(gclk));
	jdff dff_A_5iniG0Kh2_0(.dout(w_dff_A_vfGtvVCT7_0),.din(w_dff_A_5iniG0Kh2_0),.clk(gclk));
	jdff dff_A_tW67o2ko8_0(.dout(w_dff_A_5iniG0Kh2_0),.din(w_dff_A_tW67o2ko8_0),.clk(gclk));
	jdff dff_A_YI8ihUHD9_0(.dout(w_dff_A_tW67o2ko8_0),.din(w_dff_A_YI8ihUHD9_0),.clk(gclk));
	jdff dff_A_2f3bqegi4_0(.dout(w_dff_A_YI8ihUHD9_0),.din(w_dff_A_2f3bqegi4_0),.clk(gclk));
	jdff dff_A_eBanHSkz1_0(.dout(w_dff_A_2f3bqegi4_0),.din(w_dff_A_eBanHSkz1_0),.clk(gclk));
	jdff dff_A_jc5aLY4O8_0(.dout(w_dff_A_eBanHSkz1_0),.din(w_dff_A_jc5aLY4O8_0),.clk(gclk));
	jdff dff_A_2rokQqMN5_0(.dout(w_dff_A_jc5aLY4O8_0),.din(w_dff_A_2rokQqMN5_0),.clk(gclk));
	jdff dff_A_Gw2FmiMh0_0(.dout(w_dff_A_2rokQqMN5_0),.din(w_dff_A_Gw2FmiMh0_0),.clk(gclk));
	jdff dff_A_3D0cCzIt9_0(.dout(w_G176gat_0[0]),.din(w_dff_A_3D0cCzIt9_0),.clk(gclk));
	jdff dff_A_BhFxGBCj9_0(.dout(w_dff_A_3D0cCzIt9_0),.din(w_dff_A_BhFxGBCj9_0),.clk(gclk));
	jdff dff_A_HMn7Fy4c6_0(.dout(w_dff_A_BhFxGBCj9_0),.din(w_dff_A_HMn7Fy4c6_0),.clk(gclk));
	jdff dff_A_slSttrwN2_0(.dout(w_dff_A_HMn7Fy4c6_0),.din(w_dff_A_slSttrwN2_0),.clk(gclk));
	jdff dff_A_R1Hjm5YU9_0(.dout(w_dff_A_slSttrwN2_0),.din(w_dff_A_R1Hjm5YU9_0),.clk(gclk));
	jdff dff_A_wUu2E1Tg6_0(.dout(w_dff_A_R1Hjm5YU9_0),.din(w_dff_A_wUu2E1Tg6_0),.clk(gclk));
	jdff dff_A_RbKkd4CZ7_0(.dout(w_dff_A_wUu2E1Tg6_0),.din(w_dff_A_RbKkd4CZ7_0),.clk(gclk));
	jdff dff_A_JGf72LPl7_0(.dout(w_dff_A_RbKkd4CZ7_0),.din(w_dff_A_JGf72LPl7_0),.clk(gclk));
	jdff dff_A_IWKs33zr3_0(.dout(w_dff_A_JGf72LPl7_0),.din(w_dff_A_IWKs33zr3_0),.clk(gclk));
	jdff dff_A_bHvBKiqW2_0(.dout(w_G64gat_0[0]),.din(w_dff_A_bHvBKiqW2_0),.clk(gclk));
	jdff dff_A_vOk5WkIj4_0(.dout(w_dff_A_bHvBKiqW2_0),.din(w_dff_A_vOk5WkIj4_0),.clk(gclk));
	jdff dff_A_BQ855u9F3_0(.dout(w_dff_A_vOk5WkIj4_0),.din(w_dff_A_BQ855u9F3_0),.clk(gclk));
	jdff dff_A_Nq4r9eQU4_0(.dout(w_dff_A_BQ855u9F3_0),.din(w_dff_A_Nq4r9eQU4_0),.clk(gclk));
	jdff dff_A_F8juxuHs6_0(.dout(w_dff_A_Nq4r9eQU4_0),.din(w_dff_A_F8juxuHs6_0),.clk(gclk));
	jdff dff_A_7CJVnmPL8_0(.dout(w_dff_A_F8juxuHs6_0),.din(w_dff_A_7CJVnmPL8_0),.clk(gclk));
	jdff dff_A_LgLOrG210_0(.dout(w_dff_A_7CJVnmPL8_0),.din(w_dff_A_LgLOrG210_0),.clk(gclk));
	jdff dff_A_jQITJNMj2_0(.dout(w_dff_A_LgLOrG210_0),.din(w_dff_A_jQITJNMj2_0),.clk(gclk));
	jdff dff_A_O0xEvHZB4_0(.dout(w_dff_A_jQITJNMj2_0),.din(w_dff_A_O0xEvHZB4_0),.clk(gclk));
	jdff dff_A_YWECeiuH1_0(.dout(w_G57gat_0[0]),.din(w_dff_A_YWECeiuH1_0),.clk(gclk));
	jdff dff_A_K8ht5ClC1_0(.dout(w_dff_A_YWECeiuH1_0),.din(w_dff_A_K8ht5ClC1_0),.clk(gclk));
	jdff dff_A_APuOohiE9_0(.dout(w_dff_A_K8ht5ClC1_0),.din(w_dff_A_APuOohiE9_0),.clk(gclk));
	jdff dff_A_qsbhR7XD2_0(.dout(w_dff_A_APuOohiE9_0),.din(w_dff_A_qsbhR7XD2_0),.clk(gclk));
	jdff dff_A_hJCevG5D6_0(.dout(w_dff_A_qsbhR7XD2_0),.din(w_dff_A_hJCevG5D6_0),.clk(gclk));
	jdff dff_A_wfJVwl017_0(.dout(w_dff_A_hJCevG5D6_0),.din(w_dff_A_wfJVwl017_0),.clk(gclk));
	jdff dff_A_CAd6zvoO0_0(.dout(w_dff_A_wfJVwl017_0),.din(w_dff_A_CAd6zvoO0_0),.clk(gclk));
	jdff dff_A_P3d78dXh2_0(.dout(w_dff_A_CAd6zvoO0_0),.din(w_dff_A_P3d78dXh2_0),.clk(gclk));
	jdff dff_A_vUEa1tOP9_0(.dout(w_dff_A_P3d78dXh2_0),.din(w_dff_A_vUEa1tOP9_0),.clk(gclk));
	jdff dff_A_JRmpj3vW1_0(.dout(w_G78gat_0[0]),.din(w_dff_A_JRmpj3vW1_0),.clk(gclk));
	jdff dff_A_mIkq9KWc7_0(.dout(w_dff_A_JRmpj3vW1_0),.din(w_dff_A_mIkq9KWc7_0),.clk(gclk));
	jdff dff_A_kVgO0sV91_0(.dout(w_dff_A_mIkq9KWc7_0),.din(w_dff_A_kVgO0sV91_0),.clk(gclk));
	jdff dff_A_ivwwygLT0_0(.dout(w_dff_A_kVgO0sV91_0),.din(w_dff_A_ivwwygLT0_0),.clk(gclk));
	jdff dff_A_tnoy1bpI3_0(.dout(w_dff_A_ivwwygLT0_0),.din(w_dff_A_tnoy1bpI3_0),.clk(gclk));
	jdff dff_A_xl3vBmQY7_0(.dout(w_dff_A_tnoy1bpI3_0),.din(w_dff_A_xl3vBmQY7_0),.clk(gclk));
	jdff dff_A_lw9uu5et0_0(.dout(w_dff_A_xl3vBmQY7_0),.din(w_dff_A_lw9uu5et0_0),.clk(gclk));
	jdff dff_A_ApUu8QX68_0(.dout(w_dff_A_lw9uu5et0_0),.din(w_dff_A_ApUu8QX68_0),.clk(gclk));
	jdff dff_A_SyaQvzUr9_0(.dout(w_dff_A_ApUu8QX68_0),.din(w_dff_A_SyaQvzUr9_0),.clk(gclk));
	jdff dff_A_wqM4bRK39_0(.dout(w_G71gat_0[0]),.din(w_dff_A_wqM4bRK39_0),.clk(gclk));
	jdff dff_A_hmxSCtab0_0(.dout(w_dff_A_wqM4bRK39_0),.din(w_dff_A_hmxSCtab0_0),.clk(gclk));
	jdff dff_A_IiVfJ6Lt3_0(.dout(w_dff_A_hmxSCtab0_0),.din(w_dff_A_IiVfJ6Lt3_0),.clk(gclk));
	jdff dff_A_dEnjAOzf4_0(.dout(w_dff_A_IiVfJ6Lt3_0),.din(w_dff_A_dEnjAOzf4_0),.clk(gclk));
	jdff dff_A_SMsC3kwI7_0(.dout(w_dff_A_dEnjAOzf4_0),.din(w_dff_A_SMsC3kwI7_0),.clk(gclk));
	jdff dff_A_JpiXpZXw7_0(.dout(w_dff_A_SMsC3kwI7_0),.din(w_dff_A_JpiXpZXw7_0),.clk(gclk));
	jdff dff_A_Q9tQXbC02_0(.dout(w_dff_A_JpiXpZXw7_0),.din(w_dff_A_Q9tQXbC02_0),.clk(gclk));
	jdff dff_A_MrFTOFe00_0(.dout(w_dff_A_Q9tQXbC02_0),.din(w_dff_A_MrFTOFe00_0),.clk(gclk));
	jdff dff_A_bH14foRf7_0(.dout(w_dff_A_MrFTOFe00_0),.din(w_dff_A_bH14foRf7_0),.clk(gclk));
	jdff dff_A_SS3Vkgin2_0(.dout(w_G141gat_0[0]),.din(w_dff_A_SS3Vkgin2_0),.clk(gclk));
	jdff dff_A_lLV4X3S78_0(.dout(w_dff_A_SS3Vkgin2_0),.din(w_dff_A_lLV4X3S78_0),.clk(gclk));
	jdff dff_A_ErAp9cSi4_0(.dout(w_dff_A_lLV4X3S78_0),.din(w_dff_A_ErAp9cSi4_0),.clk(gclk));
	jdff dff_A_KDP32BWO9_0(.dout(w_dff_A_ErAp9cSi4_0),.din(w_dff_A_KDP32BWO9_0),.clk(gclk));
	jdff dff_A_V7QMWGL00_0(.dout(w_dff_A_KDP32BWO9_0),.din(w_dff_A_V7QMWGL00_0),.clk(gclk));
	jdff dff_A_uNJqB8J02_0(.dout(w_dff_A_V7QMWGL00_0),.din(w_dff_A_uNJqB8J02_0),.clk(gclk));
	jdff dff_A_b8JYYJic6_0(.dout(w_dff_A_uNJqB8J02_0),.din(w_dff_A_b8JYYJic6_0),.clk(gclk));
	jdff dff_A_rmSHLCRY7_0(.dout(w_dff_A_b8JYYJic6_0),.din(w_dff_A_rmSHLCRY7_0),.clk(gclk));
	jdff dff_A_i5rz0XZO0_0(.dout(w_dff_A_rmSHLCRY7_0),.din(w_dff_A_i5rz0XZO0_0),.clk(gclk));
	jdff dff_A_5xvVeZUQ1_0(.dout(w_G113gat_0[0]),.din(w_dff_A_5xvVeZUQ1_0),.clk(gclk));
	jdff dff_A_L926TgT70_0(.dout(w_dff_A_5xvVeZUQ1_0),.din(w_dff_A_L926TgT70_0),.clk(gclk));
	jdff dff_A_uGDL3LlH8_0(.dout(w_dff_A_L926TgT70_0),.din(w_dff_A_uGDL3LlH8_0),.clk(gclk));
	jdff dff_A_LQnVihV25_0(.dout(w_dff_A_uGDL3LlH8_0),.din(w_dff_A_LQnVihV25_0),.clk(gclk));
	jdff dff_A_LARyHFiL2_0(.dout(w_dff_A_LQnVihV25_0),.din(w_dff_A_LARyHFiL2_0),.clk(gclk));
	jdff dff_A_y93UQyjQ9_0(.dout(w_dff_A_LARyHFiL2_0),.din(w_dff_A_y93UQyjQ9_0),.clk(gclk));
	jdff dff_A_mgdO3aCs5_0(.dout(w_dff_A_y93UQyjQ9_0),.din(w_dff_A_mgdO3aCs5_0),.clk(gclk));
	jdff dff_A_Cds15KqZ2_0(.dout(w_dff_A_mgdO3aCs5_0),.din(w_dff_A_Cds15KqZ2_0),.clk(gclk));
	jdff dff_A_RJtrtdK02_0(.dout(w_dff_A_Cds15KqZ2_0),.din(w_dff_A_RJtrtdK02_0),.clk(gclk));
	jdff dff_A_8cZgt6PL3_0(.dout(w_G197gat_0[0]),.din(w_dff_A_8cZgt6PL3_0),.clk(gclk));
	jdff dff_A_gyWsRh5u5_0(.dout(w_dff_A_8cZgt6PL3_0),.din(w_dff_A_gyWsRh5u5_0),.clk(gclk));
	jdff dff_A_cP7XeylB5_0(.dout(w_dff_A_gyWsRh5u5_0),.din(w_dff_A_cP7XeylB5_0),.clk(gclk));
	jdff dff_A_WKBsu2kb7_0(.dout(w_dff_A_cP7XeylB5_0),.din(w_dff_A_WKBsu2kb7_0),.clk(gclk));
	jdff dff_A_yk7MLahK2_0(.dout(w_dff_A_WKBsu2kb7_0),.din(w_dff_A_yk7MLahK2_0),.clk(gclk));
	jdff dff_A_6IjGjCaJ9_0(.dout(w_dff_A_yk7MLahK2_0),.din(w_dff_A_6IjGjCaJ9_0),.clk(gclk));
	jdff dff_A_aBYOTLyX7_0(.dout(w_dff_A_6IjGjCaJ9_0),.din(w_dff_A_aBYOTLyX7_0),.clk(gclk));
	jdff dff_A_xQl0VRP72_0(.dout(w_dff_A_aBYOTLyX7_0),.din(w_dff_A_xQl0VRP72_0),.clk(gclk));
	jdff dff_A_DgsZDsXk0_0(.dout(w_dff_A_xQl0VRP72_0),.din(w_dff_A_DgsZDsXk0_0),.clk(gclk));
	jdff dff_A_8tqHFnHw5_0(.dout(w_G169gat_0[0]),.din(w_dff_A_8tqHFnHw5_0),.clk(gclk));
	jdff dff_A_gA4zrwt49_0(.dout(w_dff_A_8tqHFnHw5_0),.din(w_dff_A_gA4zrwt49_0),.clk(gclk));
	jdff dff_A_0geqOlnf9_0(.dout(w_dff_A_gA4zrwt49_0),.din(w_dff_A_0geqOlnf9_0),.clk(gclk));
	jdff dff_A_OTtH03OS3_0(.dout(w_dff_A_0geqOlnf9_0),.din(w_dff_A_OTtH03OS3_0),.clk(gclk));
	jdff dff_A_7rsDzaEd8_0(.dout(w_dff_A_OTtH03OS3_0),.din(w_dff_A_7rsDzaEd8_0),.clk(gclk));
	jdff dff_A_8msweTtN0_0(.dout(w_dff_A_7rsDzaEd8_0),.din(w_dff_A_8msweTtN0_0),.clk(gclk));
	jdff dff_A_P6twqtTa7_0(.dout(w_dff_A_8msweTtN0_0),.din(w_dff_A_P6twqtTa7_0),.clk(gclk));
	jdff dff_A_HZ4p6TmS2_0(.dout(w_dff_A_P6twqtTa7_0),.din(w_dff_A_HZ4p6TmS2_0),.clk(gclk));
	jdff dff_A_fdC9aunC4_0(.dout(w_dff_A_HZ4p6TmS2_0),.din(w_dff_A_fdC9aunC4_0),.clk(gclk));
	jdff dff_A_qxa5TtMk0_0(.dout(w_G8gat_0[0]),.din(w_dff_A_qxa5TtMk0_0),.clk(gclk));
	jdff dff_A_V76aXWiQ6_0(.dout(w_dff_A_qxa5TtMk0_0),.din(w_dff_A_V76aXWiQ6_0),.clk(gclk));
	jdff dff_A_WRnJI9Kl9_0(.dout(w_dff_A_V76aXWiQ6_0),.din(w_dff_A_WRnJI9Kl9_0),.clk(gclk));
	jdff dff_A_kDVMhmEy5_0(.dout(w_dff_A_WRnJI9Kl9_0),.din(w_dff_A_kDVMhmEy5_0),.clk(gclk));
	jdff dff_A_BvkTwHL13_0(.dout(w_dff_A_kDVMhmEy5_0),.din(w_dff_A_BvkTwHL13_0),.clk(gclk));
	jdff dff_A_7I6nZD8M5_0(.dout(w_dff_A_BvkTwHL13_0),.din(w_dff_A_7I6nZD8M5_0),.clk(gclk));
	jdff dff_A_jzEg5pm64_0(.dout(w_dff_A_7I6nZD8M5_0),.din(w_dff_A_jzEg5pm64_0),.clk(gclk));
	jdff dff_A_nCG7rUg54_0(.dout(w_dff_A_jzEg5pm64_0),.din(w_dff_A_nCG7rUg54_0),.clk(gclk));
	jdff dff_A_gBnaavUD6_0(.dout(w_dff_A_nCG7rUg54_0),.din(w_dff_A_gBnaavUD6_0),.clk(gclk));
	jdff dff_A_d6pMsqyY1_0(.dout(w_G1gat_0[0]),.din(w_dff_A_d6pMsqyY1_0),.clk(gclk));
	jdff dff_A_8XMPAys19_0(.dout(w_dff_A_d6pMsqyY1_0),.din(w_dff_A_8XMPAys19_0),.clk(gclk));
	jdff dff_A_YZJZwMlC4_0(.dout(w_dff_A_8XMPAys19_0),.din(w_dff_A_YZJZwMlC4_0),.clk(gclk));
	jdff dff_A_cMuuJ3HN3_0(.dout(w_dff_A_YZJZwMlC4_0),.din(w_dff_A_cMuuJ3HN3_0),.clk(gclk));
	jdff dff_A_YsrSFMqX9_0(.dout(w_dff_A_cMuuJ3HN3_0),.din(w_dff_A_YsrSFMqX9_0),.clk(gclk));
	jdff dff_A_aqUX2jBo3_0(.dout(w_dff_A_YsrSFMqX9_0),.din(w_dff_A_aqUX2jBo3_0),.clk(gclk));
	jdff dff_A_hQ7lpytX3_0(.dout(w_dff_A_aqUX2jBo3_0),.din(w_dff_A_hQ7lpytX3_0),.clk(gclk));
	jdff dff_A_3lu6ZQS50_0(.dout(w_dff_A_hQ7lpytX3_0),.din(w_dff_A_3lu6ZQS50_0),.clk(gclk));
	jdff dff_A_R1Kk3biT2_0(.dout(w_dff_A_3lu6ZQS50_0),.din(w_dff_A_R1Kk3biT2_0),.clk(gclk));
	jdff dff_A_z94p2JxK8_0(.dout(w_G22gat_0[0]),.din(w_dff_A_z94p2JxK8_0),.clk(gclk));
	jdff dff_A_6WvV3fa74_0(.dout(w_dff_A_z94p2JxK8_0),.din(w_dff_A_6WvV3fa74_0),.clk(gclk));
	jdff dff_A_eYngrMjt2_0(.dout(w_dff_A_6WvV3fa74_0),.din(w_dff_A_eYngrMjt2_0),.clk(gclk));
	jdff dff_A_7P5UDB3E3_0(.dout(w_dff_A_eYngrMjt2_0),.din(w_dff_A_7P5UDB3E3_0),.clk(gclk));
	jdff dff_A_8uX3ycbG4_0(.dout(w_dff_A_7P5UDB3E3_0),.din(w_dff_A_8uX3ycbG4_0),.clk(gclk));
	jdff dff_A_EGVbRc0F9_0(.dout(w_dff_A_8uX3ycbG4_0),.din(w_dff_A_EGVbRc0F9_0),.clk(gclk));
	jdff dff_A_iDYW34Zv8_0(.dout(w_dff_A_EGVbRc0F9_0),.din(w_dff_A_iDYW34Zv8_0),.clk(gclk));
	jdff dff_A_FqZZi1YR1_0(.dout(w_dff_A_iDYW34Zv8_0),.din(w_dff_A_FqZZi1YR1_0),.clk(gclk));
	jdff dff_A_stWt3Lte9_0(.dout(w_dff_A_FqZZi1YR1_0),.din(w_dff_A_stWt3Lte9_0),.clk(gclk));
	jdff dff_A_IqyTzLwR5_0(.dout(w_G15gat_0[0]),.din(w_dff_A_IqyTzLwR5_0),.clk(gclk));
	jdff dff_A_845PcrZY6_0(.dout(w_dff_A_IqyTzLwR5_0),.din(w_dff_A_845PcrZY6_0),.clk(gclk));
	jdff dff_A_eWXkWq271_0(.dout(w_dff_A_845PcrZY6_0),.din(w_dff_A_eWXkWq271_0),.clk(gclk));
	jdff dff_A_KYjcePUD0_0(.dout(w_dff_A_eWXkWq271_0),.din(w_dff_A_KYjcePUD0_0),.clk(gclk));
	jdff dff_A_izVBTHt02_0(.dout(w_dff_A_KYjcePUD0_0),.din(w_dff_A_izVBTHt02_0),.clk(gclk));
	jdff dff_A_cKHFlPhF7_0(.dout(w_dff_A_izVBTHt02_0),.din(w_dff_A_cKHFlPhF7_0),.clk(gclk));
	jdff dff_A_Ppkqod837_0(.dout(w_dff_A_cKHFlPhF7_0),.din(w_dff_A_Ppkqod837_0),.clk(gclk));
	jdff dff_A_BrXcoD0H4_0(.dout(w_dff_A_Ppkqod837_0),.din(w_dff_A_BrXcoD0H4_0),.clk(gclk));
	jdff dff_A_1aKUPuaX8_0(.dout(w_dff_A_BrXcoD0H4_0),.din(w_dff_A_1aKUPuaX8_0),.clk(gclk));
	jdff dff_A_GWzDKBZD4_1(.dout(w_n193_0[1]),.din(w_dff_A_GWzDKBZD4_1),.clk(gclk));
	jdff dff_A_btjalPWr6_1(.dout(w_dff_A_GWzDKBZD4_1),.din(w_dff_A_btjalPWr6_1),.clk(gclk));
	jdff dff_A_b8y4dfmI3_1(.dout(w_dff_A_btjalPWr6_1),.din(w_dff_A_b8y4dfmI3_1),.clk(gclk));
	jdff dff_A_mXsTGYGu8_1(.dout(w_dff_A_b8y4dfmI3_1),.din(w_dff_A_mXsTGYGu8_1),.clk(gclk));
	jdff dff_A_lNEaeZEi6_2(.dout(w_n193_0[2]),.din(w_dff_A_lNEaeZEi6_2),.clk(gclk));
	jdff dff_A_xzS7HUuI9_2(.dout(w_dff_A_lNEaeZEi6_2),.din(w_dff_A_xzS7HUuI9_2),.clk(gclk));
	jdff dff_A_3yfnbr4L1_2(.dout(w_dff_A_xzS7HUuI9_2),.din(w_dff_A_3yfnbr4L1_2),.clk(gclk));
	jdff dff_A_zHWUR9p43_2(.dout(w_dff_A_3yfnbr4L1_2),.din(w_dff_A_zHWUR9p43_2),.clk(gclk));
	jdff dff_A_ibsX1cxs4_0(.dout(w_G162gat_0[0]),.din(w_dff_A_ibsX1cxs4_0),.clk(gclk));
	jdff dff_A_tCdREcKa2_0(.dout(w_dff_A_ibsX1cxs4_0),.din(w_dff_A_tCdREcKa2_0),.clk(gclk));
	jdff dff_A_vFNQZEMZ1_0(.dout(w_dff_A_tCdREcKa2_0),.din(w_dff_A_vFNQZEMZ1_0),.clk(gclk));
	jdff dff_A_iUmeuBPm1_0(.dout(w_dff_A_vFNQZEMZ1_0),.din(w_dff_A_iUmeuBPm1_0),.clk(gclk));
	jdff dff_A_PzxzdSoV4_0(.dout(w_dff_A_iUmeuBPm1_0),.din(w_dff_A_PzxzdSoV4_0),.clk(gclk));
	jdff dff_A_rjqeuLkK5_0(.dout(w_dff_A_PzxzdSoV4_0),.din(w_dff_A_rjqeuLkK5_0),.clk(gclk));
	jdff dff_A_jUz51r6j8_0(.dout(w_dff_A_rjqeuLkK5_0),.din(w_dff_A_jUz51r6j8_0),.clk(gclk));
	jdff dff_A_Box9InxF9_0(.dout(w_dff_A_jUz51r6j8_0),.din(w_dff_A_Box9InxF9_0),.clk(gclk));
	jdff dff_A_rAX5N1mb8_0(.dout(w_dff_A_Box9InxF9_0),.din(w_dff_A_rAX5N1mb8_0),.clk(gclk));
	jdff dff_A_3BfG94Lu2_0(.dout(w_G134gat_0[0]),.din(w_dff_A_3BfG94Lu2_0),.clk(gclk));
	jdff dff_A_eHZZYIL78_0(.dout(w_dff_A_3BfG94Lu2_0),.din(w_dff_A_eHZZYIL78_0),.clk(gclk));
	jdff dff_A_uBxlZuto1_0(.dout(w_dff_A_eHZZYIL78_0),.din(w_dff_A_uBxlZuto1_0),.clk(gclk));
	jdff dff_A_jAx6sNoT5_0(.dout(w_dff_A_uBxlZuto1_0),.din(w_dff_A_jAx6sNoT5_0),.clk(gclk));
	jdff dff_A_rMxDDKKr1_0(.dout(w_dff_A_jAx6sNoT5_0),.din(w_dff_A_rMxDDKKr1_0),.clk(gclk));
	jdff dff_A_vUssrorw4_0(.dout(w_dff_A_rMxDDKKr1_0),.din(w_dff_A_vUssrorw4_0),.clk(gclk));
	jdff dff_A_sgcqp6yk5_0(.dout(w_dff_A_vUssrorw4_0),.din(w_dff_A_sgcqp6yk5_0),.clk(gclk));
	jdff dff_A_bh1PU6yV7_0(.dout(w_dff_A_sgcqp6yk5_0),.din(w_dff_A_bh1PU6yV7_0),.clk(gclk));
	jdff dff_A_R0VlCnVr4_0(.dout(w_dff_A_bh1PU6yV7_0),.din(w_dff_A_R0VlCnVr4_0),.clk(gclk));
	jdff dff_A_nh98z9qp3_0(.dout(w_G218gat_0[0]),.din(w_dff_A_nh98z9qp3_0),.clk(gclk));
	jdff dff_A_38qDdbeF7_0(.dout(w_dff_A_nh98z9qp3_0),.din(w_dff_A_38qDdbeF7_0),.clk(gclk));
	jdff dff_A_AVpyYFh75_0(.dout(w_dff_A_38qDdbeF7_0),.din(w_dff_A_AVpyYFh75_0),.clk(gclk));
	jdff dff_A_ODtt1Elw8_0(.dout(w_dff_A_AVpyYFh75_0),.din(w_dff_A_ODtt1Elw8_0),.clk(gclk));
	jdff dff_A_ybj2aDPc2_0(.dout(w_dff_A_ODtt1Elw8_0),.din(w_dff_A_ybj2aDPc2_0),.clk(gclk));
	jdff dff_A_jKvWkiT39_0(.dout(w_dff_A_ybj2aDPc2_0),.din(w_dff_A_jKvWkiT39_0),.clk(gclk));
	jdff dff_A_ui2ARFNK3_0(.dout(w_dff_A_jKvWkiT39_0),.din(w_dff_A_ui2ARFNK3_0),.clk(gclk));
	jdff dff_A_pXC3GHm42_0(.dout(w_dff_A_ui2ARFNK3_0),.din(w_dff_A_pXC3GHm42_0),.clk(gclk));
	jdff dff_A_4ix7yO1c6_0(.dout(w_dff_A_pXC3GHm42_0),.din(w_dff_A_4ix7yO1c6_0),.clk(gclk));
	jdff dff_A_u4DOqvYj9_0(.dout(w_G190gat_0[0]),.din(w_dff_A_u4DOqvYj9_0),.clk(gclk));
	jdff dff_A_mnUv4xHz2_0(.dout(w_dff_A_u4DOqvYj9_0),.din(w_dff_A_mnUv4xHz2_0),.clk(gclk));
	jdff dff_A_Zq7j6Wug3_0(.dout(w_dff_A_mnUv4xHz2_0),.din(w_dff_A_Zq7j6Wug3_0),.clk(gclk));
	jdff dff_A_7kQCIwvX5_0(.dout(w_dff_A_Zq7j6Wug3_0),.din(w_dff_A_7kQCIwvX5_0),.clk(gclk));
	jdff dff_A_cZZvKzC88_0(.dout(w_dff_A_7kQCIwvX5_0),.din(w_dff_A_cZZvKzC88_0),.clk(gclk));
	jdff dff_A_xMa23chv2_0(.dout(w_dff_A_cZZvKzC88_0),.din(w_dff_A_xMa23chv2_0),.clk(gclk));
	jdff dff_A_aLRmqX4y5_0(.dout(w_dff_A_xMa23chv2_0),.din(w_dff_A_aLRmqX4y5_0),.clk(gclk));
	jdff dff_A_0rgyHWSn3_0(.dout(w_dff_A_aLRmqX4y5_0),.din(w_dff_A_0rgyHWSn3_0),.clk(gclk));
	jdff dff_A_7bIcqB0f7_0(.dout(w_dff_A_0rgyHWSn3_0),.din(w_dff_A_7bIcqB0f7_0),.clk(gclk));
	jdff dff_A_HgIZFkTJ4_0(.dout(w_G92gat_0[0]),.din(w_dff_A_HgIZFkTJ4_0),.clk(gclk));
	jdff dff_A_S1zPxHxo4_0(.dout(w_dff_A_HgIZFkTJ4_0),.din(w_dff_A_S1zPxHxo4_0),.clk(gclk));
	jdff dff_A_N5qQfwvz4_0(.dout(w_dff_A_S1zPxHxo4_0),.din(w_dff_A_N5qQfwvz4_0),.clk(gclk));
	jdff dff_A_SbXpIhpg1_0(.dout(w_dff_A_N5qQfwvz4_0),.din(w_dff_A_SbXpIhpg1_0),.clk(gclk));
	jdff dff_A_jARsJAHT1_0(.dout(w_dff_A_SbXpIhpg1_0),.din(w_dff_A_jARsJAHT1_0),.clk(gclk));
	jdff dff_A_8bmxk5ct5_0(.dout(w_dff_A_jARsJAHT1_0),.din(w_dff_A_8bmxk5ct5_0),.clk(gclk));
	jdff dff_A_YLBSHGtv6_0(.dout(w_dff_A_8bmxk5ct5_0),.din(w_dff_A_YLBSHGtv6_0),.clk(gclk));
	jdff dff_A_Wo2KMpZw1_0(.dout(w_dff_A_YLBSHGtv6_0),.din(w_dff_A_Wo2KMpZw1_0),.clk(gclk));
	jdff dff_A_jq8KQ46T1_0(.dout(w_dff_A_Wo2KMpZw1_0),.din(w_dff_A_jq8KQ46T1_0),.clk(gclk));
	jdff dff_A_dcTQargd2_0(.dout(w_G85gat_0[0]),.din(w_dff_A_dcTQargd2_0),.clk(gclk));
	jdff dff_A_41sYUzFO3_0(.dout(w_dff_A_dcTQargd2_0),.din(w_dff_A_41sYUzFO3_0),.clk(gclk));
	jdff dff_A_sJYDNqPR5_0(.dout(w_dff_A_41sYUzFO3_0),.din(w_dff_A_sJYDNqPR5_0),.clk(gclk));
	jdff dff_A_pegcWvZv1_0(.dout(w_dff_A_sJYDNqPR5_0),.din(w_dff_A_pegcWvZv1_0),.clk(gclk));
	jdff dff_A_iweDOZN63_0(.dout(w_dff_A_pegcWvZv1_0),.din(w_dff_A_iweDOZN63_0),.clk(gclk));
	jdff dff_A_laIWXTMB6_0(.dout(w_dff_A_iweDOZN63_0),.din(w_dff_A_laIWXTMB6_0),.clk(gclk));
	jdff dff_A_uiXBeY8o9_0(.dout(w_dff_A_laIWXTMB6_0),.din(w_dff_A_uiXBeY8o9_0),.clk(gclk));
	jdff dff_A_oczNyP5o9_0(.dout(w_dff_A_uiXBeY8o9_0),.din(w_dff_A_oczNyP5o9_0),.clk(gclk));
	jdff dff_A_VwcYzyRB8_0(.dout(w_dff_A_oczNyP5o9_0),.din(w_dff_A_VwcYzyRB8_0),.clk(gclk));
	jdff dff_A_OzhPNIhy0_0(.dout(w_G106gat_0[0]),.din(w_dff_A_OzhPNIhy0_0),.clk(gclk));
	jdff dff_A_2HuVFVWt7_0(.dout(w_dff_A_OzhPNIhy0_0),.din(w_dff_A_2HuVFVWt7_0),.clk(gclk));
	jdff dff_A_KoDAHiOe0_0(.dout(w_dff_A_2HuVFVWt7_0),.din(w_dff_A_KoDAHiOe0_0),.clk(gclk));
	jdff dff_A_JCRifkk40_0(.dout(w_dff_A_KoDAHiOe0_0),.din(w_dff_A_JCRifkk40_0),.clk(gclk));
	jdff dff_A_Uhqsz52h4_0(.dout(w_dff_A_JCRifkk40_0),.din(w_dff_A_Uhqsz52h4_0),.clk(gclk));
	jdff dff_A_cldGPkuk8_0(.dout(w_dff_A_Uhqsz52h4_0),.din(w_dff_A_cldGPkuk8_0),.clk(gclk));
	jdff dff_A_N76rax1t8_0(.dout(w_dff_A_cldGPkuk8_0),.din(w_dff_A_N76rax1t8_0),.clk(gclk));
	jdff dff_A_ik88G5GF9_0(.dout(w_dff_A_N76rax1t8_0),.din(w_dff_A_ik88G5GF9_0),.clk(gclk));
	jdff dff_A_LGoqKOvX1_0(.dout(w_dff_A_ik88G5GF9_0),.din(w_dff_A_LGoqKOvX1_0),.clk(gclk));
	jdff dff_A_hjYQRhIH2_0(.dout(w_G99gat_0[0]),.din(w_dff_A_hjYQRhIH2_0),.clk(gclk));
	jdff dff_A_tNw4S6Df5_0(.dout(w_dff_A_hjYQRhIH2_0),.din(w_dff_A_tNw4S6Df5_0),.clk(gclk));
	jdff dff_A_FFLW49A00_0(.dout(w_dff_A_tNw4S6Df5_0),.din(w_dff_A_FFLW49A00_0),.clk(gclk));
	jdff dff_A_jsZlvTon1_0(.dout(w_dff_A_FFLW49A00_0),.din(w_dff_A_jsZlvTon1_0),.clk(gclk));
	jdff dff_A_j6uKOymn5_0(.dout(w_dff_A_jsZlvTon1_0),.din(w_dff_A_j6uKOymn5_0),.clk(gclk));
	jdff dff_A_rAMLe7Y78_0(.dout(w_dff_A_j6uKOymn5_0),.din(w_dff_A_rAMLe7Y78_0),.clk(gclk));
	jdff dff_A_eFPGJfq35_0(.dout(w_dff_A_rAMLe7Y78_0),.din(w_dff_A_eFPGJfq35_0),.clk(gclk));
	jdff dff_A_1rgRVts25_0(.dout(w_dff_A_eFPGJfq35_0),.din(w_dff_A_1rgRVts25_0),.clk(gclk));
	jdff dff_A_jpqv8m5G6_0(.dout(w_dff_A_1rgRVts25_0),.din(w_dff_A_jpqv8m5G6_0),.clk(gclk));
	jdff dff_B_lGXLKP903_0(.din(n191),.dout(w_dff_B_lGXLKP903_0),.clk(gclk));
	jdff dff_A_cHovN6V07_0(.dout(w_G36gat_0[0]),.din(w_dff_A_cHovN6V07_0),.clk(gclk));
	jdff dff_A_bLhCn3Y76_0(.dout(w_dff_A_cHovN6V07_0),.din(w_dff_A_bLhCn3Y76_0),.clk(gclk));
	jdff dff_A_mBEEZ1aI1_0(.dout(w_dff_A_bLhCn3Y76_0),.din(w_dff_A_mBEEZ1aI1_0),.clk(gclk));
	jdff dff_A_3jdHesJ14_0(.dout(w_dff_A_mBEEZ1aI1_0),.din(w_dff_A_3jdHesJ14_0),.clk(gclk));
	jdff dff_A_6PHoglSS2_0(.dout(w_dff_A_3jdHesJ14_0),.din(w_dff_A_6PHoglSS2_0),.clk(gclk));
	jdff dff_A_7DELWPFL7_0(.dout(w_dff_A_6PHoglSS2_0),.din(w_dff_A_7DELWPFL7_0),.clk(gclk));
	jdff dff_A_lP662Jqj8_0(.dout(w_dff_A_7DELWPFL7_0),.din(w_dff_A_lP662Jqj8_0),.clk(gclk));
	jdff dff_A_ZMWiXPVM8_0(.dout(w_dff_A_lP662Jqj8_0),.din(w_dff_A_ZMWiXPVM8_0),.clk(gclk));
	jdff dff_A_v7ED5tYc9_0(.dout(w_dff_A_ZMWiXPVM8_0),.din(w_dff_A_v7ED5tYc9_0),.clk(gclk));
	jdff dff_A_VwB4v1RI5_0(.dout(w_G29gat_0[0]),.din(w_dff_A_VwB4v1RI5_0),.clk(gclk));
	jdff dff_A_LaQyHxma8_0(.dout(w_dff_A_VwB4v1RI5_0),.din(w_dff_A_LaQyHxma8_0),.clk(gclk));
	jdff dff_A_I3KZClPs6_0(.dout(w_dff_A_LaQyHxma8_0),.din(w_dff_A_I3KZClPs6_0),.clk(gclk));
	jdff dff_A_ht4nWXRa4_0(.dout(w_dff_A_I3KZClPs6_0),.din(w_dff_A_ht4nWXRa4_0),.clk(gclk));
	jdff dff_A_FOQxKWTa0_0(.dout(w_dff_A_ht4nWXRa4_0),.din(w_dff_A_FOQxKWTa0_0),.clk(gclk));
	jdff dff_A_CbVdveOh1_0(.dout(w_dff_A_FOQxKWTa0_0),.din(w_dff_A_CbVdveOh1_0),.clk(gclk));
	jdff dff_A_Kz7moYql1_0(.dout(w_dff_A_CbVdveOh1_0),.din(w_dff_A_Kz7moYql1_0),.clk(gclk));
	jdff dff_A_50J4jW6q2_0(.dout(w_dff_A_Kz7moYql1_0),.din(w_dff_A_50J4jW6q2_0),.clk(gclk));
	jdff dff_A_SDqRMGgO8_0(.dout(w_dff_A_50J4jW6q2_0),.din(w_dff_A_SDqRMGgO8_0),.clk(gclk));
	jdff dff_A_x3xM2y5l7_0(.dout(w_G50gat_0[0]),.din(w_dff_A_x3xM2y5l7_0),.clk(gclk));
	jdff dff_A_RGLLuGf07_0(.dout(w_dff_A_x3xM2y5l7_0),.din(w_dff_A_RGLLuGf07_0),.clk(gclk));
	jdff dff_A_baFEwu9S7_0(.dout(w_dff_A_RGLLuGf07_0),.din(w_dff_A_baFEwu9S7_0),.clk(gclk));
	jdff dff_A_A8XbdSah2_0(.dout(w_dff_A_baFEwu9S7_0),.din(w_dff_A_A8XbdSah2_0),.clk(gclk));
	jdff dff_A_n2qcSHdG9_0(.dout(w_dff_A_A8XbdSah2_0),.din(w_dff_A_n2qcSHdG9_0),.clk(gclk));
	jdff dff_A_apya2kGJ1_0(.dout(w_dff_A_n2qcSHdG9_0),.din(w_dff_A_apya2kGJ1_0),.clk(gclk));
	jdff dff_A_qnaUJiEI2_0(.dout(w_dff_A_apya2kGJ1_0),.din(w_dff_A_qnaUJiEI2_0),.clk(gclk));
	jdff dff_A_eD3q2sz12_0(.dout(w_dff_A_qnaUJiEI2_0),.din(w_dff_A_eD3q2sz12_0),.clk(gclk));
	jdff dff_A_jrgtPD7H9_0(.dout(w_dff_A_eD3q2sz12_0),.din(w_dff_A_jrgtPD7H9_0),.clk(gclk));
	jdff dff_A_3pmWagUy8_0(.dout(w_G43gat_0[0]),.din(w_dff_A_3pmWagUy8_0),.clk(gclk));
	jdff dff_A_v7PwXPi94_0(.dout(w_dff_A_3pmWagUy8_0),.din(w_dff_A_v7PwXPi94_0),.clk(gclk));
	jdff dff_A_cPhaBPVu6_0(.dout(w_dff_A_v7PwXPi94_0),.din(w_dff_A_cPhaBPVu6_0),.clk(gclk));
	jdff dff_A_hxFmtyc21_0(.dout(w_dff_A_cPhaBPVu6_0),.din(w_dff_A_hxFmtyc21_0),.clk(gclk));
	jdff dff_A_nc7ErHap5_0(.dout(w_dff_A_hxFmtyc21_0),.din(w_dff_A_nc7ErHap5_0),.clk(gclk));
	jdff dff_A_oKgMuC9Y5_0(.dout(w_dff_A_nc7ErHap5_0),.din(w_dff_A_oKgMuC9Y5_0),.clk(gclk));
	jdff dff_A_UBXeWElZ8_0(.dout(w_dff_A_oKgMuC9Y5_0),.din(w_dff_A_UBXeWElZ8_0),.clk(gclk));
	jdff dff_A_7UIp3iqL5_0(.dout(w_dff_A_UBXeWElZ8_0),.din(w_dff_A_7UIp3iqL5_0),.clk(gclk));
	jdff dff_A_EHOuqmax2_0(.dout(w_dff_A_7UIp3iqL5_0),.din(w_dff_A_EHOuqmax2_0),.clk(gclk));
endmodule

