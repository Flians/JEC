/*
gf_c5315:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jdff: 6080
	jand: 606
	jor: 486

Summary:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jdff: 6080
	jand: 606
	jor: 486

The maximum logic level gap of any gate:
	gf_c5315: 22
*/

module gf_c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [1:0] w_G1_2;
	wire [2:0] w_G4_0;
	wire [1:0] w_G11_0;
	wire [1:0] w_G14_0;
	wire [1:0] w_G17_0;
	wire [1:0] w_G20_0;
	wire [1:0] w_G37_0;
	wire [1:0] w_G40_0;
	wire [1:0] w_G43_0;
	wire [1:0] w_G46_0;
	wire [1:0] w_G49_0;
	wire [2:0] w_G54_0;
	wire [1:0] w_G61_0;
	wire [1:0] w_G64_0;
	wire [1:0] w_G67_0;
	wire [1:0] w_G70_0;
	wire [1:0] w_G73_0;
	wire [1:0] w_G76_0;
	wire [1:0] w_G91_0;
	wire [1:0] w_G100_0;
	wire [1:0] w_G103_0;
	wire [1:0] w_G106_0;
	wire [1:0] w_G109_0;
	wire [1:0] w_G123_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G137_2;
	wire [2:0] w_G137_3;
	wire [2:0] w_G137_4;
	wire [2:0] w_G137_5;
	wire [2:0] w_G137_6;
	wire [2:0] w_G137_7;
	wire [2:0] w_G137_8;
	wire [1:0] w_G137_9;
	wire [2:0] w_G141_0;
	wire [2:0] w_G141_1;
	wire [2:0] w_G141_2;
	wire [1:0] w_G146_0;
	wire [1:0] w_G149_0;
	wire [1:0] w_G152_0;
	wire [1:0] w_G155_0;
	wire [1:0] w_G158_0;
	wire [1:0] w_G161_0;
	wire [1:0] w_G164_0;
	wire [1:0] w_G167_0;
	wire [1:0] w_G170_0;
	wire [1:0] w_G173_0;
	wire [1:0] w_G182_0;
	wire [1:0] w_G185_0;
	wire [1:0] w_G188_0;
	wire [1:0] w_G191_0;
	wire [1:0] w_G194_0;
	wire [1:0] w_G197_0;
	wire [1:0] w_G200_0;
	wire [1:0] w_G203_0;
	wire [2:0] w_G206_0;
	wire [2:0] w_G206_1;
	wire [2:0] w_G210_0;
	wire [2:0] w_G210_1;
	wire [1:0] w_G210_2;
	wire [2:0] w_G218_0;
	wire [2:0] w_G218_1;
	wire [1:0] w_G218_2;
	wire [2:0] w_G226_0;
	wire [2:0] w_G226_1;
	wire [1:0] w_G226_2;
	wire [2:0] w_G234_0;
	wire [2:0] w_G234_1;
	wire [1:0] w_G234_2;
	wire [2:0] w_G242_0;
	wire [1:0] w_G242_1;
	wire [1:0] w_G245_0;
	wire [2:0] w_G248_0;
	wire [2:0] w_G248_1;
	wire [2:0] w_G248_2;
	wire [2:0] w_G248_3;
	wire [2:0] w_G248_4;
	wire [2:0] w_G248_5;
	wire [2:0] w_G251_0;
	wire [2:0] w_G251_1;
	wire [2:0] w_G251_2;
	wire [2:0] w_G251_3;
	wire [2:0] w_G251_4;
	wire [1:0] w_G251_5;
	wire [2:0] w_G254_0;
	wire [1:0] w_G254_1;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [1:0] w_G257_2;
	wire [2:0] w_G265_0;
	wire [2:0] w_G265_1;
	wire [2:0] w_G273_0;
	wire [2:0] w_G273_1;
	wire [1:0] w_G273_2;
	wire [2:0] w_G281_0;
	wire [2:0] w_G281_1;
	wire [1:0] w_G281_2;
	wire [1:0] w_G289_0;
	wire [2:0] w_G293_0;
	wire [2:0] w_G299_0;
	wire [2:0] w_G302_0;
	wire [2:0] w_G308_0;
	wire [2:0] w_G308_1;
	wire [2:0] w_G316_0;
	wire [1:0] w_G316_1;
	wire [2:0] w_G324_0;
	wire [2:0] w_G324_1;
	wire [1:0] w_G331_0;
	wire [2:0] w_G332_0;
	wire [2:0] w_G332_1;
	wire [2:0] w_G332_2;
	wire [2:0] w_G332_3;
	wire [2:0] w_G335_0;
	wire [1:0] w_G338_0;
	wire [2:0] w_G341_0;
	wire [2:0] w_G341_1;
	wire [2:0] w_G341_2;
	wire [1:0] w_G348_0;
	wire [2:0] w_G351_0;
	wire [2:0] w_G351_1;
	wire [2:0] w_G351_2;
	wire [1:0] w_G358_0;
	wire [2:0] w_G361_0;
	wire [1:0] w_G361_1;
	wire [1:0] w_G366_0;
	wire [1:0] w_G369_0;
	wire [2:0] w_G374_0;
	wire [2:0] w_G374_1;
	wire [2:0] w_G389_0;
	wire [2:0] w_G389_1;
	wire [2:0] w_G400_0;
	wire [2:0] w_G400_1;
	wire [2:0] w_G411_0;
	wire [2:0] w_G411_1;
	wire [1:0] w_G411_2;
	wire [2:0] w_G422_0;
	wire [1:0] w_G422_1;
	wire [2:0] w_G435_0;
	wire [2:0] w_G435_1;
	wire [2:0] w_G446_0;
	wire [2:0] w_G446_1;
	wire [2:0] w_G457_0;
	wire [2:0] w_G457_1;
	wire [2:0] w_G468_0;
	wire [2:0] w_G468_1;
	wire [2:0] w_G479_0;
	wire [2:0] w_G490_0;
	wire [1:0] w_G490_1;
	wire [2:0] w_G503_0;
	wire [2:0] w_G503_1;
	wire [1:0] w_G503_2;
	wire [2:0] w_G514_0;
	wire [2:0] w_G514_1;
	wire [1:0] w_G514_2;
	wire [2:0] w_G523_0;
	wire [2:0] w_G523_1;
	wire [2:0] w_G534_0;
	wire [2:0] w_G534_1;
	wire [1:0] w_G534_2;
	wire [2:0] w_G545_0;
	wire [2:0] w_G549_0;
	wire [1:0] w_G552_0;
	wire [1:0] w_G559_0;
	wire [1:0] w_G562_0;
	wire [2:0] w_G1497_0;
	wire [2:0] w_G1689_0;
	wire [2:0] w_G1689_1;
	wire [2:0] w_G1689_2;
	wire [2:0] w_G1689_3;
	wire [2:0] w_G1689_4;
	wire [1:0] w_G1689_5;
	wire [2:0] w_G1690_0;
	wire [1:0] w_G1690_1;
	wire [2:0] w_G1691_0;
	wire [2:0] w_G1691_1;
	wire [2:0] w_G1691_2;
	wire [2:0] w_G1691_3;
	wire [2:0] w_G1691_4;
	wire [1:0] w_G1691_5;
	wire [2:0] w_G1694_0;
	wire [1:0] w_G1694_1;
	wire [2:0] w_G2174_0;
	wire [2:0] w_G2358_0;
	wire [2:0] w_G2358_1;
	wire [2:0] w_G2358_2;
	wire [1:0] w_G3173_0;
	wire [2:0] w_G3546_0;
	wire [2:0] w_G3546_1;
	wire [2:0] w_G3546_2;
	wire [2:0] w_G3546_3;
	wire [2:0] w_G3546_4;
	wire [1:0] w_G3546_5;
	wire [2:0] w_G3548_0;
	wire [2:0] w_G3548_1;
	wire [2:0] w_G3548_2;
	wire [2:0] w_G3548_3;
	wire [2:0] w_G3548_4;
	wire [1:0] w_G3552_0;
	wire [1:0] w_G3717_0;
	wire [2:0] w_G3724_0;
	wire [2:0] w_G4087_0;
	wire [2:0] w_G4087_1;
	wire [2:0] w_G4087_2;
	wire [2:0] w_G4087_3;
	wire [2:0] w_G4087_4;
	wire [2:0] w_G4088_0;
	wire [2:0] w_G4088_1;
	wire [2:0] w_G4088_2;
	wire [2:0] w_G4088_3;
	wire [2:0] w_G4088_4;
	wire [2:0] w_G4088_5;
	wire [2:0] w_G4088_6;
	wire [2:0] w_G4088_7;
	wire [2:0] w_G4088_8;
	wire [2:0] w_G4088_9;
	wire [2:0] w_G4089_0;
	wire [2:0] w_G4089_1;
	wire [2:0] w_G4089_2;
	wire [2:0] w_G4089_3;
	wire [2:0] w_G4089_4;
	wire [2:0] w_G4089_5;
	wire [2:0] w_G4089_6;
	wire [2:0] w_G4089_7;
	wire [2:0] w_G4089_8;
	wire [2:0] w_G4089_9;
	wire [2:0] w_G4090_0;
	wire [2:0] w_G4090_1;
	wire [2:0] w_G4090_2;
	wire [2:0] w_G4090_3;
	wire [2:0] w_G4090_4;
	wire [2:0] w_G4091_0;
	wire [2:0] w_G4091_1;
	wire [2:0] w_G4091_2;
	wire [2:0] w_G4091_3;
	wire [2:0] w_G4091_4;
	wire [2:0] w_G4091_5;
	wire [1:0] w_G4091_6;
	wire [2:0] w_G4092_0;
	wire [2:0] w_G4092_1;
	wire [2:0] w_G4092_2;
	wire [2:0] w_G4092_3;
	wire [2:0] w_G4092_4;
	wire [2:0] w_G4092_5;
	wire [2:0] w_G4092_6;
	wire [2:0] w_G4092_7;
	wire [2:0] w_G4092_8;
	wire [2:0] w_G4092_9;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire [2:0] w_G809_0;
	wire [2:0] w_G809_1;
	wire [2:0] w_G809_2;
	wire [1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G623_0;
	wire G623_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G998_0;
	wire G998_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G865_0;
	wire G865_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire [1:0] w_n316_0;
	wire [1:0] w_n318_0;
	wire [2:0] w_n326_0;
	wire [2:0] w_n326_1;
	wire [1:0] w_n326_2;
	wire [1:0] w_n333_0;
	wire [1:0] w_n336_0;
	wire [1:0] w_n361_0;
	wire [1:0] w_n365_0;
	wire [2:0] w_n366_0;
	wire [2:0] w_n366_1;
	wire [2:0] w_n369_0;
	wire [2:0] w_n369_1;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [2:0] w_n374_0;
	wire [1:0] w_n374_1;
	wire [2:0] w_n375_0;
	wire [2:0] w_n375_1;
	wire [2:0] w_n375_2;
	wire [2:0] w_n375_3;
	wire [2:0] w_n375_4;
	wire [2:0] w_n377_0;
	wire [1:0] w_n377_1;
	wire [2:0] w_n378_0;
	wire [2:0] w_n378_1;
	wire [2:0] w_n378_2;
	wire [2:0] w_n378_3;
	wire [2:0] w_n378_4;
	wire [1:0] w_n386_0;
	wire [2:0] w_n387_0;
	wire [1:0] w_n387_1;
	wire [2:0] w_n389_0;
	wire [1:0] w_n389_1;
	wire [1:0] w_n397_0;
	wire [1:0] w_n401_0;
	wire [2:0] w_n402_0;
	wire [2:0] w_n406_0;
	wire [2:0] w_n406_1;
	wire [2:0] w_n406_2;
	wire [2:0] w_n406_3;
	wire [2:0] w_n406_4;
	wire [1:0] w_n406_5;
	wire [2:0] w_n408_0;
	wire [2:0] w_n408_1;
	wire [2:0] w_n408_2;
	wire [2:0] w_n408_3;
	wire [2:0] w_n408_4;
	wire [2:0] w_n408_5;
	wire [2:0] w_n412_0;
	wire [1:0] w_n414_0;
	wire [1:0] w_n415_0;
	wire [2:0] w_n423_0;
	wire [2:0] w_n425_0;
	wire [2:0] w_n428_0;
	wire [1:0] w_n428_1;
	wire [1:0] w_n429_0;
	wire [2:0] w_n433_0;
	wire [2:0] w_n435_0;
	wire [2:0] w_n435_1;
	wire [1:0] w_n435_2;
	wire [1:0] w_n437_0;
	wire [1:0] w_n445_0;
	wire [2:0] w_n449_0;
	wire [2:0] w_n449_1;
	wire [2:0] w_n451_0;
	wire [1:0] w_n459_0;
	wire [2:0] w_n460_0;
	wire [2:0] w_n460_1;
	wire [2:0] w_n462_0;
	wire [1:0] w_n470_0;
	wire [2:0] w_n471_0;
	wire [2:0] w_n471_1;
	wire [2:0] w_n473_0;
	wire [1:0] w_n473_1;
	wire [1:0] w_n481_0;
	wire [2:0] w_n483_0;
	wire [2:0] w_n483_1;
	wire [1:0] w_n483_2;
	wire [2:0] w_n485_0;
	wire [1:0] w_n485_1;
	wire [1:0] w_n493_0;
	wire [2:0] w_n494_0;
	wire [2:0] w_n494_1;
	wire [2:0] w_n496_0;
	wire [1:0] w_n496_1;
	wire [1:0] w_n504_0;
	wire [2:0] w_n507_0;
	wire [2:0] w_n507_1;
	wire [2:0] w_n509_0;
	wire [1:0] w_n517_0;
	wire [2:0] w_n518_0;
	wire [2:0] w_n518_1;
	wire [2:0] w_n520_0;
	wire [1:0] w_n528_0;
	wire [2:0] w_n530_0;
	wire [2:0] w_n530_1;
	wire [2:0] w_n532_0;
	wire [1:0] w_n532_1;
	wire [1:0] w_n540_0;
	wire [1:0] w_n543_0;
	wire [2:0] w_n551_0;
	wire [2:0] w_n556_0;
	wire [2:0] w_n556_1;
	wire [2:0] w_n556_2;
	wire [2:0] w_n556_3;
	wire [2:0] w_n556_4;
	wire [2:0] w_n556_5;
	wire [2:0] w_n556_6;
	wire [2:0] w_n556_7;
	wire [1:0] w_n556_8;
	wire [1:0] w_n557_0;
	wire [1:0] w_n559_0;
	wire [2:0] w_n560_0;
	wire [2:0] w_n561_0;
	wire [1:0] w_n561_1;
	wire [1:0] w_n562_0;
	wire [1:0] w_n564_0;
	wire [2:0] w_n565_0;
	wire [2:0] w_n566_0;
	wire [2:0] w_n567_0;
	wire [1:0] w_n569_0;
	wire [1:0] w_n571_0;
	wire [2:0] w_n572_0;
	wire [2:0] w_n573_0;
	wire [2:0] w_n574_0;
	wire [2:0] w_n578_0;
	wire [1:0] w_n578_1;
	wire [2:0] w_n579_0;
	wire [1:0] w_n579_1;
	wire [1:0] w_n581_0;
	wire [2:0] w_n586_0;
	wire [1:0] w_n586_1;
	wire [1:0] w_n587_0;
	wire [2:0] w_n588_0;
	wire [1:0] w_n588_1;
	wire [2:0] w_n591_0;
	wire [1:0] w_n591_1;
	wire [2:0] w_n592_0;
	wire [2:0] w_n596_0;
	wire [1:0] w_n596_1;
	wire [2:0] w_n597_0;
	wire [2:0] w_n601_0;
	wire [1:0] w_n601_1;
	wire [2:0] w_n602_0;
	wire [1:0] w_n603_0;
	wire [2:0] w_n607_0;
	wire [1:0] w_n607_1;
	wire [2:0] w_n608_0;
	wire [2:0] w_n609_0;
	wire [2:0] w_n611_0;
	wire [2:0] w_n613_0;
	wire [2:0] w_n613_1;
	wire [2:0] w_n613_2;
	wire [2:0] w_n613_3;
	wire [2:0] w_n613_4;
	wire [2:0] w_n613_5;
	wire [2:0] w_n617_0;
	wire [1:0] w_n617_1;
	wire [2:0] w_n618_0;
	wire [2:0] w_n619_0;
	wire [2:0] w_n619_1;
	wire [2:0] w_n620_0;
	wire [1:0] w_n620_1;
	wire [1:0] w_n621_0;
	wire [1:0] w_n623_0;
	wire [2:0] w_n624_0;
	wire [1:0] w_n625_0;
	wire [2:0] w_n627_0;
	wire [1:0] w_n627_1;
	wire [2:0] w_n628_0;
	wire [1:0] w_n631_0;
	wire [1:0] w_n632_0;
	wire [2:0] w_n635_0;
	wire [1:0] w_n635_1;
	wire [2:0] w_n636_0;
	wire [2:0] w_n637_0;
	wire [1:0] w_n638_0;
	wire [2:0] w_n639_0;
	wire [1:0] w_n640_0;
	wire [2:0] w_n641_0;
	wire [2:0] w_n641_1;
	wire [2:0] w_n644_0;
	wire [2:0] w_n648_0;
	wire [1:0] w_n648_1;
	wire [1:0] w_n649_0;
	wire [1:0] w_n650_0;
	wire [2:0] w_n653_0;
	wire [2:0] w_n654_0;
	wire [2:0] w_n654_1;
	wire [2:0] w_n654_2;
	wire [2:0] w_n658_0;
	wire [1:0] w_n658_1;
	wire [1:0] w_n659_0;
	wire [2:0] w_n660_0;
	wire [1:0] w_n660_1;
	wire [1:0] w_n661_0;
	wire [1:0] w_n670_0;
	wire [1:0] w_n680_0;
	wire [2:0] w_n682_0;
	wire [1:0] w_n684_0;
	wire [1:0] w_n685_0;
	wire [1:0] w_n686_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n689_0;
	wire [1:0] w_n690_0;
	wire [1:0] w_n692_0;
	wire [2:0] w_n694_0;
	wire [2:0] w_n695_0;
	wire [2:0] w_n699_0;
	wire [1:0] w_n701_0;
	wire [2:0] w_n703_0;
	wire [1:0] w_n704_0;
	wire [1:0] w_n709_0;
	wire [1:0] w_n710_0;
	wire [1:0] w_n711_0;
	wire [2:0] w_n713_0;
	wire [2:0] w_n715_0;
	wire [1:0] w_n717_0;
	wire [1:0] w_n719_0;
	wire [1:0] w_n720_0;
	wire [1:0] w_n721_0;
	wire [1:0] w_n722_0;
	wire [2:0] w_n725_0;
	wire [1:0] w_n726_0;
	wire [1:0] w_n728_0;
	wire [2:0] w_n733_0;
	wire [2:0] w_n735_0;
	wire [2:0] w_n737_0;
	wire [1:0] w_n737_1;
	wire [1:0] w_n738_0;
	wire [2:0] w_n742_0;
	wire [1:0] w_n745_0;
	wire [2:0] w_n746_0;
	wire [1:0] w_n747_0;
	wire [2:0] w_n749_0;
	wire [2:0] w_n749_1;
	wire [2:0] w_n749_2;
	wire [2:0] w_n749_3;
	wire [2:0] w_n749_4;
	wire [2:0] w_n749_5;
	wire [2:0] w_n749_6;
	wire [2:0] w_n749_7;
	wire [2:0] w_n749_8;
	wire [2:0] w_n749_9;
	wire [2:0] w_n749_10;
	wire [2:0] w_n749_11;
	wire [2:0] w_n749_12;
	wire [1:0] w_n749_13;
	wire [2:0] w_n750_0;
	wire [2:0] w_n750_1;
	wire [2:0] w_n750_2;
	wire [2:0] w_n750_3;
	wire [2:0] w_n750_4;
	wire [2:0] w_n750_5;
	wire [2:0] w_n750_6;
	wire [2:0] w_n750_7;
	wire [2:0] w_n750_8;
	wire [2:0] w_n753_0;
	wire [1:0] w_n753_1;
	wire [1:0] w_n755_0;
	wire [2:0] w_n763_0;
	wire [1:0] w_n767_0;
	wire [1:0] w_n779_0;
	wire [2:0] w_n786_0;
	wire [2:0] w_n788_0;
	wire [2:0] w_n790_0;
	wire [2:0] w_n792_0;
	wire [2:0] w_n795_0;
	wire [1:0] w_n795_1;
	wire [2:0] w_n797_0;
	wire [2:0] w_n797_1;
	wire [2:0] w_n797_2;
	wire [2:0] w_n797_3;
	wire [2:0] w_n797_4;
	wire [2:0] w_n797_5;
	wire [2:0] w_n797_6;
	wire [2:0] w_n797_7;
	wire [2:0] w_n797_8;
	wire [1:0] w_n797_9;
	wire [2:0] w_n798_0;
	wire [1:0] w_n798_1;
	wire [2:0] w_n800_0;
	wire [2:0] w_n800_1;
	wire [2:0] w_n800_2;
	wire [2:0] w_n800_3;
	wire [1:0] w_n800_4;
	wire [2:0] w_n801_0;
	wire [1:0] w_n801_1;
	wire [2:0] w_n814_0;
	wire [2:0] w_n819_0;
	wire [1:0] w_n821_0;
	wire [1:0] w_n824_0;
	wire [1:0] w_n827_0;
	wire [1:0] w_n836_0;
	wire [1:0] w_n847_0;
	wire [2:0] w_n852_0;
	wire [2:0] w_n852_1;
	wire [2:0] w_n852_2;
	wire [2:0] w_n852_3;
	wire [2:0] w_n852_4;
	wire [2:0] w_n852_5;
	wire [2:0] w_n852_6;
	wire [2:0] w_n852_7;
	wire [2:0] w_n852_8;
	wire [1:0] w_n852_9;
	wire [2:0] w_n854_0;
	wire [2:0] w_n854_1;
	wire [2:0] w_n854_2;
	wire [2:0] w_n854_3;
	wire [1:0] w_n854_4;
	wire [2:0] w_n865_0;
	wire [1:0] w_n867_0;
	wire [1:0] w_n868_0;
	wire [1:0] w_n870_0;
	wire [1:0] w_n871_0;
	wire [1:0] w_n880_0;
	wire [1:0] w_n890_0;
	wire [1:0] w_n901_0;
	wire [2:0] w_n923_0;
	wire [1:0] w_n935_0;
	wire [2:0] w_n938_0;
	wire [2:0] w_n940_0;
	wire [1:0] w_n940_1;
	wire [1:0] w_n944_0;
	wire [1:0] w_n949_0;
	wire [1:0] w_n953_0;
	wire [2:0] w_n954_0;
	wire [1:0] w_n957_0;
	wire [1:0] w_n962_0;
	wire [1:0] w_n964_0;
	wire [1:0] w_n969_0;
	wire [2:0] w_n977_0;
	wire [1:0] w_n981_0;
	wire [1:0] w_n986_0;
	wire [1:0] w_n989_0;
	wire [2:0] w_n993_0;
	wire [2:0] w_n993_1;
	wire [2:0] w_n993_2;
	wire [2:0] w_n993_3;
	wire [2:0] w_n993_4;
	wire [2:0] w_n994_0;
	wire [2:0] w_n994_1;
	wire [2:0] w_n994_2;
	wire [2:0] w_n994_3;
	wire [1:0] w_n994_4;
	wire [2:0] w_n996_0;
	wire [2:0] w_n996_1;
	wire [2:0] w_n996_2;
	wire [2:0] w_n996_3;
	wire [1:0] w_n996_4;
	wire [2:0] w_n999_0;
	wire [2:0] w_n999_1;
	wire [2:0] w_n999_2;
	wire [2:0] w_n999_3;
	wire [2:0] w_n1007_0;
	wire [2:0] w_n1007_1;
	wire [2:0] w_n1007_2;
	wire [2:0] w_n1007_3;
	wire [2:0] w_n1008_0;
	wire [2:0] w_n1008_1;
	wire [2:0] w_n1008_2;
	wire [2:0] w_n1008_3;
	wire [2:0] w_n1008_4;
	wire [2:0] w_n1012_0;
	wire [2:0] w_n1012_1;
	wire [2:0] w_n1012_2;
	wire [2:0] w_n1012_3;
	wire [1:0] w_n1012_4;
	wire [2:0] w_n1014_0;
	wire [2:0] w_n1014_1;
	wire [2:0] w_n1014_2;
	wire [2:0] w_n1014_3;
	wire [1:0] w_n1014_4;
	wire [2:0] w_n1019_0;
	wire [1:0] w_n1019_1;
	wire [2:0] w_n1021_0;
	wire [1:0] w_n1021_1;
	wire [2:0] w_n1030_0;
	wire [1:0] w_n1030_1;
	wire [2:0] w_n1032_0;
	wire [1:0] w_n1032_1;
	wire [2:0] w_n1041_0;
	wire [1:0] w_n1041_1;
	wire [2:0] w_n1043_0;
	wire [1:0] w_n1043_1;
	wire [2:0] w_n1052_0;
	wire [1:0] w_n1052_1;
	wire [2:0] w_n1054_0;
	wire [1:0] w_n1054_1;
	wire [1:0] w_n1177_0;
	wire [1:0] w_n1179_0;
	wire [2:0] w_n1196_0;
	wire [2:0] w_n1196_1;
	wire [2:0] w_n1201_0;
	wire [2:0] w_n1205_0;
	wire [2:0] w_n1205_1;
	wire [2:0] w_n1213_0;
	wire [2:0] w_n1213_1;
	wire [2:0] w_n1236_0;
	wire [2:0] w_n1236_1;
	wire [2:0] w_n1251_0;
	wire [2:0] w_n1251_1;
	wire [2:0] w_n1279_0;
	wire [1:0] w_n1279_1;
	wire [2:0] w_n1297_0;
	wire [1:0] w_n1297_1;
	wire [2:0] w_n1299_0;
	wire [1:0] w_n1299_1;
	wire [2:0] w_n1410_0;
	wire [2:0] w_n1412_0;
	wire [1:0] w_n1416_0;
	wire [1:0] w_n1422_0;
	wire [1:0] w_n1425_0;
	wire [1:0] w_n1428_0;
	wire [1:0] w_n1429_0;
	wire [1:0] w_n1451_0;
	wire [1:0] w_n1503_0;
	wire [1:0] w_n1504_0;
	wire [1:0] w_n1592_0;
	wire [1:0] w_n1593_0;
	wire [1:0] w_n1596_0;
	wire [1:0] w_n1599_0;
	wire [1:0] w_n1603_0;
	wire [1:0] w_n1605_0;
	wire [1:0] w_n1609_0;
	wire [2:0] w_n1611_0;
	wire [1:0] w_n1613_0;
	wire [1:0] w_n1615_0;
	wire [1:0] w_n1618_0;
	wire [1:0] w_n1633_0;
	wire [1:0] w_n1637_0;
	wire [1:0] w_n1643_0;
	wire [1:0] w_n1652_0;
	wire [1:0] w_n1665_0;
	wire [2:0] w_n1674_0;
	wire [1:0] w_n1675_0;
	wire [2:0] w_n1679_0;
	wire [1:0] w_n1680_0;
	wire [1:0] w_n1694_0;
	wire [1:0] w_n1695_0;
	wire [1:0] w_n1698_0;
	wire w_dff_B_xJVd7vh19_1;
	wire w_dff_B_NeekBaFp4_0;
	wire w_dff_B_H5ICgJDO2_1;
	wire w_dff_B_T4h4UUWo7_1;
	wire w_dff_B_m9fN94CJ9_2;
	wire w_dff_B_FiSJvVee4_1;
	wire w_dff_B_V1WkeonP1_1;
	wire w_dff_B_dFPnBT7I9_0;
	wire w_dff_B_AUPL4UiY9_1;
	wire w_dff_B_ELkE3jRs4_1;
	wire w_dff_B_PDYKQJxI2_0;
	wire w_dff_B_u5UjHSah1_1;
	wire w_dff_A_EyYMh1gb3_0;
	wire w_dff_A_hBgOeFl60_0;
	wire w_dff_A_naU6d0v53_0;
	wire w_dff_A_G139qUXC6_0;
	wire w_dff_A_isseKvlO1_1;
	wire w_dff_A_V6aJmz8T1_1;
	wire w_dff_A_z4bRBYaS8_1;
	wire w_dff_A_9pMjfsWj9_1;
	wire w_dff_B_7UYQIOoi0_1;
	wire w_dff_B_Mo4niKpk5_0;
	wire w_dff_B_9OtLNadY3_1;
	wire w_dff_B_KSukqhV45_1;
	wire w_dff_B_kBiuCscR6_1;
	wire w_dff_B_OnyUwNWl5_1;
	wire w_dff_A_5H7xdybX2_0;
	wire w_dff_A_tmZmnfvl0_1;
	wire w_dff_A_2bn3N6YZ7_1;
	wire w_dff_A_3GYoWiuU0_1;
	wire w_dff_A_6YSjiHj03_1;
	wire w_dff_A_TU9gGnzH5_1;
	wire w_dff_A_kMWxVDrh2_2;
	wire w_dff_A_jZ6qwYt01_2;
	wire w_dff_A_bRtp74It2_2;
	wire w_dff_A_edFeGmke8_2;
	wire w_dff_B_ppgzI1QW4_1;
	wire w_dff_B_WslEtSt70_2;
	wire w_dff_B_tLzJNkdT5_2;
	wire w_dff_B_Tm0nih7h7_2;
	wire w_dff_B_QAeNhS517_2;
	wire w_dff_B_HxvTgeKW1_1;
	wire w_dff_B_MCOzTeU11_1;
	wire w_dff_B_LM8uvOAs5_1;
	wire w_dff_B_Wl4ntgBJ8_1;
	wire w_dff_B_EUhZeJeu1_1;
	wire w_dff_B_QUdYuxkV7_1;
	wire w_dff_B_0mqaafZo4_1;
	wire w_dff_B_wDUsRAim3_1;
	wire w_dff_B_0oPw1zAC4_1;
	wire w_dff_B_SWBiYy6v8_1;
	wire w_dff_B_V8QbOeQJ2_1;
	wire w_dff_A_qgprgtJz4_1;
	wire w_dff_A_27kRFvmS5_1;
	wire w_dff_B_Gk7CQZEh4_3;
	wire w_dff_B_rVPAffzR7_2;
	wire w_dff_B_pKIMdEps8_2;
	wire w_dff_B_Ug8Ns8L68_1;
	wire w_dff_B_faKqSggN7_1;
	wire w_dff_A_TUQM28mg7_0;
	wire w_dff_A_LqDBCJup0_0;
	wire w_dff_A_hOsm0uFm5_0;
	wire w_dff_A_33gZIik94_0;
	wire w_dff_A_38Pjr5fa8_0;
	wire w_dff_B_8A802oyh5_0;
	wire w_dff_B_OPIUQjYO2_0;
	wire w_dff_B_VKWfFFBw6_0;
	wire w_dff_B_3alZRvZ45_0;
	wire w_dff_B_ZsBQnEA47_0;
	wire w_dff_B_NPYzj9ey3_0;
	wire w_dff_B_SESaneVA4_0;
	wire w_dff_B_GIU1vtYK0_0;
	wire w_dff_B_5IETn2KG4_0;
	wire w_dff_B_oplNXEDL6_0;
	wire w_dff_B_1PScmEgp4_0;
	wire w_dff_A_c8nKUhZi0_1;
	wire w_dff_A_seo738dG0_1;
	wire w_dff_A_HOayV5bp4_1;
	wire w_dff_A_AjbdDBgO6_1;
	wire w_dff_A_0T4J5fkg1_1;
	wire w_dff_A_dmjpzGTR8_1;
	wire w_dff_A_EKuwZTdH8_1;
	wire w_dff_A_iOrnd5Pj3_1;
	wire w_dff_A_zISZqvFC3_1;
	wire w_dff_A_losgSMuX1_1;
	wire w_dff_B_t0Lv9bLg5_0;
	wire w_dff_B_IY6zNTzk1_0;
	wire w_dff_B_Y1Crni0n0_0;
	wire w_dff_B_2lQCkvPH6_0;
	wire w_dff_B_DwmqAbxu1_0;
	wire w_dff_B_yO2Ld9hd1_0;
	wire w_dff_B_Wm19bM8k6_0;
	wire w_dff_B_CCcAZDDj1_0;
	wire w_dff_B_IdQgVWDq7_0;
	wire w_dff_B_ka2cL7cq3_0;
	wire w_dff_B_5Pi8sLZf6_2;
	wire w_dff_B_Zj1aWoW30_0;
	wire w_dff_A_aRXDzq5t5_1;
	wire w_dff_A_54vCDj965_1;
	wire w_dff_A_Tjsbs8C07_1;
	wire w_dff_A_DjrPyRvT1_1;
	wire w_dff_A_RFF4a3Id4_1;
	wire w_dff_A_MGMIOyFU5_1;
	wire w_dff_A_SmllZ8dT6_1;
	wire w_dff_A_R7B2ihJO3_1;
	wire w_dff_A_Q5mkiUxB4_1;
	wire w_dff_A_GStFKiis3_1;
	wire w_dff_B_ifnOJc1U1_0;
	wire w_dff_B_ynuAR34F0_1;
	wire w_dff_B_bZ4GVU5u1_1;
	wire w_dff_B_nTaXBT9q0_1;
	wire w_dff_B_iqLddp8R8_0;
	wire w_dff_B_a6qgBGCl0_1;
	wire w_dff_B_cm89qgb02_1;
	wire w_dff_B_Y4rYfPA96_1;
	wire w_dff_B_qLpZPYUP7_1;
	wire w_dff_B_AxD9PwDr3_1;
	wire w_dff_B_0mYtizdg0_1;
	wire w_dff_B_CpVbdhlH2_1;
	wire w_dff_B_rpc69Qrr7_1;
	wire w_dff_B_jNILjL1c7_1;
	wire w_dff_B_M9tgOfoG7_1;
	wire w_dff_B_iFErXtgI2_1;
	wire w_dff_B_emGytDbn3_1;
	wire w_dff_B_2fWqJBgV3_1;
	wire w_dff_B_YPTvsFTT1_1;
	wire w_dff_B_xOad4M3p8_1;
	wire w_dff_B_fHaFuXNL2_1;
	wire w_dff_B_WddvAmdt9_1;
	wire w_dff_B_bIlR0n4s5_1;
	wire w_dff_B_bepvfav89_1;
	wire w_dff_B_PmBeLX548_1;
	wire w_dff_B_rzfiyyni7_1;
	wire w_dff_B_KQ2RIcrD9_1;
	wire w_dff_B_wEc3UVnu1_1;
	wire w_dff_B_oAnQ5GPc4_1;
	wire w_dff_B_3BuDIKdG0_1;
	wire w_dff_B_GQUnHn8g1_1;
	wire w_dff_B_eqL0ZiLh0_1;
	wire w_dff_B_pBC8bezt1_1;
	wire w_dff_B_zadYHcFr1_1;
	wire w_dff_B_gGhJvAVX2_0;
	wire w_dff_B_YFsucXNK3_0;
	wire w_dff_B_NX7qa5h72_0;
	wire w_dff_B_yX0JgzqU5_0;
	wire w_dff_B_P8VxAMFw6_0;
	wire w_dff_B_hu4syHSm8_0;
	wire w_dff_B_JB8MMbPs8_0;
	wire w_dff_B_LsuiAY8o2_0;
	wire w_dff_B_6zHzrdVX2_0;
	wire w_dff_B_V17nTjdJ3_0;
	wire w_dff_B_Ma1gKVog9_0;
	wire w_dff_B_s0XwuCNn0_1;
	wire w_dff_B_TEwl3wgg6_2;
	wire w_dff_B_UXYvnfD98_2;
	wire w_dff_B_cX4vbk7M7_2;
	wire w_dff_B_TH3AsybK0_1;
	wire w_dff_B_pJs3TDkA4_1;
	wire w_dff_B_PSJp4qRu8_1;
	wire w_dff_B_llc5HBxt6_1;
	wire w_dff_B_tPDLTsEY6_1;
	wire w_dff_B_X4NEc9x47_1;
	wire w_dff_B_7H31U1To0_1;
	wire w_dff_B_0fwNjf782_1;
	wire w_dff_B_kwHGDFZX7_0;
	wire w_dff_B_u9pdidx38_1;
	wire w_dff_B_3XLwB3kW2_1;
	wire w_dff_A_0kNBMird8_0;
	wire w_dff_A_qnGRR56D9_0;
	wire w_dff_B_llH03iJn7_1;
	wire w_dff_B_uWQdhYHv7_1;
	wire w_dff_B_OT9KcLqn4_1;
	wire w_dff_B_GrmjhGxS4_1;
	wire w_dff_B_Wr6GDBT12_1;
	wire w_dff_A_3ZG8IpOA9_0;
	wire w_dff_A_68n6HSoo1_0;
	wire w_dff_A_ATfgVxmz3_0;
	wire w_dff_A_pJggtBVe3_0;
	wire w_dff_A_FkQn2sEm6_0;
	wire w_dff_A_MJ8r3R6z6_0;
	wire w_dff_A_DDxqCbB22_0;
	wire w_dff_A_9lKhqlHn3_0;
	wire w_dff_A_biLyGV7G6_0;
	wire w_dff_A_HR22AKG65_0;
	wire w_dff_A_AFcJoeIn8_0;
	wire w_dff_B_VjocPBUU2_1;
	wire w_dff_B_5JNCKSIB9_1;
	wire w_dff_B_6C7xYPwX4_0;
	wire w_dff_B_6usAEpL71_0;
	wire w_dff_B_DPoBePda6_0;
	wire w_dff_B_p43uRxwh4_0;
	wire w_dff_B_PXHs6AVa0_0;
	wire w_dff_B_NCJWC3Zs6_0;
	wire w_dff_B_C9UyJnCz3_0;
	wire w_dff_B_nT9GyZhR6_0;
	wire w_dff_B_4kE6BgE56_0;
	wire w_dff_B_GmDFS35I0_0;
	wire w_dff_B_VSsnlerl0_0;
	wire w_dff_B_SCP58RGa4_0;
	wire w_dff_B_017KG9S71_0;
	wire w_dff_B_9ldMJKpa4_0;
	wire w_dff_B_qmgLwixf3_0;
	wire w_dff_B_UIq314s07_0;
	wire w_dff_B_IsG2THwt3_1;
	wire w_dff_A_TZScAyTj2_0;
	wire w_dff_A_QNrzqIJH1_0;
	wire w_dff_A_9hnClhKi8_0;
	wire w_dff_A_L0En3HXn6_0;
	wire w_dff_A_3K82hbXV2_0;
	wire w_dff_A_OpI0ot5M8_0;
	wire w_dff_A_zylMXVli7_0;
	wire w_dff_B_Po2ISzVd5_0;
	wire w_dff_B_ZRmtmCjC7_0;
	wire w_dff_B_hTIicSsr5_0;
	wire w_dff_B_mTUB5HaQ7_0;
	wire w_dff_B_7hy4n0E68_0;
	wire w_dff_B_otWUI5sG6_0;
	wire w_dff_B_XS6BAxRR8_0;
	wire w_dff_B_HaHF3kcj8_0;
	wire w_dff_B_ZyqN2vLL3_0;
	wire w_dff_B_qYCT38415_0;
	wire w_dff_B_p8auc4tf7_0;
	wire w_dff_B_fqGVN7Vg8_0;
	wire w_dff_B_DXGhJf8M6_0;
	wire w_dff_B_uKusfTFG7_0;
	wire w_dff_B_EmJXUkSS3_0;
	wire w_dff_B_QvF7cfS06_1;
	wire w_dff_B_JNeHI5JZ0_1;
	wire w_dff_A_MQEkn3ZQ3_0;
	wire w_dff_A_8JSkwwNG0_0;
	wire w_dff_A_SD5aRq3n2_0;
	wire w_dff_A_yHlDPozQ3_0;
	wire w_dff_A_KIAw0P6t3_0;
	wire w_dff_A_tJYE0Yn30_0;
	wire w_dff_A_6uxWNdtr7_0;
	wire w_dff_A_UZllMLiM0_0;
	wire w_dff_A_t1A3h8wG4_0;
	wire w_dff_A_Vrkc4mDz8_0;
	wire w_dff_A_pjGbuDnr6_0;
	wire w_dff_A_Cp83xP6V3_0;
	wire w_dff_A_Cqi6r2G91_0;
	wire w_dff_A_PyUVJ6Sk0_0;
	wire w_dff_A_p986CboN5_0;
	wire w_dff_A_6a5PsfXW0_2;
	wire w_dff_A_XA8MWyHc0_2;
	wire w_dff_A_8kFdNVLW4_2;
	wire w_dff_A_5wl5X6Qu4_2;
	wire w_dff_A_2uSKnKuM9_2;
	wire w_dff_A_OXGEE86E0_2;
	wire w_dff_A_KFXFmrLM3_2;
	wire w_dff_A_DkQQXndv4_2;
	wire w_dff_A_yxXdYlDR6_2;
	wire w_dff_A_iG2oJDo61_2;
	wire w_dff_A_uGZtE6xb4_2;
	wire w_dff_A_m8qufn2Y3_2;
	wire w_dff_A_3jfaWwH20_2;
	wire w_dff_A_W5PlwJbf8_2;
	wire w_dff_A_qaMVEAhk2_2;
	wire w_dff_A_FgbyN03F3_2;
	wire w_dff_A_VvG59TxG9_0;
	wire w_dff_A_rzUZXHyG7_0;
	wire w_dff_A_nuSZUysl8_0;
	wire w_dff_A_OadZqIXw7_0;
	wire w_dff_A_k39D8FCz7_0;
	wire w_dff_A_wQb28WFR7_0;
	wire w_dff_A_Kpw8bXjQ3_0;
	wire w_dff_A_21fj1h7t2_0;
	wire w_dff_A_OayhSrbs8_0;
	wire w_dff_A_Uj7yy23O6_0;
	wire w_dff_A_0VW1blZh0_0;
	wire w_dff_A_aBn7HYKn3_0;
	wire w_dff_A_RMKQ9xKZ3_0;
	wire w_dff_A_wMSaZ8gK4_2;
	wire w_dff_A_W6bTy4494_2;
	wire w_dff_A_lKCBf1TV2_2;
	wire w_dff_A_CIauddfq1_2;
	wire w_dff_A_6YOhI7Sq3_2;
	wire w_dff_A_IKtUNxUx4_2;
	wire w_dff_A_FrqyaWoV3_2;
	wire w_dff_A_8v3wnTHs3_2;
	wire w_dff_A_zbAwwr7D1_2;
	wire w_dff_A_3GY1SmH09_2;
	wire w_dff_A_WVYYgkO42_2;
	wire w_dff_A_h1z21ejw0_2;
	wire w_dff_A_oATnb0JV4_2;
	wire w_dff_A_yvKF8FNS8_2;
	wire w_dff_A_szCXB5hr2_2;
	wire w_dff_B_K0taASR83_0;
	wire w_dff_B_fgCIVJWI4_0;
	wire w_dff_B_Q390yZn54_0;
	wire w_dff_B_yjwzU9cr8_0;
	wire w_dff_B_t7VcwXUB3_0;
	wire w_dff_B_kDLvE5YN3_0;
	wire w_dff_B_WDpM9Pgp1_0;
	wire w_dff_B_XiOc0Asl2_0;
	wire w_dff_B_peDalsoS3_0;
	wire w_dff_B_50vjEcMR2_0;
	wire w_dff_B_E6G42R591_0;
	wire w_dff_B_7gGHSTfS2_0;
	wire w_dff_B_5cicOMT37_0;
	wire w_dff_B_wp0a28OD5_1;
	wire w_dff_A_Jo3bcgaK9_1;
	wire w_dff_A_CDwIySkN4_1;
	wire w_dff_A_OnXB51Bp8_1;
	wire w_dff_A_M7YEE43P3_1;
	wire w_dff_A_kg6GLHO41_1;
	wire w_dff_A_sddRlp4C4_1;
	wire w_dff_A_zz3pZw4u9_1;
	wire w_dff_A_4ZzXPOML7_1;
	wire w_dff_A_b2kEv4le4_1;
	wire w_dff_A_PV1fhr5j4_1;
	wire w_dff_A_ReqLpIV65_1;
	wire w_dff_A_OTCTdaMt9_1;
	wire w_dff_A_0ZF2PpQz8_1;
	wire w_dff_A_dfc0ZRY10_1;
	wire w_dff_A_wZfI1sYx5_1;
	wire w_dff_A_L00xSYiA9_1;
	wire w_dff_A_9hH4qnTQ4_1;
	wire w_dff_A_lfyjIjk33_1;
	wire w_dff_A_KwGtuKwl6_1;
	wire w_dff_A_rDygWqJN8_1;
	wire w_dff_A_S0JEouFS1_1;
	wire w_dff_A_kWWrLE427_1;
	wire w_dff_A_mipak4EX4_1;
	wire w_dff_A_z1tFrmCv4_1;
	wire w_dff_A_J40c4J9p9_1;
	wire w_dff_B_WvLGDAOl0_0;
	wire w_dff_B_OdkadJJI6_0;
	wire w_dff_B_CmNxNxjB0_0;
	wire w_dff_B_oBXown095_0;
	wire w_dff_B_cCeYb6eM9_0;
	wire w_dff_B_JQWwtTVl8_0;
	wire w_dff_B_nUqsHqs90_0;
	wire w_dff_B_ml71n9Iu4_0;
	wire w_dff_B_Y1IV97me7_0;
	wire w_dff_B_yL46Ax4v3_0;
	wire w_dff_B_fh5LHN6Z9_0;
	wire w_dff_B_yEGekuBd7_0;
	wire w_dff_B_WT21Q8Wg1_0;
	wire w_dff_B_PrVErDRB6_0;
	wire w_dff_B_pOXsZQ7t5_1;
	wire w_dff_B_TzjUy8CR7_1;
	wire w_dff_B_BkBJegN79_1;
	wire w_dff_A_foNLMS0P2_0;
	wire w_dff_A_Hu32o2cR8_2;
	wire w_dff_A_ptkvh7EA1_2;
	wire w_dff_B_3CTSQPKb8_1;
	wire w_dff_B_fijrpWob9_1;
	wire w_dff_B_cH8S5oks3_1;
	wire w_dff_B_E5l4s9jY8_1;
	wire w_dff_B_zycsE9ZW7_1;
	wire w_dff_B_7ZP9AhMz0_1;
	wire w_dff_B_a5S6kHUC3_1;
	wire w_dff_B_0YZn9x8B0_1;
	wire w_dff_B_SbA090H36_1;
	wire w_dff_B_DRl243DJ4_1;
	wire w_dff_B_SsELJ9Fa7_1;
	wire w_dff_B_JRRzcMFs5_1;
	wire w_dff_B_2xTmNc0b9_1;
	wire w_dff_B_EitWhjPr9_1;
	wire w_dff_B_sw0kQIIT5_1;
	wire w_dff_A_ebht2U5w7_0;
	wire w_dff_A_hV5J1of21_0;
	wire w_dff_A_sy4FFc0i5_0;
	wire w_dff_A_EB8dtqpN0_0;
	wire w_dff_A_4nLjo1g16_0;
	wire w_dff_A_p4UPIfMP6_0;
	wire w_dff_A_olaywdnc3_0;
	wire w_dff_A_p2PiHSc06_0;
	wire w_dff_B_KLHKgBge4_1;
	wire w_dff_B_fm2x8dKD1_1;
	wire w_dff_B_h9kxZlyU6_2;
	wire w_dff_B_fKlRZZMc0_1;
	wire w_dff_B_8ooZeVHK3_1;
	wire w_dff_B_X8ZmFST18_1;
	wire w_dff_B_krsKa70A5_1;
	wire w_dff_B_67anivFM8_1;
	wire w_dff_B_pcoQU6oO2_1;
	wire w_dff_B_qlaTCUvJ4_1;
	wire w_dff_B_iAz9VOY70_1;
	wire w_dff_B_4QN1Pk018_1;
	wire w_dff_B_eZD9rZFq6_1;
	wire w_dff_B_WIKI6WIU3_1;
	wire w_dff_B_gSEg92IP8_1;
	wire w_dff_B_1Ho6YZSd5_1;
	wire w_dff_B_R3xuKQ1A8_1;
	wire w_dff_B_3RUDA86W1_0;
	wire w_dff_B_FiZVK3de1_1;
	wire w_dff_B_dSaYggRw8_1;
	wire w_dff_A_CABZ38Nm4_1;
	wire w_dff_A_Mhpg5Sw66_1;
	wire w_dff_A_2f3ygkh53_1;
	wire w_dff_A_1pNpKMnn3_1;
	wire w_dff_A_UFtGMjOv9_1;
	wire w_dff_A_G7Upt35M5_1;
	wire w_dff_A_wHomhmqu2_1;
	wire w_dff_A_2evvlSFa6_1;
	wire w_dff_A_THPnx7fu3_1;
	wire w_dff_A_XpyDvBDb2_1;
	wire w_dff_A_svcPAzKj3_1;
	wire w_dff_A_otY84Bj83_1;
	wire w_dff_A_1xzMNccD6_1;
	wire w_dff_A_MIEN68w72_1;
	wire w_dff_A_p2KaDZoD7_1;
	wire w_dff_B_MZAmZeka7_2;
	wire w_dff_A_4gwFou728_1;
	wire w_dff_A_nDKLfZ6A8_1;
	wire w_dff_A_LVXdMjz14_1;
	wire w_dff_A_UMAllwSa6_1;
	wire w_dff_A_ZbHJusbg5_1;
	wire w_dff_A_eeUq2Ocq7_1;
	wire w_dff_A_2cVaDhVt5_1;
	wire w_dff_A_n6PN850D5_1;
	wire w_dff_A_OSHVIPAF3_1;
	wire w_dff_A_MCF6eygg6_1;
	wire w_dff_A_ATIub3M57_1;
	wire w_dff_A_cZyCyK2P3_1;
	wire w_dff_A_8MendlBx5_1;
	wire w_dff_A_4GTmbS0q8_1;
	wire w_dff_A_R5t2f0y17_1;
	wire w_dff_A_DGMxBQG38_1;
	wire w_dff_B_U62sgSUC8_1;
	wire w_dff_B_xB9NwQL76_1;
	wire w_dff_B_y19k6eIt3_1;
	wire w_dff_B_s05LFa7k9_1;
	wire w_dff_B_i3CRBM249_1;
	wire w_dff_B_S6GmqtZn9_1;
	wire w_dff_B_ul5oidY57_1;
	wire w_dff_B_fdimDfiK2_1;
	wire w_dff_B_3GWiesPE3_1;
	wire w_dff_B_AUFu4Drc0_1;
	wire w_dff_B_KDCB6Twn2_1;
	wire w_dff_B_QtbKjWVe1_1;
	wire w_dff_B_2Krg9KE16_1;
	wire w_dff_B_wsR42LE81_1;
	wire w_dff_A_AdgkasZo8_0;
	wire w_dff_A_3wMHiP440_0;
	wire w_dff_A_2CVtRpox0_0;
	wire w_dff_A_JpFHzrtN9_0;
	wire w_dff_A_4lukrovC8_0;
	wire w_dff_A_7HUDM1Yw4_0;
	wire w_dff_A_Azb8ug1R9_0;
	wire w_dff_A_Bb8YF7Ma6_0;
	wire w_dff_A_cQkQ1UbB1_0;
	wire w_dff_A_pcWhhPNn3_0;
	wire w_dff_A_fVceHLmP6_0;
	wire w_dff_A_z4pdcwoX3_0;
	wire w_dff_A_33GAKJi55_2;
	wire w_dff_A_EgB1K0cH3_2;
	wire w_dff_A_RUC4aArw9_2;
	wire w_dff_A_DunTaVRw4_2;
	wire w_dff_A_2ZDS1ZtK8_2;
	wire w_dff_A_o4Hb3cco8_2;
	wire w_dff_A_7SqNkHp28_2;
	wire w_dff_A_B21LMjTn3_2;
	wire w_dff_A_nB8D89q28_2;
	wire w_dff_A_HIX9uVYh9_2;
	wire w_dff_A_RyWzwAUx5_2;
	wire w_dff_A_98xNmKra5_2;
	wire w_dff_A_js8pimOP0_2;
	wire w_dff_B_RPIWd08X5_2;
	wire w_dff_A_H2jeIYjO1_0;
	wire w_dff_A_nrzLWmSR1_0;
	wire w_dff_A_44DkNbkz7_0;
	wire w_dff_A_m6WbrJ8L0_0;
	wire w_dff_A_lapcYyYX9_0;
	wire w_dff_A_O62LtL2A0_0;
	wire w_dff_A_5Gdr1D451_0;
	wire w_dff_A_XuHovybZ8_0;
	wire w_dff_A_Wc0Fc5UN9_0;
	wire w_dff_A_27Pe6pAY1_0;
	wire w_dff_A_pVhTbSdy7_0;
	wire w_dff_A_BUisNmyH8_0;
	wire w_dff_A_EGw3OCqi1_0;
	wire w_dff_A_oK2ZZWd80_2;
	wire w_dff_A_cbpnOs2t2_2;
	wire w_dff_A_1dQ0nBsJ4_2;
	wire w_dff_A_wnUlBMJS2_2;
	wire w_dff_A_tAIIr8Mb2_2;
	wire w_dff_A_U4VeFLT89_2;
	wire w_dff_A_0YTHVqHw1_2;
	wire w_dff_A_Uv1ru2fl1_2;
	wire w_dff_A_UYzecIFh4_2;
	wire w_dff_A_QgoiUmMT1_2;
	wire w_dff_A_TntnKZWC6_2;
	wire w_dff_A_P7p4HuS22_2;
	wire w_dff_A_6eMntC6i9_2;
	wire w_dff_A_i9DnFPfo7_2;
	wire w_dff_A_d2WmELSA3_2;
	wire w_dff_B_dwgKOCQT5_0;
	wire w_dff_B_MJXpMlSz8_0;
	wire w_dff_B_lVtnwA7P9_0;
	wire w_dff_B_q54FTbbG2_0;
	wire w_dff_B_LEZjdAOF2_0;
	wire w_dff_B_K5gxWMxw9_0;
	wire w_dff_B_jhGhSjXn1_0;
	wire w_dff_B_XXn0nBBT4_0;
	wire w_dff_B_8XvexMbO0_0;
	wire w_dff_B_k5ROGEeQ9_0;
	wire w_dff_B_dPS8gKbJ3_0;
	wire w_dff_B_Mqwo4kXx0_0;
	wire w_dff_B_tgwF8Qzt1_0;
	wire w_dff_B_fUQ7IRTy5_0;
	wire w_dff_A_YxLnYYPV2_1;
	wire w_dff_A_wZ5mTor86_2;
	wire w_dff_B_FIoheWbs5_2;
	wire w_dff_B_IGq84fdi5_1;
	wire w_dff_B_Y32ShMuw6_1;
	wire w_dff_B_hPqcY2iD9_1;
	wire w_dff_A_3W4kvWNZ3_2;
	wire w_dff_A_nMHJbxjT1_2;
	wire w_dff_B_ZVmm8MNS6_0;
	wire w_dff_B_0A3Ro9nz0_0;
	wire w_dff_B_ep9uS0Mf1_0;
	wire w_dff_B_3aDHVfrs0_0;
	wire w_dff_B_ujgqR1BA0_0;
	wire w_dff_B_Lpe4bac67_0;
	wire w_dff_B_qqefWXnl8_0;
	wire w_dff_B_2YvTkKCA9_0;
	wire w_dff_B_kWAgN8za5_0;
	wire w_dff_B_h2W2eMv27_0;
	wire w_dff_B_eYQWpjpO9_0;
	wire w_dff_B_u2gv6qbn2_0;
	wire w_dff_B_65GFBJ5i0_0;
	wire w_dff_B_1S2oHxRv6_0;
	wire w_dff_B_n4Z3kC0B8_0;
	wire w_dff_B_69LkdRe29_0;
	wire w_dff_B_BFLz6QQE7_1;
	wire w_dff_B_WEtm194H6_0;
	wire w_dff_B_7IBwxlQT2_0;
	wire w_dff_B_HnBuq4GM7_0;
	wire w_dff_B_j0gK1YOY6_0;
	wire w_dff_B_817Q2Pqi5_0;
	wire w_dff_B_J9CF1wra9_0;
	wire w_dff_B_rC1cw62D8_0;
	wire w_dff_B_xWmwhYEu5_0;
	wire w_dff_B_NAUXOCim6_0;
	wire w_dff_B_NeoQELkz9_0;
	wire w_dff_B_nsN7kUO77_0;
	wire w_dff_B_Fo0Afh4i9_0;
	wire w_dff_B_44vAecWO2_0;
	wire w_dff_B_jYDj2gId5_0;
	wire w_dff_A_sc3jI8Q69_0;
	wire w_dff_A_ojvfwOxf9_0;
	wire w_dff_A_RUcvG7n60_0;
	wire w_dff_A_ax7OvO1A0_1;
	wire w_dff_A_1tEDy0cf0_1;
	wire w_dff_A_By1RKrdX8_1;
	wire w_dff_A_DC7nCXXN2_1;
	wire w_dff_A_sjV8SmEY9_1;
	wire w_dff_A_eihDuhsQ7_1;
	wire w_dff_A_ex2SzdNi7_1;
	wire w_dff_A_xXCSNQrE9_0;
	wire w_dff_A_NbS7Alik6_0;
	wire w_dff_A_FPGa4Tmv5_0;
	wire w_dff_A_4mEEVqk35_0;
	wire w_dff_A_BNuCiqWE6_0;
	wire w_dff_A_gyXkKqaX3_1;
	wire w_dff_A_0fZTBHr02_1;
	wire w_dff_A_If7SqYPf4_1;
	wire w_dff_A_9DpGzOIF8_1;
	wire w_dff_A_mKOuAFjK0_1;
	wire w_dff_A_L7SHkB7f7_1;
	wire w_dff_A_NmeBqJej4_1;
	wire w_dff_B_DqTLLdrs8_0;
	wire w_dff_B_Hg05mqed6_0;
	wire w_dff_B_4C7GlDBG1_0;
	wire w_dff_B_O1iGWmKO3_0;
	wire w_dff_B_uIzJ5YwN7_0;
	wire w_dff_B_DWi30R3v4_0;
	wire w_dff_B_DzHoF0Ho2_0;
	wire w_dff_B_6vc9JUTF5_0;
	wire w_dff_B_ipExecNx7_0;
	wire w_dff_B_IGY9THnU3_0;
	wire w_dff_B_dvbZwwhr3_0;
	wire w_dff_B_0gPtaQdm0_0;
	wire w_dff_B_u5p460Ly0_0;
	wire w_dff_B_vv2nfHoo5_1;
	wire w_dff_A_Z1lAP6kb0_2;
	wire w_dff_A_OZ82CCvQ3_2;
	wire w_dff_A_snODAuqc6_2;
	wire w_dff_B_q1kALwgv4_0;
	wire w_dff_B_Akr5dmJX1_0;
	wire w_dff_B_voAJ6e0B4_0;
	wire w_dff_B_LbmON4d04_0;
	wire w_dff_B_czf60rpt0_0;
	wire w_dff_B_OtENGNYd1_0;
	wire w_dff_B_6pjDQfW88_0;
	wire w_dff_B_nIM3frMz3_0;
	wire w_dff_B_sumYEOPg6_0;
	wire w_dff_B_wKto22uR8_0;
	wire w_dff_B_83oAMUNY6_0;
	wire w_dff_B_0ovZIQyE8_0;
	wire w_dff_B_DHFhcBXc5_0;
	wire w_dff_B_sFCOBFKZ8_0;
	wire w_dff_A_YrGfyymj5_0;
	wire w_dff_A_gamMfp6T9_0;
	wire w_dff_A_iXDsf0Av2_1;
	wire w_dff_B_d44rBEZQ4_1;
	wire w_dff_B_hLhYhoOa3_1;
	wire w_dff_B_Kq7EokUD6_1;
	wire w_dff_B_nSl6TPh82_1;
	wire w_dff_B_dWZPMxOD5_1;
	wire w_dff_B_vhe6go5h3_1;
	wire w_dff_B_VPO1xM0b1_1;
	wire w_dff_B_xl4fjvn14_1;
	wire w_dff_B_prMlvip00_1;
	wire w_dff_B_lB19PUY14_1;
	wire w_dff_B_fW7CWBUT3_1;
	wire w_dff_B_2bYdIWHR2_1;
	wire w_dff_B_QlE12RLM6_1;
	wire w_dff_B_lc1B8HQ97_1;
	wire w_dff_B_8HXiJ17M2_1;
	wire w_dff_B_IbNvrrdT9_1;
	wire w_dff_B_4rKzi5ft5_1;
	wire w_dff_B_hr4RBaw75_1;
	wire w_dff_B_JPTkieWH6_1;
	wire w_dff_B_JFrPKMCF7_1;
	wire w_dff_B_6bJ5mfPR9_1;
	wire w_dff_B_HLYyn1f77_1;
	wire w_dff_B_7YKmGSuK7_1;
	wire w_dff_B_7lvApMHE8_1;
	wire w_dff_B_ONpsITEh0_1;
	wire w_dff_B_9P3iOI6n7_1;
	wire w_dff_B_RWnyobUg6_1;
	wire w_dff_B_KZoARXLc0_1;
	wire w_dff_B_FqkfDwMg0_1;
	wire w_dff_B_IDc6rDxQ2_1;
	wire w_dff_B_URZBSOEB9_1;
	wire w_dff_B_mgwEUQS91_1;
	wire w_dff_B_sRWC0tdv5_1;
	wire w_dff_B_dzFlQmzL4_1;
	wire w_dff_B_tuaV0hrY5_1;
	wire w_dff_B_j17Q7vPS0_1;
	wire w_dff_B_Li0bAqfx2_1;
	wire w_dff_B_4DN8KS018_1;
	wire w_dff_B_T3Kapml73_1;
	wire w_dff_B_H7MzAnXL8_1;
	wire w_dff_B_erHClltW3_1;
	wire w_dff_B_VRr48Sni9_1;
	wire w_dff_B_GjJOhlnr9_1;
	wire w_dff_B_YaNA41sQ1_1;
	wire w_dff_B_cuEdzt2S1_0;
	wire w_dff_B_LPgtyoLW5_0;
	wire w_dff_B_uYNAnF3P9_0;
	wire w_dff_B_TTI3V0c07_0;
	wire w_dff_B_0LeQCjqX9_0;
	wire w_dff_B_hGo6aE1L4_0;
	wire w_dff_B_vrHzVBPs5_1;
	wire w_dff_B_8P1YGzgQ2_1;
	wire w_dff_B_Quo6qYtP7_1;
	wire w_dff_B_oUcrpXRb4_1;
	wire w_dff_B_vAZPEblA7_1;
	wire w_dff_B_iQPIcCBI1_1;
	wire w_dff_B_qwPBKtuU9_1;
	wire w_dff_B_7ursiyCr0_1;
	wire w_dff_B_9EyVRvmn8_1;
	wire w_dff_B_DUiIQvWy4_1;
	wire w_dff_B_WTgw8wve6_1;
	wire w_dff_B_7O6ie4Ck9_1;
	wire w_dff_B_Ni0PLMRt2_1;
	wire w_dff_B_VfuJOKvu7_1;
	wire w_dff_B_ujPWr6ve6_1;
	wire w_dff_B_rbAuemPE9_1;
	wire w_dff_B_3TGk4T0w7_1;
	wire w_dff_B_ZBum0YOh9_1;
	wire w_dff_B_mRm8lSLm3_1;
	wire w_dff_B_FXetr5Jf8_0;
	wire w_dff_B_bj1sZqhK9_0;
	wire w_dff_B_ZzupltTq5_0;
	wire w_dff_B_RCQ0KC3s0_0;
	wire w_dff_B_PbjgCsSE0_0;
	wire w_dff_B_ZIzc92Bh0_0;
	wire w_dff_B_AKBIMfoM4_1;
	wire w_dff_B_VkR0RJnO3_1;
	wire w_dff_B_YoXDgICp1_1;
	wire w_dff_B_7UNUH5rp2_1;
	wire w_dff_B_o2AF7ZD13_2;
	wire w_dff_B_kgOnxlfu9_2;
	wire w_dff_B_O2epEFNI8_2;
	wire w_dff_B_zdIME7Wv5_0;
	wire w_dff_B_0t4XAYSf0_0;
	wire w_dff_B_kdRm8gLu1_0;
	wire w_dff_B_M5D640MM2_0;
	wire w_dff_B_TnHaRBC44_0;
	wire w_dff_B_2hFp0IYO8_0;
	wire w_dff_B_D4dwODuW2_0;
	wire w_dff_B_bUX2u2H59_0;
	wire w_dff_B_9KqjEjrP8_0;
	wire w_dff_B_7o2KHG086_0;
	wire w_dff_B_oQ8gKiWd9_0;
	wire w_dff_B_9vShPgtL7_0;
	wire w_dff_B_iKYzvaD16_0;
	wire w_dff_B_SJjDmDZT6_2;
	wire w_dff_B_bsAacwTI8_2;
	wire w_dff_B_K9zwZyi23_2;
	wire w_dff_B_metFiBlD4_0;
	wire w_dff_B_XEBaaWNY0_1;
	wire w_dff_B_cWW7BqkY5_1;
	wire w_dff_B_FT55muRm4_1;
	wire w_dff_B_P2bFHe5K8_1;
	wire w_dff_B_4UIEkQYb6_1;
	wire w_dff_B_VwpLRZYF3_1;
	wire w_dff_B_GtsUyFiA0_0;
	wire w_dff_B_S49bTiMW9_0;
	wire w_dff_B_RLUsb3Cv4_1;
	wire w_dff_B_z12meKbH6_1;
	wire w_dff_A_0VM845kW6_0;
	wire w_dff_A_EsAjOgU65_0;
	wire w_dff_B_eJ69Mfy49_1;
	wire w_dff_B_uLwGAIUX9_1;
	wire w_dff_B_PS2S0xBY7_1;
	wire w_dff_A_npS2ivQk8_0;
	wire w_dff_A_IqrBrl157_1;
	wire w_dff_A_U4fR8iQ06_1;
	wire w_dff_A_2xgFELTQ7_1;
	wire w_dff_A_tGcLAQFM9_1;
	wire w_dff_A_CX0tG5144_1;
	wire w_dff_A_6u7w5u6X9_1;
	wire w_dff_B_tlusE0j86_1;
	wire w_dff_B_sWwHpGJt0_1;
	wire w_dff_B_GuCnLKnr4_1;
	wire w_dff_B_4J9ddOpI5_1;
	wire w_dff_B_HlcYQuNT3_1;
	wire w_dff_B_c1L8sULW9_1;
	wire w_dff_B_p49FRbal8_1;
	wire w_dff_B_ZbyInzDL9_1;
	wire w_dff_B_iVd2sr9e1_0;
	wire w_dff_B_yRqSM7OQ3_0;
	wire w_dff_B_LoDdlt7O8_0;
	wire w_dff_B_HGmizWoM4_0;
	wire w_dff_B_oZOwAB332_1;
	wire w_dff_B_hamSiRHx7_1;
	wire w_dff_B_5IjkzF0r0_0;
	wire w_dff_B_7wNVapkp3_0;
	wire w_dff_B_kJmmPrrk2_0;
	wire w_dff_B_vFdVfgzK6_0;
	wire w_dff_A_B0xsdXZn9_0;
	wire w_dff_A_OTKIU66v7_0;
	wire w_dff_A_YV5OdHI91_0;
	wire w_dff_A_PPiBdDlg1_0;
	wire w_dff_A_xrLt9rQJ6_0;
	wire w_dff_A_TwveDcUk1_0;
	wire w_dff_A_YM1cTB718_0;
	wire w_dff_A_5cmZxVG40_0;
	wire w_dff_A_9W5ELkMv7_0;
	wire w_dff_A_xhrFUx5g6_0;
	wire w_dff_A_K8kkhlAe6_2;
	wire w_dff_A_dO3Ntust9_2;
	wire w_dff_A_2hM6Ucfa7_2;
	wire w_dff_B_tGjzBN9i0_1;
	wire w_dff_B_NJuNj2kG9_1;
	wire w_dff_A_NnsPrOqX9_1;
	wire w_dff_A_qQP3m4jI7_1;
	wire w_dff_A_0NMZDrI95_1;
	wire w_dff_A_gGGJZbzA5_1;
	wire w_dff_A_GGM1gy4q7_2;
	wire w_dff_A_D9Wcx2QM8_0;
	wire w_dff_A_vfZVX75W4_0;
	wire w_dff_A_bdDwh1Wl4_1;
	wire w_dff_A_Jw5QYtyr4_1;
	wire w_dff_B_CUT3gRE58_0;
	wire w_dff_B_bWLS9a6V2_0;
	wire w_dff_B_vI2VsaJz9_0;
	wire w_dff_B_zGKyLPLR5_0;
	wire w_dff_B_0XECho6T1_0;
	wire w_dff_B_0ZMRQjxo5_0;
	wire w_dff_B_Ce7ze7A05_0;
	wire w_dff_B_04LfTljs7_0;
	wire w_dff_B_5FLfSNxX5_0;
	wire w_dff_B_E4IgnFj56_0;
	wire w_dff_B_0spYFI720_0;
	wire w_dff_B_0FbXlvoh7_0;
	wire w_dff_B_kwmSNrEv6_0;
	wire w_dff_B_8AGxI0Mu5_2;
	wire w_dff_B_ASVoifaa9_2;
	wire w_dff_B_Ajmd820Z0_2;
	wire w_dff_B_EFBbqyKg0_1;
	wire w_dff_B_NuMGKBgK4_1;
	wire w_dff_B_fIKJ2Mgp5_1;
	wire w_dff_B_d4z54aPe4_1;
	wire w_dff_B_MylFQXjh9_1;
	wire w_dff_B_hWOXd6XA6_1;
	wire w_dff_B_Periazxo7_1;
	wire w_dff_B_9P4ED7zy1_1;
	wire w_dff_B_U8M86RnQ3_0;
	wire w_dff_B_gBzeg0a72_0;
	wire w_dff_B_I1dON0uH7_0;
	wire w_dff_B_ugITFTmU9_1;
	wire w_dff_B_ybO4WRJc4_1;
	wire w_dff_B_8U0Oim1p9_1;
	wire w_dff_B_l6Ij8nIr3_1;
	wire w_dff_B_CG8aC8g90_1;
	wire w_dff_B_onHZEBtR5_1;
	wire w_dff_B_B3Sll7g45_1;
	wire w_dff_B_HHaPyPg73_1;
	wire w_dff_B_fieNrXQD7_1;
	wire w_dff_B_BFd0Oyoi6_1;
	wire w_dff_B_Pg0Xh79Q8_1;
	wire w_dff_B_8rQ7rliv3_1;
	wire w_dff_B_LxXzK1Q48_1;
	wire w_dff_B_OEziAhiQ8_1;
	wire w_dff_B_sStGSEa44_1;
	wire w_dff_A_SwyMxSwn5_0;
	wire w_dff_A_K1FPsr598_0;
	wire w_dff_A_FL9tvQGF9_0;
	wire w_dff_A_yezpWkaN3_0;
	wire w_dff_A_3lqhmAhK7_0;
	wire w_dff_B_90WGFX200_1;
	wire w_dff_B_WTvEmP2Q3_1;
	wire w_dff_B_gCPz57zM4_1;
	wire w_dff_B_7640OupI3_1;
	wire w_dff_B_RnR6lCWr1_0;
	wire w_dff_B_bk9oqwj17_0;
	wire w_dff_B_zjR3F0PZ6_0;
	wire w_dff_B_uAVllWra0_0;
	wire w_dff_B_RU9gjels2_0;
	wire w_dff_B_vNbCm1wf4_0;
	wire w_dff_B_sczV63Oz7_0;
	wire w_dff_B_TU8pH5Wq5_0;
	wire w_dff_B_pA0nuJHF3_0;
	wire w_dff_B_iecZB5iN5_0;
	wire w_dff_B_EaveTiGR9_0;
	wire w_dff_B_I7cht51M1_0;
	wire w_dff_B_MEIhhaKH4_0;
	wire w_dff_B_l83lBKCX4_0;
	wire w_dff_B_ZI5yvDHv8_2;
	wire w_dff_B_BiHPPjJQ1_2;
	wire w_dff_B_t5CF08rg6_2;
	wire w_dff_B_UXzmJdT80_1;
	wire w_dff_B_gGE7O5iU9_1;
	wire w_dff_B_hU0SneQp0_1;
	wire w_dff_B_VzT1cfgR9_1;
	wire w_dff_B_I7I4M44f4_1;
	wire w_dff_B_3lXXAADx3_1;
	wire w_dff_B_GTMGHZwB8_1;
	wire w_dff_B_c9O17rgw7_1;
	wire w_dff_B_Ej5h7qih9_0;
	wire w_dff_B_KpAM97bC1_0;
	wire w_dff_B_h8VxbfjI7_0;
	wire w_dff_B_wazcHJKO4_0;
	wire w_dff_B_Ib7fXhQc1_1;
	wire w_dff_B_kZQ8zMyd6_1;
	wire w_dff_A_rNiPtXLH8_2;
	wire w_dff_A_3aedCEev1_2;
	wire w_dff_A_QMPVijS82_2;
	wire w_dff_A_GZeO6MGe9_0;
	wire w_dff_A_0WMH8yzG8_0;
	wire w_dff_A_cdAeYYAu1_0;
	wire w_dff_A_bIIZgxBS9_0;
	wire w_dff_A_Pp1HGQRd6_0;
	wire w_dff_A_za0xKMAC7_1;
	wire w_dff_A_7WVyANtA8_2;
	wire w_dff_A_Yv7YRBAz8_2;
	wire w_dff_B_u4wgZrrl9_1;
	wire w_dff_B_e7Aq2xOM1_1;
	wire w_dff_A_0V2656ta9_0;
	wire w_dff_A_QiqEtPaT6_0;
	wire w_dff_A_LWUS1reT6_1;
	wire w_dff_B_l3iQHOaA7_1;
	wire w_dff_B_2JDzgvY80_1;
	wire w_dff_B_X9qMtqnv1_1;
	wire w_dff_B_Y1iIcmNt6_1;
	wire w_dff_B_0f47Wv3m5_1;
	wire w_dff_B_At1YA5Vh4_1;
	wire w_dff_B_lJZSXHvj7_1;
	wire w_dff_B_m1rdW9ar1_1;
	wire w_dff_B_BQ2EQVOl9_1;
	wire w_dff_B_1iNS7Nap6_0;
	wire w_dff_B_eMTh1SQH4_0;
	wire w_dff_B_SXzXfOxQ5_0;
	wire w_dff_B_LDLs90Uk8_0;
	wire w_dff_B_heqfmxww4_0;
	wire w_dff_B_G225qpP34_0;
	wire w_dff_B_Sq3v5Xdh4_1;
	wire w_dff_A_9JjDmRhG0_0;
	wire w_dff_A_7TidQJ6G5_1;
	wire w_dff_A_Q62aijYp6_0;
	wire w_dff_A_QcqzsMkw0_2;
	wire w_dff_A_QegbFgMH0_1;
	wire w_dff_A_fI6T211y3_2;
	wire w_dff_A_ORZgCVlI8_0;
	wire w_dff_A_7suQ0XYU3_0;
	wire w_dff_A_hAkS5YAw9_0;
	wire w_dff_A_d6GDjhyS9_0;
	wire w_dff_A_97sd9oJa1_0;
	wire w_dff_A_7ThD62w13_0;
	wire w_dff_A_V7JhJi4I3_0;
	wire w_dff_A_crg4mZyX4_1;
	wire w_dff_A_Xx2je7Ng9_1;
	wire w_dff_A_segWPjME5_2;
	wire w_dff_A_yIPwBlnh7_2;
	wire w_dff_A_dJn9XU4r0_2;
	wire w_dff_A_J9WMtu723_2;
	wire w_dff_A_eCToI8218_2;
	wire w_dff_B_gMSfxgK16_3;
	wire w_dff_B_KcNeIWmv8_3;
	wire w_dff_A_1TDZkw5D4_0;
	wire w_dff_A_UmKYnHNg0_0;
	wire w_dff_A_AlWs86Wg8_0;
	wire w_dff_A_vWLEkGRQ2_0;
	wire w_dff_A_dzVduUWR0_2;
	wire w_dff_A_PWGx2d8f6_2;
	wire w_dff_A_a58CEpQU8_2;
	wire w_dff_B_mjLra52h0_1;
	wire w_dff_B_4LVBH2It6_1;
	wire w_dff_B_SJTCTUpE8_1;
	wire w_dff_B_0pq8b4099_1;
	wire w_dff_B_wP0WAYa06_1;
	wire w_dff_B_FfW8U1v00_1;
	wire w_dff_B_dw0eGgNd5_1;
	wire w_dff_B_BDi1Z0Wg1_1;
	wire w_dff_B_NK9pg6376_1;
	wire w_dff_B_gxIe1wTu2_1;
	wire w_dff_B_jhc8k3IX3_1;
	wire w_dff_B_yS83qBjv9_1;
	wire w_dff_B_JIjnueRV8_1;
	wire w_dff_B_262O5ZM97_1;
	wire w_dff_B_h34gSi9m2_1;
	wire w_dff_B_wujcZsIp8_1;
	wire w_dff_B_rzkQElNl3_1;
	wire w_dff_B_YehUqUFZ2_1;
	wire w_dff_B_yPIn38pH5_1;
	wire w_dff_B_IR1js6PY9_1;
	wire w_dff_B_p01T7xu26_1;
	wire w_dff_B_x2B1v9ul5_1;
	wire w_dff_B_9XDQ9MuK2_1;
	wire w_dff_B_6rxE4lJ27_1;
	wire w_dff_B_S5HSk2m91_1;
	wire w_dff_B_fBrT7Hht7_1;
	wire w_dff_B_LbGTneuH2_1;
	wire w_dff_B_TSoGnU751_1;
	wire w_dff_B_giGWtHgu2_1;
	wire w_dff_B_AcWpHut54_1;
	wire w_dff_B_Y2q2okYk1_0;
	wire w_dff_B_pma8W6UL3_0;
	wire w_dff_B_jifYEoLa5_0;
	wire w_dff_B_ZEnctCti8_0;
	wire w_dff_B_EmH8pxP01_0;
	wire w_dff_B_Naal926N0_0;
	wire w_dff_B_q67KMKMI6_0;
	wire w_dff_B_Gmtzc4x55_0;
	wire w_dff_B_gWjX512N1_0;
	wire w_dff_B_9K9OXY3N2_0;
	wire w_dff_B_HwYRXSb17_0;
	wire w_dff_B_8KOJ0rAh4_0;
	wire w_dff_B_aGH9xiGJ4_0;
	wire w_dff_B_oL3F66b33_0;
	wire w_dff_B_FuoDS0bO8_0;
	wire w_dff_B_REvoa9Uk5_0;
	wire w_dff_B_t6pHtrQy5_1;
	wire w_dff_B_dDzzxKxE0_1;
	wire w_dff_B_eTcQlCR77_1;
	wire w_dff_B_Txjh1bF79_1;
	wire w_dff_B_EEK85wo98_1;
	wire w_dff_B_e6rApPUh7_1;
	wire w_dff_B_0OOP1XMK4_1;
	wire w_dff_B_utxupP6v0_1;
	wire w_dff_B_fkywhnmy6_1;
	wire w_dff_A_qAfsH6ps1_0;
	wire w_dff_A_ka0Af7gB1_0;
	wire w_dff_A_Y7VtoUEM8_0;
	wire w_dff_A_vXaZmONx2_0;
	wire w_dff_A_3u8AhDZ50_0;
	wire w_dff_A_CBmTJGOR5_0;
	wire w_dff_A_2n1SrRKC7_0;
	wire w_dff_A_FdbRZcal4_0;
	wire w_dff_A_XpKbW4934_0;
	wire w_dff_A_WAbi9woj3_0;
	wire w_dff_A_q0KUU9WO9_0;
	wire w_dff_B_1JrkY8Dv8_2;
	wire w_dff_B_Ozu4KnEC0_2;
	wire w_dff_B_llg6wm2I2_2;
	wire w_dff_B_nGukN8y83_2;
	wire w_dff_B_eBuerXZk9_2;
	wire w_dff_A_yY3htEE00_0;
	wire w_dff_A_Spe8grpu6_1;
	wire w_dff_A_ce82iF9C0_2;
	wire w_dff_A_bqmsRlfN6_2;
	wire w_dff_A_iymLysLC7_2;
	wire w_dff_A_nRGnI5Q08_2;
	wire w_dff_A_faYPsANX9_0;
	wire w_dff_A_IL6xpjDa7_0;
	wire w_dff_A_Q6I6sg426_0;
	wire w_dff_A_2ESL2CEo6_0;
	wire w_dff_A_ZDO7B8j88_0;
	wire w_dff_A_zyAtjveW0_0;
	wire w_dff_A_VihzxTqh9_0;
	wire w_dff_A_l1TPZ3Kj2_0;
	wire w_dff_A_zOHvRT210_0;
	wire w_dff_A_kjwlrNqP9_0;
	wire w_dff_A_HFFMZKXC4_0;
	wire w_dff_B_2ODW0byy4_1;
	wire w_dff_B_bR5wdcvE0_1;
	wire w_dff_B_YCh1T0KM1_1;
	wire w_dff_B_WLeseU1z1_1;
	wire w_dff_B_GBcMuDia6_1;
	wire w_dff_B_9WsjWPI97_0;
	wire w_dff_B_PoXP9G9H8_0;
	wire w_dff_B_LH6zC8nH4_0;
	wire w_dff_B_N5kgZ4q98_0;
	wire w_dff_B_tam88bC02_0;
	wire w_dff_A_JmBuoIrZ9_0;
	wire w_dff_A_FtQ5RHRX1_0;
	wire w_dff_B_lwgdiKd39_0;
	wire w_dff_B_Qa0kXc944_1;
	wire w_dff_B_gv7JNX2u5_1;
	wire w_dff_B_ArBKaFRb0_1;
	wire w_dff_B_GgwDVmIk2_0;
	wire w_dff_B_xLQe94xi2_1;
	wire w_dff_B_Y91lCFsy5_0;
	wire w_dff_B_UpMQVbjd6_1;
	wire w_dff_B_jaZ47cMA7_1;
	wire w_dff_B_7xINs6mG3_1;
	wire w_dff_B_Y2yoSY4w4_0;
	wire w_dff_B_jOxmupOZ6_0;
	wire w_dff_B_yrPwA8uG8_0;
	wire w_dff_B_kSKAt8eF0_0;
	wire w_dff_B_HIzuN37p7_1;
	wire w_dff_A_J483ghBZ3_0;
	wire w_dff_A_R1I8Dhts8_0;
	wire w_dff_A_bXDUOtni8_0;
	wire w_dff_A_lTOzkCx56_0;
	wire w_dff_B_Lkz0kzL29_1;
	wire w_dff_B_FTZIdq6L0_1;
	wire w_dff_B_WMbiIHUO3_1;
	wire w_dff_B_1GSiAlF65_1;
	wire w_dff_B_KzVdmX5f1_1;
	wire w_dff_B_Eh8xcU5w1_1;
	wire w_dff_B_R6OPvu1m6_1;
	wire w_dff_B_tO5YvwMX9_1;
	wire w_dff_B_xTqVdMq19_1;
	wire w_dff_B_Yn23Ap934_1;
	wire w_dff_B_OUA70wuN8_1;
	wire w_dff_B_CHoghGGr2_1;
	wire w_dff_B_sRwG79PK9_1;
	wire w_dff_B_d0vPN1jU2_1;
	wire w_dff_B_XgTP2XRT7_1;
	wire w_dff_B_xF71wDdE2_1;
	wire w_dff_B_vUmjxWLO5_1;
	wire w_dff_B_Qv13RY871_1;
	wire w_dff_B_WLoJdSsh8_1;
	wire w_dff_B_blNbS6wX1_1;
	wire w_dff_B_Rh31UQkH5_1;
	wire w_dff_B_TT1moR132_1;
	wire w_dff_B_Ah0S6DeG2_1;
	wire w_dff_B_awItk95I5_1;
	wire w_dff_B_LVHBRYbN7_1;
	wire w_dff_B_RL3xREXt5_1;
	wire w_dff_A_bRwySmv44_2;
	wire w_dff_A_hIMjxelj8_2;
	wire w_dff_A_0YCsWJI95_2;
	wire w_dff_A_NdvFqruk6_2;
	wire w_dff_A_vBqxePfa1_2;
	wire w_dff_A_klTK2TIY7_2;
	wire w_dff_A_8gqaPvZ35_2;
	wire w_dff_A_T2fUFLh32_2;
	wire w_dff_A_eIaYIMDb1_2;
	wire w_dff_A_R2KmGRb39_2;
	wire w_dff_A_GbTFOAwC9_2;
	wire w_dff_A_Jn6agjht7_2;
	wire w_dff_A_zK74rVjF6_2;
	wire w_dff_A_WoT2ruqa0_2;
	wire w_dff_A_fgX5Exue9_2;
	wire w_dff_A_QtfeuDtX3_2;
	wire w_dff_A_NunGVhI32_2;
	wire w_dff_A_ZPlxwMdM3_2;
	wire w_dff_A_IMnj1xPy9_2;
	wire w_dff_A_5zXiPppJ4_2;
	wire w_dff_A_5VTLUQNs7_2;
	wire w_dff_A_6zJ0XKoK5_2;
	wire w_dff_A_NWM5yy8d4_2;
	wire w_dff_A_BePHHIG12_2;
	wire w_dff_A_SuyHfsP33_2;
	wire w_dff_B_WRpIyDKr5_0;
	wire w_dff_B_G6NOgQou0_0;
	wire w_dff_B_AsRt94t66_0;
	wire w_dff_B_xa0r5KoB9_0;
	wire w_dff_B_VOw4BDys5_0;
	wire w_dff_B_9tOouuU77_0;
	wire w_dff_B_GIuNXjbb3_0;
	wire w_dff_B_xoYDG25r2_0;
	wire w_dff_B_3MNhwztg4_0;
	wire w_dff_B_tooZ1f2L3_0;
	wire w_dff_B_97cH0skD7_0;
	wire w_dff_B_VZ8CXkyb1_0;
	wire w_dff_B_VFOFqvPb3_0;
	wire w_dff_B_yYWLHLHx1_0;
	wire w_dff_B_BXeoeUfm2_0;
	wire w_dff_B_G9lWqzGc2_0;
	wire w_dff_B_3VyOr7uT0_0;
	wire w_dff_B_Pdrz4BLb9_0;
	wire w_dff_B_oiuRAOfW1_0;
	wire w_dff_B_oDyragN69_0;
	wire w_dff_B_VNDVWmfp6_0;
	wire w_dff_B_ysMN1GsA7_2;
	wire w_dff_B_kPe973K11_1;
	wire w_dff_B_gFIIPHp96_1;
	wire w_dff_A_lNU0yOKL0_0;
	wire w_dff_A_5oygKVDc0_0;
	wire w_dff_A_Oj3gjdpi9_0;
	wire w_dff_A_9heJPZ8k6_0;
	wire w_dff_A_fGTiVtRK4_0;
	wire w_dff_A_nQQgaYQw0_0;
	wire w_dff_A_YLZyl7P60_0;
	wire w_dff_A_Moh6W1In2_0;
	wire w_dff_A_PMi9rjUu8_0;
	wire w_dff_A_ZKnW40b80_0;
	wire w_dff_A_Z8AzZGpY8_0;
	wire w_dff_A_gSJ0gdUE4_0;
	wire w_dff_A_YvUVRR3i0_0;
	wire w_dff_A_W1rNttzp8_0;
	wire w_dff_A_U71Wqot97_0;
	wire w_dff_A_THkQBd0N4_0;
	wire w_dff_A_sQllPZOP3_0;
	wire w_dff_A_M3Jx9hsM7_0;
	wire w_dff_A_m3CNYkjw4_0;
	wire w_dff_A_tb1vKi2D2_0;
	wire w_dff_A_ZBIkZu7l7_2;
	wire w_dff_A_6Wjp8grj5_2;
	wire w_dff_A_T3SAIYIW2_2;
	wire w_dff_A_kw7EHbiv4_2;
	wire w_dff_A_NtF6MYvO1_2;
	wire w_dff_A_6tCwbCYX8_2;
	wire w_dff_A_apcfSdi74_2;
	wire w_dff_A_ATFi6iuZ7_2;
	wire w_dff_A_xAlNmWun0_2;
	wire w_dff_A_j40pknwC0_2;
	wire w_dff_A_Ll5Z3cAM9_2;
	wire w_dff_A_xYaKMUou5_0;
	wire w_dff_A_aVDGvTBl0_0;
	wire w_dff_A_RxSHQLeR8_0;
	wire w_dff_A_Nnpg2m7N6_0;
	wire w_dff_A_Ir6YNkOk1_0;
	wire w_dff_A_bz7cpQx72_0;
	wire w_dff_A_4tC039Cp9_0;
	wire w_dff_A_3vRFSR4i9_0;
	wire w_dff_A_5vdkZwtE7_0;
	wire w_dff_A_a4OH2zoE8_0;
	wire w_dff_A_w2IaFdIS4_0;
	wire w_dff_A_XhCivb6b2_0;
	wire w_dff_A_TjHKLjft5_0;
	wire w_dff_A_CPCe5i563_0;
	wire w_dff_A_0owSNGe31_0;
	wire w_dff_A_mCWSBeBZ3_0;
	wire w_dff_A_Gop5yYRW1_0;
	wire w_dff_A_ANmvAQjt5_0;
	wire w_dff_A_EpucYBj75_0;
	wire w_dff_A_UAnolVtf5_0;
	wire w_dff_A_UL2OIh3Q1_2;
	wire w_dff_A_bHQMXbCU3_2;
	wire w_dff_A_wkO4e9Mb7_2;
	wire w_dff_A_X2obzv4Q0_2;
	wire w_dff_A_5nRUB4HX9_2;
	wire w_dff_A_OYYFGldD6_2;
	wire w_dff_A_5CJESW8C2_2;
	wire w_dff_A_Z56cqX7z9_2;
	wire w_dff_A_4nEIVHXF1_2;
	wire w_dff_A_6X6eDHsP7_2;
	wire w_dff_A_NJJxwybQ5_2;
	wire w_dff_A_HPTCquTi3_2;
	wire w_dff_A_xCSFowHo3_2;
	wire w_dff_A_ycHHp8f25_2;
	wire w_dff_B_ib0tolKH8_0;
	wire w_dff_B_ZHJTGL6T5_0;
	wire w_dff_B_rrzrgDyO1_0;
	wire w_dff_B_rZKLo1xI4_0;
	wire w_dff_B_HgiEKKdQ0_0;
	wire w_dff_B_ze0IZd1g9_0;
	wire w_dff_B_nr8ZFi4z4_0;
	wire w_dff_B_f3FXnLPP7_0;
	wire w_dff_B_UEjY8Sqi8_0;
	wire w_dff_B_CZsidcyL3_0;
	wire w_dff_B_KwH0vJ9X5_0;
	wire w_dff_B_jK4BFWzy9_0;
	wire w_dff_B_xRRWSQSy0_0;
	wire w_dff_B_zDEEEJlf7_0;
	wire w_dff_B_xj7QYRbn9_0;
	wire w_dff_B_sE56QogI2_0;
	wire w_dff_B_iMDAzPsU1_0;
	wire w_dff_B_2tifSvW78_0;
	wire w_dff_B_ydx6ld577_0;
	wire w_dff_B_EGaddTYu8_0;
	wire w_dff_B_L6RmGUHe6_1;
	wire w_dff_B_humdkuXK2_1;
	wire w_dff_A_BU7ua3pb8_1;
	wire w_dff_A_NzWahemj5_1;
	wire w_dff_A_5hpZymzW3_1;
	wire w_dff_A_50tdOzGC6_1;
	wire w_dff_A_NCM9XFF52_1;
	wire w_dff_A_jOjA4B3G5_1;
	wire w_dff_A_t6JmLTNz6_1;
	wire w_dff_A_CL7LuoBa3_1;
	wire w_dff_A_E07EwdgE8_1;
	wire w_dff_A_l26b1K5J8_1;
	wire w_dff_A_X8EoCYOa1_1;
	wire w_dff_A_Bfwzorlg8_1;
	wire w_dff_A_7dZYS9B62_1;
	wire w_dff_A_eJL18UmO4_1;
	wire w_dff_A_i4rtBFi63_1;
	wire w_dff_A_x9mLeMmb5_1;
	wire w_dff_A_AprcE3Le9_1;
	wire w_dff_A_vENDE7u71_1;
	wire w_dff_A_a30Dc9h31_1;
	wire w_dff_A_nERkjmNx0_1;
	wire w_dff_A_2B9x6Pbt1_1;
	wire w_dff_A_E1ohL8k44_1;
	wire w_dff_A_CDMp4Ikt7_1;
	wire w_dff_A_QRTRrZUQ5_1;
	wire w_dff_A_1TQ1Sbgq5_1;
	wire w_dff_A_0yJBJbhp4_1;
	wire w_dff_A_RpM7D0SV8_1;
	wire w_dff_A_fpNWQqcX6_1;
	wire w_dff_A_DnYYmT1e8_1;
	wire w_dff_A_9fTUwbFM1_1;
	wire w_dff_A_NkOUE4QV9_1;
	wire w_dff_A_KCDM5riV0_1;
	wire w_dff_A_iveCsrqg5_1;
	wire w_dff_A_enNOYNb38_1;
	wire w_dff_A_MW1Bc9OL0_1;
	wire w_dff_A_0cPIuAtG6_1;
	wire w_dff_A_qmWfOSdh2_1;
	wire w_dff_A_cevV5e9A0_1;
	wire w_dff_B_Kgrl6t8O0_0;
	wire w_dff_B_DLZeU8Xl6_0;
	wire w_dff_B_sMp9HhWS2_0;
	wire w_dff_B_g9U9IYyX3_0;
	wire w_dff_B_YwCy8oZN3_0;
	wire w_dff_B_wMXNHpyY5_0;
	wire w_dff_B_Sx8LJqTa0_0;
	wire w_dff_B_Ffcd17VR9_0;
	wire w_dff_B_IH7fL4Nm9_0;
	wire w_dff_B_IpeAaenE6_0;
	wire w_dff_B_7BFlbH6r1_0;
	wire w_dff_B_kBY2X3PQ8_0;
	wire w_dff_B_dZxcuT3S9_0;
	wire w_dff_B_pjaLm7MK4_0;
	wire w_dff_B_42xHG2kJ5_0;
	wire w_dff_B_UydGTAgU1_0;
	wire w_dff_B_c9vALxBW9_0;
	wire w_dff_B_JhodgRi09_0;
	wire w_dff_B_MLLz04vA7_0;
	wire w_dff_B_TSdQhI3G0_0;
	wire w_dff_B_IzLWxCMd6_1;
	wire w_dff_A_4tE30Vwy7_2;
	wire w_dff_B_vSewMB1y0_0;
	wire w_dff_B_K9I4zaTN6_0;
	wire w_dff_B_o2NWN9GO7_0;
	wire w_dff_B_vmfxdA4W9_0;
	wire w_dff_B_cbtK9TAa6_0;
	wire w_dff_B_7hdcCF510_0;
	wire w_dff_B_MnZpJsH21_0;
	wire w_dff_B_GLoHxRd08_0;
	wire w_dff_B_o5P7f0169_0;
	wire w_dff_B_A2ZDyqOk5_0;
	wire w_dff_B_hmoUdjim9_0;
	wire w_dff_B_H7AUu1EA1_0;
	wire w_dff_B_O1AictfI4_0;
	wire w_dff_B_HoPAZZOw6_0;
	wire w_dff_B_EcNXww7o1_0;
	wire w_dff_B_q3PBkS4d2_0;
	wire w_dff_B_Fbl7Xien0_0;
	wire w_dff_B_qn5bWogX8_0;
	wire w_dff_B_aZcDLtDG6_0;
	wire w_dff_B_Jq7OWrXU8_1;
	wire w_dff_B_ovKHhbdz1_1;
	wire w_dff_B_Q8ABeuZd7_1;
	wire w_dff_A_ki0ASF4M8_0;
	wire w_dff_A_lFomooOb5_0;
	wire w_dff_A_ZrhT11cM2_0;
	wire w_dff_A_3gcMCGJO1_0;
	wire w_dff_A_WwunhunA1_0;
	wire w_dff_A_NbYHYZhP2_0;
	wire w_dff_A_Ubr6QMM37_0;
	wire w_dff_A_KlvC5Bed3_0;
	wire w_dff_A_bpKVYhvG2_0;
	wire w_dff_A_14KvqGfs6_0;
	wire w_dff_A_dugp3Xvq2_0;
	wire w_dff_A_EfMp3gX20_0;
	wire w_dff_A_GSPtApM15_0;
	wire w_dff_A_sxe1NpZs7_0;
	wire w_dff_A_pw6QaPsH7_0;
	wire w_dff_A_QLx6BECE6_0;
	wire w_dff_A_jMObl2In7_0;
	wire w_dff_A_58dpKpKG9_0;
	wire w_dff_A_7j2i70Da2_2;
	wire w_dff_A_5saTnAlU9_2;
	wire w_dff_A_wOJZlyW08_2;
	wire w_dff_A_rW2uadle0_2;
	wire w_dff_A_QeePR53M7_2;
	wire w_dff_A_tXPiKJdB2_2;
	wire w_dff_A_HUASIeDg1_2;
	wire w_dff_A_3iIQOlkU6_2;
	wire w_dff_A_FKKUxtHb1_2;
	wire w_dff_A_BeAran7r8_2;
	wire w_dff_A_mnwn4CYJ5_2;
	wire w_dff_A_wmHjxtnJ2_2;
	wire w_dff_A_tTGgUwVC5_2;
	wire w_dff_A_0k1q2xTD9_2;
	wire w_dff_A_778z624G2_2;
	wire w_dff_A_HUKVj8fA4_2;
	wire w_dff_A_K6Iq2SXH5_2;
	wire w_dff_A_rh61vUaI2_2;
	wire w_dff_A_vwgUazEv3_2;
	wire w_dff_A_q0V7oPRS2_0;
	wire w_dff_A_JTX3UDzV4_0;
	wire w_dff_A_Iyijq3FQ7_0;
	wire w_dff_A_1kc3LsSs4_0;
	wire w_dff_A_itu51oVY4_0;
	wire w_dff_A_s6sk633O5_0;
	wire w_dff_A_VOyMETQt6_0;
	wire w_dff_A_R8iQ81MI1_0;
	wire w_dff_A_nqY2Uh666_0;
	wire w_dff_A_Z4VBhC2g9_0;
	wire w_dff_A_EGko19t43_0;
	wire w_dff_A_iT981qWw0_0;
	wire w_dff_A_xPFvLJPM0_0;
	wire w_dff_A_RBKwFwSC2_0;
	wire w_dff_A_PifznpmR9_0;
	wire w_dff_A_THl7v3H99_0;
	wire w_dff_A_jVEqA2kz8_0;
	wire w_dff_A_Jz1nKuwT1_2;
	wire w_dff_A_ZKftlHUA6_2;
	wire w_dff_A_QpGET3A94_2;
	wire w_dff_A_dpVnm63O7_2;
	wire w_dff_A_iBsoTUgp3_2;
	wire w_dff_A_pwfpBjgA7_2;
	wire w_dff_A_2heLTJ250_2;
	wire w_dff_A_DwYJ2Z3T6_2;
	wire w_dff_A_kL3I5mTA9_2;
	wire w_dff_A_On1pbqBq8_2;
	wire w_dff_A_4MEsVlrA7_2;
	wire w_dff_A_034kpSf43_2;
	wire w_dff_A_PVtJZn7T6_2;
	wire w_dff_A_44gbeMXv9_2;
	wire w_dff_A_u8NlSWp98_2;
	wire w_dff_A_pUhPiI5Q7_2;
	wire w_dff_A_iDITvLu20_2;
	wire w_dff_A_DWaEN6e94_2;
	wire w_dff_A_YEAViCjk5_2;
	wire w_dff_A_SBWxVdOH5_2;
	wire w_dff_B_n0JULlMa2_0;
	wire w_dff_B_6uClxzp97_0;
	wire w_dff_B_mASb81U03_0;
	wire w_dff_B_7u1vgKYg6_0;
	wire w_dff_B_6ZiCbqQd3_0;
	wire w_dff_B_DoasNh6g3_0;
	wire w_dff_B_ESwQ3rgW2_0;
	wire w_dff_B_LQ1ySkNK0_0;
	wire w_dff_B_4WIrFQMY0_0;
	wire w_dff_B_m5LPkm6d0_0;
	wire w_dff_B_nv4Y54bF1_0;
	wire w_dff_B_66LUithL5_0;
	wire w_dff_B_1Rt8GaNl3_0;
	wire w_dff_B_zPBW5Ady7_0;
	wire w_dff_B_NYOotvNJ2_0;
	wire w_dff_B_6hQY9w0h2_0;
	wire w_dff_B_ttaq4fJM2_0;
	wire w_dff_B_uSs6b6rw5_0;
	wire w_dff_B_htTGsVSt9_0;
	wire w_dff_B_pwxvlKCd3_0;
	wire w_dff_B_QHr4jZ8J4_2;
	wire w_dff_B_7nPZ3Rre2_1;
	wire w_dff_B_1fOuwH6L7_1;
	wire w_dff_A_XYqQI4tr2_1;
	wire w_dff_A_oq3zXX0C7_1;
	wire w_dff_A_6zqY6HDs9_1;
	wire w_dff_A_oOvmg0VM2_1;
	wire w_dff_A_cWTMDDHd3_1;
	wire w_dff_A_KmnruPb86_1;
	wire w_dff_A_UVi6WQcO4_1;
	wire w_dff_A_L0DHTAX51_1;
	wire w_dff_A_8fx1SEuP8_1;
	wire w_dff_A_uVTEgqv23_1;
	wire w_dff_A_pem9On199_1;
	wire w_dff_A_6PSyUXSh4_1;
	wire w_dff_A_w6WjhYjx1_1;
	wire w_dff_A_buocVb7d9_1;
	wire w_dff_A_Ewn4RtIF1_1;
	wire w_dff_A_5EtBrdRd7_1;
	wire w_dff_A_0lFLGziL8_1;
	wire w_dff_A_ZCrqRcRk6_1;
	wire w_dff_A_WPWSIian4_1;
	wire w_dff_A_d1MpCJDD3_2;
	wire w_dff_A_3pxIiuSN9_2;
	wire w_dff_A_YSWYsvqi3_2;
	wire w_dff_A_fyPmQcVm8_2;
	wire w_dff_A_trAjfuju2_2;
	wire w_dff_A_FvB1Qr9T2_2;
	wire w_dff_A_d94azWjj7_2;
	wire w_dff_A_dghaaWEf4_2;
	wire w_dff_A_sKsSBgEk9_2;
	wire w_dff_A_Zg41apJI9_2;
	wire w_dff_A_nL5LldgU1_2;
	wire w_dff_A_pYk34Idd7_2;
	wire w_dff_A_p2CFUgv18_2;
	wire w_dff_A_2VVTXPgh1_2;
	wire w_dff_A_IXYfh8WW7_2;
	wire w_dff_A_hQSBjLl80_2;
	wire w_dff_A_7U4jiEVr8_2;
	wire w_dff_A_GGkEp1kd8_2;
	wire w_dff_A_i8NayOmt2_2;
	wire w_dff_A_NG1cNPox5_2;
	wire w_dff_A_2T0YjRoR8_1;
	wire w_dff_A_ukj2lMYs3_1;
	wire w_dff_A_v3sMnOfD6_1;
	wire w_dff_A_GqDT4R8b0_1;
	wire w_dff_A_yTlniVR09_1;
	wire w_dff_A_xVptjahG8_1;
	wire w_dff_A_fXwbrHrn6_1;
	wire w_dff_A_p6MkiGPY8_1;
	wire w_dff_A_gTLj0d0T3_1;
	wire w_dff_A_ydVYs9g36_1;
	wire w_dff_A_3TXZKoFM6_1;
	wire w_dff_A_t7MkKv054_1;
	wire w_dff_A_cuEbSjxY8_1;
	wire w_dff_A_oVjjiMYT7_1;
	wire w_dff_A_TkRUub3H9_1;
	wire w_dff_A_nx9bvsxe4_1;
	wire w_dff_A_9HOC5UXP4_1;
	wire w_dff_A_WmhOFS8T7_1;
	wire w_dff_A_TBX5Mh469_1;
	wire w_dff_A_8JXtxRY97_2;
	wire w_dff_A_fEPr5yPk6_2;
	wire w_dff_A_2EIqdY9a5_2;
	wire w_dff_A_G1ybo0jX4_2;
	wire w_dff_A_OLvqYejf3_2;
	wire w_dff_A_SlkMDmm30_2;
	wire w_dff_A_RBqN83Ax1_2;
	wire w_dff_A_rIpBa0Ap7_2;
	wire w_dff_A_cNl0c7bd9_2;
	wire w_dff_A_OXGOCku81_2;
	wire w_dff_A_he3bOx2Q8_2;
	wire w_dff_A_vSTRQghL4_2;
	wire w_dff_A_Kv3cKQwf0_2;
	wire w_dff_A_qKsaUKEO2_2;
	wire w_dff_A_eDAwHI2u4_2;
	wire w_dff_A_P8UycJDD8_2;
	wire w_dff_A_QxwvuVAj4_2;
	wire w_dff_A_rNFC4wfo5_2;
	wire w_dff_A_kcw9hboA7_2;
	wire w_dff_A_RJWpgXXD6_2;
	wire w_dff_B_Tx3nH3oS8_0;
	wire w_dff_B_hgGxcLaZ2_0;
	wire w_dff_B_mbycB4hs9_0;
	wire w_dff_B_idaAs0Bw9_0;
	wire w_dff_B_XzBlgQAC4_0;
	wire w_dff_B_Q6RuIBFz3_0;
	wire w_dff_B_Q7Atw7ZZ3_0;
	wire w_dff_B_da2HRq8B2_0;
	wire w_dff_B_Y1Z1LecR4_0;
	wire w_dff_B_ijvYExa02_0;
	wire w_dff_B_dsWROEKM4_0;
	wire w_dff_B_AYDWcRqT7_0;
	wire w_dff_B_fegGlux16_0;
	wire w_dff_B_bLveDmSc6_0;
	wire w_dff_B_F7XzmOPd8_0;
	wire w_dff_B_F3T0l02s7_0;
	wire w_dff_B_Xtb5aoXD7_0;
	wire w_dff_B_4VDLMkRI1_0;
	wire w_dff_B_ESMV3WSY4_0;
	wire w_dff_B_GRzCDFLx2_0;
	wire w_dff_A_RHULBzFo7_2;
	wire w_dff_B_uaO0d8MK4_2;
	wire w_dff_B_T1W1r0Mi2_1;
	wire w_dff_B_hdS1Xd212_0;
	wire w_dff_B_qh3ZIsU17_0;
	wire w_dff_B_pnffsTc89_0;
	wire w_dff_B_Y2FFdj650_0;
	wire w_dff_B_PCe4hWqu0_0;
	wire w_dff_B_iIdX5ytB4_0;
	wire w_dff_B_8ru6XpIH6_0;
	wire w_dff_B_o7zdvJmS4_0;
	wire w_dff_B_jSKjCHVl7_0;
	wire w_dff_B_IPorO2iJ9_0;
	wire w_dff_B_wiAzWvOK8_0;
	wire w_dff_B_59pWEpqM0_0;
	wire w_dff_B_0NrHRDnN8_0;
	wire w_dff_B_z5Yeu1YP3_0;
	wire w_dff_B_2RxG98qb5_0;
	wire w_dff_B_evBNwruV0_0;
	wire w_dff_B_LO9JOhnI8_0;
	wire w_dff_B_LqHYB27G5_0;
	wire w_dff_B_tCYsu0WS0_0;
	wire w_dff_B_YnmLANBf9_2;
	wire w_dff_B_WKybI4lD9_1;
	wire w_dff_B_Nt5hPK6m3_1;
	wire w_dff_B_C4l1m0gX6_1;
	wire w_dff_A_vnhR8o3d4_0;
	wire w_dff_A_GEU44v5Q4_0;
	wire w_dff_A_wfZ8ZsLa1_0;
	wire w_dff_A_F5aYLFnV1_0;
	wire w_dff_A_tmBuKDQV3_0;
	wire w_dff_A_vLkJbTwn0_0;
	wire w_dff_A_1WgpBUtp3_0;
	wire w_dff_A_ilK3GIH75_0;
	wire w_dff_A_Emgmwmvm8_0;
	wire w_dff_A_MfPtqWRG0_0;
	wire w_dff_A_R9fmyxep8_0;
	wire w_dff_A_7wRx7xaG3_0;
	wire w_dff_A_cHzaRFDO4_0;
	wire w_dff_A_G4Xxnea55_0;
	wire w_dff_A_MvsB6TA38_0;
	wire w_dff_A_iA2VBYc17_0;
	wire w_dff_A_GgQ1ID3J5_0;
	wire w_dff_A_bNh4M6Ep2_0;
	wire w_dff_A_TJygGqzl7_2;
	wire w_dff_A_iU15CS426_2;
	wire w_dff_A_dpzeTCi89_2;
	wire w_dff_A_yQgaYmtb1_2;
	wire w_dff_A_cfEQ7Qna0_2;
	wire w_dff_A_E56k601s3_2;
	wire w_dff_A_jio8YAFG7_2;
	wire w_dff_A_PZrhnLXL2_2;
	wire w_dff_A_jxw9vpws8_2;
	wire w_dff_A_cJft473K6_2;
	wire w_dff_A_7PRmW6Ip6_2;
	wire w_dff_A_v5VCptiH7_2;
	wire w_dff_A_O40I5Xo73_2;
	wire w_dff_A_lsbdGSYB5_2;
	wire w_dff_A_VAJHHmLj1_2;
	wire w_dff_A_KKh4rwpx4_2;
	wire w_dff_A_HFgvA4HM3_2;
	wire w_dff_A_IPJr4FrX8_2;
	wire w_dff_A_FHS91h1n8_2;
	wire w_dff_A_HSz7qNpi9_0;
	wire w_dff_A_viGMn3QI9_0;
	wire w_dff_A_5uhSE4tk9_0;
	wire w_dff_A_yD8WmPpv2_0;
	wire w_dff_A_pFbS3kbv3_0;
	wire w_dff_A_eSWenga86_0;
	wire w_dff_A_K2qJq7z68_0;
	wire w_dff_A_JJWtZTpV4_0;
	wire w_dff_A_yc4fj2JV3_0;
	wire w_dff_A_RRimMF1z8_0;
	wire w_dff_A_g6rtoMU50_0;
	wire w_dff_A_NM2AqfPu2_0;
	wire w_dff_A_IhdNb4sX1_0;
	wire w_dff_A_lpLbDs6F4_0;
	wire w_dff_A_2neD71Vj8_0;
	wire w_dff_A_y72R2Axt7_0;
	wire w_dff_A_Hzdn82JJ8_0;
	wire w_dff_A_a1Ck1LAN9_2;
	wire w_dff_A_O6xluIb36_2;
	wire w_dff_A_GiiiFa3n3_2;
	wire w_dff_A_rAuThIDR2_2;
	wire w_dff_A_DHgXbhto7_2;
	wire w_dff_A_7XYq4DsJ4_2;
	wire w_dff_A_K5jHEDma0_2;
	wire w_dff_A_496LZMLI8_2;
	wire w_dff_A_pYJCONra7_2;
	wire w_dff_A_FyPPEUMn5_2;
	wire w_dff_A_Qtz8xAoZ2_2;
	wire w_dff_A_d4lzdykj4_2;
	wire w_dff_A_KXSTPiPM8_2;
	wire w_dff_A_ncMREv2P8_2;
	wire w_dff_A_1dAyC3bT0_2;
	wire w_dff_A_woZw5Kyi8_2;
	wire w_dff_A_4uPCxWrf1_2;
	wire w_dff_A_uif6g65M9_2;
	wire w_dff_A_XOZcIZ1n5_2;
	wire w_dff_A_8Qwl9bBz2_2;
	wire w_dff_B_yYB6TAZo9_0;
	wire w_dff_B_N9rGxIIx6_0;
	wire w_dff_B_Arf4ptQS9_0;
	wire w_dff_B_LT7gTv8j4_0;
	wire w_dff_B_PPi1ZdXw9_0;
	wire w_dff_B_1zYuoSQ24_0;
	wire w_dff_B_9ZxP1CpH4_0;
	wire w_dff_B_dYNfhZ5W5_0;
	wire w_dff_B_8Ouoy7LE7_0;
	wire w_dff_B_15p2zQ3u1_0;
	wire w_dff_B_sPD79SSp3_0;
	wire w_dff_B_THVAymhP4_0;
	wire w_dff_B_h3nGbSLd0_0;
	wire w_dff_B_MLpbz2IM5_0;
	wire w_dff_B_e4BKR3X65_0;
	wire w_dff_B_YKawyxsP8_0;
	wire w_dff_B_ylHZqwYG2_0;
	wire w_dff_B_o3U269by6_0;
	wire w_dff_B_o2lYWXg34_0;
	wire w_dff_B_QTf9ErPX5_1;
	wire w_dff_B_oWAW81qD6_1;
	wire w_dff_B_oMESUjmC8_1;
	wire w_dff_A_3K5qGB1N1_0;
	wire w_dff_A_95xPttmD4_0;
	wire w_dff_A_Di47PCmo2_0;
	wire w_dff_A_GB3lom5E6_0;
	wire w_dff_A_PKL4Ihwc6_0;
	wire w_dff_A_VOAFHszn5_0;
	wire w_dff_A_APFbucbk9_1;
	wire w_dff_A_tXUoP4lF0_0;
	wire w_dff_A_Aw6lNMMU4_0;
	wire w_dff_A_z9ivnzQ28_0;
	wire w_dff_A_wAZAh3OW7_0;
	wire w_dff_A_VYfevSgU1_1;
	wire w_dff_A_IdOvsTrc2_1;
	wire w_dff_A_2k6ktBTe1_0;
	wire w_dff_A_zT7UaD024_0;
	wire w_dff_A_hra1La5V3_0;
	wire w_dff_A_uC2OrI8W5_0;
	wire w_dff_A_Ho32hBRl7_0;
	wire w_dff_A_wEzRSUOx8_0;
	wire w_dff_A_9uvh0oUf1_1;
	wire w_dff_B_Qjq07H452_0;
	wire w_dff_B_Ijvwahbm8_0;
	wire w_dff_B_U1WfJBmg3_0;
	wire w_dff_B_npXesAWe5_0;
	wire w_dff_B_Zv8jywsV7_0;
	wire w_dff_B_RVc9EPDD6_0;
	wire w_dff_B_F2soZxR53_0;
	wire w_dff_B_6hvB721S8_0;
	wire w_dff_B_lBoNCdOZ8_0;
	wire w_dff_B_9lUh3Cp42_0;
	wire w_dff_B_WSczm8ck7_0;
	wire w_dff_B_xbporivq5_0;
	wire w_dff_B_1DElu1if2_0;
	wire w_dff_B_yu3bNiHn0_0;
	wire w_dff_B_w0Eo8hmv1_0;
	wire w_dff_B_eZzwnoab4_0;
	wire w_dff_B_myS6yNBK6_0;
	wire w_dff_B_v9gZSm0M9_0;
	wire w_dff_B_k8e4oTpX8_0;
	wire w_dff_B_YFV8slcf0_0;
	wire w_dff_B_WtmtCWCJ1_1;
	wire w_dff_B_lXMbRhuD4_1;
	wire w_dff_B_HY13YXOs5_1;
	wire w_dff_B_FonaWKoP9_1;
	wire w_dff_B_i6hooBBx6_1;
	wire w_dff_B_pPnBGupb1_1;
	wire w_dff_B_r4f2I6v88_1;
	wire w_dff_B_o77agAi46_1;
	wire w_dff_B_5ZIGr0MD4_1;
	wire w_dff_B_fug5m2Uz6_1;
	wire w_dff_B_PMrZCyXN4_1;
	wire w_dff_B_h1rIcDDy2_1;
	wire w_dff_B_cUS0QtHJ5_1;
	wire w_dff_B_vT0DQTLX3_1;
	wire w_dff_B_4RuFdNRT6_1;
	wire w_dff_B_OX8ualn71_1;
	wire w_dff_B_fKIVnX7K4_1;
	wire w_dff_B_m6W3wUY36_1;
	wire w_dff_B_7enCrB7h2_1;
	wire w_dff_B_m5sqUrVV8_1;
	wire w_dff_B_ObQwgJC15_1;
	wire w_dff_A_5xdz7XYU7_0;
	wire w_dff_A_Hpy5MfOc2_1;
	wire w_dff_B_Ym1YPgLI8_0;
	wire w_dff_B_AtolZT8F9_1;
	wire w_dff_B_pwRJUksx3_1;
	wire w_dff_B_8woNUihl2_1;
	wire w_dff_B_skGCBfp53_1;
	wire w_dff_B_ZRgVQ4vv1_1;
	wire w_dff_B_JL4i2ARc7_1;
	wire w_dff_B_zbAMYEjV6_1;
	wire w_dff_B_aHWdyLhU9_1;
	wire w_dff_B_LWqd3uZb3_1;
	wire w_dff_B_V6K2BZu84_1;
	wire w_dff_B_16LEHejr9_1;
	wire w_dff_B_0660sNOs6_1;
	wire w_dff_B_daWiL30p6_1;
	wire w_dff_B_LD59wa0H4_1;
	wire w_dff_B_RkSYgIEO4_1;
	wire w_dff_B_xxMAb5BD6_1;
	wire w_dff_B_LBvUITzk2_1;
	wire w_dff_B_gbqBUwIl1_1;
	wire w_dff_B_5ibtmSeG1_1;
	wire w_dff_B_AZuUwZqn7_1;
	wire w_dff_B_EWcgwott5_1;
	wire w_dff_A_HFPQpTJG5_0;
	wire w_dff_A_ppmNuYTf8_2;
	wire w_dff_A_eTspS4q13_0;
	wire w_dff_A_yDlvjHw96_0;
	wire w_dff_A_1hELk9MS9_1;
	wire w_dff_A_4nj4cidn5_0;
	wire w_dff_A_76uPv6W69_0;
	wire w_dff_A_OEPIWn4Y0_0;
	wire w_dff_A_rwowK5U84_0;
	wire w_dff_A_luLEJHA67_0;
	wire w_dff_A_NTrox4ME1_0;
	wire w_dff_A_oTeowHYw0_0;
	wire w_dff_A_XzEB0ILD7_0;
	wire w_dff_A_DL87QF4n7_0;
	wire w_dff_A_c9J82Jq75_0;
	wire w_dff_A_VMh60d2x4_0;
	wire w_dff_A_yBwxPKn73_1;
	wire w_dff_A_DRZzqlun9_1;
	wire w_dff_A_pFQl3gRB8_1;
	wire w_dff_A_eZp5P86f6_1;
	wire w_dff_B_FXNeghKD8_3;
	wire w_dff_B_KHVOwOSr1_3;
	wire w_dff_B_B8UBqGIR9_3;
	wire w_dff_B_6qKQzCyJ9_3;
	wire w_dff_B_3aabpeHx6_3;
	wire w_dff_B_68lGMx9Z2_3;
	wire w_dff_B_7zwlRWqY0_3;
	wire w_dff_B_VhKtsMnV0_3;
	wire w_dff_B_XHslf9w03_3;
	wire w_dff_B_KcfGaCcD5_0;
	wire w_dff_A_0vW8M7pl8_0;
	wire w_dff_B_CRtjkcmB5_0;
	wire w_dff_B_XD00l3zH0_0;
	wire w_dff_B_qQ5xfVII6_0;
	wire w_dff_B_MOeP6t8y4_0;
	wire w_dff_B_pN7XJb359_0;
	wire w_dff_B_EZtPf5V10_0;
	wire w_dff_B_6nFsEehQ2_0;
	wire w_dff_B_qsbTU6aX5_0;
	wire w_dff_B_ZRSVymbL6_0;
	wire w_dff_B_xFuDborj1_0;
	wire w_dff_B_ZP3Ou09r3_0;
	wire w_dff_B_t1GA4otx5_0;
	wire w_dff_B_TYfR1S6V5_0;
	wire w_dff_B_nOX7kZNc2_0;
	wire w_dff_B_Lwbztwl10_0;
	wire w_dff_B_F7ipmCq31_0;
	wire w_dff_B_bZvC7fT64_0;
	wire w_dff_B_XKntAtJb8_0;
	wire w_dff_B_ihjrzGeK4_0;
	wire w_dff_B_hv1i2ayl9_2;
	wire w_dff_B_r4QAimLG6_2;
	wire w_dff_B_PZmhi2Ux9_2;
	wire w_dff_B_tiUFcGwx2_1;
	wire w_dff_B_5TN3qEZ67_1;
	wire w_dff_B_6BA4nhSw3_1;
	wire w_dff_B_BtdO2gts0_1;
	wire w_dff_B_ePHP2b9y8_1;
	wire w_dff_B_fcLVQSPd9_1;
	wire w_dff_B_EB1jyn2G3_1;
	wire w_dff_B_SwwdMu4Y8_1;
	wire w_dff_B_Y0z90IVy1_1;
	wire w_dff_B_6X7uMZkU6_1;
	wire w_dff_B_Q2EHH6wW5_1;
	wire w_dff_B_GyAtbnbc1_1;
	wire w_dff_B_uBwPSrnu7_1;
	wire w_dff_B_nszbMZii6_1;
	wire w_dff_B_kOvO2zm75_1;
	wire w_dff_B_7ZKBsrZl6_1;
	wire w_dff_B_lMTC9uL96_0;
	wire w_dff_B_NaHG9NqN9_0;
	wire w_dff_B_ePknq90s6_0;
	wire w_dff_B_9zm5aosW8_0;
	wire w_dff_B_K9NaHNCa3_0;
	wire w_dff_B_xDbWoImo4_0;
	wire w_dff_B_q0elnQ2I0_0;
	wire w_dff_B_Li3oPenu2_0;
	wire w_dff_B_75NlZSdJ8_0;
	wire w_dff_B_ZXo0Ajip9_1;
	wire w_dff_B_GWbKGlHL4_1;
	wire w_dff_B_UdMAZiz87_1;
	wire w_dff_B_aljd1Jnr4_1;
	wire w_dff_A_vrU2TEnj8_0;
	wire w_dff_A_c63SQAcV4_0;
	wire w_dff_A_IhPVHmS03_0;
	wire w_dff_A_ppsnujPY6_0;
	wire w_dff_A_L3tuD2tc0_0;
	wire w_dff_A_eY1SVWxl9_0;
	wire w_dff_A_A9qC9FTc9_1;
	wire w_dff_B_wd3WBX613_1;
	wire w_dff_B_6TtA3TpS8_1;
	wire w_dff_B_5xvRDIY67_1;
	wire w_dff_B_8dNRyRnD0_1;
	wire w_dff_B_bPLbmZ3P5_1;
	wire w_dff_B_5aPzewHF4_1;
	wire w_dff_B_mUOTr4No8_1;
	wire w_dff_B_tCN1YVT29_1;
	wire w_dff_B_EHvUj70j2_1;
	wire w_dff_B_yJWGdK1H6_1;
	wire w_dff_B_J8o4nnxb3_1;
	wire w_dff_B_nhj6bx8W5_0;
	wire w_dff_B_QAm637499_0;
	wire w_dff_B_iyvZikVc5_0;
	wire w_dff_B_qxjqu7PP5_0;
	wire w_dff_B_sltbgdBD4_0;
	wire w_dff_B_Ghv57Xo84_0;
	wire w_dff_B_fx5k9FZY9_0;
	wire w_dff_A_2Oqkcr7F2_1;
	wire w_dff_A_qO258kTB7_1;
	wire w_dff_A_WqYq0zA37_1;
	wire w_dff_A_GxTLhJZx7_1;
	wire w_dff_A_wfN3sNeB6_1;
	wire w_dff_B_WcBNWtOU8_1;
	wire w_dff_B_bapi0k3s0_1;
	wire w_dff_B_e1ncb7Vw9_1;
	wire w_dff_B_ymZyGPr64_1;
	wire w_dff_B_ndtNxg8A0_1;
	wire w_dff_B_SyvHB0u91_1;
	wire w_dff_B_0RGx7qUb3_1;
	wire w_dff_B_F7iw6GAC2_1;
	wire w_dff_A_ewr4SXXH1_0;
	wire w_dff_A_atevLuvj3_0;
	wire w_dff_A_31nNRVPo0_0;
	wire w_dff_A_PTfTAvJb1_0;
	wire w_dff_A_hdUzfdID3_1;
	wire w_dff_A_vpSkG3G47_1;
	wire w_dff_B_3gObBvtq6_1;
	wire w_dff_B_7BNYNatJ7_1;
	wire w_dff_B_vWtlvFBq7_1;
	wire w_dff_B_pal9sUyi5_1;
	wire w_dff_B_sxWPdZfA4_1;
	wire w_dff_B_pd2DNL1X3_1;
	wire w_dff_B_QU100WUX8_1;
	wire w_dff_B_27yDHJjp1_1;
	wire w_dff_B_tUL6pXNC2_1;
	wire w_dff_B_quc5fPgB3_1;
	wire w_dff_B_JY4lHCv44_1;
	wire w_dff_B_uGKSFA9M9_1;
	wire w_dff_B_qZageBzx2_1;
	wire w_dff_B_Kqho8I655_1;
	wire w_dff_B_zzhyHL5h9_1;
	wire w_dff_B_xYUlCryM1_1;
	wire w_dff_B_kAxv4aJy7_1;
	wire w_dff_B_T6D8dj7o7_1;
	wire w_dff_B_jthn2JR95_1;
	wire w_dff_B_FMdVkkiS9_1;
	wire w_dff_B_RlXyN75Z2_1;
	wire w_dff_B_HffqlGeD3_1;
	wire w_dff_B_BrRlp7DK5_1;
	wire w_dff_B_HtTzx4SS0_1;
	wire w_dff_B_g4pXpyvD2_1;
	wire w_dff_B_qMC45aoi3_1;
	wire w_dff_B_Ryg6WJ9s5_1;
	wire w_dff_B_mYKFUuBt2_1;
	wire w_dff_B_ODHRcNGn0_1;
	wire w_dff_B_WB9zdLi83_1;
	wire w_dff_B_VSfgctiF3_1;
	wire w_dff_B_h15wSets3_1;
	wire w_dff_B_nA4l5icK4_1;
	wire w_dff_B_FO7cTvde1_1;
	wire w_dff_B_IQtoGsNT7_1;
	wire w_dff_B_qgl7C1FO8_1;
	wire w_dff_B_BQmwYZ0S5_1;
	wire w_dff_B_wmaGa7Tq4_1;
	wire w_dff_B_3GEBUdvs2_1;
	wire w_dff_B_txWFpU7O5_1;
	wire w_dff_B_LLRgr22f0_1;
	wire w_dff_B_8WiDnjDU1_1;
	wire w_dff_B_4zoGhQZS1_1;
	wire w_dff_B_A6XYkeE92_1;
	wire w_dff_B_poQmnGEx7_1;
	wire w_dff_B_Cp2TkbYB7_1;
	wire w_dff_B_rM69akLu3_1;
	wire w_dff_B_hhR8mnqz5_1;
	wire w_dff_B_M8GRt5Zw8_1;
	wire w_dff_B_73a9uzZc8_1;
	wire w_dff_B_GNB9tcu21_1;
	wire w_dff_B_EzmdNFix3_1;
	wire w_dff_B_eInc3zi74_1;
	wire w_dff_B_gwymAcpq4_1;
	wire w_dff_B_6atzRXp50_1;
	wire w_dff_B_0c6LfmK61_1;
	wire w_dff_B_yOGDY6he7_1;
	wire w_dff_B_DevnYb509_1;
	wire w_dff_B_3LTRgAEm6_1;
	wire w_dff_B_5P3q6PZK0_1;
	wire w_dff_B_pKYzJm8L7_1;
	wire w_dff_B_gh8tn6QU6_1;
	wire w_dff_B_pIKEtVug2_1;
	wire w_dff_B_YBUokWUn1_1;
	wire w_dff_B_UQh2oZzD2_1;
	wire w_dff_B_mLOE9ARC1_1;
	wire w_dff_B_7C5wYFeg3_1;
	wire w_dff_B_tCXuAXLT7_1;
	wire w_dff_B_D6QwLJ9m6_1;
	wire w_dff_B_VqM9cSes9_1;
	wire w_dff_B_5XZ1CRXX8_1;
	wire w_dff_B_GXFxBcp05_1;
	wire w_dff_B_QMHplCug2_1;
	wire w_dff_B_WPIHHPTY2_1;
	wire w_dff_B_kWb1quw83_1;
	wire w_dff_B_rEvkE60D6_0;
	wire w_dff_B_zINwDq7O3_0;
	wire w_dff_B_zQ9aCCvk7_0;
	wire w_dff_B_lqbikiFs9_0;
	wire w_dff_B_ikIkOiEX1_0;
	wire w_dff_B_g8HhNVks3_0;
	wire w_dff_B_hZfhGPNm0_0;
	wire w_dff_B_JHIZx4mV9_0;
	wire w_dff_B_OaAbXU2z9_0;
	wire w_dff_B_0wWjNpv39_0;
	wire w_dff_B_4kuolSpY5_1;
	wire w_dff_B_jz1Kwpoq7_1;
	wire w_dff_B_uH0ugx2r4_1;
	wire w_dff_B_YLf6kt0O4_1;
	wire w_dff_B_ygeRtY650_1;
	wire w_dff_B_RSAys7RH0_1;
	wire w_dff_B_PGwbWVVH2_1;
	wire w_dff_B_FebDitlu7_1;
	wire w_dff_B_ICYdCDT54_1;
	wire w_dff_B_pyHhzsWM4_1;
	wire w_dff_B_MyokzfJG6_1;
	wire w_dff_B_qatXc8VV6_1;
	wire w_dff_B_5f5v76gk3_1;
	wire w_dff_B_9T0J95il7_1;
	wire w_dff_B_0D9ogn6Y8_1;
	wire w_dff_B_MF9Owc8L0_1;
	wire w_dff_B_kYjK86vv1_1;
	wire w_dff_B_QCQEHJBJ9_0;
	wire w_dff_B_NwUqWdPU1_2;
	wire w_dff_B_KUr6AdJf3_2;
	wire w_dff_B_6Z1okz4h3_2;
	wire w_dff_B_yroClNli2_0;
	wire w_dff_B_zdAzHRRF8_0;
	wire w_dff_B_6UYEQL2x2_0;
	wire w_dff_B_mfpd21pw8_0;
	wire w_dff_B_udkTUowa9_0;
	wire w_dff_B_hs6jSJjl1_0;
	wire w_dff_B_AWSvcsWE1_0;
	wire w_dff_B_rz8kvVKx4_0;
	wire w_dff_B_m0Oq0xMV3_0;
	wire w_dff_B_yYVWrSDQ9_0;
	wire w_dff_B_oNLfMOBy9_0;
	wire w_dff_B_zHKFq20D8_0;
	wire w_dff_B_4W0Uptyo6_0;
	wire w_dff_B_7Iq5rWsd2_0;
	wire w_dff_B_pMCEaWye6_0;
	wire w_dff_B_RssjXhAQ3_0;
	wire w_dff_B_8hCC8MqE5_0;
	wire w_dff_B_cRRZ9vyq5_0;
	wire w_dff_B_aECCcNub3_0;
	wire w_dff_B_j1n3kkOT6_0;
	wire w_dff_B_shkYsADX0_2;
	wire w_dff_B_ForsF7Gk3_2;
	wire w_dff_B_GHXBL6V70_2;
	wire w_dff_B_SATYeYta6_1;
	wire w_dff_B_IRc6Jqif2_1;
	wire w_dff_B_SuASEOwW9_1;
	wire w_dff_B_khujN4kz9_1;
	wire w_dff_B_F3Kxm83X1_1;
	wire w_dff_B_8dQBZvQ76_1;
	wire w_dff_B_aQaHBYYT8_1;
	wire w_dff_B_tlWiEksU1_1;
	wire w_dff_B_V4g9B0Bc1_1;
	wire w_dff_B_4IMke6an4_1;
	wire w_dff_B_is8T0Zvx8_1;
	wire w_dff_B_uY0k4gIV8_1;
	wire w_dff_B_p4AXBXKC0_1;
	wire w_dff_B_NTB3WyIr9_1;
	wire w_dff_B_KGmhtZ5V7_1;
	wire w_dff_B_jXg2uAaj1_1;
	wire w_dff_B_gDMHa5dD1_0;
	wire w_dff_B_hnlt39in2_0;
	wire w_dff_B_CzjmnqsG2_0;
	wire w_dff_B_Uk6SWWo31_0;
	wire w_dff_B_amk12isJ4_0;
	wire w_dff_B_aqHn981c9_0;
	wire w_dff_B_TOhZOnpB9_0;
	wire w_dff_B_Y2HgL4gd1_0;
	wire w_dff_B_JAOvdGPG3_0;
	wire w_dff_B_Vhmy5KCT8_0;
	wire w_dff_A_HArAgng82_1;
	wire w_dff_A_M0jMOAI95_1;
	wire w_dff_A_9OEWihJg9_1;
	wire w_dff_B_2TSL03jK6_1;
	wire w_dff_B_q9Ly9YM44_3;
	wire w_dff_B_cRRncVaF6_1;
	wire w_dff_A_VoJQY4mK5_0;
	wire w_dff_A_zOK6Sc6G1_0;
	wire w_dff_A_W72xPigz0_0;
	wire w_dff_A_XUWvpTXo5_0;
	wire w_dff_A_7EGXfocg3_0;
	wire w_dff_A_jj5mAno66_0;
	wire w_dff_A_aKgZac1K6_0;
	wire w_dff_A_mDIJjcnI8_0;
	wire w_dff_A_moObGmSF6_0;
	wire w_dff_A_2m1qgmXz6_0;
	wire w_dff_A_O9OK7o6x9_0;
	wire w_dff_A_09PEiPU34_1;
	wire w_dff_A_uXdx9I4O0_1;
	wire w_dff_B_9fTv7oJp4_1;
	wire w_dff_B_c0RnFSPh6_1;
	wire w_dff_B_Wu4ANowT3_1;
	wire w_dff_B_Eq7yUAjh0_1;
	wire w_dff_B_zqJrC4xK2_1;
	wire w_dff_B_YgrLRGQT5_1;
	wire w_dff_A_yPdgnVZq1_0;
	wire w_dff_A_EQO7aPUZ7_0;
	wire w_dff_A_Sdgvmiav8_1;
	wire w_dff_A_IFemFwP97_1;
	wire w_dff_A_DB8a6sF52_1;
	wire w_dff_B_babhDdva3_1;
	wire w_dff_B_Or80r8Bu4_1;
	wire w_dff_A_bDAjTJQY5_0;
	wire w_dff_A_5i6QK7o84_1;
	wire w_dff_B_50hXFk5M3_1;
	wire w_dff_B_FFfn2ho82_1;
	wire w_dff_B_SIN1FyzY3_1;
	wire w_dff_B_Yu8UBpLi6_1;
	wire w_dff_B_xWGtZ0OT7_1;
	wire w_dff_B_Kmxdsp1M9_1;
	wire w_dff_B_R9w9evNC0_1;
	wire w_dff_B_6JhyAsAc9_1;
	wire w_dff_B_AGGg2M6Z2_1;
	wire w_dff_B_cFioTv9R6_1;
	wire w_dff_B_wFZP9U8Z9_1;
	wire w_dff_B_oMLOhkRf6_1;
	wire w_dff_B_e3JhcnfG7_1;
	wire w_dff_B_ot4T40aM7_1;
	wire w_dff_B_UZUkPoFP0_1;
	wire w_dff_B_dmjTBYiW3_1;
	wire w_dff_B_zaz4tCVY8_1;
	wire w_dff_B_neIGb0Nn7_1;
	wire w_dff_B_w0ha3GHo1_1;
	wire w_dff_B_iyvx0Osu3_1;
	wire w_dff_B_ypEKkKHu1_1;
	wire w_dff_B_1HBEN5Er7_1;
	wire w_dff_B_9orisDh76_1;
	wire w_dff_B_NwbyyCxe4_1;
	wire w_dff_B_ovtLENyn1_1;
	wire w_dff_B_TA9c7iQR3_1;
	wire w_dff_A_KpkyMcK08_0;
	wire w_dff_A_AIMvmSNJ1_0;
	wire w_dff_A_uAYq9qwW0_0;
	wire w_dff_A_sXdHsCJz1_0;
	wire w_dff_A_Sp5I7ldP9_0;
	wire w_dff_A_vqtaKSFB4_0;
	wire w_dff_A_mlYvGYp88_0;
	wire w_dff_A_BDO4lIXq1_0;
	wire w_dff_A_M55HYp4e6_0;
	wire w_dff_A_5CRQ0zB80_1;
	wire w_dff_A_jES8ImbP5_1;
	wire w_dff_A_g6TZUcjN9_1;
	wire w_dff_A_rH4vGzSu7_1;
	wire w_dff_A_l22ymRVk8_1;
	wire w_dff_A_r41c0YZ74_1;
	wire w_dff_A_tsD94GUS7_1;
	wire w_dff_A_usWIVe4r6_1;
	wire w_dff_A_VbB6nsO87_1;
	wire w_dff_A_Gm075tNU0_1;
	wire w_dff_A_8x7QodEG0_1;
	wire w_dff_A_GPQp5Te57_1;
	wire w_dff_A_MpLo72ts6_2;
	wire w_dff_A_3E1I7apd9_2;
	wire w_dff_A_gY5xpIeV8_2;
	wire w_dff_A_DFk1rNYC3_2;
	wire w_dff_A_9YSRrLIq5_2;
	wire w_dff_A_ceGm2RIz5_2;
	wire w_dff_A_khqusC305_2;
	wire w_dff_A_ZIh2Izqh5_2;
	wire w_dff_A_oOh3FEj50_2;
	wire w_dff_A_kRe9C1FU2_2;
	wire w_dff_B_2Ko6HozK1_1;
	wire w_dff_B_4nhfmZyy7_1;
	wire w_dff_A_kCA1roIz8_0;
	wire w_dff_A_Ii9nEp3G4_1;
	wire w_dff_A_Uantm8hy6_0;
	wire w_dff_A_EvlWgjHm5_0;
	wire w_dff_A_zFhXjUh34_0;
	wire w_dff_A_5SjB4z280_0;
	wire w_dff_A_GTGvGoaV3_0;
	wire w_dff_A_9SF0wWVx1_0;
	wire w_dff_A_5UICh8js7_1;
	wire w_dff_A_fvgm4vOr9_1;
	wire w_dff_A_jFoquQJb9_1;
	wire w_dff_A_rm8v5iUM7_1;
	wire w_dff_A_rqTSfhJM6_1;
	wire w_dff_A_ViVAQnti7_1;
	wire w_dff_A_z3v7vRp71_1;
	wire w_dff_B_IaT2PVUl3_0;
	wire w_dff_B_OPohOdCj5_0;
	wire w_dff_B_Sz85MPJU5_0;
	wire w_dff_B_aKXskUcH3_0;
	wire w_dff_B_9uX8harz7_0;
	wire w_dff_B_9QUziSNQ6_0;
	wire w_dff_B_dhOeJycN7_0;
	wire w_dff_B_jBhjZjjS2_0;
	wire w_dff_B_57gpdxxg8_0;
	wire w_dff_B_0MA2VM3V0_0;
	wire w_dff_B_9qarWJfO7_0;
	wire w_dff_B_ijD61zwB8_0;
	wire w_dff_B_bkfVty1l4_0;
	wire w_dff_B_5qIDoWML4_0;
	wire w_dff_B_w3f5EaIq8_0;
	wire w_dff_B_NRyAP7tH3_0;
	wire w_dff_B_fzndBmR54_0;
	wire w_dff_B_l1DuayOK1_0;
	wire w_dff_B_80SRCvM26_0;
	wire w_dff_B_E3wrtXIv4_0;
	wire w_dff_B_ZoSLA8cb9_2;
	wire w_dff_B_7uLmyHdV4_2;
	wire w_dff_B_fGuvLndO3_2;
	wire w_dff_B_V0qgLHDs2_1;
	wire w_dff_B_9KWmcCOm7_1;
	wire w_dff_B_f1VurmMl8_1;
	wire w_dff_B_N78XHgTI0_1;
	wire w_dff_B_TihVkcu21_1;
	wire w_dff_B_8gj5Y2tG9_1;
	wire w_dff_B_YJDpsx4H3_1;
	wire w_dff_B_HCH1NubT5_1;
	wire w_dff_B_XW4WyXIR5_1;
	wire w_dff_B_CelSJfSW6_1;
	wire w_dff_B_fAe2TAn28_1;
	wire w_dff_B_8qwtpWrV4_1;
	wire w_dff_B_V4Ppvtsg0_1;
	wire w_dff_B_34MWWBSD3_1;
	wire w_dff_B_G67N6VPI7_1;
	wire w_dff_B_BGM5W6S45_1;
	wire w_dff_B_GKfzRS3d7_0;
	wire w_dff_B_VzNzpOiO9_0;
	wire w_dff_B_lJ3dHqQx5_0;
	wire w_dff_B_QVsNxBfM1_0;
	wire w_dff_B_Tzipyeb02_0;
	wire w_dff_B_eD5iR0z97_0;
	wire w_dff_B_jZNhevm24_0;
	wire w_dff_B_yv72Z9yD3_0;
	wire w_dff_B_aXOr8GyN4_0;
	wire w_dff_B_VmEIurYj1_0;
	wire w_dff_B_WLwvlIPA5_0;
	wire w_dff_B_s4WOZmBm6_0;
	wire w_dff_A_BH3rsD105_1;
	wire w_dff_A_rLeApYgQ2_1;
	wire w_dff_A_nymskFp84_2;
	wire w_dff_A_Zoy8pnXB4_2;
	wire w_dff_B_7CzP2E2L3_0;
	wire w_dff_B_m8lrl0n79_0;
	wire w_dff_A_BmOSzjts1_0;
	wire w_dff_A_sGehzmu81_0;
	wire w_dff_A_Rni5PH7f7_0;
	wire w_dff_A_u0eNrmBu4_0;
	wire w_dff_A_GbWrzrA04_0;
	wire w_dff_A_dgYS5rF39_0;
	wire w_dff_A_HKIO64mQ1_0;
	wire w_dff_A_6WBjMV9a8_0;
	wire w_dff_A_IjOfffxg2_0;
	wire w_dff_A_5zH7QhnH9_1;
	wire w_dff_A_wJ3Ouuzb5_1;
	wire w_dff_A_WbcQvHDP1_1;
	wire w_dff_A_w3gOLomI2_1;
	wire w_dff_A_NxClbYBH0_0;
	wire w_dff_A_1Dx4HAHp7_2;
	wire w_dff_A_qso3eQg61_2;
	wire w_dff_A_xQg7Be0V8_2;
	wire w_dff_A_UcqKxuSJ8_2;
	wire w_dff_A_oZwZOjGH5_2;
	wire w_dff_A_xj9gEQvJ1_2;
	wire w_dff_A_eLxW5qXp5_2;
	wire w_dff_A_1CdI0S0G6_2;
	wire w_dff_A_rdRbeQpz7_2;
	wire w_dff_A_DKIsNxmh3_2;
	wire w_dff_A_tFqvLuoQ2_2;
	wire w_dff_A_nnfxkria6_2;
	wire w_dff_A_LFp7k7aZ3_2;
	wire w_dff_A_aOqhSAk29_2;
	wire w_dff_A_u5tFlz3S7_0;
	wire w_dff_A_bJ19DS6e9_0;
	wire w_dff_A_phMaxgek3_0;
	wire w_dff_A_4i0Tqhj48_2;
	wire w_dff_A_0YtcJIVr1_2;
	wire w_dff_A_5ZHG9g6R5_0;
	wire w_dff_A_wfRDHPzP8_0;
	wire w_dff_A_hD979AwS9_0;
	wire w_dff_A_9HBBF0OZ2_0;
	wire w_dff_A_kNJtKEVH1_0;
	wire w_dff_A_A93dWc351_0;
	wire w_dff_A_1fpD5eUO1_0;
	wire w_dff_A_1UH77wLh7_0;
	wire w_dff_A_H4V82B3V1_0;
	wire w_dff_A_DKLNwFK66_1;
	wire w_dff_A_u2T2DKa28_1;
	wire w_dff_B_7eAZoxY13_3;
	wire w_dff_B_CWRxvdPn2_3;
	wire w_dff_B_4g4Q6Rvf1_3;
	wire w_dff_B_7pfkPapK2_3;
	wire w_dff_B_IGDUEajs0_3;
	wire w_dff_B_wcC1iBGy8_3;
	wire w_dff_B_ylLpoCZ65_3;
	wire w_dff_B_dQiEg0El9_3;
	wire w_dff_B_sJ1C3hQo8_3;
	wire w_dff_B_gaPX4nAc7_3;
	wire w_dff_B_djOsCc3g3_3;
	wire w_dff_B_FHX8TLny0_1;
	wire w_dff_B_P19qavdH1_1;
	wire w_dff_B_ycbutOvK2_1;
	wire w_dff_B_Soo3w26k1_1;
	wire w_dff_B_7pt7jynQ8_1;
	wire w_dff_B_mZSUNb9g1_1;
	wire w_dff_B_NBxSAoRi8_1;
	wire w_dff_B_n9wQfuIa9_1;
	wire w_dff_B_njhLuD006_1;
	wire w_dff_B_SohIp7eS4_1;
	wire w_dff_B_VEGbVZ7T5_1;
	wire w_dff_B_hel2dOG81_1;
	wire w_dff_B_tX8kMrfL6_1;
	wire w_dff_B_mlc6LtcC8_1;
	wire w_dff_B_5faaRwDs5_1;
	wire w_dff_B_HTpe1VCg2_1;
	wire w_dff_B_0Z5IiwPq7_1;
	wire w_dff_B_BjCTQoto0_1;
	wire w_dff_B_VckX4ovK6_1;
	wire w_dff_B_MbvjTpVM5_1;
	wire w_dff_B_LA1x1T553_1;
	wire w_dff_B_DEk286bu7_1;
	wire w_dff_B_9V0H138A9_1;
	wire w_dff_B_Ghu6kiR09_1;
	wire w_dff_B_L9lWMhdF2_1;
	wire w_dff_B_o8GKBQRI7_1;
	wire w_dff_B_iWhCo6B03_1;
	wire w_dff_B_i48UCTAL8_1;
	wire w_dff_B_E104wsN56_1;
	wire w_dff_B_GCUTKeC38_1;
	wire w_dff_B_pdUuINJl0_1;
	wire w_dff_B_UpfYWGsR2_1;
	wire w_dff_B_K3RuSd0b4_1;
	wire w_dff_B_4gLCdTGb0_1;
	wire w_dff_B_pOTZXhRw8_1;
	wire w_dff_B_TULGqpbe4_1;
	wire w_dff_B_r2KtQKQg4_1;
	wire w_dff_B_rLWnffD82_1;
	wire w_dff_B_pJBymsxM6_1;
	wire w_dff_B_ulWuoMYT0_1;
	wire w_dff_B_1etY6Mwd5_0;
	wire w_dff_B_GEUE8hrs9_1;
	wire w_dff_B_9UXiCv0m5_1;
	wire w_dff_A_zhbpJqqR3_1;
	wire w_dff_B_Djb85jzw6_3;
	wire w_dff_B_XbMfPNC78_3;
	wire w_dff_B_kXpySNY15_3;
	wire w_dff_B_7lgsNG6L1_3;
	wire w_dff_B_3BFNaT9z0_3;
	wire w_dff_A_nshC9MZh4_0;
	wire w_dff_A_ZLrIieCK1_1;
	wire w_dff_A_Tjcoy3949_1;
	wire w_dff_B_6soiylNA4_3;
	wire w_dff_B_gaxXnFkz7_3;
	wire w_dff_B_D6GWk81n4_3;
	wire w_dff_B_hKojJ9Rp0_3;
	wire w_dff_B_KLBHPtCb3_3;
	wire w_dff_B_boVhpqj27_3;
	wire w_dff_B_x6UQqVXX7_3;
	wire w_dff_B_7XORGzGK5_3;
	wire w_dff_B_nu7RB4Nl2_3;
	wire w_dff_B_XZuJ79wq8_3;
	wire w_dff_B_TJkDqrhs3_3;
	wire w_dff_B_3PiQHyt39_3;
	wire w_dff_B_oqp7mgxB8_3;
	wire w_dff_B_G1XF9B541_3;
	wire w_dff_B_Vg4hOFcp5_3;
	wire w_dff_A_LypQKKcW0_0;
	wire w_dff_A_yXRHn23c6_0;
	wire w_dff_A_kAPst4rG7_0;
	wire w_dff_A_olHE7vfl9_0;
	wire w_dff_A_LWuJLPGe4_0;
	wire w_dff_A_93243qg33_0;
	wire w_dff_A_L9n2n8oJ8_1;
	wire w_dff_A_edaGDRxl6_1;
	wire w_dff_A_Z4Y8e3Fm2_1;
	wire w_dff_A_2jivuVoV2_1;
	wire w_dff_A_vYseTm2Q7_1;
	wire w_dff_A_N2iAANj73_1;
	wire w_dff_A_tdTttx1A4_0;
	wire w_dff_A_6TS6vlq43_0;
	wire w_dff_A_UnODfP1e7_0;
	wire w_dff_A_AA0Aec4E5_0;
	wire w_dff_A_pg1yx1tx3_0;
	wire w_dff_A_vqeYpe6u4_0;
	wire w_dff_A_T1XhDIww2_0;
	wire w_dff_A_riKcW56x8_0;
	wire w_dff_A_nmRawhVX0_0;
	wire w_dff_A_orhdBHcl5_0;
	wire w_dff_A_KUKgTNlP7_0;
	wire w_dff_A_jhT5jWgK2_0;
	wire w_dff_A_fZvtdc804_0;
	wire w_dff_A_UGEY9o3W6_0;
	wire w_dff_A_2WSEciTN5_1;
	wire w_dff_A_r6mjsyH68_1;
	wire w_dff_B_Ehju4Z324_1;
	wire w_dff_B_uKlhyMAY6_1;
	wire w_dff_B_wDrfRkwT3_0;
	wire w_dff_B_Cwc16hRW5_0;
	wire w_dff_B_vWWfOqqQ9_0;
	wire w_dff_B_D5UDEj6N8_0;
	wire w_dff_B_bzNCjmpl3_0;
	wire w_dff_B_dLbIVf7M8_0;
	wire w_dff_B_3o1tM25u3_0;
	wire w_dff_B_SOWLTAqs1_0;
	wire w_dff_B_L4TOTHkU6_0;
	wire w_dff_B_AvUsMNqQ5_0;
	wire w_dff_B_qosWfwVb2_0;
	wire w_dff_B_0EAHIAn80_0;
	wire w_dff_B_4saqOU3Y3_0;
	wire w_dff_B_Ec75XCn20_0;
	wire w_dff_B_HvZxSwsH1_0;
	wire w_dff_B_1Y5pUuUD6_0;
	wire w_dff_B_ow9X3H7R6_0;
	wire w_dff_B_us0caNch4_1;
	wire w_dff_B_OIAyBtWZ3_1;
	wire w_dff_B_qS653Y2i8_1;
	wire w_dff_B_o2XB3q0z2_0;
	wire w_dff_B_N02CtFAU5_0;
	wire w_dff_B_y3ymCFBe5_0;
	wire w_dff_B_N5YZXX2n3_0;
	wire w_dff_B_GVlPamiQ3_0;
	wire w_dff_B_BIpqgLrW3_0;
	wire w_dff_B_gFIt59JH6_0;
	wire w_dff_B_cNBuyqeU3_0;
	wire w_dff_B_t8gWkXLY8_0;
	wire w_dff_B_SPPxYmft4_0;
	wire w_dff_B_JMA2Ojso9_0;
	wire w_dff_B_bdhzgnpS6_0;
	wire w_dff_B_5yvKG2eJ0_0;
	wire w_dff_B_I2IkDyHH9_0;
	wire w_dff_B_61X5ZuyU4_0;
	wire w_dff_B_NaYOdTpP1_0;
	wire w_dff_B_9NRyjmDE9_0;
	wire w_dff_B_PBRsEGmR6_1;
	wire w_dff_B_1u8wWBmn5_1;
	wire w_dff_B_E0dWacZS0_1;
	wire w_dff_A_YlAgmg6T7_0;
	wire w_dff_A_rcfcSIjf5_0;
	wire w_dff_A_Jn97mrZK5_0;
	wire w_dff_A_C4NNP8Xo9_0;
	wire w_dff_A_5lvsBwnu3_0;
	wire w_dff_A_xfi47aKt6_1;
	wire w_dff_A_XX8s0kTl5_1;
	wire w_dff_A_wcH6QTuZ3_1;
	wire w_dff_A_R2cCntsR9_1;
	wire w_dff_A_2ThLU8My3_0;
	wire w_dff_A_PUvMD4Qh7_0;
	wire w_dff_A_0T5gnU6g4_0;
	wire w_dff_A_RIoXXCcc6_0;
	wire w_dff_A_Rcqv1pnE6_0;
	wire w_dff_A_mFeMHTtF2_1;
	wire w_dff_A_v7kFF0zp0_1;
	wire w_dff_A_KkthLwDo4_1;
	wire w_dff_A_u4fEX5Gh2_1;
	wire w_dff_A_6vxKppbj8_0;
	wire w_dff_A_Q1y0rw1J0_0;
	wire w_dff_A_MYjoLYpB8_0;
	wire w_dff_B_zEo4q6Xh3_1;
	wire w_dff_B_BJBS0wp33_1;
	wire w_dff_B_nsg6w8Jg1_1;
	wire w_dff_B_9DeTDEkl1_1;
	wire w_dff_B_eqHr8K7Z4_1;
	wire w_dff_B_m6uGQahr0_1;
	wire w_dff_B_w4OiuBEM4_1;
	wire w_dff_B_uGzj4GnF2_1;
	wire w_dff_B_Cu8AVbP31_1;
	wire w_dff_B_3T8p3AbB2_1;
	wire w_dff_B_bSBCFu0d3_1;
	wire w_dff_B_cMV8N3sX5_1;
	wire w_dff_B_8oSCkhnx1_1;
	wire w_dff_B_pvphTkoP5_1;
	wire w_dff_B_P2UAXcJf8_1;
	wire w_dff_B_d6bv0RBw7_1;
	wire w_dff_B_YPFyJM4S1_1;
	wire w_dff_B_eiqe9rVO8_1;
	wire w_dff_B_u3QlNxvx7_1;
	wire w_dff_B_tirUx62I2_1;
	wire w_dff_B_rxo2Dayk1_1;
	wire w_dff_B_DQdEZMtx8_1;
	wire w_dff_B_Xab86eH79_1;
	wire w_dff_A_hdXM7sbV1_1;
	wire w_dff_A_Z0m7DK4o2_1;
	wire w_dff_A_Q03PM3lt4_1;
	wire w_dff_A_YmGFXRcK2_1;
	wire w_dff_A_v0v4KUoW6_1;
	wire w_dff_A_lEOxaR872_1;
	wire w_dff_A_uFJdQoKg6_1;
	wire w_dff_A_hWrlshFl1_1;
	wire w_dff_A_7UY9nmdC8_1;
	wire w_dff_A_niaUuaPX1_1;
	wire w_dff_A_sKnW5gSz2_1;
	wire w_dff_A_qh4CeztD9_1;
	wire w_dff_A_ygC8iK3D9_1;
	wire w_dff_A_29YK8VA16_1;
	wire w_dff_A_FM70XG8Q0_2;
	wire w_dff_A_5HkoReu22_2;
	wire w_dff_A_8YKp4dCs0_2;
	wire w_dff_A_PdafN9kM7_2;
	wire w_dff_A_tSoASTp51_2;
	wire w_dff_A_l3SVPDTu0_2;
	wire w_dff_A_NCeIZyn30_2;
	wire w_dff_A_c33zlPMx0_2;
	wire w_dff_A_CKntm3vl8_2;
	wire w_dff_A_Pbl6qVni4_2;
	wire w_dff_A_4ukLVA8O8_1;
	wire w_dff_A_8FvYFgJ17_1;
	wire w_dff_A_cymLraMl8_1;
	wire w_dff_A_APp8NyV30_1;
	wire w_dff_A_vADtSfHk0_1;
	wire w_dff_A_iB6LAnTI1_1;
	wire w_dff_A_C60DUzXr7_1;
	wire w_dff_A_CP8EoBFH8_1;
	wire w_dff_A_L2OZaSFY0_1;
	wire w_dff_A_yp4yISs39_1;
	wire w_dff_A_ChpFXZM95_1;
	wire w_dff_A_cLxXia6N4_2;
	wire w_dff_A_BlkVTWEQ9_2;
	wire w_dff_A_WIcn31uy0_2;
	wire w_dff_A_6zlKOZOd4_2;
	wire w_dff_B_ScrxC0ex8_3;
	wire w_dff_B_bF9HSW5h6_3;
	wire w_dff_B_iV8XZhOK8_3;
	wire w_dff_B_IgwPsuVZ1_3;
	wire w_dff_B_pAHPjq7V4_3;
	wire w_dff_B_7mfdTIcv8_3;
	wire w_dff_B_bDR0fVtB4_3;
	wire w_dff_B_3WtelaWZ0_3;
	wire w_dff_B_1YMFOaP55_3;
	wire w_dff_A_uKSr5MXa6_0;
	wire w_dff_A_pPMSWfET9_1;
	wire w_dff_B_wjVMUX9z6_1;
	wire w_dff_B_F1BdJIRn7_1;
	wire w_dff_A_J7RpXy9j0_0;
	wire w_dff_A_B2b2QXRq5_0;
	wire w_dff_A_U73T2Cer5_0;
	wire w_dff_A_w39mU8Y99_0;
	wire w_dff_A_m15o0S1P9_0;
	wire w_dff_A_mcMP1zUM8_0;
	wire w_dff_A_zjECLO450_0;
	wire w_dff_A_aM0peksZ5_0;
	wire w_dff_A_FQZO09FO5_0;
	wire w_dff_A_Spd7vZn46_0;
	wire w_dff_A_bQitdwoY1_0;
	wire w_dff_A_oThGbyep6_0;
	wire w_dff_A_BZXl5qNo8_0;
	wire w_dff_A_DR3dhzZL6_0;
	wire w_dff_A_0X6f479c5_0;
	wire w_dff_A_AN4zE28N9_0;
	wire w_dff_A_M3BwlCt59_0;
	wire w_dff_A_RaZXe41y5_0;
	wire w_dff_A_ZTLypPDO1_0;
	wire w_dff_A_557w5x5b3_0;
	wire w_dff_A_70LyU2fl4_0;
	wire w_dff_A_ExNRHowj8_0;
	wire w_dff_A_9CG4UPxr9_1;
	wire w_dff_A_V1YRyjog0_1;
	wire w_dff_A_NCDTHPr95_1;
	wire w_dff_A_wIyHRV9x1_1;
	wire w_dff_A_zYyz2T3b6_1;
	wire w_dff_A_Jq3nLSms4_1;
	wire w_dff_A_SfRM7CcV4_1;
	wire w_dff_A_ouvJbN4a0_1;
	wire w_dff_A_F4a1JVaO5_1;
	wire w_dff_A_FjZ8h4rR6_1;
	wire w_dff_A_qxidpLW09_1;
	wire w_dff_A_EXoqS4CX2_2;
	wire w_dff_A_ZtjjC1cr6_1;
	wire w_dff_A_yQpYbEpp5_2;
	wire w_dff_A_stD9tdsP3_0;
	wire w_dff_A_GzQHRemz8_0;
	wire w_dff_A_q2xxL2809_0;
	wire w_dff_A_wjn5NGJL4_0;
	wire w_dff_A_3vHb5jwq0_0;
	wire w_dff_A_BxOZloTC5_0;
	wire w_dff_A_d2LAGOai2_0;
	wire w_dff_A_gKJA16UU5_0;
	wire w_dff_A_4c45Rt3G2_0;
	wire w_dff_A_7f1V6vuB5_0;
	wire w_dff_A_IdcioEF45_0;
	wire w_dff_A_NXCW0Peo0_0;
	wire w_dff_A_cKVgP91G6_0;
	wire w_dff_A_Rr3erOfF6_0;
	wire w_dff_A_I5pOKBT10_0;
	wire w_dff_A_rKht7d1D0_0;
	wire w_dff_A_EOyZ921T3_0;
	wire w_dff_A_eP5pG42G3_0;
	wire w_dff_A_m5UgHlOP8_0;
	wire w_dff_A_BIn5dbuA0_0;
	wire w_dff_A_ZrCBTGC77_0;
	wire w_dff_A_xo76DDLe0_0;
	wire w_dff_A_e2DMmeF93_0;
	wire w_dff_B_5VWJlEk10_1;
	wire w_dff_B_FKUbdl895_1;
	wire w_dff_B_GhtElLy78_1;
	wire w_dff_B_N1ppBTzP7_1;
	wire w_dff_B_qaJaVZEb7_1;
	wire w_dff_B_DPx4D44O9_1;
	wire w_dff_B_MIPrLEAQ4_1;
	wire w_dff_B_2p7NKM7G4_1;
	wire w_dff_B_W4eb44Fa9_1;
	wire w_dff_B_WueJfSvG9_1;
	wire w_dff_B_i02qVWdV5_1;
	wire w_dff_B_tz9ImYf91_1;
	wire w_dff_B_kFRza5023_1;
	wire w_dff_B_Jw1xMxJU9_1;
	wire w_dff_B_rGCXZjog7_1;
	wire w_dff_B_A6VkFRSM6_1;
	wire w_dff_B_7zLHV44n1_1;
	wire w_dff_B_vVmKJpte0_1;
	wire w_dff_B_JxXsnwWw9_1;
	wire w_dff_B_AvTLxa0U9_1;
	wire w_dff_B_0COEn1EF5_1;
	wire w_dff_B_JZhC67786_1;
	wire w_dff_B_4w8ijg4L1_1;
	wire w_dff_A_XHd2QwV55_1;
	wire w_dff_A_Ap4mMjKA8_1;
	wire w_dff_A_v0A9eA911_1;
	wire w_dff_A_ysOOM7QB4_1;
	wire w_dff_A_Ka0TaOuV2_1;
	wire w_dff_A_mmrxd1oL7_1;
	wire w_dff_A_6bNMblGB6_1;
	wire w_dff_A_xji6pgNy8_1;
	wire w_dff_A_ToTuOMhx6_1;
	wire w_dff_A_6ZjksA0e1_1;
	wire w_dff_A_bPTvEwAl5_1;
	wire w_dff_A_tUZ1kFg80_1;
	wire w_dff_A_AzxWRYBH5_1;
	wire w_dff_A_MADeFKk91_1;
	wire w_dff_A_HSeYYdKz2_2;
	wire w_dff_A_vIcfKhgF2_2;
	wire w_dff_A_lQAzILS92_2;
	wire w_dff_A_vcWsDHm01_2;
	wire w_dff_A_N3rKhFR06_2;
	wire w_dff_A_kkjVur1N4_2;
	wire w_dff_A_vpbSd4Xr2_2;
	wire w_dff_A_UbJhJIwu0_2;
	wire w_dff_A_5Lr90UL94_2;
	wire w_dff_A_cFnCmMlb6_2;
	wire w_dff_A_duCczTxM6_1;
	wire w_dff_A_vsdwndrL6_1;
	wire w_dff_A_DnrT2OXK6_1;
	wire w_dff_A_oUqq3q7g6_1;
	wire w_dff_A_BPJPEmzi0_1;
	wire w_dff_A_Ej2ttc3v6_1;
	wire w_dff_A_o4OMuCUz2_1;
	wire w_dff_A_YB9OgIea1_1;
	wire w_dff_A_3VItfUrT1_1;
	wire w_dff_A_A304rUl82_1;
	wire w_dff_A_DhjotKiY6_1;
	wire w_dff_A_BhU2XX7h7_2;
	wire w_dff_A_2niEqCLp7_2;
	wire w_dff_A_YhQiCBCf8_2;
	wire w_dff_A_8CdQoD6j4_2;
	wire w_dff_A_GJS3iESA2_2;
	wire w_dff_B_YU5aFbwY8_3;
	wire w_dff_B_mASZFfYi0_3;
	wire w_dff_B_X7VLNaWq3_3;
	wire w_dff_B_QCV7Orfh1_3;
	wire w_dff_B_v84117wn9_3;
	wire w_dff_B_KIsqCmnf9_3;
	wire w_dff_B_YNEIxzyE8_3;
	wire w_dff_B_QnYnZjV90_3;
	wire w_dff_B_LKKyFNdM0_3;
	wire w_dff_A_rTzxTR3f9_0;
	wire w_dff_A_ghHCOaPZ1_0;
	wire w_dff_A_y0stXhZv5_1;
	wire w_dff_B_6890W6Pk6_1;
	wire w_dff_B_zD5UW9OE9_1;
	wire w_dff_A_Md6L4ZLk1_0;
	wire w_dff_A_L1rL8Lnv3_0;
	wire w_dff_A_qRNKc1yt7_0;
	wire w_dff_A_ePbmOZq23_0;
	wire w_dff_A_h4WNevPM8_0;
	wire w_dff_A_4BdJor4m2_0;
	wire w_dff_A_AiDyksuY8_0;
	wire w_dff_A_LiFeRp1E3_0;
	wire w_dff_A_MccVLTGR2_0;
	wire w_dff_A_FOVAUchP1_0;
	wire w_dff_A_AMohUKfL5_0;
	wire w_dff_A_xy8G4voT8_0;
	wire w_dff_A_EOr0CDKt2_0;
	wire w_dff_A_cDeiVApS6_0;
	wire w_dff_A_7OK8rxKQ2_0;
	wire w_dff_A_8K67Gti73_0;
	wire w_dff_A_w9dg7Net7_0;
	wire w_dff_A_TEtlqzdT3_0;
	wire w_dff_A_8HZgfnTa5_0;
	wire w_dff_A_mwdF4tvc7_0;
	wire w_dff_A_hthhEKpR5_0;
	wire w_dff_A_gPRdKgN45_0;
	wire w_dff_A_wt8bNgyy7_1;
	wire w_dff_A_A6De25d65_1;
	wire w_dff_A_OdmbJE6u6_1;
	wire w_dff_A_2W0nE7DX9_1;
	wire w_dff_A_HwNHOzNl1_1;
	wire w_dff_A_VBKp2dHu3_1;
	wire w_dff_A_txW4Kzme7_1;
	wire w_dff_A_1xkcgrRy6_1;
	wire w_dff_A_y6gLe14R0_1;
	wire w_dff_B_YuQ5o83W9_2;
	wire w_dff_A_rrKM09fd4_1;
	wire w_dff_A_a1NFrYxL3_1;
	wire w_dff_A_oHlGz0YR3_2;
	wire w_dff_A_98uwd9An2_1;
	wire w_dff_A_N5K4KyUj0_2;
	wire w_dff_A_rdeyPKAs0_0;
	wire w_dff_A_rJ4BELuO9_0;
	wire w_dff_A_QsjLx9Ce7_0;
	wire w_dff_A_C9GsvAJa7_0;
	wire w_dff_A_y1xvDWAF2_0;
	wire w_dff_A_tO0Qrx1f1_0;
	wire w_dff_A_IEu0Uf5u3_0;
	wire w_dff_A_oBHPoYYs8_0;
	wire w_dff_A_k35eJEDi1_0;
	wire w_dff_A_MsesAbzI5_0;
	wire w_dff_A_TAEROzuT5_0;
	wire w_dff_A_ATy3qVdy1_0;
	wire w_dff_A_oHE4udjl1_0;
	wire w_dff_A_tAkLuTeL3_0;
	wire w_dff_A_MFrG6Vnt9_0;
	wire w_dff_A_j6HF3K6N8_0;
	wire w_dff_A_bPPJTE1Z3_0;
	wire w_dff_A_jyR1jeXn2_0;
	wire w_dff_A_rfIPd6nx3_0;
	wire w_dff_A_RSZ9pChh2_0;
	wire w_dff_A_ie7Z40Gz9_0;
	wire w_dff_A_ZPALRbNc1_0;
	wire w_dff_A_M6dwhNZe0_0;
	wire w_dff_B_bMIbFn0F5_1;
	wire w_dff_B_Oa9qd6IH4_1;
	wire w_dff_B_wGu4CYYp9_1;
	wire w_dff_B_Ue4dzxzn0_1;
	wire w_dff_B_ELSlJ2Fh7_1;
	wire w_dff_B_TnFwnLhE0_1;
	wire w_dff_B_0Mqoad4x4_1;
	wire w_dff_B_ltrxup4S5_1;
	wire w_dff_B_5LAFverN7_1;
	wire w_dff_B_JCr0poLX2_1;
	wire w_dff_B_5G8zQwIv0_1;
	wire w_dff_B_fP0jmasL8_1;
	wire w_dff_B_AB3Z6gZY9_1;
	wire w_dff_B_N9p2ONu75_1;
	wire w_dff_B_6uQeOPUq7_1;
	wire w_dff_B_uW0c6eat7_1;
	wire w_dff_B_K7gGYNGh6_1;
	wire w_dff_B_e9N9hQB34_1;
	wire w_dff_B_yBPMgex56_1;
	wire w_dff_B_EJ1vIkfj9_1;
	wire w_dff_B_3Pnvo5Wy4_1;
	wire w_dff_B_yxl5bIgC1_1;
	wire w_dff_B_OFoLb81D1_1;
	wire w_dff_B_BtjNFnQ62_1;
	wire w_dff_B_7zbOjT482_1;
	wire w_dff_B_X3Q2TPw86_1;
	wire w_dff_B_VBQ2ByaR2_1;
	wire w_dff_B_HP4pVqIo7_1;
	wire w_dff_B_szQD7lG23_1;
	wire w_dff_B_Wk9oLYPq2_1;
	wire w_dff_B_J4crlOi21_1;
	wire w_dff_B_d289MB6R7_1;
	wire w_dff_B_9qFjxQSI4_1;
	wire w_dff_B_lFXW8lHy0_1;
	wire w_dff_B_3aozawya1_1;
	wire w_dff_B_35hDRlGt3_1;
	wire w_dff_B_g8DzMmqT5_1;
	wire w_dff_B_1V2d6Ptw3_1;
	wire w_dff_B_VaCCbFQW1_1;
	wire w_dff_B_3lYlaJqe7_1;
	wire w_dff_B_vErUsyA04_1;
	wire w_dff_B_v4T5gsVC4_1;
	wire w_dff_B_0kJnOtNr6_1;
	wire w_dff_B_2cHRsFbU8_1;
	wire w_dff_B_yScOK9ru2_1;
	wire w_dff_A_SlYv8LDR1_0;
	wire w_dff_A_ItebSVhY6_0;
	wire w_dff_A_MdmZpCRp5_0;
	wire w_dff_A_F3uKWVcV2_0;
	wire w_dff_A_qhnKv03l0_0;
	wire w_dff_A_jyFXtZNu1_0;
	wire w_dff_A_a3kbefkD9_0;
	wire w_dff_A_wDfwGPd80_0;
	wire w_dff_A_jqIEugti6_0;
	wire w_dff_A_Ioz0d5Nt4_0;
	wire w_dff_A_wYl1bAxT8_0;
	wire w_dff_A_yo3MvZQ20_0;
	wire w_dff_A_CA7cmmFD8_0;
	wire w_dff_A_jAKgpXcQ3_0;
	wire w_dff_A_GY8z1wY53_0;
	wire w_dff_A_hBs0JYMO5_1;
	wire w_dff_A_E00msF9S8_1;
	wire w_dff_A_KBrCNoyH2_1;
	wire w_dff_A_hQt0O5c47_1;
	wire w_dff_A_s4HPvbzB5_1;
	wire w_dff_A_9XR28cZQ0_1;
	wire w_dff_A_SaluuUvc8_1;
	wire w_dff_A_IBgY35Ba8_1;
	wire w_dff_A_LcIc8VQ40_1;
	wire w_dff_A_0fxBTHVS6_1;
	wire w_dff_A_Sx4BI8977_1;
	wire w_dff_A_BgW4wWCA1_1;
	wire w_dff_A_zbtyXcT68_1;
	wire w_dff_A_RXC5pQLZ0_1;
	wire w_dff_A_6q7gu6kZ5_1;
	wire w_dff_A_PvgqQlK40_1;
	wire w_dff_A_krANA6Z87_1;
	wire w_dff_A_1naFaLhF2_1;
	wire w_dff_A_Ojn0kkYc3_1;
	wire w_dff_A_LJnRnScN6_1;
	wire w_dff_A_oMXIdcBD7_1;
	wire w_dff_A_DRrznnA01_1;
	wire w_dff_A_X0KzkqqW8_1;
	wire w_dff_A_q488RTdU3_1;
	wire w_dff_A_pC6vtcTT4_1;
	wire w_dff_A_oErH0m2e9_1;
	wire w_dff_A_SmdYjCkC2_1;
	wire w_dff_A_wv8LgdWo5_1;
	wire w_dff_A_vfOOW9eV1_1;
	wire w_dff_A_OmbFbeiy7_1;
	wire w_dff_A_LPoxAlm50_1;
	wire w_dff_A_1apXy0ad4_2;
	wire w_dff_A_SjCjHrU97_2;
	wire w_dff_A_y2R6h7587_2;
	wire w_dff_A_Ra9P4r6X0_2;
	wire w_dff_A_XXSDnZKZ6_2;
	wire w_dff_A_7tYfKjwv0_2;
	wire w_dff_A_fwTHRFFT7_2;
	wire w_dff_A_kes8BGOy5_2;
	wire w_dff_A_cIKV6sB89_2;
	wire w_dff_A_tBOTIIWJ7_2;
	wire w_dff_A_uO7t2O6z3_2;
	wire w_dff_A_f4Zs8oBC4_2;
	wire w_dff_A_Whe0g9Av0_2;
	wire w_dff_A_2B1qupzO7_2;
	wire w_dff_A_jG06aDOL0_2;
	wire w_dff_A_NaB2w87d7_2;
	wire w_dff_A_Twvw7lxj4_2;
	wire w_dff_A_oewqjaCp0_2;
	wire w_dff_A_Lt74J5M05_2;
	wire w_dff_A_bFcptGNJ2_2;
	wire w_dff_A_p4nLFl8q3_1;
	wire w_dff_A_EYrLqPqr0_1;
	wire w_dff_A_mBvmh2bY5_1;
	wire w_dff_A_VRP4Ngk05_1;
	wire w_dff_A_X82o1FL83_1;
	wire w_dff_A_0lDIfkg95_1;
	wire w_dff_A_IzmYZUuV3_1;
	wire w_dff_A_VGJA1fJn7_1;
	wire w_dff_A_LMANtSHB6_1;
	wire w_dff_A_ahxEezkt2_1;
	wire w_dff_A_x6JB4o569_1;
	wire w_dff_A_2QQSaOSQ2_1;
	wire w_dff_A_AZzYQT3o6_1;
	wire w_dff_A_vp6kULU05_1;
	wire w_dff_A_MJtMi19x2_1;
	wire w_dff_A_67K9j7t85_1;
	wire w_dff_A_fFSRRVgn1_1;
	wire w_dff_A_KDQYG55A6_1;
	wire w_dff_A_oLysiJcs3_2;
	wire w_dff_A_ggRoZm195_2;
	wire w_dff_A_b0G6MoTR1_2;
	wire w_dff_A_HIL9ujgO0_2;
	wire w_dff_A_6SxZoqee7_2;
	wire w_dff_A_NxmArqPE9_2;
	wire w_dff_A_FD6LLLM71_2;
	wire w_dff_A_K6hrhoON0_2;
	wire w_dff_A_1RU6fnuX6_2;
	wire w_dff_A_zpurIaVN1_2;
	wire w_dff_A_HLISzOAQ6_2;
	wire w_dff_A_oQ6hWZ8K6_1;
	wire w_dff_A_ZqQ5dgBf9_1;
	wire w_dff_A_BCD8u8gK8_1;
	wire w_dff_A_g8SwvjE69_1;
	wire w_dff_A_L21lRDsT2_1;
	wire w_dff_A_mjSB2XIM0_1;
	wire w_dff_A_Z1j81ptQ7_1;
	wire w_dff_A_2aaxuw399_1;
	wire w_dff_A_jMxfTBlk9_1;
	wire w_dff_A_poynQU1Y6_1;
	wire w_dff_A_v8Bg2hU68_1;
	wire w_dff_A_4U0l04jV0_1;
	wire w_dff_A_u4DWv6Lg0_1;
	wire w_dff_A_eIXvyG0r8_1;
	wire w_dff_A_5RWirk279_1;
	wire w_dff_A_yECbOnJk5_1;
	wire w_dff_A_c2vrPWTn6_1;
	wire w_dff_A_odjQJDVI1_1;
	wire w_dff_A_otNrD9H20_1;
	wire w_dff_A_YA7kGA5z9_1;
	wire w_dff_A_AitZwGyh9_1;
	wire w_dff_A_2UrOsUSd1_1;
	wire w_dff_A_hgNgdS730_1;
	wire w_dff_A_8q1v2Fau8_1;
	wire w_dff_A_VwzzJvf65_0;
	wire w_dff_A_ShNaac751_0;
	wire w_dff_A_5Oz4lCsW3_0;
	wire w_dff_A_ESwHyVEX2_0;
	wire w_dff_A_ji7vJUdB3_0;
	wire w_dff_A_CS8RqFnI3_0;
	wire w_dff_A_pappRIuy5_0;
	wire w_dff_A_E009sSDJ5_0;
	wire w_dff_A_DjEPVuot6_0;
	wire w_dff_A_63qojU8U2_2;
	wire w_dff_A_RfNOAa5D4_2;
	wire w_dff_A_iZPFkH8r6_2;
	wire w_dff_A_S0IfHSAp0_2;
	wire w_dff_A_Nq2xCbnW4_2;
	wire w_dff_A_crbYARKb0_2;
	wire w_dff_A_FgkZB9Mw4_2;
	wire w_dff_A_vQ3mENBJ9_2;
	wire w_dff_A_s85UEDSu3_2;
	wire w_dff_A_ibqOQKJ08_2;
	wire w_dff_A_5jt12NCG6_2;
	wire w_dff_A_VOUGfFPN2_2;
	wire w_dff_A_KbnJfHre1_2;
	wire w_dff_A_kApJddP89_2;
	wire w_dff_A_LIRcmzzV4_2;
	wire w_dff_A_DCfos2bf9_2;
	wire w_dff_A_10iNWcyt9_2;
	wire w_dff_A_iWZg5kyo0_2;
	wire w_dff_A_DKhhC6jr6_2;
	wire w_dff_A_8Bhrdh8W6_2;
	wire w_dff_A_X8tib3Xx3_2;
	wire w_dff_A_V9AeNPX94_2;
	wire w_dff_A_773q4Ajn8_1;
	wire w_dff_A_c8B6M1fH1_1;
	wire w_dff_A_QlWRPz4U7_1;
	wire w_dff_A_nnpthrqL4_1;
	wire w_dff_A_wPmKhg8A0_1;
	wire w_dff_A_cwOmZkHW5_1;
	wire w_dff_A_M4Db9nyY5_1;
	wire w_dff_A_FJJYCpmb3_1;
	wire w_dff_A_C8UCi4yX7_1;
	wire w_dff_A_eH6uomXR6_1;
	wire w_dff_A_zfQgTGRS8_1;
	wire w_dff_A_GVWeV97E2_1;
	wire w_dff_A_OUTm0v0B0_1;
	wire w_dff_A_F960wYkX9_1;
	wire w_dff_A_JCCE42rm0_1;
	wire w_dff_A_fxVNohek0_1;
	wire w_dff_A_rrl7vplS7_1;
	wire w_dff_A_gawc5Su77_1;
	wire w_dff_A_TRFWSf9o9_1;
	wire w_dff_A_2UEpnK4m7_2;
	wire w_dff_A_acpypHIp4_2;
	wire w_dff_A_3ensXNEH3_2;
	wire w_dff_A_9GgifZZj0_2;
	wire w_dff_A_SLN9LdOC7_2;
	wire w_dff_A_EuADFi455_2;
	wire w_dff_A_taIc74Ms2_2;
	wire w_dff_A_pYmkRsUp5_2;
	wire w_dff_A_BJZnq2nh9_2;
	wire w_dff_A_GwsTqavO7_2;
	wire w_dff_A_wl56k2at9_2;
	wire w_dff_A_dqC8Jl5g8_2;
	wire w_dff_A_qhYXJhut8_2;
	wire w_dff_B_fappLODQ3_1;
	wire w_dff_B_K1eSItKk0_1;
	wire w_dff_B_f4UNuX4U5_1;
	wire w_dff_B_Xe6OwQUV0_1;
	wire w_dff_B_vltlLjBs2_1;
	wire w_dff_B_ZNPbb3Je8_1;
	wire w_dff_B_LigNWl0D7_1;
	wire w_dff_B_JxbLPvAR2_1;
	wire w_dff_B_N8ynxXMk0_1;
	wire w_dff_B_84PIClfp7_1;
	wire w_dff_B_G8uzX2zx0_1;
	wire w_dff_B_a1GkaZ6l0_1;
	wire w_dff_B_jBZI8hw18_1;
	wire w_dff_B_PqLUO8oi4_1;
	wire w_dff_B_3ubxHMpQ4_1;
	wire w_dff_B_lkcI4hR56_1;
	wire w_dff_B_OYdWE7k76_1;
	wire w_dff_B_A84Spr3i9_1;
	wire w_dff_B_dG9LJPdV7_1;
	wire w_dff_B_qKANdGMn4_1;
	wire w_dff_B_x3SmIgxL6_1;
	wire w_dff_B_Zp839Tqa8_1;
	wire w_dff_B_4pl9l5DJ3_1;
	wire w_dff_B_7KxXvuiq5_1;
	wire w_dff_B_VwMv84VU3_1;
	wire w_dff_B_AztD1pwj1_1;
	wire w_dff_B_LyzQh7MP8_1;
	wire w_dff_B_dJFA7P208_1;
	wire w_dff_B_Fq43BFwN3_1;
	wire w_dff_B_G0BVtXRn7_1;
	wire w_dff_B_kn63FJ2r7_1;
	wire w_dff_B_5Zutcn3n0_1;
	wire w_dff_B_TAinSHb54_1;
	wire w_dff_B_VLJu7GQG7_1;
	wire w_dff_B_GNgU3cM99_1;
	wire w_dff_B_kIOcZ6FJ0_1;
	wire w_dff_B_3mwH3La20_1;
	wire w_dff_B_pWpPGTZd5_1;
	wire w_dff_B_tT7GL0eE8_1;
	wire w_dff_B_vevqLO3x7_1;
	wire w_dff_B_vQ9pZ3jq7_1;
	wire w_dff_B_aOWQD9044_1;
	wire w_dff_B_r5AAnhzs6_1;
	wire w_dff_B_lPnA7KxI1_1;
	wire w_dff_B_TvwtaERu1_1;
	wire w_dff_B_uMayVPtM2_0;
	wire w_dff_B_YehyMLQ18_0;
	wire w_dff_B_oyrNO1rC6_0;
	wire w_dff_B_Pzqkmj7s0_0;
	wire w_dff_B_l9nXCu7R0_0;
	wire w_dff_B_VuH0LG3Y0_0;
	wire w_dff_B_7CLkLhNS4_0;
	wire w_dff_B_dZfUUkFQ9_0;
	wire w_dff_B_R0ph8LWv6_0;
	wire w_dff_B_ihydbqsS0_0;
	wire w_dff_B_1uf5h5F70_0;
	wire w_dff_B_d88tFYTL8_0;
	wire w_dff_B_t3YGfFxZ4_0;
	wire w_dff_B_KLvwqxyX5_0;
	wire w_dff_B_seZyezCh5_0;
	wire w_dff_B_dJcJZI5n5_0;
	wire w_dff_B_wpWc3Yfc5_0;
	wire w_dff_B_AR7NSALd2_0;
	wire w_dff_B_tshotWrx4_0;
	wire w_dff_B_SX1hBGvL9_0;
	wire w_dff_B_Vu0RJXKf9_0;
	wire w_dff_B_n5BF50uh8_0;
	wire w_dff_B_Az16hyfc7_0;
	wire w_dff_B_HzbJxaAG6_0;
	wire w_dff_B_wexuEVra7_0;
	wire w_dff_B_oCa9GmqI7_0;
	wire w_dff_B_Xefk6Yl04_0;
	wire w_dff_B_LnFfZrMQ4_0;
	wire w_dff_B_vCCTPlxH9_1;
	wire w_dff_B_KY4oClPQ5_1;
	wire w_dff_B_HKApNhrR4_1;
	wire w_dff_A_ScLRp0dH0_0;
	wire w_dff_B_IuHkOkDX2_1;
	wire w_dff_B_yyfaiPDj6_1;
	wire w_dff_A_ZpN0xOKU4_1;
	wire w_dff_B_8Xf7QnmY4_0;
	wire w_dff_A_S8jCp1lV4_0;
	wire w_dff_B_4uGaUG2h6_1;
	wire w_dff_A_JMj54jpY1_0;
	wire w_dff_B_SB3eUVwo7_2;
	wire w_dff_A_bqOqBG597_0;
	wire w_dff_A_0rgalY9k1_0;
	wire w_dff_A_PXTYXeMl1_0;
	wire w_dff_B_EY5P9kkJ0_1;
	wire w_dff_B_xQ7tHhqd7_1;
	wire w_dff_B_3bgIAedx2_1;
	wire w_dff_A_F6B7u8qa1_1;
	wire w_dff_B_TnwyGcai3_1;
	wire w_dff_B_Ifi5KaPP0_1;
	wire w_dff_A_ngYc9BaC7_1;
	wire w_dff_B_z7gTYVop1_1;
	wire w_dff_A_V7FGggCU2_0;
	wire w_dff_A_yTmRByLd0_0;
	wire w_dff_A_aUEeXtDh7_0;
	wire w_dff_A_ZGbPL6sO7_1;
	wire w_dff_A_xCDea2wl3_1;
	wire w_dff_A_gJgdEIrO5_1;
	wire w_dff_A_QtdHhHKE0_1;
	wire w_dff_A_8mDJimVz1_1;
	wire w_dff_A_FCBxGdyh3_1;
	wire w_dff_A_h9R3Tg6B4_1;
	wire w_dff_A_Bn8s0z5C4_1;
	wire w_dff_A_qWGh3QJT3_1;
	wire w_dff_A_acbRl9gy2_1;
	wire w_dff_A_GpYsJDvJ6_1;
	wire w_dff_A_Y5kv7rC74_1;
	wire w_dff_B_99f1ywRJ4_0;
	wire w_dff_A_ZotBMQ0D5_0;
	wire w_dff_A_TmQHv6xl0_0;
	wire w_dff_B_KKXQIs3M6_0;
	wire w_dff_B_03kMr17E1_0;
	wire w_dff_B_c3XXmCf30_0;
	wire w_dff_B_pC6Oo3Vw3_1;
	wire w_dff_B_BwKl9oSn1_1;
	wire w_dff_B_HMWdFj7t1_1;
	wire w_dff_A_jOpFjveP9_0;
	wire w_dff_A_0WBcNEnh6_0;
	wire w_dff_A_Colzfz4w2_0;
	wire w_dff_A_2gaaYJ2z9_0;
	wire w_dff_A_pKK52SXc3_0;
	wire w_dff_A_zCWqs08e9_0;
	wire w_dff_A_ZDmExVea5_0;
	wire w_dff_A_Nh5iaij37_0;
	wire w_dff_B_gkOm9f2C8_1;
	wire w_dff_B_X7h3zKJR7_1;
	wire w_dff_B_HFXHnHTq0_0;
	wire w_dff_B_YmCA8NpP5_0;
	wire w_dff_A_fLKCUw2Z1_0;
	wire w_dff_B_CGHTI8A53_1;
	wire w_dff_A_qr3O2Jyf8_2;
	wire w_dff_A_3lMUSRFd5_2;
	wire w_dff_A_pp4HwyNl2_0;
	wire w_dff_A_hISlCyLZ4_0;
	wire w_dff_A_PUUWdHUJ7_0;
	wire w_dff_A_Jhn4XrRk4_0;
	wire w_dff_A_TizUnkPX5_1;
	wire w_dff_B_8fAdz1ZW7_3;
	wire w_dff_B_XUuxerAk5_3;
	wire w_dff_A_SYi6c45J6_1;
	wire w_dff_A_3MEM3U4V7_1;
	wire w_dff_A_3umru07q0_1;
	wire w_dff_A_NHz2SRfK7_1;
	wire w_dff_A_qHr140EL7_1;
	wire w_dff_A_GwQxQH0o0_1;
	wire w_dff_A_pu0aBU7w3_2;
	wire w_dff_A_B2AbRm9C6_2;
	wire w_dff_A_RzH3MoT43_2;
	wire w_dff_A_UnQODbXq5_2;
	wire w_dff_A_QAGcJSPV5_2;
	wire w_dff_A_fdnYTmS70_2;
	wire w_dff_A_ioamGLlq1_2;
	wire w_dff_A_4Q6uc5GK7_1;
	wire w_dff_A_dsFZ2h5H1_1;
	wire w_dff_A_JL4ZPdIW2_1;
	wire w_dff_A_NFvJFWBi9_1;
	wire w_dff_A_2ddUJsYP3_1;
	wire w_dff_A_zHayOKWN5_1;
	wire w_dff_A_3tylgieY3_2;
	wire w_dff_A_qBVbiEbx0_2;
	wire w_dff_A_XOM3sFug4_2;
	wire w_dff_A_5WLf0liM1_0;
	wire w_dff_B_T4kygeEA9_1;
	wire w_dff_A_O4Bg95WV8_0;
	wire w_dff_B_1KSxEyng2_1;
	wire w_dff_B_xjS2fJOz2_1;
	wire w_dff_B_g9698oLR9_1;
	wire w_dff_B_CXq2RJea6_1;
	wire w_dff_B_fuURMbT48_1;
	wire w_dff_A_8KmR0YJP9_2;
	wire w_dff_A_snwGPB9Z3_2;
	wire w_dff_A_E2gla9Im8_2;
	wire w_dff_A_lvIaQO0g4_2;
	wire w_dff_A_8dtaMtdk8_2;
	wire w_dff_A_L4yrxRrg8_2;
	wire w_dff_A_PLnNkKAR6_2;
	wire w_dff_A_tPGViu0P0_2;
	wire w_dff_A_LiZCO5hy1_2;
	wire w_dff_A_38fXQmRj4_2;
	wire w_dff_A_JJd7wOE12_2;
	wire w_dff_A_NSJ5nVXs1_2;
	wire w_dff_A_slkS1ByX2_2;
	wire w_dff_A_N3Gq0osR5_2;
	wire w_dff_A_68PoRUC35_2;
	wire w_dff_A_wo7kR2uM2_1;
	wire w_dff_A_yLioJ1nj9_1;
	wire w_dff_A_lBhsoe5B3_1;
	wire w_dff_A_QNWnC9vh2_1;
	wire w_dff_A_xVD02jHt7_1;
	wire w_dff_A_kgVQSWxH0_1;
	wire w_dff_A_0fIJiKcG7_1;
	wire w_dff_A_jtqU0hGe6_1;
	wire w_dff_A_54lJdxHT6_1;
	wire w_dff_A_4MuFKhJy2_1;
	wire w_dff_B_9CdaUsTE7_1;
	wire w_dff_B_IcLk55ca2_1;
	wire w_dff_B_2Y962Pvs2_1;
	wire w_dff_B_Qoa6Ht6s8_1;
	wire w_dff_B_S0q4jkJ69_1;
	wire w_dff_B_7ueIVrlP4_1;
	wire w_dff_B_mAlA7HAG8_1;
	wire w_dff_A_mfsUWL0M9_1;
	wire w_dff_B_0iqja61s8_1;
	wire w_dff_B_EKjZM2YP1_1;
	wire w_dff_B_8z1ZQthU8_1;
	wire w_dff_B_WzlzO9Pe6_1;
	wire w_dff_B_xABjFLal2_1;
	wire w_dff_B_X11dDHA70_1;
	wire w_dff_B_N0rTAIrb9_1;
	wire w_dff_A_ls8UL0Zm0_1;
	wire w_dff_A_IYJMrDp93_1;
	wire w_dff_A_iWDqtKCR1_0;
	wire w_dff_A_wS2vt67i1_0;
	wire w_dff_A_2ZtELZvn1_0;
	wire w_dff_A_12ZkINdP0_0;
	wire w_dff_A_z7p6YUjr6_1;
	wire w_dff_A_TJs1W6DT4_1;
	wire w_dff_A_Gva3RcoY4_2;
	wire w_dff_B_8YMo3sLn6_3;
	wire w_dff_A_eNIehFkN6_0;
	wire w_dff_A_9sijSR7X7_0;
	wire w_dff_A_YeTVb28I2_0;
	wire w_dff_A_uj2YxGOe0_1;
	wire w_dff_A_uacR1U299_1;
	wire w_dff_A_7rkIrt1C7_2;
	wire w_dff_B_PgG8jdQ65_3;
	wire w_dff_B_G1Da8Jhw2_3;
	wire w_dff_B_Z2ESZr7E7_3;
	wire w_dff_B_FP36ZvEP7_3;
	wire w_dff_B_H0CS5pZQ4_3;
	wire w_dff_B_3ffLWUqT4_3;
	wire w_dff_B_nUYSVcto3_3;
	wire w_dff_B_Fvxerrtk9_3;
	wire w_dff_B_sdwmjEXH9_3;
	wire w_dff_B_1mfQGzjy0_3;
	wire w_dff_A_rBMiAk2D1_0;
	wire w_dff_A_OCUCIsPn8_0;
	wire w_dff_A_Rs7jDHPV2_0;
	wire w_dff_A_GzMljIXB9_0;
	wire w_dff_A_AbNsvuMK8_0;
	wire w_dff_A_LcXRCDil6_0;
	wire w_dff_A_kBWWMt8I3_0;
	wire w_dff_A_5Rwlu8WZ7_0;
	wire w_dff_A_J0FTVxWY9_0;
	wire w_dff_A_mkjfvBAA2_0;
	wire w_dff_A_xNidbHy21_0;
	wire w_dff_A_HzJQC4BY7_0;
	wire w_dff_A_Jsb5G67L3_0;
	wire w_dff_A_3XgOyV4A3_1;
	wire w_dff_A_l5Fp4qqx5_1;
	wire w_dff_A_RpzViQAF7_1;
	wire w_dff_A_FKCEAtMd9_1;
	wire w_dff_A_4leJHROL5_1;
	wire w_dff_A_kt02p7lV7_1;
	wire w_dff_A_FcLCn6tK6_1;
	wire w_dff_A_tRzY0CQz2_1;
	wire w_dff_A_0oDtY7i71_1;
	wire w_dff_A_ibm6KBV90_1;
	wire w_dff_A_xGYv2QMQ1_0;
	wire w_dff_B_96UzNQdT7_0;
	wire w_dff_B_T4ChUrjp5_0;
	wire w_dff_A_c6y1Byqp4_0;
	wire w_dff_A_akJRuCx35_0;
	wire w_dff_A_TG9rKCVs5_0;
	wire w_dff_B_dxrmcj3p8_2;
	wire w_dff_A_BCOMpbI92_0;
	wire w_dff_A_jIE75rIy5_0;
	wire w_dff_A_DlOB61Du6_0;
	wire w_dff_A_fl2XX5NO3_1;
	wire w_dff_A_KzDCsPxR0_1;
	wire w_dff_A_CuvyOiKi4_1;
	wire w_dff_A_CseopRmD1_1;
	wire w_dff_A_DtV5yOsa7_1;
	wire w_dff_A_Av5iEvP98_1;
	wire w_dff_A_cY01WQiF5_1;
	wire w_dff_A_8SolGUlR1_1;
	wire w_dff_A_MaZmCqmi6_0;
	wire w_dff_A_7DuDT1AJ7_0;
	wire w_dff_A_y04Tg1jh5_0;
	wire w_dff_A_YnXvQpkT4_0;
	wire w_dff_A_KcQBLqEE2_2;
	wire w_dff_A_lxg9sKrs5_2;
	wire w_dff_A_ohMqcqoZ8_1;
	wire w_dff_A_IkZ0w3dF1_1;
	wire w_dff_A_LIpZI4sY9_1;
	wire w_dff_A_h9jhfxll5_1;
	wire w_dff_A_1cjKdCl93_1;
	wire w_dff_B_L78YjEUY2_1;
	wire w_dff_B_6s7BJUn44_1;
	wire w_dff_A_bMOUi0UJ9_1;
	wire w_dff_A_mU1xbz8d0_1;
	wire w_dff_A_89hbxUXa5_1;
	wire w_dff_A_9WVpNVBm1_1;
	wire w_dff_A_sinFkYgd5_1;
	wire w_dff_A_Y2fP7vZz7_1;
	wire w_dff_A_QbkPiTFN8_1;
	wire w_dff_B_asLk4WND6_0;
	wire w_dff_B_tschl8w45_1;
	wire w_dff_A_gRwoKJ1I1_2;
	wire w_dff_A_9Xax7Uze0_1;
	wire w_dff_A_WFQWTIZ04_1;
	wire w_dff_A_YhHvhUHd6_1;
	wire w_dff_A_S77Krj036_1;
	wire w_dff_A_ebeDXyY83_2;
	wire w_dff_A_D8d91TvS3_2;
	wire w_dff_A_UsOjqMgw6_2;
	wire w_dff_A_lcGgPAjg9_2;
	wire w_dff_A_xFdiiL3z1_0;
	wire w_dff_A_BrKvvSPn1_0;
	wire w_dff_B_r3BFdL1o3_3;
	wire w_dff_A_qKiqqAVL5_0;
	wire w_dff_B_xOOQgFa32_1;
	wire w_dff_B_IrD5C1yu8_1;
	wire w_dff_A_Xsngfe2U3_0;
	wire w_dff_A_f4tHy0gm6_0;
	wire w_dff_B_zrNIoY7t3_2;
	wire w_dff_A_exMnkZjk4_0;
	wire w_dff_A_fwH1ofpW3_0;
	wire w_dff_A_U2B1WQkS2_0;
	wire w_dff_A_ktMtPHfW7_1;
	wire w_dff_A_LtTTofiA0_1;
	wire w_dff_A_EbD5XZ6A1_1;
	wire w_dff_A_5E871zXd0_1;
	wire w_dff_A_jkidX6wY6_1;
	wire w_dff_A_FpBvAnXV4_1;
	wire w_dff_A_hVwjUmak5_1;
	wire w_dff_A_gEJ9SdA75_2;
	wire w_dff_A_Uo8RRHtf5_2;
	wire w_dff_A_JuVocacq3_2;
	wire w_dff_A_GgqagvSJ3_2;
	wire w_dff_A_E5nnNKxj8_2;
	wire w_dff_B_J7QSLHkv8_0;
	wire w_dff_B_G0FqcR0X5_1;
	wire w_dff_A_etQq017Q2_0;
	wire w_dff_A_kGtQubRU4_1;
	wire w_dff_B_h14bxRSR8_1;
	wire w_dff_A_UPDBQr5m9_0;
	wire w_dff_A_xmHMGbPn5_1;
	wire w_dff_A_1wofKjqD7_1;
	wire w_dff_B_Ye6HFRXg6_1;
	wire w_dff_A_MJ0ViibJ4_0;
	wire w_dff_A_ebIdPORu4_0;
	wire w_dff_A_5elyxUXx2_2;
	wire w_dff_A_HMrfA5Gf4_0;
	wire w_dff_A_pQe7xHr40_0;
	wire w_dff_A_nGDxQYAn0_0;
	wire w_dff_A_iHYFifiN4_2;
	wire w_dff_A_qeIdu1Xg2_0;
	wire w_dff_A_jmzSzmoB4_1;
	wire w_dff_A_SNlAwwOi8_2;
	wire w_dff_A_5ATc7Gsn9_0;
	wire w_dff_A_u6gIaMjr6_0;
	wire w_dff_A_LAEMmbVG5_0;
	wire w_dff_A_0Z1fpFhw9_2;
	wire w_dff_A_h2orIroB3_2;
	wire w_dff_A_uz8yns7j3_2;
	wire w_dff_A_wogrT4di4_0;
	wire w_dff_A_qDepDr3V9_0;
	wire w_dff_A_hItFPknl1_0;
	wire w_dff_A_FPSHAf153_1;
	wire w_dff_A_tpYJbV0X3_1;
	wire w_dff_A_r9ppHhem0_2;
	wire w_dff_A_vNWGVL5O1_0;
	wire w_dff_A_jcIciAi55_2;
	wire w_dff_B_43Qwqhk89_3;
	wire w_dff_A_y5zcxQJw1_0;
	wire w_dff_A_58qlD1fI5_0;
	wire w_dff_A_RzdvU1OF3_0;
	wire w_dff_A_jc1tYchS5_1;
	wire w_dff_A_lp7GHm1F6_1;
	wire w_dff_A_5oDTPYdf1_1;
	wire w_dff_A_yoxJaAYq4_1;
	wire w_dff_A_nbuYs9md5_1;
	wire w_dff_A_w06BWhO72_1;
	wire w_dff_A_toLwCWIm7_2;
	wire w_dff_A_4lpIsodn8_2;
	wire w_dff_A_jo6hae3s0_2;
	wire w_dff_A_95nW45hR3_1;
	wire w_dff_A_Ud1hYCRi0_1;
	wire w_dff_A_qV2cdtfx4_1;
	wire w_dff_A_8hthiOcC1_1;
	wire w_dff_A_mwgLu1SD4_1;
	wire w_dff_A_lCkwKWrU1_1;
	wire w_dff_A_M4yv3f1H0_1;
	wire w_dff_A_I7cHtpOf1_1;
	wire w_dff_A_XKG0JAaY6_1;
	wire w_dff_A_pdF4pMba5_1;
	wire w_dff_A_ZNLjUrh03_1;
	wire w_dff_A_RfHlSoqf7_0;
	wire w_dff_A_PQmDPWnJ9_0;
	wire w_dff_A_3n8RWLgq4_0;
	wire w_dff_A_khKlBzin5_2;
	wire w_dff_A_zBOEPcfw3_1;
	wire w_dff_A_qwX6CVHe2_1;
	wire w_dff_A_A6QyrXHa2_1;
	wire w_dff_A_p4Fayc1v9_1;
	wire w_dff_A_pbft6EN75_1;
	wire w_dff_A_v9ao2i6o1_1;
	wire w_dff_A_uqg8fGWl4_1;
	wire w_dff_A_XfTKPgdB9_1;
	wire w_dff_A_1awB07r12_1;
	wire w_dff_B_57G6NsdX4_0;
	wire w_dff_A_R1RIDmXh3_1;
	wire w_dff_A_F8Uk3U9y7_1;
	wire w_dff_A_zFfp6bVg0_2;
	wire w_dff_A_VICh85vW4_0;
	wire w_dff_A_R6CvotoX6_0;
	wire w_dff_A_jKyAwvkP8_0;
	wire w_dff_A_GN83aTc42_0;
	wire w_dff_A_10AtPci18_2;
	wire w_dff_A_NJpbWQ6H2_2;
	wire w_dff_A_EIhQxOxi1_0;
	wire w_dff_A_qJsf05Up1_0;
	wire w_dff_A_wYSDX8fS2_0;
	wire w_dff_A_VOUIoQCP5_0;
	wire w_dff_A_TAJot7FE7_0;
	wire w_dff_A_uISgwoQ22_0;
	wire w_dff_A_oTkjMKGO6_0;
	wire w_dff_A_9LdN4vs39_0;
	wire w_dff_A_kh43U5pn6_0;
	wire w_dff_A_4bJdu3ei3_0;
	wire w_dff_A_UvAzVEjK0_0;
	wire w_dff_A_djvkdCPF3_0;
	wire w_dff_A_ArpKi3J15_0;
	wire w_dff_A_opWE1Xsm3_0;
	wire w_dff_A_5H3EhhXK2_0;
	wire w_dff_A_AwplXlA05_0;
	wire w_dff_A_SvU9OCQG5_0;
	wire w_dff_A_PfGgEJzT3_0;
	wire w_dff_A_r73D5zJI9_0;
	wire w_dff_A_xXFR20xn1_0;
	wire w_dff_A_kn2ty5aY0_2;
	wire w_dff_A_4QZMshbv7_2;
	wire w_dff_A_0DjVm3660_2;
	wire w_dff_A_8AaK8aOG1_2;
	wire w_dff_B_OQgniS8Z0_0;
	wire w_dff_B_c7wDodW81_0;
	wire w_dff_B_dxlYHcWx4_0;
	wire w_dff_B_Ukh7m1Bv2_0;
	wire w_dff_B_7QClgarR9_0;
	wire w_dff_B_H1gZ39aE4_0;
	wire w_dff_B_d2uBp8jE2_0;
	wire w_dff_B_5OCG9Rsg8_0;
	wire w_dff_B_9qu58Pm82_0;
	wire w_dff_B_qKqzwTI43_0;
	wire w_dff_B_FNlDNXDC1_0;
	wire w_dff_B_RH52Fyov0_0;
	wire w_dff_B_iQyb6XoS3_0;
	wire w_dff_B_SkypU4MT0_0;
	wire w_dff_B_L8xjIghs4_0;
	wire w_dff_B_OnK7SI3H5_0;
	wire w_dff_B_WPf0bgdS4_0;
	wire w_dff_B_8UmPLGEf0_0;
	wire w_dff_B_UAoLTV0I0_0;
	wire w_dff_B_FRDYFa6S5_1;
	wire w_dff_B_vce812uo3_1;
	wire w_dff_B_qfHGV0D74_1;
	wire w_dff_B_efRlcB7r5_1;
	wire w_dff_B_LEQP3c7v9_1;
	wire w_dff_B_7dmBLewq7_1;
	wire w_dff_B_t6fAe9au6_1;
	wire w_dff_B_1X3yTzcg9_1;
	wire w_dff_B_6iQyRD5L9_1;
	wire w_dff_B_Nb21UJTq6_1;
	wire w_dff_A_xlkFGP9J9_2;
	wire w_dff_A_4SjY06lH7_2;
	wire w_dff_A_L7QMeyn52_1;
	wire w_dff_B_QoTvP5CI6_0;
	wire w_dff_B_kEmmUmCN9_1;
	wire w_dff_B_U1nnP5rN5_1;
	wire w_dff_B_WBi1Vhx51_1;
	wire w_dff_B_8IX8KGr32_1;
	wire w_dff_B_8cdrglPg3_1;
	wire w_dff_B_keaKlAXc1_1;
	wire w_dff_B_KfVMJ9oW4_1;
	wire w_dff_B_u1f4EHL35_0;
	wire w_dff_B_T8eDJLQt1_0;
	wire w_dff_A_Uws9P4kF7_1;
	wire w_dff_A_3trX53hq8_1;
	wire w_dff_A_QtIGU6nu1_1;
	wire w_dff_A_FyMgIb5q1_1;
	wire w_dff_A_oMSGCTfm4_1;
	wire w_dff_A_1f2BLEyN8_1;
	wire w_dff_A_1UZuqTSm6_1;
	wire w_dff_A_rUws5IQk5_1;
	wire w_dff_A_vvzJet7l9_1;
	wire w_dff_A_bID7jaFa3_1;
	wire w_dff_A_MTSappig0_1;
	wire w_dff_A_5r6h0yxY4_1;
	wire w_dff_A_qKtk3BAZ0_1;
	wire w_dff_B_06dA8gXU0_2;
	wire w_dff_A_moXGfcut3_2;
	wire w_dff_A_kxwH2KKG7_2;
	wire w_dff_A_4VevNxZE6_2;
	wire w_dff_A_MBniGXJD5_2;
	wire w_dff_A_GBmzx6wz4_2;
	wire w_dff_B_z6k5rTOH2_1;
	wire w_dff_B_cvGlQ0044_1;
	wire w_dff_B_bsMZhnDY2_1;
	wire w_dff_B_ttpy0CZW9_1;
	wire w_dff_B_3VKKs2DS2_1;
	wire w_dff_A_fZQ7cme07_1;
	wire w_dff_A_Aco4Rfxw7_1;
	wire w_dff_A_EUgEOsnn9_1;
	wire w_dff_A_khJRHsrT5_1;
	wire w_dff_A_OY7Q8sWP2_1;
	wire w_dff_A_9aUQXAKb9_1;
	wire w_dff_A_srQ6aHx94_1;
	wire w_dff_A_mi9eGh4F5_0;
	wire w_dff_A_rLAMROX73_0;
	wire w_dff_A_enGQamJO4_0;
	wire w_dff_A_62LuOKr94_0;
	wire w_dff_A_ji7Ssb0i9_0;
	wire w_dff_A_FHuImOqd3_0;
	wire w_dff_A_8VYSaQLh2_0;
	wire w_dff_A_F7FvTbIU6_0;
	wire w_dff_A_xXu241s53_0;
	wire w_dff_A_GPjp26wa3_0;
	wire w_dff_A_mqHihzL63_0;
	wire w_dff_A_Dp3jRNxF2_0;
	wire w_dff_A_1T9U05Yz1_0;
	wire w_dff_A_dpYbe0Vd4_0;
	wire w_dff_A_JOATgsfg6_0;
	wire w_dff_A_37apWN0E4_0;
	wire w_dff_A_LEtQZjGE5_0;
	wire w_dff_B_cPd2n3vn8_2;
	wire w_dff_B_pJnT534a4_2;
	wire w_dff_A_mirKFcdb1_1;
	wire w_dff_A_8b2e4GZU0_1;
	wire w_dff_A_1dhyPwgU6_1;
	wire w_dff_A_xHW8LyAM9_1;
	wire w_dff_A_Wjj189Lq3_1;
	wire w_dff_A_qGF3hIIh8_1;
	wire w_dff_A_oNpKmeNu2_1;
	wire w_dff_A_L83vThpW0_1;
	wire w_dff_A_PhQ3LTox0_1;
	wire w_dff_A_enWkxjoB9_1;
	wire w_dff_A_EMhCsHJR1_2;
	wire w_dff_B_EXzRqPhv9_0;
	wire w_dff_B_vbotFnb24_1;
	wire w_dff_A_Rr5OZwbN8_0;
	wire w_dff_A_4x3qatY19_2;
	wire w_dff_A_8mxpvWCz0_2;
	wire w_dff_A_Yv6kDql04_2;
	wire w_dff_A_ib9Rh1lq1_2;
	wire w_dff_B_qtKr0fpF5_1;
	wire w_dff_B_O0nRUcvV3_1;
	wire w_dff_A_fpZxkH2L2_0;
	wire w_dff_A_BmdpZ4Lh4_0;
	wire w_dff_A_4cNbMmsO6_0;
	wire w_dff_A_r3NdDLcl6_2;
	wire w_dff_A_mLhvBfUC2_2;
	wire w_dff_A_weVSCX4f8_2;
	wire w_dff_A_g4AstPkX1_2;
	wire w_dff_A_cRaF1Mbl7_2;
	wire w_dff_A_G6qPK8wB9_2;
	wire w_dff_A_xgc5JR2D4_2;
	wire w_dff_B_K5Phutoi0_2;
	wire w_dff_A_7Weigvoq1_1;
	wire w_dff_B_G1yOpguQ2_0;
	wire w_dff_B_y63hCaOL7_1;
	wire w_dff_B_Yd1FmHXW5_0;
	wire w_dff_B_8f4RVvMu5_1;
	wire w_dff_A_VySiNYam7_1;
	wire w_dff_A_BLVgBP3s8_0;
	wire w_dff_A_KaP3mLZ20_0;
	wire w_dff_B_8quRQZr08_2;
	wire w_dff_B_PGJ73wt72_2;
	wire w_dff_B_i8QFpFER7_2;
	wire w_dff_A_hyklK2l55_0;
	wire w_dff_A_B2v12AOc4_0;
	wire w_dff_A_HKTgWa7w6_0;
	wire w_dff_A_Awaqc4aS2_0;
	wire w_dff_A_2QmQ8UmM1_1;
	wire w_dff_A_0VGBal8i6_1;
	wire w_dff_A_WHOrqpLf1_1;
	wire w_dff_A_mp2OLete7_1;
	wire w_dff_A_RIzCUENo3_1;
	wire w_dff_A_Xw0QZFdE1_1;
	wire w_dff_A_MXSlLSCG9_2;
	wire w_dff_A_UexTmkzh5_2;
	wire w_dff_A_2JeTvPl28_2;
	wire w_dff_A_obhZ1qgF7_2;
	wire w_dff_A_9OxIGf3C9_2;
	wire w_dff_A_NxH4tdPn0_2;
	wire w_dff_B_kghlOlOs9_0;
	wire w_dff_B_h6UqhT4u7_0;
	wire w_dff_B_ZRUgqySz6_0;
	wire w_dff_B_cgW0hOZr8_0;
	wire w_dff_B_wcYJ1TzN1_0;
	wire w_dff_B_BrCnk7Kw2_0;
	wire w_dff_B_SmgpBJxx1_0;
	wire w_dff_B_jFPfXCOu8_0;
	wire w_dff_B_kmufscFm5_0;
	wire w_dff_B_2j0nYXVw6_0;
	wire w_dff_B_6bkGyK2w7_0;
	wire w_dff_B_NmUcLTXn0_1;
	wire w_dff_B_8COAyz5T1_1;
	wire w_dff_B_4grUwu5F0_1;
	wire w_dff_A_NxE5199g4_0;
	wire w_dff_A_c1571MWv0_0;
	wire w_dff_B_1UAZNobP5_2;
	wire w_dff_B_VNHm9cY24_2;
	wire w_dff_B_918j1l7K2_2;
	wire w_dff_B_VjbN95og9_2;
	wire w_dff_B_fivtRROq9_2;
	wire w_dff_B_ux2iu24m6_2;
	wire w_dff_B_6ape9e1y0_2;
	wire w_dff_B_7HdnSMWM1_2;
	wire w_dff_B_TWfjzTAo4_2;
	wire w_dff_B_3apDr30h5_2;
	wire w_dff_B_Ujo9Syr77_2;
	wire w_dff_B_fCBI0eF75_2;
	wire w_dff_A_Kyha9QU23_0;
	wire w_dff_A_LpLLVyIt7_0;
	wire w_dff_A_b8Zi22nb3_0;
	wire w_dff_A_G8jV60gn7_0;
	wire w_dff_A_gv9hIwzM5_0;
	wire w_dff_A_efNm6fAq4_0;
	wire w_dff_A_7lweI8Tw5_0;
	wire w_dff_A_MwC5JsDB6_0;
	wire w_dff_A_WqcEn3r81_0;
	wire w_dff_A_XuDmv30e4_0;
	wire w_dff_A_AccpODWJ0_0;
	wire w_dff_A_MVkNx5Pp9_0;
	wire w_dff_A_2UiPeyF29_0;
	wire w_dff_A_nSdn0rlr3_0;
	wire w_dff_A_USsYQNdK9_0;
	wire w_dff_A_4ouY8qtj9_1;
	wire w_dff_A_F4FUDs3M5_1;
	wire w_dff_A_TLumZ1LD0_1;
	wire w_dff_A_nq8MFM1V3_1;
	wire w_dff_A_OpuR5ybL5_1;
	wire w_dff_A_Kyfo73fF2_1;
	wire w_dff_A_OAl2Lzxh7_1;
	wire w_dff_A_D5i4tLOH4_1;
	wire w_dff_A_1Perz2kI6_1;
	wire w_dff_A_qGhmJ1uq6_1;
	wire w_dff_A_uod133Nn2_1;
	wire w_dff_A_fKRahply6_1;
	wire w_dff_B_KmuGB4Wa4_1;
	wire w_dff_B_2bHVAlJb1_1;
	wire w_dff_B_iWpnZ9fZ2_0;
	wire w_dff_B_KmjT6LZ54_0;
	wire w_dff_B_QXQtFWVM3_0;
	wire w_dff_B_KEuu4M2p9_0;
	wire w_dff_A_jmLmb4bc5_0;
	wire w_dff_A_SdXrTuRN7_0;
	wire w_dff_A_KftsghUC4_0;
	wire w_dff_A_zQUxjSjB4_0;
	wire w_dff_A_1iPsS97d8_0;
	wire w_dff_A_S4J3oz055_0;
	wire w_dff_A_tLTauKTU4_2;
	wire w_dff_A_8QoqLDaH3_2;
	wire w_dff_A_j64Xv3qz2_2;
	wire w_dff_A_i3G21l3P2_2;
	wire w_dff_A_QqAqicj04_2;
	wire w_dff_A_6POUhTop1_1;
	wire w_dff_A_uIGeh2Lg0_1;
	wire w_dff_A_Nbzwjh4j8_1;
	wire w_dff_A_oC8bNNVc9_1;
	wire w_dff_B_yCM6XrYW8_0;
	wire w_dff_B_LGHcPilM5_1;
	wire w_dff_B_eWV88eXH9_1;
	wire w_dff_B_FjYJOSeL0_1;
	wire w_dff_B_xDHxEj471_1;
	wire w_dff_B_9qF6hteK6_1;
	wire w_dff_B_RS5LCjhX5_1;
	wire w_dff_A_Z638JVzt5_1;
	wire w_dff_A_CvzPEdAw0_1;
	wire w_dff_A_5jgei4zv9_1;
	wire w_dff_A_thC6SE5m2_1;
	wire w_dff_A_v8XxsTxc9_1;
	wire w_dff_A_hur0nhdE9_1;
	wire w_dff_A_2tTVCuS14_1;
	wire w_dff_A_h5ww4nX32_0;
	wire w_dff_A_IP7kNLv53_0;
	wire w_dff_A_3drH5Idj8_1;
	wire w_dff_A_oXcb4rub9_1;
	wire w_dff_A_NVFluDeo3_2;
	wire w_dff_A_VL4FUWSr8_2;
	wire w_dff_A_vLl8KNLZ3_2;
	wire w_dff_A_apldzcTr2_2;
	wire w_dff_B_36jfe22f8_0;
	wire w_dff_B_rh2BxCzh4_1;
	wire w_dff_A_PZqyPr7U8_1;
	wire w_dff_A_ZC2bstJW3_1;
	wire w_dff_A_oMKzX95G8_0;
	wire w_dff_A_DCcBNEoT4_0;
	wire w_dff_B_UZ0RO1iU3_0;
	wire w_dff_B_xzfxRi8R7_0;
	wire w_dff_B_NbMeyCxI1_0;
	wire w_dff_A_E8RvXwhG7_0;
	wire w_dff_A_LlCKywvu0_1;
	wire w_dff_A_6f9bX2tD6_1;
	wire w_dff_B_I6rSOM260_1;
	wire w_dff_A_s88eH5Y14_0;
	wire w_dff_A_Qe9sEAx29_1;
	wire w_dff_A_NHIWFKCJ9_1;
	wire w_dff_B_hQ7pqEYK6_1;
	wire w_dff_A_2L149ccd6_0;
	wire w_dff_A_Hv98Ul3Y0_0;
	wire w_dff_A_s2LmmwUv5_1;
	wire w_dff_B_dcyVP1xp6_1;
	wire w_dff_A_zuN3zQmS5_0;
	wire w_dff_A_qDxhoPsK9_0;
	wire w_dff_A_hl6HUjuu1_0;
	wire w_dff_A_b2al5vls9_1;
	wire w_dff_B_WxmNg9VF5_1;
	wire w_dff_A_v4ndQapO6_0;
	wire w_dff_A_vm5gbBGa0_0;
	wire w_dff_A_K02QV1Jy0_0;
	wire w_dff_B_889MNSiZ3_0;
	wire w_dff_B_Q1twm8zD2_1;
	wire w_dff_B_EtmbtrLr8_1;
	wire w_dff_A_oLekoJB74_0;
	wire w_dff_A_v255Axo79_1;
	wire w_dff_A_begpvNal4_1;
	wire w_dff_B_fLnXQ0Lb0_3;
	wire w_dff_A_8eZYEhHf5_0;
	wire w_dff_A_j9NSDTOJ0_0;
	wire w_dff_A_9ln3n0g28_0;
	wire w_dff_A_ofFN2KXF6_0;
	wire w_dff_A_IvhJg8688_1;
	wire w_dff_A_Fz4uHTIG0_1;
	wire w_dff_A_L5HpIfiT5_1;
	wire w_dff_A_j1EMTddv1_1;
	wire w_dff_A_1KzzcdFs5_1;
	wire w_dff_A_y63zbw8x4_1;
	wire w_dff_A_cKOUHrFF9_2;
	wire w_dff_A_rmmWmvdv0_2;
	wire w_dff_A_YXtTpnJ03_2;
	wire w_dff_A_SfgBxLJ12_2;
	wire w_dff_A_ObGN1cyK6_2;
	wire w_dff_B_wX4VpuQn3_1;
	wire w_dff_A_5zvoiHyn4_0;
	wire w_dff_A_qvgEtbMD4_1;
	wire w_dff_A_g2ibEBXg4_1;
	wire w_dff_B_HKAzCg7R7_3;
	wire w_dff_A_ZPEVKmD71_0;
	wire w_dff_A_FkFWjuf19_0;
	wire w_dff_A_MAAjVj5D3_0;
	wire w_dff_A_A5Y9CIJd1_0;
	wire w_dff_A_6IczPJFg8_1;
	wire w_dff_A_kk6Xg4d20_1;
	wire w_dff_A_UmtnvGTW6_1;
	wire w_dff_B_d0nm04rx4_1;
	wire w_dff_A_omqAYVWi0_0;
	wire w_dff_A_dOKrPts53_1;
	wire w_dff_A_Zllgn7rC3_1;
	wire w_dff_A_M1BjK6yz4_2;
	wire w_dff_A_X80VAKJu5_2;
	wire w_dff_A_QVEhdUTm7_2;
	wire w_dff_A_C4MnImA90_2;
	wire w_dff_A_GfG3u0CN9_0;
	wire w_dff_B_Evnm23O15_1;
	wire w_dff_B_2GqOtywX5_1;
	wire w_dff_A_jKyEDYcW2_0;
	wire w_dff_A_EnrzktwJ9_2;
	wire w_dff_A_2XBEw37y9_2;
	wire w_dff_A_Kof4lzNX5_2;
	wire w_dff_B_OzpKQcnl0_3;
	wire w_dff_A_p5OtCipC7_0;
	wire w_dff_A_LtzjnPaH2_0;
	wire w_dff_A_byQV1EwN1_0;
	wire w_dff_A_67X00Ndi9_1;
	wire w_dff_A_uxQAF81y4_1;
	wire w_dff_A_sS3oEy2s3_1;
	wire w_dff_A_e1WClZRI7_2;
	wire w_dff_A_pbJw1qfz5_2;
	wire w_dff_A_U6Ikx0Vg4_2;
	wire w_dff_A_M0zNXlLG7_2;
	wire w_dff_A_gT9buK4T4_2;
	wire w_dff_B_MT3m1v0b3_1;
	wire w_dff_B_Iy94drE61_1;
	wire w_dff_B_VYw4pF030_1;
	wire w_dff_A_vMNUiQfu8_0;
	wire w_dff_A_KR7BGXZC0_0;
	wire w_dff_A_ofgL8hNt0_0;
	wire w_dff_A_PoDJRc4n1_1;
	wire w_dff_A_1GH9ejTP0_1;
	wire w_dff_A_ClsEoZwW8_1;
	wire w_dff_A_d9umcNL71_1;
	wire w_dff_A_m1ayBrvp4_1;
	wire w_dff_A_ZxaHmWHq9_1;
	wire w_dff_A_TKLUWJgi2_2;
	wire w_dff_A_77SFOBKl7_2;
	wire w_dff_A_Mmgn51Xh7_2;
	wire w_dff_A_5HCCnfVr4_0;
	wire w_dff_B_UhzF9ryi3_1;
	wire w_dff_B_wNMw5I5N0_1;
	wire w_dff_B_tRZZYgo67_1;
	wire w_dff_B_SeD0dRPb3_1;
	wire w_dff_A_IAv7bVlJ3_0;
	wire w_dff_A_k3UyB8Po6_1;
	wire w_dff_A_KZ8wSDaz2_1;
	wire w_dff_A_vrW7pce47_1;
	wire w_dff_B_d2dBaqaS5_3;
	wire w_dff_A_ixjX31sh3_0;
	wire w_dff_A_GtMqQLe60_0;
	wire w_dff_A_YbWXFDCo7_0;
	wire w_dff_A_ZOupd35Q9_0;
	wire w_dff_A_4nBuZFG15_1;
	wire w_dff_A_fZxMoYKW5_1;
	wire w_dff_A_lrnp6gFq2_1;
	wire w_dff_A_Nnii9NIS3_1;
	wire w_dff_A_a1yMwuBY3_1;
	wire w_dff_A_qaPcEWrT7_1;
	wire w_dff_A_N81RKIix8_2;
	wire w_dff_A_sFDtG4JR7_2;
	wire w_dff_A_Noi6SRXT0_2;
	wire w_dff_A_8lsHxblE7_2;
	wire w_dff_A_zJ4OzjGQ4_2;
	wire w_dff_B_m6dmyI8h8_1;
	wire w_dff_B_GsQmPUvU2_1;
	wire w_dff_A_jWHGvtCa9_0;
	wire w_dff_A_LwEQZpPG1_1;
	wire w_dff_A_SsfZd5P01_1;
	wire w_dff_B_9BYI8BGR2_3;
	wire w_dff_A_jk3Igepg2_0;
	wire w_dff_A_A3snWA4u5_0;
	wire w_dff_A_8CYTgtUW9_0;
	wire w_dff_A_SWo3DVyA2_0;
	wire w_dff_A_VxC4n2dU9_1;
	wire w_dff_A_QxBoCB4y1_1;
	wire w_dff_A_VgDuH2sX9_1;
	wire w_dff_A_McdFHEj28_1;
	wire w_dff_A_SSYCyo4y7_1;
	wire w_dff_A_RU41QhYS4_1;
	wire w_dff_A_BYPkcyG07_2;
	wire w_dff_A_SpExcGnA3_2;
	wire w_dff_A_xlgPmUFB1_2;
	wire w_dff_A_A8WUKmeI4_2;
	wire w_dff_A_CID2Snx76_2;
	wire w_dff_B_vQWbygcP6_1;
	wire w_dff_A_TJDdjxDN3_1;
	wire w_dff_A_Fq7oCxoN3_1;
	wire w_dff_A_pMW24VFp3_2;
	wire w_dff_B_5B0514A33_3;
	wire w_dff_A_0HziCBUR3_0;
	wire w_dff_A_xtl1iMlQ9_0;
	wire w_dff_A_I4r5TiI65_0;
	wire w_dff_A_PRE9t4K11_0;
	wire w_dff_A_CDgMUzjN4_1;
	wire w_dff_A_mGBU1vtR5_1;
	wire w_dff_A_BcsnzGcI1_1;
	wire w_dff_B_ii3wpd5b0_1;
	wire w_dff_A_J1GBjRnw5_0;
	wire w_dff_A_iW6HyRsz8_0;
	wire w_dff_A_3HPeGmjr0_2;
	wire w_dff_A_Xe8Fmw9H8_1;
	wire w_dff_A_poS3m5Qm4_1;
	wire w_dff_A_AsvBBfPu7_2;
	wire w_dff_A_WrXyI5iu0_2;
	wire w_dff_A_v6NM0Qup3_2;
	wire w_dff_A_OVVhrC421_2;
	wire w_dff_A_yKhhrmpy2_1;
	wire w_dff_A_c5SsxF4r5_2;
	wire w_dff_B_9eh08wkv9_1;
	wire w_dff_B_o8C3BcRH5_1;
	wire w_dff_A_YLF0ccXX5_0;
	wire w_dff_A_NuzqmZ4V1_1;
	wire w_dff_A_zxckjhqV0_1;
	wire w_dff_A_vRi5HaW28_2;
	wire w_dff_A_oEkkQGhu1_2;
	wire w_dff_B_b9meJiND4_3;
	wire w_dff_A_3BW8hfJP5_0;
	wire w_dff_A_vZMHX8wm5_0;
	wire w_dff_A_9TpVP1lK2_0;
	wire w_dff_A_oxlsLqtp8_0;
	wire w_dff_A_kYWSXtUk2_1;
	wire w_dff_A_MfbTLasS1_1;
	wire w_dff_A_pi6uTrMi7_1;
	wire w_dff_A_8d7Ye7kU8_1;
	wire w_dff_A_D5okqryN3_1;
	wire w_dff_A_MbOpF8PG8_1;
	wire w_dff_A_vRwjoFX78_2;
	wire w_dff_A_2PR6l5d35_2;
	wire w_dff_A_XbVAolyy7_2;
	wire w_dff_A_5g6MpCxj4_2;
	wire w_dff_A_YoDwKxKM6_2;
	wire w_dff_A_ObhXBezk2_0;
	wire w_dff_A_vXPYLiIZ1_1;
	wire w_dff_A_zeUXuxX64_2;
	wire w_dff_B_J9zxAP4D0_1;
	wire w_dff_B_4fm55Zox3_1;
	wire w_dff_A_CCG8Zxt41_0;
	wire w_dff_A_h7Jd0gJN0_1;
	wire w_dff_A_DQGrjRHK8_2;
	wire w_dff_A_AKrFKqE09_1;
	wire w_dff_A_fWW2UeFb7_1;
	wire w_dff_A_JRx1cu4J3_2;
	wire w_dff_A_r91G5d5d1_2;
	wire w_dff_B_2DsNOHuP7_3;
	wire w_dff_A_ijT9kB0A1_0;
	wire w_dff_A_Wwvhte7V5_0;
	wire w_dff_A_El7HS5tF9_0;
	wire w_dff_A_juiEJIiC2_0;
	wire w_dff_A_z5CTrU3b2_0;
	wire w_dff_A_MFdt46Gh2_0;
	wire w_dff_A_lge6Nse23_0;
	wire w_dff_A_kMCUL8xc2_2;
	wire w_dff_A_QctWO7aU5_2;
	wire w_dff_A_HuQwAL7r3_2;
	wire w_dff_A_AK5xYz0k8_1;
	wire w_dff_A_4imqgMe79_2;
	wire w_dff_A_OfhDr8Jr0_2;
	wire w_dff_A_XL4AbLks6_1;
	wire w_dff_A_2ZuXrpe36_1;
	wire w_dff_A_t8w2e87r8_1;
	wire w_dff_A_oPNC0mPF0_1;
	wire w_dff_A_5yGfR4rj6_1;
	wire w_dff_A_MJ6Hvoij0_1;
	wire w_dff_A_RCJMwuVo0_1;
	wire w_dff_A_VBAUcQae1_1;
	wire w_dff_A_q49p95m61_1;
	wire w_dff_A_EXDpjo6W6_1;
	wire w_dff_A_QOcUvxSe8_1;
	wire w_dff_A_T1dFYe3G1_1;
	wire w_dff_A_rmSyudrV7_1;
	wire w_dff_A_sgr2C9MX6_1;
	wire w_dff_A_HEfhdYZv6_1;
	wire w_dff_A_vd0hohDx2_1;
	wire w_dff_A_CQbw284R5_1;
	wire w_dff_A_qc0WrT8J1_2;
	wire w_dff_A_oCgrTsBV9_2;
	wire w_dff_A_HIR4MtVn9_2;
	wire w_dff_A_KO4VY6Sp8_2;
	wire w_dff_A_40Z9CLjG2_2;
	wire w_dff_A_8QOhCgk58_2;
	wire w_dff_A_YfRbn58s9_2;
	wire w_dff_A_oRDUx95A7_2;
	wire w_dff_A_xo8H0iUw2_1;
	wire w_dff_A_pU6HVoYk6_1;
	wire w_dff_A_h14ZsECt1_1;
	wire w_dff_A_WSPSDGqZ9_1;
	wire w_dff_A_9q4aPqhS1_2;
	wire w_dff_A_yHz3fP6c9_2;
	wire w_dff_A_dsMB0Ji38_2;
	wire w_dff_A_MsncRhbx1_2;
	wire w_dff_A_2uW4Q9kK5_1;
	wire w_dff_A_lYHRuC0r7_1;
	wire w_dff_A_Aur4jt7Q5_2;
	wire w_dff_A_71ICoD9D2_2;
	wire w_dff_A_dbchnsP29_2;
	wire w_dff_A_VjbP3K595_0;
	wire w_dff_A_86b8CQdR3_0;
	wire w_dff_A_IEo8tGwN3_0;
	wire w_dff_A_mljz6IqM0_0;
	wire w_dff_A_piDFrEPc8_0;
	wire w_dff_A_EitXLudL1_0;
	wire w_dff_A_QnZl4vUa2_0;
	wire w_dff_A_9Xb9cIaV5_0;
	wire w_dff_A_0E3KASNc4_0;
	wire w_dff_A_ZZv3dkAw8_0;
	wire w_dff_A_tUwb5tTI9_0;
	wire w_dff_A_sQwWNgac7_0;
	wire w_dff_A_WS9eeEtU1_0;
	wire w_dff_A_9OEWljUK9_1;
	wire w_dff_A_Wo73ayXj5_1;
	wire w_dff_A_9HeyBpws5_1;
	wire w_dff_A_8LSCkkyj2_1;
	wire w_dff_A_PIJVGkZz1_1;
	wire w_dff_A_Ss8MEqmn8_1;
	wire w_dff_A_H1SsEM2h4_1;
	wire w_dff_A_9MtcZvZE4_1;
	wire w_dff_A_KKuVZUuQ7_1;
	wire w_dff_A_yQfGyEy12_1;
	wire w_dff_A_cf86T9NH3_1;
	wire w_dff_A_VjAtKayS5_1;
	wire w_dff_A_ajbuNz1y3_1;
	wire w_dff_A_Szs7ReQ35_1;
	wire w_dff_A_UGiFwJl39_1;
	wire w_dff_A_t3Q4ZoCk4_1;
	wire w_dff_A_5QgE2dt85_1;
	wire w_dff_A_2I9ItvmN3_1;
	wire w_dff_A_XdZlMQAp8_1;
	wire w_dff_A_ZsiNco8d4_1;
	wire w_dff_A_sV38P4L49_2;
	wire w_dff_A_o1bSZhtG4_2;
	wire w_dff_A_RxDwcOHl8_2;
	wire w_dff_A_4GsiOF2g8_2;
	wire w_dff_A_id7i98L30_2;
	wire w_dff_A_z11Eld5C5_2;
	wire w_dff_A_b6se461D7_2;
	wire w_dff_A_pFqduqXp0_2;
	wire w_dff_A_r7IPFdiu7_2;
	wire w_dff_A_ugPDC4sW7_2;
	wire w_dff_A_JW7ucBXq1_2;
	wire w_dff_A_orSiVrM64_2;
	wire w_dff_A_psOsMHOR2_2;
	wire w_dff_A_tQ5rBqIt1_2;
	wire w_dff_A_TQCfDaYJ3_2;
	wire w_dff_A_WV4ki3Zp1_2;
	wire w_dff_A_hNALHbFE6_2;
	wire w_dff_A_YnuYCGgS8_2;
	wire w_dff_A_tWgS3oAK1_2;
	wire w_dff_A_WsPtK1r61_2;
	wire w_dff_A_Tvm6nn3e3_2;
	wire w_dff_A_DnTYD3nX1_2;
	wire w_dff_A_fCJhd0fm9_2;
	wire w_dff_A_UJ2Znemh6_2;
	wire w_dff_A_Ws7c9QGw6_2;
	wire w_dff_A_r7lXwKxe0_2;
	wire w_dff_A_8AcuioY74_2;
	wire w_dff_A_4gOJRDdD0_2;
	wire w_dff_A_QPoL2Yr86_1;
	wire w_dff_A_WSqycTFI7_0;
	wire w_dff_A_uUSEqkrO9_0;
	wire w_dff_A_ON0sg6aB4_0;
	wire w_dff_A_4uUDOd8n9_0;
	wire w_dff_A_ok1mW5CE9_0;
	wire w_dff_A_Qx3w1VQI2_0;
	wire w_dff_A_8f1KVLOG8_0;
	wire w_dff_A_SMf7Agkr3_0;
	wire w_dff_A_n88UjXSt9_0;
	wire w_dff_A_4EMrDtKz7_0;
	wire w_dff_A_2ZojMmEh2_0;
	wire w_dff_A_OYIlsWXH8_0;
	wire w_dff_A_qFgT65Bj9_0;
	wire w_dff_A_XCvCTKxb7_0;
	wire w_dff_A_SKWies1N4_0;
	wire w_dff_A_u3Idcy3m6_2;
	wire w_dff_A_LA10yz5M3_2;
	wire w_dff_A_TlxeCcEY4_2;
	wire w_dff_A_QQO0Bdfn3_2;
	wire w_dff_A_bSPJPTBF8_2;
	wire w_dff_A_EGyJJntq3_2;
	wire w_dff_A_D5C9xmcl9_2;
	wire w_dff_A_OQJO4pMg6_2;
	wire w_dff_A_zcNQ3ys02_2;
	wire w_dff_A_mZ86McBp3_2;
	wire w_dff_A_kSfNaV7k4_1;
	wire w_dff_A_XCW97tO20_1;
	wire w_dff_A_dsynUTGi1_1;
	wire w_dff_A_oLJktYkX3_1;
	wire w_dff_A_OhuHp5ts4_1;
	wire w_dff_A_dnfSHvyF5_1;
	wire w_dff_A_Bh0PukLk2_1;
	wire w_dff_A_Q7GQe5kG7_1;
	wire w_dff_A_VJp9CNGQ7_1;
	wire w_dff_A_Npfoxvkr2_1;
	wire w_dff_A_RRf0z1JV7_1;
	wire w_dff_A_0LDNOHWG8_1;
	wire w_dff_A_pjQgGHN08_1;
	wire w_dff_A_XJr2CE7J8_1;
	wire w_dff_A_wayGqTb63_1;
	wire w_dff_A_DYHgFZ441_1;
	wire w_dff_A_52KHvoTS2_1;
	wire w_dff_A_WR26FZwb7_1;
	wire w_dff_A_xftwfBFJ9_1;
	wire w_dff_A_QDnQbt1F5_1;
	wire w_dff_A_pQ3HAkyF6_1;
	wire w_dff_A_SIxGBBAz0_2;
	wire w_dff_A_oR8Ojy7Q8_2;
	wire w_dff_A_Fs10dkLd6_2;
	wire w_dff_A_pO8CWy865_2;
	wire w_dff_A_mP8DDIcz7_2;
	wire w_dff_A_rdAFcOJ67_2;
	wire w_dff_A_sTvDPdlT3_2;
	wire w_dff_A_bHA0pX3V9_2;
	wire w_dff_A_ZxqKzhHM7_2;
	wire w_dff_A_5LGF4Llh5_2;
	wire w_dff_A_YuYIoP734_2;
	wire w_dff_A_RMrA0vc58_2;
	wire w_dff_A_1DDlXiSl7_2;
	wire w_dff_A_A0wXchy67_2;
	wire w_dff_A_axxn571j7_2;
	wire w_dff_A_fizGF83e2_2;
	wire w_dff_A_7exSQ6oc8_2;
	wire w_dff_A_Klt8O5nc0_2;
	wire w_dff_A_AwGANxKm8_2;
	wire w_dff_A_SwhyDRds8_2;
	wire w_dff_A_joNpa7pj5_1;
	wire w_dff_A_IwgFjkYh3_1;
	wire w_dff_A_KLZFKEtw2_1;
	wire w_dff_A_7FxgQzyS8_1;
	wire w_dff_A_mKKPOxLH8_1;
	wire w_dff_A_eFGPnXsz7_1;
	wire w_dff_A_EHMk3NIn7_1;
	wire w_dff_A_NklZwVqI4_1;
	wire w_dff_A_Sv95TVcw6_1;
	wire w_dff_A_PKwUAUwU8_1;
	wire w_dff_A_oUP31tfa2_1;
	wire w_dff_A_MVYqPbwh5_1;
	wire w_dff_A_CRBbVg4z5_1;
	wire w_dff_A_8BtsdIM15_1;
	wire w_dff_A_vH45RwE30_1;
	wire w_dff_A_CBJv59lI3_1;
	wire w_dff_A_fDL2Gcz20_1;
	wire w_dff_A_b1Z1GqIh7_1;
	wire w_dff_A_gZloFhOf3_2;
	wire w_dff_A_Lu9EV3RW3_2;
	wire w_dff_A_jNxfeHUK6_2;
	wire w_dff_A_CDcBIiOV7_2;
	wire w_dff_A_HW3Sb6ig8_2;
	wire w_dff_A_C9YfbesS1_2;
	wire w_dff_A_pyMCgMEp8_2;
	wire w_dff_A_da5ylVH45_2;
	wire w_dff_A_9BWh89Fn8_2;
	wire w_dff_A_PoY3Yy488_2;
	wire w_dff_A_wtsjZLC43_2;
	wire w_dff_A_lvhsygkr0_1;
	wire w_dff_A_nGbJspLH0_1;
	wire w_dff_A_zMCP0Xa69_1;
	wire w_dff_A_Mtb30mf10_1;
	wire w_dff_A_7z7cGEbk7_1;
	wire w_dff_A_LLipclX71_1;
	wire w_dff_A_sXUPwNmt9_1;
	wire w_dff_A_GUx2y2KX8_1;
	wire w_dff_A_KCA2LkGM5_1;
	wire w_dff_B_JFNhjRj26_2;
	wire w_dff_B_SHjTvCFN8_2;
	wire w_dff_A_NrHeVJaU2_1;
	wire w_dff_A_OYuBxBoI3_1;
	wire w_dff_A_83w313hf4_1;
	wire w_dff_A_uq3IpMya7_1;
	wire w_dff_A_PndnQEq71_1;
	wire w_dff_A_tt66UUE16_1;
	wire w_dff_A_MkNfVwnp9_1;
	wire w_dff_A_6CU7N1Vx3_1;
	wire w_dff_A_HL2V6y215_1;
	wire w_dff_A_MgmqeuPb5_1;
	wire w_dff_A_R894gWeW2_1;
	wire w_dff_A_xVXb5A5Y1_1;
	wire w_dff_A_bvIW5vGo3_1;
	wire w_dff_A_aHrjlshB3_1;
	wire w_dff_A_n8pSpgXP7_1;
	wire w_dff_A_WI9PiHta0_1;
	wire w_dff_A_K8lD1TQj4_1;
	wire w_dff_A_LbbRRbec4_1;
	wire w_dff_A_veYxSZ2n8_1;
	wire w_dff_A_IR6oyroZ0_1;
	wire w_dff_A_o6R8sHul4_1;
	wire w_dff_A_rm69yGQw1_1;
	wire w_dff_A_PuJrd79y3_1;
	wire w_dff_A_dgGMwTgw5_2;
	wire w_dff_A_jez6q3ck6_0;
	wire w_dff_A_Y5Htbw501_0;
	wire w_dff_A_y1XNu93O5_0;
	wire w_dff_A_nuFK7bXb4_0;
	wire w_dff_A_EupK70Ep0_0;
	wire w_dff_A_lFRbiMll2_0;
	wire w_dff_A_rffl1DUk7_0;
	wire w_dff_A_jg5l5pMu3_0;
	wire w_dff_A_uU8WhNG28_0;
	wire w_dff_A_hKfi0Hnm4_0;
	wire w_dff_A_lmAqRxtF5_0;
	wire w_dff_A_nGpldJDP8_0;
	wire w_dff_A_OSok7hQx6_0;
	wire w_dff_A_eNq6EuQo6_0;
	wire w_dff_A_ZJRvuEij9_1;
	wire w_dff_A_DPFh9Ds93_1;
	wire w_dff_A_cnEbxqi33_1;
	wire w_dff_A_wKY5CZ829_1;
	wire w_dff_A_tSDqsGMI2_1;
	wire w_dff_A_fgD7Vqk01_1;
	wire w_dff_A_eqb7eVTU8_1;
	wire w_dff_A_6WBwahvX6_1;
	wire w_dff_A_nDzZ8UwB1_1;
	wire w_dff_A_51fD4GFb3_1;
	wire w_dff_A_MORzu4mx0_1;
	wire w_dff_A_9MzmqfIV6_1;
	wire w_dff_A_6UCJrQ7E3_1;
	wire w_dff_A_c1qCztz99_1;
	wire w_dff_A_Al4YqERy7_1;
	wire w_dff_A_XLZ3R2fU3_1;
	wire w_dff_A_ZtOT0hLB6_2;
	wire w_dff_A_pel3Qd872_2;
	wire w_dff_A_bqdsjcwZ5_2;
	wire w_dff_A_RF67uqnd0_2;
	wire w_dff_A_sLk00SdQ3_2;
	wire w_dff_A_oTAhzqlh9_2;
	wire w_dff_A_5DeqOacz4_2;
	wire w_dff_A_ApLMwgYC1_2;
	wire w_dff_A_r9sl2ikc0_2;
	wire w_dff_A_tnokxD7K6_2;
	wire w_dff_A_PKYjso3T5_2;
	wire w_dff_A_aETqB8B26_2;
	wire w_dff_A_XFia1uVj0_2;
	wire w_dff_A_e2Ael8mC2_2;
	wire w_dff_A_WtGp5k6j4_2;
	wire w_dff_A_NibZ94Xm9_2;
	wire w_dff_A_iq4YHuwO1_2;
	wire w_dff_A_GcuuUpUv0_2;
	wire w_dff_A_lnW7Jwxq5_2;
	wire w_dff_A_bf8uZ9ug9_2;
	wire w_dff_A_nfyhVbYY1_2;
	wire w_dff_A_DEUdClEX8_2;
	wire w_dff_A_uOHIpPs64_1;
	wire w_dff_A_Pe0dDGyj5_1;
	wire w_dff_A_RAB56aaU4_1;
	wire w_dff_A_HUKCjav54_1;
	wire w_dff_A_Rb6g0GMP0_1;
	wire w_dff_A_UOAqTRwi0_1;
	wire w_dff_A_RqlN2u1v4_1;
	wire w_dff_A_05hehML31_1;
	wire w_dff_A_IjBL1HG98_1;
	wire w_dff_A_lboOwYLZ3_1;
	wire w_dff_A_qlbNgzLd4_1;
	wire w_dff_A_ivzypPC02_1;
	wire w_dff_A_glX40HsQ0_1;
	wire w_dff_A_MBUqYFrl2_1;
	wire w_dff_A_wbaxU3AM2_1;
	wire w_dff_A_xAhcRo9w8_1;
	wire w_dff_A_RX3Z8UeR4_1;
	wire w_dff_A_KJeWS4oe5_1;
	wire w_dff_A_6aehFRuv9_1;
	wire w_dff_A_dMd4Dplq1_2;
	wire w_dff_A_4GLrp35o8_2;
	wire w_dff_A_WuFYFDj19_2;
	wire w_dff_A_5zI5gduW9_2;
	wire w_dff_A_JcBH96rA1_2;
	wire w_dff_A_RwUuL03E9_2;
	wire w_dff_A_qSKoB0l20_2;
	wire w_dff_A_JzZxz98o0_2;
	wire w_dff_A_KFrZBu1F1_2;
	wire w_dff_A_0RcGyH1M4_2;
	wire w_dff_A_klkUp8ao9_2;
	wire w_dff_A_dT8Ia2OZ0_2;
	wire w_dff_A_vGHTfhyW9_2;
	wire w_dff_B_AzGMDA8y8_2;
	wire w_dff_B_uy03LviU8_2;
	wire w_dff_B_8e51ZPui5_2;
	wire w_dff_B_UI1HZQrx3_2;
	wire w_dff_B_ONbC3eCq1_2;
	wire w_dff_B_lfDjGvPZ0_2;
	wire w_dff_B_CMs9GZ1y0_2;
	wire w_dff_B_4fPtujk65_2;
	wire w_dff_B_mWon9R7R9_2;
	wire w_dff_B_HuA5otXH4_2;
	wire w_dff_B_31jyz91C5_2;
	wire w_dff_B_Kj3JMYLO7_2;
	wire w_dff_B_rt2susp59_2;
	wire w_dff_B_moXigPB47_2;
	wire w_dff_B_Ey2tPuqD6_2;
	wire w_dff_B_7tL7QzxS7_2;
	wire w_dff_B_k5cSsR3t0_2;
	wire w_dff_B_4755z2Hn7_2;
	wire w_dff_B_s9yo5N0r9_2;
	wire w_dff_B_OFXG6fSg7_2;
	wire w_dff_B_CFnvvsaX4_2;
	wire w_dff_B_wk8eK7oI1_2;
	wire w_dff_B_VoyoSs4I0_2;
	wire w_dff_B_NYN7OKw15_2;
	wire w_dff_B_4ld0KiXW7_2;
	wire w_dff_B_CxtvxXxF4_2;
	wire w_dff_B_ZhlFiBiX3_2;
	wire w_dff_A_PWzSKAnh2_2;
	wire w_dff_A_pJu6TLUw5_2;
	wire w_dff_A_VaawTq0Y3_2;
	wire w_dff_A_yOYMrknm3_2;
	wire w_dff_A_s6wrYOsC1_2;
	wire w_dff_A_LsHyNQB36_2;
	wire w_dff_A_48j3K6HD4_2;
	wire w_dff_A_eqg8PPEo6_2;
	wire w_dff_A_ELQkdxmX1_2;
	wire w_dff_A_uuq7jWJm9_2;
	wire w_dff_A_LBfUyJGt2_2;
	wire w_dff_A_vnLBMEmj1_2;
	wire w_dff_A_6VPhDO5v1_2;
	wire w_dff_A_RMshaW478_2;
	wire w_dff_A_ZSAPFrF88_2;
	wire w_dff_A_vKJ96aS84_2;
	wire w_dff_A_xRPTxXmC9_2;
	wire w_dff_A_Io6h3bx43_2;
	wire w_dff_A_B9ujESKV2_2;
	wire w_dff_A_B02DsWh05_2;
	wire w_dff_A_C0zyaOhS4_2;
	wire w_dff_A_7KLxEBCn3_2;
	wire w_dff_A_6QicL7n99_2;
	wire w_dff_A_tdkmqNYI7_2;
	wire w_dff_A_JaX8JiOJ9_0;
	wire w_dff_A_DWFiqVPp2_0;
	wire w_dff_A_4Y8E3njp6_0;
	wire w_dff_A_uTKog0qp3_0;
	wire w_dff_A_Yl6sBJFe7_0;
	wire w_dff_A_vrU1h5q76_0;
	wire w_dff_A_6h6MoGTq4_0;
	wire w_dff_A_3sz47knn2_0;
	wire w_dff_A_5Z5PhRWw2_0;
	wire w_dff_A_4qQJtJNU1_0;
	wire w_dff_A_qxrKAmvh1_0;
	wire w_dff_A_8SFuhkZz4_0;
	wire w_dff_A_fLt2uriD4_0;
	wire w_dff_A_XYpH9AIa3_0;
	wire w_dff_A_8HvueTtx2_0;
	wire w_dff_A_1IJ4gebr6_0;
	wire w_dff_A_yOntMPx73_0;
	wire w_dff_A_PgPS7vHF7_1;
	wire w_dff_A_U7LGI2NW6_1;
	wire w_dff_A_5H0sIIw53_1;
	wire w_dff_A_vR1YJq4y5_1;
	wire w_dff_A_E6SiKNQJ1_1;
	wire w_dff_A_Dnlmsim40_1;
	wire w_dff_A_IfxHcgWw0_1;
	wire w_dff_A_CS1XUDc44_1;
	wire w_dff_A_lgskrCNj6_1;
	wire w_dff_A_TaMCCUBL4_1;
	wire w_dff_A_cLxrOEJU8_1;
	wire w_dff_A_BhUrfjsT4_1;
	wire w_dff_A_MyMfKrmE2_1;
	wire w_dff_A_UikOBbBR2_1;
	wire w_dff_A_fEh8IIwQ7_1;
	wire w_dff_A_3qesbko21_1;
	wire w_dff_A_rZMUeqtT1_0;
	wire w_dff_A_2xZl2LHc0_0;
	wire w_dff_A_o4hKRHkh8_0;
	wire w_dff_A_fbl2CEZY5_0;
	wire w_dff_A_LmrBxr9C2_0;
	wire w_dff_A_DOIi9s5f9_0;
	wire w_dff_A_9iYeXxQm9_0;
	wire w_dff_A_DQTCx7PV6_0;
	wire w_dff_A_9pd7nHgI1_0;
	wire w_dff_A_U7Vz4sXe9_0;
	wire w_dff_A_Rk1zU4oN8_0;
	wire w_dff_A_8EcYE1yi1_0;
	wire w_dff_A_kXzompdx0_0;
	wire w_dff_A_N1qdQRdK4_0;
	wire w_dff_A_UP7Tw7xo6_0;
	wire w_dff_A_4BObyJuZ0_0;
	wire w_dff_A_9IdfYSln5_0;
	wire w_dff_A_jdP6U8b07_0;
	wire w_dff_A_kZqzrERF1_0;
	wire w_dff_A_JS09NjOF6_0;
	wire w_dff_A_izbnWL9K6_0;
	wire w_dff_A_WgQjA4mu7_0;
	wire w_dff_A_5kcqco9f3_0;
	wire w_dff_A_PW2Da1iG2_0;
	wire w_dff_A_JFty1vSw1_0;
	wire w_dff_A_Kk4Jsm8Y5_0;
	wire w_dff_A_k5hS1sGE3_1;
	wire w_dff_A_8uWlESyb2_0;
	wire w_dff_A_ZxbXG1ZX7_0;
	wire w_dff_A_XUqMXgsB7_0;
	wire w_dff_A_Ke4YvWgH0_0;
	wire w_dff_A_jyng7xC70_0;
	wire w_dff_A_Y917uZt44_0;
	wire w_dff_A_NC2HOdeJ7_0;
	wire w_dff_A_4a5o1oev5_0;
	wire w_dff_A_cYgNx4oo5_0;
	wire w_dff_A_b7edN0jj3_0;
	wire w_dff_A_XuUOAamh3_0;
	wire w_dff_A_mZbRYjb50_0;
	wire w_dff_A_PbfIIqdM0_0;
	wire w_dff_A_7pT2pHSk2_0;
	wire w_dff_A_ROW0QVMA0_0;
	wire w_dff_A_6WUchvPs2_0;
	wire w_dff_A_P1xrhZVX1_0;
	wire w_dff_A_q4ZuV6WA7_0;
	wire w_dff_A_kKeVad1S9_0;
	wire w_dff_A_IevzEcxt4_0;
	wire w_dff_A_TeifZMw32_0;
	wire w_dff_A_Xm0W3xgQ8_0;
	wire w_dff_A_vjGNUgun3_0;
	wire w_dff_A_xCMijMMy9_0;
	wire w_dff_A_6VqqoTRR5_0;
	wire w_dff_A_bVoxBf3X7_0;
	wire w_dff_A_d6kwjLVZ0_1;
	wire w_dff_A_Zs4FhmDx9_0;
	wire w_dff_A_udvjerb55_0;
	wire w_dff_A_jHunwUCV1_0;
	wire w_dff_A_ojg6VGAY8_0;
	wire w_dff_A_twwtg2867_0;
	wire w_dff_A_QQUPyo6B3_0;
	wire w_dff_A_aKnkfTMm3_0;
	wire w_dff_A_griBH8TH1_0;
	wire w_dff_A_WkKUe34a9_0;
	wire w_dff_A_cUFSCdBl4_0;
	wire w_dff_A_jV4oyZOf2_0;
	wire w_dff_A_KWia5jN18_0;
	wire w_dff_A_FV4HJGny4_0;
	wire w_dff_A_NkiHE9p90_0;
	wire w_dff_A_hD5vSv531_0;
	wire w_dff_A_mLW3L2zd3_0;
	wire w_dff_A_gTUaK7PN3_0;
	wire w_dff_A_9GUhU2QS7_0;
	wire w_dff_A_lpMKehaN0_0;
	wire w_dff_A_tLHd8NGO8_0;
	wire w_dff_A_osog69XA8_0;
	wire w_dff_A_8Y1H6pcH4_0;
	wire w_dff_A_8MYk7QEc1_0;
	wire w_dff_A_THwqZlsa1_0;
	wire w_dff_A_fzLeF5Br9_0;
	wire w_dff_A_JfqOrBRk2_0;
	wire w_dff_A_VHpW1ILW7_1;
	wire w_dff_A_0EdNBvdh9_0;
	wire w_dff_A_D4OkyQ4G9_0;
	wire w_dff_A_QfKA9iXQ7_0;
	wire w_dff_A_wOhFogC16_0;
	wire w_dff_A_UGs0r12P4_0;
	wire w_dff_A_zaSpRqku1_0;
	wire w_dff_A_dbPsrNvz1_0;
	wire w_dff_A_HoAwRdxX7_0;
	wire w_dff_A_8QFTlGAL7_0;
	wire w_dff_A_9jFSz56R8_0;
	wire w_dff_A_urHNbyaD5_0;
	wire w_dff_A_smurInE44_0;
	wire w_dff_A_cc0bom7j3_0;
	wire w_dff_A_oZePYS4c6_0;
	wire w_dff_A_Bo94DYig0_0;
	wire w_dff_A_MErWuuNG0_0;
	wire w_dff_A_pCcJklv01_0;
	wire w_dff_A_JKooQMiB5_0;
	wire w_dff_A_KKURhmtQ4_0;
	wire w_dff_A_QmFJHWQj2_0;
	wire w_dff_A_SFC6N8698_0;
	wire w_dff_A_6rukfAPk6_0;
	wire w_dff_A_YTZ4OCzy0_0;
	wire w_dff_A_OZW0BpKb4_0;
	wire w_dff_A_Pkn8qxHJ5_0;
	wire w_dff_A_PCekqYEQ0_0;
	wire w_dff_A_2GuE02g96_1;
	wire w_dff_A_0qKeY6Yy4_0;
	wire w_dff_A_P27MWUUx8_0;
	wire w_dff_A_kllTJxuw5_0;
	wire w_dff_A_XIJ9hcLF3_0;
	wire w_dff_A_uMbhdoe53_0;
	wire w_dff_A_uVwGQOzg1_0;
	wire w_dff_A_ajn1NoHo4_0;
	wire w_dff_A_ZMYKSxSU9_0;
	wire w_dff_A_4h0mS7gB3_0;
	wire w_dff_A_RrypEcrR9_0;
	wire w_dff_A_Xjea6bvo8_0;
	wire w_dff_A_QKlP35xm6_0;
	wire w_dff_A_ce8jm6bc2_0;
	wire w_dff_A_fXEt5rXm9_0;
	wire w_dff_A_HNZ1HHDk2_0;
	wire w_dff_A_cm8vsMiB2_0;
	wire w_dff_A_mN0D8Rpu3_0;
	wire w_dff_A_Q8rV6Zat7_0;
	wire w_dff_A_t7wZdGwX1_0;
	wire w_dff_A_KJ8rTuVl5_0;
	wire w_dff_A_zlVkK4YB4_0;
	wire w_dff_A_Taqzk2LZ4_0;
	wire w_dff_A_S6zLf6W24_0;
	wire w_dff_A_7r8n76n82_0;
	wire w_dff_A_GVBvY17J3_0;
	wire w_dff_A_qZdKgzVe7_0;
	wire w_dff_A_63AobLUF2_1;
	wire w_dff_A_dAlUDEjG1_0;
	wire w_dff_A_tejdBBNT0_0;
	wire w_dff_A_xzriuna22_0;
	wire w_dff_A_Mf5s9S5i2_0;
	wire w_dff_A_phDcnlxx3_0;
	wire w_dff_A_Ld3TBmQB5_0;
	wire w_dff_A_aCUV8FGK3_0;
	wire w_dff_A_ylPMQHgv6_0;
	wire w_dff_A_18iQsGit3_0;
	wire w_dff_A_HQp5Isk29_0;
	wire w_dff_A_4pNBlFnC9_0;
	wire w_dff_A_cegTMNkz5_0;
	wire w_dff_A_LuWf17Ek6_0;
	wire w_dff_A_olEg0y025_0;
	wire w_dff_A_tmqmlhJE8_0;
	wire w_dff_A_LNVrH9Rq0_0;
	wire w_dff_A_exksNRci6_0;
	wire w_dff_A_KVigNA9U1_0;
	wire w_dff_A_dAUd8jss8_0;
	wire w_dff_A_d9VRJBek8_0;
	wire w_dff_A_n6PlnGlr2_0;
	wire w_dff_A_5wiTCPxQ0_0;
	wire w_dff_A_Ne1VqeQd2_0;
	wire w_dff_A_ToJmm2N25_0;
	wire w_dff_A_Iy23Gdq82_0;
	wire w_dff_A_A0RiMfTY7_0;
	wire w_dff_A_xSrgjd2r2_1;
	wire w_dff_A_z1MV1RVm5_0;
	wire w_dff_A_NCvQSvrP0_0;
	wire w_dff_A_31ZmXWPA6_0;
	wire w_dff_A_rzdzpzl07_0;
	wire w_dff_A_8yCoMCvI6_0;
	wire w_dff_A_YwJr4WJK3_0;
	wire w_dff_A_Ow12GLnX5_0;
	wire w_dff_A_BEeT3fNA1_0;
	wire w_dff_A_258yxaEp7_0;
	wire w_dff_A_Bea28Dpj7_0;
	wire w_dff_A_gXe7JpOF8_0;
	wire w_dff_A_rRlDJQLa1_0;
	wire w_dff_A_jyi9a2ds0_0;
	wire w_dff_A_AvGh5mxf9_0;
	wire w_dff_A_DfVOl6jg6_0;
	wire w_dff_A_W1Q5HWHK8_0;
	wire w_dff_A_9QFRuSy82_0;
	wire w_dff_A_Ljxk9B0y1_0;
	wire w_dff_A_xkJtNxKY0_0;
	wire w_dff_A_RZNQa8Zp0_0;
	wire w_dff_A_sAMT18Ip3_0;
	wire w_dff_A_FOkR76ml9_0;
	wire w_dff_A_AXurrEUk1_0;
	wire w_dff_A_HhopjXlZ5_0;
	wire w_dff_A_EnmNRsPi0_0;
	wire w_dff_A_dKQThvRv8_0;
	wire w_dff_A_FJrUYRUW2_1;
	wire w_dff_A_midEEXwi6_0;
	wire w_dff_A_nEvJflSm7_0;
	wire w_dff_A_SESSf9AI6_0;
	wire w_dff_A_YsZvdVsm1_0;
	wire w_dff_A_btPF0H3W0_0;
	wire w_dff_A_M0YggQ760_0;
	wire w_dff_A_SzLWu1io6_0;
	wire w_dff_A_dZB7ziFm4_0;
	wire w_dff_A_9XyS5e731_0;
	wire w_dff_A_r8lzG5NM2_0;
	wire w_dff_A_QPF6Efy87_0;
	wire w_dff_A_sZTpVlYA9_0;
	wire w_dff_A_BNg0veXI8_0;
	wire w_dff_A_FdehvAmM2_0;
	wire w_dff_A_fs63tjHV7_0;
	wire w_dff_A_nX1Dl57M2_0;
	wire w_dff_A_gtSoiKOo4_0;
	wire w_dff_A_RMXDH7rG7_0;
	wire w_dff_A_ymzgro2G8_0;
	wire w_dff_A_eCLMDY9V5_0;
	wire w_dff_A_JmltyGqX9_0;
	wire w_dff_A_zrdcGyY85_0;
	wire w_dff_A_LRXr5ju66_0;
	wire w_dff_A_VhDntoKw5_0;
	wire w_dff_A_oGAw2bVZ4_0;
	wire w_dff_A_zYPLqGsr8_0;
	wire w_dff_A_hsW6rtkC8_1;
	wire w_dff_A_szKiCzJS1_0;
	wire w_dff_A_yJBiMRC79_0;
	wire w_dff_A_Z9VSso8D1_0;
	wire w_dff_A_gZdKDqab3_0;
	wire w_dff_A_9RZ0kxKC1_0;
	wire w_dff_A_Tf7IENfH1_0;
	wire w_dff_A_6c6RHEE55_0;
	wire w_dff_A_Cj9JVRMP3_0;
	wire w_dff_A_TWAnU5KB2_0;
	wire w_dff_A_EYi4WWD14_0;
	wire w_dff_A_Jv1Yxix80_0;
	wire w_dff_A_GezRUYTJ9_0;
	wire w_dff_A_IbrxoSpm7_0;
	wire w_dff_A_ruY906Ta4_0;
	wire w_dff_A_irFwQcnP4_0;
	wire w_dff_A_OuKPEvKB0_0;
	wire w_dff_A_7c4ZfVoG7_0;
	wire w_dff_A_N3TJd7Gp5_0;
	wire w_dff_A_tgloV8av7_0;
	wire w_dff_A_Xets2Obk2_0;
	wire w_dff_A_RKyVqdFx5_0;
	wire w_dff_A_eXir635X9_0;
	wire w_dff_A_KPIQcHyP7_0;
	wire w_dff_A_pdkIhO8J0_0;
	wire w_dff_A_GNYTEDO03_0;
	wire w_dff_A_I2luZ5AD4_0;
	wire w_dff_A_PX3V940Q1_1;
	wire w_dff_A_Szlr61vU3_0;
	wire w_dff_A_txxwIzN43_0;
	wire w_dff_A_TcaYo2gG9_0;
	wire w_dff_A_JhxAfswL4_0;
	wire w_dff_A_57InIhXx1_0;
	wire w_dff_A_qYmlp08P4_0;
	wire w_dff_A_xxcY15o56_0;
	wire w_dff_A_SyNuU87b4_0;
	wire w_dff_A_3axgsdQM0_0;
	wire w_dff_A_CHWLo9YL9_0;
	wire w_dff_A_w6Npeprv7_0;
	wire w_dff_A_iA6SLOYw2_0;
	wire w_dff_A_VpihWe7C8_0;
	wire w_dff_A_vmXYj26E5_0;
	wire w_dff_A_Wj1A375y5_0;
	wire w_dff_A_oUPPLDIT1_0;
	wire w_dff_A_fFCFGCtw3_0;
	wire w_dff_A_gxbjnoIh6_0;
	wire w_dff_A_40w87G6r0_0;
	wire w_dff_A_7Nczw42J7_0;
	wire w_dff_A_bjmRyeJX8_0;
	wire w_dff_A_D3aERHvU1_0;
	wire w_dff_A_tsTZTo0n4_0;
	wire w_dff_A_eOrHbXe88_0;
	wire w_dff_A_bmPpN7js2_0;
	wire w_dff_A_jf8spJsC9_0;
	wire w_dff_A_FpfbrbRf3_1;
	wire w_dff_A_hWBhh0uA5_0;
	wire w_dff_A_DF2pDixM4_0;
	wire w_dff_A_uuuBjRoR1_0;
	wire w_dff_A_WohuxkYd2_0;
	wire w_dff_A_Ir2xvp0x1_0;
	wire w_dff_A_afzONmUh7_0;
	wire w_dff_A_jKnjhFfZ6_0;
	wire w_dff_A_YS4lJjbE0_0;
	wire w_dff_A_sV06MLaO8_0;
	wire w_dff_A_8K2SK2cJ2_0;
	wire w_dff_A_YJ15L2IW5_0;
	wire w_dff_A_PkL00IS48_0;
	wire w_dff_A_gBzSJv3r7_0;
	wire w_dff_A_BVzplejU9_0;
	wire w_dff_A_Zj3TXxVz6_0;
	wire w_dff_A_tsCG02bx4_0;
	wire w_dff_A_D1O1SYim5_0;
	wire w_dff_A_HGvRUoVW5_0;
	wire w_dff_A_cSJqokbd4_0;
	wire w_dff_A_nwWD9v3C3_0;
	wire w_dff_A_9P9q7ot19_0;
	wire w_dff_A_QSwPkL6k4_0;
	wire w_dff_A_eo6KGMVz7_0;
	wire w_dff_A_3prTw2Z20_0;
	wire w_dff_A_ZyehewfO2_0;
	wire w_dff_A_nCxU7v4v1_0;
	wire w_dff_A_ngtpAtsY5_1;
	wire w_dff_A_dI8qiuRa9_0;
	wire w_dff_A_XS6ojzl56_0;
	wire w_dff_A_pSpZeeOU2_0;
	wire w_dff_A_xfaVxp8y8_0;
	wire w_dff_A_SQJ3DB1P9_0;
	wire w_dff_A_uzOI3sGp8_0;
	wire w_dff_A_p3Xx526u7_0;
	wire w_dff_A_WV6L8kQ13_0;
	wire w_dff_A_uexmfjaw3_0;
	wire w_dff_A_9MXOBaWj9_0;
	wire w_dff_A_I8JayFcY4_0;
	wire w_dff_A_PAx9P8q05_0;
	wire w_dff_A_4DQmtHqt2_0;
	wire w_dff_A_88KhvHXC0_0;
	wire w_dff_A_50UI5PGD0_0;
	wire w_dff_A_GkKeEPc17_0;
	wire w_dff_A_vLElKZTm0_0;
	wire w_dff_A_HBHEkfUe2_0;
	wire w_dff_A_uCqDNxO10_0;
	wire w_dff_A_QRwZmUjI4_0;
	wire w_dff_A_chnGNUjU5_0;
	wire w_dff_A_2GV3F85s8_0;
	wire w_dff_A_dnBudaaR9_0;
	wire w_dff_A_ZQ8Rg5qF5_0;
	wire w_dff_A_lq9Bm5JV2_0;
	wire w_dff_A_9T2mPAHf9_0;
	wire w_dff_A_5cfRan3F4_2;
	wire w_dff_A_TNeGIopd8_0;
	wire w_dff_A_cliTpmkT3_0;
	wire w_dff_A_DcGSxjqq2_0;
	wire w_dff_A_FV1UWYjJ3_0;
	wire w_dff_A_QhuGMRpv6_0;
	wire w_dff_A_gvTpK0tC8_0;
	wire w_dff_A_fSPPQFY42_0;
	wire w_dff_A_C8pYUjey9_0;
	wire w_dff_A_Dq5SKNWG6_0;
	wire w_dff_A_5Qp6DBuz4_0;
	wire w_dff_A_IYpkiHMX6_0;
	wire w_dff_A_WWeMLzkC5_0;
	wire w_dff_A_6bTjRrRU4_0;
	wire w_dff_A_MYVkEitD8_0;
	wire w_dff_A_cSWIX6eW9_0;
	wire w_dff_A_KGf7Iqt45_0;
	wire w_dff_A_FoV0X4GM5_0;
	wire w_dff_A_Bty9xsM37_0;
	wire w_dff_A_JufoRDEz4_0;
	wire w_dff_A_uk2DcbNv8_0;
	wire w_dff_A_3RmbsgOM2_0;
	wire w_dff_A_soGFIDx60_0;
	wire w_dff_A_0Asvl05L1_0;
	wire w_dff_A_vG3AJPai3_0;
	wire w_dff_A_2VOakzUt5_0;
	wire w_dff_A_mJOSM8RJ0_0;
	wire w_dff_A_5t6DzlqV5_1;
	wire w_dff_A_AkO6TqAN1_0;
	wire w_dff_A_0fViiNHk7_0;
	wire w_dff_A_KMSQqxDl9_0;
	wire w_dff_A_ClQuB2hj4_0;
	wire w_dff_A_56vSMsC89_0;
	wire w_dff_A_GGQcJnL39_0;
	wire w_dff_A_Ek0i76k61_0;
	wire w_dff_A_blfsYTeX7_0;
	wire w_dff_A_SSTP5gav9_0;
	wire w_dff_A_IUJH1Rzh6_0;
	wire w_dff_A_UnpMCpFA6_0;
	wire w_dff_A_toLzv5Wz8_0;
	wire w_dff_A_9cBlObww6_0;
	wire w_dff_A_rZeDuzOa5_0;
	wire w_dff_A_jzQ6eMdj7_0;
	wire w_dff_A_DjBUioum9_0;
	wire w_dff_A_CxweOoky9_0;
	wire w_dff_A_bkcEcDCz8_0;
	wire w_dff_A_Cp66eVQd7_0;
	wire w_dff_A_eljnh0Zq4_0;
	wire w_dff_A_dWtolInX2_0;
	wire w_dff_A_J9jSSohA0_0;
	wire w_dff_A_AzGZECcC4_0;
	wire w_dff_A_s23nZGQS9_0;
	wire w_dff_A_TtBkZVw68_0;
	wire w_dff_A_oLgyeFaj7_0;
	wire w_dff_A_WU84By202_1;
	wire w_dff_A_ExbZdFft7_0;
	wire w_dff_A_LipODtBL2_0;
	wire w_dff_A_IP95x7VF3_0;
	wire w_dff_A_ohwzvEnL0_0;
	wire w_dff_A_wRzVTGBz1_0;
	wire w_dff_A_M1J9ofQx9_0;
	wire w_dff_A_XxZuVF487_0;
	wire w_dff_A_8CmjZnUN6_0;
	wire w_dff_A_en6iky532_0;
	wire w_dff_A_vdY2E7GL0_0;
	wire w_dff_A_8c4tUJNl4_0;
	wire w_dff_A_9s12XcWn3_0;
	wire w_dff_A_hKg7IygA9_0;
	wire w_dff_A_KaKR3Fko9_0;
	wire w_dff_A_Dr8oBaGF7_0;
	wire w_dff_A_SzQjdAPg7_0;
	wire w_dff_A_WIXvc3nZ4_0;
	wire w_dff_A_be6sH0uC5_0;
	wire w_dff_A_2dfySpkn9_0;
	wire w_dff_A_x9n3u7oK2_0;
	wire w_dff_A_y55xJ1ku5_0;
	wire w_dff_A_Bdq7bNDo0_0;
	wire w_dff_A_7M6NhEP52_0;
	wire w_dff_A_k2LO6yXs7_0;
	wire w_dff_A_M83EPBTI6_0;
	wire w_dff_A_ZVtp3RYb3_0;
	wire w_dff_A_00yBnyGB8_1;
	wire w_dff_A_UDlJXt8c6_0;
	wire w_dff_A_LMDyBa0b8_0;
	wire w_dff_A_JjWo0d4c7_0;
	wire w_dff_A_seqQ42bY6_0;
	wire w_dff_A_9PjKnYGS6_0;
	wire w_dff_A_6NSocSQc1_0;
	wire w_dff_A_VogwunOA4_0;
	wire w_dff_A_RWtZAbBh4_0;
	wire w_dff_A_3umFCYI50_0;
	wire w_dff_A_TnSQms2s5_0;
	wire w_dff_A_m0PwIy8J4_0;
	wire w_dff_A_zxzhDAm66_0;
	wire w_dff_A_h6FErAJP6_0;
	wire w_dff_A_Vex5MC0l7_0;
	wire w_dff_A_7AhQ1E7u2_0;
	wire w_dff_A_3zbwA3tH1_0;
	wire w_dff_A_ynQ30shl7_0;
	wire w_dff_A_NbYM2WC09_0;
	wire w_dff_A_yPhRucby9_0;
	wire w_dff_A_g9U8ADko8_0;
	wire w_dff_A_xFuGE22u5_0;
	wire w_dff_A_P4hpayBY0_0;
	wire w_dff_A_hCCATq3l4_0;
	wire w_dff_A_fIboX2j20_0;
	wire w_dff_A_DHO0Yl9L6_0;
	wire w_dff_A_W4LvPFHI2_0;
	wire w_dff_A_9O4gAV2i7_1;
	wire w_dff_A_VlzhPncD2_0;
	wire w_dff_A_mAC2MZIc1_0;
	wire w_dff_A_xNV2BHgZ1_0;
	wire w_dff_A_2yPk94W95_0;
	wire w_dff_A_wrbFE21X9_0;
	wire w_dff_A_JEXyzaBW5_0;
	wire w_dff_A_WMqTFTfS4_0;
	wire w_dff_A_L2x21T8C4_0;
	wire w_dff_A_eqxLe8Ly2_0;
	wire w_dff_A_poOSoO2I6_0;
	wire w_dff_A_dPQMv4Ly5_0;
	wire w_dff_A_UTtF3snW4_0;
	wire w_dff_A_4CIW0D9p0_0;
	wire w_dff_A_2oWqbx8g0_0;
	wire w_dff_A_eGUVLsiR1_0;
	wire w_dff_A_gFoE7tEK5_0;
	wire w_dff_A_qeXe7CHZ3_0;
	wire w_dff_A_ll7FEGeB0_0;
	wire w_dff_A_yqtzfzdn2_0;
	wire w_dff_A_cGLikj2N9_0;
	wire w_dff_A_IF9OC0EY6_0;
	wire w_dff_A_EVMxK5z23_0;
	wire w_dff_A_CJUHXIz74_0;
	wire w_dff_A_LPG7EiUM4_0;
	wire w_dff_A_wd7LoYRr0_0;
	wire w_dff_A_ed7jCAqA2_0;
	wire w_dff_A_wElPQzTe5_2;
	wire w_dff_A_4AOl2UH79_0;
	wire w_dff_A_JlKtbfur3_0;
	wire w_dff_A_DkNyWvK76_0;
	wire w_dff_A_mJmbW3Cc4_0;
	wire w_dff_A_UzGttZvD9_0;
	wire w_dff_A_YNd6SKU43_0;
	wire w_dff_A_Ov1Tvs7f5_0;
	wire w_dff_A_dA0TC0dG4_0;
	wire w_dff_A_ZBWY9wqZ4_0;
	wire w_dff_A_AR1uQiiT7_0;
	wire w_dff_A_FRkgn1Go4_0;
	wire w_dff_A_QPLO1r0R1_0;
	wire w_dff_A_UBbajyiL4_0;
	wire w_dff_A_nmLoOm7U5_0;
	wire w_dff_A_cOdwUzQW6_0;
	wire w_dff_A_QGb8wMTu9_0;
	wire w_dff_A_LXWUVEv72_0;
	wire w_dff_A_qwnZtuUh2_0;
	wire w_dff_A_EhaPn7jp7_0;
	wire w_dff_A_MuPXOk6G3_0;
	wire w_dff_A_eJuhSk0E3_0;
	wire w_dff_A_uZ8yTvPd7_0;
	wire w_dff_A_eEvjbcGu3_0;
	wire w_dff_A_hUtW2DhM9_0;
	wire w_dff_A_obxRtBkU9_0;
	wire w_dff_A_0UmWNMxX9_0;
	wire w_dff_A_5ftdZgkS7_2;
	wire w_dff_A_CMaaRmQY4_0;
	wire w_dff_A_TeZA8vRj1_0;
	wire w_dff_A_bYTk6TVq9_0;
	wire w_dff_A_JtqXfOQ52_0;
	wire w_dff_A_Gl0DGDjm2_0;
	wire w_dff_A_XBCRh5Pa5_0;
	wire w_dff_A_hXemu6u64_0;
	wire w_dff_A_7qpG2OMS7_0;
	wire w_dff_A_j2lCvmCJ4_0;
	wire w_dff_A_lTi6JReR2_0;
	wire w_dff_A_9NPOSaKl7_0;
	wire w_dff_A_BrrOSoGj3_0;
	wire w_dff_A_VfwoEhfr4_0;
	wire w_dff_A_sgMNeLux8_0;
	wire w_dff_A_tuU4C99N4_0;
	wire w_dff_A_rzzQlwH61_0;
	wire w_dff_A_iGuArtNh5_0;
	wire w_dff_A_3Qf12oSp8_0;
	wire w_dff_A_8w1NMvb74_0;
	wire w_dff_A_aDNivSHy6_0;
	wire w_dff_A_yj4CGCgA1_0;
	wire w_dff_A_WrKFg0mw8_0;
	wire w_dff_A_c0JWgtOE4_0;
	wire w_dff_A_BzV8wqwf9_0;
	wire w_dff_A_4CP3EiGh6_0;
	wire w_dff_A_nNW8Oyib6_2;
	wire w_dff_A_n2FdJ63z5_0;
	wire w_dff_A_3hoEDqA48_0;
	wire w_dff_A_sysUsWEc8_0;
	wire w_dff_A_CYim9ad56_0;
	wire w_dff_A_bbMcMkbS4_0;
	wire w_dff_A_usgfN2SQ1_0;
	wire w_dff_A_ZHwqDeh71_0;
	wire w_dff_A_23SLu1YI9_0;
	wire w_dff_A_i3VyskVW1_0;
	wire w_dff_A_dtyqkMfr6_0;
	wire w_dff_A_U7dZrVpH5_0;
	wire w_dff_A_1KddJRVb4_0;
	wire w_dff_A_9Y8SiPe14_0;
	wire w_dff_A_cNKUpofq4_0;
	wire w_dff_A_uFhzg1g85_0;
	wire w_dff_A_Im1meCHG2_0;
	wire w_dff_A_oTmKnql35_0;
	wire w_dff_A_UtBCzH9v6_0;
	wire w_dff_A_eiCgoMAU3_0;
	wire w_dff_A_6lobc3xM7_0;
	wire w_dff_A_z3VMAUdJ6_0;
	wire w_dff_A_1sDwaukh1_0;
	wire w_dff_A_jfUiw9GR5_0;
	wire w_dff_A_ubHt4fJJ2_0;
	wire w_dff_A_lshyIWXp2_0;
	wire w_dff_A_IZSXO4y19_1;
	wire w_dff_A_FdvWJKLi8_0;
	wire w_dff_A_DrzRPN2R6_0;
	wire w_dff_A_2lRx43hP9_0;
	wire w_dff_A_32fzlnBH8_0;
	wire w_dff_A_7DbEmEQ39_0;
	wire w_dff_A_n1W7Q6ga7_0;
	wire w_dff_A_nP5pYstd3_0;
	wire w_dff_A_XSXuxrB71_0;
	wire w_dff_A_QCC3DIq40_0;
	wire w_dff_A_45UY7L592_0;
	wire w_dff_A_M4L6E43p3_0;
	wire w_dff_A_vmM6rYJd2_0;
	wire w_dff_A_ACNoAteu2_0;
	wire w_dff_A_wNhRjP6A5_0;
	wire w_dff_A_S0oksRfg3_0;
	wire w_dff_A_JZIrDp5I0_0;
	wire w_dff_A_KicmJWUX2_0;
	wire w_dff_A_PgAkvC1X2_0;
	wire w_dff_A_8gATiKRr1_0;
	wire w_dff_A_pgriklao0_0;
	wire w_dff_A_X5LgeMM37_0;
	wire w_dff_A_8HS1W8TA4_0;
	wire w_dff_A_lEUlsqKZ1_0;
	wire w_dff_A_KDgHikqk8_0;
	wire w_dff_A_BoNDu9p83_0;
	wire w_dff_A_tBsHYMsf0_1;
	wire w_dff_A_Di9tBEy93_0;
	wire w_dff_A_FRrNlEBd4_0;
	wire w_dff_A_KDHxzONX2_0;
	wire w_dff_A_tb6xgNvv2_0;
	wire w_dff_A_16iSviNr2_0;
	wire w_dff_A_rlu5irWz5_0;
	wire w_dff_A_2TB6mGr13_0;
	wire w_dff_A_yIYqBvIk8_0;
	wire w_dff_A_nL8meCCM3_0;
	wire w_dff_A_fqKWxqRr2_0;
	wire w_dff_A_NUY8XYjB8_0;
	wire w_dff_A_gAw9JrmO5_0;
	wire w_dff_A_abkL6C4w1_0;
	wire w_dff_A_7fPhmR1o3_0;
	wire w_dff_A_ieokOxlL6_0;
	wire w_dff_A_xmzZY5IA8_0;
	wire w_dff_A_lL5ppykf2_0;
	wire w_dff_A_1fZ3Z1300_0;
	wire w_dff_A_A7DEkHDH2_0;
	wire w_dff_A_sdzZicac3_0;
	wire w_dff_A_vn2J0xgn3_0;
	wire w_dff_A_moB7jOxG0_0;
	wire w_dff_A_MpMlg4gU8_0;
	wire w_dff_A_E8J6kf2r8_0;
	wire w_dff_A_hyqtacLo7_0;
	wire w_dff_A_fchFTvy15_0;
	wire w_dff_A_tPCLe9f04_1;
	wire w_dff_A_APa8b5xU3_0;
	wire w_dff_A_0kTMdKbI4_0;
	wire w_dff_A_AUCit7yg7_0;
	wire w_dff_A_QZ0dxaob8_0;
	wire w_dff_A_t9fDaZFZ9_0;
	wire w_dff_A_XEpRULQ03_0;
	wire w_dff_A_66Gf8kif4_0;
	wire w_dff_A_rHx8OWQg6_0;
	wire w_dff_A_mcoIyVux9_0;
	wire w_dff_A_s69KssoD8_0;
	wire w_dff_A_NFtq4UzW4_0;
	wire w_dff_A_UHkfVC438_0;
	wire w_dff_A_w0cdKska7_0;
	wire w_dff_A_odd9nTRY5_0;
	wire w_dff_A_BQ1Z48kf7_0;
	wire w_dff_A_nvUjCZu32_0;
	wire w_dff_A_nLZSCQ2u2_0;
	wire w_dff_A_aqnbexse8_0;
	wire w_dff_A_sk1Spi356_0;
	wire w_dff_A_pb3IABQT4_0;
	wire w_dff_A_ouqLDWaW0_0;
	wire w_dff_A_01kzzUme9_0;
	wire w_dff_A_KXvKvncn6_0;
	wire w_dff_A_ClpyFt7J9_0;
	wire w_dff_A_aZQfPyvd9_0;
	wire w_dff_A_dafibjqx9_0;
	wire w_dff_A_mnbyVjQA2_1;
	wire w_dff_A_Jm13IGCP0_0;
	wire w_dff_A_fhbz7wsS6_0;
	wire w_dff_A_UlAn2Kdo1_0;
	wire w_dff_A_J3GvyTlB8_0;
	wire w_dff_A_cBNDgBw72_0;
	wire w_dff_A_5kuH9gVS2_0;
	wire w_dff_A_b052TarJ5_0;
	wire w_dff_A_NzKOpNRB5_0;
	wire w_dff_A_L5yaxj4p3_0;
	wire w_dff_A_317FVENG8_0;
	wire w_dff_A_LKKJsjVo7_0;
	wire w_dff_A_bCx5BuDl4_0;
	wire w_dff_A_6DjmhvjB9_0;
	wire w_dff_A_DWYFI0Vn2_0;
	wire w_dff_A_7e0zUIbQ6_0;
	wire w_dff_A_lOZo7eb14_0;
	wire w_dff_A_wP2WmMbE2_0;
	wire w_dff_A_mwwNQD667_0;
	wire w_dff_A_f462eIbp7_0;
	wire w_dff_A_6gt7HUvI4_0;
	wire w_dff_A_wjDFJL4O0_0;
	wire w_dff_A_vieZz9Ka5_0;
	wire w_dff_A_1qpbX8co8_0;
	wire w_dff_A_2bmp3zIS0_0;
	wire w_dff_A_RcPgZUiL4_0;
	wire w_dff_A_knvHDWqy4_0;
	wire w_dff_A_HsXSJqmW2_1;
	wire w_dff_A_OKpwcyB81_0;
	wire w_dff_A_3F3vAHQd6_0;
	wire w_dff_A_rggA0Xjo4_0;
	wire w_dff_A_vtwirMfd2_0;
	wire w_dff_A_uSiiAwV32_0;
	wire w_dff_A_MMk7vI6F0_0;
	wire w_dff_A_XJfbGET98_0;
	wire w_dff_A_enUVeP9G1_0;
	wire w_dff_A_RW2z4dJ44_0;
	wire w_dff_A_9Cm7KGQt9_0;
	wire w_dff_A_BoATiG8v7_0;
	wire w_dff_A_65ZGevFm9_0;
	wire w_dff_A_URTE9TmN8_0;
	wire w_dff_A_HfyHt0xL1_0;
	wire w_dff_A_TUWilLHJ6_0;
	wire w_dff_A_myPRZoEq7_0;
	wire w_dff_A_N51r9fdv0_0;
	wire w_dff_A_zunUBKVQ0_0;
	wire w_dff_A_NX7Px3B18_0;
	wire w_dff_A_0eb4s6Ac5_0;
	wire w_dff_A_wKPSXQ9S5_0;
	wire w_dff_A_WS8MKiuX9_0;
	wire w_dff_A_HW2uTXjD8_0;
	wire w_dff_A_01lhwsU58_0;
	wire w_dff_A_UyJWuDAO7_0;
	wire w_dff_A_mfr6wMuy6_0;
	wire w_dff_A_YrcMuZjh5_1;
	wire w_dff_A_jhEr5zGS5_0;
	wire w_dff_A_vjbUvAEs7_0;
	wire w_dff_A_yLelHxPb9_0;
	wire w_dff_A_ZDCQfVVY7_0;
	wire w_dff_A_CXROt8NI0_0;
	wire w_dff_A_u0KRek7n0_0;
	wire w_dff_A_sB0yXDSc6_0;
	wire w_dff_A_fiLpjyuf1_0;
	wire w_dff_A_rUUSTHGH2_0;
	wire w_dff_A_WLXMhlYe7_0;
	wire w_dff_A_mN1szGLP0_0;
	wire w_dff_A_kulQlXRO5_0;
	wire w_dff_A_iiseMS9g5_0;
	wire w_dff_A_q4JDALdd1_0;
	wire w_dff_A_Ld6FerP87_0;
	wire w_dff_A_rlfMbOL13_0;
	wire w_dff_A_3pIkzwlY5_0;
	wire w_dff_A_CSqsZH544_0;
	wire w_dff_A_XX0lVAs04_0;
	wire w_dff_A_5ljnhUSX1_0;
	wire w_dff_A_9wXbLuQx4_0;
	wire w_dff_A_Mj3Yn2ok4_0;
	wire w_dff_A_gKOno9Oj4_0;
	wire w_dff_A_UIzerzom4_0;
	wire w_dff_A_mSOx0lHj4_0;
	wire w_dff_A_8xdMCJWG0_0;
	wire w_dff_A_i0f25SsS5_1;
	wire w_dff_A_EaoC9uBY9_0;
	wire w_dff_A_SSYifb0q5_0;
	wire w_dff_A_fxEzwhkz5_0;
	wire w_dff_A_gImH4YvO7_0;
	wire w_dff_A_mx8rY8fB6_0;
	wire w_dff_A_BjcwPdQA4_0;
	wire w_dff_A_pPx2SNbI8_0;
	wire w_dff_A_uyXOxEBR7_0;
	wire w_dff_A_8rO5yTEq1_0;
	wire w_dff_A_w57orzIn7_0;
	wire w_dff_A_ob5EmfXZ0_0;
	wire w_dff_A_vJT2ArS15_0;
	wire w_dff_A_5iai8qls3_0;
	wire w_dff_A_UxVvbBJv4_0;
	wire w_dff_A_XRKPOS2V9_0;
	wire w_dff_A_Vcg7Vzz66_0;
	wire w_dff_A_z3FQ501J3_0;
	wire w_dff_A_wtDX4HwP1_0;
	wire w_dff_A_iR93SuQP7_0;
	wire w_dff_A_AqdjrelI3_0;
	wire w_dff_A_VHv4GM3C5_0;
	wire w_dff_A_H8DPBpjF6_0;
	wire w_dff_A_VJ3md6VJ3_0;
	wire w_dff_A_tzFXcQsT8_0;
	wire w_dff_A_3mgvfYY55_0;
	wire w_dff_A_Tt7Kreo86_0;
	wire w_dff_A_pkH3YkUJ5_2;
	wire w_dff_A_bVproxhZ1_0;
	wire w_dff_A_NnggmJRV8_0;
	wire w_dff_A_Dtng7xtL1_0;
	wire w_dff_A_VzWPLMQo1_0;
	wire w_dff_A_5peywzLZ3_0;
	wire w_dff_A_FknypKjz8_0;
	wire w_dff_A_zYJzvywN2_0;
	wire w_dff_A_8d2IWV7w7_0;
	wire w_dff_A_syANXWzw9_0;
	wire w_dff_A_mQRD1Het5_0;
	wire w_dff_A_oz7vJrKv5_0;
	wire w_dff_A_2gabycod7_0;
	wire w_dff_A_RLZewH0M7_0;
	wire w_dff_A_SQ4fMz7y7_0;
	wire w_dff_A_P9lMhNpW4_0;
	wire w_dff_A_SbWgZuYa5_0;
	wire w_dff_A_3p5gu8aV5_0;
	wire w_dff_A_XlJ7iejh3_0;
	wire w_dff_A_LyygyGZP6_0;
	wire w_dff_A_n6ByNeGz2_0;
	wire w_dff_A_4Uq4ytKh1_0;
	wire w_dff_A_C9Nwdp014_0;
	wire w_dff_A_EpQxD4l68_0;
	wire w_dff_A_LcbV2KB71_0;
	wire w_dff_A_f2GSdHvr4_2;
	wire w_dff_A_4GI2vdTM9_0;
	wire w_dff_A_9DPRFH3j1_0;
	wire w_dff_A_brnb3pLh2_0;
	wire w_dff_A_4LTPbnYX6_0;
	wire w_dff_A_432jsq1W8_0;
	wire w_dff_A_Nv5oegAo6_0;
	wire w_dff_A_l7UkE0E24_0;
	wire w_dff_A_E7QuBlZJ4_0;
	wire w_dff_A_TwXQ17uT1_0;
	wire w_dff_A_orOK3QiK0_0;
	wire w_dff_A_OqWgzCzh6_0;
	wire w_dff_A_ck27aEon9_0;
	wire w_dff_A_LlKry5MB5_0;
	wire w_dff_A_GvQS4EHy0_0;
	wire w_dff_A_k3ETe60u0_0;
	wire w_dff_A_mY05oQWp8_0;
	wire w_dff_A_txr2TGNJ1_0;
	wire w_dff_A_HhBUpIvU3_0;
	wire w_dff_A_RmNhbpNS3_0;
	wire w_dff_A_KJrxWuKz7_0;
	wire w_dff_A_ab98WgBp3_0;
	wire w_dff_A_FEs7AWUG6_0;
	wire w_dff_A_BmlfKb2Z0_0;
	wire w_dff_A_5zh3mgN75_0;
	wire w_dff_A_t57oU9fo7_0;
	wire w_dff_A_jBXFRELh6_1;
	wire w_dff_A_O4279mhi6_0;
	wire w_dff_A_gkLomz2O2_0;
	wire w_dff_A_5IO90M1b1_0;
	wire w_dff_A_w25WQnhG5_0;
	wire w_dff_A_Al5wD0XM5_0;
	wire w_dff_A_WUt9Obbs2_0;
	wire w_dff_A_IEARGc4p8_0;
	wire w_dff_A_oCdrQpEF4_0;
	wire w_dff_A_0P59qezH7_0;
	wire w_dff_A_tf3dk7eV5_0;
	wire w_dff_A_eU0hxtQK5_0;
	wire w_dff_A_J8ltMfCs6_0;
	wire w_dff_A_qO1vkvcG9_0;
	wire w_dff_A_xSu0o2Jz4_0;
	wire w_dff_A_m7EMncmL0_0;
	wire w_dff_A_rbuAS3CU6_0;
	wire w_dff_A_7Z6O8Y0J9_0;
	wire w_dff_A_WX9bIBWT6_0;
	wire w_dff_A_cIln2rmy5_0;
	wire w_dff_A_Rrj2gw9F6_0;
	wire w_dff_A_F36pxWCQ3_0;
	wire w_dff_A_kEDOBLfu4_0;
	wire w_dff_A_loYdKfFg6_0;
	wire w_dff_A_nO5ramgs1_0;
	wire w_dff_A_xxC0s3NU1_0;
	wire w_dff_A_x4ak0bCm9_0;
	wire w_dff_A_AOkWbxaA9_1;
	wire w_dff_A_UrKL7IBP3_0;
	wire w_dff_A_OCoDPrgc0_0;
	wire w_dff_A_ID8Ltcb10_0;
	wire w_dff_A_Mz87F2Wy8_0;
	wire w_dff_A_HspfVHHf7_0;
	wire w_dff_A_zX0zbdhB7_0;
	wire w_dff_A_DlXVKrQM3_0;
	wire w_dff_A_og3hDeDi0_0;
	wire w_dff_A_Y8uGbWbG4_0;
	wire w_dff_A_sTDa7OYi2_0;
	wire w_dff_A_eWh4NSQ39_0;
	wire w_dff_A_BXFX4jj31_0;
	wire w_dff_A_Jnkop36Y9_0;
	wire w_dff_A_Vmxipy6w2_0;
	wire w_dff_A_Ok8Y0cGv1_0;
	wire w_dff_A_uwv5k4xR7_0;
	wire w_dff_A_qADDLnHx0_0;
	wire w_dff_A_kgcBYuEQ4_0;
	wire w_dff_A_rAveruXr9_0;
	wire w_dff_A_uQBIO8VC7_0;
	wire w_dff_A_WFc12DKO2_0;
	wire w_dff_A_Tr9ThHPu3_0;
	wire w_dff_A_cMjBiDnC8_0;
	wire w_dff_A_e5yMkLbO6_0;
	wire w_dff_A_NvcJmCpU8_0;
	wire w_dff_A_bBfrkhR76_0;
	wire w_dff_A_8UBzqmtz1_1;
	wire w_dff_A_xAMmuwKd7_0;
	wire w_dff_A_FCy7xAyr4_0;
	wire w_dff_A_hiaAwhs56_0;
	wire w_dff_A_9aQqzs390_0;
	wire w_dff_A_V4O7HvQ07_0;
	wire w_dff_A_6dOjmLPT6_0;
	wire w_dff_A_RArkxi7X6_0;
	wire w_dff_A_lryukamR8_0;
	wire w_dff_A_a6ocVgTp5_0;
	wire w_dff_A_HnBEWdAw3_0;
	wire w_dff_A_dJ5c2YAM4_0;
	wire w_dff_A_RZhauPO90_0;
	wire w_dff_A_cFFHib127_0;
	wire w_dff_A_7QR5pUC97_0;
	wire w_dff_A_YP6GqKyh1_0;
	wire w_dff_A_Z3yLKJJr0_0;
	wire w_dff_A_n8oRfgRV9_0;
	wire w_dff_A_0l0E9Php1_0;
	wire w_dff_A_JOz6Y5zA2_0;
	wire w_dff_A_xgNSg37t8_0;
	wire w_dff_A_MDeAfenL1_0;
	wire w_dff_A_IUkC6Joo2_0;
	wire w_dff_A_b3V2Ghm33_0;
	wire w_dff_A_yvOhH7523_0;
	wire w_dff_A_t2vfrKCz6_0;
	wire w_dff_A_BoOOBYC89_0;
	wire w_dff_A_SKPLdeyi8_1;
	wire w_dff_A_2qSTzhyE9_0;
	wire w_dff_A_nucsXvpf2_0;
	wire w_dff_A_pJq5yQqh4_0;
	wire w_dff_A_wu97i3l88_0;
	wire w_dff_A_5S0JHsZ41_0;
	wire w_dff_A_z7kyIMWU7_0;
	wire w_dff_A_PDVDedOh3_0;
	wire w_dff_A_WVwJhwtm7_0;
	wire w_dff_A_YwIrpcYa1_0;
	wire w_dff_A_xHz7VYgs1_0;
	wire w_dff_A_jXAdoxY40_0;
	wire w_dff_A_OmOWHH8i7_0;
	wire w_dff_A_u15K7vWv4_0;
	wire w_dff_A_tLPxEEPG4_0;
	wire w_dff_A_SalfHBKp8_0;
	wire w_dff_A_X20frKLI7_0;
	wire w_dff_A_ZA4oBV7I1_0;
	wire w_dff_A_keFdkTBZ4_0;
	wire w_dff_A_wH64j8n76_0;
	wire w_dff_A_qrSLvkpL6_0;
	wire w_dff_A_23jIzKqa0_0;
	wire w_dff_A_xymuw4o74_0;
	wire w_dff_A_pD3W7Z586_0;
	wire w_dff_A_JFYKppkd0_0;
	wire w_dff_A_CcltRsG24_0;
	wire w_dff_A_B2DvfHSf5_0;
	wire w_dff_A_Femo9NLV5_1;
	wire w_dff_A_NlHBCzV31_0;
	wire w_dff_A_wg5gnJ2k1_0;
	wire w_dff_A_P479h9P96_0;
	wire w_dff_A_HqpFnqCb7_0;
	wire w_dff_A_PvnhAJg39_0;
	wire w_dff_A_LZll5Fm78_0;
	wire w_dff_A_0z4SIJqg6_0;
	wire w_dff_A_IFWuuGx01_0;
	wire w_dff_A_XSxmljR30_0;
	wire w_dff_A_BrKoEwES3_0;
	wire w_dff_A_rYEawTOG9_0;
	wire w_dff_A_a7fR5RQd1_0;
	wire w_dff_A_4IOJGG5X4_0;
	wire w_dff_A_W9iTcZTk2_0;
	wire w_dff_A_65rT7D2V2_0;
	wire w_dff_A_FswOCQ1x5_0;
	wire w_dff_A_rr1mzzEm5_0;
	wire w_dff_A_LzvWqzG99_0;
	wire w_dff_A_qHF1pcbb0_0;
	wire w_dff_A_OUaEY0X33_0;
	wire w_dff_A_0iAljFpq4_0;
	wire w_dff_A_YPIditjM1_0;
	wire w_dff_A_EN3CGhBf4_0;
	wire w_dff_A_W6UzBvUa9_0;
	wire w_dff_A_0gxnXOPP4_0;
	wire w_dff_A_0NxvzrgN0_0;
	wire w_dff_A_JlUsfOTy7_1;
	wire w_dff_A_3B9HwBPe0_0;
	wire w_dff_A_yStGtaew4_0;
	wire w_dff_A_jaLX8CQ02_0;
	wire w_dff_A_67wNSxP11_0;
	wire w_dff_A_GegosreC5_0;
	wire w_dff_A_XHWoNeFP3_0;
	wire w_dff_A_bLfiJvCO4_0;
	wire w_dff_A_BS0uVRY25_0;
	wire w_dff_A_kVvwKqRh3_0;
	wire w_dff_A_XGBQ3QtX9_0;
	wire w_dff_A_MMY6qRtf4_0;
	wire w_dff_A_j4alQXXo8_0;
	wire w_dff_A_riaw58ne8_0;
	wire w_dff_A_MN2uMMIk9_0;
	wire w_dff_A_XRWpcieE0_0;
	wire w_dff_A_0IZ2WCww9_0;
	wire w_dff_A_jKIJe3Cs1_0;
	wire w_dff_A_Eon0llJ00_0;
	wire w_dff_A_I302w8E71_0;
	wire w_dff_A_WbLeyYaB7_0;
	wire w_dff_A_WkftCjGB1_0;
	wire w_dff_A_mPYVDaIn7_0;
	wire w_dff_A_rzLVcdgv7_0;
	wire w_dff_A_xL5DAQUP6_0;
	wire w_dff_A_iTB1BQ4n3_0;
	wire w_dff_A_lzRGMTWg1_0;
	wire w_dff_A_ggxnG5mk7_2;
	wire w_dff_A_soGqoBSU8_0;
	wire w_dff_A_a0JslDTl1_0;
	wire w_dff_A_zpTnZla65_0;
	wire w_dff_A_tTRpNvXs0_0;
	wire w_dff_A_bjOdwmAc2_0;
	wire w_dff_A_YJ9ZAu3J6_0;
	wire w_dff_A_PixvskVl1_0;
	wire w_dff_A_p3qbVq8r3_0;
	wire w_dff_A_aW56xJAs5_0;
	wire w_dff_A_3Wlp8vE85_0;
	wire w_dff_A_E8mM1muW5_0;
	wire w_dff_A_SLFWPjY44_0;
	wire w_dff_A_J8kL7Sgt9_0;
	wire w_dff_A_sw8PUaHd1_0;
	wire w_dff_A_KIuylHh73_0;
	wire w_dff_A_sHYEi02l3_0;
	wire w_dff_A_yUvjfvIO8_0;
	wire w_dff_A_px2WHpYM5_0;
	wire w_dff_A_zRF8JdTh0_0;
	wire w_dff_A_9DUo6PBV2_0;
	wire w_dff_A_sgrLK5Oe7_0;
	wire w_dff_A_8zEUF1Kx6_0;
	wire w_dff_A_r5BCFrqL9_0;
	wire w_dff_A_9Fp90GiW7_2;
	wire w_dff_A_wkmp6lrl8_0;
	wire w_dff_A_Om9gIXYj8_0;
	wire w_dff_A_J8bKEIoc2_0;
	wire w_dff_A_1IR9LRMQ0_0;
	wire w_dff_A_Q27Pe5oZ8_0;
	wire w_dff_A_pmrRKuYQ3_0;
	wire w_dff_A_HZstU9Dd0_0;
	wire w_dff_A_3MOpmkng3_0;
	wire w_dff_A_zYDO4QhQ1_0;
	wire w_dff_A_CgGxoC2F7_0;
	wire w_dff_A_qWBRdyc79_0;
	wire w_dff_A_D1H3cY1Z2_0;
	wire w_dff_A_0l9AKiTB8_0;
	wire w_dff_A_XEqDzIra2_0;
	wire w_dff_A_SWGWLOGt5_0;
	wire w_dff_A_g2POdUbn9_0;
	wire w_dff_A_n3wg9EoG8_0;
	wire w_dff_A_tk4VvaVL2_0;
	wire w_dff_A_ViiQ19Ro7_0;
	wire w_dff_A_snizAxlQ4_0;
	wire w_dff_A_gQzsw8tX0_0;
	wire w_dff_A_ySsGHG3o4_0;
	wire w_dff_A_eJEs7m0C0_0;
	wire w_dff_A_BaD8i8TF9_2;
	wire w_dff_A_xjBKTD4I1_0;
	wire w_dff_A_6YM20goG0_0;
	wire w_dff_A_MElF77n31_0;
	wire w_dff_A_xDGqj1qa7_0;
	wire w_dff_A_gMJ0bC1b7_0;
	wire w_dff_A_OZD5cGSG7_0;
	wire w_dff_A_dgKvcHDk1_0;
	wire w_dff_A_PqCbBv3R6_0;
	wire w_dff_A_fAYB8dnB5_0;
	wire w_dff_A_JP7SyptP2_0;
	wire w_dff_A_KI5jhp3e5_0;
	wire w_dff_A_zwuUHvm75_0;
	wire w_dff_A_otvnUqrg0_0;
	wire w_dff_A_NJ3uvGoa6_0;
	wire w_dff_A_3mvlPVQ53_0;
	wire w_dff_A_DDumhluL6_0;
	wire w_dff_A_8IuzqLEW7_0;
	wire w_dff_A_boPSc9fI5_0;
	wire w_dff_A_ESwuOz9u6_0;
	wire w_dff_A_UANjooBs1_0;
	wire w_dff_A_ADvYnNf58_0;
	wire w_dff_A_1CiA6Af43_0;
	wire w_dff_A_tzjUCfjA9_0;
	wire w_dff_A_7aIGYmBt8_2;
	wire w_dff_A_fdslbe5r7_0;
	wire w_dff_A_bgmIoIfr6_0;
	wire w_dff_A_eB9DO8Xr2_0;
	wire w_dff_A_FztlOzVp5_0;
	wire w_dff_A_GKY3LsMV0_0;
	wire w_dff_A_iNwDsvSD2_0;
	wire w_dff_A_xER18dRt8_0;
	wire w_dff_A_Vw79pbN41_0;
	wire w_dff_A_eD7oyL8r7_0;
	wire w_dff_A_QnfkqptZ9_0;
	wire w_dff_A_qkJJt8qk1_0;
	wire w_dff_A_v32xaZdh5_0;
	wire w_dff_A_EpydQUZR8_0;
	wire w_dff_A_oIQ15tVM3_0;
	wire w_dff_A_FecwbBKd7_0;
	wire w_dff_A_DJp5nEX43_0;
	wire w_dff_A_fagqzMmt2_0;
	wire w_dff_A_t6mYyL5t3_0;
	wire w_dff_A_fdUuXirF3_0;
	wire w_dff_A_sc2fG96P1_0;
	wire w_dff_A_lm5H9nBY1_0;
	wire w_dff_A_adDaodPF2_0;
	wire w_dff_A_RpYPwKbW1_0;
	wire w_dff_A_22ycq4ex2_0;
	wire w_dff_A_oXh5hHFP5_2;
	wire w_dff_A_4LtYUCoT8_0;
	wire w_dff_A_4iVz71ut0_0;
	wire w_dff_A_IWIDMaw86_0;
	wire w_dff_A_XkkHFvoO4_0;
	wire w_dff_A_IaQB31nO0_0;
	wire w_dff_A_CfsQocWg1_0;
	wire w_dff_A_eHgmuEbK1_0;
	wire w_dff_A_pqbmqe2y1_0;
	wire w_dff_A_lcQfdGmx4_0;
	wire w_dff_A_8QrI6YU44_0;
	wire w_dff_A_nX2fVv7i5_0;
	wire w_dff_A_2lH3SzDG5_0;
	wire w_dff_A_JjVnmOAe2_0;
	wire w_dff_A_uWwO6c0V0_0;
	wire w_dff_A_Scr4Xdlr9_0;
	wire w_dff_A_MNmT17kz0_0;
	wire w_dff_A_4NhZrj4o5_0;
	wire w_dff_A_Z3M9vFrv1_0;
	wire w_dff_A_HweYZHgk8_0;
	wire w_dff_A_yykWYldi2_0;
	wire w_dff_A_9OoTzEzV7_0;
	wire w_dff_A_Zlckauki5_0;
	wire w_dff_A_4VBlrx7w2_2;
	wire w_dff_A_BIlgfuI73_0;
	wire w_dff_A_uXeSAsFX3_0;
	wire w_dff_A_VomWAx9P1_0;
	wire w_dff_A_sRlKKdnF4_0;
	wire w_dff_A_duknT22U1_0;
	wire w_dff_A_HALbsMQM1_0;
	wire w_dff_A_qKlXLPIF0_0;
	wire w_dff_A_VXSzI9iX9_0;
	wire w_dff_A_xcijaDCS4_0;
	wire w_dff_A_5X1gZXtG7_0;
	wire w_dff_A_lRDBTsYm8_0;
	wire w_dff_A_MYOlMxxt1_0;
	wire w_dff_A_JdmnnDJw6_0;
	wire w_dff_A_Dn4OQfkn4_0;
	wire w_dff_A_6ygsp5KJ0_0;
	wire w_dff_A_rh6YIwCc6_0;
	wire w_dff_A_S0F2NR0R8_0;
	wire w_dff_A_FwX7Takh2_0;
	wire w_dff_A_N3KcFBa32_0;
	wire w_dff_A_LoEkIqHu8_0;
	wire w_dff_A_euh4H7FH7_0;
	wire w_dff_A_McPKAUHR9_0;
	wire w_dff_A_TnyExUOt6_2;
	wire w_dff_A_m2QxoPEi7_0;
	wire w_dff_A_6DCS2fUy9_0;
	wire w_dff_A_QxOHOkW36_0;
	wire w_dff_A_jyRVJxNl4_0;
	wire w_dff_A_BUaKj3Nn2_0;
	wire w_dff_A_Ti9mOnCh1_0;
	wire w_dff_A_VuWBPtCy4_0;
	wire w_dff_A_NFPZ5n9V4_0;
	wire w_dff_A_QyhQHejV1_0;
	wire w_dff_A_HtsmvrZi3_0;
	wire w_dff_A_T4XC26Jg7_0;
	wire w_dff_A_nFvlLH8c1_0;
	wire w_dff_A_OShEDruo9_0;
	wire w_dff_A_GGdVLRBB7_0;
	wire w_dff_A_rFgGl2NK4_0;
	wire w_dff_A_VahjnZhW6_0;
	wire w_dff_A_DEaQaxxT2_0;
	wire w_dff_A_gUfDPPDN6_0;
	wire w_dff_A_8afGv2pz2_0;
	wire w_dff_A_3lv0jjFW6_0;
	wire w_dff_A_YmzDT3ym0_0;
	wire w_dff_A_IfE1XxdW2_0;
	wire w_dff_A_jviPCy004_2;
	wire w_dff_A_04uaOXrN9_0;
	wire w_dff_A_UdbLiJgG5_0;
	wire w_dff_A_MzDfdB4P0_0;
	wire w_dff_A_SxgIrgyv4_0;
	wire w_dff_A_MHWEKNgO1_0;
	wire w_dff_A_WGdGq7Ey9_0;
	wire w_dff_A_OxGqiwtK2_0;
	wire w_dff_A_y1IPsVse8_0;
	wire w_dff_A_2B6Q3m830_0;
	wire w_dff_A_LX8HlE9g4_0;
	wire w_dff_A_xk5ejCSe6_0;
	wire w_dff_A_BaoSDj0W1_0;
	wire w_dff_A_5cs0LYHE3_0;
	wire w_dff_A_Ex6JadYn8_0;
	wire w_dff_A_fTvKbmDP0_0;
	wire w_dff_A_4mydeKCB9_0;
	wire w_dff_A_0ozEw7dI5_0;
	wire w_dff_A_K9IfZtmH3_0;
	wire w_dff_A_rJ51SNR76_0;
	wire w_dff_A_4YzD4k2h4_0;
	wire w_dff_A_dYaBkdA04_0;
	wire w_dff_A_u6GnkU9e7_0;
	wire w_dff_A_FCzrs7lI1_2;
	wire w_dff_A_ahcWene33_0;
	wire w_dff_A_E4ut34AA3_0;
	wire w_dff_A_lZiDdcn39_0;
	wire w_dff_A_irKjk10M5_0;
	wire w_dff_A_7ouXLBM22_0;
	wire w_dff_A_GP3KJ3lY1_0;
	wire w_dff_A_0rpV5NER2_0;
	wire w_dff_A_M6Sqze256_0;
	wire w_dff_A_yZ8dW7Bl7_0;
	wire w_dff_A_Cbq7JKkt2_0;
	wire w_dff_A_3zy9uUce6_0;
	wire w_dff_A_gLx2fgw39_0;
	wire w_dff_A_GvvLizGC0_0;
	wire w_dff_A_MfhM0JDk7_0;
	wire w_dff_A_yLhM6FhX1_0;
	wire w_dff_A_Gvzo9Uf08_0;
	wire w_dff_A_IOssKhkH6_0;
	wire w_dff_A_h5pezWX06_0;
	wire w_dff_A_54HgQfUU5_0;
	wire w_dff_A_w6ptbcNI1_2;
	wire w_dff_A_wKcYnG6L0_0;
	wire w_dff_A_WLfds1zs2_0;
	wire w_dff_A_t8op28g67_0;
	wire w_dff_A_JHfpfx4h0_0;
	wire w_dff_A_2RMLKFdb4_0;
	wire w_dff_A_DDD1tYNc4_0;
	wire w_dff_A_s0hmulKZ0_0;
	wire w_dff_A_A9p0smSx1_0;
	wire w_dff_A_Cj9sbDPR6_0;
	wire w_dff_A_Kod3pKDV5_0;
	wire w_dff_A_7xhQmYh16_0;
	wire w_dff_A_vG0ZTohM3_0;
	wire w_dff_A_QvoG1XTB6_0;
	wire w_dff_A_e1pzCSdJ9_0;
	wire w_dff_A_CzWkz3IL9_0;
	wire w_dff_A_bhbvxTPo5_0;
	wire w_dff_A_YBZbAwDs7_0;
	wire w_dff_A_bi0nBdus6_0;
	wire w_dff_A_hjs3pf4K4_2;
	wire w_dff_A_xktMmrAI2_0;
	wire w_dff_A_B0XsbOgY5_0;
	wire w_dff_A_hSHgTJH43_0;
	wire w_dff_A_bhUEti0a3_0;
	wire w_dff_A_LFUSm4GD1_0;
	wire w_dff_A_uUDNsvUN0_0;
	wire w_dff_A_ypLymG1f1_0;
	wire w_dff_A_Wl3MkFn20_0;
	wire w_dff_A_JT2tdUVw6_0;
	wire w_dff_A_OHzqKTJu2_0;
	wire w_dff_A_Kmwsm5hn3_0;
	wire w_dff_A_1hSgZx2J6_0;
	wire w_dff_A_mtPWx4Va4_0;
	wire w_dff_A_DmnnXYYn4_0;
	wire w_dff_A_UJa8BsNY4_0;
	wire w_dff_A_l2uks8bl3_0;
	wire w_dff_A_QVvvToBY8_2;
	wire w_dff_A_r8UDSSn76_0;
	wire w_dff_A_6fgyXfer9_0;
	wire w_dff_A_zTl1PCT15_0;
	wire w_dff_A_favJvT4u8_0;
	wire w_dff_A_udDgwovk2_0;
	wire w_dff_A_fikQLPbe8_0;
	wire w_dff_A_QRgNZbL06_0;
	wire w_dff_A_A1BnklJE4_0;
	wire w_dff_A_ZOKzsVmy0_0;
	wire w_dff_A_L6JCwsmY9_0;
	wire w_dff_A_VdTOdjVu4_0;
	wire w_dff_A_1haxGdVJ2_0;
	wire w_dff_A_wZD9eGAg9_0;
	wire w_dff_A_Kvt6v9Sw6_0;
	wire w_dff_A_6Glt6atn6_0;
	wire w_dff_A_bzvNBOYj0_0;
	wire w_dff_A_6BM5FR752_0;
	wire w_dff_A_VyRNnbsR6_2;
	wire w_dff_A_8v0iwfKN0_0;
	wire w_dff_A_5c3an98c5_0;
	wire w_dff_A_eP0RgtWU9_0;
	wire w_dff_A_2lkPwFN80_0;
	wire w_dff_A_ara8B4DS4_0;
	wire w_dff_A_JkxiWNce1_0;
	wire w_dff_A_yo4P0xeu7_0;
	wire w_dff_A_5BWg8Psx7_0;
	wire w_dff_A_c08IIq7k5_0;
	wire w_dff_A_vjE7kXum4_0;
	wire w_dff_A_OACUKO5e1_0;
	wire w_dff_A_EIFAbSCw3_0;
	wire w_dff_A_Uns95WFP8_0;
	wire w_dff_A_ywLwuiAb9_0;
	wire w_dff_A_dQbOsoUn7_0;
	wire w_dff_A_y1Id65Fp3_0;
	wire w_dff_A_LwtLdMpv7_0;
	wire w_dff_A_RZ4RQ0L23_2;
	wire w_dff_A_txr7Wh484_0;
	wire w_dff_A_fn7ZApTB9_0;
	wire w_dff_A_iJ58sCCY4_0;
	wire w_dff_A_mWkPQRQa3_0;
	wire w_dff_A_WSB7tngo1_0;
	wire w_dff_A_xgaQshQA7_0;
	wire w_dff_A_BVDzHZaB2_0;
	wire w_dff_A_O1jl03pm7_0;
	wire w_dff_A_4IB0tKDg2_0;
	wire w_dff_A_iGAv61P90_0;
	wire w_dff_A_y24CL9Za1_0;
	wire w_dff_A_kZduCUAf2_0;
	wire w_dff_A_JTr66KAw8_0;
	wire w_dff_A_K6d8Q3cU9_0;
	wire w_dff_A_yoJGiT3X1_0;
	wire w_dff_A_BlRKl12i8_0;
	wire w_dff_A_lYUtd87F9_1;
	wire w_dff_A_bwbB4dfk5_0;
	wire w_dff_A_8gTHU8iS2_0;
	wire w_dff_A_BvnYNZOB3_0;
	wire w_dff_A_QyN45Ac36_0;
	wire w_dff_A_BxAN3miV1_0;
	wire w_dff_A_Too8TLhh7_0;
	wire w_dff_A_jz0cGITH3_0;
	wire w_dff_A_w6kU9sVE5_0;
	wire w_dff_A_QRrpYB9c1_0;
	wire w_dff_A_FUU9QeKu5_0;
	wire w_dff_A_TBPKl1lf1_0;
	wire w_dff_A_UYjP4O1j9_0;
	wire w_dff_A_AZEwqLtC2_0;
	wire w_dff_A_wjOrQWWf2_0;
	wire w_dff_A_rAk1AOeY4_0;
	wire w_dff_A_sV3M7dZY7_0;
	wire w_dff_A_mQ3bit1g5_0;
	wire w_dff_A_KcNSmz6o9_0;
	wire w_dff_A_hOU7wK100_0;
	wire w_dff_A_aHLi1u3A8_0;
	wire w_dff_A_DGGQpU6e9_0;
	wire w_dff_A_GVvo75fl8_0;
	wire w_dff_A_tW43U9KN1_1;
	wire w_dff_A_7s0FSjaT0_0;
	wire w_dff_A_NBBiu6xp2_0;
	wire w_dff_A_moFeEk9L8_0;
	wire w_dff_A_u35H4Nyf2_0;
	wire w_dff_A_XBD0ESze7_0;
	wire w_dff_A_6PKRrom93_0;
	wire w_dff_A_jHLZZbYD8_0;
	wire w_dff_A_3SyNmhWU4_0;
	wire w_dff_A_w04x8hvn5_0;
	wire w_dff_A_rQy1K00S9_0;
	wire w_dff_A_FTsbSBtP3_0;
	wire w_dff_A_NVQh7i3k5_0;
	wire w_dff_A_GQzo0G338_0;
	wire w_dff_A_fvr5Y7cP2_0;
	wire w_dff_A_rASdqLYY9_0;
	wire w_dff_A_ZOroC7IB1_0;
	wire w_dff_A_A3B0aA2U6_0;
	wire w_dff_A_Oo3iQI7s2_0;
	wire w_dff_A_vnD58Lnw5_0;
	wire w_dff_A_3eEVLCv52_0;
	wire w_dff_A_x4WjN8389_0;
	wire w_dff_A_DAIpVBCT2_0;
	wire w_dff_A_vKR5DkTS6_2;
	wire w_dff_A_l2Yh8SJN9_0;
	wire w_dff_A_hZpNyaxf5_0;
	wire w_dff_A_q48AADeD4_0;
	wire w_dff_A_KZ6E29cY1_0;
	wire w_dff_A_agM5eRlM2_0;
	wire w_dff_A_GTUDroBe6_0;
	wire w_dff_A_74FdOBZp5_0;
	wire w_dff_A_KQ0wm0q25_0;
	wire w_dff_A_imkArTzf6_0;
	wire w_dff_A_ylvXNnnE9_0;
	wire w_dff_A_T0qagvLT7_0;
	wire w_dff_A_MFYl9Z271_0;
	wire w_dff_A_vaK6s1wt0_0;
	wire w_dff_A_XZnSM4Bv2_2;
	wire w_dff_A_oGdPn1nK8_0;
	wire w_dff_A_5Ce3RTXV1_0;
	wire w_dff_A_lA1EDnP07_0;
	wire w_dff_A_PV3IfrPl2_0;
	wire w_dff_A_f1PNTAgp5_0;
	wire w_dff_A_wHyvzA8D8_0;
	wire w_dff_A_lo68ThQf3_0;
	wire w_dff_A_ZTqyAL0G6_0;
	wire w_dff_A_2S9IQ4Vn5_0;
	wire w_dff_A_2tJdZ4Iw1_0;
	wire w_dff_A_3Svn1WWl9_0;
	wire w_dff_A_SgNjeYdC0_0;
	wire w_dff_A_GqrtkXJw6_0;
	wire w_dff_A_BxyG4Isx5_0;
	wire w_dff_A_B0akqYdF7_2;
	wire w_dff_A_qvv5I8vh5_0;
	wire w_dff_A_Rt79gU1P5_0;
	wire w_dff_A_U7OSUIat9_0;
	wire w_dff_A_BB1WxiYa9_0;
	wire w_dff_A_Tqmo8nN45_0;
	wire w_dff_A_NrzH5RsR3_0;
	wire w_dff_A_VMqkaL9U6_0;
	wire w_dff_A_thk2pDGw4_0;
	wire w_dff_A_TAC9M9JF0_0;
	wire w_dff_A_iksfG1dY1_0;
	wire w_dff_A_UZitD0P75_0;
	wire w_dff_A_tjDiisG77_0;
	wire w_dff_A_PCsd5L9P9_0;
	wire w_dff_A_Znsu090U2_2;
	wire w_dff_A_HUDI3Dhr7_0;
	wire w_dff_A_QhGHobqZ0_0;
	wire w_dff_A_c3eQQTJu4_0;
	wire w_dff_A_hz8SHt0D4_0;
	wire w_dff_A_sh5jV3hW6_0;
	wire w_dff_A_1XTfuPD71_0;
	wire w_dff_A_hBPpjwvc4_0;
	wire w_dff_A_TfHZUdBq6_0;
	wire w_dff_A_wHMlGAhe1_0;
	wire w_dff_A_Gf2jRHr16_0;
	wire w_dff_A_sqN5JeLQ7_0;
	wire w_dff_A_hxVwygIH9_0;
	wire w_dff_A_JDnLuERo5_0;
	wire w_dff_A_QHnbNUT07_0;
	wire w_dff_A_hgFfuhYA3_1;
	wire w_dff_A_wAgdn2DK8_0;
	wire w_dff_A_8EZQGkaj3_0;
	wire w_dff_A_6HeZkhuj6_0;
	wire w_dff_A_UWlpq2183_0;
	wire w_dff_A_njN7BIqv7_0;
	wire w_dff_A_3KS7syv66_0;
	wire w_dff_A_5o9JObNK3_0;
	wire w_dff_A_6TMyAyPJ9_0;
	wire w_dff_A_Q196gJ983_0;
	wire w_dff_A_YX4Gu2rD1_0;
	wire w_dff_A_o7Y8otNz4_0;
	wire w_dff_A_J3fltsUP7_0;
	wire w_dff_A_XjWylWI51_0;
	wire w_dff_A_rGc7iKsR2_0;
	wire w_dff_A_Wd7ai7VE9_0;
	wire w_dff_A_0H6mhUGq6_0;
	wire w_dff_A_8TAhpgxJ2_0;
	wire w_dff_A_FwMUFPoV6_0;
	wire w_dff_A_kKS3FP4J0_0;
	wire w_dff_A_9ExCEcXI6_1;
	wire w_dff_A_eULcMGbE2_0;
	wire w_dff_A_5WNC0i9U5_0;
	wire w_dff_A_LOuHhHfj4_0;
	wire w_dff_A_AOIUlj3i0_0;
	wire w_dff_A_wxpy3BVI8_0;
	wire w_dff_A_pdWw09zv8_0;
	wire w_dff_A_KQP8SEZB1_0;
	wire w_dff_A_7CfHCbMw1_0;
	wire w_dff_A_tDp8novG2_0;
	wire w_dff_A_rwGFPfjV1_0;
	wire w_dff_A_CPYOVB9c5_0;
	wire w_dff_A_QEwFEsPo3_0;
	wire w_dff_A_KQ3X0ZOR6_0;
	wire w_dff_A_dv6LnonX7_0;
	wire w_dff_A_an0UBJ8I1_1;
	wire w_dff_A_gUBJuViZ4_0;
	wire w_dff_A_EG4FM7dn2_0;
	wire w_dff_A_hqKisNM08_0;
	wire w_dff_A_7m5xpbTN7_0;
	wire w_dff_A_jufIAScu7_0;
	wire w_dff_A_pAAohuZF1_0;
	wire w_dff_A_JzpEgPu87_0;
	wire w_dff_A_TKvq1jPF5_0;
	wire w_dff_A_CX8VlSlG2_0;
	wire w_dff_A_0a0JOHZa0_0;
	wire w_dff_A_QL9xJwti7_0;
	wire w_dff_A_kfqdzEDL3_0;
	wire w_dff_A_2XRKEYz92_0;
	wire w_dff_A_wSJYx65l6_0;
	wire w_dff_A_MVi9QUKQ4_0;
	wire w_dff_A_rbsSBUxY7_0;
	wire w_dff_A_6hXiobxC6_0;
	wire w_dff_A_J3A90Aak2_1;
	wire w_dff_A_095S7ZBa5_0;
	wire w_dff_A_ESVnY7PM7_0;
	wire w_dff_A_GOSnef3m9_0;
	wire w_dff_A_Vbzm2oFo6_0;
	wire w_dff_A_xxznfzh42_0;
	wire w_dff_A_oK2HLNsr3_0;
	wire w_dff_A_WhBfwYZv5_0;
	wire w_dff_A_rNfutp1c7_0;
	wire w_dff_A_TatpMFv50_0;
	wire w_dff_A_PsMfZTAJ4_2;
	wire w_dff_A_AZvzbllH8_0;
	wire w_dff_A_1LBFoYk27_0;
	wire w_dff_A_GvaxARSZ6_0;
	wire w_dff_A_RGKrigig4_0;
	wire w_dff_A_22YHxR059_0;
	wire w_dff_A_eifgiYac8_0;
	wire w_dff_A_RtUT9neU7_0;
	wire w_dff_A_oSiMinqj7_0;
	wire w_dff_A_iKvcm3a23_0;
	wire w_dff_A_nZEMvpum1_0;
	wire w_dff_A_IxD0SVC77_0;
	wire w_dff_A_HVknhIRf2_0;
	wire w_dff_A_9n7I7ANS1_0;
	wire w_dff_A_lbSS0iQn2_1;
	wire w_dff_A_sCQVAFv34_0;
	wire w_dff_A_nmGTiiY77_0;
	wire w_dff_A_Hq1NbPsd3_0;
	wire w_dff_A_zMQESlBm2_0;
	wire w_dff_A_gMPz0CsY7_0;
	wire w_dff_A_brNZPAFR7_0;
	wire w_dff_A_v6oYvakf3_0;
	wire w_dff_A_6i2p1qVP1_0;
	wire w_dff_A_uChanSAJ6_0;
	wire w_dff_A_jI2swj6e0_0;
	wire w_dff_A_UUzW6DcE1_0;
	wire w_dff_A_3qqKZWbw7_0;
	wire w_dff_A_D28W5EYA0_1;
	wire w_dff_A_p0u4xb6B4_0;
	wire w_dff_A_eFblj2Xf9_0;
	wire w_dff_A_quJ1lWA34_0;
	wire w_dff_A_C1xp1yR35_0;
	wire w_dff_A_0Lj3NiCX0_0;
	wire w_dff_A_gTNtLMVa8_0;
	wire w_dff_A_SiWz9tmd0_0;
	wire w_dff_A_3LcXvDW19_0;
	wire w_dff_A_p4evVdpo6_0;
	wire w_dff_A_KTLNCtdL9_0;
	wire w_dff_A_zOelNpH78_0;
	wire w_dff_A_NzvvGosU3_0;
	wire w_dff_A_DKQ6jBI75_0;
	wire w_dff_A_4PavxOpF1_1;
	wire w_dff_A_Qv8LXOZe8_0;
	wire w_dff_A_I4BcIiKF5_0;
	wire w_dff_A_HR1U3KUx8_0;
	wire w_dff_A_anHhA3nr4_0;
	wire w_dff_A_9Aen7PEI7_0;
	wire w_dff_A_J0I4b43A6_0;
	wire w_dff_A_uZTXq8lc1_0;
	wire w_dff_A_iIueJcY23_0;
	wire w_dff_A_GoJv94Cg9_0;
	wire w_dff_A_TVBGNKJm3_0;
	wire w_dff_A_z73FdqE16_0;
	wire w_dff_A_WbPvDGwR3_0;
	wire w_dff_A_7j605oDE4_0;
	wire w_dff_A_gfl235sD6_0;
	wire w_dff_A_XbWshpzL5_0;
	wire w_dff_A_uCgvuOjA0_2;
	wire w_dff_A_v0jJKr6S3_0;
	wire w_dff_A_XrzYRPur9_0;
	wire w_dff_A_wlbXbTYG4_0;
	wire w_dff_A_62uB0t0e8_0;
	wire w_dff_A_CwDC2akM7_0;
	wire w_dff_A_tloivukf8_0;
	wire w_dff_A_wPEG65Sn7_0;
	wire w_dff_A_W9HPife25_0;
	wire w_dff_A_1ewGm17r1_0;
	wire w_dff_A_hPvTzWf08_0;
	wire w_dff_A_8HJp41DM4_0;
	wire w_dff_A_xMM7kB9L9_0;
	wire w_dff_A_SkCjaWIe4_0;
	wire w_dff_A_PwVeE3Jp6_1;
	wire w_dff_A_vvDe9zXd5_0;
	wire w_dff_A_D7X7ut397_0;
	wire w_dff_A_l8GjwcZV4_0;
	wire w_dff_A_3rMJ9UZe3_0;
	wire w_dff_A_xgoXUh0e2_0;
	wire w_dff_A_7o2950PG1_0;
	wire w_dff_A_GQn8F1U73_0;
	wire w_dff_A_h8qWiK589_0;
	wire w_dff_A_N75vCvc63_0;
	wire w_dff_A_rZhRhsc42_0;
	wire w_dff_A_OidMD6HS4_0;
	wire w_dff_A_xk218FQj0_0;
	wire w_dff_A_ORWvyfmF9_1;
	wire w_dff_A_NTttsbUL7_0;
	wire w_dff_A_OyKzx4fv1_0;
	wire w_dff_A_bMXasXir8_0;
	wire w_dff_A_2tKugoVb1_0;
	wire w_dff_A_RcngK7Hr4_0;
	wire w_dff_A_Qo4FkX5p5_0;
	wire w_dff_A_VjyYokhV5_0;
	wire w_dff_A_52Dt3Y2q1_0;
	wire w_dff_A_Q1CVm3Fv4_0;
	wire w_dff_A_O6Qpz3XO9_0;
	wire w_dff_A_tPCvkRa59_0;
	wire w_dff_A_EPsyu48S8_0;
	wire w_dff_A_jYA1aPvp5_0;
	wire w_dff_A_4MmVsxrl7_0;
	wire w_dff_A_lkGGGKZR7_1;
	wire w_dff_A_hI1Tcukw9_0;
	wire w_dff_A_iBqs50su2_0;
	wire w_dff_A_nX7Q4mEr4_0;
	wire w_dff_A_dBjPSm9l5_0;
	wire w_dff_A_3AnIbj842_0;
	wire w_dff_A_eIEMQ4sF1_0;
	wire w_dff_A_qlFVpBF09_0;
	wire w_dff_A_deqvx5Zb0_0;
	wire w_dff_A_MkKoFrcX8_0;
	wire w_dff_A_fio9PFVt0_0;
	wire w_dff_A_iAyjbgUq2_0;
	wire w_dff_A_A9GE2VRZ3_0;
	wire w_dff_A_WVPwuZV38_0;
	wire w_dff_A_83uEDLpM4_0;
	wire w_dff_A_LYLIQECz2_0;
	wire w_dff_A_y5o85UER5_1;
	wire w_dff_A_g1MK8hkL5_0;
	wire w_dff_A_T9WIBBTr5_0;
	wire w_dff_A_eSKIkpYy0_0;
	wire w_dff_A_moeM5zwB5_0;
	wire w_dff_A_kvuU1oFX2_0;
	wire w_dff_A_CFAsKBJq7_0;
	wire w_dff_A_4EIEZhWY3_0;
	wire w_dff_A_SWEKU9a34_0;
	wire w_dff_A_Nhj46LBa6_0;
	wire w_dff_A_7hpTfjw56_0;
	wire w_dff_A_o2a6b3xQ4_0;
	wire w_dff_A_5KMMxAwb2_0;
	wire w_dff_A_pqSbxMkD1_0;
	wire w_dff_A_eEBuOLFI7_0;
	wire w_dff_A_mR46Ugkq4_0;
	wire w_dff_A_dCiS2op41_0;
	wire w_dff_A_32pOtW9D1_1;
	wire w_dff_A_XddnKyiD5_0;
	wire w_dff_A_OoJRoECC9_0;
	wire w_dff_A_nD75eIp11_0;
	wire w_dff_A_aFRatdU13_0;
	wire w_dff_A_lW3A9Ekv9_0;
	wire w_dff_A_9695fvsc5_0;
	wire w_dff_A_S3U6ijvB5_0;
	wire w_dff_A_f70mi43T6_0;
	wire w_dff_A_ESCMdPsy2_0;
	wire w_dff_A_ES9gYQ6i5_0;
	wire w_dff_A_Z7PbR7z03_0;
	wire w_dff_A_dpReoaM02_0;
	wire w_dff_A_onUMXk6V9_0;
	wire w_dff_A_Tz4jAXf56_0;
	wire w_dff_A_aIQslsMW3_0;
	wire w_dff_A_xvWGgnOV7_0;
	wire w_dff_A_cLzWTcj00_0;
	wire w_dff_A_csnrMbGv0_0;
	wire w_dff_A_cLd5Q0cP9_0;
	wire w_dff_A_DX0Mtc6R2_1;
	wire w_dff_A_nTfjI0cF2_0;
	wire w_dff_A_ryLxFFBv7_0;
	wire w_dff_A_7yPlVLkp1_0;
	wire w_dff_A_ZERoUCzr9_0;
	wire w_dff_A_JWwDsi4h2_0;
	wire w_dff_A_6ZUh4y4v1_0;
	wire w_dff_A_16vCrZbw8_0;
	wire w_dff_A_FSZwXZ276_0;
	wire w_dff_A_hK9kiUZD7_0;
	wire w_dff_A_wW4156Sl2_0;
	wire w_dff_A_6Opw3FZL5_0;
	wire w_dff_A_fxiYAWL33_0;
	wire w_dff_A_WklZoigz0_0;
	wire w_dff_A_WQgKZmDb2_0;
	wire w_dff_A_mAjVlnfA4_0;
	wire w_dff_A_Qcn33iHW0_0;
	wire w_dff_A_6WPFaNR41_0;
	wire w_dff_A_micxCBgF9_0;
	wire w_dff_A_WTTfnauU2_2;
	wire w_dff_A_qiNPFECI1_0;
	wire w_dff_A_wUORH9CY2_0;
	wire w_dff_A_N39xu8ts0_0;
	wire w_dff_A_mIlpv17y8_0;
	wire w_dff_A_qm8ipQwt3_0;
	wire w_dff_A_5Wi4odPO4_0;
	wire w_dff_A_LVK68FTZ8_0;
	wire w_dff_A_RJ18dgvy4_2;
	wire w_dff_A_ickgKFvR1_0;
	wire w_dff_A_01GTjzFh5_0;
	wire w_dff_A_pLEqq7yX9_0;
	wire w_dff_A_26apLcSj0_0;
	wire w_dff_A_csXTs7Yw4_0;
	wire w_dff_A_pmWRA6JS0_0;
	wire w_dff_A_cgdxqHwN3_2;
	wire w_dff_A_aoyZcCuj3_0;
	wire w_dff_A_6ish0ona2_0;
	wire w_dff_A_0ZF7D4nz8_0;
	wire w_dff_A_y9XzhXBi3_0;
	wire w_dff_A_JIkxsbV44_0;
	wire w_dff_A_NNzvW05A4_0;
	wire w_dff_A_ioNsIhzp4_0;
	wire w_dff_A_pekoyJtn2_0;
	wire w_dff_A_0KlY1cIq4_0;
	wire w_dff_A_pSp5ibAu8_0;
	wire w_dff_A_oMrIBUE60_0;
	wire w_dff_A_7W4GWUDP1_2;
	wire w_dff_A_xvOKcKuY6_0;
	wire w_dff_A_8kfcHEHr0_0;
	wire w_dff_A_66JR4QGx3_0;
	wire w_dff_A_qbl5jmXt5_0;
	wire w_dff_A_Rjm9jPqe8_0;
	wire w_dff_A_IdYvVSNC8_0;
	wire w_dff_A_DzCJnUyy5_0;
	wire w_dff_A_nuMBE6R39_0;
	wire w_dff_A_W8lInqRb8_0;
	wire w_dff_A_9U9Fyhuk2_0;
	wire w_dff_A_iBAJdm7G7_0;
	wire w_dff_A_GBVcLEQV9_2;
	wire w_dff_A_DWhri1bT0_0;
	wire w_dff_A_HHLtTfzI9_0;
	wire w_dff_A_EW1wDWNf1_0;
	wire w_dff_A_ppKmVk3i2_0;
	wire w_dff_A_h1qgAggJ6_0;
	wire w_dff_A_kFWA9HyF6_0;
	wire w_dff_A_chlM9X4k7_0;
	wire w_dff_A_nBX0wvip1_2;
	wire w_dff_A_Y6zRAHiT2_0;
	wire w_dff_A_gsqUxdvN0_0;
	wire w_dff_A_LN3kr5iU5_0;
	wire w_dff_A_hgH6Jr8k8_0;
	wire w_dff_A_oa1i2zPk6_0;
	wire w_dff_A_alPBq42p3_0;
	wire w_dff_A_7d2cgz226_0;
	wire w_dff_A_gvDaQNL11_0;
	wire w_dff_A_7if5Ex0z2_2;
	wire w_dff_A_AiUgCs3j2_0;
	wire w_dff_A_TwTHJyww3_0;
	wire w_dff_A_IvKZmHXa9_0;
	wire w_dff_A_pxTGSbKb4_0;
	wire w_dff_A_iB2f7KVS4_0;
	wire w_dff_A_Evi6oj1V5_0;
	wire w_dff_A_kB58hnys1_0;
	wire w_dff_A_2Rc8y7wi0_0;
	wire w_dff_A_FePXc5eJ4_0;
	wire w_dff_A_a8Qk4bxx1_0;
	wire w_dff_A_esKhrEUJ8_2;
	wire w_dff_A_5DTFfIwR9_0;
	wire w_dff_A_0vWcoYRv3_0;
	wire w_dff_A_TvWaKho87_0;
	wire w_dff_A_SGB4ZzDu8_0;
	wire w_dff_A_wydLsCJt6_0;
	wire w_dff_A_qg0TwOd41_0;
	wire w_dff_A_titBxf2B9_0;
	wire w_dff_A_kXSjycLt2_0;
	wire w_dff_A_7YUUNSrQ2_0;
	wire w_dff_A_Zo2KDTfC2_2;
	wire w_dff_A_Sz9vAu1E6_0;
	wire w_dff_A_3CMRcvsG8_0;
	wire w_dff_A_guSCZ5V70_0;
	wire w_dff_A_utjEpEXv7_0;
	wire w_dff_A_07LDldsB9_0;
	wire w_dff_A_8AryYicP2_0;
	wire w_dff_A_5kDxmMZn0_0;
	wire w_dff_A_AdHQiQye7_2;
	wire w_dff_A_AhJMBAbg8_0;
	wire w_dff_A_I6U6F1X47_0;
	wire w_dff_A_WRvWehwM1_0;
	wire w_dff_A_FOVkeETD8_0;
	wire w_dff_A_8PdqdZtj4_0;
	wire w_dff_A_LBw97b4V0_0;
	wire w_dff_A_XcBEXdFK7_0;
	wire w_dff_A_R7He8G2k5_0;
	wire w_dff_A_JuenzXYu0_2;
	wire w_dff_A_M3DLpiA72_0;
	wire w_dff_A_PmQtesJW5_0;
	wire w_dff_A_uWF7OVIf0_0;
	wire w_dff_A_5orXmOyV5_0;
	wire w_dff_A_IS7AgNOe9_0;
	wire w_dff_A_ylGy2fok4_0;
	wire w_dff_A_eq05BWI14_0;
	wire w_dff_A_Zr4QqwU15_0;
	wire w_dff_A_zrmWGPMr4_0;
	wire w_dff_A_qu9L4y1s5_0;
	wire w_dff_A_Oq5Agr8v8_2;
	wire w_dff_A_zfoHNcgE4_0;
	wire w_dff_A_LlrZNhX42_0;
	wire w_dff_A_53MU5xUe5_0;
	wire w_dff_A_oG3gG4hH5_0;
	wire w_dff_A_H6Wft9bg2_0;
	wire w_dff_A_CBOLz7UP0_0;
	wire w_dff_A_atVMBKUE6_0;
	wire w_dff_A_AoKy7gAF3_0;
	wire w_dff_A_QVX67lTB4_0;
	wire w_dff_A_oXtvQCRh0_2;
	wire w_dff_A_AFy31fML3_0;
	wire w_dff_A_yLTkF0KQ9_0;
	wire w_dff_A_UZ72JWAY2_0;
	wire w_dff_A_9pnHBrWs3_0;
	wire w_dff_A_zry6GCFm8_0;
	wire w_dff_A_h9veY0Y49_0;
	wire w_dff_A_kmX7ykt16_2;
	wire w_dff_A_8c1TUqnO7_0;
	wire w_dff_A_eKQkdrWr5_0;
	wire w_dff_A_LYkqClVd5_0;
	wire w_dff_A_5YXDiOFk2_0;
	wire w_dff_A_MjXwIlmF3_0;
	wire w_dff_A_LoHZeWOW8_0;
	wire w_dff_A_yyGcsfkC2_0;
	wire w_dff_A_65IWDiCl7_0;
	wire w_dff_A_cytpHSzO3_0;
	wire w_dff_A_hZ4sVGkq1_2;
	wire w_dff_A_udKfIzWQ4_0;
	wire w_dff_A_vejniamN9_0;
	wire w_dff_A_neo7xxPE8_0;
	wire w_dff_A_YHclVrpf8_0;
	wire w_dff_A_ceJUF5kM6_0;
	wire w_dff_A_bUP0NYwP1_0;
	wire w_dff_A_ucfcjsAp5_0;
	wire w_dff_A_TRamPBMB1_0;
	wire w_dff_A_11QVwRVB7_0;
	wire w_dff_A_IObyZMPk5_2;
	wire w_dff_A_4QyUmgVw0_0;
	wire w_dff_A_StUcGH4c1_0;
	wire w_dff_A_MSnstR2G4_0;
	wire w_dff_A_CWFexcX38_0;
	wire w_dff_A_J7X7YSBc0_0;
	wire w_dff_A_lEPF0NfB0_0;
	wire w_dff_A_T75FYnvw5_0;
	wire w_dff_A_uS2qjpmo0_0;
	wire w_dff_A_GYTpg0iA4_2;
	wire w_dff_A_qr71TKgs6_0;
	wire w_dff_A_fCCOpQyt7_0;
	wire w_dff_A_JvJfqCJj5_0;
	wire w_dff_A_hYM606gy2_0;
	wire w_dff_A_jCghNv7G4_0;
	wire w_dff_A_8eEJ4Fst4_2;
	wire w_dff_A_z29pUF2q2_0;
	wire w_dff_A_ABvZrmUz6_0;
	wire w_dff_A_9gxXs9RW4_0;
	wire w_dff_A_ZR5Hs4fi9_0;
	wire w_dff_A_VbV0U5Qh2_0;
	wire w_dff_A_Otgs3z9w2_0;
	wire w_dff_A_OjxKfTJd9_0;
	wire w_dff_A_3TeE7m7O3_0;
	wire w_dff_A_P5M5q3K66_0;
	wire w_dff_A_2N0KkA108_2;
	wire w_dff_A_DeXEoGm77_0;
	wire w_dff_A_jRRsxoCY2_0;
	wire w_dff_A_jMVx26Eo7_0;
	wire w_dff_A_u7lIUA0f9_0;
	wire w_dff_A_OXHogqZl0_0;
	wire w_dff_A_aFDQzf0f6_0;
	wire w_dff_A_Pe7egUoa6_0;
	wire w_dff_A_YuQ5v5OO5_0;
	wire w_dff_A_CF9Du5FX7_0;
	wire w_dff_A_gyEHSMrf9_2;
	wire w_dff_A_nUEvxDSH5_0;
	wire w_dff_A_6gwONjtW0_0;
	wire w_dff_A_p98PBW9Q3_0;
	wire w_dff_A_MG9fIiLi9_0;
	wire w_dff_A_xScfjUXN6_0;
	wire w_dff_A_n5ZA8VPH5_0;
	wire w_dff_A_tuWa77KN8_0;
	wire w_dff_A_ubA97bsl7_0;
	wire w_dff_A_6D6rviAx0_2;
	wire w_dff_A_go1YCpUD8_0;
	wire w_dff_A_d0mWpsIG6_0;
	wire w_dff_A_d1AauKi04_0;
	wire w_dff_A_VnZF5srs2_0;
	wire w_dff_A_tsj9VRhx1_0;
	wire w_dff_A_8ZQBge4d2_0;
	wire w_dff_A_yfUFm8z19_2;
	wire w_dff_A_ipkVkOPj4_0;
	wire w_dff_A_nktSdCDh8_0;
	wire w_dff_A_WdVzl2oX6_0;
	wire w_dff_A_DsKGo98l7_0;
	wire w_dff_A_rNDqtyMM3_0;
	wire w_dff_A_ARy93q053_0;
	wire w_dff_A_pkJbzM3e8_0;
	wire w_dff_A_61roVGaG6_0;
	wire w_dff_A_uaOdc2z75_0;
	wire w_dff_A_JP0ztOG01_1;
	wire w_dff_A_XteXsbNS7_0;
	wire w_dff_A_3J3C8zlF7_0;
	wire w_dff_A_IbKSO0nV9_0;
	wire w_dff_A_0i01aeYu0_0;
	wire w_dff_A_mHR4cvL27_0;
	wire w_dff_A_gHpjmiQs1_0;
	wire w_dff_A_BfQNuq0O6_1;
	wire w_dff_A_XBmdcbDl4_0;
	wire w_dff_A_KFbpGayW2_0;
	wire w_dff_A_K8ITLv3f5_0;
	wire w_dff_A_MqXftXCi9_0;
	wire w_dff_A_QVQFkG3y9_0;
	wire w_dff_A_JlobzhOr4_0;
	wire w_dff_A_U2IuuViG0_0;
	wire w_dff_A_EMYGxBMS3_1;
	wire w_dff_A_2JoAGth54_0;
	wire w_dff_A_U3tmic7N8_0;
	wire w_dff_A_BP2h6ADM8_0;
	wire w_dff_A_hm9aLquT5_0;
	wire w_dff_A_MdeDkIKL4_0;
	wire w_dff_A_PC2vSuin3_0;
	wire w_dff_A_lO1QpRnm5_1;
	wire w_dff_A_gSlZSXwH6_0;
	wire w_dff_A_4oM9h1By1_0;
	wire w_dff_A_602QKs9Q0_0;
	wire w_dff_A_SdQ38IQz7_0;
	wire w_dff_A_HT0lfgmT0_0;
	wire w_dff_A_sJPm82kd9_0;
	wire w_dff_A_3NYxN2fx2_0;
	wire w_dff_A_rrEDsG667_0;
	wire w_dff_A_jRoTd1a24_0;
	wire w_dff_A_ElkFPYjj3_0;
	wire w_dff_A_bVfZZB9E3_0;
	wire w_dff_A_895FGv130_2;
	wire w_dff_A_iYY8G84B7_0;
	wire w_dff_A_wAm89jr86_0;
	wire w_dff_A_onCEKMEY6_0;
	wire w_dff_A_ofDz5DV79_0;
	wire w_dff_A_64wp8i3q5_0;
	wire w_dff_A_XJybgXKZ4_0;
	wire w_dff_A_8JSSzpdP3_0;
	wire w_dff_A_NqzCJA5O3_0;
	wire w_dff_A_K4j0spcf0_0;
	wire w_dff_A_GcND7V5D3_0;
	wire w_dff_A_JgKoGoOG6_0;
	wire w_dff_A_0OuHfazO0_0;
	wire w_dff_A_7qxCi5Hh4_0;
	wire w_dff_A_9g95h1Z50_0;
	wire w_dff_A_Pop8U8747_0;
	wire w_dff_A_HT2ozZiF6_0;
	wire w_dff_A_6KcRPZEY1_1;
	wire w_dff_A_VL4u1syn8_0;
	wire w_dff_A_qq8TKOja5_0;
	wire w_dff_A_ovPhs7Em2_0;
	wire w_dff_A_TZKGaMGi8_0;
	wire w_dff_A_XuaPGdcM1_0;
	wire w_dff_A_8HK7cpkl2_1;
	wire w_dff_A_XHwCdkcM9_0;
	wire w_dff_A_RMCiEWdP1_0;
	wire w_dff_A_ndgumlmq8_0;
	wire w_dff_A_JKwEgMNF6_0;
	wire w_dff_A_8y39fQ1n8_0;
	wire w_dff_A_qwXK7NWB1_0;
	wire w_dff_A_N9gBLWNS1_0;
	wire w_dff_A_T9EiKK7U8_0;
	wire w_dff_A_ybOm80nJ7_1;
	wire w_dff_A_pllF5Uob6_0;
	wire w_dff_A_H5JPP1089_0;
	wire w_dff_A_g4zNuHiz0_0;
	wire w_dff_A_tNXXiEgG1_0;
	wire w_dff_A_NGxlt3pd2_0;
	wire w_dff_A_N2KlKkZ48_0;
	wire w_dff_A_YxXv40kT5_1;
	wire w_dff_A_nr5st40n4_0;
	wire w_dff_A_lEjOuwSH1_0;
	wire w_dff_A_eopy3nFu1_0;
	wire w_dff_A_2mUDQUYi4_0;
	wire w_dff_A_eJneS3RH0_0;
	wire w_dff_A_TOixvbg22_0;
	wire w_dff_A_oERts3xA4_0;
	wire w_dff_A_aSH3WLwF9_0;
	wire w_dff_A_UA3c6uSj0_0;
	wire w_dff_A_9sxuK1rx0_2;
	wire w_dff_A_8Vbysi9b2_0;
	wire w_dff_A_WpWKO3K38_0;
	wire w_dff_A_0LeTCrT14_0;
	wire w_dff_A_9ZseDTY54_2;
	wire w_dff_A_HVf0SUn03_0;
	wire w_dff_A_dizJkHxB8_0;
	wire w_dff_A_1o2NTLEO3_2;
	wire w_dff_A_wmaiJ6M16_0;
	wire w_dff_A_oJAdkQg52_0;
	wire w_dff_A_ejDAC4ma8_0;
	wire w_dff_A_UFCuDxvQ5_2;
	wire w_dff_A_nwSLAHCZ1_0;
	wire w_dff_A_UsCiql2t9_0;
	wire w_dff_A_cfobi81r2_0;
	wire w_dff_A_LJKa69Qm9_2;
	wire w_dff_A_6DDb7pdb3_0;
	wire w_dff_A_u4CHBI0j2_0;
	wire w_dff_A_jXQAFSfX9_0;
	wire w_dff_A_ur4sohGn4_0;
	wire w_dff_A_YNkz6Tgg6_2;
	wire w_dff_A_mukuAoNM5_0;
	wire w_dff_A_pycDjWzk1_0;
	wire w_dff_A_6IPccs4l1_0;
	wire w_dff_A_iVlpqlh74_2;
	wire w_dff_A_c6sjhufo6_0;
	wire w_dff_A_elfhUkaj9_0;
	wire w_dff_A_lnSRuheC9_0;
	wire w_dff_A_8lfa568n2_2;
	wire w_dff_A_L4953zrj5_0;
	wire w_dff_A_tvjJ54RO0_0;
	wire w_dff_A_p0FFlBzA3_0;
	wire w_dff_A_xSGnrJLD0_0;
	wire w_dff_A_iUpifcdH2_2;
	wire w_dff_A_lQAtOq602_0;
	wire w_dff_A_44bWtlZI3_0;
	wire w_dff_A_qSB0BDZw9_0;
	wire w_dff_A_2tJJd17T5_2;
	wire w_dff_A_lCoSCkNt9_0;
	wire w_dff_A_xk7Cz47b9_0;
	wire w_dff_A_8Et3bTWw1_2;
	wire w_dff_A_q80xYIbs9_0;
	wire w_dff_A_hEQsiTAf9_0;
	wire w_dff_A_W8e3w3NF5_2;
	wire w_dff_A_iFsWFNfO5_0;
	wire w_dff_A_JhrkJhl39_2;
	wire w_dff_A_lkCp01sO9_0;
	wire w_dff_A_XYb04rwh0_0;
	wire w_dff_A_FsMUJCpF2_0;
	wire w_dff_A_EU9AjEys6_2;
	wire w_dff_A_gBeoBIe98_0;
	wire w_dff_A_Agly4Fzj9_0;
	wire w_dff_A_BvotNGEA0_2;
	wire w_dff_A_Kib1mxWx5_0;
	wire w_dff_A_Bbj03Fq73_0;
	wire w_dff_A_et8vM2y52_2;
	wire w_dff_A_5Kjw3Tkd6_0;
	wire w_dff_A_LMlsjDrx1_0;
	wire w_dff_A_EMPb80Xy4_2;
	wire w_dff_A_LzkmumMs1_0;
	wire w_dff_A_sTH0gPWI1_0;
	wire w_dff_A_cmeWtwhA1_0;
	wire w_dff_A_RaE1t2gH7_0;
	wire w_dff_A_qhYBnWPj1_0;
	wire w_dff_A_d5yH2TQb2_2;
	wire w_dff_A_0DNiYuTX8_0;
	wire w_dff_A_z297T3Oe8_0;
	wire w_dff_A_o0pkMQJ63_0;
	wire w_dff_A_KtDh1uLu6_0;
	wire w_dff_A_Z6lxaLEo3_0;
	wire w_dff_A_uayLeJHg8_2;
	wire w_dff_A_Y9j4iuZu8_2;
	jnot g0000(.din(w_G545_0[2]),.dout(w_dff_A_VHpW1ILW7_1),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(w_G366_0[1]),.dout(w_dff_A_63AobLUF2_1),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(w_dff_A_FJrUYRUW2_1),.clk(gclk));
	jnot g0005(.din(w_G338_0[1]),.dout(w_dff_A_FpfbrbRf3_1),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(w_dff_A_5cfRan3F4_2),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(w_dff_A_5t6DzlqV5_1),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(w_dff_A_WU84By202_1),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(w_dff_A_00yBnyGB8_1),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(w_dff_A_9O4gAV2i7_1),.clk(gclk));
	jand g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(w_dff_A_wElPQzTe5_2),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_xJVd7vh19_1),.dout(w_dff_A_5ftdZgkS7_2),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jor g0016(.dina(w_dff_B_NeekBaFp4_0),.dinb(w_n316_0[1]),.dout(w_dff_A_nNW8Oyib6_2),.clk(gclk));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(w_dff_A_IZSXO4y19_1),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jor g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_),.clk(gclk));
	jor g0022(.dina(w_G809_3[1]),.dinb(w_dff_B_H5ICgJDO2_1),.dout(w_dff_A_pkH3YkUJ5_2),.clk(gclk));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jor g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330),.clk(gclk));
	jor g0030(.dina(n330),.dinb(w_dff_B_T4h4UUWo7_1),.dout(w_dff_A_ggxnG5mk7_2),.clk(gclk));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jor g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336),.clk(gclk));
	jor g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(w_dff_A_9Fp90GiW7_2),.clk(gclk));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jor g0038(.dina(w_G809_2[1]),.dinb(w_dff_B_FiSJvVee4_1),.dout(w_dff_A_7aIGYmBt8_2),.clk(gclk));
	jand g0039(.dina(w_n326_1[2]),.dinb(w_dff_B_AUPL4UiY9_1),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jor g0041(.dina(w_dff_B_dFPnBT7I9_0),.dinb(w_G809_2[0]),.dout(n342),.clk(gclk));
	jor g0042(.dina(n342),.dinb(w_dff_B_V1WkeonP1_1),.dout(n343),.clk(gclk));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(w_dff_A_oXh5hHFP5_2),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(w_dff_B_u5UjHSah1_1),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jor g0046(.dina(w_dff_B_PDYKQJxI2_0),.dinb(w_G809_1[2]),.dout(n347),.clk(gclk));
	jor g0047(.dina(n347),.dinb(w_dff_B_ELkE3jRs4_1),.dout(n348),.clk(gclk));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(w_dff_A_4VBlrx7w2_2),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(w_dff_B_9OtLNadY3_1),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jor g0051(.dina(w_dff_B_Mo4niKpk5_0),.dinb(w_G809_1[1]),.dout(n352),.clk(gclk));
	jor g0052(.dina(n352),.dinb(w_dff_B_7UYQIOoi0_1),.dout(n353),.clk(gclk));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(w_dff_A_TnyExUOt6_2),.clk(gclk));
	jand g0054(.dina(w_G2358_0[2]),.dinb(G80),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_n326_0[2]),.dinb(w_dff_B_OnyUwNWl5_1),.dout(n356),.clk(gclk));
	jor g0056(.dina(n356),.dinb(w_G809_1[0]),.dout(n357),.clk(gclk));
	jor g0057(.dina(n357),.dinb(w_dff_B_kBiuCscR6_1),.dout(n358),.clk(gclk));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(w_dff_A_jviPCy004_2),.clk(gclk));
	jand g0059(.dina(w_G3552_0[1]),.dinb(w_G514_2[1]),.dout(n360),.clk(gclk));
	jnot g0060(.din(w_G514_2[0]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G3546_5[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(n362),.dinb(w_n361_0[1]),.dout(n363),.clk(gclk));
	jor g0063(.dina(n363),.dinb(w_dff_B_Sq3v5Xdh4_1),.dout(n364),.clk(gclk));
	jnot g0064(.din(n364),.dout(n365),.clk(gclk));
	jnot g0065(.din(w_G251_5[1]),.dout(n366),.clk(gclk));
	jnot g0066(.din(w_G361_1[1]),.dout(n367),.clk(gclk));
	jand g0067(.dina(n367),.dinb(w_n366_1[2]),.dout(n368),.clk(gclk));
	jnot g0068(.din(w_G248_5[2]),.dout(n369),.clk(gclk));
	jand g0069(.dina(w_G361_1[0]),.dinb(w_n369_1[2]),.dout(n370),.clk(gclk));
	jor g0070(.dina(n370),.dinb(n368),.dout(n371),.clk(gclk));
	jnot g0071(.din(w_n371_0[1]),.dout(n372),.clk(gclk));
	jand g0072(.dina(w_n372_0[1]),.dinb(w_n365_0[1]),.dout(n373),.clk(gclk));
	jnot g0073(.din(w_G351_2[2]),.dout(n374),.clk(gclk));
	jnot g0074(.din(G3550),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_n375_4[2]),.dinb(w_n374_1[1]),.dout(n376),.clk(gclk));
	jnot g0076(.din(w_G534_2[1]),.dout(n377),.clk(gclk));
	jnot g0077(.din(w_G3552_0[0]),.dout(n378),.clk(gclk));
	jand g0078(.dina(w_n378_4[2]),.dinb(w_G351_2[1]),.dout(n379),.clk(gclk));
	jor g0079(.dina(n379),.dinb(w_n377_1[1]),.dout(n380),.clk(gclk));
	jor g0080(.dina(n380),.dinb(w_dff_B_hamSiRHx7_1),.dout(n381),.clk(gclk));
	jand g0081(.dina(w_G3546_5[0]),.dinb(w_G351_2[0]),.dout(n382),.clk(gclk));
	jand g0082(.dina(w_G3548_4[2]),.dinb(w_n374_1[0]),.dout(n383),.clk(gclk));
	jor g0083(.dina(n383),.dinb(w_dff_B_oZOwAB332_1),.dout(n384),.clk(gclk));
	jor g0084(.dina(n384),.dinb(w_G534_2[0]),.dout(n385),.clk(gclk));
	jand g0085(.dina(n385),.dinb(n381),.dout(n386),.clk(gclk));
	jnot g0086(.din(w_G341_2[2]),.dout(n387),.clk(gclk));
	jand g0087(.dina(w_n375_4[1]),.dinb(w_n387_1[1]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G523_1[2]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n378_4[1]),.dinb(w_G341_2[1]),.dout(n390),.clk(gclk));
	jor g0090(.dina(n390),.dinb(w_n389_1[1]),.dout(n391),.clk(gclk));
	jor g0091(.dina(n391),.dinb(w_dff_B_WTvEmP2Q3_1),.dout(n392),.clk(gclk));
	jand g0092(.dina(w_G3546_4[2]),.dinb(w_G341_2[0]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3548_4[1]),.dinb(w_n387_1[0]),.dout(n394),.clk(gclk));
	jor g0094(.dina(n394),.dinb(w_dff_B_90WGFX200_1),.dout(n395),.clk(gclk));
	jor g0095(.dina(n395),.dinb(w_G523_1[1]),.dout(n396),.clk(gclk));
	jand g0096(.dina(n396),.dinb(n392),.dout(n397),.clk(gclk));
	jand g0097(.dina(w_n397_0[1]),.dinb(w_n386_0[1]),.dout(n398),.clk(gclk));
	jand g0098(.dina(n398),.dinb(w_dff_B_ppgzI1QW4_1),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G316_1[1]),.dinb(w_G248_5[1]),.dout(n400),.clk(gclk));
	jnot g0100(.din(w_G490_1[1]),.dout(n401),.clk(gclk));
	jnot g0101(.din(w_G316_1[0]),.dout(n402),.clk(gclk));
	jand g0102(.dina(w_n402_0[2]),.dinb(w_G251_5[0]),.dout(n403),.clk(gclk));
	jor g0103(.dina(n403),.dinb(w_n401_0[1]),.dout(n404),.clk(gclk));
	jor g0104(.dina(n404),.dinb(w_dff_B_yyfaiPDj6_1),.dout(n405),.clk(gclk));
	jnot g0105(.din(w_G254_1[1]),.dout(n406),.clk(gclk));
	jand g0106(.dina(w_n402_0[1]),.dinb(w_n406_5[1]),.dout(n407),.clk(gclk));
	jnot g0107(.din(w_G242_1[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_G316_0[2]),.dinb(w_n408_5[2]),.dout(n409),.clk(gclk));
	jor g0109(.dina(n409),.dinb(n407),.dout(n410),.clk(gclk));
	jor g0110(.dina(n410),.dinb(w_G490_1[0]),.dout(n411),.clk(gclk));
	jand g0111(.dina(n411),.dinb(n405),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G308_1[2]),.dinb(w_G248_5[0]),.dout(n413),.clk(gclk));
	jnot g0113(.din(w_G479_0[2]),.dout(n414),.clk(gclk));
	jnot g0114(.din(w_G308_1[1]),.dout(n415),.clk(gclk));
	jand g0115(.dina(w_n415_0[1]),.dinb(w_G251_4[2]),.dout(n416),.clk(gclk));
	jor g0116(.dina(n416),.dinb(w_n414_0[1]),.dout(n417),.clk(gclk));
	jor g0117(.dina(n417),.dinb(w_dff_B_HKApNhrR4_1),.dout(n418),.clk(gclk));
	jand g0118(.dina(w_n415_0[0]),.dinb(w_n406_5[0]),.dout(n419),.clk(gclk));
	jand g0119(.dina(w_G308_1[0]),.dinb(w_n408_5[1]),.dout(n420),.clk(gclk));
	jor g0120(.dina(n420),.dinb(n419),.dout(n421),.clk(gclk));
	jor g0121(.dina(n421),.dinb(w_G479_0[1]),.dout(n422),.clk(gclk));
	jand g0122(.dina(n422),.dinb(n418),.dout(n423),.clk(gclk));
	jand g0123(.dina(w_n423_0[2]),.dinb(w_n412_0[2]),.dout(n424),.clk(gclk));
	jnot g0124(.din(w_G293_0[2]),.dout(n425),.clk(gclk));
	jand g0125(.dina(w_n425_0[2]),.dinb(w_n406_4[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_G293_0[1]),.dinb(w_n408_5[0]),.dout(n427),.clk(gclk));
	jor g0127(.dina(n427),.dinb(n426),.dout(n428),.clk(gclk));
	jnot g0128(.din(w_G302_0[2]),.dout(n429),.clk(gclk));
	jand g0129(.dina(w_n429_0[1]),.dinb(w_n366_1[1]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G302_0[1]),.dinb(w_n369_1[1]),.dout(n431),.clk(gclk));
	jor g0131(.dina(n431),.dinb(n430),.dout(n432),.clk(gclk));
	jnot g0132(.din(n432),.dout(n433),.clk(gclk));
	jand g0133(.dina(w_n433_0[2]),.dinb(w_n428_1[1]),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G324_1[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n375_4[0]),.dinb(w_n435_2[1]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G503_2[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n378_4[0]),.dinb(w_G324_1[1]),.dout(n438),.clk(gclk));
	jor g0138(.dina(n438),.dinb(w_n437_0[1]),.dout(n439),.clk(gclk));
	jor g0139(.dina(n439),.dinb(w_dff_B_8P1YGzgQ2_1),.dout(n440),.clk(gclk));
	jand g0140(.dina(w_G3546_4[1]),.dinb(w_G324_1[0]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3548_4[0]),.dinb(w_n435_2[0]),.dout(n442),.clk(gclk));
	jor g0142(.dina(n442),.dinb(w_dff_B_vrHzVBPs5_1),.dout(n443),.clk(gclk));
	jor g0143(.dina(n443),.dinb(w_G503_2[0]),.dout(n444),.clk(gclk));
	jand g0144(.dina(n444),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(n434),.dout(n446),.clk(gclk));
	jand g0146(.dina(n446),.dinb(n424),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(n399),.dout(w_dff_A_FCzrs7lI1_2),.clk(gclk));
	jnot g0148(.din(w_G210_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n375_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G457_1[2]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n378_3[2]),.dinb(w_G210_2[0]),.dout(n452),.clk(gclk));
	jor g0152(.dina(n452),.dinb(w_n451_0[2]),.dout(n453),.clk(gclk));
	jor g0153(.dina(n453),.dinb(w_dff_B_cRRncVaF6_1),.dout(n454),.clk(gclk));
	jand g0154(.dina(w_G3546_4[0]),.dinb(w_G210_1[2]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n456),.clk(gclk));
	jor g0156(.dina(n456),.dinb(w_dff_B_2TSL03jK6_1),.dout(n457),.clk(gclk));
	jor g0157(.dina(n457),.dinb(w_G457_1[1]),.dout(n458),.clk(gclk));
	jand g0158(.dina(n458),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n375_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n378_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jor g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464),.clk(gclk));
	jor g0164(.dina(n464),.dinb(w_dff_B_VkR0RJnO3_1),.dout(n465),.clk(gclk));
	jand g0165(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n467),.clk(gclk));
	jor g0167(.dina(n467),.dinb(w_dff_B_AKBIMfoM4_1),.dout(n468),.clk(gclk));
	jor g0168(.dina(n468),.dinb(w_G435_1[1]),.dout(n469),.clk(gclk));
	jand g0169(.dina(n469),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G273_2[1]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n375_3[0]),.dinb(w_n471_1[2]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G411_2[1]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n378_3[0]),.dinb(w_G273_2[0]),.dout(n474),.clk(gclk));
	jor g0174(.dina(n474),.dinb(w_n473_1[1]),.dout(n475),.clk(gclk));
	jor g0175(.dina(n475),.dinb(w_dff_B_z12meKbH6_1),.dout(n476),.clk(gclk));
	jand g0176(.dina(w_G3546_3[1]),.dinb(w_G273_1[2]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3548_3[0]),.dinb(w_n471_1[1]),.dout(n478),.clk(gclk));
	jor g0178(.dina(n478),.dinb(w_dff_B_RLUsb3Cv4_1),.dout(n479),.clk(gclk));
	jor g0179(.dina(n479),.dinb(w_G411_2[0]),.dout(n480),.clk(gclk));
	jand g0180(.dina(n480),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jnot g0182(.din(w_G265_1[2]),.dout(n483),.clk(gclk));
	jand g0183(.dina(w_n375_2[2]),.dinb(w_n483_2[1]),.dout(n484),.clk(gclk));
	jnot g0184(.din(w_G400_1[2]),.dout(n485),.clk(gclk));
	jand g0185(.dina(w_n378_2[2]),.dinb(w_G265_1[1]),.dout(n486),.clk(gclk));
	jor g0186(.dina(n486),.dinb(w_n485_1[1]),.dout(n487),.clk(gclk));
	jor g0187(.dina(n487),.dinb(w_dff_B_ybO4WRJc4_1),.dout(n488),.clk(gclk));
	jand g0188(.dina(w_G3546_3[0]),.dinb(w_G265_1[0]),.dout(n489),.clk(gclk));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n483_2[0]),.dout(n490),.clk(gclk));
	jor g0190(.dina(n490),.dinb(w_dff_B_ugITFTmU9_1),.dout(n491),.clk(gclk));
	jor g0191(.dina(n491),.dinb(w_G400_1[1]),.dout(n492),.clk(gclk));
	jand g0192(.dina(n492),.dinb(n488),.dout(n493),.clk(gclk));
	jnot g0193(.din(w_G226_2[1]),.dout(n494),.clk(gclk));
	jand g0194(.dina(w_n375_2[1]),.dinb(w_n494_1[2]),.dout(n495),.clk(gclk));
	jnot g0195(.din(w_G422_1[1]),.dout(n496),.clk(gclk));
	jand g0196(.dina(w_n378_2[1]),.dinb(w_G226_2[0]),.dout(n497),.clk(gclk));
	jor g0197(.dina(n497),.dinb(w_n496_1[1]),.dout(n498),.clk(gclk));
	jor g0198(.dina(n498),.dinb(w_dff_B_GWbKGlHL4_1),.dout(n499),.clk(gclk));
	jand g0199(.dina(w_G3546_2[2]),.dinb(w_G226_1[2]),.dout(n500),.clk(gclk));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n494_1[1]),.dout(n501),.clk(gclk));
	jor g0201(.dina(n501),.dinb(w_dff_B_ZXo0Ajip9_1),.dout(n502),.clk(gclk));
	jor g0202(.dina(n502),.dinb(w_G422_1[0]),.dout(n503),.clk(gclk));
	jand g0203(.dina(n503),.dinb(n499),.dout(n504),.clk(gclk));
	jand g0204(.dina(w_n504_0[1]),.dinb(w_n493_0[1]),.dout(n505),.clk(gclk));
	jand g0205(.dina(n505),.dinb(n482),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[1]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n375_2[0]),.dinb(w_n507_1[2]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n378_2[0]),.dinb(w_G218_2[0]),.dout(n510),.clk(gclk));
	jor g0210(.dina(n510),.dinb(w_n509_0[2]),.dout(n511),.clk(gclk));
	jor g0211(.dina(n511),.dinb(w_dff_B_yOGDY6he7_1),.dout(n512),.clk(gclk));
	jand g0212(.dina(w_G3546_2[1]),.dinb(w_G218_1[2]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3548_2[0]),.dinb(w_n507_1[1]),.dout(n514),.clk(gclk));
	jor g0214(.dina(n514),.dinb(w_dff_B_0c6LfmK61_1),.dout(n515),.clk(gclk));
	jor g0215(.dina(n515),.dinb(w_G468_1[1]),.dout(n516),.clk(gclk));
	jand g0216(.dina(n516),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G257_2[1]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_n375_1[2]),.dinb(w_n518_1[2]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G389_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_n378_1[2]),.dinb(w_G257_2[0]),.dout(n521),.clk(gclk));
	jor g0221(.dina(n521),.dinb(w_n520_0[2]),.dout(n522),.clk(gclk));
	jor g0222(.dina(n522),.dinb(w_dff_B_kZQ8zMyd6_1),.dout(n523),.clk(gclk));
	jand g0223(.dina(w_G3546_2[0]),.dinb(w_G257_1[2]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_G3548_1[2]),.dinb(w_n518_1[1]),.dout(n525),.clk(gclk));
	jor g0225(.dina(n525),.dinb(w_dff_B_Ib7fXhQc1_1),.dout(n526),.clk(gclk));
	jor g0226(.dina(n526),.dinb(w_G389_1[1]),.dout(n527),.clk(gclk));
	jand g0227(.dina(n527),.dinb(n523),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[1]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G281_2[1]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n375_1[1]),.dinb(w_n530_1[2]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G374_1[2]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n378_1[1]),.dinb(w_G281_2[0]),.dout(n533),.clk(gclk));
	jor g0233(.dina(n533),.dinb(w_n532_1[1]),.dout(n534),.clk(gclk));
	jor g0234(.dina(n534),.dinb(w_dff_B_3XLwB3kW2_1),.dout(n535),.clk(gclk));
	jand g0235(.dina(w_G3546_1[2]),.dinb(w_G281_1[2]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3548_1[1]),.dinb(w_n530_1[1]),.dout(n537),.clk(gclk));
	jor g0237(.dina(n537),.dinb(w_dff_B_u9pdidx38_1),.dout(n538),.clk(gclk));
	jor g0238(.dina(n538),.dinb(w_G374_1[1]),.dout(n539),.clk(gclk));
	jand g0239(.dina(n539),.dinb(n535),.dout(n540),.clk(gclk));
	jand g0240(.dina(w_G248_4[2]),.dinb(w_G206_1[2]),.dout(n541),.clk(gclk));
	jnot g0241(.din(w_G446_1[2]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G206_1[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_G251_4[1]),.dinb(w_n543_0[1]),.dout(n544),.clk(gclk));
	jor g0244(.dina(n544),.dinb(w_dff_B_VYw4pF030_1),.dout(n545),.clk(gclk));
	jor g0245(.dina(n545),.dinb(w_dff_B_Iy94drE61_1),.dout(n546),.clk(gclk));
	jand g0246(.dina(w_n406_4[1]),.dinb(w_n543_0[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_n408_4[2]),.dinb(w_G206_1[0]),.dout(n548),.clk(gclk));
	jor g0248(.dina(n548),.dinb(n547),.dout(n549),.clk(gclk));
	jor g0249(.dina(n549),.dinb(w_G446_1[1]),.dout(n550),.clk(gclk));
	jand g0250(.dina(n550),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[2]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(n506),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_n459_0[1]),.dout(w_dff_A_w6ptbcNI1_2),.clk(gclk));
	jnot g0255(.din(w_G335_0[2]),.dout(n556),.clk(gclk));
	jand g0256(.dina(w_n556_8[1]),.dinb(w_n530_1[0]),.dout(n557),.clk(gclk));
	jnot g0257(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jor g0258(.dina(w_n556_8[0]),.dinb(w_dff_B_dcyVP1xp6_1),.dout(n559),.clk(gclk));
	jand g0259(.dina(w_n559_0[1]),.dinb(n558),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_0[2]),.dinb(w_G374_1[0]),.dout(n561),.clk(gclk));
	jand g0261(.dina(w_n556_7[2]),.dinb(w_n471_1[0]),.dout(n562),.clk(gclk));
	jnot g0262(.din(w_n562_0[1]),.dout(n563),.clk(gclk));
	jor g0263(.dina(w_n556_7[1]),.dinb(w_dff_B_hQ7pqEYK6_1),.dout(n564),.clk(gclk));
	jand g0264(.dina(w_n564_0[1]),.dinb(n563),.dout(n565),.clk(gclk));
	jxor g0265(.dina(w_n565_0[2]),.dinb(w_G411_1[2]),.dout(n566),.clk(gclk));
	jand g0266(.dina(w_n566_0[2]),.dinb(w_n561_1[1]),.dout(n567),.clk(gclk));
	jnot g0267(.din(w_n567_0[2]),.dout(n568),.clk(gclk));
	jand g0268(.dina(w_n556_7[0]),.dinb(w_n483_1[2]),.dout(n569),.clk(gclk));
	jnot g0269(.din(w_n569_0[1]),.dout(n570),.clk(gclk));
	jor g0270(.dina(w_n556_6[2]),.dinb(w_dff_B_WxmNg9VF5_1),.dout(n571),.clk(gclk));
	jand g0271(.dina(w_n571_0[1]),.dinb(n570),.dout(n572),.clk(gclk));
	jxor g0272(.dina(w_n572_0[2]),.dinb(w_G400_1[0]),.dout(n573),.clk(gclk));
	jnot g0273(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jand g0274(.dina(w_n556_6[1]),.dinb(w_n518_1[0]),.dout(n575),.clk(gclk));
	jnot g0275(.din(n575),.dout(n576),.clk(gclk));
	jor g0276(.dina(w_n556_6[0]),.dinb(w_dff_B_rh2BxCzh4_1),.dout(n577),.clk(gclk));
	jand g0277(.dina(w_dff_B_36jfe22f8_0),.dinb(n576),.dout(n578),.clk(gclk));
	jxor g0278(.dina(w_n578_1[1]),.dinb(w_n520_0[1]),.dout(n579),.clk(gclk));
	jor g0279(.dina(w_n579_1[1]),.dinb(w_n574_0[2]),.dout(n580),.clk(gclk));
	jor g0280(.dina(n580),.dinb(n568),.dout(n581),.clk(gclk));
	jnot g0281(.din(w_n581_0[1]),.dout(n582),.clk(gclk));
	jand g0282(.dina(w_n556_5[2]),.dinb(w_n460_1[0]),.dout(n583),.clk(gclk));
	jnot g0283(.din(n583),.dout(n584),.clk(gclk));
	jor g0284(.dina(w_n556_5[1]),.dinb(w_dff_B_LGHcPilM5_1),.dout(n585),.clk(gclk));
	jand g0285(.dina(w_dff_B_yCM6XrYW8_0),.dinb(n584),.dout(n586),.clk(gclk));
	jxor g0286(.dina(w_n586_1[1]),.dinb(w_G435_1[0]),.dout(n587),.clk(gclk));
	jand g0287(.dina(w_n587_0[1]),.dinb(n582),.dout(n588),.clk(gclk));
	jor g0288(.dina(w_G335_0[1]),.dinb(w_G206_0[2]),.dout(n589),.clk(gclk));
	jor g0289(.dina(w_n556_5[0]),.dinb(w_dff_B_O0nRUcvV3_1),.dout(n590),.clk(gclk));
	jand g0290(.dina(n590),.dinb(w_dff_B_qtKr0fpF5_1),.dout(n591),.clk(gclk));
	jxor g0291(.dina(w_n591_1[1]),.dinb(w_G446_1[0]),.dout(n592),.clk(gclk));
	jand g0292(.dina(w_n556_4[2]),.dinb(w_n494_1[0]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jor g0294(.dina(w_n556_4[1]),.dinb(w_dff_B_8f4RVvMu5_1),.dout(n595),.clk(gclk));
	jand g0295(.dina(w_dff_B_Yd1FmHXW5_0),.dinb(n594),.dout(n596),.clk(gclk));
	jxor g0296(.dina(w_n596_1[1]),.dinb(w_n496_1[0]),.dout(n597),.clk(gclk));
	jand g0297(.dina(w_n556_4[0]),.dinb(w_n507_1[0]),.dout(n598),.clk(gclk));
	jnot g0298(.din(n598),.dout(n599),.clk(gclk));
	jor g0299(.dina(w_n556_3[2]),.dinb(w_dff_B_y63hCaOL7_1),.dout(n600),.clk(gclk));
	jand g0300(.dina(w_dff_B_G1yOpguQ2_0),.dinb(n599),.dout(n601),.clk(gclk));
	jxor g0301(.dina(w_n601_1[1]),.dinb(w_n509_0[1]),.dout(n602),.clk(gclk));
	jor g0302(.dina(w_n602_0[2]),.dinb(w_n597_0[2]),.dout(n603),.clk(gclk));
	jand g0303(.dina(w_n556_3[1]),.dinb(w_n449_1[0]),.dout(n604),.clk(gclk));
	jnot g0304(.din(n604),.dout(n605),.clk(gclk));
	jor g0305(.dina(w_n556_3[0]),.dinb(w_dff_B_vbotFnb24_1),.dout(n606),.clk(gclk));
	jand g0306(.dina(w_dff_B_EXzRqPhv9_0),.dinb(n605),.dout(n607),.clk(gclk));
	jxor g0307(.dina(w_n607_1[1]),.dinb(w_n451_0[1]),.dout(n608),.clk(gclk));
	jor g0308(.dina(w_n608_0[2]),.dinb(w_n603_0[1]),.dout(n609),.clk(gclk));
	jnot g0309(.din(w_n609_0[2]),.dout(n610),.clk(gclk));
	jand g0310(.dina(n610),.dinb(w_n592_0[2]),.dout(n611),.clk(gclk));
	jand g0311(.dina(w_n611_0[2]),.dinb(w_n588_1[1]),.dout(w_dff_A_hjs3pf4K4_2),.clk(gclk));
	jnot g0312(.din(w_G332_3[2]),.dout(n613),.clk(gclk));
	jand g0313(.dina(w_n613_5[2]),.dinb(w_n435_1[2]),.dout(n614),.clk(gclk));
	jnot g0314(.din(n614),.dout(n615),.clk(gclk));
	jor g0315(.dina(w_n613_5[1]),.dinb(w_G331_0[1]),.dout(n616),.clk(gclk));
	jand g0316(.dina(w_dff_B_57G6NsdX4_0),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_G503_1[2]),.dout(n618),.clk(gclk));
	jor g0318(.dina(w_G338_0[0]),.dinb(w_n613_5[0]),.dout(n619),.clk(gclk));
	jxor g0319(.dina(w_n619_1[2]),.dinb(w_G514_1[2]),.dout(n620),.clk(gclk));
	jor g0320(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n621),.clk(gclk));
	jor g0321(.dina(w_G348_0[0]),.dinb(w_n613_4[2]),.dout(n622),.clk(gclk));
	jand g0322(.dina(n622),.dinb(w_n621_0[1]),.dout(n623),.clk(gclk));
	jxor g0323(.dina(w_n623_0[1]),.dinb(w_G523_1[0]),.dout(n624),.clk(gclk));
	jor g0324(.dina(w_G351_1[2]),.dinb(w_G332_3[0]),.dout(n625),.clk(gclk));
	jor g0325(.dina(w_G358_0[0]),.dinb(w_n613_4[1]),.dout(n626),.clk(gclk));
	jand g0326(.dina(n626),.dinb(w_n625_0[1]),.dout(n627),.clk(gclk));
	jor g0327(.dina(w_n627_1[1]),.dinb(w_G534_1[2]),.dout(n628),.clk(gclk));
	jnot g0328(.din(w_n625_0[0]),.dout(n629),.clk(gclk));
	jand g0329(.dina(w_G612_0),.dinb(w_G332_2[2]),.dout(n630),.clk(gclk));
	jor g0330(.dina(n630),.dinb(n629),.dout(n631),.clk(gclk));
	jor g0331(.dina(w_n631_0[1]),.dinb(w_n377_1[0]),.dout(n632),.clk(gclk));
	jor g0332(.dina(w_G361_0[2]),.dinb(w_G332_2[1]),.dout(n633),.clk(gclk));
	jor g0333(.dina(w_G366_0[0]),.dinb(w_n613_4[0]),.dout(n634),.clk(gclk));
	jand g0334(.dina(n634),.dinb(w_dff_B_Ye6HFRXg6_1),.dout(n635),.clk(gclk));
	jnot g0335(.din(w_n635_1[1]),.dout(n636),.clk(gclk));
	jand g0336(.dina(w_n636_0[2]),.dinb(w_n632_0[1]),.dout(n637),.clk(gclk));
	jand g0337(.dina(w_n637_0[2]),.dinb(w_n628_0[2]),.dout(n638),.clk(gclk));
	jand g0338(.dina(w_n638_0[1]),.dinb(w_n624_0[2]),.dout(n639),.clk(gclk));
	jand g0339(.dina(w_n639_0[2]),.dinb(w_n620_1[1]),.dout(n640),.clk(gclk));
	jand g0340(.dina(w_n640_0[1]),.dinb(w_n618_0[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n613_3[2]),.dinb(w_n425_0[1]),.dout(n642),.clk(gclk));
	jand g0342(.dina(w_G332_2[0]),.dinb(w_G593_0),.dout(n643),.clk(gclk));
	jor g0343(.dina(n643),.dinb(n642),.dout(n644),.clk(gclk));
	jand g0344(.dina(w_n613_3[1]),.dinb(w_n429_0[0]),.dout(n645),.clk(gclk));
	jnot g0345(.din(n645),.dout(n646),.clk(gclk));
	jor g0346(.dina(w_n613_3[0]),.dinb(w_dff_B_G0FqcR0X5_1),.dout(n647),.clk(gclk));
	jand g0347(.dina(w_dff_B_J7QSLHkv8_0),.dinb(n646),.dout(n648),.clk(gclk));
	jnot g0348(.din(w_n648_1[1]),.dout(n649),.clk(gclk));
	jand g0349(.dina(w_n649_0[1]),.dinb(w_n644_0[2]),.dout(n650),.clk(gclk));
	jor g0350(.dina(w_G332_1[2]),.dinb(w_G308_0[2]),.dout(n651),.clk(gclk));
	jor g0351(.dina(w_n613_2[2]),.dinb(w_dff_B_IrD5C1yu8_1),.dout(n652),.clk(gclk));
	jand g0352(.dina(n652),.dinb(w_dff_B_xOOQgFa32_1),.dout(n653),.clk(gclk));
	jxor g0353(.dina(w_n653_0[2]),.dinb(w_G479_0[0]),.dout(n654),.clk(gclk));
	jand g0354(.dina(w_n613_2[1]),.dinb(w_n402_0[0]),.dout(n655),.clk(gclk));
	jnot g0355(.din(n655),.dout(n656),.clk(gclk));
	jor g0356(.dina(w_n613_2[0]),.dinb(w_dff_B_tschl8w45_1),.dout(n657),.clk(gclk));
	jand g0357(.dina(w_dff_B_asLk4WND6_0),.dinb(n656),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_n658_1[1]),.dinb(w_G490_0[2]),.dout(n659),.clk(gclk));
	jand g0359(.dina(w_n659_0[1]),.dinb(w_n654_2[2]),.dout(n660),.clk(gclk));
	jand g0360(.dina(w_n660_1[1]),.dinb(w_n650_0[1]),.dout(n661),.clk(gclk));
	jand g0361(.dina(w_n661_0[1]),.dinb(w_n641_1[2]),.dout(w_dff_A_QVvvToBY8_2),.clk(gclk));
	jxor g0362(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G302_0[0]),.dinb(w_n425_0[0]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(w_dff_B_Qa0kXc944_1),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G369_0[1]),.dinb(w_G361_0[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(n666),.dinb(w_n435_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n668),.clk(gclk));
	jxor g0368(.dina(w_dff_B_lwgdiKd39_0),.dinb(n667),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n665),.dout(n670),.clk(gclk));
	jnot g0370(.din(w_n670_0[1]),.dout(w_dff_A_lYUtd87F9_1),.clk(gclk));
	jxor g0371(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n672),.clk(gclk));
	jxor g0372(.dina(w_G273_1[1]),.dinb(w_n483_1[1]),.dout(n673),.clk(gclk));
	jxor g0373(.dina(n673),.dinb(w_dff_B_HIzuN37p7_1),.dout(n674),.clk(gclk));
	jxor g0374(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n675),.clk(gclk));
	jxor g0375(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n676),.clk(gclk));
	jxor g0376(.dina(n676),.dinb(n675),.dout(n677),.clk(gclk));
	jxor g0377(.dina(w_G210_1[1]),.dinb(w_G206_0[1]),.dout(n678),.clk(gclk));
	jxor g0378(.dina(w_dff_B_kSKAt8eF0_0),.dinb(n677),.dout(n679),.clk(gclk));
	jxor g0379(.dina(n679),.dinb(n674),.dout(n680),.clk(gclk));
	jnot g0380(.din(w_n680_0[1]),.dout(w_dff_A_tW43U9KN1_1),.clk(gclk));
	jand g0381(.dina(w_n586_1[0]),.dinb(w_G435_0[2]),.dout(n682),.clk(gclk));
	jnot g0382(.din(w_n586_0[2]),.dout(n683),.clk(gclk));
	jand g0383(.dina(n683),.dinb(w_n462_0[1]),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n684_0[1]),.dout(n685),.clk(gclk));
	jand g0385(.dina(w_n578_1[0]),.dinb(w_G389_1[0]),.dout(n686),.clk(gclk));
	jor g0386(.dina(w_n578_0[2]),.dinb(w_G389_0[2]),.dout(n687),.clk(gclk));
	jnot g0387(.din(w_n571_0[0]),.dout(n688),.clk(gclk));
	jor g0388(.dina(n688),.dinb(w_n569_0[0]),.dout(n689),.clk(gclk));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n485_1[0]),.dout(n690),.clk(gclk));
	jnot g0390(.din(w_n690_0[1]),.dout(n691),.clk(gclk));
	jand g0391(.dina(w_n560_0[1]),.dinb(w_G374_0[2]),.dout(n692),.clk(gclk));
	jor g0392(.dina(w_n565_0[1]),.dinb(w_G411_1[1]),.dout(n693),.clk(gclk));
	jand g0393(.dina(n693),.dinb(w_n692_0[1]),.dout(n694),.clk(gclk));
	jand g0394(.dina(w_n565_0[0]),.dinb(w_G411_1[0]),.dout(n695),.clk(gclk));
	jand g0395(.dina(w_n572_0[1]),.dinb(w_G400_0[2]),.dout(n696),.clk(gclk));
	jor g0396(.dina(n696),.dinb(w_n695_0[2]),.dout(n697),.clk(gclk));
	jor g0397(.dina(n697),.dinb(w_n694_0[2]),.dout(n698),.clk(gclk));
	jand g0398(.dina(n698),.dinb(w_dff_B_I6rSOM260_1),.dout(n699),.clk(gclk));
	jand g0399(.dina(w_n699_0[2]),.dinb(w_n687_0[1]),.dout(n700),.clk(gclk));
	jor g0400(.dina(n700),.dinb(w_n686_0[1]),.dout(n701),.clk(gclk));
	jand g0401(.dina(w_n701_0[1]),.dinb(w_n685_0[1]),.dout(n702),.clk(gclk));
	jor g0402(.dina(n702),.dinb(w_n682_0[2]),.dout(n703),.clk(gclk));
	jand g0403(.dina(w_n703_0[2]),.dinb(w_n611_0[1]),.dout(n704),.clk(gclk));
	jand g0404(.dina(w_n591_1[0]),.dinb(w_G446_0[2]),.dout(n705),.clk(gclk));
	jor g0405(.dina(w_n591_0[2]),.dinb(w_G446_0[1]),.dout(n706),.clk(gclk));
	jand g0406(.dina(w_n607_1[0]),.dinb(w_G457_1[0]),.dout(n707),.clk(gclk));
	jor g0407(.dina(w_n607_0[2]),.dinb(w_G457_0[2]),.dout(n708),.clk(gclk));
	jand g0408(.dina(w_n601_1[0]),.dinb(w_G468_1[0]),.dout(n709),.clk(gclk));
	jand g0409(.dina(w_n596_1[0]),.dinb(w_G422_0[2]),.dout(n710),.clk(gclk));
	jor g0410(.dina(w_n601_0[2]),.dinb(w_G468_0[2]),.dout(n711),.clk(gclk));
	jand g0411(.dina(w_n711_0[1]),.dinb(w_n710_0[1]),.dout(n712),.clk(gclk));
	jor g0412(.dina(n712),.dinb(w_n709_0[1]),.dout(n713),.clk(gclk));
	jand g0413(.dina(w_n713_0[2]),.dinb(w_dff_B_3VKKs2DS2_1),.dout(n714),.clk(gclk));
	jor g0414(.dina(n714),.dinb(w_dff_B_bsMZhnDY2_1),.dout(n715),.clk(gclk));
	jand g0415(.dina(w_n715_0[2]),.dinb(w_dff_B_V8QbOeQJ2_1),.dout(n716),.clk(gclk));
	jor g0416(.dina(n716),.dinb(w_dff_B_QUdYuxkV7_1),.dout(n717),.clk(gclk));
	jor g0417(.dina(w_n717_0[1]),.dinb(w_n704_0[1]),.dout(w_dff_A_vKR5DkTS6_2),.clk(gclk));
	jand g0418(.dina(w_n617_1[0]),.dinb(w_G503_1[1]),.dout(n719),.clk(gclk));
	jor g0419(.dina(w_n617_0[2]),.dinb(w_G503_1[0]),.dout(n720),.clk(gclk));
	jor g0420(.dina(w_n619_1[1]),.dinb(w_G514_1[1]),.dout(n721),.clk(gclk));
	jand g0421(.dina(w_n619_1[0]),.dinb(w_G514_1[0]),.dout(n722),.clk(gclk));
	jnot g0422(.din(w_n621_0[0]),.dout(n723),.clk(gclk));
	jand g0423(.dina(w_G599_0),.dinb(w_G332_1[1]),.dout(n724),.clk(gclk));
	jor g0424(.dina(n724),.dinb(n723),.dout(n725),.clk(gclk));
	jand g0425(.dina(w_n725_0[2]),.dinb(w_n389_1[0]),.dout(n726),.clk(gclk));
	jnot g0426(.din(w_n726_0[1]),.dout(n727),.clk(gclk));
	jand g0427(.dina(w_n635_1[0]),.dinb(w_n628_0[1]),.dout(n728),.clk(gclk));
	jand g0428(.dina(w_n623_0[0]),.dinb(w_G523_0[2]),.dout(n729),.clk(gclk));
	jand g0429(.dina(w_n627_1[0]),.dinb(w_G534_1[1]),.dout(n730),.clk(gclk));
	jor g0430(.dina(n730),.dinb(n729),.dout(n731),.clk(gclk));
	jor g0431(.dina(n731),.dinb(w_n728_0[1]),.dout(n732),.clk(gclk));
	jand g0432(.dina(n732),.dinb(w_dff_B_h14bxRSR8_1),.dout(n733),.clk(gclk));
	jor g0433(.dina(w_n733_0[2]),.dinb(w_n722_0[1]),.dout(n734),.clk(gclk));
	jand g0434(.dina(n734),.dinb(w_n721_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[2]),.dinb(w_n720_0[1]),.dout(n736),.clk(gclk));
	jor g0436(.dina(n736),.dinb(w_n719_0[1]),.dout(n737),.clk(gclk));
	jand g0437(.dina(w_n737_1[1]),.dinb(w_n660_1[0]),.dout(n738),.clk(gclk));
	jnot g0438(.din(w_n650_0[0]),.dout(n739),.clk(gclk));
	jnot g0439(.din(w_n653_0[1]),.dout(n740),.clk(gclk));
	jor g0440(.dina(n740),.dinb(w_n414_0[0]),.dout(n741),.clk(gclk));
	jand g0441(.dina(w_n658_1[0]),.dinb(w_G490_0[1]),.dout(n742),.clk(gclk));
	jand g0442(.dina(w_n742_0[2]),.dinb(w_n654_2[1]),.dout(n743),.clk(gclk));
	jnot g0443(.din(n743),.dout(n744),.clk(gclk));
	jand g0444(.dina(n744),.dinb(w_dff_B_6s7BJUn44_1),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_n745_0[1]),.dout(n746),.clk(gclk));
	jor g0446(.dina(w_n746_0[2]),.dinb(w_dff_B_faKqSggN7_1),.dout(n747),.clk(gclk));
	jor g0447(.dina(w_n747_0[1]),.dinb(w_n738_0[1]),.dout(w_dff_A_XZnSM4Bv2_2),.clk(gclk));
	jnot g0448(.din(w_G4091_6[1]),.dout(n749),.clk(gclk));
	jand g0449(.dina(w_G4092_9[2]),.dinb(w_n749_13[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n750_8[2]),.dinb(w_dff_B_5JNCKSIB9_1),.dout(n751),.clk(gclk));
	jnot g0451(.din(n751),.dout(n752),.clk(gclk));
	jnot g0452(.din(w_G54_0[2]),.dout(n753),.clk(gclk));
	jxor g0453(.dina(w_n635_0[2]),.dinb(w_n753_1[1]),.dout(n754),.clk(gclk));
	jnot g0454(.din(n754),.dout(n755),.clk(gclk));
	jand g0455(.dina(w_n755_0[1]),.dinb(w_G4091_6[0]),.dout(n756),.clk(gclk));
	jand g0456(.dina(w_n372_0[0]),.dinb(w_n749_13[0]),.dout(n757),.clk(gclk));
	jor g0457(.dina(n757),.dinb(w_G4092_9[1]),.dout(n758),.clk(gclk));
	jor g0458(.dina(n758),.dinb(n756),.dout(n759),.clk(gclk));
	jand g0459(.dina(n759),.dinb(w_dff_B_Wr6GDBT12_1),.dout(G822_fa_),.clk(gclk));
	jand g0460(.dina(w_n750_8[1]),.dinb(w_dff_B_NJuNj2kG9_1),.dout(n761),.clk(gclk));
	jnot g0461(.din(n761),.dout(n762),.clk(gclk));
	jxor g0462(.dina(w_n627_0[2]),.dinb(w_G534_1[0]),.dout(n763),.clk(gclk));
	jnot g0463(.din(w_n763_0[2]),.dout(n764),.clk(gclk));
	jand g0464(.dina(n764),.dinb(w_n635_0[1]),.dout(n765),.clk(gclk));
	jor g0465(.dina(n765),.dinb(w_n638_0[0]),.dout(n766),.clk(gclk));
	jnot g0466(.din(n766),.dout(n767),.clk(gclk));
	jand g0467(.dina(w_n767_0[1]),.dinb(w_n753_1[0]),.dout(n768),.clk(gclk));
	jand g0468(.dina(w_n763_0[1]),.dinb(w_G54_0[1]),.dout(n769),.clk(gclk));
	jor g0469(.dina(w_dff_B_vFdVfgzK6_0),.dinb(n768),.dout(n770),.clk(gclk));
	jand g0470(.dina(n770),.dinb(w_G4091_5[2]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n386_0[0]),.dinb(w_n749_12[2]),.dout(n772),.clk(gclk));
	jor g0472(.dina(n772),.dinb(w_G4092_9[0]),.dout(n773),.clk(gclk));
	jor g0473(.dina(w_dff_B_HGmizWoM4_0),.dinb(n771),.dout(n774),.clk(gclk));
	jand g0474(.dina(n774),.dinb(w_dff_B_ZbyInzDL9_1),.dout(G838_fa_),.clk(gclk));
	jand g0475(.dina(w_n750_8[0]),.dinb(w_dff_B_uWQdhYHv7_1),.dout(n776),.clk(gclk));
	jnot g0476(.din(n776),.dout(n777),.clk(gclk));
	jxor g0477(.dina(w_n561_1[0]),.dinb(w_G4_0[2]),.dout(n778),.clk(gclk));
	jnot g0478(.din(n778),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n779_0[1]),.dinb(w_G4091_5[1]),.dout(n780),.clk(gclk));
	jand g0480(.dina(w_n540_0[0]),.dinb(w_n749_12[1]),.dout(n781),.clk(gclk));
	jor g0481(.dina(n781),.dinb(w_G4092_8[2]),.dout(n782),.clk(gclk));
	jor g0482(.dina(w_dff_B_kwHGDFZX7_0),.dinb(n780),.dout(n783),.clk(gclk));
	jand g0483(.dina(n783),.dinb(w_dff_B_0fwNjf782_1),.dout(G861_fa_),.clk(gclk));
	jand g0484(.dina(w_n641_1[1]),.dinb(w_G54_0[0]),.dout(n785),.clk(gclk));
	jor g0485(.dina(w_dff_B_m8lrl0n79_0),.dinb(w_n737_1[0]),.dout(n786),.clk(gclk));
	jand g0486(.dina(w_n786_0[2]),.dinb(w_n660_0[2]),.dout(n787),.clk(gclk));
	jor g0487(.dina(n787),.dinb(w_n746_0[1]),.dout(n788),.clk(gclk));
	jnot g0488(.din(w_n788_0[2]),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n644_0[1]),.dout(n790),.clk(gclk));
	jxor g0490(.dina(w_n648_1[0]),.dinb(w_n790_0[2]),.dout(n791),.clk(gclk));
	jnot g0491(.din(n791),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_n792_0[2]),.dinb(n789),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n788_0[1]),.dinb(w_n790_0[1]),.dout(n794),.clk(gclk));
	jor g0494(.dina(w_dff_B_7CzP2E2L3_0),.dinb(n793),.dout(n795),.clk(gclk));
	jnot g0495(.din(w_n795_1[1]),.dout(G623_fa_),.clk(gclk));
	jnot g0496(.din(w_G4088_9[2]),.dout(n797),.clk(gclk));
	jnot g0497(.din(w_G861_0),.dout(n798),.clk(gclk));
	jor g0498(.dina(w_n798_1[1]),.dinb(w_n797_9[1]),.dout(n799),.clk(gclk));
	jnot g0499(.din(w_G4087_4[2]),.dout(n800),.clk(gclk));
	jnot g0500(.din(w_G822_0),.dout(n801),.clk(gclk));
	jor g0501(.dina(w_n801_1[1]),.dinb(w_G4088_9[1]),.dout(n802),.clk(gclk));
	jand g0502(.dina(n802),.dinb(w_n800_4[1]),.dout(n803),.clk(gclk));
	jand g0503(.dina(w_dff_B_1PScmEgp4_0),.dinb(n799),.dout(n804),.clk(gclk));
	jor g0504(.dina(w_n797_9[0]),.dinb(w_G61_0[1]),.dout(n805),.clk(gclk));
	jor g0505(.dina(w_G4088_9[0]),.dinb(w_G11_0[1]),.dout(n806),.clk(gclk));
	jand g0506(.dina(n806),.dinb(w_G4087_4[1]),.dout(n807),.clk(gclk));
	jand g0507(.dina(n807),.dinb(n805),.dout(n808),.clk(gclk));
	jor g0508(.dina(w_dff_B_oplNXEDL6_0),.dinb(n804),.dout(w_dff_A_PsMfZTAJ4_2),.clk(gclk));
	jand g0509(.dina(w_n750_7[2]),.dinb(w_dff_B_9EyVRvmn8_1),.dout(n810),.clk(gclk));
	jnot g0510(.din(n810),.dout(n811),.clk(gclk));
	jnot g0511(.din(w_n721_0[0]),.dout(n812),.clk(gclk));
	jnot g0512(.din(w_n722_0[0]),.dout(n813),.clk(gclk));
	jand g0513(.dina(w_n631_0[0]),.dinb(w_n377_0[2]),.dout(n814),.clk(gclk));
	jor g0514(.dina(w_n636_0[1]),.dinb(w_n814_0[2]),.dout(n815),.clk(gclk));
	jor g0515(.dina(w_n725_0[1]),.dinb(w_n389_0[2]),.dout(n816),.clk(gclk));
	jand g0516(.dina(w_n632_0[0]),.dinb(n816),.dout(n817),.clk(gclk));
	jand g0517(.dina(n817),.dinb(n815),.dout(n818),.clk(gclk));
	jor g0518(.dina(n818),.dinb(w_n726_0[0]),.dout(n819),.clk(gclk));
	jand g0519(.dina(w_n819_0[2]),.dinb(w_dff_B_N0rTAIrb9_1),.dout(n820),.clk(gclk));
	jor g0520(.dina(n820),.dinb(w_dff_B_WzlzO9Pe6_1),.dout(n821),.clk(gclk));
	jnot g0521(.din(w_n620_1[0]),.dout(n822),.clk(gclk));
	jnot g0522(.din(w_n639_0[1]),.dout(n823),.clk(gclk));
	jor g0523(.dina(n823),.dinb(w_n753_0[2]),.dout(n824),.clk(gclk));
	jor g0524(.dina(w_n824_0[1]),.dinb(w_dff_B_qwPBKtuU9_1),.dout(n825),.clk(gclk));
	jand g0525(.dina(n825),.dinb(w_n821_0[1]),.dout(n826),.clk(gclk));
	jxor g0526(.dina(n826),.dinb(w_n618_0[1]),.dout(n827),.clk(gclk));
	jand g0527(.dina(w_n827_0[1]),.dinb(w_G4091_5[0]),.dout(n828),.clk(gclk));
	jand g0528(.dina(w_n445_0[0]),.dinb(w_n749_12[0]),.dout(n829),.clk(gclk));
	jor g0529(.dina(n829),.dinb(w_G4092_8[1]),.dout(n830),.clk(gclk));
	jor g0530(.dina(w_dff_B_hGo6aE1L4_0),.dinb(n828),.dout(n831),.clk(gclk));
	jand g0531(.dina(n831),.dinb(w_dff_B_YaNA41sQ1_1),.dout(G832_fa_),.clk(gclk));
	jand g0532(.dina(w_n750_7[1]),.dinb(w_dff_B_4LVBH2It6_1),.dout(n833),.clk(gclk));
	jnot g0533(.din(n833),.dout(n834),.clk(gclk));
	jand g0534(.dina(w_n824_0[0]),.dinb(w_n819_0[1]),.dout(n835),.clk(gclk));
	jxor g0535(.dina(n835),.dinb(w_n620_0[2]),.dout(n836),.clk(gclk));
	jand g0536(.dina(w_n836_0[1]),.dinb(w_G4091_4[2]),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_n365_0[0]),.dinb(w_n749_11[2]),.dout(n838),.clk(gclk));
	jor g0538(.dina(n838),.dinb(w_G4092_8[0]),.dout(n839),.clk(gclk));
	jor g0539(.dina(w_dff_B_G225qpP34_0),.dinb(n837),.dout(n840),.clk(gclk));
	jand g0540(.dina(n840),.dinb(w_dff_B_BQ2EQVOl9_1),.dout(G834_fa_),.clk(gclk));
	jand g0541(.dina(w_n750_7[0]),.dinb(w_dff_B_7640OupI3_1),.dout(n842),.clk(gclk));
	jnot g0542(.din(n842),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n397_0[0]),.dinb(w_n749_11[1]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_n637_0[1]),.dinb(w_n753_0[1]),.dout(n845),.clk(gclk));
	jor g0545(.dina(n845),.dinb(w_n814_0[1]),.dout(n846),.clk(gclk));
	jxor g0546(.dina(n846),.dinb(w_n624_0[1]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_0[1]),.dinb(w_G4091_4[1]),.dout(n848),.clk(gclk));
	jor g0548(.dina(n848),.dinb(w_G4092_7[2]),.dout(n849),.clk(gclk));
	jor g0549(.dina(n849),.dinb(w_dff_B_sStGSEa44_1),.dout(n850),.clk(gclk));
	jand g0550(.dina(n850),.dinb(w_dff_B_Pg0Xh79Q8_1),.dout(G836_fa_),.clk(gclk));
	jnot g0551(.din(w_G4089_9[2]),.dout(n852),.clk(gclk));
	jor g0552(.dina(w_n798_1[0]),.dinb(w_n852_9[1]),.dout(n853),.clk(gclk));
	jnot g0553(.din(w_G4090_4[2]),.dout(n854),.clk(gclk));
	jor g0554(.dina(w_n801_1[0]),.dinb(w_G4089_9[1]),.dout(n855),.clk(gclk));
	jand g0555(.dina(n855),.dinb(w_n854_4[1]),.dout(n856),.clk(gclk));
	jand g0556(.dina(w_dff_B_Zj1aWoW30_0),.dinb(n853),.dout(n857),.clk(gclk));
	jor g0557(.dina(w_n852_9[0]),.dinb(w_G61_0[0]),.dout(n858),.clk(gclk));
	jor g0558(.dina(w_G4089_9[0]),.dinb(w_G11_0[0]),.dout(n859),.clk(gclk));
	jand g0559(.dina(n859),.dinb(w_G4090_4[1]),.dout(n860),.clk(gclk));
	jand g0560(.dina(n860),.dinb(n858),.dout(n861),.clk(gclk));
	jor g0561(.dina(w_dff_B_ka2cL7cq3_0),.dinb(n857),.dout(w_dff_A_uCgvuOjA0_2),.clk(gclk));
	jand g0562(.dina(w_n750_6[2]),.dinb(w_dff_B_7UNUH5rp2_1),.dout(n863),.clk(gclk));
	jnot g0563(.din(n863),.dout(n864),.clk(gclk));
	jnot g0564(.din(w_n587_0[0]),.dout(n865),.clk(gclk));
	jnot g0565(.din(w_n579_1[0]),.dout(n866),.clk(gclk));
	jand g0566(.dina(w_n567_0[1]),.dinb(w_G4_0[1]),.dout(n867),.clk(gclk));
	jand g0567(.dina(w_n867_0[1]),.dinb(w_n573_0[1]),.dout(n868),.clk(gclk));
	jand g0568(.dina(w_n868_0[1]),.dinb(w_dff_B_9UXiCv0m5_1),.dout(n869),.clk(gclk));
	jor g0569(.dina(w_dff_B_1etY6Mwd5_0),.dinb(w_n701_0[0]),.dout(n870),.clk(gclk));
	jxor g0570(.dina(w_n870_0[1]),.dinb(w_n865_0[2]),.dout(n871),.clk(gclk));
	jand g0571(.dina(w_n871_0[1]),.dinb(w_G4091_4[0]),.dout(n872),.clk(gclk));
	jand g0572(.dina(w_n470_0[0]),.dinb(w_n749_11[0]),.dout(n873),.clk(gclk));
	jor g0573(.dina(n873),.dinb(w_G4092_7[1]),.dout(n874),.clk(gclk));
	jor g0574(.dina(w_dff_B_ZIzc92Bh0_0),.dinb(n872),.dout(n875),.clk(gclk));
	jand g0575(.dina(n875),.dinb(w_dff_B_mRm8lSLm3_1),.dout(G871_fa_),.clk(gclk));
	jand g0576(.dina(w_n750_6[1]),.dinb(w_dff_B_e7Aq2xOM1_1),.dout(n877),.clk(gclk));
	jnot g0577(.din(n877),.dout(n878),.clk(gclk));
	jor g0578(.dina(w_n868_0[0]),.dinb(w_n699_0[1]),.dout(n879),.clk(gclk));
	jxor g0579(.dina(n879),.dinb(w_n579_0[2]),.dout(n880),.clk(gclk));
	jand g0580(.dina(w_n880_0[1]),.dinb(w_G4091_3[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n528_0[0]),.dinb(w_n749_10[2]),.dout(n882),.clk(gclk));
	jor g0582(.dina(n882),.dinb(w_G4092_7[0]),.dout(n883),.clk(gclk));
	jor g0583(.dina(w_dff_B_wazcHJKO4_0),.dinb(n881),.dout(n884),.clk(gclk));
	jand g0584(.dina(n884),.dinb(w_dff_B_c9O17rgw7_1),.dout(G873_fa_),.clk(gclk));
	jand g0585(.dina(w_n750_6[0]),.dinb(w_dff_B_l6Ij8nIr3_1),.dout(n886),.clk(gclk));
	jnot g0586(.din(n886),.dout(n887),.clk(gclk));
	jor g0587(.dina(w_n694_0[1]),.dinb(w_n695_0[1]),.dout(n888),.clk(gclk));
	jor g0588(.dina(n888),.dinb(w_n867_0[0]),.dout(n889),.clk(gclk));
	jxor g0589(.dina(n889),.dinb(w_n574_0[1]),.dout(n890),.clk(gclk));
	jand g0590(.dina(w_n890_0[1]),.dinb(w_G4091_3[1]),.dout(n891),.clk(gclk));
	jand g0591(.dina(w_n493_0[0]),.dinb(w_n749_10[1]),.dout(n892),.clk(gclk));
	jor g0592(.dina(n892),.dinb(w_G4092_6[2]),.dout(n893),.clk(gclk));
	jor g0593(.dina(w_dff_B_I1dON0uH7_0),.dinb(n891),.dout(n894),.clk(gclk));
	jand g0594(.dina(n894),.dinb(w_dff_B_9P4ED7zy1_1),.dout(G875_fa_),.clk(gclk));
	jand g0595(.dina(w_n750_5[2]),.dinb(w_dff_B_PS2S0xBY7_1),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jnot g0597(.din(w_n566_0[1]),.dout(n898),.clk(gclk));
	jand g0598(.dina(w_n561_0[2]),.dinb(w_G4_0[0]),.dout(n899),.clk(gclk));
	jor g0599(.dina(n899),.dinb(w_n692_0[0]),.dout(n900),.clk(gclk));
	jxor g0600(.dina(n900),.dinb(w_dff_B_eJ69Mfy49_1),.dout(n901),.clk(gclk));
	jand g0601(.dina(w_n901_0[1]),.dinb(w_G4091_3[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_n481_0[0]),.dinb(w_n749_10[0]),.dout(n903),.clk(gclk));
	jor g0603(.dina(n903),.dinb(w_G4092_6[1]),.dout(n904),.clk(gclk));
	jor g0604(.dina(w_dff_B_S49bTiMW9_0),.dinb(n902),.dout(n905),.clk(gclk));
	jand g0605(.dina(n905),.dinb(w_dff_B_VwpLRZYF3_1),.dout(G877_fa_),.clk(gclk));
	jnot g0606(.din(w_G331_0[0]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_n619_0[2]),.dout(n908),.clk(gclk));
	jand g0608(.dina(n908),.dinb(w_dff_B_7xINs6mG3_1),.dout(n909),.clk(gclk));
	jand g0609(.dina(w_n619_0[1]),.dinb(w_n617_0[1]),.dout(n910),.clk(gclk));
	jor g0610(.dina(n910),.dinb(w_dff_B_UpMQVbjd6_1),.dout(n911),.clk(gclk));
	jxor g0611(.dina(n911),.dinb(w_n792_0[1]),.dout(n912),.clk(gclk));
	jor g0612(.dina(w_G369_0[0]),.dinb(w_G332_1[0]),.dout(n913),.clk(gclk));
	jor g0613(.dina(w_dff_B_Y91lCFsy5_0),.dinb(w_n613_1[2]),.dout(n914),.clk(gclk));
	jand g0614(.dina(n914),.dinb(w_dff_B_xLQe94xi2_1),.dout(n915),.clk(gclk));
	jxor g0615(.dina(w_dff_B_GgwDVmIk2_0),.dinb(w_n636_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n627_0[1]),.dinb(w_n725_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(w_n658_0[2]),.dinb(w_n653_0[0]),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_dff_B_ArBKaFRb0_1),.dout(n919),.clk(gclk));
	jxor g0619(.dina(n919),.dinb(w_dff_B_gv7JNX2u5_1),.dout(n920),.clk(gclk));
	jxor g0620(.dina(n920),.dinb(n912),.dout(G998_fa_),.clk(gclk));
	jnot g0621(.din(w_n564_0[0]),.dout(n922),.clk(gclk));
	jor g0622(.dina(n922),.dinb(w_n562_0[0]),.dout(n923),.clk(gclk));
	jxor g0623(.dina(w_n578_0[1]),.dinb(w_n923_0[2]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n572_0[0]),.dinb(w_n560_0[0]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jor g0626(.dina(w_G335_0[0]),.dinb(w_G289_0[0]),.dout(n927),.clk(gclk));
	jor g0627(.dina(w_n556_2[2]),.dinb(w_dff_B_KzVdmX5f1_1),.dout(n928),.clk(gclk));
	jand g0628(.dina(n928),.dinb(w_dff_B_1GSiAlF65_1),.dout(n929),.clk(gclk));
	jxor g0629(.dina(n929),.dinb(w_n591_0[1]),.dout(n930),.clk(gclk));
	jxor g0630(.dina(w_n596_0[2]),.dinb(w_n586_0[1]),.dout(n931),.clk(gclk));
	jxor g0631(.dina(w_n607_0[1]),.dinb(w_n601_0[1]),.dout(n932),.clk(gclk));
	jxor g0632(.dina(n932),.dinb(n931),.dout(n933),.clk(gclk));
	jxor g0633(.dina(n933),.dinb(w_dff_B_WMbiIHUO3_1),.dout(n934),.clk(gclk));
	jxor g0634(.dina(n934),.dinb(w_dff_B_Lkz0kzL29_1),.dout(n935),.clk(gclk));
	jnot g0635(.din(w_n935_0[1]),.dout(w_dff_A_DX0Mtc6R2_1),.clk(gclk));
	jnot g0636(.din(w_n592_0[1]),.dout(n937),.clk(gclk));
	jnot g0637(.din(w_n715_0[1]),.dout(n938),.clk(gclk));
	jor g0638(.dina(w_n870_0[0]),.dinb(w_n682_0[1]),.dout(n939),.clk(gclk));
	jand g0639(.dina(n939),.dinb(w_n685_0[0]),.dout(n940),.clk(gclk));
	jnot g0640(.din(w_n940_1[1]),.dout(n941),.clk(gclk));
	jor g0641(.dina(n941),.dinb(w_n609_0[1]),.dout(n942),.clk(gclk));
	jand g0642(.dina(n942),.dinb(w_n938_0[2]),.dout(n943),.clk(gclk));
	jxor g0643(.dina(n943),.dinb(w_dff_B_ulWuoMYT0_1),.dout(n944),.clk(gclk));
	jnot g0644(.din(w_n944_0[1]),.dout(n945),.clk(gclk));
	jnot g0645(.din(w_n603_0[0]),.dout(n946),.clk(gclk));
	jand g0646(.dina(w_n940_1[0]),.dinb(w_dff_B_YgrLRGQT5_1),.dout(n947),.clk(gclk));
	jor g0647(.dina(n947),.dinb(w_n713_0[1]),.dout(n948),.clk(gclk));
	jxor g0648(.dina(n948),.dinb(w_n608_0[1]),.dout(n949),.clk(gclk));
	jand g0649(.dina(w_n949_0[1]),.dinb(n945),.dout(n950),.clk(gclk));
	jnot g0650(.din(w_n602_0[1]),.dout(n951),.clk(gclk));
	jnot g0651(.din(w_n596_0[1]),.dout(n952),.clk(gclk));
	jand g0652(.dina(n952),.dinb(w_n496_0[2]),.dout(n953),.clk(gclk));
	jnot g0653(.din(w_n953_0[1]),.dout(n954),.clk(gclk));
	jor g0654(.dina(w_n940_0[2]),.dinb(w_n710_0[0]),.dout(n955),.clk(gclk));
	jand g0655(.dina(n955),.dinb(w_n954_0[2]),.dout(n956),.clk(gclk));
	jxor g0656(.dina(n956),.dinb(w_dff_B_6atzRXp50_1),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n957_0[1]),.dout(n958),.clk(gclk));
	jand g0658(.dina(w_n890_0[0]),.dinb(w_n779_0[0]),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(w_n901_0[0]),.dout(n960),.clk(gclk));
	jand g0660(.dina(w_dff_B_iqLddp8R8_0),.dinb(w_n871_0[0]),.dout(n961),.clk(gclk));
	jnot g0661(.din(w_n597_0[1]),.dout(n962),.clk(gclk));
	jxor g0662(.dina(w_n940_0[1]),.dinb(w_n962_0[1]),.dout(n963),.clk(gclk));
	jnot g0663(.din(n963),.dout(n964),.clk(gclk));
	jand g0664(.dina(w_n964_0[1]),.dinb(w_n880_0[0]),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(w_dff_B_nTaXBT9q0_1),.dout(n966),.clk(gclk));
	jand g0666(.dina(n966),.dinb(n958),.dout(n967),.clk(gclk));
	jand g0667(.dina(w_dff_B_ifnOJc1U1_0),.dinb(n950),.dout(w_dff_A_WTTfnauU2_2),.clk(gclk));
	jxor g0668(.dina(w_n788_0[0]),.dinb(w_n649_0[0]),.dout(n969),.clk(gclk));
	jnot g0669(.din(w_n969_0[1]),.dout(n970),.clk(gclk));
	jand g0670(.dina(n970),.dinb(w_n755_0[0]),.dout(n971),.clk(gclk));
	jand g0671(.dina(w_n836_0[0]),.dinb(w_G623_0),.dout(n972),.clk(gclk));
	jand g0672(.dina(n972),.dinb(w_dff_B_CpVbdhlH2_1),.dout(n973),.clk(gclk));
	jand g0673(.dina(w_n827_0[0]),.dinb(w_n763_0[0]),.dout(n974),.clk(gclk));
	jand g0674(.dina(n974),.dinb(w_n847_0[0]),.dout(n975),.clk(gclk));
	jnot g0675(.din(w_n658_0[1]),.dout(n976),.clk(gclk));
	jand g0676(.dina(n976),.dinb(w_n401_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(w_n977_0[2]),.dinb(w_n654_2[0]),.dout(n978),.clk(gclk));
	jor g0678(.dina(w_n977_0[1]),.dinb(w_n654_1[2]),.dout(n979),.clk(gclk));
	jnot g0679(.din(n979),.dout(n980),.clk(gclk));
	jor g0680(.dina(w_n786_0[1]),.dinb(w_n742_0[1]),.dout(n981),.clk(gclk));
	jand g0681(.dina(w_n981_0[1]),.dinb(w_dff_B_0D9ogn6Y8_1),.dout(n982),.clk(gclk));
	jnot g0682(.din(w_n981_0[0]),.dout(n983),.clk(gclk));
	jand g0683(.dina(n983),.dinb(w_n654_1[1]),.dout(n984),.clk(gclk));
	jor g0684(.dina(n984),.dinb(w_dff_B_pyHhzsWM4_1),.dout(n985),.clk(gclk));
	jor g0685(.dina(n985),.dinb(w_dff_B_ICYdCDT54_1),.dout(n986),.clk(gclk));
	jnot g0686(.din(w_n986_0[1]),.dout(n987),.clk(gclk));
	jnot g0687(.din(w_n659_0[0]),.dout(n988),.clk(gclk));
	jxor g0688(.dina(w_n786_0[0]),.dinb(w_dff_B_SyvHB0u91_1),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_n989_0[1]),.dinb(n987),.dout(n990),.clk(gclk));
	jand g0690(.dina(n990),.dinb(w_dff_B_AxD9PwDr3_1),.dout(n991),.clk(gclk));
	jand g0691(.dina(n991),.dinb(n973),.dout(w_dff_A_RJ18dgvy4_2),.clk(gclk));
	jnot g0692(.din(w_G1689_5[1]),.dout(n993),.clk(gclk));
	jand g0693(.dina(w_G1690_1[1]),.dinb(w_n993_4[2]),.dout(n994),.clk(gclk));
	jand g0694(.dina(w_n994_4[1]),.dinb(w_G182_0[1]),.dout(n995),.clk(gclk));
	jand g0695(.dina(w_G1690_1[0]),.dinb(w_G1689_5[0]),.dout(n996),.clk(gclk));
	jand g0696(.dina(w_n996_4[1]),.dinb(w_G185_0[1]),.dout(n997),.clk(gclk));
	jor g0697(.dina(w_n798_0[2]),.dinb(w_n993_4[1]),.dout(n998),.clk(gclk));
	jnot g0698(.din(w_G1690_0[2]),.dout(n999),.clk(gclk));
	jor g0699(.dina(w_n801_0[2]),.dinb(w_G1689_4[2]),.dout(n1000),.clk(gclk));
	jand g0700(.dina(n1000),.dinb(w_n999_3[2]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_dff_B_gGhJvAVX2_0),.dinb(n998),.dout(n1002),.clk(gclk));
	jor g0702(.dina(n1002),.dinb(w_dff_B_zadYHcFr1_1),.dout(n1003),.clk(gclk));
	jor g0703(.dina(n1003),.dinb(w_dff_B_bIlR0n4s5_1),.dout(n1004),.clk(gclk));
	jand g0704(.dina(n1004),.dinb(w_G137_9[1]),.dout(w_dff_A_cgdxqHwN3_2),.clk(gclk));
	jor g0705(.dina(w_n801_0[1]),.dinb(w_G1691_5[1]),.dout(n1006),.clk(gclk));
	jnot g0706(.din(w_G1694_1[1]),.dout(n1007),.clk(gclk));
	jnot g0707(.din(w_G1691_5[0]),.dout(n1008),.clk(gclk));
	jor g0708(.dina(w_n798_0[1]),.dinb(w_n1008_4[2]),.dout(n1009),.clk(gclk));
	jand g0709(.dina(n1009),.dinb(w_n1007_3[2]),.dout(n1010),.clk(gclk));
	jand g0710(.dina(n1010),.dinb(w_dff_B_PSJp4qRu8_1),.dout(n1011),.clk(gclk));
	jand g0711(.dina(w_G1694_1[0]),.dinb(w_G1691_4[2]),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_4[1]),.dinb(w_G185_0[0]),.dout(n1013),.clk(gclk));
	jand g0713(.dina(w_G1694_0[2]),.dinb(w_n1008_4[1]),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_4[1]),.dinb(w_G182_0[0]),.dout(n1015),.clk(gclk));
	jor g0715(.dina(n1015),.dinb(w_dff_B_s0XwuCNn0_1),.dout(n1016),.clk(gclk));
	jor g0716(.dina(w_dff_B_Ma1gKVog9_0),.dinb(n1011),.dout(n1017),.clk(gclk));
	jand g0717(.dina(n1017),.dinb(w_G137_9[0]),.dout(w_dff_A_7W4GWUDP1_2),.clk(gclk));
	jnot g0718(.din(w_G871_0),.dout(n1019),.clk(gclk));
	jor g0719(.dina(w_n1019_1[1]),.dinb(w_n797_8[2]),.dout(n1020),.clk(gclk));
	jnot g0720(.din(w_G832_0),.dout(n1021),.clk(gclk));
	jor g0721(.dina(w_n1021_1[1]),.dinb(w_G4088_8[2]),.dout(n1022),.clk(gclk));
	jand g0722(.dina(n1022),.dinb(w_n800_4[0]),.dout(n1023),.clk(gclk));
	jand g0723(.dina(n1023),.dinb(w_dff_B_IsG2THwt3_1),.dout(n1024),.clk(gclk));
	jor g0724(.dina(w_n797_8[1]),.dinb(w_G37_0[1]),.dout(n1025),.clk(gclk));
	jor g0725(.dina(w_G4088_8[1]),.dinb(w_G43_0[1]),.dout(n1026),.clk(gclk));
	jand g0726(.dina(n1026),.dinb(w_G4087_4[0]),.dout(n1027),.clk(gclk));
	jand g0727(.dina(n1027),.dinb(n1025),.dout(n1028),.clk(gclk));
	jor g0728(.dina(w_dff_B_UIq314s07_0),.dinb(n1024),.dout(w_dff_A_GBVcLEQV9_2),.clk(gclk));
	jnot g0729(.din(w_G873_0),.dout(n1030),.clk(gclk));
	jor g0730(.dina(w_n1030_1[1]),.dinb(w_n797_8[0]),.dout(n1031),.clk(gclk));
	jnot g0731(.din(w_G834_0),.dout(n1032),.clk(gclk));
	jor g0732(.dina(w_n1032_1[1]),.dinb(w_G4088_8[0]),.dout(n1033),.clk(gclk));
	jand g0733(.dina(n1033),.dinb(w_n800_3[2]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(n1034),.dinb(w_dff_B_JNeHI5JZ0_1),.dout(n1035),.clk(gclk));
	jor g0735(.dina(w_n797_7[2]),.dinb(w_G20_0[1]),.dout(n1036),.clk(gclk));
	jor g0736(.dina(w_G4088_7[2]),.dinb(w_G76_0[1]),.dout(n1037),.clk(gclk));
	jand g0737(.dina(n1037),.dinb(w_G4087_3[2]),.dout(n1038),.clk(gclk));
	jand g0738(.dina(n1038),.dinb(n1036),.dout(n1039),.clk(gclk));
	jor g0739(.dina(w_dff_B_EmJXUkSS3_0),.dinb(n1035),.dout(w_dff_A_nBX0wvip1_2),.clk(gclk));
	jnot g0740(.din(w_G836_0),.dout(n1041),.clk(gclk));
	jor g0741(.dina(w_n1041_1[1]),.dinb(w_G4088_7[1]),.dout(n1042),.clk(gclk));
	jnot g0742(.din(w_G875_0),.dout(n1043),.clk(gclk));
	jor g0743(.dina(w_n1043_1[1]),.dinb(w_n797_7[1]),.dout(n1044),.clk(gclk));
	jand g0744(.dina(n1044),.dinb(w_n800_3[1]),.dout(n1045),.clk(gclk));
	jand g0745(.dina(n1045),.dinb(w_dff_B_wp0a28OD5_1),.dout(n1046),.clk(gclk));
	jor g0746(.dina(w_n797_7[0]),.dinb(w_G17_0[1]),.dout(n1047),.clk(gclk));
	jor g0747(.dina(w_G4088_7[0]),.dinb(w_G73_0[1]),.dout(n1048),.clk(gclk));
	jand g0748(.dina(n1048),.dinb(w_G4087_3[1]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(n1049),.dinb(n1047),.dout(n1050),.clk(gclk));
	jor g0750(.dina(w_dff_B_5cicOMT37_0),.dinb(n1046),.dout(w_dff_A_7if5Ex0z2_2),.clk(gclk));
	jnot g0751(.din(w_G877_0),.dout(n1052),.clk(gclk));
	jor g0752(.dina(w_n1052_1[1]),.dinb(w_n797_6[2]),.dout(n1053),.clk(gclk));
	jnot g0753(.din(w_G838_0),.dout(n1054),.clk(gclk));
	jor g0754(.dina(w_n1054_1[1]),.dinb(w_G4088_6[2]),.dout(n1055),.clk(gclk));
	jand g0755(.dina(n1055),.dinb(w_n800_3[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(n1056),.dinb(w_dff_B_BkBJegN79_1),.dout(n1057),.clk(gclk));
	jor g0757(.dina(w_n797_6[1]),.dinb(w_G70_0[1]),.dout(n1058),.clk(gclk));
	jor g0758(.dina(w_G4088_6[1]),.dinb(w_G67_0[1]),.dout(n1059),.clk(gclk));
	jand g0759(.dina(n1059),.dinb(w_G4087_3[0]),.dout(n1060),.clk(gclk));
	jand g0760(.dina(n1060),.dinb(n1058),.dout(n1061),.clk(gclk));
	jor g0761(.dina(w_dff_B_PrVErDRB6_0),.dinb(n1057),.dout(w_dff_A_esKhrEUJ8_2),.clk(gclk));
	jor g0762(.dina(w_G4089_8[2]),.dinb(w_G43_0[0]),.dout(n1063),.clk(gclk));
	jor g0763(.dina(w_n852_8[2]),.dinb(w_G37_0[0]),.dout(n1064),.clk(gclk));
	jand g0764(.dina(n1064),.dinb(w_G4090_4[0]),.dout(n1065),.clk(gclk));
	jand g0765(.dina(n1065),.dinb(w_dff_B_fm2x8dKD1_1),.dout(n1066),.clk(gclk));
	jor g0766(.dina(w_n1021_1[0]),.dinb(w_G4089_8[1]),.dout(n1067),.clk(gclk));
	jor g0767(.dina(w_n1019_1[0]),.dinb(w_n852_8[1]),.dout(n1068),.clk(gclk));
	jand g0768(.dina(n1068),.dinb(n1067),.dout(n1069),.clk(gclk));
	jand g0769(.dina(n1069),.dinb(w_n854_4[0]),.dout(n1070),.clk(gclk));
	jor g0770(.dina(n1070),.dinb(w_dff_B_sw0kQIIT5_1),.dout(w_dff_A_Zo2KDTfC2_2),.clk(gclk));
	jor g0771(.dina(w_G4089_8[0]),.dinb(w_G76_0[0]),.dout(n1072),.clk(gclk));
	jor g0772(.dina(w_n852_8[0]),.dinb(w_G20_0[0]),.dout(n1073),.clk(gclk));
	jand g0773(.dina(n1073),.dinb(w_G4090_3[2]),.dout(n1074),.clk(gclk));
	jand g0774(.dina(n1074),.dinb(w_dff_B_dSaYggRw8_1),.dout(n1075),.clk(gclk));
	jor g0775(.dina(w_n1032_1[0]),.dinb(w_G4089_7[2]),.dout(n1076),.clk(gclk));
	jor g0776(.dina(w_n1030_1[0]),.dinb(w_n852_7[2]),.dout(n1077),.clk(gclk));
	jand g0777(.dina(w_dff_B_3RUDA86W1_0),.dinb(n1076),.dout(n1078),.clk(gclk));
	jand g0778(.dina(n1078),.dinb(w_n854_3[2]),.dout(n1079),.clk(gclk));
	jor g0779(.dina(n1079),.dinb(w_dff_B_R3xuKQ1A8_1),.dout(w_dff_A_AdHQiQye7_2),.clk(gclk));
	jor g0780(.dina(w_G4089_7[1]),.dinb(w_G73_0[0]),.dout(n1081),.clk(gclk));
	jor g0781(.dina(w_n852_7[1]),.dinb(w_G17_0[0]),.dout(n1082),.clk(gclk));
	jand g0782(.dina(n1082),.dinb(w_G4090_3[1]),.dout(n1083),.clk(gclk));
	jand g0783(.dina(n1083),.dinb(w_dff_B_wsR42LE81_1),.dout(n1084),.clk(gclk));
	jor g0784(.dina(w_n1043_1[0]),.dinb(w_n852_7[0]),.dout(n1085),.clk(gclk));
	jor g0785(.dina(w_n1041_1[0]),.dinb(w_G4089_7[0]),.dout(n1086),.clk(gclk));
	jand g0786(.dina(n1086),.dinb(n1085),.dout(n1087),.clk(gclk));
	jand g0787(.dina(n1087),.dinb(w_n854_3[1]),.dout(n1088),.clk(gclk));
	jor g0788(.dina(n1088),.dinb(w_dff_B_QtbKjWVe1_1),.dout(w_dff_A_JuenzXYu0_2),.clk(gclk));
	jor g0789(.dina(w_n1052_1[0]),.dinb(w_n852_6[2]),.dout(n1090),.clk(gclk));
	jor g0790(.dina(w_n1054_1[0]),.dinb(w_G4089_6[2]),.dout(n1091),.clk(gclk));
	jand g0791(.dina(n1091),.dinb(w_n854_3[0]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(n1092),.dinb(w_dff_B_hPqcY2iD9_1),.dout(n1093),.clk(gclk));
	jor g0793(.dina(w_n852_6[1]),.dinb(w_G70_0[0]),.dout(n1094),.clk(gclk));
	jor g0794(.dina(w_G4089_6[1]),.dinb(w_G67_0[0]),.dout(n1095),.clk(gclk));
	jand g0795(.dina(n1095),.dinb(w_G4090_3[0]),.dout(n1096),.clk(gclk));
	jand g0796(.dina(n1096),.dinb(n1094),.dout(n1097),.clk(gclk));
	jor g0797(.dina(w_dff_B_fUQ7IRTy5_0),.dinb(n1093),.dout(w_dff_A_Oq5Agr8v8_2),.clk(gclk));
	jor g0798(.dina(w_n1021_0[2]),.dinb(w_G1689_4[1]),.dout(n1099),.clk(gclk));
	jor g0799(.dina(w_n1019_0[2]),.dinb(w_n993_4[0]),.dout(n1100),.clk(gclk));
	jand g0800(.dina(n1100),.dinb(w_n999_3[1]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(n1101),.dinb(w_dff_B_BFLz6QQE7_1),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n994_4[0]),.dinb(w_G200_0[1]),.dout(n1103),.clk(gclk));
	jand g0803(.dina(w_n996_4[0]),.dinb(w_G170_0[1]),.dout(n1104),.clk(gclk));
	jor g0804(.dina(w_dff_B_69LkdRe29_0),.dinb(n1103),.dout(n1105),.clk(gclk));
	jor g0805(.dina(w_dff_B_n4Z3kC0B8_0),.dinb(n1102),.dout(n1106),.clk(gclk));
	jand g0806(.dina(n1106),.dinb(w_G137_8[2]),.dout(w_dff_A_oXtvQCRh0_2),.clk(gclk));
	jor g0807(.dina(w_n1054_0[2]),.dinb(w_G1689_4[0]),.dout(n1108),.clk(gclk));
	jor g0808(.dina(w_n1052_0[2]),.dinb(w_n993_3[2]),.dout(n1109),.clk(gclk));
	jand g0809(.dina(n1109),.dinb(w_n999_3[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(w_dff_B_jYDj2gId5_0),.dinb(n1108),.dout(n1111),.clk(gclk));
	jand g0811(.dina(w_n994_3[2]),.dinb(w_G188_0[1]),.dout(n1112),.clk(gclk));
	jand g0812(.dina(w_n996_3[2]),.dinb(w_G158_0[1]),.dout(n1113),.clk(gclk));
	jor g0813(.dina(w_dff_B_44vAecWO2_0),.dinb(n1112),.dout(n1114),.clk(gclk));
	jor g0814(.dina(w_dff_B_Fo0Afh4i9_0),.dinb(n1111),.dout(n1115),.clk(gclk));
	jand g0815(.dina(n1115),.dinb(w_G137_8[1]),.dout(w_dff_A_kmX7ykt16_2),.clk(gclk));
	jor g0816(.dina(w_n1041_0[2]),.dinb(w_G1689_3[2]),.dout(n1117),.clk(gclk));
	jor g0817(.dina(w_n1043_0[2]),.dinb(w_n993_3[1]),.dout(n1118),.clk(gclk));
	jand g0818(.dina(n1118),.dinb(w_n999_2[2]),.dout(n1119),.clk(gclk));
	jand g0819(.dina(n1119),.dinb(w_dff_B_vv2nfHoo5_1),.dout(n1120),.clk(gclk));
	jand g0820(.dina(w_n994_3[1]),.dinb(w_G155_0[1]),.dout(n1121),.clk(gclk));
	jand g0821(.dina(w_n996_3[1]),.dinb(w_G152_0[1]),.dout(n1122),.clk(gclk));
	jor g0822(.dina(w_dff_B_u5p460Ly0_0),.dinb(n1121),.dout(n1123),.clk(gclk));
	jor g0823(.dina(w_dff_B_0gPtaQdm0_0),.dinb(n1120),.dout(n1124),.clk(gclk));
	jand g0824(.dina(n1124),.dinb(w_G137_8[0]),.dout(w_dff_A_hZ4sVGkq1_2),.clk(gclk));
	jor g0825(.dina(w_n1032_0[2]),.dinb(w_G1689_3[1]),.dout(n1126),.clk(gclk));
	jor g0826(.dina(w_n1030_0[2]),.dinb(w_n993_3[0]),.dout(n1127),.clk(gclk));
	jand g0827(.dina(n1127),.dinb(w_n999_2[1]),.dout(n1128),.clk(gclk));
	jand g0828(.dina(n1128),.dinb(n1126),.dout(n1129),.clk(gclk));
	jand g0829(.dina(w_n994_3[0]),.dinb(w_G149_0[1]),.dout(n1130),.clk(gclk));
	jand g0830(.dina(w_n996_3[0]),.dinb(w_G146_0[1]),.dout(n1131),.clk(gclk));
	jor g0831(.dina(w_dff_B_sFCOBFKZ8_0),.dinb(n1130),.dout(n1132),.clk(gclk));
	jor g0832(.dina(w_dff_B_DHFhcBXc5_0),.dinb(n1129),.dout(n1133),.clk(gclk));
	jand g0833(.dina(n1133),.dinb(w_G137_7[2]),.dout(w_dff_A_IObyZMPk5_2),.clk(gclk));
	jand g0834(.dina(w_n1014_4[0]),.dinb(w_G200_0[0]),.dout(n1135),.clk(gclk));
	jand g0835(.dina(w_n1012_4[0]),.dinb(w_G170_0[0]),.dout(n1136),.clk(gclk));
	jor g0836(.dina(w_n1019_0[1]),.dinb(w_n1008_4[0]),.dout(n1137),.clk(gclk));
	jor g0837(.dina(w_n1021_0[1]),.dinb(w_G1691_4[1]),.dout(n1138),.clk(gclk));
	jand g0838(.dina(n1138),.dinb(n1137),.dout(n1139),.clk(gclk));
	jand g0839(.dina(n1139),.dinb(w_n1007_3[1]),.dout(n1140),.clk(gclk));
	jor g0840(.dina(n1140),.dinb(w_dff_B_dzFlQmzL4_1),.dout(n1141),.clk(gclk));
	jor g0841(.dina(n1141),.dinb(w_dff_B_4rKzi5ft5_1),.dout(n1142),.clk(gclk));
	jand g0842(.dina(n1142),.dinb(w_G137_7[1]),.dout(w_dff_A_GYTpg0iA4_2),.clk(gclk));
	jor g0843(.dina(w_n1054_0[1]),.dinb(w_G1691_4[0]),.dout(n1144),.clk(gclk));
	jor g0844(.dina(w_n1052_0[1]),.dinb(w_n1008_3[2]),.dout(n1145),.clk(gclk));
	jand g0845(.dina(n1145),.dinb(w_n1007_3[0]),.dout(n1146),.clk(gclk));
	jand g0846(.dina(w_dff_B_metFiBlD4_0),.dinb(n1144),.dout(n1147),.clk(gclk));
	jand g0847(.dina(w_n1014_3[2]),.dinb(w_G188_0[0]),.dout(n1148),.clk(gclk));
	jand g0848(.dina(w_n1012_3[2]),.dinb(w_G158_0[0]),.dout(n1149),.clk(gclk));
	jor g0849(.dina(w_dff_B_iKYzvaD16_0),.dinb(n1148),.dout(n1150),.clk(gclk));
	jor g0850(.dina(w_dff_B_9vShPgtL7_0),.dinb(n1147),.dout(n1151),.clk(gclk));
	jand g0851(.dina(n1151),.dinb(w_G137_7[0]),.dout(w_dff_A_8eEJ4Fst4_2),.clk(gclk));
	jor g0852(.dina(w_n1041_0[1]),.dinb(w_G1691_3[2]),.dout(n1153),.clk(gclk));
	jor g0853(.dina(w_n1043_0[1]),.dinb(w_n1008_3[1]),.dout(n1154),.clk(gclk));
	jand g0854(.dina(n1154),.dinb(w_n1007_2[2]),.dout(n1155),.clk(gclk));
	jand g0855(.dina(n1155),.dinb(w_dff_B_EFBbqyKg0_1),.dout(n1156),.clk(gclk));
	jand g0856(.dina(w_n1014_3[1]),.dinb(w_G155_0[0]),.dout(n1157),.clk(gclk));
	jand g0857(.dina(w_n1012_3[1]),.dinb(w_G152_0[0]),.dout(n1158),.clk(gclk));
	jor g0858(.dina(w_dff_B_kwmSNrEv6_0),.dinb(n1157),.dout(n1159),.clk(gclk));
	jor g0859(.dina(w_dff_B_0FbXlvoh7_0),.dinb(n1156),.dout(n1160),.clk(gclk));
	jand g0860(.dina(n1160),.dinb(w_G137_6[2]),.dout(w_dff_A_2N0KkA108_2),.clk(gclk));
	jor g0861(.dina(w_n1032_0[1]),.dinb(w_G1691_3[1]),.dout(n1162),.clk(gclk));
	jor g0862(.dina(w_n1030_0[1]),.dinb(w_n1008_3[0]),.dout(n1163),.clk(gclk));
	jand g0863(.dina(n1163),.dinb(w_n1007_2[1]),.dout(n1164),.clk(gclk));
	jand g0864(.dina(n1164),.dinb(n1162),.dout(n1165),.clk(gclk));
	jand g0865(.dina(w_n1014_3[0]),.dinb(w_G149_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n1012_3[0]),.dinb(w_G146_0[0]),.dout(n1167),.clk(gclk));
	jor g0867(.dina(w_dff_B_l83lBKCX4_0),.dinb(n1166),.dout(n1168),.clk(gclk));
	jor g0868(.dina(w_dff_B_MEIhhaKH4_0),.dinb(n1165),.dout(n1169),.clk(gclk));
	jand g0869(.dina(n1169),.dinb(w_G137_6[1]),.dout(w_dff_A_gyEHSMrf9_2),.clk(gclk));
	jnot g0870(.din(G135),.dout(n1171),.clk(gclk));
	jnot g0871(.din(G4115),.dout(n1172),.clk(gclk));
	jor g0872(.dina(n1172),.dinb(n1171),.dout(n1173),.clk(gclk));
	jnot g0873(.din(w_n428_1[0]),.dout(n1174),.clk(gclk));
	jor g0874(.dina(n1174),.dinb(w_G3724_0[2]),.dout(n1175),.clk(gclk));
	jnot g0875(.din(w_G3717_0[1]),.dout(n1176),.clk(gclk));
	jnot g0876(.din(w_G3724_0[1]),.dout(n1177),.clk(gclk));
	jxor g0877(.dina(w_n790_0[0]),.dinb(w_dff_B_WLeseU1z1_1),.dout(n1178),.clk(gclk));
	jnot g0878(.din(n1178),.dout(n1179),.clk(gclk));
	jor g0879(.dina(w_n1179_0[1]),.dinb(w_n1177_0[1]),.dout(n1180),.clk(gclk));
	jand g0880(.dina(n1180),.dinb(w_dff_B_fkywhnmy6_1),.dout(n1181),.clk(gclk));
	jand g0881(.dina(n1181),.dinb(w_dff_B_eTcQlCR77_1),.dout(n1182),.clk(gclk));
	jor g0882(.dina(w_n795_1[0]),.dinb(w_n1177_0[0]),.dout(n1183),.clk(gclk));
	jor g0883(.dina(w_G3724_0[0]),.dinb(w_G123_0[1]),.dout(n1184),.clk(gclk));
	jand g0884(.dina(n1184),.dinb(w_G3717_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(w_dff_B_REvoa9Uk5_0),.dinb(n1183),.dout(n1186),.clk(gclk));
	jor g0886(.dina(n1186),.dinb(w_dff_B_AcWpHut54_1),.dout(n1187),.clk(gclk));
	jand g0887(.dina(n1187),.dinb(w_dff_B_IR1js6PY9_1),.dout(w_dff_A_6D6rviAx0_2),.clk(gclk));
	jxor g0888(.dina(w_n1179_0[0]),.dinb(w_n795_0[2]),.dout(w_dff_A_yfUFm8z19_2),.clk(gclk));
	jand g0889(.dina(w_n750_5[1]),.dinb(w_G123_0[0]),.dout(n1190),.clk(gclk));
	jor g0890(.dina(w_n795_0[1]),.dinb(w_n749_9[2]),.dout(n1191),.clk(gclk));
	jand g0891(.dina(w_n428_0[2]),.dinb(w_n749_9[1]),.dout(n1192),.clk(gclk));
	jor g0892(.dina(n1192),.dinb(w_G4092_6[0]),.dout(n1193),.clk(gclk));
	jnot g0893(.din(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_dff_B_s4WOZmBm6_0),.dinb(n1191),.dout(n1195),.clk(gclk));
	jor g0895(.dina(n1195),.dinb(w_dff_B_BGM5W6S45_1),.dout(n1196),.clk(gclk));
	jnot g0896(.din(w_n1196_1[2]),.dout(w_dff_A_JP0ztOG01_1),.clk(gclk));
	jand g0897(.dina(w_n750_5[0]),.dinb(w_dff_B_4nhfmZyy7_1),.dout(n1198),.clk(gclk));
	jand g0898(.dina(w_n433_0[1]),.dinb(w_n749_9[0]),.dout(n1199),.clk(gclk));
	jnot g0899(.din(n1199),.dout(n1200),.clk(gclk));
	jnot g0900(.din(w_G4092_5[2]),.dout(n1201),.clk(gclk));
	jor g0901(.dina(w_n969_0[0]),.dinb(w_n749_8[2]),.dout(n1202),.clk(gclk));
	jand g0902(.dina(n1202),.dinb(w_n1201_0[2]),.dout(n1203),.clk(gclk));
	jand g0903(.dina(n1203),.dinb(w_dff_B_TA9c7iQR3_1),.dout(n1204),.clk(gclk));
	jor g0904(.dina(n1204),.dinb(w_dff_B_UZUkPoFP0_1),.dout(n1205),.clk(gclk));
	jnot g0905(.din(w_n1205_1[2]),.dout(w_dff_A_BfQNuq0O6_1),.clk(gclk));
	jand g0906(.dina(w_n750_4[2]),.dinb(w_dff_B_kYjK86vv1_1),.dout(n1207),.clk(gclk));
	jor g0907(.dina(w_n986_0[0]),.dinb(w_n749_8[1]),.dout(n1208),.clk(gclk));
	jand g0908(.dina(w_n423_0[1]),.dinb(w_n749_8[0]),.dout(n1209),.clk(gclk));
	jor g0909(.dina(n1209),.dinb(w_G4092_5[1]),.dout(n1210),.clk(gclk));
	jnot g0910(.din(n1210),.dout(n1211),.clk(gclk));
	jand g0911(.dina(w_dff_B_0wWjNpv39_0),.dinb(n1208),.dout(n1212),.clk(gclk));
	jor g0912(.dina(n1212),.dinb(w_dff_B_kWb1quw83_1),.dout(n1213),.clk(gclk));
	jnot g0913(.din(w_n1213_1[2]),.dout(w_dff_A_EMYGxBMS3_1),.clk(gclk));
	jand g0914(.dina(w_n750_4[1]),.dinb(w_dff_B_F7iw6GAC2_1),.dout(n1215),.clk(gclk));
	jnot g0915(.din(n1215),.dout(n1216),.clk(gclk));
	jand g0916(.dina(w_n989_0[0]),.dinb(w_G4091_2[2]),.dout(n1217),.clk(gclk));
	jand g0917(.dina(w_n412_0[1]),.dinb(w_n749_7[2]),.dout(n1218),.clk(gclk));
	jor g0918(.dina(n1218),.dinb(w_G4092_5[0]),.dout(n1219),.clk(gclk));
	jor g0919(.dina(w_dff_B_fx5k9FZY9_0),.dinb(n1217),.dout(n1220),.clk(gclk));
	jand g0920(.dina(n1220),.dinb(w_dff_B_J8o4nnxb3_1),.dout(G830_fa_),.clk(gclk));
	jand g0921(.dina(w_n680_0[0]),.dinb(w_G245_0[0]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(w_dff_B_yrPwA8uG8_0),.dinb(w_n935_0[0]),.dout(n1223),.clk(gclk));
	jnot g0923(.din(w_G998_0),.dout(n1224),.clk(gclk));
	jand g0924(.dina(w_n318_0[0]),.dinb(w_G601_0),.dout(n1225),.clk(gclk));
	jand g0925(.dina(n1225),.dinb(w_G559_0[0]),.dout(n1226),.clk(gclk));
	jand g0926(.dina(w_dff_B_tam88bC02_0),.dinb(w_n670_0[0]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_dff_B_N5kgZ4q98_0),.dinb(n1224),.dout(n1228),.clk(gclk));
	jand g0928(.dina(n1228),.dinb(w_dff_B_GBcMuDia6_1),.dout(w_dff_A_895FGv130_2),.clk(gclk));
	jand g0929(.dina(w_n750_4[0]),.dinb(w_dff_B_uKlhyMAY6_1),.dout(n1230),.clk(gclk));
	jand g0930(.dina(w_n551_0[1]),.dinb(w_n749_7[1]),.dout(n1231),.clk(gclk));
	jnot g0931(.din(n1231),.dout(n1232),.clk(gclk));
	jor g0932(.dina(w_n944_0[0]),.dinb(w_n749_7[0]),.dout(n1233),.clk(gclk));
	jand g0933(.dina(n1233),.dinb(w_n1201_0[1]),.dout(n1234),.clk(gclk));
	jand g0934(.dina(n1234),.dinb(w_dff_B_E104wsN56_1),.dout(n1235),.clk(gclk));
	jor g0935(.dina(n1235),.dinb(w_dff_B_0Z5IiwPq7_1),.dout(n1236),.clk(gclk));
	jnot g0936(.din(w_n1236_1[2]),.dout(w_dff_A_6KcRPZEY1_1),.clk(gclk));
	jand g0937(.dina(w_n750_3[2]),.dinb(w_dff_B_Or80r8Bu4_1),.dout(n1238),.clk(gclk));
	jnot g0938(.din(n1238),.dout(n1239),.clk(gclk));
	jand g0939(.dina(w_n949_0[0]),.dinb(w_G4091_2[1]),.dout(n1240),.clk(gclk));
	jand g0940(.dina(w_n459_0[0]),.dinb(w_n749_6[2]),.dout(n1241),.clk(gclk));
	jor g0941(.dina(n1241),.dinb(w_G4092_4[2]),.dout(n1242),.clk(gclk));
	jor g0942(.dina(w_dff_B_Vhmy5KCT8_0),.dinb(n1240),.dout(n1243),.clk(gclk));
	jand g0943(.dina(n1243),.dinb(w_dff_B_jXg2uAaj1_1),.dout(G865_fa_),.clk(gclk));
	jand g0944(.dina(w_n750_3[1]),.dinb(w_dff_B_3LTRgAEm6_1),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n517_0[0]),.dinb(w_n749_6[1]),.dout(n1246),.clk(gclk));
	jnot g0946(.din(n1246),.dout(n1247),.clk(gclk));
	jor g0947(.dina(w_n957_0[0]),.dinb(w_n749_6[0]),.dout(n1248),.clk(gclk));
	jand g0948(.dina(n1248),.dinb(w_n1201_0[0]),.dout(n1249),.clk(gclk));
	jand g0949(.dina(n1249),.dinb(w_dff_B_Cp2TkbYB7_1),.dout(n1250),.clk(gclk));
	jor g0950(.dina(n1250),.dinb(w_dff_B_IQtoGsNT7_1),.dout(n1251),.clk(gclk));
	jnot g0951(.din(w_n1251_1[2]),.dout(w_dff_A_ybOm80nJ7_1),.clk(gclk));
	jand g0952(.dina(w_n750_3[0]),.dinb(w_dff_B_aljd1Jnr4_1),.dout(n1253),.clk(gclk));
	jnot g0953(.din(n1253),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n964_0[0]),.dinb(w_G4091_2[0]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n504_0[0]),.dinb(w_n749_5[2]),.dout(n1256),.clk(gclk));
	jor g0956(.dina(n1256),.dinb(w_G4092_4[1]),.dout(n1257),.clk(gclk));
	jor g0957(.dina(w_dff_B_75NlZSdJ8_0),.dinb(n1255),.dout(n1258),.clk(gclk));
	jand g0958(.dina(n1258),.dinb(w_dff_B_7ZKBsrZl6_1),.dout(G869_fa_),.clk(gclk));
	jor g0959(.dina(w_G4089_6[0]),.dinb(w_G109_0[1]),.dout(n1260),.clk(gclk));
	jor g0960(.dina(w_n852_6[0]),.dinb(w_G106_0[1]),.dout(n1261),.clk(gclk));
	jand g0961(.dina(n1261),.dinb(w_G4090_2[2]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(n1262),.dinb(w_dff_B_RL3xREXt5_1),.dout(n1263),.clk(gclk));
	jor g0963(.dina(w_n1236_1[1]),.dinb(w_n852_5[2]),.dout(n1264),.clk(gclk));
	jor g0964(.dina(w_n1196_1[1]),.dinb(w_G4089_5[2]),.dout(n1265),.clk(gclk));
	jand g0965(.dina(n1265),.dinb(w_n854_2[2]),.dout(n1266),.clk(gclk));
	jand g0966(.dina(n1266),.dinb(n1264),.dout(n1267),.clk(gclk));
	jor g0967(.dina(n1267),.dinb(w_dff_B_awItk95I5_1),.dout(w_dff_A_9sxuK1rx0_2),.clk(gclk));
	jor g0968(.dina(w_n1196_1[0]),.dinb(w_G4088_6[0]),.dout(n1269),.clk(gclk));
	jor g0969(.dina(w_n1236_1[0]),.dinb(w_n797_6[0]),.dout(n1270),.clk(gclk));
	jand g0970(.dina(n1270),.dinb(w_n800_2[2]),.dout(n1271),.clk(gclk));
	jand g0971(.dina(n1271),.dinb(w_dff_B_gFIIPHp96_1),.dout(n1272),.clk(gclk));
	jor g0972(.dina(w_n797_5[2]),.dinb(w_G106_0[0]),.dout(n1273),.clk(gclk));
	jor g0973(.dina(w_G4088_5[2]),.dinb(w_G109_0[0]),.dout(n1274),.clk(gclk));
	jand g0974(.dina(n1274),.dinb(w_G4087_2[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(n1275),.dinb(n1273),.dout(n1276),.clk(gclk));
	jor g0976(.dina(w_dff_B_VNDVWmfp6_0),.dinb(n1272),.dout(w_dff_A_9ZseDTY54_2),.clk(gclk));
	jor g0977(.dina(w_n1205_1[1]),.dinb(w_G4088_5[1]),.dout(n1278),.clk(gclk));
	jnot g0978(.din(w_G865_0),.dout(n1279),.clk(gclk));
	jor g0979(.dina(w_n1279_1[1]),.dinb(w_n797_5[1]),.dout(n1280),.clk(gclk));
	jand g0980(.dina(n1280),.dinb(w_n800_2[1]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(n1281),.dinb(w_dff_B_humdkuXK2_1),.dout(n1282),.clk(gclk));
	jor g0982(.dina(w_n797_5[0]),.dinb(w_G49_0[1]),.dout(n1283),.clk(gclk));
	jor g0983(.dina(w_G4088_5[0]),.dinb(w_G46_0[1]),.dout(n1284),.clk(gclk));
	jand g0984(.dina(n1284),.dinb(w_G4087_2[1]),.dout(n1285),.clk(gclk));
	jand g0985(.dina(n1285),.dinb(n1283),.dout(n1286),.clk(gclk));
	jor g0986(.dina(w_dff_B_EGaddTYu8_0),.dinb(n1282),.dout(w_dff_A_1o2NTLEO3_2),.clk(gclk));
	jor g0987(.dina(w_n1213_1[1]),.dinb(w_G4088_4[2]),.dout(n1288),.clk(gclk));
	jor g0988(.dina(w_n1251_1[1]),.dinb(w_n797_4[2]),.dout(n1289),.clk(gclk));
	jand g0989(.dina(n1289),.dinb(w_n800_2[0]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(n1290),.dinb(w_dff_B_IzLWxCMd6_1),.dout(n1291),.clk(gclk));
	jor g0991(.dina(w_n797_4[1]),.dinb(w_G103_0[1]),.dout(n1292),.clk(gclk));
	jor g0992(.dina(w_G4088_4[1]),.dinb(w_G100_0[1]),.dout(n1293),.clk(gclk));
	jand g0993(.dina(n1293),.dinb(w_G4087_2[0]),.dout(n1294),.clk(gclk));
	jand g0994(.dina(n1294),.dinb(n1292),.dout(n1295),.clk(gclk));
	jor g0995(.dina(w_dff_B_TSdQhI3G0_0),.dinb(n1291),.dout(w_dff_A_UFCuDxvQ5_2),.clk(gclk));
	jnot g0996(.din(w_G830_0),.dout(n1297),.clk(gclk));
	jor g0997(.dina(w_n1297_1[1]),.dinb(w_G4088_4[0]),.dout(n1298),.clk(gclk));
	jnot g0998(.din(w_G869_0),.dout(n1299),.clk(gclk));
	jor g0999(.dina(w_n1299_1[1]),.dinb(w_n797_4[0]),.dout(n1300),.clk(gclk));
	jand g1000(.dina(n1300),.dinb(w_n800_1[2]),.dout(n1301),.clk(gclk));
	jand g1001(.dina(n1301),.dinb(w_dff_B_Q8ABeuZd7_1),.dout(n1302),.clk(gclk));
	jor g1002(.dina(w_n797_3[2]),.dinb(w_G40_0[1]),.dout(n1303),.clk(gclk));
	jor g1003(.dina(w_G4088_3[2]),.dinb(w_G91_0[1]),.dout(n1304),.clk(gclk));
	jand g1004(.dina(n1304),.dinb(w_G4087_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(n1305),.dinb(n1303),.dout(n1306),.clk(gclk));
	jor g1006(.dina(w_dff_B_aZcDLtDG6_0),.dinb(n1302),.dout(w_dff_A_LJKa69Qm9_2),.clk(gclk));
	jor g1007(.dina(w_n1205_1[0]),.dinb(w_G4089_5[1]),.dout(n1308),.clk(gclk));
	jor g1008(.dina(w_n1279_1[0]),.dinb(w_n852_5[1]),.dout(n1309),.clk(gclk));
	jand g1009(.dina(n1309),.dinb(w_n854_2[1]),.dout(n1310),.clk(gclk));
	jand g1010(.dina(n1310),.dinb(w_dff_B_1fOuwH6L7_1),.dout(n1311),.clk(gclk));
	jor g1011(.dina(w_n852_5[0]),.dinb(w_G49_0[0]),.dout(n1312),.clk(gclk));
	jor g1012(.dina(w_G4089_5[0]),.dinb(w_G46_0[0]),.dout(n1313),.clk(gclk));
	jand g1013(.dina(n1313),.dinb(w_G4090_2[1]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(n1314),.dinb(n1312),.dout(n1315),.clk(gclk));
	jor g1015(.dina(w_dff_B_pwxvlKCd3_0),.dinb(n1311),.dout(w_dff_A_YNkz6Tgg6_2),.clk(gclk));
	jor g1016(.dina(w_n1213_1[0]),.dinb(w_G4089_4[2]),.dout(n1317),.clk(gclk));
	jor g1017(.dina(w_n1251_1[0]),.dinb(w_n852_4[2]),.dout(n1318),.clk(gclk));
	jand g1018(.dina(n1318),.dinb(w_n854_2[0]),.dout(n1319),.clk(gclk));
	jand g1019(.dina(n1319),.dinb(w_dff_B_T1W1r0Mi2_1),.dout(n1320),.clk(gclk));
	jor g1020(.dina(w_n852_4[1]),.dinb(w_G103_0[0]),.dout(n1321),.clk(gclk));
	jor g1021(.dina(w_G4089_4[1]),.dinb(w_G100_0[0]),.dout(n1322),.clk(gclk));
	jand g1022(.dina(n1322),.dinb(w_G4090_2[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(n1323),.dinb(n1321),.dout(n1324),.clk(gclk));
	jor g1024(.dina(w_dff_B_GRzCDFLx2_0),.dinb(n1320),.dout(w_dff_A_iVlpqlh74_2),.clk(gclk));
	jor g1025(.dina(w_n1297_1[0]),.dinb(w_G4089_4[0]),.dout(n1326),.clk(gclk));
	jor g1026(.dina(w_n1299_1[0]),.dinb(w_n852_4[0]),.dout(n1327),.clk(gclk));
	jand g1027(.dina(n1327),.dinb(w_n854_1[2]),.dout(n1328),.clk(gclk));
	jand g1028(.dina(n1328),.dinb(w_dff_B_C4l1m0gX6_1),.dout(n1329),.clk(gclk));
	jor g1029(.dina(w_n852_3[2]),.dinb(w_G40_0[0]),.dout(n1330),.clk(gclk));
	jor g1030(.dina(w_G4089_3[2]),.dinb(w_G91_0[0]),.dout(n1331),.clk(gclk));
	jand g1031(.dina(n1331),.dinb(w_G4090_1[2]),.dout(n1332),.clk(gclk));
	jand g1032(.dina(n1332),.dinb(n1330),.dout(n1333),.clk(gclk));
	jor g1033(.dina(w_dff_B_tCYsu0WS0_0),.dinb(n1329),.dout(w_dff_A_8lfa568n2_2),.clk(gclk));
	jor g1034(.dina(w_n1297_0[2]),.dinb(w_G1689_3[0]),.dout(n1335),.clk(gclk));
	jor g1035(.dina(w_n1299_0[2]),.dinb(w_n993_2[2]),.dout(n1336),.clk(gclk));
	jand g1036(.dina(n1336),.dinb(w_n999_2[0]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(n1337),.dinb(w_dff_B_oMESUjmC8_1),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n994_2[2]),.dinb(w_G203_0[1]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n996_2[2]),.dinb(w_G173_0[1]),.dout(n1340),.clk(gclk));
	jor g1040(.dina(w_dff_B_o2lYWXg34_0),.dinb(n1339),.dout(n1341),.clk(gclk));
	jor g1041(.dina(w_dff_B_o3U269by6_0),.dinb(n1338),.dout(n1342),.clk(gclk));
	jand g1042(.dina(n1342),.dinb(w_G137_6[0]),.dout(w_dff_A_iUpifcdH2_2),.clk(gclk));
	jor g1043(.dina(w_n1251_0[2]),.dinb(w_n993_2[1]),.dout(n1344),.clk(gclk));
	jor g1044(.dina(w_n1213_0[2]),.dinb(w_G1689_2[2]),.dout(n1345),.clk(gclk));
	jand g1045(.dina(n1345),.dinb(w_n999_1[2]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(n1346),.dinb(w_dff_B_WtmtCWCJ1_1),.dout(n1347),.clk(gclk));
	jand g1047(.dina(w_n994_2[1]),.dinb(w_G197_0[1]),.dout(n1348),.clk(gclk));
	jand g1048(.dina(w_n996_2[1]),.dinb(w_G167_0[1]),.dout(n1349),.clk(gclk));
	jor g1049(.dina(w_dff_B_YFV8slcf0_0),.dinb(n1348),.dout(n1350),.clk(gclk));
	jor g1050(.dina(w_dff_B_k8e4oTpX8_0),.dinb(n1347),.dout(n1351),.clk(gclk));
	jand g1051(.dina(n1351),.dinb(w_G137_5[2]),.dout(w_dff_A_2tJJd17T5_2),.clk(gclk));
	jand g1052(.dina(w_n994_2[0]),.dinb(w_G194_0[1]),.dout(n1353),.clk(gclk));
	jand g1053(.dina(w_n996_2[0]),.dinb(w_G164_0[1]),.dout(n1354),.clk(gclk));
	jor g1054(.dina(w_dff_B_Ym1YPgLI8_0),.dinb(n1353),.dout(n1355),.clk(gclk));
	jor g1055(.dina(w_n1205_0[2]),.dinb(w_G1689_2[1]),.dout(n1356),.clk(gclk));
	jor g1056(.dina(w_n1279_0[2]),.dinb(w_n993_2[0]),.dout(n1357),.clk(gclk));
	jand g1057(.dina(n1357),.dinb(w_dff_B_ObQwgJC15_1),.dout(n1358),.clk(gclk));
	jand g1058(.dina(n1358),.dinb(w_n999_1[1]),.dout(n1359),.clk(gclk));
	jor g1059(.dina(n1359),.dinb(w_dff_B_m5sqUrVV8_1),.dout(n1360),.clk(gclk));
	jand g1060(.dina(n1360),.dinb(w_G137_5[1]),.dout(w_dff_A_8Et3bTWw1_2),.clk(gclk));
	jand g1061(.dina(w_n994_1[2]),.dinb(w_G191_0[1]),.dout(n1362),.clk(gclk));
	jand g1062(.dina(w_n996_1[2]),.dinb(w_G161_0[1]),.dout(n1363),.clk(gclk));
	jor g1063(.dina(w_dff_B_KcfGaCcD5_0),.dinb(n1362),.dout(n1364),.clk(gclk));
	jor g1064(.dina(w_n1196_0[2]),.dinb(w_G1689_2[0]),.dout(n1365),.clk(gclk));
	jor g1065(.dina(w_n1236_0[2]),.dinb(w_n993_1[2]),.dout(n1366),.clk(gclk));
	jand g1066(.dina(n1366),.dinb(w_dff_B_EWcgwott5_1),.dout(n1367),.clk(gclk));
	jand g1067(.dina(n1367),.dinb(w_n999_1[0]),.dout(n1368),.clk(gclk));
	jor g1068(.dina(n1368),.dinb(w_dff_B_AZuUwZqn7_1),.dout(n1369),.clk(gclk));
	jand g1069(.dina(n1369),.dinb(w_G137_5[0]),.dout(w_dff_A_W8e3w3NF5_2),.clk(gclk));
	jor g1070(.dina(w_n1297_0[1]),.dinb(w_G1691_3[0]),.dout(n1371),.clk(gclk));
	jor g1071(.dina(w_n1299_0[1]),.dinb(w_n1008_2[2]),.dout(n1372),.clk(gclk));
	jand g1072(.dina(n1372),.dinb(w_n1007_2[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(n1373),.dinb(w_dff_B_6BA4nhSw3_1),.dout(n1374),.clk(gclk));
	jand g1074(.dina(w_n1014_2[2]),.dinb(w_G203_0[0]),.dout(n1375),.clk(gclk));
	jand g1075(.dina(w_n1012_2[2]),.dinb(w_G173_0[0]),.dout(n1376),.clk(gclk));
	jor g1076(.dina(w_dff_B_ihjrzGeK4_0),.dinb(n1375),.dout(n1377),.clk(gclk));
	jor g1077(.dina(w_dff_B_XKntAtJb8_0),.dinb(n1374),.dout(n1378),.clk(gclk));
	jand g1078(.dina(n1378),.dinb(w_G137_4[2]),.dout(w_dff_A_JhrkJhl39_2),.clk(gclk));
	jand g1079(.dina(w_n1014_2[1]),.dinb(w_G197_0[0]),.dout(n1380),.clk(gclk));
	jand g1080(.dina(w_n1012_2[1]),.dinb(w_G167_0[0]),.dout(n1381),.clk(gclk));
	jor g1081(.dina(w_dff_B_QCQEHJBJ9_0),.dinb(n1380),.dout(n1382),.clk(gclk));
	jor g1082(.dina(w_n1213_0[1]),.dinb(w_G1691_2[2]),.dout(n1383),.clk(gclk));
	jor g1083(.dina(w_n1251_0[1]),.dinb(w_n1008_2[1]),.dout(n1384),.clk(gclk));
	jand g1084(.dina(n1384),.dinb(n1383),.dout(n1385),.clk(gclk));
	jand g1085(.dina(n1385),.dinb(w_n1007_1[2]),.dout(n1386),.clk(gclk));
	jor g1086(.dina(n1386),.dinb(w_dff_B_jthn2JR95_1),.dout(n1387),.clk(gclk));
	jand g1087(.dina(n1387),.dinb(w_G137_4[1]),.dout(w_dff_A_EU9AjEys6_2),.clk(gclk));
	jor g1088(.dina(w_n1205_0[1]),.dinb(w_G1691_2[1]),.dout(n1389),.clk(gclk));
	jor g1089(.dina(w_n1279_0[1]),.dinb(w_n1008_2[0]),.dout(n1390),.clk(gclk));
	jand g1090(.dina(n1390),.dinb(w_n1007_1[1]),.dout(n1391),.clk(gclk));
	jand g1091(.dina(n1391),.dinb(w_dff_B_IRc6Jqif2_1),.dout(n1392),.clk(gclk));
	jand g1092(.dina(w_n1014_2[0]),.dinb(w_G194_0[0]),.dout(n1393),.clk(gclk));
	jand g1093(.dina(w_n1012_2[0]),.dinb(w_G164_0[0]),.dout(n1394),.clk(gclk));
	jor g1094(.dina(w_dff_B_j1n3kkOT6_0),.dinb(n1393),.dout(n1395),.clk(gclk));
	jor g1095(.dina(w_dff_B_aECCcNub3_0),.dinb(n1392),.dout(n1396),.clk(gclk));
	jand g1096(.dina(n1396),.dinb(w_G137_4[0]),.dout(w_dff_A_BvotNGEA0_2),.clk(gclk));
	jor g1097(.dina(w_n1236_0[1]),.dinb(w_n1008_1[2]),.dout(n1398),.clk(gclk));
	jor g1098(.dina(w_n1196_0[1]),.dinb(w_G1691_2[0]),.dout(n1399),.clk(gclk));
	jand g1099(.dina(n1399),.dinb(w_n1007_1[0]),.dout(n1400),.clk(gclk));
	jand g1100(.dina(n1400),.dinb(n1398),.dout(n1401),.clk(gclk));
	jand g1101(.dina(w_n1014_1[2]),.dinb(w_G191_0[0]),.dout(n1402),.clk(gclk));
	jand g1102(.dina(w_n1012_1[2]),.dinb(w_G161_0[0]),.dout(n1403),.clk(gclk));
	jor g1103(.dina(w_dff_B_E3wrtXIv4_0),.dinb(n1402),.dout(n1404),.clk(gclk));
	jor g1104(.dina(w_dff_B_80SRCvM26_0),.dinb(n1401),.dout(n1405),.clk(gclk));
	jand g1105(.dina(n1405),.dinb(w_G137_3[2]),.dout(w_dff_A_et8vM2y52_2),.clk(gclk));
	jand g1106(.dina(w_n746_0[0]),.dinb(w_n648_0[2]),.dout(n1407),.clk(gclk));
	jxor g1107(.dina(w_n977_0[0]),.dinb(w_n654_1[0]),.dout(n1408),.clk(gclk));
	jxor g1108(.dina(n1408),.dinb(w_n644_0[0]),.dout(n1409),.clk(gclk));
	jxor g1109(.dina(w_dff_B_T4ChUrjp5_0),.dinb(n1407),.dout(n1410),.clk(gclk));
	jor g1110(.dina(w_n1410_0[2]),.dinb(w_n737_0[2]),.dout(n1411),.clk(gclk));
	jnot g1111(.din(w_G2174_0[2]),.dout(n1412),.clk(gclk));
	jnot g1112(.din(w_n719_0[0]),.dout(n1413),.clk(gclk));
	jnot g1113(.din(w_n720_0[0]),.dout(n1414),.clk(gclk));
	jor g1114(.dina(w_n821_0[0]),.dinb(w_dff_B_mAlA7HAG8_1),.dout(n1415),.clk(gclk));
	jand g1115(.dina(n1415),.dinb(w_dff_B_Qoa6Ht6s8_1),.dout(n1416),.clk(gclk));
	jxor g1116(.dina(w_n742_0[0]),.dinb(w_n654_0[2]),.dout(n1417),.clk(gclk));
	jxor g1117(.dina(n1417),.dinb(w_n792_0[0]),.dout(n1418),.clk(gclk));
	jnot g1118(.din(w_n660_0[1]),.dout(n1419),.clk(gclk));
	jand g1119(.dina(w_n745_0[0]),.dinb(w_n648_0[1]),.dout(n1420),.clk(gclk));
	jand g1120(.dina(n1420),.dinb(w_dff_B_fuURMbT48_1),.dout(n1421),.clk(gclk));
	jxor g1121(.dina(n1421),.dinb(w_dff_B_g9698oLR9_1),.dout(n1422),.clk(gclk));
	jor g1122(.dina(w_n1422_0[1]),.dinb(w_n1416_0[1]),.dout(n1423),.clk(gclk));
	jand g1123(.dina(n1423),.dinb(w_n1412_0[2]),.dout(n1424),.clk(gclk));
	jand g1124(.dina(n1424),.dinb(w_dff_B_T4kygeEA9_1),.dout(n1425),.clk(gclk));
	jnot g1125(.din(w_n1425_0[1]),.dout(n1426),.clk(gclk));
	jnot g1126(.din(w_n641_1[0]),.dout(n1427),.clk(gclk));
	jand g1127(.dina(w_n1416_0[0]),.dinb(w_dff_B_CGHTI8A53_1),.dout(n1428),.clk(gclk));
	jor g1128(.dina(w_n1428_0[1]),.dinb(w_n1422_0[0]),.dout(n1429),.clk(gclk));
	jnot g1129(.din(w_n1429_0[1]),.dout(n1430),.clk(gclk));
	jnot g1130(.din(w_n1410_0[1]),.dout(n1431),.clk(gclk));
	jand g1131(.dina(w_n1428_0[0]),.dinb(n1431),.dout(n1432),.clk(gclk));
	jor g1132(.dina(n1432),.dinb(w_n1412_0[1]),.dout(n1433),.clk(gclk));
	jor g1133(.dina(n1433),.dinb(n1430),.dout(n1434),.clk(gclk));
	jand g1134(.dina(n1434),.dinb(n1426),.dout(n1435),.clk(gclk));
	jor g1135(.dina(w_n728_0[0]),.dinb(w_n637_0[0]),.dout(n1436),.clk(gclk));
	jxor g1136(.dina(w_dff_B_YmCA8NpP5_0),.dinb(w_n733_0[1]),.dout(n1437),.clk(gclk));
	jxor g1137(.dina(w_dff_B_HFXHnHTq0_0),.dinb(w_n735_0[1]),.dout(n1438),.clk(gclk));
	jor g1138(.dina(n1438),.dinb(w_G2174_0[1]),.dout(n1439),.clk(gclk));
	jor g1139(.dina(w_n735_0[0]),.dinb(w_n640_0[0]),.dout(n1440),.clk(gclk));
	jor g1140(.dina(w_n819_0[0]),.dinb(w_n628_0[0]),.dout(n1441),.clk(gclk));
	jor g1141(.dina(w_n733_0[0]),.dinb(w_n814_0[0]),.dout(n1442),.clk(gclk));
	jor g1142(.dina(n1442),.dinb(w_n639_0[0]),.dout(n1443),.clk(gclk));
	jand g1143(.dina(n1443),.dinb(w_dff_B_X7h3zKJR7_1),.dout(n1444),.clk(gclk));
	jxor g1144(.dina(n1444),.dinb(n1440),.dout(n1445),.clk(gclk));
	jor g1145(.dina(n1445),.dinb(w_n1412_0[0]),.dout(n1446),.clk(gclk));
	jand g1146(.dina(n1446),.dinb(w_dff_B_gkOm9f2C8_1),.dout(n1447),.clk(gclk));
	jxor g1147(.dina(w_n620_0[1]),.dinb(w_n618_0[0]),.dout(n1448),.clk(gclk));
	jxor g1148(.dina(w_n767_0[0]),.dinb(w_n624_0[0]),.dout(n1449),.clk(gclk));
	jxor g1149(.dina(n1449),.dinb(w_dff_B_HMWdFj7t1_1),.dout(n1450),.clk(gclk));
	jxor g1150(.dina(w_dff_B_c3XXmCf30_0),.dinb(n1447),.dout(n1451),.clk(gclk));
	jnot g1151(.din(w_n1451_0[1]),.dout(n1452),.clk(gclk));
	jand g1152(.dina(w_dff_B_99f1ywRJ4_0),.dinb(n1435),.dout(n1453),.clk(gclk));
	jor g1153(.dina(w_n737_0[1]),.dinb(w_n641_0[2]),.dout(n1454),.clk(gclk));
	jor g1154(.dina(n1454),.dinb(w_n1410_0[0]),.dout(n1455),.clk(gclk));
	jand g1155(.dina(n1455),.dinb(w_G2174_0[0]),.dout(n1456),.clk(gclk));
	jand g1156(.dina(n1456),.dinb(w_n1429_0[0]),.dout(n1457),.clk(gclk));
	jor g1157(.dina(n1457),.dinb(w_n1425_0[0]),.dout(n1458),.clk(gclk));
	jand g1158(.dina(w_n1451_0[0]),.dinb(n1458),.dout(n1459),.clk(gclk));
	jor g1159(.dina(n1459),.dinb(w_n749_5[1]),.dout(n1460),.clk(gclk));
	jor g1160(.dina(n1460),.dinb(w_dff_B_z7gTYVop1_1),.dout(n1461),.clk(gclk));
	jand g1161(.dina(w_G351_1[0]),.dinb(w_G248_4[1]),.dout(n1462),.clk(gclk));
	jand g1162(.dina(w_n374_0[2]),.dinb(w_G251_4[0]),.dout(n1463),.clk(gclk));
	jor g1163(.dina(n1463),.dinb(w_n377_0[1]),.dout(n1464),.clk(gclk));
	jor g1164(.dina(n1464),.dinb(w_dff_B_Ifi5KaPP0_1),.dout(n1465),.clk(gclk));
	jand g1165(.dina(w_n374_0[1]),.dinb(w_n406_4[0]),.dout(n1466),.clk(gclk));
	jand g1166(.dina(w_G351_0[2]),.dinb(w_n408_4[1]),.dout(n1467),.clk(gclk));
	jor g1167(.dina(n1467),.dinb(n1466),.dout(n1468),.clk(gclk));
	jor g1168(.dina(n1468),.dinb(w_G534_0[2]),.dout(n1469),.clk(gclk));
	jand g1169(.dina(n1469),.dinb(n1465),.dout(n1470),.clk(gclk));
	jand g1170(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1471),.clk(gclk));
	jand g1171(.dina(w_n387_0[2]),.dinb(w_G251_3[2]),.dout(n1472),.clk(gclk));
	jor g1172(.dina(n1472),.dinb(w_n389_0[1]),.dout(n1473),.clk(gclk));
	jor g1173(.dina(n1473),.dinb(w_dff_B_3bgIAedx2_1),.dout(n1474),.clk(gclk));
	jand g1174(.dina(w_n387_0[1]),.dinb(w_n406_3[2]),.dout(n1475),.clk(gclk));
	jand g1175(.dina(w_G341_0[2]),.dinb(w_n408_4[0]),.dout(n1476),.clk(gclk));
	jor g1176(.dina(n1476),.dinb(n1475),.dout(n1477),.clk(gclk));
	jor g1177(.dina(n1477),.dinb(w_G523_0[1]),.dout(n1478),.clk(gclk));
	jand g1178(.dina(n1478),.dinb(n1474),.dout(n1479),.clk(gclk));
	jxor g1179(.dina(n1479),.dinb(n1470),.dout(n1480),.clk(gclk));
	jor g1180(.dina(w_n435_1[0]),.dinb(w_n369_1[0]),.dout(n1481),.clk(gclk));
	jor g1181(.dina(w_G324_0[2]),.dinb(w_n366_1[0]),.dout(n1482),.clk(gclk));
	jand g1182(.dina(n1482),.dinb(w_G503_0[2]),.dout(n1483),.clk(gclk));
	jand g1183(.dina(n1483),.dinb(w_dff_B_EY5P9kkJ0_1),.dout(n1484),.clk(gclk));
	jor g1184(.dina(w_G324_0[1]),.dinb(w_G254_1[0]),.dout(n1485),.clk(gclk));
	jor g1185(.dina(w_n435_0[2]),.dinb(w_G242_1[0]),.dout(n1486),.clk(gclk));
	jand g1186(.dina(n1486),.dinb(w_dff_B_4uGaUG2h6_1),.dout(n1487),.clk(gclk));
	jand g1187(.dina(n1487),.dinb(w_n437_0[0]),.dout(n1488),.clk(gclk));
	jor g1188(.dina(n1488),.dinb(n1484),.dout(n1489),.clk(gclk));
	jor g1189(.dina(w_G514_0[2]),.dinb(w_n408_3[2]),.dout(n1490),.clk(gclk));
	jor g1190(.dina(w_n361_0[0]),.dinb(w_G248_3[2]),.dout(n1491),.clk(gclk));
	jand g1191(.dina(n1491),.dinb(n1490),.dout(n1492),.clk(gclk));
	jxor g1192(.dina(n1492),.dinb(w_n371_0[0]),.dout(n1493),.clk(gclk));
	jxor g1193(.dina(w_dff_B_8Xf7QnmY4_0),.dinb(n1489),.dout(n1494),.clk(gclk));
	jxor g1194(.dina(n1494),.dinb(n1480),.dout(n1495),.clk(gclk));
	jxor g1195(.dina(w_n433_0[0]),.dinb(w_n428_0[1]),.dout(n1496),.clk(gclk));
	jxor g1196(.dina(w_n423_0[0]),.dinb(w_n412_0[0]),.dout(n1497),.clk(gclk));
	jxor g1197(.dina(n1497),.dinb(w_dff_B_vCCTPlxH9_1),.dout(n1498),.clk(gclk));
	jxor g1198(.dina(n1498),.dinb(n1495),.dout(n1499),.clk(gclk));
	jand g1199(.dina(n1499),.dinb(w_n749_5[0]),.dout(n1500),.clk(gclk));
	jnot g1200(.din(n1500),.dout(n1501),.clk(gclk));
	jand g1201(.dina(w_dff_B_LnFfZrMQ4_0),.dinb(n1461),.dout(n1502),.clk(gclk));
	jor g1202(.dina(n1502),.dinb(w_G4092_4[0]),.dout(n1503),.clk(gclk));
	jnot g1203(.din(w_n750_2[2]),.dout(n1504),.clk(gclk));
	jor g1204(.dina(w_n1504_0[1]),.dinb(w_dff_B_qS653Y2i8_1),.dout(n1505),.clk(gclk));
	jand g1205(.dina(w_dff_B_ow9X3H7R6_0),.dinb(w_n1503_0[1]),.dout(w_dff_A_EMPb80Xy4_2),.clk(gclk));
	jand g1206(.dina(w_G273_1[0]),.dinb(w_G248_3[1]),.dout(n1507),.clk(gclk));
	jand g1207(.dina(w_n471_0[2]),.dinb(w_G251_3[1]),.dout(n1508),.clk(gclk));
	jor g1208(.dina(n1508),.dinb(w_n473_1[0]),.dout(n1509),.clk(gclk));
	jor g1209(.dina(n1509),.dinb(w_dff_B_4fm55Zox3_1),.dout(n1510),.clk(gclk));
	jand g1210(.dina(w_n471_0[1]),.dinb(w_n406_3[1]),.dout(n1511),.clk(gclk));
	jand g1211(.dina(w_G273_0[2]),.dinb(w_n408_3[1]),.dout(n1512),.clk(gclk));
	jor g1212(.dina(n1512),.dinb(n1511),.dout(n1513),.clk(gclk));
	jor g1213(.dina(n1513),.dinb(w_G411_0[2]),.dout(n1514),.clk(gclk));
	jand g1214(.dina(n1514),.dinb(n1510),.dout(n1515),.clk(gclk));
	jand g1215(.dina(w_G281_1[0]),.dinb(w_G248_3[0]),.dout(n1516),.clk(gclk));
	jand g1216(.dina(w_n530_0[2]),.dinb(w_G251_3[0]),.dout(n1517),.clk(gclk));
	jor g1217(.dina(n1517),.dinb(w_n532_1[0]),.dout(n1518),.clk(gclk));
	jor g1218(.dina(n1518),.dinb(w_dff_B_o8C3BcRH5_1),.dout(n1519),.clk(gclk));
	jand g1219(.dina(w_n530_0[1]),.dinb(w_n406_3[0]),.dout(n1520),.clk(gclk));
	jand g1220(.dina(w_G281_0[2]),.dinb(w_n408_3[0]),.dout(n1521),.clk(gclk));
	jor g1221(.dina(n1521),.dinb(n1520),.dout(n1522),.clk(gclk));
	jor g1222(.dina(n1522),.dinb(w_G374_0[1]),.dout(n1523),.clk(gclk));
	jand g1223(.dina(n1523),.dinb(n1519),.dout(n1524),.clk(gclk));
	jxor g1224(.dina(n1524),.dinb(n1515),.dout(n1525),.clk(gclk));
	jor g1225(.dina(w_n483_1[0]),.dinb(w_n369_0[2]),.dout(n1526),.clk(gclk));
	jor g1226(.dina(w_G265_0[2]),.dinb(w_n366_0[2]),.dout(n1527),.clk(gclk));
	jand g1227(.dina(n1527),.dinb(w_G400_0[1]),.dout(n1528),.clk(gclk));
	jand g1228(.dina(n1528),.dinb(w_dff_B_ii3wpd5b0_1),.dout(n1529),.clk(gclk));
	jor g1229(.dina(w_G265_0[1]),.dinb(w_G254_0[2]),.dout(n1530),.clk(gclk));
	jor g1230(.dina(w_n483_0[2]),.dinb(w_G242_0[2]),.dout(n1531),.clk(gclk));
	jand g1231(.dina(n1531),.dinb(w_dff_B_vQWbygcP6_1),.dout(n1532),.clk(gclk));
	jand g1232(.dina(n1532),.dinb(w_n485_0[2]),.dout(n1533),.clk(gclk));
	jor g1233(.dina(n1533),.dinb(n1529),.dout(n1534),.clk(gclk));
	jand g1234(.dina(w_G257_1[0]),.dinb(w_G248_2[2]),.dout(n1535),.clk(gclk));
	jand g1235(.dina(w_n518_0[2]),.dinb(w_G251_2[2]),.dout(n1536),.clk(gclk));
	jor g1236(.dina(n1536),.dinb(w_n520_0[0]),.dout(n1537),.clk(gclk));
	jor g1237(.dina(n1537),.dinb(w_dff_B_GsQmPUvU2_1),.dout(n1538),.clk(gclk));
	jand g1238(.dina(w_n518_0[1]),.dinb(w_n406_2[2]),.dout(n1539),.clk(gclk));
	jand g1239(.dina(w_G257_0[2]),.dinb(w_n408_2[2]),.dout(n1540),.clk(gclk));
	jor g1240(.dina(n1540),.dinb(n1539),.dout(n1541),.clk(gclk));
	jor g1241(.dina(n1541),.dinb(w_G389_0[1]),.dout(n1542),.clk(gclk));
	jand g1242(.dina(n1542),.dinb(n1538),.dout(n1543),.clk(gclk));
	jand g1243(.dina(w_G248_2[1]),.dinb(w_G234_1[0]),.dout(n1544),.clk(gclk));
	jand g1244(.dina(w_G251_2[1]),.dinb(w_n460_0[2]),.dout(n1545),.clk(gclk));
	jor g1245(.dina(n1545),.dinb(w_n462_0[0]),.dout(n1546),.clk(gclk));
	jor g1246(.dina(n1546),.dinb(w_dff_B_SeD0dRPb3_1),.dout(n1547),.clk(gclk));
	jand g1247(.dina(w_n406_2[1]),.dinb(w_n460_0[1]),.dout(n1548),.clk(gclk));
	jand g1248(.dina(w_n408_2[1]),.dinb(w_G234_0[2]),.dout(n1549),.clk(gclk));
	jor g1249(.dina(n1549),.dinb(n1548),.dout(n1550),.clk(gclk));
	jor g1250(.dina(n1550),.dinb(w_G435_0[1]),.dout(n1551),.clk(gclk));
	jand g1251(.dina(n1551),.dinb(n1547),.dout(n1552),.clk(gclk));
	jxor g1252(.dina(n1552),.dinb(n1543),.dout(n1553),.clk(gclk));
	jxor g1253(.dina(n1553),.dinb(w_dff_B_wNMw5I5N0_1),.dout(n1554),.clk(gclk));
	jxor g1254(.dina(n1554),.dinb(w_dff_B_UhzF9ryi3_1),.dout(n1555),.clk(gclk));
	jand g1255(.dina(w_G248_2[0]),.dinb(w_G226_1[0]),.dout(n1556),.clk(gclk));
	jand g1256(.dina(w_G251_2[0]),.dinb(w_n494_0[2]),.dout(n1557),.clk(gclk));
	jor g1257(.dina(n1557),.dinb(w_n496_0[1]),.dout(n1558),.clk(gclk));
	jor g1258(.dina(n1558),.dinb(w_dff_B_2GqOtywX5_1),.dout(n1559),.clk(gclk));
	jand g1259(.dina(w_n406_2[0]),.dinb(w_n494_0[1]),.dout(n1560),.clk(gclk));
	jand g1260(.dina(w_n408_2[0]),.dinb(w_G226_0[2]),.dout(n1561),.clk(gclk));
	jor g1261(.dina(n1561),.dinb(n1560),.dout(n1562),.clk(gclk));
	jor g1262(.dina(n1562),.dinb(w_G422_0[1]),.dout(n1563),.clk(gclk));
	jand g1263(.dina(n1563),.dinb(n1559),.dout(n1564),.clk(gclk));
	jxor g1264(.dina(n1564),.dinb(w_n551_0[0]),.dout(n1565),.clk(gclk));
	jor g1265(.dina(w_n369_0[1]),.dinb(w_n507_0[2]),.dout(n1566),.clk(gclk));
	jor g1266(.dina(w_n366_0[1]),.dinb(w_G218_1[0]),.dout(n1567),.clk(gclk));
	jand g1267(.dina(n1567),.dinb(w_G468_0[1]),.dout(n1568),.clk(gclk));
	jand g1268(.dina(n1568),.dinb(w_dff_B_d0nm04rx4_1),.dout(n1569),.clk(gclk));
	jor g1269(.dina(w_G254_0[1]),.dinb(w_G218_0[2]),.dout(n1570),.clk(gclk));
	jor g1270(.dina(w_G242_0[1]),.dinb(w_n507_0[1]),.dout(n1571),.clk(gclk));
	jand g1271(.dina(n1571),.dinb(w_dff_B_wX4VpuQn3_1),.dout(n1572),.clk(gclk));
	jand g1272(.dina(n1572),.dinb(w_n509_0[0]),.dout(n1573),.clk(gclk));
	jor g1273(.dina(n1573),.dinb(n1569),.dout(n1574),.clk(gclk));
	jand g1274(.dina(w_G248_1[2]),.dinb(w_G210_1[0]),.dout(n1575),.clk(gclk));
	jand g1275(.dina(w_G251_1[2]),.dinb(w_n449_0[2]),.dout(n1576),.clk(gclk));
	jor g1276(.dina(n1576),.dinb(w_n451_0[0]),.dout(n1577),.clk(gclk));
	jor g1277(.dina(n1577),.dinb(w_dff_B_EtmbtrLr8_1),.dout(n1578),.clk(gclk));
	jand g1278(.dina(w_n406_1[2]),.dinb(w_n449_0[1]),.dout(n1579),.clk(gclk));
	jand g1279(.dina(w_n408_1[2]),.dinb(w_G210_0[2]),.dout(n1580),.clk(gclk));
	jor g1280(.dina(n1580),.dinb(n1579),.dout(n1581),.clk(gclk));
	jor g1281(.dina(n1581),.dinb(w_G457_0[1]),.dout(n1582),.clk(gclk));
	jand g1282(.dina(n1582),.dinb(n1578),.dout(n1583),.clk(gclk));
	jxor g1283(.dina(n1583),.dinb(n1574),.dout(n1584),.clk(gclk));
	jxor g1284(.dina(n1584),.dinb(n1565),.dout(n1585),.clk(gclk));
	jxor g1285(.dina(w_dff_B_889MNSiZ3_0),.dinb(n1555),.dout(n1586),.clk(gclk));
	jand g1286(.dina(n1586),.dinb(w_n749_4[2]),.dout(n1587),.clk(gclk));
	jnot g1287(.din(n1587),.dout(n1588),.clk(gclk));
	jand g1288(.dina(w_n573_0[0]),.dinb(w_n567_0[0]),.dout(n1589),.clk(gclk));
	jor g1289(.dina(w_dff_B_NbMeyCxI1_0),.dinb(w_n699_0[0]),.dout(n1590),.clk(gclk));
	jnot g1290(.din(w_n559_0[0]),.dout(n1591),.clk(gclk));
	jor g1291(.dina(n1591),.dinb(w_n557_0[0]),.dout(n1592),.clk(gclk));
	jand g1292(.dina(w_n1592_0[1]),.dinb(w_n532_0[2]),.dout(n1593),.clk(gclk));
	jnot g1293(.din(w_n1593_0[1]),.dout(n1594),.clk(gclk));
	jor g1294(.dina(w_n695_0[0]),.dinb(n1594),.dout(n1595),.clk(gclk));
	jand g1295(.dina(w_n923_0[1]),.dinb(w_n473_0[2]),.dout(n1596),.clk(gclk));
	jor g1296(.dina(w_n1596_0[1]),.dinb(w_n1593_0[0]),.dout(n1597),.clk(gclk));
	jand g1297(.dina(w_dff_B_xzfxRi8R7_0),.dinb(n1595),.dout(n1598),.clk(gclk));
	jxor g1298(.dina(w_dff_B_UZ0RO1iU3_0),.dinb(n1590),.dout(n1599),.clk(gclk));
	jnot g1299(.din(w_n1599_0[1]),.dout(n1600),.clk(gclk));
	jnot g1300(.din(w_n686_0[0]),.dout(n1601),.clk(gclk));
	jnot g1301(.din(w_n687_0[0]),.dout(n1602),.clk(gclk));
	jor g1302(.dina(w_n1592_0[0]),.dinb(w_n532_0[1]),.dout(n1603),.clk(gclk));
	jor g1303(.dina(w_n1596_0[0]),.dinb(w_n1603_0[1]),.dout(n1604),.clk(gclk));
	jor g1304(.dina(w_n923_0[0]),.dinb(w_n473_0[1]),.dout(n1605),.clk(gclk));
	jor g1305(.dina(w_n689_0[0]),.dinb(w_n485_0[1]),.dout(n1606),.clk(gclk));
	jand g1306(.dina(n1606),.dinb(w_n1605_0[1]),.dout(n1607),.clk(gclk));
	jand g1307(.dina(n1607),.dinb(n1604),.dout(n1608),.clk(gclk));
	jor g1308(.dina(n1608),.dinb(w_n690_0[0]),.dout(n1609),.clk(gclk));
	jor g1309(.dina(w_n1609_0[1]),.dinb(w_dff_B_RS5LCjhX5_1),.dout(n1610),.clk(gclk));
	jand g1310(.dina(n1610),.dinb(w_dff_B_xDHxEj471_1),.dout(n1611),.clk(gclk));
	jand g1311(.dina(w_n1611_0[2]),.dinb(w_n581_0[0]),.dout(n1612),.clk(gclk));
	jxor g1312(.dina(w_n566_0[0]),.dinb(w_n561_0[1]),.dout(n1613),.clk(gclk));
	jxor g1313(.dina(w_n1613_0[1]),.dinb(w_n865_0[1]),.dout(n1614),.clk(gclk));
	jxor g1314(.dina(w_dff_B_KEuu4M2p9_0),.dinb(n1612),.dout(n1615),.clk(gclk));
	jnot g1315(.din(w_n1615_0[1]),.dout(n1616),.clk(gclk));
	jand g1316(.dina(n1616),.dinb(w_dff_B_2bHVAlJb1_1),.dout(n1617),.clk(gclk));
	jnot g1317(.din(w_G1497_0[2]),.dout(n1618),.clk(gclk));
	jand g1318(.dina(w_n1615_0[0]),.dinb(w_n1599_0[0]),.dout(n1619),.clk(gclk));
	jor g1319(.dina(n1619),.dinb(w_n1618_0[1]),.dout(n1620),.clk(gclk));
	jor g1320(.dina(n1620),.dinb(n1617),.dout(n1621),.clk(gclk));
	jand g1321(.dina(w_n1605_0[0]),.dinb(w_n1603_0[0]),.dout(n1622),.clk(gclk));
	jor g1322(.dina(n1622),.dinb(w_n694_0[0]),.dout(n1623),.clk(gclk));
	jxor g1323(.dina(w_n1613_0[0]),.dinb(w_n1609_0[0]),.dout(n1624),.clk(gclk));
	jxor g1324(.dina(n1624),.dinb(w_dff_B_4grUwu5F0_1),.dout(n1625),.clk(gclk));
	jxor g1325(.dina(w_n1611_0[1]),.dinb(w_n865_0[0]),.dout(n1626),.clk(gclk));
	jxor g1326(.dina(n1626),.dinb(w_dff_B_NmUcLTXn0_1),.dout(n1627),.clk(gclk));
	jor g1327(.dina(n1627),.dinb(w_G1497_0[1]),.dout(n1628),.clk(gclk));
	jand g1328(.dina(w_dff_B_6bkGyK2w7_0),.dinb(n1621),.dout(n1629),.clk(gclk));
	jxor g1329(.dina(w_n579_0[1]),.dinb(w_n574_0[0]),.dout(n1630),.clk(gclk));
	jxor g1330(.dina(w_dff_B_kmufscFm5_0),.dinb(n1629),.dout(n1631),.clk(gclk));
	jnot g1331(.din(w_n709_0[0]),.dout(n1632),.clk(gclk));
	jand g1332(.dina(n1632),.dinb(w_n953_0[0]),.dout(n1633),.clk(gclk));
	jand g1333(.dina(w_n711_0[0]),.dinb(w_n954_0[1]),.dout(n1634),.clk(gclk));
	jor g1334(.dina(n1634),.dinb(w_n1633_0[1]),.dout(n1635),.clk(gclk));
	jxor g1335(.dina(w_n608_0[0]),.dinb(w_n592_0[0]),.dout(n1636),.clk(gclk));
	jxor g1336(.dina(n1636),.dinb(w_n602_0[0]),.dout(n1637),.clk(gclk));
	jxor g1337(.dina(w_n1637_0[1]),.dinb(n1635),.dout(n1638),.clk(gclk));
	jor g1338(.dina(w_n938_0[1]),.dinb(w_n597_0[0]),.dout(n1639),.clk(gclk));
	jand g1339(.dina(w_n609_0[0]),.dinb(w_n962_0[0]),.dout(n1640),.clk(gclk));
	jor g1340(.dina(w_dff_B_T8eDJLQt1_0),.dinb(w_n715_0[0]),.dout(n1641),.clk(gclk));
	jand g1341(.dina(w_dff_B_u1f4EHL35_0),.dinb(n1639),.dout(n1642),.clk(gclk));
	jxor g1342(.dina(n1642),.dinb(w_dff_B_KfVMJ9oW4_1),.dout(n1643),.clk(gclk));
	jand g1343(.dina(w_n1643_0[1]),.dinb(w_n703_0[1]),.dout(n1644),.clk(gclk));
	jnot g1344(.din(w_n682_0[0]),.dout(n1645),.clk(gclk));
	jor g1345(.dina(w_n1611_0[0]),.dinb(w_n684_0[0]),.dout(n1646),.clk(gclk));
	jand g1346(.dina(n1646),.dinb(w_dff_B_8cdrglPg3_1),.dout(n1647),.clk(gclk));
	jand g1347(.dina(w_n713_0[0]),.dinb(w_n954_0[0]),.dout(n1648),.clk(gclk));
	jor g1348(.dina(n1648),.dinb(w_n1633_0[0]),.dout(n1649),.clk(gclk));
	jxor g1349(.dina(w_dff_B_QoTvP5CI6_0),.dinb(w_n938_0[0]),.dout(n1650),.clk(gclk));
	jxor g1350(.dina(n1650),.dinb(w_n1637_0[0]),.dout(n1651),.clk(gclk));
	jand g1351(.dina(n1651),.dinb(n1647),.dout(n1652),.clk(gclk));
	jor g1352(.dina(w_n1652_0[1]),.dinb(n1644),.dout(n1653),.clk(gclk));
	jor g1353(.dina(n1653),.dinb(w_G1497_0[0]),.dout(n1654),.clk(gclk));
	jnot g1354(.din(w_n588_1[0]),.dout(n1655),.clk(gclk));
	jand g1355(.dina(w_n1652_0[0]),.dinb(w_dff_B_Nb21UJTq6_1),.dout(n1656),.clk(gclk));
	jor g1356(.dina(w_n703_0[0]),.dinb(w_n588_0[2]),.dout(n1657),.clk(gclk));
	jand g1357(.dina(n1657),.dinb(w_n1643_0[0]),.dout(n1658),.clk(gclk));
	jor g1358(.dina(n1658),.dinb(n1656),.dout(n1659),.clk(gclk));
	jor g1359(.dina(n1659),.dinb(w_n1618_0[0]),.dout(n1660),.clk(gclk));
	jand g1360(.dina(n1660),.dinb(n1654),.dout(n1661),.clk(gclk));
	jxor g1361(.dina(n1661),.dinb(n1631),.dout(n1662),.clk(gclk));
	jor g1362(.dina(n1662),.dinb(w_n749_4[1]),.dout(n1663),.clk(gclk));
	jand g1363(.dina(n1663),.dinb(w_dff_B_1X3yTzcg9_1),.dout(n1664),.clk(gclk));
	jor g1364(.dina(n1664),.dinb(w_G4092_3[2]),.dout(n1665),.clk(gclk));
	jor g1365(.dina(w_n1504_0[0]),.dinb(w_dff_B_E0dWacZS0_1),.dout(n1666),.clk(gclk));
	jand g1366(.dina(w_dff_B_9NRyjmDE9_0),.dinb(w_n1665_0[1]),.dout(w_dff_A_d5yH2TQb2_2),.clk(gclk));
	jor g1367(.dina(w_G4088_3[1]),.dinb(w_G14_0[1]),.dout(n1668),.clk(gclk));
	jor g1368(.dina(w_n797_3[1]),.dinb(w_G64_0[1]),.dout(n1669),.clk(gclk));
	jand g1369(.dina(n1669),.dinb(w_G4087_1[1]),.dout(n1670),.clk(gclk));
	jand g1370(.dina(n1670),.dinb(w_dff_B_F1BdJIRn7_1),.dout(n1671),.clk(gclk));
	jand g1371(.dina(w_G4092_3[1]),.dinb(G97),.dout(n1672),.clk(gclk));
	jnot g1372(.din(n1672),.dout(n1673),.clk(gclk));
	jand g1373(.dina(w_dff_B_UAoLTV0I0_0),.dinb(w_n1665_0[0]),.dout(n1674),.clk(gclk));
	jnot g1374(.din(w_n1674_0[2]),.dout(n1675),.clk(gclk));
	jor g1375(.dina(w_n1675_0[1]),.dinb(w_n797_3[0]),.dout(n1676),.clk(gclk));
	jand g1376(.dina(w_G4092_3[0]),.dinb(G94),.dout(n1677),.clk(gclk));
	jnot g1377(.din(n1677),.dout(n1678),.clk(gclk));
	jand g1378(.dina(w_dff_B_tshotWrx4_0),.dinb(w_n1503_0[0]),.dout(n1679),.clk(gclk));
	jnot g1379(.din(w_n1679_0[2]),.dout(n1680),.clk(gclk));
	jor g1380(.dina(w_n1680_0[1]),.dinb(w_G4088_3[0]),.dout(n1681),.clk(gclk));
	jand g1381(.dina(n1681),.dinb(w_n800_1[1]),.dout(n1682),.clk(gclk));
	jand g1382(.dina(n1682),.dinb(w_dff_B_Xab86eH79_1),.dout(n1683),.clk(gclk));
	jor g1383(.dina(n1683),.dinb(w_dff_B_DQdEZMtx8_1),.dout(w_dff_A_uayLeJHg8_2),.clk(gclk));
	jor g1384(.dina(w_G4089_3[1]),.dinb(w_G14_0[0]),.dout(n1685),.clk(gclk));
	jor g1385(.dina(w_n852_3[1]),.dinb(w_G64_0[0]),.dout(n1686),.clk(gclk));
	jand g1386(.dina(n1686),.dinb(w_G4090_1[1]),.dout(n1687),.clk(gclk));
	jand g1387(.dina(n1687),.dinb(w_dff_B_zD5UW9OE9_1),.dout(n1688),.clk(gclk));
	jor g1388(.dina(w_n1675_0[0]),.dinb(w_n852_3[0]),.dout(n1689),.clk(gclk));
	jor g1389(.dina(w_n1680_0[0]),.dinb(w_G4089_3[0]),.dout(n1690),.clk(gclk));
	jand g1390(.dina(n1690),.dinb(w_n854_1[1]),.dout(n1691),.clk(gclk));
	jand g1391(.dina(n1691),.dinb(w_dff_B_4w8ijg4L1_1),.dout(n1692),.clk(gclk));
	jor g1392(.dina(n1692),.dinb(w_dff_B_JZhC67786_1),.dout(w_dff_A_Y9j4iuZu8_2),.clk(gclk));
	jnot g1393(.din(w_G137_3[1]),.dout(n1694),.clk(gclk));
	jnot g1394(.din(G179),.dout(n1695),.clk(gclk));
	jnot g1395(.din(w_n996_1[1]),.dout(n1696),.clk(gclk));
	jor g1396(.dina(n1696),.dinb(w_n1695_0[1]),.dout(n1697),.clk(gclk));
	jnot g1397(.din(G176),.dout(n1698),.clk(gclk));
	jnot g1398(.din(w_n994_1[1]),.dout(n1699),.clk(gclk));
	jor g1399(.dina(n1699),.dinb(w_n1698_0[1]),.dout(n1700),.clk(gclk));
	jand g1400(.dina(w_n1674_0[1]),.dinb(w_G1689_1[2]),.dout(n1701),.clk(gclk));
	jand g1401(.dina(w_n1679_0[1]),.dinb(w_n993_1[1]),.dout(n1702),.clk(gclk));
	jor g1402(.dina(n1702),.dinb(w_G1690_0[1]),.dout(n1703),.clk(gclk));
	jor g1403(.dina(n1703),.dinb(w_dff_B_yScOK9ru2_1),.dout(n1704),.clk(gclk));
	jand g1404(.dina(n1704),.dinb(w_dff_B_2cHRsFbU8_1),.dout(n1705),.clk(gclk));
	jand g1405(.dina(n1705),.dinb(w_dff_B_OFoLb81D1_1),.dout(n1706),.clk(gclk));
	jor g1406(.dina(n1706),.dinb(w_n1694_0[1]),.dout(G658),.clk(gclk));
	jnot g1407(.din(w_n1012_1[1]),.dout(n1708),.clk(gclk));
	jor g1408(.dina(n1708),.dinb(w_n1695_0[0]),.dout(n1709),.clk(gclk));
	jnot g1409(.din(w_n1014_1[1]),.dout(n1710),.clk(gclk));
	jor g1410(.dina(n1710),.dinb(w_n1698_0[0]),.dout(n1711),.clk(gclk));
	jand g1411(.dina(w_n1674_0[0]),.dinb(w_G1691_1[2]),.dout(n1712),.clk(gclk));
	jand g1412(.dina(w_n1679_0[0]),.dinb(w_n1008_1[1]),.dout(n1713),.clk(gclk));
	jor g1413(.dina(n1713),.dinb(w_G1694_0[1]),.dout(n1714),.clk(gclk));
	jor g1414(.dina(n1714),.dinb(w_dff_B_TvwtaERu1_1),.dout(n1715),.clk(gclk));
	jand g1415(.dina(n1715),.dinb(w_dff_B_lPnA7KxI1_1),.dout(n1716),.clk(gclk));
	jand g1416(.dina(n1716),.dinb(w_dff_B_4pl9l5DJ3_1),.dout(n1717),.clk(gclk));
	jor g1417(.dina(n1717),.dinb(w_n1694_0[0]),.dout(G690),.clk(gclk));
	jdff g1418(.din(w_G141_1[0]),.dout(w_dff_A_3qesbko21_1),.clk(gclk));
	jdff g1419(.din(w_G293_0[0]),.dout(w_dff_A_k5hS1sGE3_1),.clk(gclk));
	jdff g1420(.din(w_G3173_0[0]),.dout(w_dff_A_d6kwjLVZ0_1),.clk(gclk));
	jnot g1421(.din(w_G545_0[1]),.dout(w_dff_A_hsW6rtkC8_1),.clk(gclk));
	jnot g1422(.din(w_G545_0[0]),.dout(w_dff_A_PX3V940Q1_1),.clk(gclk));
	jdff g1423(.din(w_G137_3[0]),.dout(w_dff_A_tBsHYMsf0_1),.clk(gclk));
	jdff g1424(.din(w_G141_0[2]),.dout(w_dff_A_tPCLe9f04_1),.clk(gclk));
	jdff g1425(.din(w_G1_2[0]),.dout(w_dff_A_mnbyVjQA2_1),.clk(gclk));
	jdff g1426(.din(w_G549_0[1]),.dout(w_dff_A_HsXSJqmW2_1),.clk(gclk));
	jdff g1427(.din(w_G299_0[1]),.dout(w_dff_A_YrcMuZjh5_1),.clk(gclk));
	jnot g1428(.din(w_G549_0[0]),.dout(w_dff_A_i0f25SsS5_1),.clk(gclk));
	jdff g1429(.din(w_G1_1[2]),.dout(w_dff_A_jBXFRELh6_1),.clk(gclk));
	jdff g1430(.din(w_G1_1[1]),.dout(w_dff_A_AOkWbxaA9_1),.clk(gclk));
	jdff g1431(.din(w_G1_1[0]),.dout(w_dff_A_8UBzqmtz1_1),.clk(gclk));
	jdff g1432(.din(w_G1_0[2]),.dout(w_dff_A_SKPLdeyi8_1),.clk(gclk));
	jdff g1433(.din(w_G299_0[0]),.dout(w_dff_A_Femo9NLV5_1),.clk(gclk));
	jor g1434(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(w_dff_A_BaD8i8TF9_2),.clk(gclk));
	jand g1435(.dina(w_n661_0[0]),.dinb(w_n641_0[1]),.dout(w_dff_A_VyRNnbsR6_2),.clk(gclk));
	jand g1436(.dina(w_n611_0[0]),.dinb(w_n588_0[1]),.dout(w_dff_A_RZ4RQ0L23_2),.clk(gclk));
	jor g1437(.dina(w_n717_0[0]),.dinb(w_n704_0[0]),.dout(w_dff_A_B0akqYdF7_2),.clk(gclk));
	jor g1438(.dina(w_n747_0[0]),.dinb(w_n738_0[0]),.dout(w_dff_A_Znsu090U2_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_dff_A_zhbpJqqR3_1),.doutc(w_G4_0[2]),.din(w_dff_B_3BFNaT9z0_3));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(G11));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(G14));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(w_dff_B_RPIWd08X5_2));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(w_dff_B_MZAmZeka7_2));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(w_dff_B_h9kxZlyU6_2));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(w_dff_B_YnmLANBf9_2));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(G43));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(G46));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(w_dff_B_QHr4jZ8J4_2));
	jspl3 jspl3_w_G54_0(.douta(w_dff_A_IjOfffxg2_0),.doutb(w_dff_A_w3gOLomI2_1),.doutc(w_G54_0[2]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(w_dff_B_5Pi8sLZf6_2));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(w_dff_B_YuQ5o83W9_2));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(G67));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(w_dff_B_FIoheWbs5_2));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(G73));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(G76));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(G91));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(G100));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(w_dff_B_uaO0d8MK4_2));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(w_dff_B_ysMN1GsA7_2));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(G109));
	jspl jspl_w_G123_0(.douta(w_dff_A_bJ19DS6e9_0),.doutb(w_G123_0[1]),.din(G123));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_yOntMPx73_0),.doutb(w_dff_A_fEh8IIwQ7_1),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_9SF0wWVx1_0),.doutb(w_dff_A_z3v7vRp71_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_vfZVX75W4_0),.doutb(w_dff_A_Jw5QYtyr4_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_dff_A_tdkmqNYI7_2),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_dff_A_kCA1roIz8_0),.doutb(w_dff_A_Ii9nEp3G4_1),.doutc(w_G137_4[2]),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_dff_A_0vW8M7pl8_0),.doutb(w_G137_5[1]),.doutc(w_G137_5[2]),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_wEzRSUOx8_0),.doutb(w_dff_A_9uvh0oUf1_1),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_gGGJZbzA5_1),.doutc(w_dff_A_GGM1gy4q7_2),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_G137_8[0]),.doutb(w_G137_8[1]),.doutc(w_dff_A_snODAuqc6_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_G137_9[0]),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_TU9gGnzH5_1),.doutc(w_dff_A_edFeGmke8_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_G139qUXC6_0),.doutb(w_dff_A_9pMjfsWj9_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(w_dff_B_ZI5yvDHv8_2));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(w_dff_B_t5CF08rg6_2));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(w_dff_B_8AGxI0Mu5_2));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(w_dff_B_Ajmd820Z0_2));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(w_dff_B_SJjDmDZT6_2));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(w_dff_B_ZoSLA8cb9_2));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(w_dff_B_shkYsADX0_2));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(w_dff_B_NwUqWdPU1_2));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(w_dff_B_o2AF7ZD13_2));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(w_dff_B_hv1i2ayl9_2));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(w_dff_B_UXYvnfD98_2));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(w_dff_B_cX4vbk7M7_2));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(w_dff_B_K9zwZyi23_2));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(w_dff_B_fGuvLndO3_2));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(w_dff_B_GHXBL6V70_2));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(w_dff_B_6Z1okz4h3_2));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(w_dff_B_O2epEFNI8_2));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(w_dff_B_PZmhi2Ux9_2));
	jspl3 jspl3_w_G206_0(.douta(w_G206_0[0]),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G206_1(.douta(w_dff_A_5HCCnfVr4_0),.doutb(w_G206_1[1]),.doutc(w_G206_1[2]),.din(w_G206_0[0]));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_dff_A_ObGN1cyK6_2),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_G210_1[1]),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl jspl_w_G210_2(.douta(w_dff_A_oLekoJB74_0),.doutb(w_G210_2[1]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_dff_A_omqAYVWi0_0),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl jspl_w_G218_2(.douta(w_dff_A_GfG3u0CN9_0),.doutb(w_G218_2[1]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_dff_A_gT9buK4T4_2),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_G226_1[0]),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl jspl_w_G226_2(.douta(w_dff_A_jKyEDYcW2_0),.doutb(w_G226_2[1]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_dff_A_zJ4OzjGQ4_2),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_dff_A_IAv7bVlJ3_0),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_dff_A_vXPYLiIZ1_1),.doutc(w_dff_A_zeUXuxX64_2),.din(G242));
	jspl jspl_w_G242_1(.douta(w_dff_A_ObhXBezk2_0),.doutb(w_G242_1[1]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_dff_A_lTOzkCx56_0),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_dff_A_OfhDr8Jr0_2),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl3 jspl3_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.doutc(w_G248_5[2]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_dff_A_h7Jd0gJN0_1),.doutc(w_dff_A_DQGrjRHK8_2),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_dff_A_iW6HyRsz8_0),.doutb(w_G251_1[1]),.doutc(w_dff_A_3HPeGmjr0_2),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_G251_4[1]),.doutc(w_G251_4[2]),.din(w_G251_1[0]));
	jspl jspl_w_G251_5(.douta(w_dff_A_J1GBjRnw5_0),.doutb(w_G251_5[1]),.din(w_G251_1[1]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl jspl_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_dff_A_CID2Snx76_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_G257_1[0]),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl jspl_w_G257_2(.douta(w_dff_A_jWHGvtCa9_0),.doutb(w_G257_2[1]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_dff_A_c5SsxF4r5_2),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_dff_A_yKhhrmpy2_1),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_dff_A_4imqgMe79_2),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_dff_A_AK5xYz0k8_1),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl jspl_w_G273_2(.douta(w_dff_A_CCG8Zxt41_0),.doutb(w_G273_2[1]),.din(w_G273_0[1]));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_dff_A_YoDwKxKM6_2),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_dff_A_YLF0ccXX5_0),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_G289_0[0]),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_dff_A_ohMqcqoZ8_1),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_dff_A_etQq017Q2_0),.doutb(w_dff_A_kGtQubRU4_1),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_dff_A_ScLRp0dH0_0),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_dff_A_gRwoKJ1I1_2),.din(G316));
	jspl jspl_w_G316_1(.douta(w_G316_1[0]),.doutb(w_G316_1[1]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_G324_0[1]),.doutc(w_dff_A_zFfp6bVg0_2),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_dff_A_F8Uk3U9y7_1),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_dff_A_R1RIDmXh3_1),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_dff_A_FPSHAf153_1),.doutc(w_G332_1[2]),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_dff_A_ebIdPORu4_0),.doutb(w_G332_2[1]),.doutc(w_dff_A_5elyxUXx2_2),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_G332_3[0]),.doutb(w_G332_3[1]),.doutc(w_G332_3[2]),.din(w_G332_0[2]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl jspl_w_G338_0(.douta(w_dff_A_RfHlSoqf7_0),.doutb(w_G338_0[1]),.din(G338));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_dff_A_r9ppHhem0_2),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_dff_A_F6B7u8qa1_1),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_dff_A_hItFPknl1_0),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_dff_A_SNlAwwOi8_2),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_G351_1[0]),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_dff_A_ngYc9BaC7_1),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_dff_A_qeIdu1Xg2_0),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_G361_0[1]),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G361_1(.douta(w_dff_A_S8jCp1lV4_0),.doutb(w_G361_1[1]),.din(w_G361_0[0]));
	jspl jspl_w_G366_0(.douta(w_dff_A_MJ0ViibJ4_0),.doutb(w_G366_0[1]),.din(G366));
	jspl jspl_w_G369_0(.douta(w_G369_0[0]),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_G374_0[0]),.doutb(w_dff_A_MbOpF8PG8_1),.doutc(w_dff_A_5g6MpCxj4_2),.din(G374));
	jspl3 jspl3_w_G374_1(.douta(w_dff_A_oxlsLqtp8_0),.doutb(w_dff_A_pi6uTrMi7_1),.doutc(w_G374_1[2]),.din(w_G374_0[0]));
	jspl3 jspl3_w_G389_0(.douta(w_G389_0[0]),.doutb(w_dff_A_RU41QhYS4_1),.doutc(w_dff_A_A8WUKmeI4_2),.din(G389));
	jspl3 jspl3_w_G389_1(.douta(w_dff_A_SWo3DVyA2_0),.doutb(w_dff_A_VgDuH2sX9_1),.doutc(w_G389_1[2]),.din(w_G389_0[0]));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_dff_A_poS3m5Qm4_1),.doutc(w_dff_A_OVVhrC421_2),.din(G400));
	jspl3 jspl3_w_G400_1(.douta(w_dff_A_PRE9t4K11_0),.doutb(w_dff_A_BcsnzGcI1_1),.doutc(w_G400_1[2]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_dff_A_lge6Nse23_0),.doutb(w_G411_0[1]),.doutc(w_dff_A_HuQwAL7r3_2),.din(G411));
	jspl3 jspl3_w_G411_1(.douta(w_G411_1[0]),.doutb(w_G411_1[1]),.doutc(w_G411_1[2]),.din(w_G411_0[0]));
	jspl jspl_w_G411_2(.douta(w_dff_A_El7HS5tF9_0),.doutb(w_G411_2[1]),.din(w_G411_0[1]));
	jspl3 jspl3_w_G422_0(.douta(w_G422_0[0]),.doutb(w_dff_A_sS3oEy2s3_1),.doutc(w_dff_A_M0zNXlLG7_2),.din(G422));
	jspl jspl_w_G422_1(.douta(w_dff_A_byQV1EwN1_0),.doutb(w_G422_1[1]),.din(w_G422_0[0]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_dff_A_qaPcEWrT7_1),.doutc(w_dff_A_8lsHxblE7_2),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_dff_A_ZOupd35Q9_0),.doutb(w_dff_A_lrnp6gFq2_1),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_dff_A_ZxaHmWHq9_1),.doutc(w_dff_A_Mmgn51Xh7_2),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_dff_A_ofgL8hNt0_0),.doutb(w_dff_A_ClsEoZwW8_1),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_G457_0[0]),.doutb(w_dff_A_y63zbw8x4_1),.doutc(w_dff_A_SfgBxLJ12_2),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_dff_A_ofFN2KXF6_0),.doutb(w_dff_A_L5HpIfiT5_1),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_dff_A_Zllgn7rC3_1),.doutc(w_dff_A_C4MnImA90_2),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_dff_A_A5Y9CIJd1_0),.doutb(w_dff_A_UmtnvGTW6_1),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_dff_A_U2B1WQkS2_0),.doutb(w_dff_A_EbD5XZ6A1_1),.doutc(w_G479_0[2]),.din(G479));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_dff_A_S77Krj036_1),.doutc(w_dff_A_lcGgPAjg9_2),.din(G490));
	jspl jspl_w_G490_1(.douta(w_dff_A_DlOB61Du6_0),.doutb(w_G490_1[1]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_dff_A_GN83aTc42_0),.doutb(w_G503_0[1]),.doutc(w_dff_A_NJpbWQ6H2_2),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_G503_1[0]),.doutb(w_G503_1[1]),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl jspl_w_G503_2(.douta(w_dff_A_PXTYXeMl1_0),.doutb(w_G503_2[1]),.din(w_G503_0[1]));
	jspl3 jspl3_w_G514_0(.douta(w_dff_A_3n8RWLgq4_0),.doutb(w_G514_0[1]),.doutc(w_dff_A_khKlBzin5_2),.din(G514));
	jspl3 jspl3_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.doutc(w_G514_1[2]),.din(w_G514_0[0]));
	jspl jspl_w_G514_2(.douta(w_G514_2[0]),.doutb(w_G514_2[1]),.din(w_G514_0[1]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_dff_A_w06BWhO72_1),.doutc(w_dff_A_jo6hae3s0_2),.din(G523));
	jspl3 jspl3_w_G523_1(.douta(w_dff_A_RzdvU1OF3_0),.doutb(w_dff_A_5oDTPYdf1_1),.doutc(w_G523_1[2]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_dff_A_LAEMmbVG5_0),.doutb(w_G534_0[1]),.doutc(w_dff_A_uz8yns7j3_2),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_G534_1[0]),.doutb(w_G534_1[1]),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl jspl_w_G534_2(.douta(w_dff_A_YeTVb28I2_0),.doutb(w_G534_2[1]),.din(w_G534_0[1]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_dff_A_FtQ5RHRX1_0),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_dff_A_USsYQNdK9_0),.doutb(w_dff_A_fKRahply6_1),.doutc(w_G1497_0[2]),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_dff_A_TRFWSf9o9_1),.doutc(w_dff_A_qhYXJhut8_2),.din(G1689));
	jspl3 jspl3_w_G1689_1(.douta(w_dff_A_DjEPVuot6_0),.doutb(w_G1689_1[1]),.doutc(w_dff_A_V9AeNPX94_2),.din(w_G1689_0[0]));
	jspl3 jspl3_w_G1689_2(.douta(w_dff_A_HFPQpTJG5_0),.doutb(w_G1689_2[1]),.doutc(w_dff_A_ppmNuYTf8_2),.din(w_G1689_0[1]));
	jspl3 jspl3_w_G1689_3(.douta(w_dff_A_wAZAh3OW7_0),.doutb(w_dff_A_IdOvsTrc2_1),.doutc(w_G1689_3[2]),.din(w_G1689_0[2]));
	jspl3 jspl3_w_G1689_4(.douta(w_dff_A_BNuCiqWE6_0),.doutb(w_dff_A_NmeBqJej4_1),.doutc(w_G1689_4[2]),.din(w_G1689_1[0]));
	jspl jspl_w_G1689_5(.douta(w_G1689_5[0]),.doutb(w_G1689_5[1]),.din(w_G1689_1[1]));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_dff_A_8q1v2Fau8_1),.doutc(w_G1690_0[2]),.din(G1690));
	jspl jspl_w_G1690_1(.douta(w_G1690_1[0]),.doutb(w_dff_A_oQ6hWZ8K6_1),.din(w_G1690_0[0]));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_dff_A_6aehFRuv9_1),.doutc(w_dff_A_vGHTfhyW9_2),.din(G1691));
	jspl3 jspl3_w_G1691_1(.douta(w_G1691_1[0]),.doutb(w_G1691_1[1]),.doutc(w_dff_A_DEUdClEX8_2),.din(w_G1691_0[0]));
	jspl3 jspl3_w_G1691_2(.douta(w_dff_A_phMaxgek3_0),.doutb(w_G1691_2[1]),.doutc(w_dff_A_4i0Tqhj48_2),.din(w_G1691_0[1]));
	jspl3 jspl3_w_G1691_3(.douta(w_dff_A_PTfTAvJb1_0),.doutb(w_dff_A_vpSkG3G47_1),.doutc(w_G1691_3[2]),.din(w_G1691_0[2]));
	jspl3 jspl3_w_G1691_4(.douta(w_dff_A_eNq6EuQo6_0),.doutb(w_dff_A_XLZ3R2fU3_1),.doutc(w_G1691_4[2]),.din(w_G1691_1[0]));
	jspl jspl_w_G1691_5(.douta(w_G1691_5[0]),.doutb(w_dff_A_KCA2LkGM5_1),.din(w_G1691_1[1]));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_dff_A_PuJrd79y3_1),.doutc(w_dff_A_dgGMwTgw5_2),.din(G1694));
	jspl jspl_w_G1694_1(.douta(w_G1694_1[0]),.doutb(w_G1694_1[1]),.din(w_G1694_0[0]));
	jspl3 jspl3_w_G2174_0(.douta(w_dff_A_Jsb5G67L3_0),.doutb(w_dff_A_ibm6KBV90_1),.doutc(w_G2174_0[2]),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_dff_A_5H7xdybX2_0),.doutb(w_dff_A_tmZmnfvl0_1),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(w_dff_B_q9Ly9YM44_3));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_dff_A_yY3htEE00_0),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_G3724_0[0]),.doutb(w_G3724_0[1]),.doutc(w_dff_A_nRGnI5Q08_2),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_dff_A_ZtjjC1cr6_1),.doutc(w_dff_A_yQpYbEpp5_2),.din(G4087));
	jspl3 jspl3_w_G4087_1(.douta(w_G4087_1[0]),.doutb(w_dff_A_qxidpLW09_1),.doutc(w_dff_A_EXoqS4CX2_2),.din(w_G4087_0[0]));
	jspl3 jspl3_w_G4087_2(.douta(w_G4087_2[0]),.doutb(w_G4087_2[1]),.doutc(w_G4087_2[2]),.din(w_G4087_0[1]));
	jspl3 jspl3_w_G4087_3(.douta(w_G4087_3[0]),.doutb(w_G4087_3[1]),.doutc(w_G4087_3[2]),.din(w_G4087_0[2]));
	jspl3 jspl3_w_G4087_4(.douta(w_dff_A_uKSr5MXa6_0),.doutb(w_dff_A_pPMSWfET9_1),.doutc(w_G4087_4[2]),.din(w_G4087_1[0]));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_G4088_0[2]),.din(G4088));
	jspl3 jspl3_w_G4088_1(.douta(w_G4088_1[0]),.doutb(w_G4088_1[1]),.doutc(w_G4088_1[2]),.din(w_G4088_0[0]));
	jspl3 jspl3_w_G4088_2(.douta(w_G4088_2[0]),.doutb(w_G4088_2[1]),.doutc(w_G4088_2[2]),.din(w_G4088_0[1]));
	jspl3 jspl3_w_G4088_3(.douta(w_dff_A_e2DMmeF93_0),.doutb(w_G4088_3[1]),.doutc(w_G4088_3[2]),.din(w_G4088_0[2]));
	jspl3 jspl3_w_G4088_4(.douta(w_dff_A_jVEqA2kz8_0),.doutb(w_G4088_4[1]),.doutc(w_dff_A_SBWxVdOH5_2),.din(w_G4088_1[0]));
	jspl3 jspl3_w_G4088_5(.douta(w_G4088_5[0]),.doutb(w_dff_A_cevV5e9A0_1),.doutc(w_G4088_5[2]),.din(w_G4088_1[1]));
	jspl3 jspl3_w_G4088_6(.douta(w_dff_A_UAnolVtf5_0),.doutb(w_G4088_6[1]),.doutc(w_dff_A_ycHHp8f25_2),.din(w_G4088_1[2]));
	jspl3 jspl3_w_G4088_7(.douta(w_G4088_7[0]),.doutb(w_dff_A_J40c4J9p9_1),.doutc(w_G4088_7[2]),.din(w_G4088_2[0]));
	jspl3 jspl3_w_G4088_8(.douta(w_dff_A_p986CboN5_0),.doutb(w_G4088_8[1]),.doutc(w_dff_A_FgbyN03F3_2),.din(w_G4088_2[1]));
	jspl3 jspl3_w_G4088_9(.douta(w_G4088_9[0]),.doutb(w_dff_A_F4a1JVaO5_1),.doutc(w_G4088_9[2]),.din(w_G4088_2[2]));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_G4089_0[2]),.din(G4089));
	jspl3 jspl3_w_G4089_1(.douta(w_G4089_1[0]),.doutb(w_G4089_1[1]),.doutc(w_G4089_1[2]),.din(w_G4089_0[0]));
	jspl3 jspl3_w_G4089_2(.douta(w_G4089_2[0]),.doutb(w_G4089_2[1]),.doutc(w_G4089_2[2]),.din(w_G4089_0[1]));
	jspl3 jspl3_w_G4089_3(.douta(w_dff_A_M6dwhNZe0_0),.doutb(w_G4089_3[1]),.doutc(w_G4089_3[2]),.din(w_G4089_0[2]));
	jspl3 jspl3_w_G4089_4(.douta(w_dff_A_Hzdn82JJ8_0),.doutb(w_G4089_4[1]),.doutc(w_dff_A_8Qwl9bBz2_2),.din(w_G4089_1[0]));
	jspl3 jspl3_w_G4089_5(.douta(w_G4089_5[0]),.doutb(w_dff_A_TBX5Mh469_1),.doutc(w_dff_A_RJWpgXXD6_2),.din(w_G4089_1[1]));
	jspl3 jspl3_w_G4089_6(.douta(w_G4089_6[0]),.doutb(w_G4089_6[1]),.doutc(w_dff_A_SuyHfsP33_2),.din(w_G4089_1[2]));
	jspl3 jspl3_w_G4089_7(.douta(w_dff_A_EGw3OCqi1_0),.doutb(w_G4089_7[1]),.doutc(w_dff_A_d2WmELSA3_2),.din(w_G4089_2[0]));
	jspl3 jspl3_w_G4089_8(.douta(w_G4089_8[0]),.doutb(w_dff_A_DGMxBQG38_1),.doutc(w_G4089_8[2]),.din(w_G4089_2[1]));
	jspl3 jspl3_w_G4089_9(.douta(w_G4089_9[0]),.doutb(w_dff_A_y6gLe14R0_1),.doutc(w_G4089_9[2]),.din(w_G4089_2[2]));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_dff_A_98uwd9An2_1),.doutc(w_dff_A_N5K4KyUj0_2),.din(G4090));
	jspl3 jspl3_w_G4090_1(.douta(w_G4090_1[0]),.doutb(w_dff_A_a1NFrYxL3_1),.doutc(w_dff_A_oHlGz0YR3_2),.din(w_G4090_0[0]));
	jspl3 jspl3_w_G4090_2(.douta(w_G4090_2[0]),.doutb(w_G4090_2[1]),.doutc(w_dff_A_RHULBzFo7_2),.din(w_G4090_0[1]));
	jspl3 jspl3_w_G4090_3(.douta(w_G4090_3[0]),.doutb(w_dff_A_YxLnYYPV2_1),.doutc(w_dff_A_wZ5mTor86_2),.din(w_G4090_0[2]));
	jspl3 jspl3_w_G4090_4(.douta(w_dff_A_ghHCOaPZ1_0),.doutb(w_dff_A_y0stXhZv5_1),.doutc(w_G4090_4[2]),.din(w_G4090_1[0]));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_dff_A_ZsiNco8d4_1),.doutc(w_dff_A_pFqduqXp0_2),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_dff_A_WS9eeEtU1_0),.doutb(w_dff_A_H1SsEM2h4_1),.doutc(w_G4091_1[2]),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_dff_A_EQO7aPUZ7_0),.doutb(w_dff_A_DB8a6sF52_1),.doutc(w_G4091_2[2]),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4091_3(.douta(w_G4091_3[0]),.doutb(w_dff_A_za0xKMAC7_1),.doutc(w_dff_A_Yv7YRBAz8_2),.din(w_G4091_0[2]));
	jspl3 jspl3_w_G4091_4(.douta(w_dff_A_vWLEkGRQ2_0),.doutb(w_G4091_4[1]),.doutc(w_dff_A_a58CEpQU8_2),.din(w_G4091_1[0]));
	jspl3 jspl3_w_G4091_5(.douta(w_dff_A_xhrFUx5g6_0),.doutb(w_G4091_5[1]),.doutc(w_dff_A_2hM6Ucfa7_2),.din(w_G4091_1[1]));
	jspl jspl_w_G4091_6(.douta(w_dff_A_piDFrEPc8_0),.doutb(w_G4091_6[1]),.din(w_G4091_1[2]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_dff_A_QPoL2Yr86_1),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_dff_A_xXFR20xn1_0),.doutb(w_G4092_1[1]),.doutc(w_dff_A_8AaK8aOG1_2),.din(w_G4092_0[0]));
	jspl3 jspl3_w_G4092_2(.douta(w_dff_A_Rcqv1pnE6_0),.doutb(w_dff_A_u4fEX5Gh2_1),.doutc(w_G4092_2[2]),.din(w_G4092_0[1]));
	jspl3 jspl3_w_G4092_3(.douta(w_G4092_3[0]),.doutb(w_G4092_3[1]),.doutc(w_dff_A_4gOJRDdD0_2),.din(w_G4092_0[2]));
	jspl3 jspl3_w_G4092_4(.douta(w_dff_A_opWE1Xsm3_0),.doutb(w_G4092_4[1]),.doutc(w_G4092_4[2]),.din(w_G4092_1[0]));
	jspl3 jspl3_w_G4092_5(.douta(w_dff_A_93243qg33_0),.doutb(w_dff_A_N2iAANj73_1),.doutc(w_G4092_5[2]),.din(w_G4092_1[1]));
	jspl3 jspl3_w_G4092_6(.douta(w_G4092_6[0]),.doutb(w_dff_A_rLeApYgQ2_1),.doutc(w_dff_A_Zoy8pnXB4_2),.din(w_G4092_1[2]));
	jspl3 jspl3_w_G4092_7(.douta(w_G4092_7[0]),.doutb(w_G4092_7[1]),.doutc(w_dff_A_QMPVijS82_2),.din(w_G4092_2[0]));
	jspl3 jspl3_w_G4092_8(.douta(w_G4092_8[0]),.doutb(w_dff_A_QegbFgMH0_1),.doutc(w_dff_A_fI6T211y3_2),.din(w_G4092_2[1]));
	jspl3 jspl3_w_G4092_9(.douta(w_dff_A_5lvsBwnu3_0),.doutb(w_dff_A_R2cCntsR9_1),.doutc(w_G4092_9[2]),.din(w_G4092_2[2]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(w_dff_A_2GuE02g96_1),.din(G599_fa_));
	jspl jspl_w_G601_0(.douta(w_G601_0),.doutb(w_dff_A_xSrgjd2r2_1),.din(G601_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(w_dff_A_ngtpAtsY5_1),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_G809_1[0]),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_G809_2[2]),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_G809_3[0]),.doutb(w_G809_3[1]),.doutc(w_dff_A_f2GSdHvr4_2),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(w_dff_A_JlUsfOTy7_1),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(w_dff_A_hgFfuhYA3_1),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(w_dff_A_9ExCEcXI6_1),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(w_dff_A_an0UBJ8I1_1),.din(G861_fa_));
	jspl jspl_w_G623_0(.douta(w_G623_0),.doutb(w_dff_A_J3A90Aak2_1),.din(G623_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(w_dff_A_lbSS0iQn2_1),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(w_dff_A_D28W5EYA0_1),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(w_dff_A_4PavxOpF1_1),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(w_dff_A_PwVeE3Jp6_1),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(w_dff_A_ORWvyfmF9_1),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(w_dff_A_lkGGGKZR7_1),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(w_dff_A_y5o85UER5_1),.din(G877_fa_));
	jspl jspl_w_G998_0(.douta(w_G998_0),.doutb(w_dff_A_32pOtW9D1_1),.din(G998_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(w_dff_A_lO1QpRnm5_1),.din(G830_fa_));
	jspl jspl_w_G865_0(.douta(w_G865_0),.doutb(w_dff_A_8HK7cpkl2_1),.din(G865_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(w_dff_A_YxXv40kT5_1),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(w_dff_B_m9fN94CJ9_2));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.doutc(w_n369_0[2]),.din(n369));
	jspl3 jspl3_w_n369_1(.douta(w_n369_1[0]),.doutb(w_n369_1[1]),.doutc(w_n369_1[2]),.din(w_n369_0[0]));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl3 jspl3_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.doutc(w_n374_0[2]),.din(n374));
	jspl jspl_w_n374_1(.douta(w_n374_1[0]),.doutb(w_n374_1[1]),.din(w_n374_0[0]));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl3 jspl3_w_n375_1(.douta(w_n375_1[0]),.doutb(w_n375_1[1]),.doutc(w_n375_1[2]),.din(w_n375_0[0]));
	jspl3 jspl3_w_n375_2(.douta(w_n375_2[0]),.doutb(w_n375_2[1]),.doutc(w_n375_2[2]),.din(w_n375_0[1]));
	jspl3 jspl3_w_n375_3(.douta(w_n375_3[0]),.doutb(w_n375_3[1]),.doutc(w_n375_3[2]),.din(w_n375_0[2]));
	jspl3 jspl3_w_n375_4(.douta(w_n375_4[0]),.doutb(w_n375_4[1]),.doutc(w_n375_4[2]),.din(w_n375_1[0]));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_dff_A_Gva3RcoY4_2),.din(w_dff_B_8YMo3sLn6_3));
	jspl jspl_w_n377_1(.douta(w_dff_A_iWDqtKCR1_0),.doutb(w_n377_1[1]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.doutc(w_n378_0[2]),.din(n378));
	jspl3 jspl3_w_n378_1(.douta(w_n378_1[0]),.doutb(w_n378_1[1]),.doutc(w_n378_1[2]),.din(w_n378_0[0]));
	jspl3 jspl3_w_n378_2(.douta(w_n378_2[0]),.doutb(w_n378_2[1]),.doutc(w_n378_2[2]),.din(w_n378_0[1]));
	jspl3 jspl3_w_n378_3(.douta(w_n378_3[0]),.doutb(w_n378_3[1]),.doutc(w_n378_3[2]),.din(w_n378_0[2]));
	jspl3 jspl3_w_n378_4(.douta(w_n378_4[0]),.doutb(w_n378_4[1]),.doutc(w_n378_4[2]),.din(w_n378_1[0]));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_dff_A_jcIciAi55_2),.din(w_dff_B_43Qwqhk89_3));
	jspl jspl_w_n389_1(.douta(w_dff_A_vNWGVL5O1_0),.doutb(w_n389_1[1]),.din(w_n389_0[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n401_0(.douta(w_dff_A_TG9rKCVs5_0),.doutb(w_n401_0[1]),.din(w_dff_B_dxrmcj3p8_2));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.doutc(w_n406_0[2]),.din(n406));
	jspl3 jspl3_w_n406_1(.douta(w_n406_1[0]),.doutb(w_n406_1[1]),.doutc(w_n406_1[2]),.din(w_n406_0[0]));
	jspl3 jspl3_w_n406_2(.douta(w_n406_2[0]),.doutb(w_n406_2[1]),.doutc(w_n406_2[2]),.din(w_n406_0[1]));
	jspl3 jspl3_w_n406_3(.douta(w_n406_3[0]),.doutb(w_n406_3[1]),.doutc(w_n406_3[2]),.din(w_n406_0[2]));
	jspl3 jspl3_w_n406_4(.douta(w_n406_4[0]),.doutb(w_n406_4[1]),.doutc(w_n406_4[2]),.din(w_n406_1[0]));
	jspl jspl_w_n406_5(.douta(w_n406_5[0]),.doutb(w_n406_5[1]),.din(w_n406_1[1]));
	jspl3 jspl3_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.doutc(w_n408_0[2]),.din(n408));
	jspl3 jspl3_w_n408_1(.douta(w_n408_1[0]),.doutb(w_n408_1[1]),.doutc(w_n408_1[2]),.din(w_n408_0[0]));
	jspl3 jspl3_w_n408_2(.douta(w_n408_2[0]),.doutb(w_n408_2[1]),.doutc(w_n408_2[2]),.din(w_n408_0[1]));
	jspl3 jspl3_w_n408_3(.douta(w_n408_3[0]),.doutb(w_n408_3[1]),.doutc(w_n408_3[2]),.din(w_n408_0[2]));
	jspl3 jspl3_w_n408_4(.douta(w_n408_4[0]),.doutb(w_n408_4[1]),.doutc(w_n408_4[2]),.din(w_n408_1[0]));
	jspl3 jspl3_w_n408_5(.douta(w_n408_5[0]),.doutb(w_n408_5[1]),.doutc(w_n408_5[2]),.din(w_n408_1[1]));
	jspl3 jspl3_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.doutc(w_n412_0[2]),.din(n412));
	jspl jspl_w_n414_0(.douta(w_dff_A_f4tHy0gm6_0),.doutb(w_n414_0[1]),.din(w_dff_B_zrNIoY7t3_2));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl3 jspl3_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.doutc(w_n423_0[2]),.din(n423));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_n425_0[2]),.din(n425));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_dff_A_ZpN0xOKU4_1),.doutc(w_n428_0[2]),.din(n428));
	jspl jspl_w_n428_1(.douta(w_n428_1[0]),.doutb(w_dff_A_Spe8grpu6_1),.din(w_n428_0[0]));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl3 jspl3_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.doutc(w_n433_0[2]),.din(n433));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl jspl_w_n435_2(.douta(w_n435_2[0]),.doutb(w_n435_2[1]),.din(w_n435_0[1]));
	jspl jspl_w_n437_0(.douta(w_dff_A_JMj54jpY1_0),.doutb(w_n437_0[1]),.din(w_dff_B_SB3eUVwo7_2));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_dff_A_begpvNal4_1),.doutc(w_n451_0[2]),.din(w_dff_B_fLnXQ0Lb0_3));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_dff_A_9OEWihJg9_1),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_vrW7pce47_1),.doutc(w_n462_0[2]),.din(w_dff_B_d2dBaqaS5_3));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl3 jspl3_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.doutc(w_n471_1[2]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_dff_A_fWW2UeFb7_1),.doutc(w_dff_A_r91G5d5d1_2),.din(w_dff_B_2DsNOHuP7_3));
	jspl jspl_w_n473_1(.douta(w_n473_1[0]),.doutb(w_n473_1[1]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.doutc(w_n483_0[2]),.din(n483));
	jspl3 jspl3_w_n483_1(.douta(w_n483_1[0]),.doutb(w_n483_1[1]),.doutc(w_n483_1[2]),.din(w_n483_0[0]));
	jspl jspl_w_n483_2(.douta(w_n483_2[0]),.doutb(w_n483_2[1]),.din(w_n483_0[1]));
	jspl3 jspl3_w_n485_0(.douta(w_n485_0[0]),.doutb(w_dff_A_Fq7oCxoN3_1),.doutc(w_dff_A_pMW24VFp3_2),.din(w_dff_B_5B0514A33_3));
	jspl jspl_w_n485_1(.douta(w_dff_A_K02QV1Jy0_0),.doutb(w_n485_1[1]),.din(w_n485_0[0]));
	jspl jspl_w_n493_0(.douta(w_n493_0[0]),.doutb(w_n493_0[1]),.din(n493));
	jspl3 jspl3_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.doutc(w_n494_0[2]),.din(n494));
	jspl3 jspl3_w_n494_1(.douta(w_n494_1[0]),.doutb(w_n494_1[1]),.doutc(w_n494_1[2]),.din(w_n494_0[0]));
	jspl3 jspl3_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.doutc(w_dff_A_Kof4lzNX5_2),.din(w_dff_B_OzpKQcnl0_3));
	jspl jspl_w_n496_1(.douta(w_dff_A_JOATgsfg6_0),.doutb(w_n496_1[1]),.din(w_n496_0[0]));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl3 jspl3_w_n509_0(.douta(w_dff_A_5zvoiHyn4_0),.doutb(w_dff_A_g2ibEBXg4_1),.doutc(w_n509_0[2]),.din(w_dff_B_HKAzCg7R7_3));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl3 jspl3_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.doutc(w_n518_1[2]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n520_0(.douta(w_n520_0[0]),.doutb(w_dff_A_SsfZd5P01_1),.doutc(w_n520_0[2]),.din(w_dff_B_9BYI8BGR2_3));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl3 jspl3_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.doutc(w_n530_1[2]),.din(w_n530_0[0]));
	jspl3 jspl3_w_n532_0(.douta(w_n532_0[0]),.doutb(w_dff_A_zxckjhqV0_1),.doutc(w_dff_A_oEkkQGhu1_2),.din(w_dff_B_b9meJiND4_3));
	jspl jspl_w_n532_1(.douta(w_n532_1[0]),.doutb(w_n532_1[1]),.din(w_n532_0[0]));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.doutc(w_n551_0[2]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl3 jspl3_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.doutc(w_n556_5[2]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n556_6(.douta(w_n556_6[0]),.doutb(w_n556_6[1]),.doutc(w_n556_6[2]),.din(w_n556_1[2]));
	jspl3 jspl3_w_n556_7(.douta(w_n556_7[0]),.doutb(w_n556_7[1]),.doutc(w_n556_7[2]),.din(w_n556_2[0]));
	jspl jspl_w_n556_8(.douta(w_n556_8[0]),.doutb(w_n556_8[1]),.din(w_n556_2[1]));
	jspl jspl_w_n557_0(.douta(w_dff_A_zuN3zQmS5_0),.doutb(w_n557_0[1]),.din(n557));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_dff_A_s2LmmwUv5_1),.din(n559));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n561_1(.douta(w_n561_1[0]),.doutb(w_n561_1[1]),.din(w_n561_0[0]));
	jspl jspl_w_n562_0(.douta(w_dff_A_2L149ccd6_0),.doutb(w_n562_0[1]),.din(n562));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_NHIWFKCJ9_1),.din(n564));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n569_0(.douta(w_dff_A_v4ndQapO6_0),.doutb(w_n569_0[1]),.din(n569));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_dff_A_b2al5vls9_1),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_dff_A_E8RvXwhG7_0),.doutb(w_dff_A_6f9bX2tD6_1),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_dff_A_ZC2bstJW3_1),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.doutc(w_n578_0[2]),.din(n578));
	jspl jspl_w_n578_1(.douta(w_n578_1[0]),.doutb(w_n578_1[1]),.din(w_n578_0[0]));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_dff_A_oXcb4rub9_1),.doutc(w_dff_A_apldzcTr2_2),.din(n579));
	jspl jspl_w_n579_1(.douta(w_n579_1[0]),.doutb(w_dff_A_3drH5Idj8_1),.din(w_n579_0[0]));
	jspl jspl_w_n581_0(.douta(w_dff_A_IP7kNLv53_0),.doutb(w_n581_0[1]),.din(n581));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n586_1(.douta(w_n586_1[0]),.doutb(w_n586_1[1]),.din(w_n586_0[0]));
	jspl jspl_w_n587_0(.douta(w_n587_0[0]),.doutb(w_dff_A_oC8bNNVc9_1),.din(n587));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_dff_A_4SjY06lH7_2),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.doutc(w_n591_0[2]),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_dff_A_Rr5OZwbN8_0),.doutb(w_n592_0[1]),.doutc(w_dff_A_ib9Rh1lq1_2),.din(n592));
	jspl3 jspl3_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl jspl_w_n596_1(.douta(w_n596_1[0]),.doutb(w_n596_1[1]),.din(w_n596_0[0]));
	jspl3 jspl3_w_n597_0(.douta(w_dff_A_1T9U05Yz1_0),.doutb(w_n597_0[1]),.doutc(w_n597_0[2]),.din(n597));
	jspl3 jspl3_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.doutc(w_n601_0[2]),.din(n601));
	jspl jspl_w_n601_1(.douta(w_n601_1[0]),.doutb(w_n601_1[1]),.din(w_n601_0[0]));
	jspl3 jspl3_w_n602_0(.douta(w_dff_A_fpZxkH2L2_0),.doutb(w_n602_0[1]),.doutc(w_n602_0[2]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n607_1(.douta(w_n607_1[0]),.doutb(w_n607_1[1]),.din(w_n607_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_dff_A_enWkxjoB9_1),.doutc(w_dff_A_EMhCsHJR1_2),.din(n608));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_dff_A_1UZuqTSm6_1),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n611_0(.douta(w_n611_0[0]),.doutb(w_dff_A_27kRFvmS5_1),.doutc(w_n611_0[2]),.din(w_dff_B_Gk7CQZEh4_3));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.doutc(w_n613_1[2]),.din(w_n613_0[0]));
	jspl3 jspl3_w_n613_2(.douta(w_n613_2[0]),.doutb(w_n613_2[1]),.doutc(w_n613_2[2]),.din(w_n613_0[1]));
	jspl3 jspl3_w_n613_3(.douta(w_n613_3[0]),.doutb(w_n613_3[1]),.doutc(w_n613_3[2]),.din(w_n613_0[2]));
	jspl3 jspl3_w_n613_4(.douta(w_n613_4[0]),.doutb(w_n613_4[1]),.doutc(w_n613_4[2]),.din(w_n613_1[0]));
	jspl3 jspl3_w_n613_5(.douta(w_n613_5[0]),.doutb(w_n613_5[1]),.doutc(w_n613_5[2]),.din(w_n613_1[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_dff_A_zHayOKWN5_1),.doutc(w_dff_A_XOM3sFug4_2),.din(n618));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_dff_A_ZNLjUrh03_1),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n619_1(.douta(w_n619_1[0]),.doutb(w_n619_1[1]),.doutc(w_n619_1[2]),.din(w_n619_0[0]));
	jspl3 jspl3_w_n620_0(.douta(w_n620_0[0]),.doutb(w_dff_A_GwQxQH0o0_1),.doutc(w_dff_A_ioamGLlq1_2),.din(n620));
	jspl jspl_w_n620_1(.douta(w_n620_1[0]),.doutb(w_dff_A_NHz2SRfK7_1),.din(w_n620_0[0]));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_dff_A_tpYJbV0X3_1),.din(n621));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_dff_A_Jhn4XrRk4_0),.doutb(w_dff_A_TizUnkPX5_1),.doutc(w_n624_0[2]),.din(w_dff_B_XUuxerAk5_3));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_dff_A_jmzSzmoB4_1),.din(n625));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl jspl_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n628_0(.douta(w_dff_A_nGDxQYAn0_0),.doutb(w_n628_0[1]),.doutc(w_dff_A_iHYFifiN4_2),.din(n628));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_dff_A_1wofKjqD7_1),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n635_1(.douta(w_dff_A_UPDBQr5m9_0),.doutb(w_n635_1[1]),.din(w_n635_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.doutc(w_n637_0[2]),.din(n637));
	jspl jspl_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.din(n638));
	jspl3 jspl3_w_n639_0(.douta(w_dff_A_hISlCyLZ4_0),.doutb(w_n639_0[1]),.doutc(w_n639_0[2]),.din(n639));
	jspl jspl_w_n640_0(.douta(w_dff_A_pp4HwyNl2_0),.doutb(w_n640_0[1]),.din(n640));
	jspl3 jspl3_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.doutc(w_dff_A_3lMUSRFd5_2),.din(n641));
	jspl3 jspl3_w_n641_1(.douta(w_n641_1[0]),.doutb(w_n641_1[1]),.doutc(w_n641_1[2]),.din(w_n641_0[0]));
	jspl3 jspl3_w_n644_0(.douta(w_dff_A_YnXvQpkT4_0),.doutb(w_n644_0[1]),.doutc(w_dff_A_lxg9sKrs5_2),.din(n644));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_dff_A_hVwjUmak5_1),.doutc(w_dff_A_E5nnNKxj8_2),.din(n648));
	jspl jspl_w_n648_1(.douta(w_n648_1[0]),.doutb(w_n648_1[1]),.din(w_n648_0[0]));
	jspl jspl_w_n649_0(.douta(w_dff_A_M55HYp4e6_0),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n653_0(.douta(w_dff_A_qKiqqAVL5_0),.doutb(w_n653_0[1]),.doutc(w_n653_0[2]),.din(n653));
	jspl3 jspl3_w_n654_0(.douta(w_dff_A_BrKvvSPn1_0),.doutb(w_n654_0[1]),.doutc(w_n654_0[2]),.din(w_dff_B_r3BFdL1o3_3));
	jspl3 jspl3_w_n654_1(.douta(w_n654_1[0]),.doutb(w_dff_A_8SolGUlR1_1),.doutc(w_n654_1[2]),.din(w_n654_0[0]));
	jspl3 jspl3_w_n654_2(.douta(w_dff_A_xFdiiL3z1_0),.doutb(w_n654_2[1]),.doutc(w_n654_2[2]),.din(w_n654_0[1]));
	jspl3 jspl3_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.doutc(w_n658_0[2]),.din(n658));
	jspl jspl_w_n658_1(.douta(w_n658_1[0]),.doutb(w_n658_1[1]),.din(w_n658_0[0]));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_dff_A_L4yrxRrg8_2),.din(n660));
	jspl jspl_w_n660_1(.douta(w_dff_A_38Pjr5fa8_0),.doutb(w_n660_1[1]),.din(w_n660_0[0]));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(w_dff_B_tLzJNkdT5_2));
	jspl jspl_w_n670_0(.douta(w_n670_0[0]),.doutb(w_n670_0[1]),.din(n670));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl3 jspl3_w_n682_0(.douta(w_n682_0[0]),.doutb(w_dff_A_Xw0QZFdE1_1),.doutc(w_dff_A_NxH4tdPn0_2),.din(n682));
	jspl jspl_w_n684_0(.douta(w_dff_A_Awaqc4aS2_0),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_dff_A_KaP3mLZ20_0),.doutb(w_n685_0[1]),.din(w_dff_B_i8QFpFER7_2));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_dff_A_2tTVCuS14_1),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_dff_A_5jgei4zv9_1),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_dff_A_hl6HUjuu1_0),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n692_0(.douta(w_dff_A_Hv98Ul3Y0_0),.doutb(w_n692_0[1]),.din(n692));
	jspl3 jspl3_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.doutc(w_n694_0[2]),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_dff_A_s88eH5Y14_0),.doutb(w_dff_A_Qe9sEAx29_1),.doutc(w_n695_0[2]),.din(n695));
	jspl3 jspl3_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.doutc(w_n699_0[2]),.din(n699));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_dff_A_VySiNYam7_1),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_dff_A_7Weigvoq1_1),.din(n709));
	jspl jspl_w_n710_0(.douta(w_dff_A_F7FvTbIU6_0),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_dff_A_4cNbMmsO6_0),.doutb(w_n711_0[1]),.din(n711));
	jspl3 jspl3_w_n713_0(.douta(w_n713_0[0]),.doutb(w_dff_A_srQ6aHx94_1),.doutc(w_n713_0[2]),.din(n713));
	jspl3 jspl3_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.doutc(w_n715_0[2]),.din(n715));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(w_dff_B_QAeNhS517_2));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_dff_A_1awB07r12_1),.din(n719));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_dff_A_p4Fayc1v9_1),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_dff_A_XKG0JAaY6_1),.din(n721));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_dff_A_8hthiOcC1_1),.din(n722));
	jspl3 jspl3_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.doutc(w_n725_0[2]),.din(n725));
	jspl jspl_w_n726_0(.douta(w_dff_A_qDepDr3V9_0),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.doutc(w_n733_0[2]),.din(n733));
	jspl3 jspl3_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.doutc(w_n735_0[2]),.din(n735));
	jspl3 jspl3_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl jspl_w_n737_1(.douta(w_n737_1[0]),.doutb(w_n737_1[1]),.din(w_n737_0[0]));
	jspl jspl_w_n738_0(.douta(w_n738_0[0]),.doutb(w_n738_0[1]),.din(n738));
	jspl3 jspl3_w_n742_0(.douta(w_n742_0[0]),.doutb(w_dff_A_QbkPiTFN8_1),.doutc(w_n742_0[2]),.din(n742));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_dff_A_1cjKdCl93_1),.doutc(w_n746_0[2]),.din(n746));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(w_dff_B_pKIMdEps8_2));
	jspl3 jspl3_w_n749_0(.douta(w_n749_0[0]),.doutb(w_dff_A_lYHRuC0r7_1),.doutc(w_dff_A_dbchnsP29_2),.din(n749));
	jspl3 jspl3_w_n749_1(.douta(w_n749_1[0]),.doutb(w_dff_A_WSPSDGqZ9_1),.doutc(w_dff_A_MsncRhbx1_2),.din(w_n749_0[0]));
	jspl3 jspl3_w_n749_2(.douta(w_dff_A_UGEY9o3W6_0),.doutb(w_dff_A_r6mjsyH68_1),.doutc(w_n749_2[2]),.din(w_n749_0[1]));
	jspl3 jspl3_w_n749_3(.douta(w_dff_A_Q62aijYp6_0),.doutb(w_n749_3[1]),.doutc(w_dff_A_QcqzsMkw0_2),.din(w_n749_0[2]));
	jspl3 jspl3_w_n749_4(.douta(w_n749_4[0]),.doutb(w_dff_A_CQbw284R5_1),.doutc(w_dff_A_oRDUx95A7_2),.din(w_n749_1[0]));
	jspl3 jspl3_w_n749_5(.douta(w_dff_A_aUEeXtDh7_0),.doutb(w_dff_A_Y5kv7rC74_1),.doutc(w_n749_5[2]),.din(w_n749_1[1]));
	jspl3 jspl3_w_n749_6(.douta(w_dff_A_O9OK7o6x9_0),.doutb(w_n749_6[1]),.doutc(w_n749_6[2]),.din(w_n749_1[2]));
	jspl3 jspl3_w_n749_7(.douta(w_dff_A_jhT5jWgK2_0),.doutb(w_n749_7[1]),.doutc(w_n749_7[2]),.din(w_n749_2[0]));
	jspl3 jspl3_w_n749_8(.douta(w_n749_8[0]),.doutb(w_dff_A_GPQp5Te57_1),.doutc(w_dff_A_kRe9C1FU2_2),.din(w_n749_2[1]));
	jspl3 jspl3_w_n749_9(.douta(w_dff_A_NxClbYBH0_0),.doutb(w_n749_9[1]),.doutc(w_dff_A_aOqhSAk29_2),.din(w_n749_2[2]));
	jspl3 jspl3_w_n749_10(.douta(w_n749_10[0]),.doutb(w_n749_10[1]),.doutc(w_n749_10[2]),.din(w_n749_3[0]));
	jspl3 jspl3_w_n749_11(.douta(w_dff_A_9JjDmRhG0_0),.doutb(w_dff_A_7TidQJ6G5_1),.doutc(w_n749_11[2]),.din(w_n749_3[1]));
	jspl3 jspl3_w_n749_12(.douta(w_n749_12[0]),.doutb(w_n749_12[1]),.doutc(w_n749_12[2]),.din(w_n749_3[2]));
	jspl jspl_w_n749_13(.douta(w_dff_A_MYjoLYpB8_0),.doutb(w_n749_13[1]),.din(w_n749_4[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.doutc(w_n750_0[2]),.din(n750));
	jspl3 jspl3_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.doutc(w_n750_1[2]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n750_2(.douta(w_n750_2[0]),.doutb(w_n750_2[1]),.doutc(w_n750_2[2]),.din(w_n750_0[1]));
	jspl3 jspl3_w_n750_3(.douta(w_n750_3[0]),.doutb(w_n750_3[1]),.doutc(w_n750_3[2]),.din(w_n750_0[2]));
	jspl3 jspl3_w_n750_4(.douta(w_n750_4[0]),.doutb(w_n750_4[1]),.doutc(w_n750_4[2]),.din(w_n750_1[0]));
	jspl3 jspl3_w_n750_5(.douta(w_n750_5[0]),.doutb(w_n750_5[1]),.doutc(w_n750_5[2]),.din(w_n750_1[1]));
	jspl3 jspl3_w_n750_6(.douta(w_n750_6[0]),.doutb(w_n750_6[1]),.doutc(w_n750_6[2]),.din(w_n750_1[2]));
	jspl3 jspl3_w_n750_7(.douta(w_n750_7[0]),.doutb(w_n750_7[1]),.doutc(w_n750_7[2]),.din(w_n750_2[0]));
	jspl3 jspl3_w_n750_8(.douta(w_n750_8[0]),.doutb(w_n750_8[1]),.doutc(w_n750_8[2]),.din(w_n750_2[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_dff_A_Xx2je7Ng9_1),.doutc(w_dff_A_eCToI8218_2),.din(w_dff_B_KcNeIWmv8_3));
	jspl jspl_w_n753_1(.douta(w_dff_A_xrLt9rQJ6_0),.doutb(w_n753_1[1]),.din(w_n753_0[0]));
	jspl jspl_w_n755_0(.douta(w_dff_A_AFcJoeIn8_0),.doutb(w_n755_0[1]),.din(n755));
	jspl3 jspl3_w_n763_0(.douta(w_dff_A_Nh5iaij37_0),.doutb(w_n763_0[1]),.doutc(w_n763_0[2]),.din(n763));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl jspl_w_n779_0(.douta(w_dff_A_qnGRR56D9_0),.doutb(w_n779_0[1]),.din(n779));
	jspl3 jspl3_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.doutc(w_n786_0[2]),.din(n786));
	jspl3 jspl3_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.doutc(w_n788_0[2]),.din(n788));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_dff_A_4MuFKhJy2_1),.doutc(w_n790_0[2]),.din(n790));
	jspl3 jspl3_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.doutc(w_dff_A_68PoRUC35_2),.din(n792));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_n797_1[1]),.doutc(w_n797_1[2]),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_n797_2[2]),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_dff_A_ExNRHowj8_0),.doutb(w_n797_3[1]),.doutc(w_n797_3[2]),.din(w_n797_0[2]));
	jspl3 jspl3_w_n797_4(.douta(w_dff_A_58dpKpKG9_0),.doutb(w_n797_4[1]),.doutc(w_dff_A_vwgUazEv3_2),.din(w_n797_1[0]));
	jspl3 jspl3_w_n797_5(.douta(w_n797_5[0]),.doutb(w_dff_A_a30Dc9h31_1),.doutc(w_n797_5[2]),.din(w_n797_1[1]));
	jspl3 jspl3_w_n797_6(.douta(w_dff_A_tb1vKi2D2_0),.doutb(w_n797_6[1]),.doutc(w_dff_A_Ll5Z3cAM9_2),.din(w_n797_1[2]));
	jspl3 jspl3_w_n797_7(.douta(w_n797_7[0]),.doutb(w_dff_A_OTCTdaMt9_1),.doutc(w_n797_7[2]),.din(w_n797_2[0]));
	jspl3 jspl3_w_n797_8(.douta(w_dff_A_RMKQ9xKZ3_0),.doutb(w_n797_8[1]),.doutc(w_dff_A_szCXB5hr2_2),.din(w_n797_2[1]));
	jspl jspl_w_n797_9(.douta(w_n797_9[0]),.doutb(w_dff_A_losgSMuX1_1),.din(w_n797_2[2]));
	jspl3 jspl3_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.doutc(w_n798_0[2]),.din(n798));
	jspl jspl_w_n798_1(.douta(w_n798_1[0]),.doutb(w_n798_1[1]),.din(w_n798_0[0]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_dff_A_ChpFXZM95_1),.doutc(w_dff_A_6zlKOZOd4_2),.din(w_dff_B_1YMFOaP55_3));
	jspl3 jspl3_w_n800_1(.douta(w_n800_1[0]),.doutb(w_dff_A_29YK8VA16_1),.doutc(w_dff_A_Pbl6qVni4_2),.din(w_n800_0[0]));
	jspl3 jspl3_w_n800_2(.douta(w_n800_2[0]),.doutb(w_n800_2[1]),.doutc(w_dff_A_4tE30Vwy7_2),.din(w_n800_0[1]));
	jspl3 jspl3_w_n800_3(.douta(w_dff_A_foNLMS0P2_0),.doutb(w_n800_3[1]),.doutc(w_dff_A_ptkvh7EA1_2),.din(w_n800_0[2]));
	jspl jspl_w_n800_4(.douta(w_dff_A_zylMXVli7_0),.doutb(w_n800_4[1]),.din(w_n800_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl jspl_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n814_0(.douta(w_dff_A_12ZkINdP0_0),.doutb(w_dff_A_TJs1W6DT4_1),.doutc(w_n814_0[2]),.din(n814));
	jspl3 jspl3_w_n819_0(.douta(w_n819_0[0]),.doutb(w_dff_A_IYJMrDp93_1),.doutc(w_n819_0[2]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_dff_A_mfsUWL0M9_1),.din(n821));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n836_0(.douta(w_dff_A_V7JhJi4I3_0),.doutb(w_n836_0[1]),.din(n836));
	jspl jspl_w_n847_0(.douta(w_dff_A_3lqhmAhK7_0),.doutb(w_n847_0[1]),.din(n847));
	jspl3 jspl3_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.doutc(w_n852_0[2]),.din(n852));
	jspl3 jspl3_w_n852_1(.douta(w_n852_1[0]),.doutb(w_n852_1[1]),.doutc(w_n852_1[2]),.din(w_n852_0[0]));
	jspl3 jspl3_w_n852_2(.douta(w_n852_2[0]),.doutb(w_n852_2[1]),.doutc(w_n852_2[2]),.din(w_n852_0[1]));
	jspl3 jspl3_w_n852_3(.douta(w_dff_A_gPRdKgN45_0),.doutb(w_n852_3[1]),.doutc(w_n852_3[2]),.din(w_n852_0[2]));
	jspl3 jspl3_w_n852_4(.douta(w_dff_A_bNh4M6Ep2_0),.doutb(w_n852_4[1]),.doutc(w_dff_A_FHS91h1n8_2),.din(w_n852_1[0]));
	jspl3 jspl3_w_n852_5(.douta(w_n852_5[0]),.doutb(w_dff_A_WPWSIian4_1),.doutc(w_dff_A_NG1cNPox5_2),.din(w_n852_1[1]));
	jspl3 jspl3_w_n852_6(.douta(w_n852_6[0]),.doutb(w_n852_6[1]),.doutc(w_dff_A_GbTFOAwC9_2),.din(w_n852_1[2]));
	jspl3 jspl3_w_n852_7(.douta(w_dff_A_z4pdcwoX3_0),.doutb(w_n852_7[1]),.doutc(w_dff_A_js8pimOP0_2),.din(w_n852_2[0]));
	jspl3 jspl3_w_n852_8(.douta(w_n852_8[0]),.doutb(w_dff_A_p2KaDZoD7_1),.doutc(w_n852_8[2]),.din(w_n852_2[1]));
	jspl jspl_w_n852_9(.douta(w_n852_9[0]),.doutb(w_dff_A_GStFKiis3_1),.din(w_n852_2[2]));
	jspl3 jspl3_w_n854_0(.douta(w_n854_0[0]),.doutb(w_dff_A_DhjotKiY6_1),.doutc(w_dff_A_GJS3iESA2_2),.din(w_dff_B_LKKyFNdM0_3));
	jspl3 jspl3_w_n854_1(.douta(w_n854_1[0]),.doutb(w_dff_A_MADeFKk91_1),.doutc(w_dff_A_cFnCmMlb6_2),.din(w_n854_0[0]));
	jspl3 jspl3_w_n854_2(.douta(w_n854_2[0]),.doutb(w_n854_2[1]),.doutc(w_n854_2[2]),.din(w_n854_0[1]));
	jspl3 jspl3_w_n854_3(.douta(w_n854_3[0]),.doutb(w_n854_3[1]),.doutc(w_dff_A_nMHJbxjT1_2),.din(w_n854_0[2]));
	jspl jspl_w_n854_4(.douta(w_dff_A_p2PiHSc06_0),.doutb(w_n854_4[1]),.din(w_n854_1[0]));
	jspl3 jspl3_w_n865_0(.douta(w_dff_A_S4J3oz055_0),.doutb(w_n865_0[1]),.doutc(w_dff_A_QqAqicj04_2),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n868_0(.douta(w_n868_0[0]),.doutb(w_n868_0[1]),.din(n868));
	jspl jspl_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.din(n870));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl jspl_w_n880_0(.douta(w_dff_A_Pp1HGQRd6_0),.doutb(w_n880_0[1]),.din(n880));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(n890));
	jspl jspl_w_n901_0(.douta(w_dff_A_EsAjOgU65_0),.doutb(w_n901_0[1]),.din(n901));
	jspl3 jspl3_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.doutc(w_n923_0[2]),.din(n923));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl3 jspl3_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.doutc(w_dff_A_GBmzx6wz4_2),.din(n938));
	jspl3 jspl3_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.doutc(w_n940_0[2]),.din(n940));
	jspl jspl_w_n940_1(.douta(w_n940_1[0]),.doutb(w_n940_1[1]),.din(w_n940_0[0]));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(n944));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_dff_A_uXdx9I4O0_1),.din(n949));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl3 jspl3_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.doutc(w_dff_A_xgc5JR2D4_2),.din(n954));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_dff_A_qKtk3BAZ0_1),.din(w_dff_B_06dA8gXU0_2));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl3 jspl3_w_n977_0(.douta(w_n977_0[0]),.doutb(w_n977_0[1]),.doutc(w_n977_0[2]),.din(n977));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_dff_A_wfN3sNeB6_1),.din(n989));
	jspl3 jspl3_w_n993_0(.douta(w_n993_0[0]),.doutb(w_dff_A_KDQYG55A6_1),.doutc(w_dff_A_HLISzOAQ6_2),.din(n993));
	jspl3 jspl3_w_n993_1(.douta(w_n993_1[0]),.doutb(w_dff_A_LPoxAlm50_1),.doutc(w_dff_A_bFcptGNJ2_2),.din(w_n993_0[0]));
	jspl3 jspl3_w_n993_2(.douta(w_dff_A_5xdz7XYU7_0),.doutb(w_dff_A_Hpy5MfOc2_1),.doutc(w_n993_2[2]),.din(w_n993_0[1]));
	jspl3 jspl3_w_n993_3(.douta(w_dff_A_gamMfp6T9_0),.doutb(w_dff_A_iXDsf0Av2_1),.doutc(w_n993_3[2]),.din(w_n993_0[2]));
	jspl3 jspl3_w_n993_4(.douta(w_dff_A_GY8z1wY53_0),.doutb(w_dff_A_0fxBTHVS6_1),.doutc(w_n993_4[2]),.din(w_n993_1[0]));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n994_1(.douta(w_n994_1[0]),.doutb(w_n994_1[1]),.doutc(w_n994_1[2]),.din(w_n994_0[0]));
	jspl3 jspl3_w_n994_2(.douta(w_n994_2[0]),.doutb(w_n994_2[1]),.doutc(w_n994_2[2]),.din(w_n994_0[1]));
	jspl3 jspl3_w_n994_3(.douta(w_n994_3[0]),.doutb(w_n994_3[1]),.doutc(w_n994_3[2]),.din(w_n994_0[2]));
	jspl jspl_w_n994_4(.douta(w_n994_4[0]),.doutb(w_n994_4[1]),.din(w_n994_1[0]));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl3 jspl3_w_n996_1(.douta(w_n996_1[0]),.doutb(w_n996_1[1]),.doutc(w_n996_1[2]),.din(w_n996_0[0]));
	jspl3 jspl3_w_n996_2(.douta(w_n996_2[0]),.doutb(w_n996_2[1]),.doutc(w_n996_2[2]),.din(w_n996_0[1]));
	jspl3 jspl3_w_n996_3(.douta(w_n996_3[0]),.doutb(w_n996_3[1]),.doutc(w_n996_3[2]),.din(w_n996_0[2]));
	jspl jspl_w_n996_4(.douta(w_n996_4[0]),.doutb(w_n996_4[1]),.din(w_n996_1[0]));
	jspl3 jspl3_w_n999_0(.douta(w_dff_A_VMh60d2x4_0),.doutb(w_dff_A_eZp5P86f6_1),.doutc(w_n999_0[2]),.din(w_dff_B_XHslf9w03_3));
	jspl3 jspl3_w_n999_1(.douta(w_dff_A_yDlvjHw96_0),.doutb(w_dff_A_1hELk9MS9_1),.doutc(w_n999_1[2]),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_dff_A_VOAFHszn5_0),.doutb(w_dff_A_APFbucbk9_1),.doutc(w_n999_2[2]),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_dff_A_RUcvG7n60_0),.doutb(w_dff_A_ex2SzdNi7_1),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl3 jspl3_w_n1007_0(.douta(w_dff_A_H4V82B3V1_0),.doutb(w_dff_A_u2T2DKa28_1),.doutc(w_n1007_0[2]),.din(w_dff_B_djOsCc3g3_3));
	jspl3 jspl3_w_n1007_1(.douta(w_n1007_1[0]),.doutb(w_n1007_1[1]),.doutc(w_dff_A_0YtcJIVr1_2),.din(w_n1007_0[0]));
	jspl3 jspl3_w_n1007_2(.douta(w_dff_A_eY1SVWxl9_0),.doutb(w_dff_A_A9qC9FTc9_1),.doutc(w_n1007_2[2]),.din(w_n1007_0[1]));
	jspl3 jspl3_w_n1007_3(.douta(w_dff_A_npS2ivQk8_0),.doutb(w_dff_A_6u7w5u6X9_1),.doutc(w_n1007_3[2]),.din(w_n1007_0[2]));
	jspl3 jspl3_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_dff_A_b1Z1GqIh7_1),.doutc(w_dff_A_wtsjZLC43_2),.din(n1008));
	jspl3 jspl3_w_n1008_1(.douta(w_n1008_1[0]),.doutb(w_dff_A_pQ3HAkyF6_1),.doutc(w_dff_A_SwhyDRds8_2),.din(w_n1008_0[0]));
	jspl3 jspl3_w_n1008_2(.douta(w_dff_A_bDAjTJQY5_0),.doutb(w_dff_A_5i6QK7o84_1),.doutc(w_n1008_2[2]),.din(w_n1008_0[1]));
	jspl3 jspl3_w_n1008_3(.douta(w_dff_A_QiqEtPaT6_0),.doutb(w_dff_A_LWUS1reT6_1),.doutc(w_n1008_3[2]),.din(w_n1008_0[2]));
	jspl3 jspl3_w_n1008_4(.douta(w_dff_A_SKWies1N4_0),.doutb(w_n1008_4[1]),.doutc(w_dff_A_mZ86McBp3_2),.din(w_n1008_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl3 jspl3_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.doutc(w_n1012_1[2]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1012_2(.douta(w_n1012_2[0]),.doutb(w_n1012_2[1]),.doutc(w_n1012_2[2]),.din(w_n1012_0[1]));
	jspl3 jspl3_w_n1012_3(.douta(w_n1012_3[0]),.doutb(w_n1012_3[1]),.doutc(w_n1012_3[2]),.din(w_n1012_0[2]));
	jspl jspl_w_n1012_4(.douta(w_n1012_4[0]),.doutb(w_n1012_4[1]),.din(w_n1012_1[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl3 jspl3_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.doutc(w_n1014_1[2]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1014_2(.douta(w_n1014_2[0]),.doutb(w_n1014_2[1]),.doutc(w_n1014_2[2]),.din(w_n1014_0[1]));
	jspl3 jspl3_w_n1014_3(.douta(w_n1014_3[0]),.doutb(w_n1014_3[1]),.doutc(w_n1014_3[2]),.din(w_n1014_0[2]));
	jspl jspl_w_n1014_4(.douta(w_n1014_4[0]),.doutb(w_n1014_4[1]),.din(w_n1014_1[0]));
	jspl3 jspl3_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.doutc(w_n1019_0[2]),.din(n1019));
	jspl jspl_w_n1019_1(.douta(w_n1019_1[0]),.doutb(w_n1019_1[1]),.din(w_n1019_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl3 jspl3_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.doutc(w_n1043_0[2]),.din(n1043));
	jspl jspl_w_n1043_1(.douta(w_n1043_1[0]),.doutb(w_n1043_1[1]),.din(w_n1043_0[0]));
	jspl3 jspl3_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.doutc(w_n1052_0[2]),.din(n1052));
	jspl jspl_w_n1052_1(.douta(w_n1052_1[0]),.doutb(w_n1052_1[1]),.din(w_n1052_0[0]));
	jspl3 jspl3_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.doutc(w_n1054_0[2]),.din(n1054));
	jspl jspl_w_n1054_1(.douta(w_n1054_1[0]),.doutb(w_n1054_1[1]),.din(w_n1054_0[0]));
	jspl jspl_w_n1177_0(.douta(w_dff_A_q0KUU9WO9_0),.doutb(w_n1177_0[1]),.din(w_dff_B_eBuerXZk9_2));
	jspl jspl_w_n1179_0(.douta(w_dff_A_HFFMZKXC4_0),.doutb(w_n1179_0[1]),.din(n1179));
	jspl3 jspl3_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.doutc(w_n1196_0[2]),.din(n1196));
	jspl3 jspl3_w_n1196_1(.douta(w_n1196_1[0]),.doutb(w_n1196_1[1]),.doutc(w_n1196_1[2]),.din(w_n1196_0[0]));
	jspl3 jspl3_w_n1201_0(.douta(w_dff_A_nshC9MZh4_0),.doutb(w_dff_A_Tjcoy3949_1),.doutc(w_n1201_0[2]),.din(w_dff_B_Vg4hOFcp5_3));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.doutc(w_n1213_0[2]),.din(n1213));
	jspl3 jspl3_w_n1213_1(.douta(w_n1213_1[0]),.doutb(w_n1213_1[1]),.doutc(w_n1213_1[2]),.din(w_n1213_0[0]));
	jspl3 jspl3_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.doutc(w_n1236_0[2]),.din(n1236));
	jspl3 jspl3_w_n1236_1(.douta(w_n1236_1[0]),.doutb(w_n1236_1[1]),.doutc(w_n1236_1[2]),.din(w_n1236_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl3 jspl3_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.doutc(w_n1251_1[2]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.doutc(w_n1279_0[2]),.din(n1279));
	jspl jspl_w_n1279_1(.douta(w_n1279_1[0]),.doutb(w_n1279_1[1]),.din(w_n1279_0[0]));
	jspl3 jspl3_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.doutc(w_n1297_0[2]),.din(n1297));
	jspl jspl_w_n1297_1(.douta(w_n1297_1[0]),.doutb(w_n1297_1[1]),.din(w_n1297_0[0]));
	jspl3 jspl3_w_n1299_0(.douta(w_n1299_0[0]),.doutb(w_n1299_0[1]),.doutc(w_n1299_0[2]),.din(n1299));
	jspl jspl_w_n1299_1(.douta(w_n1299_1[0]),.doutb(w_n1299_1[1]),.din(w_n1299_0[0]));
	jspl3 jspl3_w_n1410_0(.douta(w_dff_A_xGYv2QMQ1_0),.doutb(w_n1410_0[1]),.doutc(w_n1410_0[2]),.din(n1410));
	jspl3 jspl3_w_n1412_0(.douta(w_n1412_0[0]),.doutb(w_dff_A_uacR1U299_1),.doutc(w_dff_A_7rkIrt1C7_2),.din(w_dff_B_1mfQGzjy0_3));
	jspl jspl_w_n1416_0(.douta(w_n1416_0[0]),.doutb(w_n1416_0[1]),.din(n1416));
	jspl jspl_w_n1422_0(.douta(w_dff_A_O4Bg95WV8_0),.doutb(w_n1422_0[1]),.din(n1422));
	jspl jspl_w_n1425_0(.douta(w_dff_A_5WLf0liM1_0),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(n1428));
	jspl jspl_w_n1429_0(.douta(w_dff_A_fLKCUw2Z1_0),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1451_0(.douta(w_dff_A_TmQHv6xl0_0),.doutb(w_n1451_0[1]),.din(n1451));
	jspl jspl_w_n1503_0(.douta(w_n1503_0[0]),.doutb(w_n1503_0[1]),.din(n1503));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1592_0(.douta(w_n1592_0[0]),.doutb(w_n1592_0[1]),.din(n1592));
	jspl jspl_w_n1593_0(.douta(w_n1593_0[0]),.doutb(w_n1593_0[1]),.din(n1593));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1599_0(.douta(w_dff_A_DCcBNEoT4_0),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_n1603_0[1]),.din(n1603));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl3 jspl3_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.doutc(w_n1611_0[2]),.din(n1611));
	jspl jspl_w_n1613_0(.douta(w_dff_A_SdXrTuRN7_0),.doutb(w_n1613_0[1]),.din(n1613));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(n1615));
	jspl jspl_w_n1618_0(.douta(w_dff_A_c1571MWv0_0),.doutb(w_n1618_0[1]),.din(w_dff_B_fCBI0eF75_2));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(w_dff_B_K5Phutoi0_2));
	jspl jspl_w_n1637_0(.douta(w_dff_A_LEtQZjGE5_0),.doutb(w_n1637_0[1]),.din(w_dff_B_pJnT534a4_2));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(n1643));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_dff_A_L7QMeyn52_1),.din(n1652));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl3 jspl3_w_n1674_0(.douta(w_n1674_0[0]),.doutb(w_n1674_0[1]),.doutc(w_n1674_0[2]),.din(n1674));
	jspl jspl_w_n1675_0(.douta(w_n1675_0[0]),.doutb(w_n1675_0[1]),.din(n1675));
	jspl3 jspl3_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.doutc(w_n1679_0[2]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(w_dff_B_ZhlFiBiX3_2));
	jspl jspl_w_n1695_0(.douta(w_n1695_0[0]),.doutb(w_n1695_0[1]),.din(w_dff_B_AzGMDA8y8_2));
	jspl jspl_w_n1698_0(.douta(w_n1698_0[0]),.doutb(w_n1698_0[1]),.din(w_dff_B_SHjTvCFN8_2));
	jdff dff_B_xJVd7vh19_1(.din(G136),.dout(w_dff_B_xJVd7vh19_1),.clk(gclk));
	jdff dff_B_NeekBaFp4_0(.din(G2824),.dout(w_dff_B_NeekBaFp4_0),.clk(gclk));
	jdff dff_B_H5ICgJDO2_1(.din(n320),.dout(w_dff_B_H5ICgJDO2_1),.clk(gclk));
	jdff dff_B_T4h4UUWo7_1(.din(n327),.dout(w_dff_B_T4h4UUWo7_1),.clk(gclk));
	jdff dff_B_m9fN94CJ9_2(.din(n333),.dout(w_dff_B_m9fN94CJ9_2),.clk(gclk));
	jdff dff_B_FiSJvVee4_1(.din(n338),.dout(w_dff_B_FiSJvVee4_1),.clk(gclk));
	jdff dff_B_V1WkeonP1_1(.din(n340),.dout(w_dff_B_V1WkeonP1_1),.clk(gclk));
	jdff dff_B_dFPnBT7I9_0(.din(n341),.dout(w_dff_B_dFPnBT7I9_0),.clk(gclk));
	jdff dff_B_AUPL4UiY9_1(.din(G24),.dout(w_dff_B_AUPL4UiY9_1),.clk(gclk));
	jdff dff_B_ELkE3jRs4_1(.din(n345),.dout(w_dff_B_ELkE3jRs4_1),.clk(gclk));
	jdff dff_B_PDYKQJxI2_0(.din(n346),.dout(w_dff_B_PDYKQJxI2_0),.clk(gclk));
	jdff dff_B_u5UjHSah1_1(.din(G26),.dout(w_dff_B_u5UjHSah1_1),.clk(gclk));
	jdff dff_A_EyYMh1gb3_0(.dout(w_G141_2[0]),.din(w_dff_A_EyYMh1gb3_0),.clk(gclk));
	jdff dff_A_hBgOeFl60_0(.dout(w_dff_A_EyYMh1gb3_0),.din(w_dff_A_hBgOeFl60_0),.clk(gclk));
	jdff dff_A_naU6d0v53_0(.dout(w_dff_A_hBgOeFl60_0),.din(w_dff_A_naU6d0v53_0),.clk(gclk));
	jdff dff_A_G139qUXC6_0(.dout(w_dff_A_naU6d0v53_0),.din(w_dff_A_G139qUXC6_0),.clk(gclk));
	jdff dff_A_isseKvlO1_1(.dout(w_G141_2[1]),.din(w_dff_A_isseKvlO1_1),.clk(gclk));
	jdff dff_A_V6aJmz8T1_1(.dout(w_dff_A_isseKvlO1_1),.din(w_dff_A_V6aJmz8T1_1),.clk(gclk));
	jdff dff_A_z4bRBYaS8_1(.dout(w_dff_A_V6aJmz8T1_1),.din(w_dff_A_z4bRBYaS8_1),.clk(gclk));
	jdff dff_A_9pMjfsWj9_1(.dout(w_dff_A_z4bRBYaS8_1),.din(w_dff_A_9pMjfsWj9_1),.clk(gclk));
	jdff dff_B_7UYQIOoi0_1(.din(n350),.dout(w_dff_B_7UYQIOoi0_1),.clk(gclk));
	jdff dff_B_Mo4niKpk5_0(.din(n351),.dout(w_dff_B_Mo4niKpk5_0),.clk(gclk));
	jdff dff_B_9OtLNadY3_1(.din(G79),.dout(w_dff_B_9OtLNadY3_1),.clk(gclk));
	jdff dff_B_KSukqhV45_1(.din(n355),.dout(w_dff_B_KSukqhV45_1),.clk(gclk));
	jdff dff_B_kBiuCscR6_1(.din(w_dff_B_KSukqhV45_1),.dout(w_dff_B_kBiuCscR6_1),.clk(gclk));
	jdff dff_B_OnyUwNWl5_1(.din(G82),.dout(w_dff_B_OnyUwNWl5_1),.clk(gclk));
	jdff dff_A_5H7xdybX2_0(.dout(w_G2358_2[0]),.din(w_dff_A_5H7xdybX2_0),.clk(gclk));
	jdff dff_A_tmZmnfvl0_1(.dout(w_G2358_2[1]),.din(w_dff_A_tmZmnfvl0_1),.clk(gclk));
	jdff dff_A_2bn3N6YZ7_1(.dout(w_G141_1[1]),.din(w_dff_A_2bn3N6YZ7_1),.clk(gclk));
	jdff dff_A_3GYoWiuU0_1(.dout(w_dff_A_2bn3N6YZ7_1),.din(w_dff_A_3GYoWiuU0_1),.clk(gclk));
	jdff dff_A_6YSjiHj03_1(.dout(w_dff_A_3GYoWiuU0_1),.din(w_dff_A_6YSjiHj03_1),.clk(gclk));
	jdff dff_A_TU9gGnzH5_1(.dout(w_dff_A_6YSjiHj03_1),.din(w_dff_A_TU9gGnzH5_1),.clk(gclk));
	jdff dff_A_kMWxVDrh2_2(.dout(w_G141_1[2]),.din(w_dff_A_kMWxVDrh2_2),.clk(gclk));
	jdff dff_A_jZ6qwYt01_2(.dout(w_dff_A_kMWxVDrh2_2),.din(w_dff_A_jZ6qwYt01_2),.clk(gclk));
	jdff dff_A_bRtp74It2_2(.dout(w_dff_A_jZ6qwYt01_2),.din(w_dff_A_bRtp74It2_2),.clk(gclk));
	jdff dff_A_edFeGmke8_2(.dout(w_dff_A_bRtp74It2_2),.din(w_dff_A_edFeGmke8_2),.clk(gclk));
	jdff dff_B_ppgzI1QW4_1(.din(n373),.dout(w_dff_B_ppgzI1QW4_1),.clk(gclk));
	jdff dff_B_WslEtSt70_2(.din(n661),.dout(w_dff_B_WslEtSt70_2),.clk(gclk));
	jdff dff_B_tLzJNkdT5_2(.din(w_dff_B_WslEtSt70_2),.dout(w_dff_B_tLzJNkdT5_2),.clk(gclk));
	jdff dff_B_Tm0nih7h7_2(.din(n717),.dout(w_dff_B_Tm0nih7h7_2),.clk(gclk));
	jdff dff_B_QAeNhS517_2(.din(w_dff_B_Tm0nih7h7_2),.dout(w_dff_B_QAeNhS517_2),.clk(gclk));
	jdff dff_B_HxvTgeKW1_1(.din(n705),.dout(w_dff_B_HxvTgeKW1_1),.clk(gclk));
	jdff dff_B_MCOzTeU11_1(.din(w_dff_B_HxvTgeKW1_1),.dout(w_dff_B_MCOzTeU11_1),.clk(gclk));
	jdff dff_B_LM8uvOAs5_1(.din(w_dff_B_MCOzTeU11_1),.dout(w_dff_B_LM8uvOAs5_1),.clk(gclk));
	jdff dff_B_Wl4ntgBJ8_1(.din(w_dff_B_LM8uvOAs5_1),.dout(w_dff_B_Wl4ntgBJ8_1),.clk(gclk));
	jdff dff_B_EUhZeJeu1_1(.din(w_dff_B_Wl4ntgBJ8_1),.dout(w_dff_B_EUhZeJeu1_1),.clk(gclk));
	jdff dff_B_QUdYuxkV7_1(.din(w_dff_B_EUhZeJeu1_1),.dout(w_dff_B_QUdYuxkV7_1),.clk(gclk));
	jdff dff_B_0mqaafZo4_1(.din(n706),.dout(w_dff_B_0mqaafZo4_1),.clk(gclk));
	jdff dff_B_wDUsRAim3_1(.din(w_dff_B_0mqaafZo4_1),.dout(w_dff_B_wDUsRAim3_1),.clk(gclk));
	jdff dff_B_0oPw1zAC4_1(.din(w_dff_B_wDUsRAim3_1),.dout(w_dff_B_0oPw1zAC4_1),.clk(gclk));
	jdff dff_B_SWBiYy6v8_1(.din(w_dff_B_0oPw1zAC4_1),.dout(w_dff_B_SWBiYy6v8_1),.clk(gclk));
	jdff dff_B_V8QbOeQJ2_1(.din(w_dff_B_SWBiYy6v8_1),.dout(w_dff_B_V8QbOeQJ2_1),.clk(gclk));
	jdff dff_A_qgprgtJz4_1(.dout(w_n611_0[1]),.din(w_dff_A_qgprgtJz4_1),.clk(gclk));
	jdff dff_A_27kRFvmS5_1(.dout(w_dff_A_qgprgtJz4_1),.din(w_dff_A_27kRFvmS5_1),.clk(gclk));
	jdff dff_B_Gk7CQZEh4_3(.din(n611),.dout(w_dff_B_Gk7CQZEh4_3),.clk(gclk));
	jdff dff_B_rVPAffzR7_2(.din(n747),.dout(w_dff_B_rVPAffzR7_2),.clk(gclk));
	jdff dff_B_pKIMdEps8_2(.din(w_dff_B_rVPAffzR7_2),.dout(w_dff_B_pKIMdEps8_2),.clk(gclk));
	jdff dff_B_Ug8Ns8L68_1(.din(n739),.dout(w_dff_B_Ug8Ns8L68_1),.clk(gclk));
	jdff dff_B_faKqSggN7_1(.din(w_dff_B_Ug8Ns8L68_1),.dout(w_dff_B_faKqSggN7_1),.clk(gclk));
	jdff dff_A_TUQM28mg7_0(.dout(w_n660_1[0]),.din(w_dff_A_TUQM28mg7_0),.clk(gclk));
	jdff dff_A_LqDBCJup0_0(.dout(w_dff_A_TUQM28mg7_0),.din(w_dff_A_LqDBCJup0_0),.clk(gclk));
	jdff dff_A_hOsm0uFm5_0(.dout(w_dff_A_LqDBCJup0_0),.din(w_dff_A_hOsm0uFm5_0),.clk(gclk));
	jdff dff_A_33gZIik94_0(.dout(w_dff_A_hOsm0uFm5_0),.din(w_dff_A_33gZIik94_0),.clk(gclk));
	jdff dff_A_38Pjr5fa8_0(.dout(w_dff_A_33gZIik94_0),.din(w_dff_A_38Pjr5fa8_0),.clk(gclk));
	jdff dff_B_8A802oyh5_0(.din(n808),.dout(w_dff_B_8A802oyh5_0),.clk(gclk));
	jdff dff_B_OPIUQjYO2_0(.din(w_dff_B_8A802oyh5_0),.dout(w_dff_B_OPIUQjYO2_0),.clk(gclk));
	jdff dff_B_VKWfFFBw6_0(.din(w_dff_B_OPIUQjYO2_0),.dout(w_dff_B_VKWfFFBw6_0),.clk(gclk));
	jdff dff_B_3alZRvZ45_0(.din(w_dff_B_VKWfFFBw6_0),.dout(w_dff_B_3alZRvZ45_0),.clk(gclk));
	jdff dff_B_ZsBQnEA47_0(.din(w_dff_B_3alZRvZ45_0),.dout(w_dff_B_ZsBQnEA47_0),.clk(gclk));
	jdff dff_B_NPYzj9ey3_0(.din(w_dff_B_ZsBQnEA47_0),.dout(w_dff_B_NPYzj9ey3_0),.clk(gclk));
	jdff dff_B_SESaneVA4_0(.din(w_dff_B_NPYzj9ey3_0),.dout(w_dff_B_SESaneVA4_0),.clk(gclk));
	jdff dff_B_GIU1vtYK0_0(.din(w_dff_B_SESaneVA4_0),.dout(w_dff_B_GIU1vtYK0_0),.clk(gclk));
	jdff dff_B_5IETn2KG4_0(.din(w_dff_B_GIU1vtYK0_0),.dout(w_dff_B_5IETn2KG4_0),.clk(gclk));
	jdff dff_B_oplNXEDL6_0(.din(w_dff_B_5IETn2KG4_0),.dout(w_dff_B_oplNXEDL6_0),.clk(gclk));
	jdff dff_B_1PScmEgp4_0(.din(n803),.dout(w_dff_B_1PScmEgp4_0),.clk(gclk));
	jdff dff_A_c8nKUhZi0_1(.dout(w_n797_9[1]),.din(w_dff_A_c8nKUhZi0_1),.clk(gclk));
	jdff dff_A_seo738dG0_1(.dout(w_dff_A_c8nKUhZi0_1),.din(w_dff_A_seo738dG0_1),.clk(gclk));
	jdff dff_A_HOayV5bp4_1(.dout(w_dff_A_seo738dG0_1),.din(w_dff_A_HOayV5bp4_1),.clk(gclk));
	jdff dff_A_AjbdDBgO6_1(.dout(w_dff_A_HOayV5bp4_1),.din(w_dff_A_AjbdDBgO6_1),.clk(gclk));
	jdff dff_A_0T4J5fkg1_1(.dout(w_dff_A_AjbdDBgO6_1),.din(w_dff_A_0T4J5fkg1_1),.clk(gclk));
	jdff dff_A_dmjpzGTR8_1(.dout(w_dff_A_0T4J5fkg1_1),.din(w_dff_A_dmjpzGTR8_1),.clk(gclk));
	jdff dff_A_EKuwZTdH8_1(.dout(w_dff_A_dmjpzGTR8_1),.din(w_dff_A_EKuwZTdH8_1),.clk(gclk));
	jdff dff_A_iOrnd5Pj3_1(.dout(w_dff_A_EKuwZTdH8_1),.din(w_dff_A_iOrnd5Pj3_1),.clk(gclk));
	jdff dff_A_zISZqvFC3_1(.dout(w_dff_A_iOrnd5Pj3_1),.din(w_dff_A_zISZqvFC3_1),.clk(gclk));
	jdff dff_A_losgSMuX1_1(.dout(w_dff_A_zISZqvFC3_1),.din(w_dff_A_losgSMuX1_1),.clk(gclk));
	jdff dff_B_t0Lv9bLg5_0(.din(n861),.dout(w_dff_B_t0Lv9bLg5_0),.clk(gclk));
	jdff dff_B_IY6zNTzk1_0(.din(w_dff_B_t0Lv9bLg5_0),.dout(w_dff_B_IY6zNTzk1_0),.clk(gclk));
	jdff dff_B_Y1Crni0n0_0(.din(w_dff_B_IY6zNTzk1_0),.dout(w_dff_B_Y1Crni0n0_0),.clk(gclk));
	jdff dff_B_2lQCkvPH6_0(.din(w_dff_B_Y1Crni0n0_0),.dout(w_dff_B_2lQCkvPH6_0),.clk(gclk));
	jdff dff_B_DwmqAbxu1_0(.din(w_dff_B_2lQCkvPH6_0),.dout(w_dff_B_DwmqAbxu1_0),.clk(gclk));
	jdff dff_B_yO2Ld9hd1_0(.din(w_dff_B_DwmqAbxu1_0),.dout(w_dff_B_yO2Ld9hd1_0),.clk(gclk));
	jdff dff_B_Wm19bM8k6_0(.din(w_dff_B_yO2Ld9hd1_0),.dout(w_dff_B_Wm19bM8k6_0),.clk(gclk));
	jdff dff_B_CCcAZDDj1_0(.din(w_dff_B_Wm19bM8k6_0),.dout(w_dff_B_CCcAZDDj1_0),.clk(gclk));
	jdff dff_B_IdQgVWDq7_0(.din(w_dff_B_CCcAZDDj1_0),.dout(w_dff_B_IdQgVWDq7_0),.clk(gclk));
	jdff dff_B_ka2cL7cq3_0(.din(w_dff_B_IdQgVWDq7_0),.dout(w_dff_B_ka2cL7cq3_0),.clk(gclk));
	jdff dff_B_5Pi8sLZf6_2(.din(G61),.dout(w_dff_B_5Pi8sLZf6_2),.clk(gclk));
	jdff dff_B_Zj1aWoW30_0(.din(n856),.dout(w_dff_B_Zj1aWoW30_0),.clk(gclk));
	jdff dff_A_aRXDzq5t5_1(.dout(w_n852_9[1]),.din(w_dff_A_aRXDzq5t5_1),.clk(gclk));
	jdff dff_A_54vCDj965_1(.dout(w_dff_A_aRXDzq5t5_1),.din(w_dff_A_54vCDj965_1),.clk(gclk));
	jdff dff_A_Tjsbs8C07_1(.dout(w_dff_A_54vCDj965_1),.din(w_dff_A_Tjsbs8C07_1),.clk(gclk));
	jdff dff_A_DjrPyRvT1_1(.dout(w_dff_A_Tjsbs8C07_1),.din(w_dff_A_DjrPyRvT1_1),.clk(gclk));
	jdff dff_A_RFF4a3Id4_1(.dout(w_dff_A_DjrPyRvT1_1),.din(w_dff_A_RFF4a3Id4_1),.clk(gclk));
	jdff dff_A_MGMIOyFU5_1(.dout(w_dff_A_RFF4a3Id4_1),.din(w_dff_A_MGMIOyFU5_1),.clk(gclk));
	jdff dff_A_SmllZ8dT6_1(.dout(w_dff_A_MGMIOyFU5_1),.din(w_dff_A_SmllZ8dT6_1),.clk(gclk));
	jdff dff_A_R7B2ihJO3_1(.dout(w_dff_A_SmllZ8dT6_1),.din(w_dff_A_R7B2ihJO3_1),.clk(gclk));
	jdff dff_A_Q5mkiUxB4_1(.dout(w_dff_A_R7B2ihJO3_1),.din(w_dff_A_Q5mkiUxB4_1),.clk(gclk));
	jdff dff_A_GStFKiis3_1(.dout(w_dff_A_Q5mkiUxB4_1),.din(w_dff_A_GStFKiis3_1),.clk(gclk));
	jdff dff_B_ifnOJc1U1_0(.din(n967),.dout(w_dff_B_ifnOJc1U1_0),.clk(gclk));
	jdff dff_B_ynuAR34F0_1(.din(n961),.dout(w_dff_B_ynuAR34F0_1),.clk(gclk));
	jdff dff_B_bZ4GVU5u1_1(.din(w_dff_B_ynuAR34F0_1),.dout(w_dff_B_bZ4GVU5u1_1),.clk(gclk));
	jdff dff_B_nTaXBT9q0_1(.din(w_dff_B_bZ4GVU5u1_1),.dout(w_dff_B_nTaXBT9q0_1),.clk(gclk));
	jdff dff_B_iqLddp8R8_0(.din(n960),.dout(w_dff_B_iqLddp8R8_0),.clk(gclk));
	jdff dff_B_a6qgBGCl0_1(.din(n975),.dout(w_dff_B_a6qgBGCl0_1),.clk(gclk));
	jdff dff_B_cm89qgb02_1(.din(w_dff_B_a6qgBGCl0_1),.dout(w_dff_B_cm89qgb02_1),.clk(gclk));
	jdff dff_B_Y4rYfPA96_1(.din(w_dff_B_cm89qgb02_1),.dout(w_dff_B_Y4rYfPA96_1),.clk(gclk));
	jdff dff_B_qLpZPYUP7_1(.din(w_dff_B_Y4rYfPA96_1),.dout(w_dff_B_qLpZPYUP7_1),.clk(gclk));
	jdff dff_B_AxD9PwDr3_1(.din(w_dff_B_qLpZPYUP7_1),.dout(w_dff_B_AxD9PwDr3_1),.clk(gclk));
	jdff dff_B_0mYtizdg0_1(.din(n971),.dout(w_dff_B_0mYtizdg0_1),.clk(gclk));
	jdff dff_B_CpVbdhlH2_1(.din(w_dff_B_0mYtizdg0_1),.dout(w_dff_B_CpVbdhlH2_1),.clk(gclk));
	jdff dff_B_rpc69Qrr7_1(.din(n995),.dout(w_dff_B_rpc69Qrr7_1),.clk(gclk));
	jdff dff_B_jNILjL1c7_1(.din(w_dff_B_rpc69Qrr7_1),.dout(w_dff_B_jNILjL1c7_1),.clk(gclk));
	jdff dff_B_M9tgOfoG7_1(.din(w_dff_B_jNILjL1c7_1),.dout(w_dff_B_M9tgOfoG7_1),.clk(gclk));
	jdff dff_B_iFErXtgI2_1(.din(w_dff_B_M9tgOfoG7_1),.dout(w_dff_B_iFErXtgI2_1),.clk(gclk));
	jdff dff_B_emGytDbn3_1(.din(w_dff_B_iFErXtgI2_1),.dout(w_dff_B_emGytDbn3_1),.clk(gclk));
	jdff dff_B_2fWqJBgV3_1(.din(w_dff_B_emGytDbn3_1),.dout(w_dff_B_2fWqJBgV3_1),.clk(gclk));
	jdff dff_B_YPTvsFTT1_1(.din(w_dff_B_2fWqJBgV3_1),.dout(w_dff_B_YPTvsFTT1_1),.clk(gclk));
	jdff dff_B_xOad4M3p8_1(.din(w_dff_B_YPTvsFTT1_1),.dout(w_dff_B_xOad4M3p8_1),.clk(gclk));
	jdff dff_B_fHaFuXNL2_1(.din(w_dff_B_xOad4M3p8_1),.dout(w_dff_B_fHaFuXNL2_1),.clk(gclk));
	jdff dff_B_WddvAmdt9_1(.din(w_dff_B_fHaFuXNL2_1),.dout(w_dff_B_WddvAmdt9_1),.clk(gclk));
	jdff dff_B_bIlR0n4s5_1(.din(w_dff_B_WddvAmdt9_1),.dout(w_dff_B_bIlR0n4s5_1),.clk(gclk));
	jdff dff_B_bepvfav89_1(.din(n997),.dout(w_dff_B_bepvfav89_1),.clk(gclk));
	jdff dff_B_PmBeLX548_1(.din(w_dff_B_bepvfav89_1),.dout(w_dff_B_PmBeLX548_1),.clk(gclk));
	jdff dff_B_rzfiyyni7_1(.din(w_dff_B_PmBeLX548_1),.dout(w_dff_B_rzfiyyni7_1),.clk(gclk));
	jdff dff_B_KQ2RIcrD9_1(.din(w_dff_B_rzfiyyni7_1),.dout(w_dff_B_KQ2RIcrD9_1),.clk(gclk));
	jdff dff_B_wEc3UVnu1_1(.din(w_dff_B_KQ2RIcrD9_1),.dout(w_dff_B_wEc3UVnu1_1),.clk(gclk));
	jdff dff_B_oAnQ5GPc4_1(.din(w_dff_B_wEc3UVnu1_1),.dout(w_dff_B_oAnQ5GPc4_1),.clk(gclk));
	jdff dff_B_3BuDIKdG0_1(.din(w_dff_B_oAnQ5GPc4_1),.dout(w_dff_B_3BuDIKdG0_1),.clk(gclk));
	jdff dff_B_GQUnHn8g1_1(.din(w_dff_B_3BuDIKdG0_1),.dout(w_dff_B_GQUnHn8g1_1),.clk(gclk));
	jdff dff_B_eqL0ZiLh0_1(.din(w_dff_B_GQUnHn8g1_1),.dout(w_dff_B_eqL0ZiLh0_1),.clk(gclk));
	jdff dff_B_pBC8bezt1_1(.din(w_dff_B_eqL0ZiLh0_1),.dout(w_dff_B_pBC8bezt1_1),.clk(gclk));
	jdff dff_B_zadYHcFr1_1(.din(w_dff_B_pBC8bezt1_1),.dout(w_dff_B_zadYHcFr1_1),.clk(gclk));
	jdff dff_B_gGhJvAVX2_0(.din(n1001),.dout(w_dff_B_gGhJvAVX2_0),.clk(gclk));
	jdff dff_B_YFsucXNK3_0(.din(n1016),.dout(w_dff_B_YFsucXNK3_0),.clk(gclk));
	jdff dff_B_NX7qa5h72_0(.din(w_dff_B_YFsucXNK3_0),.dout(w_dff_B_NX7qa5h72_0),.clk(gclk));
	jdff dff_B_yX0JgzqU5_0(.din(w_dff_B_NX7qa5h72_0),.dout(w_dff_B_yX0JgzqU5_0),.clk(gclk));
	jdff dff_B_P8VxAMFw6_0(.din(w_dff_B_yX0JgzqU5_0),.dout(w_dff_B_P8VxAMFw6_0),.clk(gclk));
	jdff dff_B_hu4syHSm8_0(.din(w_dff_B_P8VxAMFw6_0),.dout(w_dff_B_hu4syHSm8_0),.clk(gclk));
	jdff dff_B_JB8MMbPs8_0(.din(w_dff_B_hu4syHSm8_0),.dout(w_dff_B_JB8MMbPs8_0),.clk(gclk));
	jdff dff_B_LsuiAY8o2_0(.din(w_dff_B_JB8MMbPs8_0),.dout(w_dff_B_LsuiAY8o2_0),.clk(gclk));
	jdff dff_B_6zHzrdVX2_0(.din(w_dff_B_LsuiAY8o2_0),.dout(w_dff_B_6zHzrdVX2_0),.clk(gclk));
	jdff dff_B_V17nTjdJ3_0(.din(w_dff_B_6zHzrdVX2_0),.dout(w_dff_B_V17nTjdJ3_0),.clk(gclk));
	jdff dff_B_Ma1gKVog9_0(.din(w_dff_B_V17nTjdJ3_0),.dout(w_dff_B_Ma1gKVog9_0),.clk(gclk));
	jdff dff_B_s0XwuCNn0_1(.din(n1013),.dout(w_dff_B_s0XwuCNn0_1),.clk(gclk));
	jdff dff_B_TEwl3wgg6_2(.din(G182),.dout(w_dff_B_TEwl3wgg6_2),.clk(gclk));
	jdff dff_B_UXYvnfD98_2(.din(w_dff_B_TEwl3wgg6_2),.dout(w_dff_B_UXYvnfD98_2),.clk(gclk));
	jdff dff_B_cX4vbk7M7_2(.din(G185),.dout(w_dff_B_cX4vbk7M7_2),.clk(gclk));
	jdff dff_B_TH3AsybK0_1(.din(n1006),.dout(w_dff_B_TH3AsybK0_1),.clk(gclk));
	jdff dff_B_pJs3TDkA4_1(.din(w_dff_B_TH3AsybK0_1),.dout(w_dff_B_pJs3TDkA4_1),.clk(gclk));
	jdff dff_B_PSJp4qRu8_1(.din(w_dff_B_pJs3TDkA4_1),.dout(w_dff_B_PSJp4qRu8_1),.clk(gclk));
	jdff dff_B_llc5HBxt6_1(.din(n777),.dout(w_dff_B_llc5HBxt6_1),.clk(gclk));
	jdff dff_B_tPDLTsEY6_1(.din(w_dff_B_llc5HBxt6_1),.dout(w_dff_B_tPDLTsEY6_1),.clk(gclk));
	jdff dff_B_X4NEc9x47_1(.din(w_dff_B_tPDLTsEY6_1),.dout(w_dff_B_X4NEc9x47_1),.clk(gclk));
	jdff dff_B_7H31U1To0_1(.din(w_dff_B_X4NEc9x47_1),.dout(w_dff_B_7H31U1To0_1),.clk(gclk));
	jdff dff_B_0fwNjf782_1(.din(w_dff_B_7H31U1To0_1),.dout(w_dff_B_0fwNjf782_1),.clk(gclk));
	jdff dff_B_kwHGDFZX7_0(.din(n782),.dout(w_dff_B_kwHGDFZX7_0),.clk(gclk));
	jdff dff_B_u9pdidx38_1(.din(n536),.dout(w_dff_B_u9pdidx38_1),.clk(gclk));
	jdff dff_B_3XLwB3kW2_1(.din(n531),.dout(w_dff_B_3XLwB3kW2_1),.clk(gclk));
	jdff dff_A_0kNBMird8_0(.dout(w_n779_0[0]),.din(w_dff_A_0kNBMird8_0),.clk(gclk));
	jdff dff_A_qnGRR56D9_0(.dout(w_dff_A_0kNBMird8_0),.din(w_dff_A_qnGRR56D9_0),.clk(gclk));
	jdff dff_B_llH03iJn7_1(.din(G117),.dout(w_dff_B_llH03iJn7_1),.clk(gclk));
	jdff dff_B_uWQdhYHv7_1(.din(w_dff_B_llH03iJn7_1),.dout(w_dff_B_uWQdhYHv7_1),.clk(gclk));
	jdff dff_B_OT9KcLqn4_1(.din(n752),.dout(w_dff_B_OT9KcLqn4_1),.clk(gclk));
	jdff dff_B_GrmjhGxS4_1(.din(w_dff_B_OT9KcLqn4_1),.dout(w_dff_B_GrmjhGxS4_1),.clk(gclk));
	jdff dff_B_Wr6GDBT12_1(.din(w_dff_B_GrmjhGxS4_1),.dout(w_dff_B_Wr6GDBT12_1),.clk(gclk));
	jdff dff_A_3ZG8IpOA9_0(.dout(w_n755_0[0]),.din(w_dff_A_3ZG8IpOA9_0),.clk(gclk));
	jdff dff_A_68n6HSoo1_0(.dout(w_dff_A_3ZG8IpOA9_0),.din(w_dff_A_68n6HSoo1_0),.clk(gclk));
	jdff dff_A_ATfgVxmz3_0(.dout(w_dff_A_68n6HSoo1_0),.din(w_dff_A_ATfgVxmz3_0),.clk(gclk));
	jdff dff_A_pJggtBVe3_0(.dout(w_dff_A_ATfgVxmz3_0),.din(w_dff_A_pJggtBVe3_0),.clk(gclk));
	jdff dff_A_FkQn2sEm6_0(.dout(w_dff_A_pJggtBVe3_0),.din(w_dff_A_FkQn2sEm6_0),.clk(gclk));
	jdff dff_A_MJ8r3R6z6_0(.dout(w_dff_A_FkQn2sEm6_0),.din(w_dff_A_MJ8r3R6z6_0),.clk(gclk));
	jdff dff_A_DDxqCbB22_0(.dout(w_dff_A_MJ8r3R6z6_0),.din(w_dff_A_DDxqCbB22_0),.clk(gclk));
	jdff dff_A_9lKhqlHn3_0(.dout(w_dff_A_DDxqCbB22_0),.din(w_dff_A_9lKhqlHn3_0),.clk(gclk));
	jdff dff_A_biLyGV7G6_0(.dout(w_dff_A_9lKhqlHn3_0),.din(w_dff_A_biLyGV7G6_0),.clk(gclk));
	jdff dff_A_HR22AKG65_0(.dout(w_dff_A_biLyGV7G6_0),.din(w_dff_A_HR22AKG65_0),.clk(gclk));
	jdff dff_A_AFcJoeIn8_0(.dout(w_dff_A_HR22AKG65_0),.din(w_dff_A_AFcJoeIn8_0),.clk(gclk));
	jdff dff_B_VjocPBUU2_1(.din(G131),.dout(w_dff_B_VjocPBUU2_1),.clk(gclk));
	jdff dff_B_5JNCKSIB9_1(.din(w_dff_B_VjocPBUU2_1),.dout(w_dff_B_5JNCKSIB9_1),.clk(gclk));
	jdff dff_B_6C7xYPwX4_0(.din(n1028),.dout(w_dff_B_6C7xYPwX4_0),.clk(gclk));
	jdff dff_B_6usAEpL71_0(.din(w_dff_B_6C7xYPwX4_0),.dout(w_dff_B_6usAEpL71_0),.clk(gclk));
	jdff dff_B_DPoBePda6_0(.din(w_dff_B_6usAEpL71_0),.dout(w_dff_B_DPoBePda6_0),.clk(gclk));
	jdff dff_B_p43uRxwh4_0(.din(w_dff_B_DPoBePda6_0),.dout(w_dff_B_p43uRxwh4_0),.clk(gclk));
	jdff dff_B_PXHs6AVa0_0(.din(w_dff_B_p43uRxwh4_0),.dout(w_dff_B_PXHs6AVa0_0),.clk(gclk));
	jdff dff_B_NCJWC3Zs6_0(.din(w_dff_B_PXHs6AVa0_0),.dout(w_dff_B_NCJWC3Zs6_0),.clk(gclk));
	jdff dff_B_C9UyJnCz3_0(.din(w_dff_B_NCJWC3Zs6_0),.dout(w_dff_B_C9UyJnCz3_0),.clk(gclk));
	jdff dff_B_nT9GyZhR6_0(.din(w_dff_B_C9UyJnCz3_0),.dout(w_dff_B_nT9GyZhR6_0),.clk(gclk));
	jdff dff_B_4kE6BgE56_0(.din(w_dff_B_nT9GyZhR6_0),.dout(w_dff_B_4kE6BgE56_0),.clk(gclk));
	jdff dff_B_GmDFS35I0_0(.din(w_dff_B_4kE6BgE56_0),.dout(w_dff_B_GmDFS35I0_0),.clk(gclk));
	jdff dff_B_VSsnlerl0_0(.din(w_dff_B_GmDFS35I0_0),.dout(w_dff_B_VSsnlerl0_0),.clk(gclk));
	jdff dff_B_SCP58RGa4_0(.din(w_dff_B_VSsnlerl0_0),.dout(w_dff_B_SCP58RGa4_0),.clk(gclk));
	jdff dff_B_017KG9S71_0(.din(w_dff_B_SCP58RGa4_0),.dout(w_dff_B_017KG9S71_0),.clk(gclk));
	jdff dff_B_9ldMJKpa4_0(.din(w_dff_B_017KG9S71_0),.dout(w_dff_B_9ldMJKpa4_0),.clk(gclk));
	jdff dff_B_qmgLwixf3_0(.din(w_dff_B_9ldMJKpa4_0),.dout(w_dff_B_qmgLwixf3_0),.clk(gclk));
	jdff dff_B_UIq314s07_0(.din(w_dff_B_qmgLwixf3_0),.dout(w_dff_B_UIq314s07_0),.clk(gclk));
	jdff dff_B_IsG2THwt3_1(.din(n1020),.dout(w_dff_B_IsG2THwt3_1),.clk(gclk));
	jdff dff_A_TZScAyTj2_0(.dout(w_n800_4[0]),.din(w_dff_A_TZScAyTj2_0),.clk(gclk));
	jdff dff_A_QNrzqIJH1_0(.dout(w_dff_A_TZScAyTj2_0),.din(w_dff_A_QNrzqIJH1_0),.clk(gclk));
	jdff dff_A_9hnClhKi8_0(.dout(w_dff_A_QNrzqIJH1_0),.din(w_dff_A_9hnClhKi8_0),.clk(gclk));
	jdff dff_A_L0En3HXn6_0(.dout(w_dff_A_9hnClhKi8_0),.din(w_dff_A_L0En3HXn6_0),.clk(gclk));
	jdff dff_A_3K82hbXV2_0(.dout(w_dff_A_L0En3HXn6_0),.din(w_dff_A_3K82hbXV2_0),.clk(gclk));
	jdff dff_A_OpI0ot5M8_0(.dout(w_dff_A_3K82hbXV2_0),.din(w_dff_A_OpI0ot5M8_0),.clk(gclk));
	jdff dff_A_zylMXVli7_0(.dout(w_dff_A_OpI0ot5M8_0),.din(w_dff_A_zylMXVli7_0),.clk(gclk));
	jdff dff_B_Po2ISzVd5_0(.din(n1039),.dout(w_dff_B_Po2ISzVd5_0),.clk(gclk));
	jdff dff_B_ZRmtmCjC7_0(.din(w_dff_B_Po2ISzVd5_0),.dout(w_dff_B_ZRmtmCjC7_0),.clk(gclk));
	jdff dff_B_hTIicSsr5_0(.din(w_dff_B_ZRmtmCjC7_0),.dout(w_dff_B_hTIicSsr5_0),.clk(gclk));
	jdff dff_B_mTUB5HaQ7_0(.din(w_dff_B_hTIicSsr5_0),.dout(w_dff_B_mTUB5HaQ7_0),.clk(gclk));
	jdff dff_B_7hy4n0E68_0(.din(w_dff_B_mTUB5HaQ7_0),.dout(w_dff_B_7hy4n0E68_0),.clk(gclk));
	jdff dff_B_otWUI5sG6_0(.din(w_dff_B_7hy4n0E68_0),.dout(w_dff_B_otWUI5sG6_0),.clk(gclk));
	jdff dff_B_XS6BAxRR8_0(.din(w_dff_B_otWUI5sG6_0),.dout(w_dff_B_XS6BAxRR8_0),.clk(gclk));
	jdff dff_B_HaHF3kcj8_0(.din(w_dff_B_XS6BAxRR8_0),.dout(w_dff_B_HaHF3kcj8_0),.clk(gclk));
	jdff dff_B_ZyqN2vLL3_0(.din(w_dff_B_HaHF3kcj8_0),.dout(w_dff_B_ZyqN2vLL3_0),.clk(gclk));
	jdff dff_B_qYCT38415_0(.din(w_dff_B_ZyqN2vLL3_0),.dout(w_dff_B_qYCT38415_0),.clk(gclk));
	jdff dff_B_p8auc4tf7_0(.din(w_dff_B_qYCT38415_0),.dout(w_dff_B_p8auc4tf7_0),.clk(gclk));
	jdff dff_B_fqGVN7Vg8_0(.din(w_dff_B_p8auc4tf7_0),.dout(w_dff_B_fqGVN7Vg8_0),.clk(gclk));
	jdff dff_B_DXGhJf8M6_0(.din(w_dff_B_fqGVN7Vg8_0),.dout(w_dff_B_DXGhJf8M6_0),.clk(gclk));
	jdff dff_B_uKusfTFG7_0(.din(w_dff_B_DXGhJf8M6_0),.dout(w_dff_B_uKusfTFG7_0),.clk(gclk));
	jdff dff_B_EmJXUkSS3_0(.din(w_dff_B_uKusfTFG7_0),.dout(w_dff_B_EmJXUkSS3_0),.clk(gclk));
	jdff dff_B_QvF7cfS06_1(.din(n1031),.dout(w_dff_B_QvF7cfS06_1),.clk(gclk));
	jdff dff_B_JNeHI5JZ0_1(.din(w_dff_B_QvF7cfS06_1),.dout(w_dff_B_JNeHI5JZ0_1),.clk(gclk));
	jdff dff_A_MQEkn3ZQ3_0(.dout(w_G4088_8[0]),.din(w_dff_A_MQEkn3ZQ3_0),.clk(gclk));
	jdff dff_A_8JSkwwNG0_0(.dout(w_dff_A_MQEkn3ZQ3_0),.din(w_dff_A_8JSkwwNG0_0),.clk(gclk));
	jdff dff_A_SD5aRq3n2_0(.dout(w_dff_A_8JSkwwNG0_0),.din(w_dff_A_SD5aRq3n2_0),.clk(gclk));
	jdff dff_A_yHlDPozQ3_0(.dout(w_dff_A_SD5aRq3n2_0),.din(w_dff_A_yHlDPozQ3_0),.clk(gclk));
	jdff dff_A_KIAw0P6t3_0(.dout(w_dff_A_yHlDPozQ3_0),.din(w_dff_A_KIAw0P6t3_0),.clk(gclk));
	jdff dff_A_tJYE0Yn30_0(.dout(w_dff_A_KIAw0P6t3_0),.din(w_dff_A_tJYE0Yn30_0),.clk(gclk));
	jdff dff_A_6uxWNdtr7_0(.dout(w_dff_A_tJYE0Yn30_0),.din(w_dff_A_6uxWNdtr7_0),.clk(gclk));
	jdff dff_A_UZllMLiM0_0(.dout(w_dff_A_6uxWNdtr7_0),.din(w_dff_A_UZllMLiM0_0),.clk(gclk));
	jdff dff_A_t1A3h8wG4_0(.dout(w_dff_A_UZllMLiM0_0),.din(w_dff_A_t1A3h8wG4_0),.clk(gclk));
	jdff dff_A_Vrkc4mDz8_0(.dout(w_dff_A_t1A3h8wG4_0),.din(w_dff_A_Vrkc4mDz8_0),.clk(gclk));
	jdff dff_A_pjGbuDnr6_0(.dout(w_dff_A_Vrkc4mDz8_0),.din(w_dff_A_pjGbuDnr6_0),.clk(gclk));
	jdff dff_A_Cp83xP6V3_0(.dout(w_dff_A_pjGbuDnr6_0),.din(w_dff_A_Cp83xP6V3_0),.clk(gclk));
	jdff dff_A_Cqi6r2G91_0(.dout(w_dff_A_Cp83xP6V3_0),.din(w_dff_A_Cqi6r2G91_0),.clk(gclk));
	jdff dff_A_PyUVJ6Sk0_0(.dout(w_dff_A_Cqi6r2G91_0),.din(w_dff_A_PyUVJ6Sk0_0),.clk(gclk));
	jdff dff_A_p986CboN5_0(.dout(w_dff_A_PyUVJ6Sk0_0),.din(w_dff_A_p986CboN5_0),.clk(gclk));
	jdff dff_A_6a5PsfXW0_2(.dout(w_G4088_8[2]),.din(w_dff_A_6a5PsfXW0_2),.clk(gclk));
	jdff dff_A_XA8MWyHc0_2(.dout(w_dff_A_6a5PsfXW0_2),.din(w_dff_A_XA8MWyHc0_2),.clk(gclk));
	jdff dff_A_8kFdNVLW4_2(.dout(w_dff_A_XA8MWyHc0_2),.din(w_dff_A_8kFdNVLW4_2),.clk(gclk));
	jdff dff_A_5wl5X6Qu4_2(.dout(w_dff_A_8kFdNVLW4_2),.din(w_dff_A_5wl5X6Qu4_2),.clk(gclk));
	jdff dff_A_2uSKnKuM9_2(.dout(w_dff_A_5wl5X6Qu4_2),.din(w_dff_A_2uSKnKuM9_2),.clk(gclk));
	jdff dff_A_OXGEE86E0_2(.dout(w_dff_A_2uSKnKuM9_2),.din(w_dff_A_OXGEE86E0_2),.clk(gclk));
	jdff dff_A_KFXFmrLM3_2(.dout(w_dff_A_OXGEE86E0_2),.din(w_dff_A_KFXFmrLM3_2),.clk(gclk));
	jdff dff_A_DkQQXndv4_2(.dout(w_dff_A_KFXFmrLM3_2),.din(w_dff_A_DkQQXndv4_2),.clk(gclk));
	jdff dff_A_yxXdYlDR6_2(.dout(w_dff_A_DkQQXndv4_2),.din(w_dff_A_yxXdYlDR6_2),.clk(gclk));
	jdff dff_A_iG2oJDo61_2(.dout(w_dff_A_yxXdYlDR6_2),.din(w_dff_A_iG2oJDo61_2),.clk(gclk));
	jdff dff_A_uGZtE6xb4_2(.dout(w_dff_A_iG2oJDo61_2),.din(w_dff_A_uGZtE6xb4_2),.clk(gclk));
	jdff dff_A_m8qufn2Y3_2(.dout(w_dff_A_uGZtE6xb4_2),.din(w_dff_A_m8qufn2Y3_2),.clk(gclk));
	jdff dff_A_3jfaWwH20_2(.dout(w_dff_A_m8qufn2Y3_2),.din(w_dff_A_3jfaWwH20_2),.clk(gclk));
	jdff dff_A_W5PlwJbf8_2(.dout(w_dff_A_3jfaWwH20_2),.din(w_dff_A_W5PlwJbf8_2),.clk(gclk));
	jdff dff_A_qaMVEAhk2_2(.dout(w_dff_A_W5PlwJbf8_2),.din(w_dff_A_qaMVEAhk2_2),.clk(gclk));
	jdff dff_A_FgbyN03F3_2(.dout(w_dff_A_qaMVEAhk2_2),.din(w_dff_A_FgbyN03F3_2),.clk(gclk));
	jdff dff_A_VvG59TxG9_0(.dout(w_n797_8[0]),.din(w_dff_A_VvG59TxG9_0),.clk(gclk));
	jdff dff_A_rzUZXHyG7_0(.dout(w_dff_A_VvG59TxG9_0),.din(w_dff_A_rzUZXHyG7_0),.clk(gclk));
	jdff dff_A_nuSZUysl8_0(.dout(w_dff_A_rzUZXHyG7_0),.din(w_dff_A_nuSZUysl8_0),.clk(gclk));
	jdff dff_A_OadZqIXw7_0(.dout(w_dff_A_nuSZUysl8_0),.din(w_dff_A_OadZqIXw7_0),.clk(gclk));
	jdff dff_A_k39D8FCz7_0(.dout(w_dff_A_OadZqIXw7_0),.din(w_dff_A_k39D8FCz7_0),.clk(gclk));
	jdff dff_A_wQb28WFR7_0(.dout(w_dff_A_k39D8FCz7_0),.din(w_dff_A_wQb28WFR7_0),.clk(gclk));
	jdff dff_A_Kpw8bXjQ3_0(.dout(w_dff_A_wQb28WFR7_0),.din(w_dff_A_Kpw8bXjQ3_0),.clk(gclk));
	jdff dff_A_21fj1h7t2_0(.dout(w_dff_A_Kpw8bXjQ3_0),.din(w_dff_A_21fj1h7t2_0),.clk(gclk));
	jdff dff_A_OayhSrbs8_0(.dout(w_dff_A_21fj1h7t2_0),.din(w_dff_A_OayhSrbs8_0),.clk(gclk));
	jdff dff_A_Uj7yy23O6_0(.dout(w_dff_A_OayhSrbs8_0),.din(w_dff_A_Uj7yy23O6_0),.clk(gclk));
	jdff dff_A_0VW1blZh0_0(.dout(w_dff_A_Uj7yy23O6_0),.din(w_dff_A_0VW1blZh0_0),.clk(gclk));
	jdff dff_A_aBn7HYKn3_0(.dout(w_dff_A_0VW1blZh0_0),.din(w_dff_A_aBn7HYKn3_0),.clk(gclk));
	jdff dff_A_RMKQ9xKZ3_0(.dout(w_dff_A_aBn7HYKn3_0),.din(w_dff_A_RMKQ9xKZ3_0),.clk(gclk));
	jdff dff_A_wMSaZ8gK4_2(.dout(w_n797_8[2]),.din(w_dff_A_wMSaZ8gK4_2),.clk(gclk));
	jdff dff_A_W6bTy4494_2(.dout(w_dff_A_wMSaZ8gK4_2),.din(w_dff_A_W6bTy4494_2),.clk(gclk));
	jdff dff_A_lKCBf1TV2_2(.dout(w_dff_A_W6bTy4494_2),.din(w_dff_A_lKCBf1TV2_2),.clk(gclk));
	jdff dff_A_CIauddfq1_2(.dout(w_dff_A_lKCBf1TV2_2),.din(w_dff_A_CIauddfq1_2),.clk(gclk));
	jdff dff_A_6YOhI7Sq3_2(.dout(w_dff_A_CIauddfq1_2),.din(w_dff_A_6YOhI7Sq3_2),.clk(gclk));
	jdff dff_A_IKtUNxUx4_2(.dout(w_dff_A_6YOhI7Sq3_2),.din(w_dff_A_IKtUNxUx4_2),.clk(gclk));
	jdff dff_A_FrqyaWoV3_2(.dout(w_dff_A_IKtUNxUx4_2),.din(w_dff_A_FrqyaWoV3_2),.clk(gclk));
	jdff dff_A_8v3wnTHs3_2(.dout(w_dff_A_FrqyaWoV3_2),.din(w_dff_A_8v3wnTHs3_2),.clk(gclk));
	jdff dff_A_zbAwwr7D1_2(.dout(w_dff_A_8v3wnTHs3_2),.din(w_dff_A_zbAwwr7D1_2),.clk(gclk));
	jdff dff_A_3GY1SmH09_2(.dout(w_dff_A_zbAwwr7D1_2),.din(w_dff_A_3GY1SmH09_2),.clk(gclk));
	jdff dff_A_WVYYgkO42_2(.dout(w_dff_A_3GY1SmH09_2),.din(w_dff_A_WVYYgkO42_2),.clk(gclk));
	jdff dff_A_h1z21ejw0_2(.dout(w_dff_A_WVYYgkO42_2),.din(w_dff_A_h1z21ejw0_2),.clk(gclk));
	jdff dff_A_oATnb0JV4_2(.dout(w_dff_A_h1z21ejw0_2),.din(w_dff_A_oATnb0JV4_2),.clk(gclk));
	jdff dff_A_yvKF8FNS8_2(.dout(w_dff_A_oATnb0JV4_2),.din(w_dff_A_yvKF8FNS8_2),.clk(gclk));
	jdff dff_A_szCXB5hr2_2(.dout(w_dff_A_yvKF8FNS8_2),.din(w_dff_A_szCXB5hr2_2),.clk(gclk));
	jdff dff_B_K0taASR83_0(.din(n1050),.dout(w_dff_B_K0taASR83_0),.clk(gclk));
	jdff dff_B_fgCIVJWI4_0(.din(w_dff_B_K0taASR83_0),.dout(w_dff_B_fgCIVJWI4_0),.clk(gclk));
	jdff dff_B_Q390yZn54_0(.din(w_dff_B_fgCIVJWI4_0),.dout(w_dff_B_Q390yZn54_0),.clk(gclk));
	jdff dff_B_yjwzU9cr8_0(.din(w_dff_B_Q390yZn54_0),.dout(w_dff_B_yjwzU9cr8_0),.clk(gclk));
	jdff dff_B_t7VcwXUB3_0(.din(w_dff_B_yjwzU9cr8_0),.dout(w_dff_B_t7VcwXUB3_0),.clk(gclk));
	jdff dff_B_kDLvE5YN3_0(.din(w_dff_B_t7VcwXUB3_0),.dout(w_dff_B_kDLvE5YN3_0),.clk(gclk));
	jdff dff_B_WDpM9Pgp1_0(.din(w_dff_B_kDLvE5YN3_0),.dout(w_dff_B_WDpM9Pgp1_0),.clk(gclk));
	jdff dff_B_XiOc0Asl2_0(.din(w_dff_B_WDpM9Pgp1_0),.dout(w_dff_B_XiOc0Asl2_0),.clk(gclk));
	jdff dff_B_peDalsoS3_0(.din(w_dff_B_XiOc0Asl2_0),.dout(w_dff_B_peDalsoS3_0),.clk(gclk));
	jdff dff_B_50vjEcMR2_0(.din(w_dff_B_peDalsoS3_0),.dout(w_dff_B_50vjEcMR2_0),.clk(gclk));
	jdff dff_B_E6G42R591_0(.din(w_dff_B_50vjEcMR2_0),.dout(w_dff_B_E6G42R591_0),.clk(gclk));
	jdff dff_B_7gGHSTfS2_0(.din(w_dff_B_E6G42R591_0),.dout(w_dff_B_7gGHSTfS2_0),.clk(gclk));
	jdff dff_B_5cicOMT37_0(.din(w_dff_B_7gGHSTfS2_0),.dout(w_dff_B_5cicOMT37_0),.clk(gclk));
	jdff dff_B_wp0a28OD5_1(.din(n1042),.dout(w_dff_B_wp0a28OD5_1),.clk(gclk));
	jdff dff_A_Jo3bcgaK9_1(.dout(w_n797_7[1]),.din(w_dff_A_Jo3bcgaK9_1),.clk(gclk));
	jdff dff_A_CDwIySkN4_1(.dout(w_dff_A_Jo3bcgaK9_1),.din(w_dff_A_CDwIySkN4_1),.clk(gclk));
	jdff dff_A_OnXB51Bp8_1(.dout(w_dff_A_CDwIySkN4_1),.din(w_dff_A_OnXB51Bp8_1),.clk(gclk));
	jdff dff_A_M7YEE43P3_1(.dout(w_dff_A_OnXB51Bp8_1),.din(w_dff_A_M7YEE43P3_1),.clk(gclk));
	jdff dff_A_kg6GLHO41_1(.dout(w_dff_A_M7YEE43P3_1),.din(w_dff_A_kg6GLHO41_1),.clk(gclk));
	jdff dff_A_sddRlp4C4_1(.dout(w_dff_A_kg6GLHO41_1),.din(w_dff_A_sddRlp4C4_1),.clk(gclk));
	jdff dff_A_zz3pZw4u9_1(.dout(w_dff_A_sddRlp4C4_1),.din(w_dff_A_zz3pZw4u9_1),.clk(gclk));
	jdff dff_A_4ZzXPOML7_1(.dout(w_dff_A_zz3pZw4u9_1),.din(w_dff_A_4ZzXPOML7_1),.clk(gclk));
	jdff dff_A_b2kEv4le4_1(.dout(w_dff_A_4ZzXPOML7_1),.din(w_dff_A_b2kEv4le4_1),.clk(gclk));
	jdff dff_A_PV1fhr5j4_1(.dout(w_dff_A_b2kEv4le4_1),.din(w_dff_A_PV1fhr5j4_1),.clk(gclk));
	jdff dff_A_ReqLpIV65_1(.dout(w_dff_A_PV1fhr5j4_1),.din(w_dff_A_ReqLpIV65_1),.clk(gclk));
	jdff dff_A_OTCTdaMt9_1(.dout(w_dff_A_ReqLpIV65_1),.din(w_dff_A_OTCTdaMt9_1),.clk(gclk));
	jdff dff_A_0ZF2PpQz8_1(.dout(w_G4088_7[1]),.din(w_dff_A_0ZF2PpQz8_1),.clk(gclk));
	jdff dff_A_dfc0ZRY10_1(.dout(w_dff_A_0ZF2PpQz8_1),.din(w_dff_A_dfc0ZRY10_1),.clk(gclk));
	jdff dff_A_wZfI1sYx5_1(.dout(w_dff_A_dfc0ZRY10_1),.din(w_dff_A_wZfI1sYx5_1),.clk(gclk));
	jdff dff_A_L00xSYiA9_1(.dout(w_dff_A_wZfI1sYx5_1),.din(w_dff_A_L00xSYiA9_1),.clk(gclk));
	jdff dff_A_9hH4qnTQ4_1(.dout(w_dff_A_L00xSYiA9_1),.din(w_dff_A_9hH4qnTQ4_1),.clk(gclk));
	jdff dff_A_lfyjIjk33_1(.dout(w_dff_A_9hH4qnTQ4_1),.din(w_dff_A_lfyjIjk33_1),.clk(gclk));
	jdff dff_A_KwGtuKwl6_1(.dout(w_dff_A_lfyjIjk33_1),.din(w_dff_A_KwGtuKwl6_1),.clk(gclk));
	jdff dff_A_rDygWqJN8_1(.dout(w_dff_A_KwGtuKwl6_1),.din(w_dff_A_rDygWqJN8_1),.clk(gclk));
	jdff dff_A_S0JEouFS1_1(.dout(w_dff_A_rDygWqJN8_1),.din(w_dff_A_S0JEouFS1_1),.clk(gclk));
	jdff dff_A_kWWrLE427_1(.dout(w_dff_A_S0JEouFS1_1),.din(w_dff_A_kWWrLE427_1),.clk(gclk));
	jdff dff_A_mipak4EX4_1(.dout(w_dff_A_kWWrLE427_1),.din(w_dff_A_mipak4EX4_1),.clk(gclk));
	jdff dff_A_z1tFrmCv4_1(.dout(w_dff_A_mipak4EX4_1),.din(w_dff_A_z1tFrmCv4_1),.clk(gclk));
	jdff dff_A_J40c4J9p9_1(.dout(w_dff_A_z1tFrmCv4_1),.din(w_dff_A_J40c4J9p9_1),.clk(gclk));
	jdff dff_B_WvLGDAOl0_0(.din(n1061),.dout(w_dff_B_WvLGDAOl0_0),.clk(gclk));
	jdff dff_B_OdkadJJI6_0(.din(w_dff_B_WvLGDAOl0_0),.dout(w_dff_B_OdkadJJI6_0),.clk(gclk));
	jdff dff_B_CmNxNxjB0_0(.din(w_dff_B_OdkadJJI6_0),.dout(w_dff_B_CmNxNxjB0_0),.clk(gclk));
	jdff dff_B_oBXown095_0(.din(w_dff_B_CmNxNxjB0_0),.dout(w_dff_B_oBXown095_0),.clk(gclk));
	jdff dff_B_cCeYb6eM9_0(.din(w_dff_B_oBXown095_0),.dout(w_dff_B_cCeYb6eM9_0),.clk(gclk));
	jdff dff_B_JQWwtTVl8_0(.din(w_dff_B_cCeYb6eM9_0),.dout(w_dff_B_JQWwtTVl8_0),.clk(gclk));
	jdff dff_B_nUqsHqs90_0(.din(w_dff_B_JQWwtTVl8_0),.dout(w_dff_B_nUqsHqs90_0),.clk(gclk));
	jdff dff_B_ml71n9Iu4_0(.din(w_dff_B_nUqsHqs90_0),.dout(w_dff_B_ml71n9Iu4_0),.clk(gclk));
	jdff dff_B_Y1IV97me7_0(.din(w_dff_B_ml71n9Iu4_0),.dout(w_dff_B_Y1IV97me7_0),.clk(gclk));
	jdff dff_B_yL46Ax4v3_0(.din(w_dff_B_Y1IV97me7_0),.dout(w_dff_B_yL46Ax4v3_0),.clk(gclk));
	jdff dff_B_fh5LHN6Z9_0(.din(w_dff_B_yL46Ax4v3_0),.dout(w_dff_B_fh5LHN6Z9_0),.clk(gclk));
	jdff dff_B_yEGekuBd7_0(.din(w_dff_B_fh5LHN6Z9_0),.dout(w_dff_B_yEGekuBd7_0),.clk(gclk));
	jdff dff_B_WT21Q8Wg1_0(.din(w_dff_B_yEGekuBd7_0),.dout(w_dff_B_WT21Q8Wg1_0),.clk(gclk));
	jdff dff_B_PrVErDRB6_0(.din(w_dff_B_WT21Q8Wg1_0),.dout(w_dff_B_PrVErDRB6_0),.clk(gclk));
	jdff dff_B_pOXsZQ7t5_1(.din(n1053),.dout(w_dff_B_pOXsZQ7t5_1),.clk(gclk));
	jdff dff_B_TzjUy8CR7_1(.din(w_dff_B_pOXsZQ7t5_1),.dout(w_dff_B_TzjUy8CR7_1),.clk(gclk));
	jdff dff_B_BkBJegN79_1(.din(w_dff_B_TzjUy8CR7_1),.dout(w_dff_B_BkBJegN79_1),.clk(gclk));
	jdff dff_A_foNLMS0P2_0(.dout(w_n800_3[0]),.din(w_dff_A_foNLMS0P2_0),.clk(gclk));
	jdff dff_A_Hu32o2cR8_2(.dout(w_n800_3[2]),.din(w_dff_A_Hu32o2cR8_2),.clk(gclk));
	jdff dff_A_ptkvh7EA1_2(.dout(w_dff_A_Hu32o2cR8_2),.din(w_dff_A_ptkvh7EA1_2),.clk(gclk));
	jdff dff_B_3CTSQPKb8_1(.din(n1066),.dout(w_dff_B_3CTSQPKb8_1),.clk(gclk));
	jdff dff_B_fijrpWob9_1(.din(w_dff_B_3CTSQPKb8_1),.dout(w_dff_B_fijrpWob9_1),.clk(gclk));
	jdff dff_B_cH8S5oks3_1(.din(w_dff_B_fijrpWob9_1),.dout(w_dff_B_cH8S5oks3_1),.clk(gclk));
	jdff dff_B_E5l4s9jY8_1(.din(w_dff_B_cH8S5oks3_1),.dout(w_dff_B_E5l4s9jY8_1),.clk(gclk));
	jdff dff_B_zycsE9ZW7_1(.din(w_dff_B_E5l4s9jY8_1),.dout(w_dff_B_zycsE9ZW7_1),.clk(gclk));
	jdff dff_B_7ZP9AhMz0_1(.din(w_dff_B_zycsE9ZW7_1),.dout(w_dff_B_7ZP9AhMz0_1),.clk(gclk));
	jdff dff_B_a5S6kHUC3_1(.din(w_dff_B_7ZP9AhMz0_1),.dout(w_dff_B_a5S6kHUC3_1),.clk(gclk));
	jdff dff_B_0YZn9x8B0_1(.din(w_dff_B_a5S6kHUC3_1),.dout(w_dff_B_0YZn9x8B0_1),.clk(gclk));
	jdff dff_B_SbA090H36_1(.din(w_dff_B_0YZn9x8B0_1),.dout(w_dff_B_SbA090H36_1),.clk(gclk));
	jdff dff_B_DRl243DJ4_1(.din(w_dff_B_SbA090H36_1),.dout(w_dff_B_DRl243DJ4_1),.clk(gclk));
	jdff dff_B_SsELJ9Fa7_1(.din(w_dff_B_DRl243DJ4_1),.dout(w_dff_B_SsELJ9Fa7_1),.clk(gclk));
	jdff dff_B_JRRzcMFs5_1(.din(w_dff_B_SsELJ9Fa7_1),.dout(w_dff_B_JRRzcMFs5_1),.clk(gclk));
	jdff dff_B_2xTmNc0b9_1(.din(w_dff_B_JRRzcMFs5_1),.dout(w_dff_B_2xTmNc0b9_1),.clk(gclk));
	jdff dff_B_EitWhjPr9_1(.din(w_dff_B_2xTmNc0b9_1),.dout(w_dff_B_EitWhjPr9_1),.clk(gclk));
	jdff dff_B_sw0kQIIT5_1(.din(w_dff_B_EitWhjPr9_1),.dout(w_dff_B_sw0kQIIT5_1),.clk(gclk));
	jdff dff_A_ebht2U5w7_0(.dout(w_n854_4[0]),.din(w_dff_A_ebht2U5w7_0),.clk(gclk));
	jdff dff_A_hV5J1of21_0(.dout(w_dff_A_ebht2U5w7_0),.din(w_dff_A_hV5J1of21_0),.clk(gclk));
	jdff dff_A_sy4FFc0i5_0(.dout(w_dff_A_hV5J1of21_0),.din(w_dff_A_sy4FFc0i5_0),.clk(gclk));
	jdff dff_A_EB8dtqpN0_0(.dout(w_dff_A_sy4FFc0i5_0),.din(w_dff_A_EB8dtqpN0_0),.clk(gclk));
	jdff dff_A_4nLjo1g16_0(.dout(w_dff_A_EB8dtqpN0_0),.din(w_dff_A_4nLjo1g16_0),.clk(gclk));
	jdff dff_A_p4UPIfMP6_0(.dout(w_dff_A_4nLjo1g16_0),.din(w_dff_A_p4UPIfMP6_0),.clk(gclk));
	jdff dff_A_olaywdnc3_0(.dout(w_dff_A_p4UPIfMP6_0),.din(w_dff_A_olaywdnc3_0),.clk(gclk));
	jdff dff_A_p2PiHSc06_0(.dout(w_dff_A_olaywdnc3_0),.din(w_dff_A_p2PiHSc06_0),.clk(gclk));
	jdff dff_B_KLHKgBge4_1(.din(n1063),.dout(w_dff_B_KLHKgBge4_1),.clk(gclk));
	jdff dff_B_fm2x8dKD1_1(.din(w_dff_B_KLHKgBge4_1),.dout(w_dff_B_fm2x8dKD1_1),.clk(gclk));
	jdff dff_B_h9kxZlyU6_2(.din(G37),.dout(w_dff_B_h9kxZlyU6_2),.clk(gclk));
	jdff dff_B_fKlRZZMc0_1(.din(n1075),.dout(w_dff_B_fKlRZZMc0_1),.clk(gclk));
	jdff dff_B_8ooZeVHK3_1(.din(w_dff_B_fKlRZZMc0_1),.dout(w_dff_B_8ooZeVHK3_1),.clk(gclk));
	jdff dff_B_X8ZmFST18_1(.din(w_dff_B_8ooZeVHK3_1),.dout(w_dff_B_X8ZmFST18_1),.clk(gclk));
	jdff dff_B_krsKa70A5_1(.din(w_dff_B_X8ZmFST18_1),.dout(w_dff_B_krsKa70A5_1),.clk(gclk));
	jdff dff_B_67anivFM8_1(.din(w_dff_B_krsKa70A5_1),.dout(w_dff_B_67anivFM8_1),.clk(gclk));
	jdff dff_B_pcoQU6oO2_1(.din(w_dff_B_67anivFM8_1),.dout(w_dff_B_pcoQU6oO2_1),.clk(gclk));
	jdff dff_B_qlaTCUvJ4_1(.din(w_dff_B_pcoQU6oO2_1),.dout(w_dff_B_qlaTCUvJ4_1),.clk(gclk));
	jdff dff_B_iAz9VOY70_1(.din(w_dff_B_qlaTCUvJ4_1),.dout(w_dff_B_iAz9VOY70_1),.clk(gclk));
	jdff dff_B_4QN1Pk018_1(.din(w_dff_B_iAz9VOY70_1),.dout(w_dff_B_4QN1Pk018_1),.clk(gclk));
	jdff dff_B_eZD9rZFq6_1(.din(w_dff_B_4QN1Pk018_1),.dout(w_dff_B_eZD9rZFq6_1),.clk(gclk));
	jdff dff_B_WIKI6WIU3_1(.din(w_dff_B_eZD9rZFq6_1),.dout(w_dff_B_WIKI6WIU3_1),.clk(gclk));
	jdff dff_B_gSEg92IP8_1(.din(w_dff_B_WIKI6WIU3_1),.dout(w_dff_B_gSEg92IP8_1),.clk(gclk));
	jdff dff_B_1Ho6YZSd5_1(.din(w_dff_B_gSEg92IP8_1),.dout(w_dff_B_1Ho6YZSd5_1),.clk(gclk));
	jdff dff_B_R3xuKQ1A8_1(.din(w_dff_B_1Ho6YZSd5_1),.dout(w_dff_B_R3xuKQ1A8_1),.clk(gclk));
	jdff dff_B_3RUDA86W1_0(.din(n1077),.dout(w_dff_B_3RUDA86W1_0),.clk(gclk));
	jdff dff_B_FiZVK3de1_1(.din(n1072),.dout(w_dff_B_FiZVK3de1_1),.clk(gclk));
	jdff dff_B_dSaYggRw8_1(.din(w_dff_B_FiZVK3de1_1),.dout(w_dff_B_dSaYggRw8_1),.clk(gclk));
	jdff dff_A_CABZ38Nm4_1(.dout(w_n852_8[1]),.din(w_dff_A_CABZ38Nm4_1),.clk(gclk));
	jdff dff_A_Mhpg5Sw66_1(.dout(w_dff_A_CABZ38Nm4_1),.din(w_dff_A_Mhpg5Sw66_1),.clk(gclk));
	jdff dff_A_2f3ygkh53_1(.dout(w_dff_A_Mhpg5Sw66_1),.din(w_dff_A_2f3ygkh53_1),.clk(gclk));
	jdff dff_A_1pNpKMnn3_1(.dout(w_dff_A_2f3ygkh53_1),.din(w_dff_A_1pNpKMnn3_1),.clk(gclk));
	jdff dff_A_UFtGMjOv9_1(.dout(w_dff_A_1pNpKMnn3_1),.din(w_dff_A_UFtGMjOv9_1),.clk(gclk));
	jdff dff_A_G7Upt35M5_1(.dout(w_dff_A_UFtGMjOv9_1),.din(w_dff_A_G7Upt35M5_1),.clk(gclk));
	jdff dff_A_wHomhmqu2_1(.dout(w_dff_A_G7Upt35M5_1),.din(w_dff_A_wHomhmqu2_1),.clk(gclk));
	jdff dff_A_2evvlSFa6_1(.dout(w_dff_A_wHomhmqu2_1),.din(w_dff_A_2evvlSFa6_1),.clk(gclk));
	jdff dff_A_THPnx7fu3_1(.dout(w_dff_A_2evvlSFa6_1),.din(w_dff_A_THPnx7fu3_1),.clk(gclk));
	jdff dff_A_XpyDvBDb2_1(.dout(w_dff_A_THPnx7fu3_1),.din(w_dff_A_XpyDvBDb2_1),.clk(gclk));
	jdff dff_A_svcPAzKj3_1(.dout(w_dff_A_XpyDvBDb2_1),.din(w_dff_A_svcPAzKj3_1),.clk(gclk));
	jdff dff_A_otY84Bj83_1(.dout(w_dff_A_svcPAzKj3_1),.din(w_dff_A_otY84Bj83_1),.clk(gclk));
	jdff dff_A_1xzMNccD6_1(.dout(w_dff_A_otY84Bj83_1),.din(w_dff_A_1xzMNccD6_1),.clk(gclk));
	jdff dff_A_MIEN68w72_1(.dout(w_dff_A_1xzMNccD6_1),.din(w_dff_A_MIEN68w72_1),.clk(gclk));
	jdff dff_A_p2KaDZoD7_1(.dout(w_dff_A_MIEN68w72_1),.din(w_dff_A_p2KaDZoD7_1),.clk(gclk));
	jdff dff_B_MZAmZeka7_2(.din(G20),.dout(w_dff_B_MZAmZeka7_2),.clk(gclk));
	jdff dff_A_4gwFou728_1(.dout(w_G4089_8[1]),.din(w_dff_A_4gwFou728_1),.clk(gclk));
	jdff dff_A_nDKLfZ6A8_1(.dout(w_dff_A_4gwFou728_1),.din(w_dff_A_nDKLfZ6A8_1),.clk(gclk));
	jdff dff_A_LVXdMjz14_1(.dout(w_dff_A_nDKLfZ6A8_1),.din(w_dff_A_LVXdMjz14_1),.clk(gclk));
	jdff dff_A_UMAllwSa6_1(.dout(w_dff_A_LVXdMjz14_1),.din(w_dff_A_UMAllwSa6_1),.clk(gclk));
	jdff dff_A_ZbHJusbg5_1(.dout(w_dff_A_UMAllwSa6_1),.din(w_dff_A_ZbHJusbg5_1),.clk(gclk));
	jdff dff_A_eeUq2Ocq7_1(.dout(w_dff_A_ZbHJusbg5_1),.din(w_dff_A_eeUq2Ocq7_1),.clk(gclk));
	jdff dff_A_2cVaDhVt5_1(.dout(w_dff_A_eeUq2Ocq7_1),.din(w_dff_A_2cVaDhVt5_1),.clk(gclk));
	jdff dff_A_n6PN850D5_1(.dout(w_dff_A_2cVaDhVt5_1),.din(w_dff_A_n6PN850D5_1),.clk(gclk));
	jdff dff_A_OSHVIPAF3_1(.dout(w_dff_A_n6PN850D5_1),.din(w_dff_A_OSHVIPAF3_1),.clk(gclk));
	jdff dff_A_MCF6eygg6_1(.dout(w_dff_A_OSHVIPAF3_1),.din(w_dff_A_MCF6eygg6_1),.clk(gclk));
	jdff dff_A_ATIub3M57_1(.dout(w_dff_A_MCF6eygg6_1),.din(w_dff_A_ATIub3M57_1),.clk(gclk));
	jdff dff_A_cZyCyK2P3_1(.dout(w_dff_A_ATIub3M57_1),.din(w_dff_A_cZyCyK2P3_1),.clk(gclk));
	jdff dff_A_8MendlBx5_1(.dout(w_dff_A_cZyCyK2P3_1),.din(w_dff_A_8MendlBx5_1),.clk(gclk));
	jdff dff_A_4GTmbS0q8_1(.dout(w_dff_A_8MendlBx5_1),.din(w_dff_A_4GTmbS0q8_1),.clk(gclk));
	jdff dff_A_R5t2f0y17_1(.dout(w_dff_A_4GTmbS0q8_1),.din(w_dff_A_R5t2f0y17_1),.clk(gclk));
	jdff dff_A_DGMxBQG38_1(.dout(w_dff_A_R5t2f0y17_1),.din(w_dff_A_DGMxBQG38_1),.clk(gclk));
	jdff dff_B_U62sgSUC8_1(.din(n1084),.dout(w_dff_B_U62sgSUC8_1),.clk(gclk));
	jdff dff_B_xB9NwQL76_1(.din(w_dff_B_U62sgSUC8_1),.dout(w_dff_B_xB9NwQL76_1),.clk(gclk));
	jdff dff_B_y19k6eIt3_1(.din(w_dff_B_xB9NwQL76_1),.dout(w_dff_B_y19k6eIt3_1),.clk(gclk));
	jdff dff_B_s05LFa7k9_1(.din(w_dff_B_y19k6eIt3_1),.dout(w_dff_B_s05LFa7k9_1),.clk(gclk));
	jdff dff_B_i3CRBM249_1(.din(w_dff_B_s05LFa7k9_1),.dout(w_dff_B_i3CRBM249_1),.clk(gclk));
	jdff dff_B_S6GmqtZn9_1(.din(w_dff_B_i3CRBM249_1),.dout(w_dff_B_S6GmqtZn9_1),.clk(gclk));
	jdff dff_B_ul5oidY57_1(.din(w_dff_B_S6GmqtZn9_1),.dout(w_dff_B_ul5oidY57_1),.clk(gclk));
	jdff dff_B_fdimDfiK2_1(.din(w_dff_B_ul5oidY57_1),.dout(w_dff_B_fdimDfiK2_1),.clk(gclk));
	jdff dff_B_3GWiesPE3_1(.din(w_dff_B_fdimDfiK2_1),.dout(w_dff_B_3GWiesPE3_1),.clk(gclk));
	jdff dff_B_AUFu4Drc0_1(.din(w_dff_B_3GWiesPE3_1),.dout(w_dff_B_AUFu4Drc0_1),.clk(gclk));
	jdff dff_B_KDCB6Twn2_1(.din(w_dff_B_AUFu4Drc0_1),.dout(w_dff_B_KDCB6Twn2_1),.clk(gclk));
	jdff dff_B_QtbKjWVe1_1(.din(w_dff_B_KDCB6Twn2_1),.dout(w_dff_B_QtbKjWVe1_1),.clk(gclk));
	jdff dff_B_2Krg9KE16_1(.din(n1081),.dout(w_dff_B_2Krg9KE16_1),.clk(gclk));
	jdff dff_B_wsR42LE81_1(.din(w_dff_B_2Krg9KE16_1),.dout(w_dff_B_wsR42LE81_1),.clk(gclk));
	jdff dff_A_AdgkasZo8_0(.dout(w_n852_7[0]),.din(w_dff_A_AdgkasZo8_0),.clk(gclk));
	jdff dff_A_3wMHiP440_0(.dout(w_dff_A_AdgkasZo8_0),.din(w_dff_A_3wMHiP440_0),.clk(gclk));
	jdff dff_A_2CVtRpox0_0(.dout(w_dff_A_3wMHiP440_0),.din(w_dff_A_2CVtRpox0_0),.clk(gclk));
	jdff dff_A_JpFHzrtN9_0(.dout(w_dff_A_2CVtRpox0_0),.din(w_dff_A_JpFHzrtN9_0),.clk(gclk));
	jdff dff_A_4lukrovC8_0(.dout(w_dff_A_JpFHzrtN9_0),.din(w_dff_A_4lukrovC8_0),.clk(gclk));
	jdff dff_A_7HUDM1Yw4_0(.dout(w_dff_A_4lukrovC8_0),.din(w_dff_A_7HUDM1Yw4_0),.clk(gclk));
	jdff dff_A_Azb8ug1R9_0(.dout(w_dff_A_7HUDM1Yw4_0),.din(w_dff_A_Azb8ug1R9_0),.clk(gclk));
	jdff dff_A_Bb8YF7Ma6_0(.dout(w_dff_A_Azb8ug1R9_0),.din(w_dff_A_Bb8YF7Ma6_0),.clk(gclk));
	jdff dff_A_cQkQ1UbB1_0(.dout(w_dff_A_Bb8YF7Ma6_0),.din(w_dff_A_cQkQ1UbB1_0),.clk(gclk));
	jdff dff_A_pcWhhPNn3_0(.dout(w_dff_A_cQkQ1UbB1_0),.din(w_dff_A_pcWhhPNn3_0),.clk(gclk));
	jdff dff_A_fVceHLmP6_0(.dout(w_dff_A_pcWhhPNn3_0),.din(w_dff_A_fVceHLmP6_0),.clk(gclk));
	jdff dff_A_z4pdcwoX3_0(.dout(w_dff_A_fVceHLmP6_0),.din(w_dff_A_z4pdcwoX3_0),.clk(gclk));
	jdff dff_A_33GAKJi55_2(.dout(w_n852_7[2]),.din(w_dff_A_33GAKJi55_2),.clk(gclk));
	jdff dff_A_EgB1K0cH3_2(.dout(w_dff_A_33GAKJi55_2),.din(w_dff_A_EgB1K0cH3_2),.clk(gclk));
	jdff dff_A_RUC4aArw9_2(.dout(w_dff_A_EgB1K0cH3_2),.din(w_dff_A_RUC4aArw9_2),.clk(gclk));
	jdff dff_A_DunTaVRw4_2(.dout(w_dff_A_RUC4aArw9_2),.din(w_dff_A_DunTaVRw4_2),.clk(gclk));
	jdff dff_A_2ZDS1ZtK8_2(.dout(w_dff_A_DunTaVRw4_2),.din(w_dff_A_2ZDS1ZtK8_2),.clk(gclk));
	jdff dff_A_o4Hb3cco8_2(.dout(w_dff_A_2ZDS1ZtK8_2),.din(w_dff_A_o4Hb3cco8_2),.clk(gclk));
	jdff dff_A_7SqNkHp28_2(.dout(w_dff_A_o4Hb3cco8_2),.din(w_dff_A_7SqNkHp28_2),.clk(gclk));
	jdff dff_A_B21LMjTn3_2(.dout(w_dff_A_7SqNkHp28_2),.din(w_dff_A_B21LMjTn3_2),.clk(gclk));
	jdff dff_A_nB8D89q28_2(.dout(w_dff_A_B21LMjTn3_2),.din(w_dff_A_nB8D89q28_2),.clk(gclk));
	jdff dff_A_HIX9uVYh9_2(.dout(w_dff_A_nB8D89q28_2),.din(w_dff_A_HIX9uVYh9_2),.clk(gclk));
	jdff dff_A_RyWzwAUx5_2(.dout(w_dff_A_HIX9uVYh9_2),.din(w_dff_A_RyWzwAUx5_2),.clk(gclk));
	jdff dff_A_98xNmKra5_2(.dout(w_dff_A_RyWzwAUx5_2),.din(w_dff_A_98xNmKra5_2),.clk(gclk));
	jdff dff_A_js8pimOP0_2(.dout(w_dff_A_98xNmKra5_2),.din(w_dff_A_js8pimOP0_2),.clk(gclk));
	jdff dff_B_RPIWd08X5_2(.din(G17),.dout(w_dff_B_RPIWd08X5_2),.clk(gclk));
	jdff dff_A_H2jeIYjO1_0(.dout(w_G4089_7[0]),.din(w_dff_A_H2jeIYjO1_0),.clk(gclk));
	jdff dff_A_nrzLWmSR1_0(.dout(w_dff_A_H2jeIYjO1_0),.din(w_dff_A_nrzLWmSR1_0),.clk(gclk));
	jdff dff_A_44DkNbkz7_0(.dout(w_dff_A_nrzLWmSR1_0),.din(w_dff_A_44DkNbkz7_0),.clk(gclk));
	jdff dff_A_m6WbrJ8L0_0(.dout(w_dff_A_44DkNbkz7_0),.din(w_dff_A_m6WbrJ8L0_0),.clk(gclk));
	jdff dff_A_lapcYyYX9_0(.dout(w_dff_A_m6WbrJ8L0_0),.din(w_dff_A_lapcYyYX9_0),.clk(gclk));
	jdff dff_A_O62LtL2A0_0(.dout(w_dff_A_lapcYyYX9_0),.din(w_dff_A_O62LtL2A0_0),.clk(gclk));
	jdff dff_A_5Gdr1D451_0(.dout(w_dff_A_O62LtL2A0_0),.din(w_dff_A_5Gdr1D451_0),.clk(gclk));
	jdff dff_A_XuHovybZ8_0(.dout(w_dff_A_5Gdr1D451_0),.din(w_dff_A_XuHovybZ8_0),.clk(gclk));
	jdff dff_A_Wc0Fc5UN9_0(.dout(w_dff_A_XuHovybZ8_0),.din(w_dff_A_Wc0Fc5UN9_0),.clk(gclk));
	jdff dff_A_27Pe6pAY1_0(.dout(w_dff_A_Wc0Fc5UN9_0),.din(w_dff_A_27Pe6pAY1_0),.clk(gclk));
	jdff dff_A_pVhTbSdy7_0(.dout(w_dff_A_27Pe6pAY1_0),.din(w_dff_A_pVhTbSdy7_0),.clk(gclk));
	jdff dff_A_BUisNmyH8_0(.dout(w_dff_A_pVhTbSdy7_0),.din(w_dff_A_BUisNmyH8_0),.clk(gclk));
	jdff dff_A_EGw3OCqi1_0(.dout(w_dff_A_BUisNmyH8_0),.din(w_dff_A_EGw3OCqi1_0),.clk(gclk));
	jdff dff_A_oK2ZZWd80_2(.dout(w_G4089_7[2]),.din(w_dff_A_oK2ZZWd80_2),.clk(gclk));
	jdff dff_A_cbpnOs2t2_2(.dout(w_dff_A_oK2ZZWd80_2),.din(w_dff_A_cbpnOs2t2_2),.clk(gclk));
	jdff dff_A_1dQ0nBsJ4_2(.dout(w_dff_A_cbpnOs2t2_2),.din(w_dff_A_1dQ0nBsJ4_2),.clk(gclk));
	jdff dff_A_wnUlBMJS2_2(.dout(w_dff_A_1dQ0nBsJ4_2),.din(w_dff_A_wnUlBMJS2_2),.clk(gclk));
	jdff dff_A_tAIIr8Mb2_2(.dout(w_dff_A_wnUlBMJS2_2),.din(w_dff_A_tAIIr8Mb2_2),.clk(gclk));
	jdff dff_A_U4VeFLT89_2(.dout(w_dff_A_tAIIr8Mb2_2),.din(w_dff_A_U4VeFLT89_2),.clk(gclk));
	jdff dff_A_0YTHVqHw1_2(.dout(w_dff_A_U4VeFLT89_2),.din(w_dff_A_0YTHVqHw1_2),.clk(gclk));
	jdff dff_A_Uv1ru2fl1_2(.dout(w_dff_A_0YTHVqHw1_2),.din(w_dff_A_Uv1ru2fl1_2),.clk(gclk));
	jdff dff_A_UYzecIFh4_2(.dout(w_dff_A_Uv1ru2fl1_2),.din(w_dff_A_UYzecIFh4_2),.clk(gclk));
	jdff dff_A_QgoiUmMT1_2(.dout(w_dff_A_UYzecIFh4_2),.din(w_dff_A_QgoiUmMT1_2),.clk(gclk));
	jdff dff_A_TntnKZWC6_2(.dout(w_dff_A_QgoiUmMT1_2),.din(w_dff_A_TntnKZWC6_2),.clk(gclk));
	jdff dff_A_P7p4HuS22_2(.dout(w_dff_A_TntnKZWC6_2),.din(w_dff_A_P7p4HuS22_2),.clk(gclk));
	jdff dff_A_6eMntC6i9_2(.dout(w_dff_A_P7p4HuS22_2),.din(w_dff_A_6eMntC6i9_2),.clk(gclk));
	jdff dff_A_i9DnFPfo7_2(.dout(w_dff_A_6eMntC6i9_2),.din(w_dff_A_i9DnFPfo7_2),.clk(gclk));
	jdff dff_A_d2WmELSA3_2(.dout(w_dff_A_i9DnFPfo7_2),.din(w_dff_A_d2WmELSA3_2),.clk(gclk));
	jdff dff_B_dwgKOCQT5_0(.din(n1097),.dout(w_dff_B_dwgKOCQT5_0),.clk(gclk));
	jdff dff_B_MJXpMlSz8_0(.din(w_dff_B_dwgKOCQT5_0),.dout(w_dff_B_MJXpMlSz8_0),.clk(gclk));
	jdff dff_B_lVtnwA7P9_0(.din(w_dff_B_MJXpMlSz8_0),.dout(w_dff_B_lVtnwA7P9_0),.clk(gclk));
	jdff dff_B_q54FTbbG2_0(.din(w_dff_B_lVtnwA7P9_0),.dout(w_dff_B_q54FTbbG2_0),.clk(gclk));
	jdff dff_B_LEZjdAOF2_0(.din(w_dff_B_q54FTbbG2_0),.dout(w_dff_B_LEZjdAOF2_0),.clk(gclk));
	jdff dff_B_K5gxWMxw9_0(.din(w_dff_B_LEZjdAOF2_0),.dout(w_dff_B_K5gxWMxw9_0),.clk(gclk));
	jdff dff_B_jhGhSjXn1_0(.din(w_dff_B_K5gxWMxw9_0),.dout(w_dff_B_jhGhSjXn1_0),.clk(gclk));
	jdff dff_B_XXn0nBBT4_0(.din(w_dff_B_jhGhSjXn1_0),.dout(w_dff_B_XXn0nBBT4_0),.clk(gclk));
	jdff dff_B_8XvexMbO0_0(.din(w_dff_B_XXn0nBBT4_0),.dout(w_dff_B_8XvexMbO0_0),.clk(gclk));
	jdff dff_B_k5ROGEeQ9_0(.din(w_dff_B_8XvexMbO0_0),.dout(w_dff_B_k5ROGEeQ9_0),.clk(gclk));
	jdff dff_B_dPS8gKbJ3_0(.din(w_dff_B_k5ROGEeQ9_0),.dout(w_dff_B_dPS8gKbJ3_0),.clk(gclk));
	jdff dff_B_Mqwo4kXx0_0(.din(w_dff_B_dPS8gKbJ3_0),.dout(w_dff_B_Mqwo4kXx0_0),.clk(gclk));
	jdff dff_B_tgwF8Qzt1_0(.din(w_dff_B_Mqwo4kXx0_0),.dout(w_dff_B_tgwF8Qzt1_0),.clk(gclk));
	jdff dff_B_fUQ7IRTy5_0(.din(w_dff_B_tgwF8Qzt1_0),.dout(w_dff_B_fUQ7IRTy5_0),.clk(gclk));
	jdff dff_A_YxLnYYPV2_1(.dout(w_G4090_3[1]),.din(w_dff_A_YxLnYYPV2_1),.clk(gclk));
	jdff dff_A_wZ5mTor86_2(.dout(w_G4090_3[2]),.din(w_dff_A_wZ5mTor86_2),.clk(gclk));
	jdff dff_B_FIoheWbs5_2(.din(G70),.dout(w_dff_B_FIoheWbs5_2),.clk(gclk));
	jdff dff_B_IGq84fdi5_1(.din(n1090),.dout(w_dff_B_IGq84fdi5_1),.clk(gclk));
	jdff dff_B_Y32ShMuw6_1(.din(w_dff_B_IGq84fdi5_1),.dout(w_dff_B_Y32ShMuw6_1),.clk(gclk));
	jdff dff_B_hPqcY2iD9_1(.din(w_dff_B_Y32ShMuw6_1),.dout(w_dff_B_hPqcY2iD9_1),.clk(gclk));
	jdff dff_A_3W4kvWNZ3_2(.dout(w_n854_3[2]),.din(w_dff_A_3W4kvWNZ3_2),.clk(gclk));
	jdff dff_A_nMHJbxjT1_2(.dout(w_dff_A_3W4kvWNZ3_2),.din(w_dff_A_nMHJbxjT1_2),.clk(gclk));
	jdff dff_B_ZVmm8MNS6_0(.din(n1105),.dout(w_dff_B_ZVmm8MNS6_0),.clk(gclk));
	jdff dff_B_0A3Ro9nz0_0(.din(w_dff_B_ZVmm8MNS6_0),.dout(w_dff_B_0A3Ro9nz0_0),.clk(gclk));
	jdff dff_B_ep9uS0Mf1_0(.din(w_dff_B_0A3Ro9nz0_0),.dout(w_dff_B_ep9uS0Mf1_0),.clk(gclk));
	jdff dff_B_3aDHVfrs0_0(.din(w_dff_B_ep9uS0Mf1_0),.dout(w_dff_B_3aDHVfrs0_0),.clk(gclk));
	jdff dff_B_ujgqR1BA0_0(.din(w_dff_B_3aDHVfrs0_0),.dout(w_dff_B_ujgqR1BA0_0),.clk(gclk));
	jdff dff_B_Lpe4bac67_0(.din(w_dff_B_ujgqR1BA0_0),.dout(w_dff_B_Lpe4bac67_0),.clk(gclk));
	jdff dff_B_qqefWXnl8_0(.din(w_dff_B_Lpe4bac67_0),.dout(w_dff_B_qqefWXnl8_0),.clk(gclk));
	jdff dff_B_2YvTkKCA9_0(.din(w_dff_B_qqefWXnl8_0),.dout(w_dff_B_2YvTkKCA9_0),.clk(gclk));
	jdff dff_B_kWAgN8za5_0(.din(w_dff_B_2YvTkKCA9_0),.dout(w_dff_B_kWAgN8za5_0),.clk(gclk));
	jdff dff_B_h2W2eMv27_0(.din(w_dff_B_kWAgN8za5_0),.dout(w_dff_B_h2W2eMv27_0),.clk(gclk));
	jdff dff_B_eYQWpjpO9_0(.din(w_dff_B_h2W2eMv27_0),.dout(w_dff_B_eYQWpjpO9_0),.clk(gclk));
	jdff dff_B_u2gv6qbn2_0(.din(w_dff_B_eYQWpjpO9_0),.dout(w_dff_B_u2gv6qbn2_0),.clk(gclk));
	jdff dff_B_65GFBJ5i0_0(.din(w_dff_B_u2gv6qbn2_0),.dout(w_dff_B_65GFBJ5i0_0),.clk(gclk));
	jdff dff_B_1S2oHxRv6_0(.din(w_dff_B_65GFBJ5i0_0),.dout(w_dff_B_1S2oHxRv6_0),.clk(gclk));
	jdff dff_B_n4Z3kC0B8_0(.din(w_dff_B_1S2oHxRv6_0),.dout(w_dff_B_n4Z3kC0B8_0),.clk(gclk));
	jdff dff_B_69LkdRe29_0(.din(n1104),.dout(w_dff_B_69LkdRe29_0),.clk(gclk));
	jdff dff_B_BFLz6QQE7_1(.din(n1099),.dout(w_dff_B_BFLz6QQE7_1),.clk(gclk));
	jdff dff_B_WEtm194H6_0(.din(n1114),.dout(w_dff_B_WEtm194H6_0),.clk(gclk));
	jdff dff_B_7IBwxlQT2_0(.din(w_dff_B_WEtm194H6_0),.dout(w_dff_B_7IBwxlQT2_0),.clk(gclk));
	jdff dff_B_HnBuq4GM7_0(.din(w_dff_B_7IBwxlQT2_0),.dout(w_dff_B_HnBuq4GM7_0),.clk(gclk));
	jdff dff_B_j0gK1YOY6_0(.din(w_dff_B_HnBuq4GM7_0),.dout(w_dff_B_j0gK1YOY6_0),.clk(gclk));
	jdff dff_B_817Q2Pqi5_0(.din(w_dff_B_j0gK1YOY6_0),.dout(w_dff_B_817Q2Pqi5_0),.clk(gclk));
	jdff dff_B_J9CF1wra9_0(.din(w_dff_B_817Q2Pqi5_0),.dout(w_dff_B_J9CF1wra9_0),.clk(gclk));
	jdff dff_B_rC1cw62D8_0(.din(w_dff_B_J9CF1wra9_0),.dout(w_dff_B_rC1cw62D8_0),.clk(gclk));
	jdff dff_B_xWmwhYEu5_0(.din(w_dff_B_rC1cw62D8_0),.dout(w_dff_B_xWmwhYEu5_0),.clk(gclk));
	jdff dff_B_NAUXOCim6_0(.din(w_dff_B_xWmwhYEu5_0),.dout(w_dff_B_NAUXOCim6_0),.clk(gclk));
	jdff dff_B_NeoQELkz9_0(.din(w_dff_B_NAUXOCim6_0),.dout(w_dff_B_NeoQELkz9_0),.clk(gclk));
	jdff dff_B_nsN7kUO77_0(.din(w_dff_B_NeoQELkz9_0),.dout(w_dff_B_nsN7kUO77_0),.clk(gclk));
	jdff dff_B_Fo0Afh4i9_0(.din(w_dff_B_nsN7kUO77_0),.dout(w_dff_B_Fo0Afh4i9_0),.clk(gclk));
	jdff dff_B_44vAecWO2_0(.din(n1113),.dout(w_dff_B_44vAecWO2_0),.clk(gclk));
	jdff dff_B_jYDj2gId5_0(.din(n1110),.dout(w_dff_B_jYDj2gId5_0),.clk(gclk));
	jdff dff_A_sc3jI8Q69_0(.dout(w_n999_3[0]),.din(w_dff_A_sc3jI8Q69_0),.clk(gclk));
	jdff dff_A_ojvfwOxf9_0(.dout(w_dff_A_sc3jI8Q69_0),.din(w_dff_A_ojvfwOxf9_0),.clk(gclk));
	jdff dff_A_RUcvG7n60_0(.dout(w_dff_A_ojvfwOxf9_0),.din(w_dff_A_RUcvG7n60_0),.clk(gclk));
	jdff dff_A_ax7OvO1A0_1(.dout(w_n999_3[1]),.din(w_dff_A_ax7OvO1A0_1),.clk(gclk));
	jdff dff_A_1tEDy0cf0_1(.dout(w_dff_A_ax7OvO1A0_1),.din(w_dff_A_1tEDy0cf0_1),.clk(gclk));
	jdff dff_A_By1RKrdX8_1(.dout(w_dff_A_1tEDy0cf0_1),.din(w_dff_A_By1RKrdX8_1),.clk(gclk));
	jdff dff_A_DC7nCXXN2_1(.dout(w_dff_A_By1RKrdX8_1),.din(w_dff_A_DC7nCXXN2_1),.clk(gclk));
	jdff dff_A_sjV8SmEY9_1(.dout(w_dff_A_DC7nCXXN2_1),.din(w_dff_A_sjV8SmEY9_1),.clk(gclk));
	jdff dff_A_eihDuhsQ7_1(.dout(w_dff_A_sjV8SmEY9_1),.din(w_dff_A_eihDuhsQ7_1),.clk(gclk));
	jdff dff_A_ex2SzdNi7_1(.dout(w_dff_A_eihDuhsQ7_1),.din(w_dff_A_ex2SzdNi7_1),.clk(gclk));
	jdff dff_A_xXCSNQrE9_0(.dout(w_G1689_4[0]),.din(w_dff_A_xXCSNQrE9_0),.clk(gclk));
	jdff dff_A_NbS7Alik6_0(.dout(w_dff_A_xXCSNQrE9_0),.din(w_dff_A_NbS7Alik6_0),.clk(gclk));
	jdff dff_A_FPGa4Tmv5_0(.dout(w_dff_A_NbS7Alik6_0),.din(w_dff_A_FPGa4Tmv5_0),.clk(gclk));
	jdff dff_A_4mEEVqk35_0(.dout(w_dff_A_FPGa4Tmv5_0),.din(w_dff_A_4mEEVqk35_0),.clk(gclk));
	jdff dff_A_BNuCiqWE6_0(.dout(w_dff_A_4mEEVqk35_0),.din(w_dff_A_BNuCiqWE6_0),.clk(gclk));
	jdff dff_A_gyXkKqaX3_1(.dout(w_G1689_4[1]),.din(w_dff_A_gyXkKqaX3_1),.clk(gclk));
	jdff dff_A_0fZTBHr02_1(.dout(w_dff_A_gyXkKqaX3_1),.din(w_dff_A_0fZTBHr02_1),.clk(gclk));
	jdff dff_A_If7SqYPf4_1(.dout(w_dff_A_0fZTBHr02_1),.din(w_dff_A_If7SqYPf4_1),.clk(gclk));
	jdff dff_A_9DpGzOIF8_1(.dout(w_dff_A_If7SqYPf4_1),.din(w_dff_A_9DpGzOIF8_1),.clk(gclk));
	jdff dff_A_mKOuAFjK0_1(.dout(w_dff_A_9DpGzOIF8_1),.din(w_dff_A_mKOuAFjK0_1),.clk(gclk));
	jdff dff_A_L7SHkB7f7_1(.dout(w_dff_A_mKOuAFjK0_1),.din(w_dff_A_L7SHkB7f7_1),.clk(gclk));
	jdff dff_A_NmeBqJej4_1(.dout(w_dff_A_L7SHkB7f7_1),.din(w_dff_A_NmeBqJej4_1),.clk(gclk));
	jdff dff_B_DqTLLdrs8_0(.din(n1123),.dout(w_dff_B_DqTLLdrs8_0),.clk(gclk));
	jdff dff_B_Hg05mqed6_0(.din(w_dff_B_DqTLLdrs8_0),.dout(w_dff_B_Hg05mqed6_0),.clk(gclk));
	jdff dff_B_4C7GlDBG1_0(.din(w_dff_B_Hg05mqed6_0),.dout(w_dff_B_4C7GlDBG1_0),.clk(gclk));
	jdff dff_B_O1iGWmKO3_0(.din(w_dff_B_4C7GlDBG1_0),.dout(w_dff_B_O1iGWmKO3_0),.clk(gclk));
	jdff dff_B_uIzJ5YwN7_0(.din(w_dff_B_O1iGWmKO3_0),.dout(w_dff_B_uIzJ5YwN7_0),.clk(gclk));
	jdff dff_B_DWi30R3v4_0(.din(w_dff_B_uIzJ5YwN7_0),.dout(w_dff_B_DWi30R3v4_0),.clk(gclk));
	jdff dff_B_DzHoF0Ho2_0(.din(w_dff_B_DWi30R3v4_0),.dout(w_dff_B_DzHoF0Ho2_0),.clk(gclk));
	jdff dff_B_6vc9JUTF5_0(.din(w_dff_B_DzHoF0Ho2_0),.dout(w_dff_B_6vc9JUTF5_0),.clk(gclk));
	jdff dff_B_ipExecNx7_0(.din(w_dff_B_6vc9JUTF5_0),.dout(w_dff_B_ipExecNx7_0),.clk(gclk));
	jdff dff_B_IGY9THnU3_0(.din(w_dff_B_ipExecNx7_0),.dout(w_dff_B_IGY9THnU3_0),.clk(gclk));
	jdff dff_B_dvbZwwhr3_0(.din(w_dff_B_IGY9THnU3_0),.dout(w_dff_B_dvbZwwhr3_0),.clk(gclk));
	jdff dff_B_0gPtaQdm0_0(.din(w_dff_B_dvbZwwhr3_0),.dout(w_dff_B_0gPtaQdm0_0),.clk(gclk));
	jdff dff_B_u5p460Ly0_0(.din(n1122),.dout(w_dff_B_u5p460Ly0_0),.clk(gclk));
	jdff dff_B_vv2nfHoo5_1(.din(n1117),.dout(w_dff_B_vv2nfHoo5_1),.clk(gclk));
	jdff dff_A_Z1lAP6kb0_2(.dout(w_G137_8[2]),.din(w_dff_A_Z1lAP6kb0_2),.clk(gclk));
	jdff dff_A_OZ82CCvQ3_2(.dout(w_dff_A_Z1lAP6kb0_2),.din(w_dff_A_OZ82CCvQ3_2),.clk(gclk));
	jdff dff_A_snODAuqc6_2(.dout(w_dff_A_OZ82CCvQ3_2),.din(w_dff_A_snODAuqc6_2),.clk(gclk));
	jdff dff_B_q1kALwgv4_0(.din(n1132),.dout(w_dff_B_q1kALwgv4_0),.clk(gclk));
	jdff dff_B_Akr5dmJX1_0(.din(w_dff_B_q1kALwgv4_0),.dout(w_dff_B_Akr5dmJX1_0),.clk(gclk));
	jdff dff_B_voAJ6e0B4_0(.din(w_dff_B_Akr5dmJX1_0),.dout(w_dff_B_voAJ6e0B4_0),.clk(gclk));
	jdff dff_B_LbmON4d04_0(.din(w_dff_B_voAJ6e0B4_0),.dout(w_dff_B_LbmON4d04_0),.clk(gclk));
	jdff dff_B_czf60rpt0_0(.din(w_dff_B_LbmON4d04_0),.dout(w_dff_B_czf60rpt0_0),.clk(gclk));
	jdff dff_B_OtENGNYd1_0(.din(w_dff_B_czf60rpt0_0),.dout(w_dff_B_OtENGNYd1_0),.clk(gclk));
	jdff dff_B_6pjDQfW88_0(.din(w_dff_B_OtENGNYd1_0),.dout(w_dff_B_6pjDQfW88_0),.clk(gclk));
	jdff dff_B_nIM3frMz3_0(.din(w_dff_B_6pjDQfW88_0),.dout(w_dff_B_nIM3frMz3_0),.clk(gclk));
	jdff dff_B_sumYEOPg6_0(.din(w_dff_B_nIM3frMz3_0),.dout(w_dff_B_sumYEOPg6_0),.clk(gclk));
	jdff dff_B_wKto22uR8_0(.din(w_dff_B_sumYEOPg6_0),.dout(w_dff_B_wKto22uR8_0),.clk(gclk));
	jdff dff_B_83oAMUNY6_0(.din(w_dff_B_wKto22uR8_0),.dout(w_dff_B_83oAMUNY6_0),.clk(gclk));
	jdff dff_B_0ovZIQyE8_0(.din(w_dff_B_83oAMUNY6_0),.dout(w_dff_B_0ovZIQyE8_0),.clk(gclk));
	jdff dff_B_DHFhcBXc5_0(.din(w_dff_B_0ovZIQyE8_0),.dout(w_dff_B_DHFhcBXc5_0),.clk(gclk));
	jdff dff_B_sFCOBFKZ8_0(.din(n1131),.dout(w_dff_B_sFCOBFKZ8_0),.clk(gclk));
	jdff dff_A_YrGfyymj5_0(.dout(w_n993_3[0]),.din(w_dff_A_YrGfyymj5_0),.clk(gclk));
	jdff dff_A_gamMfp6T9_0(.dout(w_dff_A_YrGfyymj5_0),.din(w_dff_A_gamMfp6T9_0),.clk(gclk));
	jdff dff_A_iXDsf0Av2_1(.dout(w_n993_3[1]),.din(w_dff_A_iXDsf0Av2_1),.clk(gclk));
	jdff dff_B_d44rBEZQ4_1(.din(n1135),.dout(w_dff_B_d44rBEZQ4_1),.clk(gclk));
	jdff dff_B_hLhYhoOa3_1(.din(w_dff_B_d44rBEZQ4_1),.dout(w_dff_B_hLhYhoOa3_1),.clk(gclk));
	jdff dff_B_Kq7EokUD6_1(.din(w_dff_B_hLhYhoOa3_1),.dout(w_dff_B_Kq7EokUD6_1),.clk(gclk));
	jdff dff_B_nSl6TPh82_1(.din(w_dff_B_Kq7EokUD6_1),.dout(w_dff_B_nSl6TPh82_1),.clk(gclk));
	jdff dff_B_dWZPMxOD5_1(.din(w_dff_B_nSl6TPh82_1),.dout(w_dff_B_dWZPMxOD5_1),.clk(gclk));
	jdff dff_B_vhe6go5h3_1(.din(w_dff_B_dWZPMxOD5_1),.dout(w_dff_B_vhe6go5h3_1),.clk(gclk));
	jdff dff_B_VPO1xM0b1_1(.din(w_dff_B_vhe6go5h3_1),.dout(w_dff_B_VPO1xM0b1_1),.clk(gclk));
	jdff dff_B_xl4fjvn14_1(.din(w_dff_B_VPO1xM0b1_1),.dout(w_dff_B_xl4fjvn14_1),.clk(gclk));
	jdff dff_B_prMlvip00_1(.din(w_dff_B_xl4fjvn14_1),.dout(w_dff_B_prMlvip00_1),.clk(gclk));
	jdff dff_B_lB19PUY14_1(.din(w_dff_B_prMlvip00_1),.dout(w_dff_B_lB19PUY14_1),.clk(gclk));
	jdff dff_B_fW7CWBUT3_1(.din(w_dff_B_lB19PUY14_1),.dout(w_dff_B_fW7CWBUT3_1),.clk(gclk));
	jdff dff_B_2bYdIWHR2_1(.din(w_dff_B_fW7CWBUT3_1),.dout(w_dff_B_2bYdIWHR2_1),.clk(gclk));
	jdff dff_B_QlE12RLM6_1(.din(w_dff_B_2bYdIWHR2_1),.dout(w_dff_B_QlE12RLM6_1),.clk(gclk));
	jdff dff_B_lc1B8HQ97_1(.din(w_dff_B_QlE12RLM6_1),.dout(w_dff_B_lc1B8HQ97_1),.clk(gclk));
	jdff dff_B_8HXiJ17M2_1(.din(w_dff_B_lc1B8HQ97_1),.dout(w_dff_B_8HXiJ17M2_1),.clk(gclk));
	jdff dff_B_IbNvrrdT9_1(.din(w_dff_B_8HXiJ17M2_1),.dout(w_dff_B_IbNvrrdT9_1),.clk(gclk));
	jdff dff_B_4rKzi5ft5_1(.din(w_dff_B_IbNvrrdT9_1),.dout(w_dff_B_4rKzi5ft5_1),.clk(gclk));
	jdff dff_B_hr4RBaw75_1(.din(n1136),.dout(w_dff_B_hr4RBaw75_1),.clk(gclk));
	jdff dff_B_JPTkieWH6_1(.din(w_dff_B_hr4RBaw75_1),.dout(w_dff_B_JPTkieWH6_1),.clk(gclk));
	jdff dff_B_JFrPKMCF7_1(.din(w_dff_B_JPTkieWH6_1),.dout(w_dff_B_JFrPKMCF7_1),.clk(gclk));
	jdff dff_B_6bJ5mfPR9_1(.din(w_dff_B_JFrPKMCF7_1),.dout(w_dff_B_6bJ5mfPR9_1),.clk(gclk));
	jdff dff_B_HLYyn1f77_1(.din(w_dff_B_6bJ5mfPR9_1),.dout(w_dff_B_HLYyn1f77_1),.clk(gclk));
	jdff dff_B_7YKmGSuK7_1(.din(w_dff_B_HLYyn1f77_1),.dout(w_dff_B_7YKmGSuK7_1),.clk(gclk));
	jdff dff_B_7lvApMHE8_1(.din(w_dff_B_7YKmGSuK7_1),.dout(w_dff_B_7lvApMHE8_1),.clk(gclk));
	jdff dff_B_ONpsITEh0_1(.din(w_dff_B_7lvApMHE8_1),.dout(w_dff_B_ONpsITEh0_1),.clk(gclk));
	jdff dff_B_9P3iOI6n7_1(.din(w_dff_B_ONpsITEh0_1),.dout(w_dff_B_9P3iOI6n7_1),.clk(gclk));
	jdff dff_B_RWnyobUg6_1(.din(w_dff_B_9P3iOI6n7_1),.dout(w_dff_B_RWnyobUg6_1),.clk(gclk));
	jdff dff_B_KZoARXLc0_1(.din(w_dff_B_RWnyobUg6_1),.dout(w_dff_B_KZoARXLc0_1),.clk(gclk));
	jdff dff_B_FqkfDwMg0_1(.din(w_dff_B_KZoARXLc0_1),.dout(w_dff_B_FqkfDwMg0_1),.clk(gclk));
	jdff dff_B_IDc6rDxQ2_1(.din(w_dff_B_FqkfDwMg0_1),.dout(w_dff_B_IDc6rDxQ2_1),.clk(gclk));
	jdff dff_B_URZBSOEB9_1(.din(w_dff_B_IDc6rDxQ2_1),.dout(w_dff_B_URZBSOEB9_1),.clk(gclk));
	jdff dff_B_mgwEUQS91_1(.din(w_dff_B_URZBSOEB9_1),.dout(w_dff_B_mgwEUQS91_1),.clk(gclk));
	jdff dff_B_sRWC0tdv5_1(.din(w_dff_B_mgwEUQS91_1),.dout(w_dff_B_sRWC0tdv5_1),.clk(gclk));
	jdff dff_B_dzFlQmzL4_1(.din(w_dff_B_sRWC0tdv5_1),.dout(w_dff_B_dzFlQmzL4_1),.clk(gclk));
	jdff dff_B_tuaV0hrY5_1(.din(n811),.dout(w_dff_B_tuaV0hrY5_1),.clk(gclk));
	jdff dff_B_j17Q7vPS0_1(.din(w_dff_B_tuaV0hrY5_1),.dout(w_dff_B_j17Q7vPS0_1),.clk(gclk));
	jdff dff_B_Li0bAqfx2_1(.din(w_dff_B_j17Q7vPS0_1),.dout(w_dff_B_Li0bAqfx2_1),.clk(gclk));
	jdff dff_B_4DN8KS018_1(.din(w_dff_B_Li0bAqfx2_1),.dout(w_dff_B_4DN8KS018_1),.clk(gclk));
	jdff dff_B_T3Kapml73_1(.din(w_dff_B_4DN8KS018_1),.dout(w_dff_B_T3Kapml73_1),.clk(gclk));
	jdff dff_B_H7MzAnXL8_1(.din(w_dff_B_T3Kapml73_1),.dout(w_dff_B_H7MzAnXL8_1),.clk(gclk));
	jdff dff_B_erHClltW3_1(.din(w_dff_B_H7MzAnXL8_1),.dout(w_dff_B_erHClltW3_1),.clk(gclk));
	jdff dff_B_VRr48Sni9_1(.din(w_dff_B_erHClltW3_1),.dout(w_dff_B_VRr48Sni9_1),.clk(gclk));
	jdff dff_B_GjJOhlnr9_1(.din(w_dff_B_VRr48Sni9_1),.dout(w_dff_B_GjJOhlnr9_1),.clk(gclk));
	jdff dff_B_YaNA41sQ1_1(.din(w_dff_B_GjJOhlnr9_1),.dout(w_dff_B_YaNA41sQ1_1),.clk(gclk));
	jdff dff_B_cuEdzt2S1_0(.din(n830),.dout(w_dff_B_cuEdzt2S1_0),.clk(gclk));
	jdff dff_B_LPgtyoLW5_0(.din(w_dff_B_cuEdzt2S1_0),.dout(w_dff_B_LPgtyoLW5_0),.clk(gclk));
	jdff dff_B_uYNAnF3P9_0(.din(w_dff_B_LPgtyoLW5_0),.dout(w_dff_B_uYNAnF3P9_0),.clk(gclk));
	jdff dff_B_TTI3V0c07_0(.din(w_dff_B_uYNAnF3P9_0),.dout(w_dff_B_TTI3V0c07_0),.clk(gclk));
	jdff dff_B_0LeQCjqX9_0(.din(w_dff_B_TTI3V0c07_0),.dout(w_dff_B_0LeQCjqX9_0),.clk(gclk));
	jdff dff_B_hGo6aE1L4_0(.din(w_dff_B_0LeQCjqX9_0),.dout(w_dff_B_hGo6aE1L4_0),.clk(gclk));
	jdff dff_B_vrHzVBPs5_1(.din(n441),.dout(w_dff_B_vrHzVBPs5_1),.clk(gclk));
	jdff dff_B_8P1YGzgQ2_1(.din(n436),.dout(w_dff_B_8P1YGzgQ2_1),.clk(gclk));
	jdff dff_B_Quo6qYtP7_1(.din(n822),.dout(w_dff_B_Quo6qYtP7_1),.clk(gclk));
	jdff dff_B_oUcrpXRb4_1(.din(w_dff_B_Quo6qYtP7_1),.dout(w_dff_B_oUcrpXRb4_1),.clk(gclk));
	jdff dff_B_vAZPEblA7_1(.din(w_dff_B_oUcrpXRb4_1),.dout(w_dff_B_vAZPEblA7_1),.clk(gclk));
	jdff dff_B_iQPIcCBI1_1(.din(w_dff_B_vAZPEblA7_1),.dout(w_dff_B_iQPIcCBI1_1),.clk(gclk));
	jdff dff_B_qwPBKtuU9_1(.din(w_dff_B_iQPIcCBI1_1),.dout(w_dff_B_qwPBKtuU9_1),.clk(gclk));
	jdff dff_B_7ursiyCr0_1(.din(G52),.dout(w_dff_B_7ursiyCr0_1),.clk(gclk));
	jdff dff_B_9EyVRvmn8_1(.din(w_dff_B_7ursiyCr0_1),.dout(w_dff_B_9EyVRvmn8_1),.clk(gclk));
	jdff dff_B_DUiIQvWy4_1(.din(n864),.dout(w_dff_B_DUiIQvWy4_1),.clk(gclk));
	jdff dff_B_WTgw8wve6_1(.din(w_dff_B_DUiIQvWy4_1),.dout(w_dff_B_WTgw8wve6_1),.clk(gclk));
	jdff dff_B_7O6ie4Ck9_1(.din(w_dff_B_WTgw8wve6_1),.dout(w_dff_B_7O6ie4Ck9_1),.clk(gclk));
	jdff dff_B_Ni0PLMRt2_1(.din(w_dff_B_7O6ie4Ck9_1),.dout(w_dff_B_Ni0PLMRt2_1),.clk(gclk));
	jdff dff_B_VfuJOKvu7_1(.din(w_dff_B_Ni0PLMRt2_1),.dout(w_dff_B_VfuJOKvu7_1),.clk(gclk));
	jdff dff_B_ujPWr6ve6_1(.din(w_dff_B_VfuJOKvu7_1),.dout(w_dff_B_ujPWr6ve6_1),.clk(gclk));
	jdff dff_B_rbAuemPE9_1(.din(w_dff_B_ujPWr6ve6_1),.dout(w_dff_B_rbAuemPE9_1),.clk(gclk));
	jdff dff_B_3TGk4T0w7_1(.din(w_dff_B_rbAuemPE9_1),.dout(w_dff_B_3TGk4T0w7_1),.clk(gclk));
	jdff dff_B_ZBum0YOh9_1(.din(w_dff_B_3TGk4T0w7_1),.dout(w_dff_B_ZBum0YOh9_1),.clk(gclk));
	jdff dff_B_mRm8lSLm3_1(.din(w_dff_B_ZBum0YOh9_1),.dout(w_dff_B_mRm8lSLm3_1),.clk(gclk));
	jdff dff_B_FXetr5Jf8_0(.din(n874),.dout(w_dff_B_FXetr5Jf8_0),.clk(gclk));
	jdff dff_B_bj1sZqhK9_0(.din(w_dff_B_FXetr5Jf8_0),.dout(w_dff_B_bj1sZqhK9_0),.clk(gclk));
	jdff dff_B_ZzupltTq5_0(.din(w_dff_B_bj1sZqhK9_0),.dout(w_dff_B_ZzupltTq5_0),.clk(gclk));
	jdff dff_B_RCQ0KC3s0_0(.din(w_dff_B_ZzupltTq5_0),.dout(w_dff_B_RCQ0KC3s0_0),.clk(gclk));
	jdff dff_B_PbjgCsSE0_0(.din(w_dff_B_RCQ0KC3s0_0),.dout(w_dff_B_PbjgCsSE0_0),.clk(gclk));
	jdff dff_B_ZIzc92Bh0_0(.din(w_dff_B_PbjgCsSE0_0),.dout(w_dff_B_ZIzc92Bh0_0),.clk(gclk));
	jdff dff_B_AKBIMfoM4_1(.din(n466),.dout(w_dff_B_AKBIMfoM4_1),.clk(gclk));
	jdff dff_B_VkR0RJnO3_1(.din(n461),.dout(w_dff_B_VkR0RJnO3_1),.clk(gclk));
	jdff dff_B_YoXDgICp1_1(.din(G122),.dout(w_dff_B_YoXDgICp1_1),.clk(gclk));
	jdff dff_B_7UNUH5rp2_1(.din(w_dff_B_YoXDgICp1_1),.dout(w_dff_B_7UNUH5rp2_1),.clk(gclk));
	jdff dff_B_o2AF7ZD13_2(.din(G170),.dout(w_dff_B_o2AF7ZD13_2),.clk(gclk));
	jdff dff_B_kgOnxlfu9_2(.din(G200),.dout(w_dff_B_kgOnxlfu9_2),.clk(gclk));
	jdff dff_B_O2epEFNI8_2(.din(w_dff_B_kgOnxlfu9_2),.dout(w_dff_B_O2epEFNI8_2),.clk(gclk));
	jdff dff_B_zdIME7Wv5_0(.din(n1150),.dout(w_dff_B_zdIME7Wv5_0),.clk(gclk));
	jdff dff_B_0t4XAYSf0_0(.din(w_dff_B_zdIME7Wv5_0),.dout(w_dff_B_0t4XAYSf0_0),.clk(gclk));
	jdff dff_B_kdRm8gLu1_0(.din(w_dff_B_0t4XAYSf0_0),.dout(w_dff_B_kdRm8gLu1_0),.clk(gclk));
	jdff dff_B_M5D640MM2_0(.din(w_dff_B_kdRm8gLu1_0),.dout(w_dff_B_M5D640MM2_0),.clk(gclk));
	jdff dff_B_TnHaRBC44_0(.din(w_dff_B_M5D640MM2_0),.dout(w_dff_B_TnHaRBC44_0),.clk(gclk));
	jdff dff_B_2hFp0IYO8_0(.din(w_dff_B_TnHaRBC44_0),.dout(w_dff_B_2hFp0IYO8_0),.clk(gclk));
	jdff dff_B_D4dwODuW2_0(.din(w_dff_B_2hFp0IYO8_0),.dout(w_dff_B_D4dwODuW2_0),.clk(gclk));
	jdff dff_B_bUX2u2H59_0(.din(w_dff_B_D4dwODuW2_0),.dout(w_dff_B_bUX2u2H59_0),.clk(gclk));
	jdff dff_B_9KqjEjrP8_0(.din(w_dff_B_bUX2u2H59_0),.dout(w_dff_B_9KqjEjrP8_0),.clk(gclk));
	jdff dff_B_7o2KHG086_0(.din(w_dff_B_9KqjEjrP8_0),.dout(w_dff_B_7o2KHG086_0),.clk(gclk));
	jdff dff_B_oQ8gKiWd9_0(.din(w_dff_B_7o2KHG086_0),.dout(w_dff_B_oQ8gKiWd9_0),.clk(gclk));
	jdff dff_B_9vShPgtL7_0(.din(w_dff_B_oQ8gKiWd9_0),.dout(w_dff_B_9vShPgtL7_0),.clk(gclk));
	jdff dff_B_iKYzvaD16_0(.din(n1149),.dout(w_dff_B_iKYzvaD16_0),.clk(gclk));
	jdff dff_B_SJjDmDZT6_2(.din(G158),.dout(w_dff_B_SJjDmDZT6_2),.clk(gclk));
	jdff dff_B_bsAacwTI8_2(.din(G188),.dout(w_dff_B_bsAacwTI8_2),.clk(gclk));
	jdff dff_B_K9zwZyi23_2(.din(w_dff_B_bsAacwTI8_2),.dout(w_dff_B_K9zwZyi23_2),.clk(gclk));
	jdff dff_B_metFiBlD4_0(.din(n1146),.dout(w_dff_B_metFiBlD4_0),.clk(gclk));
	jdff dff_B_XEBaaWNY0_1(.din(n897),.dout(w_dff_B_XEBaaWNY0_1),.clk(gclk));
	jdff dff_B_cWW7BqkY5_1(.din(w_dff_B_XEBaaWNY0_1),.dout(w_dff_B_cWW7BqkY5_1),.clk(gclk));
	jdff dff_B_FT55muRm4_1(.din(w_dff_B_cWW7BqkY5_1),.dout(w_dff_B_FT55muRm4_1),.clk(gclk));
	jdff dff_B_P2bFHe5K8_1(.din(w_dff_B_FT55muRm4_1),.dout(w_dff_B_P2bFHe5K8_1),.clk(gclk));
	jdff dff_B_4UIEkQYb6_1(.din(w_dff_B_P2bFHe5K8_1),.dout(w_dff_B_4UIEkQYb6_1),.clk(gclk));
	jdff dff_B_VwpLRZYF3_1(.din(w_dff_B_4UIEkQYb6_1),.dout(w_dff_B_VwpLRZYF3_1),.clk(gclk));
	jdff dff_B_GtsUyFiA0_0(.din(n904),.dout(w_dff_B_GtsUyFiA0_0),.clk(gclk));
	jdff dff_B_S49bTiMW9_0(.din(w_dff_B_GtsUyFiA0_0),.dout(w_dff_B_S49bTiMW9_0),.clk(gclk));
	jdff dff_B_RLUsb3Cv4_1(.din(n477),.dout(w_dff_B_RLUsb3Cv4_1),.clk(gclk));
	jdff dff_B_z12meKbH6_1(.din(n472),.dout(w_dff_B_z12meKbH6_1),.clk(gclk));
	jdff dff_A_0VM845kW6_0(.dout(w_n901_0[0]),.din(w_dff_A_0VM845kW6_0),.clk(gclk));
	jdff dff_A_EsAjOgU65_0(.dout(w_dff_A_0VM845kW6_0),.din(w_dff_A_EsAjOgU65_0),.clk(gclk));
	jdff dff_B_eJ69Mfy49_1(.din(n898),.dout(w_dff_B_eJ69Mfy49_1),.clk(gclk));
	jdff dff_B_uLwGAIUX9_1(.din(G126),.dout(w_dff_B_uLwGAIUX9_1),.clk(gclk));
	jdff dff_B_PS2S0xBY7_1(.din(w_dff_B_uLwGAIUX9_1),.dout(w_dff_B_PS2S0xBY7_1),.clk(gclk));
	jdff dff_A_npS2ivQk8_0(.dout(w_n1007_3[0]),.din(w_dff_A_npS2ivQk8_0),.clk(gclk));
	jdff dff_A_IqrBrl157_1(.dout(w_n1007_3[1]),.din(w_dff_A_IqrBrl157_1),.clk(gclk));
	jdff dff_A_U4fR8iQ06_1(.dout(w_dff_A_IqrBrl157_1),.din(w_dff_A_U4fR8iQ06_1),.clk(gclk));
	jdff dff_A_2xgFELTQ7_1(.dout(w_dff_A_U4fR8iQ06_1),.din(w_dff_A_2xgFELTQ7_1),.clk(gclk));
	jdff dff_A_tGcLAQFM9_1(.dout(w_dff_A_2xgFELTQ7_1),.din(w_dff_A_tGcLAQFM9_1),.clk(gclk));
	jdff dff_A_CX0tG5144_1(.dout(w_dff_A_tGcLAQFM9_1),.din(w_dff_A_CX0tG5144_1),.clk(gclk));
	jdff dff_A_6u7w5u6X9_1(.dout(w_dff_A_CX0tG5144_1),.din(w_dff_A_6u7w5u6X9_1),.clk(gclk));
	jdff dff_B_tlusE0j86_1(.din(n762),.dout(w_dff_B_tlusE0j86_1),.clk(gclk));
	jdff dff_B_sWwHpGJt0_1(.din(w_dff_B_tlusE0j86_1),.dout(w_dff_B_sWwHpGJt0_1),.clk(gclk));
	jdff dff_B_GuCnLKnr4_1(.din(w_dff_B_sWwHpGJt0_1),.dout(w_dff_B_GuCnLKnr4_1),.clk(gclk));
	jdff dff_B_4J9ddOpI5_1(.din(w_dff_B_GuCnLKnr4_1),.dout(w_dff_B_4J9ddOpI5_1),.clk(gclk));
	jdff dff_B_HlcYQuNT3_1(.din(w_dff_B_4J9ddOpI5_1),.dout(w_dff_B_HlcYQuNT3_1),.clk(gclk));
	jdff dff_B_c1L8sULW9_1(.din(w_dff_B_HlcYQuNT3_1),.dout(w_dff_B_c1L8sULW9_1),.clk(gclk));
	jdff dff_B_p49FRbal8_1(.din(w_dff_B_c1L8sULW9_1),.dout(w_dff_B_p49FRbal8_1),.clk(gclk));
	jdff dff_B_ZbyInzDL9_1(.din(w_dff_B_p49FRbal8_1),.dout(w_dff_B_ZbyInzDL9_1),.clk(gclk));
	jdff dff_B_iVd2sr9e1_0(.din(n773),.dout(w_dff_B_iVd2sr9e1_0),.clk(gclk));
	jdff dff_B_yRqSM7OQ3_0(.din(w_dff_B_iVd2sr9e1_0),.dout(w_dff_B_yRqSM7OQ3_0),.clk(gclk));
	jdff dff_B_LoDdlt7O8_0(.din(w_dff_B_yRqSM7OQ3_0),.dout(w_dff_B_LoDdlt7O8_0),.clk(gclk));
	jdff dff_B_HGmizWoM4_0(.din(w_dff_B_LoDdlt7O8_0),.dout(w_dff_B_HGmizWoM4_0),.clk(gclk));
	jdff dff_B_oZOwAB332_1(.din(n382),.dout(w_dff_B_oZOwAB332_1),.clk(gclk));
	jdff dff_B_hamSiRHx7_1(.din(n376),.dout(w_dff_B_hamSiRHx7_1),.clk(gclk));
	jdff dff_B_5IjkzF0r0_0(.din(n769),.dout(w_dff_B_5IjkzF0r0_0),.clk(gclk));
	jdff dff_B_7wNVapkp3_0(.din(w_dff_B_5IjkzF0r0_0),.dout(w_dff_B_7wNVapkp3_0),.clk(gclk));
	jdff dff_B_kJmmPrrk2_0(.din(w_dff_B_7wNVapkp3_0),.dout(w_dff_B_kJmmPrrk2_0),.clk(gclk));
	jdff dff_B_vFdVfgzK6_0(.din(w_dff_B_kJmmPrrk2_0),.dout(w_dff_B_vFdVfgzK6_0),.clk(gclk));
	jdff dff_A_B0xsdXZn9_0(.dout(w_n753_1[0]),.din(w_dff_A_B0xsdXZn9_0),.clk(gclk));
	jdff dff_A_OTKIU66v7_0(.dout(w_dff_A_B0xsdXZn9_0),.din(w_dff_A_OTKIU66v7_0),.clk(gclk));
	jdff dff_A_YV5OdHI91_0(.dout(w_dff_A_OTKIU66v7_0),.din(w_dff_A_YV5OdHI91_0),.clk(gclk));
	jdff dff_A_PPiBdDlg1_0(.dout(w_dff_A_YV5OdHI91_0),.din(w_dff_A_PPiBdDlg1_0),.clk(gclk));
	jdff dff_A_xrLt9rQJ6_0(.dout(w_dff_A_PPiBdDlg1_0),.din(w_dff_A_xrLt9rQJ6_0),.clk(gclk));
	jdff dff_A_TwveDcUk1_0(.dout(w_G4091_5[0]),.din(w_dff_A_TwveDcUk1_0),.clk(gclk));
	jdff dff_A_YM1cTB718_0(.dout(w_dff_A_TwveDcUk1_0),.din(w_dff_A_YM1cTB718_0),.clk(gclk));
	jdff dff_A_5cmZxVG40_0(.dout(w_dff_A_YM1cTB718_0),.din(w_dff_A_5cmZxVG40_0),.clk(gclk));
	jdff dff_A_9W5ELkMv7_0(.dout(w_dff_A_5cmZxVG40_0),.din(w_dff_A_9W5ELkMv7_0),.clk(gclk));
	jdff dff_A_xhrFUx5g6_0(.dout(w_dff_A_9W5ELkMv7_0),.din(w_dff_A_xhrFUx5g6_0),.clk(gclk));
	jdff dff_A_K8kkhlAe6_2(.dout(w_G4091_5[2]),.din(w_dff_A_K8kkhlAe6_2),.clk(gclk));
	jdff dff_A_dO3Ntust9_2(.dout(w_dff_A_K8kkhlAe6_2),.din(w_dff_A_dO3Ntust9_2),.clk(gclk));
	jdff dff_A_2hM6Ucfa7_2(.dout(w_dff_A_dO3Ntust9_2),.din(w_dff_A_2hM6Ucfa7_2),.clk(gclk));
	jdff dff_B_tGjzBN9i0_1(.din(G129),.dout(w_dff_B_tGjzBN9i0_1),.clk(gclk));
	jdff dff_B_NJuNj2kG9_1(.din(w_dff_B_tGjzBN9i0_1),.dout(w_dff_B_NJuNj2kG9_1),.clk(gclk));
	jdff dff_A_NnsPrOqX9_1(.dout(w_G137_7[1]),.din(w_dff_A_NnsPrOqX9_1),.clk(gclk));
	jdff dff_A_qQP3m4jI7_1(.dout(w_dff_A_NnsPrOqX9_1),.din(w_dff_A_qQP3m4jI7_1),.clk(gclk));
	jdff dff_A_0NMZDrI95_1(.dout(w_dff_A_qQP3m4jI7_1),.din(w_dff_A_0NMZDrI95_1),.clk(gclk));
	jdff dff_A_gGGJZbzA5_1(.dout(w_dff_A_0NMZDrI95_1),.din(w_dff_A_gGGJZbzA5_1),.clk(gclk));
	jdff dff_A_GGM1gy4q7_2(.dout(w_G137_7[2]),.din(w_dff_A_GGM1gy4q7_2),.clk(gclk));
	jdff dff_A_D9Wcx2QM8_0(.dout(w_G137_2[0]),.din(w_dff_A_D9Wcx2QM8_0),.clk(gclk));
	jdff dff_A_vfZVX75W4_0(.dout(w_dff_A_D9Wcx2QM8_0),.din(w_dff_A_vfZVX75W4_0),.clk(gclk));
	jdff dff_A_bdDwh1Wl4_1(.dout(w_G137_2[1]),.din(w_dff_A_bdDwh1Wl4_1),.clk(gclk));
	jdff dff_A_Jw5QYtyr4_1(.dout(w_dff_A_bdDwh1Wl4_1),.din(w_dff_A_Jw5QYtyr4_1),.clk(gclk));
	jdff dff_B_CUT3gRE58_0(.din(n1159),.dout(w_dff_B_CUT3gRE58_0),.clk(gclk));
	jdff dff_B_bWLS9a6V2_0(.din(w_dff_B_CUT3gRE58_0),.dout(w_dff_B_bWLS9a6V2_0),.clk(gclk));
	jdff dff_B_vI2VsaJz9_0(.din(w_dff_B_bWLS9a6V2_0),.dout(w_dff_B_vI2VsaJz9_0),.clk(gclk));
	jdff dff_B_zGKyLPLR5_0(.din(w_dff_B_vI2VsaJz9_0),.dout(w_dff_B_zGKyLPLR5_0),.clk(gclk));
	jdff dff_B_0XECho6T1_0(.din(w_dff_B_zGKyLPLR5_0),.dout(w_dff_B_0XECho6T1_0),.clk(gclk));
	jdff dff_B_0ZMRQjxo5_0(.din(w_dff_B_0XECho6T1_0),.dout(w_dff_B_0ZMRQjxo5_0),.clk(gclk));
	jdff dff_B_Ce7ze7A05_0(.din(w_dff_B_0ZMRQjxo5_0),.dout(w_dff_B_Ce7ze7A05_0),.clk(gclk));
	jdff dff_B_04LfTljs7_0(.din(w_dff_B_Ce7ze7A05_0),.dout(w_dff_B_04LfTljs7_0),.clk(gclk));
	jdff dff_B_5FLfSNxX5_0(.din(w_dff_B_04LfTljs7_0),.dout(w_dff_B_5FLfSNxX5_0),.clk(gclk));
	jdff dff_B_E4IgnFj56_0(.din(w_dff_B_5FLfSNxX5_0),.dout(w_dff_B_E4IgnFj56_0),.clk(gclk));
	jdff dff_B_0spYFI720_0(.din(w_dff_B_E4IgnFj56_0),.dout(w_dff_B_0spYFI720_0),.clk(gclk));
	jdff dff_B_0FbXlvoh7_0(.din(w_dff_B_0spYFI720_0),.dout(w_dff_B_0FbXlvoh7_0),.clk(gclk));
	jdff dff_B_kwmSNrEv6_0(.din(n1158),.dout(w_dff_B_kwmSNrEv6_0),.clk(gclk));
	jdff dff_B_8AGxI0Mu5_2(.din(G152),.dout(w_dff_B_8AGxI0Mu5_2),.clk(gclk));
	jdff dff_B_ASVoifaa9_2(.din(G155),.dout(w_dff_B_ASVoifaa9_2),.clk(gclk));
	jdff dff_B_Ajmd820Z0_2(.din(w_dff_B_ASVoifaa9_2),.dout(w_dff_B_Ajmd820Z0_2),.clk(gclk));
	jdff dff_B_EFBbqyKg0_1(.din(n1153),.dout(w_dff_B_EFBbqyKg0_1),.clk(gclk));
	jdff dff_B_NuMGKBgK4_1(.din(n887),.dout(w_dff_B_NuMGKBgK4_1),.clk(gclk));
	jdff dff_B_fIKJ2Mgp5_1(.din(w_dff_B_NuMGKBgK4_1),.dout(w_dff_B_fIKJ2Mgp5_1),.clk(gclk));
	jdff dff_B_d4z54aPe4_1(.din(w_dff_B_fIKJ2Mgp5_1),.dout(w_dff_B_d4z54aPe4_1),.clk(gclk));
	jdff dff_B_MylFQXjh9_1(.din(w_dff_B_d4z54aPe4_1),.dout(w_dff_B_MylFQXjh9_1),.clk(gclk));
	jdff dff_B_hWOXd6XA6_1(.din(w_dff_B_MylFQXjh9_1),.dout(w_dff_B_hWOXd6XA6_1),.clk(gclk));
	jdff dff_B_Periazxo7_1(.din(w_dff_B_hWOXd6XA6_1),.dout(w_dff_B_Periazxo7_1),.clk(gclk));
	jdff dff_B_9P4ED7zy1_1(.din(w_dff_B_Periazxo7_1),.dout(w_dff_B_9P4ED7zy1_1),.clk(gclk));
	jdff dff_B_U8M86RnQ3_0(.din(n893),.dout(w_dff_B_U8M86RnQ3_0),.clk(gclk));
	jdff dff_B_gBzeg0a72_0(.din(w_dff_B_U8M86RnQ3_0),.dout(w_dff_B_gBzeg0a72_0),.clk(gclk));
	jdff dff_B_I1dON0uH7_0(.din(w_dff_B_gBzeg0a72_0),.dout(w_dff_B_I1dON0uH7_0),.clk(gclk));
	jdff dff_B_ugITFTmU9_1(.din(n489),.dout(w_dff_B_ugITFTmU9_1),.clk(gclk));
	jdff dff_B_ybO4WRJc4_1(.din(n484),.dout(w_dff_B_ybO4WRJc4_1),.clk(gclk));
	jdff dff_B_8U0Oim1p9_1(.din(G127),.dout(w_dff_B_8U0Oim1p9_1),.clk(gclk));
	jdff dff_B_l6Ij8nIr3_1(.din(w_dff_B_8U0Oim1p9_1),.dout(w_dff_B_l6Ij8nIr3_1),.clk(gclk));
	jdff dff_B_CG8aC8g90_1(.din(n843),.dout(w_dff_B_CG8aC8g90_1),.clk(gclk));
	jdff dff_B_onHZEBtR5_1(.din(w_dff_B_CG8aC8g90_1),.dout(w_dff_B_onHZEBtR5_1),.clk(gclk));
	jdff dff_B_B3Sll7g45_1(.din(w_dff_B_onHZEBtR5_1),.dout(w_dff_B_B3Sll7g45_1),.clk(gclk));
	jdff dff_B_HHaPyPg73_1(.din(w_dff_B_B3Sll7g45_1),.dout(w_dff_B_HHaPyPg73_1),.clk(gclk));
	jdff dff_B_fieNrXQD7_1(.din(w_dff_B_HHaPyPg73_1),.dout(w_dff_B_fieNrXQD7_1),.clk(gclk));
	jdff dff_B_BFd0Oyoi6_1(.din(w_dff_B_fieNrXQD7_1),.dout(w_dff_B_BFd0Oyoi6_1),.clk(gclk));
	jdff dff_B_Pg0Xh79Q8_1(.din(w_dff_B_BFd0Oyoi6_1),.dout(w_dff_B_Pg0Xh79Q8_1),.clk(gclk));
	jdff dff_B_8rQ7rliv3_1(.din(n844),.dout(w_dff_B_8rQ7rliv3_1),.clk(gclk));
	jdff dff_B_LxXzK1Q48_1(.din(w_dff_B_8rQ7rliv3_1),.dout(w_dff_B_LxXzK1Q48_1),.clk(gclk));
	jdff dff_B_OEziAhiQ8_1(.din(w_dff_B_LxXzK1Q48_1),.dout(w_dff_B_OEziAhiQ8_1),.clk(gclk));
	jdff dff_B_sStGSEa44_1(.din(w_dff_B_OEziAhiQ8_1),.dout(w_dff_B_sStGSEa44_1),.clk(gclk));
	jdff dff_A_SwyMxSwn5_0(.dout(w_n847_0[0]),.din(w_dff_A_SwyMxSwn5_0),.clk(gclk));
	jdff dff_A_K1FPsr598_0(.dout(w_dff_A_SwyMxSwn5_0),.din(w_dff_A_K1FPsr598_0),.clk(gclk));
	jdff dff_A_FL9tvQGF9_0(.dout(w_dff_A_K1FPsr598_0),.din(w_dff_A_FL9tvQGF9_0),.clk(gclk));
	jdff dff_A_yezpWkaN3_0(.dout(w_dff_A_FL9tvQGF9_0),.din(w_dff_A_yezpWkaN3_0),.clk(gclk));
	jdff dff_A_3lqhmAhK7_0(.dout(w_dff_A_yezpWkaN3_0),.din(w_dff_A_3lqhmAhK7_0),.clk(gclk));
	jdff dff_B_90WGFX200_1(.din(n393),.dout(w_dff_B_90WGFX200_1),.clk(gclk));
	jdff dff_B_WTvEmP2Q3_1(.din(n388),.dout(w_dff_B_WTvEmP2Q3_1),.clk(gclk));
	jdff dff_B_gCPz57zM4_1(.din(G119),.dout(w_dff_B_gCPz57zM4_1),.clk(gclk));
	jdff dff_B_7640OupI3_1(.din(w_dff_B_gCPz57zM4_1),.dout(w_dff_B_7640OupI3_1),.clk(gclk));
	jdff dff_B_RnR6lCWr1_0(.din(n1168),.dout(w_dff_B_RnR6lCWr1_0),.clk(gclk));
	jdff dff_B_bk9oqwj17_0(.din(w_dff_B_RnR6lCWr1_0),.dout(w_dff_B_bk9oqwj17_0),.clk(gclk));
	jdff dff_B_zjR3F0PZ6_0(.din(w_dff_B_bk9oqwj17_0),.dout(w_dff_B_zjR3F0PZ6_0),.clk(gclk));
	jdff dff_B_uAVllWra0_0(.din(w_dff_B_zjR3F0PZ6_0),.dout(w_dff_B_uAVllWra0_0),.clk(gclk));
	jdff dff_B_RU9gjels2_0(.din(w_dff_B_uAVllWra0_0),.dout(w_dff_B_RU9gjels2_0),.clk(gclk));
	jdff dff_B_vNbCm1wf4_0(.din(w_dff_B_RU9gjels2_0),.dout(w_dff_B_vNbCm1wf4_0),.clk(gclk));
	jdff dff_B_sczV63Oz7_0(.din(w_dff_B_vNbCm1wf4_0),.dout(w_dff_B_sczV63Oz7_0),.clk(gclk));
	jdff dff_B_TU8pH5Wq5_0(.din(w_dff_B_sczV63Oz7_0),.dout(w_dff_B_TU8pH5Wq5_0),.clk(gclk));
	jdff dff_B_pA0nuJHF3_0(.din(w_dff_B_TU8pH5Wq5_0),.dout(w_dff_B_pA0nuJHF3_0),.clk(gclk));
	jdff dff_B_iecZB5iN5_0(.din(w_dff_B_pA0nuJHF3_0),.dout(w_dff_B_iecZB5iN5_0),.clk(gclk));
	jdff dff_B_EaveTiGR9_0(.din(w_dff_B_iecZB5iN5_0),.dout(w_dff_B_EaveTiGR9_0),.clk(gclk));
	jdff dff_B_I7cht51M1_0(.din(w_dff_B_EaveTiGR9_0),.dout(w_dff_B_I7cht51M1_0),.clk(gclk));
	jdff dff_B_MEIhhaKH4_0(.din(w_dff_B_I7cht51M1_0),.dout(w_dff_B_MEIhhaKH4_0),.clk(gclk));
	jdff dff_B_l83lBKCX4_0(.din(n1167),.dout(w_dff_B_l83lBKCX4_0),.clk(gclk));
	jdff dff_B_ZI5yvDHv8_2(.din(G146),.dout(w_dff_B_ZI5yvDHv8_2),.clk(gclk));
	jdff dff_B_BiHPPjJQ1_2(.din(G149),.dout(w_dff_B_BiHPPjJQ1_2),.clk(gclk));
	jdff dff_B_t5CF08rg6_2(.din(w_dff_B_BiHPPjJQ1_2),.dout(w_dff_B_t5CF08rg6_2),.clk(gclk));
	jdff dff_B_UXzmJdT80_1(.din(n878),.dout(w_dff_B_UXzmJdT80_1),.clk(gclk));
	jdff dff_B_gGE7O5iU9_1(.din(w_dff_B_UXzmJdT80_1),.dout(w_dff_B_gGE7O5iU9_1),.clk(gclk));
	jdff dff_B_hU0SneQp0_1(.din(w_dff_B_gGE7O5iU9_1),.dout(w_dff_B_hU0SneQp0_1),.clk(gclk));
	jdff dff_B_VzT1cfgR9_1(.din(w_dff_B_hU0SneQp0_1),.dout(w_dff_B_VzT1cfgR9_1),.clk(gclk));
	jdff dff_B_I7I4M44f4_1(.din(w_dff_B_VzT1cfgR9_1),.dout(w_dff_B_I7I4M44f4_1),.clk(gclk));
	jdff dff_B_3lXXAADx3_1(.din(w_dff_B_I7I4M44f4_1),.dout(w_dff_B_3lXXAADx3_1),.clk(gclk));
	jdff dff_B_GTMGHZwB8_1(.din(w_dff_B_3lXXAADx3_1),.dout(w_dff_B_GTMGHZwB8_1),.clk(gclk));
	jdff dff_B_c9O17rgw7_1(.din(w_dff_B_GTMGHZwB8_1),.dout(w_dff_B_c9O17rgw7_1),.clk(gclk));
	jdff dff_B_Ej5h7qih9_0(.din(n883),.dout(w_dff_B_Ej5h7qih9_0),.clk(gclk));
	jdff dff_B_KpAM97bC1_0(.din(w_dff_B_Ej5h7qih9_0),.dout(w_dff_B_KpAM97bC1_0),.clk(gclk));
	jdff dff_B_h8VxbfjI7_0(.din(w_dff_B_KpAM97bC1_0),.dout(w_dff_B_h8VxbfjI7_0),.clk(gclk));
	jdff dff_B_wazcHJKO4_0(.din(w_dff_B_h8VxbfjI7_0),.dout(w_dff_B_wazcHJKO4_0),.clk(gclk));
	jdff dff_B_Ib7fXhQc1_1(.din(n524),.dout(w_dff_B_Ib7fXhQc1_1),.clk(gclk));
	jdff dff_B_kZQ8zMyd6_1(.din(n519),.dout(w_dff_B_kZQ8zMyd6_1),.clk(gclk));
	jdff dff_A_rNiPtXLH8_2(.dout(w_G4092_7[2]),.din(w_dff_A_rNiPtXLH8_2),.clk(gclk));
	jdff dff_A_3aedCEev1_2(.dout(w_dff_A_rNiPtXLH8_2),.din(w_dff_A_3aedCEev1_2),.clk(gclk));
	jdff dff_A_QMPVijS82_2(.dout(w_dff_A_3aedCEev1_2),.din(w_dff_A_QMPVijS82_2),.clk(gclk));
	jdff dff_A_GZeO6MGe9_0(.dout(w_n880_0[0]),.din(w_dff_A_GZeO6MGe9_0),.clk(gclk));
	jdff dff_A_0WMH8yzG8_0(.dout(w_dff_A_GZeO6MGe9_0),.din(w_dff_A_0WMH8yzG8_0),.clk(gclk));
	jdff dff_A_cdAeYYAu1_0(.dout(w_dff_A_0WMH8yzG8_0),.din(w_dff_A_cdAeYYAu1_0),.clk(gclk));
	jdff dff_A_bIIZgxBS9_0(.dout(w_dff_A_cdAeYYAu1_0),.din(w_dff_A_bIIZgxBS9_0),.clk(gclk));
	jdff dff_A_Pp1HGQRd6_0(.dout(w_dff_A_bIIZgxBS9_0),.din(w_dff_A_Pp1HGQRd6_0),.clk(gclk));
	jdff dff_A_za0xKMAC7_1(.dout(w_G4091_3[1]),.din(w_dff_A_za0xKMAC7_1),.clk(gclk));
	jdff dff_A_7WVyANtA8_2(.dout(w_G4091_3[2]),.din(w_dff_A_7WVyANtA8_2),.clk(gclk));
	jdff dff_A_Yv7YRBAz8_2(.dout(w_dff_A_7WVyANtA8_2),.din(w_dff_A_Yv7YRBAz8_2),.clk(gclk));
	jdff dff_B_u4wgZrrl9_1(.din(G128),.dout(w_dff_B_u4wgZrrl9_1),.clk(gclk));
	jdff dff_B_e7Aq2xOM1_1(.din(w_dff_B_u4wgZrrl9_1),.dout(w_dff_B_e7Aq2xOM1_1),.clk(gclk));
	jdff dff_A_0V2656ta9_0(.dout(w_n1008_3[0]),.din(w_dff_A_0V2656ta9_0),.clk(gclk));
	jdff dff_A_QiqEtPaT6_0(.dout(w_dff_A_0V2656ta9_0),.din(w_dff_A_QiqEtPaT6_0),.clk(gclk));
	jdff dff_A_LWUS1reT6_1(.dout(w_n1008_3[1]),.din(w_dff_A_LWUS1reT6_1),.clk(gclk));
	jdff dff_B_l3iQHOaA7_1(.din(n834),.dout(w_dff_B_l3iQHOaA7_1),.clk(gclk));
	jdff dff_B_2JDzgvY80_1(.din(w_dff_B_l3iQHOaA7_1),.dout(w_dff_B_2JDzgvY80_1),.clk(gclk));
	jdff dff_B_X9qMtqnv1_1(.din(w_dff_B_2JDzgvY80_1),.dout(w_dff_B_X9qMtqnv1_1),.clk(gclk));
	jdff dff_B_Y1iIcmNt6_1(.din(w_dff_B_X9qMtqnv1_1),.dout(w_dff_B_Y1iIcmNt6_1),.clk(gclk));
	jdff dff_B_0f47Wv3m5_1(.din(w_dff_B_Y1iIcmNt6_1),.dout(w_dff_B_0f47Wv3m5_1),.clk(gclk));
	jdff dff_B_At1YA5Vh4_1(.din(w_dff_B_0f47Wv3m5_1),.dout(w_dff_B_At1YA5Vh4_1),.clk(gclk));
	jdff dff_B_lJZSXHvj7_1(.din(w_dff_B_At1YA5Vh4_1),.dout(w_dff_B_lJZSXHvj7_1),.clk(gclk));
	jdff dff_B_m1rdW9ar1_1(.din(w_dff_B_lJZSXHvj7_1),.dout(w_dff_B_m1rdW9ar1_1),.clk(gclk));
	jdff dff_B_BQ2EQVOl9_1(.din(w_dff_B_m1rdW9ar1_1),.dout(w_dff_B_BQ2EQVOl9_1),.clk(gclk));
	jdff dff_B_1iNS7Nap6_0(.din(n839),.dout(w_dff_B_1iNS7Nap6_0),.clk(gclk));
	jdff dff_B_eMTh1SQH4_0(.din(w_dff_B_1iNS7Nap6_0),.dout(w_dff_B_eMTh1SQH4_0),.clk(gclk));
	jdff dff_B_SXzXfOxQ5_0(.din(w_dff_B_eMTh1SQH4_0),.dout(w_dff_B_SXzXfOxQ5_0),.clk(gclk));
	jdff dff_B_LDLs90Uk8_0(.din(w_dff_B_SXzXfOxQ5_0),.dout(w_dff_B_LDLs90Uk8_0),.clk(gclk));
	jdff dff_B_heqfmxww4_0(.din(w_dff_B_LDLs90Uk8_0),.dout(w_dff_B_heqfmxww4_0),.clk(gclk));
	jdff dff_B_G225qpP34_0(.din(w_dff_B_heqfmxww4_0),.dout(w_dff_B_G225qpP34_0),.clk(gclk));
	jdff dff_B_Sq3v5Xdh4_1(.din(n360),.dout(w_dff_B_Sq3v5Xdh4_1),.clk(gclk));
	jdff dff_A_9JjDmRhG0_0(.dout(w_n749_11[0]),.din(w_dff_A_9JjDmRhG0_0),.clk(gclk));
	jdff dff_A_7TidQJ6G5_1(.dout(w_n749_11[1]),.din(w_dff_A_7TidQJ6G5_1),.clk(gclk));
	jdff dff_A_Q62aijYp6_0(.dout(w_n749_3[0]),.din(w_dff_A_Q62aijYp6_0),.clk(gclk));
	jdff dff_A_QcqzsMkw0_2(.dout(w_n749_3[2]),.din(w_dff_A_QcqzsMkw0_2),.clk(gclk));
	jdff dff_A_QegbFgMH0_1(.dout(w_G4092_8[1]),.din(w_dff_A_QegbFgMH0_1),.clk(gclk));
	jdff dff_A_fI6T211y3_2(.dout(w_G4092_8[2]),.din(w_dff_A_fI6T211y3_2),.clk(gclk));
	jdff dff_A_ORZgCVlI8_0(.dout(w_n836_0[0]),.din(w_dff_A_ORZgCVlI8_0),.clk(gclk));
	jdff dff_A_7suQ0XYU3_0(.dout(w_dff_A_ORZgCVlI8_0),.din(w_dff_A_7suQ0XYU3_0),.clk(gclk));
	jdff dff_A_hAkS5YAw9_0(.dout(w_dff_A_7suQ0XYU3_0),.din(w_dff_A_hAkS5YAw9_0),.clk(gclk));
	jdff dff_A_d6GDjhyS9_0(.dout(w_dff_A_hAkS5YAw9_0),.din(w_dff_A_d6GDjhyS9_0),.clk(gclk));
	jdff dff_A_97sd9oJa1_0(.dout(w_dff_A_d6GDjhyS9_0),.din(w_dff_A_97sd9oJa1_0),.clk(gclk));
	jdff dff_A_7ThD62w13_0(.dout(w_dff_A_97sd9oJa1_0),.din(w_dff_A_7ThD62w13_0),.clk(gclk));
	jdff dff_A_V7JhJi4I3_0(.dout(w_dff_A_7ThD62w13_0),.din(w_dff_A_V7JhJi4I3_0),.clk(gclk));
	jdff dff_A_crg4mZyX4_1(.dout(w_n753_0[1]),.din(w_dff_A_crg4mZyX4_1),.clk(gclk));
	jdff dff_A_Xx2je7Ng9_1(.dout(w_dff_A_crg4mZyX4_1),.din(w_dff_A_Xx2je7Ng9_1),.clk(gclk));
	jdff dff_A_segWPjME5_2(.dout(w_n753_0[2]),.din(w_dff_A_segWPjME5_2),.clk(gclk));
	jdff dff_A_yIPwBlnh7_2(.dout(w_dff_A_segWPjME5_2),.din(w_dff_A_yIPwBlnh7_2),.clk(gclk));
	jdff dff_A_dJn9XU4r0_2(.dout(w_dff_A_yIPwBlnh7_2),.din(w_dff_A_dJn9XU4r0_2),.clk(gclk));
	jdff dff_A_J9WMtu723_2(.dout(w_dff_A_dJn9XU4r0_2),.din(w_dff_A_J9WMtu723_2),.clk(gclk));
	jdff dff_A_eCToI8218_2(.dout(w_dff_A_J9WMtu723_2),.din(w_dff_A_eCToI8218_2),.clk(gclk));
	jdff dff_B_gMSfxgK16_3(.din(n753),.dout(w_dff_B_gMSfxgK16_3),.clk(gclk));
	jdff dff_B_KcNeIWmv8_3(.din(w_dff_B_gMSfxgK16_3),.dout(w_dff_B_KcNeIWmv8_3),.clk(gclk));
	jdff dff_A_1TDZkw5D4_0(.dout(w_G4091_4[0]),.din(w_dff_A_1TDZkw5D4_0),.clk(gclk));
	jdff dff_A_UmKYnHNg0_0(.dout(w_dff_A_1TDZkw5D4_0),.din(w_dff_A_UmKYnHNg0_0),.clk(gclk));
	jdff dff_A_AlWs86Wg8_0(.dout(w_dff_A_UmKYnHNg0_0),.din(w_dff_A_AlWs86Wg8_0),.clk(gclk));
	jdff dff_A_vWLEkGRQ2_0(.dout(w_dff_A_AlWs86Wg8_0),.din(w_dff_A_vWLEkGRQ2_0),.clk(gclk));
	jdff dff_A_dzVduUWR0_2(.dout(w_G4091_4[2]),.din(w_dff_A_dzVduUWR0_2),.clk(gclk));
	jdff dff_A_PWGx2d8f6_2(.dout(w_dff_A_dzVduUWR0_2),.din(w_dff_A_PWGx2d8f6_2),.clk(gclk));
	jdff dff_A_a58CEpQU8_2(.dout(w_dff_A_PWGx2d8f6_2),.din(w_dff_A_a58CEpQU8_2),.clk(gclk));
	jdff dff_B_mjLra52h0_1(.din(G130),.dout(w_dff_B_mjLra52h0_1),.clk(gclk));
	jdff dff_B_4LVBH2It6_1(.din(w_dff_B_mjLra52h0_1),.dout(w_dff_B_4LVBH2It6_1),.clk(gclk));
	jdff dff_B_SJTCTUpE8_1(.din(n1173),.dout(w_dff_B_SJTCTUpE8_1),.clk(gclk));
	jdff dff_B_0pq8b4099_1(.din(w_dff_B_SJTCTUpE8_1),.dout(w_dff_B_0pq8b4099_1),.clk(gclk));
	jdff dff_B_wP0WAYa06_1(.din(w_dff_B_0pq8b4099_1),.dout(w_dff_B_wP0WAYa06_1),.clk(gclk));
	jdff dff_B_FfW8U1v00_1(.din(w_dff_B_wP0WAYa06_1),.dout(w_dff_B_FfW8U1v00_1),.clk(gclk));
	jdff dff_B_dw0eGgNd5_1(.din(w_dff_B_FfW8U1v00_1),.dout(w_dff_B_dw0eGgNd5_1),.clk(gclk));
	jdff dff_B_BDi1Z0Wg1_1(.din(w_dff_B_dw0eGgNd5_1),.dout(w_dff_B_BDi1Z0Wg1_1),.clk(gclk));
	jdff dff_B_NK9pg6376_1(.din(w_dff_B_BDi1Z0Wg1_1),.dout(w_dff_B_NK9pg6376_1),.clk(gclk));
	jdff dff_B_gxIe1wTu2_1(.din(w_dff_B_NK9pg6376_1),.dout(w_dff_B_gxIe1wTu2_1),.clk(gclk));
	jdff dff_B_jhc8k3IX3_1(.din(w_dff_B_gxIe1wTu2_1),.dout(w_dff_B_jhc8k3IX3_1),.clk(gclk));
	jdff dff_B_yS83qBjv9_1(.din(w_dff_B_jhc8k3IX3_1),.dout(w_dff_B_yS83qBjv9_1),.clk(gclk));
	jdff dff_B_JIjnueRV8_1(.din(w_dff_B_yS83qBjv9_1),.dout(w_dff_B_JIjnueRV8_1),.clk(gclk));
	jdff dff_B_262O5ZM97_1(.din(w_dff_B_JIjnueRV8_1),.dout(w_dff_B_262O5ZM97_1),.clk(gclk));
	jdff dff_B_h34gSi9m2_1(.din(w_dff_B_262O5ZM97_1),.dout(w_dff_B_h34gSi9m2_1),.clk(gclk));
	jdff dff_B_wujcZsIp8_1(.din(w_dff_B_h34gSi9m2_1),.dout(w_dff_B_wujcZsIp8_1),.clk(gclk));
	jdff dff_B_rzkQElNl3_1(.din(w_dff_B_wujcZsIp8_1),.dout(w_dff_B_rzkQElNl3_1),.clk(gclk));
	jdff dff_B_YehUqUFZ2_1(.din(w_dff_B_rzkQElNl3_1),.dout(w_dff_B_YehUqUFZ2_1),.clk(gclk));
	jdff dff_B_yPIn38pH5_1(.din(w_dff_B_YehUqUFZ2_1),.dout(w_dff_B_yPIn38pH5_1),.clk(gclk));
	jdff dff_B_IR1js6PY9_1(.din(w_dff_B_yPIn38pH5_1),.dout(w_dff_B_IR1js6PY9_1),.clk(gclk));
	jdff dff_B_p01T7xu26_1(.din(n1182),.dout(w_dff_B_p01T7xu26_1),.clk(gclk));
	jdff dff_B_x2B1v9ul5_1(.din(w_dff_B_p01T7xu26_1),.dout(w_dff_B_x2B1v9ul5_1),.clk(gclk));
	jdff dff_B_9XDQ9MuK2_1(.din(w_dff_B_x2B1v9ul5_1),.dout(w_dff_B_9XDQ9MuK2_1),.clk(gclk));
	jdff dff_B_6rxE4lJ27_1(.din(w_dff_B_9XDQ9MuK2_1),.dout(w_dff_B_6rxE4lJ27_1),.clk(gclk));
	jdff dff_B_S5HSk2m91_1(.din(w_dff_B_6rxE4lJ27_1),.dout(w_dff_B_S5HSk2m91_1),.clk(gclk));
	jdff dff_B_fBrT7Hht7_1(.din(w_dff_B_S5HSk2m91_1),.dout(w_dff_B_fBrT7Hht7_1),.clk(gclk));
	jdff dff_B_LbGTneuH2_1(.din(w_dff_B_fBrT7Hht7_1),.dout(w_dff_B_LbGTneuH2_1),.clk(gclk));
	jdff dff_B_TSoGnU751_1(.din(w_dff_B_LbGTneuH2_1),.dout(w_dff_B_TSoGnU751_1),.clk(gclk));
	jdff dff_B_giGWtHgu2_1(.din(w_dff_B_TSoGnU751_1),.dout(w_dff_B_giGWtHgu2_1),.clk(gclk));
	jdff dff_B_AcWpHut54_1(.din(w_dff_B_giGWtHgu2_1),.dout(w_dff_B_AcWpHut54_1),.clk(gclk));
	jdff dff_B_Y2q2okYk1_0(.din(n1185),.dout(w_dff_B_Y2q2okYk1_0),.clk(gclk));
	jdff dff_B_pma8W6UL3_0(.din(w_dff_B_Y2q2okYk1_0),.dout(w_dff_B_pma8W6UL3_0),.clk(gclk));
	jdff dff_B_jifYEoLa5_0(.din(w_dff_B_pma8W6UL3_0),.dout(w_dff_B_jifYEoLa5_0),.clk(gclk));
	jdff dff_B_ZEnctCti8_0(.din(w_dff_B_jifYEoLa5_0),.dout(w_dff_B_ZEnctCti8_0),.clk(gclk));
	jdff dff_B_EmH8pxP01_0(.din(w_dff_B_ZEnctCti8_0),.dout(w_dff_B_EmH8pxP01_0),.clk(gclk));
	jdff dff_B_Naal926N0_0(.din(w_dff_B_EmH8pxP01_0),.dout(w_dff_B_Naal926N0_0),.clk(gclk));
	jdff dff_B_q67KMKMI6_0(.din(w_dff_B_Naal926N0_0),.dout(w_dff_B_q67KMKMI6_0),.clk(gclk));
	jdff dff_B_Gmtzc4x55_0(.din(w_dff_B_q67KMKMI6_0),.dout(w_dff_B_Gmtzc4x55_0),.clk(gclk));
	jdff dff_B_gWjX512N1_0(.din(w_dff_B_Gmtzc4x55_0),.dout(w_dff_B_gWjX512N1_0),.clk(gclk));
	jdff dff_B_9K9OXY3N2_0(.din(w_dff_B_gWjX512N1_0),.dout(w_dff_B_9K9OXY3N2_0),.clk(gclk));
	jdff dff_B_HwYRXSb17_0(.din(w_dff_B_9K9OXY3N2_0),.dout(w_dff_B_HwYRXSb17_0),.clk(gclk));
	jdff dff_B_8KOJ0rAh4_0(.din(w_dff_B_HwYRXSb17_0),.dout(w_dff_B_8KOJ0rAh4_0),.clk(gclk));
	jdff dff_B_aGH9xiGJ4_0(.din(w_dff_B_8KOJ0rAh4_0),.dout(w_dff_B_aGH9xiGJ4_0),.clk(gclk));
	jdff dff_B_oL3F66b33_0(.din(w_dff_B_aGH9xiGJ4_0),.dout(w_dff_B_oL3F66b33_0),.clk(gclk));
	jdff dff_B_FuoDS0bO8_0(.din(w_dff_B_oL3F66b33_0),.dout(w_dff_B_FuoDS0bO8_0),.clk(gclk));
	jdff dff_B_REvoa9Uk5_0(.din(w_dff_B_FuoDS0bO8_0),.dout(w_dff_B_REvoa9Uk5_0),.clk(gclk));
	jdff dff_B_t6pHtrQy5_1(.din(n1175),.dout(w_dff_B_t6pHtrQy5_1),.clk(gclk));
	jdff dff_B_dDzzxKxE0_1(.din(w_dff_B_t6pHtrQy5_1),.dout(w_dff_B_dDzzxKxE0_1),.clk(gclk));
	jdff dff_B_eTcQlCR77_1(.din(w_dff_B_dDzzxKxE0_1),.dout(w_dff_B_eTcQlCR77_1),.clk(gclk));
	jdff dff_B_Txjh1bF79_1(.din(n1176),.dout(w_dff_B_Txjh1bF79_1),.clk(gclk));
	jdff dff_B_EEK85wo98_1(.din(w_dff_B_Txjh1bF79_1),.dout(w_dff_B_EEK85wo98_1),.clk(gclk));
	jdff dff_B_e6rApPUh7_1(.din(w_dff_B_EEK85wo98_1),.dout(w_dff_B_e6rApPUh7_1),.clk(gclk));
	jdff dff_B_0OOP1XMK4_1(.din(w_dff_B_e6rApPUh7_1),.dout(w_dff_B_0OOP1XMK4_1),.clk(gclk));
	jdff dff_B_utxupP6v0_1(.din(w_dff_B_0OOP1XMK4_1),.dout(w_dff_B_utxupP6v0_1),.clk(gclk));
	jdff dff_B_fkywhnmy6_1(.din(w_dff_B_utxupP6v0_1),.dout(w_dff_B_fkywhnmy6_1),.clk(gclk));
	jdff dff_A_qAfsH6ps1_0(.dout(w_n1177_0[0]),.din(w_dff_A_qAfsH6ps1_0),.clk(gclk));
	jdff dff_A_ka0Af7gB1_0(.dout(w_dff_A_qAfsH6ps1_0),.din(w_dff_A_ka0Af7gB1_0),.clk(gclk));
	jdff dff_A_Y7VtoUEM8_0(.dout(w_dff_A_ka0Af7gB1_0),.din(w_dff_A_Y7VtoUEM8_0),.clk(gclk));
	jdff dff_A_vXaZmONx2_0(.dout(w_dff_A_Y7VtoUEM8_0),.din(w_dff_A_vXaZmONx2_0),.clk(gclk));
	jdff dff_A_3u8AhDZ50_0(.dout(w_dff_A_vXaZmONx2_0),.din(w_dff_A_3u8AhDZ50_0),.clk(gclk));
	jdff dff_A_CBmTJGOR5_0(.dout(w_dff_A_3u8AhDZ50_0),.din(w_dff_A_CBmTJGOR5_0),.clk(gclk));
	jdff dff_A_2n1SrRKC7_0(.dout(w_dff_A_CBmTJGOR5_0),.din(w_dff_A_2n1SrRKC7_0),.clk(gclk));
	jdff dff_A_FdbRZcal4_0(.dout(w_dff_A_2n1SrRKC7_0),.din(w_dff_A_FdbRZcal4_0),.clk(gclk));
	jdff dff_A_XpKbW4934_0(.dout(w_dff_A_FdbRZcal4_0),.din(w_dff_A_XpKbW4934_0),.clk(gclk));
	jdff dff_A_WAbi9woj3_0(.dout(w_dff_A_XpKbW4934_0),.din(w_dff_A_WAbi9woj3_0),.clk(gclk));
	jdff dff_A_q0KUU9WO9_0(.dout(w_dff_A_WAbi9woj3_0),.din(w_dff_A_q0KUU9WO9_0),.clk(gclk));
	jdff dff_B_1JrkY8Dv8_2(.din(n1177),.dout(w_dff_B_1JrkY8Dv8_2),.clk(gclk));
	jdff dff_B_Ozu4KnEC0_2(.din(w_dff_B_1JrkY8Dv8_2),.dout(w_dff_B_Ozu4KnEC0_2),.clk(gclk));
	jdff dff_B_llg6wm2I2_2(.din(w_dff_B_Ozu4KnEC0_2),.dout(w_dff_B_llg6wm2I2_2),.clk(gclk));
	jdff dff_B_nGukN8y83_2(.din(w_dff_B_llg6wm2I2_2),.dout(w_dff_B_nGukN8y83_2),.clk(gclk));
	jdff dff_B_eBuerXZk9_2(.din(w_dff_B_nGukN8y83_2),.dout(w_dff_B_eBuerXZk9_2),.clk(gclk));
	jdff dff_A_yY3htEE00_0(.dout(w_G3717_0[0]),.din(w_dff_A_yY3htEE00_0),.clk(gclk));
	jdff dff_A_Spe8grpu6_1(.dout(w_n428_1[1]),.din(w_dff_A_Spe8grpu6_1),.clk(gclk));
	jdff dff_A_ce82iF9C0_2(.dout(w_G3724_0[2]),.din(w_dff_A_ce82iF9C0_2),.clk(gclk));
	jdff dff_A_bqmsRlfN6_2(.dout(w_dff_A_ce82iF9C0_2),.din(w_dff_A_bqmsRlfN6_2),.clk(gclk));
	jdff dff_A_iymLysLC7_2(.dout(w_dff_A_bqmsRlfN6_2),.din(w_dff_A_iymLysLC7_2),.clk(gclk));
	jdff dff_A_nRGnI5Q08_2(.dout(w_dff_A_iymLysLC7_2),.din(w_dff_A_nRGnI5Q08_2),.clk(gclk));
	jdff dff_A_faYPsANX9_0(.dout(w_n1179_0[0]),.din(w_dff_A_faYPsANX9_0),.clk(gclk));
	jdff dff_A_IL6xpjDa7_0(.dout(w_dff_A_faYPsANX9_0),.din(w_dff_A_IL6xpjDa7_0),.clk(gclk));
	jdff dff_A_Q6I6sg426_0(.dout(w_dff_A_IL6xpjDa7_0),.din(w_dff_A_Q6I6sg426_0),.clk(gclk));
	jdff dff_A_2ESL2CEo6_0(.dout(w_dff_A_Q6I6sg426_0),.din(w_dff_A_2ESL2CEo6_0),.clk(gclk));
	jdff dff_A_ZDO7B8j88_0(.dout(w_dff_A_2ESL2CEo6_0),.din(w_dff_A_ZDO7B8j88_0),.clk(gclk));
	jdff dff_A_zyAtjveW0_0(.dout(w_dff_A_ZDO7B8j88_0),.din(w_dff_A_zyAtjveW0_0),.clk(gclk));
	jdff dff_A_VihzxTqh9_0(.dout(w_dff_A_zyAtjveW0_0),.din(w_dff_A_VihzxTqh9_0),.clk(gclk));
	jdff dff_A_l1TPZ3Kj2_0(.dout(w_dff_A_VihzxTqh9_0),.din(w_dff_A_l1TPZ3Kj2_0),.clk(gclk));
	jdff dff_A_zOHvRT210_0(.dout(w_dff_A_l1TPZ3Kj2_0),.din(w_dff_A_zOHvRT210_0),.clk(gclk));
	jdff dff_A_kjwlrNqP9_0(.dout(w_dff_A_zOHvRT210_0),.din(w_dff_A_kjwlrNqP9_0),.clk(gclk));
	jdff dff_A_HFFMZKXC4_0(.dout(w_dff_A_kjwlrNqP9_0),.din(w_dff_A_HFFMZKXC4_0),.clk(gclk));
	jdff dff_B_2ODW0byy4_1(.din(G132),.dout(w_dff_B_2ODW0byy4_1),.clk(gclk));
	jdff dff_B_bR5wdcvE0_1(.din(w_dff_B_2ODW0byy4_1),.dout(w_dff_B_bR5wdcvE0_1),.clk(gclk));
	jdff dff_B_YCh1T0KM1_1(.din(w_dff_B_bR5wdcvE0_1),.dout(w_dff_B_YCh1T0KM1_1),.clk(gclk));
	jdff dff_B_WLeseU1z1_1(.din(w_dff_B_YCh1T0KM1_1),.dout(w_dff_B_WLeseU1z1_1),.clk(gclk));
	jdff dff_B_GBcMuDia6_1(.din(n1223),.dout(w_dff_B_GBcMuDia6_1),.clk(gclk));
	jdff dff_B_9WsjWPI97_0(.din(n1227),.dout(w_dff_B_9WsjWPI97_0),.clk(gclk));
	jdff dff_B_PoXP9G9H8_0(.din(w_dff_B_9WsjWPI97_0),.dout(w_dff_B_PoXP9G9H8_0),.clk(gclk));
	jdff dff_B_LH6zC8nH4_0(.din(w_dff_B_PoXP9G9H8_0),.dout(w_dff_B_LH6zC8nH4_0),.clk(gclk));
	jdff dff_B_N5kgZ4q98_0(.din(w_dff_B_LH6zC8nH4_0),.dout(w_dff_B_N5kgZ4q98_0),.clk(gclk));
	jdff dff_B_tam88bC02_0(.din(n1226),.dout(w_dff_B_tam88bC02_0),.clk(gclk));
	jdff dff_A_JmBuoIrZ9_0(.dout(w_G559_0[0]),.din(w_dff_A_JmBuoIrZ9_0),.clk(gclk));
	jdff dff_A_FtQ5RHRX1_0(.dout(w_dff_A_JmBuoIrZ9_0),.din(w_dff_A_FtQ5RHRX1_0),.clk(gclk));
	jdff dff_B_lwgdiKd39_0(.din(n668),.dout(w_dff_B_lwgdiKd39_0),.clk(gclk));
	jdff dff_B_Qa0kXc944_1(.din(n663),.dout(w_dff_B_Qa0kXc944_1),.clk(gclk));
	jdff dff_B_gv7JNX2u5_1(.din(n916),.dout(w_dff_B_gv7JNX2u5_1),.clk(gclk));
	jdff dff_B_ArBKaFRb0_1(.din(n917),.dout(w_dff_B_ArBKaFRb0_1),.clk(gclk));
	jdff dff_B_GgwDVmIk2_0(.din(n915),.dout(w_dff_B_GgwDVmIk2_0),.clk(gclk));
	jdff dff_B_xLQe94xi2_1(.din(n913),.dout(w_dff_B_xLQe94xi2_1),.clk(gclk));
	jdff dff_B_Y91lCFsy5_0(.din(G372),.dout(w_dff_B_Y91lCFsy5_0),.clk(gclk));
	jdff dff_B_UpMQVbjd6_1(.din(n909),.dout(w_dff_B_UpMQVbjd6_1),.clk(gclk));
	jdff dff_B_jaZ47cMA7_1(.din(n907),.dout(w_dff_B_jaZ47cMA7_1),.clk(gclk));
	jdff dff_B_7xINs6mG3_1(.din(w_dff_B_jaZ47cMA7_1),.dout(w_dff_B_7xINs6mG3_1),.clk(gclk));
	jdff dff_B_Y2yoSY4w4_0(.din(n1222),.dout(w_dff_B_Y2yoSY4w4_0),.clk(gclk));
	jdff dff_B_jOxmupOZ6_0(.din(w_dff_B_Y2yoSY4w4_0),.dout(w_dff_B_jOxmupOZ6_0),.clk(gclk));
	jdff dff_B_yrPwA8uG8_0(.din(w_dff_B_jOxmupOZ6_0),.dout(w_dff_B_yrPwA8uG8_0),.clk(gclk));
	jdff dff_B_kSKAt8eF0_0(.din(n678),.dout(w_dff_B_kSKAt8eF0_0),.clk(gclk));
	jdff dff_B_HIzuN37p7_1(.din(n672),.dout(w_dff_B_HIzuN37p7_1),.clk(gclk));
	jdff dff_A_J483ghBZ3_0(.dout(w_G245_0[0]),.din(w_dff_A_J483ghBZ3_0),.clk(gclk));
	jdff dff_A_R1I8Dhts8_0(.dout(w_dff_A_J483ghBZ3_0),.din(w_dff_A_R1I8Dhts8_0),.clk(gclk));
	jdff dff_A_bXDUOtni8_0(.dout(w_dff_A_R1I8Dhts8_0),.din(w_dff_A_bXDUOtni8_0),.clk(gclk));
	jdff dff_A_lTOzkCx56_0(.dout(w_dff_A_bXDUOtni8_0),.din(w_dff_A_lTOzkCx56_0),.clk(gclk));
	jdff dff_B_Lkz0kzL29_1(.din(n926),.dout(w_dff_B_Lkz0kzL29_1),.clk(gclk));
	jdff dff_B_FTZIdq6L0_1(.din(n930),.dout(w_dff_B_FTZIdq6L0_1),.clk(gclk));
	jdff dff_B_WMbiIHUO3_1(.din(w_dff_B_FTZIdq6L0_1),.dout(w_dff_B_WMbiIHUO3_1),.clk(gclk));
	jdff dff_B_1GSiAlF65_1(.din(n927),.dout(w_dff_B_1GSiAlF65_1),.clk(gclk));
	jdff dff_B_KzVdmX5f1_1(.din(G292),.dout(w_dff_B_KzVdmX5f1_1),.clk(gclk));
	jdff dff_B_Eh8xcU5w1_1(.din(n1263),.dout(w_dff_B_Eh8xcU5w1_1),.clk(gclk));
	jdff dff_B_R6OPvu1m6_1(.din(w_dff_B_Eh8xcU5w1_1),.dout(w_dff_B_R6OPvu1m6_1),.clk(gclk));
	jdff dff_B_tO5YvwMX9_1(.din(w_dff_B_R6OPvu1m6_1),.dout(w_dff_B_tO5YvwMX9_1),.clk(gclk));
	jdff dff_B_xTqVdMq19_1(.din(w_dff_B_tO5YvwMX9_1),.dout(w_dff_B_xTqVdMq19_1),.clk(gclk));
	jdff dff_B_Yn23Ap934_1(.din(w_dff_B_xTqVdMq19_1),.dout(w_dff_B_Yn23Ap934_1),.clk(gclk));
	jdff dff_B_OUA70wuN8_1(.din(w_dff_B_Yn23Ap934_1),.dout(w_dff_B_OUA70wuN8_1),.clk(gclk));
	jdff dff_B_CHoghGGr2_1(.din(w_dff_B_OUA70wuN8_1),.dout(w_dff_B_CHoghGGr2_1),.clk(gclk));
	jdff dff_B_sRwG79PK9_1(.din(w_dff_B_CHoghGGr2_1),.dout(w_dff_B_sRwG79PK9_1),.clk(gclk));
	jdff dff_B_d0vPN1jU2_1(.din(w_dff_B_sRwG79PK9_1),.dout(w_dff_B_d0vPN1jU2_1),.clk(gclk));
	jdff dff_B_XgTP2XRT7_1(.din(w_dff_B_d0vPN1jU2_1),.dout(w_dff_B_XgTP2XRT7_1),.clk(gclk));
	jdff dff_B_xF71wDdE2_1(.din(w_dff_B_XgTP2XRT7_1),.dout(w_dff_B_xF71wDdE2_1),.clk(gclk));
	jdff dff_B_vUmjxWLO5_1(.din(w_dff_B_xF71wDdE2_1),.dout(w_dff_B_vUmjxWLO5_1),.clk(gclk));
	jdff dff_B_Qv13RY871_1(.din(w_dff_B_vUmjxWLO5_1),.dout(w_dff_B_Qv13RY871_1),.clk(gclk));
	jdff dff_B_WLoJdSsh8_1(.din(w_dff_B_Qv13RY871_1),.dout(w_dff_B_WLoJdSsh8_1),.clk(gclk));
	jdff dff_B_blNbS6wX1_1(.din(w_dff_B_WLoJdSsh8_1),.dout(w_dff_B_blNbS6wX1_1),.clk(gclk));
	jdff dff_B_Rh31UQkH5_1(.din(w_dff_B_blNbS6wX1_1),.dout(w_dff_B_Rh31UQkH5_1),.clk(gclk));
	jdff dff_B_TT1moR132_1(.din(w_dff_B_Rh31UQkH5_1),.dout(w_dff_B_TT1moR132_1),.clk(gclk));
	jdff dff_B_Ah0S6DeG2_1(.din(w_dff_B_TT1moR132_1),.dout(w_dff_B_Ah0S6DeG2_1),.clk(gclk));
	jdff dff_B_awItk95I5_1(.din(w_dff_B_Ah0S6DeG2_1),.dout(w_dff_B_awItk95I5_1),.clk(gclk));
	jdff dff_B_LVHBRYbN7_1(.din(n1260),.dout(w_dff_B_LVHBRYbN7_1),.clk(gclk));
	jdff dff_B_RL3xREXt5_1(.din(w_dff_B_LVHBRYbN7_1),.dout(w_dff_B_RL3xREXt5_1),.clk(gclk));
	jdff dff_A_bRwySmv44_2(.dout(w_n852_6[2]),.din(w_dff_A_bRwySmv44_2),.clk(gclk));
	jdff dff_A_hIMjxelj8_2(.dout(w_dff_A_bRwySmv44_2),.din(w_dff_A_hIMjxelj8_2),.clk(gclk));
	jdff dff_A_0YCsWJI95_2(.dout(w_dff_A_hIMjxelj8_2),.din(w_dff_A_0YCsWJI95_2),.clk(gclk));
	jdff dff_A_NdvFqruk6_2(.dout(w_dff_A_0YCsWJI95_2),.din(w_dff_A_NdvFqruk6_2),.clk(gclk));
	jdff dff_A_vBqxePfa1_2(.dout(w_dff_A_NdvFqruk6_2),.din(w_dff_A_vBqxePfa1_2),.clk(gclk));
	jdff dff_A_klTK2TIY7_2(.dout(w_dff_A_vBqxePfa1_2),.din(w_dff_A_klTK2TIY7_2),.clk(gclk));
	jdff dff_A_8gqaPvZ35_2(.dout(w_dff_A_klTK2TIY7_2),.din(w_dff_A_8gqaPvZ35_2),.clk(gclk));
	jdff dff_A_T2fUFLh32_2(.dout(w_dff_A_8gqaPvZ35_2),.din(w_dff_A_T2fUFLh32_2),.clk(gclk));
	jdff dff_A_eIaYIMDb1_2(.dout(w_dff_A_T2fUFLh32_2),.din(w_dff_A_eIaYIMDb1_2),.clk(gclk));
	jdff dff_A_R2KmGRb39_2(.dout(w_dff_A_eIaYIMDb1_2),.din(w_dff_A_R2KmGRb39_2),.clk(gclk));
	jdff dff_A_GbTFOAwC9_2(.dout(w_dff_A_R2KmGRb39_2),.din(w_dff_A_GbTFOAwC9_2),.clk(gclk));
	jdff dff_A_Jn6agjht7_2(.dout(w_G4089_6[2]),.din(w_dff_A_Jn6agjht7_2),.clk(gclk));
	jdff dff_A_zK74rVjF6_2(.dout(w_dff_A_Jn6agjht7_2),.din(w_dff_A_zK74rVjF6_2),.clk(gclk));
	jdff dff_A_WoT2ruqa0_2(.dout(w_dff_A_zK74rVjF6_2),.din(w_dff_A_WoT2ruqa0_2),.clk(gclk));
	jdff dff_A_fgX5Exue9_2(.dout(w_dff_A_WoT2ruqa0_2),.din(w_dff_A_fgX5Exue9_2),.clk(gclk));
	jdff dff_A_QtfeuDtX3_2(.dout(w_dff_A_fgX5Exue9_2),.din(w_dff_A_QtfeuDtX3_2),.clk(gclk));
	jdff dff_A_NunGVhI32_2(.dout(w_dff_A_QtfeuDtX3_2),.din(w_dff_A_NunGVhI32_2),.clk(gclk));
	jdff dff_A_ZPlxwMdM3_2(.dout(w_dff_A_NunGVhI32_2),.din(w_dff_A_ZPlxwMdM3_2),.clk(gclk));
	jdff dff_A_IMnj1xPy9_2(.dout(w_dff_A_ZPlxwMdM3_2),.din(w_dff_A_IMnj1xPy9_2),.clk(gclk));
	jdff dff_A_5zXiPppJ4_2(.dout(w_dff_A_IMnj1xPy9_2),.din(w_dff_A_5zXiPppJ4_2),.clk(gclk));
	jdff dff_A_5VTLUQNs7_2(.dout(w_dff_A_5zXiPppJ4_2),.din(w_dff_A_5VTLUQNs7_2),.clk(gclk));
	jdff dff_A_6zJ0XKoK5_2(.dout(w_dff_A_5VTLUQNs7_2),.din(w_dff_A_6zJ0XKoK5_2),.clk(gclk));
	jdff dff_A_NWM5yy8d4_2(.dout(w_dff_A_6zJ0XKoK5_2),.din(w_dff_A_NWM5yy8d4_2),.clk(gclk));
	jdff dff_A_BePHHIG12_2(.dout(w_dff_A_NWM5yy8d4_2),.din(w_dff_A_BePHHIG12_2),.clk(gclk));
	jdff dff_A_SuyHfsP33_2(.dout(w_dff_A_BePHHIG12_2),.din(w_dff_A_SuyHfsP33_2),.clk(gclk));
	jdff dff_B_WRpIyDKr5_0(.din(n1276),.dout(w_dff_B_WRpIyDKr5_0),.clk(gclk));
	jdff dff_B_G6NOgQou0_0(.din(w_dff_B_WRpIyDKr5_0),.dout(w_dff_B_G6NOgQou0_0),.clk(gclk));
	jdff dff_B_AsRt94t66_0(.din(w_dff_B_G6NOgQou0_0),.dout(w_dff_B_AsRt94t66_0),.clk(gclk));
	jdff dff_B_xa0r5KoB9_0(.din(w_dff_B_AsRt94t66_0),.dout(w_dff_B_xa0r5KoB9_0),.clk(gclk));
	jdff dff_B_VOw4BDys5_0(.din(w_dff_B_xa0r5KoB9_0),.dout(w_dff_B_VOw4BDys5_0),.clk(gclk));
	jdff dff_B_9tOouuU77_0(.din(w_dff_B_VOw4BDys5_0),.dout(w_dff_B_9tOouuU77_0),.clk(gclk));
	jdff dff_B_GIuNXjbb3_0(.din(w_dff_B_9tOouuU77_0),.dout(w_dff_B_GIuNXjbb3_0),.clk(gclk));
	jdff dff_B_xoYDG25r2_0(.din(w_dff_B_GIuNXjbb3_0),.dout(w_dff_B_xoYDG25r2_0),.clk(gclk));
	jdff dff_B_3MNhwztg4_0(.din(w_dff_B_xoYDG25r2_0),.dout(w_dff_B_3MNhwztg4_0),.clk(gclk));
	jdff dff_B_tooZ1f2L3_0(.din(w_dff_B_3MNhwztg4_0),.dout(w_dff_B_tooZ1f2L3_0),.clk(gclk));
	jdff dff_B_97cH0skD7_0(.din(w_dff_B_tooZ1f2L3_0),.dout(w_dff_B_97cH0skD7_0),.clk(gclk));
	jdff dff_B_VZ8CXkyb1_0(.din(w_dff_B_97cH0skD7_0),.dout(w_dff_B_VZ8CXkyb1_0),.clk(gclk));
	jdff dff_B_VFOFqvPb3_0(.din(w_dff_B_VZ8CXkyb1_0),.dout(w_dff_B_VFOFqvPb3_0),.clk(gclk));
	jdff dff_B_yYWLHLHx1_0(.din(w_dff_B_VFOFqvPb3_0),.dout(w_dff_B_yYWLHLHx1_0),.clk(gclk));
	jdff dff_B_BXeoeUfm2_0(.din(w_dff_B_yYWLHLHx1_0),.dout(w_dff_B_BXeoeUfm2_0),.clk(gclk));
	jdff dff_B_G9lWqzGc2_0(.din(w_dff_B_BXeoeUfm2_0),.dout(w_dff_B_G9lWqzGc2_0),.clk(gclk));
	jdff dff_B_3VyOr7uT0_0(.din(w_dff_B_G9lWqzGc2_0),.dout(w_dff_B_3VyOr7uT0_0),.clk(gclk));
	jdff dff_B_Pdrz4BLb9_0(.din(w_dff_B_3VyOr7uT0_0),.dout(w_dff_B_Pdrz4BLb9_0),.clk(gclk));
	jdff dff_B_oiuRAOfW1_0(.din(w_dff_B_Pdrz4BLb9_0),.dout(w_dff_B_oiuRAOfW1_0),.clk(gclk));
	jdff dff_B_oDyragN69_0(.din(w_dff_B_oiuRAOfW1_0),.dout(w_dff_B_oDyragN69_0),.clk(gclk));
	jdff dff_B_VNDVWmfp6_0(.din(w_dff_B_oDyragN69_0),.dout(w_dff_B_VNDVWmfp6_0),.clk(gclk));
	jdff dff_B_ysMN1GsA7_2(.din(G106),.dout(w_dff_B_ysMN1GsA7_2),.clk(gclk));
	jdff dff_B_kPe973K11_1(.din(n1269),.dout(w_dff_B_kPe973K11_1),.clk(gclk));
	jdff dff_B_gFIIPHp96_1(.din(w_dff_B_kPe973K11_1),.dout(w_dff_B_gFIIPHp96_1),.clk(gclk));
	jdff dff_A_lNU0yOKL0_0(.dout(w_n797_6[0]),.din(w_dff_A_lNU0yOKL0_0),.clk(gclk));
	jdff dff_A_5oygKVDc0_0(.dout(w_dff_A_lNU0yOKL0_0),.din(w_dff_A_5oygKVDc0_0),.clk(gclk));
	jdff dff_A_Oj3gjdpi9_0(.dout(w_dff_A_5oygKVDc0_0),.din(w_dff_A_Oj3gjdpi9_0),.clk(gclk));
	jdff dff_A_9heJPZ8k6_0(.dout(w_dff_A_Oj3gjdpi9_0),.din(w_dff_A_9heJPZ8k6_0),.clk(gclk));
	jdff dff_A_fGTiVtRK4_0(.dout(w_dff_A_9heJPZ8k6_0),.din(w_dff_A_fGTiVtRK4_0),.clk(gclk));
	jdff dff_A_nQQgaYQw0_0(.dout(w_dff_A_fGTiVtRK4_0),.din(w_dff_A_nQQgaYQw0_0),.clk(gclk));
	jdff dff_A_YLZyl7P60_0(.dout(w_dff_A_nQQgaYQw0_0),.din(w_dff_A_YLZyl7P60_0),.clk(gclk));
	jdff dff_A_Moh6W1In2_0(.dout(w_dff_A_YLZyl7P60_0),.din(w_dff_A_Moh6W1In2_0),.clk(gclk));
	jdff dff_A_PMi9rjUu8_0(.dout(w_dff_A_Moh6W1In2_0),.din(w_dff_A_PMi9rjUu8_0),.clk(gclk));
	jdff dff_A_ZKnW40b80_0(.dout(w_dff_A_PMi9rjUu8_0),.din(w_dff_A_ZKnW40b80_0),.clk(gclk));
	jdff dff_A_Z8AzZGpY8_0(.dout(w_dff_A_ZKnW40b80_0),.din(w_dff_A_Z8AzZGpY8_0),.clk(gclk));
	jdff dff_A_gSJ0gdUE4_0(.dout(w_dff_A_Z8AzZGpY8_0),.din(w_dff_A_gSJ0gdUE4_0),.clk(gclk));
	jdff dff_A_YvUVRR3i0_0(.dout(w_dff_A_gSJ0gdUE4_0),.din(w_dff_A_YvUVRR3i0_0),.clk(gclk));
	jdff dff_A_W1rNttzp8_0(.dout(w_dff_A_YvUVRR3i0_0),.din(w_dff_A_W1rNttzp8_0),.clk(gclk));
	jdff dff_A_U71Wqot97_0(.dout(w_dff_A_W1rNttzp8_0),.din(w_dff_A_U71Wqot97_0),.clk(gclk));
	jdff dff_A_THkQBd0N4_0(.dout(w_dff_A_U71Wqot97_0),.din(w_dff_A_THkQBd0N4_0),.clk(gclk));
	jdff dff_A_sQllPZOP3_0(.dout(w_dff_A_THkQBd0N4_0),.din(w_dff_A_sQllPZOP3_0),.clk(gclk));
	jdff dff_A_M3Jx9hsM7_0(.dout(w_dff_A_sQllPZOP3_0),.din(w_dff_A_M3Jx9hsM7_0),.clk(gclk));
	jdff dff_A_m3CNYkjw4_0(.dout(w_dff_A_M3Jx9hsM7_0),.din(w_dff_A_m3CNYkjw4_0),.clk(gclk));
	jdff dff_A_tb1vKi2D2_0(.dout(w_dff_A_m3CNYkjw4_0),.din(w_dff_A_tb1vKi2D2_0),.clk(gclk));
	jdff dff_A_ZBIkZu7l7_2(.dout(w_n797_6[2]),.din(w_dff_A_ZBIkZu7l7_2),.clk(gclk));
	jdff dff_A_6Wjp8grj5_2(.dout(w_dff_A_ZBIkZu7l7_2),.din(w_dff_A_6Wjp8grj5_2),.clk(gclk));
	jdff dff_A_T3SAIYIW2_2(.dout(w_dff_A_6Wjp8grj5_2),.din(w_dff_A_T3SAIYIW2_2),.clk(gclk));
	jdff dff_A_kw7EHbiv4_2(.dout(w_dff_A_T3SAIYIW2_2),.din(w_dff_A_kw7EHbiv4_2),.clk(gclk));
	jdff dff_A_NtF6MYvO1_2(.dout(w_dff_A_kw7EHbiv4_2),.din(w_dff_A_NtF6MYvO1_2),.clk(gclk));
	jdff dff_A_6tCwbCYX8_2(.dout(w_dff_A_NtF6MYvO1_2),.din(w_dff_A_6tCwbCYX8_2),.clk(gclk));
	jdff dff_A_apcfSdi74_2(.dout(w_dff_A_6tCwbCYX8_2),.din(w_dff_A_apcfSdi74_2),.clk(gclk));
	jdff dff_A_ATFi6iuZ7_2(.dout(w_dff_A_apcfSdi74_2),.din(w_dff_A_ATFi6iuZ7_2),.clk(gclk));
	jdff dff_A_xAlNmWun0_2(.dout(w_dff_A_ATFi6iuZ7_2),.din(w_dff_A_xAlNmWun0_2),.clk(gclk));
	jdff dff_A_j40pknwC0_2(.dout(w_dff_A_xAlNmWun0_2),.din(w_dff_A_j40pknwC0_2),.clk(gclk));
	jdff dff_A_Ll5Z3cAM9_2(.dout(w_dff_A_j40pknwC0_2),.din(w_dff_A_Ll5Z3cAM9_2),.clk(gclk));
	jdff dff_A_xYaKMUou5_0(.dout(w_G4088_6[0]),.din(w_dff_A_xYaKMUou5_0),.clk(gclk));
	jdff dff_A_aVDGvTBl0_0(.dout(w_dff_A_xYaKMUou5_0),.din(w_dff_A_aVDGvTBl0_0),.clk(gclk));
	jdff dff_A_RxSHQLeR8_0(.dout(w_dff_A_aVDGvTBl0_0),.din(w_dff_A_RxSHQLeR8_0),.clk(gclk));
	jdff dff_A_Nnpg2m7N6_0(.dout(w_dff_A_RxSHQLeR8_0),.din(w_dff_A_Nnpg2m7N6_0),.clk(gclk));
	jdff dff_A_Ir6YNkOk1_0(.dout(w_dff_A_Nnpg2m7N6_0),.din(w_dff_A_Ir6YNkOk1_0),.clk(gclk));
	jdff dff_A_bz7cpQx72_0(.dout(w_dff_A_Ir6YNkOk1_0),.din(w_dff_A_bz7cpQx72_0),.clk(gclk));
	jdff dff_A_4tC039Cp9_0(.dout(w_dff_A_bz7cpQx72_0),.din(w_dff_A_4tC039Cp9_0),.clk(gclk));
	jdff dff_A_3vRFSR4i9_0(.dout(w_dff_A_4tC039Cp9_0),.din(w_dff_A_3vRFSR4i9_0),.clk(gclk));
	jdff dff_A_5vdkZwtE7_0(.dout(w_dff_A_3vRFSR4i9_0),.din(w_dff_A_5vdkZwtE7_0),.clk(gclk));
	jdff dff_A_a4OH2zoE8_0(.dout(w_dff_A_5vdkZwtE7_0),.din(w_dff_A_a4OH2zoE8_0),.clk(gclk));
	jdff dff_A_w2IaFdIS4_0(.dout(w_dff_A_a4OH2zoE8_0),.din(w_dff_A_w2IaFdIS4_0),.clk(gclk));
	jdff dff_A_XhCivb6b2_0(.dout(w_dff_A_w2IaFdIS4_0),.din(w_dff_A_XhCivb6b2_0),.clk(gclk));
	jdff dff_A_TjHKLjft5_0(.dout(w_dff_A_XhCivb6b2_0),.din(w_dff_A_TjHKLjft5_0),.clk(gclk));
	jdff dff_A_CPCe5i563_0(.dout(w_dff_A_TjHKLjft5_0),.din(w_dff_A_CPCe5i563_0),.clk(gclk));
	jdff dff_A_0owSNGe31_0(.dout(w_dff_A_CPCe5i563_0),.din(w_dff_A_0owSNGe31_0),.clk(gclk));
	jdff dff_A_mCWSBeBZ3_0(.dout(w_dff_A_0owSNGe31_0),.din(w_dff_A_mCWSBeBZ3_0),.clk(gclk));
	jdff dff_A_Gop5yYRW1_0(.dout(w_dff_A_mCWSBeBZ3_0),.din(w_dff_A_Gop5yYRW1_0),.clk(gclk));
	jdff dff_A_ANmvAQjt5_0(.dout(w_dff_A_Gop5yYRW1_0),.din(w_dff_A_ANmvAQjt5_0),.clk(gclk));
	jdff dff_A_EpucYBj75_0(.dout(w_dff_A_ANmvAQjt5_0),.din(w_dff_A_EpucYBj75_0),.clk(gclk));
	jdff dff_A_UAnolVtf5_0(.dout(w_dff_A_EpucYBj75_0),.din(w_dff_A_UAnolVtf5_0),.clk(gclk));
	jdff dff_A_UL2OIh3Q1_2(.dout(w_G4088_6[2]),.din(w_dff_A_UL2OIh3Q1_2),.clk(gclk));
	jdff dff_A_bHQMXbCU3_2(.dout(w_dff_A_UL2OIh3Q1_2),.din(w_dff_A_bHQMXbCU3_2),.clk(gclk));
	jdff dff_A_wkO4e9Mb7_2(.dout(w_dff_A_bHQMXbCU3_2),.din(w_dff_A_wkO4e9Mb7_2),.clk(gclk));
	jdff dff_A_X2obzv4Q0_2(.dout(w_dff_A_wkO4e9Mb7_2),.din(w_dff_A_X2obzv4Q0_2),.clk(gclk));
	jdff dff_A_5nRUB4HX9_2(.dout(w_dff_A_X2obzv4Q0_2),.din(w_dff_A_5nRUB4HX9_2),.clk(gclk));
	jdff dff_A_OYYFGldD6_2(.dout(w_dff_A_5nRUB4HX9_2),.din(w_dff_A_OYYFGldD6_2),.clk(gclk));
	jdff dff_A_5CJESW8C2_2(.dout(w_dff_A_OYYFGldD6_2),.din(w_dff_A_5CJESW8C2_2),.clk(gclk));
	jdff dff_A_Z56cqX7z9_2(.dout(w_dff_A_5CJESW8C2_2),.din(w_dff_A_Z56cqX7z9_2),.clk(gclk));
	jdff dff_A_4nEIVHXF1_2(.dout(w_dff_A_Z56cqX7z9_2),.din(w_dff_A_4nEIVHXF1_2),.clk(gclk));
	jdff dff_A_6X6eDHsP7_2(.dout(w_dff_A_4nEIVHXF1_2),.din(w_dff_A_6X6eDHsP7_2),.clk(gclk));
	jdff dff_A_NJJxwybQ5_2(.dout(w_dff_A_6X6eDHsP7_2),.din(w_dff_A_NJJxwybQ5_2),.clk(gclk));
	jdff dff_A_HPTCquTi3_2(.dout(w_dff_A_NJJxwybQ5_2),.din(w_dff_A_HPTCquTi3_2),.clk(gclk));
	jdff dff_A_xCSFowHo3_2(.dout(w_dff_A_HPTCquTi3_2),.din(w_dff_A_xCSFowHo3_2),.clk(gclk));
	jdff dff_A_ycHHp8f25_2(.dout(w_dff_A_xCSFowHo3_2),.din(w_dff_A_ycHHp8f25_2),.clk(gclk));
	jdff dff_B_ib0tolKH8_0(.din(n1286),.dout(w_dff_B_ib0tolKH8_0),.clk(gclk));
	jdff dff_B_ZHJTGL6T5_0(.din(w_dff_B_ib0tolKH8_0),.dout(w_dff_B_ZHJTGL6T5_0),.clk(gclk));
	jdff dff_B_rrzrgDyO1_0(.din(w_dff_B_ZHJTGL6T5_0),.dout(w_dff_B_rrzrgDyO1_0),.clk(gclk));
	jdff dff_B_rZKLo1xI4_0(.din(w_dff_B_rrzrgDyO1_0),.dout(w_dff_B_rZKLo1xI4_0),.clk(gclk));
	jdff dff_B_HgiEKKdQ0_0(.din(w_dff_B_rZKLo1xI4_0),.dout(w_dff_B_HgiEKKdQ0_0),.clk(gclk));
	jdff dff_B_ze0IZd1g9_0(.din(w_dff_B_HgiEKKdQ0_0),.dout(w_dff_B_ze0IZd1g9_0),.clk(gclk));
	jdff dff_B_nr8ZFi4z4_0(.din(w_dff_B_ze0IZd1g9_0),.dout(w_dff_B_nr8ZFi4z4_0),.clk(gclk));
	jdff dff_B_f3FXnLPP7_0(.din(w_dff_B_nr8ZFi4z4_0),.dout(w_dff_B_f3FXnLPP7_0),.clk(gclk));
	jdff dff_B_UEjY8Sqi8_0(.din(w_dff_B_f3FXnLPP7_0),.dout(w_dff_B_UEjY8Sqi8_0),.clk(gclk));
	jdff dff_B_CZsidcyL3_0(.din(w_dff_B_UEjY8Sqi8_0),.dout(w_dff_B_CZsidcyL3_0),.clk(gclk));
	jdff dff_B_KwH0vJ9X5_0(.din(w_dff_B_CZsidcyL3_0),.dout(w_dff_B_KwH0vJ9X5_0),.clk(gclk));
	jdff dff_B_jK4BFWzy9_0(.din(w_dff_B_KwH0vJ9X5_0),.dout(w_dff_B_jK4BFWzy9_0),.clk(gclk));
	jdff dff_B_xRRWSQSy0_0(.din(w_dff_B_jK4BFWzy9_0),.dout(w_dff_B_xRRWSQSy0_0),.clk(gclk));
	jdff dff_B_zDEEEJlf7_0(.din(w_dff_B_xRRWSQSy0_0),.dout(w_dff_B_zDEEEJlf7_0),.clk(gclk));
	jdff dff_B_xj7QYRbn9_0(.din(w_dff_B_zDEEEJlf7_0),.dout(w_dff_B_xj7QYRbn9_0),.clk(gclk));
	jdff dff_B_sE56QogI2_0(.din(w_dff_B_xj7QYRbn9_0),.dout(w_dff_B_sE56QogI2_0),.clk(gclk));
	jdff dff_B_iMDAzPsU1_0(.din(w_dff_B_sE56QogI2_0),.dout(w_dff_B_iMDAzPsU1_0),.clk(gclk));
	jdff dff_B_2tifSvW78_0(.din(w_dff_B_iMDAzPsU1_0),.dout(w_dff_B_2tifSvW78_0),.clk(gclk));
	jdff dff_B_ydx6ld577_0(.din(w_dff_B_2tifSvW78_0),.dout(w_dff_B_ydx6ld577_0),.clk(gclk));
	jdff dff_B_EGaddTYu8_0(.din(w_dff_B_ydx6ld577_0),.dout(w_dff_B_EGaddTYu8_0),.clk(gclk));
	jdff dff_B_L6RmGUHe6_1(.din(n1278),.dout(w_dff_B_L6RmGUHe6_1),.clk(gclk));
	jdff dff_B_humdkuXK2_1(.din(w_dff_B_L6RmGUHe6_1),.dout(w_dff_B_humdkuXK2_1),.clk(gclk));
	jdff dff_A_BU7ua3pb8_1(.dout(w_n797_5[1]),.din(w_dff_A_BU7ua3pb8_1),.clk(gclk));
	jdff dff_A_NzWahemj5_1(.dout(w_dff_A_BU7ua3pb8_1),.din(w_dff_A_NzWahemj5_1),.clk(gclk));
	jdff dff_A_5hpZymzW3_1(.dout(w_dff_A_NzWahemj5_1),.din(w_dff_A_5hpZymzW3_1),.clk(gclk));
	jdff dff_A_50tdOzGC6_1(.dout(w_dff_A_5hpZymzW3_1),.din(w_dff_A_50tdOzGC6_1),.clk(gclk));
	jdff dff_A_NCM9XFF52_1(.dout(w_dff_A_50tdOzGC6_1),.din(w_dff_A_NCM9XFF52_1),.clk(gclk));
	jdff dff_A_jOjA4B3G5_1(.dout(w_dff_A_NCM9XFF52_1),.din(w_dff_A_jOjA4B3G5_1),.clk(gclk));
	jdff dff_A_t6JmLTNz6_1(.dout(w_dff_A_jOjA4B3G5_1),.din(w_dff_A_t6JmLTNz6_1),.clk(gclk));
	jdff dff_A_CL7LuoBa3_1(.dout(w_dff_A_t6JmLTNz6_1),.din(w_dff_A_CL7LuoBa3_1),.clk(gclk));
	jdff dff_A_E07EwdgE8_1(.dout(w_dff_A_CL7LuoBa3_1),.din(w_dff_A_E07EwdgE8_1),.clk(gclk));
	jdff dff_A_l26b1K5J8_1(.dout(w_dff_A_E07EwdgE8_1),.din(w_dff_A_l26b1K5J8_1),.clk(gclk));
	jdff dff_A_X8EoCYOa1_1(.dout(w_dff_A_l26b1K5J8_1),.din(w_dff_A_X8EoCYOa1_1),.clk(gclk));
	jdff dff_A_Bfwzorlg8_1(.dout(w_dff_A_X8EoCYOa1_1),.din(w_dff_A_Bfwzorlg8_1),.clk(gclk));
	jdff dff_A_7dZYS9B62_1(.dout(w_dff_A_Bfwzorlg8_1),.din(w_dff_A_7dZYS9B62_1),.clk(gclk));
	jdff dff_A_eJL18UmO4_1(.dout(w_dff_A_7dZYS9B62_1),.din(w_dff_A_eJL18UmO4_1),.clk(gclk));
	jdff dff_A_i4rtBFi63_1(.dout(w_dff_A_eJL18UmO4_1),.din(w_dff_A_i4rtBFi63_1),.clk(gclk));
	jdff dff_A_x9mLeMmb5_1(.dout(w_dff_A_i4rtBFi63_1),.din(w_dff_A_x9mLeMmb5_1),.clk(gclk));
	jdff dff_A_AprcE3Le9_1(.dout(w_dff_A_x9mLeMmb5_1),.din(w_dff_A_AprcE3Le9_1),.clk(gclk));
	jdff dff_A_vENDE7u71_1(.dout(w_dff_A_AprcE3Le9_1),.din(w_dff_A_vENDE7u71_1),.clk(gclk));
	jdff dff_A_a30Dc9h31_1(.dout(w_dff_A_vENDE7u71_1),.din(w_dff_A_a30Dc9h31_1),.clk(gclk));
	jdff dff_A_nERkjmNx0_1(.dout(w_G4088_5[1]),.din(w_dff_A_nERkjmNx0_1),.clk(gclk));
	jdff dff_A_2B9x6Pbt1_1(.dout(w_dff_A_nERkjmNx0_1),.din(w_dff_A_2B9x6Pbt1_1),.clk(gclk));
	jdff dff_A_E1ohL8k44_1(.dout(w_dff_A_2B9x6Pbt1_1),.din(w_dff_A_E1ohL8k44_1),.clk(gclk));
	jdff dff_A_CDMp4Ikt7_1(.dout(w_dff_A_E1ohL8k44_1),.din(w_dff_A_CDMp4Ikt7_1),.clk(gclk));
	jdff dff_A_QRTRrZUQ5_1(.dout(w_dff_A_CDMp4Ikt7_1),.din(w_dff_A_QRTRrZUQ5_1),.clk(gclk));
	jdff dff_A_1TQ1Sbgq5_1(.dout(w_dff_A_QRTRrZUQ5_1),.din(w_dff_A_1TQ1Sbgq5_1),.clk(gclk));
	jdff dff_A_0yJBJbhp4_1(.dout(w_dff_A_1TQ1Sbgq5_1),.din(w_dff_A_0yJBJbhp4_1),.clk(gclk));
	jdff dff_A_RpM7D0SV8_1(.dout(w_dff_A_0yJBJbhp4_1),.din(w_dff_A_RpM7D0SV8_1),.clk(gclk));
	jdff dff_A_fpNWQqcX6_1(.dout(w_dff_A_RpM7D0SV8_1),.din(w_dff_A_fpNWQqcX6_1),.clk(gclk));
	jdff dff_A_DnYYmT1e8_1(.dout(w_dff_A_fpNWQqcX6_1),.din(w_dff_A_DnYYmT1e8_1),.clk(gclk));
	jdff dff_A_9fTUwbFM1_1(.dout(w_dff_A_DnYYmT1e8_1),.din(w_dff_A_9fTUwbFM1_1),.clk(gclk));
	jdff dff_A_NkOUE4QV9_1(.dout(w_dff_A_9fTUwbFM1_1),.din(w_dff_A_NkOUE4QV9_1),.clk(gclk));
	jdff dff_A_KCDM5riV0_1(.dout(w_dff_A_NkOUE4QV9_1),.din(w_dff_A_KCDM5riV0_1),.clk(gclk));
	jdff dff_A_iveCsrqg5_1(.dout(w_dff_A_KCDM5riV0_1),.din(w_dff_A_iveCsrqg5_1),.clk(gclk));
	jdff dff_A_enNOYNb38_1(.dout(w_dff_A_iveCsrqg5_1),.din(w_dff_A_enNOYNb38_1),.clk(gclk));
	jdff dff_A_MW1Bc9OL0_1(.dout(w_dff_A_enNOYNb38_1),.din(w_dff_A_MW1Bc9OL0_1),.clk(gclk));
	jdff dff_A_0cPIuAtG6_1(.dout(w_dff_A_MW1Bc9OL0_1),.din(w_dff_A_0cPIuAtG6_1),.clk(gclk));
	jdff dff_A_qmWfOSdh2_1(.dout(w_dff_A_0cPIuAtG6_1),.din(w_dff_A_qmWfOSdh2_1),.clk(gclk));
	jdff dff_A_cevV5e9A0_1(.dout(w_dff_A_qmWfOSdh2_1),.din(w_dff_A_cevV5e9A0_1),.clk(gclk));
	jdff dff_B_Kgrl6t8O0_0(.din(n1295),.dout(w_dff_B_Kgrl6t8O0_0),.clk(gclk));
	jdff dff_B_DLZeU8Xl6_0(.din(w_dff_B_Kgrl6t8O0_0),.dout(w_dff_B_DLZeU8Xl6_0),.clk(gclk));
	jdff dff_B_sMp9HhWS2_0(.din(w_dff_B_DLZeU8Xl6_0),.dout(w_dff_B_sMp9HhWS2_0),.clk(gclk));
	jdff dff_B_g9U9IYyX3_0(.din(w_dff_B_sMp9HhWS2_0),.dout(w_dff_B_g9U9IYyX3_0),.clk(gclk));
	jdff dff_B_YwCy8oZN3_0(.din(w_dff_B_g9U9IYyX3_0),.dout(w_dff_B_YwCy8oZN3_0),.clk(gclk));
	jdff dff_B_wMXNHpyY5_0(.din(w_dff_B_YwCy8oZN3_0),.dout(w_dff_B_wMXNHpyY5_0),.clk(gclk));
	jdff dff_B_Sx8LJqTa0_0(.din(w_dff_B_wMXNHpyY5_0),.dout(w_dff_B_Sx8LJqTa0_0),.clk(gclk));
	jdff dff_B_Ffcd17VR9_0(.din(w_dff_B_Sx8LJqTa0_0),.dout(w_dff_B_Ffcd17VR9_0),.clk(gclk));
	jdff dff_B_IH7fL4Nm9_0(.din(w_dff_B_Ffcd17VR9_0),.dout(w_dff_B_IH7fL4Nm9_0),.clk(gclk));
	jdff dff_B_IpeAaenE6_0(.din(w_dff_B_IH7fL4Nm9_0),.dout(w_dff_B_IpeAaenE6_0),.clk(gclk));
	jdff dff_B_7BFlbH6r1_0(.din(w_dff_B_IpeAaenE6_0),.dout(w_dff_B_7BFlbH6r1_0),.clk(gclk));
	jdff dff_B_kBY2X3PQ8_0(.din(w_dff_B_7BFlbH6r1_0),.dout(w_dff_B_kBY2X3PQ8_0),.clk(gclk));
	jdff dff_B_dZxcuT3S9_0(.din(w_dff_B_kBY2X3PQ8_0),.dout(w_dff_B_dZxcuT3S9_0),.clk(gclk));
	jdff dff_B_pjaLm7MK4_0(.din(w_dff_B_dZxcuT3S9_0),.dout(w_dff_B_pjaLm7MK4_0),.clk(gclk));
	jdff dff_B_42xHG2kJ5_0(.din(w_dff_B_pjaLm7MK4_0),.dout(w_dff_B_42xHG2kJ5_0),.clk(gclk));
	jdff dff_B_UydGTAgU1_0(.din(w_dff_B_42xHG2kJ5_0),.dout(w_dff_B_UydGTAgU1_0),.clk(gclk));
	jdff dff_B_c9vALxBW9_0(.din(w_dff_B_UydGTAgU1_0),.dout(w_dff_B_c9vALxBW9_0),.clk(gclk));
	jdff dff_B_JhodgRi09_0(.din(w_dff_B_c9vALxBW9_0),.dout(w_dff_B_JhodgRi09_0),.clk(gclk));
	jdff dff_B_MLLz04vA7_0(.din(w_dff_B_JhodgRi09_0),.dout(w_dff_B_MLLz04vA7_0),.clk(gclk));
	jdff dff_B_TSdQhI3G0_0(.din(w_dff_B_MLLz04vA7_0),.dout(w_dff_B_TSdQhI3G0_0),.clk(gclk));
	jdff dff_B_IzLWxCMd6_1(.din(n1288),.dout(w_dff_B_IzLWxCMd6_1),.clk(gclk));
	jdff dff_A_4tE30Vwy7_2(.dout(w_n800_2[2]),.din(w_dff_A_4tE30Vwy7_2),.clk(gclk));
	jdff dff_B_vSewMB1y0_0(.din(n1306),.dout(w_dff_B_vSewMB1y0_0),.clk(gclk));
	jdff dff_B_K9I4zaTN6_0(.din(w_dff_B_vSewMB1y0_0),.dout(w_dff_B_K9I4zaTN6_0),.clk(gclk));
	jdff dff_B_o2NWN9GO7_0(.din(w_dff_B_K9I4zaTN6_0),.dout(w_dff_B_o2NWN9GO7_0),.clk(gclk));
	jdff dff_B_vmfxdA4W9_0(.din(w_dff_B_o2NWN9GO7_0),.dout(w_dff_B_vmfxdA4W9_0),.clk(gclk));
	jdff dff_B_cbtK9TAa6_0(.din(w_dff_B_vmfxdA4W9_0),.dout(w_dff_B_cbtK9TAa6_0),.clk(gclk));
	jdff dff_B_7hdcCF510_0(.din(w_dff_B_cbtK9TAa6_0),.dout(w_dff_B_7hdcCF510_0),.clk(gclk));
	jdff dff_B_MnZpJsH21_0(.din(w_dff_B_7hdcCF510_0),.dout(w_dff_B_MnZpJsH21_0),.clk(gclk));
	jdff dff_B_GLoHxRd08_0(.din(w_dff_B_MnZpJsH21_0),.dout(w_dff_B_GLoHxRd08_0),.clk(gclk));
	jdff dff_B_o5P7f0169_0(.din(w_dff_B_GLoHxRd08_0),.dout(w_dff_B_o5P7f0169_0),.clk(gclk));
	jdff dff_B_A2ZDyqOk5_0(.din(w_dff_B_o5P7f0169_0),.dout(w_dff_B_A2ZDyqOk5_0),.clk(gclk));
	jdff dff_B_hmoUdjim9_0(.din(w_dff_B_A2ZDyqOk5_0),.dout(w_dff_B_hmoUdjim9_0),.clk(gclk));
	jdff dff_B_H7AUu1EA1_0(.din(w_dff_B_hmoUdjim9_0),.dout(w_dff_B_H7AUu1EA1_0),.clk(gclk));
	jdff dff_B_O1AictfI4_0(.din(w_dff_B_H7AUu1EA1_0),.dout(w_dff_B_O1AictfI4_0),.clk(gclk));
	jdff dff_B_HoPAZZOw6_0(.din(w_dff_B_O1AictfI4_0),.dout(w_dff_B_HoPAZZOw6_0),.clk(gclk));
	jdff dff_B_EcNXww7o1_0(.din(w_dff_B_HoPAZZOw6_0),.dout(w_dff_B_EcNXww7o1_0),.clk(gclk));
	jdff dff_B_q3PBkS4d2_0(.din(w_dff_B_EcNXww7o1_0),.dout(w_dff_B_q3PBkS4d2_0),.clk(gclk));
	jdff dff_B_Fbl7Xien0_0(.din(w_dff_B_q3PBkS4d2_0),.dout(w_dff_B_Fbl7Xien0_0),.clk(gclk));
	jdff dff_B_qn5bWogX8_0(.din(w_dff_B_Fbl7Xien0_0),.dout(w_dff_B_qn5bWogX8_0),.clk(gclk));
	jdff dff_B_aZcDLtDG6_0(.din(w_dff_B_qn5bWogX8_0),.dout(w_dff_B_aZcDLtDG6_0),.clk(gclk));
	jdff dff_B_Jq7OWrXU8_1(.din(n1298),.dout(w_dff_B_Jq7OWrXU8_1),.clk(gclk));
	jdff dff_B_ovKHhbdz1_1(.din(w_dff_B_Jq7OWrXU8_1),.dout(w_dff_B_ovKHhbdz1_1),.clk(gclk));
	jdff dff_B_Q8ABeuZd7_1(.din(w_dff_B_ovKHhbdz1_1),.dout(w_dff_B_Q8ABeuZd7_1),.clk(gclk));
	jdff dff_A_ki0ASF4M8_0(.dout(w_n797_4[0]),.din(w_dff_A_ki0ASF4M8_0),.clk(gclk));
	jdff dff_A_lFomooOb5_0(.dout(w_dff_A_ki0ASF4M8_0),.din(w_dff_A_lFomooOb5_0),.clk(gclk));
	jdff dff_A_ZrhT11cM2_0(.dout(w_dff_A_lFomooOb5_0),.din(w_dff_A_ZrhT11cM2_0),.clk(gclk));
	jdff dff_A_3gcMCGJO1_0(.dout(w_dff_A_ZrhT11cM2_0),.din(w_dff_A_3gcMCGJO1_0),.clk(gclk));
	jdff dff_A_WwunhunA1_0(.dout(w_dff_A_3gcMCGJO1_0),.din(w_dff_A_WwunhunA1_0),.clk(gclk));
	jdff dff_A_NbYHYZhP2_0(.dout(w_dff_A_WwunhunA1_0),.din(w_dff_A_NbYHYZhP2_0),.clk(gclk));
	jdff dff_A_Ubr6QMM37_0(.dout(w_dff_A_NbYHYZhP2_0),.din(w_dff_A_Ubr6QMM37_0),.clk(gclk));
	jdff dff_A_KlvC5Bed3_0(.dout(w_dff_A_Ubr6QMM37_0),.din(w_dff_A_KlvC5Bed3_0),.clk(gclk));
	jdff dff_A_bpKVYhvG2_0(.dout(w_dff_A_KlvC5Bed3_0),.din(w_dff_A_bpKVYhvG2_0),.clk(gclk));
	jdff dff_A_14KvqGfs6_0(.dout(w_dff_A_bpKVYhvG2_0),.din(w_dff_A_14KvqGfs6_0),.clk(gclk));
	jdff dff_A_dugp3Xvq2_0(.dout(w_dff_A_14KvqGfs6_0),.din(w_dff_A_dugp3Xvq2_0),.clk(gclk));
	jdff dff_A_EfMp3gX20_0(.dout(w_dff_A_dugp3Xvq2_0),.din(w_dff_A_EfMp3gX20_0),.clk(gclk));
	jdff dff_A_GSPtApM15_0(.dout(w_dff_A_EfMp3gX20_0),.din(w_dff_A_GSPtApM15_0),.clk(gclk));
	jdff dff_A_sxe1NpZs7_0(.dout(w_dff_A_GSPtApM15_0),.din(w_dff_A_sxe1NpZs7_0),.clk(gclk));
	jdff dff_A_pw6QaPsH7_0(.dout(w_dff_A_sxe1NpZs7_0),.din(w_dff_A_pw6QaPsH7_0),.clk(gclk));
	jdff dff_A_QLx6BECE6_0(.dout(w_dff_A_pw6QaPsH7_0),.din(w_dff_A_QLx6BECE6_0),.clk(gclk));
	jdff dff_A_jMObl2In7_0(.dout(w_dff_A_QLx6BECE6_0),.din(w_dff_A_jMObl2In7_0),.clk(gclk));
	jdff dff_A_58dpKpKG9_0(.dout(w_dff_A_jMObl2In7_0),.din(w_dff_A_58dpKpKG9_0),.clk(gclk));
	jdff dff_A_7j2i70Da2_2(.dout(w_n797_4[2]),.din(w_dff_A_7j2i70Da2_2),.clk(gclk));
	jdff dff_A_5saTnAlU9_2(.dout(w_dff_A_7j2i70Da2_2),.din(w_dff_A_5saTnAlU9_2),.clk(gclk));
	jdff dff_A_wOJZlyW08_2(.dout(w_dff_A_5saTnAlU9_2),.din(w_dff_A_wOJZlyW08_2),.clk(gclk));
	jdff dff_A_rW2uadle0_2(.dout(w_dff_A_wOJZlyW08_2),.din(w_dff_A_rW2uadle0_2),.clk(gclk));
	jdff dff_A_QeePR53M7_2(.dout(w_dff_A_rW2uadle0_2),.din(w_dff_A_QeePR53M7_2),.clk(gclk));
	jdff dff_A_tXPiKJdB2_2(.dout(w_dff_A_QeePR53M7_2),.din(w_dff_A_tXPiKJdB2_2),.clk(gclk));
	jdff dff_A_HUASIeDg1_2(.dout(w_dff_A_tXPiKJdB2_2),.din(w_dff_A_HUASIeDg1_2),.clk(gclk));
	jdff dff_A_3iIQOlkU6_2(.dout(w_dff_A_HUASIeDg1_2),.din(w_dff_A_3iIQOlkU6_2),.clk(gclk));
	jdff dff_A_FKKUxtHb1_2(.dout(w_dff_A_3iIQOlkU6_2),.din(w_dff_A_FKKUxtHb1_2),.clk(gclk));
	jdff dff_A_BeAran7r8_2(.dout(w_dff_A_FKKUxtHb1_2),.din(w_dff_A_BeAran7r8_2),.clk(gclk));
	jdff dff_A_mnwn4CYJ5_2(.dout(w_dff_A_BeAran7r8_2),.din(w_dff_A_mnwn4CYJ5_2),.clk(gclk));
	jdff dff_A_wmHjxtnJ2_2(.dout(w_dff_A_mnwn4CYJ5_2),.din(w_dff_A_wmHjxtnJ2_2),.clk(gclk));
	jdff dff_A_tTGgUwVC5_2(.dout(w_dff_A_wmHjxtnJ2_2),.din(w_dff_A_tTGgUwVC5_2),.clk(gclk));
	jdff dff_A_0k1q2xTD9_2(.dout(w_dff_A_tTGgUwVC5_2),.din(w_dff_A_0k1q2xTD9_2),.clk(gclk));
	jdff dff_A_778z624G2_2(.dout(w_dff_A_0k1q2xTD9_2),.din(w_dff_A_778z624G2_2),.clk(gclk));
	jdff dff_A_HUKVj8fA4_2(.dout(w_dff_A_778z624G2_2),.din(w_dff_A_HUKVj8fA4_2),.clk(gclk));
	jdff dff_A_K6Iq2SXH5_2(.dout(w_dff_A_HUKVj8fA4_2),.din(w_dff_A_K6Iq2SXH5_2),.clk(gclk));
	jdff dff_A_rh61vUaI2_2(.dout(w_dff_A_K6Iq2SXH5_2),.din(w_dff_A_rh61vUaI2_2),.clk(gclk));
	jdff dff_A_vwgUazEv3_2(.dout(w_dff_A_rh61vUaI2_2),.din(w_dff_A_vwgUazEv3_2),.clk(gclk));
	jdff dff_A_q0V7oPRS2_0(.dout(w_G4088_4[0]),.din(w_dff_A_q0V7oPRS2_0),.clk(gclk));
	jdff dff_A_JTX3UDzV4_0(.dout(w_dff_A_q0V7oPRS2_0),.din(w_dff_A_JTX3UDzV4_0),.clk(gclk));
	jdff dff_A_Iyijq3FQ7_0(.dout(w_dff_A_JTX3UDzV4_0),.din(w_dff_A_Iyijq3FQ7_0),.clk(gclk));
	jdff dff_A_1kc3LsSs4_0(.dout(w_dff_A_Iyijq3FQ7_0),.din(w_dff_A_1kc3LsSs4_0),.clk(gclk));
	jdff dff_A_itu51oVY4_0(.dout(w_dff_A_1kc3LsSs4_0),.din(w_dff_A_itu51oVY4_0),.clk(gclk));
	jdff dff_A_s6sk633O5_0(.dout(w_dff_A_itu51oVY4_0),.din(w_dff_A_s6sk633O5_0),.clk(gclk));
	jdff dff_A_VOyMETQt6_0(.dout(w_dff_A_s6sk633O5_0),.din(w_dff_A_VOyMETQt6_0),.clk(gclk));
	jdff dff_A_R8iQ81MI1_0(.dout(w_dff_A_VOyMETQt6_0),.din(w_dff_A_R8iQ81MI1_0),.clk(gclk));
	jdff dff_A_nqY2Uh666_0(.dout(w_dff_A_R8iQ81MI1_0),.din(w_dff_A_nqY2Uh666_0),.clk(gclk));
	jdff dff_A_Z4VBhC2g9_0(.dout(w_dff_A_nqY2Uh666_0),.din(w_dff_A_Z4VBhC2g9_0),.clk(gclk));
	jdff dff_A_EGko19t43_0(.dout(w_dff_A_Z4VBhC2g9_0),.din(w_dff_A_EGko19t43_0),.clk(gclk));
	jdff dff_A_iT981qWw0_0(.dout(w_dff_A_EGko19t43_0),.din(w_dff_A_iT981qWw0_0),.clk(gclk));
	jdff dff_A_xPFvLJPM0_0(.dout(w_dff_A_iT981qWw0_0),.din(w_dff_A_xPFvLJPM0_0),.clk(gclk));
	jdff dff_A_RBKwFwSC2_0(.dout(w_dff_A_xPFvLJPM0_0),.din(w_dff_A_RBKwFwSC2_0),.clk(gclk));
	jdff dff_A_PifznpmR9_0(.dout(w_dff_A_RBKwFwSC2_0),.din(w_dff_A_PifznpmR9_0),.clk(gclk));
	jdff dff_A_THl7v3H99_0(.dout(w_dff_A_PifznpmR9_0),.din(w_dff_A_THl7v3H99_0),.clk(gclk));
	jdff dff_A_jVEqA2kz8_0(.dout(w_dff_A_THl7v3H99_0),.din(w_dff_A_jVEqA2kz8_0),.clk(gclk));
	jdff dff_A_Jz1nKuwT1_2(.dout(w_G4088_4[2]),.din(w_dff_A_Jz1nKuwT1_2),.clk(gclk));
	jdff dff_A_ZKftlHUA6_2(.dout(w_dff_A_Jz1nKuwT1_2),.din(w_dff_A_ZKftlHUA6_2),.clk(gclk));
	jdff dff_A_QpGET3A94_2(.dout(w_dff_A_ZKftlHUA6_2),.din(w_dff_A_QpGET3A94_2),.clk(gclk));
	jdff dff_A_dpVnm63O7_2(.dout(w_dff_A_QpGET3A94_2),.din(w_dff_A_dpVnm63O7_2),.clk(gclk));
	jdff dff_A_iBsoTUgp3_2(.dout(w_dff_A_dpVnm63O7_2),.din(w_dff_A_iBsoTUgp3_2),.clk(gclk));
	jdff dff_A_pwfpBjgA7_2(.dout(w_dff_A_iBsoTUgp3_2),.din(w_dff_A_pwfpBjgA7_2),.clk(gclk));
	jdff dff_A_2heLTJ250_2(.dout(w_dff_A_pwfpBjgA7_2),.din(w_dff_A_2heLTJ250_2),.clk(gclk));
	jdff dff_A_DwYJ2Z3T6_2(.dout(w_dff_A_2heLTJ250_2),.din(w_dff_A_DwYJ2Z3T6_2),.clk(gclk));
	jdff dff_A_kL3I5mTA9_2(.dout(w_dff_A_DwYJ2Z3T6_2),.din(w_dff_A_kL3I5mTA9_2),.clk(gclk));
	jdff dff_A_On1pbqBq8_2(.dout(w_dff_A_kL3I5mTA9_2),.din(w_dff_A_On1pbqBq8_2),.clk(gclk));
	jdff dff_A_4MEsVlrA7_2(.dout(w_dff_A_On1pbqBq8_2),.din(w_dff_A_4MEsVlrA7_2),.clk(gclk));
	jdff dff_A_034kpSf43_2(.dout(w_dff_A_4MEsVlrA7_2),.din(w_dff_A_034kpSf43_2),.clk(gclk));
	jdff dff_A_PVtJZn7T6_2(.dout(w_dff_A_034kpSf43_2),.din(w_dff_A_PVtJZn7T6_2),.clk(gclk));
	jdff dff_A_44gbeMXv9_2(.dout(w_dff_A_PVtJZn7T6_2),.din(w_dff_A_44gbeMXv9_2),.clk(gclk));
	jdff dff_A_u8NlSWp98_2(.dout(w_dff_A_44gbeMXv9_2),.din(w_dff_A_u8NlSWp98_2),.clk(gclk));
	jdff dff_A_pUhPiI5Q7_2(.dout(w_dff_A_u8NlSWp98_2),.din(w_dff_A_pUhPiI5Q7_2),.clk(gclk));
	jdff dff_A_iDITvLu20_2(.dout(w_dff_A_pUhPiI5Q7_2),.din(w_dff_A_iDITvLu20_2),.clk(gclk));
	jdff dff_A_DWaEN6e94_2(.dout(w_dff_A_iDITvLu20_2),.din(w_dff_A_DWaEN6e94_2),.clk(gclk));
	jdff dff_A_YEAViCjk5_2(.dout(w_dff_A_DWaEN6e94_2),.din(w_dff_A_YEAViCjk5_2),.clk(gclk));
	jdff dff_A_SBWxVdOH5_2(.dout(w_dff_A_YEAViCjk5_2),.din(w_dff_A_SBWxVdOH5_2),.clk(gclk));
	jdff dff_B_n0JULlMa2_0(.din(n1315),.dout(w_dff_B_n0JULlMa2_0),.clk(gclk));
	jdff dff_B_6uClxzp97_0(.din(w_dff_B_n0JULlMa2_0),.dout(w_dff_B_6uClxzp97_0),.clk(gclk));
	jdff dff_B_mASb81U03_0(.din(w_dff_B_6uClxzp97_0),.dout(w_dff_B_mASb81U03_0),.clk(gclk));
	jdff dff_B_7u1vgKYg6_0(.din(w_dff_B_mASb81U03_0),.dout(w_dff_B_7u1vgKYg6_0),.clk(gclk));
	jdff dff_B_6ZiCbqQd3_0(.din(w_dff_B_7u1vgKYg6_0),.dout(w_dff_B_6ZiCbqQd3_0),.clk(gclk));
	jdff dff_B_DoasNh6g3_0(.din(w_dff_B_6ZiCbqQd3_0),.dout(w_dff_B_DoasNh6g3_0),.clk(gclk));
	jdff dff_B_ESwQ3rgW2_0(.din(w_dff_B_DoasNh6g3_0),.dout(w_dff_B_ESwQ3rgW2_0),.clk(gclk));
	jdff dff_B_LQ1ySkNK0_0(.din(w_dff_B_ESwQ3rgW2_0),.dout(w_dff_B_LQ1ySkNK0_0),.clk(gclk));
	jdff dff_B_4WIrFQMY0_0(.din(w_dff_B_LQ1ySkNK0_0),.dout(w_dff_B_4WIrFQMY0_0),.clk(gclk));
	jdff dff_B_m5LPkm6d0_0(.din(w_dff_B_4WIrFQMY0_0),.dout(w_dff_B_m5LPkm6d0_0),.clk(gclk));
	jdff dff_B_nv4Y54bF1_0(.din(w_dff_B_m5LPkm6d0_0),.dout(w_dff_B_nv4Y54bF1_0),.clk(gclk));
	jdff dff_B_66LUithL5_0(.din(w_dff_B_nv4Y54bF1_0),.dout(w_dff_B_66LUithL5_0),.clk(gclk));
	jdff dff_B_1Rt8GaNl3_0(.din(w_dff_B_66LUithL5_0),.dout(w_dff_B_1Rt8GaNl3_0),.clk(gclk));
	jdff dff_B_zPBW5Ady7_0(.din(w_dff_B_1Rt8GaNl3_0),.dout(w_dff_B_zPBW5Ady7_0),.clk(gclk));
	jdff dff_B_NYOotvNJ2_0(.din(w_dff_B_zPBW5Ady7_0),.dout(w_dff_B_NYOotvNJ2_0),.clk(gclk));
	jdff dff_B_6hQY9w0h2_0(.din(w_dff_B_NYOotvNJ2_0),.dout(w_dff_B_6hQY9w0h2_0),.clk(gclk));
	jdff dff_B_ttaq4fJM2_0(.din(w_dff_B_6hQY9w0h2_0),.dout(w_dff_B_ttaq4fJM2_0),.clk(gclk));
	jdff dff_B_uSs6b6rw5_0(.din(w_dff_B_ttaq4fJM2_0),.dout(w_dff_B_uSs6b6rw5_0),.clk(gclk));
	jdff dff_B_htTGsVSt9_0(.din(w_dff_B_uSs6b6rw5_0),.dout(w_dff_B_htTGsVSt9_0),.clk(gclk));
	jdff dff_B_pwxvlKCd3_0(.din(w_dff_B_htTGsVSt9_0),.dout(w_dff_B_pwxvlKCd3_0),.clk(gclk));
	jdff dff_B_QHr4jZ8J4_2(.din(G49),.dout(w_dff_B_QHr4jZ8J4_2),.clk(gclk));
	jdff dff_B_7nPZ3Rre2_1(.din(n1308),.dout(w_dff_B_7nPZ3Rre2_1),.clk(gclk));
	jdff dff_B_1fOuwH6L7_1(.din(w_dff_B_7nPZ3Rre2_1),.dout(w_dff_B_1fOuwH6L7_1),.clk(gclk));
	jdff dff_A_XYqQI4tr2_1(.dout(w_n852_5[1]),.din(w_dff_A_XYqQI4tr2_1),.clk(gclk));
	jdff dff_A_oq3zXX0C7_1(.dout(w_dff_A_XYqQI4tr2_1),.din(w_dff_A_oq3zXX0C7_1),.clk(gclk));
	jdff dff_A_6zqY6HDs9_1(.dout(w_dff_A_oq3zXX0C7_1),.din(w_dff_A_6zqY6HDs9_1),.clk(gclk));
	jdff dff_A_oOvmg0VM2_1(.dout(w_dff_A_6zqY6HDs9_1),.din(w_dff_A_oOvmg0VM2_1),.clk(gclk));
	jdff dff_A_cWTMDDHd3_1(.dout(w_dff_A_oOvmg0VM2_1),.din(w_dff_A_cWTMDDHd3_1),.clk(gclk));
	jdff dff_A_KmnruPb86_1(.dout(w_dff_A_cWTMDDHd3_1),.din(w_dff_A_KmnruPb86_1),.clk(gclk));
	jdff dff_A_UVi6WQcO4_1(.dout(w_dff_A_KmnruPb86_1),.din(w_dff_A_UVi6WQcO4_1),.clk(gclk));
	jdff dff_A_L0DHTAX51_1(.dout(w_dff_A_UVi6WQcO4_1),.din(w_dff_A_L0DHTAX51_1),.clk(gclk));
	jdff dff_A_8fx1SEuP8_1(.dout(w_dff_A_L0DHTAX51_1),.din(w_dff_A_8fx1SEuP8_1),.clk(gclk));
	jdff dff_A_uVTEgqv23_1(.dout(w_dff_A_8fx1SEuP8_1),.din(w_dff_A_uVTEgqv23_1),.clk(gclk));
	jdff dff_A_pem9On199_1(.dout(w_dff_A_uVTEgqv23_1),.din(w_dff_A_pem9On199_1),.clk(gclk));
	jdff dff_A_6PSyUXSh4_1(.dout(w_dff_A_pem9On199_1),.din(w_dff_A_6PSyUXSh4_1),.clk(gclk));
	jdff dff_A_w6WjhYjx1_1(.dout(w_dff_A_6PSyUXSh4_1),.din(w_dff_A_w6WjhYjx1_1),.clk(gclk));
	jdff dff_A_buocVb7d9_1(.dout(w_dff_A_w6WjhYjx1_1),.din(w_dff_A_buocVb7d9_1),.clk(gclk));
	jdff dff_A_Ewn4RtIF1_1(.dout(w_dff_A_buocVb7d9_1),.din(w_dff_A_Ewn4RtIF1_1),.clk(gclk));
	jdff dff_A_5EtBrdRd7_1(.dout(w_dff_A_Ewn4RtIF1_1),.din(w_dff_A_5EtBrdRd7_1),.clk(gclk));
	jdff dff_A_0lFLGziL8_1(.dout(w_dff_A_5EtBrdRd7_1),.din(w_dff_A_0lFLGziL8_1),.clk(gclk));
	jdff dff_A_ZCrqRcRk6_1(.dout(w_dff_A_0lFLGziL8_1),.din(w_dff_A_ZCrqRcRk6_1),.clk(gclk));
	jdff dff_A_WPWSIian4_1(.dout(w_dff_A_ZCrqRcRk6_1),.din(w_dff_A_WPWSIian4_1),.clk(gclk));
	jdff dff_A_d1MpCJDD3_2(.dout(w_n852_5[2]),.din(w_dff_A_d1MpCJDD3_2),.clk(gclk));
	jdff dff_A_3pxIiuSN9_2(.dout(w_dff_A_d1MpCJDD3_2),.din(w_dff_A_3pxIiuSN9_2),.clk(gclk));
	jdff dff_A_YSWYsvqi3_2(.dout(w_dff_A_3pxIiuSN9_2),.din(w_dff_A_YSWYsvqi3_2),.clk(gclk));
	jdff dff_A_fyPmQcVm8_2(.dout(w_dff_A_YSWYsvqi3_2),.din(w_dff_A_fyPmQcVm8_2),.clk(gclk));
	jdff dff_A_trAjfuju2_2(.dout(w_dff_A_fyPmQcVm8_2),.din(w_dff_A_trAjfuju2_2),.clk(gclk));
	jdff dff_A_FvB1Qr9T2_2(.dout(w_dff_A_trAjfuju2_2),.din(w_dff_A_FvB1Qr9T2_2),.clk(gclk));
	jdff dff_A_d94azWjj7_2(.dout(w_dff_A_FvB1Qr9T2_2),.din(w_dff_A_d94azWjj7_2),.clk(gclk));
	jdff dff_A_dghaaWEf4_2(.dout(w_dff_A_d94azWjj7_2),.din(w_dff_A_dghaaWEf4_2),.clk(gclk));
	jdff dff_A_sKsSBgEk9_2(.dout(w_dff_A_dghaaWEf4_2),.din(w_dff_A_sKsSBgEk9_2),.clk(gclk));
	jdff dff_A_Zg41apJI9_2(.dout(w_dff_A_sKsSBgEk9_2),.din(w_dff_A_Zg41apJI9_2),.clk(gclk));
	jdff dff_A_nL5LldgU1_2(.dout(w_dff_A_Zg41apJI9_2),.din(w_dff_A_nL5LldgU1_2),.clk(gclk));
	jdff dff_A_pYk34Idd7_2(.dout(w_dff_A_nL5LldgU1_2),.din(w_dff_A_pYk34Idd7_2),.clk(gclk));
	jdff dff_A_p2CFUgv18_2(.dout(w_dff_A_pYk34Idd7_2),.din(w_dff_A_p2CFUgv18_2),.clk(gclk));
	jdff dff_A_2VVTXPgh1_2(.dout(w_dff_A_p2CFUgv18_2),.din(w_dff_A_2VVTXPgh1_2),.clk(gclk));
	jdff dff_A_IXYfh8WW7_2(.dout(w_dff_A_2VVTXPgh1_2),.din(w_dff_A_IXYfh8WW7_2),.clk(gclk));
	jdff dff_A_hQSBjLl80_2(.dout(w_dff_A_IXYfh8WW7_2),.din(w_dff_A_hQSBjLl80_2),.clk(gclk));
	jdff dff_A_7U4jiEVr8_2(.dout(w_dff_A_hQSBjLl80_2),.din(w_dff_A_7U4jiEVr8_2),.clk(gclk));
	jdff dff_A_GGkEp1kd8_2(.dout(w_dff_A_7U4jiEVr8_2),.din(w_dff_A_GGkEp1kd8_2),.clk(gclk));
	jdff dff_A_i8NayOmt2_2(.dout(w_dff_A_GGkEp1kd8_2),.din(w_dff_A_i8NayOmt2_2),.clk(gclk));
	jdff dff_A_NG1cNPox5_2(.dout(w_dff_A_i8NayOmt2_2),.din(w_dff_A_NG1cNPox5_2),.clk(gclk));
	jdff dff_A_2T0YjRoR8_1(.dout(w_G4089_5[1]),.din(w_dff_A_2T0YjRoR8_1),.clk(gclk));
	jdff dff_A_ukj2lMYs3_1(.dout(w_dff_A_2T0YjRoR8_1),.din(w_dff_A_ukj2lMYs3_1),.clk(gclk));
	jdff dff_A_v3sMnOfD6_1(.dout(w_dff_A_ukj2lMYs3_1),.din(w_dff_A_v3sMnOfD6_1),.clk(gclk));
	jdff dff_A_GqDT4R8b0_1(.dout(w_dff_A_v3sMnOfD6_1),.din(w_dff_A_GqDT4R8b0_1),.clk(gclk));
	jdff dff_A_yTlniVR09_1(.dout(w_dff_A_GqDT4R8b0_1),.din(w_dff_A_yTlniVR09_1),.clk(gclk));
	jdff dff_A_xVptjahG8_1(.dout(w_dff_A_yTlniVR09_1),.din(w_dff_A_xVptjahG8_1),.clk(gclk));
	jdff dff_A_fXwbrHrn6_1(.dout(w_dff_A_xVptjahG8_1),.din(w_dff_A_fXwbrHrn6_1),.clk(gclk));
	jdff dff_A_p6MkiGPY8_1(.dout(w_dff_A_fXwbrHrn6_1),.din(w_dff_A_p6MkiGPY8_1),.clk(gclk));
	jdff dff_A_gTLj0d0T3_1(.dout(w_dff_A_p6MkiGPY8_1),.din(w_dff_A_gTLj0d0T3_1),.clk(gclk));
	jdff dff_A_ydVYs9g36_1(.dout(w_dff_A_gTLj0d0T3_1),.din(w_dff_A_ydVYs9g36_1),.clk(gclk));
	jdff dff_A_3TXZKoFM6_1(.dout(w_dff_A_ydVYs9g36_1),.din(w_dff_A_3TXZKoFM6_1),.clk(gclk));
	jdff dff_A_t7MkKv054_1(.dout(w_dff_A_3TXZKoFM6_1),.din(w_dff_A_t7MkKv054_1),.clk(gclk));
	jdff dff_A_cuEbSjxY8_1(.dout(w_dff_A_t7MkKv054_1),.din(w_dff_A_cuEbSjxY8_1),.clk(gclk));
	jdff dff_A_oVjjiMYT7_1(.dout(w_dff_A_cuEbSjxY8_1),.din(w_dff_A_oVjjiMYT7_1),.clk(gclk));
	jdff dff_A_TkRUub3H9_1(.dout(w_dff_A_oVjjiMYT7_1),.din(w_dff_A_TkRUub3H9_1),.clk(gclk));
	jdff dff_A_nx9bvsxe4_1(.dout(w_dff_A_TkRUub3H9_1),.din(w_dff_A_nx9bvsxe4_1),.clk(gclk));
	jdff dff_A_9HOC5UXP4_1(.dout(w_dff_A_nx9bvsxe4_1),.din(w_dff_A_9HOC5UXP4_1),.clk(gclk));
	jdff dff_A_WmhOFS8T7_1(.dout(w_dff_A_9HOC5UXP4_1),.din(w_dff_A_WmhOFS8T7_1),.clk(gclk));
	jdff dff_A_TBX5Mh469_1(.dout(w_dff_A_WmhOFS8T7_1),.din(w_dff_A_TBX5Mh469_1),.clk(gclk));
	jdff dff_A_8JXtxRY97_2(.dout(w_G4089_5[2]),.din(w_dff_A_8JXtxRY97_2),.clk(gclk));
	jdff dff_A_fEPr5yPk6_2(.dout(w_dff_A_8JXtxRY97_2),.din(w_dff_A_fEPr5yPk6_2),.clk(gclk));
	jdff dff_A_2EIqdY9a5_2(.dout(w_dff_A_fEPr5yPk6_2),.din(w_dff_A_2EIqdY9a5_2),.clk(gclk));
	jdff dff_A_G1ybo0jX4_2(.dout(w_dff_A_2EIqdY9a5_2),.din(w_dff_A_G1ybo0jX4_2),.clk(gclk));
	jdff dff_A_OLvqYejf3_2(.dout(w_dff_A_G1ybo0jX4_2),.din(w_dff_A_OLvqYejf3_2),.clk(gclk));
	jdff dff_A_SlkMDmm30_2(.dout(w_dff_A_OLvqYejf3_2),.din(w_dff_A_SlkMDmm30_2),.clk(gclk));
	jdff dff_A_RBqN83Ax1_2(.dout(w_dff_A_SlkMDmm30_2),.din(w_dff_A_RBqN83Ax1_2),.clk(gclk));
	jdff dff_A_rIpBa0Ap7_2(.dout(w_dff_A_RBqN83Ax1_2),.din(w_dff_A_rIpBa0Ap7_2),.clk(gclk));
	jdff dff_A_cNl0c7bd9_2(.dout(w_dff_A_rIpBa0Ap7_2),.din(w_dff_A_cNl0c7bd9_2),.clk(gclk));
	jdff dff_A_OXGOCku81_2(.dout(w_dff_A_cNl0c7bd9_2),.din(w_dff_A_OXGOCku81_2),.clk(gclk));
	jdff dff_A_he3bOx2Q8_2(.dout(w_dff_A_OXGOCku81_2),.din(w_dff_A_he3bOx2Q8_2),.clk(gclk));
	jdff dff_A_vSTRQghL4_2(.dout(w_dff_A_he3bOx2Q8_2),.din(w_dff_A_vSTRQghL4_2),.clk(gclk));
	jdff dff_A_Kv3cKQwf0_2(.dout(w_dff_A_vSTRQghL4_2),.din(w_dff_A_Kv3cKQwf0_2),.clk(gclk));
	jdff dff_A_qKsaUKEO2_2(.dout(w_dff_A_Kv3cKQwf0_2),.din(w_dff_A_qKsaUKEO2_2),.clk(gclk));
	jdff dff_A_eDAwHI2u4_2(.dout(w_dff_A_qKsaUKEO2_2),.din(w_dff_A_eDAwHI2u4_2),.clk(gclk));
	jdff dff_A_P8UycJDD8_2(.dout(w_dff_A_eDAwHI2u4_2),.din(w_dff_A_P8UycJDD8_2),.clk(gclk));
	jdff dff_A_QxwvuVAj4_2(.dout(w_dff_A_P8UycJDD8_2),.din(w_dff_A_QxwvuVAj4_2),.clk(gclk));
	jdff dff_A_rNFC4wfo5_2(.dout(w_dff_A_QxwvuVAj4_2),.din(w_dff_A_rNFC4wfo5_2),.clk(gclk));
	jdff dff_A_kcw9hboA7_2(.dout(w_dff_A_rNFC4wfo5_2),.din(w_dff_A_kcw9hboA7_2),.clk(gclk));
	jdff dff_A_RJWpgXXD6_2(.dout(w_dff_A_kcw9hboA7_2),.din(w_dff_A_RJWpgXXD6_2),.clk(gclk));
	jdff dff_B_Tx3nH3oS8_0(.din(n1324),.dout(w_dff_B_Tx3nH3oS8_0),.clk(gclk));
	jdff dff_B_hgGxcLaZ2_0(.din(w_dff_B_Tx3nH3oS8_0),.dout(w_dff_B_hgGxcLaZ2_0),.clk(gclk));
	jdff dff_B_mbycB4hs9_0(.din(w_dff_B_hgGxcLaZ2_0),.dout(w_dff_B_mbycB4hs9_0),.clk(gclk));
	jdff dff_B_idaAs0Bw9_0(.din(w_dff_B_mbycB4hs9_0),.dout(w_dff_B_idaAs0Bw9_0),.clk(gclk));
	jdff dff_B_XzBlgQAC4_0(.din(w_dff_B_idaAs0Bw9_0),.dout(w_dff_B_XzBlgQAC4_0),.clk(gclk));
	jdff dff_B_Q6RuIBFz3_0(.din(w_dff_B_XzBlgQAC4_0),.dout(w_dff_B_Q6RuIBFz3_0),.clk(gclk));
	jdff dff_B_Q7Atw7ZZ3_0(.din(w_dff_B_Q6RuIBFz3_0),.dout(w_dff_B_Q7Atw7ZZ3_0),.clk(gclk));
	jdff dff_B_da2HRq8B2_0(.din(w_dff_B_Q7Atw7ZZ3_0),.dout(w_dff_B_da2HRq8B2_0),.clk(gclk));
	jdff dff_B_Y1Z1LecR4_0(.din(w_dff_B_da2HRq8B2_0),.dout(w_dff_B_Y1Z1LecR4_0),.clk(gclk));
	jdff dff_B_ijvYExa02_0(.din(w_dff_B_Y1Z1LecR4_0),.dout(w_dff_B_ijvYExa02_0),.clk(gclk));
	jdff dff_B_dsWROEKM4_0(.din(w_dff_B_ijvYExa02_0),.dout(w_dff_B_dsWROEKM4_0),.clk(gclk));
	jdff dff_B_AYDWcRqT7_0(.din(w_dff_B_dsWROEKM4_0),.dout(w_dff_B_AYDWcRqT7_0),.clk(gclk));
	jdff dff_B_fegGlux16_0(.din(w_dff_B_AYDWcRqT7_0),.dout(w_dff_B_fegGlux16_0),.clk(gclk));
	jdff dff_B_bLveDmSc6_0(.din(w_dff_B_fegGlux16_0),.dout(w_dff_B_bLveDmSc6_0),.clk(gclk));
	jdff dff_B_F7XzmOPd8_0(.din(w_dff_B_bLveDmSc6_0),.dout(w_dff_B_F7XzmOPd8_0),.clk(gclk));
	jdff dff_B_F3T0l02s7_0(.din(w_dff_B_F7XzmOPd8_0),.dout(w_dff_B_F3T0l02s7_0),.clk(gclk));
	jdff dff_B_Xtb5aoXD7_0(.din(w_dff_B_F3T0l02s7_0),.dout(w_dff_B_Xtb5aoXD7_0),.clk(gclk));
	jdff dff_B_4VDLMkRI1_0(.din(w_dff_B_Xtb5aoXD7_0),.dout(w_dff_B_4VDLMkRI1_0),.clk(gclk));
	jdff dff_B_ESMV3WSY4_0(.din(w_dff_B_4VDLMkRI1_0),.dout(w_dff_B_ESMV3WSY4_0),.clk(gclk));
	jdff dff_B_GRzCDFLx2_0(.din(w_dff_B_ESMV3WSY4_0),.dout(w_dff_B_GRzCDFLx2_0),.clk(gclk));
	jdff dff_A_RHULBzFo7_2(.dout(w_G4090_2[2]),.din(w_dff_A_RHULBzFo7_2),.clk(gclk));
	jdff dff_B_uaO0d8MK4_2(.din(G103),.dout(w_dff_B_uaO0d8MK4_2),.clk(gclk));
	jdff dff_B_T1W1r0Mi2_1(.din(n1317),.dout(w_dff_B_T1W1r0Mi2_1),.clk(gclk));
	jdff dff_B_hdS1Xd212_0(.din(n1333),.dout(w_dff_B_hdS1Xd212_0),.clk(gclk));
	jdff dff_B_qh3ZIsU17_0(.din(w_dff_B_hdS1Xd212_0),.dout(w_dff_B_qh3ZIsU17_0),.clk(gclk));
	jdff dff_B_pnffsTc89_0(.din(w_dff_B_qh3ZIsU17_0),.dout(w_dff_B_pnffsTc89_0),.clk(gclk));
	jdff dff_B_Y2FFdj650_0(.din(w_dff_B_pnffsTc89_0),.dout(w_dff_B_Y2FFdj650_0),.clk(gclk));
	jdff dff_B_PCe4hWqu0_0(.din(w_dff_B_Y2FFdj650_0),.dout(w_dff_B_PCe4hWqu0_0),.clk(gclk));
	jdff dff_B_iIdX5ytB4_0(.din(w_dff_B_PCe4hWqu0_0),.dout(w_dff_B_iIdX5ytB4_0),.clk(gclk));
	jdff dff_B_8ru6XpIH6_0(.din(w_dff_B_iIdX5ytB4_0),.dout(w_dff_B_8ru6XpIH6_0),.clk(gclk));
	jdff dff_B_o7zdvJmS4_0(.din(w_dff_B_8ru6XpIH6_0),.dout(w_dff_B_o7zdvJmS4_0),.clk(gclk));
	jdff dff_B_jSKjCHVl7_0(.din(w_dff_B_o7zdvJmS4_0),.dout(w_dff_B_jSKjCHVl7_0),.clk(gclk));
	jdff dff_B_IPorO2iJ9_0(.din(w_dff_B_jSKjCHVl7_0),.dout(w_dff_B_IPorO2iJ9_0),.clk(gclk));
	jdff dff_B_wiAzWvOK8_0(.din(w_dff_B_IPorO2iJ9_0),.dout(w_dff_B_wiAzWvOK8_0),.clk(gclk));
	jdff dff_B_59pWEpqM0_0(.din(w_dff_B_wiAzWvOK8_0),.dout(w_dff_B_59pWEpqM0_0),.clk(gclk));
	jdff dff_B_0NrHRDnN8_0(.din(w_dff_B_59pWEpqM0_0),.dout(w_dff_B_0NrHRDnN8_0),.clk(gclk));
	jdff dff_B_z5Yeu1YP3_0(.din(w_dff_B_0NrHRDnN8_0),.dout(w_dff_B_z5Yeu1YP3_0),.clk(gclk));
	jdff dff_B_2RxG98qb5_0(.din(w_dff_B_z5Yeu1YP3_0),.dout(w_dff_B_2RxG98qb5_0),.clk(gclk));
	jdff dff_B_evBNwruV0_0(.din(w_dff_B_2RxG98qb5_0),.dout(w_dff_B_evBNwruV0_0),.clk(gclk));
	jdff dff_B_LO9JOhnI8_0(.din(w_dff_B_evBNwruV0_0),.dout(w_dff_B_LO9JOhnI8_0),.clk(gclk));
	jdff dff_B_LqHYB27G5_0(.din(w_dff_B_LO9JOhnI8_0),.dout(w_dff_B_LqHYB27G5_0),.clk(gclk));
	jdff dff_B_tCYsu0WS0_0(.din(w_dff_B_LqHYB27G5_0),.dout(w_dff_B_tCYsu0WS0_0),.clk(gclk));
	jdff dff_B_YnmLANBf9_2(.din(G40),.dout(w_dff_B_YnmLANBf9_2),.clk(gclk));
	jdff dff_B_WKybI4lD9_1(.din(n1326),.dout(w_dff_B_WKybI4lD9_1),.clk(gclk));
	jdff dff_B_Nt5hPK6m3_1(.din(w_dff_B_WKybI4lD9_1),.dout(w_dff_B_Nt5hPK6m3_1),.clk(gclk));
	jdff dff_B_C4l1m0gX6_1(.din(w_dff_B_Nt5hPK6m3_1),.dout(w_dff_B_C4l1m0gX6_1),.clk(gclk));
	jdff dff_A_vnhR8o3d4_0(.dout(w_n852_4[0]),.din(w_dff_A_vnhR8o3d4_0),.clk(gclk));
	jdff dff_A_GEU44v5Q4_0(.dout(w_dff_A_vnhR8o3d4_0),.din(w_dff_A_GEU44v5Q4_0),.clk(gclk));
	jdff dff_A_wfZ8ZsLa1_0(.dout(w_dff_A_GEU44v5Q4_0),.din(w_dff_A_wfZ8ZsLa1_0),.clk(gclk));
	jdff dff_A_F5aYLFnV1_0(.dout(w_dff_A_wfZ8ZsLa1_0),.din(w_dff_A_F5aYLFnV1_0),.clk(gclk));
	jdff dff_A_tmBuKDQV3_0(.dout(w_dff_A_F5aYLFnV1_0),.din(w_dff_A_tmBuKDQV3_0),.clk(gclk));
	jdff dff_A_vLkJbTwn0_0(.dout(w_dff_A_tmBuKDQV3_0),.din(w_dff_A_vLkJbTwn0_0),.clk(gclk));
	jdff dff_A_1WgpBUtp3_0(.dout(w_dff_A_vLkJbTwn0_0),.din(w_dff_A_1WgpBUtp3_0),.clk(gclk));
	jdff dff_A_ilK3GIH75_0(.dout(w_dff_A_1WgpBUtp3_0),.din(w_dff_A_ilK3GIH75_0),.clk(gclk));
	jdff dff_A_Emgmwmvm8_0(.dout(w_dff_A_ilK3GIH75_0),.din(w_dff_A_Emgmwmvm8_0),.clk(gclk));
	jdff dff_A_MfPtqWRG0_0(.dout(w_dff_A_Emgmwmvm8_0),.din(w_dff_A_MfPtqWRG0_0),.clk(gclk));
	jdff dff_A_R9fmyxep8_0(.dout(w_dff_A_MfPtqWRG0_0),.din(w_dff_A_R9fmyxep8_0),.clk(gclk));
	jdff dff_A_7wRx7xaG3_0(.dout(w_dff_A_R9fmyxep8_0),.din(w_dff_A_7wRx7xaG3_0),.clk(gclk));
	jdff dff_A_cHzaRFDO4_0(.dout(w_dff_A_7wRx7xaG3_0),.din(w_dff_A_cHzaRFDO4_0),.clk(gclk));
	jdff dff_A_G4Xxnea55_0(.dout(w_dff_A_cHzaRFDO4_0),.din(w_dff_A_G4Xxnea55_0),.clk(gclk));
	jdff dff_A_MvsB6TA38_0(.dout(w_dff_A_G4Xxnea55_0),.din(w_dff_A_MvsB6TA38_0),.clk(gclk));
	jdff dff_A_iA2VBYc17_0(.dout(w_dff_A_MvsB6TA38_0),.din(w_dff_A_iA2VBYc17_0),.clk(gclk));
	jdff dff_A_GgQ1ID3J5_0(.dout(w_dff_A_iA2VBYc17_0),.din(w_dff_A_GgQ1ID3J5_0),.clk(gclk));
	jdff dff_A_bNh4M6Ep2_0(.dout(w_dff_A_GgQ1ID3J5_0),.din(w_dff_A_bNh4M6Ep2_0),.clk(gclk));
	jdff dff_A_TJygGqzl7_2(.dout(w_n852_4[2]),.din(w_dff_A_TJygGqzl7_2),.clk(gclk));
	jdff dff_A_iU15CS426_2(.dout(w_dff_A_TJygGqzl7_2),.din(w_dff_A_iU15CS426_2),.clk(gclk));
	jdff dff_A_dpzeTCi89_2(.dout(w_dff_A_iU15CS426_2),.din(w_dff_A_dpzeTCi89_2),.clk(gclk));
	jdff dff_A_yQgaYmtb1_2(.dout(w_dff_A_dpzeTCi89_2),.din(w_dff_A_yQgaYmtb1_2),.clk(gclk));
	jdff dff_A_cfEQ7Qna0_2(.dout(w_dff_A_yQgaYmtb1_2),.din(w_dff_A_cfEQ7Qna0_2),.clk(gclk));
	jdff dff_A_E56k601s3_2(.dout(w_dff_A_cfEQ7Qna0_2),.din(w_dff_A_E56k601s3_2),.clk(gclk));
	jdff dff_A_jio8YAFG7_2(.dout(w_dff_A_E56k601s3_2),.din(w_dff_A_jio8YAFG7_2),.clk(gclk));
	jdff dff_A_PZrhnLXL2_2(.dout(w_dff_A_jio8YAFG7_2),.din(w_dff_A_PZrhnLXL2_2),.clk(gclk));
	jdff dff_A_jxw9vpws8_2(.dout(w_dff_A_PZrhnLXL2_2),.din(w_dff_A_jxw9vpws8_2),.clk(gclk));
	jdff dff_A_cJft473K6_2(.dout(w_dff_A_jxw9vpws8_2),.din(w_dff_A_cJft473K6_2),.clk(gclk));
	jdff dff_A_7PRmW6Ip6_2(.dout(w_dff_A_cJft473K6_2),.din(w_dff_A_7PRmW6Ip6_2),.clk(gclk));
	jdff dff_A_v5VCptiH7_2(.dout(w_dff_A_7PRmW6Ip6_2),.din(w_dff_A_v5VCptiH7_2),.clk(gclk));
	jdff dff_A_O40I5Xo73_2(.dout(w_dff_A_v5VCptiH7_2),.din(w_dff_A_O40I5Xo73_2),.clk(gclk));
	jdff dff_A_lsbdGSYB5_2(.dout(w_dff_A_O40I5Xo73_2),.din(w_dff_A_lsbdGSYB5_2),.clk(gclk));
	jdff dff_A_VAJHHmLj1_2(.dout(w_dff_A_lsbdGSYB5_2),.din(w_dff_A_VAJHHmLj1_2),.clk(gclk));
	jdff dff_A_KKh4rwpx4_2(.dout(w_dff_A_VAJHHmLj1_2),.din(w_dff_A_KKh4rwpx4_2),.clk(gclk));
	jdff dff_A_HFgvA4HM3_2(.dout(w_dff_A_KKh4rwpx4_2),.din(w_dff_A_HFgvA4HM3_2),.clk(gclk));
	jdff dff_A_IPJr4FrX8_2(.dout(w_dff_A_HFgvA4HM3_2),.din(w_dff_A_IPJr4FrX8_2),.clk(gclk));
	jdff dff_A_FHS91h1n8_2(.dout(w_dff_A_IPJr4FrX8_2),.din(w_dff_A_FHS91h1n8_2),.clk(gclk));
	jdff dff_A_HSz7qNpi9_0(.dout(w_G4089_4[0]),.din(w_dff_A_HSz7qNpi9_0),.clk(gclk));
	jdff dff_A_viGMn3QI9_0(.dout(w_dff_A_HSz7qNpi9_0),.din(w_dff_A_viGMn3QI9_0),.clk(gclk));
	jdff dff_A_5uhSE4tk9_0(.dout(w_dff_A_viGMn3QI9_0),.din(w_dff_A_5uhSE4tk9_0),.clk(gclk));
	jdff dff_A_yD8WmPpv2_0(.dout(w_dff_A_5uhSE4tk9_0),.din(w_dff_A_yD8WmPpv2_0),.clk(gclk));
	jdff dff_A_pFbS3kbv3_0(.dout(w_dff_A_yD8WmPpv2_0),.din(w_dff_A_pFbS3kbv3_0),.clk(gclk));
	jdff dff_A_eSWenga86_0(.dout(w_dff_A_pFbS3kbv3_0),.din(w_dff_A_eSWenga86_0),.clk(gclk));
	jdff dff_A_K2qJq7z68_0(.dout(w_dff_A_eSWenga86_0),.din(w_dff_A_K2qJq7z68_0),.clk(gclk));
	jdff dff_A_JJWtZTpV4_0(.dout(w_dff_A_K2qJq7z68_0),.din(w_dff_A_JJWtZTpV4_0),.clk(gclk));
	jdff dff_A_yc4fj2JV3_0(.dout(w_dff_A_JJWtZTpV4_0),.din(w_dff_A_yc4fj2JV3_0),.clk(gclk));
	jdff dff_A_RRimMF1z8_0(.dout(w_dff_A_yc4fj2JV3_0),.din(w_dff_A_RRimMF1z8_0),.clk(gclk));
	jdff dff_A_g6rtoMU50_0(.dout(w_dff_A_RRimMF1z8_0),.din(w_dff_A_g6rtoMU50_0),.clk(gclk));
	jdff dff_A_NM2AqfPu2_0(.dout(w_dff_A_g6rtoMU50_0),.din(w_dff_A_NM2AqfPu2_0),.clk(gclk));
	jdff dff_A_IhdNb4sX1_0(.dout(w_dff_A_NM2AqfPu2_0),.din(w_dff_A_IhdNb4sX1_0),.clk(gclk));
	jdff dff_A_lpLbDs6F4_0(.dout(w_dff_A_IhdNb4sX1_0),.din(w_dff_A_lpLbDs6F4_0),.clk(gclk));
	jdff dff_A_2neD71Vj8_0(.dout(w_dff_A_lpLbDs6F4_0),.din(w_dff_A_2neD71Vj8_0),.clk(gclk));
	jdff dff_A_y72R2Axt7_0(.dout(w_dff_A_2neD71Vj8_0),.din(w_dff_A_y72R2Axt7_0),.clk(gclk));
	jdff dff_A_Hzdn82JJ8_0(.dout(w_dff_A_y72R2Axt7_0),.din(w_dff_A_Hzdn82JJ8_0),.clk(gclk));
	jdff dff_A_a1Ck1LAN9_2(.dout(w_G4089_4[2]),.din(w_dff_A_a1Ck1LAN9_2),.clk(gclk));
	jdff dff_A_O6xluIb36_2(.dout(w_dff_A_a1Ck1LAN9_2),.din(w_dff_A_O6xluIb36_2),.clk(gclk));
	jdff dff_A_GiiiFa3n3_2(.dout(w_dff_A_O6xluIb36_2),.din(w_dff_A_GiiiFa3n3_2),.clk(gclk));
	jdff dff_A_rAuThIDR2_2(.dout(w_dff_A_GiiiFa3n3_2),.din(w_dff_A_rAuThIDR2_2),.clk(gclk));
	jdff dff_A_DHgXbhto7_2(.dout(w_dff_A_rAuThIDR2_2),.din(w_dff_A_DHgXbhto7_2),.clk(gclk));
	jdff dff_A_7XYq4DsJ4_2(.dout(w_dff_A_DHgXbhto7_2),.din(w_dff_A_7XYq4DsJ4_2),.clk(gclk));
	jdff dff_A_K5jHEDma0_2(.dout(w_dff_A_7XYq4DsJ4_2),.din(w_dff_A_K5jHEDma0_2),.clk(gclk));
	jdff dff_A_496LZMLI8_2(.dout(w_dff_A_K5jHEDma0_2),.din(w_dff_A_496LZMLI8_2),.clk(gclk));
	jdff dff_A_pYJCONra7_2(.dout(w_dff_A_496LZMLI8_2),.din(w_dff_A_pYJCONra7_2),.clk(gclk));
	jdff dff_A_FyPPEUMn5_2(.dout(w_dff_A_pYJCONra7_2),.din(w_dff_A_FyPPEUMn5_2),.clk(gclk));
	jdff dff_A_Qtz8xAoZ2_2(.dout(w_dff_A_FyPPEUMn5_2),.din(w_dff_A_Qtz8xAoZ2_2),.clk(gclk));
	jdff dff_A_d4lzdykj4_2(.dout(w_dff_A_Qtz8xAoZ2_2),.din(w_dff_A_d4lzdykj4_2),.clk(gclk));
	jdff dff_A_KXSTPiPM8_2(.dout(w_dff_A_d4lzdykj4_2),.din(w_dff_A_KXSTPiPM8_2),.clk(gclk));
	jdff dff_A_ncMREv2P8_2(.dout(w_dff_A_KXSTPiPM8_2),.din(w_dff_A_ncMREv2P8_2),.clk(gclk));
	jdff dff_A_1dAyC3bT0_2(.dout(w_dff_A_ncMREv2P8_2),.din(w_dff_A_1dAyC3bT0_2),.clk(gclk));
	jdff dff_A_woZw5Kyi8_2(.dout(w_dff_A_1dAyC3bT0_2),.din(w_dff_A_woZw5Kyi8_2),.clk(gclk));
	jdff dff_A_4uPCxWrf1_2(.dout(w_dff_A_woZw5Kyi8_2),.din(w_dff_A_4uPCxWrf1_2),.clk(gclk));
	jdff dff_A_uif6g65M9_2(.dout(w_dff_A_4uPCxWrf1_2),.din(w_dff_A_uif6g65M9_2),.clk(gclk));
	jdff dff_A_XOZcIZ1n5_2(.dout(w_dff_A_uif6g65M9_2),.din(w_dff_A_XOZcIZ1n5_2),.clk(gclk));
	jdff dff_A_8Qwl9bBz2_2(.dout(w_dff_A_XOZcIZ1n5_2),.din(w_dff_A_8Qwl9bBz2_2),.clk(gclk));
	jdff dff_B_yYB6TAZo9_0(.din(n1341),.dout(w_dff_B_yYB6TAZo9_0),.clk(gclk));
	jdff dff_B_N9rGxIIx6_0(.din(w_dff_B_yYB6TAZo9_0),.dout(w_dff_B_N9rGxIIx6_0),.clk(gclk));
	jdff dff_B_Arf4ptQS9_0(.din(w_dff_B_N9rGxIIx6_0),.dout(w_dff_B_Arf4ptQS9_0),.clk(gclk));
	jdff dff_B_LT7gTv8j4_0(.din(w_dff_B_Arf4ptQS9_0),.dout(w_dff_B_LT7gTv8j4_0),.clk(gclk));
	jdff dff_B_PPi1ZdXw9_0(.din(w_dff_B_LT7gTv8j4_0),.dout(w_dff_B_PPi1ZdXw9_0),.clk(gclk));
	jdff dff_B_1zYuoSQ24_0(.din(w_dff_B_PPi1ZdXw9_0),.dout(w_dff_B_1zYuoSQ24_0),.clk(gclk));
	jdff dff_B_9ZxP1CpH4_0(.din(w_dff_B_1zYuoSQ24_0),.dout(w_dff_B_9ZxP1CpH4_0),.clk(gclk));
	jdff dff_B_dYNfhZ5W5_0(.din(w_dff_B_9ZxP1CpH4_0),.dout(w_dff_B_dYNfhZ5W5_0),.clk(gclk));
	jdff dff_B_8Ouoy7LE7_0(.din(w_dff_B_dYNfhZ5W5_0),.dout(w_dff_B_8Ouoy7LE7_0),.clk(gclk));
	jdff dff_B_15p2zQ3u1_0(.din(w_dff_B_8Ouoy7LE7_0),.dout(w_dff_B_15p2zQ3u1_0),.clk(gclk));
	jdff dff_B_sPD79SSp3_0(.din(w_dff_B_15p2zQ3u1_0),.dout(w_dff_B_sPD79SSp3_0),.clk(gclk));
	jdff dff_B_THVAymhP4_0(.din(w_dff_B_sPD79SSp3_0),.dout(w_dff_B_THVAymhP4_0),.clk(gclk));
	jdff dff_B_h3nGbSLd0_0(.din(w_dff_B_THVAymhP4_0),.dout(w_dff_B_h3nGbSLd0_0),.clk(gclk));
	jdff dff_B_MLpbz2IM5_0(.din(w_dff_B_h3nGbSLd0_0),.dout(w_dff_B_MLpbz2IM5_0),.clk(gclk));
	jdff dff_B_e4BKR3X65_0(.din(w_dff_B_MLpbz2IM5_0),.dout(w_dff_B_e4BKR3X65_0),.clk(gclk));
	jdff dff_B_YKawyxsP8_0(.din(w_dff_B_e4BKR3X65_0),.dout(w_dff_B_YKawyxsP8_0),.clk(gclk));
	jdff dff_B_ylHZqwYG2_0(.din(w_dff_B_YKawyxsP8_0),.dout(w_dff_B_ylHZqwYG2_0),.clk(gclk));
	jdff dff_B_o3U269by6_0(.din(w_dff_B_ylHZqwYG2_0),.dout(w_dff_B_o3U269by6_0),.clk(gclk));
	jdff dff_B_o2lYWXg34_0(.din(n1340),.dout(w_dff_B_o2lYWXg34_0),.clk(gclk));
	jdff dff_B_QTf9ErPX5_1(.din(n1335),.dout(w_dff_B_QTf9ErPX5_1),.clk(gclk));
	jdff dff_B_oWAW81qD6_1(.din(w_dff_B_QTf9ErPX5_1),.dout(w_dff_B_oWAW81qD6_1),.clk(gclk));
	jdff dff_B_oMESUjmC8_1(.din(w_dff_B_oWAW81qD6_1),.dout(w_dff_B_oMESUjmC8_1),.clk(gclk));
	jdff dff_A_3K5qGB1N1_0(.dout(w_n999_2[0]),.din(w_dff_A_3K5qGB1N1_0),.clk(gclk));
	jdff dff_A_95xPttmD4_0(.dout(w_dff_A_3K5qGB1N1_0),.din(w_dff_A_95xPttmD4_0),.clk(gclk));
	jdff dff_A_Di47PCmo2_0(.dout(w_dff_A_95xPttmD4_0),.din(w_dff_A_Di47PCmo2_0),.clk(gclk));
	jdff dff_A_GB3lom5E6_0(.dout(w_dff_A_Di47PCmo2_0),.din(w_dff_A_GB3lom5E6_0),.clk(gclk));
	jdff dff_A_PKL4Ihwc6_0(.dout(w_dff_A_GB3lom5E6_0),.din(w_dff_A_PKL4Ihwc6_0),.clk(gclk));
	jdff dff_A_VOAFHszn5_0(.dout(w_dff_A_PKL4Ihwc6_0),.din(w_dff_A_VOAFHszn5_0),.clk(gclk));
	jdff dff_A_APFbucbk9_1(.dout(w_n999_2[1]),.din(w_dff_A_APFbucbk9_1),.clk(gclk));
	jdff dff_A_tXUoP4lF0_0(.dout(w_G1689_3[0]),.din(w_dff_A_tXUoP4lF0_0),.clk(gclk));
	jdff dff_A_Aw6lNMMU4_0(.dout(w_dff_A_tXUoP4lF0_0),.din(w_dff_A_Aw6lNMMU4_0),.clk(gclk));
	jdff dff_A_z9ivnzQ28_0(.dout(w_dff_A_Aw6lNMMU4_0),.din(w_dff_A_z9ivnzQ28_0),.clk(gclk));
	jdff dff_A_wAZAh3OW7_0(.dout(w_dff_A_z9ivnzQ28_0),.din(w_dff_A_wAZAh3OW7_0),.clk(gclk));
	jdff dff_A_VYfevSgU1_1(.dout(w_G1689_3[1]),.din(w_dff_A_VYfevSgU1_1),.clk(gclk));
	jdff dff_A_IdOvsTrc2_1(.dout(w_dff_A_VYfevSgU1_1),.din(w_dff_A_IdOvsTrc2_1),.clk(gclk));
	jdff dff_A_2k6ktBTe1_0(.dout(w_G137_6[0]),.din(w_dff_A_2k6ktBTe1_0),.clk(gclk));
	jdff dff_A_zT7UaD024_0(.dout(w_dff_A_2k6ktBTe1_0),.din(w_dff_A_zT7UaD024_0),.clk(gclk));
	jdff dff_A_hra1La5V3_0(.dout(w_dff_A_zT7UaD024_0),.din(w_dff_A_hra1La5V3_0),.clk(gclk));
	jdff dff_A_uC2OrI8W5_0(.dout(w_dff_A_hra1La5V3_0),.din(w_dff_A_uC2OrI8W5_0),.clk(gclk));
	jdff dff_A_Ho32hBRl7_0(.dout(w_dff_A_uC2OrI8W5_0),.din(w_dff_A_Ho32hBRl7_0),.clk(gclk));
	jdff dff_A_wEzRSUOx8_0(.dout(w_dff_A_Ho32hBRl7_0),.din(w_dff_A_wEzRSUOx8_0),.clk(gclk));
	jdff dff_A_9uvh0oUf1_1(.dout(w_G137_6[1]),.din(w_dff_A_9uvh0oUf1_1),.clk(gclk));
	jdff dff_B_Qjq07H452_0(.din(n1350),.dout(w_dff_B_Qjq07H452_0),.clk(gclk));
	jdff dff_B_Ijvwahbm8_0(.din(w_dff_B_Qjq07H452_0),.dout(w_dff_B_Ijvwahbm8_0),.clk(gclk));
	jdff dff_B_U1WfJBmg3_0(.din(w_dff_B_Ijvwahbm8_0),.dout(w_dff_B_U1WfJBmg3_0),.clk(gclk));
	jdff dff_B_npXesAWe5_0(.din(w_dff_B_U1WfJBmg3_0),.dout(w_dff_B_npXesAWe5_0),.clk(gclk));
	jdff dff_B_Zv8jywsV7_0(.din(w_dff_B_npXesAWe5_0),.dout(w_dff_B_Zv8jywsV7_0),.clk(gclk));
	jdff dff_B_RVc9EPDD6_0(.din(w_dff_B_Zv8jywsV7_0),.dout(w_dff_B_RVc9EPDD6_0),.clk(gclk));
	jdff dff_B_F2soZxR53_0(.din(w_dff_B_RVc9EPDD6_0),.dout(w_dff_B_F2soZxR53_0),.clk(gclk));
	jdff dff_B_6hvB721S8_0(.din(w_dff_B_F2soZxR53_0),.dout(w_dff_B_6hvB721S8_0),.clk(gclk));
	jdff dff_B_lBoNCdOZ8_0(.din(w_dff_B_6hvB721S8_0),.dout(w_dff_B_lBoNCdOZ8_0),.clk(gclk));
	jdff dff_B_9lUh3Cp42_0(.din(w_dff_B_lBoNCdOZ8_0),.dout(w_dff_B_9lUh3Cp42_0),.clk(gclk));
	jdff dff_B_WSczm8ck7_0(.din(w_dff_B_9lUh3Cp42_0),.dout(w_dff_B_WSczm8ck7_0),.clk(gclk));
	jdff dff_B_xbporivq5_0(.din(w_dff_B_WSczm8ck7_0),.dout(w_dff_B_xbporivq5_0),.clk(gclk));
	jdff dff_B_1DElu1if2_0(.din(w_dff_B_xbporivq5_0),.dout(w_dff_B_1DElu1if2_0),.clk(gclk));
	jdff dff_B_yu3bNiHn0_0(.din(w_dff_B_1DElu1if2_0),.dout(w_dff_B_yu3bNiHn0_0),.clk(gclk));
	jdff dff_B_w0Eo8hmv1_0(.din(w_dff_B_yu3bNiHn0_0),.dout(w_dff_B_w0Eo8hmv1_0),.clk(gclk));
	jdff dff_B_eZzwnoab4_0(.din(w_dff_B_w0Eo8hmv1_0),.dout(w_dff_B_eZzwnoab4_0),.clk(gclk));
	jdff dff_B_myS6yNBK6_0(.din(w_dff_B_eZzwnoab4_0),.dout(w_dff_B_myS6yNBK6_0),.clk(gclk));
	jdff dff_B_v9gZSm0M9_0(.din(w_dff_B_myS6yNBK6_0),.dout(w_dff_B_v9gZSm0M9_0),.clk(gclk));
	jdff dff_B_k8e4oTpX8_0(.din(w_dff_B_v9gZSm0M9_0),.dout(w_dff_B_k8e4oTpX8_0),.clk(gclk));
	jdff dff_B_YFV8slcf0_0(.din(n1349),.dout(w_dff_B_YFV8slcf0_0),.clk(gclk));
	jdff dff_B_WtmtCWCJ1_1(.din(n1344),.dout(w_dff_B_WtmtCWCJ1_1),.clk(gclk));
	jdff dff_B_lXMbRhuD4_1(.din(n1355),.dout(w_dff_B_lXMbRhuD4_1),.clk(gclk));
	jdff dff_B_HY13YXOs5_1(.din(w_dff_B_lXMbRhuD4_1),.dout(w_dff_B_HY13YXOs5_1),.clk(gclk));
	jdff dff_B_FonaWKoP9_1(.din(w_dff_B_HY13YXOs5_1),.dout(w_dff_B_FonaWKoP9_1),.clk(gclk));
	jdff dff_B_i6hooBBx6_1(.din(w_dff_B_FonaWKoP9_1),.dout(w_dff_B_i6hooBBx6_1),.clk(gclk));
	jdff dff_B_pPnBGupb1_1(.din(w_dff_B_i6hooBBx6_1),.dout(w_dff_B_pPnBGupb1_1),.clk(gclk));
	jdff dff_B_r4f2I6v88_1(.din(w_dff_B_pPnBGupb1_1),.dout(w_dff_B_r4f2I6v88_1),.clk(gclk));
	jdff dff_B_o77agAi46_1(.din(w_dff_B_r4f2I6v88_1),.dout(w_dff_B_o77agAi46_1),.clk(gclk));
	jdff dff_B_5ZIGr0MD4_1(.din(w_dff_B_o77agAi46_1),.dout(w_dff_B_5ZIGr0MD4_1),.clk(gclk));
	jdff dff_B_fug5m2Uz6_1(.din(w_dff_B_5ZIGr0MD4_1),.dout(w_dff_B_fug5m2Uz6_1),.clk(gclk));
	jdff dff_B_PMrZCyXN4_1(.din(w_dff_B_fug5m2Uz6_1),.dout(w_dff_B_PMrZCyXN4_1),.clk(gclk));
	jdff dff_B_h1rIcDDy2_1(.din(w_dff_B_PMrZCyXN4_1),.dout(w_dff_B_h1rIcDDy2_1),.clk(gclk));
	jdff dff_B_cUS0QtHJ5_1(.din(w_dff_B_h1rIcDDy2_1),.dout(w_dff_B_cUS0QtHJ5_1),.clk(gclk));
	jdff dff_B_vT0DQTLX3_1(.din(w_dff_B_cUS0QtHJ5_1),.dout(w_dff_B_vT0DQTLX3_1),.clk(gclk));
	jdff dff_B_4RuFdNRT6_1(.din(w_dff_B_vT0DQTLX3_1),.dout(w_dff_B_4RuFdNRT6_1),.clk(gclk));
	jdff dff_B_OX8ualn71_1(.din(w_dff_B_4RuFdNRT6_1),.dout(w_dff_B_OX8ualn71_1),.clk(gclk));
	jdff dff_B_fKIVnX7K4_1(.din(w_dff_B_OX8ualn71_1),.dout(w_dff_B_fKIVnX7K4_1),.clk(gclk));
	jdff dff_B_m6W3wUY36_1(.din(w_dff_B_fKIVnX7K4_1),.dout(w_dff_B_m6W3wUY36_1),.clk(gclk));
	jdff dff_B_7enCrB7h2_1(.din(w_dff_B_m6W3wUY36_1),.dout(w_dff_B_7enCrB7h2_1),.clk(gclk));
	jdff dff_B_m5sqUrVV8_1(.din(w_dff_B_7enCrB7h2_1),.dout(w_dff_B_m5sqUrVV8_1),.clk(gclk));
	jdff dff_B_ObQwgJC15_1(.din(n1356),.dout(w_dff_B_ObQwgJC15_1),.clk(gclk));
	jdff dff_A_5xdz7XYU7_0(.dout(w_n993_2[0]),.din(w_dff_A_5xdz7XYU7_0),.clk(gclk));
	jdff dff_A_Hpy5MfOc2_1(.dout(w_n993_2[1]),.din(w_dff_A_Hpy5MfOc2_1),.clk(gclk));
	jdff dff_B_Ym1YPgLI8_0(.din(n1354),.dout(w_dff_B_Ym1YPgLI8_0),.clk(gclk));
	jdff dff_B_AtolZT8F9_1(.din(n1364),.dout(w_dff_B_AtolZT8F9_1),.clk(gclk));
	jdff dff_B_pwRJUksx3_1(.din(w_dff_B_AtolZT8F9_1),.dout(w_dff_B_pwRJUksx3_1),.clk(gclk));
	jdff dff_B_8woNUihl2_1(.din(w_dff_B_pwRJUksx3_1),.dout(w_dff_B_8woNUihl2_1),.clk(gclk));
	jdff dff_B_skGCBfp53_1(.din(w_dff_B_8woNUihl2_1),.dout(w_dff_B_skGCBfp53_1),.clk(gclk));
	jdff dff_B_ZRgVQ4vv1_1(.din(w_dff_B_skGCBfp53_1),.dout(w_dff_B_ZRgVQ4vv1_1),.clk(gclk));
	jdff dff_B_JL4i2ARc7_1(.din(w_dff_B_ZRgVQ4vv1_1),.dout(w_dff_B_JL4i2ARc7_1),.clk(gclk));
	jdff dff_B_zbAMYEjV6_1(.din(w_dff_B_JL4i2ARc7_1),.dout(w_dff_B_zbAMYEjV6_1),.clk(gclk));
	jdff dff_B_aHWdyLhU9_1(.din(w_dff_B_zbAMYEjV6_1),.dout(w_dff_B_aHWdyLhU9_1),.clk(gclk));
	jdff dff_B_LWqd3uZb3_1(.din(w_dff_B_aHWdyLhU9_1),.dout(w_dff_B_LWqd3uZb3_1),.clk(gclk));
	jdff dff_B_V6K2BZu84_1(.din(w_dff_B_LWqd3uZb3_1),.dout(w_dff_B_V6K2BZu84_1),.clk(gclk));
	jdff dff_B_16LEHejr9_1(.din(w_dff_B_V6K2BZu84_1),.dout(w_dff_B_16LEHejr9_1),.clk(gclk));
	jdff dff_B_0660sNOs6_1(.din(w_dff_B_16LEHejr9_1),.dout(w_dff_B_0660sNOs6_1),.clk(gclk));
	jdff dff_B_daWiL30p6_1(.din(w_dff_B_0660sNOs6_1),.dout(w_dff_B_daWiL30p6_1),.clk(gclk));
	jdff dff_B_LD59wa0H4_1(.din(w_dff_B_daWiL30p6_1),.dout(w_dff_B_LD59wa0H4_1),.clk(gclk));
	jdff dff_B_RkSYgIEO4_1(.din(w_dff_B_LD59wa0H4_1),.dout(w_dff_B_RkSYgIEO4_1),.clk(gclk));
	jdff dff_B_xxMAb5BD6_1(.din(w_dff_B_RkSYgIEO4_1),.dout(w_dff_B_xxMAb5BD6_1),.clk(gclk));
	jdff dff_B_LBvUITzk2_1(.din(w_dff_B_xxMAb5BD6_1),.dout(w_dff_B_LBvUITzk2_1),.clk(gclk));
	jdff dff_B_gbqBUwIl1_1(.din(w_dff_B_LBvUITzk2_1),.dout(w_dff_B_gbqBUwIl1_1),.clk(gclk));
	jdff dff_B_5ibtmSeG1_1(.din(w_dff_B_gbqBUwIl1_1),.dout(w_dff_B_5ibtmSeG1_1),.clk(gclk));
	jdff dff_B_AZuUwZqn7_1(.din(w_dff_B_5ibtmSeG1_1),.dout(w_dff_B_AZuUwZqn7_1),.clk(gclk));
	jdff dff_B_EWcgwott5_1(.din(n1365),.dout(w_dff_B_EWcgwott5_1),.clk(gclk));
	jdff dff_A_HFPQpTJG5_0(.dout(w_G1689_2[0]),.din(w_dff_A_HFPQpTJG5_0),.clk(gclk));
	jdff dff_A_ppmNuYTf8_2(.dout(w_G1689_2[2]),.din(w_dff_A_ppmNuYTf8_2),.clk(gclk));
	jdff dff_A_eTspS4q13_0(.dout(w_n999_1[0]),.din(w_dff_A_eTspS4q13_0),.clk(gclk));
	jdff dff_A_yDlvjHw96_0(.dout(w_dff_A_eTspS4q13_0),.din(w_dff_A_yDlvjHw96_0),.clk(gclk));
	jdff dff_A_1hELk9MS9_1(.dout(w_n999_1[1]),.din(w_dff_A_1hELk9MS9_1),.clk(gclk));
	jdff dff_A_4nj4cidn5_0(.dout(w_n999_0[0]),.din(w_dff_A_4nj4cidn5_0),.clk(gclk));
	jdff dff_A_76uPv6W69_0(.dout(w_dff_A_4nj4cidn5_0),.din(w_dff_A_76uPv6W69_0),.clk(gclk));
	jdff dff_A_OEPIWn4Y0_0(.dout(w_dff_A_76uPv6W69_0),.din(w_dff_A_OEPIWn4Y0_0),.clk(gclk));
	jdff dff_A_rwowK5U84_0(.dout(w_dff_A_OEPIWn4Y0_0),.din(w_dff_A_rwowK5U84_0),.clk(gclk));
	jdff dff_A_luLEJHA67_0(.dout(w_dff_A_rwowK5U84_0),.din(w_dff_A_luLEJHA67_0),.clk(gclk));
	jdff dff_A_NTrox4ME1_0(.dout(w_dff_A_luLEJHA67_0),.din(w_dff_A_NTrox4ME1_0),.clk(gclk));
	jdff dff_A_oTeowHYw0_0(.dout(w_dff_A_NTrox4ME1_0),.din(w_dff_A_oTeowHYw0_0),.clk(gclk));
	jdff dff_A_XzEB0ILD7_0(.dout(w_dff_A_oTeowHYw0_0),.din(w_dff_A_XzEB0ILD7_0),.clk(gclk));
	jdff dff_A_DL87QF4n7_0(.dout(w_dff_A_XzEB0ILD7_0),.din(w_dff_A_DL87QF4n7_0),.clk(gclk));
	jdff dff_A_c9J82Jq75_0(.dout(w_dff_A_DL87QF4n7_0),.din(w_dff_A_c9J82Jq75_0),.clk(gclk));
	jdff dff_A_VMh60d2x4_0(.dout(w_dff_A_c9J82Jq75_0),.din(w_dff_A_VMh60d2x4_0),.clk(gclk));
	jdff dff_A_yBwxPKn73_1(.dout(w_n999_0[1]),.din(w_dff_A_yBwxPKn73_1),.clk(gclk));
	jdff dff_A_DRZzqlun9_1(.dout(w_dff_A_yBwxPKn73_1),.din(w_dff_A_DRZzqlun9_1),.clk(gclk));
	jdff dff_A_pFQl3gRB8_1(.dout(w_dff_A_DRZzqlun9_1),.din(w_dff_A_pFQl3gRB8_1),.clk(gclk));
	jdff dff_A_eZp5P86f6_1(.dout(w_dff_A_pFQl3gRB8_1),.din(w_dff_A_eZp5P86f6_1),.clk(gclk));
	jdff dff_B_FXNeghKD8_3(.din(n999),.dout(w_dff_B_FXNeghKD8_3),.clk(gclk));
	jdff dff_B_KHVOwOSr1_3(.din(w_dff_B_FXNeghKD8_3),.dout(w_dff_B_KHVOwOSr1_3),.clk(gclk));
	jdff dff_B_B8UBqGIR9_3(.din(w_dff_B_KHVOwOSr1_3),.dout(w_dff_B_B8UBqGIR9_3),.clk(gclk));
	jdff dff_B_6qKQzCyJ9_3(.din(w_dff_B_B8UBqGIR9_3),.dout(w_dff_B_6qKQzCyJ9_3),.clk(gclk));
	jdff dff_B_3aabpeHx6_3(.din(w_dff_B_6qKQzCyJ9_3),.dout(w_dff_B_3aabpeHx6_3),.clk(gclk));
	jdff dff_B_68lGMx9Z2_3(.din(w_dff_B_3aabpeHx6_3),.dout(w_dff_B_68lGMx9Z2_3),.clk(gclk));
	jdff dff_B_7zwlRWqY0_3(.din(w_dff_B_68lGMx9Z2_3),.dout(w_dff_B_7zwlRWqY0_3),.clk(gclk));
	jdff dff_B_VhKtsMnV0_3(.din(w_dff_B_7zwlRWqY0_3),.dout(w_dff_B_VhKtsMnV0_3),.clk(gclk));
	jdff dff_B_XHslf9w03_3(.din(w_dff_B_VhKtsMnV0_3),.dout(w_dff_B_XHslf9w03_3),.clk(gclk));
	jdff dff_B_KcfGaCcD5_0(.din(n1363),.dout(w_dff_B_KcfGaCcD5_0),.clk(gclk));
	jdff dff_A_0vW8M7pl8_0(.dout(w_G137_5[0]),.din(w_dff_A_0vW8M7pl8_0),.clk(gclk));
	jdff dff_B_CRtjkcmB5_0(.din(n1377),.dout(w_dff_B_CRtjkcmB5_0),.clk(gclk));
	jdff dff_B_XD00l3zH0_0(.din(w_dff_B_CRtjkcmB5_0),.dout(w_dff_B_XD00l3zH0_0),.clk(gclk));
	jdff dff_B_qQ5xfVII6_0(.din(w_dff_B_XD00l3zH0_0),.dout(w_dff_B_qQ5xfVII6_0),.clk(gclk));
	jdff dff_B_MOeP6t8y4_0(.din(w_dff_B_qQ5xfVII6_0),.dout(w_dff_B_MOeP6t8y4_0),.clk(gclk));
	jdff dff_B_pN7XJb359_0(.din(w_dff_B_MOeP6t8y4_0),.dout(w_dff_B_pN7XJb359_0),.clk(gclk));
	jdff dff_B_EZtPf5V10_0(.din(w_dff_B_pN7XJb359_0),.dout(w_dff_B_EZtPf5V10_0),.clk(gclk));
	jdff dff_B_6nFsEehQ2_0(.din(w_dff_B_EZtPf5V10_0),.dout(w_dff_B_6nFsEehQ2_0),.clk(gclk));
	jdff dff_B_qsbTU6aX5_0(.din(w_dff_B_6nFsEehQ2_0),.dout(w_dff_B_qsbTU6aX5_0),.clk(gclk));
	jdff dff_B_ZRSVymbL6_0(.din(w_dff_B_qsbTU6aX5_0),.dout(w_dff_B_ZRSVymbL6_0),.clk(gclk));
	jdff dff_B_xFuDborj1_0(.din(w_dff_B_ZRSVymbL6_0),.dout(w_dff_B_xFuDborj1_0),.clk(gclk));
	jdff dff_B_ZP3Ou09r3_0(.din(w_dff_B_xFuDborj1_0),.dout(w_dff_B_ZP3Ou09r3_0),.clk(gclk));
	jdff dff_B_t1GA4otx5_0(.din(w_dff_B_ZP3Ou09r3_0),.dout(w_dff_B_t1GA4otx5_0),.clk(gclk));
	jdff dff_B_TYfR1S6V5_0(.din(w_dff_B_t1GA4otx5_0),.dout(w_dff_B_TYfR1S6V5_0),.clk(gclk));
	jdff dff_B_nOX7kZNc2_0(.din(w_dff_B_TYfR1S6V5_0),.dout(w_dff_B_nOX7kZNc2_0),.clk(gclk));
	jdff dff_B_Lwbztwl10_0(.din(w_dff_B_nOX7kZNc2_0),.dout(w_dff_B_Lwbztwl10_0),.clk(gclk));
	jdff dff_B_F7ipmCq31_0(.din(w_dff_B_Lwbztwl10_0),.dout(w_dff_B_F7ipmCq31_0),.clk(gclk));
	jdff dff_B_bZvC7fT64_0(.din(w_dff_B_F7ipmCq31_0),.dout(w_dff_B_bZvC7fT64_0),.clk(gclk));
	jdff dff_B_XKntAtJb8_0(.din(w_dff_B_bZvC7fT64_0),.dout(w_dff_B_XKntAtJb8_0),.clk(gclk));
	jdff dff_B_ihjrzGeK4_0(.din(n1376),.dout(w_dff_B_ihjrzGeK4_0),.clk(gclk));
	jdff dff_B_hv1i2ayl9_2(.din(G173),.dout(w_dff_B_hv1i2ayl9_2),.clk(gclk));
	jdff dff_B_r4QAimLG6_2(.din(G203),.dout(w_dff_B_r4QAimLG6_2),.clk(gclk));
	jdff dff_B_PZmhi2Ux9_2(.din(w_dff_B_r4QAimLG6_2),.dout(w_dff_B_PZmhi2Ux9_2),.clk(gclk));
	jdff dff_B_tiUFcGwx2_1(.din(n1371),.dout(w_dff_B_tiUFcGwx2_1),.clk(gclk));
	jdff dff_B_5TN3qEZ67_1(.din(w_dff_B_tiUFcGwx2_1),.dout(w_dff_B_5TN3qEZ67_1),.clk(gclk));
	jdff dff_B_6BA4nhSw3_1(.din(w_dff_B_5TN3qEZ67_1),.dout(w_dff_B_6BA4nhSw3_1),.clk(gclk));
	jdff dff_B_BtdO2gts0_1(.din(n1254),.dout(w_dff_B_BtdO2gts0_1),.clk(gclk));
	jdff dff_B_ePHP2b9y8_1(.din(w_dff_B_BtdO2gts0_1),.dout(w_dff_B_ePHP2b9y8_1),.clk(gclk));
	jdff dff_B_fcLVQSPd9_1(.din(w_dff_B_ePHP2b9y8_1),.dout(w_dff_B_fcLVQSPd9_1),.clk(gclk));
	jdff dff_B_EB1jyn2G3_1(.din(w_dff_B_fcLVQSPd9_1),.dout(w_dff_B_EB1jyn2G3_1),.clk(gclk));
	jdff dff_B_SwwdMu4Y8_1(.din(w_dff_B_EB1jyn2G3_1),.dout(w_dff_B_SwwdMu4Y8_1),.clk(gclk));
	jdff dff_B_Y0z90IVy1_1(.din(w_dff_B_SwwdMu4Y8_1),.dout(w_dff_B_Y0z90IVy1_1),.clk(gclk));
	jdff dff_B_6X7uMZkU6_1(.din(w_dff_B_Y0z90IVy1_1),.dout(w_dff_B_6X7uMZkU6_1),.clk(gclk));
	jdff dff_B_Q2EHH6wW5_1(.din(w_dff_B_6X7uMZkU6_1),.dout(w_dff_B_Q2EHH6wW5_1),.clk(gclk));
	jdff dff_B_GyAtbnbc1_1(.din(w_dff_B_Q2EHH6wW5_1),.dout(w_dff_B_GyAtbnbc1_1),.clk(gclk));
	jdff dff_B_uBwPSrnu7_1(.din(w_dff_B_GyAtbnbc1_1),.dout(w_dff_B_uBwPSrnu7_1),.clk(gclk));
	jdff dff_B_nszbMZii6_1(.din(w_dff_B_uBwPSrnu7_1),.dout(w_dff_B_nszbMZii6_1),.clk(gclk));
	jdff dff_B_kOvO2zm75_1(.din(w_dff_B_nszbMZii6_1),.dout(w_dff_B_kOvO2zm75_1),.clk(gclk));
	jdff dff_B_7ZKBsrZl6_1(.din(w_dff_B_kOvO2zm75_1),.dout(w_dff_B_7ZKBsrZl6_1),.clk(gclk));
	jdff dff_B_lMTC9uL96_0(.din(n1257),.dout(w_dff_B_lMTC9uL96_0),.clk(gclk));
	jdff dff_B_NaHG9NqN9_0(.din(w_dff_B_lMTC9uL96_0),.dout(w_dff_B_NaHG9NqN9_0),.clk(gclk));
	jdff dff_B_ePknq90s6_0(.din(w_dff_B_NaHG9NqN9_0),.dout(w_dff_B_ePknq90s6_0),.clk(gclk));
	jdff dff_B_9zm5aosW8_0(.din(w_dff_B_ePknq90s6_0),.dout(w_dff_B_9zm5aosW8_0),.clk(gclk));
	jdff dff_B_K9NaHNCa3_0(.din(w_dff_B_9zm5aosW8_0),.dout(w_dff_B_K9NaHNCa3_0),.clk(gclk));
	jdff dff_B_xDbWoImo4_0(.din(w_dff_B_K9NaHNCa3_0),.dout(w_dff_B_xDbWoImo4_0),.clk(gclk));
	jdff dff_B_q0elnQ2I0_0(.din(w_dff_B_xDbWoImo4_0),.dout(w_dff_B_q0elnQ2I0_0),.clk(gclk));
	jdff dff_B_Li3oPenu2_0(.din(w_dff_B_q0elnQ2I0_0),.dout(w_dff_B_Li3oPenu2_0),.clk(gclk));
	jdff dff_B_75NlZSdJ8_0(.din(w_dff_B_Li3oPenu2_0),.dout(w_dff_B_75NlZSdJ8_0),.clk(gclk));
	jdff dff_B_ZXo0Ajip9_1(.din(n500),.dout(w_dff_B_ZXo0Ajip9_1),.clk(gclk));
	jdff dff_B_GWbKGlHL4_1(.din(n495),.dout(w_dff_B_GWbKGlHL4_1),.clk(gclk));
	jdff dff_B_UdMAZiz87_1(.din(G113),.dout(w_dff_B_UdMAZiz87_1),.clk(gclk));
	jdff dff_B_aljd1Jnr4_1(.din(w_dff_B_UdMAZiz87_1),.dout(w_dff_B_aljd1Jnr4_1),.clk(gclk));
	jdff dff_A_vrU2TEnj8_0(.dout(w_n1007_2[0]),.din(w_dff_A_vrU2TEnj8_0),.clk(gclk));
	jdff dff_A_c63SQAcV4_0(.dout(w_dff_A_vrU2TEnj8_0),.din(w_dff_A_c63SQAcV4_0),.clk(gclk));
	jdff dff_A_IhPVHmS03_0(.dout(w_dff_A_c63SQAcV4_0),.din(w_dff_A_IhPVHmS03_0),.clk(gclk));
	jdff dff_A_ppsnujPY6_0(.dout(w_dff_A_IhPVHmS03_0),.din(w_dff_A_ppsnujPY6_0),.clk(gclk));
	jdff dff_A_L3tuD2tc0_0(.dout(w_dff_A_ppsnujPY6_0),.din(w_dff_A_L3tuD2tc0_0),.clk(gclk));
	jdff dff_A_eY1SVWxl9_0(.dout(w_dff_A_L3tuD2tc0_0),.din(w_dff_A_eY1SVWxl9_0),.clk(gclk));
	jdff dff_A_A9qC9FTc9_1(.dout(w_n1007_2[1]),.din(w_dff_A_A9qC9FTc9_1),.clk(gclk));
	jdff dff_B_wd3WBX613_1(.din(n1216),.dout(w_dff_B_wd3WBX613_1),.clk(gclk));
	jdff dff_B_6TtA3TpS8_1(.din(w_dff_B_wd3WBX613_1),.dout(w_dff_B_6TtA3TpS8_1),.clk(gclk));
	jdff dff_B_5xvRDIY67_1(.din(w_dff_B_6TtA3TpS8_1),.dout(w_dff_B_5xvRDIY67_1),.clk(gclk));
	jdff dff_B_8dNRyRnD0_1(.din(w_dff_B_5xvRDIY67_1),.dout(w_dff_B_8dNRyRnD0_1),.clk(gclk));
	jdff dff_B_bPLbmZ3P5_1(.din(w_dff_B_8dNRyRnD0_1),.dout(w_dff_B_bPLbmZ3P5_1),.clk(gclk));
	jdff dff_B_5aPzewHF4_1(.din(w_dff_B_bPLbmZ3P5_1),.dout(w_dff_B_5aPzewHF4_1),.clk(gclk));
	jdff dff_B_mUOTr4No8_1(.din(w_dff_B_5aPzewHF4_1),.dout(w_dff_B_mUOTr4No8_1),.clk(gclk));
	jdff dff_B_tCN1YVT29_1(.din(w_dff_B_mUOTr4No8_1),.dout(w_dff_B_tCN1YVT29_1),.clk(gclk));
	jdff dff_B_EHvUj70j2_1(.din(w_dff_B_tCN1YVT29_1),.dout(w_dff_B_EHvUj70j2_1),.clk(gclk));
	jdff dff_B_yJWGdK1H6_1(.din(w_dff_B_EHvUj70j2_1),.dout(w_dff_B_yJWGdK1H6_1),.clk(gclk));
	jdff dff_B_J8o4nnxb3_1(.din(w_dff_B_yJWGdK1H6_1),.dout(w_dff_B_J8o4nnxb3_1),.clk(gclk));
	jdff dff_B_nhj6bx8W5_0(.din(n1219),.dout(w_dff_B_nhj6bx8W5_0),.clk(gclk));
	jdff dff_B_QAm637499_0(.din(w_dff_B_nhj6bx8W5_0),.dout(w_dff_B_QAm637499_0),.clk(gclk));
	jdff dff_B_iyvZikVc5_0(.din(w_dff_B_QAm637499_0),.dout(w_dff_B_iyvZikVc5_0),.clk(gclk));
	jdff dff_B_qxjqu7PP5_0(.din(w_dff_B_iyvZikVc5_0),.dout(w_dff_B_qxjqu7PP5_0),.clk(gclk));
	jdff dff_B_sltbgdBD4_0(.din(w_dff_B_qxjqu7PP5_0),.dout(w_dff_B_sltbgdBD4_0),.clk(gclk));
	jdff dff_B_Ghv57Xo84_0(.din(w_dff_B_sltbgdBD4_0),.dout(w_dff_B_Ghv57Xo84_0),.clk(gclk));
	jdff dff_B_fx5k9FZY9_0(.din(w_dff_B_Ghv57Xo84_0),.dout(w_dff_B_fx5k9FZY9_0),.clk(gclk));
	jdff dff_A_2Oqkcr7F2_1(.dout(w_n989_0[1]),.din(w_dff_A_2Oqkcr7F2_1),.clk(gclk));
	jdff dff_A_qO258kTB7_1(.dout(w_dff_A_2Oqkcr7F2_1),.din(w_dff_A_qO258kTB7_1),.clk(gclk));
	jdff dff_A_WqYq0zA37_1(.dout(w_dff_A_qO258kTB7_1),.din(w_dff_A_WqYq0zA37_1),.clk(gclk));
	jdff dff_A_GxTLhJZx7_1(.dout(w_dff_A_WqYq0zA37_1),.din(w_dff_A_GxTLhJZx7_1),.clk(gclk));
	jdff dff_A_wfN3sNeB6_1(.dout(w_dff_A_GxTLhJZx7_1),.din(w_dff_A_wfN3sNeB6_1),.clk(gclk));
	jdff dff_B_WcBNWtOU8_1(.din(n988),.dout(w_dff_B_WcBNWtOU8_1),.clk(gclk));
	jdff dff_B_bapi0k3s0_1(.din(w_dff_B_WcBNWtOU8_1),.dout(w_dff_B_bapi0k3s0_1),.clk(gclk));
	jdff dff_B_e1ncb7Vw9_1(.din(w_dff_B_bapi0k3s0_1),.dout(w_dff_B_e1ncb7Vw9_1),.clk(gclk));
	jdff dff_B_ymZyGPr64_1(.din(w_dff_B_e1ncb7Vw9_1),.dout(w_dff_B_ymZyGPr64_1),.clk(gclk));
	jdff dff_B_ndtNxg8A0_1(.din(w_dff_B_ymZyGPr64_1),.dout(w_dff_B_ndtNxg8A0_1),.clk(gclk));
	jdff dff_B_SyvHB0u91_1(.din(w_dff_B_ndtNxg8A0_1),.dout(w_dff_B_SyvHB0u91_1),.clk(gclk));
	jdff dff_B_0RGx7qUb3_1(.din(G112),.dout(w_dff_B_0RGx7qUb3_1),.clk(gclk));
	jdff dff_B_F7iw6GAC2_1(.din(w_dff_B_0RGx7qUb3_1),.dout(w_dff_B_F7iw6GAC2_1),.clk(gclk));
	jdff dff_A_ewr4SXXH1_0(.dout(w_G1691_3[0]),.din(w_dff_A_ewr4SXXH1_0),.clk(gclk));
	jdff dff_A_atevLuvj3_0(.dout(w_dff_A_ewr4SXXH1_0),.din(w_dff_A_atevLuvj3_0),.clk(gclk));
	jdff dff_A_31nNRVPo0_0(.dout(w_dff_A_atevLuvj3_0),.din(w_dff_A_31nNRVPo0_0),.clk(gclk));
	jdff dff_A_PTfTAvJb1_0(.dout(w_dff_A_31nNRVPo0_0),.din(w_dff_A_PTfTAvJb1_0),.clk(gclk));
	jdff dff_A_hdUzfdID3_1(.dout(w_G1691_3[1]),.din(w_dff_A_hdUzfdID3_1),.clk(gclk));
	jdff dff_A_vpSkG3G47_1(.dout(w_dff_A_hdUzfdID3_1),.din(w_dff_A_vpSkG3G47_1),.clk(gclk));
	jdff dff_B_3gObBvtq6_1(.din(n1382),.dout(w_dff_B_3gObBvtq6_1),.clk(gclk));
	jdff dff_B_7BNYNatJ7_1(.din(w_dff_B_3gObBvtq6_1),.dout(w_dff_B_7BNYNatJ7_1),.clk(gclk));
	jdff dff_B_vWtlvFBq7_1(.din(w_dff_B_7BNYNatJ7_1),.dout(w_dff_B_vWtlvFBq7_1),.clk(gclk));
	jdff dff_B_pal9sUyi5_1(.din(w_dff_B_vWtlvFBq7_1),.dout(w_dff_B_pal9sUyi5_1),.clk(gclk));
	jdff dff_B_sxWPdZfA4_1(.din(w_dff_B_pal9sUyi5_1),.dout(w_dff_B_sxWPdZfA4_1),.clk(gclk));
	jdff dff_B_pd2DNL1X3_1(.din(w_dff_B_sxWPdZfA4_1),.dout(w_dff_B_pd2DNL1X3_1),.clk(gclk));
	jdff dff_B_QU100WUX8_1(.din(w_dff_B_pd2DNL1X3_1),.dout(w_dff_B_QU100WUX8_1),.clk(gclk));
	jdff dff_B_27yDHJjp1_1(.din(w_dff_B_QU100WUX8_1),.dout(w_dff_B_27yDHJjp1_1),.clk(gclk));
	jdff dff_B_tUL6pXNC2_1(.din(w_dff_B_27yDHJjp1_1),.dout(w_dff_B_tUL6pXNC2_1),.clk(gclk));
	jdff dff_B_quc5fPgB3_1(.din(w_dff_B_tUL6pXNC2_1),.dout(w_dff_B_quc5fPgB3_1),.clk(gclk));
	jdff dff_B_JY4lHCv44_1(.din(w_dff_B_quc5fPgB3_1),.dout(w_dff_B_JY4lHCv44_1),.clk(gclk));
	jdff dff_B_uGKSFA9M9_1(.din(w_dff_B_JY4lHCv44_1),.dout(w_dff_B_uGKSFA9M9_1),.clk(gclk));
	jdff dff_B_qZageBzx2_1(.din(w_dff_B_uGKSFA9M9_1),.dout(w_dff_B_qZageBzx2_1),.clk(gclk));
	jdff dff_B_Kqho8I655_1(.din(w_dff_B_qZageBzx2_1),.dout(w_dff_B_Kqho8I655_1),.clk(gclk));
	jdff dff_B_zzhyHL5h9_1(.din(w_dff_B_Kqho8I655_1),.dout(w_dff_B_zzhyHL5h9_1),.clk(gclk));
	jdff dff_B_xYUlCryM1_1(.din(w_dff_B_zzhyHL5h9_1),.dout(w_dff_B_xYUlCryM1_1),.clk(gclk));
	jdff dff_B_kAxv4aJy7_1(.din(w_dff_B_xYUlCryM1_1),.dout(w_dff_B_kAxv4aJy7_1),.clk(gclk));
	jdff dff_B_T6D8dj7o7_1(.din(w_dff_B_kAxv4aJy7_1),.dout(w_dff_B_T6D8dj7o7_1),.clk(gclk));
	jdff dff_B_jthn2JR95_1(.din(w_dff_B_T6D8dj7o7_1),.dout(w_dff_B_jthn2JR95_1),.clk(gclk));
	jdff dff_B_FMdVkkiS9_1(.din(n1245),.dout(w_dff_B_FMdVkkiS9_1),.clk(gclk));
	jdff dff_B_RlXyN75Z2_1(.din(w_dff_B_FMdVkkiS9_1),.dout(w_dff_B_RlXyN75Z2_1),.clk(gclk));
	jdff dff_B_HffqlGeD3_1(.din(w_dff_B_RlXyN75Z2_1),.dout(w_dff_B_HffqlGeD3_1),.clk(gclk));
	jdff dff_B_BrRlp7DK5_1(.din(w_dff_B_HffqlGeD3_1),.dout(w_dff_B_BrRlp7DK5_1),.clk(gclk));
	jdff dff_B_HtTzx4SS0_1(.din(w_dff_B_BrRlp7DK5_1),.dout(w_dff_B_HtTzx4SS0_1),.clk(gclk));
	jdff dff_B_g4pXpyvD2_1(.din(w_dff_B_HtTzx4SS0_1),.dout(w_dff_B_g4pXpyvD2_1),.clk(gclk));
	jdff dff_B_qMC45aoi3_1(.din(w_dff_B_g4pXpyvD2_1),.dout(w_dff_B_qMC45aoi3_1),.clk(gclk));
	jdff dff_B_Ryg6WJ9s5_1(.din(w_dff_B_qMC45aoi3_1),.dout(w_dff_B_Ryg6WJ9s5_1),.clk(gclk));
	jdff dff_B_mYKFUuBt2_1(.din(w_dff_B_Ryg6WJ9s5_1),.dout(w_dff_B_mYKFUuBt2_1),.clk(gclk));
	jdff dff_B_ODHRcNGn0_1(.din(w_dff_B_mYKFUuBt2_1),.dout(w_dff_B_ODHRcNGn0_1),.clk(gclk));
	jdff dff_B_WB9zdLi83_1(.din(w_dff_B_ODHRcNGn0_1),.dout(w_dff_B_WB9zdLi83_1),.clk(gclk));
	jdff dff_B_VSfgctiF3_1(.din(w_dff_B_WB9zdLi83_1),.dout(w_dff_B_VSfgctiF3_1),.clk(gclk));
	jdff dff_B_h15wSets3_1(.din(w_dff_B_VSfgctiF3_1),.dout(w_dff_B_h15wSets3_1),.clk(gclk));
	jdff dff_B_nA4l5icK4_1(.din(w_dff_B_h15wSets3_1),.dout(w_dff_B_nA4l5icK4_1),.clk(gclk));
	jdff dff_B_FO7cTvde1_1(.din(w_dff_B_nA4l5icK4_1),.dout(w_dff_B_FO7cTvde1_1),.clk(gclk));
	jdff dff_B_IQtoGsNT7_1(.din(w_dff_B_FO7cTvde1_1),.dout(w_dff_B_IQtoGsNT7_1),.clk(gclk));
	jdff dff_B_qgl7C1FO8_1(.din(n1247),.dout(w_dff_B_qgl7C1FO8_1),.clk(gclk));
	jdff dff_B_BQmwYZ0S5_1(.din(w_dff_B_qgl7C1FO8_1),.dout(w_dff_B_BQmwYZ0S5_1),.clk(gclk));
	jdff dff_B_wmaGa7Tq4_1(.din(w_dff_B_BQmwYZ0S5_1),.dout(w_dff_B_wmaGa7Tq4_1),.clk(gclk));
	jdff dff_B_3GEBUdvs2_1(.din(w_dff_B_wmaGa7Tq4_1),.dout(w_dff_B_3GEBUdvs2_1),.clk(gclk));
	jdff dff_B_txWFpU7O5_1(.din(w_dff_B_3GEBUdvs2_1),.dout(w_dff_B_txWFpU7O5_1),.clk(gclk));
	jdff dff_B_LLRgr22f0_1(.din(w_dff_B_txWFpU7O5_1),.dout(w_dff_B_LLRgr22f0_1),.clk(gclk));
	jdff dff_B_8WiDnjDU1_1(.din(w_dff_B_LLRgr22f0_1),.dout(w_dff_B_8WiDnjDU1_1),.clk(gclk));
	jdff dff_B_4zoGhQZS1_1(.din(w_dff_B_8WiDnjDU1_1),.dout(w_dff_B_4zoGhQZS1_1),.clk(gclk));
	jdff dff_B_A6XYkeE92_1(.din(w_dff_B_4zoGhQZS1_1),.dout(w_dff_B_A6XYkeE92_1),.clk(gclk));
	jdff dff_B_poQmnGEx7_1(.din(w_dff_B_A6XYkeE92_1),.dout(w_dff_B_poQmnGEx7_1),.clk(gclk));
	jdff dff_B_Cp2TkbYB7_1(.din(w_dff_B_poQmnGEx7_1),.dout(w_dff_B_Cp2TkbYB7_1),.clk(gclk));
	jdff dff_B_rM69akLu3_1(.din(n951),.dout(w_dff_B_rM69akLu3_1),.clk(gclk));
	jdff dff_B_hhR8mnqz5_1(.din(w_dff_B_rM69akLu3_1),.dout(w_dff_B_hhR8mnqz5_1),.clk(gclk));
	jdff dff_B_M8GRt5Zw8_1(.din(w_dff_B_hhR8mnqz5_1),.dout(w_dff_B_M8GRt5Zw8_1),.clk(gclk));
	jdff dff_B_73a9uzZc8_1(.din(w_dff_B_M8GRt5Zw8_1),.dout(w_dff_B_73a9uzZc8_1),.clk(gclk));
	jdff dff_B_GNB9tcu21_1(.din(w_dff_B_73a9uzZc8_1),.dout(w_dff_B_GNB9tcu21_1),.clk(gclk));
	jdff dff_B_EzmdNFix3_1(.din(w_dff_B_GNB9tcu21_1),.dout(w_dff_B_EzmdNFix3_1),.clk(gclk));
	jdff dff_B_eInc3zi74_1(.din(w_dff_B_EzmdNFix3_1),.dout(w_dff_B_eInc3zi74_1),.clk(gclk));
	jdff dff_B_gwymAcpq4_1(.din(w_dff_B_eInc3zi74_1),.dout(w_dff_B_gwymAcpq4_1),.clk(gclk));
	jdff dff_B_6atzRXp50_1(.din(w_dff_B_gwymAcpq4_1),.dout(w_dff_B_6atzRXp50_1),.clk(gclk));
	jdff dff_B_0c6LfmK61_1(.din(n513),.dout(w_dff_B_0c6LfmK61_1),.clk(gclk));
	jdff dff_B_yOGDY6he7_1(.din(n508),.dout(w_dff_B_yOGDY6he7_1),.clk(gclk));
	jdff dff_B_DevnYb509_1(.din(G53),.dout(w_dff_B_DevnYb509_1),.clk(gclk));
	jdff dff_B_3LTRgAEm6_1(.din(w_dff_B_DevnYb509_1),.dout(w_dff_B_3LTRgAEm6_1),.clk(gclk));
	jdff dff_B_5P3q6PZK0_1(.din(n1207),.dout(w_dff_B_5P3q6PZK0_1),.clk(gclk));
	jdff dff_B_pKYzJm8L7_1(.din(w_dff_B_5P3q6PZK0_1),.dout(w_dff_B_pKYzJm8L7_1),.clk(gclk));
	jdff dff_B_gh8tn6QU6_1(.din(w_dff_B_pKYzJm8L7_1),.dout(w_dff_B_gh8tn6QU6_1),.clk(gclk));
	jdff dff_B_pIKEtVug2_1(.din(w_dff_B_gh8tn6QU6_1),.dout(w_dff_B_pIKEtVug2_1),.clk(gclk));
	jdff dff_B_YBUokWUn1_1(.din(w_dff_B_pIKEtVug2_1),.dout(w_dff_B_YBUokWUn1_1),.clk(gclk));
	jdff dff_B_UQh2oZzD2_1(.din(w_dff_B_YBUokWUn1_1),.dout(w_dff_B_UQh2oZzD2_1),.clk(gclk));
	jdff dff_B_mLOE9ARC1_1(.din(w_dff_B_UQh2oZzD2_1),.dout(w_dff_B_mLOE9ARC1_1),.clk(gclk));
	jdff dff_B_7C5wYFeg3_1(.din(w_dff_B_mLOE9ARC1_1),.dout(w_dff_B_7C5wYFeg3_1),.clk(gclk));
	jdff dff_B_tCXuAXLT7_1(.din(w_dff_B_7C5wYFeg3_1),.dout(w_dff_B_tCXuAXLT7_1),.clk(gclk));
	jdff dff_B_D6QwLJ9m6_1(.din(w_dff_B_tCXuAXLT7_1),.dout(w_dff_B_D6QwLJ9m6_1),.clk(gclk));
	jdff dff_B_VqM9cSes9_1(.din(w_dff_B_D6QwLJ9m6_1),.dout(w_dff_B_VqM9cSes9_1),.clk(gclk));
	jdff dff_B_5XZ1CRXX8_1(.din(w_dff_B_VqM9cSes9_1),.dout(w_dff_B_5XZ1CRXX8_1),.clk(gclk));
	jdff dff_B_GXFxBcp05_1(.din(w_dff_B_5XZ1CRXX8_1),.dout(w_dff_B_GXFxBcp05_1),.clk(gclk));
	jdff dff_B_QMHplCug2_1(.din(w_dff_B_GXFxBcp05_1),.dout(w_dff_B_QMHplCug2_1),.clk(gclk));
	jdff dff_B_WPIHHPTY2_1(.din(w_dff_B_QMHplCug2_1),.dout(w_dff_B_WPIHHPTY2_1),.clk(gclk));
	jdff dff_B_kWb1quw83_1(.din(w_dff_B_WPIHHPTY2_1),.dout(w_dff_B_kWb1quw83_1),.clk(gclk));
	jdff dff_B_rEvkE60D6_0(.din(n1211),.dout(w_dff_B_rEvkE60D6_0),.clk(gclk));
	jdff dff_B_zINwDq7O3_0(.din(w_dff_B_rEvkE60D6_0),.dout(w_dff_B_zINwDq7O3_0),.clk(gclk));
	jdff dff_B_zQ9aCCvk7_0(.din(w_dff_B_zINwDq7O3_0),.dout(w_dff_B_zQ9aCCvk7_0),.clk(gclk));
	jdff dff_B_lqbikiFs9_0(.din(w_dff_B_zQ9aCCvk7_0),.dout(w_dff_B_lqbikiFs9_0),.clk(gclk));
	jdff dff_B_ikIkOiEX1_0(.din(w_dff_B_lqbikiFs9_0),.dout(w_dff_B_ikIkOiEX1_0),.clk(gclk));
	jdff dff_B_g8HhNVks3_0(.din(w_dff_B_ikIkOiEX1_0),.dout(w_dff_B_g8HhNVks3_0),.clk(gclk));
	jdff dff_B_hZfhGPNm0_0(.din(w_dff_B_g8HhNVks3_0),.dout(w_dff_B_hZfhGPNm0_0),.clk(gclk));
	jdff dff_B_JHIZx4mV9_0(.din(w_dff_B_hZfhGPNm0_0),.dout(w_dff_B_JHIZx4mV9_0),.clk(gclk));
	jdff dff_B_OaAbXU2z9_0(.din(w_dff_B_JHIZx4mV9_0),.dout(w_dff_B_OaAbXU2z9_0),.clk(gclk));
	jdff dff_B_0wWjNpv39_0(.din(w_dff_B_OaAbXU2z9_0),.dout(w_dff_B_0wWjNpv39_0),.clk(gclk));
	jdff dff_B_4kuolSpY5_1(.din(n978),.dout(w_dff_B_4kuolSpY5_1),.clk(gclk));
	jdff dff_B_jz1Kwpoq7_1(.din(w_dff_B_4kuolSpY5_1),.dout(w_dff_B_jz1Kwpoq7_1),.clk(gclk));
	jdff dff_B_uH0ugx2r4_1(.din(w_dff_B_jz1Kwpoq7_1),.dout(w_dff_B_uH0ugx2r4_1),.clk(gclk));
	jdff dff_B_YLf6kt0O4_1(.din(w_dff_B_uH0ugx2r4_1),.dout(w_dff_B_YLf6kt0O4_1),.clk(gclk));
	jdff dff_B_ygeRtY650_1(.din(w_dff_B_YLf6kt0O4_1),.dout(w_dff_B_ygeRtY650_1),.clk(gclk));
	jdff dff_B_RSAys7RH0_1(.din(w_dff_B_ygeRtY650_1),.dout(w_dff_B_RSAys7RH0_1),.clk(gclk));
	jdff dff_B_PGwbWVVH2_1(.din(w_dff_B_RSAys7RH0_1),.dout(w_dff_B_PGwbWVVH2_1),.clk(gclk));
	jdff dff_B_FebDitlu7_1(.din(w_dff_B_PGwbWVVH2_1),.dout(w_dff_B_FebDitlu7_1),.clk(gclk));
	jdff dff_B_ICYdCDT54_1(.din(w_dff_B_FebDitlu7_1),.dout(w_dff_B_ICYdCDT54_1),.clk(gclk));
	jdff dff_B_pyHhzsWM4_1(.din(n982),.dout(w_dff_B_pyHhzsWM4_1),.clk(gclk));
	jdff dff_B_MyokzfJG6_1(.din(n980),.dout(w_dff_B_MyokzfJG6_1),.clk(gclk));
	jdff dff_B_qatXc8VV6_1(.din(w_dff_B_MyokzfJG6_1),.dout(w_dff_B_qatXc8VV6_1),.clk(gclk));
	jdff dff_B_5f5v76gk3_1(.din(w_dff_B_qatXc8VV6_1),.dout(w_dff_B_5f5v76gk3_1),.clk(gclk));
	jdff dff_B_9T0J95il7_1(.din(w_dff_B_5f5v76gk3_1),.dout(w_dff_B_9T0J95il7_1),.clk(gclk));
	jdff dff_B_0D9ogn6Y8_1(.din(w_dff_B_9T0J95il7_1),.dout(w_dff_B_0D9ogn6Y8_1),.clk(gclk));
	jdff dff_B_MF9Owc8L0_1(.din(G116),.dout(w_dff_B_MF9Owc8L0_1),.clk(gclk));
	jdff dff_B_kYjK86vv1_1(.din(w_dff_B_MF9Owc8L0_1),.dout(w_dff_B_kYjK86vv1_1),.clk(gclk));
	jdff dff_B_QCQEHJBJ9_0(.din(n1381),.dout(w_dff_B_QCQEHJBJ9_0),.clk(gclk));
	jdff dff_B_NwUqWdPU1_2(.din(G167),.dout(w_dff_B_NwUqWdPU1_2),.clk(gclk));
	jdff dff_B_KUr6AdJf3_2(.din(G197),.dout(w_dff_B_KUr6AdJf3_2),.clk(gclk));
	jdff dff_B_6Z1okz4h3_2(.din(w_dff_B_KUr6AdJf3_2),.dout(w_dff_B_6Z1okz4h3_2),.clk(gclk));
	jdff dff_B_yroClNli2_0(.din(n1395),.dout(w_dff_B_yroClNli2_0),.clk(gclk));
	jdff dff_B_zdAzHRRF8_0(.din(w_dff_B_yroClNli2_0),.dout(w_dff_B_zdAzHRRF8_0),.clk(gclk));
	jdff dff_B_6UYEQL2x2_0(.din(w_dff_B_zdAzHRRF8_0),.dout(w_dff_B_6UYEQL2x2_0),.clk(gclk));
	jdff dff_B_mfpd21pw8_0(.din(w_dff_B_6UYEQL2x2_0),.dout(w_dff_B_mfpd21pw8_0),.clk(gclk));
	jdff dff_B_udkTUowa9_0(.din(w_dff_B_mfpd21pw8_0),.dout(w_dff_B_udkTUowa9_0),.clk(gclk));
	jdff dff_B_hs6jSJjl1_0(.din(w_dff_B_udkTUowa9_0),.dout(w_dff_B_hs6jSJjl1_0),.clk(gclk));
	jdff dff_B_AWSvcsWE1_0(.din(w_dff_B_hs6jSJjl1_0),.dout(w_dff_B_AWSvcsWE1_0),.clk(gclk));
	jdff dff_B_rz8kvVKx4_0(.din(w_dff_B_AWSvcsWE1_0),.dout(w_dff_B_rz8kvVKx4_0),.clk(gclk));
	jdff dff_B_m0Oq0xMV3_0(.din(w_dff_B_rz8kvVKx4_0),.dout(w_dff_B_m0Oq0xMV3_0),.clk(gclk));
	jdff dff_B_yYVWrSDQ9_0(.din(w_dff_B_m0Oq0xMV3_0),.dout(w_dff_B_yYVWrSDQ9_0),.clk(gclk));
	jdff dff_B_oNLfMOBy9_0(.din(w_dff_B_yYVWrSDQ9_0),.dout(w_dff_B_oNLfMOBy9_0),.clk(gclk));
	jdff dff_B_zHKFq20D8_0(.din(w_dff_B_oNLfMOBy9_0),.dout(w_dff_B_zHKFq20D8_0),.clk(gclk));
	jdff dff_B_4W0Uptyo6_0(.din(w_dff_B_zHKFq20D8_0),.dout(w_dff_B_4W0Uptyo6_0),.clk(gclk));
	jdff dff_B_7Iq5rWsd2_0(.din(w_dff_B_4W0Uptyo6_0),.dout(w_dff_B_7Iq5rWsd2_0),.clk(gclk));
	jdff dff_B_pMCEaWye6_0(.din(w_dff_B_7Iq5rWsd2_0),.dout(w_dff_B_pMCEaWye6_0),.clk(gclk));
	jdff dff_B_RssjXhAQ3_0(.din(w_dff_B_pMCEaWye6_0),.dout(w_dff_B_RssjXhAQ3_0),.clk(gclk));
	jdff dff_B_8hCC8MqE5_0(.din(w_dff_B_RssjXhAQ3_0),.dout(w_dff_B_8hCC8MqE5_0),.clk(gclk));
	jdff dff_B_cRRZ9vyq5_0(.din(w_dff_B_8hCC8MqE5_0),.dout(w_dff_B_cRRZ9vyq5_0),.clk(gclk));
	jdff dff_B_aECCcNub3_0(.din(w_dff_B_cRRZ9vyq5_0),.dout(w_dff_B_aECCcNub3_0),.clk(gclk));
	jdff dff_B_j1n3kkOT6_0(.din(n1394),.dout(w_dff_B_j1n3kkOT6_0),.clk(gclk));
	jdff dff_B_shkYsADX0_2(.din(G164),.dout(w_dff_B_shkYsADX0_2),.clk(gclk));
	jdff dff_B_ForsF7Gk3_2(.din(G194),.dout(w_dff_B_ForsF7Gk3_2),.clk(gclk));
	jdff dff_B_GHXBL6V70_2(.din(w_dff_B_ForsF7Gk3_2),.dout(w_dff_B_GHXBL6V70_2),.clk(gclk));
	jdff dff_B_SATYeYta6_1(.din(n1389),.dout(w_dff_B_SATYeYta6_1),.clk(gclk));
	jdff dff_B_IRc6Jqif2_1(.din(w_dff_B_SATYeYta6_1),.dout(w_dff_B_IRc6Jqif2_1),.clk(gclk));
	jdff dff_B_SuASEOwW9_1(.din(n1239),.dout(w_dff_B_SuASEOwW9_1),.clk(gclk));
	jdff dff_B_khujN4kz9_1(.din(w_dff_B_SuASEOwW9_1),.dout(w_dff_B_khujN4kz9_1),.clk(gclk));
	jdff dff_B_F3Kxm83X1_1(.din(w_dff_B_khujN4kz9_1),.dout(w_dff_B_F3Kxm83X1_1),.clk(gclk));
	jdff dff_B_8dQBZvQ76_1(.din(w_dff_B_F3Kxm83X1_1),.dout(w_dff_B_8dQBZvQ76_1),.clk(gclk));
	jdff dff_B_aQaHBYYT8_1(.din(w_dff_B_8dQBZvQ76_1),.dout(w_dff_B_aQaHBYYT8_1),.clk(gclk));
	jdff dff_B_tlWiEksU1_1(.din(w_dff_B_aQaHBYYT8_1),.dout(w_dff_B_tlWiEksU1_1),.clk(gclk));
	jdff dff_B_V4g9B0Bc1_1(.din(w_dff_B_tlWiEksU1_1),.dout(w_dff_B_V4g9B0Bc1_1),.clk(gclk));
	jdff dff_B_4IMke6an4_1(.din(w_dff_B_V4g9B0Bc1_1),.dout(w_dff_B_4IMke6an4_1),.clk(gclk));
	jdff dff_B_is8T0Zvx8_1(.din(w_dff_B_4IMke6an4_1),.dout(w_dff_B_is8T0Zvx8_1),.clk(gclk));
	jdff dff_B_uY0k4gIV8_1(.din(w_dff_B_is8T0Zvx8_1),.dout(w_dff_B_uY0k4gIV8_1),.clk(gclk));
	jdff dff_B_p4AXBXKC0_1(.din(w_dff_B_uY0k4gIV8_1),.dout(w_dff_B_p4AXBXKC0_1),.clk(gclk));
	jdff dff_B_NTB3WyIr9_1(.din(w_dff_B_p4AXBXKC0_1),.dout(w_dff_B_NTB3WyIr9_1),.clk(gclk));
	jdff dff_B_KGmhtZ5V7_1(.din(w_dff_B_NTB3WyIr9_1),.dout(w_dff_B_KGmhtZ5V7_1),.clk(gclk));
	jdff dff_B_jXg2uAaj1_1(.din(w_dff_B_KGmhtZ5V7_1),.dout(w_dff_B_jXg2uAaj1_1),.clk(gclk));
	jdff dff_B_gDMHa5dD1_0(.din(n1242),.dout(w_dff_B_gDMHa5dD1_0),.clk(gclk));
	jdff dff_B_hnlt39in2_0(.din(w_dff_B_gDMHa5dD1_0),.dout(w_dff_B_hnlt39in2_0),.clk(gclk));
	jdff dff_B_CzjmnqsG2_0(.din(w_dff_B_hnlt39in2_0),.dout(w_dff_B_CzjmnqsG2_0),.clk(gclk));
	jdff dff_B_Uk6SWWo31_0(.din(w_dff_B_CzjmnqsG2_0),.dout(w_dff_B_Uk6SWWo31_0),.clk(gclk));
	jdff dff_B_amk12isJ4_0(.din(w_dff_B_Uk6SWWo31_0),.dout(w_dff_B_amk12isJ4_0),.clk(gclk));
	jdff dff_B_aqHn981c9_0(.din(w_dff_B_amk12isJ4_0),.dout(w_dff_B_aqHn981c9_0),.clk(gclk));
	jdff dff_B_TOhZOnpB9_0(.din(w_dff_B_aqHn981c9_0),.dout(w_dff_B_TOhZOnpB9_0),.clk(gclk));
	jdff dff_B_Y2HgL4gd1_0(.din(w_dff_B_TOhZOnpB9_0),.dout(w_dff_B_Y2HgL4gd1_0),.clk(gclk));
	jdff dff_B_JAOvdGPG3_0(.din(w_dff_B_Y2HgL4gd1_0),.dout(w_dff_B_JAOvdGPG3_0),.clk(gclk));
	jdff dff_B_Vhmy5KCT8_0(.din(w_dff_B_JAOvdGPG3_0),.dout(w_dff_B_Vhmy5KCT8_0),.clk(gclk));
	jdff dff_A_HArAgng82_1(.dout(w_n459_0[1]),.din(w_dff_A_HArAgng82_1),.clk(gclk));
	jdff dff_A_M0jMOAI95_1(.dout(w_dff_A_HArAgng82_1),.din(w_dff_A_M0jMOAI95_1),.clk(gclk));
	jdff dff_A_9OEWihJg9_1(.dout(w_dff_A_M0jMOAI95_1),.din(w_dff_A_9OEWihJg9_1),.clk(gclk));
	jdff dff_B_2TSL03jK6_1(.din(n455),.dout(w_dff_B_2TSL03jK6_1),.clk(gclk));
	jdff dff_B_q9Ly9YM44_3(.din(G3548),.dout(w_dff_B_q9Ly9YM44_3),.clk(gclk));
	jdff dff_B_cRRncVaF6_1(.din(n450),.dout(w_dff_B_cRRncVaF6_1),.clk(gclk));
	jdff dff_A_VoJQY4mK5_0(.dout(w_n749_6[0]),.din(w_dff_A_VoJQY4mK5_0),.clk(gclk));
	jdff dff_A_zOK6Sc6G1_0(.dout(w_dff_A_VoJQY4mK5_0),.din(w_dff_A_zOK6Sc6G1_0),.clk(gclk));
	jdff dff_A_W72xPigz0_0(.dout(w_dff_A_zOK6Sc6G1_0),.din(w_dff_A_W72xPigz0_0),.clk(gclk));
	jdff dff_A_XUWvpTXo5_0(.dout(w_dff_A_W72xPigz0_0),.din(w_dff_A_XUWvpTXo5_0),.clk(gclk));
	jdff dff_A_7EGXfocg3_0(.dout(w_dff_A_XUWvpTXo5_0),.din(w_dff_A_7EGXfocg3_0),.clk(gclk));
	jdff dff_A_jj5mAno66_0(.dout(w_dff_A_7EGXfocg3_0),.din(w_dff_A_jj5mAno66_0),.clk(gclk));
	jdff dff_A_aKgZac1K6_0(.dout(w_dff_A_jj5mAno66_0),.din(w_dff_A_aKgZac1K6_0),.clk(gclk));
	jdff dff_A_mDIJjcnI8_0(.dout(w_dff_A_aKgZac1K6_0),.din(w_dff_A_mDIJjcnI8_0),.clk(gclk));
	jdff dff_A_moObGmSF6_0(.dout(w_dff_A_mDIJjcnI8_0),.din(w_dff_A_moObGmSF6_0),.clk(gclk));
	jdff dff_A_2m1qgmXz6_0(.dout(w_dff_A_moObGmSF6_0),.din(w_dff_A_2m1qgmXz6_0),.clk(gclk));
	jdff dff_A_O9OK7o6x9_0(.dout(w_dff_A_2m1qgmXz6_0),.din(w_dff_A_O9OK7o6x9_0),.clk(gclk));
	jdff dff_A_09PEiPU34_1(.dout(w_n949_0[1]),.din(w_dff_A_09PEiPU34_1),.clk(gclk));
	jdff dff_A_uXdx9I4O0_1(.dout(w_dff_A_09PEiPU34_1),.din(w_dff_A_uXdx9I4O0_1),.clk(gclk));
	jdff dff_B_9fTv7oJp4_1(.din(n946),.dout(w_dff_B_9fTv7oJp4_1),.clk(gclk));
	jdff dff_B_c0RnFSPh6_1(.din(w_dff_B_9fTv7oJp4_1),.dout(w_dff_B_c0RnFSPh6_1),.clk(gclk));
	jdff dff_B_Wu4ANowT3_1(.din(w_dff_B_c0RnFSPh6_1),.dout(w_dff_B_Wu4ANowT3_1),.clk(gclk));
	jdff dff_B_Eq7yUAjh0_1(.din(w_dff_B_Wu4ANowT3_1),.dout(w_dff_B_Eq7yUAjh0_1),.clk(gclk));
	jdff dff_B_zqJrC4xK2_1(.din(w_dff_B_Eq7yUAjh0_1),.dout(w_dff_B_zqJrC4xK2_1),.clk(gclk));
	jdff dff_B_YgrLRGQT5_1(.din(w_dff_B_zqJrC4xK2_1),.dout(w_dff_B_YgrLRGQT5_1),.clk(gclk));
	jdff dff_A_yPdgnVZq1_0(.dout(w_G4091_2[0]),.din(w_dff_A_yPdgnVZq1_0),.clk(gclk));
	jdff dff_A_EQO7aPUZ7_0(.dout(w_dff_A_yPdgnVZq1_0),.din(w_dff_A_EQO7aPUZ7_0),.clk(gclk));
	jdff dff_A_Sdgvmiav8_1(.dout(w_G4091_2[1]),.din(w_dff_A_Sdgvmiav8_1),.clk(gclk));
	jdff dff_A_IFemFwP97_1(.dout(w_dff_A_Sdgvmiav8_1),.din(w_dff_A_IFemFwP97_1),.clk(gclk));
	jdff dff_A_DB8a6sF52_1(.dout(w_dff_A_IFemFwP97_1),.din(w_dff_A_DB8a6sF52_1),.clk(gclk));
	jdff dff_B_babhDdva3_1(.din(G114),.dout(w_dff_B_babhDdva3_1),.clk(gclk));
	jdff dff_B_Or80r8Bu4_1(.din(w_dff_B_babhDdva3_1),.dout(w_dff_B_Or80r8Bu4_1),.clk(gclk));
	jdff dff_A_bDAjTJQY5_0(.dout(w_n1008_2[0]),.din(w_dff_A_bDAjTJQY5_0),.clk(gclk));
	jdff dff_A_5i6QK7o84_1(.dout(w_n1008_2[1]),.din(w_dff_A_5i6QK7o84_1),.clk(gclk));
	jdff dff_B_50hXFk5M3_1(.din(n1198),.dout(w_dff_B_50hXFk5M3_1),.clk(gclk));
	jdff dff_B_FFfn2ho82_1(.din(w_dff_B_50hXFk5M3_1),.dout(w_dff_B_FFfn2ho82_1),.clk(gclk));
	jdff dff_B_SIN1FyzY3_1(.din(w_dff_B_FFfn2ho82_1),.dout(w_dff_B_SIN1FyzY3_1),.clk(gclk));
	jdff dff_B_Yu8UBpLi6_1(.din(w_dff_B_SIN1FyzY3_1),.dout(w_dff_B_Yu8UBpLi6_1),.clk(gclk));
	jdff dff_B_xWGtZ0OT7_1(.din(w_dff_B_Yu8UBpLi6_1),.dout(w_dff_B_xWGtZ0OT7_1),.clk(gclk));
	jdff dff_B_Kmxdsp1M9_1(.din(w_dff_B_xWGtZ0OT7_1),.dout(w_dff_B_Kmxdsp1M9_1),.clk(gclk));
	jdff dff_B_R9w9evNC0_1(.din(w_dff_B_Kmxdsp1M9_1),.dout(w_dff_B_R9w9evNC0_1),.clk(gclk));
	jdff dff_B_6JhyAsAc9_1(.din(w_dff_B_R9w9evNC0_1),.dout(w_dff_B_6JhyAsAc9_1),.clk(gclk));
	jdff dff_B_AGGg2M6Z2_1(.din(w_dff_B_6JhyAsAc9_1),.dout(w_dff_B_AGGg2M6Z2_1),.clk(gclk));
	jdff dff_B_cFioTv9R6_1(.din(w_dff_B_AGGg2M6Z2_1),.dout(w_dff_B_cFioTv9R6_1),.clk(gclk));
	jdff dff_B_wFZP9U8Z9_1(.din(w_dff_B_cFioTv9R6_1),.dout(w_dff_B_wFZP9U8Z9_1),.clk(gclk));
	jdff dff_B_oMLOhkRf6_1(.din(w_dff_B_wFZP9U8Z9_1),.dout(w_dff_B_oMLOhkRf6_1),.clk(gclk));
	jdff dff_B_e3JhcnfG7_1(.din(w_dff_B_oMLOhkRf6_1),.dout(w_dff_B_e3JhcnfG7_1),.clk(gclk));
	jdff dff_B_ot4T40aM7_1(.din(w_dff_B_e3JhcnfG7_1),.dout(w_dff_B_ot4T40aM7_1),.clk(gclk));
	jdff dff_B_UZUkPoFP0_1(.din(w_dff_B_ot4T40aM7_1),.dout(w_dff_B_UZUkPoFP0_1),.clk(gclk));
	jdff dff_B_dmjTBYiW3_1(.din(n1200),.dout(w_dff_B_dmjTBYiW3_1),.clk(gclk));
	jdff dff_B_zaz4tCVY8_1(.din(w_dff_B_dmjTBYiW3_1),.dout(w_dff_B_zaz4tCVY8_1),.clk(gclk));
	jdff dff_B_neIGb0Nn7_1(.din(w_dff_B_zaz4tCVY8_1),.dout(w_dff_B_neIGb0Nn7_1),.clk(gclk));
	jdff dff_B_w0ha3GHo1_1(.din(w_dff_B_neIGb0Nn7_1),.dout(w_dff_B_w0ha3GHo1_1),.clk(gclk));
	jdff dff_B_iyvx0Osu3_1(.din(w_dff_B_w0ha3GHo1_1),.dout(w_dff_B_iyvx0Osu3_1),.clk(gclk));
	jdff dff_B_ypEKkKHu1_1(.din(w_dff_B_iyvx0Osu3_1),.dout(w_dff_B_ypEKkKHu1_1),.clk(gclk));
	jdff dff_B_1HBEN5Er7_1(.din(w_dff_B_ypEKkKHu1_1),.dout(w_dff_B_1HBEN5Er7_1),.clk(gclk));
	jdff dff_B_9orisDh76_1(.din(w_dff_B_1HBEN5Er7_1),.dout(w_dff_B_9orisDh76_1),.clk(gclk));
	jdff dff_B_NwbyyCxe4_1(.din(w_dff_B_9orisDh76_1),.dout(w_dff_B_NwbyyCxe4_1),.clk(gclk));
	jdff dff_B_ovtLENyn1_1(.din(w_dff_B_NwbyyCxe4_1),.dout(w_dff_B_ovtLENyn1_1),.clk(gclk));
	jdff dff_B_TA9c7iQR3_1(.din(w_dff_B_ovtLENyn1_1),.dout(w_dff_B_TA9c7iQR3_1),.clk(gclk));
	jdff dff_A_KpkyMcK08_0(.dout(w_n649_0[0]),.din(w_dff_A_KpkyMcK08_0),.clk(gclk));
	jdff dff_A_AIMvmSNJ1_0(.dout(w_dff_A_KpkyMcK08_0),.din(w_dff_A_AIMvmSNJ1_0),.clk(gclk));
	jdff dff_A_uAYq9qwW0_0(.dout(w_dff_A_AIMvmSNJ1_0),.din(w_dff_A_uAYq9qwW0_0),.clk(gclk));
	jdff dff_A_sXdHsCJz1_0(.dout(w_dff_A_uAYq9qwW0_0),.din(w_dff_A_sXdHsCJz1_0),.clk(gclk));
	jdff dff_A_Sp5I7ldP9_0(.dout(w_dff_A_sXdHsCJz1_0),.din(w_dff_A_Sp5I7ldP9_0),.clk(gclk));
	jdff dff_A_vqtaKSFB4_0(.dout(w_dff_A_Sp5I7ldP9_0),.din(w_dff_A_vqtaKSFB4_0),.clk(gclk));
	jdff dff_A_mlYvGYp88_0(.dout(w_dff_A_vqtaKSFB4_0),.din(w_dff_A_mlYvGYp88_0),.clk(gclk));
	jdff dff_A_BDO4lIXq1_0(.dout(w_dff_A_mlYvGYp88_0),.din(w_dff_A_BDO4lIXq1_0),.clk(gclk));
	jdff dff_A_M55HYp4e6_0(.dout(w_dff_A_BDO4lIXq1_0),.din(w_dff_A_M55HYp4e6_0),.clk(gclk));
	jdff dff_A_5CRQ0zB80_1(.dout(w_n749_8[1]),.din(w_dff_A_5CRQ0zB80_1),.clk(gclk));
	jdff dff_A_jES8ImbP5_1(.dout(w_dff_A_5CRQ0zB80_1),.din(w_dff_A_jES8ImbP5_1),.clk(gclk));
	jdff dff_A_g6TZUcjN9_1(.dout(w_dff_A_jES8ImbP5_1),.din(w_dff_A_g6TZUcjN9_1),.clk(gclk));
	jdff dff_A_rH4vGzSu7_1(.dout(w_dff_A_g6TZUcjN9_1),.din(w_dff_A_rH4vGzSu7_1),.clk(gclk));
	jdff dff_A_l22ymRVk8_1(.dout(w_dff_A_rH4vGzSu7_1),.din(w_dff_A_l22ymRVk8_1),.clk(gclk));
	jdff dff_A_r41c0YZ74_1(.dout(w_dff_A_l22ymRVk8_1),.din(w_dff_A_r41c0YZ74_1),.clk(gclk));
	jdff dff_A_tsD94GUS7_1(.dout(w_dff_A_r41c0YZ74_1),.din(w_dff_A_tsD94GUS7_1),.clk(gclk));
	jdff dff_A_usWIVe4r6_1(.dout(w_dff_A_tsD94GUS7_1),.din(w_dff_A_usWIVe4r6_1),.clk(gclk));
	jdff dff_A_VbB6nsO87_1(.dout(w_dff_A_usWIVe4r6_1),.din(w_dff_A_VbB6nsO87_1),.clk(gclk));
	jdff dff_A_Gm075tNU0_1(.dout(w_dff_A_VbB6nsO87_1),.din(w_dff_A_Gm075tNU0_1),.clk(gclk));
	jdff dff_A_8x7QodEG0_1(.dout(w_dff_A_Gm075tNU0_1),.din(w_dff_A_8x7QodEG0_1),.clk(gclk));
	jdff dff_A_GPQp5Te57_1(.dout(w_dff_A_8x7QodEG0_1),.din(w_dff_A_GPQp5Te57_1),.clk(gclk));
	jdff dff_A_MpLo72ts6_2(.dout(w_n749_8[2]),.din(w_dff_A_MpLo72ts6_2),.clk(gclk));
	jdff dff_A_3E1I7apd9_2(.dout(w_dff_A_MpLo72ts6_2),.din(w_dff_A_3E1I7apd9_2),.clk(gclk));
	jdff dff_A_gY5xpIeV8_2(.dout(w_dff_A_3E1I7apd9_2),.din(w_dff_A_gY5xpIeV8_2),.clk(gclk));
	jdff dff_A_DFk1rNYC3_2(.dout(w_dff_A_gY5xpIeV8_2),.din(w_dff_A_DFk1rNYC3_2),.clk(gclk));
	jdff dff_A_9YSRrLIq5_2(.dout(w_dff_A_DFk1rNYC3_2),.din(w_dff_A_9YSRrLIq5_2),.clk(gclk));
	jdff dff_A_ceGm2RIz5_2(.dout(w_dff_A_9YSRrLIq5_2),.din(w_dff_A_ceGm2RIz5_2),.clk(gclk));
	jdff dff_A_khqusC305_2(.dout(w_dff_A_ceGm2RIz5_2),.din(w_dff_A_khqusC305_2),.clk(gclk));
	jdff dff_A_ZIh2Izqh5_2(.dout(w_dff_A_khqusC305_2),.din(w_dff_A_ZIh2Izqh5_2),.clk(gclk));
	jdff dff_A_oOh3FEj50_2(.dout(w_dff_A_ZIh2Izqh5_2),.din(w_dff_A_oOh3FEj50_2),.clk(gclk));
	jdff dff_A_kRe9C1FU2_2(.dout(w_dff_A_oOh3FEj50_2),.din(w_dff_A_kRe9C1FU2_2),.clk(gclk));
	jdff dff_B_2Ko6HozK1_1(.din(G121),.dout(w_dff_B_2Ko6HozK1_1),.clk(gclk));
	jdff dff_B_4nhfmZyy7_1(.din(w_dff_B_2Ko6HozK1_1),.dout(w_dff_B_4nhfmZyy7_1),.clk(gclk));
	jdff dff_A_kCA1roIz8_0(.dout(w_G137_4[0]),.din(w_dff_A_kCA1roIz8_0),.clk(gclk));
	jdff dff_A_Ii9nEp3G4_1(.dout(w_G137_4[1]),.din(w_dff_A_Ii9nEp3G4_1),.clk(gclk));
	jdff dff_A_Uantm8hy6_0(.dout(w_G137_1[0]),.din(w_dff_A_Uantm8hy6_0),.clk(gclk));
	jdff dff_A_EvlWgjHm5_0(.dout(w_dff_A_Uantm8hy6_0),.din(w_dff_A_EvlWgjHm5_0),.clk(gclk));
	jdff dff_A_zFhXjUh34_0(.dout(w_dff_A_EvlWgjHm5_0),.din(w_dff_A_zFhXjUh34_0),.clk(gclk));
	jdff dff_A_5SjB4z280_0(.dout(w_dff_A_zFhXjUh34_0),.din(w_dff_A_5SjB4z280_0),.clk(gclk));
	jdff dff_A_GTGvGoaV3_0(.dout(w_dff_A_5SjB4z280_0),.din(w_dff_A_GTGvGoaV3_0),.clk(gclk));
	jdff dff_A_9SF0wWVx1_0(.dout(w_dff_A_GTGvGoaV3_0),.din(w_dff_A_9SF0wWVx1_0),.clk(gclk));
	jdff dff_A_5UICh8js7_1(.dout(w_G137_1[1]),.din(w_dff_A_5UICh8js7_1),.clk(gclk));
	jdff dff_A_fvgm4vOr9_1(.dout(w_dff_A_5UICh8js7_1),.din(w_dff_A_fvgm4vOr9_1),.clk(gclk));
	jdff dff_A_jFoquQJb9_1(.dout(w_dff_A_fvgm4vOr9_1),.din(w_dff_A_jFoquQJb9_1),.clk(gclk));
	jdff dff_A_rm8v5iUM7_1(.dout(w_dff_A_jFoquQJb9_1),.din(w_dff_A_rm8v5iUM7_1),.clk(gclk));
	jdff dff_A_rqTSfhJM6_1(.dout(w_dff_A_rm8v5iUM7_1),.din(w_dff_A_rqTSfhJM6_1),.clk(gclk));
	jdff dff_A_ViVAQnti7_1(.dout(w_dff_A_rqTSfhJM6_1),.din(w_dff_A_ViVAQnti7_1),.clk(gclk));
	jdff dff_A_z3v7vRp71_1(.dout(w_dff_A_ViVAQnti7_1),.din(w_dff_A_z3v7vRp71_1),.clk(gclk));
	jdff dff_B_IaT2PVUl3_0(.din(n1404),.dout(w_dff_B_IaT2PVUl3_0),.clk(gclk));
	jdff dff_B_OPohOdCj5_0(.din(w_dff_B_IaT2PVUl3_0),.dout(w_dff_B_OPohOdCj5_0),.clk(gclk));
	jdff dff_B_Sz85MPJU5_0(.din(w_dff_B_OPohOdCj5_0),.dout(w_dff_B_Sz85MPJU5_0),.clk(gclk));
	jdff dff_B_aKXskUcH3_0(.din(w_dff_B_Sz85MPJU5_0),.dout(w_dff_B_aKXskUcH3_0),.clk(gclk));
	jdff dff_B_9uX8harz7_0(.din(w_dff_B_aKXskUcH3_0),.dout(w_dff_B_9uX8harz7_0),.clk(gclk));
	jdff dff_B_9QUziSNQ6_0(.din(w_dff_B_9uX8harz7_0),.dout(w_dff_B_9QUziSNQ6_0),.clk(gclk));
	jdff dff_B_dhOeJycN7_0(.din(w_dff_B_9QUziSNQ6_0),.dout(w_dff_B_dhOeJycN7_0),.clk(gclk));
	jdff dff_B_jBhjZjjS2_0(.din(w_dff_B_dhOeJycN7_0),.dout(w_dff_B_jBhjZjjS2_0),.clk(gclk));
	jdff dff_B_57gpdxxg8_0(.din(w_dff_B_jBhjZjjS2_0),.dout(w_dff_B_57gpdxxg8_0),.clk(gclk));
	jdff dff_B_0MA2VM3V0_0(.din(w_dff_B_57gpdxxg8_0),.dout(w_dff_B_0MA2VM3V0_0),.clk(gclk));
	jdff dff_B_9qarWJfO7_0(.din(w_dff_B_0MA2VM3V0_0),.dout(w_dff_B_9qarWJfO7_0),.clk(gclk));
	jdff dff_B_ijD61zwB8_0(.din(w_dff_B_9qarWJfO7_0),.dout(w_dff_B_ijD61zwB8_0),.clk(gclk));
	jdff dff_B_bkfVty1l4_0(.din(w_dff_B_ijD61zwB8_0),.dout(w_dff_B_bkfVty1l4_0),.clk(gclk));
	jdff dff_B_5qIDoWML4_0(.din(w_dff_B_bkfVty1l4_0),.dout(w_dff_B_5qIDoWML4_0),.clk(gclk));
	jdff dff_B_w3f5EaIq8_0(.din(w_dff_B_5qIDoWML4_0),.dout(w_dff_B_w3f5EaIq8_0),.clk(gclk));
	jdff dff_B_NRyAP7tH3_0(.din(w_dff_B_w3f5EaIq8_0),.dout(w_dff_B_NRyAP7tH3_0),.clk(gclk));
	jdff dff_B_fzndBmR54_0(.din(w_dff_B_NRyAP7tH3_0),.dout(w_dff_B_fzndBmR54_0),.clk(gclk));
	jdff dff_B_l1DuayOK1_0(.din(w_dff_B_fzndBmR54_0),.dout(w_dff_B_l1DuayOK1_0),.clk(gclk));
	jdff dff_B_80SRCvM26_0(.din(w_dff_B_l1DuayOK1_0),.dout(w_dff_B_80SRCvM26_0),.clk(gclk));
	jdff dff_B_E3wrtXIv4_0(.din(n1403),.dout(w_dff_B_E3wrtXIv4_0),.clk(gclk));
	jdff dff_B_ZoSLA8cb9_2(.din(G161),.dout(w_dff_B_ZoSLA8cb9_2),.clk(gclk));
	jdff dff_B_7uLmyHdV4_2(.din(G191),.dout(w_dff_B_7uLmyHdV4_2),.clk(gclk));
	jdff dff_B_fGuvLndO3_2(.din(w_dff_B_7uLmyHdV4_2),.dout(w_dff_B_fGuvLndO3_2),.clk(gclk));
	jdff dff_B_V0qgLHDs2_1(.din(n1190),.dout(w_dff_B_V0qgLHDs2_1),.clk(gclk));
	jdff dff_B_9KWmcCOm7_1(.din(w_dff_B_V0qgLHDs2_1),.dout(w_dff_B_9KWmcCOm7_1),.clk(gclk));
	jdff dff_B_f1VurmMl8_1(.din(w_dff_B_9KWmcCOm7_1),.dout(w_dff_B_f1VurmMl8_1),.clk(gclk));
	jdff dff_B_N78XHgTI0_1(.din(w_dff_B_f1VurmMl8_1),.dout(w_dff_B_N78XHgTI0_1),.clk(gclk));
	jdff dff_B_TihVkcu21_1(.din(w_dff_B_N78XHgTI0_1),.dout(w_dff_B_TihVkcu21_1),.clk(gclk));
	jdff dff_B_8gj5Y2tG9_1(.din(w_dff_B_TihVkcu21_1),.dout(w_dff_B_8gj5Y2tG9_1),.clk(gclk));
	jdff dff_B_YJDpsx4H3_1(.din(w_dff_B_8gj5Y2tG9_1),.dout(w_dff_B_YJDpsx4H3_1),.clk(gclk));
	jdff dff_B_HCH1NubT5_1(.din(w_dff_B_YJDpsx4H3_1),.dout(w_dff_B_HCH1NubT5_1),.clk(gclk));
	jdff dff_B_XW4WyXIR5_1(.din(w_dff_B_HCH1NubT5_1),.dout(w_dff_B_XW4WyXIR5_1),.clk(gclk));
	jdff dff_B_CelSJfSW6_1(.din(w_dff_B_XW4WyXIR5_1),.dout(w_dff_B_CelSJfSW6_1),.clk(gclk));
	jdff dff_B_fAe2TAn28_1(.din(w_dff_B_CelSJfSW6_1),.dout(w_dff_B_fAe2TAn28_1),.clk(gclk));
	jdff dff_B_8qwtpWrV4_1(.din(w_dff_B_fAe2TAn28_1),.dout(w_dff_B_8qwtpWrV4_1),.clk(gclk));
	jdff dff_B_V4Ppvtsg0_1(.din(w_dff_B_8qwtpWrV4_1),.dout(w_dff_B_V4Ppvtsg0_1),.clk(gclk));
	jdff dff_B_34MWWBSD3_1(.din(w_dff_B_V4Ppvtsg0_1),.dout(w_dff_B_34MWWBSD3_1),.clk(gclk));
	jdff dff_B_G67N6VPI7_1(.din(w_dff_B_34MWWBSD3_1),.dout(w_dff_B_G67N6VPI7_1),.clk(gclk));
	jdff dff_B_BGM5W6S45_1(.din(w_dff_B_G67N6VPI7_1),.dout(w_dff_B_BGM5W6S45_1),.clk(gclk));
	jdff dff_B_GKfzRS3d7_0(.din(n1194),.dout(w_dff_B_GKfzRS3d7_0),.clk(gclk));
	jdff dff_B_VzNzpOiO9_0(.din(w_dff_B_GKfzRS3d7_0),.dout(w_dff_B_VzNzpOiO9_0),.clk(gclk));
	jdff dff_B_lJ3dHqQx5_0(.din(w_dff_B_VzNzpOiO9_0),.dout(w_dff_B_lJ3dHqQx5_0),.clk(gclk));
	jdff dff_B_QVsNxBfM1_0(.din(w_dff_B_lJ3dHqQx5_0),.dout(w_dff_B_QVsNxBfM1_0),.clk(gclk));
	jdff dff_B_Tzipyeb02_0(.din(w_dff_B_QVsNxBfM1_0),.dout(w_dff_B_Tzipyeb02_0),.clk(gclk));
	jdff dff_B_eD5iR0z97_0(.din(w_dff_B_Tzipyeb02_0),.dout(w_dff_B_eD5iR0z97_0),.clk(gclk));
	jdff dff_B_jZNhevm24_0(.din(w_dff_B_eD5iR0z97_0),.dout(w_dff_B_jZNhevm24_0),.clk(gclk));
	jdff dff_B_yv72Z9yD3_0(.din(w_dff_B_jZNhevm24_0),.dout(w_dff_B_yv72Z9yD3_0),.clk(gclk));
	jdff dff_B_aXOr8GyN4_0(.din(w_dff_B_yv72Z9yD3_0),.dout(w_dff_B_aXOr8GyN4_0),.clk(gclk));
	jdff dff_B_VmEIurYj1_0(.din(w_dff_B_aXOr8GyN4_0),.dout(w_dff_B_VmEIurYj1_0),.clk(gclk));
	jdff dff_B_WLwvlIPA5_0(.din(w_dff_B_VmEIurYj1_0),.dout(w_dff_B_WLwvlIPA5_0),.clk(gclk));
	jdff dff_B_s4WOZmBm6_0(.din(w_dff_B_WLwvlIPA5_0),.dout(w_dff_B_s4WOZmBm6_0),.clk(gclk));
	jdff dff_A_BH3rsD105_1(.dout(w_G4092_6[1]),.din(w_dff_A_BH3rsD105_1),.clk(gclk));
	jdff dff_A_rLeApYgQ2_1(.dout(w_dff_A_BH3rsD105_1),.din(w_dff_A_rLeApYgQ2_1),.clk(gclk));
	jdff dff_A_nymskFp84_2(.dout(w_G4092_6[2]),.din(w_dff_A_nymskFp84_2),.clk(gclk));
	jdff dff_A_Zoy8pnXB4_2(.dout(w_dff_A_nymskFp84_2),.din(w_dff_A_Zoy8pnXB4_2),.clk(gclk));
	jdff dff_B_7CzP2E2L3_0(.din(n794),.dout(w_dff_B_7CzP2E2L3_0),.clk(gclk));
	jdff dff_B_m8lrl0n79_0(.din(n785),.dout(w_dff_B_m8lrl0n79_0),.clk(gclk));
	jdff dff_A_BmOSzjts1_0(.dout(w_G54_0[0]),.din(w_dff_A_BmOSzjts1_0),.clk(gclk));
	jdff dff_A_sGehzmu81_0(.dout(w_dff_A_BmOSzjts1_0),.din(w_dff_A_sGehzmu81_0),.clk(gclk));
	jdff dff_A_Rni5PH7f7_0(.dout(w_dff_A_sGehzmu81_0),.din(w_dff_A_Rni5PH7f7_0),.clk(gclk));
	jdff dff_A_u0eNrmBu4_0(.dout(w_dff_A_Rni5PH7f7_0),.din(w_dff_A_u0eNrmBu4_0),.clk(gclk));
	jdff dff_A_GbWrzrA04_0(.dout(w_dff_A_u0eNrmBu4_0),.din(w_dff_A_GbWrzrA04_0),.clk(gclk));
	jdff dff_A_dgYS5rF39_0(.dout(w_dff_A_GbWrzrA04_0),.din(w_dff_A_dgYS5rF39_0),.clk(gclk));
	jdff dff_A_HKIO64mQ1_0(.dout(w_dff_A_dgYS5rF39_0),.din(w_dff_A_HKIO64mQ1_0),.clk(gclk));
	jdff dff_A_6WBjMV9a8_0(.dout(w_dff_A_HKIO64mQ1_0),.din(w_dff_A_6WBjMV9a8_0),.clk(gclk));
	jdff dff_A_IjOfffxg2_0(.dout(w_dff_A_6WBjMV9a8_0),.din(w_dff_A_IjOfffxg2_0),.clk(gclk));
	jdff dff_A_5zH7QhnH9_1(.dout(w_G54_0[1]),.din(w_dff_A_5zH7QhnH9_1),.clk(gclk));
	jdff dff_A_wJ3Ouuzb5_1(.dout(w_dff_A_5zH7QhnH9_1),.din(w_dff_A_wJ3Ouuzb5_1),.clk(gclk));
	jdff dff_A_WbcQvHDP1_1(.dout(w_dff_A_wJ3Ouuzb5_1),.din(w_dff_A_WbcQvHDP1_1),.clk(gclk));
	jdff dff_A_w3gOLomI2_1(.dout(w_dff_A_WbcQvHDP1_1),.din(w_dff_A_w3gOLomI2_1),.clk(gclk));
	jdff dff_A_NxClbYBH0_0(.dout(w_n749_9[0]),.din(w_dff_A_NxClbYBH0_0),.clk(gclk));
	jdff dff_A_1Dx4HAHp7_2(.dout(w_n749_9[2]),.din(w_dff_A_1Dx4HAHp7_2),.clk(gclk));
	jdff dff_A_qso3eQg61_2(.dout(w_dff_A_1Dx4HAHp7_2),.din(w_dff_A_qso3eQg61_2),.clk(gclk));
	jdff dff_A_xQg7Be0V8_2(.dout(w_dff_A_qso3eQg61_2),.din(w_dff_A_xQg7Be0V8_2),.clk(gclk));
	jdff dff_A_UcqKxuSJ8_2(.dout(w_dff_A_xQg7Be0V8_2),.din(w_dff_A_UcqKxuSJ8_2),.clk(gclk));
	jdff dff_A_oZwZOjGH5_2(.dout(w_dff_A_UcqKxuSJ8_2),.din(w_dff_A_oZwZOjGH5_2),.clk(gclk));
	jdff dff_A_xj9gEQvJ1_2(.dout(w_dff_A_oZwZOjGH5_2),.din(w_dff_A_xj9gEQvJ1_2),.clk(gclk));
	jdff dff_A_eLxW5qXp5_2(.dout(w_dff_A_xj9gEQvJ1_2),.din(w_dff_A_eLxW5qXp5_2),.clk(gclk));
	jdff dff_A_1CdI0S0G6_2(.dout(w_dff_A_eLxW5qXp5_2),.din(w_dff_A_1CdI0S0G6_2),.clk(gclk));
	jdff dff_A_rdRbeQpz7_2(.dout(w_dff_A_1CdI0S0G6_2),.din(w_dff_A_rdRbeQpz7_2),.clk(gclk));
	jdff dff_A_DKIsNxmh3_2(.dout(w_dff_A_rdRbeQpz7_2),.din(w_dff_A_DKIsNxmh3_2),.clk(gclk));
	jdff dff_A_tFqvLuoQ2_2(.dout(w_dff_A_DKIsNxmh3_2),.din(w_dff_A_tFqvLuoQ2_2),.clk(gclk));
	jdff dff_A_nnfxkria6_2(.dout(w_dff_A_tFqvLuoQ2_2),.din(w_dff_A_nnfxkria6_2),.clk(gclk));
	jdff dff_A_LFp7k7aZ3_2(.dout(w_dff_A_nnfxkria6_2),.din(w_dff_A_LFp7k7aZ3_2),.clk(gclk));
	jdff dff_A_aOqhSAk29_2(.dout(w_dff_A_LFp7k7aZ3_2),.din(w_dff_A_aOqhSAk29_2),.clk(gclk));
	jdff dff_A_u5tFlz3S7_0(.dout(w_G123_0[0]),.din(w_dff_A_u5tFlz3S7_0),.clk(gclk));
	jdff dff_A_bJ19DS6e9_0(.dout(w_dff_A_u5tFlz3S7_0),.din(w_dff_A_bJ19DS6e9_0),.clk(gclk));
	jdff dff_A_phMaxgek3_0(.dout(w_G1691_2[0]),.din(w_dff_A_phMaxgek3_0),.clk(gclk));
	jdff dff_A_4i0Tqhj48_2(.dout(w_G1691_2[2]),.din(w_dff_A_4i0Tqhj48_2),.clk(gclk));
	jdff dff_A_0YtcJIVr1_2(.dout(w_n1007_1[2]),.din(w_dff_A_0YtcJIVr1_2),.clk(gclk));
	jdff dff_A_5ZHG9g6R5_0(.dout(w_n1007_0[0]),.din(w_dff_A_5ZHG9g6R5_0),.clk(gclk));
	jdff dff_A_wfRDHPzP8_0(.dout(w_dff_A_5ZHG9g6R5_0),.din(w_dff_A_wfRDHPzP8_0),.clk(gclk));
	jdff dff_A_hD979AwS9_0(.dout(w_dff_A_wfRDHPzP8_0),.din(w_dff_A_hD979AwS9_0),.clk(gclk));
	jdff dff_A_9HBBF0OZ2_0(.dout(w_dff_A_hD979AwS9_0),.din(w_dff_A_9HBBF0OZ2_0),.clk(gclk));
	jdff dff_A_kNJtKEVH1_0(.dout(w_dff_A_9HBBF0OZ2_0),.din(w_dff_A_kNJtKEVH1_0),.clk(gclk));
	jdff dff_A_A93dWc351_0(.dout(w_dff_A_kNJtKEVH1_0),.din(w_dff_A_A93dWc351_0),.clk(gclk));
	jdff dff_A_1fpD5eUO1_0(.dout(w_dff_A_A93dWc351_0),.din(w_dff_A_1fpD5eUO1_0),.clk(gclk));
	jdff dff_A_1UH77wLh7_0(.dout(w_dff_A_1fpD5eUO1_0),.din(w_dff_A_1UH77wLh7_0),.clk(gclk));
	jdff dff_A_H4V82B3V1_0(.dout(w_dff_A_1UH77wLh7_0),.din(w_dff_A_H4V82B3V1_0),.clk(gclk));
	jdff dff_A_DKLNwFK66_1(.dout(w_n1007_0[1]),.din(w_dff_A_DKLNwFK66_1),.clk(gclk));
	jdff dff_A_u2T2DKa28_1(.dout(w_dff_A_DKLNwFK66_1),.din(w_dff_A_u2T2DKa28_1),.clk(gclk));
	jdff dff_B_7eAZoxY13_3(.din(n1007),.dout(w_dff_B_7eAZoxY13_3),.clk(gclk));
	jdff dff_B_CWRxvdPn2_3(.din(w_dff_B_7eAZoxY13_3),.dout(w_dff_B_CWRxvdPn2_3),.clk(gclk));
	jdff dff_B_4g4Q6Rvf1_3(.din(w_dff_B_CWRxvdPn2_3),.dout(w_dff_B_4g4Q6Rvf1_3),.clk(gclk));
	jdff dff_B_7pfkPapK2_3(.din(w_dff_B_4g4Q6Rvf1_3),.dout(w_dff_B_7pfkPapK2_3),.clk(gclk));
	jdff dff_B_IGDUEajs0_3(.din(w_dff_B_7pfkPapK2_3),.dout(w_dff_B_IGDUEajs0_3),.clk(gclk));
	jdff dff_B_wcC1iBGy8_3(.din(w_dff_B_IGDUEajs0_3),.dout(w_dff_B_wcC1iBGy8_3),.clk(gclk));
	jdff dff_B_ylLpoCZ65_3(.din(w_dff_B_wcC1iBGy8_3),.dout(w_dff_B_ylLpoCZ65_3),.clk(gclk));
	jdff dff_B_dQiEg0El9_3(.din(w_dff_B_ylLpoCZ65_3),.dout(w_dff_B_dQiEg0El9_3),.clk(gclk));
	jdff dff_B_sJ1C3hQo8_3(.din(w_dff_B_dQiEg0El9_3),.dout(w_dff_B_sJ1C3hQo8_3),.clk(gclk));
	jdff dff_B_gaPX4nAc7_3(.din(w_dff_B_sJ1C3hQo8_3),.dout(w_dff_B_gaPX4nAc7_3),.clk(gclk));
	jdff dff_B_djOsCc3g3_3(.din(w_dff_B_gaPX4nAc7_3),.dout(w_dff_B_djOsCc3g3_3),.clk(gclk));
	jdff dff_B_FHX8TLny0_1(.din(n1230),.dout(w_dff_B_FHX8TLny0_1),.clk(gclk));
	jdff dff_B_P19qavdH1_1(.din(w_dff_B_FHX8TLny0_1),.dout(w_dff_B_P19qavdH1_1),.clk(gclk));
	jdff dff_B_ycbutOvK2_1(.din(w_dff_B_P19qavdH1_1),.dout(w_dff_B_ycbutOvK2_1),.clk(gclk));
	jdff dff_B_Soo3w26k1_1(.din(w_dff_B_ycbutOvK2_1),.dout(w_dff_B_Soo3w26k1_1),.clk(gclk));
	jdff dff_B_7pt7jynQ8_1(.din(w_dff_B_Soo3w26k1_1),.dout(w_dff_B_7pt7jynQ8_1),.clk(gclk));
	jdff dff_B_mZSUNb9g1_1(.din(w_dff_B_7pt7jynQ8_1),.dout(w_dff_B_mZSUNb9g1_1),.clk(gclk));
	jdff dff_B_NBxSAoRi8_1(.din(w_dff_B_mZSUNb9g1_1),.dout(w_dff_B_NBxSAoRi8_1),.clk(gclk));
	jdff dff_B_n9wQfuIa9_1(.din(w_dff_B_NBxSAoRi8_1),.dout(w_dff_B_n9wQfuIa9_1),.clk(gclk));
	jdff dff_B_njhLuD006_1(.din(w_dff_B_n9wQfuIa9_1),.dout(w_dff_B_njhLuD006_1),.clk(gclk));
	jdff dff_B_SohIp7eS4_1(.din(w_dff_B_njhLuD006_1),.dout(w_dff_B_SohIp7eS4_1),.clk(gclk));
	jdff dff_B_VEGbVZ7T5_1(.din(w_dff_B_SohIp7eS4_1),.dout(w_dff_B_VEGbVZ7T5_1),.clk(gclk));
	jdff dff_B_hel2dOG81_1(.din(w_dff_B_VEGbVZ7T5_1),.dout(w_dff_B_hel2dOG81_1),.clk(gclk));
	jdff dff_B_tX8kMrfL6_1(.din(w_dff_B_hel2dOG81_1),.dout(w_dff_B_tX8kMrfL6_1),.clk(gclk));
	jdff dff_B_mlc6LtcC8_1(.din(w_dff_B_tX8kMrfL6_1),.dout(w_dff_B_mlc6LtcC8_1),.clk(gclk));
	jdff dff_B_5faaRwDs5_1(.din(w_dff_B_mlc6LtcC8_1),.dout(w_dff_B_5faaRwDs5_1),.clk(gclk));
	jdff dff_B_HTpe1VCg2_1(.din(w_dff_B_5faaRwDs5_1),.dout(w_dff_B_HTpe1VCg2_1),.clk(gclk));
	jdff dff_B_0Z5IiwPq7_1(.din(w_dff_B_HTpe1VCg2_1),.dout(w_dff_B_0Z5IiwPq7_1),.clk(gclk));
	jdff dff_B_BjCTQoto0_1(.din(n1232),.dout(w_dff_B_BjCTQoto0_1),.clk(gclk));
	jdff dff_B_VckX4ovK6_1(.din(w_dff_B_BjCTQoto0_1),.dout(w_dff_B_VckX4ovK6_1),.clk(gclk));
	jdff dff_B_MbvjTpVM5_1(.din(w_dff_B_VckX4ovK6_1),.dout(w_dff_B_MbvjTpVM5_1),.clk(gclk));
	jdff dff_B_LA1x1T553_1(.din(w_dff_B_MbvjTpVM5_1),.dout(w_dff_B_LA1x1T553_1),.clk(gclk));
	jdff dff_B_DEk286bu7_1(.din(w_dff_B_LA1x1T553_1),.dout(w_dff_B_DEk286bu7_1),.clk(gclk));
	jdff dff_B_9V0H138A9_1(.din(w_dff_B_DEk286bu7_1),.dout(w_dff_B_9V0H138A9_1),.clk(gclk));
	jdff dff_B_Ghu6kiR09_1(.din(w_dff_B_9V0H138A9_1),.dout(w_dff_B_Ghu6kiR09_1),.clk(gclk));
	jdff dff_B_L9lWMhdF2_1(.din(w_dff_B_Ghu6kiR09_1),.dout(w_dff_B_L9lWMhdF2_1),.clk(gclk));
	jdff dff_B_o8GKBQRI7_1(.din(w_dff_B_L9lWMhdF2_1),.dout(w_dff_B_o8GKBQRI7_1),.clk(gclk));
	jdff dff_B_iWhCo6B03_1(.din(w_dff_B_o8GKBQRI7_1),.dout(w_dff_B_iWhCo6B03_1),.clk(gclk));
	jdff dff_B_i48UCTAL8_1(.din(w_dff_B_iWhCo6B03_1),.dout(w_dff_B_i48UCTAL8_1),.clk(gclk));
	jdff dff_B_E104wsN56_1(.din(w_dff_B_i48UCTAL8_1),.dout(w_dff_B_E104wsN56_1),.clk(gclk));
	jdff dff_B_GCUTKeC38_1(.din(n937),.dout(w_dff_B_GCUTKeC38_1),.clk(gclk));
	jdff dff_B_pdUuINJl0_1(.din(w_dff_B_GCUTKeC38_1),.dout(w_dff_B_pdUuINJl0_1),.clk(gclk));
	jdff dff_B_UpfYWGsR2_1(.din(w_dff_B_pdUuINJl0_1),.dout(w_dff_B_UpfYWGsR2_1),.clk(gclk));
	jdff dff_B_K3RuSd0b4_1(.din(w_dff_B_UpfYWGsR2_1),.dout(w_dff_B_K3RuSd0b4_1),.clk(gclk));
	jdff dff_B_4gLCdTGb0_1(.din(w_dff_B_K3RuSd0b4_1),.dout(w_dff_B_4gLCdTGb0_1),.clk(gclk));
	jdff dff_B_pOTZXhRw8_1(.din(w_dff_B_4gLCdTGb0_1),.dout(w_dff_B_pOTZXhRw8_1),.clk(gclk));
	jdff dff_B_TULGqpbe4_1(.din(w_dff_B_pOTZXhRw8_1),.dout(w_dff_B_TULGqpbe4_1),.clk(gclk));
	jdff dff_B_r2KtQKQg4_1(.din(w_dff_B_TULGqpbe4_1),.dout(w_dff_B_r2KtQKQg4_1),.clk(gclk));
	jdff dff_B_rLWnffD82_1(.din(w_dff_B_r2KtQKQg4_1),.dout(w_dff_B_rLWnffD82_1),.clk(gclk));
	jdff dff_B_pJBymsxM6_1(.din(w_dff_B_rLWnffD82_1),.dout(w_dff_B_pJBymsxM6_1),.clk(gclk));
	jdff dff_B_ulWuoMYT0_1(.din(w_dff_B_pJBymsxM6_1),.dout(w_dff_B_ulWuoMYT0_1),.clk(gclk));
	jdff dff_B_1etY6Mwd5_0(.din(n869),.dout(w_dff_B_1etY6Mwd5_0),.clk(gclk));
	jdff dff_B_GEUE8hrs9_1(.din(n866),.dout(w_dff_B_GEUE8hrs9_1),.clk(gclk));
	jdff dff_B_9UXiCv0m5_1(.din(w_dff_B_GEUE8hrs9_1),.dout(w_dff_B_9UXiCv0m5_1),.clk(gclk));
	jdff dff_A_zhbpJqqR3_1(.dout(w_G4_0[1]),.din(w_dff_A_zhbpJqqR3_1),.clk(gclk));
	jdff dff_B_Djb85jzw6_3(.din(G4),.dout(w_dff_B_Djb85jzw6_3),.clk(gclk));
	jdff dff_B_XbMfPNC78_3(.din(w_dff_B_Djb85jzw6_3),.dout(w_dff_B_XbMfPNC78_3),.clk(gclk));
	jdff dff_B_kXpySNY15_3(.din(w_dff_B_XbMfPNC78_3),.dout(w_dff_B_kXpySNY15_3),.clk(gclk));
	jdff dff_B_7lgsNG6L1_3(.din(w_dff_B_kXpySNY15_3),.dout(w_dff_B_7lgsNG6L1_3),.clk(gclk));
	jdff dff_B_3BFNaT9z0_3(.din(w_dff_B_7lgsNG6L1_3),.dout(w_dff_B_3BFNaT9z0_3),.clk(gclk));
	jdff dff_A_nshC9MZh4_0(.dout(w_n1201_0[0]),.din(w_dff_A_nshC9MZh4_0),.clk(gclk));
	jdff dff_A_ZLrIieCK1_1(.dout(w_n1201_0[1]),.din(w_dff_A_ZLrIieCK1_1),.clk(gclk));
	jdff dff_A_Tjcoy3949_1(.dout(w_dff_A_ZLrIieCK1_1),.din(w_dff_A_Tjcoy3949_1),.clk(gclk));
	jdff dff_B_6soiylNA4_3(.din(n1201),.dout(w_dff_B_6soiylNA4_3),.clk(gclk));
	jdff dff_B_gaxXnFkz7_3(.din(w_dff_B_6soiylNA4_3),.dout(w_dff_B_gaxXnFkz7_3),.clk(gclk));
	jdff dff_B_D6GWk81n4_3(.din(w_dff_B_gaxXnFkz7_3),.dout(w_dff_B_D6GWk81n4_3),.clk(gclk));
	jdff dff_B_hKojJ9Rp0_3(.din(w_dff_B_D6GWk81n4_3),.dout(w_dff_B_hKojJ9Rp0_3),.clk(gclk));
	jdff dff_B_KLBHPtCb3_3(.din(w_dff_B_hKojJ9Rp0_3),.dout(w_dff_B_KLBHPtCb3_3),.clk(gclk));
	jdff dff_B_boVhpqj27_3(.din(w_dff_B_KLBHPtCb3_3),.dout(w_dff_B_boVhpqj27_3),.clk(gclk));
	jdff dff_B_x6UQqVXX7_3(.din(w_dff_B_boVhpqj27_3),.dout(w_dff_B_x6UQqVXX7_3),.clk(gclk));
	jdff dff_B_7XORGzGK5_3(.din(w_dff_B_x6UQqVXX7_3),.dout(w_dff_B_7XORGzGK5_3),.clk(gclk));
	jdff dff_B_nu7RB4Nl2_3(.din(w_dff_B_7XORGzGK5_3),.dout(w_dff_B_nu7RB4Nl2_3),.clk(gclk));
	jdff dff_B_XZuJ79wq8_3(.din(w_dff_B_nu7RB4Nl2_3),.dout(w_dff_B_XZuJ79wq8_3),.clk(gclk));
	jdff dff_B_TJkDqrhs3_3(.din(w_dff_B_XZuJ79wq8_3),.dout(w_dff_B_TJkDqrhs3_3),.clk(gclk));
	jdff dff_B_3PiQHyt39_3(.din(w_dff_B_TJkDqrhs3_3),.dout(w_dff_B_3PiQHyt39_3),.clk(gclk));
	jdff dff_B_oqp7mgxB8_3(.din(w_dff_B_3PiQHyt39_3),.dout(w_dff_B_oqp7mgxB8_3),.clk(gclk));
	jdff dff_B_G1XF9B541_3(.din(w_dff_B_oqp7mgxB8_3),.dout(w_dff_B_G1XF9B541_3),.clk(gclk));
	jdff dff_B_Vg4hOFcp5_3(.din(w_dff_B_G1XF9B541_3),.dout(w_dff_B_Vg4hOFcp5_3),.clk(gclk));
	jdff dff_A_LypQKKcW0_0(.dout(w_G4092_5[0]),.din(w_dff_A_LypQKKcW0_0),.clk(gclk));
	jdff dff_A_yXRHn23c6_0(.dout(w_dff_A_LypQKKcW0_0),.din(w_dff_A_yXRHn23c6_0),.clk(gclk));
	jdff dff_A_kAPst4rG7_0(.dout(w_dff_A_yXRHn23c6_0),.din(w_dff_A_kAPst4rG7_0),.clk(gclk));
	jdff dff_A_olHE7vfl9_0(.dout(w_dff_A_kAPst4rG7_0),.din(w_dff_A_olHE7vfl9_0),.clk(gclk));
	jdff dff_A_LWuJLPGe4_0(.dout(w_dff_A_olHE7vfl9_0),.din(w_dff_A_LWuJLPGe4_0),.clk(gclk));
	jdff dff_A_93243qg33_0(.dout(w_dff_A_LWuJLPGe4_0),.din(w_dff_A_93243qg33_0),.clk(gclk));
	jdff dff_A_L9n2n8oJ8_1(.dout(w_G4092_5[1]),.din(w_dff_A_L9n2n8oJ8_1),.clk(gclk));
	jdff dff_A_edaGDRxl6_1(.dout(w_dff_A_L9n2n8oJ8_1),.din(w_dff_A_edaGDRxl6_1),.clk(gclk));
	jdff dff_A_Z4Y8e3Fm2_1(.dout(w_dff_A_edaGDRxl6_1),.din(w_dff_A_Z4Y8e3Fm2_1),.clk(gclk));
	jdff dff_A_2jivuVoV2_1(.dout(w_dff_A_Z4Y8e3Fm2_1),.din(w_dff_A_2jivuVoV2_1),.clk(gclk));
	jdff dff_A_vYseTm2Q7_1(.dout(w_dff_A_2jivuVoV2_1),.din(w_dff_A_vYseTm2Q7_1),.clk(gclk));
	jdff dff_A_N2iAANj73_1(.dout(w_dff_A_vYseTm2Q7_1),.din(w_dff_A_N2iAANj73_1),.clk(gclk));
	jdff dff_A_tdTttx1A4_0(.dout(w_n749_7[0]),.din(w_dff_A_tdTttx1A4_0),.clk(gclk));
	jdff dff_A_6TS6vlq43_0(.dout(w_dff_A_tdTttx1A4_0),.din(w_dff_A_6TS6vlq43_0),.clk(gclk));
	jdff dff_A_UnODfP1e7_0(.dout(w_dff_A_6TS6vlq43_0),.din(w_dff_A_UnODfP1e7_0),.clk(gclk));
	jdff dff_A_AA0Aec4E5_0(.dout(w_dff_A_UnODfP1e7_0),.din(w_dff_A_AA0Aec4E5_0),.clk(gclk));
	jdff dff_A_pg1yx1tx3_0(.dout(w_dff_A_AA0Aec4E5_0),.din(w_dff_A_pg1yx1tx3_0),.clk(gclk));
	jdff dff_A_vqeYpe6u4_0(.dout(w_dff_A_pg1yx1tx3_0),.din(w_dff_A_vqeYpe6u4_0),.clk(gclk));
	jdff dff_A_T1XhDIww2_0(.dout(w_dff_A_vqeYpe6u4_0),.din(w_dff_A_T1XhDIww2_0),.clk(gclk));
	jdff dff_A_riKcW56x8_0(.dout(w_dff_A_T1XhDIww2_0),.din(w_dff_A_riKcW56x8_0),.clk(gclk));
	jdff dff_A_nmRawhVX0_0(.dout(w_dff_A_riKcW56x8_0),.din(w_dff_A_nmRawhVX0_0),.clk(gclk));
	jdff dff_A_orhdBHcl5_0(.dout(w_dff_A_nmRawhVX0_0),.din(w_dff_A_orhdBHcl5_0),.clk(gclk));
	jdff dff_A_KUKgTNlP7_0(.dout(w_dff_A_orhdBHcl5_0),.din(w_dff_A_KUKgTNlP7_0),.clk(gclk));
	jdff dff_A_jhT5jWgK2_0(.dout(w_dff_A_KUKgTNlP7_0),.din(w_dff_A_jhT5jWgK2_0),.clk(gclk));
	jdff dff_A_fZvtdc804_0(.dout(w_n749_2[0]),.din(w_dff_A_fZvtdc804_0),.clk(gclk));
	jdff dff_A_UGEY9o3W6_0(.dout(w_dff_A_fZvtdc804_0),.din(w_dff_A_UGEY9o3W6_0),.clk(gclk));
	jdff dff_A_2WSEciTN5_1(.dout(w_n749_2[1]),.din(w_dff_A_2WSEciTN5_1),.clk(gclk));
	jdff dff_A_r6mjsyH68_1(.dout(w_dff_A_2WSEciTN5_1),.din(w_dff_A_r6mjsyH68_1),.clk(gclk));
	jdff dff_B_Ehju4Z324_1(.din(G115),.dout(w_dff_B_Ehju4Z324_1),.clk(gclk));
	jdff dff_B_uKlhyMAY6_1(.din(w_dff_B_Ehju4Z324_1),.dout(w_dff_B_uKlhyMAY6_1),.clk(gclk));
	jdff dff_B_wDrfRkwT3_0(.din(n1505),.dout(w_dff_B_wDrfRkwT3_0),.clk(gclk));
	jdff dff_B_Cwc16hRW5_0(.din(w_dff_B_wDrfRkwT3_0),.dout(w_dff_B_Cwc16hRW5_0),.clk(gclk));
	jdff dff_B_vWWfOqqQ9_0(.din(w_dff_B_Cwc16hRW5_0),.dout(w_dff_B_vWWfOqqQ9_0),.clk(gclk));
	jdff dff_B_D5UDEj6N8_0(.din(w_dff_B_vWWfOqqQ9_0),.dout(w_dff_B_D5UDEj6N8_0),.clk(gclk));
	jdff dff_B_bzNCjmpl3_0(.din(w_dff_B_D5UDEj6N8_0),.dout(w_dff_B_bzNCjmpl3_0),.clk(gclk));
	jdff dff_B_dLbIVf7M8_0(.din(w_dff_B_bzNCjmpl3_0),.dout(w_dff_B_dLbIVf7M8_0),.clk(gclk));
	jdff dff_B_3o1tM25u3_0(.din(w_dff_B_dLbIVf7M8_0),.dout(w_dff_B_3o1tM25u3_0),.clk(gclk));
	jdff dff_B_SOWLTAqs1_0(.din(w_dff_B_3o1tM25u3_0),.dout(w_dff_B_SOWLTAqs1_0),.clk(gclk));
	jdff dff_B_L4TOTHkU6_0(.din(w_dff_B_SOWLTAqs1_0),.dout(w_dff_B_L4TOTHkU6_0),.clk(gclk));
	jdff dff_B_AvUsMNqQ5_0(.din(w_dff_B_L4TOTHkU6_0),.dout(w_dff_B_AvUsMNqQ5_0),.clk(gclk));
	jdff dff_B_qosWfwVb2_0(.din(w_dff_B_AvUsMNqQ5_0),.dout(w_dff_B_qosWfwVb2_0),.clk(gclk));
	jdff dff_B_0EAHIAn80_0(.din(w_dff_B_qosWfwVb2_0),.dout(w_dff_B_0EAHIAn80_0),.clk(gclk));
	jdff dff_B_4saqOU3Y3_0(.din(w_dff_B_0EAHIAn80_0),.dout(w_dff_B_4saqOU3Y3_0),.clk(gclk));
	jdff dff_B_Ec75XCn20_0(.din(w_dff_B_4saqOU3Y3_0),.dout(w_dff_B_Ec75XCn20_0),.clk(gclk));
	jdff dff_B_HvZxSwsH1_0(.din(w_dff_B_Ec75XCn20_0),.dout(w_dff_B_HvZxSwsH1_0),.clk(gclk));
	jdff dff_B_1Y5pUuUD6_0(.din(w_dff_B_HvZxSwsH1_0),.dout(w_dff_B_1Y5pUuUD6_0),.clk(gclk));
	jdff dff_B_ow9X3H7R6_0(.din(w_dff_B_1Y5pUuUD6_0),.dout(w_dff_B_ow9X3H7R6_0),.clk(gclk));
	jdff dff_B_us0caNch4_1(.din(G120),.dout(w_dff_B_us0caNch4_1),.clk(gclk));
	jdff dff_B_OIAyBtWZ3_1(.din(w_dff_B_us0caNch4_1),.dout(w_dff_B_OIAyBtWZ3_1),.clk(gclk));
	jdff dff_B_qS653Y2i8_1(.din(w_dff_B_OIAyBtWZ3_1),.dout(w_dff_B_qS653Y2i8_1),.clk(gclk));
	jdff dff_B_o2XB3q0z2_0(.din(n1666),.dout(w_dff_B_o2XB3q0z2_0),.clk(gclk));
	jdff dff_B_N02CtFAU5_0(.din(w_dff_B_o2XB3q0z2_0),.dout(w_dff_B_N02CtFAU5_0),.clk(gclk));
	jdff dff_B_y3ymCFBe5_0(.din(w_dff_B_N02CtFAU5_0),.dout(w_dff_B_y3ymCFBe5_0),.clk(gclk));
	jdff dff_B_N5YZXX2n3_0(.din(w_dff_B_y3ymCFBe5_0),.dout(w_dff_B_N5YZXX2n3_0),.clk(gclk));
	jdff dff_B_GVlPamiQ3_0(.din(w_dff_B_N5YZXX2n3_0),.dout(w_dff_B_GVlPamiQ3_0),.clk(gclk));
	jdff dff_B_BIpqgLrW3_0(.din(w_dff_B_GVlPamiQ3_0),.dout(w_dff_B_BIpqgLrW3_0),.clk(gclk));
	jdff dff_B_gFIt59JH6_0(.din(w_dff_B_BIpqgLrW3_0),.dout(w_dff_B_gFIt59JH6_0),.clk(gclk));
	jdff dff_B_cNBuyqeU3_0(.din(w_dff_B_gFIt59JH6_0),.dout(w_dff_B_cNBuyqeU3_0),.clk(gclk));
	jdff dff_B_t8gWkXLY8_0(.din(w_dff_B_cNBuyqeU3_0),.dout(w_dff_B_t8gWkXLY8_0),.clk(gclk));
	jdff dff_B_SPPxYmft4_0(.din(w_dff_B_t8gWkXLY8_0),.dout(w_dff_B_SPPxYmft4_0),.clk(gclk));
	jdff dff_B_JMA2Ojso9_0(.din(w_dff_B_SPPxYmft4_0),.dout(w_dff_B_JMA2Ojso9_0),.clk(gclk));
	jdff dff_B_bdhzgnpS6_0(.din(w_dff_B_JMA2Ojso9_0),.dout(w_dff_B_bdhzgnpS6_0),.clk(gclk));
	jdff dff_B_5yvKG2eJ0_0(.din(w_dff_B_bdhzgnpS6_0),.dout(w_dff_B_5yvKG2eJ0_0),.clk(gclk));
	jdff dff_B_I2IkDyHH9_0(.din(w_dff_B_5yvKG2eJ0_0),.dout(w_dff_B_I2IkDyHH9_0),.clk(gclk));
	jdff dff_B_61X5ZuyU4_0(.din(w_dff_B_I2IkDyHH9_0),.dout(w_dff_B_61X5ZuyU4_0),.clk(gclk));
	jdff dff_B_NaYOdTpP1_0(.din(w_dff_B_61X5ZuyU4_0),.dout(w_dff_B_NaYOdTpP1_0),.clk(gclk));
	jdff dff_B_9NRyjmDE9_0(.din(w_dff_B_NaYOdTpP1_0),.dout(w_dff_B_9NRyjmDE9_0),.clk(gclk));
	jdff dff_B_PBRsEGmR6_1(.din(G118),.dout(w_dff_B_PBRsEGmR6_1),.clk(gclk));
	jdff dff_B_1u8wWBmn5_1(.din(w_dff_B_PBRsEGmR6_1),.dout(w_dff_B_1u8wWBmn5_1),.clk(gclk));
	jdff dff_B_E0dWacZS0_1(.din(w_dff_B_1u8wWBmn5_1),.dout(w_dff_B_E0dWacZS0_1),.clk(gclk));
	jdff dff_A_YlAgmg6T7_0(.dout(w_G4092_9[0]),.din(w_dff_A_YlAgmg6T7_0),.clk(gclk));
	jdff dff_A_rcfcSIjf5_0(.dout(w_dff_A_YlAgmg6T7_0),.din(w_dff_A_rcfcSIjf5_0),.clk(gclk));
	jdff dff_A_Jn97mrZK5_0(.dout(w_dff_A_rcfcSIjf5_0),.din(w_dff_A_Jn97mrZK5_0),.clk(gclk));
	jdff dff_A_C4NNP8Xo9_0(.dout(w_dff_A_Jn97mrZK5_0),.din(w_dff_A_C4NNP8Xo9_0),.clk(gclk));
	jdff dff_A_5lvsBwnu3_0(.dout(w_dff_A_C4NNP8Xo9_0),.din(w_dff_A_5lvsBwnu3_0),.clk(gclk));
	jdff dff_A_xfi47aKt6_1(.dout(w_G4092_9[1]),.din(w_dff_A_xfi47aKt6_1),.clk(gclk));
	jdff dff_A_XX8s0kTl5_1(.dout(w_dff_A_xfi47aKt6_1),.din(w_dff_A_XX8s0kTl5_1),.clk(gclk));
	jdff dff_A_wcH6QTuZ3_1(.dout(w_dff_A_XX8s0kTl5_1),.din(w_dff_A_wcH6QTuZ3_1),.clk(gclk));
	jdff dff_A_R2cCntsR9_1(.dout(w_dff_A_wcH6QTuZ3_1),.din(w_dff_A_R2cCntsR9_1),.clk(gclk));
	jdff dff_A_2ThLU8My3_0(.dout(w_G4092_2[0]),.din(w_dff_A_2ThLU8My3_0),.clk(gclk));
	jdff dff_A_PUvMD4Qh7_0(.dout(w_dff_A_2ThLU8My3_0),.din(w_dff_A_PUvMD4Qh7_0),.clk(gclk));
	jdff dff_A_0T5gnU6g4_0(.dout(w_dff_A_PUvMD4Qh7_0),.din(w_dff_A_0T5gnU6g4_0),.clk(gclk));
	jdff dff_A_RIoXXCcc6_0(.dout(w_dff_A_0T5gnU6g4_0),.din(w_dff_A_RIoXXCcc6_0),.clk(gclk));
	jdff dff_A_Rcqv1pnE6_0(.dout(w_dff_A_RIoXXCcc6_0),.din(w_dff_A_Rcqv1pnE6_0),.clk(gclk));
	jdff dff_A_mFeMHTtF2_1(.dout(w_G4092_2[1]),.din(w_dff_A_mFeMHTtF2_1),.clk(gclk));
	jdff dff_A_v7kFF0zp0_1(.dout(w_dff_A_mFeMHTtF2_1),.din(w_dff_A_v7kFF0zp0_1),.clk(gclk));
	jdff dff_A_KkthLwDo4_1(.dout(w_dff_A_v7kFF0zp0_1),.din(w_dff_A_KkthLwDo4_1),.clk(gclk));
	jdff dff_A_u4fEX5Gh2_1(.dout(w_dff_A_KkthLwDo4_1),.din(w_dff_A_u4fEX5Gh2_1),.clk(gclk));
	jdff dff_A_6vxKppbj8_0(.dout(w_n749_13[0]),.din(w_dff_A_6vxKppbj8_0),.clk(gclk));
	jdff dff_A_Q1y0rw1J0_0(.dout(w_dff_A_6vxKppbj8_0),.din(w_dff_A_Q1y0rw1J0_0),.clk(gclk));
	jdff dff_A_MYjoLYpB8_0(.dout(w_dff_A_Q1y0rw1J0_0),.din(w_dff_A_MYjoLYpB8_0),.clk(gclk));
	jdff dff_B_zEo4q6Xh3_1(.din(n1671),.dout(w_dff_B_zEo4q6Xh3_1),.clk(gclk));
	jdff dff_B_BJBS0wp33_1(.din(w_dff_B_zEo4q6Xh3_1),.dout(w_dff_B_BJBS0wp33_1),.clk(gclk));
	jdff dff_B_nsg6w8Jg1_1(.din(w_dff_B_BJBS0wp33_1),.dout(w_dff_B_nsg6w8Jg1_1),.clk(gclk));
	jdff dff_B_9DeTDEkl1_1(.din(w_dff_B_nsg6w8Jg1_1),.dout(w_dff_B_9DeTDEkl1_1),.clk(gclk));
	jdff dff_B_eqHr8K7Z4_1(.din(w_dff_B_9DeTDEkl1_1),.dout(w_dff_B_eqHr8K7Z4_1),.clk(gclk));
	jdff dff_B_m6uGQahr0_1(.din(w_dff_B_eqHr8K7Z4_1),.dout(w_dff_B_m6uGQahr0_1),.clk(gclk));
	jdff dff_B_w4OiuBEM4_1(.din(w_dff_B_m6uGQahr0_1),.dout(w_dff_B_w4OiuBEM4_1),.clk(gclk));
	jdff dff_B_uGzj4GnF2_1(.din(w_dff_B_w4OiuBEM4_1),.dout(w_dff_B_uGzj4GnF2_1),.clk(gclk));
	jdff dff_B_Cu8AVbP31_1(.din(w_dff_B_uGzj4GnF2_1),.dout(w_dff_B_Cu8AVbP31_1),.clk(gclk));
	jdff dff_B_3T8p3AbB2_1(.din(w_dff_B_Cu8AVbP31_1),.dout(w_dff_B_3T8p3AbB2_1),.clk(gclk));
	jdff dff_B_bSBCFu0d3_1(.din(w_dff_B_3T8p3AbB2_1),.dout(w_dff_B_bSBCFu0d3_1),.clk(gclk));
	jdff dff_B_cMV8N3sX5_1(.din(w_dff_B_bSBCFu0d3_1),.dout(w_dff_B_cMV8N3sX5_1),.clk(gclk));
	jdff dff_B_8oSCkhnx1_1(.din(w_dff_B_cMV8N3sX5_1),.dout(w_dff_B_8oSCkhnx1_1),.clk(gclk));
	jdff dff_B_pvphTkoP5_1(.din(w_dff_B_8oSCkhnx1_1),.dout(w_dff_B_pvphTkoP5_1),.clk(gclk));
	jdff dff_B_P2UAXcJf8_1(.din(w_dff_B_pvphTkoP5_1),.dout(w_dff_B_P2UAXcJf8_1),.clk(gclk));
	jdff dff_B_d6bv0RBw7_1(.din(w_dff_B_P2UAXcJf8_1),.dout(w_dff_B_d6bv0RBw7_1),.clk(gclk));
	jdff dff_B_YPFyJM4S1_1(.din(w_dff_B_d6bv0RBw7_1),.dout(w_dff_B_YPFyJM4S1_1),.clk(gclk));
	jdff dff_B_eiqe9rVO8_1(.din(w_dff_B_YPFyJM4S1_1),.dout(w_dff_B_eiqe9rVO8_1),.clk(gclk));
	jdff dff_B_u3QlNxvx7_1(.din(w_dff_B_eiqe9rVO8_1),.dout(w_dff_B_u3QlNxvx7_1),.clk(gclk));
	jdff dff_B_tirUx62I2_1(.din(w_dff_B_u3QlNxvx7_1),.dout(w_dff_B_tirUx62I2_1),.clk(gclk));
	jdff dff_B_rxo2Dayk1_1(.din(w_dff_B_tirUx62I2_1),.dout(w_dff_B_rxo2Dayk1_1),.clk(gclk));
	jdff dff_B_DQdEZMtx8_1(.din(w_dff_B_rxo2Dayk1_1),.dout(w_dff_B_DQdEZMtx8_1),.clk(gclk));
	jdff dff_B_Xab86eH79_1(.din(n1676),.dout(w_dff_B_Xab86eH79_1),.clk(gclk));
	jdff dff_A_hdXM7sbV1_1(.dout(w_n800_1[1]),.din(w_dff_A_hdXM7sbV1_1),.clk(gclk));
	jdff dff_A_Z0m7DK4o2_1(.dout(w_dff_A_hdXM7sbV1_1),.din(w_dff_A_Z0m7DK4o2_1),.clk(gclk));
	jdff dff_A_Q03PM3lt4_1(.dout(w_dff_A_Z0m7DK4o2_1),.din(w_dff_A_Q03PM3lt4_1),.clk(gclk));
	jdff dff_A_YmGFXRcK2_1(.dout(w_dff_A_Q03PM3lt4_1),.din(w_dff_A_YmGFXRcK2_1),.clk(gclk));
	jdff dff_A_v0v4KUoW6_1(.dout(w_dff_A_YmGFXRcK2_1),.din(w_dff_A_v0v4KUoW6_1),.clk(gclk));
	jdff dff_A_lEOxaR872_1(.dout(w_dff_A_v0v4KUoW6_1),.din(w_dff_A_lEOxaR872_1),.clk(gclk));
	jdff dff_A_uFJdQoKg6_1(.dout(w_dff_A_lEOxaR872_1),.din(w_dff_A_uFJdQoKg6_1),.clk(gclk));
	jdff dff_A_hWrlshFl1_1(.dout(w_dff_A_uFJdQoKg6_1),.din(w_dff_A_hWrlshFl1_1),.clk(gclk));
	jdff dff_A_7UY9nmdC8_1(.dout(w_dff_A_hWrlshFl1_1),.din(w_dff_A_7UY9nmdC8_1),.clk(gclk));
	jdff dff_A_niaUuaPX1_1(.dout(w_dff_A_7UY9nmdC8_1),.din(w_dff_A_niaUuaPX1_1),.clk(gclk));
	jdff dff_A_sKnW5gSz2_1(.dout(w_dff_A_niaUuaPX1_1),.din(w_dff_A_sKnW5gSz2_1),.clk(gclk));
	jdff dff_A_qh4CeztD9_1(.dout(w_dff_A_sKnW5gSz2_1),.din(w_dff_A_qh4CeztD9_1),.clk(gclk));
	jdff dff_A_ygC8iK3D9_1(.dout(w_dff_A_qh4CeztD9_1),.din(w_dff_A_ygC8iK3D9_1),.clk(gclk));
	jdff dff_A_29YK8VA16_1(.dout(w_dff_A_ygC8iK3D9_1),.din(w_dff_A_29YK8VA16_1),.clk(gclk));
	jdff dff_A_FM70XG8Q0_2(.dout(w_n800_1[2]),.din(w_dff_A_FM70XG8Q0_2),.clk(gclk));
	jdff dff_A_5HkoReu22_2(.dout(w_dff_A_FM70XG8Q0_2),.din(w_dff_A_5HkoReu22_2),.clk(gclk));
	jdff dff_A_8YKp4dCs0_2(.dout(w_dff_A_5HkoReu22_2),.din(w_dff_A_8YKp4dCs0_2),.clk(gclk));
	jdff dff_A_PdafN9kM7_2(.dout(w_dff_A_8YKp4dCs0_2),.din(w_dff_A_PdafN9kM7_2),.clk(gclk));
	jdff dff_A_tSoASTp51_2(.dout(w_dff_A_PdafN9kM7_2),.din(w_dff_A_tSoASTp51_2),.clk(gclk));
	jdff dff_A_l3SVPDTu0_2(.dout(w_dff_A_tSoASTp51_2),.din(w_dff_A_l3SVPDTu0_2),.clk(gclk));
	jdff dff_A_NCeIZyn30_2(.dout(w_dff_A_l3SVPDTu0_2),.din(w_dff_A_NCeIZyn30_2),.clk(gclk));
	jdff dff_A_c33zlPMx0_2(.dout(w_dff_A_NCeIZyn30_2),.din(w_dff_A_c33zlPMx0_2),.clk(gclk));
	jdff dff_A_CKntm3vl8_2(.dout(w_dff_A_c33zlPMx0_2),.din(w_dff_A_CKntm3vl8_2),.clk(gclk));
	jdff dff_A_Pbl6qVni4_2(.dout(w_dff_A_CKntm3vl8_2),.din(w_dff_A_Pbl6qVni4_2),.clk(gclk));
	jdff dff_A_4ukLVA8O8_1(.dout(w_n800_0[1]),.din(w_dff_A_4ukLVA8O8_1),.clk(gclk));
	jdff dff_A_8FvYFgJ17_1(.dout(w_dff_A_4ukLVA8O8_1),.din(w_dff_A_8FvYFgJ17_1),.clk(gclk));
	jdff dff_A_cymLraMl8_1(.dout(w_dff_A_8FvYFgJ17_1),.din(w_dff_A_cymLraMl8_1),.clk(gclk));
	jdff dff_A_APp8NyV30_1(.dout(w_dff_A_cymLraMl8_1),.din(w_dff_A_APp8NyV30_1),.clk(gclk));
	jdff dff_A_vADtSfHk0_1(.dout(w_dff_A_APp8NyV30_1),.din(w_dff_A_vADtSfHk0_1),.clk(gclk));
	jdff dff_A_iB6LAnTI1_1(.dout(w_dff_A_vADtSfHk0_1),.din(w_dff_A_iB6LAnTI1_1),.clk(gclk));
	jdff dff_A_C60DUzXr7_1(.dout(w_dff_A_iB6LAnTI1_1),.din(w_dff_A_C60DUzXr7_1),.clk(gclk));
	jdff dff_A_CP8EoBFH8_1(.dout(w_dff_A_C60DUzXr7_1),.din(w_dff_A_CP8EoBFH8_1),.clk(gclk));
	jdff dff_A_L2OZaSFY0_1(.dout(w_dff_A_CP8EoBFH8_1),.din(w_dff_A_L2OZaSFY0_1),.clk(gclk));
	jdff dff_A_yp4yISs39_1(.dout(w_dff_A_L2OZaSFY0_1),.din(w_dff_A_yp4yISs39_1),.clk(gclk));
	jdff dff_A_ChpFXZM95_1(.dout(w_dff_A_yp4yISs39_1),.din(w_dff_A_ChpFXZM95_1),.clk(gclk));
	jdff dff_A_cLxXia6N4_2(.dout(w_n800_0[2]),.din(w_dff_A_cLxXia6N4_2),.clk(gclk));
	jdff dff_A_BlkVTWEQ9_2(.dout(w_dff_A_cLxXia6N4_2),.din(w_dff_A_BlkVTWEQ9_2),.clk(gclk));
	jdff dff_A_WIcn31uy0_2(.dout(w_dff_A_BlkVTWEQ9_2),.din(w_dff_A_WIcn31uy0_2),.clk(gclk));
	jdff dff_A_6zlKOZOd4_2(.dout(w_dff_A_WIcn31uy0_2),.din(w_dff_A_6zlKOZOd4_2),.clk(gclk));
	jdff dff_B_ScrxC0ex8_3(.din(n800),.dout(w_dff_B_ScrxC0ex8_3),.clk(gclk));
	jdff dff_B_bF9HSW5h6_3(.din(w_dff_B_ScrxC0ex8_3),.dout(w_dff_B_bF9HSW5h6_3),.clk(gclk));
	jdff dff_B_iV8XZhOK8_3(.din(w_dff_B_bF9HSW5h6_3),.dout(w_dff_B_iV8XZhOK8_3),.clk(gclk));
	jdff dff_B_IgwPsuVZ1_3(.din(w_dff_B_iV8XZhOK8_3),.dout(w_dff_B_IgwPsuVZ1_3),.clk(gclk));
	jdff dff_B_pAHPjq7V4_3(.din(w_dff_B_IgwPsuVZ1_3),.dout(w_dff_B_pAHPjq7V4_3),.clk(gclk));
	jdff dff_B_7mfdTIcv8_3(.din(w_dff_B_pAHPjq7V4_3),.dout(w_dff_B_7mfdTIcv8_3),.clk(gclk));
	jdff dff_B_bDR0fVtB4_3(.din(w_dff_B_7mfdTIcv8_3),.dout(w_dff_B_bDR0fVtB4_3),.clk(gclk));
	jdff dff_B_3WtelaWZ0_3(.din(w_dff_B_bDR0fVtB4_3),.dout(w_dff_B_3WtelaWZ0_3),.clk(gclk));
	jdff dff_B_1YMFOaP55_3(.din(w_dff_B_3WtelaWZ0_3),.dout(w_dff_B_1YMFOaP55_3),.clk(gclk));
	jdff dff_A_uKSr5MXa6_0(.dout(w_G4087_4[0]),.din(w_dff_A_uKSr5MXa6_0),.clk(gclk));
	jdff dff_A_pPMSWfET9_1(.dout(w_G4087_4[1]),.din(w_dff_A_pPMSWfET9_1),.clk(gclk));
	jdff dff_B_wjVMUX9z6_1(.din(n1668),.dout(w_dff_B_wjVMUX9z6_1),.clk(gclk));
	jdff dff_B_F1BdJIRn7_1(.din(w_dff_B_wjVMUX9z6_1),.dout(w_dff_B_F1BdJIRn7_1),.clk(gclk));
	jdff dff_A_J7RpXy9j0_0(.dout(w_n797_3[0]),.din(w_dff_A_J7RpXy9j0_0),.clk(gclk));
	jdff dff_A_B2b2QXRq5_0(.dout(w_dff_A_J7RpXy9j0_0),.din(w_dff_A_B2b2QXRq5_0),.clk(gclk));
	jdff dff_A_U73T2Cer5_0(.dout(w_dff_A_B2b2QXRq5_0),.din(w_dff_A_U73T2Cer5_0),.clk(gclk));
	jdff dff_A_w39mU8Y99_0(.dout(w_dff_A_U73T2Cer5_0),.din(w_dff_A_w39mU8Y99_0),.clk(gclk));
	jdff dff_A_m15o0S1P9_0(.dout(w_dff_A_w39mU8Y99_0),.din(w_dff_A_m15o0S1P9_0),.clk(gclk));
	jdff dff_A_mcMP1zUM8_0(.dout(w_dff_A_m15o0S1P9_0),.din(w_dff_A_mcMP1zUM8_0),.clk(gclk));
	jdff dff_A_zjECLO450_0(.dout(w_dff_A_mcMP1zUM8_0),.din(w_dff_A_zjECLO450_0),.clk(gclk));
	jdff dff_A_aM0peksZ5_0(.dout(w_dff_A_zjECLO450_0),.din(w_dff_A_aM0peksZ5_0),.clk(gclk));
	jdff dff_A_FQZO09FO5_0(.dout(w_dff_A_aM0peksZ5_0),.din(w_dff_A_FQZO09FO5_0),.clk(gclk));
	jdff dff_A_Spd7vZn46_0(.dout(w_dff_A_FQZO09FO5_0),.din(w_dff_A_Spd7vZn46_0),.clk(gclk));
	jdff dff_A_bQitdwoY1_0(.dout(w_dff_A_Spd7vZn46_0),.din(w_dff_A_bQitdwoY1_0),.clk(gclk));
	jdff dff_A_oThGbyep6_0(.dout(w_dff_A_bQitdwoY1_0),.din(w_dff_A_oThGbyep6_0),.clk(gclk));
	jdff dff_A_BZXl5qNo8_0(.dout(w_dff_A_oThGbyep6_0),.din(w_dff_A_BZXl5qNo8_0),.clk(gclk));
	jdff dff_A_DR3dhzZL6_0(.dout(w_dff_A_BZXl5qNo8_0),.din(w_dff_A_DR3dhzZL6_0),.clk(gclk));
	jdff dff_A_0X6f479c5_0(.dout(w_dff_A_DR3dhzZL6_0),.din(w_dff_A_0X6f479c5_0),.clk(gclk));
	jdff dff_A_AN4zE28N9_0(.dout(w_dff_A_0X6f479c5_0),.din(w_dff_A_AN4zE28N9_0),.clk(gclk));
	jdff dff_A_M3BwlCt59_0(.dout(w_dff_A_AN4zE28N9_0),.din(w_dff_A_M3BwlCt59_0),.clk(gclk));
	jdff dff_A_RaZXe41y5_0(.dout(w_dff_A_M3BwlCt59_0),.din(w_dff_A_RaZXe41y5_0),.clk(gclk));
	jdff dff_A_ZTLypPDO1_0(.dout(w_dff_A_RaZXe41y5_0),.din(w_dff_A_ZTLypPDO1_0),.clk(gclk));
	jdff dff_A_557w5x5b3_0(.dout(w_dff_A_ZTLypPDO1_0),.din(w_dff_A_557w5x5b3_0),.clk(gclk));
	jdff dff_A_70LyU2fl4_0(.dout(w_dff_A_557w5x5b3_0),.din(w_dff_A_70LyU2fl4_0),.clk(gclk));
	jdff dff_A_ExNRHowj8_0(.dout(w_dff_A_70LyU2fl4_0),.din(w_dff_A_ExNRHowj8_0),.clk(gclk));
	jdff dff_A_9CG4UPxr9_1(.dout(w_G4088_9[1]),.din(w_dff_A_9CG4UPxr9_1),.clk(gclk));
	jdff dff_A_V1YRyjog0_1(.dout(w_dff_A_9CG4UPxr9_1),.din(w_dff_A_V1YRyjog0_1),.clk(gclk));
	jdff dff_A_NCDTHPr95_1(.dout(w_dff_A_V1YRyjog0_1),.din(w_dff_A_NCDTHPr95_1),.clk(gclk));
	jdff dff_A_wIyHRV9x1_1(.dout(w_dff_A_NCDTHPr95_1),.din(w_dff_A_wIyHRV9x1_1),.clk(gclk));
	jdff dff_A_zYyz2T3b6_1(.dout(w_dff_A_wIyHRV9x1_1),.din(w_dff_A_zYyz2T3b6_1),.clk(gclk));
	jdff dff_A_Jq3nLSms4_1(.dout(w_dff_A_zYyz2T3b6_1),.din(w_dff_A_Jq3nLSms4_1),.clk(gclk));
	jdff dff_A_SfRM7CcV4_1(.dout(w_dff_A_Jq3nLSms4_1),.din(w_dff_A_SfRM7CcV4_1),.clk(gclk));
	jdff dff_A_ouvJbN4a0_1(.dout(w_dff_A_SfRM7CcV4_1),.din(w_dff_A_ouvJbN4a0_1),.clk(gclk));
	jdff dff_A_F4a1JVaO5_1(.dout(w_dff_A_ouvJbN4a0_1),.din(w_dff_A_F4a1JVaO5_1),.clk(gclk));
	jdff dff_A_FjZ8h4rR6_1(.dout(w_G4087_1[1]),.din(w_dff_A_FjZ8h4rR6_1),.clk(gclk));
	jdff dff_A_qxidpLW09_1(.dout(w_dff_A_FjZ8h4rR6_1),.din(w_dff_A_qxidpLW09_1),.clk(gclk));
	jdff dff_A_EXoqS4CX2_2(.dout(w_G4087_1[2]),.din(w_dff_A_EXoqS4CX2_2),.clk(gclk));
	jdff dff_A_ZtjjC1cr6_1(.dout(w_G4087_0[1]),.din(w_dff_A_ZtjjC1cr6_1),.clk(gclk));
	jdff dff_A_yQpYbEpp5_2(.dout(w_G4087_0[2]),.din(w_dff_A_yQpYbEpp5_2),.clk(gclk));
	jdff dff_A_stD9tdsP3_0(.dout(w_G4088_3[0]),.din(w_dff_A_stD9tdsP3_0),.clk(gclk));
	jdff dff_A_GzQHRemz8_0(.dout(w_dff_A_stD9tdsP3_0),.din(w_dff_A_GzQHRemz8_0),.clk(gclk));
	jdff dff_A_q2xxL2809_0(.dout(w_dff_A_GzQHRemz8_0),.din(w_dff_A_q2xxL2809_0),.clk(gclk));
	jdff dff_A_wjn5NGJL4_0(.dout(w_dff_A_q2xxL2809_0),.din(w_dff_A_wjn5NGJL4_0),.clk(gclk));
	jdff dff_A_3vHb5jwq0_0(.dout(w_dff_A_wjn5NGJL4_0),.din(w_dff_A_3vHb5jwq0_0),.clk(gclk));
	jdff dff_A_BxOZloTC5_0(.dout(w_dff_A_3vHb5jwq0_0),.din(w_dff_A_BxOZloTC5_0),.clk(gclk));
	jdff dff_A_d2LAGOai2_0(.dout(w_dff_A_BxOZloTC5_0),.din(w_dff_A_d2LAGOai2_0),.clk(gclk));
	jdff dff_A_gKJA16UU5_0(.dout(w_dff_A_d2LAGOai2_0),.din(w_dff_A_gKJA16UU5_0),.clk(gclk));
	jdff dff_A_4c45Rt3G2_0(.dout(w_dff_A_gKJA16UU5_0),.din(w_dff_A_4c45Rt3G2_0),.clk(gclk));
	jdff dff_A_7f1V6vuB5_0(.dout(w_dff_A_4c45Rt3G2_0),.din(w_dff_A_7f1V6vuB5_0),.clk(gclk));
	jdff dff_A_IdcioEF45_0(.dout(w_dff_A_7f1V6vuB5_0),.din(w_dff_A_IdcioEF45_0),.clk(gclk));
	jdff dff_A_NXCW0Peo0_0(.dout(w_dff_A_IdcioEF45_0),.din(w_dff_A_NXCW0Peo0_0),.clk(gclk));
	jdff dff_A_cKVgP91G6_0(.dout(w_dff_A_NXCW0Peo0_0),.din(w_dff_A_cKVgP91G6_0),.clk(gclk));
	jdff dff_A_Rr3erOfF6_0(.dout(w_dff_A_cKVgP91G6_0),.din(w_dff_A_Rr3erOfF6_0),.clk(gclk));
	jdff dff_A_I5pOKBT10_0(.dout(w_dff_A_Rr3erOfF6_0),.din(w_dff_A_I5pOKBT10_0),.clk(gclk));
	jdff dff_A_rKht7d1D0_0(.dout(w_dff_A_I5pOKBT10_0),.din(w_dff_A_rKht7d1D0_0),.clk(gclk));
	jdff dff_A_EOyZ921T3_0(.dout(w_dff_A_rKht7d1D0_0),.din(w_dff_A_EOyZ921T3_0),.clk(gclk));
	jdff dff_A_eP5pG42G3_0(.dout(w_dff_A_EOyZ921T3_0),.din(w_dff_A_eP5pG42G3_0),.clk(gclk));
	jdff dff_A_m5UgHlOP8_0(.dout(w_dff_A_eP5pG42G3_0),.din(w_dff_A_m5UgHlOP8_0),.clk(gclk));
	jdff dff_A_BIn5dbuA0_0(.dout(w_dff_A_m5UgHlOP8_0),.din(w_dff_A_BIn5dbuA0_0),.clk(gclk));
	jdff dff_A_ZrCBTGC77_0(.dout(w_dff_A_BIn5dbuA0_0),.din(w_dff_A_ZrCBTGC77_0),.clk(gclk));
	jdff dff_A_xo76DDLe0_0(.dout(w_dff_A_ZrCBTGC77_0),.din(w_dff_A_xo76DDLe0_0),.clk(gclk));
	jdff dff_A_e2DMmeF93_0(.dout(w_dff_A_xo76DDLe0_0),.din(w_dff_A_e2DMmeF93_0),.clk(gclk));
	jdff dff_B_5VWJlEk10_1(.din(n1688),.dout(w_dff_B_5VWJlEk10_1),.clk(gclk));
	jdff dff_B_FKUbdl895_1(.din(w_dff_B_5VWJlEk10_1),.dout(w_dff_B_FKUbdl895_1),.clk(gclk));
	jdff dff_B_GhtElLy78_1(.din(w_dff_B_FKUbdl895_1),.dout(w_dff_B_GhtElLy78_1),.clk(gclk));
	jdff dff_B_N1ppBTzP7_1(.din(w_dff_B_GhtElLy78_1),.dout(w_dff_B_N1ppBTzP7_1),.clk(gclk));
	jdff dff_B_qaJaVZEb7_1(.din(w_dff_B_N1ppBTzP7_1),.dout(w_dff_B_qaJaVZEb7_1),.clk(gclk));
	jdff dff_B_DPx4D44O9_1(.din(w_dff_B_qaJaVZEb7_1),.dout(w_dff_B_DPx4D44O9_1),.clk(gclk));
	jdff dff_B_MIPrLEAQ4_1(.din(w_dff_B_DPx4D44O9_1),.dout(w_dff_B_MIPrLEAQ4_1),.clk(gclk));
	jdff dff_B_2p7NKM7G4_1(.din(w_dff_B_MIPrLEAQ4_1),.dout(w_dff_B_2p7NKM7G4_1),.clk(gclk));
	jdff dff_B_W4eb44Fa9_1(.din(w_dff_B_2p7NKM7G4_1),.dout(w_dff_B_W4eb44Fa9_1),.clk(gclk));
	jdff dff_B_WueJfSvG9_1(.din(w_dff_B_W4eb44Fa9_1),.dout(w_dff_B_WueJfSvG9_1),.clk(gclk));
	jdff dff_B_i02qVWdV5_1(.din(w_dff_B_WueJfSvG9_1),.dout(w_dff_B_i02qVWdV5_1),.clk(gclk));
	jdff dff_B_tz9ImYf91_1(.din(w_dff_B_i02qVWdV5_1),.dout(w_dff_B_tz9ImYf91_1),.clk(gclk));
	jdff dff_B_kFRza5023_1(.din(w_dff_B_tz9ImYf91_1),.dout(w_dff_B_kFRza5023_1),.clk(gclk));
	jdff dff_B_Jw1xMxJU9_1(.din(w_dff_B_kFRza5023_1),.dout(w_dff_B_Jw1xMxJU9_1),.clk(gclk));
	jdff dff_B_rGCXZjog7_1(.din(w_dff_B_Jw1xMxJU9_1),.dout(w_dff_B_rGCXZjog7_1),.clk(gclk));
	jdff dff_B_A6VkFRSM6_1(.din(w_dff_B_rGCXZjog7_1),.dout(w_dff_B_A6VkFRSM6_1),.clk(gclk));
	jdff dff_B_7zLHV44n1_1(.din(w_dff_B_A6VkFRSM6_1),.dout(w_dff_B_7zLHV44n1_1),.clk(gclk));
	jdff dff_B_vVmKJpte0_1(.din(w_dff_B_7zLHV44n1_1),.dout(w_dff_B_vVmKJpte0_1),.clk(gclk));
	jdff dff_B_JxXsnwWw9_1(.din(w_dff_B_vVmKJpte0_1),.dout(w_dff_B_JxXsnwWw9_1),.clk(gclk));
	jdff dff_B_AvTLxa0U9_1(.din(w_dff_B_JxXsnwWw9_1),.dout(w_dff_B_AvTLxa0U9_1),.clk(gclk));
	jdff dff_B_0COEn1EF5_1(.din(w_dff_B_AvTLxa0U9_1),.dout(w_dff_B_0COEn1EF5_1),.clk(gclk));
	jdff dff_B_JZhC67786_1(.din(w_dff_B_0COEn1EF5_1),.dout(w_dff_B_JZhC67786_1),.clk(gclk));
	jdff dff_B_4w8ijg4L1_1(.din(n1689),.dout(w_dff_B_4w8ijg4L1_1),.clk(gclk));
	jdff dff_A_XHd2QwV55_1(.dout(w_n854_1[1]),.din(w_dff_A_XHd2QwV55_1),.clk(gclk));
	jdff dff_A_Ap4mMjKA8_1(.dout(w_dff_A_XHd2QwV55_1),.din(w_dff_A_Ap4mMjKA8_1),.clk(gclk));
	jdff dff_A_v0A9eA911_1(.dout(w_dff_A_Ap4mMjKA8_1),.din(w_dff_A_v0A9eA911_1),.clk(gclk));
	jdff dff_A_ysOOM7QB4_1(.dout(w_dff_A_v0A9eA911_1),.din(w_dff_A_ysOOM7QB4_1),.clk(gclk));
	jdff dff_A_Ka0TaOuV2_1(.dout(w_dff_A_ysOOM7QB4_1),.din(w_dff_A_Ka0TaOuV2_1),.clk(gclk));
	jdff dff_A_mmrxd1oL7_1(.dout(w_dff_A_Ka0TaOuV2_1),.din(w_dff_A_mmrxd1oL7_1),.clk(gclk));
	jdff dff_A_6bNMblGB6_1(.dout(w_dff_A_mmrxd1oL7_1),.din(w_dff_A_6bNMblGB6_1),.clk(gclk));
	jdff dff_A_xji6pgNy8_1(.dout(w_dff_A_6bNMblGB6_1),.din(w_dff_A_xji6pgNy8_1),.clk(gclk));
	jdff dff_A_ToTuOMhx6_1(.dout(w_dff_A_xji6pgNy8_1),.din(w_dff_A_ToTuOMhx6_1),.clk(gclk));
	jdff dff_A_6ZjksA0e1_1(.dout(w_dff_A_ToTuOMhx6_1),.din(w_dff_A_6ZjksA0e1_1),.clk(gclk));
	jdff dff_A_bPTvEwAl5_1(.dout(w_dff_A_6ZjksA0e1_1),.din(w_dff_A_bPTvEwAl5_1),.clk(gclk));
	jdff dff_A_tUZ1kFg80_1(.dout(w_dff_A_bPTvEwAl5_1),.din(w_dff_A_tUZ1kFg80_1),.clk(gclk));
	jdff dff_A_AzxWRYBH5_1(.dout(w_dff_A_tUZ1kFg80_1),.din(w_dff_A_AzxWRYBH5_1),.clk(gclk));
	jdff dff_A_MADeFKk91_1(.dout(w_dff_A_AzxWRYBH5_1),.din(w_dff_A_MADeFKk91_1),.clk(gclk));
	jdff dff_A_HSeYYdKz2_2(.dout(w_n854_1[2]),.din(w_dff_A_HSeYYdKz2_2),.clk(gclk));
	jdff dff_A_vIcfKhgF2_2(.dout(w_dff_A_HSeYYdKz2_2),.din(w_dff_A_vIcfKhgF2_2),.clk(gclk));
	jdff dff_A_lQAzILS92_2(.dout(w_dff_A_vIcfKhgF2_2),.din(w_dff_A_lQAzILS92_2),.clk(gclk));
	jdff dff_A_vcWsDHm01_2(.dout(w_dff_A_lQAzILS92_2),.din(w_dff_A_vcWsDHm01_2),.clk(gclk));
	jdff dff_A_N3rKhFR06_2(.dout(w_dff_A_vcWsDHm01_2),.din(w_dff_A_N3rKhFR06_2),.clk(gclk));
	jdff dff_A_kkjVur1N4_2(.dout(w_dff_A_N3rKhFR06_2),.din(w_dff_A_kkjVur1N4_2),.clk(gclk));
	jdff dff_A_vpbSd4Xr2_2(.dout(w_dff_A_kkjVur1N4_2),.din(w_dff_A_vpbSd4Xr2_2),.clk(gclk));
	jdff dff_A_UbJhJIwu0_2(.dout(w_dff_A_vpbSd4Xr2_2),.din(w_dff_A_UbJhJIwu0_2),.clk(gclk));
	jdff dff_A_5Lr90UL94_2(.dout(w_dff_A_UbJhJIwu0_2),.din(w_dff_A_5Lr90UL94_2),.clk(gclk));
	jdff dff_A_cFnCmMlb6_2(.dout(w_dff_A_5Lr90UL94_2),.din(w_dff_A_cFnCmMlb6_2),.clk(gclk));
	jdff dff_A_duCczTxM6_1(.dout(w_n854_0[1]),.din(w_dff_A_duCczTxM6_1),.clk(gclk));
	jdff dff_A_vsdwndrL6_1(.dout(w_dff_A_duCczTxM6_1),.din(w_dff_A_vsdwndrL6_1),.clk(gclk));
	jdff dff_A_DnrT2OXK6_1(.dout(w_dff_A_vsdwndrL6_1),.din(w_dff_A_DnrT2OXK6_1),.clk(gclk));
	jdff dff_A_oUqq3q7g6_1(.dout(w_dff_A_DnrT2OXK6_1),.din(w_dff_A_oUqq3q7g6_1),.clk(gclk));
	jdff dff_A_BPJPEmzi0_1(.dout(w_dff_A_oUqq3q7g6_1),.din(w_dff_A_BPJPEmzi0_1),.clk(gclk));
	jdff dff_A_Ej2ttc3v6_1(.dout(w_dff_A_BPJPEmzi0_1),.din(w_dff_A_Ej2ttc3v6_1),.clk(gclk));
	jdff dff_A_o4OMuCUz2_1(.dout(w_dff_A_Ej2ttc3v6_1),.din(w_dff_A_o4OMuCUz2_1),.clk(gclk));
	jdff dff_A_YB9OgIea1_1(.dout(w_dff_A_o4OMuCUz2_1),.din(w_dff_A_YB9OgIea1_1),.clk(gclk));
	jdff dff_A_3VItfUrT1_1(.dout(w_dff_A_YB9OgIea1_1),.din(w_dff_A_3VItfUrT1_1),.clk(gclk));
	jdff dff_A_A304rUl82_1(.dout(w_dff_A_3VItfUrT1_1),.din(w_dff_A_A304rUl82_1),.clk(gclk));
	jdff dff_A_DhjotKiY6_1(.dout(w_dff_A_A304rUl82_1),.din(w_dff_A_DhjotKiY6_1),.clk(gclk));
	jdff dff_A_BhU2XX7h7_2(.dout(w_n854_0[2]),.din(w_dff_A_BhU2XX7h7_2),.clk(gclk));
	jdff dff_A_2niEqCLp7_2(.dout(w_dff_A_BhU2XX7h7_2),.din(w_dff_A_2niEqCLp7_2),.clk(gclk));
	jdff dff_A_YhQiCBCf8_2(.dout(w_dff_A_2niEqCLp7_2),.din(w_dff_A_YhQiCBCf8_2),.clk(gclk));
	jdff dff_A_8CdQoD6j4_2(.dout(w_dff_A_YhQiCBCf8_2),.din(w_dff_A_8CdQoD6j4_2),.clk(gclk));
	jdff dff_A_GJS3iESA2_2(.dout(w_dff_A_8CdQoD6j4_2),.din(w_dff_A_GJS3iESA2_2),.clk(gclk));
	jdff dff_B_YU5aFbwY8_3(.din(n854),.dout(w_dff_B_YU5aFbwY8_3),.clk(gclk));
	jdff dff_B_mASZFfYi0_3(.din(w_dff_B_YU5aFbwY8_3),.dout(w_dff_B_mASZFfYi0_3),.clk(gclk));
	jdff dff_B_X7VLNaWq3_3(.din(w_dff_B_mASZFfYi0_3),.dout(w_dff_B_X7VLNaWq3_3),.clk(gclk));
	jdff dff_B_QCV7Orfh1_3(.din(w_dff_B_X7VLNaWq3_3),.dout(w_dff_B_QCV7Orfh1_3),.clk(gclk));
	jdff dff_B_v84117wn9_3(.din(w_dff_B_QCV7Orfh1_3),.dout(w_dff_B_v84117wn9_3),.clk(gclk));
	jdff dff_B_KIsqCmnf9_3(.din(w_dff_B_v84117wn9_3),.dout(w_dff_B_KIsqCmnf9_3),.clk(gclk));
	jdff dff_B_YNEIxzyE8_3(.din(w_dff_B_KIsqCmnf9_3),.dout(w_dff_B_YNEIxzyE8_3),.clk(gclk));
	jdff dff_B_QnYnZjV90_3(.din(w_dff_B_YNEIxzyE8_3),.dout(w_dff_B_QnYnZjV90_3),.clk(gclk));
	jdff dff_B_LKKyFNdM0_3(.din(w_dff_B_QnYnZjV90_3),.dout(w_dff_B_LKKyFNdM0_3),.clk(gclk));
	jdff dff_A_rTzxTR3f9_0(.dout(w_G4090_4[0]),.din(w_dff_A_rTzxTR3f9_0),.clk(gclk));
	jdff dff_A_ghHCOaPZ1_0(.dout(w_dff_A_rTzxTR3f9_0),.din(w_dff_A_ghHCOaPZ1_0),.clk(gclk));
	jdff dff_A_y0stXhZv5_1(.dout(w_G4090_4[1]),.din(w_dff_A_y0stXhZv5_1),.clk(gclk));
	jdff dff_B_6890W6Pk6_1(.din(n1685),.dout(w_dff_B_6890W6Pk6_1),.clk(gclk));
	jdff dff_B_zD5UW9OE9_1(.din(w_dff_B_6890W6Pk6_1),.dout(w_dff_B_zD5UW9OE9_1),.clk(gclk));
	jdff dff_A_Md6L4ZLk1_0(.dout(w_n852_3[0]),.din(w_dff_A_Md6L4ZLk1_0),.clk(gclk));
	jdff dff_A_L1rL8Lnv3_0(.dout(w_dff_A_Md6L4ZLk1_0),.din(w_dff_A_L1rL8Lnv3_0),.clk(gclk));
	jdff dff_A_qRNKc1yt7_0(.dout(w_dff_A_L1rL8Lnv3_0),.din(w_dff_A_qRNKc1yt7_0),.clk(gclk));
	jdff dff_A_ePbmOZq23_0(.dout(w_dff_A_qRNKc1yt7_0),.din(w_dff_A_ePbmOZq23_0),.clk(gclk));
	jdff dff_A_h4WNevPM8_0(.dout(w_dff_A_ePbmOZq23_0),.din(w_dff_A_h4WNevPM8_0),.clk(gclk));
	jdff dff_A_4BdJor4m2_0(.dout(w_dff_A_h4WNevPM8_0),.din(w_dff_A_4BdJor4m2_0),.clk(gclk));
	jdff dff_A_AiDyksuY8_0(.dout(w_dff_A_4BdJor4m2_0),.din(w_dff_A_AiDyksuY8_0),.clk(gclk));
	jdff dff_A_LiFeRp1E3_0(.dout(w_dff_A_AiDyksuY8_0),.din(w_dff_A_LiFeRp1E3_0),.clk(gclk));
	jdff dff_A_MccVLTGR2_0(.dout(w_dff_A_LiFeRp1E3_0),.din(w_dff_A_MccVLTGR2_0),.clk(gclk));
	jdff dff_A_FOVAUchP1_0(.dout(w_dff_A_MccVLTGR2_0),.din(w_dff_A_FOVAUchP1_0),.clk(gclk));
	jdff dff_A_AMohUKfL5_0(.dout(w_dff_A_FOVAUchP1_0),.din(w_dff_A_AMohUKfL5_0),.clk(gclk));
	jdff dff_A_xy8G4voT8_0(.dout(w_dff_A_AMohUKfL5_0),.din(w_dff_A_xy8G4voT8_0),.clk(gclk));
	jdff dff_A_EOr0CDKt2_0(.dout(w_dff_A_xy8G4voT8_0),.din(w_dff_A_EOr0CDKt2_0),.clk(gclk));
	jdff dff_A_cDeiVApS6_0(.dout(w_dff_A_EOr0CDKt2_0),.din(w_dff_A_cDeiVApS6_0),.clk(gclk));
	jdff dff_A_7OK8rxKQ2_0(.dout(w_dff_A_cDeiVApS6_0),.din(w_dff_A_7OK8rxKQ2_0),.clk(gclk));
	jdff dff_A_8K67Gti73_0(.dout(w_dff_A_7OK8rxKQ2_0),.din(w_dff_A_8K67Gti73_0),.clk(gclk));
	jdff dff_A_w9dg7Net7_0(.dout(w_dff_A_8K67Gti73_0),.din(w_dff_A_w9dg7Net7_0),.clk(gclk));
	jdff dff_A_TEtlqzdT3_0(.dout(w_dff_A_w9dg7Net7_0),.din(w_dff_A_TEtlqzdT3_0),.clk(gclk));
	jdff dff_A_8HZgfnTa5_0(.dout(w_dff_A_TEtlqzdT3_0),.din(w_dff_A_8HZgfnTa5_0),.clk(gclk));
	jdff dff_A_mwdF4tvc7_0(.dout(w_dff_A_8HZgfnTa5_0),.din(w_dff_A_mwdF4tvc7_0),.clk(gclk));
	jdff dff_A_hthhEKpR5_0(.dout(w_dff_A_mwdF4tvc7_0),.din(w_dff_A_hthhEKpR5_0),.clk(gclk));
	jdff dff_A_gPRdKgN45_0(.dout(w_dff_A_hthhEKpR5_0),.din(w_dff_A_gPRdKgN45_0),.clk(gclk));
	jdff dff_A_wt8bNgyy7_1(.dout(w_G4089_9[1]),.din(w_dff_A_wt8bNgyy7_1),.clk(gclk));
	jdff dff_A_A6De25d65_1(.dout(w_dff_A_wt8bNgyy7_1),.din(w_dff_A_A6De25d65_1),.clk(gclk));
	jdff dff_A_OdmbJE6u6_1(.dout(w_dff_A_A6De25d65_1),.din(w_dff_A_OdmbJE6u6_1),.clk(gclk));
	jdff dff_A_2W0nE7DX9_1(.dout(w_dff_A_OdmbJE6u6_1),.din(w_dff_A_2W0nE7DX9_1),.clk(gclk));
	jdff dff_A_HwNHOzNl1_1(.dout(w_dff_A_2W0nE7DX9_1),.din(w_dff_A_HwNHOzNl1_1),.clk(gclk));
	jdff dff_A_VBKp2dHu3_1(.dout(w_dff_A_HwNHOzNl1_1),.din(w_dff_A_VBKp2dHu3_1),.clk(gclk));
	jdff dff_A_txW4Kzme7_1(.dout(w_dff_A_VBKp2dHu3_1),.din(w_dff_A_txW4Kzme7_1),.clk(gclk));
	jdff dff_A_1xkcgrRy6_1(.dout(w_dff_A_txW4Kzme7_1),.din(w_dff_A_1xkcgrRy6_1),.clk(gclk));
	jdff dff_A_y6gLe14R0_1(.dout(w_dff_A_1xkcgrRy6_1),.din(w_dff_A_y6gLe14R0_1),.clk(gclk));
	jdff dff_B_YuQ5o83W9_2(.din(G64),.dout(w_dff_B_YuQ5o83W9_2),.clk(gclk));
	jdff dff_A_rrKM09fd4_1(.dout(w_G4090_1[1]),.din(w_dff_A_rrKM09fd4_1),.clk(gclk));
	jdff dff_A_a1NFrYxL3_1(.dout(w_dff_A_rrKM09fd4_1),.din(w_dff_A_a1NFrYxL3_1),.clk(gclk));
	jdff dff_A_oHlGz0YR3_2(.dout(w_G4090_1[2]),.din(w_dff_A_oHlGz0YR3_2),.clk(gclk));
	jdff dff_A_98uwd9An2_1(.dout(w_G4090_0[1]),.din(w_dff_A_98uwd9An2_1),.clk(gclk));
	jdff dff_A_N5K4KyUj0_2(.dout(w_G4090_0[2]),.din(w_dff_A_N5K4KyUj0_2),.clk(gclk));
	jdff dff_A_rdeyPKAs0_0(.dout(w_G4089_3[0]),.din(w_dff_A_rdeyPKAs0_0),.clk(gclk));
	jdff dff_A_rJ4BELuO9_0(.dout(w_dff_A_rdeyPKAs0_0),.din(w_dff_A_rJ4BELuO9_0),.clk(gclk));
	jdff dff_A_QsjLx9Ce7_0(.dout(w_dff_A_rJ4BELuO9_0),.din(w_dff_A_QsjLx9Ce7_0),.clk(gclk));
	jdff dff_A_C9GsvAJa7_0(.dout(w_dff_A_QsjLx9Ce7_0),.din(w_dff_A_C9GsvAJa7_0),.clk(gclk));
	jdff dff_A_y1xvDWAF2_0(.dout(w_dff_A_C9GsvAJa7_0),.din(w_dff_A_y1xvDWAF2_0),.clk(gclk));
	jdff dff_A_tO0Qrx1f1_0(.dout(w_dff_A_y1xvDWAF2_0),.din(w_dff_A_tO0Qrx1f1_0),.clk(gclk));
	jdff dff_A_IEu0Uf5u3_0(.dout(w_dff_A_tO0Qrx1f1_0),.din(w_dff_A_IEu0Uf5u3_0),.clk(gclk));
	jdff dff_A_oBHPoYYs8_0(.dout(w_dff_A_IEu0Uf5u3_0),.din(w_dff_A_oBHPoYYs8_0),.clk(gclk));
	jdff dff_A_k35eJEDi1_0(.dout(w_dff_A_oBHPoYYs8_0),.din(w_dff_A_k35eJEDi1_0),.clk(gclk));
	jdff dff_A_MsesAbzI5_0(.dout(w_dff_A_k35eJEDi1_0),.din(w_dff_A_MsesAbzI5_0),.clk(gclk));
	jdff dff_A_TAEROzuT5_0(.dout(w_dff_A_MsesAbzI5_0),.din(w_dff_A_TAEROzuT5_0),.clk(gclk));
	jdff dff_A_ATy3qVdy1_0(.dout(w_dff_A_TAEROzuT5_0),.din(w_dff_A_ATy3qVdy1_0),.clk(gclk));
	jdff dff_A_oHE4udjl1_0(.dout(w_dff_A_ATy3qVdy1_0),.din(w_dff_A_oHE4udjl1_0),.clk(gclk));
	jdff dff_A_tAkLuTeL3_0(.dout(w_dff_A_oHE4udjl1_0),.din(w_dff_A_tAkLuTeL3_0),.clk(gclk));
	jdff dff_A_MFrG6Vnt9_0(.dout(w_dff_A_tAkLuTeL3_0),.din(w_dff_A_MFrG6Vnt9_0),.clk(gclk));
	jdff dff_A_j6HF3K6N8_0(.dout(w_dff_A_MFrG6Vnt9_0),.din(w_dff_A_j6HF3K6N8_0),.clk(gclk));
	jdff dff_A_bPPJTE1Z3_0(.dout(w_dff_A_j6HF3K6N8_0),.din(w_dff_A_bPPJTE1Z3_0),.clk(gclk));
	jdff dff_A_jyR1jeXn2_0(.dout(w_dff_A_bPPJTE1Z3_0),.din(w_dff_A_jyR1jeXn2_0),.clk(gclk));
	jdff dff_A_rfIPd6nx3_0(.dout(w_dff_A_jyR1jeXn2_0),.din(w_dff_A_rfIPd6nx3_0),.clk(gclk));
	jdff dff_A_RSZ9pChh2_0(.dout(w_dff_A_rfIPd6nx3_0),.din(w_dff_A_RSZ9pChh2_0),.clk(gclk));
	jdff dff_A_ie7Z40Gz9_0(.dout(w_dff_A_RSZ9pChh2_0),.din(w_dff_A_ie7Z40Gz9_0),.clk(gclk));
	jdff dff_A_ZPALRbNc1_0(.dout(w_dff_A_ie7Z40Gz9_0),.din(w_dff_A_ZPALRbNc1_0),.clk(gclk));
	jdff dff_A_M6dwhNZe0_0(.dout(w_dff_A_ZPALRbNc1_0),.din(w_dff_A_M6dwhNZe0_0),.clk(gclk));
	jdff dff_B_bMIbFn0F5_1(.din(n1697),.dout(w_dff_B_bMIbFn0F5_1),.clk(gclk));
	jdff dff_B_Oa9qd6IH4_1(.din(w_dff_B_bMIbFn0F5_1),.dout(w_dff_B_Oa9qd6IH4_1),.clk(gclk));
	jdff dff_B_wGu4CYYp9_1(.din(w_dff_B_Oa9qd6IH4_1),.dout(w_dff_B_wGu4CYYp9_1),.clk(gclk));
	jdff dff_B_Ue4dzxzn0_1(.din(w_dff_B_wGu4CYYp9_1),.dout(w_dff_B_Ue4dzxzn0_1),.clk(gclk));
	jdff dff_B_ELSlJ2Fh7_1(.din(w_dff_B_Ue4dzxzn0_1),.dout(w_dff_B_ELSlJ2Fh7_1),.clk(gclk));
	jdff dff_B_TnFwnLhE0_1(.din(w_dff_B_ELSlJ2Fh7_1),.dout(w_dff_B_TnFwnLhE0_1),.clk(gclk));
	jdff dff_B_0Mqoad4x4_1(.din(w_dff_B_TnFwnLhE0_1),.dout(w_dff_B_0Mqoad4x4_1),.clk(gclk));
	jdff dff_B_ltrxup4S5_1(.din(w_dff_B_0Mqoad4x4_1),.dout(w_dff_B_ltrxup4S5_1),.clk(gclk));
	jdff dff_B_5LAFverN7_1(.din(w_dff_B_ltrxup4S5_1),.dout(w_dff_B_5LAFverN7_1),.clk(gclk));
	jdff dff_B_JCr0poLX2_1(.din(w_dff_B_5LAFverN7_1),.dout(w_dff_B_JCr0poLX2_1),.clk(gclk));
	jdff dff_B_5G8zQwIv0_1(.din(w_dff_B_JCr0poLX2_1),.dout(w_dff_B_5G8zQwIv0_1),.clk(gclk));
	jdff dff_B_fP0jmasL8_1(.din(w_dff_B_5G8zQwIv0_1),.dout(w_dff_B_fP0jmasL8_1),.clk(gclk));
	jdff dff_B_AB3Z6gZY9_1(.din(w_dff_B_fP0jmasL8_1),.dout(w_dff_B_AB3Z6gZY9_1),.clk(gclk));
	jdff dff_B_N9p2ONu75_1(.din(w_dff_B_AB3Z6gZY9_1),.dout(w_dff_B_N9p2ONu75_1),.clk(gclk));
	jdff dff_B_6uQeOPUq7_1(.din(w_dff_B_N9p2ONu75_1),.dout(w_dff_B_6uQeOPUq7_1),.clk(gclk));
	jdff dff_B_uW0c6eat7_1(.din(w_dff_B_6uQeOPUq7_1),.dout(w_dff_B_uW0c6eat7_1),.clk(gclk));
	jdff dff_B_K7gGYNGh6_1(.din(w_dff_B_uW0c6eat7_1),.dout(w_dff_B_K7gGYNGh6_1),.clk(gclk));
	jdff dff_B_e9N9hQB34_1(.din(w_dff_B_K7gGYNGh6_1),.dout(w_dff_B_e9N9hQB34_1),.clk(gclk));
	jdff dff_B_yBPMgex56_1(.din(w_dff_B_e9N9hQB34_1),.dout(w_dff_B_yBPMgex56_1),.clk(gclk));
	jdff dff_B_EJ1vIkfj9_1(.din(w_dff_B_yBPMgex56_1),.dout(w_dff_B_EJ1vIkfj9_1),.clk(gclk));
	jdff dff_B_3Pnvo5Wy4_1(.din(w_dff_B_EJ1vIkfj9_1),.dout(w_dff_B_3Pnvo5Wy4_1),.clk(gclk));
	jdff dff_B_yxl5bIgC1_1(.din(w_dff_B_3Pnvo5Wy4_1),.dout(w_dff_B_yxl5bIgC1_1),.clk(gclk));
	jdff dff_B_OFoLb81D1_1(.din(w_dff_B_yxl5bIgC1_1),.dout(w_dff_B_OFoLb81D1_1),.clk(gclk));
	jdff dff_B_BtjNFnQ62_1(.din(n1700),.dout(w_dff_B_BtjNFnQ62_1),.clk(gclk));
	jdff dff_B_7zbOjT482_1(.din(w_dff_B_BtjNFnQ62_1),.dout(w_dff_B_7zbOjT482_1),.clk(gclk));
	jdff dff_B_X3Q2TPw86_1(.din(w_dff_B_7zbOjT482_1),.dout(w_dff_B_X3Q2TPw86_1),.clk(gclk));
	jdff dff_B_VBQ2ByaR2_1(.din(w_dff_B_X3Q2TPw86_1),.dout(w_dff_B_VBQ2ByaR2_1),.clk(gclk));
	jdff dff_B_HP4pVqIo7_1(.din(w_dff_B_VBQ2ByaR2_1),.dout(w_dff_B_HP4pVqIo7_1),.clk(gclk));
	jdff dff_B_szQD7lG23_1(.din(w_dff_B_HP4pVqIo7_1),.dout(w_dff_B_szQD7lG23_1),.clk(gclk));
	jdff dff_B_Wk9oLYPq2_1(.din(w_dff_B_szQD7lG23_1),.dout(w_dff_B_Wk9oLYPq2_1),.clk(gclk));
	jdff dff_B_J4crlOi21_1(.din(w_dff_B_Wk9oLYPq2_1),.dout(w_dff_B_J4crlOi21_1),.clk(gclk));
	jdff dff_B_d289MB6R7_1(.din(w_dff_B_J4crlOi21_1),.dout(w_dff_B_d289MB6R7_1),.clk(gclk));
	jdff dff_B_9qFjxQSI4_1(.din(w_dff_B_d289MB6R7_1),.dout(w_dff_B_9qFjxQSI4_1),.clk(gclk));
	jdff dff_B_lFXW8lHy0_1(.din(w_dff_B_9qFjxQSI4_1),.dout(w_dff_B_lFXW8lHy0_1),.clk(gclk));
	jdff dff_B_3aozawya1_1(.din(w_dff_B_lFXW8lHy0_1),.dout(w_dff_B_3aozawya1_1),.clk(gclk));
	jdff dff_B_35hDRlGt3_1(.din(w_dff_B_3aozawya1_1),.dout(w_dff_B_35hDRlGt3_1),.clk(gclk));
	jdff dff_B_g8DzMmqT5_1(.din(w_dff_B_35hDRlGt3_1),.dout(w_dff_B_g8DzMmqT5_1),.clk(gclk));
	jdff dff_B_1V2d6Ptw3_1(.din(w_dff_B_g8DzMmqT5_1),.dout(w_dff_B_1V2d6Ptw3_1),.clk(gclk));
	jdff dff_B_VaCCbFQW1_1(.din(w_dff_B_1V2d6Ptw3_1),.dout(w_dff_B_VaCCbFQW1_1),.clk(gclk));
	jdff dff_B_3lYlaJqe7_1(.din(w_dff_B_VaCCbFQW1_1),.dout(w_dff_B_3lYlaJqe7_1),.clk(gclk));
	jdff dff_B_vErUsyA04_1(.din(w_dff_B_3lYlaJqe7_1),.dout(w_dff_B_vErUsyA04_1),.clk(gclk));
	jdff dff_B_v4T5gsVC4_1(.din(w_dff_B_vErUsyA04_1),.dout(w_dff_B_v4T5gsVC4_1),.clk(gclk));
	jdff dff_B_0kJnOtNr6_1(.din(w_dff_B_v4T5gsVC4_1),.dout(w_dff_B_0kJnOtNr6_1),.clk(gclk));
	jdff dff_B_2cHRsFbU8_1(.din(w_dff_B_0kJnOtNr6_1),.dout(w_dff_B_2cHRsFbU8_1),.clk(gclk));
	jdff dff_B_yScOK9ru2_1(.din(n1701),.dout(w_dff_B_yScOK9ru2_1),.clk(gclk));
	jdff dff_A_SlYv8LDR1_0(.dout(w_n993_4[0]),.din(w_dff_A_SlYv8LDR1_0),.clk(gclk));
	jdff dff_A_ItebSVhY6_0(.dout(w_dff_A_SlYv8LDR1_0),.din(w_dff_A_ItebSVhY6_0),.clk(gclk));
	jdff dff_A_MdmZpCRp5_0(.dout(w_dff_A_ItebSVhY6_0),.din(w_dff_A_MdmZpCRp5_0),.clk(gclk));
	jdff dff_A_F3uKWVcV2_0(.dout(w_dff_A_MdmZpCRp5_0),.din(w_dff_A_F3uKWVcV2_0),.clk(gclk));
	jdff dff_A_qhnKv03l0_0(.dout(w_dff_A_F3uKWVcV2_0),.din(w_dff_A_qhnKv03l0_0),.clk(gclk));
	jdff dff_A_jyFXtZNu1_0(.dout(w_dff_A_qhnKv03l0_0),.din(w_dff_A_jyFXtZNu1_0),.clk(gclk));
	jdff dff_A_a3kbefkD9_0(.dout(w_dff_A_jyFXtZNu1_0),.din(w_dff_A_a3kbefkD9_0),.clk(gclk));
	jdff dff_A_wDfwGPd80_0(.dout(w_dff_A_a3kbefkD9_0),.din(w_dff_A_wDfwGPd80_0),.clk(gclk));
	jdff dff_A_jqIEugti6_0(.dout(w_dff_A_wDfwGPd80_0),.din(w_dff_A_jqIEugti6_0),.clk(gclk));
	jdff dff_A_Ioz0d5Nt4_0(.dout(w_dff_A_jqIEugti6_0),.din(w_dff_A_Ioz0d5Nt4_0),.clk(gclk));
	jdff dff_A_wYl1bAxT8_0(.dout(w_dff_A_Ioz0d5Nt4_0),.din(w_dff_A_wYl1bAxT8_0),.clk(gclk));
	jdff dff_A_yo3MvZQ20_0(.dout(w_dff_A_wYl1bAxT8_0),.din(w_dff_A_yo3MvZQ20_0),.clk(gclk));
	jdff dff_A_CA7cmmFD8_0(.dout(w_dff_A_yo3MvZQ20_0),.din(w_dff_A_CA7cmmFD8_0),.clk(gclk));
	jdff dff_A_jAKgpXcQ3_0(.dout(w_dff_A_CA7cmmFD8_0),.din(w_dff_A_jAKgpXcQ3_0),.clk(gclk));
	jdff dff_A_GY8z1wY53_0(.dout(w_dff_A_jAKgpXcQ3_0),.din(w_dff_A_GY8z1wY53_0),.clk(gclk));
	jdff dff_A_hBs0JYMO5_1(.dout(w_n993_4[1]),.din(w_dff_A_hBs0JYMO5_1),.clk(gclk));
	jdff dff_A_E00msF9S8_1(.dout(w_dff_A_hBs0JYMO5_1),.din(w_dff_A_E00msF9S8_1),.clk(gclk));
	jdff dff_A_KBrCNoyH2_1(.dout(w_dff_A_E00msF9S8_1),.din(w_dff_A_KBrCNoyH2_1),.clk(gclk));
	jdff dff_A_hQt0O5c47_1(.dout(w_dff_A_KBrCNoyH2_1),.din(w_dff_A_hQt0O5c47_1),.clk(gclk));
	jdff dff_A_s4HPvbzB5_1(.dout(w_dff_A_hQt0O5c47_1),.din(w_dff_A_s4HPvbzB5_1),.clk(gclk));
	jdff dff_A_9XR28cZQ0_1(.dout(w_dff_A_s4HPvbzB5_1),.din(w_dff_A_9XR28cZQ0_1),.clk(gclk));
	jdff dff_A_SaluuUvc8_1(.dout(w_dff_A_9XR28cZQ0_1),.din(w_dff_A_SaluuUvc8_1),.clk(gclk));
	jdff dff_A_IBgY35Ba8_1(.dout(w_dff_A_SaluuUvc8_1),.din(w_dff_A_IBgY35Ba8_1),.clk(gclk));
	jdff dff_A_LcIc8VQ40_1(.dout(w_dff_A_IBgY35Ba8_1),.din(w_dff_A_LcIc8VQ40_1),.clk(gclk));
	jdff dff_A_0fxBTHVS6_1(.dout(w_dff_A_LcIc8VQ40_1),.din(w_dff_A_0fxBTHVS6_1),.clk(gclk));
	jdff dff_A_Sx4BI8977_1(.dout(w_n993_1[1]),.din(w_dff_A_Sx4BI8977_1),.clk(gclk));
	jdff dff_A_BgW4wWCA1_1(.dout(w_dff_A_Sx4BI8977_1),.din(w_dff_A_BgW4wWCA1_1),.clk(gclk));
	jdff dff_A_zbtyXcT68_1(.dout(w_dff_A_BgW4wWCA1_1),.din(w_dff_A_zbtyXcT68_1),.clk(gclk));
	jdff dff_A_RXC5pQLZ0_1(.dout(w_dff_A_zbtyXcT68_1),.din(w_dff_A_RXC5pQLZ0_1),.clk(gclk));
	jdff dff_A_6q7gu6kZ5_1(.dout(w_dff_A_RXC5pQLZ0_1),.din(w_dff_A_6q7gu6kZ5_1),.clk(gclk));
	jdff dff_A_PvgqQlK40_1(.dout(w_dff_A_6q7gu6kZ5_1),.din(w_dff_A_PvgqQlK40_1),.clk(gclk));
	jdff dff_A_krANA6Z87_1(.dout(w_dff_A_PvgqQlK40_1),.din(w_dff_A_krANA6Z87_1),.clk(gclk));
	jdff dff_A_1naFaLhF2_1(.dout(w_dff_A_krANA6Z87_1),.din(w_dff_A_1naFaLhF2_1),.clk(gclk));
	jdff dff_A_Ojn0kkYc3_1(.dout(w_dff_A_1naFaLhF2_1),.din(w_dff_A_Ojn0kkYc3_1),.clk(gclk));
	jdff dff_A_LJnRnScN6_1(.dout(w_dff_A_Ojn0kkYc3_1),.din(w_dff_A_LJnRnScN6_1),.clk(gclk));
	jdff dff_A_oMXIdcBD7_1(.dout(w_dff_A_LJnRnScN6_1),.din(w_dff_A_oMXIdcBD7_1),.clk(gclk));
	jdff dff_A_DRrznnA01_1(.dout(w_dff_A_oMXIdcBD7_1),.din(w_dff_A_DRrznnA01_1),.clk(gclk));
	jdff dff_A_X0KzkqqW8_1(.dout(w_dff_A_DRrznnA01_1),.din(w_dff_A_X0KzkqqW8_1),.clk(gclk));
	jdff dff_A_q488RTdU3_1(.dout(w_dff_A_X0KzkqqW8_1),.din(w_dff_A_q488RTdU3_1),.clk(gclk));
	jdff dff_A_pC6vtcTT4_1(.dout(w_dff_A_q488RTdU3_1),.din(w_dff_A_pC6vtcTT4_1),.clk(gclk));
	jdff dff_A_oErH0m2e9_1(.dout(w_dff_A_pC6vtcTT4_1),.din(w_dff_A_oErH0m2e9_1),.clk(gclk));
	jdff dff_A_SmdYjCkC2_1(.dout(w_dff_A_oErH0m2e9_1),.din(w_dff_A_SmdYjCkC2_1),.clk(gclk));
	jdff dff_A_wv8LgdWo5_1(.dout(w_dff_A_SmdYjCkC2_1),.din(w_dff_A_wv8LgdWo5_1),.clk(gclk));
	jdff dff_A_vfOOW9eV1_1(.dout(w_dff_A_wv8LgdWo5_1),.din(w_dff_A_vfOOW9eV1_1),.clk(gclk));
	jdff dff_A_OmbFbeiy7_1(.dout(w_dff_A_vfOOW9eV1_1),.din(w_dff_A_OmbFbeiy7_1),.clk(gclk));
	jdff dff_A_LPoxAlm50_1(.dout(w_dff_A_OmbFbeiy7_1),.din(w_dff_A_LPoxAlm50_1),.clk(gclk));
	jdff dff_A_1apXy0ad4_2(.dout(w_n993_1[2]),.din(w_dff_A_1apXy0ad4_2),.clk(gclk));
	jdff dff_A_SjCjHrU97_2(.dout(w_dff_A_1apXy0ad4_2),.din(w_dff_A_SjCjHrU97_2),.clk(gclk));
	jdff dff_A_y2R6h7587_2(.dout(w_dff_A_SjCjHrU97_2),.din(w_dff_A_y2R6h7587_2),.clk(gclk));
	jdff dff_A_Ra9P4r6X0_2(.dout(w_dff_A_y2R6h7587_2),.din(w_dff_A_Ra9P4r6X0_2),.clk(gclk));
	jdff dff_A_XXSDnZKZ6_2(.dout(w_dff_A_Ra9P4r6X0_2),.din(w_dff_A_XXSDnZKZ6_2),.clk(gclk));
	jdff dff_A_7tYfKjwv0_2(.dout(w_dff_A_XXSDnZKZ6_2),.din(w_dff_A_7tYfKjwv0_2),.clk(gclk));
	jdff dff_A_fwTHRFFT7_2(.dout(w_dff_A_7tYfKjwv0_2),.din(w_dff_A_fwTHRFFT7_2),.clk(gclk));
	jdff dff_A_kes8BGOy5_2(.dout(w_dff_A_fwTHRFFT7_2),.din(w_dff_A_kes8BGOy5_2),.clk(gclk));
	jdff dff_A_cIKV6sB89_2(.dout(w_dff_A_kes8BGOy5_2),.din(w_dff_A_cIKV6sB89_2),.clk(gclk));
	jdff dff_A_tBOTIIWJ7_2(.dout(w_dff_A_cIKV6sB89_2),.din(w_dff_A_tBOTIIWJ7_2),.clk(gclk));
	jdff dff_A_uO7t2O6z3_2(.dout(w_dff_A_tBOTIIWJ7_2),.din(w_dff_A_uO7t2O6z3_2),.clk(gclk));
	jdff dff_A_f4Zs8oBC4_2(.dout(w_dff_A_uO7t2O6z3_2),.din(w_dff_A_f4Zs8oBC4_2),.clk(gclk));
	jdff dff_A_Whe0g9Av0_2(.dout(w_dff_A_f4Zs8oBC4_2),.din(w_dff_A_Whe0g9Av0_2),.clk(gclk));
	jdff dff_A_2B1qupzO7_2(.dout(w_dff_A_Whe0g9Av0_2),.din(w_dff_A_2B1qupzO7_2),.clk(gclk));
	jdff dff_A_jG06aDOL0_2(.dout(w_dff_A_2B1qupzO7_2),.din(w_dff_A_jG06aDOL0_2),.clk(gclk));
	jdff dff_A_NaB2w87d7_2(.dout(w_dff_A_jG06aDOL0_2),.din(w_dff_A_NaB2w87d7_2),.clk(gclk));
	jdff dff_A_Twvw7lxj4_2(.dout(w_dff_A_NaB2w87d7_2),.din(w_dff_A_Twvw7lxj4_2),.clk(gclk));
	jdff dff_A_oewqjaCp0_2(.dout(w_dff_A_Twvw7lxj4_2),.din(w_dff_A_oewqjaCp0_2),.clk(gclk));
	jdff dff_A_Lt74J5M05_2(.dout(w_dff_A_oewqjaCp0_2),.din(w_dff_A_Lt74J5M05_2),.clk(gclk));
	jdff dff_A_bFcptGNJ2_2(.dout(w_dff_A_Lt74J5M05_2),.din(w_dff_A_bFcptGNJ2_2),.clk(gclk));
	jdff dff_A_p4nLFl8q3_1(.dout(w_n993_0[1]),.din(w_dff_A_p4nLFl8q3_1),.clk(gclk));
	jdff dff_A_EYrLqPqr0_1(.dout(w_dff_A_p4nLFl8q3_1),.din(w_dff_A_EYrLqPqr0_1),.clk(gclk));
	jdff dff_A_mBvmh2bY5_1(.dout(w_dff_A_EYrLqPqr0_1),.din(w_dff_A_mBvmh2bY5_1),.clk(gclk));
	jdff dff_A_VRP4Ngk05_1(.dout(w_dff_A_mBvmh2bY5_1),.din(w_dff_A_VRP4Ngk05_1),.clk(gclk));
	jdff dff_A_X82o1FL83_1(.dout(w_dff_A_VRP4Ngk05_1),.din(w_dff_A_X82o1FL83_1),.clk(gclk));
	jdff dff_A_0lDIfkg95_1(.dout(w_dff_A_X82o1FL83_1),.din(w_dff_A_0lDIfkg95_1),.clk(gclk));
	jdff dff_A_IzmYZUuV3_1(.dout(w_dff_A_0lDIfkg95_1),.din(w_dff_A_IzmYZUuV3_1),.clk(gclk));
	jdff dff_A_VGJA1fJn7_1(.dout(w_dff_A_IzmYZUuV3_1),.din(w_dff_A_VGJA1fJn7_1),.clk(gclk));
	jdff dff_A_LMANtSHB6_1(.dout(w_dff_A_VGJA1fJn7_1),.din(w_dff_A_LMANtSHB6_1),.clk(gclk));
	jdff dff_A_ahxEezkt2_1(.dout(w_dff_A_LMANtSHB6_1),.din(w_dff_A_ahxEezkt2_1),.clk(gclk));
	jdff dff_A_x6JB4o569_1(.dout(w_dff_A_ahxEezkt2_1),.din(w_dff_A_x6JB4o569_1),.clk(gclk));
	jdff dff_A_2QQSaOSQ2_1(.dout(w_dff_A_x6JB4o569_1),.din(w_dff_A_2QQSaOSQ2_1),.clk(gclk));
	jdff dff_A_AZzYQT3o6_1(.dout(w_dff_A_2QQSaOSQ2_1),.din(w_dff_A_AZzYQT3o6_1),.clk(gclk));
	jdff dff_A_vp6kULU05_1(.dout(w_dff_A_AZzYQT3o6_1),.din(w_dff_A_vp6kULU05_1),.clk(gclk));
	jdff dff_A_MJtMi19x2_1(.dout(w_dff_A_vp6kULU05_1),.din(w_dff_A_MJtMi19x2_1),.clk(gclk));
	jdff dff_A_67K9j7t85_1(.dout(w_dff_A_MJtMi19x2_1),.din(w_dff_A_67K9j7t85_1),.clk(gclk));
	jdff dff_A_fFSRRVgn1_1(.dout(w_dff_A_67K9j7t85_1),.din(w_dff_A_fFSRRVgn1_1),.clk(gclk));
	jdff dff_A_KDQYG55A6_1(.dout(w_dff_A_fFSRRVgn1_1),.din(w_dff_A_KDQYG55A6_1),.clk(gclk));
	jdff dff_A_oLysiJcs3_2(.dout(w_n993_0[2]),.din(w_dff_A_oLysiJcs3_2),.clk(gclk));
	jdff dff_A_ggRoZm195_2(.dout(w_dff_A_oLysiJcs3_2),.din(w_dff_A_ggRoZm195_2),.clk(gclk));
	jdff dff_A_b0G6MoTR1_2(.dout(w_dff_A_ggRoZm195_2),.din(w_dff_A_b0G6MoTR1_2),.clk(gclk));
	jdff dff_A_HIL9ujgO0_2(.dout(w_dff_A_b0G6MoTR1_2),.din(w_dff_A_HIL9ujgO0_2),.clk(gclk));
	jdff dff_A_6SxZoqee7_2(.dout(w_dff_A_HIL9ujgO0_2),.din(w_dff_A_6SxZoqee7_2),.clk(gclk));
	jdff dff_A_NxmArqPE9_2(.dout(w_dff_A_6SxZoqee7_2),.din(w_dff_A_NxmArqPE9_2),.clk(gclk));
	jdff dff_A_FD6LLLM71_2(.dout(w_dff_A_NxmArqPE9_2),.din(w_dff_A_FD6LLLM71_2),.clk(gclk));
	jdff dff_A_K6hrhoON0_2(.dout(w_dff_A_FD6LLLM71_2),.din(w_dff_A_K6hrhoON0_2),.clk(gclk));
	jdff dff_A_1RU6fnuX6_2(.dout(w_dff_A_K6hrhoON0_2),.din(w_dff_A_1RU6fnuX6_2),.clk(gclk));
	jdff dff_A_zpurIaVN1_2(.dout(w_dff_A_1RU6fnuX6_2),.din(w_dff_A_zpurIaVN1_2),.clk(gclk));
	jdff dff_A_HLISzOAQ6_2(.dout(w_dff_A_zpurIaVN1_2),.din(w_dff_A_HLISzOAQ6_2),.clk(gclk));
	jdff dff_A_oQ6hWZ8K6_1(.dout(w_G1690_1[1]),.din(w_dff_A_oQ6hWZ8K6_1),.clk(gclk));
	jdff dff_A_ZqQ5dgBf9_1(.dout(w_G1690_0[1]),.din(w_dff_A_ZqQ5dgBf9_1),.clk(gclk));
	jdff dff_A_BCD8u8gK8_1(.dout(w_dff_A_ZqQ5dgBf9_1),.din(w_dff_A_BCD8u8gK8_1),.clk(gclk));
	jdff dff_A_g8SwvjE69_1(.dout(w_dff_A_BCD8u8gK8_1),.din(w_dff_A_g8SwvjE69_1),.clk(gclk));
	jdff dff_A_L21lRDsT2_1(.dout(w_dff_A_g8SwvjE69_1),.din(w_dff_A_L21lRDsT2_1),.clk(gclk));
	jdff dff_A_mjSB2XIM0_1(.dout(w_dff_A_L21lRDsT2_1),.din(w_dff_A_mjSB2XIM0_1),.clk(gclk));
	jdff dff_A_Z1j81ptQ7_1(.dout(w_dff_A_mjSB2XIM0_1),.din(w_dff_A_Z1j81ptQ7_1),.clk(gclk));
	jdff dff_A_2aaxuw399_1(.dout(w_dff_A_Z1j81ptQ7_1),.din(w_dff_A_2aaxuw399_1),.clk(gclk));
	jdff dff_A_jMxfTBlk9_1(.dout(w_dff_A_2aaxuw399_1),.din(w_dff_A_jMxfTBlk9_1),.clk(gclk));
	jdff dff_A_poynQU1Y6_1(.dout(w_dff_A_jMxfTBlk9_1),.din(w_dff_A_poynQU1Y6_1),.clk(gclk));
	jdff dff_A_v8Bg2hU68_1(.dout(w_dff_A_poynQU1Y6_1),.din(w_dff_A_v8Bg2hU68_1),.clk(gclk));
	jdff dff_A_4U0l04jV0_1(.dout(w_dff_A_v8Bg2hU68_1),.din(w_dff_A_4U0l04jV0_1),.clk(gclk));
	jdff dff_A_u4DWv6Lg0_1(.dout(w_dff_A_4U0l04jV0_1),.din(w_dff_A_u4DWv6Lg0_1),.clk(gclk));
	jdff dff_A_eIXvyG0r8_1(.dout(w_dff_A_u4DWv6Lg0_1),.din(w_dff_A_eIXvyG0r8_1),.clk(gclk));
	jdff dff_A_5RWirk279_1(.dout(w_dff_A_eIXvyG0r8_1),.din(w_dff_A_5RWirk279_1),.clk(gclk));
	jdff dff_A_yECbOnJk5_1(.dout(w_dff_A_5RWirk279_1),.din(w_dff_A_yECbOnJk5_1),.clk(gclk));
	jdff dff_A_c2vrPWTn6_1(.dout(w_dff_A_yECbOnJk5_1),.din(w_dff_A_c2vrPWTn6_1),.clk(gclk));
	jdff dff_A_odjQJDVI1_1(.dout(w_dff_A_c2vrPWTn6_1),.din(w_dff_A_odjQJDVI1_1),.clk(gclk));
	jdff dff_A_otNrD9H20_1(.dout(w_dff_A_odjQJDVI1_1),.din(w_dff_A_otNrD9H20_1),.clk(gclk));
	jdff dff_A_YA7kGA5z9_1(.dout(w_dff_A_otNrD9H20_1),.din(w_dff_A_YA7kGA5z9_1),.clk(gclk));
	jdff dff_A_AitZwGyh9_1(.dout(w_dff_A_YA7kGA5z9_1),.din(w_dff_A_AitZwGyh9_1),.clk(gclk));
	jdff dff_A_2UrOsUSd1_1(.dout(w_dff_A_AitZwGyh9_1),.din(w_dff_A_2UrOsUSd1_1),.clk(gclk));
	jdff dff_A_hgNgdS730_1(.dout(w_dff_A_2UrOsUSd1_1),.din(w_dff_A_hgNgdS730_1),.clk(gclk));
	jdff dff_A_8q1v2Fau8_1(.dout(w_dff_A_hgNgdS730_1),.din(w_dff_A_8q1v2Fau8_1),.clk(gclk));
	jdff dff_A_VwzzJvf65_0(.dout(w_G1689_1[0]),.din(w_dff_A_VwzzJvf65_0),.clk(gclk));
	jdff dff_A_ShNaac751_0(.dout(w_dff_A_VwzzJvf65_0),.din(w_dff_A_ShNaac751_0),.clk(gclk));
	jdff dff_A_5Oz4lCsW3_0(.dout(w_dff_A_ShNaac751_0),.din(w_dff_A_5Oz4lCsW3_0),.clk(gclk));
	jdff dff_A_ESwHyVEX2_0(.dout(w_dff_A_5Oz4lCsW3_0),.din(w_dff_A_ESwHyVEX2_0),.clk(gclk));
	jdff dff_A_ji7vJUdB3_0(.dout(w_dff_A_ESwHyVEX2_0),.din(w_dff_A_ji7vJUdB3_0),.clk(gclk));
	jdff dff_A_CS8RqFnI3_0(.dout(w_dff_A_ji7vJUdB3_0),.din(w_dff_A_CS8RqFnI3_0),.clk(gclk));
	jdff dff_A_pappRIuy5_0(.dout(w_dff_A_CS8RqFnI3_0),.din(w_dff_A_pappRIuy5_0),.clk(gclk));
	jdff dff_A_E009sSDJ5_0(.dout(w_dff_A_pappRIuy5_0),.din(w_dff_A_E009sSDJ5_0),.clk(gclk));
	jdff dff_A_DjEPVuot6_0(.dout(w_dff_A_E009sSDJ5_0),.din(w_dff_A_DjEPVuot6_0),.clk(gclk));
	jdff dff_A_63qojU8U2_2(.dout(w_G1689_1[2]),.din(w_dff_A_63qojU8U2_2),.clk(gclk));
	jdff dff_A_RfNOAa5D4_2(.dout(w_dff_A_63qojU8U2_2),.din(w_dff_A_RfNOAa5D4_2),.clk(gclk));
	jdff dff_A_iZPFkH8r6_2(.dout(w_dff_A_RfNOAa5D4_2),.din(w_dff_A_iZPFkH8r6_2),.clk(gclk));
	jdff dff_A_S0IfHSAp0_2(.dout(w_dff_A_iZPFkH8r6_2),.din(w_dff_A_S0IfHSAp0_2),.clk(gclk));
	jdff dff_A_Nq2xCbnW4_2(.dout(w_dff_A_S0IfHSAp0_2),.din(w_dff_A_Nq2xCbnW4_2),.clk(gclk));
	jdff dff_A_crbYARKb0_2(.dout(w_dff_A_Nq2xCbnW4_2),.din(w_dff_A_crbYARKb0_2),.clk(gclk));
	jdff dff_A_FgkZB9Mw4_2(.dout(w_dff_A_crbYARKb0_2),.din(w_dff_A_FgkZB9Mw4_2),.clk(gclk));
	jdff dff_A_vQ3mENBJ9_2(.dout(w_dff_A_FgkZB9Mw4_2),.din(w_dff_A_vQ3mENBJ9_2),.clk(gclk));
	jdff dff_A_s85UEDSu3_2(.dout(w_dff_A_vQ3mENBJ9_2),.din(w_dff_A_s85UEDSu3_2),.clk(gclk));
	jdff dff_A_ibqOQKJ08_2(.dout(w_dff_A_s85UEDSu3_2),.din(w_dff_A_ibqOQKJ08_2),.clk(gclk));
	jdff dff_A_5jt12NCG6_2(.dout(w_dff_A_ibqOQKJ08_2),.din(w_dff_A_5jt12NCG6_2),.clk(gclk));
	jdff dff_A_VOUGfFPN2_2(.dout(w_dff_A_5jt12NCG6_2),.din(w_dff_A_VOUGfFPN2_2),.clk(gclk));
	jdff dff_A_KbnJfHre1_2(.dout(w_dff_A_VOUGfFPN2_2),.din(w_dff_A_KbnJfHre1_2),.clk(gclk));
	jdff dff_A_kApJddP89_2(.dout(w_dff_A_KbnJfHre1_2),.din(w_dff_A_kApJddP89_2),.clk(gclk));
	jdff dff_A_LIRcmzzV4_2(.dout(w_dff_A_kApJddP89_2),.din(w_dff_A_LIRcmzzV4_2),.clk(gclk));
	jdff dff_A_DCfos2bf9_2(.dout(w_dff_A_LIRcmzzV4_2),.din(w_dff_A_DCfos2bf9_2),.clk(gclk));
	jdff dff_A_10iNWcyt9_2(.dout(w_dff_A_DCfos2bf9_2),.din(w_dff_A_10iNWcyt9_2),.clk(gclk));
	jdff dff_A_iWZg5kyo0_2(.dout(w_dff_A_10iNWcyt9_2),.din(w_dff_A_iWZg5kyo0_2),.clk(gclk));
	jdff dff_A_DKhhC6jr6_2(.dout(w_dff_A_iWZg5kyo0_2),.din(w_dff_A_DKhhC6jr6_2),.clk(gclk));
	jdff dff_A_8Bhrdh8W6_2(.dout(w_dff_A_DKhhC6jr6_2),.din(w_dff_A_8Bhrdh8W6_2),.clk(gclk));
	jdff dff_A_X8tib3Xx3_2(.dout(w_dff_A_8Bhrdh8W6_2),.din(w_dff_A_X8tib3Xx3_2),.clk(gclk));
	jdff dff_A_V9AeNPX94_2(.dout(w_dff_A_X8tib3Xx3_2),.din(w_dff_A_V9AeNPX94_2),.clk(gclk));
	jdff dff_A_773q4Ajn8_1(.dout(w_G1689_0[1]),.din(w_dff_A_773q4Ajn8_1),.clk(gclk));
	jdff dff_A_c8B6M1fH1_1(.dout(w_dff_A_773q4Ajn8_1),.din(w_dff_A_c8B6M1fH1_1),.clk(gclk));
	jdff dff_A_QlWRPz4U7_1(.dout(w_dff_A_c8B6M1fH1_1),.din(w_dff_A_QlWRPz4U7_1),.clk(gclk));
	jdff dff_A_nnpthrqL4_1(.dout(w_dff_A_QlWRPz4U7_1),.din(w_dff_A_nnpthrqL4_1),.clk(gclk));
	jdff dff_A_wPmKhg8A0_1(.dout(w_dff_A_nnpthrqL4_1),.din(w_dff_A_wPmKhg8A0_1),.clk(gclk));
	jdff dff_A_cwOmZkHW5_1(.dout(w_dff_A_wPmKhg8A0_1),.din(w_dff_A_cwOmZkHW5_1),.clk(gclk));
	jdff dff_A_M4Db9nyY5_1(.dout(w_dff_A_cwOmZkHW5_1),.din(w_dff_A_M4Db9nyY5_1),.clk(gclk));
	jdff dff_A_FJJYCpmb3_1(.dout(w_dff_A_M4Db9nyY5_1),.din(w_dff_A_FJJYCpmb3_1),.clk(gclk));
	jdff dff_A_C8UCi4yX7_1(.dout(w_dff_A_FJJYCpmb3_1),.din(w_dff_A_C8UCi4yX7_1),.clk(gclk));
	jdff dff_A_eH6uomXR6_1(.dout(w_dff_A_C8UCi4yX7_1),.din(w_dff_A_eH6uomXR6_1),.clk(gclk));
	jdff dff_A_zfQgTGRS8_1(.dout(w_dff_A_eH6uomXR6_1),.din(w_dff_A_zfQgTGRS8_1),.clk(gclk));
	jdff dff_A_GVWeV97E2_1(.dout(w_dff_A_zfQgTGRS8_1),.din(w_dff_A_GVWeV97E2_1),.clk(gclk));
	jdff dff_A_OUTm0v0B0_1(.dout(w_dff_A_GVWeV97E2_1),.din(w_dff_A_OUTm0v0B0_1),.clk(gclk));
	jdff dff_A_F960wYkX9_1(.dout(w_dff_A_OUTm0v0B0_1),.din(w_dff_A_F960wYkX9_1),.clk(gclk));
	jdff dff_A_JCCE42rm0_1(.dout(w_dff_A_F960wYkX9_1),.din(w_dff_A_JCCE42rm0_1),.clk(gclk));
	jdff dff_A_fxVNohek0_1(.dout(w_dff_A_JCCE42rm0_1),.din(w_dff_A_fxVNohek0_1),.clk(gclk));
	jdff dff_A_rrl7vplS7_1(.dout(w_dff_A_fxVNohek0_1),.din(w_dff_A_rrl7vplS7_1),.clk(gclk));
	jdff dff_A_gawc5Su77_1(.dout(w_dff_A_rrl7vplS7_1),.din(w_dff_A_gawc5Su77_1),.clk(gclk));
	jdff dff_A_TRFWSf9o9_1(.dout(w_dff_A_gawc5Su77_1),.din(w_dff_A_TRFWSf9o9_1),.clk(gclk));
	jdff dff_A_2UEpnK4m7_2(.dout(w_G1689_0[2]),.din(w_dff_A_2UEpnK4m7_2),.clk(gclk));
	jdff dff_A_acpypHIp4_2(.dout(w_dff_A_2UEpnK4m7_2),.din(w_dff_A_acpypHIp4_2),.clk(gclk));
	jdff dff_A_3ensXNEH3_2(.dout(w_dff_A_acpypHIp4_2),.din(w_dff_A_3ensXNEH3_2),.clk(gclk));
	jdff dff_A_9GgifZZj0_2(.dout(w_dff_A_3ensXNEH3_2),.din(w_dff_A_9GgifZZj0_2),.clk(gclk));
	jdff dff_A_SLN9LdOC7_2(.dout(w_dff_A_9GgifZZj0_2),.din(w_dff_A_SLN9LdOC7_2),.clk(gclk));
	jdff dff_A_EuADFi455_2(.dout(w_dff_A_SLN9LdOC7_2),.din(w_dff_A_EuADFi455_2),.clk(gclk));
	jdff dff_A_taIc74Ms2_2(.dout(w_dff_A_EuADFi455_2),.din(w_dff_A_taIc74Ms2_2),.clk(gclk));
	jdff dff_A_pYmkRsUp5_2(.dout(w_dff_A_taIc74Ms2_2),.din(w_dff_A_pYmkRsUp5_2),.clk(gclk));
	jdff dff_A_BJZnq2nh9_2(.dout(w_dff_A_pYmkRsUp5_2),.din(w_dff_A_BJZnq2nh9_2),.clk(gclk));
	jdff dff_A_GwsTqavO7_2(.dout(w_dff_A_BJZnq2nh9_2),.din(w_dff_A_GwsTqavO7_2),.clk(gclk));
	jdff dff_A_wl56k2at9_2(.dout(w_dff_A_GwsTqavO7_2),.din(w_dff_A_wl56k2at9_2),.clk(gclk));
	jdff dff_A_dqC8Jl5g8_2(.dout(w_dff_A_wl56k2at9_2),.din(w_dff_A_dqC8Jl5g8_2),.clk(gclk));
	jdff dff_A_qhYXJhut8_2(.dout(w_dff_A_dqC8Jl5g8_2),.din(w_dff_A_qhYXJhut8_2),.clk(gclk));
	jdff dff_B_fappLODQ3_1(.din(n1709),.dout(w_dff_B_fappLODQ3_1),.clk(gclk));
	jdff dff_B_K1eSItKk0_1(.din(w_dff_B_fappLODQ3_1),.dout(w_dff_B_K1eSItKk0_1),.clk(gclk));
	jdff dff_B_f4UNuX4U5_1(.din(w_dff_B_K1eSItKk0_1),.dout(w_dff_B_f4UNuX4U5_1),.clk(gclk));
	jdff dff_B_Xe6OwQUV0_1(.din(w_dff_B_f4UNuX4U5_1),.dout(w_dff_B_Xe6OwQUV0_1),.clk(gclk));
	jdff dff_B_vltlLjBs2_1(.din(w_dff_B_Xe6OwQUV0_1),.dout(w_dff_B_vltlLjBs2_1),.clk(gclk));
	jdff dff_B_ZNPbb3Je8_1(.din(w_dff_B_vltlLjBs2_1),.dout(w_dff_B_ZNPbb3Je8_1),.clk(gclk));
	jdff dff_B_LigNWl0D7_1(.din(w_dff_B_ZNPbb3Je8_1),.dout(w_dff_B_LigNWl0D7_1),.clk(gclk));
	jdff dff_B_JxbLPvAR2_1(.din(w_dff_B_LigNWl0D7_1),.dout(w_dff_B_JxbLPvAR2_1),.clk(gclk));
	jdff dff_B_N8ynxXMk0_1(.din(w_dff_B_JxbLPvAR2_1),.dout(w_dff_B_N8ynxXMk0_1),.clk(gclk));
	jdff dff_B_84PIClfp7_1(.din(w_dff_B_N8ynxXMk0_1),.dout(w_dff_B_84PIClfp7_1),.clk(gclk));
	jdff dff_B_G8uzX2zx0_1(.din(w_dff_B_84PIClfp7_1),.dout(w_dff_B_G8uzX2zx0_1),.clk(gclk));
	jdff dff_B_a1GkaZ6l0_1(.din(w_dff_B_G8uzX2zx0_1),.dout(w_dff_B_a1GkaZ6l0_1),.clk(gclk));
	jdff dff_B_jBZI8hw18_1(.din(w_dff_B_a1GkaZ6l0_1),.dout(w_dff_B_jBZI8hw18_1),.clk(gclk));
	jdff dff_B_PqLUO8oi4_1(.din(w_dff_B_jBZI8hw18_1),.dout(w_dff_B_PqLUO8oi4_1),.clk(gclk));
	jdff dff_B_3ubxHMpQ4_1(.din(w_dff_B_PqLUO8oi4_1),.dout(w_dff_B_3ubxHMpQ4_1),.clk(gclk));
	jdff dff_B_lkcI4hR56_1(.din(w_dff_B_3ubxHMpQ4_1),.dout(w_dff_B_lkcI4hR56_1),.clk(gclk));
	jdff dff_B_OYdWE7k76_1(.din(w_dff_B_lkcI4hR56_1),.dout(w_dff_B_OYdWE7k76_1),.clk(gclk));
	jdff dff_B_A84Spr3i9_1(.din(w_dff_B_OYdWE7k76_1),.dout(w_dff_B_A84Spr3i9_1),.clk(gclk));
	jdff dff_B_dG9LJPdV7_1(.din(w_dff_B_A84Spr3i9_1),.dout(w_dff_B_dG9LJPdV7_1),.clk(gclk));
	jdff dff_B_qKANdGMn4_1(.din(w_dff_B_dG9LJPdV7_1),.dout(w_dff_B_qKANdGMn4_1),.clk(gclk));
	jdff dff_B_x3SmIgxL6_1(.din(w_dff_B_qKANdGMn4_1),.dout(w_dff_B_x3SmIgxL6_1),.clk(gclk));
	jdff dff_B_Zp839Tqa8_1(.din(w_dff_B_x3SmIgxL6_1),.dout(w_dff_B_Zp839Tqa8_1),.clk(gclk));
	jdff dff_B_4pl9l5DJ3_1(.din(w_dff_B_Zp839Tqa8_1),.dout(w_dff_B_4pl9l5DJ3_1),.clk(gclk));
	jdff dff_B_7KxXvuiq5_1(.din(n1711),.dout(w_dff_B_7KxXvuiq5_1),.clk(gclk));
	jdff dff_B_VwMv84VU3_1(.din(w_dff_B_7KxXvuiq5_1),.dout(w_dff_B_VwMv84VU3_1),.clk(gclk));
	jdff dff_B_AztD1pwj1_1(.din(w_dff_B_VwMv84VU3_1),.dout(w_dff_B_AztD1pwj1_1),.clk(gclk));
	jdff dff_B_LyzQh7MP8_1(.din(w_dff_B_AztD1pwj1_1),.dout(w_dff_B_LyzQh7MP8_1),.clk(gclk));
	jdff dff_B_dJFA7P208_1(.din(w_dff_B_LyzQh7MP8_1),.dout(w_dff_B_dJFA7P208_1),.clk(gclk));
	jdff dff_B_Fq43BFwN3_1(.din(w_dff_B_dJFA7P208_1),.dout(w_dff_B_Fq43BFwN3_1),.clk(gclk));
	jdff dff_B_G0BVtXRn7_1(.din(w_dff_B_Fq43BFwN3_1),.dout(w_dff_B_G0BVtXRn7_1),.clk(gclk));
	jdff dff_B_kn63FJ2r7_1(.din(w_dff_B_G0BVtXRn7_1),.dout(w_dff_B_kn63FJ2r7_1),.clk(gclk));
	jdff dff_B_5Zutcn3n0_1(.din(w_dff_B_kn63FJ2r7_1),.dout(w_dff_B_5Zutcn3n0_1),.clk(gclk));
	jdff dff_B_TAinSHb54_1(.din(w_dff_B_5Zutcn3n0_1),.dout(w_dff_B_TAinSHb54_1),.clk(gclk));
	jdff dff_B_VLJu7GQG7_1(.din(w_dff_B_TAinSHb54_1),.dout(w_dff_B_VLJu7GQG7_1),.clk(gclk));
	jdff dff_B_GNgU3cM99_1(.din(w_dff_B_VLJu7GQG7_1),.dout(w_dff_B_GNgU3cM99_1),.clk(gclk));
	jdff dff_B_kIOcZ6FJ0_1(.din(w_dff_B_GNgU3cM99_1),.dout(w_dff_B_kIOcZ6FJ0_1),.clk(gclk));
	jdff dff_B_3mwH3La20_1(.din(w_dff_B_kIOcZ6FJ0_1),.dout(w_dff_B_3mwH3La20_1),.clk(gclk));
	jdff dff_B_pWpPGTZd5_1(.din(w_dff_B_3mwH3La20_1),.dout(w_dff_B_pWpPGTZd5_1),.clk(gclk));
	jdff dff_B_tT7GL0eE8_1(.din(w_dff_B_pWpPGTZd5_1),.dout(w_dff_B_tT7GL0eE8_1),.clk(gclk));
	jdff dff_B_vevqLO3x7_1(.din(w_dff_B_tT7GL0eE8_1),.dout(w_dff_B_vevqLO3x7_1),.clk(gclk));
	jdff dff_B_vQ9pZ3jq7_1(.din(w_dff_B_vevqLO3x7_1),.dout(w_dff_B_vQ9pZ3jq7_1),.clk(gclk));
	jdff dff_B_aOWQD9044_1(.din(w_dff_B_vQ9pZ3jq7_1),.dout(w_dff_B_aOWQD9044_1),.clk(gclk));
	jdff dff_B_r5AAnhzs6_1(.din(w_dff_B_aOWQD9044_1),.dout(w_dff_B_r5AAnhzs6_1),.clk(gclk));
	jdff dff_B_lPnA7KxI1_1(.din(w_dff_B_r5AAnhzs6_1),.dout(w_dff_B_lPnA7KxI1_1),.clk(gclk));
	jdff dff_B_TvwtaERu1_1(.din(n1712),.dout(w_dff_B_TvwtaERu1_1),.clk(gclk));
	jdff dff_B_uMayVPtM2_0(.din(n1678),.dout(w_dff_B_uMayVPtM2_0),.clk(gclk));
	jdff dff_B_YehyMLQ18_0(.din(w_dff_B_uMayVPtM2_0),.dout(w_dff_B_YehyMLQ18_0),.clk(gclk));
	jdff dff_B_oyrNO1rC6_0(.din(w_dff_B_YehyMLQ18_0),.dout(w_dff_B_oyrNO1rC6_0),.clk(gclk));
	jdff dff_B_Pzqkmj7s0_0(.din(w_dff_B_oyrNO1rC6_0),.dout(w_dff_B_Pzqkmj7s0_0),.clk(gclk));
	jdff dff_B_l9nXCu7R0_0(.din(w_dff_B_Pzqkmj7s0_0),.dout(w_dff_B_l9nXCu7R0_0),.clk(gclk));
	jdff dff_B_VuH0LG3Y0_0(.din(w_dff_B_l9nXCu7R0_0),.dout(w_dff_B_VuH0LG3Y0_0),.clk(gclk));
	jdff dff_B_7CLkLhNS4_0(.din(w_dff_B_VuH0LG3Y0_0),.dout(w_dff_B_7CLkLhNS4_0),.clk(gclk));
	jdff dff_B_dZfUUkFQ9_0(.din(w_dff_B_7CLkLhNS4_0),.dout(w_dff_B_dZfUUkFQ9_0),.clk(gclk));
	jdff dff_B_R0ph8LWv6_0(.din(w_dff_B_dZfUUkFQ9_0),.dout(w_dff_B_R0ph8LWv6_0),.clk(gclk));
	jdff dff_B_ihydbqsS0_0(.din(w_dff_B_R0ph8LWv6_0),.dout(w_dff_B_ihydbqsS0_0),.clk(gclk));
	jdff dff_B_1uf5h5F70_0(.din(w_dff_B_ihydbqsS0_0),.dout(w_dff_B_1uf5h5F70_0),.clk(gclk));
	jdff dff_B_d88tFYTL8_0(.din(w_dff_B_1uf5h5F70_0),.dout(w_dff_B_d88tFYTL8_0),.clk(gclk));
	jdff dff_B_t3YGfFxZ4_0(.din(w_dff_B_d88tFYTL8_0),.dout(w_dff_B_t3YGfFxZ4_0),.clk(gclk));
	jdff dff_B_KLvwqxyX5_0(.din(w_dff_B_t3YGfFxZ4_0),.dout(w_dff_B_KLvwqxyX5_0),.clk(gclk));
	jdff dff_B_seZyezCh5_0(.din(w_dff_B_KLvwqxyX5_0),.dout(w_dff_B_seZyezCh5_0),.clk(gclk));
	jdff dff_B_dJcJZI5n5_0(.din(w_dff_B_seZyezCh5_0),.dout(w_dff_B_dJcJZI5n5_0),.clk(gclk));
	jdff dff_B_wpWc3Yfc5_0(.din(w_dff_B_dJcJZI5n5_0),.dout(w_dff_B_wpWc3Yfc5_0),.clk(gclk));
	jdff dff_B_AR7NSALd2_0(.din(w_dff_B_wpWc3Yfc5_0),.dout(w_dff_B_AR7NSALd2_0),.clk(gclk));
	jdff dff_B_tshotWrx4_0(.din(w_dff_B_AR7NSALd2_0),.dout(w_dff_B_tshotWrx4_0),.clk(gclk));
	jdff dff_B_SX1hBGvL9_0(.din(n1501),.dout(w_dff_B_SX1hBGvL9_0),.clk(gclk));
	jdff dff_B_Vu0RJXKf9_0(.din(w_dff_B_SX1hBGvL9_0),.dout(w_dff_B_Vu0RJXKf9_0),.clk(gclk));
	jdff dff_B_n5BF50uh8_0(.din(w_dff_B_Vu0RJXKf9_0),.dout(w_dff_B_n5BF50uh8_0),.clk(gclk));
	jdff dff_B_Az16hyfc7_0(.din(w_dff_B_n5BF50uh8_0),.dout(w_dff_B_Az16hyfc7_0),.clk(gclk));
	jdff dff_B_HzbJxaAG6_0(.din(w_dff_B_Az16hyfc7_0),.dout(w_dff_B_HzbJxaAG6_0),.clk(gclk));
	jdff dff_B_wexuEVra7_0(.din(w_dff_B_HzbJxaAG6_0),.dout(w_dff_B_wexuEVra7_0),.clk(gclk));
	jdff dff_B_oCa9GmqI7_0(.din(w_dff_B_wexuEVra7_0),.dout(w_dff_B_oCa9GmqI7_0),.clk(gclk));
	jdff dff_B_Xefk6Yl04_0(.din(w_dff_B_oCa9GmqI7_0),.dout(w_dff_B_Xefk6Yl04_0),.clk(gclk));
	jdff dff_B_LnFfZrMQ4_0(.din(w_dff_B_Xefk6Yl04_0),.dout(w_dff_B_LnFfZrMQ4_0),.clk(gclk));
	jdff dff_B_vCCTPlxH9_1(.din(n1496),.dout(w_dff_B_vCCTPlxH9_1),.clk(gclk));
	jdff dff_B_KY4oClPQ5_1(.din(n413),.dout(w_dff_B_KY4oClPQ5_1),.clk(gclk));
	jdff dff_B_HKApNhrR4_1(.din(w_dff_B_KY4oClPQ5_1),.dout(w_dff_B_HKApNhrR4_1),.clk(gclk));
	jdff dff_A_ScLRp0dH0_0(.dout(w_G308_1[0]),.din(w_dff_A_ScLRp0dH0_0),.clk(gclk));
	jdff dff_B_IuHkOkDX2_1(.din(n400),.dout(w_dff_B_IuHkOkDX2_1),.clk(gclk));
	jdff dff_B_yyfaiPDj6_1(.din(w_dff_B_IuHkOkDX2_1),.dout(w_dff_B_yyfaiPDj6_1),.clk(gclk));
	jdff dff_A_ZpN0xOKU4_1(.dout(w_n428_0[1]),.din(w_dff_A_ZpN0xOKU4_1),.clk(gclk));
	jdff dff_B_8Xf7QnmY4_0(.din(n1493),.dout(w_dff_B_8Xf7QnmY4_0),.clk(gclk));
	jdff dff_A_S8jCp1lV4_0(.dout(w_G361_1[0]),.din(w_dff_A_S8jCp1lV4_0),.clk(gclk));
	jdff dff_B_4uGaUG2h6_1(.din(n1485),.dout(w_dff_B_4uGaUG2h6_1),.clk(gclk));
	jdff dff_A_JMj54jpY1_0(.dout(w_n437_0[0]),.din(w_dff_A_JMj54jpY1_0),.clk(gclk));
	jdff dff_B_SB3eUVwo7_2(.din(n437),.dout(w_dff_B_SB3eUVwo7_2),.clk(gclk));
	jdff dff_A_bqOqBG597_0(.dout(w_G503_2[0]),.din(w_dff_A_bqOqBG597_0),.clk(gclk));
	jdff dff_A_0rgalY9k1_0(.dout(w_dff_A_bqOqBG597_0),.din(w_dff_A_0rgalY9k1_0),.clk(gclk));
	jdff dff_A_PXTYXeMl1_0(.dout(w_dff_A_0rgalY9k1_0),.din(w_dff_A_PXTYXeMl1_0),.clk(gclk));
	jdff dff_B_EY5P9kkJ0_1(.din(n1481),.dout(w_dff_B_EY5P9kkJ0_1),.clk(gclk));
	jdff dff_B_xQ7tHhqd7_1(.din(n1471),.dout(w_dff_B_xQ7tHhqd7_1),.clk(gclk));
	jdff dff_B_3bgIAedx2_1(.din(w_dff_B_xQ7tHhqd7_1),.dout(w_dff_B_3bgIAedx2_1),.clk(gclk));
	jdff dff_A_F6B7u8qa1_1(.dout(w_G341_2[1]),.din(w_dff_A_F6B7u8qa1_1),.clk(gclk));
	jdff dff_B_TnwyGcai3_1(.din(n1462),.dout(w_dff_B_TnwyGcai3_1),.clk(gclk));
	jdff dff_B_Ifi5KaPP0_1(.din(w_dff_B_TnwyGcai3_1),.dout(w_dff_B_Ifi5KaPP0_1),.clk(gclk));
	jdff dff_A_ngYc9BaC7_1(.dout(w_G351_2[1]),.din(w_dff_A_ngYc9BaC7_1),.clk(gclk));
	jdff dff_B_z7gTYVop1_1(.din(n1453),.dout(w_dff_B_z7gTYVop1_1),.clk(gclk));
	jdff dff_A_V7FGggCU2_0(.dout(w_n749_5[0]),.din(w_dff_A_V7FGggCU2_0),.clk(gclk));
	jdff dff_A_yTmRByLd0_0(.dout(w_dff_A_V7FGggCU2_0),.din(w_dff_A_yTmRByLd0_0),.clk(gclk));
	jdff dff_A_aUEeXtDh7_0(.dout(w_dff_A_yTmRByLd0_0),.din(w_dff_A_aUEeXtDh7_0),.clk(gclk));
	jdff dff_A_ZGbPL6sO7_1(.dout(w_n749_5[1]),.din(w_dff_A_ZGbPL6sO7_1),.clk(gclk));
	jdff dff_A_xCDea2wl3_1(.dout(w_dff_A_ZGbPL6sO7_1),.din(w_dff_A_xCDea2wl3_1),.clk(gclk));
	jdff dff_A_gJgdEIrO5_1(.dout(w_dff_A_xCDea2wl3_1),.din(w_dff_A_gJgdEIrO5_1),.clk(gclk));
	jdff dff_A_QtdHhHKE0_1(.dout(w_dff_A_gJgdEIrO5_1),.din(w_dff_A_QtdHhHKE0_1),.clk(gclk));
	jdff dff_A_8mDJimVz1_1(.dout(w_dff_A_QtdHhHKE0_1),.din(w_dff_A_8mDJimVz1_1),.clk(gclk));
	jdff dff_A_FCBxGdyh3_1(.dout(w_dff_A_8mDJimVz1_1),.din(w_dff_A_FCBxGdyh3_1),.clk(gclk));
	jdff dff_A_h9R3Tg6B4_1(.dout(w_dff_A_FCBxGdyh3_1),.din(w_dff_A_h9R3Tg6B4_1),.clk(gclk));
	jdff dff_A_Bn8s0z5C4_1(.dout(w_dff_A_h9R3Tg6B4_1),.din(w_dff_A_Bn8s0z5C4_1),.clk(gclk));
	jdff dff_A_qWGh3QJT3_1(.dout(w_dff_A_Bn8s0z5C4_1),.din(w_dff_A_qWGh3QJT3_1),.clk(gclk));
	jdff dff_A_acbRl9gy2_1(.dout(w_dff_A_qWGh3QJT3_1),.din(w_dff_A_acbRl9gy2_1),.clk(gclk));
	jdff dff_A_GpYsJDvJ6_1(.dout(w_dff_A_acbRl9gy2_1),.din(w_dff_A_GpYsJDvJ6_1),.clk(gclk));
	jdff dff_A_Y5kv7rC74_1(.dout(w_dff_A_GpYsJDvJ6_1),.din(w_dff_A_Y5kv7rC74_1),.clk(gclk));
	jdff dff_B_99f1ywRJ4_0(.din(n1452),.dout(w_dff_B_99f1ywRJ4_0),.clk(gclk));
	jdff dff_A_ZotBMQ0D5_0(.dout(w_n1451_0[0]),.din(w_dff_A_ZotBMQ0D5_0),.clk(gclk));
	jdff dff_A_TmQHv6xl0_0(.dout(w_dff_A_ZotBMQ0D5_0),.din(w_dff_A_TmQHv6xl0_0),.clk(gclk));
	jdff dff_B_KKXQIs3M6_0(.din(n1450),.dout(w_dff_B_KKXQIs3M6_0),.clk(gclk));
	jdff dff_B_03kMr17E1_0(.din(w_dff_B_KKXQIs3M6_0),.dout(w_dff_B_03kMr17E1_0),.clk(gclk));
	jdff dff_B_c3XXmCf30_0(.din(w_dff_B_03kMr17E1_0),.dout(w_dff_B_c3XXmCf30_0),.clk(gclk));
	jdff dff_B_pC6Oo3Vw3_1(.din(n1448),.dout(w_dff_B_pC6Oo3Vw3_1),.clk(gclk));
	jdff dff_B_BwKl9oSn1_1(.din(w_dff_B_pC6Oo3Vw3_1),.dout(w_dff_B_BwKl9oSn1_1),.clk(gclk));
	jdff dff_B_HMWdFj7t1_1(.din(w_dff_B_BwKl9oSn1_1),.dout(w_dff_B_HMWdFj7t1_1),.clk(gclk));
	jdff dff_A_jOpFjveP9_0(.dout(w_n763_0[0]),.din(w_dff_A_jOpFjveP9_0),.clk(gclk));
	jdff dff_A_0WBcNEnh6_0(.dout(w_dff_A_jOpFjveP9_0),.din(w_dff_A_0WBcNEnh6_0),.clk(gclk));
	jdff dff_A_Colzfz4w2_0(.dout(w_dff_A_0WBcNEnh6_0),.din(w_dff_A_Colzfz4w2_0),.clk(gclk));
	jdff dff_A_2gaaYJ2z9_0(.dout(w_dff_A_Colzfz4w2_0),.din(w_dff_A_2gaaYJ2z9_0),.clk(gclk));
	jdff dff_A_pKK52SXc3_0(.dout(w_dff_A_2gaaYJ2z9_0),.din(w_dff_A_pKK52SXc3_0),.clk(gclk));
	jdff dff_A_zCWqs08e9_0(.dout(w_dff_A_pKK52SXc3_0),.din(w_dff_A_zCWqs08e9_0),.clk(gclk));
	jdff dff_A_ZDmExVea5_0(.dout(w_dff_A_zCWqs08e9_0),.din(w_dff_A_ZDmExVea5_0),.clk(gclk));
	jdff dff_A_Nh5iaij37_0(.dout(w_dff_A_ZDmExVea5_0),.din(w_dff_A_Nh5iaij37_0),.clk(gclk));
	jdff dff_B_gkOm9f2C8_1(.din(n1439),.dout(w_dff_B_gkOm9f2C8_1),.clk(gclk));
	jdff dff_B_X7h3zKJR7_1(.din(n1441),.dout(w_dff_B_X7h3zKJR7_1),.clk(gclk));
	jdff dff_B_HFXHnHTq0_0(.din(n1437),.dout(w_dff_B_HFXHnHTq0_0),.clk(gclk));
	jdff dff_B_YmCA8NpP5_0(.din(n1436),.dout(w_dff_B_YmCA8NpP5_0),.clk(gclk));
	jdff dff_A_fLKCUw2Z1_0(.dout(w_n1429_0[0]),.din(w_dff_A_fLKCUw2Z1_0),.clk(gclk));
	jdff dff_B_CGHTI8A53_1(.din(n1427),.dout(w_dff_B_CGHTI8A53_1),.clk(gclk));
	jdff dff_A_qr3O2Jyf8_2(.dout(w_n641_0[2]),.din(w_dff_A_qr3O2Jyf8_2),.clk(gclk));
	jdff dff_A_3lMUSRFd5_2(.dout(w_dff_A_qr3O2Jyf8_2),.din(w_dff_A_3lMUSRFd5_2),.clk(gclk));
	jdff dff_A_pp4HwyNl2_0(.dout(w_n640_0[0]),.din(w_dff_A_pp4HwyNl2_0),.clk(gclk));
	jdff dff_A_hISlCyLZ4_0(.dout(w_n639_0[0]),.din(w_dff_A_hISlCyLZ4_0),.clk(gclk));
	jdff dff_A_PUUWdHUJ7_0(.dout(w_n624_0[0]),.din(w_dff_A_PUUWdHUJ7_0),.clk(gclk));
	jdff dff_A_Jhn4XrRk4_0(.dout(w_dff_A_PUUWdHUJ7_0),.din(w_dff_A_Jhn4XrRk4_0),.clk(gclk));
	jdff dff_A_TizUnkPX5_1(.dout(w_n624_0[1]),.din(w_dff_A_TizUnkPX5_1),.clk(gclk));
	jdff dff_B_8fAdz1ZW7_3(.din(n624),.dout(w_dff_B_8fAdz1ZW7_3),.clk(gclk));
	jdff dff_B_XUuxerAk5_3(.din(w_dff_B_8fAdz1ZW7_3),.dout(w_dff_B_XUuxerAk5_3),.clk(gclk));
	jdff dff_A_SYi6c45J6_1(.dout(w_n620_1[1]),.din(w_dff_A_SYi6c45J6_1),.clk(gclk));
	jdff dff_A_3MEM3U4V7_1(.dout(w_dff_A_SYi6c45J6_1),.din(w_dff_A_3MEM3U4V7_1),.clk(gclk));
	jdff dff_A_3umru07q0_1(.dout(w_dff_A_3MEM3U4V7_1),.din(w_dff_A_3umru07q0_1),.clk(gclk));
	jdff dff_A_NHz2SRfK7_1(.dout(w_dff_A_3umru07q0_1),.din(w_dff_A_NHz2SRfK7_1),.clk(gclk));
	jdff dff_A_qHr140EL7_1(.dout(w_n620_0[1]),.din(w_dff_A_qHr140EL7_1),.clk(gclk));
	jdff dff_A_GwQxQH0o0_1(.dout(w_dff_A_qHr140EL7_1),.din(w_dff_A_GwQxQH0o0_1),.clk(gclk));
	jdff dff_A_pu0aBU7w3_2(.dout(w_n620_0[2]),.din(w_dff_A_pu0aBU7w3_2),.clk(gclk));
	jdff dff_A_B2AbRm9C6_2(.dout(w_dff_A_pu0aBU7w3_2),.din(w_dff_A_B2AbRm9C6_2),.clk(gclk));
	jdff dff_A_RzH3MoT43_2(.dout(w_dff_A_B2AbRm9C6_2),.din(w_dff_A_RzH3MoT43_2),.clk(gclk));
	jdff dff_A_UnQODbXq5_2(.dout(w_dff_A_RzH3MoT43_2),.din(w_dff_A_UnQODbXq5_2),.clk(gclk));
	jdff dff_A_QAGcJSPV5_2(.dout(w_dff_A_UnQODbXq5_2),.din(w_dff_A_QAGcJSPV5_2),.clk(gclk));
	jdff dff_A_fdnYTmS70_2(.dout(w_dff_A_QAGcJSPV5_2),.din(w_dff_A_fdnYTmS70_2),.clk(gclk));
	jdff dff_A_ioamGLlq1_2(.dout(w_dff_A_fdnYTmS70_2),.din(w_dff_A_ioamGLlq1_2),.clk(gclk));
	jdff dff_A_4Q6uc5GK7_1(.dout(w_n618_0[1]),.din(w_dff_A_4Q6uc5GK7_1),.clk(gclk));
	jdff dff_A_dsFZ2h5H1_1(.dout(w_dff_A_4Q6uc5GK7_1),.din(w_dff_A_dsFZ2h5H1_1),.clk(gclk));
	jdff dff_A_JL4ZPdIW2_1(.dout(w_dff_A_dsFZ2h5H1_1),.din(w_dff_A_JL4ZPdIW2_1),.clk(gclk));
	jdff dff_A_NFvJFWBi9_1(.dout(w_dff_A_JL4ZPdIW2_1),.din(w_dff_A_NFvJFWBi9_1),.clk(gclk));
	jdff dff_A_2ddUJsYP3_1(.dout(w_dff_A_NFvJFWBi9_1),.din(w_dff_A_2ddUJsYP3_1),.clk(gclk));
	jdff dff_A_zHayOKWN5_1(.dout(w_dff_A_2ddUJsYP3_1),.din(w_dff_A_zHayOKWN5_1),.clk(gclk));
	jdff dff_A_3tylgieY3_2(.dout(w_n618_0[2]),.din(w_dff_A_3tylgieY3_2),.clk(gclk));
	jdff dff_A_qBVbiEbx0_2(.dout(w_dff_A_3tylgieY3_2),.din(w_dff_A_qBVbiEbx0_2),.clk(gclk));
	jdff dff_A_XOM3sFug4_2(.dout(w_dff_A_qBVbiEbx0_2),.din(w_dff_A_XOM3sFug4_2),.clk(gclk));
	jdff dff_A_5WLf0liM1_0(.dout(w_n1425_0[0]),.din(w_dff_A_5WLf0liM1_0),.clk(gclk));
	jdff dff_B_T4kygeEA9_1(.din(n1411),.dout(w_dff_B_T4kygeEA9_1),.clk(gclk));
	jdff dff_A_O4Bg95WV8_0(.dout(w_n1422_0[0]),.din(w_dff_A_O4Bg95WV8_0),.clk(gclk));
	jdff dff_B_1KSxEyng2_1(.din(n1418),.dout(w_dff_B_1KSxEyng2_1),.clk(gclk));
	jdff dff_B_xjS2fJOz2_1(.din(w_dff_B_1KSxEyng2_1),.dout(w_dff_B_xjS2fJOz2_1),.clk(gclk));
	jdff dff_B_g9698oLR9_1(.din(w_dff_B_xjS2fJOz2_1),.dout(w_dff_B_g9698oLR9_1),.clk(gclk));
	jdff dff_B_CXq2RJea6_1(.din(n1419),.dout(w_dff_B_CXq2RJea6_1),.clk(gclk));
	jdff dff_B_fuURMbT48_1(.din(w_dff_B_CXq2RJea6_1),.dout(w_dff_B_fuURMbT48_1),.clk(gclk));
	jdff dff_A_8KmR0YJP9_2(.dout(w_n660_0[2]),.din(w_dff_A_8KmR0YJP9_2),.clk(gclk));
	jdff dff_A_snwGPB9Z3_2(.dout(w_dff_A_8KmR0YJP9_2),.din(w_dff_A_snwGPB9Z3_2),.clk(gclk));
	jdff dff_A_E2gla9Im8_2(.dout(w_dff_A_snwGPB9Z3_2),.din(w_dff_A_E2gla9Im8_2),.clk(gclk));
	jdff dff_A_lvIaQO0g4_2(.dout(w_dff_A_E2gla9Im8_2),.din(w_dff_A_lvIaQO0g4_2),.clk(gclk));
	jdff dff_A_8dtaMtdk8_2(.dout(w_dff_A_lvIaQO0g4_2),.din(w_dff_A_8dtaMtdk8_2),.clk(gclk));
	jdff dff_A_L4yrxRrg8_2(.dout(w_dff_A_8dtaMtdk8_2),.din(w_dff_A_L4yrxRrg8_2),.clk(gclk));
	jdff dff_A_PLnNkKAR6_2(.dout(w_n792_0[2]),.din(w_dff_A_PLnNkKAR6_2),.clk(gclk));
	jdff dff_A_tPGViu0P0_2(.dout(w_dff_A_PLnNkKAR6_2),.din(w_dff_A_tPGViu0P0_2),.clk(gclk));
	jdff dff_A_LiZCO5hy1_2(.dout(w_dff_A_tPGViu0P0_2),.din(w_dff_A_LiZCO5hy1_2),.clk(gclk));
	jdff dff_A_38fXQmRj4_2(.dout(w_dff_A_LiZCO5hy1_2),.din(w_dff_A_38fXQmRj4_2),.clk(gclk));
	jdff dff_A_JJd7wOE12_2(.dout(w_dff_A_38fXQmRj4_2),.din(w_dff_A_JJd7wOE12_2),.clk(gclk));
	jdff dff_A_NSJ5nVXs1_2(.dout(w_dff_A_JJd7wOE12_2),.din(w_dff_A_NSJ5nVXs1_2),.clk(gclk));
	jdff dff_A_slkS1ByX2_2(.dout(w_dff_A_NSJ5nVXs1_2),.din(w_dff_A_slkS1ByX2_2),.clk(gclk));
	jdff dff_A_N3Gq0osR5_2(.dout(w_dff_A_slkS1ByX2_2),.din(w_dff_A_N3Gq0osR5_2),.clk(gclk));
	jdff dff_A_68PoRUC35_2(.dout(w_dff_A_N3Gq0osR5_2),.din(w_dff_A_68PoRUC35_2),.clk(gclk));
	jdff dff_A_wo7kR2uM2_1(.dout(w_n790_0[1]),.din(w_dff_A_wo7kR2uM2_1),.clk(gclk));
	jdff dff_A_yLioJ1nj9_1(.dout(w_dff_A_wo7kR2uM2_1),.din(w_dff_A_yLioJ1nj9_1),.clk(gclk));
	jdff dff_A_lBhsoe5B3_1(.dout(w_dff_A_yLioJ1nj9_1),.din(w_dff_A_lBhsoe5B3_1),.clk(gclk));
	jdff dff_A_QNWnC9vh2_1(.dout(w_dff_A_lBhsoe5B3_1),.din(w_dff_A_QNWnC9vh2_1),.clk(gclk));
	jdff dff_A_xVD02jHt7_1(.dout(w_dff_A_QNWnC9vh2_1),.din(w_dff_A_xVD02jHt7_1),.clk(gclk));
	jdff dff_A_kgVQSWxH0_1(.dout(w_dff_A_xVD02jHt7_1),.din(w_dff_A_kgVQSWxH0_1),.clk(gclk));
	jdff dff_A_0fIJiKcG7_1(.dout(w_dff_A_kgVQSWxH0_1),.din(w_dff_A_0fIJiKcG7_1),.clk(gclk));
	jdff dff_A_jtqU0hGe6_1(.dout(w_dff_A_0fIJiKcG7_1),.din(w_dff_A_jtqU0hGe6_1),.clk(gclk));
	jdff dff_A_54lJdxHT6_1(.dout(w_dff_A_jtqU0hGe6_1),.din(w_dff_A_54lJdxHT6_1),.clk(gclk));
	jdff dff_A_4MuFKhJy2_1(.dout(w_dff_A_54lJdxHT6_1),.din(w_dff_A_4MuFKhJy2_1),.clk(gclk));
	jdff dff_B_9CdaUsTE7_1(.din(n1413),.dout(w_dff_B_9CdaUsTE7_1),.clk(gclk));
	jdff dff_B_IcLk55ca2_1(.din(w_dff_B_9CdaUsTE7_1),.dout(w_dff_B_IcLk55ca2_1),.clk(gclk));
	jdff dff_B_2Y962Pvs2_1(.din(w_dff_B_IcLk55ca2_1),.dout(w_dff_B_2Y962Pvs2_1),.clk(gclk));
	jdff dff_B_Qoa6Ht6s8_1(.din(w_dff_B_2Y962Pvs2_1),.dout(w_dff_B_Qoa6Ht6s8_1),.clk(gclk));
	jdff dff_B_S0q4jkJ69_1(.din(n1414),.dout(w_dff_B_S0q4jkJ69_1),.clk(gclk));
	jdff dff_B_7ueIVrlP4_1(.din(w_dff_B_S0q4jkJ69_1),.dout(w_dff_B_7ueIVrlP4_1),.clk(gclk));
	jdff dff_B_mAlA7HAG8_1(.din(w_dff_B_7ueIVrlP4_1),.dout(w_dff_B_mAlA7HAG8_1),.clk(gclk));
	jdff dff_A_mfsUWL0M9_1(.dout(w_n821_0[1]),.din(w_dff_A_mfsUWL0M9_1),.clk(gclk));
	jdff dff_B_0iqja61s8_1(.din(n812),.dout(w_dff_B_0iqja61s8_1),.clk(gclk));
	jdff dff_B_EKjZM2YP1_1(.din(w_dff_B_0iqja61s8_1),.dout(w_dff_B_EKjZM2YP1_1),.clk(gclk));
	jdff dff_B_8z1ZQthU8_1(.din(w_dff_B_EKjZM2YP1_1),.dout(w_dff_B_8z1ZQthU8_1),.clk(gclk));
	jdff dff_B_WzlzO9Pe6_1(.din(w_dff_B_8z1ZQthU8_1),.dout(w_dff_B_WzlzO9Pe6_1),.clk(gclk));
	jdff dff_B_xABjFLal2_1(.din(n813),.dout(w_dff_B_xABjFLal2_1),.clk(gclk));
	jdff dff_B_X11dDHA70_1(.din(w_dff_B_xABjFLal2_1),.dout(w_dff_B_X11dDHA70_1),.clk(gclk));
	jdff dff_B_N0rTAIrb9_1(.din(w_dff_B_X11dDHA70_1),.dout(w_dff_B_N0rTAIrb9_1),.clk(gclk));
	jdff dff_A_ls8UL0Zm0_1(.dout(w_n819_0[1]),.din(w_dff_A_ls8UL0Zm0_1),.clk(gclk));
	jdff dff_A_IYJMrDp93_1(.dout(w_dff_A_ls8UL0Zm0_1),.din(w_dff_A_IYJMrDp93_1),.clk(gclk));
	jdff dff_A_iWDqtKCR1_0(.dout(w_n377_1[0]),.din(w_dff_A_iWDqtKCR1_0),.clk(gclk));
	jdff dff_A_wS2vt67i1_0(.dout(w_n814_0[0]),.din(w_dff_A_wS2vt67i1_0),.clk(gclk));
	jdff dff_A_2ZtELZvn1_0(.dout(w_dff_A_wS2vt67i1_0),.din(w_dff_A_2ZtELZvn1_0),.clk(gclk));
	jdff dff_A_12ZkINdP0_0(.dout(w_dff_A_2ZtELZvn1_0),.din(w_dff_A_12ZkINdP0_0),.clk(gclk));
	jdff dff_A_z7p6YUjr6_1(.dout(w_n814_0[1]),.din(w_dff_A_z7p6YUjr6_1),.clk(gclk));
	jdff dff_A_TJs1W6DT4_1(.dout(w_dff_A_z7p6YUjr6_1),.din(w_dff_A_TJs1W6DT4_1),.clk(gclk));
	jdff dff_A_Gva3RcoY4_2(.dout(w_n377_0[2]),.din(w_dff_A_Gva3RcoY4_2),.clk(gclk));
	jdff dff_B_8YMo3sLn6_3(.din(n377),.dout(w_dff_B_8YMo3sLn6_3),.clk(gclk));
	jdff dff_A_eNIehFkN6_0(.dout(w_G534_2[0]),.din(w_dff_A_eNIehFkN6_0),.clk(gclk));
	jdff dff_A_9sijSR7X7_0(.dout(w_dff_A_eNIehFkN6_0),.din(w_dff_A_9sijSR7X7_0),.clk(gclk));
	jdff dff_A_YeTVb28I2_0(.dout(w_dff_A_9sijSR7X7_0),.din(w_dff_A_YeTVb28I2_0),.clk(gclk));
	jdff dff_A_uj2YxGOe0_1(.dout(w_n1412_0[1]),.din(w_dff_A_uj2YxGOe0_1),.clk(gclk));
	jdff dff_A_uacR1U299_1(.dout(w_dff_A_uj2YxGOe0_1),.din(w_dff_A_uacR1U299_1),.clk(gclk));
	jdff dff_A_7rkIrt1C7_2(.dout(w_n1412_0[2]),.din(w_dff_A_7rkIrt1C7_2),.clk(gclk));
	jdff dff_B_PgG8jdQ65_3(.din(n1412),.dout(w_dff_B_PgG8jdQ65_3),.clk(gclk));
	jdff dff_B_G1Da8Jhw2_3(.din(w_dff_B_PgG8jdQ65_3),.dout(w_dff_B_G1Da8Jhw2_3),.clk(gclk));
	jdff dff_B_Z2ESZr7E7_3(.din(w_dff_B_G1Da8Jhw2_3),.dout(w_dff_B_Z2ESZr7E7_3),.clk(gclk));
	jdff dff_B_FP36ZvEP7_3(.din(w_dff_B_Z2ESZr7E7_3),.dout(w_dff_B_FP36ZvEP7_3),.clk(gclk));
	jdff dff_B_H0CS5pZQ4_3(.din(w_dff_B_FP36ZvEP7_3),.dout(w_dff_B_H0CS5pZQ4_3),.clk(gclk));
	jdff dff_B_3ffLWUqT4_3(.din(w_dff_B_H0CS5pZQ4_3),.dout(w_dff_B_3ffLWUqT4_3),.clk(gclk));
	jdff dff_B_nUYSVcto3_3(.din(w_dff_B_3ffLWUqT4_3),.dout(w_dff_B_nUYSVcto3_3),.clk(gclk));
	jdff dff_B_Fvxerrtk9_3(.din(w_dff_B_nUYSVcto3_3),.dout(w_dff_B_Fvxerrtk9_3),.clk(gclk));
	jdff dff_B_sdwmjEXH9_3(.din(w_dff_B_Fvxerrtk9_3),.dout(w_dff_B_sdwmjEXH9_3),.clk(gclk));
	jdff dff_B_1mfQGzjy0_3(.din(w_dff_B_sdwmjEXH9_3),.dout(w_dff_B_1mfQGzjy0_3),.clk(gclk));
	jdff dff_A_rBMiAk2D1_0(.dout(w_G2174_0[0]),.din(w_dff_A_rBMiAk2D1_0),.clk(gclk));
	jdff dff_A_OCUCIsPn8_0(.dout(w_dff_A_rBMiAk2D1_0),.din(w_dff_A_OCUCIsPn8_0),.clk(gclk));
	jdff dff_A_Rs7jDHPV2_0(.dout(w_dff_A_OCUCIsPn8_0),.din(w_dff_A_Rs7jDHPV2_0),.clk(gclk));
	jdff dff_A_GzMljIXB9_0(.dout(w_dff_A_Rs7jDHPV2_0),.din(w_dff_A_GzMljIXB9_0),.clk(gclk));
	jdff dff_A_AbNsvuMK8_0(.dout(w_dff_A_GzMljIXB9_0),.din(w_dff_A_AbNsvuMK8_0),.clk(gclk));
	jdff dff_A_LcXRCDil6_0(.dout(w_dff_A_AbNsvuMK8_0),.din(w_dff_A_LcXRCDil6_0),.clk(gclk));
	jdff dff_A_kBWWMt8I3_0(.dout(w_dff_A_LcXRCDil6_0),.din(w_dff_A_kBWWMt8I3_0),.clk(gclk));
	jdff dff_A_5Rwlu8WZ7_0(.dout(w_dff_A_kBWWMt8I3_0),.din(w_dff_A_5Rwlu8WZ7_0),.clk(gclk));
	jdff dff_A_J0FTVxWY9_0(.dout(w_dff_A_5Rwlu8WZ7_0),.din(w_dff_A_J0FTVxWY9_0),.clk(gclk));
	jdff dff_A_mkjfvBAA2_0(.dout(w_dff_A_J0FTVxWY9_0),.din(w_dff_A_mkjfvBAA2_0),.clk(gclk));
	jdff dff_A_xNidbHy21_0(.dout(w_dff_A_mkjfvBAA2_0),.din(w_dff_A_xNidbHy21_0),.clk(gclk));
	jdff dff_A_HzJQC4BY7_0(.dout(w_dff_A_xNidbHy21_0),.din(w_dff_A_HzJQC4BY7_0),.clk(gclk));
	jdff dff_A_Jsb5G67L3_0(.dout(w_dff_A_HzJQC4BY7_0),.din(w_dff_A_Jsb5G67L3_0),.clk(gclk));
	jdff dff_A_3XgOyV4A3_1(.dout(w_G2174_0[1]),.din(w_dff_A_3XgOyV4A3_1),.clk(gclk));
	jdff dff_A_l5Fp4qqx5_1(.dout(w_dff_A_3XgOyV4A3_1),.din(w_dff_A_l5Fp4qqx5_1),.clk(gclk));
	jdff dff_A_RpzViQAF7_1(.dout(w_dff_A_l5Fp4qqx5_1),.din(w_dff_A_RpzViQAF7_1),.clk(gclk));
	jdff dff_A_FKCEAtMd9_1(.dout(w_dff_A_RpzViQAF7_1),.din(w_dff_A_FKCEAtMd9_1),.clk(gclk));
	jdff dff_A_4leJHROL5_1(.dout(w_dff_A_FKCEAtMd9_1),.din(w_dff_A_4leJHROL5_1),.clk(gclk));
	jdff dff_A_kt02p7lV7_1(.dout(w_dff_A_4leJHROL5_1),.din(w_dff_A_kt02p7lV7_1),.clk(gclk));
	jdff dff_A_FcLCn6tK6_1(.dout(w_dff_A_kt02p7lV7_1),.din(w_dff_A_FcLCn6tK6_1),.clk(gclk));
	jdff dff_A_tRzY0CQz2_1(.dout(w_dff_A_FcLCn6tK6_1),.din(w_dff_A_tRzY0CQz2_1),.clk(gclk));
	jdff dff_A_0oDtY7i71_1(.dout(w_dff_A_tRzY0CQz2_1),.din(w_dff_A_0oDtY7i71_1),.clk(gclk));
	jdff dff_A_ibm6KBV90_1(.dout(w_dff_A_0oDtY7i71_1),.din(w_dff_A_ibm6KBV90_1),.clk(gclk));
	jdff dff_A_xGYv2QMQ1_0(.dout(w_n1410_0[0]),.din(w_dff_A_xGYv2QMQ1_0),.clk(gclk));
	jdff dff_B_96UzNQdT7_0(.din(n1409),.dout(w_dff_B_96UzNQdT7_0),.clk(gclk));
	jdff dff_B_T4ChUrjp5_0(.din(w_dff_B_96UzNQdT7_0),.dout(w_dff_B_T4ChUrjp5_0),.clk(gclk));
	jdff dff_A_c6y1Byqp4_0(.dout(w_n401_0[0]),.din(w_dff_A_c6y1Byqp4_0),.clk(gclk));
	jdff dff_A_akJRuCx35_0(.dout(w_dff_A_c6y1Byqp4_0),.din(w_dff_A_akJRuCx35_0),.clk(gclk));
	jdff dff_A_TG9rKCVs5_0(.dout(w_dff_A_akJRuCx35_0),.din(w_dff_A_TG9rKCVs5_0),.clk(gclk));
	jdff dff_B_dxrmcj3p8_2(.din(n401),.dout(w_dff_B_dxrmcj3p8_2),.clk(gclk));
	jdff dff_A_BCOMpbI92_0(.dout(w_G490_1[0]),.din(w_dff_A_BCOMpbI92_0),.clk(gclk));
	jdff dff_A_jIE75rIy5_0(.dout(w_dff_A_BCOMpbI92_0),.din(w_dff_A_jIE75rIy5_0),.clk(gclk));
	jdff dff_A_DlOB61Du6_0(.dout(w_dff_A_jIE75rIy5_0),.din(w_dff_A_DlOB61Du6_0),.clk(gclk));
	jdff dff_A_fl2XX5NO3_1(.dout(w_n654_1[1]),.din(w_dff_A_fl2XX5NO3_1),.clk(gclk));
	jdff dff_A_KzDCsPxR0_1(.dout(w_dff_A_fl2XX5NO3_1),.din(w_dff_A_KzDCsPxR0_1),.clk(gclk));
	jdff dff_A_CuvyOiKi4_1(.dout(w_dff_A_KzDCsPxR0_1),.din(w_dff_A_CuvyOiKi4_1),.clk(gclk));
	jdff dff_A_CseopRmD1_1(.dout(w_dff_A_CuvyOiKi4_1),.din(w_dff_A_CseopRmD1_1),.clk(gclk));
	jdff dff_A_DtV5yOsa7_1(.dout(w_dff_A_CseopRmD1_1),.din(w_dff_A_DtV5yOsa7_1),.clk(gclk));
	jdff dff_A_Av5iEvP98_1(.dout(w_dff_A_DtV5yOsa7_1),.din(w_dff_A_Av5iEvP98_1),.clk(gclk));
	jdff dff_A_cY01WQiF5_1(.dout(w_dff_A_Av5iEvP98_1),.din(w_dff_A_cY01WQiF5_1),.clk(gclk));
	jdff dff_A_8SolGUlR1_1(.dout(w_dff_A_cY01WQiF5_1),.din(w_dff_A_8SolGUlR1_1),.clk(gclk));
	jdff dff_A_MaZmCqmi6_0(.dout(w_n644_0[0]),.din(w_dff_A_MaZmCqmi6_0),.clk(gclk));
	jdff dff_A_7DuDT1AJ7_0(.dout(w_dff_A_MaZmCqmi6_0),.din(w_dff_A_7DuDT1AJ7_0),.clk(gclk));
	jdff dff_A_y04Tg1jh5_0(.dout(w_dff_A_7DuDT1AJ7_0),.din(w_dff_A_y04Tg1jh5_0),.clk(gclk));
	jdff dff_A_YnXvQpkT4_0(.dout(w_dff_A_y04Tg1jh5_0),.din(w_dff_A_YnXvQpkT4_0),.clk(gclk));
	jdff dff_A_KcQBLqEE2_2(.dout(w_n644_0[2]),.din(w_dff_A_KcQBLqEE2_2),.clk(gclk));
	jdff dff_A_lxg9sKrs5_2(.dout(w_dff_A_KcQBLqEE2_2),.din(w_dff_A_lxg9sKrs5_2),.clk(gclk));
	jdff dff_A_ohMqcqoZ8_1(.dout(w_G293_0[1]),.din(w_dff_A_ohMqcqoZ8_1),.clk(gclk));
	jdff dff_A_IkZ0w3dF1_1(.dout(w_n746_0[1]),.din(w_dff_A_IkZ0w3dF1_1),.clk(gclk));
	jdff dff_A_LIpZI4sY9_1(.dout(w_dff_A_IkZ0w3dF1_1),.din(w_dff_A_LIpZI4sY9_1),.clk(gclk));
	jdff dff_A_h9jhfxll5_1(.dout(w_dff_A_LIpZI4sY9_1),.din(w_dff_A_h9jhfxll5_1),.clk(gclk));
	jdff dff_A_1cjKdCl93_1(.dout(w_dff_A_h9jhfxll5_1),.din(w_dff_A_1cjKdCl93_1),.clk(gclk));
	jdff dff_B_L78YjEUY2_1(.din(n741),.dout(w_dff_B_L78YjEUY2_1),.clk(gclk));
	jdff dff_B_6s7BJUn44_1(.din(w_dff_B_L78YjEUY2_1),.dout(w_dff_B_6s7BJUn44_1),.clk(gclk));
	jdff dff_A_bMOUi0UJ9_1(.dout(w_n742_0[1]),.din(w_dff_A_bMOUi0UJ9_1),.clk(gclk));
	jdff dff_A_mU1xbz8d0_1(.dout(w_dff_A_bMOUi0UJ9_1),.din(w_dff_A_mU1xbz8d0_1),.clk(gclk));
	jdff dff_A_89hbxUXa5_1(.dout(w_dff_A_mU1xbz8d0_1),.din(w_dff_A_89hbxUXa5_1),.clk(gclk));
	jdff dff_A_9WVpNVBm1_1(.dout(w_dff_A_89hbxUXa5_1),.din(w_dff_A_9WVpNVBm1_1),.clk(gclk));
	jdff dff_A_sinFkYgd5_1(.dout(w_dff_A_9WVpNVBm1_1),.din(w_dff_A_sinFkYgd5_1),.clk(gclk));
	jdff dff_A_Y2fP7vZz7_1(.dout(w_dff_A_sinFkYgd5_1),.din(w_dff_A_Y2fP7vZz7_1),.clk(gclk));
	jdff dff_A_QbkPiTFN8_1(.dout(w_dff_A_Y2fP7vZz7_1),.din(w_dff_A_QbkPiTFN8_1),.clk(gclk));
	jdff dff_B_asLk4WND6_0(.din(n657),.dout(w_dff_B_asLk4WND6_0),.clk(gclk));
	jdff dff_B_tschl8w45_1(.din(G323),.dout(w_dff_B_tschl8w45_1),.clk(gclk));
	jdff dff_A_gRwoKJ1I1_2(.dout(w_G316_0[2]),.din(w_dff_A_gRwoKJ1I1_2),.clk(gclk));
	jdff dff_A_9Xax7Uze0_1(.dout(w_G490_0[1]),.din(w_dff_A_9Xax7Uze0_1),.clk(gclk));
	jdff dff_A_WFQWTIZ04_1(.dout(w_dff_A_9Xax7Uze0_1),.din(w_dff_A_WFQWTIZ04_1),.clk(gclk));
	jdff dff_A_YhHvhUHd6_1(.dout(w_dff_A_WFQWTIZ04_1),.din(w_dff_A_YhHvhUHd6_1),.clk(gclk));
	jdff dff_A_S77Krj036_1(.dout(w_dff_A_YhHvhUHd6_1),.din(w_dff_A_S77Krj036_1),.clk(gclk));
	jdff dff_A_ebeDXyY83_2(.dout(w_G490_0[2]),.din(w_dff_A_ebeDXyY83_2),.clk(gclk));
	jdff dff_A_D8d91TvS3_2(.dout(w_dff_A_ebeDXyY83_2),.din(w_dff_A_D8d91TvS3_2),.clk(gclk));
	jdff dff_A_UsOjqMgw6_2(.dout(w_dff_A_D8d91TvS3_2),.din(w_dff_A_UsOjqMgw6_2),.clk(gclk));
	jdff dff_A_lcGgPAjg9_2(.dout(w_dff_A_UsOjqMgw6_2),.din(w_dff_A_lcGgPAjg9_2),.clk(gclk));
	jdff dff_A_xFdiiL3z1_0(.dout(w_n654_2[0]),.din(w_dff_A_xFdiiL3z1_0),.clk(gclk));
	jdff dff_A_BrKvvSPn1_0(.dout(w_n654_0[0]),.din(w_dff_A_BrKvvSPn1_0),.clk(gclk));
	jdff dff_B_r3BFdL1o3_3(.din(n654),.dout(w_dff_B_r3BFdL1o3_3),.clk(gclk));
	jdff dff_A_qKiqqAVL5_0(.dout(w_n653_0[0]),.din(w_dff_A_qKiqqAVL5_0),.clk(gclk));
	jdff dff_B_xOOQgFa32_1(.din(n651),.dout(w_dff_B_xOOQgFa32_1),.clk(gclk));
	jdff dff_B_IrD5C1yu8_1(.din(G315),.dout(w_dff_B_IrD5C1yu8_1),.clk(gclk));
	jdff dff_A_Xsngfe2U3_0(.dout(w_n414_0[0]),.din(w_dff_A_Xsngfe2U3_0),.clk(gclk));
	jdff dff_A_f4tHy0gm6_0(.dout(w_dff_A_Xsngfe2U3_0),.din(w_dff_A_f4tHy0gm6_0),.clk(gclk));
	jdff dff_B_zrNIoY7t3_2(.din(n414),.dout(w_dff_B_zrNIoY7t3_2),.clk(gclk));
	jdff dff_A_exMnkZjk4_0(.dout(w_G479_0[0]),.din(w_dff_A_exMnkZjk4_0),.clk(gclk));
	jdff dff_A_fwH1ofpW3_0(.dout(w_dff_A_exMnkZjk4_0),.din(w_dff_A_fwH1ofpW3_0),.clk(gclk));
	jdff dff_A_U2B1WQkS2_0(.dout(w_dff_A_fwH1ofpW3_0),.din(w_dff_A_U2B1WQkS2_0),.clk(gclk));
	jdff dff_A_ktMtPHfW7_1(.dout(w_G479_0[1]),.din(w_dff_A_ktMtPHfW7_1),.clk(gclk));
	jdff dff_A_LtTTofiA0_1(.dout(w_dff_A_ktMtPHfW7_1),.din(w_dff_A_LtTTofiA0_1),.clk(gclk));
	jdff dff_A_EbD5XZ6A1_1(.dout(w_dff_A_LtTTofiA0_1),.din(w_dff_A_EbD5XZ6A1_1),.clk(gclk));
	jdff dff_A_5E871zXd0_1(.dout(w_n648_0[1]),.din(w_dff_A_5E871zXd0_1),.clk(gclk));
	jdff dff_A_jkidX6wY6_1(.dout(w_dff_A_5E871zXd0_1),.din(w_dff_A_jkidX6wY6_1),.clk(gclk));
	jdff dff_A_FpBvAnXV4_1(.dout(w_dff_A_jkidX6wY6_1),.din(w_dff_A_FpBvAnXV4_1),.clk(gclk));
	jdff dff_A_hVwjUmak5_1(.dout(w_dff_A_FpBvAnXV4_1),.din(w_dff_A_hVwjUmak5_1),.clk(gclk));
	jdff dff_A_gEJ9SdA75_2(.dout(w_n648_0[2]),.din(w_dff_A_gEJ9SdA75_2),.clk(gclk));
	jdff dff_A_Uo8RRHtf5_2(.dout(w_dff_A_gEJ9SdA75_2),.din(w_dff_A_Uo8RRHtf5_2),.clk(gclk));
	jdff dff_A_JuVocacq3_2(.dout(w_dff_A_Uo8RRHtf5_2),.din(w_dff_A_JuVocacq3_2),.clk(gclk));
	jdff dff_A_GgqagvSJ3_2(.dout(w_dff_A_JuVocacq3_2),.din(w_dff_A_GgqagvSJ3_2),.clk(gclk));
	jdff dff_A_E5nnNKxj8_2(.dout(w_dff_A_GgqagvSJ3_2),.din(w_dff_A_E5nnNKxj8_2),.clk(gclk));
	jdff dff_B_J7QSLHkv8_0(.din(n647),.dout(w_dff_B_J7QSLHkv8_0),.clk(gclk));
	jdff dff_B_G0FqcR0X5_1(.din(G307),.dout(w_dff_B_G0FqcR0X5_1),.clk(gclk));
	jdff dff_A_etQq017Q2_0(.dout(w_G302_0[0]),.din(w_dff_A_etQq017Q2_0),.clk(gclk));
	jdff dff_A_kGtQubRU4_1(.dout(w_G302_0[1]),.din(w_dff_A_kGtQubRU4_1),.clk(gclk));
	jdff dff_B_h14bxRSR8_1(.din(n727),.dout(w_dff_B_h14bxRSR8_1),.clk(gclk));
	jdff dff_A_UPDBQr5m9_0(.dout(w_n635_1[0]),.din(w_dff_A_UPDBQr5m9_0),.clk(gclk));
	jdff dff_A_xmHMGbPn5_1(.dout(w_n635_0[1]),.din(w_dff_A_xmHMGbPn5_1),.clk(gclk));
	jdff dff_A_1wofKjqD7_1(.dout(w_dff_A_xmHMGbPn5_1),.din(w_dff_A_1wofKjqD7_1),.clk(gclk));
	jdff dff_B_Ye6HFRXg6_1(.din(n633),.dout(w_dff_B_Ye6HFRXg6_1),.clk(gclk));
	jdff dff_A_MJ0ViibJ4_0(.dout(w_G366_0[0]),.din(w_dff_A_MJ0ViibJ4_0),.clk(gclk));
	jdff dff_A_ebIdPORu4_0(.dout(w_G332_2[0]),.din(w_dff_A_ebIdPORu4_0),.clk(gclk));
	jdff dff_A_5elyxUXx2_2(.dout(w_G332_2[2]),.din(w_dff_A_5elyxUXx2_2),.clk(gclk));
	jdff dff_A_HMrfA5Gf4_0(.dout(w_n628_0[0]),.din(w_dff_A_HMrfA5Gf4_0),.clk(gclk));
	jdff dff_A_pQe7xHr40_0(.dout(w_dff_A_HMrfA5Gf4_0),.din(w_dff_A_pQe7xHr40_0),.clk(gclk));
	jdff dff_A_nGDxQYAn0_0(.dout(w_dff_A_pQe7xHr40_0),.din(w_dff_A_nGDxQYAn0_0),.clk(gclk));
	jdff dff_A_iHYFifiN4_2(.dout(w_n628_0[2]),.din(w_dff_A_iHYFifiN4_2),.clk(gclk));
	jdff dff_A_qeIdu1Xg2_0(.dout(w_G358_0[0]),.din(w_dff_A_qeIdu1Xg2_0),.clk(gclk));
	jdff dff_A_jmzSzmoB4_1(.dout(w_n625_0[1]),.din(w_dff_A_jmzSzmoB4_1),.clk(gclk));
	jdff dff_A_SNlAwwOi8_2(.dout(w_G351_0[2]),.din(w_dff_A_SNlAwwOi8_2),.clk(gclk));
	jdff dff_A_5ATc7Gsn9_0(.dout(w_G534_0[0]),.din(w_dff_A_5ATc7Gsn9_0),.clk(gclk));
	jdff dff_A_u6gIaMjr6_0(.dout(w_dff_A_5ATc7Gsn9_0),.din(w_dff_A_u6gIaMjr6_0),.clk(gclk));
	jdff dff_A_LAEMmbVG5_0(.dout(w_dff_A_u6gIaMjr6_0),.din(w_dff_A_LAEMmbVG5_0),.clk(gclk));
	jdff dff_A_0Z1fpFhw9_2(.dout(w_G534_0[2]),.din(w_dff_A_0Z1fpFhw9_2),.clk(gclk));
	jdff dff_A_h2orIroB3_2(.dout(w_dff_A_0Z1fpFhw9_2),.din(w_dff_A_h2orIroB3_2),.clk(gclk));
	jdff dff_A_uz8yns7j3_2(.dout(w_dff_A_h2orIroB3_2),.din(w_dff_A_uz8yns7j3_2),.clk(gclk));
	jdff dff_A_wogrT4di4_0(.dout(w_n726_0[0]),.din(w_dff_A_wogrT4di4_0),.clk(gclk));
	jdff dff_A_qDepDr3V9_0(.dout(w_dff_A_wogrT4di4_0),.din(w_dff_A_qDepDr3V9_0),.clk(gclk));
	jdff dff_A_hItFPknl1_0(.dout(w_G348_0[0]),.din(w_dff_A_hItFPknl1_0),.clk(gclk));
	jdff dff_A_FPSHAf153_1(.dout(w_G332_1[1]),.din(w_dff_A_FPSHAf153_1),.clk(gclk));
	jdff dff_A_tpYJbV0X3_1(.dout(w_n621_0[1]),.din(w_dff_A_tpYJbV0X3_1),.clk(gclk));
	jdff dff_A_r9ppHhem0_2(.dout(w_G341_0[2]),.din(w_dff_A_r9ppHhem0_2),.clk(gclk));
	jdff dff_A_vNWGVL5O1_0(.dout(w_n389_1[0]),.din(w_dff_A_vNWGVL5O1_0),.clk(gclk));
	jdff dff_A_jcIciAi55_2(.dout(w_n389_0[2]),.din(w_dff_A_jcIciAi55_2),.clk(gclk));
	jdff dff_B_43Qwqhk89_3(.din(n389),.dout(w_dff_B_43Qwqhk89_3),.clk(gclk));
	jdff dff_A_y5zcxQJw1_0(.dout(w_G523_1[0]),.din(w_dff_A_y5zcxQJw1_0),.clk(gclk));
	jdff dff_A_58qlD1fI5_0(.dout(w_dff_A_y5zcxQJw1_0),.din(w_dff_A_58qlD1fI5_0),.clk(gclk));
	jdff dff_A_RzdvU1OF3_0(.dout(w_dff_A_58qlD1fI5_0),.din(w_dff_A_RzdvU1OF3_0),.clk(gclk));
	jdff dff_A_jc1tYchS5_1(.dout(w_G523_1[1]),.din(w_dff_A_jc1tYchS5_1),.clk(gclk));
	jdff dff_A_lp7GHm1F6_1(.dout(w_dff_A_jc1tYchS5_1),.din(w_dff_A_lp7GHm1F6_1),.clk(gclk));
	jdff dff_A_5oDTPYdf1_1(.dout(w_dff_A_lp7GHm1F6_1),.din(w_dff_A_5oDTPYdf1_1),.clk(gclk));
	jdff dff_A_yoxJaAYq4_1(.dout(w_G523_0[1]),.din(w_dff_A_yoxJaAYq4_1),.clk(gclk));
	jdff dff_A_nbuYs9md5_1(.dout(w_dff_A_yoxJaAYq4_1),.din(w_dff_A_nbuYs9md5_1),.clk(gclk));
	jdff dff_A_w06BWhO72_1(.dout(w_dff_A_nbuYs9md5_1),.din(w_dff_A_w06BWhO72_1),.clk(gclk));
	jdff dff_A_toLwCWIm7_2(.dout(w_G523_0[2]),.din(w_dff_A_toLwCWIm7_2),.clk(gclk));
	jdff dff_A_4lpIsodn8_2(.dout(w_dff_A_toLwCWIm7_2),.din(w_dff_A_4lpIsodn8_2),.clk(gclk));
	jdff dff_A_jo6hae3s0_2(.dout(w_dff_A_4lpIsodn8_2),.din(w_dff_A_jo6hae3s0_2),.clk(gclk));
	jdff dff_A_95nW45hR3_1(.dout(w_n722_0[1]),.din(w_dff_A_95nW45hR3_1),.clk(gclk));
	jdff dff_A_Ud1hYCRi0_1(.dout(w_dff_A_95nW45hR3_1),.din(w_dff_A_Ud1hYCRi0_1),.clk(gclk));
	jdff dff_A_qV2cdtfx4_1(.dout(w_dff_A_Ud1hYCRi0_1),.din(w_dff_A_qV2cdtfx4_1),.clk(gclk));
	jdff dff_A_8hthiOcC1_1(.dout(w_dff_A_qV2cdtfx4_1),.din(w_dff_A_8hthiOcC1_1),.clk(gclk));
	jdff dff_A_mwgLu1SD4_1(.dout(w_n721_0[1]),.din(w_dff_A_mwgLu1SD4_1),.clk(gclk));
	jdff dff_A_lCkwKWrU1_1(.dout(w_dff_A_mwgLu1SD4_1),.din(w_dff_A_lCkwKWrU1_1),.clk(gclk));
	jdff dff_A_M4yv3f1H0_1(.dout(w_dff_A_lCkwKWrU1_1),.din(w_dff_A_M4yv3f1H0_1),.clk(gclk));
	jdff dff_A_I7cHtpOf1_1(.dout(w_dff_A_M4yv3f1H0_1),.din(w_dff_A_I7cHtpOf1_1),.clk(gclk));
	jdff dff_A_XKG0JAaY6_1(.dout(w_dff_A_I7cHtpOf1_1),.din(w_dff_A_XKG0JAaY6_1),.clk(gclk));
	jdff dff_A_pdF4pMba5_1(.dout(w_n619_0[1]),.din(w_dff_A_pdF4pMba5_1),.clk(gclk));
	jdff dff_A_ZNLjUrh03_1(.dout(w_dff_A_pdF4pMba5_1),.din(w_dff_A_ZNLjUrh03_1),.clk(gclk));
	jdff dff_A_RfHlSoqf7_0(.dout(w_G338_0[0]),.din(w_dff_A_RfHlSoqf7_0),.clk(gclk));
	jdff dff_A_PQmDPWnJ9_0(.dout(w_G514_0[0]),.din(w_dff_A_PQmDPWnJ9_0),.clk(gclk));
	jdff dff_A_3n8RWLgq4_0(.dout(w_dff_A_PQmDPWnJ9_0),.din(w_dff_A_3n8RWLgq4_0),.clk(gclk));
	jdff dff_A_khKlBzin5_2(.dout(w_G514_0[2]),.din(w_dff_A_khKlBzin5_2),.clk(gclk));
	jdff dff_A_zBOEPcfw3_1(.dout(w_n720_0[1]),.din(w_dff_A_zBOEPcfw3_1),.clk(gclk));
	jdff dff_A_qwX6CVHe2_1(.dout(w_dff_A_zBOEPcfw3_1),.din(w_dff_A_qwX6CVHe2_1),.clk(gclk));
	jdff dff_A_A6QyrXHa2_1(.dout(w_dff_A_qwX6CVHe2_1),.din(w_dff_A_A6QyrXHa2_1),.clk(gclk));
	jdff dff_A_p4Fayc1v9_1(.dout(w_dff_A_A6QyrXHa2_1),.din(w_dff_A_p4Fayc1v9_1),.clk(gclk));
	jdff dff_A_pbft6EN75_1(.dout(w_n719_0[1]),.din(w_dff_A_pbft6EN75_1),.clk(gclk));
	jdff dff_A_v9ao2i6o1_1(.dout(w_dff_A_pbft6EN75_1),.din(w_dff_A_v9ao2i6o1_1),.clk(gclk));
	jdff dff_A_uqg8fGWl4_1(.dout(w_dff_A_v9ao2i6o1_1),.din(w_dff_A_uqg8fGWl4_1),.clk(gclk));
	jdff dff_A_XfTKPgdB9_1(.dout(w_dff_A_uqg8fGWl4_1),.din(w_dff_A_XfTKPgdB9_1),.clk(gclk));
	jdff dff_A_1awB07r12_1(.dout(w_dff_A_XfTKPgdB9_1),.din(w_dff_A_1awB07r12_1),.clk(gclk));
	jdff dff_B_57G6NsdX4_0(.din(n616),.dout(w_dff_B_57G6NsdX4_0),.clk(gclk));
	jdff dff_A_R1RIDmXh3_1(.dout(w_G331_0[1]),.din(w_dff_A_R1RIDmXh3_1),.clk(gclk));
	jdff dff_A_F8Uk3U9y7_1(.dout(w_G324_1[1]),.din(w_dff_A_F8Uk3U9y7_1),.clk(gclk));
	jdff dff_A_zFfp6bVg0_2(.dout(w_G324_0[2]),.din(w_dff_A_zFfp6bVg0_2),.clk(gclk));
	jdff dff_A_VICh85vW4_0(.dout(w_G503_0[0]),.din(w_dff_A_VICh85vW4_0),.clk(gclk));
	jdff dff_A_R6CvotoX6_0(.dout(w_dff_A_VICh85vW4_0),.din(w_dff_A_R6CvotoX6_0),.clk(gclk));
	jdff dff_A_jKyAwvkP8_0(.dout(w_dff_A_R6CvotoX6_0),.din(w_dff_A_jKyAwvkP8_0),.clk(gclk));
	jdff dff_A_GN83aTc42_0(.dout(w_dff_A_jKyAwvkP8_0),.din(w_dff_A_GN83aTc42_0),.clk(gclk));
	jdff dff_A_10AtPci18_2(.dout(w_G503_0[2]),.din(w_dff_A_10AtPci18_2),.clk(gclk));
	jdff dff_A_NJpbWQ6H2_2(.dout(w_dff_A_10AtPci18_2),.din(w_dff_A_NJpbWQ6H2_2),.clk(gclk));
	jdff dff_A_EIhQxOxi1_0(.dout(w_G4092_4[0]),.din(w_dff_A_EIhQxOxi1_0),.clk(gclk));
	jdff dff_A_qJsf05Up1_0(.dout(w_dff_A_EIhQxOxi1_0),.din(w_dff_A_qJsf05Up1_0),.clk(gclk));
	jdff dff_A_wYSDX8fS2_0(.dout(w_dff_A_qJsf05Up1_0),.din(w_dff_A_wYSDX8fS2_0),.clk(gclk));
	jdff dff_A_VOUIoQCP5_0(.dout(w_dff_A_wYSDX8fS2_0),.din(w_dff_A_VOUIoQCP5_0),.clk(gclk));
	jdff dff_A_TAJot7FE7_0(.dout(w_dff_A_VOUIoQCP5_0),.din(w_dff_A_TAJot7FE7_0),.clk(gclk));
	jdff dff_A_uISgwoQ22_0(.dout(w_dff_A_TAJot7FE7_0),.din(w_dff_A_uISgwoQ22_0),.clk(gclk));
	jdff dff_A_oTkjMKGO6_0(.dout(w_dff_A_uISgwoQ22_0),.din(w_dff_A_oTkjMKGO6_0),.clk(gclk));
	jdff dff_A_9LdN4vs39_0(.dout(w_dff_A_oTkjMKGO6_0),.din(w_dff_A_9LdN4vs39_0),.clk(gclk));
	jdff dff_A_kh43U5pn6_0(.dout(w_dff_A_9LdN4vs39_0),.din(w_dff_A_kh43U5pn6_0),.clk(gclk));
	jdff dff_A_4bJdu3ei3_0(.dout(w_dff_A_kh43U5pn6_0),.din(w_dff_A_4bJdu3ei3_0),.clk(gclk));
	jdff dff_A_UvAzVEjK0_0(.dout(w_dff_A_4bJdu3ei3_0),.din(w_dff_A_UvAzVEjK0_0),.clk(gclk));
	jdff dff_A_djvkdCPF3_0(.dout(w_dff_A_UvAzVEjK0_0),.din(w_dff_A_djvkdCPF3_0),.clk(gclk));
	jdff dff_A_ArpKi3J15_0(.dout(w_dff_A_djvkdCPF3_0),.din(w_dff_A_ArpKi3J15_0),.clk(gclk));
	jdff dff_A_opWE1Xsm3_0(.dout(w_dff_A_ArpKi3J15_0),.din(w_dff_A_opWE1Xsm3_0),.clk(gclk));
	jdff dff_A_5H3EhhXK2_0(.dout(w_G4092_1[0]),.din(w_dff_A_5H3EhhXK2_0),.clk(gclk));
	jdff dff_A_AwplXlA05_0(.dout(w_dff_A_5H3EhhXK2_0),.din(w_dff_A_AwplXlA05_0),.clk(gclk));
	jdff dff_A_SvU9OCQG5_0(.dout(w_dff_A_AwplXlA05_0),.din(w_dff_A_SvU9OCQG5_0),.clk(gclk));
	jdff dff_A_PfGgEJzT3_0(.dout(w_dff_A_SvU9OCQG5_0),.din(w_dff_A_PfGgEJzT3_0),.clk(gclk));
	jdff dff_A_r73D5zJI9_0(.dout(w_dff_A_PfGgEJzT3_0),.din(w_dff_A_r73D5zJI9_0),.clk(gclk));
	jdff dff_A_xXFR20xn1_0(.dout(w_dff_A_r73D5zJI9_0),.din(w_dff_A_xXFR20xn1_0),.clk(gclk));
	jdff dff_A_kn2ty5aY0_2(.dout(w_G4092_1[2]),.din(w_dff_A_kn2ty5aY0_2),.clk(gclk));
	jdff dff_A_4QZMshbv7_2(.dout(w_dff_A_kn2ty5aY0_2),.din(w_dff_A_4QZMshbv7_2),.clk(gclk));
	jdff dff_A_0DjVm3660_2(.dout(w_dff_A_4QZMshbv7_2),.din(w_dff_A_0DjVm3660_2),.clk(gclk));
	jdff dff_A_8AaK8aOG1_2(.dout(w_dff_A_0DjVm3660_2),.din(w_dff_A_8AaK8aOG1_2),.clk(gclk));
	jdff dff_B_OQgniS8Z0_0(.din(n1673),.dout(w_dff_B_OQgniS8Z0_0),.clk(gclk));
	jdff dff_B_c7wDodW81_0(.din(w_dff_B_OQgniS8Z0_0),.dout(w_dff_B_c7wDodW81_0),.clk(gclk));
	jdff dff_B_dxlYHcWx4_0(.din(w_dff_B_c7wDodW81_0),.dout(w_dff_B_dxlYHcWx4_0),.clk(gclk));
	jdff dff_B_Ukh7m1Bv2_0(.din(w_dff_B_dxlYHcWx4_0),.dout(w_dff_B_Ukh7m1Bv2_0),.clk(gclk));
	jdff dff_B_7QClgarR9_0(.din(w_dff_B_Ukh7m1Bv2_0),.dout(w_dff_B_7QClgarR9_0),.clk(gclk));
	jdff dff_B_H1gZ39aE4_0(.din(w_dff_B_7QClgarR9_0),.dout(w_dff_B_H1gZ39aE4_0),.clk(gclk));
	jdff dff_B_d2uBp8jE2_0(.din(w_dff_B_H1gZ39aE4_0),.dout(w_dff_B_d2uBp8jE2_0),.clk(gclk));
	jdff dff_B_5OCG9Rsg8_0(.din(w_dff_B_d2uBp8jE2_0),.dout(w_dff_B_5OCG9Rsg8_0),.clk(gclk));
	jdff dff_B_9qu58Pm82_0(.din(w_dff_B_5OCG9Rsg8_0),.dout(w_dff_B_9qu58Pm82_0),.clk(gclk));
	jdff dff_B_qKqzwTI43_0(.din(w_dff_B_9qu58Pm82_0),.dout(w_dff_B_qKqzwTI43_0),.clk(gclk));
	jdff dff_B_FNlDNXDC1_0(.din(w_dff_B_qKqzwTI43_0),.dout(w_dff_B_FNlDNXDC1_0),.clk(gclk));
	jdff dff_B_RH52Fyov0_0(.din(w_dff_B_FNlDNXDC1_0),.dout(w_dff_B_RH52Fyov0_0),.clk(gclk));
	jdff dff_B_iQyb6XoS3_0(.din(w_dff_B_RH52Fyov0_0),.dout(w_dff_B_iQyb6XoS3_0),.clk(gclk));
	jdff dff_B_SkypU4MT0_0(.din(w_dff_B_iQyb6XoS3_0),.dout(w_dff_B_SkypU4MT0_0),.clk(gclk));
	jdff dff_B_L8xjIghs4_0(.din(w_dff_B_SkypU4MT0_0),.dout(w_dff_B_L8xjIghs4_0),.clk(gclk));
	jdff dff_B_OnK7SI3H5_0(.din(w_dff_B_L8xjIghs4_0),.dout(w_dff_B_OnK7SI3H5_0),.clk(gclk));
	jdff dff_B_WPf0bgdS4_0(.din(w_dff_B_OnK7SI3H5_0),.dout(w_dff_B_WPf0bgdS4_0),.clk(gclk));
	jdff dff_B_8UmPLGEf0_0(.din(w_dff_B_WPf0bgdS4_0),.dout(w_dff_B_8UmPLGEf0_0),.clk(gclk));
	jdff dff_B_UAoLTV0I0_0(.din(w_dff_B_8UmPLGEf0_0),.dout(w_dff_B_UAoLTV0I0_0),.clk(gclk));
	jdff dff_B_FRDYFa6S5_1(.din(n1588),.dout(w_dff_B_FRDYFa6S5_1),.clk(gclk));
	jdff dff_B_vce812uo3_1(.din(w_dff_B_FRDYFa6S5_1),.dout(w_dff_B_vce812uo3_1),.clk(gclk));
	jdff dff_B_qfHGV0D74_1(.din(w_dff_B_vce812uo3_1),.dout(w_dff_B_qfHGV0D74_1),.clk(gclk));
	jdff dff_B_efRlcB7r5_1(.din(w_dff_B_qfHGV0D74_1),.dout(w_dff_B_efRlcB7r5_1),.clk(gclk));
	jdff dff_B_LEQP3c7v9_1(.din(w_dff_B_efRlcB7r5_1),.dout(w_dff_B_LEQP3c7v9_1),.clk(gclk));
	jdff dff_B_7dmBLewq7_1(.din(w_dff_B_LEQP3c7v9_1),.dout(w_dff_B_7dmBLewq7_1),.clk(gclk));
	jdff dff_B_t6fAe9au6_1(.din(w_dff_B_7dmBLewq7_1),.dout(w_dff_B_t6fAe9au6_1),.clk(gclk));
	jdff dff_B_1X3yTzcg9_1(.din(w_dff_B_t6fAe9au6_1),.dout(w_dff_B_1X3yTzcg9_1),.clk(gclk));
	jdff dff_B_6iQyRD5L9_1(.din(n1655),.dout(w_dff_B_6iQyRD5L9_1),.clk(gclk));
	jdff dff_B_Nb21UJTq6_1(.din(w_dff_B_6iQyRD5L9_1),.dout(w_dff_B_Nb21UJTq6_1),.clk(gclk));
	jdff dff_A_xlkFGP9J9_2(.dout(w_n588_0[2]),.din(w_dff_A_xlkFGP9J9_2),.clk(gclk));
	jdff dff_A_4SjY06lH7_2(.dout(w_dff_A_xlkFGP9J9_2),.din(w_dff_A_4SjY06lH7_2),.clk(gclk));
	jdff dff_A_L7QMeyn52_1(.dout(w_n1652_0[1]),.din(w_dff_A_L7QMeyn52_1),.clk(gclk));
	jdff dff_B_QoTvP5CI6_0(.din(n1649),.dout(w_dff_B_QoTvP5CI6_0),.clk(gclk));
	jdff dff_B_kEmmUmCN9_1(.din(n1645),.dout(w_dff_B_kEmmUmCN9_1),.clk(gclk));
	jdff dff_B_U1nnP5rN5_1(.din(w_dff_B_kEmmUmCN9_1),.dout(w_dff_B_U1nnP5rN5_1),.clk(gclk));
	jdff dff_B_WBi1Vhx51_1(.din(w_dff_B_U1nnP5rN5_1),.dout(w_dff_B_WBi1Vhx51_1),.clk(gclk));
	jdff dff_B_8IX8KGr32_1(.din(w_dff_B_WBi1Vhx51_1),.dout(w_dff_B_8IX8KGr32_1),.clk(gclk));
	jdff dff_B_8cdrglPg3_1(.din(w_dff_B_8IX8KGr32_1),.dout(w_dff_B_8cdrglPg3_1),.clk(gclk));
	jdff dff_B_keaKlAXc1_1(.din(n1638),.dout(w_dff_B_keaKlAXc1_1),.clk(gclk));
	jdff dff_B_KfVMJ9oW4_1(.din(w_dff_B_keaKlAXc1_1),.dout(w_dff_B_KfVMJ9oW4_1),.clk(gclk));
	jdff dff_B_u1f4EHL35_0(.din(n1641),.dout(w_dff_B_u1f4EHL35_0),.clk(gclk));
	jdff dff_B_T8eDJLQt1_0(.din(n1640),.dout(w_dff_B_T8eDJLQt1_0),.clk(gclk));
	jdff dff_A_Uws9P4kF7_1(.dout(w_n609_0[1]),.din(w_dff_A_Uws9P4kF7_1),.clk(gclk));
	jdff dff_A_3trX53hq8_1(.dout(w_dff_A_Uws9P4kF7_1),.din(w_dff_A_3trX53hq8_1),.clk(gclk));
	jdff dff_A_QtIGU6nu1_1(.dout(w_dff_A_3trX53hq8_1),.din(w_dff_A_QtIGU6nu1_1),.clk(gclk));
	jdff dff_A_FyMgIb5q1_1(.dout(w_dff_A_QtIGU6nu1_1),.din(w_dff_A_FyMgIb5q1_1),.clk(gclk));
	jdff dff_A_oMSGCTfm4_1(.dout(w_dff_A_FyMgIb5q1_1),.din(w_dff_A_oMSGCTfm4_1),.clk(gclk));
	jdff dff_A_1f2BLEyN8_1(.dout(w_dff_A_oMSGCTfm4_1),.din(w_dff_A_1f2BLEyN8_1),.clk(gclk));
	jdff dff_A_1UZuqTSm6_1(.dout(w_dff_A_1f2BLEyN8_1),.din(w_dff_A_1UZuqTSm6_1),.clk(gclk));
	jdff dff_A_rUws5IQk5_1(.dout(w_n962_0[1]),.din(w_dff_A_rUws5IQk5_1),.clk(gclk));
	jdff dff_A_vvzJet7l9_1(.dout(w_dff_A_rUws5IQk5_1),.din(w_dff_A_vvzJet7l9_1),.clk(gclk));
	jdff dff_A_bID7jaFa3_1(.dout(w_dff_A_vvzJet7l9_1),.din(w_dff_A_bID7jaFa3_1),.clk(gclk));
	jdff dff_A_MTSappig0_1(.dout(w_dff_A_bID7jaFa3_1),.din(w_dff_A_MTSappig0_1),.clk(gclk));
	jdff dff_A_5r6h0yxY4_1(.dout(w_dff_A_MTSappig0_1),.din(w_dff_A_5r6h0yxY4_1),.clk(gclk));
	jdff dff_A_qKtk3BAZ0_1(.dout(w_dff_A_5r6h0yxY4_1),.din(w_dff_A_qKtk3BAZ0_1),.clk(gclk));
	jdff dff_B_06dA8gXU0_2(.din(n962),.dout(w_dff_B_06dA8gXU0_2),.clk(gclk));
	jdff dff_A_moXGfcut3_2(.dout(w_n938_0[2]),.din(w_dff_A_moXGfcut3_2),.clk(gclk));
	jdff dff_A_kxwH2KKG7_2(.dout(w_dff_A_moXGfcut3_2),.din(w_dff_A_kxwH2KKG7_2),.clk(gclk));
	jdff dff_A_4VevNxZE6_2(.dout(w_dff_A_kxwH2KKG7_2),.din(w_dff_A_4VevNxZE6_2),.clk(gclk));
	jdff dff_A_MBniGXJD5_2(.dout(w_dff_A_4VevNxZE6_2),.din(w_dff_A_MBniGXJD5_2),.clk(gclk));
	jdff dff_A_GBmzx6wz4_2(.dout(w_dff_A_MBniGXJD5_2),.din(w_dff_A_GBmzx6wz4_2),.clk(gclk));
	jdff dff_B_z6k5rTOH2_1(.din(n707),.dout(w_dff_B_z6k5rTOH2_1),.clk(gclk));
	jdff dff_B_cvGlQ0044_1(.din(w_dff_B_z6k5rTOH2_1),.dout(w_dff_B_cvGlQ0044_1),.clk(gclk));
	jdff dff_B_bsMZhnDY2_1(.din(w_dff_B_cvGlQ0044_1),.dout(w_dff_B_bsMZhnDY2_1),.clk(gclk));
	jdff dff_B_ttpy0CZW9_1(.din(n708),.dout(w_dff_B_ttpy0CZW9_1),.clk(gclk));
	jdff dff_B_3VKKs2DS2_1(.din(w_dff_B_ttpy0CZW9_1),.dout(w_dff_B_3VKKs2DS2_1),.clk(gclk));
	jdff dff_A_fZQ7cme07_1(.dout(w_n713_0[1]),.din(w_dff_A_fZQ7cme07_1),.clk(gclk));
	jdff dff_A_Aco4Rfxw7_1(.dout(w_dff_A_fZQ7cme07_1),.din(w_dff_A_Aco4Rfxw7_1),.clk(gclk));
	jdff dff_A_EUgEOsnn9_1(.dout(w_dff_A_Aco4Rfxw7_1),.din(w_dff_A_EUgEOsnn9_1),.clk(gclk));
	jdff dff_A_khJRHsrT5_1(.dout(w_dff_A_EUgEOsnn9_1),.din(w_dff_A_khJRHsrT5_1),.clk(gclk));
	jdff dff_A_OY7Q8sWP2_1(.dout(w_dff_A_khJRHsrT5_1),.din(w_dff_A_OY7Q8sWP2_1),.clk(gclk));
	jdff dff_A_9aUQXAKb9_1(.dout(w_dff_A_OY7Q8sWP2_1),.din(w_dff_A_9aUQXAKb9_1),.clk(gclk));
	jdff dff_A_srQ6aHx94_1(.dout(w_dff_A_9aUQXAKb9_1),.din(w_dff_A_srQ6aHx94_1),.clk(gclk));
	jdff dff_A_mi9eGh4F5_0(.dout(w_n710_0[0]),.din(w_dff_A_mi9eGh4F5_0),.clk(gclk));
	jdff dff_A_rLAMROX73_0(.dout(w_dff_A_mi9eGh4F5_0),.din(w_dff_A_rLAMROX73_0),.clk(gclk));
	jdff dff_A_enGQamJO4_0(.dout(w_dff_A_rLAMROX73_0),.din(w_dff_A_enGQamJO4_0),.clk(gclk));
	jdff dff_A_62LuOKr94_0(.dout(w_dff_A_enGQamJO4_0),.din(w_dff_A_62LuOKr94_0),.clk(gclk));
	jdff dff_A_ji7Ssb0i9_0(.dout(w_dff_A_62LuOKr94_0),.din(w_dff_A_ji7Ssb0i9_0),.clk(gclk));
	jdff dff_A_FHuImOqd3_0(.dout(w_dff_A_ji7Ssb0i9_0),.din(w_dff_A_FHuImOqd3_0),.clk(gclk));
	jdff dff_A_8VYSaQLh2_0(.dout(w_dff_A_FHuImOqd3_0),.din(w_dff_A_8VYSaQLh2_0),.clk(gclk));
	jdff dff_A_F7FvTbIU6_0(.dout(w_dff_A_8VYSaQLh2_0),.din(w_dff_A_F7FvTbIU6_0),.clk(gclk));
	jdff dff_A_xXu241s53_0(.dout(w_n597_0[0]),.din(w_dff_A_xXu241s53_0),.clk(gclk));
	jdff dff_A_GPjp26wa3_0(.dout(w_dff_A_xXu241s53_0),.din(w_dff_A_GPjp26wa3_0),.clk(gclk));
	jdff dff_A_mqHihzL63_0(.dout(w_dff_A_GPjp26wa3_0),.din(w_dff_A_mqHihzL63_0),.clk(gclk));
	jdff dff_A_Dp3jRNxF2_0(.dout(w_dff_A_mqHihzL63_0),.din(w_dff_A_Dp3jRNxF2_0),.clk(gclk));
	jdff dff_A_1T9U05Yz1_0(.dout(w_dff_A_Dp3jRNxF2_0),.din(w_dff_A_1T9U05Yz1_0),.clk(gclk));
	jdff dff_A_dpYbe0Vd4_0(.dout(w_n496_1[0]),.din(w_dff_A_dpYbe0Vd4_0),.clk(gclk));
	jdff dff_A_JOATgsfg6_0(.dout(w_dff_A_dpYbe0Vd4_0),.din(w_dff_A_JOATgsfg6_0),.clk(gclk));
	jdff dff_A_37apWN0E4_0(.dout(w_n1637_0[0]),.din(w_dff_A_37apWN0E4_0),.clk(gclk));
	jdff dff_A_LEtQZjGE5_0(.dout(w_dff_A_37apWN0E4_0),.din(w_dff_A_LEtQZjGE5_0),.clk(gclk));
	jdff dff_B_cPd2n3vn8_2(.din(n1637),.dout(w_dff_B_cPd2n3vn8_2),.clk(gclk));
	jdff dff_B_pJnT534a4_2(.din(w_dff_B_cPd2n3vn8_2),.dout(w_dff_B_pJnT534a4_2),.clk(gclk));
	jdff dff_A_mirKFcdb1_1(.dout(w_n608_0[1]),.din(w_dff_A_mirKFcdb1_1),.clk(gclk));
	jdff dff_A_8b2e4GZU0_1(.dout(w_dff_A_mirKFcdb1_1),.din(w_dff_A_8b2e4GZU0_1),.clk(gclk));
	jdff dff_A_1dhyPwgU6_1(.dout(w_dff_A_8b2e4GZU0_1),.din(w_dff_A_1dhyPwgU6_1),.clk(gclk));
	jdff dff_A_xHW8LyAM9_1(.dout(w_dff_A_1dhyPwgU6_1),.din(w_dff_A_xHW8LyAM9_1),.clk(gclk));
	jdff dff_A_Wjj189Lq3_1(.dout(w_dff_A_xHW8LyAM9_1),.din(w_dff_A_Wjj189Lq3_1),.clk(gclk));
	jdff dff_A_qGF3hIIh8_1(.dout(w_dff_A_Wjj189Lq3_1),.din(w_dff_A_qGF3hIIh8_1),.clk(gclk));
	jdff dff_A_oNpKmeNu2_1(.dout(w_dff_A_qGF3hIIh8_1),.din(w_dff_A_oNpKmeNu2_1),.clk(gclk));
	jdff dff_A_L83vThpW0_1(.dout(w_dff_A_oNpKmeNu2_1),.din(w_dff_A_L83vThpW0_1),.clk(gclk));
	jdff dff_A_PhQ3LTox0_1(.dout(w_dff_A_L83vThpW0_1),.din(w_dff_A_PhQ3LTox0_1),.clk(gclk));
	jdff dff_A_enWkxjoB9_1(.dout(w_dff_A_PhQ3LTox0_1),.din(w_dff_A_enWkxjoB9_1),.clk(gclk));
	jdff dff_A_EMhCsHJR1_2(.dout(w_n608_0[2]),.din(w_dff_A_EMhCsHJR1_2),.clk(gclk));
	jdff dff_B_EXzRqPhv9_0(.din(n606),.dout(w_dff_B_EXzRqPhv9_0),.clk(gclk));
	jdff dff_B_vbotFnb24_1(.din(G217),.dout(w_dff_B_vbotFnb24_1),.clk(gclk));
	jdff dff_A_Rr5OZwbN8_0(.dout(w_n592_0[0]),.din(w_dff_A_Rr5OZwbN8_0),.clk(gclk));
	jdff dff_A_4x3qatY19_2(.dout(w_n592_0[2]),.din(w_dff_A_4x3qatY19_2),.clk(gclk));
	jdff dff_A_8mxpvWCz0_2(.dout(w_dff_A_4x3qatY19_2),.din(w_dff_A_8mxpvWCz0_2),.clk(gclk));
	jdff dff_A_Yv6kDql04_2(.dout(w_dff_A_8mxpvWCz0_2),.din(w_dff_A_Yv6kDql04_2),.clk(gclk));
	jdff dff_A_ib9Rh1lq1_2(.dout(w_dff_A_Yv6kDql04_2),.din(w_dff_A_ib9Rh1lq1_2),.clk(gclk));
	jdff dff_B_qtKr0fpF5_1(.din(n589),.dout(w_dff_B_qtKr0fpF5_1),.clk(gclk));
	jdff dff_B_O0nRUcvV3_1(.din(G209),.dout(w_dff_B_O0nRUcvV3_1),.clk(gclk));
	jdff dff_A_fpZxkH2L2_0(.dout(w_n602_0[0]),.din(w_dff_A_fpZxkH2L2_0),.clk(gclk));
	jdff dff_A_BmdpZ4Lh4_0(.dout(w_n711_0[0]),.din(w_dff_A_BmdpZ4Lh4_0),.clk(gclk));
	jdff dff_A_4cNbMmsO6_0(.dout(w_dff_A_BmdpZ4Lh4_0),.din(w_dff_A_4cNbMmsO6_0),.clk(gclk));
	jdff dff_A_r3NdDLcl6_2(.dout(w_n954_0[2]),.din(w_dff_A_r3NdDLcl6_2),.clk(gclk));
	jdff dff_A_mLhvBfUC2_2(.dout(w_dff_A_r3NdDLcl6_2),.din(w_dff_A_mLhvBfUC2_2),.clk(gclk));
	jdff dff_A_weVSCX4f8_2(.dout(w_dff_A_mLhvBfUC2_2),.din(w_dff_A_weVSCX4f8_2),.clk(gclk));
	jdff dff_A_g4AstPkX1_2(.dout(w_dff_A_weVSCX4f8_2),.din(w_dff_A_g4AstPkX1_2),.clk(gclk));
	jdff dff_A_cRaF1Mbl7_2(.dout(w_dff_A_g4AstPkX1_2),.din(w_dff_A_cRaF1Mbl7_2),.clk(gclk));
	jdff dff_A_G6qPK8wB9_2(.dout(w_dff_A_cRaF1Mbl7_2),.din(w_dff_A_G6qPK8wB9_2),.clk(gclk));
	jdff dff_A_xgc5JR2D4_2(.dout(w_dff_A_G6qPK8wB9_2),.din(w_dff_A_xgc5JR2D4_2),.clk(gclk));
	jdff dff_B_K5Phutoi0_2(.din(n1633),.dout(w_dff_B_K5Phutoi0_2),.clk(gclk));
	jdff dff_A_7Weigvoq1_1(.dout(w_n709_0[1]),.din(w_dff_A_7Weigvoq1_1),.clk(gclk));
	jdff dff_B_G1yOpguQ2_0(.din(n600),.dout(w_dff_B_G1yOpguQ2_0),.clk(gclk));
	jdff dff_B_y63hCaOL7_1(.din(G225),.dout(w_dff_B_y63hCaOL7_1),.clk(gclk));
	jdff dff_B_Yd1FmHXW5_0(.din(n595),.dout(w_dff_B_Yd1FmHXW5_0),.clk(gclk));
	jdff dff_B_8f4RVvMu5_1(.din(G233),.dout(w_dff_B_8f4RVvMu5_1),.clk(gclk));
	jdff dff_A_VySiNYam7_1(.dout(w_n703_0[1]),.din(w_dff_A_VySiNYam7_1),.clk(gclk));
	jdff dff_A_BLVgBP3s8_0(.dout(w_n685_0[0]),.din(w_dff_A_BLVgBP3s8_0),.clk(gclk));
	jdff dff_A_KaP3mLZ20_0(.dout(w_dff_A_BLVgBP3s8_0),.din(w_dff_A_KaP3mLZ20_0),.clk(gclk));
	jdff dff_B_8quRQZr08_2(.din(n685),.dout(w_dff_B_8quRQZr08_2),.clk(gclk));
	jdff dff_B_PGJ73wt72_2(.din(w_dff_B_8quRQZr08_2),.dout(w_dff_B_PGJ73wt72_2),.clk(gclk));
	jdff dff_B_i8QFpFER7_2(.din(w_dff_B_PGJ73wt72_2),.dout(w_dff_B_i8QFpFER7_2),.clk(gclk));
	jdff dff_A_hyklK2l55_0(.dout(w_n684_0[0]),.din(w_dff_A_hyklK2l55_0),.clk(gclk));
	jdff dff_A_B2v12AOc4_0(.dout(w_dff_A_hyklK2l55_0),.din(w_dff_A_B2v12AOc4_0),.clk(gclk));
	jdff dff_A_HKTgWa7w6_0(.dout(w_dff_A_B2v12AOc4_0),.din(w_dff_A_HKTgWa7w6_0),.clk(gclk));
	jdff dff_A_Awaqc4aS2_0(.dout(w_dff_A_HKTgWa7w6_0),.din(w_dff_A_Awaqc4aS2_0),.clk(gclk));
	jdff dff_A_2QmQ8UmM1_1(.dout(w_n682_0[1]),.din(w_dff_A_2QmQ8UmM1_1),.clk(gclk));
	jdff dff_A_0VGBal8i6_1(.dout(w_dff_A_2QmQ8UmM1_1),.din(w_dff_A_0VGBal8i6_1),.clk(gclk));
	jdff dff_A_WHOrqpLf1_1(.dout(w_dff_A_0VGBal8i6_1),.din(w_dff_A_WHOrqpLf1_1),.clk(gclk));
	jdff dff_A_mp2OLete7_1(.dout(w_dff_A_WHOrqpLf1_1),.din(w_dff_A_mp2OLete7_1),.clk(gclk));
	jdff dff_A_RIzCUENo3_1(.dout(w_dff_A_mp2OLete7_1),.din(w_dff_A_RIzCUENo3_1),.clk(gclk));
	jdff dff_A_Xw0QZFdE1_1(.dout(w_dff_A_RIzCUENo3_1),.din(w_dff_A_Xw0QZFdE1_1),.clk(gclk));
	jdff dff_A_MXSlLSCG9_2(.dout(w_n682_0[2]),.din(w_dff_A_MXSlLSCG9_2),.clk(gclk));
	jdff dff_A_UexTmkzh5_2(.dout(w_dff_A_MXSlLSCG9_2),.din(w_dff_A_UexTmkzh5_2),.clk(gclk));
	jdff dff_A_2JeTvPl28_2(.dout(w_dff_A_UexTmkzh5_2),.din(w_dff_A_2JeTvPl28_2),.clk(gclk));
	jdff dff_A_obhZ1qgF7_2(.dout(w_dff_A_2JeTvPl28_2),.din(w_dff_A_obhZ1qgF7_2),.clk(gclk));
	jdff dff_A_9OxIGf3C9_2(.dout(w_dff_A_obhZ1qgF7_2),.din(w_dff_A_9OxIGf3C9_2),.clk(gclk));
	jdff dff_A_NxH4tdPn0_2(.dout(w_dff_A_9OxIGf3C9_2),.din(w_dff_A_NxH4tdPn0_2),.clk(gclk));
	jdff dff_B_kghlOlOs9_0(.din(n1630),.dout(w_dff_B_kghlOlOs9_0),.clk(gclk));
	jdff dff_B_h6UqhT4u7_0(.din(w_dff_B_kghlOlOs9_0),.dout(w_dff_B_h6UqhT4u7_0),.clk(gclk));
	jdff dff_B_ZRUgqySz6_0(.din(w_dff_B_h6UqhT4u7_0),.dout(w_dff_B_ZRUgqySz6_0),.clk(gclk));
	jdff dff_B_cgW0hOZr8_0(.din(w_dff_B_ZRUgqySz6_0),.dout(w_dff_B_cgW0hOZr8_0),.clk(gclk));
	jdff dff_B_wcYJ1TzN1_0(.din(w_dff_B_cgW0hOZr8_0),.dout(w_dff_B_wcYJ1TzN1_0),.clk(gclk));
	jdff dff_B_BrCnk7Kw2_0(.din(w_dff_B_wcYJ1TzN1_0),.dout(w_dff_B_BrCnk7Kw2_0),.clk(gclk));
	jdff dff_B_SmgpBJxx1_0(.din(w_dff_B_BrCnk7Kw2_0),.dout(w_dff_B_SmgpBJxx1_0),.clk(gclk));
	jdff dff_B_jFPfXCOu8_0(.din(w_dff_B_SmgpBJxx1_0),.dout(w_dff_B_jFPfXCOu8_0),.clk(gclk));
	jdff dff_B_kmufscFm5_0(.din(w_dff_B_jFPfXCOu8_0),.dout(w_dff_B_kmufscFm5_0),.clk(gclk));
	jdff dff_B_2j0nYXVw6_0(.din(n1628),.dout(w_dff_B_2j0nYXVw6_0),.clk(gclk));
	jdff dff_B_6bkGyK2w7_0(.din(w_dff_B_2j0nYXVw6_0),.dout(w_dff_B_6bkGyK2w7_0),.clk(gclk));
	jdff dff_B_NmUcLTXn0_1(.din(n1625),.dout(w_dff_B_NmUcLTXn0_1),.clk(gclk));
	jdff dff_B_8COAyz5T1_1(.din(n1623),.dout(w_dff_B_8COAyz5T1_1),.clk(gclk));
	jdff dff_B_4grUwu5F0_1(.din(w_dff_B_8COAyz5T1_1),.dout(w_dff_B_4grUwu5F0_1),.clk(gclk));
	jdff dff_A_NxE5199g4_0(.dout(w_n1618_0[0]),.din(w_dff_A_NxE5199g4_0),.clk(gclk));
	jdff dff_A_c1571MWv0_0(.dout(w_dff_A_NxE5199g4_0),.din(w_dff_A_c1571MWv0_0),.clk(gclk));
	jdff dff_B_1UAZNobP5_2(.din(n1618),.dout(w_dff_B_1UAZNobP5_2),.clk(gclk));
	jdff dff_B_VNHm9cY24_2(.din(w_dff_B_1UAZNobP5_2),.dout(w_dff_B_VNHm9cY24_2),.clk(gclk));
	jdff dff_B_918j1l7K2_2(.din(w_dff_B_VNHm9cY24_2),.dout(w_dff_B_918j1l7K2_2),.clk(gclk));
	jdff dff_B_VjbN95og9_2(.din(w_dff_B_918j1l7K2_2),.dout(w_dff_B_VjbN95og9_2),.clk(gclk));
	jdff dff_B_fivtRROq9_2(.din(w_dff_B_VjbN95og9_2),.dout(w_dff_B_fivtRROq9_2),.clk(gclk));
	jdff dff_B_ux2iu24m6_2(.din(w_dff_B_fivtRROq9_2),.dout(w_dff_B_ux2iu24m6_2),.clk(gclk));
	jdff dff_B_6ape9e1y0_2(.din(w_dff_B_ux2iu24m6_2),.dout(w_dff_B_6ape9e1y0_2),.clk(gclk));
	jdff dff_B_7HdnSMWM1_2(.din(w_dff_B_6ape9e1y0_2),.dout(w_dff_B_7HdnSMWM1_2),.clk(gclk));
	jdff dff_B_TWfjzTAo4_2(.din(w_dff_B_7HdnSMWM1_2),.dout(w_dff_B_TWfjzTAo4_2),.clk(gclk));
	jdff dff_B_3apDr30h5_2(.din(w_dff_B_TWfjzTAo4_2),.dout(w_dff_B_3apDr30h5_2),.clk(gclk));
	jdff dff_B_Ujo9Syr77_2(.din(w_dff_B_3apDr30h5_2),.dout(w_dff_B_Ujo9Syr77_2),.clk(gclk));
	jdff dff_B_fCBI0eF75_2(.din(w_dff_B_Ujo9Syr77_2),.dout(w_dff_B_fCBI0eF75_2),.clk(gclk));
	jdff dff_A_Kyha9QU23_0(.dout(w_G1497_0[0]),.din(w_dff_A_Kyha9QU23_0),.clk(gclk));
	jdff dff_A_LpLLVyIt7_0(.dout(w_dff_A_Kyha9QU23_0),.din(w_dff_A_LpLLVyIt7_0),.clk(gclk));
	jdff dff_A_b8Zi22nb3_0(.dout(w_dff_A_LpLLVyIt7_0),.din(w_dff_A_b8Zi22nb3_0),.clk(gclk));
	jdff dff_A_G8jV60gn7_0(.dout(w_dff_A_b8Zi22nb3_0),.din(w_dff_A_G8jV60gn7_0),.clk(gclk));
	jdff dff_A_gv9hIwzM5_0(.dout(w_dff_A_G8jV60gn7_0),.din(w_dff_A_gv9hIwzM5_0),.clk(gclk));
	jdff dff_A_efNm6fAq4_0(.dout(w_dff_A_gv9hIwzM5_0),.din(w_dff_A_efNm6fAq4_0),.clk(gclk));
	jdff dff_A_7lweI8Tw5_0(.dout(w_dff_A_efNm6fAq4_0),.din(w_dff_A_7lweI8Tw5_0),.clk(gclk));
	jdff dff_A_MwC5JsDB6_0(.dout(w_dff_A_7lweI8Tw5_0),.din(w_dff_A_MwC5JsDB6_0),.clk(gclk));
	jdff dff_A_WqcEn3r81_0(.dout(w_dff_A_MwC5JsDB6_0),.din(w_dff_A_WqcEn3r81_0),.clk(gclk));
	jdff dff_A_XuDmv30e4_0(.dout(w_dff_A_WqcEn3r81_0),.din(w_dff_A_XuDmv30e4_0),.clk(gclk));
	jdff dff_A_AccpODWJ0_0(.dout(w_dff_A_XuDmv30e4_0),.din(w_dff_A_AccpODWJ0_0),.clk(gclk));
	jdff dff_A_MVkNx5Pp9_0(.dout(w_dff_A_AccpODWJ0_0),.din(w_dff_A_MVkNx5Pp9_0),.clk(gclk));
	jdff dff_A_2UiPeyF29_0(.dout(w_dff_A_MVkNx5Pp9_0),.din(w_dff_A_2UiPeyF29_0),.clk(gclk));
	jdff dff_A_nSdn0rlr3_0(.dout(w_dff_A_2UiPeyF29_0),.din(w_dff_A_nSdn0rlr3_0),.clk(gclk));
	jdff dff_A_USsYQNdK9_0(.dout(w_dff_A_nSdn0rlr3_0),.din(w_dff_A_USsYQNdK9_0),.clk(gclk));
	jdff dff_A_4ouY8qtj9_1(.dout(w_G1497_0[1]),.din(w_dff_A_4ouY8qtj9_1),.clk(gclk));
	jdff dff_A_F4FUDs3M5_1(.dout(w_dff_A_4ouY8qtj9_1),.din(w_dff_A_F4FUDs3M5_1),.clk(gclk));
	jdff dff_A_TLumZ1LD0_1(.dout(w_dff_A_F4FUDs3M5_1),.din(w_dff_A_TLumZ1LD0_1),.clk(gclk));
	jdff dff_A_nq8MFM1V3_1(.dout(w_dff_A_TLumZ1LD0_1),.din(w_dff_A_nq8MFM1V3_1),.clk(gclk));
	jdff dff_A_OpuR5ybL5_1(.dout(w_dff_A_nq8MFM1V3_1),.din(w_dff_A_OpuR5ybL5_1),.clk(gclk));
	jdff dff_A_Kyfo73fF2_1(.dout(w_dff_A_OpuR5ybL5_1),.din(w_dff_A_Kyfo73fF2_1),.clk(gclk));
	jdff dff_A_OAl2Lzxh7_1(.dout(w_dff_A_Kyfo73fF2_1),.din(w_dff_A_OAl2Lzxh7_1),.clk(gclk));
	jdff dff_A_D5i4tLOH4_1(.dout(w_dff_A_OAl2Lzxh7_1),.din(w_dff_A_D5i4tLOH4_1),.clk(gclk));
	jdff dff_A_1Perz2kI6_1(.dout(w_dff_A_D5i4tLOH4_1),.din(w_dff_A_1Perz2kI6_1),.clk(gclk));
	jdff dff_A_qGhmJ1uq6_1(.dout(w_dff_A_1Perz2kI6_1),.din(w_dff_A_qGhmJ1uq6_1),.clk(gclk));
	jdff dff_A_uod133Nn2_1(.dout(w_dff_A_qGhmJ1uq6_1),.din(w_dff_A_uod133Nn2_1),.clk(gclk));
	jdff dff_A_fKRahply6_1(.dout(w_dff_A_uod133Nn2_1),.din(w_dff_A_fKRahply6_1),.clk(gclk));
	jdff dff_B_KmuGB4Wa4_1(.din(n1600),.dout(w_dff_B_KmuGB4Wa4_1),.clk(gclk));
	jdff dff_B_2bHVAlJb1_1(.din(w_dff_B_KmuGB4Wa4_1),.dout(w_dff_B_2bHVAlJb1_1),.clk(gclk));
	jdff dff_B_iWpnZ9fZ2_0(.din(n1614),.dout(w_dff_B_iWpnZ9fZ2_0),.clk(gclk));
	jdff dff_B_KmjT6LZ54_0(.din(w_dff_B_iWpnZ9fZ2_0),.dout(w_dff_B_KmjT6LZ54_0),.clk(gclk));
	jdff dff_B_QXQtFWVM3_0(.din(w_dff_B_KmjT6LZ54_0),.dout(w_dff_B_QXQtFWVM3_0),.clk(gclk));
	jdff dff_B_KEuu4M2p9_0(.din(w_dff_B_QXQtFWVM3_0),.dout(w_dff_B_KEuu4M2p9_0),.clk(gclk));
	jdff dff_A_jmLmb4bc5_0(.dout(w_n1613_0[0]),.din(w_dff_A_jmLmb4bc5_0),.clk(gclk));
	jdff dff_A_SdXrTuRN7_0(.dout(w_dff_A_jmLmb4bc5_0),.din(w_dff_A_SdXrTuRN7_0),.clk(gclk));
	jdff dff_A_KftsghUC4_0(.dout(w_n865_0[0]),.din(w_dff_A_KftsghUC4_0),.clk(gclk));
	jdff dff_A_zQUxjSjB4_0(.dout(w_dff_A_KftsghUC4_0),.din(w_dff_A_zQUxjSjB4_0),.clk(gclk));
	jdff dff_A_1iPsS97d8_0(.dout(w_dff_A_zQUxjSjB4_0),.din(w_dff_A_1iPsS97d8_0),.clk(gclk));
	jdff dff_A_S4J3oz055_0(.dout(w_dff_A_1iPsS97d8_0),.din(w_dff_A_S4J3oz055_0),.clk(gclk));
	jdff dff_A_tLTauKTU4_2(.dout(w_n865_0[2]),.din(w_dff_A_tLTauKTU4_2),.clk(gclk));
	jdff dff_A_8QoqLDaH3_2(.dout(w_dff_A_tLTauKTU4_2),.din(w_dff_A_8QoqLDaH3_2),.clk(gclk));
	jdff dff_A_j64Xv3qz2_2(.dout(w_dff_A_8QoqLDaH3_2),.din(w_dff_A_j64Xv3qz2_2),.clk(gclk));
	jdff dff_A_i3G21l3P2_2(.dout(w_dff_A_j64Xv3qz2_2),.din(w_dff_A_i3G21l3P2_2),.clk(gclk));
	jdff dff_A_QqAqicj04_2(.dout(w_dff_A_i3G21l3P2_2),.din(w_dff_A_QqAqicj04_2),.clk(gclk));
	jdff dff_A_6POUhTop1_1(.dout(w_n587_0[1]),.din(w_dff_A_6POUhTop1_1),.clk(gclk));
	jdff dff_A_uIGeh2Lg0_1(.dout(w_dff_A_6POUhTop1_1),.din(w_dff_A_uIGeh2Lg0_1),.clk(gclk));
	jdff dff_A_Nbzwjh4j8_1(.dout(w_dff_A_uIGeh2Lg0_1),.din(w_dff_A_Nbzwjh4j8_1),.clk(gclk));
	jdff dff_A_oC8bNNVc9_1(.dout(w_dff_A_Nbzwjh4j8_1),.din(w_dff_A_oC8bNNVc9_1),.clk(gclk));
	jdff dff_B_yCM6XrYW8_0(.din(n585),.dout(w_dff_B_yCM6XrYW8_0),.clk(gclk));
	jdff dff_B_LGHcPilM5_1(.din(G241),.dout(w_dff_B_LGHcPilM5_1),.clk(gclk));
	jdff dff_B_eWV88eXH9_1(.din(n1601),.dout(w_dff_B_eWV88eXH9_1),.clk(gclk));
	jdff dff_B_FjYJOSeL0_1(.din(w_dff_B_eWV88eXH9_1),.dout(w_dff_B_FjYJOSeL0_1),.clk(gclk));
	jdff dff_B_xDHxEj471_1(.din(w_dff_B_FjYJOSeL0_1),.dout(w_dff_B_xDHxEj471_1),.clk(gclk));
	jdff dff_B_9qF6hteK6_1(.din(n1602),.dout(w_dff_B_9qF6hteK6_1),.clk(gclk));
	jdff dff_B_RS5LCjhX5_1(.din(w_dff_B_9qF6hteK6_1),.dout(w_dff_B_RS5LCjhX5_1),.clk(gclk));
	jdff dff_A_Z638JVzt5_1(.dout(w_n687_0[1]),.din(w_dff_A_Z638JVzt5_1),.clk(gclk));
	jdff dff_A_CvzPEdAw0_1(.dout(w_dff_A_Z638JVzt5_1),.din(w_dff_A_CvzPEdAw0_1),.clk(gclk));
	jdff dff_A_5jgei4zv9_1(.dout(w_dff_A_CvzPEdAw0_1),.din(w_dff_A_5jgei4zv9_1),.clk(gclk));
	jdff dff_A_thC6SE5m2_1(.dout(w_n686_0[1]),.din(w_dff_A_thC6SE5m2_1),.clk(gclk));
	jdff dff_A_v8XxsTxc9_1(.dout(w_dff_A_thC6SE5m2_1),.din(w_dff_A_v8XxsTxc9_1),.clk(gclk));
	jdff dff_A_hur0nhdE9_1(.dout(w_dff_A_v8XxsTxc9_1),.din(w_dff_A_hur0nhdE9_1),.clk(gclk));
	jdff dff_A_2tTVCuS14_1(.dout(w_dff_A_hur0nhdE9_1),.din(w_dff_A_2tTVCuS14_1),.clk(gclk));
	jdff dff_A_h5ww4nX32_0(.dout(w_n581_0[0]),.din(w_dff_A_h5ww4nX32_0),.clk(gclk));
	jdff dff_A_IP7kNLv53_0(.dout(w_dff_A_h5ww4nX32_0),.din(w_dff_A_IP7kNLv53_0),.clk(gclk));
	jdff dff_A_3drH5Idj8_1(.dout(w_n579_1[1]),.din(w_dff_A_3drH5Idj8_1),.clk(gclk));
	jdff dff_A_oXcb4rub9_1(.dout(w_n579_0[1]),.din(w_dff_A_oXcb4rub9_1),.clk(gclk));
	jdff dff_A_NVFluDeo3_2(.dout(w_n579_0[2]),.din(w_dff_A_NVFluDeo3_2),.clk(gclk));
	jdff dff_A_VL4FUWSr8_2(.dout(w_dff_A_NVFluDeo3_2),.din(w_dff_A_VL4FUWSr8_2),.clk(gclk));
	jdff dff_A_vLl8KNLZ3_2(.dout(w_dff_A_VL4FUWSr8_2),.din(w_dff_A_vLl8KNLZ3_2),.clk(gclk));
	jdff dff_A_apldzcTr2_2(.dout(w_dff_A_vLl8KNLZ3_2),.din(w_dff_A_apldzcTr2_2),.clk(gclk));
	jdff dff_B_36jfe22f8_0(.din(n577),.dout(w_dff_B_36jfe22f8_0),.clk(gclk));
	jdff dff_B_rh2BxCzh4_1(.din(G264),.dout(w_dff_B_rh2BxCzh4_1),.clk(gclk));
	jdff dff_A_PZqyPr7U8_1(.dout(w_n574_0[1]),.din(w_dff_A_PZqyPr7U8_1),.clk(gclk));
	jdff dff_A_ZC2bstJW3_1(.dout(w_dff_A_PZqyPr7U8_1),.din(w_dff_A_ZC2bstJW3_1),.clk(gclk));
	jdff dff_A_oMKzX95G8_0(.dout(w_n1599_0[0]),.din(w_dff_A_oMKzX95G8_0),.clk(gclk));
	jdff dff_A_DCcBNEoT4_0(.dout(w_dff_A_oMKzX95G8_0),.din(w_dff_A_DCcBNEoT4_0),.clk(gclk));
	jdff dff_B_UZ0RO1iU3_0(.din(n1598),.dout(w_dff_B_UZ0RO1iU3_0),.clk(gclk));
	jdff dff_B_xzfxRi8R7_0(.din(n1597),.dout(w_dff_B_xzfxRi8R7_0),.clk(gclk));
	jdff dff_B_NbMeyCxI1_0(.din(n1589),.dout(w_dff_B_NbMeyCxI1_0),.clk(gclk));
	jdff dff_A_E8RvXwhG7_0(.dout(w_n573_0[0]),.din(w_dff_A_E8RvXwhG7_0),.clk(gclk));
	jdff dff_A_LlCKywvu0_1(.dout(w_n573_0[1]),.din(w_dff_A_LlCKywvu0_1),.clk(gclk));
	jdff dff_A_6f9bX2tD6_1(.dout(w_dff_A_LlCKywvu0_1),.din(w_dff_A_6f9bX2tD6_1),.clk(gclk));
	jdff dff_B_I6rSOM260_1(.din(n691),.dout(w_dff_B_I6rSOM260_1),.clk(gclk));
	jdff dff_A_s88eH5Y14_0(.dout(w_n695_0[0]),.din(w_dff_A_s88eH5Y14_0),.clk(gclk));
	jdff dff_A_Qe9sEAx29_1(.dout(w_n695_0[1]),.din(w_dff_A_Qe9sEAx29_1),.clk(gclk));
	jdff dff_A_NHIWFKCJ9_1(.dout(w_n564_0[1]),.din(w_dff_A_NHIWFKCJ9_1),.clk(gclk));
	jdff dff_B_hQ7pqEYK6_1(.din(G280),.dout(w_dff_B_hQ7pqEYK6_1),.clk(gclk));
	jdff dff_A_2L149ccd6_0(.dout(w_n562_0[0]),.din(w_dff_A_2L149ccd6_0),.clk(gclk));
	jdff dff_A_Hv98Ul3Y0_0(.dout(w_n692_0[0]),.din(w_dff_A_Hv98Ul3Y0_0),.clk(gclk));
	jdff dff_A_s2LmmwUv5_1(.dout(w_n559_0[1]),.din(w_dff_A_s2LmmwUv5_1),.clk(gclk));
	jdff dff_B_dcyVP1xp6_1(.din(G288),.dout(w_dff_B_dcyVP1xp6_1),.clk(gclk));
	jdff dff_A_zuN3zQmS5_0(.dout(w_n557_0[0]),.din(w_dff_A_zuN3zQmS5_0),.clk(gclk));
	jdff dff_A_qDxhoPsK9_0(.dout(w_n690_0[0]),.din(w_dff_A_qDxhoPsK9_0),.clk(gclk));
	jdff dff_A_hl6HUjuu1_0(.dout(w_dff_A_qDxhoPsK9_0),.din(w_dff_A_hl6HUjuu1_0),.clk(gclk));
	jdff dff_A_b2al5vls9_1(.dout(w_n571_0[1]),.din(w_dff_A_b2al5vls9_1),.clk(gclk));
	jdff dff_B_WxmNg9VF5_1(.din(G272),.dout(w_dff_B_WxmNg9VF5_1),.clk(gclk));
	jdff dff_A_v4ndQapO6_0(.dout(w_n569_0[0]),.din(w_dff_A_v4ndQapO6_0),.clk(gclk));
	jdff dff_A_vm5gbBGa0_0(.dout(w_n485_1[0]),.din(w_dff_A_vm5gbBGa0_0),.clk(gclk));
	jdff dff_A_K02QV1Jy0_0(.dout(w_dff_A_vm5gbBGa0_0),.din(w_dff_A_K02QV1Jy0_0),.clk(gclk));
	jdff dff_B_889MNSiZ3_0(.din(n1585),.dout(w_dff_B_889MNSiZ3_0),.clk(gclk));
	jdff dff_B_Q1twm8zD2_1(.din(n1575),.dout(w_dff_B_Q1twm8zD2_1),.clk(gclk));
	jdff dff_B_EtmbtrLr8_1(.din(w_dff_B_Q1twm8zD2_1),.dout(w_dff_B_EtmbtrLr8_1),.clk(gclk));
	jdff dff_A_oLekoJB74_0(.dout(w_G210_2[0]),.din(w_dff_A_oLekoJB74_0),.clk(gclk));
	jdff dff_A_v255Axo79_1(.dout(w_n451_0[1]),.din(w_dff_A_v255Axo79_1),.clk(gclk));
	jdff dff_A_begpvNal4_1(.dout(w_dff_A_v255Axo79_1),.din(w_dff_A_begpvNal4_1),.clk(gclk));
	jdff dff_B_fLnXQ0Lb0_3(.din(n451),.dout(w_dff_B_fLnXQ0Lb0_3),.clk(gclk));
	jdff dff_A_8eZYEhHf5_0(.dout(w_G457_1[0]),.din(w_dff_A_8eZYEhHf5_0),.clk(gclk));
	jdff dff_A_j9NSDTOJ0_0(.dout(w_dff_A_8eZYEhHf5_0),.din(w_dff_A_j9NSDTOJ0_0),.clk(gclk));
	jdff dff_A_9ln3n0g28_0(.dout(w_dff_A_j9NSDTOJ0_0),.din(w_dff_A_9ln3n0g28_0),.clk(gclk));
	jdff dff_A_ofFN2KXF6_0(.dout(w_dff_A_9ln3n0g28_0),.din(w_dff_A_ofFN2KXF6_0),.clk(gclk));
	jdff dff_A_IvhJg8688_1(.dout(w_G457_1[1]),.din(w_dff_A_IvhJg8688_1),.clk(gclk));
	jdff dff_A_Fz4uHTIG0_1(.dout(w_dff_A_IvhJg8688_1),.din(w_dff_A_Fz4uHTIG0_1),.clk(gclk));
	jdff dff_A_L5HpIfiT5_1(.dout(w_dff_A_Fz4uHTIG0_1),.din(w_dff_A_L5HpIfiT5_1),.clk(gclk));
	jdff dff_A_j1EMTddv1_1(.dout(w_G457_0[1]),.din(w_dff_A_j1EMTddv1_1),.clk(gclk));
	jdff dff_A_1KzzcdFs5_1(.dout(w_dff_A_j1EMTddv1_1),.din(w_dff_A_1KzzcdFs5_1),.clk(gclk));
	jdff dff_A_y63zbw8x4_1(.dout(w_dff_A_1KzzcdFs5_1),.din(w_dff_A_y63zbw8x4_1),.clk(gclk));
	jdff dff_A_cKOUHrFF9_2(.dout(w_G457_0[2]),.din(w_dff_A_cKOUHrFF9_2),.clk(gclk));
	jdff dff_A_rmmWmvdv0_2(.dout(w_dff_A_cKOUHrFF9_2),.din(w_dff_A_rmmWmvdv0_2),.clk(gclk));
	jdff dff_A_YXtTpnJ03_2(.dout(w_dff_A_rmmWmvdv0_2),.din(w_dff_A_YXtTpnJ03_2),.clk(gclk));
	jdff dff_A_SfgBxLJ12_2(.dout(w_dff_A_YXtTpnJ03_2),.din(w_dff_A_SfgBxLJ12_2),.clk(gclk));
	jdff dff_A_ObGN1cyK6_2(.dout(w_G210_0[2]),.din(w_dff_A_ObGN1cyK6_2),.clk(gclk));
	jdff dff_B_wX4VpuQn3_1(.din(n1570),.dout(w_dff_B_wX4VpuQn3_1),.clk(gclk));
	jdff dff_A_5zvoiHyn4_0(.dout(w_n509_0[0]),.din(w_dff_A_5zvoiHyn4_0),.clk(gclk));
	jdff dff_A_qvgEtbMD4_1(.dout(w_n509_0[1]),.din(w_dff_A_qvgEtbMD4_1),.clk(gclk));
	jdff dff_A_g2ibEBXg4_1(.dout(w_dff_A_qvgEtbMD4_1),.din(w_dff_A_g2ibEBXg4_1),.clk(gclk));
	jdff dff_B_HKAzCg7R7_3(.din(n509),.dout(w_dff_B_HKAzCg7R7_3),.clk(gclk));
	jdff dff_A_ZPEVKmD71_0(.dout(w_G468_1[0]),.din(w_dff_A_ZPEVKmD71_0),.clk(gclk));
	jdff dff_A_FkFWjuf19_0(.dout(w_dff_A_ZPEVKmD71_0),.din(w_dff_A_FkFWjuf19_0),.clk(gclk));
	jdff dff_A_MAAjVj5D3_0(.dout(w_dff_A_FkFWjuf19_0),.din(w_dff_A_MAAjVj5D3_0),.clk(gclk));
	jdff dff_A_A5Y9CIJd1_0(.dout(w_dff_A_MAAjVj5D3_0),.din(w_dff_A_A5Y9CIJd1_0),.clk(gclk));
	jdff dff_A_6IczPJFg8_1(.dout(w_G468_1[1]),.din(w_dff_A_6IczPJFg8_1),.clk(gclk));
	jdff dff_A_kk6Xg4d20_1(.dout(w_dff_A_6IczPJFg8_1),.din(w_dff_A_kk6Xg4d20_1),.clk(gclk));
	jdff dff_A_UmtnvGTW6_1(.dout(w_dff_A_kk6Xg4d20_1),.din(w_dff_A_UmtnvGTW6_1),.clk(gclk));
	jdff dff_B_d0nm04rx4_1(.din(n1566),.dout(w_dff_B_d0nm04rx4_1),.clk(gclk));
	jdff dff_A_omqAYVWi0_0(.dout(w_G218_1[0]),.din(w_dff_A_omqAYVWi0_0),.clk(gclk));
	jdff dff_A_dOKrPts53_1(.dout(w_G468_0[1]),.din(w_dff_A_dOKrPts53_1),.clk(gclk));
	jdff dff_A_Zllgn7rC3_1(.dout(w_dff_A_dOKrPts53_1),.din(w_dff_A_Zllgn7rC3_1),.clk(gclk));
	jdff dff_A_M1BjK6yz4_2(.dout(w_G468_0[2]),.din(w_dff_A_M1BjK6yz4_2),.clk(gclk));
	jdff dff_A_X80VAKJu5_2(.dout(w_dff_A_M1BjK6yz4_2),.din(w_dff_A_X80VAKJu5_2),.clk(gclk));
	jdff dff_A_QVEhdUTm7_2(.dout(w_dff_A_X80VAKJu5_2),.din(w_dff_A_QVEhdUTm7_2),.clk(gclk));
	jdff dff_A_C4MnImA90_2(.dout(w_dff_A_QVEhdUTm7_2),.din(w_dff_A_C4MnImA90_2),.clk(gclk));
	jdff dff_A_GfG3u0CN9_0(.dout(w_G218_2[0]),.din(w_dff_A_GfG3u0CN9_0),.clk(gclk));
	jdff dff_B_Evnm23O15_1(.din(n1556),.dout(w_dff_B_Evnm23O15_1),.clk(gclk));
	jdff dff_B_2GqOtywX5_1(.din(w_dff_B_Evnm23O15_1),.dout(w_dff_B_2GqOtywX5_1),.clk(gclk));
	jdff dff_A_jKyEDYcW2_0(.dout(w_G226_2[0]),.din(w_dff_A_jKyEDYcW2_0),.clk(gclk));
	jdff dff_A_EnrzktwJ9_2(.dout(w_n496_0[2]),.din(w_dff_A_EnrzktwJ9_2),.clk(gclk));
	jdff dff_A_2XBEw37y9_2(.dout(w_dff_A_EnrzktwJ9_2),.din(w_dff_A_2XBEw37y9_2),.clk(gclk));
	jdff dff_A_Kof4lzNX5_2(.dout(w_dff_A_2XBEw37y9_2),.din(w_dff_A_Kof4lzNX5_2),.clk(gclk));
	jdff dff_B_OzpKQcnl0_3(.din(n496),.dout(w_dff_B_OzpKQcnl0_3),.clk(gclk));
	jdff dff_A_p5OtCipC7_0(.dout(w_G422_1[0]),.din(w_dff_A_p5OtCipC7_0),.clk(gclk));
	jdff dff_A_LtzjnPaH2_0(.dout(w_dff_A_p5OtCipC7_0),.din(w_dff_A_LtzjnPaH2_0),.clk(gclk));
	jdff dff_A_byQV1EwN1_0(.dout(w_dff_A_LtzjnPaH2_0),.din(w_dff_A_byQV1EwN1_0),.clk(gclk));
	jdff dff_A_67X00Ndi9_1(.dout(w_G422_0[1]),.din(w_dff_A_67X00Ndi9_1),.clk(gclk));
	jdff dff_A_uxQAF81y4_1(.dout(w_dff_A_67X00Ndi9_1),.din(w_dff_A_uxQAF81y4_1),.clk(gclk));
	jdff dff_A_sS3oEy2s3_1(.dout(w_dff_A_uxQAF81y4_1),.din(w_dff_A_sS3oEy2s3_1),.clk(gclk));
	jdff dff_A_e1WClZRI7_2(.dout(w_G422_0[2]),.din(w_dff_A_e1WClZRI7_2),.clk(gclk));
	jdff dff_A_pbJw1qfz5_2(.dout(w_dff_A_e1WClZRI7_2),.din(w_dff_A_pbJw1qfz5_2),.clk(gclk));
	jdff dff_A_U6Ikx0Vg4_2(.dout(w_dff_A_pbJw1qfz5_2),.din(w_dff_A_U6Ikx0Vg4_2),.clk(gclk));
	jdff dff_A_M0zNXlLG7_2(.dout(w_dff_A_U6Ikx0Vg4_2),.din(w_dff_A_M0zNXlLG7_2),.clk(gclk));
	jdff dff_A_gT9buK4T4_2(.dout(w_G226_0[2]),.din(w_dff_A_gT9buK4T4_2),.clk(gclk));
	jdff dff_B_MT3m1v0b3_1(.din(n541),.dout(w_dff_B_MT3m1v0b3_1),.clk(gclk));
	jdff dff_B_Iy94drE61_1(.din(w_dff_B_MT3m1v0b3_1),.dout(w_dff_B_Iy94drE61_1),.clk(gclk));
	jdff dff_B_VYw4pF030_1(.din(n542),.dout(w_dff_B_VYw4pF030_1),.clk(gclk));
	jdff dff_A_vMNUiQfu8_0(.dout(w_G446_1[0]),.din(w_dff_A_vMNUiQfu8_0),.clk(gclk));
	jdff dff_A_KR7BGXZC0_0(.dout(w_dff_A_vMNUiQfu8_0),.din(w_dff_A_KR7BGXZC0_0),.clk(gclk));
	jdff dff_A_ofgL8hNt0_0(.dout(w_dff_A_KR7BGXZC0_0),.din(w_dff_A_ofgL8hNt0_0),.clk(gclk));
	jdff dff_A_PoDJRc4n1_1(.dout(w_G446_1[1]),.din(w_dff_A_PoDJRc4n1_1),.clk(gclk));
	jdff dff_A_1GH9ejTP0_1(.dout(w_dff_A_PoDJRc4n1_1),.din(w_dff_A_1GH9ejTP0_1),.clk(gclk));
	jdff dff_A_ClsEoZwW8_1(.dout(w_dff_A_1GH9ejTP0_1),.din(w_dff_A_ClsEoZwW8_1),.clk(gclk));
	jdff dff_A_d9umcNL71_1(.dout(w_G446_0[1]),.din(w_dff_A_d9umcNL71_1),.clk(gclk));
	jdff dff_A_m1ayBrvp4_1(.dout(w_dff_A_d9umcNL71_1),.din(w_dff_A_m1ayBrvp4_1),.clk(gclk));
	jdff dff_A_ZxaHmWHq9_1(.dout(w_dff_A_m1ayBrvp4_1),.din(w_dff_A_ZxaHmWHq9_1),.clk(gclk));
	jdff dff_A_TKLUWJgi2_2(.dout(w_G446_0[2]),.din(w_dff_A_TKLUWJgi2_2),.clk(gclk));
	jdff dff_A_77SFOBKl7_2(.dout(w_dff_A_TKLUWJgi2_2),.din(w_dff_A_77SFOBKl7_2),.clk(gclk));
	jdff dff_A_Mmgn51Xh7_2(.dout(w_dff_A_77SFOBKl7_2),.din(w_dff_A_Mmgn51Xh7_2),.clk(gclk));
	jdff dff_A_5HCCnfVr4_0(.dout(w_G206_1[0]),.din(w_dff_A_5HCCnfVr4_0),.clk(gclk));
	jdff dff_B_UhzF9ryi3_1(.din(n1525),.dout(w_dff_B_UhzF9ryi3_1),.clk(gclk));
	jdff dff_B_wNMw5I5N0_1(.din(n1534),.dout(w_dff_B_wNMw5I5N0_1),.clk(gclk));
	jdff dff_B_tRZZYgo67_1(.din(n1544),.dout(w_dff_B_tRZZYgo67_1),.clk(gclk));
	jdff dff_B_SeD0dRPb3_1(.din(w_dff_B_tRZZYgo67_1),.dout(w_dff_B_SeD0dRPb3_1),.clk(gclk));
	jdff dff_A_IAv7bVlJ3_0(.dout(w_G234_2[0]),.din(w_dff_A_IAv7bVlJ3_0),.clk(gclk));
	jdff dff_A_k3UyB8Po6_1(.dout(w_n462_0[1]),.din(w_dff_A_k3UyB8Po6_1),.clk(gclk));
	jdff dff_A_KZ8wSDaz2_1(.dout(w_dff_A_k3UyB8Po6_1),.din(w_dff_A_KZ8wSDaz2_1),.clk(gclk));
	jdff dff_A_vrW7pce47_1(.dout(w_dff_A_KZ8wSDaz2_1),.din(w_dff_A_vrW7pce47_1),.clk(gclk));
	jdff dff_B_d2dBaqaS5_3(.din(n462),.dout(w_dff_B_d2dBaqaS5_3),.clk(gclk));
	jdff dff_A_ixjX31sh3_0(.dout(w_G435_1[0]),.din(w_dff_A_ixjX31sh3_0),.clk(gclk));
	jdff dff_A_GtMqQLe60_0(.dout(w_dff_A_ixjX31sh3_0),.din(w_dff_A_GtMqQLe60_0),.clk(gclk));
	jdff dff_A_YbWXFDCo7_0(.dout(w_dff_A_GtMqQLe60_0),.din(w_dff_A_YbWXFDCo7_0),.clk(gclk));
	jdff dff_A_ZOupd35Q9_0(.dout(w_dff_A_YbWXFDCo7_0),.din(w_dff_A_ZOupd35Q9_0),.clk(gclk));
	jdff dff_A_4nBuZFG15_1(.dout(w_G435_1[1]),.din(w_dff_A_4nBuZFG15_1),.clk(gclk));
	jdff dff_A_fZxMoYKW5_1(.dout(w_dff_A_4nBuZFG15_1),.din(w_dff_A_fZxMoYKW5_1),.clk(gclk));
	jdff dff_A_lrnp6gFq2_1(.dout(w_dff_A_fZxMoYKW5_1),.din(w_dff_A_lrnp6gFq2_1),.clk(gclk));
	jdff dff_A_Nnii9NIS3_1(.dout(w_G435_0[1]),.din(w_dff_A_Nnii9NIS3_1),.clk(gclk));
	jdff dff_A_a1yMwuBY3_1(.dout(w_dff_A_Nnii9NIS3_1),.din(w_dff_A_a1yMwuBY3_1),.clk(gclk));
	jdff dff_A_qaPcEWrT7_1(.dout(w_dff_A_a1yMwuBY3_1),.din(w_dff_A_qaPcEWrT7_1),.clk(gclk));
	jdff dff_A_N81RKIix8_2(.dout(w_G435_0[2]),.din(w_dff_A_N81RKIix8_2),.clk(gclk));
	jdff dff_A_sFDtG4JR7_2(.dout(w_dff_A_N81RKIix8_2),.din(w_dff_A_sFDtG4JR7_2),.clk(gclk));
	jdff dff_A_Noi6SRXT0_2(.dout(w_dff_A_sFDtG4JR7_2),.din(w_dff_A_Noi6SRXT0_2),.clk(gclk));
	jdff dff_A_8lsHxblE7_2(.dout(w_dff_A_Noi6SRXT0_2),.din(w_dff_A_8lsHxblE7_2),.clk(gclk));
	jdff dff_A_zJ4OzjGQ4_2(.dout(w_G234_0[2]),.din(w_dff_A_zJ4OzjGQ4_2),.clk(gclk));
	jdff dff_B_m6dmyI8h8_1(.din(n1535),.dout(w_dff_B_m6dmyI8h8_1),.clk(gclk));
	jdff dff_B_GsQmPUvU2_1(.din(w_dff_B_m6dmyI8h8_1),.dout(w_dff_B_GsQmPUvU2_1),.clk(gclk));
	jdff dff_A_jWHGvtCa9_0(.dout(w_G257_2[0]),.din(w_dff_A_jWHGvtCa9_0),.clk(gclk));
	jdff dff_A_LwEQZpPG1_1(.dout(w_n520_0[1]),.din(w_dff_A_LwEQZpPG1_1),.clk(gclk));
	jdff dff_A_SsfZd5P01_1(.dout(w_dff_A_LwEQZpPG1_1),.din(w_dff_A_SsfZd5P01_1),.clk(gclk));
	jdff dff_B_9BYI8BGR2_3(.din(n520),.dout(w_dff_B_9BYI8BGR2_3),.clk(gclk));
	jdff dff_A_jk3Igepg2_0(.dout(w_G389_1[0]),.din(w_dff_A_jk3Igepg2_0),.clk(gclk));
	jdff dff_A_A3snWA4u5_0(.dout(w_dff_A_jk3Igepg2_0),.din(w_dff_A_A3snWA4u5_0),.clk(gclk));
	jdff dff_A_8CYTgtUW9_0(.dout(w_dff_A_A3snWA4u5_0),.din(w_dff_A_8CYTgtUW9_0),.clk(gclk));
	jdff dff_A_SWo3DVyA2_0(.dout(w_dff_A_8CYTgtUW9_0),.din(w_dff_A_SWo3DVyA2_0),.clk(gclk));
	jdff dff_A_VxC4n2dU9_1(.dout(w_G389_1[1]),.din(w_dff_A_VxC4n2dU9_1),.clk(gclk));
	jdff dff_A_QxBoCB4y1_1(.dout(w_dff_A_VxC4n2dU9_1),.din(w_dff_A_QxBoCB4y1_1),.clk(gclk));
	jdff dff_A_VgDuH2sX9_1(.dout(w_dff_A_QxBoCB4y1_1),.din(w_dff_A_VgDuH2sX9_1),.clk(gclk));
	jdff dff_A_McdFHEj28_1(.dout(w_G389_0[1]),.din(w_dff_A_McdFHEj28_1),.clk(gclk));
	jdff dff_A_SSYCyo4y7_1(.dout(w_dff_A_McdFHEj28_1),.din(w_dff_A_SSYCyo4y7_1),.clk(gclk));
	jdff dff_A_RU41QhYS4_1(.dout(w_dff_A_SSYCyo4y7_1),.din(w_dff_A_RU41QhYS4_1),.clk(gclk));
	jdff dff_A_BYPkcyG07_2(.dout(w_G389_0[2]),.din(w_dff_A_BYPkcyG07_2),.clk(gclk));
	jdff dff_A_SpExcGnA3_2(.dout(w_dff_A_BYPkcyG07_2),.din(w_dff_A_SpExcGnA3_2),.clk(gclk));
	jdff dff_A_xlgPmUFB1_2(.dout(w_dff_A_SpExcGnA3_2),.din(w_dff_A_xlgPmUFB1_2),.clk(gclk));
	jdff dff_A_A8WUKmeI4_2(.dout(w_dff_A_xlgPmUFB1_2),.din(w_dff_A_A8WUKmeI4_2),.clk(gclk));
	jdff dff_A_CID2Snx76_2(.dout(w_G257_0[2]),.din(w_dff_A_CID2Snx76_2),.clk(gclk));
	jdff dff_B_vQWbygcP6_1(.din(n1530),.dout(w_dff_B_vQWbygcP6_1),.clk(gclk));
	jdff dff_A_TJDdjxDN3_1(.dout(w_n485_0[1]),.din(w_dff_A_TJDdjxDN3_1),.clk(gclk));
	jdff dff_A_Fq7oCxoN3_1(.dout(w_dff_A_TJDdjxDN3_1),.din(w_dff_A_Fq7oCxoN3_1),.clk(gclk));
	jdff dff_A_pMW24VFp3_2(.dout(w_n485_0[2]),.din(w_dff_A_pMW24VFp3_2),.clk(gclk));
	jdff dff_B_5B0514A33_3(.din(n485),.dout(w_dff_B_5B0514A33_3),.clk(gclk));
	jdff dff_A_0HziCBUR3_0(.dout(w_G400_1[0]),.din(w_dff_A_0HziCBUR3_0),.clk(gclk));
	jdff dff_A_xtl1iMlQ9_0(.dout(w_dff_A_0HziCBUR3_0),.din(w_dff_A_xtl1iMlQ9_0),.clk(gclk));
	jdff dff_A_I4r5TiI65_0(.dout(w_dff_A_xtl1iMlQ9_0),.din(w_dff_A_I4r5TiI65_0),.clk(gclk));
	jdff dff_A_PRE9t4K11_0(.dout(w_dff_A_I4r5TiI65_0),.din(w_dff_A_PRE9t4K11_0),.clk(gclk));
	jdff dff_A_CDgMUzjN4_1(.dout(w_G400_1[1]),.din(w_dff_A_CDgMUzjN4_1),.clk(gclk));
	jdff dff_A_mGBU1vtR5_1(.dout(w_dff_A_CDgMUzjN4_1),.din(w_dff_A_mGBU1vtR5_1),.clk(gclk));
	jdff dff_A_BcsnzGcI1_1(.dout(w_dff_A_mGBU1vtR5_1),.din(w_dff_A_BcsnzGcI1_1),.clk(gclk));
	jdff dff_B_ii3wpd5b0_1(.din(n1526),.dout(w_dff_B_ii3wpd5b0_1),.clk(gclk));
	jdff dff_A_J1GBjRnw5_0(.dout(w_G251_5[0]),.din(w_dff_A_J1GBjRnw5_0),.clk(gclk));
	jdff dff_A_iW6HyRsz8_0(.dout(w_G251_1[0]),.din(w_dff_A_iW6HyRsz8_0),.clk(gclk));
	jdff dff_A_3HPeGmjr0_2(.dout(w_G251_1[2]),.din(w_dff_A_3HPeGmjr0_2),.clk(gclk));
	jdff dff_A_Xe8Fmw9H8_1(.dout(w_G400_0[1]),.din(w_dff_A_Xe8Fmw9H8_1),.clk(gclk));
	jdff dff_A_poS3m5Qm4_1(.dout(w_dff_A_Xe8Fmw9H8_1),.din(w_dff_A_poS3m5Qm4_1),.clk(gclk));
	jdff dff_A_AsvBBfPu7_2(.dout(w_G400_0[2]),.din(w_dff_A_AsvBBfPu7_2),.clk(gclk));
	jdff dff_A_WrXyI5iu0_2(.dout(w_dff_A_AsvBBfPu7_2),.din(w_dff_A_WrXyI5iu0_2),.clk(gclk));
	jdff dff_A_v6NM0Qup3_2(.dout(w_dff_A_WrXyI5iu0_2),.din(w_dff_A_v6NM0Qup3_2),.clk(gclk));
	jdff dff_A_OVVhrC421_2(.dout(w_dff_A_v6NM0Qup3_2),.din(w_dff_A_OVVhrC421_2),.clk(gclk));
	jdff dff_A_yKhhrmpy2_1(.dout(w_G265_1[1]),.din(w_dff_A_yKhhrmpy2_1),.clk(gclk));
	jdff dff_A_c5SsxF4r5_2(.dout(w_G265_0[2]),.din(w_dff_A_c5SsxF4r5_2),.clk(gclk));
	jdff dff_B_9eh08wkv9_1(.din(n1516),.dout(w_dff_B_9eh08wkv9_1),.clk(gclk));
	jdff dff_B_o8C3BcRH5_1(.din(w_dff_B_9eh08wkv9_1),.dout(w_dff_B_o8C3BcRH5_1),.clk(gclk));
	jdff dff_A_YLF0ccXX5_0(.dout(w_G281_2[0]),.din(w_dff_A_YLF0ccXX5_0),.clk(gclk));
	jdff dff_A_NuzqmZ4V1_1(.dout(w_n532_0[1]),.din(w_dff_A_NuzqmZ4V1_1),.clk(gclk));
	jdff dff_A_zxckjhqV0_1(.dout(w_dff_A_NuzqmZ4V1_1),.din(w_dff_A_zxckjhqV0_1),.clk(gclk));
	jdff dff_A_vRi5HaW28_2(.dout(w_n532_0[2]),.din(w_dff_A_vRi5HaW28_2),.clk(gclk));
	jdff dff_A_oEkkQGhu1_2(.dout(w_dff_A_vRi5HaW28_2),.din(w_dff_A_oEkkQGhu1_2),.clk(gclk));
	jdff dff_B_b9meJiND4_3(.din(n532),.dout(w_dff_B_b9meJiND4_3),.clk(gclk));
	jdff dff_A_3BW8hfJP5_0(.dout(w_G374_1[0]),.din(w_dff_A_3BW8hfJP5_0),.clk(gclk));
	jdff dff_A_vZMHX8wm5_0(.dout(w_dff_A_3BW8hfJP5_0),.din(w_dff_A_vZMHX8wm5_0),.clk(gclk));
	jdff dff_A_9TpVP1lK2_0(.dout(w_dff_A_vZMHX8wm5_0),.din(w_dff_A_9TpVP1lK2_0),.clk(gclk));
	jdff dff_A_oxlsLqtp8_0(.dout(w_dff_A_9TpVP1lK2_0),.din(w_dff_A_oxlsLqtp8_0),.clk(gclk));
	jdff dff_A_kYWSXtUk2_1(.dout(w_G374_1[1]),.din(w_dff_A_kYWSXtUk2_1),.clk(gclk));
	jdff dff_A_MfbTLasS1_1(.dout(w_dff_A_kYWSXtUk2_1),.din(w_dff_A_MfbTLasS1_1),.clk(gclk));
	jdff dff_A_pi6uTrMi7_1(.dout(w_dff_A_MfbTLasS1_1),.din(w_dff_A_pi6uTrMi7_1),.clk(gclk));
	jdff dff_A_8d7Ye7kU8_1(.dout(w_G374_0[1]),.din(w_dff_A_8d7Ye7kU8_1),.clk(gclk));
	jdff dff_A_D5okqryN3_1(.dout(w_dff_A_8d7Ye7kU8_1),.din(w_dff_A_D5okqryN3_1),.clk(gclk));
	jdff dff_A_MbOpF8PG8_1(.dout(w_dff_A_D5okqryN3_1),.din(w_dff_A_MbOpF8PG8_1),.clk(gclk));
	jdff dff_A_vRwjoFX78_2(.dout(w_G374_0[2]),.din(w_dff_A_vRwjoFX78_2),.clk(gclk));
	jdff dff_A_2PR6l5d35_2(.dout(w_dff_A_vRwjoFX78_2),.din(w_dff_A_2PR6l5d35_2),.clk(gclk));
	jdff dff_A_XbVAolyy7_2(.dout(w_dff_A_2PR6l5d35_2),.din(w_dff_A_XbVAolyy7_2),.clk(gclk));
	jdff dff_A_5g6MpCxj4_2(.dout(w_dff_A_XbVAolyy7_2),.din(w_dff_A_5g6MpCxj4_2),.clk(gclk));
	jdff dff_A_YoDwKxKM6_2(.dout(w_G281_0[2]),.din(w_dff_A_YoDwKxKM6_2),.clk(gclk));
	jdff dff_A_ObhXBezk2_0(.dout(w_G242_1[0]),.din(w_dff_A_ObhXBezk2_0),.clk(gclk));
	jdff dff_A_vXPYLiIZ1_1(.dout(w_G242_0[1]),.din(w_dff_A_vXPYLiIZ1_1),.clk(gclk));
	jdff dff_A_zeUXuxX64_2(.dout(w_G242_0[2]),.din(w_dff_A_zeUXuxX64_2),.clk(gclk));
	jdff dff_B_J9zxAP4D0_1(.din(n1507),.dout(w_dff_B_J9zxAP4D0_1),.clk(gclk));
	jdff dff_B_4fm55Zox3_1(.din(w_dff_B_J9zxAP4D0_1),.dout(w_dff_B_4fm55Zox3_1),.clk(gclk));
	jdff dff_A_CCG8Zxt41_0(.dout(w_G273_2[0]),.din(w_dff_A_CCG8Zxt41_0),.clk(gclk));
	jdff dff_A_h7Jd0gJN0_1(.dout(w_G251_0[1]),.din(w_dff_A_h7Jd0gJN0_1),.clk(gclk));
	jdff dff_A_DQGrjRHK8_2(.dout(w_G251_0[2]),.din(w_dff_A_DQGrjRHK8_2),.clk(gclk));
	jdff dff_A_AKrFKqE09_1(.dout(w_n473_0[1]),.din(w_dff_A_AKrFKqE09_1),.clk(gclk));
	jdff dff_A_fWW2UeFb7_1(.dout(w_dff_A_AKrFKqE09_1),.din(w_dff_A_fWW2UeFb7_1),.clk(gclk));
	jdff dff_A_JRx1cu4J3_2(.dout(w_n473_0[2]),.din(w_dff_A_JRx1cu4J3_2),.clk(gclk));
	jdff dff_A_r91G5d5d1_2(.dout(w_dff_A_JRx1cu4J3_2),.din(w_dff_A_r91G5d5d1_2),.clk(gclk));
	jdff dff_B_2DsNOHuP7_3(.din(n473),.dout(w_dff_B_2DsNOHuP7_3),.clk(gclk));
	jdff dff_A_ijT9kB0A1_0(.dout(w_G411_2[0]),.din(w_dff_A_ijT9kB0A1_0),.clk(gclk));
	jdff dff_A_Wwvhte7V5_0(.dout(w_dff_A_ijT9kB0A1_0),.din(w_dff_A_Wwvhte7V5_0),.clk(gclk));
	jdff dff_A_El7HS5tF9_0(.dout(w_dff_A_Wwvhte7V5_0),.din(w_dff_A_El7HS5tF9_0),.clk(gclk));
	jdff dff_A_juiEJIiC2_0(.dout(w_G411_0[0]),.din(w_dff_A_juiEJIiC2_0),.clk(gclk));
	jdff dff_A_z5CTrU3b2_0(.dout(w_dff_A_juiEJIiC2_0),.din(w_dff_A_z5CTrU3b2_0),.clk(gclk));
	jdff dff_A_MFdt46Gh2_0(.dout(w_dff_A_z5CTrU3b2_0),.din(w_dff_A_MFdt46Gh2_0),.clk(gclk));
	jdff dff_A_lge6Nse23_0(.dout(w_dff_A_MFdt46Gh2_0),.din(w_dff_A_lge6Nse23_0),.clk(gclk));
	jdff dff_A_kMCUL8xc2_2(.dout(w_G411_0[2]),.din(w_dff_A_kMCUL8xc2_2),.clk(gclk));
	jdff dff_A_QctWO7aU5_2(.dout(w_dff_A_kMCUL8xc2_2),.din(w_dff_A_QctWO7aU5_2),.clk(gclk));
	jdff dff_A_HuQwAL7r3_2(.dout(w_dff_A_QctWO7aU5_2),.din(w_dff_A_HuQwAL7r3_2),.clk(gclk));
	jdff dff_A_AK5xYz0k8_1(.dout(w_G273_1[1]),.din(w_dff_A_AK5xYz0k8_1),.clk(gclk));
	jdff dff_A_4imqgMe79_2(.dout(w_G273_0[2]),.din(w_dff_A_4imqgMe79_2),.clk(gclk));
	jdff dff_A_OfhDr8Jr0_2(.dout(w_G248_3[2]),.din(w_dff_A_OfhDr8Jr0_2),.clk(gclk));
	jdff dff_A_XL4AbLks6_1(.dout(w_n749_4[1]),.din(w_dff_A_XL4AbLks6_1),.clk(gclk));
	jdff dff_A_2ZuXrpe36_1(.dout(w_dff_A_XL4AbLks6_1),.din(w_dff_A_2ZuXrpe36_1),.clk(gclk));
	jdff dff_A_t8w2e87r8_1(.dout(w_dff_A_2ZuXrpe36_1),.din(w_dff_A_t8w2e87r8_1),.clk(gclk));
	jdff dff_A_oPNC0mPF0_1(.dout(w_dff_A_t8w2e87r8_1),.din(w_dff_A_oPNC0mPF0_1),.clk(gclk));
	jdff dff_A_5yGfR4rj6_1(.dout(w_dff_A_oPNC0mPF0_1),.din(w_dff_A_5yGfR4rj6_1),.clk(gclk));
	jdff dff_A_MJ6Hvoij0_1(.dout(w_dff_A_5yGfR4rj6_1),.din(w_dff_A_MJ6Hvoij0_1),.clk(gclk));
	jdff dff_A_RCJMwuVo0_1(.dout(w_dff_A_MJ6Hvoij0_1),.din(w_dff_A_RCJMwuVo0_1),.clk(gclk));
	jdff dff_A_VBAUcQae1_1(.dout(w_dff_A_RCJMwuVo0_1),.din(w_dff_A_VBAUcQae1_1),.clk(gclk));
	jdff dff_A_q49p95m61_1(.dout(w_dff_A_VBAUcQae1_1),.din(w_dff_A_q49p95m61_1),.clk(gclk));
	jdff dff_A_EXDpjo6W6_1(.dout(w_dff_A_q49p95m61_1),.din(w_dff_A_EXDpjo6W6_1),.clk(gclk));
	jdff dff_A_QOcUvxSe8_1(.dout(w_dff_A_EXDpjo6W6_1),.din(w_dff_A_QOcUvxSe8_1),.clk(gclk));
	jdff dff_A_T1dFYe3G1_1(.dout(w_dff_A_QOcUvxSe8_1),.din(w_dff_A_T1dFYe3G1_1),.clk(gclk));
	jdff dff_A_rmSyudrV7_1(.dout(w_dff_A_T1dFYe3G1_1),.din(w_dff_A_rmSyudrV7_1),.clk(gclk));
	jdff dff_A_sgr2C9MX6_1(.dout(w_dff_A_rmSyudrV7_1),.din(w_dff_A_sgr2C9MX6_1),.clk(gclk));
	jdff dff_A_HEfhdYZv6_1(.dout(w_dff_A_sgr2C9MX6_1),.din(w_dff_A_HEfhdYZv6_1),.clk(gclk));
	jdff dff_A_vd0hohDx2_1(.dout(w_dff_A_HEfhdYZv6_1),.din(w_dff_A_vd0hohDx2_1),.clk(gclk));
	jdff dff_A_CQbw284R5_1(.dout(w_dff_A_vd0hohDx2_1),.din(w_dff_A_CQbw284R5_1),.clk(gclk));
	jdff dff_A_qc0WrT8J1_2(.dout(w_n749_4[2]),.din(w_dff_A_qc0WrT8J1_2),.clk(gclk));
	jdff dff_A_oCgrTsBV9_2(.dout(w_dff_A_qc0WrT8J1_2),.din(w_dff_A_oCgrTsBV9_2),.clk(gclk));
	jdff dff_A_HIR4MtVn9_2(.dout(w_dff_A_oCgrTsBV9_2),.din(w_dff_A_HIR4MtVn9_2),.clk(gclk));
	jdff dff_A_KO4VY6Sp8_2(.dout(w_dff_A_HIR4MtVn9_2),.din(w_dff_A_KO4VY6Sp8_2),.clk(gclk));
	jdff dff_A_40Z9CLjG2_2(.dout(w_dff_A_KO4VY6Sp8_2),.din(w_dff_A_40Z9CLjG2_2),.clk(gclk));
	jdff dff_A_8QOhCgk58_2(.dout(w_dff_A_40Z9CLjG2_2),.din(w_dff_A_8QOhCgk58_2),.clk(gclk));
	jdff dff_A_YfRbn58s9_2(.dout(w_dff_A_8QOhCgk58_2),.din(w_dff_A_YfRbn58s9_2),.clk(gclk));
	jdff dff_A_oRDUx95A7_2(.dout(w_dff_A_YfRbn58s9_2),.din(w_dff_A_oRDUx95A7_2),.clk(gclk));
	jdff dff_A_xo8H0iUw2_1(.dout(w_n749_1[1]),.din(w_dff_A_xo8H0iUw2_1),.clk(gclk));
	jdff dff_A_pU6HVoYk6_1(.dout(w_dff_A_xo8H0iUw2_1),.din(w_dff_A_pU6HVoYk6_1),.clk(gclk));
	jdff dff_A_h14ZsECt1_1(.dout(w_dff_A_pU6HVoYk6_1),.din(w_dff_A_h14ZsECt1_1),.clk(gclk));
	jdff dff_A_WSPSDGqZ9_1(.dout(w_dff_A_h14ZsECt1_1),.din(w_dff_A_WSPSDGqZ9_1),.clk(gclk));
	jdff dff_A_9q4aPqhS1_2(.dout(w_n749_1[2]),.din(w_dff_A_9q4aPqhS1_2),.clk(gclk));
	jdff dff_A_yHz3fP6c9_2(.dout(w_dff_A_9q4aPqhS1_2),.din(w_dff_A_yHz3fP6c9_2),.clk(gclk));
	jdff dff_A_dsMB0Ji38_2(.dout(w_dff_A_yHz3fP6c9_2),.din(w_dff_A_dsMB0Ji38_2),.clk(gclk));
	jdff dff_A_MsncRhbx1_2(.dout(w_dff_A_dsMB0Ji38_2),.din(w_dff_A_MsncRhbx1_2),.clk(gclk));
	jdff dff_A_2uW4Q9kK5_1(.dout(w_n749_0[1]),.din(w_dff_A_2uW4Q9kK5_1),.clk(gclk));
	jdff dff_A_lYHRuC0r7_1(.dout(w_dff_A_2uW4Q9kK5_1),.din(w_dff_A_lYHRuC0r7_1),.clk(gclk));
	jdff dff_A_Aur4jt7Q5_2(.dout(w_n749_0[2]),.din(w_dff_A_Aur4jt7Q5_2),.clk(gclk));
	jdff dff_A_71ICoD9D2_2(.dout(w_dff_A_Aur4jt7Q5_2),.din(w_dff_A_71ICoD9D2_2),.clk(gclk));
	jdff dff_A_dbchnsP29_2(.dout(w_dff_A_71ICoD9D2_2),.din(w_dff_A_dbchnsP29_2),.clk(gclk));
	jdff dff_A_VjbP3K595_0(.dout(w_G4091_6[0]),.din(w_dff_A_VjbP3K595_0),.clk(gclk));
	jdff dff_A_86b8CQdR3_0(.dout(w_dff_A_VjbP3K595_0),.din(w_dff_A_86b8CQdR3_0),.clk(gclk));
	jdff dff_A_IEo8tGwN3_0(.dout(w_dff_A_86b8CQdR3_0),.din(w_dff_A_IEo8tGwN3_0),.clk(gclk));
	jdff dff_A_mljz6IqM0_0(.dout(w_dff_A_IEo8tGwN3_0),.din(w_dff_A_mljz6IqM0_0),.clk(gclk));
	jdff dff_A_piDFrEPc8_0(.dout(w_dff_A_mljz6IqM0_0),.din(w_dff_A_piDFrEPc8_0),.clk(gclk));
	jdff dff_A_EitXLudL1_0(.dout(w_G4091_1[0]),.din(w_dff_A_EitXLudL1_0),.clk(gclk));
	jdff dff_A_QnZl4vUa2_0(.dout(w_dff_A_EitXLudL1_0),.din(w_dff_A_QnZl4vUa2_0),.clk(gclk));
	jdff dff_A_9Xb9cIaV5_0(.dout(w_dff_A_QnZl4vUa2_0),.din(w_dff_A_9Xb9cIaV5_0),.clk(gclk));
	jdff dff_A_0E3KASNc4_0(.dout(w_dff_A_9Xb9cIaV5_0),.din(w_dff_A_0E3KASNc4_0),.clk(gclk));
	jdff dff_A_ZZv3dkAw8_0(.dout(w_dff_A_0E3KASNc4_0),.din(w_dff_A_ZZv3dkAw8_0),.clk(gclk));
	jdff dff_A_tUwb5tTI9_0(.dout(w_dff_A_ZZv3dkAw8_0),.din(w_dff_A_tUwb5tTI9_0),.clk(gclk));
	jdff dff_A_sQwWNgac7_0(.dout(w_dff_A_tUwb5tTI9_0),.din(w_dff_A_sQwWNgac7_0),.clk(gclk));
	jdff dff_A_WS9eeEtU1_0(.dout(w_dff_A_sQwWNgac7_0),.din(w_dff_A_WS9eeEtU1_0),.clk(gclk));
	jdff dff_A_9OEWljUK9_1(.dout(w_G4091_1[1]),.din(w_dff_A_9OEWljUK9_1),.clk(gclk));
	jdff dff_A_Wo73ayXj5_1(.dout(w_dff_A_9OEWljUK9_1),.din(w_dff_A_Wo73ayXj5_1),.clk(gclk));
	jdff dff_A_9HeyBpws5_1(.dout(w_dff_A_Wo73ayXj5_1),.din(w_dff_A_9HeyBpws5_1),.clk(gclk));
	jdff dff_A_8LSCkkyj2_1(.dout(w_dff_A_9HeyBpws5_1),.din(w_dff_A_8LSCkkyj2_1),.clk(gclk));
	jdff dff_A_PIJVGkZz1_1(.dout(w_dff_A_8LSCkkyj2_1),.din(w_dff_A_PIJVGkZz1_1),.clk(gclk));
	jdff dff_A_Ss8MEqmn8_1(.dout(w_dff_A_PIJVGkZz1_1),.din(w_dff_A_Ss8MEqmn8_1),.clk(gclk));
	jdff dff_A_H1SsEM2h4_1(.dout(w_dff_A_Ss8MEqmn8_1),.din(w_dff_A_H1SsEM2h4_1),.clk(gclk));
	jdff dff_A_9MtcZvZE4_1(.dout(w_G4091_0[1]),.din(w_dff_A_9MtcZvZE4_1),.clk(gclk));
	jdff dff_A_KKuVZUuQ7_1(.dout(w_dff_A_9MtcZvZE4_1),.din(w_dff_A_KKuVZUuQ7_1),.clk(gclk));
	jdff dff_A_yQfGyEy12_1(.dout(w_dff_A_KKuVZUuQ7_1),.din(w_dff_A_yQfGyEy12_1),.clk(gclk));
	jdff dff_A_cf86T9NH3_1(.dout(w_dff_A_yQfGyEy12_1),.din(w_dff_A_cf86T9NH3_1),.clk(gclk));
	jdff dff_A_VjAtKayS5_1(.dout(w_dff_A_cf86T9NH3_1),.din(w_dff_A_VjAtKayS5_1),.clk(gclk));
	jdff dff_A_ajbuNz1y3_1(.dout(w_dff_A_VjAtKayS5_1),.din(w_dff_A_ajbuNz1y3_1),.clk(gclk));
	jdff dff_A_Szs7ReQ35_1(.dout(w_dff_A_ajbuNz1y3_1),.din(w_dff_A_Szs7ReQ35_1),.clk(gclk));
	jdff dff_A_UGiFwJl39_1(.dout(w_dff_A_Szs7ReQ35_1),.din(w_dff_A_UGiFwJl39_1),.clk(gclk));
	jdff dff_A_t3Q4ZoCk4_1(.dout(w_dff_A_UGiFwJl39_1),.din(w_dff_A_t3Q4ZoCk4_1),.clk(gclk));
	jdff dff_A_5QgE2dt85_1(.dout(w_dff_A_t3Q4ZoCk4_1),.din(w_dff_A_5QgE2dt85_1),.clk(gclk));
	jdff dff_A_2I9ItvmN3_1(.dout(w_dff_A_5QgE2dt85_1),.din(w_dff_A_2I9ItvmN3_1),.clk(gclk));
	jdff dff_A_XdZlMQAp8_1(.dout(w_dff_A_2I9ItvmN3_1),.din(w_dff_A_XdZlMQAp8_1),.clk(gclk));
	jdff dff_A_ZsiNco8d4_1(.dout(w_dff_A_XdZlMQAp8_1),.din(w_dff_A_ZsiNco8d4_1),.clk(gclk));
	jdff dff_A_sV38P4L49_2(.dout(w_G4091_0[2]),.din(w_dff_A_sV38P4L49_2),.clk(gclk));
	jdff dff_A_o1bSZhtG4_2(.dout(w_dff_A_sV38P4L49_2),.din(w_dff_A_o1bSZhtG4_2),.clk(gclk));
	jdff dff_A_RxDwcOHl8_2(.dout(w_dff_A_o1bSZhtG4_2),.din(w_dff_A_RxDwcOHl8_2),.clk(gclk));
	jdff dff_A_4GsiOF2g8_2(.dout(w_dff_A_RxDwcOHl8_2),.din(w_dff_A_4GsiOF2g8_2),.clk(gclk));
	jdff dff_A_id7i98L30_2(.dout(w_dff_A_4GsiOF2g8_2),.din(w_dff_A_id7i98L30_2),.clk(gclk));
	jdff dff_A_z11Eld5C5_2(.dout(w_dff_A_id7i98L30_2),.din(w_dff_A_z11Eld5C5_2),.clk(gclk));
	jdff dff_A_b6se461D7_2(.dout(w_dff_A_z11Eld5C5_2),.din(w_dff_A_b6se461D7_2),.clk(gclk));
	jdff dff_A_pFqduqXp0_2(.dout(w_dff_A_b6se461D7_2),.din(w_dff_A_pFqduqXp0_2),.clk(gclk));
	jdff dff_A_r7IPFdiu7_2(.dout(w_G4092_3[2]),.din(w_dff_A_r7IPFdiu7_2),.clk(gclk));
	jdff dff_A_ugPDC4sW7_2(.dout(w_dff_A_r7IPFdiu7_2),.din(w_dff_A_ugPDC4sW7_2),.clk(gclk));
	jdff dff_A_JW7ucBXq1_2(.dout(w_dff_A_ugPDC4sW7_2),.din(w_dff_A_JW7ucBXq1_2),.clk(gclk));
	jdff dff_A_orSiVrM64_2(.dout(w_dff_A_JW7ucBXq1_2),.din(w_dff_A_orSiVrM64_2),.clk(gclk));
	jdff dff_A_psOsMHOR2_2(.dout(w_dff_A_orSiVrM64_2),.din(w_dff_A_psOsMHOR2_2),.clk(gclk));
	jdff dff_A_tQ5rBqIt1_2(.dout(w_dff_A_psOsMHOR2_2),.din(w_dff_A_tQ5rBqIt1_2),.clk(gclk));
	jdff dff_A_TQCfDaYJ3_2(.dout(w_dff_A_tQ5rBqIt1_2),.din(w_dff_A_TQCfDaYJ3_2),.clk(gclk));
	jdff dff_A_WV4ki3Zp1_2(.dout(w_dff_A_TQCfDaYJ3_2),.din(w_dff_A_WV4ki3Zp1_2),.clk(gclk));
	jdff dff_A_hNALHbFE6_2(.dout(w_dff_A_WV4ki3Zp1_2),.din(w_dff_A_hNALHbFE6_2),.clk(gclk));
	jdff dff_A_YnuYCGgS8_2(.dout(w_dff_A_hNALHbFE6_2),.din(w_dff_A_YnuYCGgS8_2),.clk(gclk));
	jdff dff_A_tWgS3oAK1_2(.dout(w_dff_A_YnuYCGgS8_2),.din(w_dff_A_tWgS3oAK1_2),.clk(gclk));
	jdff dff_A_WsPtK1r61_2(.dout(w_dff_A_tWgS3oAK1_2),.din(w_dff_A_WsPtK1r61_2),.clk(gclk));
	jdff dff_A_Tvm6nn3e3_2(.dout(w_dff_A_WsPtK1r61_2),.din(w_dff_A_Tvm6nn3e3_2),.clk(gclk));
	jdff dff_A_DnTYD3nX1_2(.dout(w_dff_A_Tvm6nn3e3_2),.din(w_dff_A_DnTYD3nX1_2),.clk(gclk));
	jdff dff_A_fCJhd0fm9_2(.dout(w_dff_A_DnTYD3nX1_2),.din(w_dff_A_fCJhd0fm9_2),.clk(gclk));
	jdff dff_A_UJ2Znemh6_2(.dout(w_dff_A_fCJhd0fm9_2),.din(w_dff_A_UJ2Znemh6_2),.clk(gclk));
	jdff dff_A_Ws7c9QGw6_2(.dout(w_dff_A_UJ2Znemh6_2),.din(w_dff_A_Ws7c9QGw6_2),.clk(gclk));
	jdff dff_A_r7lXwKxe0_2(.dout(w_dff_A_Ws7c9QGw6_2),.din(w_dff_A_r7lXwKxe0_2),.clk(gclk));
	jdff dff_A_8AcuioY74_2(.dout(w_dff_A_r7lXwKxe0_2),.din(w_dff_A_8AcuioY74_2),.clk(gclk));
	jdff dff_A_4gOJRDdD0_2(.dout(w_dff_A_8AcuioY74_2),.din(w_dff_A_4gOJRDdD0_2),.clk(gclk));
	jdff dff_A_QPoL2Yr86_1(.dout(w_G4092_0[1]),.din(w_dff_A_QPoL2Yr86_1),.clk(gclk));
	jdff dff_A_WSqycTFI7_0(.dout(w_n1008_4[0]),.din(w_dff_A_WSqycTFI7_0),.clk(gclk));
	jdff dff_A_uUSEqkrO9_0(.dout(w_dff_A_WSqycTFI7_0),.din(w_dff_A_uUSEqkrO9_0),.clk(gclk));
	jdff dff_A_ON0sg6aB4_0(.dout(w_dff_A_uUSEqkrO9_0),.din(w_dff_A_ON0sg6aB4_0),.clk(gclk));
	jdff dff_A_4uUDOd8n9_0(.dout(w_dff_A_ON0sg6aB4_0),.din(w_dff_A_4uUDOd8n9_0),.clk(gclk));
	jdff dff_A_ok1mW5CE9_0(.dout(w_dff_A_4uUDOd8n9_0),.din(w_dff_A_ok1mW5CE9_0),.clk(gclk));
	jdff dff_A_Qx3w1VQI2_0(.dout(w_dff_A_ok1mW5CE9_0),.din(w_dff_A_Qx3w1VQI2_0),.clk(gclk));
	jdff dff_A_8f1KVLOG8_0(.dout(w_dff_A_Qx3w1VQI2_0),.din(w_dff_A_8f1KVLOG8_0),.clk(gclk));
	jdff dff_A_SMf7Agkr3_0(.dout(w_dff_A_8f1KVLOG8_0),.din(w_dff_A_SMf7Agkr3_0),.clk(gclk));
	jdff dff_A_n88UjXSt9_0(.dout(w_dff_A_SMf7Agkr3_0),.din(w_dff_A_n88UjXSt9_0),.clk(gclk));
	jdff dff_A_4EMrDtKz7_0(.dout(w_dff_A_n88UjXSt9_0),.din(w_dff_A_4EMrDtKz7_0),.clk(gclk));
	jdff dff_A_2ZojMmEh2_0(.dout(w_dff_A_4EMrDtKz7_0),.din(w_dff_A_2ZojMmEh2_0),.clk(gclk));
	jdff dff_A_OYIlsWXH8_0(.dout(w_dff_A_2ZojMmEh2_0),.din(w_dff_A_OYIlsWXH8_0),.clk(gclk));
	jdff dff_A_qFgT65Bj9_0(.dout(w_dff_A_OYIlsWXH8_0),.din(w_dff_A_qFgT65Bj9_0),.clk(gclk));
	jdff dff_A_XCvCTKxb7_0(.dout(w_dff_A_qFgT65Bj9_0),.din(w_dff_A_XCvCTKxb7_0),.clk(gclk));
	jdff dff_A_SKWies1N4_0(.dout(w_dff_A_XCvCTKxb7_0),.din(w_dff_A_SKWies1N4_0),.clk(gclk));
	jdff dff_A_u3Idcy3m6_2(.dout(w_n1008_4[2]),.din(w_dff_A_u3Idcy3m6_2),.clk(gclk));
	jdff dff_A_LA10yz5M3_2(.dout(w_dff_A_u3Idcy3m6_2),.din(w_dff_A_LA10yz5M3_2),.clk(gclk));
	jdff dff_A_TlxeCcEY4_2(.dout(w_dff_A_LA10yz5M3_2),.din(w_dff_A_TlxeCcEY4_2),.clk(gclk));
	jdff dff_A_QQO0Bdfn3_2(.dout(w_dff_A_TlxeCcEY4_2),.din(w_dff_A_QQO0Bdfn3_2),.clk(gclk));
	jdff dff_A_bSPJPTBF8_2(.dout(w_dff_A_QQO0Bdfn3_2),.din(w_dff_A_bSPJPTBF8_2),.clk(gclk));
	jdff dff_A_EGyJJntq3_2(.dout(w_dff_A_bSPJPTBF8_2),.din(w_dff_A_EGyJJntq3_2),.clk(gclk));
	jdff dff_A_D5C9xmcl9_2(.dout(w_dff_A_EGyJJntq3_2),.din(w_dff_A_D5C9xmcl9_2),.clk(gclk));
	jdff dff_A_OQJO4pMg6_2(.dout(w_dff_A_D5C9xmcl9_2),.din(w_dff_A_OQJO4pMg6_2),.clk(gclk));
	jdff dff_A_zcNQ3ys02_2(.dout(w_dff_A_OQJO4pMg6_2),.din(w_dff_A_zcNQ3ys02_2),.clk(gclk));
	jdff dff_A_mZ86McBp3_2(.dout(w_dff_A_zcNQ3ys02_2),.din(w_dff_A_mZ86McBp3_2),.clk(gclk));
	jdff dff_A_kSfNaV7k4_1(.dout(w_n1008_1[1]),.din(w_dff_A_kSfNaV7k4_1),.clk(gclk));
	jdff dff_A_XCW97tO20_1(.dout(w_dff_A_kSfNaV7k4_1),.din(w_dff_A_XCW97tO20_1),.clk(gclk));
	jdff dff_A_dsynUTGi1_1(.dout(w_dff_A_XCW97tO20_1),.din(w_dff_A_dsynUTGi1_1),.clk(gclk));
	jdff dff_A_oLJktYkX3_1(.dout(w_dff_A_dsynUTGi1_1),.din(w_dff_A_oLJktYkX3_1),.clk(gclk));
	jdff dff_A_OhuHp5ts4_1(.dout(w_dff_A_oLJktYkX3_1),.din(w_dff_A_OhuHp5ts4_1),.clk(gclk));
	jdff dff_A_dnfSHvyF5_1(.dout(w_dff_A_OhuHp5ts4_1),.din(w_dff_A_dnfSHvyF5_1),.clk(gclk));
	jdff dff_A_Bh0PukLk2_1(.dout(w_dff_A_dnfSHvyF5_1),.din(w_dff_A_Bh0PukLk2_1),.clk(gclk));
	jdff dff_A_Q7GQe5kG7_1(.dout(w_dff_A_Bh0PukLk2_1),.din(w_dff_A_Q7GQe5kG7_1),.clk(gclk));
	jdff dff_A_VJp9CNGQ7_1(.dout(w_dff_A_Q7GQe5kG7_1),.din(w_dff_A_VJp9CNGQ7_1),.clk(gclk));
	jdff dff_A_Npfoxvkr2_1(.dout(w_dff_A_VJp9CNGQ7_1),.din(w_dff_A_Npfoxvkr2_1),.clk(gclk));
	jdff dff_A_RRf0z1JV7_1(.dout(w_dff_A_Npfoxvkr2_1),.din(w_dff_A_RRf0z1JV7_1),.clk(gclk));
	jdff dff_A_0LDNOHWG8_1(.dout(w_dff_A_RRf0z1JV7_1),.din(w_dff_A_0LDNOHWG8_1),.clk(gclk));
	jdff dff_A_pjQgGHN08_1(.dout(w_dff_A_0LDNOHWG8_1),.din(w_dff_A_pjQgGHN08_1),.clk(gclk));
	jdff dff_A_XJr2CE7J8_1(.dout(w_dff_A_pjQgGHN08_1),.din(w_dff_A_XJr2CE7J8_1),.clk(gclk));
	jdff dff_A_wayGqTb63_1(.dout(w_dff_A_XJr2CE7J8_1),.din(w_dff_A_wayGqTb63_1),.clk(gclk));
	jdff dff_A_DYHgFZ441_1(.dout(w_dff_A_wayGqTb63_1),.din(w_dff_A_DYHgFZ441_1),.clk(gclk));
	jdff dff_A_52KHvoTS2_1(.dout(w_dff_A_DYHgFZ441_1),.din(w_dff_A_52KHvoTS2_1),.clk(gclk));
	jdff dff_A_WR26FZwb7_1(.dout(w_dff_A_52KHvoTS2_1),.din(w_dff_A_WR26FZwb7_1),.clk(gclk));
	jdff dff_A_xftwfBFJ9_1(.dout(w_dff_A_WR26FZwb7_1),.din(w_dff_A_xftwfBFJ9_1),.clk(gclk));
	jdff dff_A_QDnQbt1F5_1(.dout(w_dff_A_xftwfBFJ9_1),.din(w_dff_A_QDnQbt1F5_1),.clk(gclk));
	jdff dff_A_pQ3HAkyF6_1(.dout(w_dff_A_QDnQbt1F5_1),.din(w_dff_A_pQ3HAkyF6_1),.clk(gclk));
	jdff dff_A_SIxGBBAz0_2(.dout(w_n1008_1[2]),.din(w_dff_A_SIxGBBAz0_2),.clk(gclk));
	jdff dff_A_oR8Ojy7Q8_2(.dout(w_dff_A_SIxGBBAz0_2),.din(w_dff_A_oR8Ojy7Q8_2),.clk(gclk));
	jdff dff_A_Fs10dkLd6_2(.dout(w_dff_A_oR8Ojy7Q8_2),.din(w_dff_A_Fs10dkLd6_2),.clk(gclk));
	jdff dff_A_pO8CWy865_2(.dout(w_dff_A_Fs10dkLd6_2),.din(w_dff_A_pO8CWy865_2),.clk(gclk));
	jdff dff_A_mP8DDIcz7_2(.dout(w_dff_A_pO8CWy865_2),.din(w_dff_A_mP8DDIcz7_2),.clk(gclk));
	jdff dff_A_rdAFcOJ67_2(.dout(w_dff_A_mP8DDIcz7_2),.din(w_dff_A_rdAFcOJ67_2),.clk(gclk));
	jdff dff_A_sTvDPdlT3_2(.dout(w_dff_A_rdAFcOJ67_2),.din(w_dff_A_sTvDPdlT3_2),.clk(gclk));
	jdff dff_A_bHA0pX3V9_2(.dout(w_dff_A_sTvDPdlT3_2),.din(w_dff_A_bHA0pX3V9_2),.clk(gclk));
	jdff dff_A_ZxqKzhHM7_2(.dout(w_dff_A_bHA0pX3V9_2),.din(w_dff_A_ZxqKzhHM7_2),.clk(gclk));
	jdff dff_A_5LGF4Llh5_2(.dout(w_dff_A_ZxqKzhHM7_2),.din(w_dff_A_5LGF4Llh5_2),.clk(gclk));
	jdff dff_A_YuYIoP734_2(.dout(w_dff_A_5LGF4Llh5_2),.din(w_dff_A_YuYIoP734_2),.clk(gclk));
	jdff dff_A_RMrA0vc58_2(.dout(w_dff_A_YuYIoP734_2),.din(w_dff_A_RMrA0vc58_2),.clk(gclk));
	jdff dff_A_1DDlXiSl7_2(.dout(w_dff_A_RMrA0vc58_2),.din(w_dff_A_1DDlXiSl7_2),.clk(gclk));
	jdff dff_A_A0wXchy67_2(.dout(w_dff_A_1DDlXiSl7_2),.din(w_dff_A_A0wXchy67_2),.clk(gclk));
	jdff dff_A_axxn571j7_2(.dout(w_dff_A_A0wXchy67_2),.din(w_dff_A_axxn571j7_2),.clk(gclk));
	jdff dff_A_fizGF83e2_2(.dout(w_dff_A_axxn571j7_2),.din(w_dff_A_fizGF83e2_2),.clk(gclk));
	jdff dff_A_7exSQ6oc8_2(.dout(w_dff_A_fizGF83e2_2),.din(w_dff_A_7exSQ6oc8_2),.clk(gclk));
	jdff dff_A_Klt8O5nc0_2(.dout(w_dff_A_7exSQ6oc8_2),.din(w_dff_A_Klt8O5nc0_2),.clk(gclk));
	jdff dff_A_AwGANxKm8_2(.dout(w_dff_A_Klt8O5nc0_2),.din(w_dff_A_AwGANxKm8_2),.clk(gclk));
	jdff dff_A_SwhyDRds8_2(.dout(w_dff_A_AwGANxKm8_2),.din(w_dff_A_SwhyDRds8_2),.clk(gclk));
	jdff dff_A_joNpa7pj5_1(.dout(w_n1008_0[1]),.din(w_dff_A_joNpa7pj5_1),.clk(gclk));
	jdff dff_A_IwgFjkYh3_1(.dout(w_dff_A_joNpa7pj5_1),.din(w_dff_A_IwgFjkYh3_1),.clk(gclk));
	jdff dff_A_KLZFKEtw2_1(.dout(w_dff_A_IwgFjkYh3_1),.din(w_dff_A_KLZFKEtw2_1),.clk(gclk));
	jdff dff_A_7FxgQzyS8_1(.dout(w_dff_A_KLZFKEtw2_1),.din(w_dff_A_7FxgQzyS8_1),.clk(gclk));
	jdff dff_A_mKKPOxLH8_1(.dout(w_dff_A_7FxgQzyS8_1),.din(w_dff_A_mKKPOxLH8_1),.clk(gclk));
	jdff dff_A_eFGPnXsz7_1(.dout(w_dff_A_mKKPOxLH8_1),.din(w_dff_A_eFGPnXsz7_1),.clk(gclk));
	jdff dff_A_EHMk3NIn7_1(.dout(w_dff_A_eFGPnXsz7_1),.din(w_dff_A_EHMk3NIn7_1),.clk(gclk));
	jdff dff_A_NklZwVqI4_1(.dout(w_dff_A_EHMk3NIn7_1),.din(w_dff_A_NklZwVqI4_1),.clk(gclk));
	jdff dff_A_Sv95TVcw6_1(.dout(w_dff_A_NklZwVqI4_1),.din(w_dff_A_Sv95TVcw6_1),.clk(gclk));
	jdff dff_A_PKwUAUwU8_1(.dout(w_dff_A_Sv95TVcw6_1),.din(w_dff_A_PKwUAUwU8_1),.clk(gclk));
	jdff dff_A_oUP31tfa2_1(.dout(w_dff_A_PKwUAUwU8_1),.din(w_dff_A_oUP31tfa2_1),.clk(gclk));
	jdff dff_A_MVYqPbwh5_1(.dout(w_dff_A_oUP31tfa2_1),.din(w_dff_A_MVYqPbwh5_1),.clk(gclk));
	jdff dff_A_CRBbVg4z5_1(.dout(w_dff_A_MVYqPbwh5_1),.din(w_dff_A_CRBbVg4z5_1),.clk(gclk));
	jdff dff_A_8BtsdIM15_1(.dout(w_dff_A_CRBbVg4z5_1),.din(w_dff_A_8BtsdIM15_1),.clk(gclk));
	jdff dff_A_vH45RwE30_1(.dout(w_dff_A_8BtsdIM15_1),.din(w_dff_A_vH45RwE30_1),.clk(gclk));
	jdff dff_A_CBJv59lI3_1(.dout(w_dff_A_vH45RwE30_1),.din(w_dff_A_CBJv59lI3_1),.clk(gclk));
	jdff dff_A_fDL2Gcz20_1(.dout(w_dff_A_CBJv59lI3_1),.din(w_dff_A_fDL2Gcz20_1),.clk(gclk));
	jdff dff_A_b1Z1GqIh7_1(.dout(w_dff_A_fDL2Gcz20_1),.din(w_dff_A_b1Z1GqIh7_1),.clk(gclk));
	jdff dff_A_gZloFhOf3_2(.dout(w_n1008_0[2]),.din(w_dff_A_gZloFhOf3_2),.clk(gclk));
	jdff dff_A_Lu9EV3RW3_2(.dout(w_dff_A_gZloFhOf3_2),.din(w_dff_A_Lu9EV3RW3_2),.clk(gclk));
	jdff dff_A_jNxfeHUK6_2(.dout(w_dff_A_Lu9EV3RW3_2),.din(w_dff_A_jNxfeHUK6_2),.clk(gclk));
	jdff dff_A_CDcBIiOV7_2(.dout(w_dff_A_jNxfeHUK6_2),.din(w_dff_A_CDcBIiOV7_2),.clk(gclk));
	jdff dff_A_HW3Sb6ig8_2(.dout(w_dff_A_CDcBIiOV7_2),.din(w_dff_A_HW3Sb6ig8_2),.clk(gclk));
	jdff dff_A_C9YfbesS1_2(.dout(w_dff_A_HW3Sb6ig8_2),.din(w_dff_A_C9YfbesS1_2),.clk(gclk));
	jdff dff_A_pyMCgMEp8_2(.dout(w_dff_A_C9YfbesS1_2),.din(w_dff_A_pyMCgMEp8_2),.clk(gclk));
	jdff dff_A_da5ylVH45_2(.dout(w_dff_A_pyMCgMEp8_2),.din(w_dff_A_da5ylVH45_2),.clk(gclk));
	jdff dff_A_9BWh89Fn8_2(.dout(w_dff_A_da5ylVH45_2),.din(w_dff_A_9BWh89Fn8_2),.clk(gclk));
	jdff dff_A_PoY3Yy488_2(.dout(w_dff_A_9BWh89Fn8_2),.din(w_dff_A_PoY3Yy488_2),.clk(gclk));
	jdff dff_A_wtsjZLC43_2(.dout(w_dff_A_PoY3Yy488_2),.din(w_dff_A_wtsjZLC43_2),.clk(gclk));
	jdff dff_A_lvhsygkr0_1(.dout(w_G1691_5[1]),.din(w_dff_A_lvhsygkr0_1),.clk(gclk));
	jdff dff_A_nGbJspLH0_1(.dout(w_dff_A_lvhsygkr0_1),.din(w_dff_A_nGbJspLH0_1),.clk(gclk));
	jdff dff_A_zMCP0Xa69_1(.dout(w_dff_A_nGbJspLH0_1),.din(w_dff_A_zMCP0Xa69_1),.clk(gclk));
	jdff dff_A_Mtb30mf10_1(.dout(w_dff_A_zMCP0Xa69_1),.din(w_dff_A_Mtb30mf10_1),.clk(gclk));
	jdff dff_A_7z7cGEbk7_1(.dout(w_dff_A_Mtb30mf10_1),.din(w_dff_A_7z7cGEbk7_1),.clk(gclk));
	jdff dff_A_LLipclX71_1(.dout(w_dff_A_7z7cGEbk7_1),.din(w_dff_A_LLipclX71_1),.clk(gclk));
	jdff dff_A_sXUPwNmt9_1(.dout(w_dff_A_LLipclX71_1),.din(w_dff_A_sXUPwNmt9_1),.clk(gclk));
	jdff dff_A_GUx2y2KX8_1(.dout(w_dff_A_sXUPwNmt9_1),.din(w_dff_A_GUx2y2KX8_1),.clk(gclk));
	jdff dff_A_KCA2LkGM5_1(.dout(w_dff_A_GUx2y2KX8_1),.din(w_dff_A_KCA2LkGM5_1),.clk(gclk));
	jdff dff_B_JFNhjRj26_2(.din(n1698),.dout(w_dff_B_JFNhjRj26_2),.clk(gclk));
	jdff dff_B_SHjTvCFN8_2(.din(w_dff_B_JFNhjRj26_2),.dout(w_dff_B_SHjTvCFN8_2),.clk(gclk));
	jdff dff_A_NrHeVJaU2_1(.dout(w_G1694_0[1]),.din(w_dff_A_NrHeVJaU2_1),.clk(gclk));
	jdff dff_A_OYuBxBoI3_1(.dout(w_dff_A_NrHeVJaU2_1),.din(w_dff_A_OYuBxBoI3_1),.clk(gclk));
	jdff dff_A_83w313hf4_1(.dout(w_dff_A_OYuBxBoI3_1),.din(w_dff_A_83w313hf4_1),.clk(gclk));
	jdff dff_A_uq3IpMya7_1(.dout(w_dff_A_83w313hf4_1),.din(w_dff_A_uq3IpMya7_1),.clk(gclk));
	jdff dff_A_PndnQEq71_1(.dout(w_dff_A_uq3IpMya7_1),.din(w_dff_A_PndnQEq71_1),.clk(gclk));
	jdff dff_A_tt66UUE16_1(.dout(w_dff_A_PndnQEq71_1),.din(w_dff_A_tt66UUE16_1),.clk(gclk));
	jdff dff_A_MkNfVwnp9_1(.dout(w_dff_A_tt66UUE16_1),.din(w_dff_A_MkNfVwnp9_1),.clk(gclk));
	jdff dff_A_6CU7N1Vx3_1(.dout(w_dff_A_MkNfVwnp9_1),.din(w_dff_A_6CU7N1Vx3_1),.clk(gclk));
	jdff dff_A_HL2V6y215_1(.dout(w_dff_A_6CU7N1Vx3_1),.din(w_dff_A_HL2V6y215_1),.clk(gclk));
	jdff dff_A_MgmqeuPb5_1(.dout(w_dff_A_HL2V6y215_1),.din(w_dff_A_MgmqeuPb5_1),.clk(gclk));
	jdff dff_A_R894gWeW2_1(.dout(w_dff_A_MgmqeuPb5_1),.din(w_dff_A_R894gWeW2_1),.clk(gclk));
	jdff dff_A_xVXb5A5Y1_1(.dout(w_dff_A_R894gWeW2_1),.din(w_dff_A_xVXb5A5Y1_1),.clk(gclk));
	jdff dff_A_bvIW5vGo3_1(.dout(w_dff_A_xVXb5A5Y1_1),.din(w_dff_A_bvIW5vGo3_1),.clk(gclk));
	jdff dff_A_aHrjlshB3_1(.dout(w_dff_A_bvIW5vGo3_1),.din(w_dff_A_aHrjlshB3_1),.clk(gclk));
	jdff dff_A_n8pSpgXP7_1(.dout(w_dff_A_aHrjlshB3_1),.din(w_dff_A_n8pSpgXP7_1),.clk(gclk));
	jdff dff_A_WI9PiHta0_1(.dout(w_dff_A_n8pSpgXP7_1),.din(w_dff_A_WI9PiHta0_1),.clk(gclk));
	jdff dff_A_K8lD1TQj4_1(.dout(w_dff_A_WI9PiHta0_1),.din(w_dff_A_K8lD1TQj4_1),.clk(gclk));
	jdff dff_A_LbbRRbec4_1(.dout(w_dff_A_K8lD1TQj4_1),.din(w_dff_A_LbbRRbec4_1),.clk(gclk));
	jdff dff_A_veYxSZ2n8_1(.dout(w_dff_A_LbbRRbec4_1),.din(w_dff_A_veYxSZ2n8_1),.clk(gclk));
	jdff dff_A_IR6oyroZ0_1(.dout(w_dff_A_veYxSZ2n8_1),.din(w_dff_A_IR6oyroZ0_1),.clk(gclk));
	jdff dff_A_o6R8sHul4_1(.dout(w_dff_A_IR6oyroZ0_1),.din(w_dff_A_o6R8sHul4_1),.clk(gclk));
	jdff dff_A_rm69yGQw1_1(.dout(w_dff_A_o6R8sHul4_1),.din(w_dff_A_rm69yGQw1_1),.clk(gclk));
	jdff dff_A_PuJrd79y3_1(.dout(w_dff_A_rm69yGQw1_1),.din(w_dff_A_PuJrd79y3_1),.clk(gclk));
	jdff dff_A_dgGMwTgw5_2(.dout(w_G1694_0[2]),.din(w_dff_A_dgGMwTgw5_2),.clk(gclk));
	jdff dff_A_jez6q3ck6_0(.dout(w_G1691_4[0]),.din(w_dff_A_jez6q3ck6_0),.clk(gclk));
	jdff dff_A_Y5Htbw501_0(.dout(w_dff_A_jez6q3ck6_0),.din(w_dff_A_Y5Htbw501_0),.clk(gclk));
	jdff dff_A_y1XNu93O5_0(.dout(w_dff_A_Y5Htbw501_0),.din(w_dff_A_y1XNu93O5_0),.clk(gclk));
	jdff dff_A_nuFK7bXb4_0(.dout(w_dff_A_y1XNu93O5_0),.din(w_dff_A_nuFK7bXb4_0),.clk(gclk));
	jdff dff_A_EupK70Ep0_0(.dout(w_dff_A_nuFK7bXb4_0),.din(w_dff_A_EupK70Ep0_0),.clk(gclk));
	jdff dff_A_lFRbiMll2_0(.dout(w_dff_A_EupK70Ep0_0),.din(w_dff_A_lFRbiMll2_0),.clk(gclk));
	jdff dff_A_rffl1DUk7_0(.dout(w_dff_A_lFRbiMll2_0),.din(w_dff_A_rffl1DUk7_0),.clk(gclk));
	jdff dff_A_jg5l5pMu3_0(.dout(w_dff_A_rffl1DUk7_0),.din(w_dff_A_jg5l5pMu3_0),.clk(gclk));
	jdff dff_A_uU8WhNG28_0(.dout(w_dff_A_jg5l5pMu3_0),.din(w_dff_A_uU8WhNG28_0),.clk(gclk));
	jdff dff_A_hKfi0Hnm4_0(.dout(w_dff_A_uU8WhNG28_0),.din(w_dff_A_hKfi0Hnm4_0),.clk(gclk));
	jdff dff_A_lmAqRxtF5_0(.dout(w_dff_A_hKfi0Hnm4_0),.din(w_dff_A_lmAqRxtF5_0),.clk(gclk));
	jdff dff_A_nGpldJDP8_0(.dout(w_dff_A_lmAqRxtF5_0),.din(w_dff_A_nGpldJDP8_0),.clk(gclk));
	jdff dff_A_OSok7hQx6_0(.dout(w_dff_A_nGpldJDP8_0),.din(w_dff_A_OSok7hQx6_0),.clk(gclk));
	jdff dff_A_eNq6EuQo6_0(.dout(w_dff_A_OSok7hQx6_0),.din(w_dff_A_eNq6EuQo6_0),.clk(gclk));
	jdff dff_A_ZJRvuEij9_1(.dout(w_G1691_4[1]),.din(w_dff_A_ZJRvuEij9_1),.clk(gclk));
	jdff dff_A_DPFh9Ds93_1(.dout(w_dff_A_ZJRvuEij9_1),.din(w_dff_A_DPFh9Ds93_1),.clk(gclk));
	jdff dff_A_cnEbxqi33_1(.dout(w_dff_A_DPFh9Ds93_1),.din(w_dff_A_cnEbxqi33_1),.clk(gclk));
	jdff dff_A_wKY5CZ829_1(.dout(w_dff_A_cnEbxqi33_1),.din(w_dff_A_wKY5CZ829_1),.clk(gclk));
	jdff dff_A_tSDqsGMI2_1(.dout(w_dff_A_wKY5CZ829_1),.din(w_dff_A_tSDqsGMI2_1),.clk(gclk));
	jdff dff_A_fgD7Vqk01_1(.dout(w_dff_A_tSDqsGMI2_1),.din(w_dff_A_fgD7Vqk01_1),.clk(gclk));
	jdff dff_A_eqb7eVTU8_1(.dout(w_dff_A_fgD7Vqk01_1),.din(w_dff_A_eqb7eVTU8_1),.clk(gclk));
	jdff dff_A_6WBwahvX6_1(.dout(w_dff_A_eqb7eVTU8_1),.din(w_dff_A_6WBwahvX6_1),.clk(gclk));
	jdff dff_A_nDzZ8UwB1_1(.dout(w_dff_A_6WBwahvX6_1),.din(w_dff_A_nDzZ8UwB1_1),.clk(gclk));
	jdff dff_A_51fD4GFb3_1(.dout(w_dff_A_nDzZ8UwB1_1),.din(w_dff_A_51fD4GFb3_1),.clk(gclk));
	jdff dff_A_MORzu4mx0_1(.dout(w_dff_A_51fD4GFb3_1),.din(w_dff_A_MORzu4mx0_1),.clk(gclk));
	jdff dff_A_9MzmqfIV6_1(.dout(w_dff_A_MORzu4mx0_1),.din(w_dff_A_9MzmqfIV6_1),.clk(gclk));
	jdff dff_A_6UCJrQ7E3_1(.dout(w_dff_A_9MzmqfIV6_1),.din(w_dff_A_6UCJrQ7E3_1),.clk(gclk));
	jdff dff_A_c1qCztz99_1(.dout(w_dff_A_6UCJrQ7E3_1),.din(w_dff_A_c1qCztz99_1),.clk(gclk));
	jdff dff_A_Al4YqERy7_1(.dout(w_dff_A_c1qCztz99_1),.din(w_dff_A_Al4YqERy7_1),.clk(gclk));
	jdff dff_A_XLZ3R2fU3_1(.dout(w_dff_A_Al4YqERy7_1),.din(w_dff_A_XLZ3R2fU3_1),.clk(gclk));
	jdff dff_A_ZtOT0hLB6_2(.dout(w_G1691_1[2]),.din(w_dff_A_ZtOT0hLB6_2),.clk(gclk));
	jdff dff_A_pel3Qd872_2(.dout(w_dff_A_ZtOT0hLB6_2),.din(w_dff_A_pel3Qd872_2),.clk(gclk));
	jdff dff_A_bqdsjcwZ5_2(.dout(w_dff_A_pel3Qd872_2),.din(w_dff_A_bqdsjcwZ5_2),.clk(gclk));
	jdff dff_A_RF67uqnd0_2(.dout(w_dff_A_bqdsjcwZ5_2),.din(w_dff_A_RF67uqnd0_2),.clk(gclk));
	jdff dff_A_sLk00SdQ3_2(.dout(w_dff_A_RF67uqnd0_2),.din(w_dff_A_sLk00SdQ3_2),.clk(gclk));
	jdff dff_A_oTAhzqlh9_2(.dout(w_dff_A_sLk00SdQ3_2),.din(w_dff_A_oTAhzqlh9_2),.clk(gclk));
	jdff dff_A_5DeqOacz4_2(.dout(w_dff_A_oTAhzqlh9_2),.din(w_dff_A_5DeqOacz4_2),.clk(gclk));
	jdff dff_A_ApLMwgYC1_2(.dout(w_dff_A_5DeqOacz4_2),.din(w_dff_A_ApLMwgYC1_2),.clk(gclk));
	jdff dff_A_r9sl2ikc0_2(.dout(w_dff_A_ApLMwgYC1_2),.din(w_dff_A_r9sl2ikc0_2),.clk(gclk));
	jdff dff_A_tnokxD7K6_2(.dout(w_dff_A_r9sl2ikc0_2),.din(w_dff_A_tnokxD7K6_2),.clk(gclk));
	jdff dff_A_PKYjso3T5_2(.dout(w_dff_A_tnokxD7K6_2),.din(w_dff_A_PKYjso3T5_2),.clk(gclk));
	jdff dff_A_aETqB8B26_2(.dout(w_dff_A_PKYjso3T5_2),.din(w_dff_A_aETqB8B26_2),.clk(gclk));
	jdff dff_A_XFia1uVj0_2(.dout(w_dff_A_aETqB8B26_2),.din(w_dff_A_XFia1uVj0_2),.clk(gclk));
	jdff dff_A_e2Ael8mC2_2(.dout(w_dff_A_XFia1uVj0_2),.din(w_dff_A_e2Ael8mC2_2),.clk(gclk));
	jdff dff_A_WtGp5k6j4_2(.dout(w_dff_A_e2Ael8mC2_2),.din(w_dff_A_WtGp5k6j4_2),.clk(gclk));
	jdff dff_A_NibZ94Xm9_2(.dout(w_dff_A_WtGp5k6j4_2),.din(w_dff_A_NibZ94Xm9_2),.clk(gclk));
	jdff dff_A_iq4YHuwO1_2(.dout(w_dff_A_NibZ94Xm9_2),.din(w_dff_A_iq4YHuwO1_2),.clk(gclk));
	jdff dff_A_GcuuUpUv0_2(.dout(w_dff_A_iq4YHuwO1_2),.din(w_dff_A_GcuuUpUv0_2),.clk(gclk));
	jdff dff_A_lnW7Jwxq5_2(.dout(w_dff_A_GcuuUpUv0_2),.din(w_dff_A_lnW7Jwxq5_2),.clk(gclk));
	jdff dff_A_bf8uZ9ug9_2(.dout(w_dff_A_lnW7Jwxq5_2),.din(w_dff_A_bf8uZ9ug9_2),.clk(gclk));
	jdff dff_A_nfyhVbYY1_2(.dout(w_dff_A_bf8uZ9ug9_2),.din(w_dff_A_nfyhVbYY1_2),.clk(gclk));
	jdff dff_A_DEUdClEX8_2(.dout(w_dff_A_nfyhVbYY1_2),.din(w_dff_A_DEUdClEX8_2),.clk(gclk));
	jdff dff_A_uOHIpPs64_1(.dout(w_G1691_0[1]),.din(w_dff_A_uOHIpPs64_1),.clk(gclk));
	jdff dff_A_Pe0dDGyj5_1(.dout(w_dff_A_uOHIpPs64_1),.din(w_dff_A_Pe0dDGyj5_1),.clk(gclk));
	jdff dff_A_RAB56aaU4_1(.dout(w_dff_A_Pe0dDGyj5_1),.din(w_dff_A_RAB56aaU4_1),.clk(gclk));
	jdff dff_A_HUKCjav54_1(.dout(w_dff_A_RAB56aaU4_1),.din(w_dff_A_HUKCjav54_1),.clk(gclk));
	jdff dff_A_Rb6g0GMP0_1(.dout(w_dff_A_HUKCjav54_1),.din(w_dff_A_Rb6g0GMP0_1),.clk(gclk));
	jdff dff_A_UOAqTRwi0_1(.dout(w_dff_A_Rb6g0GMP0_1),.din(w_dff_A_UOAqTRwi0_1),.clk(gclk));
	jdff dff_A_RqlN2u1v4_1(.dout(w_dff_A_UOAqTRwi0_1),.din(w_dff_A_RqlN2u1v4_1),.clk(gclk));
	jdff dff_A_05hehML31_1(.dout(w_dff_A_RqlN2u1v4_1),.din(w_dff_A_05hehML31_1),.clk(gclk));
	jdff dff_A_IjBL1HG98_1(.dout(w_dff_A_05hehML31_1),.din(w_dff_A_IjBL1HG98_1),.clk(gclk));
	jdff dff_A_lboOwYLZ3_1(.dout(w_dff_A_IjBL1HG98_1),.din(w_dff_A_lboOwYLZ3_1),.clk(gclk));
	jdff dff_A_qlbNgzLd4_1(.dout(w_dff_A_lboOwYLZ3_1),.din(w_dff_A_qlbNgzLd4_1),.clk(gclk));
	jdff dff_A_ivzypPC02_1(.dout(w_dff_A_qlbNgzLd4_1),.din(w_dff_A_ivzypPC02_1),.clk(gclk));
	jdff dff_A_glX40HsQ0_1(.dout(w_dff_A_ivzypPC02_1),.din(w_dff_A_glX40HsQ0_1),.clk(gclk));
	jdff dff_A_MBUqYFrl2_1(.dout(w_dff_A_glX40HsQ0_1),.din(w_dff_A_MBUqYFrl2_1),.clk(gclk));
	jdff dff_A_wbaxU3AM2_1(.dout(w_dff_A_MBUqYFrl2_1),.din(w_dff_A_wbaxU3AM2_1),.clk(gclk));
	jdff dff_A_xAhcRo9w8_1(.dout(w_dff_A_wbaxU3AM2_1),.din(w_dff_A_xAhcRo9w8_1),.clk(gclk));
	jdff dff_A_RX3Z8UeR4_1(.dout(w_dff_A_xAhcRo9w8_1),.din(w_dff_A_RX3Z8UeR4_1),.clk(gclk));
	jdff dff_A_KJeWS4oe5_1(.dout(w_dff_A_RX3Z8UeR4_1),.din(w_dff_A_KJeWS4oe5_1),.clk(gclk));
	jdff dff_A_6aehFRuv9_1(.dout(w_dff_A_KJeWS4oe5_1),.din(w_dff_A_6aehFRuv9_1),.clk(gclk));
	jdff dff_A_dMd4Dplq1_2(.dout(w_G1691_0[2]),.din(w_dff_A_dMd4Dplq1_2),.clk(gclk));
	jdff dff_A_4GLrp35o8_2(.dout(w_dff_A_dMd4Dplq1_2),.din(w_dff_A_4GLrp35o8_2),.clk(gclk));
	jdff dff_A_WuFYFDj19_2(.dout(w_dff_A_4GLrp35o8_2),.din(w_dff_A_WuFYFDj19_2),.clk(gclk));
	jdff dff_A_5zI5gduW9_2(.dout(w_dff_A_WuFYFDj19_2),.din(w_dff_A_5zI5gduW9_2),.clk(gclk));
	jdff dff_A_JcBH96rA1_2(.dout(w_dff_A_5zI5gduW9_2),.din(w_dff_A_JcBH96rA1_2),.clk(gclk));
	jdff dff_A_RwUuL03E9_2(.dout(w_dff_A_JcBH96rA1_2),.din(w_dff_A_RwUuL03E9_2),.clk(gclk));
	jdff dff_A_qSKoB0l20_2(.dout(w_dff_A_RwUuL03E9_2),.din(w_dff_A_qSKoB0l20_2),.clk(gclk));
	jdff dff_A_JzZxz98o0_2(.dout(w_dff_A_qSKoB0l20_2),.din(w_dff_A_JzZxz98o0_2),.clk(gclk));
	jdff dff_A_KFrZBu1F1_2(.dout(w_dff_A_JzZxz98o0_2),.din(w_dff_A_KFrZBu1F1_2),.clk(gclk));
	jdff dff_A_0RcGyH1M4_2(.dout(w_dff_A_KFrZBu1F1_2),.din(w_dff_A_0RcGyH1M4_2),.clk(gclk));
	jdff dff_A_klkUp8ao9_2(.dout(w_dff_A_0RcGyH1M4_2),.din(w_dff_A_klkUp8ao9_2),.clk(gclk));
	jdff dff_A_dT8Ia2OZ0_2(.dout(w_dff_A_klkUp8ao9_2),.din(w_dff_A_dT8Ia2OZ0_2),.clk(gclk));
	jdff dff_A_vGHTfhyW9_2(.dout(w_dff_A_dT8Ia2OZ0_2),.din(w_dff_A_vGHTfhyW9_2),.clk(gclk));
	jdff dff_B_AzGMDA8y8_2(.din(n1695),.dout(w_dff_B_AzGMDA8y8_2),.clk(gclk));
	jdff dff_B_uy03LviU8_2(.din(n1694),.dout(w_dff_B_uy03LviU8_2),.clk(gclk));
	jdff dff_B_8e51ZPui5_2(.din(w_dff_B_uy03LviU8_2),.dout(w_dff_B_8e51ZPui5_2),.clk(gclk));
	jdff dff_B_UI1HZQrx3_2(.din(w_dff_B_8e51ZPui5_2),.dout(w_dff_B_UI1HZQrx3_2),.clk(gclk));
	jdff dff_B_ONbC3eCq1_2(.din(w_dff_B_UI1HZQrx3_2),.dout(w_dff_B_ONbC3eCq1_2),.clk(gclk));
	jdff dff_B_lfDjGvPZ0_2(.din(w_dff_B_ONbC3eCq1_2),.dout(w_dff_B_lfDjGvPZ0_2),.clk(gclk));
	jdff dff_B_CMs9GZ1y0_2(.din(w_dff_B_lfDjGvPZ0_2),.dout(w_dff_B_CMs9GZ1y0_2),.clk(gclk));
	jdff dff_B_4fPtujk65_2(.din(w_dff_B_CMs9GZ1y0_2),.dout(w_dff_B_4fPtujk65_2),.clk(gclk));
	jdff dff_B_mWon9R7R9_2(.din(w_dff_B_4fPtujk65_2),.dout(w_dff_B_mWon9R7R9_2),.clk(gclk));
	jdff dff_B_HuA5otXH4_2(.din(w_dff_B_mWon9R7R9_2),.dout(w_dff_B_HuA5otXH4_2),.clk(gclk));
	jdff dff_B_31jyz91C5_2(.din(w_dff_B_HuA5otXH4_2),.dout(w_dff_B_31jyz91C5_2),.clk(gclk));
	jdff dff_B_Kj3JMYLO7_2(.din(w_dff_B_31jyz91C5_2),.dout(w_dff_B_Kj3JMYLO7_2),.clk(gclk));
	jdff dff_B_rt2susp59_2(.din(w_dff_B_Kj3JMYLO7_2),.dout(w_dff_B_rt2susp59_2),.clk(gclk));
	jdff dff_B_moXigPB47_2(.din(w_dff_B_rt2susp59_2),.dout(w_dff_B_moXigPB47_2),.clk(gclk));
	jdff dff_B_Ey2tPuqD6_2(.din(w_dff_B_moXigPB47_2),.dout(w_dff_B_Ey2tPuqD6_2),.clk(gclk));
	jdff dff_B_7tL7QzxS7_2(.din(w_dff_B_Ey2tPuqD6_2),.dout(w_dff_B_7tL7QzxS7_2),.clk(gclk));
	jdff dff_B_k5cSsR3t0_2(.din(w_dff_B_7tL7QzxS7_2),.dout(w_dff_B_k5cSsR3t0_2),.clk(gclk));
	jdff dff_B_4755z2Hn7_2(.din(w_dff_B_k5cSsR3t0_2),.dout(w_dff_B_4755z2Hn7_2),.clk(gclk));
	jdff dff_B_s9yo5N0r9_2(.din(w_dff_B_4755z2Hn7_2),.dout(w_dff_B_s9yo5N0r9_2),.clk(gclk));
	jdff dff_B_OFXG6fSg7_2(.din(w_dff_B_s9yo5N0r9_2),.dout(w_dff_B_OFXG6fSg7_2),.clk(gclk));
	jdff dff_B_CFnvvsaX4_2(.din(w_dff_B_OFXG6fSg7_2),.dout(w_dff_B_CFnvvsaX4_2),.clk(gclk));
	jdff dff_B_wk8eK7oI1_2(.din(w_dff_B_CFnvvsaX4_2),.dout(w_dff_B_wk8eK7oI1_2),.clk(gclk));
	jdff dff_B_VoyoSs4I0_2(.din(w_dff_B_wk8eK7oI1_2),.dout(w_dff_B_VoyoSs4I0_2),.clk(gclk));
	jdff dff_B_NYN7OKw15_2(.din(w_dff_B_VoyoSs4I0_2),.dout(w_dff_B_NYN7OKw15_2),.clk(gclk));
	jdff dff_B_4ld0KiXW7_2(.din(w_dff_B_NYN7OKw15_2),.dout(w_dff_B_4ld0KiXW7_2),.clk(gclk));
	jdff dff_B_CxtvxXxF4_2(.din(w_dff_B_4ld0KiXW7_2),.dout(w_dff_B_CxtvxXxF4_2),.clk(gclk));
	jdff dff_B_ZhlFiBiX3_2(.din(w_dff_B_CxtvxXxF4_2),.dout(w_dff_B_ZhlFiBiX3_2),.clk(gclk));
	jdff dff_A_PWzSKAnh2_2(.dout(w_G137_3[2]),.din(w_dff_A_PWzSKAnh2_2),.clk(gclk));
	jdff dff_A_pJu6TLUw5_2(.dout(w_dff_A_PWzSKAnh2_2),.din(w_dff_A_pJu6TLUw5_2),.clk(gclk));
	jdff dff_A_VaawTq0Y3_2(.dout(w_dff_A_pJu6TLUw5_2),.din(w_dff_A_VaawTq0Y3_2),.clk(gclk));
	jdff dff_A_yOYMrknm3_2(.dout(w_dff_A_VaawTq0Y3_2),.din(w_dff_A_yOYMrknm3_2),.clk(gclk));
	jdff dff_A_s6wrYOsC1_2(.dout(w_dff_A_yOYMrknm3_2),.din(w_dff_A_s6wrYOsC1_2),.clk(gclk));
	jdff dff_A_LsHyNQB36_2(.dout(w_dff_A_s6wrYOsC1_2),.din(w_dff_A_LsHyNQB36_2),.clk(gclk));
	jdff dff_A_48j3K6HD4_2(.dout(w_dff_A_LsHyNQB36_2),.din(w_dff_A_48j3K6HD4_2),.clk(gclk));
	jdff dff_A_eqg8PPEo6_2(.dout(w_dff_A_48j3K6HD4_2),.din(w_dff_A_eqg8PPEo6_2),.clk(gclk));
	jdff dff_A_ELQkdxmX1_2(.dout(w_dff_A_eqg8PPEo6_2),.din(w_dff_A_ELQkdxmX1_2),.clk(gclk));
	jdff dff_A_uuq7jWJm9_2(.dout(w_dff_A_ELQkdxmX1_2),.din(w_dff_A_uuq7jWJm9_2),.clk(gclk));
	jdff dff_A_LBfUyJGt2_2(.dout(w_dff_A_uuq7jWJm9_2),.din(w_dff_A_LBfUyJGt2_2),.clk(gclk));
	jdff dff_A_vnLBMEmj1_2(.dout(w_dff_A_LBfUyJGt2_2),.din(w_dff_A_vnLBMEmj1_2),.clk(gclk));
	jdff dff_A_6VPhDO5v1_2(.dout(w_dff_A_vnLBMEmj1_2),.din(w_dff_A_6VPhDO5v1_2),.clk(gclk));
	jdff dff_A_RMshaW478_2(.dout(w_dff_A_6VPhDO5v1_2),.din(w_dff_A_RMshaW478_2),.clk(gclk));
	jdff dff_A_ZSAPFrF88_2(.dout(w_dff_A_RMshaW478_2),.din(w_dff_A_ZSAPFrF88_2),.clk(gclk));
	jdff dff_A_vKJ96aS84_2(.dout(w_dff_A_ZSAPFrF88_2),.din(w_dff_A_vKJ96aS84_2),.clk(gclk));
	jdff dff_A_xRPTxXmC9_2(.dout(w_dff_A_vKJ96aS84_2),.din(w_dff_A_xRPTxXmC9_2),.clk(gclk));
	jdff dff_A_Io6h3bx43_2(.dout(w_dff_A_xRPTxXmC9_2),.din(w_dff_A_Io6h3bx43_2),.clk(gclk));
	jdff dff_A_B9ujESKV2_2(.dout(w_dff_A_Io6h3bx43_2),.din(w_dff_A_B9ujESKV2_2),.clk(gclk));
	jdff dff_A_B02DsWh05_2(.dout(w_dff_A_B9ujESKV2_2),.din(w_dff_A_B02DsWh05_2),.clk(gclk));
	jdff dff_A_C0zyaOhS4_2(.dout(w_dff_A_B02DsWh05_2),.din(w_dff_A_C0zyaOhS4_2),.clk(gclk));
	jdff dff_A_7KLxEBCn3_2(.dout(w_dff_A_C0zyaOhS4_2),.din(w_dff_A_7KLxEBCn3_2),.clk(gclk));
	jdff dff_A_6QicL7n99_2(.dout(w_dff_A_7KLxEBCn3_2),.din(w_dff_A_6QicL7n99_2),.clk(gclk));
	jdff dff_A_tdkmqNYI7_2(.dout(w_dff_A_6QicL7n99_2),.din(w_dff_A_tdkmqNYI7_2),.clk(gclk));
	jdff dff_A_JaX8JiOJ9_0(.dout(w_G137_0[0]),.din(w_dff_A_JaX8JiOJ9_0),.clk(gclk));
	jdff dff_A_DWFiqVPp2_0(.dout(w_dff_A_JaX8JiOJ9_0),.din(w_dff_A_DWFiqVPp2_0),.clk(gclk));
	jdff dff_A_4Y8E3njp6_0(.dout(w_dff_A_DWFiqVPp2_0),.din(w_dff_A_4Y8E3njp6_0),.clk(gclk));
	jdff dff_A_uTKog0qp3_0(.dout(w_dff_A_4Y8E3njp6_0),.din(w_dff_A_uTKog0qp3_0),.clk(gclk));
	jdff dff_A_Yl6sBJFe7_0(.dout(w_dff_A_uTKog0qp3_0),.din(w_dff_A_Yl6sBJFe7_0),.clk(gclk));
	jdff dff_A_vrU1h5q76_0(.dout(w_dff_A_Yl6sBJFe7_0),.din(w_dff_A_vrU1h5q76_0),.clk(gclk));
	jdff dff_A_6h6MoGTq4_0(.dout(w_dff_A_vrU1h5q76_0),.din(w_dff_A_6h6MoGTq4_0),.clk(gclk));
	jdff dff_A_3sz47knn2_0(.dout(w_dff_A_6h6MoGTq4_0),.din(w_dff_A_3sz47knn2_0),.clk(gclk));
	jdff dff_A_5Z5PhRWw2_0(.dout(w_dff_A_3sz47knn2_0),.din(w_dff_A_5Z5PhRWw2_0),.clk(gclk));
	jdff dff_A_4qQJtJNU1_0(.dout(w_dff_A_5Z5PhRWw2_0),.din(w_dff_A_4qQJtJNU1_0),.clk(gclk));
	jdff dff_A_qxrKAmvh1_0(.dout(w_dff_A_4qQJtJNU1_0),.din(w_dff_A_qxrKAmvh1_0),.clk(gclk));
	jdff dff_A_8SFuhkZz4_0(.dout(w_dff_A_qxrKAmvh1_0),.din(w_dff_A_8SFuhkZz4_0),.clk(gclk));
	jdff dff_A_fLt2uriD4_0(.dout(w_dff_A_8SFuhkZz4_0),.din(w_dff_A_fLt2uriD4_0),.clk(gclk));
	jdff dff_A_XYpH9AIa3_0(.dout(w_dff_A_fLt2uriD4_0),.din(w_dff_A_XYpH9AIa3_0),.clk(gclk));
	jdff dff_A_8HvueTtx2_0(.dout(w_dff_A_XYpH9AIa3_0),.din(w_dff_A_8HvueTtx2_0),.clk(gclk));
	jdff dff_A_1IJ4gebr6_0(.dout(w_dff_A_8HvueTtx2_0),.din(w_dff_A_1IJ4gebr6_0),.clk(gclk));
	jdff dff_A_yOntMPx73_0(.dout(w_dff_A_1IJ4gebr6_0),.din(w_dff_A_yOntMPx73_0),.clk(gclk));
	jdff dff_A_PgPS7vHF7_1(.dout(w_G137_0[1]),.din(w_dff_A_PgPS7vHF7_1),.clk(gclk));
	jdff dff_A_U7LGI2NW6_1(.dout(w_dff_A_PgPS7vHF7_1),.din(w_dff_A_U7LGI2NW6_1),.clk(gclk));
	jdff dff_A_5H0sIIw53_1(.dout(w_dff_A_U7LGI2NW6_1),.din(w_dff_A_5H0sIIw53_1),.clk(gclk));
	jdff dff_A_vR1YJq4y5_1(.dout(w_dff_A_5H0sIIw53_1),.din(w_dff_A_vR1YJq4y5_1),.clk(gclk));
	jdff dff_A_E6SiKNQJ1_1(.dout(w_dff_A_vR1YJq4y5_1),.din(w_dff_A_E6SiKNQJ1_1),.clk(gclk));
	jdff dff_A_Dnlmsim40_1(.dout(w_dff_A_E6SiKNQJ1_1),.din(w_dff_A_Dnlmsim40_1),.clk(gclk));
	jdff dff_A_IfxHcgWw0_1(.dout(w_dff_A_Dnlmsim40_1),.din(w_dff_A_IfxHcgWw0_1),.clk(gclk));
	jdff dff_A_CS1XUDc44_1(.dout(w_dff_A_IfxHcgWw0_1),.din(w_dff_A_CS1XUDc44_1),.clk(gclk));
	jdff dff_A_lgskrCNj6_1(.dout(w_dff_A_CS1XUDc44_1),.din(w_dff_A_lgskrCNj6_1),.clk(gclk));
	jdff dff_A_TaMCCUBL4_1(.dout(w_dff_A_lgskrCNj6_1),.din(w_dff_A_TaMCCUBL4_1),.clk(gclk));
	jdff dff_A_cLxrOEJU8_1(.dout(w_dff_A_TaMCCUBL4_1),.din(w_dff_A_cLxrOEJU8_1),.clk(gclk));
	jdff dff_A_BhUrfjsT4_1(.dout(w_dff_A_cLxrOEJU8_1),.din(w_dff_A_BhUrfjsT4_1),.clk(gclk));
	jdff dff_A_MyMfKrmE2_1(.dout(w_dff_A_BhUrfjsT4_1),.din(w_dff_A_MyMfKrmE2_1),.clk(gclk));
	jdff dff_A_UikOBbBR2_1(.dout(w_dff_A_MyMfKrmE2_1),.din(w_dff_A_UikOBbBR2_1),.clk(gclk));
	jdff dff_A_fEh8IIwQ7_1(.dout(w_dff_A_UikOBbBR2_1),.din(w_dff_A_fEh8IIwQ7_1),.clk(gclk));
	jdff dff_A_3qesbko21_1(.dout(w_dff_A_rZMUeqtT1_0),.din(w_dff_A_3qesbko21_1),.clk(gclk));
	jdff dff_A_rZMUeqtT1_0(.dout(w_dff_A_2xZl2LHc0_0),.din(w_dff_A_rZMUeqtT1_0),.clk(gclk));
	jdff dff_A_2xZl2LHc0_0(.dout(w_dff_A_o4hKRHkh8_0),.din(w_dff_A_2xZl2LHc0_0),.clk(gclk));
	jdff dff_A_o4hKRHkh8_0(.dout(w_dff_A_fbl2CEZY5_0),.din(w_dff_A_o4hKRHkh8_0),.clk(gclk));
	jdff dff_A_fbl2CEZY5_0(.dout(w_dff_A_LmrBxr9C2_0),.din(w_dff_A_fbl2CEZY5_0),.clk(gclk));
	jdff dff_A_LmrBxr9C2_0(.dout(w_dff_A_DOIi9s5f9_0),.din(w_dff_A_LmrBxr9C2_0),.clk(gclk));
	jdff dff_A_DOIi9s5f9_0(.dout(w_dff_A_9iYeXxQm9_0),.din(w_dff_A_DOIi9s5f9_0),.clk(gclk));
	jdff dff_A_9iYeXxQm9_0(.dout(w_dff_A_DQTCx7PV6_0),.din(w_dff_A_9iYeXxQm9_0),.clk(gclk));
	jdff dff_A_DQTCx7PV6_0(.dout(w_dff_A_9pd7nHgI1_0),.din(w_dff_A_DQTCx7PV6_0),.clk(gclk));
	jdff dff_A_9pd7nHgI1_0(.dout(w_dff_A_U7Vz4sXe9_0),.din(w_dff_A_9pd7nHgI1_0),.clk(gclk));
	jdff dff_A_U7Vz4sXe9_0(.dout(w_dff_A_Rk1zU4oN8_0),.din(w_dff_A_U7Vz4sXe9_0),.clk(gclk));
	jdff dff_A_Rk1zU4oN8_0(.dout(w_dff_A_8EcYE1yi1_0),.din(w_dff_A_Rk1zU4oN8_0),.clk(gclk));
	jdff dff_A_8EcYE1yi1_0(.dout(w_dff_A_kXzompdx0_0),.din(w_dff_A_8EcYE1yi1_0),.clk(gclk));
	jdff dff_A_kXzompdx0_0(.dout(w_dff_A_N1qdQRdK4_0),.din(w_dff_A_kXzompdx0_0),.clk(gclk));
	jdff dff_A_N1qdQRdK4_0(.dout(w_dff_A_UP7Tw7xo6_0),.din(w_dff_A_N1qdQRdK4_0),.clk(gclk));
	jdff dff_A_UP7Tw7xo6_0(.dout(w_dff_A_4BObyJuZ0_0),.din(w_dff_A_UP7Tw7xo6_0),.clk(gclk));
	jdff dff_A_4BObyJuZ0_0(.dout(w_dff_A_9IdfYSln5_0),.din(w_dff_A_4BObyJuZ0_0),.clk(gclk));
	jdff dff_A_9IdfYSln5_0(.dout(w_dff_A_jdP6U8b07_0),.din(w_dff_A_9IdfYSln5_0),.clk(gclk));
	jdff dff_A_jdP6U8b07_0(.dout(w_dff_A_kZqzrERF1_0),.din(w_dff_A_jdP6U8b07_0),.clk(gclk));
	jdff dff_A_kZqzrERF1_0(.dout(w_dff_A_JS09NjOF6_0),.din(w_dff_A_kZqzrERF1_0),.clk(gclk));
	jdff dff_A_JS09NjOF6_0(.dout(w_dff_A_izbnWL9K6_0),.din(w_dff_A_JS09NjOF6_0),.clk(gclk));
	jdff dff_A_izbnWL9K6_0(.dout(w_dff_A_WgQjA4mu7_0),.din(w_dff_A_izbnWL9K6_0),.clk(gclk));
	jdff dff_A_WgQjA4mu7_0(.dout(w_dff_A_5kcqco9f3_0),.din(w_dff_A_WgQjA4mu7_0),.clk(gclk));
	jdff dff_A_5kcqco9f3_0(.dout(w_dff_A_PW2Da1iG2_0),.din(w_dff_A_5kcqco9f3_0),.clk(gclk));
	jdff dff_A_PW2Da1iG2_0(.dout(w_dff_A_JFty1vSw1_0),.din(w_dff_A_PW2Da1iG2_0),.clk(gclk));
	jdff dff_A_JFty1vSw1_0(.dout(w_dff_A_Kk4Jsm8Y5_0),.din(w_dff_A_JFty1vSw1_0),.clk(gclk));
	jdff dff_A_Kk4Jsm8Y5_0(.dout(G144),.din(w_dff_A_Kk4Jsm8Y5_0),.clk(gclk));
	jdff dff_A_k5hS1sGE3_1(.dout(w_dff_A_8uWlESyb2_0),.din(w_dff_A_k5hS1sGE3_1),.clk(gclk));
	jdff dff_A_8uWlESyb2_0(.dout(w_dff_A_ZxbXG1ZX7_0),.din(w_dff_A_8uWlESyb2_0),.clk(gclk));
	jdff dff_A_ZxbXG1ZX7_0(.dout(w_dff_A_XUqMXgsB7_0),.din(w_dff_A_ZxbXG1ZX7_0),.clk(gclk));
	jdff dff_A_XUqMXgsB7_0(.dout(w_dff_A_Ke4YvWgH0_0),.din(w_dff_A_XUqMXgsB7_0),.clk(gclk));
	jdff dff_A_Ke4YvWgH0_0(.dout(w_dff_A_jyng7xC70_0),.din(w_dff_A_Ke4YvWgH0_0),.clk(gclk));
	jdff dff_A_jyng7xC70_0(.dout(w_dff_A_Y917uZt44_0),.din(w_dff_A_jyng7xC70_0),.clk(gclk));
	jdff dff_A_Y917uZt44_0(.dout(w_dff_A_NC2HOdeJ7_0),.din(w_dff_A_Y917uZt44_0),.clk(gclk));
	jdff dff_A_NC2HOdeJ7_0(.dout(w_dff_A_4a5o1oev5_0),.din(w_dff_A_NC2HOdeJ7_0),.clk(gclk));
	jdff dff_A_4a5o1oev5_0(.dout(w_dff_A_cYgNx4oo5_0),.din(w_dff_A_4a5o1oev5_0),.clk(gclk));
	jdff dff_A_cYgNx4oo5_0(.dout(w_dff_A_b7edN0jj3_0),.din(w_dff_A_cYgNx4oo5_0),.clk(gclk));
	jdff dff_A_b7edN0jj3_0(.dout(w_dff_A_XuUOAamh3_0),.din(w_dff_A_b7edN0jj3_0),.clk(gclk));
	jdff dff_A_XuUOAamh3_0(.dout(w_dff_A_mZbRYjb50_0),.din(w_dff_A_XuUOAamh3_0),.clk(gclk));
	jdff dff_A_mZbRYjb50_0(.dout(w_dff_A_PbfIIqdM0_0),.din(w_dff_A_mZbRYjb50_0),.clk(gclk));
	jdff dff_A_PbfIIqdM0_0(.dout(w_dff_A_7pT2pHSk2_0),.din(w_dff_A_PbfIIqdM0_0),.clk(gclk));
	jdff dff_A_7pT2pHSk2_0(.dout(w_dff_A_ROW0QVMA0_0),.din(w_dff_A_7pT2pHSk2_0),.clk(gclk));
	jdff dff_A_ROW0QVMA0_0(.dout(w_dff_A_6WUchvPs2_0),.din(w_dff_A_ROW0QVMA0_0),.clk(gclk));
	jdff dff_A_6WUchvPs2_0(.dout(w_dff_A_P1xrhZVX1_0),.din(w_dff_A_6WUchvPs2_0),.clk(gclk));
	jdff dff_A_P1xrhZVX1_0(.dout(w_dff_A_q4ZuV6WA7_0),.din(w_dff_A_P1xrhZVX1_0),.clk(gclk));
	jdff dff_A_q4ZuV6WA7_0(.dout(w_dff_A_kKeVad1S9_0),.din(w_dff_A_q4ZuV6WA7_0),.clk(gclk));
	jdff dff_A_kKeVad1S9_0(.dout(w_dff_A_IevzEcxt4_0),.din(w_dff_A_kKeVad1S9_0),.clk(gclk));
	jdff dff_A_IevzEcxt4_0(.dout(w_dff_A_TeifZMw32_0),.din(w_dff_A_IevzEcxt4_0),.clk(gclk));
	jdff dff_A_TeifZMw32_0(.dout(w_dff_A_Xm0W3xgQ8_0),.din(w_dff_A_TeifZMw32_0),.clk(gclk));
	jdff dff_A_Xm0W3xgQ8_0(.dout(w_dff_A_vjGNUgun3_0),.din(w_dff_A_Xm0W3xgQ8_0),.clk(gclk));
	jdff dff_A_vjGNUgun3_0(.dout(w_dff_A_xCMijMMy9_0),.din(w_dff_A_vjGNUgun3_0),.clk(gclk));
	jdff dff_A_xCMijMMy9_0(.dout(w_dff_A_6VqqoTRR5_0),.din(w_dff_A_xCMijMMy9_0),.clk(gclk));
	jdff dff_A_6VqqoTRR5_0(.dout(w_dff_A_bVoxBf3X7_0),.din(w_dff_A_6VqqoTRR5_0),.clk(gclk));
	jdff dff_A_bVoxBf3X7_0(.dout(G298),.din(w_dff_A_bVoxBf3X7_0),.clk(gclk));
	jdff dff_A_d6kwjLVZ0_1(.dout(w_dff_A_Zs4FhmDx9_0),.din(w_dff_A_d6kwjLVZ0_1),.clk(gclk));
	jdff dff_A_Zs4FhmDx9_0(.dout(w_dff_A_udvjerb55_0),.din(w_dff_A_Zs4FhmDx9_0),.clk(gclk));
	jdff dff_A_udvjerb55_0(.dout(w_dff_A_jHunwUCV1_0),.din(w_dff_A_udvjerb55_0),.clk(gclk));
	jdff dff_A_jHunwUCV1_0(.dout(w_dff_A_ojg6VGAY8_0),.din(w_dff_A_jHunwUCV1_0),.clk(gclk));
	jdff dff_A_ojg6VGAY8_0(.dout(w_dff_A_twwtg2867_0),.din(w_dff_A_ojg6VGAY8_0),.clk(gclk));
	jdff dff_A_twwtg2867_0(.dout(w_dff_A_QQUPyo6B3_0),.din(w_dff_A_twwtg2867_0),.clk(gclk));
	jdff dff_A_QQUPyo6B3_0(.dout(w_dff_A_aKnkfTMm3_0),.din(w_dff_A_QQUPyo6B3_0),.clk(gclk));
	jdff dff_A_aKnkfTMm3_0(.dout(w_dff_A_griBH8TH1_0),.din(w_dff_A_aKnkfTMm3_0),.clk(gclk));
	jdff dff_A_griBH8TH1_0(.dout(w_dff_A_WkKUe34a9_0),.din(w_dff_A_griBH8TH1_0),.clk(gclk));
	jdff dff_A_WkKUe34a9_0(.dout(w_dff_A_cUFSCdBl4_0),.din(w_dff_A_WkKUe34a9_0),.clk(gclk));
	jdff dff_A_cUFSCdBl4_0(.dout(w_dff_A_jV4oyZOf2_0),.din(w_dff_A_cUFSCdBl4_0),.clk(gclk));
	jdff dff_A_jV4oyZOf2_0(.dout(w_dff_A_KWia5jN18_0),.din(w_dff_A_jV4oyZOf2_0),.clk(gclk));
	jdff dff_A_KWia5jN18_0(.dout(w_dff_A_FV4HJGny4_0),.din(w_dff_A_KWia5jN18_0),.clk(gclk));
	jdff dff_A_FV4HJGny4_0(.dout(w_dff_A_NkiHE9p90_0),.din(w_dff_A_FV4HJGny4_0),.clk(gclk));
	jdff dff_A_NkiHE9p90_0(.dout(w_dff_A_hD5vSv531_0),.din(w_dff_A_NkiHE9p90_0),.clk(gclk));
	jdff dff_A_hD5vSv531_0(.dout(w_dff_A_mLW3L2zd3_0),.din(w_dff_A_hD5vSv531_0),.clk(gclk));
	jdff dff_A_mLW3L2zd3_0(.dout(w_dff_A_gTUaK7PN3_0),.din(w_dff_A_mLW3L2zd3_0),.clk(gclk));
	jdff dff_A_gTUaK7PN3_0(.dout(w_dff_A_9GUhU2QS7_0),.din(w_dff_A_gTUaK7PN3_0),.clk(gclk));
	jdff dff_A_9GUhU2QS7_0(.dout(w_dff_A_lpMKehaN0_0),.din(w_dff_A_9GUhU2QS7_0),.clk(gclk));
	jdff dff_A_lpMKehaN0_0(.dout(w_dff_A_tLHd8NGO8_0),.din(w_dff_A_lpMKehaN0_0),.clk(gclk));
	jdff dff_A_tLHd8NGO8_0(.dout(w_dff_A_osog69XA8_0),.din(w_dff_A_tLHd8NGO8_0),.clk(gclk));
	jdff dff_A_osog69XA8_0(.dout(w_dff_A_8Y1H6pcH4_0),.din(w_dff_A_osog69XA8_0),.clk(gclk));
	jdff dff_A_8Y1H6pcH4_0(.dout(w_dff_A_8MYk7QEc1_0),.din(w_dff_A_8Y1H6pcH4_0),.clk(gclk));
	jdff dff_A_8MYk7QEc1_0(.dout(w_dff_A_THwqZlsa1_0),.din(w_dff_A_8MYk7QEc1_0),.clk(gclk));
	jdff dff_A_THwqZlsa1_0(.dout(w_dff_A_fzLeF5Br9_0),.din(w_dff_A_THwqZlsa1_0),.clk(gclk));
	jdff dff_A_fzLeF5Br9_0(.dout(w_dff_A_JfqOrBRk2_0),.din(w_dff_A_fzLeF5Br9_0),.clk(gclk));
	jdff dff_A_JfqOrBRk2_0(.dout(G973),.din(w_dff_A_JfqOrBRk2_0),.clk(gclk));
	jdff dff_A_VHpW1ILW7_1(.dout(w_dff_A_0EdNBvdh9_0),.din(w_dff_A_VHpW1ILW7_1),.clk(gclk));
	jdff dff_A_0EdNBvdh9_0(.dout(w_dff_A_D4OkyQ4G9_0),.din(w_dff_A_0EdNBvdh9_0),.clk(gclk));
	jdff dff_A_D4OkyQ4G9_0(.dout(w_dff_A_QfKA9iXQ7_0),.din(w_dff_A_D4OkyQ4G9_0),.clk(gclk));
	jdff dff_A_QfKA9iXQ7_0(.dout(w_dff_A_wOhFogC16_0),.din(w_dff_A_QfKA9iXQ7_0),.clk(gclk));
	jdff dff_A_wOhFogC16_0(.dout(w_dff_A_UGs0r12P4_0),.din(w_dff_A_wOhFogC16_0),.clk(gclk));
	jdff dff_A_UGs0r12P4_0(.dout(w_dff_A_zaSpRqku1_0),.din(w_dff_A_UGs0r12P4_0),.clk(gclk));
	jdff dff_A_zaSpRqku1_0(.dout(w_dff_A_dbPsrNvz1_0),.din(w_dff_A_zaSpRqku1_0),.clk(gclk));
	jdff dff_A_dbPsrNvz1_0(.dout(w_dff_A_HoAwRdxX7_0),.din(w_dff_A_dbPsrNvz1_0),.clk(gclk));
	jdff dff_A_HoAwRdxX7_0(.dout(w_dff_A_8QFTlGAL7_0),.din(w_dff_A_HoAwRdxX7_0),.clk(gclk));
	jdff dff_A_8QFTlGAL7_0(.dout(w_dff_A_9jFSz56R8_0),.din(w_dff_A_8QFTlGAL7_0),.clk(gclk));
	jdff dff_A_9jFSz56R8_0(.dout(w_dff_A_urHNbyaD5_0),.din(w_dff_A_9jFSz56R8_0),.clk(gclk));
	jdff dff_A_urHNbyaD5_0(.dout(w_dff_A_smurInE44_0),.din(w_dff_A_urHNbyaD5_0),.clk(gclk));
	jdff dff_A_smurInE44_0(.dout(w_dff_A_cc0bom7j3_0),.din(w_dff_A_smurInE44_0),.clk(gclk));
	jdff dff_A_cc0bom7j3_0(.dout(w_dff_A_oZePYS4c6_0),.din(w_dff_A_cc0bom7j3_0),.clk(gclk));
	jdff dff_A_oZePYS4c6_0(.dout(w_dff_A_Bo94DYig0_0),.din(w_dff_A_oZePYS4c6_0),.clk(gclk));
	jdff dff_A_Bo94DYig0_0(.dout(w_dff_A_MErWuuNG0_0),.din(w_dff_A_Bo94DYig0_0),.clk(gclk));
	jdff dff_A_MErWuuNG0_0(.dout(w_dff_A_pCcJklv01_0),.din(w_dff_A_MErWuuNG0_0),.clk(gclk));
	jdff dff_A_pCcJklv01_0(.dout(w_dff_A_JKooQMiB5_0),.din(w_dff_A_pCcJklv01_0),.clk(gclk));
	jdff dff_A_JKooQMiB5_0(.dout(w_dff_A_KKURhmtQ4_0),.din(w_dff_A_JKooQMiB5_0),.clk(gclk));
	jdff dff_A_KKURhmtQ4_0(.dout(w_dff_A_QmFJHWQj2_0),.din(w_dff_A_KKURhmtQ4_0),.clk(gclk));
	jdff dff_A_QmFJHWQj2_0(.dout(w_dff_A_SFC6N8698_0),.din(w_dff_A_QmFJHWQj2_0),.clk(gclk));
	jdff dff_A_SFC6N8698_0(.dout(w_dff_A_6rukfAPk6_0),.din(w_dff_A_SFC6N8698_0),.clk(gclk));
	jdff dff_A_6rukfAPk6_0(.dout(w_dff_A_YTZ4OCzy0_0),.din(w_dff_A_6rukfAPk6_0),.clk(gclk));
	jdff dff_A_YTZ4OCzy0_0(.dout(w_dff_A_OZW0BpKb4_0),.din(w_dff_A_YTZ4OCzy0_0),.clk(gclk));
	jdff dff_A_OZW0BpKb4_0(.dout(w_dff_A_Pkn8qxHJ5_0),.din(w_dff_A_OZW0BpKb4_0),.clk(gclk));
	jdff dff_A_Pkn8qxHJ5_0(.dout(w_dff_A_PCekqYEQ0_0),.din(w_dff_A_Pkn8qxHJ5_0),.clk(gclk));
	jdff dff_A_PCekqYEQ0_0(.dout(G594),.din(w_dff_A_PCekqYEQ0_0),.clk(gclk));
	jdff dff_A_2GuE02g96_1(.dout(w_dff_A_0qKeY6Yy4_0),.din(w_dff_A_2GuE02g96_1),.clk(gclk));
	jdff dff_A_0qKeY6Yy4_0(.dout(w_dff_A_P27MWUUx8_0),.din(w_dff_A_0qKeY6Yy4_0),.clk(gclk));
	jdff dff_A_P27MWUUx8_0(.dout(w_dff_A_kllTJxuw5_0),.din(w_dff_A_P27MWUUx8_0),.clk(gclk));
	jdff dff_A_kllTJxuw5_0(.dout(w_dff_A_XIJ9hcLF3_0),.din(w_dff_A_kllTJxuw5_0),.clk(gclk));
	jdff dff_A_XIJ9hcLF3_0(.dout(w_dff_A_uMbhdoe53_0),.din(w_dff_A_XIJ9hcLF3_0),.clk(gclk));
	jdff dff_A_uMbhdoe53_0(.dout(w_dff_A_uVwGQOzg1_0),.din(w_dff_A_uMbhdoe53_0),.clk(gclk));
	jdff dff_A_uVwGQOzg1_0(.dout(w_dff_A_ajn1NoHo4_0),.din(w_dff_A_uVwGQOzg1_0),.clk(gclk));
	jdff dff_A_ajn1NoHo4_0(.dout(w_dff_A_ZMYKSxSU9_0),.din(w_dff_A_ajn1NoHo4_0),.clk(gclk));
	jdff dff_A_ZMYKSxSU9_0(.dout(w_dff_A_4h0mS7gB3_0),.din(w_dff_A_ZMYKSxSU9_0),.clk(gclk));
	jdff dff_A_4h0mS7gB3_0(.dout(w_dff_A_RrypEcrR9_0),.din(w_dff_A_4h0mS7gB3_0),.clk(gclk));
	jdff dff_A_RrypEcrR9_0(.dout(w_dff_A_Xjea6bvo8_0),.din(w_dff_A_RrypEcrR9_0),.clk(gclk));
	jdff dff_A_Xjea6bvo8_0(.dout(w_dff_A_QKlP35xm6_0),.din(w_dff_A_Xjea6bvo8_0),.clk(gclk));
	jdff dff_A_QKlP35xm6_0(.dout(w_dff_A_ce8jm6bc2_0),.din(w_dff_A_QKlP35xm6_0),.clk(gclk));
	jdff dff_A_ce8jm6bc2_0(.dout(w_dff_A_fXEt5rXm9_0),.din(w_dff_A_ce8jm6bc2_0),.clk(gclk));
	jdff dff_A_fXEt5rXm9_0(.dout(w_dff_A_HNZ1HHDk2_0),.din(w_dff_A_fXEt5rXm9_0),.clk(gclk));
	jdff dff_A_HNZ1HHDk2_0(.dout(w_dff_A_cm8vsMiB2_0),.din(w_dff_A_HNZ1HHDk2_0),.clk(gclk));
	jdff dff_A_cm8vsMiB2_0(.dout(w_dff_A_mN0D8Rpu3_0),.din(w_dff_A_cm8vsMiB2_0),.clk(gclk));
	jdff dff_A_mN0D8Rpu3_0(.dout(w_dff_A_Q8rV6Zat7_0),.din(w_dff_A_mN0D8Rpu3_0),.clk(gclk));
	jdff dff_A_Q8rV6Zat7_0(.dout(w_dff_A_t7wZdGwX1_0),.din(w_dff_A_Q8rV6Zat7_0),.clk(gclk));
	jdff dff_A_t7wZdGwX1_0(.dout(w_dff_A_KJ8rTuVl5_0),.din(w_dff_A_t7wZdGwX1_0),.clk(gclk));
	jdff dff_A_KJ8rTuVl5_0(.dout(w_dff_A_zlVkK4YB4_0),.din(w_dff_A_KJ8rTuVl5_0),.clk(gclk));
	jdff dff_A_zlVkK4YB4_0(.dout(w_dff_A_Taqzk2LZ4_0),.din(w_dff_A_zlVkK4YB4_0),.clk(gclk));
	jdff dff_A_Taqzk2LZ4_0(.dout(w_dff_A_S6zLf6W24_0),.din(w_dff_A_Taqzk2LZ4_0),.clk(gclk));
	jdff dff_A_S6zLf6W24_0(.dout(w_dff_A_7r8n76n82_0),.din(w_dff_A_S6zLf6W24_0),.clk(gclk));
	jdff dff_A_7r8n76n82_0(.dout(w_dff_A_GVBvY17J3_0),.din(w_dff_A_7r8n76n82_0),.clk(gclk));
	jdff dff_A_GVBvY17J3_0(.dout(w_dff_A_qZdKgzVe7_0),.din(w_dff_A_GVBvY17J3_0),.clk(gclk));
	jdff dff_A_qZdKgzVe7_0(.dout(G599),.din(w_dff_A_qZdKgzVe7_0),.clk(gclk));
	jdff dff_A_63AobLUF2_1(.dout(w_dff_A_dAlUDEjG1_0),.din(w_dff_A_63AobLUF2_1),.clk(gclk));
	jdff dff_A_dAlUDEjG1_0(.dout(w_dff_A_tejdBBNT0_0),.din(w_dff_A_dAlUDEjG1_0),.clk(gclk));
	jdff dff_A_tejdBBNT0_0(.dout(w_dff_A_xzriuna22_0),.din(w_dff_A_tejdBBNT0_0),.clk(gclk));
	jdff dff_A_xzriuna22_0(.dout(w_dff_A_Mf5s9S5i2_0),.din(w_dff_A_xzriuna22_0),.clk(gclk));
	jdff dff_A_Mf5s9S5i2_0(.dout(w_dff_A_phDcnlxx3_0),.din(w_dff_A_Mf5s9S5i2_0),.clk(gclk));
	jdff dff_A_phDcnlxx3_0(.dout(w_dff_A_Ld3TBmQB5_0),.din(w_dff_A_phDcnlxx3_0),.clk(gclk));
	jdff dff_A_Ld3TBmQB5_0(.dout(w_dff_A_aCUV8FGK3_0),.din(w_dff_A_Ld3TBmQB5_0),.clk(gclk));
	jdff dff_A_aCUV8FGK3_0(.dout(w_dff_A_ylPMQHgv6_0),.din(w_dff_A_aCUV8FGK3_0),.clk(gclk));
	jdff dff_A_ylPMQHgv6_0(.dout(w_dff_A_18iQsGit3_0),.din(w_dff_A_ylPMQHgv6_0),.clk(gclk));
	jdff dff_A_18iQsGit3_0(.dout(w_dff_A_HQp5Isk29_0),.din(w_dff_A_18iQsGit3_0),.clk(gclk));
	jdff dff_A_HQp5Isk29_0(.dout(w_dff_A_4pNBlFnC9_0),.din(w_dff_A_HQp5Isk29_0),.clk(gclk));
	jdff dff_A_4pNBlFnC9_0(.dout(w_dff_A_cegTMNkz5_0),.din(w_dff_A_4pNBlFnC9_0),.clk(gclk));
	jdff dff_A_cegTMNkz5_0(.dout(w_dff_A_LuWf17Ek6_0),.din(w_dff_A_cegTMNkz5_0),.clk(gclk));
	jdff dff_A_LuWf17Ek6_0(.dout(w_dff_A_olEg0y025_0),.din(w_dff_A_LuWf17Ek6_0),.clk(gclk));
	jdff dff_A_olEg0y025_0(.dout(w_dff_A_tmqmlhJE8_0),.din(w_dff_A_olEg0y025_0),.clk(gclk));
	jdff dff_A_tmqmlhJE8_0(.dout(w_dff_A_LNVrH9Rq0_0),.din(w_dff_A_tmqmlhJE8_0),.clk(gclk));
	jdff dff_A_LNVrH9Rq0_0(.dout(w_dff_A_exksNRci6_0),.din(w_dff_A_LNVrH9Rq0_0),.clk(gclk));
	jdff dff_A_exksNRci6_0(.dout(w_dff_A_KVigNA9U1_0),.din(w_dff_A_exksNRci6_0),.clk(gclk));
	jdff dff_A_KVigNA9U1_0(.dout(w_dff_A_dAUd8jss8_0),.din(w_dff_A_KVigNA9U1_0),.clk(gclk));
	jdff dff_A_dAUd8jss8_0(.dout(w_dff_A_d9VRJBek8_0),.din(w_dff_A_dAUd8jss8_0),.clk(gclk));
	jdff dff_A_d9VRJBek8_0(.dout(w_dff_A_n6PlnGlr2_0),.din(w_dff_A_d9VRJBek8_0),.clk(gclk));
	jdff dff_A_n6PlnGlr2_0(.dout(w_dff_A_5wiTCPxQ0_0),.din(w_dff_A_n6PlnGlr2_0),.clk(gclk));
	jdff dff_A_5wiTCPxQ0_0(.dout(w_dff_A_Ne1VqeQd2_0),.din(w_dff_A_5wiTCPxQ0_0),.clk(gclk));
	jdff dff_A_Ne1VqeQd2_0(.dout(w_dff_A_ToJmm2N25_0),.din(w_dff_A_Ne1VqeQd2_0),.clk(gclk));
	jdff dff_A_ToJmm2N25_0(.dout(w_dff_A_Iy23Gdq82_0),.din(w_dff_A_ToJmm2N25_0),.clk(gclk));
	jdff dff_A_Iy23Gdq82_0(.dout(w_dff_A_A0RiMfTY7_0),.din(w_dff_A_Iy23Gdq82_0),.clk(gclk));
	jdff dff_A_A0RiMfTY7_0(.dout(G600),.din(w_dff_A_A0RiMfTY7_0),.clk(gclk));
	jdff dff_A_xSrgjd2r2_1(.dout(w_dff_A_z1MV1RVm5_0),.din(w_dff_A_xSrgjd2r2_1),.clk(gclk));
	jdff dff_A_z1MV1RVm5_0(.dout(w_dff_A_NCvQSvrP0_0),.din(w_dff_A_z1MV1RVm5_0),.clk(gclk));
	jdff dff_A_NCvQSvrP0_0(.dout(w_dff_A_31ZmXWPA6_0),.din(w_dff_A_NCvQSvrP0_0),.clk(gclk));
	jdff dff_A_31ZmXWPA6_0(.dout(w_dff_A_rzdzpzl07_0),.din(w_dff_A_31ZmXWPA6_0),.clk(gclk));
	jdff dff_A_rzdzpzl07_0(.dout(w_dff_A_8yCoMCvI6_0),.din(w_dff_A_rzdzpzl07_0),.clk(gclk));
	jdff dff_A_8yCoMCvI6_0(.dout(w_dff_A_YwJr4WJK3_0),.din(w_dff_A_8yCoMCvI6_0),.clk(gclk));
	jdff dff_A_YwJr4WJK3_0(.dout(w_dff_A_Ow12GLnX5_0),.din(w_dff_A_YwJr4WJK3_0),.clk(gclk));
	jdff dff_A_Ow12GLnX5_0(.dout(w_dff_A_BEeT3fNA1_0),.din(w_dff_A_Ow12GLnX5_0),.clk(gclk));
	jdff dff_A_BEeT3fNA1_0(.dout(w_dff_A_258yxaEp7_0),.din(w_dff_A_BEeT3fNA1_0),.clk(gclk));
	jdff dff_A_258yxaEp7_0(.dout(w_dff_A_Bea28Dpj7_0),.din(w_dff_A_258yxaEp7_0),.clk(gclk));
	jdff dff_A_Bea28Dpj7_0(.dout(w_dff_A_gXe7JpOF8_0),.din(w_dff_A_Bea28Dpj7_0),.clk(gclk));
	jdff dff_A_gXe7JpOF8_0(.dout(w_dff_A_rRlDJQLa1_0),.din(w_dff_A_gXe7JpOF8_0),.clk(gclk));
	jdff dff_A_rRlDJQLa1_0(.dout(w_dff_A_jyi9a2ds0_0),.din(w_dff_A_rRlDJQLa1_0),.clk(gclk));
	jdff dff_A_jyi9a2ds0_0(.dout(w_dff_A_AvGh5mxf9_0),.din(w_dff_A_jyi9a2ds0_0),.clk(gclk));
	jdff dff_A_AvGh5mxf9_0(.dout(w_dff_A_DfVOl6jg6_0),.din(w_dff_A_AvGh5mxf9_0),.clk(gclk));
	jdff dff_A_DfVOl6jg6_0(.dout(w_dff_A_W1Q5HWHK8_0),.din(w_dff_A_DfVOl6jg6_0),.clk(gclk));
	jdff dff_A_W1Q5HWHK8_0(.dout(w_dff_A_9QFRuSy82_0),.din(w_dff_A_W1Q5HWHK8_0),.clk(gclk));
	jdff dff_A_9QFRuSy82_0(.dout(w_dff_A_Ljxk9B0y1_0),.din(w_dff_A_9QFRuSy82_0),.clk(gclk));
	jdff dff_A_Ljxk9B0y1_0(.dout(w_dff_A_xkJtNxKY0_0),.din(w_dff_A_Ljxk9B0y1_0),.clk(gclk));
	jdff dff_A_xkJtNxKY0_0(.dout(w_dff_A_RZNQa8Zp0_0),.din(w_dff_A_xkJtNxKY0_0),.clk(gclk));
	jdff dff_A_RZNQa8Zp0_0(.dout(w_dff_A_sAMT18Ip3_0),.din(w_dff_A_RZNQa8Zp0_0),.clk(gclk));
	jdff dff_A_sAMT18Ip3_0(.dout(w_dff_A_FOkR76ml9_0),.din(w_dff_A_sAMT18Ip3_0),.clk(gclk));
	jdff dff_A_FOkR76ml9_0(.dout(w_dff_A_AXurrEUk1_0),.din(w_dff_A_FOkR76ml9_0),.clk(gclk));
	jdff dff_A_AXurrEUk1_0(.dout(w_dff_A_HhopjXlZ5_0),.din(w_dff_A_AXurrEUk1_0),.clk(gclk));
	jdff dff_A_HhopjXlZ5_0(.dout(w_dff_A_EnmNRsPi0_0),.din(w_dff_A_HhopjXlZ5_0),.clk(gclk));
	jdff dff_A_EnmNRsPi0_0(.dout(w_dff_A_dKQThvRv8_0),.din(w_dff_A_EnmNRsPi0_0),.clk(gclk));
	jdff dff_A_dKQThvRv8_0(.dout(G601),.din(w_dff_A_dKQThvRv8_0),.clk(gclk));
	jdff dff_A_FJrUYRUW2_1(.dout(w_dff_A_midEEXwi6_0),.din(w_dff_A_FJrUYRUW2_1),.clk(gclk));
	jdff dff_A_midEEXwi6_0(.dout(w_dff_A_nEvJflSm7_0),.din(w_dff_A_midEEXwi6_0),.clk(gclk));
	jdff dff_A_nEvJflSm7_0(.dout(w_dff_A_SESSf9AI6_0),.din(w_dff_A_nEvJflSm7_0),.clk(gclk));
	jdff dff_A_SESSf9AI6_0(.dout(w_dff_A_YsZvdVsm1_0),.din(w_dff_A_SESSf9AI6_0),.clk(gclk));
	jdff dff_A_YsZvdVsm1_0(.dout(w_dff_A_btPF0H3W0_0),.din(w_dff_A_YsZvdVsm1_0),.clk(gclk));
	jdff dff_A_btPF0H3W0_0(.dout(w_dff_A_M0YggQ760_0),.din(w_dff_A_btPF0H3W0_0),.clk(gclk));
	jdff dff_A_M0YggQ760_0(.dout(w_dff_A_SzLWu1io6_0),.din(w_dff_A_M0YggQ760_0),.clk(gclk));
	jdff dff_A_SzLWu1io6_0(.dout(w_dff_A_dZB7ziFm4_0),.din(w_dff_A_SzLWu1io6_0),.clk(gclk));
	jdff dff_A_dZB7ziFm4_0(.dout(w_dff_A_9XyS5e731_0),.din(w_dff_A_dZB7ziFm4_0),.clk(gclk));
	jdff dff_A_9XyS5e731_0(.dout(w_dff_A_r8lzG5NM2_0),.din(w_dff_A_9XyS5e731_0),.clk(gclk));
	jdff dff_A_r8lzG5NM2_0(.dout(w_dff_A_QPF6Efy87_0),.din(w_dff_A_r8lzG5NM2_0),.clk(gclk));
	jdff dff_A_QPF6Efy87_0(.dout(w_dff_A_sZTpVlYA9_0),.din(w_dff_A_QPF6Efy87_0),.clk(gclk));
	jdff dff_A_sZTpVlYA9_0(.dout(w_dff_A_BNg0veXI8_0),.din(w_dff_A_sZTpVlYA9_0),.clk(gclk));
	jdff dff_A_BNg0veXI8_0(.dout(w_dff_A_FdehvAmM2_0),.din(w_dff_A_BNg0veXI8_0),.clk(gclk));
	jdff dff_A_FdehvAmM2_0(.dout(w_dff_A_fs63tjHV7_0),.din(w_dff_A_FdehvAmM2_0),.clk(gclk));
	jdff dff_A_fs63tjHV7_0(.dout(w_dff_A_nX1Dl57M2_0),.din(w_dff_A_fs63tjHV7_0),.clk(gclk));
	jdff dff_A_nX1Dl57M2_0(.dout(w_dff_A_gtSoiKOo4_0),.din(w_dff_A_nX1Dl57M2_0),.clk(gclk));
	jdff dff_A_gtSoiKOo4_0(.dout(w_dff_A_RMXDH7rG7_0),.din(w_dff_A_gtSoiKOo4_0),.clk(gclk));
	jdff dff_A_RMXDH7rG7_0(.dout(w_dff_A_ymzgro2G8_0),.din(w_dff_A_RMXDH7rG7_0),.clk(gclk));
	jdff dff_A_ymzgro2G8_0(.dout(w_dff_A_eCLMDY9V5_0),.din(w_dff_A_ymzgro2G8_0),.clk(gclk));
	jdff dff_A_eCLMDY9V5_0(.dout(w_dff_A_JmltyGqX9_0),.din(w_dff_A_eCLMDY9V5_0),.clk(gclk));
	jdff dff_A_JmltyGqX9_0(.dout(w_dff_A_zrdcGyY85_0),.din(w_dff_A_JmltyGqX9_0),.clk(gclk));
	jdff dff_A_zrdcGyY85_0(.dout(w_dff_A_LRXr5ju66_0),.din(w_dff_A_zrdcGyY85_0),.clk(gclk));
	jdff dff_A_LRXr5ju66_0(.dout(w_dff_A_VhDntoKw5_0),.din(w_dff_A_LRXr5ju66_0),.clk(gclk));
	jdff dff_A_VhDntoKw5_0(.dout(w_dff_A_oGAw2bVZ4_0),.din(w_dff_A_VhDntoKw5_0),.clk(gclk));
	jdff dff_A_oGAw2bVZ4_0(.dout(w_dff_A_zYPLqGsr8_0),.din(w_dff_A_oGAw2bVZ4_0),.clk(gclk));
	jdff dff_A_zYPLqGsr8_0(.dout(G602),.din(w_dff_A_zYPLqGsr8_0),.clk(gclk));
	jdff dff_A_hsW6rtkC8_1(.dout(w_dff_A_szKiCzJS1_0),.din(w_dff_A_hsW6rtkC8_1),.clk(gclk));
	jdff dff_A_szKiCzJS1_0(.dout(w_dff_A_yJBiMRC79_0),.din(w_dff_A_szKiCzJS1_0),.clk(gclk));
	jdff dff_A_yJBiMRC79_0(.dout(w_dff_A_Z9VSso8D1_0),.din(w_dff_A_yJBiMRC79_0),.clk(gclk));
	jdff dff_A_Z9VSso8D1_0(.dout(w_dff_A_gZdKDqab3_0),.din(w_dff_A_Z9VSso8D1_0),.clk(gclk));
	jdff dff_A_gZdKDqab3_0(.dout(w_dff_A_9RZ0kxKC1_0),.din(w_dff_A_gZdKDqab3_0),.clk(gclk));
	jdff dff_A_9RZ0kxKC1_0(.dout(w_dff_A_Tf7IENfH1_0),.din(w_dff_A_9RZ0kxKC1_0),.clk(gclk));
	jdff dff_A_Tf7IENfH1_0(.dout(w_dff_A_6c6RHEE55_0),.din(w_dff_A_Tf7IENfH1_0),.clk(gclk));
	jdff dff_A_6c6RHEE55_0(.dout(w_dff_A_Cj9JVRMP3_0),.din(w_dff_A_6c6RHEE55_0),.clk(gclk));
	jdff dff_A_Cj9JVRMP3_0(.dout(w_dff_A_TWAnU5KB2_0),.din(w_dff_A_Cj9JVRMP3_0),.clk(gclk));
	jdff dff_A_TWAnU5KB2_0(.dout(w_dff_A_EYi4WWD14_0),.din(w_dff_A_TWAnU5KB2_0),.clk(gclk));
	jdff dff_A_EYi4WWD14_0(.dout(w_dff_A_Jv1Yxix80_0),.din(w_dff_A_EYi4WWD14_0),.clk(gclk));
	jdff dff_A_Jv1Yxix80_0(.dout(w_dff_A_GezRUYTJ9_0),.din(w_dff_A_Jv1Yxix80_0),.clk(gclk));
	jdff dff_A_GezRUYTJ9_0(.dout(w_dff_A_IbrxoSpm7_0),.din(w_dff_A_GezRUYTJ9_0),.clk(gclk));
	jdff dff_A_IbrxoSpm7_0(.dout(w_dff_A_ruY906Ta4_0),.din(w_dff_A_IbrxoSpm7_0),.clk(gclk));
	jdff dff_A_ruY906Ta4_0(.dout(w_dff_A_irFwQcnP4_0),.din(w_dff_A_ruY906Ta4_0),.clk(gclk));
	jdff dff_A_irFwQcnP4_0(.dout(w_dff_A_OuKPEvKB0_0),.din(w_dff_A_irFwQcnP4_0),.clk(gclk));
	jdff dff_A_OuKPEvKB0_0(.dout(w_dff_A_7c4ZfVoG7_0),.din(w_dff_A_OuKPEvKB0_0),.clk(gclk));
	jdff dff_A_7c4ZfVoG7_0(.dout(w_dff_A_N3TJd7Gp5_0),.din(w_dff_A_7c4ZfVoG7_0),.clk(gclk));
	jdff dff_A_N3TJd7Gp5_0(.dout(w_dff_A_tgloV8av7_0),.din(w_dff_A_N3TJd7Gp5_0),.clk(gclk));
	jdff dff_A_tgloV8av7_0(.dout(w_dff_A_Xets2Obk2_0),.din(w_dff_A_tgloV8av7_0),.clk(gclk));
	jdff dff_A_Xets2Obk2_0(.dout(w_dff_A_RKyVqdFx5_0),.din(w_dff_A_Xets2Obk2_0),.clk(gclk));
	jdff dff_A_RKyVqdFx5_0(.dout(w_dff_A_eXir635X9_0),.din(w_dff_A_RKyVqdFx5_0),.clk(gclk));
	jdff dff_A_eXir635X9_0(.dout(w_dff_A_KPIQcHyP7_0),.din(w_dff_A_eXir635X9_0),.clk(gclk));
	jdff dff_A_KPIQcHyP7_0(.dout(w_dff_A_pdkIhO8J0_0),.din(w_dff_A_KPIQcHyP7_0),.clk(gclk));
	jdff dff_A_pdkIhO8J0_0(.dout(w_dff_A_GNYTEDO03_0),.din(w_dff_A_pdkIhO8J0_0),.clk(gclk));
	jdff dff_A_GNYTEDO03_0(.dout(w_dff_A_I2luZ5AD4_0),.din(w_dff_A_GNYTEDO03_0),.clk(gclk));
	jdff dff_A_I2luZ5AD4_0(.dout(G603),.din(w_dff_A_I2luZ5AD4_0),.clk(gclk));
	jdff dff_A_PX3V940Q1_1(.dout(w_dff_A_Szlr61vU3_0),.din(w_dff_A_PX3V940Q1_1),.clk(gclk));
	jdff dff_A_Szlr61vU3_0(.dout(w_dff_A_txxwIzN43_0),.din(w_dff_A_Szlr61vU3_0),.clk(gclk));
	jdff dff_A_txxwIzN43_0(.dout(w_dff_A_TcaYo2gG9_0),.din(w_dff_A_txxwIzN43_0),.clk(gclk));
	jdff dff_A_TcaYo2gG9_0(.dout(w_dff_A_JhxAfswL4_0),.din(w_dff_A_TcaYo2gG9_0),.clk(gclk));
	jdff dff_A_JhxAfswL4_0(.dout(w_dff_A_57InIhXx1_0),.din(w_dff_A_JhxAfswL4_0),.clk(gclk));
	jdff dff_A_57InIhXx1_0(.dout(w_dff_A_qYmlp08P4_0),.din(w_dff_A_57InIhXx1_0),.clk(gclk));
	jdff dff_A_qYmlp08P4_0(.dout(w_dff_A_xxcY15o56_0),.din(w_dff_A_qYmlp08P4_0),.clk(gclk));
	jdff dff_A_xxcY15o56_0(.dout(w_dff_A_SyNuU87b4_0),.din(w_dff_A_xxcY15o56_0),.clk(gclk));
	jdff dff_A_SyNuU87b4_0(.dout(w_dff_A_3axgsdQM0_0),.din(w_dff_A_SyNuU87b4_0),.clk(gclk));
	jdff dff_A_3axgsdQM0_0(.dout(w_dff_A_CHWLo9YL9_0),.din(w_dff_A_3axgsdQM0_0),.clk(gclk));
	jdff dff_A_CHWLo9YL9_0(.dout(w_dff_A_w6Npeprv7_0),.din(w_dff_A_CHWLo9YL9_0),.clk(gclk));
	jdff dff_A_w6Npeprv7_0(.dout(w_dff_A_iA6SLOYw2_0),.din(w_dff_A_w6Npeprv7_0),.clk(gclk));
	jdff dff_A_iA6SLOYw2_0(.dout(w_dff_A_VpihWe7C8_0),.din(w_dff_A_iA6SLOYw2_0),.clk(gclk));
	jdff dff_A_VpihWe7C8_0(.dout(w_dff_A_vmXYj26E5_0),.din(w_dff_A_VpihWe7C8_0),.clk(gclk));
	jdff dff_A_vmXYj26E5_0(.dout(w_dff_A_Wj1A375y5_0),.din(w_dff_A_vmXYj26E5_0),.clk(gclk));
	jdff dff_A_Wj1A375y5_0(.dout(w_dff_A_oUPPLDIT1_0),.din(w_dff_A_Wj1A375y5_0),.clk(gclk));
	jdff dff_A_oUPPLDIT1_0(.dout(w_dff_A_fFCFGCtw3_0),.din(w_dff_A_oUPPLDIT1_0),.clk(gclk));
	jdff dff_A_fFCFGCtw3_0(.dout(w_dff_A_gxbjnoIh6_0),.din(w_dff_A_fFCFGCtw3_0),.clk(gclk));
	jdff dff_A_gxbjnoIh6_0(.dout(w_dff_A_40w87G6r0_0),.din(w_dff_A_gxbjnoIh6_0),.clk(gclk));
	jdff dff_A_40w87G6r0_0(.dout(w_dff_A_7Nczw42J7_0),.din(w_dff_A_40w87G6r0_0),.clk(gclk));
	jdff dff_A_7Nczw42J7_0(.dout(w_dff_A_bjmRyeJX8_0),.din(w_dff_A_7Nczw42J7_0),.clk(gclk));
	jdff dff_A_bjmRyeJX8_0(.dout(w_dff_A_D3aERHvU1_0),.din(w_dff_A_bjmRyeJX8_0),.clk(gclk));
	jdff dff_A_D3aERHvU1_0(.dout(w_dff_A_tsTZTo0n4_0),.din(w_dff_A_D3aERHvU1_0),.clk(gclk));
	jdff dff_A_tsTZTo0n4_0(.dout(w_dff_A_eOrHbXe88_0),.din(w_dff_A_tsTZTo0n4_0),.clk(gclk));
	jdff dff_A_eOrHbXe88_0(.dout(w_dff_A_bmPpN7js2_0),.din(w_dff_A_eOrHbXe88_0),.clk(gclk));
	jdff dff_A_bmPpN7js2_0(.dout(w_dff_A_jf8spJsC9_0),.din(w_dff_A_bmPpN7js2_0),.clk(gclk));
	jdff dff_A_jf8spJsC9_0(.dout(G604),.din(w_dff_A_jf8spJsC9_0),.clk(gclk));
	jdff dff_A_FpfbrbRf3_1(.dout(w_dff_A_hWBhh0uA5_0),.din(w_dff_A_FpfbrbRf3_1),.clk(gclk));
	jdff dff_A_hWBhh0uA5_0(.dout(w_dff_A_DF2pDixM4_0),.din(w_dff_A_hWBhh0uA5_0),.clk(gclk));
	jdff dff_A_DF2pDixM4_0(.dout(w_dff_A_uuuBjRoR1_0),.din(w_dff_A_DF2pDixM4_0),.clk(gclk));
	jdff dff_A_uuuBjRoR1_0(.dout(w_dff_A_WohuxkYd2_0),.din(w_dff_A_uuuBjRoR1_0),.clk(gclk));
	jdff dff_A_WohuxkYd2_0(.dout(w_dff_A_Ir2xvp0x1_0),.din(w_dff_A_WohuxkYd2_0),.clk(gclk));
	jdff dff_A_Ir2xvp0x1_0(.dout(w_dff_A_afzONmUh7_0),.din(w_dff_A_Ir2xvp0x1_0),.clk(gclk));
	jdff dff_A_afzONmUh7_0(.dout(w_dff_A_jKnjhFfZ6_0),.din(w_dff_A_afzONmUh7_0),.clk(gclk));
	jdff dff_A_jKnjhFfZ6_0(.dout(w_dff_A_YS4lJjbE0_0),.din(w_dff_A_jKnjhFfZ6_0),.clk(gclk));
	jdff dff_A_YS4lJjbE0_0(.dout(w_dff_A_sV06MLaO8_0),.din(w_dff_A_YS4lJjbE0_0),.clk(gclk));
	jdff dff_A_sV06MLaO8_0(.dout(w_dff_A_8K2SK2cJ2_0),.din(w_dff_A_sV06MLaO8_0),.clk(gclk));
	jdff dff_A_8K2SK2cJ2_0(.dout(w_dff_A_YJ15L2IW5_0),.din(w_dff_A_8K2SK2cJ2_0),.clk(gclk));
	jdff dff_A_YJ15L2IW5_0(.dout(w_dff_A_PkL00IS48_0),.din(w_dff_A_YJ15L2IW5_0),.clk(gclk));
	jdff dff_A_PkL00IS48_0(.dout(w_dff_A_gBzSJv3r7_0),.din(w_dff_A_PkL00IS48_0),.clk(gclk));
	jdff dff_A_gBzSJv3r7_0(.dout(w_dff_A_BVzplejU9_0),.din(w_dff_A_gBzSJv3r7_0),.clk(gclk));
	jdff dff_A_BVzplejU9_0(.dout(w_dff_A_Zj3TXxVz6_0),.din(w_dff_A_BVzplejU9_0),.clk(gclk));
	jdff dff_A_Zj3TXxVz6_0(.dout(w_dff_A_tsCG02bx4_0),.din(w_dff_A_Zj3TXxVz6_0),.clk(gclk));
	jdff dff_A_tsCG02bx4_0(.dout(w_dff_A_D1O1SYim5_0),.din(w_dff_A_tsCG02bx4_0),.clk(gclk));
	jdff dff_A_D1O1SYim5_0(.dout(w_dff_A_HGvRUoVW5_0),.din(w_dff_A_D1O1SYim5_0),.clk(gclk));
	jdff dff_A_HGvRUoVW5_0(.dout(w_dff_A_cSJqokbd4_0),.din(w_dff_A_HGvRUoVW5_0),.clk(gclk));
	jdff dff_A_cSJqokbd4_0(.dout(w_dff_A_nwWD9v3C3_0),.din(w_dff_A_cSJqokbd4_0),.clk(gclk));
	jdff dff_A_nwWD9v3C3_0(.dout(w_dff_A_9P9q7ot19_0),.din(w_dff_A_nwWD9v3C3_0),.clk(gclk));
	jdff dff_A_9P9q7ot19_0(.dout(w_dff_A_QSwPkL6k4_0),.din(w_dff_A_9P9q7ot19_0),.clk(gclk));
	jdff dff_A_QSwPkL6k4_0(.dout(w_dff_A_eo6KGMVz7_0),.din(w_dff_A_QSwPkL6k4_0),.clk(gclk));
	jdff dff_A_eo6KGMVz7_0(.dout(w_dff_A_3prTw2Z20_0),.din(w_dff_A_eo6KGMVz7_0),.clk(gclk));
	jdff dff_A_3prTw2Z20_0(.dout(w_dff_A_ZyehewfO2_0),.din(w_dff_A_3prTw2Z20_0),.clk(gclk));
	jdff dff_A_ZyehewfO2_0(.dout(w_dff_A_nCxU7v4v1_0),.din(w_dff_A_ZyehewfO2_0),.clk(gclk));
	jdff dff_A_nCxU7v4v1_0(.dout(G611),.din(w_dff_A_nCxU7v4v1_0),.clk(gclk));
	jdff dff_A_ngtpAtsY5_1(.dout(w_dff_A_dI8qiuRa9_0),.din(w_dff_A_ngtpAtsY5_1),.clk(gclk));
	jdff dff_A_dI8qiuRa9_0(.dout(w_dff_A_XS6ojzl56_0),.din(w_dff_A_dI8qiuRa9_0),.clk(gclk));
	jdff dff_A_XS6ojzl56_0(.dout(w_dff_A_pSpZeeOU2_0),.din(w_dff_A_XS6ojzl56_0),.clk(gclk));
	jdff dff_A_pSpZeeOU2_0(.dout(w_dff_A_xfaVxp8y8_0),.din(w_dff_A_pSpZeeOU2_0),.clk(gclk));
	jdff dff_A_xfaVxp8y8_0(.dout(w_dff_A_SQJ3DB1P9_0),.din(w_dff_A_xfaVxp8y8_0),.clk(gclk));
	jdff dff_A_SQJ3DB1P9_0(.dout(w_dff_A_uzOI3sGp8_0),.din(w_dff_A_SQJ3DB1P9_0),.clk(gclk));
	jdff dff_A_uzOI3sGp8_0(.dout(w_dff_A_p3Xx526u7_0),.din(w_dff_A_uzOI3sGp8_0),.clk(gclk));
	jdff dff_A_p3Xx526u7_0(.dout(w_dff_A_WV6L8kQ13_0),.din(w_dff_A_p3Xx526u7_0),.clk(gclk));
	jdff dff_A_WV6L8kQ13_0(.dout(w_dff_A_uexmfjaw3_0),.din(w_dff_A_WV6L8kQ13_0),.clk(gclk));
	jdff dff_A_uexmfjaw3_0(.dout(w_dff_A_9MXOBaWj9_0),.din(w_dff_A_uexmfjaw3_0),.clk(gclk));
	jdff dff_A_9MXOBaWj9_0(.dout(w_dff_A_I8JayFcY4_0),.din(w_dff_A_9MXOBaWj9_0),.clk(gclk));
	jdff dff_A_I8JayFcY4_0(.dout(w_dff_A_PAx9P8q05_0),.din(w_dff_A_I8JayFcY4_0),.clk(gclk));
	jdff dff_A_PAx9P8q05_0(.dout(w_dff_A_4DQmtHqt2_0),.din(w_dff_A_PAx9P8q05_0),.clk(gclk));
	jdff dff_A_4DQmtHqt2_0(.dout(w_dff_A_88KhvHXC0_0),.din(w_dff_A_4DQmtHqt2_0),.clk(gclk));
	jdff dff_A_88KhvHXC0_0(.dout(w_dff_A_50UI5PGD0_0),.din(w_dff_A_88KhvHXC0_0),.clk(gclk));
	jdff dff_A_50UI5PGD0_0(.dout(w_dff_A_GkKeEPc17_0),.din(w_dff_A_50UI5PGD0_0),.clk(gclk));
	jdff dff_A_GkKeEPc17_0(.dout(w_dff_A_vLElKZTm0_0),.din(w_dff_A_GkKeEPc17_0),.clk(gclk));
	jdff dff_A_vLElKZTm0_0(.dout(w_dff_A_HBHEkfUe2_0),.din(w_dff_A_vLElKZTm0_0),.clk(gclk));
	jdff dff_A_HBHEkfUe2_0(.dout(w_dff_A_uCqDNxO10_0),.din(w_dff_A_HBHEkfUe2_0),.clk(gclk));
	jdff dff_A_uCqDNxO10_0(.dout(w_dff_A_QRwZmUjI4_0),.din(w_dff_A_uCqDNxO10_0),.clk(gclk));
	jdff dff_A_QRwZmUjI4_0(.dout(w_dff_A_chnGNUjU5_0),.din(w_dff_A_QRwZmUjI4_0),.clk(gclk));
	jdff dff_A_chnGNUjU5_0(.dout(w_dff_A_2GV3F85s8_0),.din(w_dff_A_chnGNUjU5_0),.clk(gclk));
	jdff dff_A_2GV3F85s8_0(.dout(w_dff_A_dnBudaaR9_0),.din(w_dff_A_2GV3F85s8_0),.clk(gclk));
	jdff dff_A_dnBudaaR9_0(.dout(w_dff_A_ZQ8Rg5qF5_0),.din(w_dff_A_dnBudaaR9_0),.clk(gclk));
	jdff dff_A_ZQ8Rg5qF5_0(.dout(w_dff_A_lq9Bm5JV2_0),.din(w_dff_A_ZQ8Rg5qF5_0),.clk(gclk));
	jdff dff_A_lq9Bm5JV2_0(.dout(w_dff_A_9T2mPAHf9_0),.din(w_dff_A_lq9Bm5JV2_0),.clk(gclk));
	jdff dff_A_9T2mPAHf9_0(.dout(G612),.din(w_dff_A_9T2mPAHf9_0),.clk(gclk));
	jdff dff_A_5cfRan3F4_2(.dout(w_dff_A_TNeGIopd8_0),.din(w_dff_A_5cfRan3F4_2),.clk(gclk));
	jdff dff_A_TNeGIopd8_0(.dout(w_dff_A_cliTpmkT3_0),.din(w_dff_A_TNeGIopd8_0),.clk(gclk));
	jdff dff_A_cliTpmkT3_0(.dout(w_dff_A_DcGSxjqq2_0),.din(w_dff_A_cliTpmkT3_0),.clk(gclk));
	jdff dff_A_DcGSxjqq2_0(.dout(w_dff_A_FV1UWYjJ3_0),.din(w_dff_A_DcGSxjqq2_0),.clk(gclk));
	jdff dff_A_FV1UWYjJ3_0(.dout(w_dff_A_QhuGMRpv6_0),.din(w_dff_A_FV1UWYjJ3_0),.clk(gclk));
	jdff dff_A_QhuGMRpv6_0(.dout(w_dff_A_gvTpK0tC8_0),.din(w_dff_A_QhuGMRpv6_0),.clk(gclk));
	jdff dff_A_gvTpK0tC8_0(.dout(w_dff_A_fSPPQFY42_0),.din(w_dff_A_gvTpK0tC8_0),.clk(gclk));
	jdff dff_A_fSPPQFY42_0(.dout(w_dff_A_C8pYUjey9_0),.din(w_dff_A_fSPPQFY42_0),.clk(gclk));
	jdff dff_A_C8pYUjey9_0(.dout(w_dff_A_Dq5SKNWG6_0),.din(w_dff_A_C8pYUjey9_0),.clk(gclk));
	jdff dff_A_Dq5SKNWG6_0(.dout(w_dff_A_5Qp6DBuz4_0),.din(w_dff_A_Dq5SKNWG6_0),.clk(gclk));
	jdff dff_A_5Qp6DBuz4_0(.dout(w_dff_A_IYpkiHMX6_0),.din(w_dff_A_5Qp6DBuz4_0),.clk(gclk));
	jdff dff_A_IYpkiHMX6_0(.dout(w_dff_A_WWeMLzkC5_0),.din(w_dff_A_IYpkiHMX6_0),.clk(gclk));
	jdff dff_A_WWeMLzkC5_0(.dout(w_dff_A_6bTjRrRU4_0),.din(w_dff_A_WWeMLzkC5_0),.clk(gclk));
	jdff dff_A_6bTjRrRU4_0(.dout(w_dff_A_MYVkEitD8_0),.din(w_dff_A_6bTjRrRU4_0),.clk(gclk));
	jdff dff_A_MYVkEitD8_0(.dout(w_dff_A_cSWIX6eW9_0),.din(w_dff_A_MYVkEitD8_0),.clk(gclk));
	jdff dff_A_cSWIX6eW9_0(.dout(w_dff_A_KGf7Iqt45_0),.din(w_dff_A_cSWIX6eW9_0),.clk(gclk));
	jdff dff_A_KGf7Iqt45_0(.dout(w_dff_A_FoV0X4GM5_0),.din(w_dff_A_KGf7Iqt45_0),.clk(gclk));
	jdff dff_A_FoV0X4GM5_0(.dout(w_dff_A_Bty9xsM37_0),.din(w_dff_A_FoV0X4GM5_0),.clk(gclk));
	jdff dff_A_Bty9xsM37_0(.dout(w_dff_A_JufoRDEz4_0),.din(w_dff_A_Bty9xsM37_0),.clk(gclk));
	jdff dff_A_JufoRDEz4_0(.dout(w_dff_A_uk2DcbNv8_0),.din(w_dff_A_JufoRDEz4_0),.clk(gclk));
	jdff dff_A_uk2DcbNv8_0(.dout(w_dff_A_3RmbsgOM2_0),.din(w_dff_A_uk2DcbNv8_0),.clk(gclk));
	jdff dff_A_3RmbsgOM2_0(.dout(w_dff_A_soGFIDx60_0),.din(w_dff_A_3RmbsgOM2_0),.clk(gclk));
	jdff dff_A_soGFIDx60_0(.dout(w_dff_A_0Asvl05L1_0),.din(w_dff_A_soGFIDx60_0),.clk(gclk));
	jdff dff_A_0Asvl05L1_0(.dout(w_dff_A_vG3AJPai3_0),.din(w_dff_A_0Asvl05L1_0),.clk(gclk));
	jdff dff_A_vG3AJPai3_0(.dout(w_dff_A_2VOakzUt5_0),.din(w_dff_A_vG3AJPai3_0),.clk(gclk));
	jdff dff_A_2VOakzUt5_0(.dout(w_dff_A_mJOSM8RJ0_0),.din(w_dff_A_2VOakzUt5_0),.clk(gclk));
	jdff dff_A_mJOSM8RJ0_0(.dout(G810),.din(w_dff_A_mJOSM8RJ0_0),.clk(gclk));
	jdff dff_A_5t6DzlqV5_1(.dout(w_dff_A_AkO6TqAN1_0),.din(w_dff_A_5t6DzlqV5_1),.clk(gclk));
	jdff dff_A_AkO6TqAN1_0(.dout(w_dff_A_0fViiNHk7_0),.din(w_dff_A_AkO6TqAN1_0),.clk(gclk));
	jdff dff_A_0fViiNHk7_0(.dout(w_dff_A_KMSQqxDl9_0),.din(w_dff_A_0fViiNHk7_0),.clk(gclk));
	jdff dff_A_KMSQqxDl9_0(.dout(w_dff_A_ClQuB2hj4_0),.din(w_dff_A_KMSQqxDl9_0),.clk(gclk));
	jdff dff_A_ClQuB2hj4_0(.dout(w_dff_A_56vSMsC89_0),.din(w_dff_A_ClQuB2hj4_0),.clk(gclk));
	jdff dff_A_56vSMsC89_0(.dout(w_dff_A_GGQcJnL39_0),.din(w_dff_A_56vSMsC89_0),.clk(gclk));
	jdff dff_A_GGQcJnL39_0(.dout(w_dff_A_Ek0i76k61_0),.din(w_dff_A_GGQcJnL39_0),.clk(gclk));
	jdff dff_A_Ek0i76k61_0(.dout(w_dff_A_blfsYTeX7_0),.din(w_dff_A_Ek0i76k61_0),.clk(gclk));
	jdff dff_A_blfsYTeX7_0(.dout(w_dff_A_SSTP5gav9_0),.din(w_dff_A_blfsYTeX7_0),.clk(gclk));
	jdff dff_A_SSTP5gav9_0(.dout(w_dff_A_IUJH1Rzh6_0),.din(w_dff_A_SSTP5gav9_0),.clk(gclk));
	jdff dff_A_IUJH1Rzh6_0(.dout(w_dff_A_UnpMCpFA6_0),.din(w_dff_A_IUJH1Rzh6_0),.clk(gclk));
	jdff dff_A_UnpMCpFA6_0(.dout(w_dff_A_toLzv5Wz8_0),.din(w_dff_A_UnpMCpFA6_0),.clk(gclk));
	jdff dff_A_toLzv5Wz8_0(.dout(w_dff_A_9cBlObww6_0),.din(w_dff_A_toLzv5Wz8_0),.clk(gclk));
	jdff dff_A_9cBlObww6_0(.dout(w_dff_A_rZeDuzOa5_0),.din(w_dff_A_9cBlObww6_0),.clk(gclk));
	jdff dff_A_rZeDuzOa5_0(.dout(w_dff_A_jzQ6eMdj7_0),.din(w_dff_A_rZeDuzOa5_0),.clk(gclk));
	jdff dff_A_jzQ6eMdj7_0(.dout(w_dff_A_DjBUioum9_0),.din(w_dff_A_jzQ6eMdj7_0),.clk(gclk));
	jdff dff_A_DjBUioum9_0(.dout(w_dff_A_CxweOoky9_0),.din(w_dff_A_DjBUioum9_0),.clk(gclk));
	jdff dff_A_CxweOoky9_0(.dout(w_dff_A_bkcEcDCz8_0),.din(w_dff_A_CxweOoky9_0),.clk(gclk));
	jdff dff_A_bkcEcDCz8_0(.dout(w_dff_A_Cp66eVQd7_0),.din(w_dff_A_bkcEcDCz8_0),.clk(gclk));
	jdff dff_A_Cp66eVQd7_0(.dout(w_dff_A_eljnh0Zq4_0),.din(w_dff_A_Cp66eVQd7_0),.clk(gclk));
	jdff dff_A_eljnh0Zq4_0(.dout(w_dff_A_dWtolInX2_0),.din(w_dff_A_eljnh0Zq4_0),.clk(gclk));
	jdff dff_A_dWtolInX2_0(.dout(w_dff_A_J9jSSohA0_0),.din(w_dff_A_dWtolInX2_0),.clk(gclk));
	jdff dff_A_J9jSSohA0_0(.dout(w_dff_A_AzGZECcC4_0),.din(w_dff_A_J9jSSohA0_0),.clk(gclk));
	jdff dff_A_AzGZECcC4_0(.dout(w_dff_A_s23nZGQS9_0),.din(w_dff_A_AzGZECcC4_0),.clk(gclk));
	jdff dff_A_s23nZGQS9_0(.dout(w_dff_A_TtBkZVw68_0),.din(w_dff_A_s23nZGQS9_0),.clk(gclk));
	jdff dff_A_TtBkZVw68_0(.dout(w_dff_A_oLgyeFaj7_0),.din(w_dff_A_TtBkZVw68_0),.clk(gclk));
	jdff dff_A_oLgyeFaj7_0(.dout(G848),.din(w_dff_A_oLgyeFaj7_0),.clk(gclk));
	jdff dff_A_WU84By202_1(.dout(w_dff_A_ExbZdFft7_0),.din(w_dff_A_WU84By202_1),.clk(gclk));
	jdff dff_A_ExbZdFft7_0(.dout(w_dff_A_LipODtBL2_0),.din(w_dff_A_ExbZdFft7_0),.clk(gclk));
	jdff dff_A_LipODtBL2_0(.dout(w_dff_A_IP95x7VF3_0),.din(w_dff_A_LipODtBL2_0),.clk(gclk));
	jdff dff_A_IP95x7VF3_0(.dout(w_dff_A_ohwzvEnL0_0),.din(w_dff_A_IP95x7VF3_0),.clk(gclk));
	jdff dff_A_ohwzvEnL0_0(.dout(w_dff_A_wRzVTGBz1_0),.din(w_dff_A_ohwzvEnL0_0),.clk(gclk));
	jdff dff_A_wRzVTGBz1_0(.dout(w_dff_A_M1J9ofQx9_0),.din(w_dff_A_wRzVTGBz1_0),.clk(gclk));
	jdff dff_A_M1J9ofQx9_0(.dout(w_dff_A_XxZuVF487_0),.din(w_dff_A_M1J9ofQx9_0),.clk(gclk));
	jdff dff_A_XxZuVF487_0(.dout(w_dff_A_8CmjZnUN6_0),.din(w_dff_A_XxZuVF487_0),.clk(gclk));
	jdff dff_A_8CmjZnUN6_0(.dout(w_dff_A_en6iky532_0),.din(w_dff_A_8CmjZnUN6_0),.clk(gclk));
	jdff dff_A_en6iky532_0(.dout(w_dff_A_vdY2E7GL0_0),.din(w_dff_A_en6iky532_0),.clk(gclk));
	jdff dff_A_vdY2E7GL0_0(.dout(w_dff_A_8c4tUJNl4_0),.din(w_dff_A_vdY2E7GL0_0),.clk(gclk));
	jdff dff_A_8c4tUJNl4_0(.dout(w_dff_A_9s12XcWn3_0),.din(w_dff_A_8c4tUJNl4_0),.clk(gclk));
	jdff dff_A_9s12XcWn3_0(.dout(w_dff_A_hKg7IygA9_0),.din(w_dff_A_9s12XcWn3_0),.clk(gclk));
	jdff dff_A_hKg7IygA9_0(.dout(w_dff_A_KaKR3Fko9_0),.din(w_dff_A_hKg7IygA9_0),.clk(gclk));
	jdff dff_A_KaKR3Fko9_0(.dout(w_dff_A_Dr8oBaGF7_0),.din(w_dff_A_KaKR3Fko9_0),.clk(gclk));
	jdff dff_A_Dr8oBaGF7_0(.dout(w_dff_A_SzQjdAPg7_0),.din(w_dff_A_Dr8oBaGF7_0),.clk(gclk));
	jdff dff_A_SzQjdAPg7_0(.dout(w_dff_A_WIXvc3nZ4_0),.din(w_dff_A_SzQjdAPg7_0),.clk(gclk));
	jdff dff_A_WIXvc3nZ4_0(.dout(w_dff_A_be6sH0uC5_0),.din(w_dff_A_WIXvc3nZ4_0),.clk(gclk));
	jdff dff_A_be6sH0uC5_0(.dout(w_dff_A_2dfySpkn9_0),.din(w_dff_A_be6sH0uC5_0),.clk(gclk));
	jdff dff_A_2dfySpkn9_0(.dout(w_dff_A_x9n3u7oK2_0),.din(w_dff_A_2dfySpkn9_0),.clk(gclk));
	jdff dff_A_x9n3u7oK2_0(.dout(w_dff_A_y55xJ1ku5_0),.din(w_dff_A_x9n3u7oK2_0),.clk(gclk));
	jdff dff_A_y55xJ1ku5_0(.dout(w_dff_A_Bdq7bNDo0_0),.din(w_dff_A_y55xJ1ku5_0),.clk(gclk));
	jdff dff_A_Bdq7bNDo0_0(.dout(w_dff_A_7M6NhEP52_0),.din(w_dff_A_Bdq7bNDo0_0),.clk(gclk));
	jdff dff_A_7M6NhEP52_0(.dout(w_dff_A_k2LO6yXs7_0),.din(w_dff_A_7M6NhEP52_0),.clk(gclk));
	jdff dff_A_k2LO6yXs7_0(.dout(w_dff_A_M83EPBTI6_0),.din(w_dff_A_k2LO6yXs7_0),.clk(gclk));
	jdff dff_A_M83EPBTI6_0(.dout(w_dff_A_ZVtp3RYb3_0),.din(w_dff_A_M83EPBTI6_0),.clk(gclk));
	jdff dff_A_ZVtp3RYb3_0(.dout(G849),.din(w_dff_A_ZVtp3RYb3_0),.clk(gclk));
	jdff dff_A_00yBnyGB8_1(.dout(w_dff_A_UDlJXt8c6_0),.din(w_dff_A_00yBnyGB8_1),.clk(gclk));
	jdff dff_A_UDlJXt8c6_0(.dout(w_dff_A_LMDyBa0b8_0),.din(w_dff_A_UDlJXt8c6_0),.clk(gclk));
	jdff dff_A_LMDyBa0b8_0(.dout(w_dff_A_JjWo0d4c7_0),.din(w_dff_A_LMDyBa0b8_0),.clk(gclk));
	jdff dff_A_JjWo0d4c7_0(.dout(w_dff_A_seqQ42bY6_0),.din(w_dff_A_JjWo0d4c7_0),.clk(gclk));
	jdff dff_A_seqQ42bY6_0(.dout(w_dff_A_9PjKnYGS6_0),.din(w_dff_A_seqQ42bY6_0),.clk(gclk));
	jdff dff_A_9PjKnYGS6_0(.dout(w_dff_A_6NSocSQc1_0),.din(w_dff_A_9PjKnYGS6_0),.clk(gclk));
	jdff dff_A_6NSocSQc1_0(.dout(w_dff_A_VogwunOA4_0),.din(w_dff_A_6NSocSQc1_0),.clk(gclk));
	jdff dff_A_VogwunOA4_0(.dout(w_dff_A_RWtZAbBh4_0),.din(w_dff_A_VogwunOA4_0),.clk(gclk));
	jdff dff_A_RWtZAbBh4_0(.dout(w_dff_A_3umFCYI50_0),.din(w_dff_A_RWtZAbBh4_0),.clk(gclk));
	jdff dff_A_3umFCYI50_0(.dout(w_dff_A_TnSQms2s5_0),.din(w_dff_A_3umFCYI50_0),.clk(gclk));
	jdff dff_A_TnSQms2s5_0(.dout(w_dff_A_m0PwIy8J4_0),.din(w_dff_A_TnSQms2s5_0),.clk(gclk));
	jdff dff_A_m0PwIy8J4_0(.dout(w_dff_A_zxzhDAm66_0),.din(w_dff_A_m0PwIy8J4_0),.clk(gclk));
	jdff dff_A_zxzhDAm66_0(.dout(w_dff_A_h6FErAJP6_0),.din(w_dff_A_zxzhDAm66_0),.clk(gclk));
	jdff dff_A_h6FErAJP6_0(.dout(w_dff_A_Vex5MC0l7_0),.din(w_dff_A_h6FErAJP6_0),.clk(gclk));
	jdff dff_A_Vex5MC0l7_0(.dout(w_dff_A_7AhQ1E7u2_0),.din(w_dff_A_Vex5MC0l7_0),.clk(gclk));
	jdff dff_A_7AhQ1E7u2_0(.dout(w_dff_A_3zbwA3tH1_0),.din(w_dff_A_7AhQ1E7u2_0),.clk(gclk));
	jdff dff_A_3zbwA3tH1_0(.dout(w_dff_A_ynQ30shl7_0),.din(w_dff_A_3zbwA3tH1_0),.clk(gclk));
	jdff dff_A_ynQ30shl7_0(.dout(w_dff_A_NbYM2WC09_0),.din(w_dff_A_ynQ30shl7_0),.clk(gclk));
	jdff dff_A_NbYM2WC09_0(.dout(w_dff_A_yPhRucby9_0),.din(w_dff_A_NbYM2WC09_0),.clk(gclk));
	jdff dff_A_yPhRucby9_0(.dout(w_dff_A_g9U8ADko8_0),.din(w_dff_A_yPhRucby9_0),.clk(gclk));
	jdff dff_A_g9U8ADko8_0(.dout(w_dff_A_xFuGE22u5_0),.din(w_dff_A_g9U8ADko8_0),.clk(gclk));
	jdff dff_A_xFuGE22u5_0(.dout(w_dff_A_P4hpayBY0_0),.din(w_dff_A_xFuGE22u5_0),.clk(gclk));
	jdff dff_A_P4hpayBY0_0(.dout(w_dff_A_hCCATq3l4_0),.din(w_dff_A_P4hpayBY0_0),.clk(gclk));
	jdff dff_A_hCCATq3l4_0(.dout(w_dff_A_fIboX2j20_0),.din(w_dff_A_hCCATq3l4_0),.clk(gclk));
	jdff dff_A_fIboX2j20_0(.dout(w_dff_A_DHO0Yl9L6_0),.din(w_dff_A_fIboX2j20_0),.clk(gclk));
	jdff dff_A_DHO0Yl9L6_0(.dout(w_dff_A_W4LvPFHI2_0),.din(w_dff_A_DHO0Yl9L6_0),.clk(gclk));
	jdff dff_A_W4LvPFHI2_0(.dout(G850),.din(w_dff_A_W4LvPFHI2_0),.clk(gclk));
	jdff dff_A_9O4gAV2i7_1(.dout(w_dff_A_VlzhPncD2_0),.din(w_dff_A_9O4gAV2i7_1),.clk(gclk));
	jdff dff_A_VlzhPncD2_0(.dout(w_dff_A_mAC2MZIc1_0),.din(w_dff_A_VlzhPncD2_0),.clk(gclk));
	jdff dff_A_mAC2MZIc1_0(.dout(w_dff_A_xNV2BHgZ1_0),.din(w_dff_A_mAC2MZIc1_0),.clk(gclk));
	jdff dff_A_xNV2BHgZ1_0(.dout(w_dff_A_2yPk94W95_0),.din(w_dff_A_xNV2BHgZ1_0),.clk(gclk));
	jdff dff_A_2yPk94W95_0(.dout(w_dff_A_wrbFE21X9_0),.din(w_dff_A_2yPk94W95_0),.clk(gclk));
	jdff dff_A_wrbFE21X9_0(.dout(w_dff_A_JEXyzaBW5_0),.din(w_dff_A_wrbFE21X9_0),.clk(gclk));
	jdff dff_A_JEXyzaBW5_0(.dout(w_dff_A_WMqTFTfS4_0),.din(w_dff_A_JEXyzaBW5_0),.clk(gclk));
	jdff dff_A_WMqTFTfS4_0(.dout(w_dff_A_L2x21T8C4_0),.din(w_dff_A_WMqTFTfS4_0),.clk(gclk));
	jdff dff_A_L2x21T8C4_0(.dout(w_dff_A_eqxLe8Ly2_0),.din(w_dff_A_L2x21T8C4_0),.clk(gclk));
	jdff dff_A_eqxLe8Ly2_0(.dout(w_dff_A_poOSoO2I6_0),.din(w_dff_A_eqxLe8Ly2_0),.clk(gclk));
	jdff dff_A_poOSoO2I6_0(.dout(w_dff_A_dPQMv4Ly5_0),.din(w_dff_A_poOSoO2I6_0),.clk(gclk));
	jdff dff_A_dPQMv4Ly5_0(.dout(w_dff_A_UTtF3snW4_0),.din(w_dff_A_dPQMv4Ly5_0),.clk(gclk));
	jdff dff_A_UTtF3snW4_0(.dout(w_dff_A_4CIW0D9p0_0),.din(w_dff_A_UTtF3snW4_0),.clk(gclk));
	jdff dff_A_4CIW0D9p0_0(.dout(w_dff_A_2oWqbx8g0_0),.din(w_dff_A_4CIW0D9p0_0),.clk(gclk));
	jdff dff_A_2oWqbx8g0_0(.dout(w_dff_A_eGUVLsiR1_0),.din(w_dff_A_2oWqbx8g0_0),.clk(gclk));
	jdff dff_A_eGUVLsiR1_0(.dout(w_dff_A_gFoE7tEK5_0),.din(w_dff_A_eGUVLsiR1_0),.clk(gclk));
	jdff dff_A_gFoE7tEK5_0(.dout(w_dff_A_qeXe7CHZ3_0),.din(w_dff_A_gFoE7tEK5_0),.clk(gclk));
	jdff dff_A_qeXe7CHZ3_0(.dout(w_dff_A_ll7FEGeB0_0),.din(w_dff_A_qeXe7CHZ3_0),.clk(gclk));
	jdff dff_A_ll7FEGeB0_0(.dout(w_dff_A_yqtzfzdn2_0),.din(w_dff_A_ll7FEGeB0_0),.clk(gclk));
	jdff dff_A_yqtzfzdn2_0(.dout(w_dff_A_cGLikj2N9_0),.din(w_dff_A_yqtzfzdn2_0),.clk(gclk));
	jdff dff_A_cGLikj2N9_0(.dout(w_dff_A_IF9OC0EY6_0),.din(w_dff_A_cGLikj2N9_0),.clk(gclk));
	jdff dff_A_IF9OC0EY6_0(.dout(w_dff_A_EVMxK5z23_0),.din(w_dff_A_IF9OC0EY6_0),.clk(gclk));
	jdff dff_A_EVMxK5z23_0(.dout(w_dff_A_CJUHXIz74_0),.din(w_dff_A_EVMxK5z23_0),.clk(gclk));
	jdff dff_A_CJUHXIz74_0(.dout(w_dff_A_LPG7EiUM4_0),.din(w_dff_A_CJUHXIz74_0),.clk(gclk));
	jdff dff_A_LPG7EiUM4_0(.dout(w_dff_A_wd7LoYRr0_0),.din(w_dff_A_LPG7EiUM4_0),.clk(gclk));
	jdff dff_A_wd7LoYRr0_0(.dout(w_dff_A_ed7jCAqA2_0),.din(w_dff_A_wd7LoYRr0_0),.clk(gclk));
	jdff dff_A_ed7jCAqA2_0(.dout(G851),.din(w_dff_A_ed7jCAqA2_0),.clk(gclk));
	jdff dff_A_wElPQzTe5_2(.dout(w_dff_A_4AOl2UH79_0),.din(w_dff_A_wElPQzTe5_2),.clk(gclk));
	jdff dff_A_4AOl2UH79_0(.dout(w_dff_A_JlKtbfur3_0),.din(w_dff_A_4AOl2UH79_0),.clk(gclk));
	jdff dff_A_JlKtbfur3_0(.dout(w_dff_A_DkNyWvK76_0),.din(w_dff_A_JlKtbfur3_0),.clk(gclk));
	jdff dff_A_DkNyWvK76_0(.dout(w_dff_A_mJmbW3Cc4_0),.din(w_dff_A_DkNyWvK76_0),.clk(gclk));
	jdff dff_A_mJmbW3Cc4_0(.dout(w_dff_A_UzGttZvD9_0),.din(w_dff_A_mJmbW3Cc4_0),.clk(gclk));
	jdff dff_A_UzGttZvD9_0(.dout(w_dff_A_YNd6SKU43_0),.din(w_dff_A_UzGttZvD9_0),.clk(gclk));
	jdff dff_A_YNd6SKU43_0(.dout(w_dff_A_Ov1Tvs7f5_0),.din(w_dff_A_YNd6SKU43_0),.clk(gclk));
	jdff dff_A_Ov1Tvs7f5_0(.dout(w_dff_A_dA0TC0dG4_0),.din(w_dff_A_Ov1Tvs7f5_0),.clk(gclk));
	jdff dff_A_dA0TC0dG4_0(.dout(w_dff_A_ZBWY9wqZ4_0),.din(w_dff_A_dA0TC0dG4_0),.clk(gclk));
	jdff dff_A_ZBWY9wqZ4_0(.dout(w_dff_A_AR1uQiiT7_0),.din(w_dff_A_ZBWY9wqZ4_0),.clk(gclk));
	jdff dff_A_AR1uQiiT7_0(.dout(w_dff_A_FRkgn1Go4_0),.din(w_dff_A_AR1uQiiT7_0),.clk(gclk));
	jdff dff_A_FRkgn1Go4_0(.dout(w_dff_A_QPLO1r0R1_0),.din(w_dff_A_FRkgn1Go4_0),.clk(gclk));
	jdff dff_A_QPLO1r0R1_0(.dout(w_dff_A_UBbajyiL4_0),.din(w_dff_A_QPLO1r0R1_0),.clk(gclk));
	jdff dff_A_UBbajyiL4_0(.dout(w_dff_A_nmLoOm7U5_0),.din(w_dff_A_UBbajyiL4_0),.clk(gclk));
	jdff dff_A_nmLoOm7U5_0(.dout(w_dff_A_cOdwUzQW6_0),.din(w_dff_A_nmLoOm7U5_0),.clk(gclk));
	jdff dff_A_cOdwUzQW6_0(.dout(w_dff_A_QGb8wMTu9_0),.din(w_dff_A_cOdwUzQW6_0),.clk(gclk));
	jdff dff_A_QGb8wMTu9_0(.dout(w_dff_A_LXWUVEv72_0),.din(w_dff_A_QGb8wMTu9_0),.clk(gclk));
	jdff dff_A_LXWUVEv72_0(.dout(w_dff_A_qwnZtuUh2_0),.din(w_dff_A_LXWUVEv72_0),.clk(gclk));
	jdff dff_A_qwnZtuUh2_0(.dout(w_dff_A_EhaPn7jp7_0),.din(w_dff_A_qwnZtuUh2_0),.clk(gclk));
	jdff dff_A_EhaPn7jp7_0(.dout(w_dff_A_MuPXOk6G3_0),.din(w_dff_A_EhaPn7jp7_0),.clk(gclk));
	jdff dff_A_MuPXOk6G3_0(.dout(w_dff_A_eJuhSk0E3_0),.din(w_dff_A_MuPXOk6G3_0),.clk(gclk));
	jdff dff_A_eJuhSk0E3_0(.dout(w_dff_A_uZ8yTvPd7_0),.din(w_dff_A_eJuhSk0E3_0),.clk(gclk));
	jdff dff_A_uZ8yTvPd7_0(.dout(w_dff_A_eEvjbcGu3_0),.din(w_dff_A_uZ8yTvPd7_0),.clk(gclk));
	jdff dff_A_eEvjbcGu3_0(.dout(w_dff_A_hUtW2DhM9_0),.din(w_dff_A_eEvjbcGu3_0),.clk(gclk));
	jdff dff_A_hUtW2DhM9_0(.dout(w_dff_A_obxRtBkU9_0),.din(w_dff_A_hUtW2DhM9_0),.clk(gclk));
	jdff dff_A_obxRtBkU9_0(.dout(w_dff_A_0UmWNMxX9_0),.din(w_dff_A_obxRtBkU9_0),.clk(gclk));
	jdff dff_A_0UmWNMxX9_0(.dout(G634),.din(w_dff_A_0UmWNMxX9_0),.clk(gclk));
	jdff dff_A_5ftdZgkS7_2(.dout(w_dff_A_CMaaRmQY4_0),.din(w_dff_A_5ftdZgkS7_2),.clk(gclk));
	jdff dff_A_CMaaRmQY4_0(.dout(w_dff_A_TeZA8vRj1_0),.din(w_dff_A_CMaaRmQY4_0),.clk(gclk));
	jdff dff_A_TeZA8vRj1_0(.dout(w_dff_A_bYTk6TVq9_0),.din(w_dff_A_TeZA8vRj1_0),.clk(gclk));
	jdff dff_A_bYTk6TVq9_0(.dout(w_dff_A_JtqXfOQ52_0),.din(w_dff_A_bYTk6TVq9_0),.clk(gclk));
	jdff dff_A_JtqXfOQ52_0(.dout(w_dff_A_Gl0DGDjm2_0),.din(w_dff_A_JtqXfOQ52_0),.clk(gclk));
	jdff dff_A_Gl0DGDjm2_0(.dout(w_dff_A_XBCRh5Pa5_0),.din(w_dff_A_Gl0DGDjm2_0),.clk(gclk));
	jdff dff_A_XBCRh5Pa5_0(.dout(w_dff_A_hXemu6u64_0),.din(w_dff_A_XBCRh5Pa5_0),.clk(gclk));
	jdff dff_A_hXemu6u64_0(.dout(w_dff_A_7qpG2OMS7_0),.din(w_dff_A_hXemu6u64_0),.clk(gclk));
	jdff dff_A_7qpG2OMS7_0(.dout(w_dff_A_j2lCvmCJ4_0),.din(w_dff_A_7qpG2OMS7_0),.clk(gclk));
	jdff dff_A_j2lCvmCJ4_0(.dout(w_dff_A_lTi6JReR2_0),.din(w_dff_A_j2lCvmCJ4_0),.clk(gclk));
	jdff dff_A_lTi6JReR2_0(.dout(w_dff_A_9NPOSaKl7_0),.din(w_dff_A_lTi6JReR2_0),.clk(gclk));
	jdff dff_A_9NPOSaKl7_0(.dout(w_dff_A_BrrOSoGj3_0),.din(w_dff_A_9NPOSaKl7_0),.clk(gclk));
	jdff dff_A_BrrOSoGj3_0(.dout(w_dff_A_VfwoEhfr4_0),.din(w_dff_A_BrrOSoGj3_0),.clk(gclk));
	jdff dff_A_VfwoEhfr4_0(.dout(w_dff_A_sgMNeLux8_0),.din(w_dff_A_VfwoEhfr4_0),.clk(gclk));
	jdff dff_A_sgMNeLux8_0(.dout(w_dff_A_tuU4C99N4_0),.din(w_dff_A_sgMNeLux8_0),.clk(gclk));
	jdff dff_A_tuU4C99N4_0(.dout(w_dff_A_rzzQlwH61_0),.din(w_dff_A_tuU4C99N4_0),.clk(gclk));
	jdff dff_A_rzzQlwH61_0(.dout(w_dff_A_iGuArtNh5_0),.din(w_dff_A_rzzQlwH61_0),.clk(gclk));
	jdff dff_A_iGuArtNh5_0(.dout(w_dff_A_3Qf12oSp8_0),.din(w_dff_A_iGuArtNh5_0),.clk(gclk));
	jdff dff_A_3Qf12oSp8_0(.dout(w_dff_A_8w1NMvb74_0),.din(w_dff_A_3Qf12oSp8_0),.clk(gclk));
	jdff dff_A_8w1NMvb74_0(.dout(w_dff_A_aDNivSHy6_0),.din(w_dff_A_8w1NMvb74_0),.clk(gclk));
	jdff dff_A_aDNivSHy6_0(.dout(w_dff_A_yj4CGCgA1_0),.din(w_dff_A_aDNivSHy6_0),.clk(gclk));
	jdff dff_A_yj4CGCgA1_0(.dout(w_dff_A_WrKFg0mw8_0),.din(w_dff_A_yj4CGCgA1_0),.clk(gclk));
	jdff dff_A_WrKFg0mw8_0(.dout(w_dff_A_c0JWgtOE4_0),.din(w_dff_A_WrKFg0mw8_0),.clk(gclk));
	jdff dff_A_c0JWgtOE4_0(.dout(w_dff_A_BzV8wqwf9_0),.din(w_dff_A_c0JWgtOE4_0),.clk(gclk));
	jdff dff_A_BzV8wqwf9_0(.dout(w_dff_A_4CP3EiGh6_0),.din(w_dff_A_BzV8wqwf9_0),.clk(gclk));
	jdff dff_A_4CP3EiGh6_0(.dout(G815),.din(w_dff_A_4CP3EiGh6_0),.clk(gclk));
	jdff dff_A_nNW8Oyib6_2(.dout(w_dff_A_n2FdJ63z5_0),.din(w_dff_A_nNW8Oyib6_2),.clk(gclk));
	jdff dff_A_n2FdJ63z5_0(.dout(w_dff_A_3hoEDqA48_0),.din(w_dff_A_n2FdJ63z5_0),.clk(gclk));
	jdff dff_A_3hoEDqA48_0(.dout(w_dff_A_sysUsWEc8_0),.din(w_dff_A_3hoEDqA48_0),.clk(gclk));
	jdff dff_A_sysUsWEc8_0(.dout(w_dff_A_CYim9ad56_0),.din(w_dff_A_sysUsWEc8_0),.clk(gclk));
	jdff dff_A_CYim9ad56_0(.dout(w_dff_A_bbMcMkbS4_0),.din(w_dff_A_CYim9ad56_0),.clk(gclk));
	jdff dff_A_bbMcMkbS4_0(.dout(w_dff_A_usgfN2SQ1_0),.din(w_dff_A_bbMcMkbS4_0),.clk(gclk));
	jdff dff_A_usgfN2SQ1_0(.dout(w_dff_A_ZHwqDeh71_0),.din(w_dff_A_usgfN2SQ1_0),.clk(gclk));
	jdff dff_A_ZHwqDeh71_0(.dout(w_dff_A_23SLu1YI9_0),.din(w_dff_A_ZHwqDeh71_0),.clk(gclk));
	jdff dff_A_23SLu1YI9_0(.dout(w_dff_A_i3VyskVW1_0),.din(w_dff_A_23SLu1YI9_0),.clk(gclk));
	jdff dff_A_i3VyskVW1_0(.dout(w_dff_A_dtyqkMfr6_0),.din(w_dff_A_i3VyskVW1_0),.clk(gclk));
	jdff dff_A_dtyqkMfr6_0(.dout(w_dff_A_U7dZrVpH5_0),.din(w_dff_A_dtyqkMfr6_0),.clk(gclk));
	jdff dff_A_U7dZrVpH5_0(.dout(w_dff_A_1KddJRVb4_0),.din(w_dff_A_U7dZrVpH5_0),.clk(gclk));
	jdff dff_A_1KddJRVb4_0(.dout(w_dff_A_9Y8SiPe14_0),.din(w_dff_A_1KddJRVb4_0),.clk(gclk));
	jdff dff_A_9Y8SiPe14_0(.dout(w_dff_A_cNKUpofq4_0),.din(w_dff_A_9Y8SiPe14_0),.clk(gclk));
	jdff dff_A_cNKUpofq4_0(.dout(w_dff_A_uFhzg1g85_0),.din(w_dff_A_cNKUpofq4_0),.clk(gclk));
	jdff dff_A_uFhzg1g85_0(.dout(w_dff_A_Im1meCHG2_0),.din(w_dff_A_uFhzg1g85_0),.clk(gclk));
	jdff dff_A_Im1meCHG2_0(.dout(w_dff_A_oTmKnql35_0),.din(w_dff_A_Im1meCHG2_0),.clk(gclk));
	jdff dff_A_oTmKnql35_0(.dout(w_dff_A_UtBCzH9v6_0),.din(w_dff_A_oTmKnql35_0),.clk(gclk));
	jdff dff_A_UtBCzH9v6_0(.dout(w_dff_A_eiCgoMAU3_0),.din(w_dff_A_UtBCzH9v6_0),.clk(gclk));
	jdff dff_A_eiCgoMAU3_0(.dout(w_dff_A_6lobc3xM7_0),.din(w_dff_A_eiCgoMAU3_0),.clk(gclk));
	jdff dff_A_6lobc3xM7_0(.dout(w_dff_A_z3VMAUdJ6_0),.din(w_dff_A_6lobc3xM7_0),.clk(gclk));
	jdff dff_A_z3VMAUdJ6_0(.dout(w_dff_A_1sDwaukh1_0),.din(w_dff_A_z3VMAUdJ6_0),.clk(gclk));
	jdff dff_A_1sDwaukh1_0(.dout(w_dff_A_jfUiw9GR5_0),.din(w_dff_A_1sDwaukh1_0),.clk(gclk));
	jdff dff_A_jfUiw9GR5_0(.dout(w_dff_A_ubHt4fJJ2_0),.din(w_dff_A_jfUiw9GR5_0),.clk(gclk));
	jdff dff_A_ubHt4fJJ2_0(.dout(w_dff_A_lshyIWXp2_0),.din(w_dff_A_ubHt4fJJ2_0),.clk(gclk));
	jdff dff_A_lshyIWXp2_0(.dout(G845),.din(w_dff_A_lshyIWXp2_0),.clk(gclk));
	jdff dff_A_IZSXO4y19_1(.dout(w_dff_A_FdvWJKLi8_0),.din(w_dff_A_IZSXO4y19_1),.clk(gclk));
	jdff dff_A_FdvWJKLi8_0(.dout(w_dff_A_DrzRPN2R6_0),.din(w_dff_A_FdvWJKLi8_0),.clk(gclk));
	jdff dff_A_DrzRPN2R6_0(.dout(w_dff_A_2lRx43hP9_0),.din(w_dff_A_DrzRPN2R6_0),.clk(gclk));
	jdff dff_A_2lRx43hP9_0(.dout(w_dff_A_32fzlnBH8_0),.din(w_dff_A_2lRx43hP9_0),.clk(gclk));
	jdff dff_A_32fzlnBH8_0(.dout(w_dff_A_7DbEmEQ39_0),.din(w_dff_A_32fzlnBH8_0),.clk(gclk));
	jdff dff_A_7DbEmEQ39_0(.dout(w_dff_A_n1W7Q6ga7_0),.din(w_dff_A_7DbEmEQ39_0),.clk(gclk));
	jdff dff_A_n1W7Q6ga7_0(.dout(w_dff_A_nP5pYstd3_0),.din(w_dff_A_n1W7Q6ga7_0),.clk(gclk));
	jdff dff_A_nP5pYstd3_0(.dout(w_dff_A_XSXuxrB71_0),.din(w_dff_A_nP5pYstd3_0),.clk(gclk));
	jdff dff_A_XSXuxrB71_0(.dout(w_dff_A_QCC3DIq40_0),.din(w_dff_A_XSXuxrB71_0),.clk(gclk));
	jdff dff_A_QCC3DIq40_0(.dout(w_dff_A_45UY7L592_0),.din(w_dff_A_QCC3DIq40_0),.clk(gclk));
	jdff dff_A_45UY7L592_0(.dout(w_dff_A_M4L6E43p3_0),.din(w_dff_A_45UY7L592_0),.clk(gclk));
	jdff dff_A_M4L6E43p3_0(.dout(w_dff_A_vmM6rYJd2_0),.din(w_dff_A_M4L6E43p3_0),.clk(gclk));
	jdff dff_A_vmM6rYJd2_0(.dout(w_dff_A_ACNoAteu2_0),.din(w_dff_A_vmM6rYJd2_0),.clk(gclk));
	jdff dff_A_ACNoAteu2_0(.dout(w_dff_A_wNhRjP6A5_0),.din(w_dff_A_ACNoAteu2_0),.clk(gclk));
	jdff dff_A_wNhRjP6A5_0(.dout(w_dff_A_S0oksRfg3_0),.din(w_dff_A_wNhRjP6A5_0),.clk(gclk));
	jdff dff_A_S0oksRfg3_0(.dout(w_dff_A_JZIrDp5I0_0),.din(w_dff_A_S0oksRfg3_0),.clk(gclk));
	jdff dff_A_JZIrDp5I0_0(.dout(w_dff_A_KicmJWUX2_0),.din(w_dff_A_JZIrDp5I0_0),.clk(gclk));
	jdff dff_A_KicmJWUX2_0(.dout(w_dff_A_PgAkvC1X2_0),.din(w_dff_A_KicmJWUX2_0),.clk(gclk));
	jdff dff_A_PgAkvC1X2_0(.dout(w_dff_A_8gATiKRr1_0),.din(w_dff_A_PgAkvC1X2_0),.clk(gclk));
	jdff dff_A_8gATiKRr1_0(.dout(w_dff_A_pgriklao0_0),.din(w_dff_A_8gATiKRr1_0),.clk(gclk));
	jdff dff_A_pgriklao0_0(.dout(w_dff_A_X5LgeMM37_0),.din(w_dff_A_pgriklao0_0),.clk(gclk));
	jdff dff_A_X5LgeMM37_0(.dout(w_dff_A_8HS1W8TA4_0),.din(w_dff_A_X5LgeMM37_0),.clk(gclk));
	jdff dff_A_8HS1W8TA4_0(.dout(w_dff_A_lEUlsqKZ1_0),.din(w_dff_A_8HS1W8TA4_0),.clk(gclk));
	jdff dff_A_lEUlsqKZ1_0(.dout(w_dff_A_KDgHikqk8_0),.din(w_dff_A_lEUlsqKZ1_0),.clk(gclk));
	jdff dff_A_KDgHikqk8_0(.dout(w_dff_A_BoNDu9p83_0),.din(w_dff_A_KDgHikqk8_0),.clk(gclk));
	jdff dff_A_BoNDu9p83_0(.dout(G847),.din(w_dff_A_BoNDu9p83_0),.clk(gclk));
	jdff dff_A_tBsHYMsf0_1(.dout(w_dff_A_Di9tBEy93_0),.din(w_dff_A_tBsHYMsf0_1),.clk(gclk));
	jdff dff_A_Di9tBEy93_0(.dout(w_dff_A_FRrNlEBd4_0),.din(w_dff_A_Di9tBEy93_0),.clk(gclk));
	jdff dff_A_FRrNlEBd4_0(.dout(w_dff_A_KDHxzONX2_0),.din(w_dff_A_FRrNlEBd4_0),.clk(gclk));
	jdff dff_A_KDHxzONX2_0(.dout(w_dff_A_tb6xgNvv2_0),.din(w_dff_A_KDHxzONX2_0),.clk(gclk));
	jdff dff_A_tb6xgNvv2_0(.dout(w_dff_A_16iSviNr2_0),.din(w_dff_A_tb6xgNvv2_0),.clk(gclk));
	jdff dff_A_16iSviNr2_0(.dout(w_dff_A_rlu5irWz5_0),.din(w_dff_A_16iSviNr2_0),.clk(gclk));
	jdff dff_A_rlu5irWz5_0(.dout(w_dff_A_2TB6mGr13_0),.din(w_dff_A_rlu5irWz5_0),.clk(gclk));
	jdff dff_A_2TB6mGr13_0(.dout(w_dff_A_yIYqBvIk8_0),.din(w_dff_A_2TB6mGr13_0),.clk(gclk));
	jdff dff_A_yIYqBvIk8_0(.dout(w_dff_A_nL8meCCM3_0),.din(w_dff_A_yIYqBvIk8_0),.clk(gclk));
	jdff dff_A_nL8meCCM3_0(.dout(w_dff_A_fqKWxqRr2_0),.din(w_dff_A_nL8meCCM3_0),.clk(gclk));
	jdff dff_A_fqKWxqRr2_0(.dout(w_dff_A_NUY8XYjB8_0),.din(w_dff_A_fqKWxqRr2_0),.clk(gclk));
	jdff dff_A_NUY8XYjB8_0(.dout(w_dff_A_gAw9JrmO5_0),.din(w_dff_A_NUY8XYjB8_0),.clk(gclk));
	jdff dff_A_gAw9JrmO5_0(.dout(w_dff_A_abkL6C4w1_0),.din(w_dff_A_gAw9JrmO5_0),.clk(gclk));
	jdff dff_A_abkL6C4w1_0(.dout(w_dff_A_7fPhmR1o3_0),.din(w_dff_A_abkL6C4w1_0),.clk(gclk));
	jdff dff_A_7fPhmR1o3_0(.dout(w_dff_A_ieokOxlL6_0),.din(w_dff_A_7fPhmR1o3_0),.clk(gclk));
	jdff dff_A_ieokOxlL6_0(.dout(w_dff_A_xmzZY5IA8_0),.din(w_dff_A_ieokOxlL6_0),.clk(gclk));
	jdff dff_A_xmzZY5IA8_0(.dout(w_dff_A_lL5ppykf2_0),.din(w_dff_A_xmzZY5IA8_0),.clk(gclk));
	jdff dff_A_lL5ppykf2_0(.dout(w_dff_A_1fZ3Z1300_0),.din(w_dff_A_lL5ppykf2_0),.clk(gclk));
	jdff dff_A_1fZ3Z1300_0(.dout(w_dff_A_A7DEkHDH2_0),.din(w_dff_A_1fZ3Z1300_0),.clk(gclk));
	jdff dff_A_A7DEkHDH2_0(.dout(w_dff_A_sdzZicac3_0),.din(w_dff_A_A7DEkHDH2_0),.clk(gclk));
	jdff dff_A_sdzZicac3_0(.dout(w_dff_A_vn2J0xgn3_0),.din(w_dff_A_sdzZicac3_0),.clk(gclk));
	jdff dff_A_vn2J0xgn3_0(.dout(w_dff_A_moB7jOxG0_0),.din(w_dff_A_vn2J0xgn3_0),.clk(gclk));
	jdff dff_A_moB7jOxG0_0(.dout(w_dff_A_MpMlg4gU8_0),.din(w_dff_A_moB7jOxG0_0),.clk(gclk));
	jdff dff_A_MpMlg4gU8_0(.dout(w_dff_A_E8J6kf2r8_0),.din(w_dff_A_MpMlg4gU8_0),.clk(gclk));
	jdff dff_A_E8J6kf2r8_0(.dout(w_dff_A_hyqtacLo7_0),.din(w_dff_A_E8J6kf2r8_0),.clk(gclk));
	jdff dff_A_hyqtacLo7_0(.dout(w_dff_A_fchFTvy15_0),.din(w_dff_A_hyqtacLo7_0),.clk(gclk));
	jdff dff_A_fchFTvy15_0(.dout(G926),.din(w_dff_A_fchFTvy15_0),.clk(gclk));
	jdff dff_A_tPCLe9f04_1(.dout(w_dff_A_APa8b5xU3_0),.din(w_dff_A_tPCLe9f04_1),.clk(gclk));
	jdff dff_A_APa8b5xU3_0(.dout(w_dff_A_0kTMdKbI4_0),.din(w_dff_A_APa8b5xU3_0),.clk(gclk));
	jdff dff_A_0kTMdKbI4_0(.dout(w_dff_A_AUCit7yg7_0),.din(w_dff_A_0kTMdKbI4_0),.clk(gclk));
	jdff dff_A_AUCit7yg7_0(.dout(w_dff_A_QZ0dxaob8_0),.din(w_dff_A_AUCit7yg7_0),.clk(gclk));
	jdff dff_A_QZ0dxaob8_0(.dout(w_dff_A_t9fDaZFZ9_0),.din(w_dff_A_QZ0dxaob8_0),.clk(gclk));
	jdff dff_A_t9fDaZFZ9_0(.dout(w_dff_A_XEpRULQ03_0),.din(w_dff_A_t9fDaZFZ9_0),.clk(gclk));
	jdff dff_A_XEpRULQ03_0(.dout(w_dff_A_66Gf8kif4_0),.din(w_dff_A_XEpRULQ03_0),.clk(gclk));
	jdff dff_A_66Gf8kif4_0(.dout(w_dff_A_rHx8OWQg6_0),.din(w_dff_A_66Gf8kif4_0),.clk(gclk));
	jdff dff_A_rHx8OWQg6_0(.dout(w_dff_A_mcoIyVux9_0),.din(w_dff_A_rHx8OWQg6_0),.clk(gclk));
	jdff dff_A_mcoIyVux9_0(.dout(w_dff_A_s69KssoD8_0),.din(w_dff_A_mcoIyVux9_0),.clk(gclk));
	jdff dff_A_s69KssoD8_0(.dout(w_dff_A_NFtq4UzW4_0),.din(w_dff_A_s69KssoD8_0),.clk(gclk));
	jdff dff_A_NFtq4UzW4_0(.dout(w_dff_A_UHkfVC438_0),.din(w_dff_A_NFtq4UzW4_0),.clk(gclk));
	jdff dff_A_UHkfVC438_0(.dout(w_dff_A_w0cdKska7_0),.din(w_dff_A_UHkfVC438_0),.clk(gclk));
	jdff dff_A_w0cdKska7_0(.dout(w_dff_A_odd9nTRY5_0),.din(w_dff_A_w0cdKska7_0),.clk(gclk));
	jdff dff_A_odd9nTRY5_0(.dout(w_dff_A_BQ1Z48kf7_0),.din(w_dff_A_odd9nTRY5_0),.clk(gclk));
	jdff dff_A_BQ1Z48kf7_0(.dout(w_dff_A_nvUjCZu32_0),.din(w_dff_A_BQ1Z48kf7_0),.clk(gclk));
	jdff dff_A_nvUjCZu32_0(.dout(w_dff_A_nLZSCQ2u2_0),.din(w_dff_A_nvUjCZu32_0),.clk(gclk));
	jdff dff_A_nLZSCQ2u2_0(.dout(w_dff_A_aqnbexse8_0),.din(w_dff_A_nLZSCQ2u2_0),.clk(gclk));
	jdff dff_A_aqnbexse8_0(.dout(w_dff_A_sk1Spi356_0),.din(w_dff_A_aqnbexse8_0),.clk(gclk));
	jdff dff_A_sk1Spi356_0(.dout(w_dff_A_pb3IABQT4_0),.din(w_dff_A_sk1Spi356_0),.clk(gclk));
	jdff dff_A_pb3IABQT4_0(.dout(w_dff_A_ouqLDWaW0_0),.din(w_dff_A_pb3IABQT4_0),.clk(gclk));
	jdff dff_A_ouqLDWaW0_0(.dout(w_dff_A_01kzzUme9_0),.din(w_dff_A_ouqLDWaW0_0),.clk(gclk));
	jdff dff_A_01kzzUme9_0(.dout(w_dff_A_KXvKvncn6_0),.din(w_dff_A_01kzzUme9_0),.clk(gclk));
	jdff dff_A_KXvKvncn6_0(.dout(w_dff_A_ClpyFt7J9_0),.din(w_dff_A_KXvKvncn6_0),.clk(gclk));
	jdff dff_A_ClpyFt7J9_0(.dout(w_dff_A_aZQfPyvd9_0),.din(w_dff_A_ClpyFt7J9_0),.clk(gclk));
	jdff dff_A_aZQfPyvd9_0(.dout(w_dff_A_dafibjqx9_0),.din(w_dff_A_aZQfPyvd9_0),.clk(gclk));
	jdff dff_A_dafibjqx9_0(.dout(G923),.din(w_dff_A_dafibjqx9_0),.clk(gclk));
	jdff dff_A_mnbyVjQA2_1(.dout(w_dff_A_Jm13IGCP0_0),.din(w_dff_A_mnbyVjQA2_1),.clk(gclk));
	jdff dff_A_Jm13IGCP0_0(.dout(w_dff_A_fhbz7wsS6_0),.din(w_dff_A_Jm13IGCP0_0),.clk(gclk));
	jdff dff_A_fhbz7wsS6_0(.dout(w_dff_A_UlAn2Kdo1_0),.din(w_dff_A_fhbz7wsS6_0),.clk(gclk));
	jdff dff_A_UlAn2Kdo1_0(.dout(w_dff_A_J3GvyTlB8_0),.din(w_dff_A_UlAn2Kdo1_0),.clk(gclk));
	jdff dff_A_J3GvyTlB8_0(.dout(w_dff_A_cBNDgBw72_0),.din(w_dff_A_J3GvyTlB8_0),.clk(gclk));
	jdff dff_A_cBNDgBw72_0(.dout(w_dff_A_5kuH9gVS2_0),.din(w_dff_A_cBNDgBw72_0),.clk(gclk));
	jdff dff_A_5kuH9gVS2_0(.dout(w_dff_A_b052TarJ5_0),.din(w_dff_A_5kuH9gVS2_0),.clk(gclk));
	jdff dff_A_b052TarJ5_0(.dout(w_dff_A_NzKOpNRB5_0),.din(w_dff_A_b052TarJ5_0),.clk(gclk));
	jdff dff_A_NzKOpNRB5_0(.dout(w_dff_A_L5yaxj4p3_0),.din(w_dff_A_NzKOpNRB5_0),.clk(gclk));
	jdff dff_A_L5yaxj4p3_0(.dout(w_dff_A_317FVENG8_0),.din(w_dff_A_L5yaxj4p3_0),.clk(gclk));
	jdff dff_A_317FVENG8_0(.dout(w_dff_A_LKKJsjVo7_0),.din(w_dff_A_317FVENG8_0),.clk(gclk));
	jdff dff_A_LKKJsjVo7_0(.dout(w_dff_A_bCx5BuDl4_0),.din(w_dff_A_LKKJsjVo7_0),.clk(gclk));
	jdff dff_A_bCx5BuDl4_0(.dout(w_dff_A_6DjmhvjB9_0),.din(w_dff_A_bCx5BuDl4_0),.clk(gclk));
	jdff dff_A_6DjmhvjB9_0(.dout(w_dff_A_DWYFI0Vn2_0),.din(w_dff_A_6DjmhvjB9_0),.clk(gclk));
	jdff dff_A_DWYFI0Vn2_0(.dout(w_dff_A_7e0zUIbQ6_0),.din(w_dff_A_DWYFI0Vn2_0),.clk(gclk));
	jdff dff_A_7e0zUIbQ6_0(.dout(w_dff_A_lOZo7eb14_0),.din(w_dff_A_7e0zUIbQ6_0),.clk(gclk));
	jdff dff_A_lOZo7eb14_0(.dout(w_dff_A_wP2WmMbE2_0),.din(w_dff_A_lOZo7eb14_0),.clk(gclk));
	jdff dff_A_wP2WmMbE2_0(.dout(w_dff_A_mwwNQD667_0),.din(w_dff_A_wP2WmMbE2_0),.clk(gclk));
	jdff dff_A_mwwNQD667_0(.dout(w_dff_A_f462eIbp7_0),.din(w_dff_A_mwwNQD667_0),.clk(gclk));
	jdff dff_A_f462eIbp7_0(.dout(w_dff_A_6gt7HUvI4_0),.din(w_dff_A_f462eIbp7_0),.clk(gclk));
	jdff dff_A_6gt7HUvI4_0(.dout(w_dff_A_wjDFJL4O0_0),.din(w_dff_A_6gt7HUvI4_0),.clk(gclk));
	jdff dff_A_wjDFJL4O0_0(.dout(w_dff_A_vieZz9Ka5_0),.din(w_dff_A_wjDFJL4O0_0),.clk(gclk));
	jdff dff_A_vieZz9Ka5_0(.dout(w_dff_A_1qpbX8co8_0),.din(w_dff_A_vieZz9Ka5_0),.clk(gclk));
	jdff dff_A_1qpbX8co8_0(.dout(w_dff_A_2bmp3zIS0_0),.din(w_dff_A_1qpbX8co8_0),.clk(gclk));
	jdff dff_A_2bmp3zIS0_0(.dout(w_dff_A_RcPgZUiL4_0),.din(w_dff_A_2bmp3zIS0_0),.clk(gclk));
	jdff dff_A_RcPgZUiL4_0(.dout(w_dff_A_knvHDWqy4_0),.din(w_dff_A_RcPgZUiL4_0),.clk(gclk));
	jdff dff_A_knvHDWqy4_0(.dout(G921),.din(w_dff_A_knvHDWqy4_0),.clk(gclk));
	jdff dff_A_HsXSJqmW2_1(.dout(w_dff_A_OKpwcyB81_0),.din(w_dff_A_HsXSJqmW2_1),.clk(gclk));
	jdff dff_A_OKpwcyB81_0(.dout(w_dff_A_3F3vAHQd6_0),.din(w_dff_A_OKpwcyB81_0),.clk(gclk));
	jdff dff_A_3F3vAHQd6_0(.dout(w_dff_A_rggA0Xjo4_0),.din(w_dff_A_3F3vAHQd6_0),.clk(gclk));
	jdff dff_A_rggA0Xjo4_0(.dout(w_dff_A_vtwirMfd2_0),.din(w_dff_A_rggA0Xjo4_0),.clk(gclk));
	jdff dff_A_vtwirMfd2_0(.dout(w_dff_A_uSiiAwV32_0),.din(w_dff_A_vtwirMfd2_0),.clk(gclk));
	jdff dff_A_uSiiAwV32_0(.dout(w_dff_A_MMk7vI6F0_0),.din(w_dff_A_uSiiAwV32_0),.clk(gclk));
	jdff dff_A_MMk7vI6F0_0(.dout(w_dff_A_XJfbGET98_0),.din(w_dff_A_MMk7vI6F0_0),.clk(gclk));
	jdff dff_A_XJfbGET98_0(.dout(w_dff_A_enUVeP9G1_0),.din(w_dff_A_XJfbGET98_0),.clk(gclk));
	jdff dff_A_enUVeP9G1_0(.dout(w_dff_A_RW2z4dJ44_0),.din(w_dff_A_enUVeP9G1_0),.clk(gclk));
	jdff dff_A_RW2z4dJ44_0(.dout(w_dff_A_9Cm7KGQt9_0),.din(w_dff_A_RW2z4dJ44_0),.clk(gclk));
	jdff dff_A_9Cm7KGQt9_0(.dout(w_dff_A_BoATiG8v7_0),.din(w_dff_A_9Cm7KGQt9_0),.clk(gclk));
	jdff dff_A_BoATiG8v7_0(.dout(w_dff_A_65ZGevFm9_0),.din(w_dff_A_BoATiG8v7_0),.clk(gclk));
	jdff dff_A_65ZGevFm9_0(.dout(w_dff_A_URTE9TmN8_0),.din(w_dff_A_65ZGevFm9_0),.clk(gclk));
	jdff dff_A_URTE9TmN8_0(.dout(w_dff_A_HfyHt0xL1_0),.din(w_dff_A_URTE9TmN8_0),.clk(gclk));
	jdff dff_A_HfyHt0xL1_0(.dout(w_dff_A_TUWilLHJ6_0),.din(w_dff_A_HfyHt0xL1_0),.clk(gclk));
	jdff dff_A_TUWilLHJ6_0(.dout(w_dff_A_myPRZoEq7_0),.din(w_dff_A_TUWilLHJ6_0),.clk(gclk));
	jdff dff_A_myPRZoEq7_0(.dout(w_dff_A_N51r9fdv0_0),.din(w_dff_A_myPRZoEq7_0),.clk(gclk));
	jdff dff_A_N51r9fdv0_0(.dout(w_dff_A_zunUBKVQ0_0),.din(w_dff_A_N51r9fdv0_0),.clk(gclk));
	jdff dff_A_zunUBKVQ0_0(.dout(w_dff_A_NX7Px3B18_0),.din(w_dff_A_zunUBKVQ0_0),.clk(gclk));
	jdff dff_A_NX7Px3B18_0(.dout(w_dff_A_0eb4s6Ac5_0),.din(w_dff_A_NX7Px3B18_0),.clk(gclk));
	jdff dff_A_0eb4s6Ac5_0(.dout(w_dff_A_wKPSXQ9S5_0),.din(w_dff_A_0eb4s6Ac5_0),.clk(gclk));
	jdff dff_A_wKPSXQ9S5_0(.dout(w_dff_A_WS8MKiuX9_0),.din(w_dff_A_wKPSXQ9S5_0),.clk(gclk));
	jdff dff_A_WS8MKiuX9_0(.dout(w_dff_A_HW2uTXjD8_0),.din(w_dff_A_WS8MKiuX9_0),.clk(gclk));
	jdff dff_A_HW2uTXjD8_0(.dout(w_dff_A_01lhwsU58_0),.din(w_dff_A_HW2uTXjD8_0),.clk(gclk));
	jdff dff_A_01lhwsU58_0(.dout(w_dff_A_UyJWuDAO7_0),.din(w_dff_A_01lhwsU58_0),.clk(gclk));
	jdff dff_A_UyJWuDAO7_0(.dout(w_dff_A_mfr6wMuy6_0),.din(w_dff_A_UyJWuDAO7_0),.clk(gclk));
	jdff dff_A_mfr6wMuy6_0(.dout(G892),.din(w_dff_A_mfr6wMuy6_0),.clk(gclk));
	jdff dff_A_YrcMuZjh5_1(.dout(w_dff_A_jhEr5zGS5_0),.din(w_dff_A_YrcMuZjh5_1),.clk(gclk));
	jdff dff_A_jhEr5zGS5_0(.dout(w_dff_A_vjbUvAEs7_0),.din(w_dff_A_jhEr5zGS5_0),.clk(gclk));
	jdff dff_A_vjbUvAEs7_0(.dout(w_dff_A_yLelHxPb9_0),.din(w_dff_A_vjbUvAEs7_0),.clk(gclk));
	jdff dff_A_yLelHxPb9_0(.dout(w_dff_A_ZDCQfVVY7_0),.din(w_dff_A_yLelHxPb9_0),.clk(gclk));
	jdff dff_A_ZDCQfVVY7_0(.dout(w_dff_A_CXROt8NI0_0),.din(w_dff_A_ZDCQfVVY7_0),.clk(gclk));
	jdff dff_A_CXROt8NI0_0(.dout(w_dff_A_u0KRek7n0_0),.din(w_dff_A_CXROt8NI0_0),.clk(gclk));
	jdff dff_A_u0KRek7n0_0(.dout(w_dff_A_sB0yXDSc6_0),.din(w_dff_A_u0KRek7n0_0),.clk(gclk));
	jdff dff_A_sB0yXDSc6_0(.dout(w_dff_A_fiLpjyuf1_0),.din(w_dff_A_sB0yXDSc6_0),.clk(gclk));
	jdff dff_A_fiLpjyuf1_0(.dout(w_dff_A_rUUSTHGH2_0),.din(w_dff_A_fiLpjyuf1_0),.clk(gclk));
	jdff dff_A_rUUSTHGH2_0(.dout(w_dff_A_WLXMhlYe7_0),.din(w_dff_A_rUUSTHGH2_0),.clk(gclk));
	jdff dff_A_WLXMhlYe7_0(.dout(w_dff_A_mN1szGLP0_0),.din(w_dff_A_WLXMhlYe7_0),.clk(gclk));
	jdff dff_A_mN1szGLP0_0(.dout(w_dff_A_kulQlXRO5_0),.din(w_dff_A_mN1szGLP0_0),.clk(gclk));
	jdff dff_A_kulQlXRO5_0(.dout(w_dff_A_iiseMS9g5_0),.din(w_dff_A_kulQlXRO5_0),.clk(gclk));
	jdff dff_A_iiseMS9g5_0(.dout(w_dff_A_q4JDALdd1_0),.din(w_dff_A_iiseMS9g5_0),.clk(gclk));
	jdff dff_A_q4JDALdd1_0(.dout(w_dff_A_Ld6FerP87_0),.din(w_dff_A_q4JDALdd1_0),.clk(gclk));
	jdff dff_A_Ld6FerP87_0(.dout(w_dff_A_rlfMbOL13_0),.din(w_dff_A_Ld6FerP87_0),.clk(gclk));
	jdff dff_A_rlfMbOL13_0(.dout(w_dff_A_3pIkzwlY5_0),.din(w_dff_A_rlfMbOL13_0),.clk(gclk));
	jdff dff_A_3pIkzwlY5_0(.dout(w_dff_A_CSqsZH544_0),.din(w_dff_A_3pIkzwlY5_0),.clk(gclk));
	jdff dff_A_CSqsZH544_0(.dout(w_dff_A_XX0lVAs04_0),.din(w_dff_A_CSqsZH544_0),.clk(gclk));
	jdff dff_A_XX0lVAs04_0(.dout(w_dff_A_5ljnhUSX1_0),.din(w_dff_A_XX0lVAs04_0),.clk(gclk));
	jdff dff_A_5ljnhUSX1_0(.dout(w_dff_A_9wXbLuQx4_0),.din(w_dff_A_5ljnhUSX1_0),.clk(gclk));
	jdff dff_A_9wXbLuQx4_0(.dout(w_dff_A_Mj3Yn2ok4_0),.din(w_dff_A_9wXbLuQx4_0),.clk(gclk));
	jdff dff_A_Mj3Yn2ok4_0(.dout(w_dff_A_gKOno9Oj4_0),.din(w_dff_A_Mj3Yn2ok4_0),.clk(gclk));
	jdff dff_A_gKOno9Oj4_0(.dout(w_dff_A_UIzerzom4_0),.din(w_dff_A_gKOno9Oj4_0),.clk(gclk));
	jdff dff_A_UIzerzom4_0(.dout(w_dff_A_mSOx0lHj4_0),.din(w_dff_A_UIzerzom4_0),.clk(gclk));
	jdff dff_A_mSOx0lHj4_0(.dout(w_dff_A_8xdMCJWG0_0),.din(w_dff_A_mSOx0lHj4_0),.clk(gclk));
	jdff dff_A_8xdMCJWG0_0(.dout(G887),.din(w_dff_A_8xdMCJWG0_0),.clk(gclk));
	jdff dff_A_i0f25SsS5_1(.dout(w_dff_A_EaoC9uBY9_0),.din(w_dff_A_i0f25SsS5_1),.clk(gclk));
	jdff dff_A_EaoC9uBY9_0(.dout(w_dff_A_SSYifb0q5_0),.din(w_dff_A_EaoC9uBY9_0),.clk(gclk));
	jdff dff_A_SSYifb0q5_0(.dout(w_dff_A_fxEzwhkz5_0),.din(w_dff_A_SSYifb0q5_0),.clk(gclk));
	jdff dff_A_fxEzwhkz5_0(.dout(w_dff_A_gImH4YvO7_0),.din(w_dff_A_fxEzwhkz5_0),.clk(gclk));
	jdff dff_A_gImH4YvO7_0(.dout(w_dff_A_mx8rY8fB6_0),.din(w_dff_A_gImH4YvO7_0),.clk(gclk));
	jdff dff_A_mx8rY8fB6_0(.dout(w_dff_A_BjcwPdQA4_0),.din(w_dff_A_mx8rY8fB6_0),.clk(gclk));
	jdff dff_A_BjcwPdQA4_0(.dout(w_dff_A_pPx2SNbI8_0),.din(w_dff_A_BjcwPdQA4_0),.clk(gclk));
	jdff dff_A_pPx2SNbI8_0(.dout(w_dff_A_uyXOxEBR7_0),.din(w_dff_A_pPx2SNbI8_0),.clk(gclk));
	jdff dff_A_uyXOxEBR7_0(.dout(w_dff_A_8rO5yTEq1_0),.din(w_dff_A_uyXOxEBR7_0),.clk(gclk));
	jdff dff_A_8rO5yTEq1_0(.dout(w_dff_A_w57orzIn7_0),.din(w_dff_A_8rO5yTEq1_0),.clk(gclk));
	jdff dff_A_w57orzIn7_0(.dout(w_dff_A_ob5EmfXZ0_0),.din(w_dff_A_w57orzIn7_0),.clk(gclk));
	jdff dff_A_ob5EmfXZ0_0(.dout(w_dff_A_vJT2ArS15_0),.din(w_dff_A_ob5EmfXZ0_0),.clk(gclk));
	jdff dff_A_vJT2ArS15_0(.dout(w_dff_A_5iai8qls3_0),.din(w_dff_A_vJT2ArS15_0),.clk(gclk));
	jdff dff_A_5iai8qls3_0(.dout(w_dff_A_UxVvbBJv4_0),.din(w_dff_A_5iai8qls3_0),.clk(gclk));
	jdff dff_A_UxVvbBJv4_0(.dout(w_dff_A_XRKPOS2V9_0),.din(w_dff_A_UxVvbBJv4_0),.clk(gclk));
	jdff dff_A_XRKPOS2V9_0(.dout(w_dff_A_Vcg7Vzz66_0),.din(w_dff_A_XRKPOS2V9_0),.clk(gclk));
	jdff dff_A_Vcg7Vzz66_0(.dout(w_dff_A_z3FQ501J3_0),.din(w_dff_A_Vcg7Vzz66_0),.clk(gclk));
	jdff dff_A_z3FQ501J3_0(.dout(w_dff_A_wtDX4HwP1_0),.din(w_dff_A_z3FQ501J3_0),.clk(gclk));
	jdff dff_A_wtDX4HwP1_0(.dout(w_dff_A_iR93SuQP7_0),.din(w_dff_A_wtDX4HwP1_0),.clk(gclk));
	jdff dff_A_iR93SuQP7_0(.dout(w_dff_A_AqdjrelI3_0),.din(w_dff_A_iR93SuQP7_0),.clk(gclk));
	jdff dff_A_AqdjrelI3_0(.dout(w_dff_A_VHv4GM3C5_0),.din(w_dff_A_AqdjrelI3_0),.clk(gclk));
	jdff dff_A_VHv4GM3C5_0(.dout(w_dff_A_H8DPBpjF6_0),.din(w_dff_A_VHv4GM3C5_0),.clk(gclk));
	jdff dff_A_H8DPBpjF6_0(.dout(w_dff_A_VJ3md6VJ3_0),.din(w_dff_A_H8DPBpjF6_0),.clk(gclk));
	jdff dff_A_VJ3md6VJ3_0(.dout(w_dff_A_tzFXcQsT8_0),.din(w_dff_A_VJ3md6VJ3_0),.clk(gclk));
	jdff dff_A_tzFXcQsT8_0(.dout(w_dff_A_3mgvfYY55_0),.din(w_dff_A_tzFXcQsT8_0),.clk(gclk));
	jdff dff_A_3mgvfYY55_0(.dout(w_dff_A_Tt7Kreo86_0),.din(w_dff_A_3mgvfYY55_0),.clk(gclk));
	jdff dff_A_Tt7Kreo86_0(.dout(G606),.din(w_dff_A_Tt7Kreo86_0),.clk(gclk));
	jdff dff_A_pkH3YkUJ5_2(.dout(w_dff_A_bVproxhZ1_0),.din(w_dff_A_pkH3YkUJ5_2),.clk(gclk));
	jdff dff_A_bVproxhZ1_0(.dout(w_dff_A_NnggmJRV8_0),.din(w_dff_A_bVproxhZ1_0),.clk(gclk));
	jdff dff_A_NnggmJRV8_0(.dout(w_dff_A_Dtng7xtL1_0),.din(w_dff_A_NnggmJRV8_0),.clk(gclk));
	jdff dff_A_Dtng7xtL1_0(.dout(w_dff_A_VzWPLMQo1_0),.din(w_dff_A_Dtng7xtL1_0),.clk(gclk));
	jdff dff_A_VzWPLMQo1_0(.dout(w_dff_A_5peywzLZ3_0),.din(w_dff_A_VzWPLMQo1_0),.clk(gclk));
	jdff dff_A_5peywzLZ3_0(.dout(w_dff_A_FknypKjz8_0),.din(w_dff_A_5peywzLZ3_0),.clk(gclk));
	jdff dff_A_FknypKjz8_0(.dout(w_dff_A_zYJzvywN2_0),.din(w_dff_A_FknypKjz8_0),.clk(gclk));
	jdff dff_A_zYJzvywN2_0(.dout(w_dff_A_8d2IWV7w7_0),.din(w_dff_A_zYJzvywN2_0),.clk(gclk));
	jdff dff_A_8d2IWV7w7_0(.dout(w_dff_A_syANXWzw9_0),.din(w_dff_A_8d2IWV7w7_0),.clk(gclk));
	jdff dff_A_syANXWzw9_0(.dout(w_dff_A_mQRD1Het5_0),.din(w_dff_A_syANXWzw9_0),.clk(gclk));
	jdff dff_A_mQRD1Het5_0(.dout(w_dff_A_oz7vJrKv5_0),.din(w_dff_A_mQRD1Het5_0),.clk(gclk));
	jdff dff_A_oz7vJrKv5_0(.dout(w_dff_A_2gabycod7_0),.din(w_dff_A_oz7vJrKv5_0),.clk(gclk));
	jdff dff_A_2gabycod7_0(.dout(w_dff_A_RLZewH0M7_0),.din(w_dff_A_2gabycod7_0),.clk(gclk));
	jdff dff_A_RLZewH0M7_0(.dout(w_dff_A_SQ4fMz7y7_0),.din(w_dff_A_RLZewH0M7_0),.clk(gclk));
	jdff dff_A_SQ4fMz7y7_0(.dout(w_dff_A_P9lMhNpW4_0),.din(w_dff_A_SQ4fMz7y7_0),.clk(gclk));
	jdff dff_A_P9lMhNpW4_0(.dout(w_dff_A_SbWgZuYa5_0),.din(w_dff_A_P9lMhNpW4_0),.clk(gclk));
	jdff dff_A_SbWgZuYa5_0(.dout(w_dff_A_3p5gu8aV5_0),.din(w_dff_A_SbWgZuYa5_0),.clk(gclk));
	jdff dff_A_3p5gu8aV5_0(.dout(w_dff_A_XlJ7iejh3_0),.din(w_dff_A_3p5gu8aV5_0),.clk(gclk));
	jdff dff_A_XlJ7iejh3_0(.dout(w_dff_A_LyygyGZP6_0),.din(w_dff_A_XlJ7iejh3_0),.clk(gclk));
	jdff dff_A_LyygyGZP6_0(.dout(w_dff_A_n6ByNeGz2_0),.din(w_dff_A_LyygyGZP6_0),.clk(gclk));
	jdff dff_A_n6ByNeGz2_0(.dout(w_dff_A_4Uq4ytKh1_0),.din(w_dff_A_n6ByNeGz2_0),.clk(gclk));
	jdff dff_A_4Uq4ytKh1_0(.dout(w_dff_A_C9Nwdp014_0),.din(w_dff_A_4Uq4ytKh1_0),.clk(gclk));
	jdff dff_A_C9Nwdp014_0(.dout(w_dff_A_EpQxD4l68_0),.din(w_dff_A_C9Nwdp014_0),.clk(gclk));
	jdff dff_A_EpQxD4l68_0(.dout(w_dff_A_LcbV2KB71_0),.din(w_dff_A_EpQxD4l68_0),.clk(gclk));
	jdff dff_A_LcbV2KB71_0(.dout(G656),.din(w_dff_A_LcbV2KB71_0),.clk(gclk));
	jdff dff_A_f2GSdHvr4_2(.dout(w_dff_A_4GI2vdTM9_0),.din(w_dff_A_f2GSdHvr4_2),.clk(gclk));
	jdff dff_A_4GI2vdTM9_0(.dout(w_dff_A_9DPRFH3j1_0),.din(w_dff_A_4GI2vdTM9_0),.clk(gclk));
	jdff dff_A_9DPRFH3j1_0(.dout(w_dff_A_brnb3pLh2_0),.din(w_dff_A_9DPRFH3j1_0),.clk(gclk));
	jdff dff_A_brnb3pLh2_0(.dout(w_dff_A_4LTPbnYX6_0),.din(w_dff_A_brnb3pLh2_0),.clk(gclk));
	jdff dff_A_4LTPbnYX6_0(.dout(w_dff_A_432jsq1W8_0),.din(w_dff_A_4LTPbnYX6_0),.clk(gclk));
	jdff dff_A_432jsq1W8_0(.dout(w_dff_A_Nv5oegAo6_0),.din(w_dff_A_432jsq1W8_0),.clk(gclk));
	jdff dff_A_Nv5oegAo6_0(.dout(w_dff_A_l7UkE0E24_0),.din(w_dff_A_Nv5oegAo6_0),.clk(gclk));
	jdff dff_A_l7UkE0E24_0(.dout(w_dff_A_E7QuBlZJ4_0),.din(w_dff_A_l7UkE0E24_0),.clk(gclk));
	jdff dff_A_E7QuBlZJ4_0(.dout(w_dff_A_TwXQ17uT1_0),.din(w_dff_A_E7QuBlZJ4_0),.clk(gclk));
	jdff dff_A_TwXQ17uT1_0(.dout(w_dff_A_orOK3QiK0_0),.din(w_dff_A_TwXQ17uT1_0),.clk(gclk));
	jdff dff_A_orOK3QiK0_0(.dout(w_dff_A_OqWgzCzh6_0),.din(w_dff_A_orOK3QiK0_0),.clk(gclk));
	jdff dff_A_OqWgzCzh6_0(.dout(w_dff_A_ck27aEon9_0),.din(w_dff_A_OqWgzCzh6_0),.clk(gclk));
	jdff dff_A_ck27aEon9_0(.dout(w_dff_A_LlKry5MB5_0),.din(w_dff_A_ck27aEon9_0),.clk(gclk));
	jdff dff_A_LlKry5MB5_0(.dout(w_dff_A_GvQS4EHy0_0),.din(w_dff_A_LlKry5MB5_0),.clk(gclk));
	jdff dff_A_GvQS4EHy0_0(.dout(w_dff_A_k3ETe60u0_0),.din(w_dff_A_GvQS4EHy0_0),.clk(gclk));
	jdff dff_A_k3ETe60u0_0(.dout(w_dff_A_mY05oQWp8_0),.din(w_dff_A_k3ETe60u0_0),.clk(gclk));
	jdff dff_A_mY05oQWp8_0(.dout(w_dff_A_txr2TGNJ1_0),.din(w_dff_A_mY05oQWp8_0),.clk(gclk));
	jdff dff_A_txr2TGNJ1_0(.dout(w_dff_A_HhBUpIvU3_0),.din(w_dff_A_txr2TGNJ1_0),.clk(gclk));
	jdff dff_A_HhBUpIvU3_0(.dout(w_dff_A_RmNhbpNS3_0),.din(w_dff_A_HhBUpIvU3_0),.clk(gclk));
	jdff dff_A_RmNhbpNS3_0(.dout(w_dff_A_KJrxWuKz7_0),.din(w_dff_A_RmNhbpNS3_0),.clk(gclk));
	jdff dff_A_KJrxWuKz7_0(.dout(w_dff_A_ab98WgBp3_0),.din(w_dff_A_KJrxWuKz7_0),.clk(gclk));
	jdff dff_A_ab98WgBp3_0(.dout(w_dff_A_FEs7AWUG6_0),.din(w_dff_A_ab98WgBp3_0),.clk(gclk));
	jdff dff_A_FEs7AWUG6_0(.dout(w_dff_A_BmlfKb2Z0_0),.din(w_dff_A_FEs7AWUG6_0),.clk(gclk));
	jdff dff_A_BmlfKb2Z0_0(.dout(w_dff_A_5zh3mgN75_0),.din(w_dff_A_BmlfKb2Z0_0),.clk(gclk));
	jdff dff_A_5zh3mgN75_0(.dout(w_dff_A_t57oU9fo7_0),.din(w_dff_A_5zh3mgN75_0),.clk(gclk));
	jdff dff_A_t57oU9fo7_0(.dout(G809),.din(w_dff_A_t57oU9fo7_0),.clk(gclk));
	jdff dff_A_jBXFRELh6_1(.dout(w_dff_A_O4279mhi6_0),.din(w_dff_A_jBXFRELh6_1),.clk(gclk));
	jdff dff_A_O4279mhi6_0(.dout(w_dff_A_gkLomz2O2_0),.din(w_dff_A_O4279mhi6_0),.clk(gclk));
	jdff dff_A_gkLomz2O2_0(.dout(w_dff_A_5IO90M1b1_0),.din(w_dff_A_gkLomz2O2_0),.clk(gclk));
	jdff dff_A_5IO90M1b1_0(.dout(w_dff_A_w25WQnhG5_0),.din(w_dff_A_5IO90M1b1_0),.clk(gclk));
	jdff dff_A_w25WQnhG5_0(.dout(w_dff_A_Al5wD0XM5_0),.din(w_dff_A_w25WQnhG5_0),.clk(gclk));
	jdff dff_A_Al5wD0XM5_0(.dout(w_dff_A_WUt9Obbs2_0),.din(w_dff_A_Al5wD0XM5_0),.clk(gclk));
	jdff dff_A_WUt9Obbs2_0(.dout(w_dff_A_IEARGc4p8_0),.din(w_dff_A_WUt9Obbs2_0),.clk(gclk));
	jdff dff_A_IEARGc4p8_0(.dout(w_dff_A_oCdrQpEF4_0),.din(w_dff_A_IEARGc4p8_0),.clk(gclk));
	jdff dff_A_oCdrQpEF4_0(.dout(w_dff_A_0P59qezH7_0),.din(w_dff_A_oCdrQpEF4_0),.clk(gclk));
	jdff dff_A_0P59qezH7_0(.dout(w_dff_A_tf3dk7eV5_0),.din(w_dff_A_0P59qezH7_0),.clk(gclk));
	jdff dff_A_tf3dk7eV5_0(.dout(w_dff_A_eU0hxtQK5_0),.din(w_dff_A_tf3dk7eV5_0),.clk(gclk));
	jdff dff_A_eU0hxtQK5_0(.dout(w_dff_A_J8ltMfCs6_0),.din(w_dff_A_eU0hxtQK5_0),.clk(gclk));
	jdff dff_A_J8ltMfCs6_0(.dout(w_dff_A_qO1vkvcG9_0),.din(w_dff_A_J8ltMfCs6_0),.clk(gclk));
	jdff dff_A_qO1vkvcG9_0(.dout(w_dff_A_xSu0o2Jz4_0),.din(w_dff_A_qO1vkvcG9_0),.clk(gclk));
	jdff dff_A_xSu0o2Jz4_0(.dout(w_dff_A_m7EMncmL0_0),.din(w_dff_A_xSu0o2Jz4_0),.clk(gclk));
	jdff dff_A_m7EMncmL0_0(.dout(w_dff_A_rbuAS3CU6_0),.din(w_dff_A_m7EMncmL0_0),.clk(gclk));
	jdff dff_A_rbuAS3CU6_0(.dout(w_dff_A_7Z6O8Y0J9_0),.din(w_dff_A_rbuAS3CU6_0),.clk(gclk));
	jdff dff_A_7Z6O8Y0J9_0(.dout(w_dff_A_WX9bIBWT6_0),.din(w_dff_A_7Z6O8Y0J9_0),.clk(gclk));
	jdff dff_A_WX9bIBWT6_0(.dout(w_dff_A_cIln2rmy5_0),.din(w_dff_A_WX9bIBWT6_0),.clk(gclk));
	jdff dff_A_cIln2rmy5_0(.dout(w_dff_A_Rrj2gw9F6_0),.din(w_dff_A_cIln2rmy5_0),.clk(gclk));
	jdff dff_A_Rrj2gw9F6_0(.dout(w_dff_A_F36pxWCQ3_0),.din(w_dff_A_Rrj2gw9F6_0),.clk(gclk));
	jdff dff_A_F36pxWCQ3_0(.dout(w_dff_A_kEDOBLfu4_0),.din(w_dff_A_F36pxWCQ3_0),.clk(gclk));
	jdff dff_A_kEDOBLfu4_0(.dout(w_dff_A_loYdKfFg6_0),.din(w_dff_A_kEDOBLfu4_0),.clk(gclk));
	jdff dff_A_loYdKfFg6_0(.dout(w_dff_A_nO5ramgs1_0),.din(w_dff_A_loYdKfFg6_0),.clk(gclk));
	jdff dff_A_nO5ramgs1_0(.dout(w_dff_A_xxC0s3NU1_0),.din(w_dff_A_nO5ramgs1_0),.clk(gclk));
	jdff dff_A_xxC0s3NU1_0(.dout(w_dff_A_x4ak0bCm9_0),.din(w_dff_A_xxC0s3NU1_0),.clk(gclk));
	jdff dff_A_x4ak0bCm9_0(.dout(G993),.din(w_dff_A_x4ak0bCm9_0),.clk(gclk));
	jdff dff_A_AOkWbxaA9_1(.dout(w_dff_A_UrKL7IBP3_0),.din(w_dff_A_AOkWbxaA9_1),.clk(gclk));
	jdff dff_A_UrKL7IBP3_0(.dout(w_dff_A_OCoDPrgc0_0),.din(w_dff_A_UrKL7IBP3_0),.clk(gclk));
	jdff dff_A_OCoDPrgc0_0(.dout(w_dff_A_ID8Ltcb10_0),.din(w_dff_A_OCoDPrgc0_0),.clk(gclk));
	jdff dff_A_ID8Ltcb10_0(.dout(w_dff_A_Mz87F2Wy8_0),.din(w_dff_A_ID8Ltcb10_0),.clk(gclk));
	jdff dff_A_Mz87F2Wy8_0(.dout(w_dff_A_HspfVHHf7_0),.din(w_dff_A_Mz87F2Wy8_0),.clk(gclk));
	jdff dff_A_HspfVHHf7_0(.dout(w_dff_A_zX0zbdhB7_0),.din(w_dff_A_HspfVHHf7_0),.clk(gclk));
	jdff dff_A_zX0zbdhB7_0(.dout(w_dff_A_DlXVKrQM3_0),.din(w_dff_A_zX0zbdhB7_0),.clk(gclk));
	jdff dff_A_DlXVKrQM3_0(.dout(w_dff_A_og3hDeDi0_0),.din(w_dff_A_DlXVKrQM3_0),.clk(gclk));
	jdff dff_A_og3hDeDi0_0(.dout(w_dff_A_Y8uGbWbG4_0),.din(w_dff_A_og3hDeDi0_0),.clk(gclk));
	jdff dff_A_Y8uGbWbG4_0(.dout(w_dff_A_sTDa7OYi2_0),.din(w_dff_A_Y8uGbWbG4_0),.clk(gclk));
	jdff dff_A_sTDa7OYi2_0(.dout(w_dff_A_eWh4NSQ39_0),.din(w_dff_A_sTDa7OYi2_0),.clk(gclk));
	jdff dff_A_eWh4NSQ39_0(.dout(w_dff_A_BXFX4jj31_0),.din(w_dff_A_eWh4NSQ39_0),.clk(gclk));
	jdff dff_A_BXFX4jj31_0(.dout(w_dff_A_Jnkop36Y9_0),.din(w_dff_A_BXFX4jj31_0),.clk(gclk));
	jdff dff_A_Jnkop36Y9_0(.dout(w_dff_A_Vmxipy6w2_0),.din(w_dff_A_Jnkop36Y9_0),.clk(gclk));
	jdff dff_A_Vmxipy6w2_0(.dout(w_dff_A_Ok8Y0cGv1_0),.din(w_dff_A_Vmxipy6w2_0),.clk(gclk));
	jdff dff_A_Ok8Y0cGv1_0(.dout(w_dff_A_uwv5k4xR7_0),.din(w_dff_A_Ok8Y0cGv1_0),.clk(gclk));
	jdff dff_A_uwv5k4xR7_0(.dout(w_dff_A_qADDLnHx0_0),.din(w_dff_A_uwv5k4xR7_0),.clk(gclk));
	jdff dff_A_qADDLnHx0_0(.dout(w_dff_A_kgcBYuEQ4_0),.din(w_dff_A_qADDLnHx0_0),.clk(gclk));
	jdff dff_A_kgcBYuEQ4_0(.dout(w_dff_A_rAveruXr9_0),.din(w_dff_A_kgcBYuEQ4_0),.clk(gclk));
	jdff dff_A_rAveruXr9_0(.dout(w_dff_A_uQBIO8VC7_0),.din(w_dff_A_rAveruXr9_0),.clk(gclk));
	jdff dff_A_uQBIO8VC7_0(.dout(w_dff_A_WFc12DKO2_0),.din(w_dff_A_uQBIO8VC7_0),.clk(gclk));
	jdff dff_A_WFc12DKO2_0(.dout(w_dff_A_Tr9ThHPu3_0),.din(w_dff_A_WFc12DKO2_0),.clk(gclk));
	jdff dff_A_Tr9ThHPu3_0(.dout(w_dff_A_cMjBiDnC8_0),.din(w_dff_A_Tr9ThHPu3_0),.clk(gclk));
	jdff dff_A_cMjBiDnC8_0(.dout(w_dff_A_e5yMkLbO6_0),.din(w_dff_A_cMjBiDnC8_0),.clk(gclk));
	jdff dff_A_e5yMkLbO6_0(.dout(w_dff_A_NvcJmCpU8_0),.din(w_dff_A_e5yMkLbO6_0),.clk(gclk));
	jdff dff_A_NvcJmCpU8_0(.dout(w_dff_A_bBfrkhR76_0),.din(w_dff_A_NvcJmCpU8_0),.clk(gclk));
	jdff dff_A_bBfrkhR76_0(.dout(G978),.din(w_dff_A_bBfrkhR76_0),.clk(gclk));
	jdff dff_A_8UBzqmtz1_1(.dout(w_dff_A_xAMmuwKd7_0),.din(w_dff_A_8UBzqmtz1_1),.clk(gclk));
	jdff dff_A_xAMmuwKd7_0(.dout(w_dff_A_FCy7xAyr4_0),.din(w_dff_A_xAMmuwKd7_0),.clk(gclk));
	jdff dff_A_FCy7xAyr4_0(.dout(w_dff_A_hiaAwhs56_0),.din(w_dff_A_FCy7xAyr4_0),.clk(gclk));
	jdff dff_A_hiaAwhs56_0(.dout(w_dff_A_9aQqzs390_0),.din(w_dff_A_hiaAwhs56_0),.clk(gclk));
	jdff dff_A_9aQqzs390_0(.dout(w_dff_A_V4O7HvQ07_0),.din(w_dff_A_9aQqzs390_0),.clk(gclk));
	jdff dff_A_V4O7HvQ07_0(.dout(w_dff_A_6dOjmLPT6_0),.din(w_dff_A_V4O7HvQ07_0),.clk(gclk));
	jdff dff_A_6dOjmLPT6_0(.dout(w_dff_A_RArkxi7X6_0),.din(w_dff_A_6dOjmLPT6_0),.clk(gclk));
	jdff dff_A_RArkxi7X6_0(.dout(w_dff_A_lryukamR8_0),.din(w_dff_A_RArkxi7X6_0),.clk(gclk));
	jdff dff_A_lryukamR8_0(.dout(w_dff_A_a6ocVgTp5_0),.din(w_dff_A_lryukamR8_0),.clk(gclk));
	jdff dff_A_a6ocVgTp5_0(.dout(w_dff_A_HnBEWdAw3_0),.din(w_dff_A_a6ocVgTp5_0),.clk(gclk));
	jdff dff_A_HnBEWdAw3_0(.dout(w_dff_A_dJ5c2YAM4_0),.din(w_dff_A_HnBEWdAw3_0),.clk(gclk));
	jdff dff_A_dJ5c2YAM4_0(.dout(w_dff_A_RZhauPO90_0),.din(w_dff_A_dJ5c2YAM4_0),.clk(gclk));
	jdff dff_A_RZhauPO90_0(.dout(w_dff_A_cFFHib127_0),.din(w_dff_A_RZhauPO90_0),.clk(gclk));
	jdff dff_A_cFFHib127_0(.dout(w_dff_A_7QR5pUC97_0),.din(w_dff_A_cFFHib127_0),.clk(gclk));
	jdff dff_A_7QR5pUC97_0(.dout(w_dff_A_YP6GqKyh1_0),.din(w_dff_A_7QR5pUC97_0),.clk(gclk));
	jdff dff_A_YP6GqKyh1_0(.dout(w_dff_A_Z3yLKJJr0_0),.din(w_dff_A_YP6GqKyh1_0),.clk(gclk));
	jdff dff_A_Z3yLKJJr0_0(.dout(w_dff_A_n8oRfgRV9_0),.din(w_dff_A_Z3yLKJJr0_0),.clk(gclk));
	jdff dff_A_n8oRfgRV9_0(.dout(w_dff_A_0l0E9Php1_0),.din(w_dff_A_n8oRfgRV9_0),.clk(gclk));
	jdff dff_A_0l0E9Php1_0(.dout(w_dff_A_JOz6Y5zA2_0),.din(w_dff_A_0l0E9Php1_0),.clk(gclk));
	jdff dff_A_JOz6Y5zA2_0(.dout(w_dff_A_xgNSg37t8_0),.din(w_dff_A_JOz6Y5zA2_0),.clk(gclk));
	jdff dff_A_xgNSg37t8_0(.dout(w_dff_A_MDeAfenL1_0),.din(w_dff_A_xgNSg37t8_0),.clk(gclk));
	jdff dff_A_MDeAfenL1_0(.dout(w_dff_A_IUkC6Joo2_0),.din(w_dff_A_MDeAfenL1_0),.clk(gclk));
	jdff dff_A_IUkC6Joo2_0(.dout(w_dff_A_b3V2Ghm33_0),.din(w_dff_A_IUkC6Joo2_0),.clk(gclk));
	jdff dff_A_b3V2Ghm33_0(.dout(w_dff_A_yvOhH7523_0),.din(w_dff_A_b3V2Ghm33_0),.clk(gclk));
	jdff dff_A_yvOhH7523_0(.dout(w_dff_A_t2vfrKCz6_0),.din(w_dff_A_yvOhH7523_0),.clk(gclk));
	jdff dff_A_t2vfrKCz6_0(.dout(w_dff_A_BoOOBYC89_0),.din(w_dff_A_t2vfrKCz6_0),.clk(gclk));
	jdff dff_A_BoOOBYC89_0(.dout(G949),.din(w_dff_A_BoOOBYC89_0),.clk(gclk));
	jdff dff_A_SKPLdeyi8_1(.dout(w_dff_A_2qSTzhyE9_0),.din(w_dff_A_SKPLdeyi8_1),.clk(gclk));
	jdff dff_A_2qSTzhyE9_0(.dout(w_dff_A_nucsXvpf2_0),.din(w_dff_A_2qSTzhyE9_0),.clk(gclk));
	jdff dff_A_nucsXvpf2_0(.dout(w_dff_A_pJq5yQqh4_0),.din(w_dff_A_nucsXvpf2_0),.clk(gclk));
	jdff dff_A_pJq5yQqh4_0(.dout(w_dff_A_wu97i3l88_0),.din(w_dff_A_pJq5yQqh4_0),.clk(gclk));
	jdff dff_A_wu97i3l88_0(.dout(w_dff_A_5S0JHsZ41_0),.din(w_dff_A_wu97i3l88_0),.clk(gclk));
	jdff dff_A_5S0JHsZ41_0(.dout(w_dff_A_z7kyIMWU7_0),.din(w_dff_A_5S0JHsZ41_0),.clk(gclk));
	jdff dff_A_z7kyIMWU7_0(.dout(w_dff_A_PDVDedOh3_0),.din(w_dff_A_z7kyIMWU7_0),.clk(gclk));
	jdff dff_A_PDVDedOh3_0(.dout(w_dff_A_WVwJhwtm7_0),.din(w_dff_A_PDVDedOh3_0),.clk(gclk));
	jdff dff_A_WVwJhwtm7_0(.dout(w_dff_A_YwIrpcYa1_0),.din(w_dff_A_WVwJhwtm7_0),.clk(gclk));
	jdff dff_A_YwIrpcYa1_0(.dout(w_dff_A_xHz7VYgs1_0),.din(w_dff_A_YwIrpcYa1_0),.clk(gclk));
	jdff dff_A_xHz7VYgs1_0(.dout(w_dff_A_jXAdoxY40_0),.din(w_dff_A_xHz7VYgs1_0),.clk(gclk));
	jdff dff_A_jXAdoxY40_0(.dout(w_dff_A_OmOWHH8i7_0),.din(w_dff_A_jXAdoxY40_0),.clk(gclk));
	jdff dff_A_OmOWHH8i7_0(.dout(w_dff_A_u15K7vWv4_0),.din(w_dff_A_OmOWHH8i7_0),.clk(gclk));
	jdff dff_A_u15K7vWv4_0(.dout(w_dff_A_tLPxEEPG4_0),.din(w_dff_A_u15K7vWv4_0),.clk(gclk));
	jdff dff_A_tLPxEEPG4_0(.dout(w_dff_A_SalfHBKp8_0),.din(w_dff_A_tLPxEEPG4_0),.clk(gclk));
	jdff dff_A_SalfHBKp8_0(.dout(w_dff_A_X20frKLI7_0),.din(w_dff_A_SalfHBKp8_0),.clk(gclk));
	jdff dff_A_X20frKLI7_0(.dout(w_dff_A_ZA4oBV7I1_0),.din(w_dff_A_X20frKLI7_0),.clk(gclk));
	jdff dff_A_ZA4oBV7I1_0(.dout(w_dff_A_keFdkTBZ4_0),.din(w_dff_A_ZA4oBV7I1_0),.clk(gclk));
	jdff dff_A_keFdkTBZ4_0(.dout(w_dff_A_wH64j8n76_0),.din(w_dff_A_keFdkTBZ4_0),.clk(gclk));
	jdff dff_A_wH64j8n76_0(.dout(w_dff_A_qrSLvkpL6_0),.din(w_dff_A_wH64j8n76_0),.clk(gclk));
	jdff dff_A_qrSLvkpL6_0(.dout(w_dff_A_23jIzKqa0_0),.din(w_dff_A_qrSLvkpL6_0),.clk(gclk));
	jdff dff_A_23jIzKqa0_0(.dout(w_dff_A_xymuw4o74_0),.din(w_dff_A_23jIzKqa0_0),.clk(gclk));
	jdff dff_A_xymuw4o74_0(.dout(w_dff_A_pD3W7Z586_0),.din(w_dff_A_xymuw4o74_0),.clk(gclk));
	jdff dff_A_pD3W7Z586_0(.dout(w_dff_A_JFYKppkd0_0),.din(w_dff_A_pD3W7Z586_0),.clk(gclk));
	jdff dff_A_JFYKppkd0_0(.dout(w_dff_A_CcltRsG24_0),.din(w_dff_A_JFYKppkd0_0),.clk(gclk));
	jdff dff_A_CcltRsG24_0(.dout(w_dff_A_B2DvfHSf5_0),.din(w_dff_A_CcltRsG24_0),.clk(gclk));
	jdff dff_A_B2DvfHSf5_0(.dout(G939),.din(w_dff_A_B2DvfHSf5_0),.clk(gclk));
	jdff dff_A_Femo9NLV5_1(.dout(w_dff_A_NlHBCzV31_0),.din(w_dff_A_Femo9NLV5_1),.clk(gclk));
	jdff dff_A_NlHBCzV31_0(.dout(w_dff_A_wg5gnJ2k1_0),.din(w_dff_A_NlHBCzV31_0),.clk(gclk));
	jdff dff_A_wg5gnJ2k1_0(.dout(w_dff_A_P479h9P96_0),.din(w_dff_A_wg5gnJ2k1_0),.clk(gclk));
	jdff dff_A_P479h9P96_0(.dout(w_dff_A_HqpFnqCb7_0),.din(w_dff_A_P479h9P96_0),.clk(gclk));
	jdff dff_A_HqpFnqCb7_0(.dout(w_dff_A_PvnhAJg39_0),.din(w_dff_A_HqpFnqCb7_0),.clk(gclk));
	jdff dff_A_PvnhAJg39_0(.dout(w_dff_A_LZll5Fm78_0),.din(w_dff_A_PvnhAJg39_0),.clk(gclk));
	jdff dff_A_LZll5Fm78_0(.dout(w_dff_A_0z4SIJqg6_0),.din(w_dff_A_LZll5Fm78_0),.clk(gclk));
	jdff dff_A_0z4SIJqg6_0(.dout(w_dff_A_IFWuuGx01_0),.din(w_dff_A_0z4SIJqg6_0),.clk(gclk));
	jdff dff_A_IFWuuGx01_0(.dout(w_dff_A_XSxmljR30_0),.din(w_dff_A_IFWuuGx01_0),.clk(gclk));
	jdff dff_A_XSxmljR30_0(.dout(w_dff_A_BrKoEwES3_0),.din(w_dff_A_XSxmljR30_0),.clk(gclk));
	jdff dff_A_BrKoEwES3_0(.dout(w_dff_A_rYEawTOG9_0),.din(w_dff_A_BrKoEwES3_0),.clk(gclk));
	jdff dff_A_rYEawTOG9_0(.dout(w_dff_A_a7fR5RQd1_0),.din(w_dff_A_rYEawTOG9_0),.clk(gclk));
	jdff dff_A_a7fR5RQd1_0(.dout(w_dff_A_4IOJGG5X4_0),.din(w_dff_A_a7fR5RQd1_0),.clk(gclk));
	jdff dff_A_4IOJGG5X4_0(.dout(w_dff_A_W9iTcZTk2_0),.din(w_dff_A_4IOJGG5X4_0),.clk(gclk));
	jdff dff_A_W9iTcZTk2_0(.dout(w_dff_A_65rT7D2V2_0),.din(w_dff_A_W9iTcZTk2_0),.clk(gclk));
	jdff dff_A_65rT7D2V2_0(.dout(w_dff_A_FswOCQ1x5_0),.din(w_dff_A_65rT7D2V2_0),.clk(gclk));
	jdff dff_A_FswOCQ1x5_0(.dout(w_dff_A_rr1mzzEm5_0),.din(w_dff_A_FswOCQ1x5_0),.clk(gclk));
	jdff dff_A_rr1mzzEm5_0(.dout(w_dff_A_LzvWqzG99_0),.din(w_dff_A_rr1mzzEm5_0),.clk(gclk));
	jdff dff_A_LzvWqzG99_0(.dout(w_dff_A_qHF1pcbb0_0),.din(w_dff_A_LzvWqzG99_0),.clk(gclk));
	jdff dff_A_qHF1pcbb0_0(.dout(w_dff_A_OUaEY0X33_0),.din(w_dff_A_qHF1pcbb0_0),.clk(gclk));
	jdff dff_A_OUaEY0X33_0(.dout(w_dff_A_0iAljFpq4_0),.din(w_dff_A_OUaEY0X33_0),.clk(gclk));
	jdff dff_A_0iAljFpq4_0(.dout(w_dff_A_YPIditjM1_0),.din(w_dff_A_0iAljFpq4_0),.clk(gclk));
	jdff dff_A_YPIditjM1_0(.dout(w_dff_A_EN3CGhBf4_0),.din(w_dff_A_YPIditjM1_0),.clk(gclk));
	jdff dff_A_EN3CGhBf4_0(.dout(w_dff_A_W6UzBvUa9_0),.din(w_dff_A_EN3CGhBf4_0),.clk(gclk));
	jdff dff_A_W6UzBvUa9_0(.dout(w_dff_A_0gxnXOPP4_0),.din(w_dff_A_W6UzBvUa9_0),.clk(gclk));
	jdff dff_A_0gxnXOPP4_0(.dout(w_dff_A_0NxvzrgN0_0),.din(w_dff_A_0gxnXOPP4_0),.clk(gclk));
	jdff dff_A_0NxvzrgN0_0(.dout(G889),.din(w_dff_A_0NxvzrgN0_0),.clk(gclk));
	jdff dff_A_JlUsfOTy7_1(.dout(w_dff_A_3B9HwBPe0_0),.din(w_dff_A_JlUsfOTy7_1),.clk(gclk));
	jdff dff_A_3B9HwBPe0_0(.dout(w_dff_A_yStGtaew4_0),.din(w_dff_A_3B9HwBPe0_0),.clk(gclk));
	jdff dff_A_yStGtaew4_0(.dout(w_dff_A_jaLX8CQ02_0),.din(w_dff_A_yStGtaew4_0),.clk(gclk));
	jdff dff_A_jaLX8CQ02_0(.dout(w_dff_A_67wNSxP11_0),.din(w_dff_A_jaLX8CQ02_0),.clk(gclk));
	jdff dff_A_67wNSxP11_0(.dout(w_dff_A_GegosreC5_0),.din(w_dff_A_67wNSxP11_0),.clk(gclk));
	jdff dff_A_GegosreC5_0(.dout(w_dff_A_XHWoNeFP3_0),.din(w_dff_A_GegosreC5_0),.clk(gclk));
	jdff dff_A_XHWoNeFP3_0(.dout(w_dff_A_bLfiJvCO4_0),.din(w_dff_A_XHWoNeFP3_0),.clk(gclk));
	jdff dff_A_bLfiJvCO4_0(.dout(w_dff_A_BS0uVRY25_0),.din(w_dff_A_bLfiJvCO4_0),.clk(gclk));
	jdff dff_A_BS0uVRY25_0(.dout(w_dff_A_kVvwKqRh3_0),.din(w_dff_A_BS0uVRY25_0),.clk(gclk));
	jdff dff_A_kVvwKqRh3_0(.dout(w_dff_A_XGBQ3QtX9_0),.din(w_dff_A_kVvwKqRh3_0),.clk(gclk));
	jdff dff_A_XGBQ3QtX9_0(.dout(w_dff_A_MMY6qRtf4_0),.din(w_dff_A_XGBQ3QtX9_0),.clk(gclk));
	jdff dff_A_MMY6qRtf4_0(.dout(w_dff_A_j4alQXXo8_0),.din(w_dff_A_MMY6qRtf4_0),.clk(gclk));
	jdff dff_A_j4alQXXo8_0(.dout(w_dff_A_riaw58ne8_0),.din(w_dff_A_j4alQXXo8_0),.clk(gclk));
	jdff dff_A_riaw58ne8_0(.dout(w_dff_A_MN2uMMIk9_0),.din(w_dff_A_riaw58ne8_0),.clk(gclk));
	jdff dff_A_MN2uMMIk9_0(.dout(w_dff_A_XRWpcieE0_0),.din(w_dff_A_MN2uMMIk9_0),.clk(gclk));
	jdff dff_A_XRWpcieE0_0(.dout(w_dff_A_0IZ2WCww9_0),.din(w_dff_A_XRWpcieE0_0),.clk(gclk));
	jdff dff_A_0IZ2WCww9_0(.dout(w_dff_A_jKIJe3Cs1_0),.din(w_dff_A_0IZ2WCww9_0),.clk(gclk));
	jdff dff_A_jKIJe3Cs1_0(.dout(w_dff_A_Eon0llJ00_0),.din(w_dff_A_jKIJe3Cs1_0),.clk(gclk));
	jdff dff_A_Eon0llJ00_0(.dout(w_dff_A_I302w8E71_0),.din(w_dff_A_Eon0llJ00_0),.clk(gclk));
	jdff dff_A_I302w8E71_0(.dout(w_dff_A_WbLeyYaB7_0),.din(w_dff_A_I302w8E71_0),.clk(gclk));
	jdff dff_A_WbLeyYaB7_0(.dout(w_dff_A_WkftCjGB1_0),.din(w_dff_A_WbLeyYaB7_0),.clk(gclk));
	jdff dff_A_WkftCjGB1_0(.dout(w_dff_A_mPYVDaIn7_0),.din(w_dff_A_WkftCjGB1_0),.clk(gclk));
	jdff dff_A_mPYVDaIn7_0(.dout(w_dff_A_rzLVcdgv7_0),.din(w_dff_A_mPYVDaIn7_0),.clk(gclk));
	jdff dff_A_rzLVcdgv7_0(.dout(w_dff_A_xL5DAQUP6_0),.din(w_dff_A_rzLVcdgv7_0),.clk(gclk));
	jdff dff_A_xL5DAQUP6_0(.dout(w_dff_A_iTB1BQ4n3_0),.din(w_dff_A_xL5DAQUP6_0),.clk(gclk));
	jdff dff_A_iTB1BQ4n3_0(.dout(w_dff_A_lzRGMTWg1_0),.din(w_dff_A_iTB1BQ4n3_0),.clk(gclk));
	jdff dff_A_lzRGMTWg1_0(.dout(G593),.din(w_dff_A_lzRGMTWg1_0),.clk(gclk));
	jdff dff_A_ggxnG5mk7_2(.dout(w_dff_A_soGqoBSU8_0),.din(w_dff_A_ggxnG5mk7_2),.clk(gclk));
	jdff dff_A_soGqoBSU8_0(.dout(w_dff_A_a0JslDTl1_0),.din(w_dff_A_soGqoBSU8_0),.clk(gclk));
	jdff dff_A_a0JslDTl1_0(.dout(w_dff_A_zpTnZla65_0),.din(w_dff_A_a0JslDTl1_0),.clk(gclk));
	jdff dff_A_zpTnZla65_0(.dout(w_dff_A_tTRpNvXs0_0),.din(w_dff_A_zpTnZla65_0),.clk(gclk));
	jdff dff_A_tTRpNvXs0_0(.dout(w_dff_A_bjOdwmAc2_0),.din(w_dff_A_tTRpNvXs0_0),.clk(gclk));
	jdff dff_A_bjOdwmAc2_0(.dout(w_dff_A_YJ9ZAu3J6_0),.din(w_dff_A_bjOdwmAc2_0),.clk(gclk));
	jdff dff_A_YJ9ZAu3J6_0(.dout(w_dff_A_PixvskVl1_0),.din(w_dff_A_YJ9ZAu3J6_0),.clk(gclk));
	jdff dff_A_PixvskVl1_0(.dout(w_dff_A_p3qbVq8r3_0),.din(w_dff_A_PixvskVl1_0),.clk(gclk));
	jdff dff_A_p3qbVq8r3_0(.dout(w_dff_A_aW56xJAs5_0),.din(w_dff_A_p3qbVq8r3_0),.clk(gclk));
	jdff dff_A_aW56xJAs5_0(.dout(w_dff_A_3Wlp8vE85_0),.din(w_dff_A_aW56xJAs5_0),.clk(gclk));
	jdff dff_A_3Wlp8vE85_0(.dout(w_dff_A_E8mM1muW5_0),.din(w_dff_A_3Wlp8vE85_0),.clk(gclk));
	jdff dff_A_E8mM1muW5_0(.dout(w_dff_A_SLFWPjY44_0),.din(w_dff_A_E8mM1muW5_0),.clk(gclk));
	jdff dff_A_SLFWPjY44_0(.dout(w_dff_A_J8kL7Sgt9_0),.din(w_dff_A_SLFWPjY44_0),.clk(gclk));
	jdff dff_A_J8kL7Sgt9_0(.dout(w_dff_A_sw8PUaHd1_0),.din(w_dff_A_J8kL7Sgt9_0),.clk(gclk));
	jdff dff_A_sw8PUaHd1_0(.dout(w_dff_A_KIuylHh73_0),.din(w_dff_A_sw8PUaHd1_0),.clk(gclk));
	jdff dff_A_KIuylHh73_0(.dout(w_dff_A_sHYEi02l3_0),.din(w_dff_A_KIuylHh73_0),.clk(gclk));
	jdff dff_A_sHYEi02l3_0(.dout(w_dff_A_yUvjfvIO8_0),.din(w_dff_A_sHYEi02l3_0),.clk(gclk));
	jdff dff_A_yUvjfvIO8_0(.dout(w_dff_A_px2WHpYM5_0),.din(w_dff_A_yUvjfvIO8_0),.clk(gclk));
	jdff dff_A_px2WHpYM5_0(.dout(w_dff_A_zRF8JdTh0_0),.din(w_dff_A_px2WHpYM5_0),.clk(gclk));
	jdff dff_A_zRF8JdTh0_0(.dout(w_dff_A_9DUo6PBV2_0),.din(w_dff_A_zRF8JdTh0_0),.clk(gclk));
	jdff dff_A_9DUo6PBV2_0(.dout(w_dff_A_sgrLK5Oe7_0),.din(w_dff_A_9DUo6PBV2_0),.clk(gclk));
	jdff dff_A_sgrLK5Oe7_0(.dout(w_dff_A_8zEUF1Kx6_0),.din(w_dff_A_sgrLK5Oe7_0),.clk(gclk));
	jdff dff_A_8zEUF1Kx6_0(.dout(w_dff_A_r5BCFrqL9_0),.din(w_dff_A_8zEUF1Kx6_0),.clk(gclk));
	jdff dff_A_r5BCFrqL9_0(.dout(G636),.din(w_dff_A_r5BCFrqL9_0),.clk(gclk));
	jdff dff_A_9Fp90GiW7_2(.dout(w_dff_A_wkmp6lrl8_0),.din(w_dff_A_9Fp90GiW7_2),.clk(gclk));
	jdff dff_A_wkmp6lrl8_0(.dout(w_dff_A_Om9gIXYj8_0),.din(w_dff_A_wkmp6lrl8_0),.clk(gclk));
	jdff dff_A_Om9gIXYj8_0(.dout(w_dff_A_J8bKEIoc2_0),.din(w_dff_A_Om9gIXYj8_0),.clk(gclk));
	jdff dff_A_J8bKEIoc2_0(.dout(w_dff_A_1IR9LRMQ0_0),.din(w_dff_A_J8bKEIoc2_0),.clk(gclk));
	jdff dff_A_1IR9LRMQ0_0(.dout(w_dff_A_Q27Pe5oZ8_0),.din(w_dff_A_1IR9LRMQ0_0),.clk(gclk));
	jdff dff_A_Q27Pe5oZ8_0(.dout(w_dff_A_pmrRKuYQ3_0),.din(w_dff_A_Q27Pe5oZ8_0),.clk(gclk));
	jdff dff_A_pmrRKuYQ3_0(.dout(w_dff_A_HZstU9Dd0_0),.din(w_dff_A_pmrRKuYQ3_0),.clk(gclk));
	jdff dff_A_HZstU9Dd0_0(.dout(w_dff_A_3MOpmkng3_0),.din(w_dff_A_HZstU9Dd0_0),.clk(gclk));
	jdff dff_A_3MOpmkng3_0(.dout(w_dff_A_zYDO4QhQ1_0),.din(w_dff_A_3MOpmkng3_0),.clk(gclk));
	jdff dff_A_zYDO4QhQ1_0(.dout(w_dff_A_CgGxoC2F7_0),.din(w_dff_A_zYDO4QhQ1_0),.clk(gclk));
	jdff dff_A_CgGxoC2F7_0(.dout(w_dff_A_qWBRdyc79_0),.din(w_dff_A_CgGxoC2F7_0),.clk(gclk));
	jdff dff_A_qWBRdyc79_0(.dout(w_dff_A_D1H3cY1Z2_0),.din(w_dff_A_qWBRdyc79_0),.clk(gclk));
	jdff dff_A_D1H3cY1Z2_0(.dout(w_dff_A_0l9AKiTB8_0),.din(w_dff_A_D1H3cY1Z2_0),.clk(gclk));
	jdff dff_A_0l9AKiTB8_0(.dout(w_dff_A_XEqDzIra2_0),.din(w_dff_A_0l9AKiTB8_0),.clk(gclk));
	jdff dff_A_XEqDzIra2_0(.dout(w_dff_A_SWGWLOGt5_0),.din(w_dff_A_XEqDzIra2_0),.clk(gclk));
	jdff dff_A_SWGWLOGt5_0(.dout(w_dff_A_g2POdUbn9_0),.din(w_dff_A_SWGWLOGt5_0),.clk(gclk));
	jdff dff_A_g2POdUbn9_0(.dout(w_dff_A_n3wg9EoG8_0),.din(w_dff_A_g2POdUbn9_0),.clk(gclk));
	jdff dff_A_n3wg9EoG8_0(.dout(w_dff_A_tk4VvaVL2_0),.din(w_dff_A_n3wg9EoG8_0),.clk(gclk));
	jdff dff_A_tk4VvaVL2_0(.dout(w_dff_A_ViiQ19Ro7_0),.din(w_dff_A_tk4VvaVL2_0),.clk(gclk));
	jdff dff_A_ViiQ19Ro7_0(.dout(w_dff_A_snizAxlQ4_0),.din(w_dff_A_ViiQ19Ro7_0),.clk(gclk));
	jdff dff_A_snizAxlQ4_0(.dout(w_dff_A_gQzsw8tX0_0),.din(w_dff_A_snizAxlQ4_0),.clk(gclk));
	jdff dff_A_gQzsw8tX0_0(.dout(w_dff_A_ySsGHG3o4_0),.din(w_dff_A_gQzsw8tX0_0),.clk(gclk));
	jdff dff_A_ySsGHG3o4_0(.dout(w_dff_A_eJEs7m0C0_0),.din(w_dff_A_ySsGHG3o4_0),.clk(gclk));
	jdff dff_A_eJEs7m0C0_0(.dout(G704),.din(w_dff_A_eJEs7m0C0_0),.clk(gclk));
	jdff dff_A_BaD8i8TF9_2(.dout(w_dff_A_xjBKTD4I1_0),.din(w_dff_A_BaD8i8TF9_2),.clk(gclk));
	jdff dff_A_xjBKTD4I1_0(.dout(w_dff_A_6YM20goG0_0),.din(w_dff_A_xjBKTD4I1_0),.clk(gclk));
	jdff dff_A_6YM20goG0_0(.dout(w_dff_A_MElF77n31_0),.din(w_dff_A_6YM20goG0_0),.clk(gclk));
	jdff dff_A_MElF77n31_0(.dout(w_dff_A_xDGqj1qa7_0),.din(w_dff_A_MElF77n31_0),.clk(gclk));
	jdff dff_A_xDGqj1qa7_0(.dout(w_dff_A_gMJ0bC1b7_0),.din(w_dff_A_xDGqj1qa7_0),.clk(gclk));
	jdff dff_A_gMJ0bC1b7_0(.dout(w_dff_A_OZD5cGSG7_0),.din(w_dff_A_gMJ0bC1b7_0),.clk(gclk));
	jdff dff_A_OZD5cGSG7_0(.dout(w_dff_A_dgKvcHDk1_0),.din(w_dff_A_OZD5cGSG7_0),.clk(gclk));
	jdff dff_A_dgKvcHDk1_0(.dout(w_dff_A_PqCbBv3R6_0),.din(w_dff_A_dgKvcHDk1_0),.clk(gclk));
	jdff dff_A_PqCbBv3R6_0(.dout(w_dff_A_fAYB8dnB5_0),.din(w_dff_A_PqCbBv3R6_0),.clk(gclk));
	jdff dff_A_fAYB8dnB5_0(.dout(w_dff_A_JP7SyptP2_0),.din(w_dff_A_fAYB8dnB5_0),.clk(gclk));
	jdff dff_A_JP7SyptP2_0(.dout(w_dff_A_KI5jhp3e5_0),.din(w_dff_A_JP7SyptP2_0),.clk(gclk));
	jdff dff_A_KI5jhp3e5_0(.dout(w_dff_A_zwuUHvm75_0),.din(w_dff_A_KI5jhp3e5_0),.clk(gclk));
	jdff dff_A_zwuUHvm75_0(.dout(w_dff_A_otvnUqrg0_0),.din(w_dff_A_zwuUHvm75_0),.clk(gclk));
	jdff dff_A_otvnUqrg0_0(.dout(w_dff_A_NJ3uvGoa6_0),.din(w_dff_A_otvnUqrg0_0),.clk(gclk));
	jdff dff_A_NJ3uvGoa6_0(.dout(w_dff_A_3mvlPVQ53_0),.din(w_dff_A_NJ3uvGoa6_0),.clk(gclk));
	jdff dff_A_3mvlPVQ53_0(.dout(w_dff_A_DDumhluL6_0),.din(w_dff_A_3mvlPVQ53_0),.clk(gclk));
	jdff dff_A_DDumhluL6_0(.dout(w_dff_A_8IuzqLEW7_0),.din(w_dff_A_DDumhluL6_0),.clk(gclk));
	jdff dff_A_8IuzqLEW7_0(.dout(w_dff_A_boPSc9fI5_0),.din(w_dff_A_8IuzqLEW7_0),.clk(gclk));
	jdff dff_A_boPSc9fI5_0(.dout(w_dff_A_ESwuOz9u6_0),.din(w_dff_A_boPSc9fI5_0),.clk(gclk));
	jdff dff_A_ESwuOz9u6_0(.dout(w_dff_A_UANjooBs1_0),.din(w_dff_A_ESwuOz9u6_0),.clk(gclk));
	jdff dff_A_UANjooBs1_0(.dout(w_dff_A_ADvYnNf58_0),.din(w_dff_A_UANjooBs1_0),.clk(gclk));
	jdff dff_A_ADvYnNf58_0(.dout(w_dff_A_1CiA6Af43_0),.din(w_dff_A_ADvYnNf58_0),.clk(gclk));
	jdff dff_A_1CiA6Af43_0(.dout(w_dff_A_tzjUCfjA9_0),.din(w_dff_A_1CiA6Af43_0),.clk(gclk));
	jdff dff_A_tzjUCfjA9_0(.dout(G717),.din(w_dff_A_tzjUCfjA9_0),.clk(gclk));
	jdff dff_A_7aIGYmBt8_2(.dout(w_dff_A_fdslbe5r7_0),.din(w_dff_A_7aIGYmBt8_2),.clk(gclk));
	jdff dff_A_fdslbe5r7_0(.dout(w_dff_A_bgmIoIfr6_0),.din(w_dff_A_fdslbe5r7_0),.clk(gclk));
	jdff dff_A_bgmIoIfr6_0(.dout(w_dff_A_eB9DO8Xr2_0),.din(w_dff_A_bgmIoIfr6_0),.clk(gclk));
	jdff dff_A_eB9DO8Xr2_0(.dout(w_dff_A_FztlOzVp5_0),.din(w_dff_A_eB9DO8Xr2_0),.clk(gclk));
	jdff dff_A_FztlOzVp5_0(.dout(w_dff_A_GKY3LsMV0_0),.din(w_dff_A_FztlOzVp5_0),.clk(gclk));
	jdff dff_A_GKY3LsMV0_0(.dout(w_dff_A_iNwDsvSD2_0),.din(w_dff_A_GKY3LsMV0_0),.clk(gclk));
	jdff dff_A_iNwDsvSD2_0(.dout(w_dff_A_xER18dRt8_0),.din(w_dff_A_iNwDsvSD2_0),.clk(gclk));
	jdff dff_A_xER18dRt8_0(.dout(w_dff_A_Vw79pbN41_0),.din(w_dff_A_xER18dRt8_0),.clk(gclk));
	jdff dff_A_Vw79pbN41_0(.dout(w_dff_A_eD7oyL8r7_0),.din(w_dff_A_Vw79pbN41_0),.clk(gclk));
	jdff dff_A_eD7oyL8r7_0(.dout(w_dff_A_QnfkqptZ9_0),.din(w_dff_A_eD7oyL8r7_0),.clk(gclk));
	jdff dff_A_QnfkqptZ9_0(.dout(w_dff_A_qkJJt8qk1_0),.din(w_dff_A_QnfkqptZ9_0),.clk(gclk));
	jdff dff_A_qkJJt8qk1_0(.dout(w_dff_A_v32xaZdh5_0),.din(w_dff_A_qkJJt8qk1_0),.clk(gclk));
	jdff dff_A_v32xaZdh5_0(.dout(w_dff_A_EpydQUZR8_0),.din(w_dff_A_v32xaZdh5_0),.clk(gclk));
	jdff dff_A_EpydQUZR8_0(.dout(w_dff_A_oIQ15tVM3_0),.din(w_dff_A_EpydQUZR8_0),.clk(gclk));
	jdff dff_A_oIQ15tVM3_0(.dout(w_dff_A_FecwbBKd7_0),.din(w_dff_A_oIQ15tVM3_0),.clk(gclk));
	jdff dff_A_FecwbBKd7_0(.dout(w_dff_A_DJp5nEX43_0),.din(w_dff_A_FecwbBKd7_0),.clk(gclk));
	jdff dff_A_DJp5nEX43_0(.dout(w_dff_A_fagqzMmt2_0),.din(w_dff_A_DJp5nEX43_0),.clk(gclk));
	jdff dff_A_fagqzMmt2_0(.dout(w_dff_A_t6mYyL5t3_0),.din(w_dff_A_fagqzMmt2_0),.clk(gclk));
	jdff dff_A_t6mYyL5t3_0(.dout(w_dff_A_fdUuXirF3_0),.din(w_dff_A_t6mYyL5t3_0),.clk(gclk));
	jdff dff_A_fdUuXirF3_0(.dout(w_dff_A_sc2fG96P1_0),.din(w_dff_A_fdUuXirF3_0),.clk(gclk));
	jdff dff_A_sc2fG96P1_0(.dout(w_dff_A_lm5H9nBY1_0),.din(w_dff_A_sc2fG96P1_0),.clk(gclk));
	jdff dff_A_lm5H9nBY1_0(.dout(w_dff_A_adDaodPF2_0),.din(w_dff_A_lm5H9nBY1_0),.clk(gclk));
	jdff dff_A_adDaodPF2_0(.dout(w_dff_A_RpYPwKbW1_0),.din(w_dff_A_adDaodPF2_0),.clk(gclk));
	jdff dff_A_RpYPwKbW1_0(.dout(w_dff_A_22ycq4ex2_0),.din(w_dff_A_RpYPwKbW1_0),.clk(gclk));
	jdff dff_A_22ycq4ex2_0(.dout(G820),.din(w_dff_A_22ycq4ex2_0),.clk(gclk));
	jdff dff_A_oXh5hHFP5_2(.dout(w_dff_A_4LtYUCoT8_0),.din(w_dff_A_oXh5hHFP5_2),.clk(gclk));
	jdff dff_A_4LtYUCoT8_0(.dout(w_dff_A_4iVz71ut0_0),.din(w_dff_A_4LtYUCoT8_0),.clk(gclk));
	jdff dff_A_4iVz71ut0_0(.dout(w_dff_A_IWIDMaw86_0),.din(w_dff_A_4iVz71ut0_0),.clk(gclk));
	jdff dff_A_IWIDMaw86_0(.dout(w_dff_A_XkkHFvoO4_0),.din(w_dff_A_IWIDMaw86_0),.clk(gclk));
	jdff dff_A_XkkHFvoO4_0(.dout(w_dff_A_IaQB31nO0_0),.din(w_dff_A_XkkHFvoO4_0),.clk(gclk));
	jdff dff_A_IaQB31nO0_0(.dout(w_dff_A_CfsQocWg1_0),.din(w_dff_A_IaQB31nO0_0),.clk(gclk));
	jdff dff_A_CfsQocWg1_0(.dout(w_dff_A_eHgmuEbK1_0),.din(w_dff_A_CfsQocWg1_0),.clk(gclk));
	jdff dff_A_eHgmuEbK1_0(.dout(w_dff_A_pqbmqe2y1_0),.din(w_dff_A_eHgmuEbK1_0),.clk(gclk));
	jdff dff_A_pqbmqe2y1_0(.dout(w_dff_A_lcQfdGmx4_0),.din(w_dff_A_pqbmqe2y1_0),.clk(gclk));
	jdff dff_A_lcQfdGmx4_0(.dout(w_dff_A_8QrI6YU44_0),.din(w_dff_A_lcQfdGmx4_0),.clk(gclk));
	jdff dff_A_8QrI6YU44_0(.dout(w_dff_A_nX2fVv7i5_0),.din(w_dff_A_8QrI6YU44_0),.clk(gclk));
	jdff dff_A_nX2fVv7i5_0(.dout(w_dff_A_2lH3SzDG5_0),.din(w_dff_A_nX2fVv7i5_0),.clk(gclk));
	jdff dff_A_2lH3SzDG5_0(.dout(w_dff_A_JjVnmOAe2_0),.din(w_dff_A_2lH3SzDG5_0),.clk(gclk));
	jdff dff_A_JjVnmOAe2_0(.dout(w_dff_A_uWwO6c0V0_0),.din(w_dff_A_JjVnmOAe2_0),.clk(gclk));
	jdff dff_A_uWwO6c0V0_0(.dout(w_dff_A_Scr4Xdlr9_0),.din(w_dff_A_uWwO6c0V0_0),.clk(gclk));
	jdff dff_A_Scr4Xdlr9_0(.dout(w_dff_A_MNmT17kz0_0),.din(w_dff_A_Scr4Xdlr9_0),.clk(gclk));
	jdff dff_A_MNmT17kz0_0(.dout(w_dff_A_4NhZrj4o5_0),.din(w_dff_A_MNmT17kz0_0),.clk(gclk));
	jdff dff_A_4NhZrj4o5_0(.dout(w_dff_A_Z3M9vFrv1_0),.din(w_dff_A_4NhZrj4o5_0),.clk(gclk));
	jdff dff_A_Z3M9vFrv1_0(.dout(w_dff_A_HweYZHgk8_0),.din(w_dff_A_Z3M9vFrv1_0),.clk(gclk));
	jdff dff_A_HweYZHgk8_0(.dout(w_dff_A_yykWYldi2_0),.din(w_dff_A_HweYZHgk8_0),.clk(gclk));
	jdff dff_A_yykWYldi2_0(.dout(w_dff_A_9OoTzEzV7_0),.din(w_dff_A_yykWYldi2_0),.clk(gclk));
	jdff dff_A_9OoTzEzV7_0(.dout(w_dff_A_Zlckauki5_0),.din(w_dff_A_9OoTzEzV7_0),.clk(gclk));
	jdff dff_A_Zlckauki5_0(.dout(G639),.din(w_dff_A_Zlckauki5_0),.clk(gclk));
	jdff dff_A_4VBlrx7w2_2(.dout(w_dff_A_BIlgfuI73_0),.din(w_dff_A_4VBlrx7w2_2),.clk(gclk));
	jdff dff_A_BIlgfuI73_0(.dout(w_dff_A_uXeSAsFX3_0),.din(w_dff_A_BIlgfuI73_0),.clk(gclk));
	jdff dff_A_uXeSAsFX3_0(.dout(w_dff_A_VomWAx9P1_0),.din(w_dff_A_uXeSAsFX3_0),.clk(gclk));
	jdff dff_A_VomWAx9P1_0(.dout(w_dff_A_sRlKKdnF4_0),.din(w_dff_A_VomWAx9P1_0),.clk(gclk));
	jdff dff_A_sRlKKdnF4_0(.dout(w_dff_A_duknT22U1_0),.din(w_dff_A_sRlKKdnF4_0),.clk(gclk));
	jdff dff_A_duknT22U1_0(.dout(w_dff_A_HALbsMQM1_0),.din(w_dff_A_duknT22U1_0),.clk(gclk));
	jdff dff_A_HALbsMQM1_0(.dout(w_dff_A_qKlXLPIF0_0),.din(w_dff_A_HALbsMQM1_0),.clk(gclk));
	jdff dff_A_qKlXLPIF0_0(.dout(w_dff_A_VXSzI9iX9_0),.din(w_dff_A_qKlXLPIF0_0),.clk(gclk));
	jdff dff_A_VXSzI9iX9_0(.dout(w_dff_A_xcijaDCS4_0),.din(w_dff_A_VXSzI9iX9_0),.clk(gclk));
	jdff dff_A_xcijaDCS4_0(.dout(w_dff_A_5X1gZXtG7_0),.din(w_dff_A_xcijaDCS4_0),.clk(gclk));
	jdff dff_A_5X1gZXtG7_0(.dout(w_dff_A_lRDBTsYm8_0),.din(w_dff_A_5X1gZXtG7_0),.clk(gclk));
	jdff dff_A_lRDBTsYm8_0(.dout(w_dff_A_MYOlMxxt1_0),.din(w_dff_A_lRDBTsYm8_0),.clk(gclk));
	jdff dff_A_MYOlMxxt1_0(.dout(w_dff_A_JdmnnDJw6_0),.din(w_dff_A_MYOlMxxt1_0),.clk(gclk));
	jdff dff_A_JdmnnDJw6_0(.dout(w_dff_A_Dn4OQfkn4_0),.din(w_dff_A_JdmnnDJw6_0),.clk(gclk));
	jdff dff_A_Dn4OQfkn4_0(.dout(w_dff_A_6ygsp5KJ0_0),.din(w_dff_A_Dn4OQfkn4_0),.clk(gclk));
	jdff dff_A_6ygsp5KJ0_0(.dout(w_dff_A_rh6YIwCc6_0),.din(w_dff_A_6ygsp5KJ0_0),.clk(gclk));
	jdff dff_A_rh6YIwCc6_0(.dout(w_dff_A_S0F2NR0R8_0),.din(w_dff_A_rh6YIwCc6_0),.clk(gclk));
	jdff dff_A_S0F2NR0R8_0(.dout(w_dff_A_FwX7Takh2_0),.din(w_dff_A_S0F2NR0R8_0),.clk(gclk));
	jdff dff_A_FwX7Takh2_0(.dout(w_dff_A_N3KcFBa32_0),.din(w_dff_A_FwX7Takh2_0),.clk(gclk));
	jdff dff_A_N3KcFBa32_0(.dout(w_dff_A_LoEkIqHu8_0),.din(w_dff_A_N3KcFBa32_0),.clk(gclk));
	jdff dff_A_LoEkIqHu8_0(.dout(w_dff_A_euh4H7FH7_0),.din(w_dff_A_LoEkIqHu8_0),.clk(gclk));
	jdff dff_A_euh4H7FH7_0(.dout(w_dff_A_McPKAUHR9_0),.din(w_dff_A_euh4H7FH7_0),.clk(gclk));
	jdff dff_A_McPKAUHR9_0(.dout(G673),.din(w_dff_A_McPKAUHR9_0),.clk(gclk));
	jdff dff_A_TnyExUOt6_2(.dout(w_dff_A_m2QxoPEi7_0),.din(w_dff_A_TnyExUOt6_2),.clk(gclk));
	jdff dff_A_m2QxoPEi7_0(.dout(w_dff_A_6DCS2fUy9_0),.din(w_dff_A_m2QxoPEi7_0),.clk(gclk));
	jdff dff_A_6DCS2fUy9_0(.dout(w_dff_A_QxOHOkW36_0),.din(w_dff_A_6DCS2fUy9_0),.clk(gclk));
	jdff dff_A_QxOHOkW36_0(.dout(w_dff_A_jyRVJxNl4_0),.din(w_dff_A_QxOHOkW36_0),.clk(gclk));
	jdff dff_A_jyRVJxNl4_0(.dout(w_dff_A_BUaKj3Nn2_0),.din(w_dff_A_jyRVJxNl4_0),.clk(gclk));
	jdff dff_A_BUaKj3Nn2_0(.dout(w_dff_A_Ti9mOnCh1_0),.din(w_dff_A_BUaKj3Nn2_0),.clk(gclk));
	jdff dff_A_Ti9mOnCh1_0(.dout(w_dff_A_VuWBPtCy4_0),.din(w_dff_A_Ti9mOnCh1_0),.clk(gclk));
	jdff dff_A_VuWBPtCy4_0(.dout(w_dff_A_NFPZ5n9V4_0),.din(w_dff_A_VuWBPtCy4_0),.clk(gclk));
	jdff dff_A_NFPZ5n9V4_0(.dout(w_dff_A_QyhQHejV1_0),.din(w_dff_A_NFPZ5n9V4_0),.clk(gclk));
	jdff dff_A_QyhQHejV1_0(.dout(w_dff_A_HtsmvrZi3_0),.din(w_dff_A_QyhQHejV1_0),.clk(gclk));
	jdff dff_A_HtsmvrZi3_0(.dout(w_dff_A_T4XC26Jg7_0),.din(w_dff_A_HtsmvrZi3_0),.clk(gclk));
	jdff dff_A_T4XC26Jg7_0(.dout(w_dff_A_nFvlLH8c1_0),.din(w_dff_A_T4XC26Jg7_0),.clk(gclk));
	jdff dff_A_nFvlLH8c1_0(.dout(w_dff_A_OShEDruo9_0),.din(w_dff_A_nFvlLH8c1_0),.clk(gclk));
	jdff dff_A_OShEDruo9_0(.dout(w_dff_A_GGdVLRBB7_0),.din(w_dff_A_OShEDruo9_0),.clk(gclk));
	jdff dff_A_GGdVLRBB7_0(.dout(w_dff_A_rFgGl2NK4_0),.din(w_dff_A_GGdVLRBB7_0),.clk(gclk));
	jdff dff_A_rFgGl2NK4_0(.dout(w_dff_A_VahjnZhW6_0),.din(w_dff_A_rFgGl2NK4_0),.clk(gclk));
	jdff dff_A_VahjnZhW6_0(.dout(w_dff_A_DEaQaxxT2_0),.din(w_dff_A_VahjnZhW6_0),.clk(gclk));
	jdff dff_A_DEaQaxxT2_0(.dout(w_dff_A_gUfDPPDN6_0),.din(w_dff_A_DEaQaxxT2_0),.clk(gclk));
	jdff dff_A_gUfDPPDN6_0(.dout(w_dff_A_8afGv2pz2_0),.din(w_dff_A_gUfDPPDN6_0),.clk(gclk));
	jdff dff_A_8afGv2pz2_0(.dout(w_dff_A_3lv0jjFW6_0),.din(w_dff_A_8afGv2pz2_0),.clk(gclk));
	jdff dff_A_3lv0jjFW6_0(.dout(w_dff_A_YmzDT3ym0_0),.din(w_dff_A_3lv0jjFW6_0),.clk(gclk));
	jdff dff_A_YmzDT3ym0_0(.dout(w_dff_A_IfE1XxdW2_0),.din(w_dff_A_YmzDT3ym0_0),.clk(gclk));
	jdff dff_A_IfE1XxdW2_0(.dout(G707),.din(w_dff_A_IfE1XxdW2_0),.clk(gclk));
	jdff dff_A_jviPCy004_2(.dout(w_dff_A_04uaOXrN9_0),.din(w_dff_A_jviPCy004_2),.clk(gclk));
	jdff dff_A_04uaOXrN9_0(.dout(w_dff_A_UdbLiJgG5_0),.din(w_dff_A_04uaOXrN9_0),.clk(gclk));
	jdff dff_A_UdbLiJgG5_0(.dout(w_dff_A_MzDfdB4P0_0),.din(w_dff_A_UdbLiJgG5_0),.clk(gclk));
	jdff dff_A_MzDfdB4P0_0(.dout(w_dff_A_SxgIrgyv4_0),.din(w_dff_A_MzDfdB4P0_0),.clk(gclk));
	jdff dff_A_SxgIrgyv4_0(.dout(w_dff_A_MHWEKNgO1_0),.din(w_dff_A_SxgIrgyv4_0),.clk(gclk));
	jdff dff_A_MHWEKNgO1_0(.dout(w_dff_A_WGdGq7Ey9_0),.din(w_dff_A_MHWEKNgO1_0),.clk(gclk));
	jdff dff_A_WGdGq7Ey9_0(.dout(w_dff_A_OxGqiwtK2_0),.din(w_dff_A_WGdGq7Ey9_0),.clk(gclk));
	jdff dff_A_OxGqiwtK2_0(.dout(w_dff_A_y1IPsVse8_0),.din(w_dff_A_OxGqiwtK2_0),.clk(gclk));
	jdff dff_A_y1IPsVse8_0(.dout(w_dff_A_2B6Q3m830_0),.din(w_dff_A_y1IPsVse8_0),.clk(gclk));
	jdff dff_A_2B6Q3m830_0(.dout(w_dff_A_LX8HlE9g4_0),.din(w_dff_A_2B6Q3m830_0),.clk(gclk));
	jdff dff_A_LX8HlE9g4_0(.dout(w_dff_A_xk5ejCSe6_0),.din(w_dff_A_LX8HlE9g4_0),.clk(gclk));
	jdff dff_A_xk5ejCSe6_0(.dout(w_dff_A_BaoSDj0W1_0),.din(w_dff_A_xk5ejCSe6_0),.clk(gclk));
	jdff dff_A_BaoSDj0W1_0(.dout(w_dff_A_5cs0LYHE3_0),.din(w_dff_A_BaoSDj0W1_0),.clk(gclk));
	jdff dff_A_5cs0LYHE3_0(.dout(w_dff_A_Ex6JadYn8_0),.din(w_dff_A_5cs0LYHE3_0),.clk(gclk));
	jdff dff_A_Ex6JadYn8_0(.dout(w_dff_A_fTvKbmDP0_0),.din(w_dff_A_Ex6JadYn8_0),.clk(gclk));
	jdff dff_A_fTvKbmDP0_0(.dout(w_dff_A_4mydeKCB9_0),.din(w_dff_A_fTvKbmDP0_0),.clk(gclk));
	jdff dff_A_4mydeKCB9_0(.dout(w_dff_A_0ozEw7dI5_0),.din(w_dff_A_4mydeKCB9_0),.clk(gclk));
	jdff dff_A_0ozEw7dI5_0(.dout(w_dff_A_K9IfZtmH3_0),.din(w_dff_A_0ozEw7dI5_0),.clk(gclk));
	jdff dff_A_K9IfZtmH3_0(.dout(w_dff_A_rJ51SNR76_0),.din(w_dff_A_K9IfZtmH3_0),.clk(gclk));
	jdff dff_A_rJ51SNR76_0(.dout(w_dff_A_4YzD4k2h4_0),.din(w_dff_A_rJ51SNR76_0),.clk(gclk));
	jdff dff_A_4YzD4k2h4_0(.dout(w_dff_A_dYaBkdA04_0),.din(w_dff_A_4YzD4k2h4_0),.clk(gclk));
	jdff dff_A_dYaBkdA04_0(.dout(w_dff_A_u6GnkU9e7_0),.din(w_dff_A_dYaBkdA04_0),.clk(gclk));
	jdff dff_A_u6GnkU9e7_0(.dout(G715),.din(w_dff_A_u6GnkU9e7_0),.clk(gclk));
	jdff dff_A_FCzrs7lI1_2(.dout(w_dff_A_ahcWene33_0),.din(w_dff_A_FCzrs7lI1_2),.clk(gclk));
	jdff dff_A_ahcWene33_0(.dout(w_dff_A_E4ut34AA3_0),.din(w_dff_A_ahcWene33_0),.clk(gclk));
	jdff dff_A_E4ut34AA3_0(.dout(w_dff_A_lZiDdcn39_0),.din(w_dff_A_E4ut34AA3_0),.clk(gclk));
	jdff dff_A_lZiDdcn39_0(.dout(w_dff_A_irKjk10M5_0),.din(w_dff_A_lZiDdcn39_0),.clk(gclk));
	jdff dff_A_irKjk10M5_0(.dout(w_dff_A_7ouXLBM22_0),.din(w_dff_A_irKjk10M5_0),.clk(gclk));
	jdff dff_A_7ouXLBM22_0(.dout(w_dff_A_GP3KJ3lY1_0),.din(w_dff_A_7ouXLBM22_0),.clk(gclk));
	jdff dff_A_GP3KJ3lY1_0(.dout(w_dff_A_0rpV5NER2_0),.din(w_dff_A_GP3KJ3lY1_0),.clk(gclk));
	jdff dff_A_0rpV5NER2_0(.dout(w_dff_A_M6Sqze256_0),.din(w_dff_A_0rpV5NER2_0),.clk(gclk));
	jdff dff_A_M6Sqze256_0(.dout(w_dff_A_yZ8dW7Bl7_0),.din(w_dff_A_M6Sqze256_0),.clk(gclk));
	jdff dff_A_yZ8dW7Bl7_0(.dout(w_dff_A_Cbq7JKkt2_0),.din(w_dff_A_yZ8dW7Bl7_0),.clk(gclk));
	jdff dff_A_Cbq7JKkt2_0(.dout(w_dff_A_3zy9uUce6_0),.din(w_dff_A_Cbq7JKkt2_0),.clk(gclk));
	jdff dff_A_3zy9uUce6_0(.dout(w_dff_A_gLx2fgw39_0),.din(w_dff_A_3zy9uUce6_0),.clk(gclk));
	jdff dff_A_gLx2fgw39_0(.dout(w_dff_A_GvvLizGC0_0),.din(w_dff_A_gLx2fgw39_0),.clk(gclk));
	jdff dff_A_GvvLizGC0_0(.dout(w_dff_A_MfhM0JDk7_0),.din(w_dff_A_GvvLizGC0_0),.clk(gclk));
	jdff dff_A_MfhM0JDk7_0(.dout(w_dff_A_yLhM6FhX1_0),.din(w_dff_A_MfhM0JDk7_0),.clk(gclk));
	jdff dff_A_yLhM6FhX1_0(.dout(w_dff_A_Gvzo9Uf08_0),.din(w_dff_A_yLhM6FhX1_0),.clk(gclk));
	jdff dff_A_Gvzo9Uf08_0(.dout(w_dff_A_IOssKhkH6_0),.din(w_dff_A_Gvzo9Uf08_0),.clk(gclk));
	jdff dff_A_IOssKhkH6_0(.dout(w_dff_A_h5pezWX06_0),.din(w_dff_A_IOssKhkH6_0),.clk(gclk));
	jdff dff_A_h5pezWX06_0(.dout(w_dff_A_54HgQfUU5_0),.din(w_dff_A_h5pezWX06_0),.clk(gclk));
	jdff dff_A_54HgQfUU5_0(.dout(G598),.din(w_dff_A_54HgQfUU5_0),.clk(gclk));
	jdff dff_A_w6ptbcNI1_2(.dout(w_dff_A_wKcYnG6L0_0),.din(w_dff_A_w6ptbcNI1_2),.clk(gclk));
	jdff dff_A_wKcYnG6L0_0(.dout(w_dff_A_WLfds1zs2_0),.din(w_dff_A_wKcYnG6L0_0),.clk(gclk));
	jdff dff_A_WLfds1zs2_0(.dout(w_dff_A_t8op28g67_0),.din(w_dff_A_WLfds1zs2_0),.clk(gclk));
	jdff dff_A_t8op28g67_0(.dout(w_dff_A_JHfpfx4h0_0),.din(w_dff_A_t8op28g67_0),.clk(gclk));
	jdff dff_A_JHfpfx4h0_0(.dout(w_dff_A_2RMLKFdb4_0),.din(w_dff_A_JHfpfx4h0_0),.clk(gclk));
	jdff dff_A_2RMLKFdb4_0(.dout(w_dff_A_DDD1tYNc4_0),.din(w_dff_A_2RMLKFdb4_0),.clk(gclk));
	jdff dff_A_DDD1tYNc4_0(.dout(w_dff_A_s0hmulKZ0_0),.din(w_dff_A_DDD1tYNc4_0),.clk(gclk));
	jdff dff_A_s0hmulKZ0_0(.dout(w_dff_A_A9p0smSx1_0),.din(w_dff_A_s0hmulKZ0_0),.clk(gclk));
	jdff dff_A_A9p0smSx1_0(.dout(w_dff_A_Cj9sbDPR6_0),.din(w_dff_A_A9p0smSx1_0),.clk(gclk));
	jdff dff_A_Cj9sbDPR6_0(.dout(w_dff_A_Kod3pKDV5_0),.din(w_dff_A_Cj9sbDPR6_0),.clk(gclk));
	jdff dff_A_Kod3pKDV5_0(.dout(w_dff_A_7xhQmYh16_0),.din(w_dff_A_Kod3pKDV5_0),.clk(gclk));
	jdff dff_A_7xhQmYh16_0(.dout(w_dff_A_vG0ZTohM3_0),.din(w_dff_A_7xhQmYh16_0),.clk(gclk));
	jdff dff_A_vG0ZTohM3_0(.dout(w_dff_A_QvoG1XTB6_0),.din(w_dff_A_vG0ZTohM3_0),.clk(gclk));
	jdff dff_A_QvoG1XTB6_0(.dout(w_dff_A_e1pzCSdJ9_0),.din(w_dff_A_QvoG1XTB6_0),.clk(gclk));
	jdff dff_A_e1pzCSdJ9_0(.dout(w_dff_A_CzWkz3IL9_0),.din(w_dff_A_e1pzCSdJ9_0),.clk(gclk));
	jdff dff_A_CzWkz3IL9_0(.dout(w_dff_A_bhbvxTPo5_0),.din(w_dff_A_CzWkz3IL9_0),.clk(gclk));
	jdff dff_A_bhbvxTPo5_0(.dout(w_dff_A_YBZbAwDs7_0),.din(w_dff_A_bhbvxTPo5_0),.clk(gclk));
	jdff dff_A_YBZbAwDs7_0(.dout(w_dff_A_bi0nBdus6_0),.din(w_dff_A_YBZbAwDs7_0),.clk(gclk));
	jdff dff_A_bi0nBdus6_0(.dout(G610),.din(w_dff_A_bi0nBdus6_0),.clk(gclk));
	jdff dff_A_hjs3pf4K4_2(.dout(w_dff_A_xktMmrAI2_0),.din(w_dff_A_hjs3pf4K4_2),.clk(gclk));
	jdff dff_A_xktMmrAI2_0(.dout(w_dff_A_B0XsbOgY5_0),.din(w_dff_A_xktMmrAI2_0),.clk(gclk));
	jdff dff_A_B0XsbOgY5_0(.dout(w_dff_A_hSHgTJH43_0),.din(w_dff_A_B0XsbOgY5_0),.clk(gclk));
	jdff dff_A_hSHgTJH43_0(.dout(w_dff_A_bhUEti0a3_0),.din(w_dff_A_hSHgTJH43_0),.clk(gclk));
	jdff dff_A_bhUEti0a3_0(.dout(w_dff_A_LFUSm4GD1_0),.din(w_dff_A_bhUEti0a3_0),.clk(gclk));
	jdff dff_A_LFUSm4GD1_0(.dout(w_dff_A_uUDNsvUN0_0),.din(w_dff_A_LFUSm4GD1_0),.clk(gclk));
	jdff dff_A_uUDNsvUN0_0(.dout(w_dff_A_ypLymG1f1_0),.din(w_dff_A_uUDNsvUN0_0),.clk(gclk));
	jdff dff_A_ypLymG1f1_0(.dout(w_dff_A_Wl3MkFn20_0),.din(w_dff_A_ypLymG1f1_0),.clk(gclk));
	jdff dff_A_Wl3MkFn20_0(.dout(w_dff_A_JT2tdUVw6_0),.din(w_dff_A_Wl3MkFn20_0),.clk(gclk));
	jdff dff_A_JT2tdUVw6_0(.dout(w_dff_A_OHzqKTJu2_0),.din(w_dff_A_JT2tdUVw6_0),.clk(gclk));
	jdff dff_A_OHzqKTJu2_0(.dout(w_dff_A_Kmwsm5hn3_0),.din(w_dff_A_OHzqKTJu2_0),.clk(gclk));
	jdff dff_A_Kmwsm5hn3_0(.dout(w_dff_A_1hSgZx2J6_0),.din(w_dff_A_Kmwsm5hn3_0),.clk(gclk));
	jdff dff_A_1hSgZx2J6_0(.dout(w_dff_A_mtPWx4Va4_0),.din(w_dff_A_1hSgZx2J6_0),.clk(gclk));
	jdff dff_A_mtPWx4Va4_0(.dout(w_dff_A_DmnnXYYn4_0),.din(w_dff_A_mtPWx4Va4_0),.clk(gclk));
	jdff dff_A_DmnnXYYn4_0(.dout(w_dff_A_UJa8BsNY4_0),.din(w_dff_A_DmnnXYYn4_0),.clk(gclk));
	jdff dff_A_UJa8BsNY4_0(.dout(w_dff_A_l2uks8bl3_0),.din(w_dff_A_UJa8BsNY4_0),.clk(gclk));
	jdff dff_A_l2uks8bl3_0(.dout(G588),.din(w_dff_A_l2uks8bl3_0),.clk(gclk));
	jdff dff_A_QVvvToBY8_2(.dout(w_dff_A_r8UDSSn76_0),.din(w_dff_A_QVvvToBY8_2),.clk(gclk));
	jdff dff_A_r8UDSSn76_0(.dout(w_dff_A_6fgyXfer9_0),.din(w_dff_A_r8UDSSn76_0),.clk(gclk));
	jdff dff_A_6fgyXfer9_0(.dout(w_dff_A_zTl1PCT15_0),.din(w_dff_A_6fgyXfer9_0),.clk(gclk));
	jdff dff_A_zTl1PCT15_0(.dout(w_dff_A_favJvT4u8_0),.din(w_dff_A_zTl1PCT15_0),.clk(gclk));
	jdff dff_A_favJvT4u8_0(.dout(w_dff_A_udDgwovk2_0),.din(w_dff_A_favJvT4u8_0),.clk(gclk));
	jdff dff_A_udDgwovk2_0(.dout(w_dff_A_fikQLPbe8_0),.din(w_dff_A_udDgwovk2_0),.clk(gclk));
	jdff dff_A_fikQLPbe8_0(.dout(w_dff_A_QRgNZbL06_0),.din(w_dff_A_fikQLPbe8_0),.clk(gclk));
	jdff dff_A_QRgNZbL06_0(.dout(w_dff_A_A1BnklJE4_0),.din(w_dff_A_QRgNZbL06_0),.clk(gclk));
	jdff dff_A_A1BnklJE4_0(.dout(w_dff_A_ZOKzsVmy0_0),.din(w_dff_A_A1BnklJE4_0),.clk(gclk));
	jdff dff_A_ZOKzsVmy0_0(.dout(w_dff_A_L6JCwsmY9_0),.din(w_dff_A_ZOKzsVmy0_0),.clk(gclk));
	jdff dff_A_L6JCwsmY9_0(.dout(w_dff_A_VdTOdjVu4_0),.din(w_dff_A_L6JCwsmY9_0),.clk(gclk));
	jdff dff_A_VdTOdjVu4_0(.dout(w_dff_A_1haxGdVJ2_0),.din(w_dff_A_VdTOdjVu4_0),.clk(gclk));
	jdff dff_A_1haxGdVJ2_0(.dout(w_dff_A_wZD9eGAg9_0),.din(w_dff_A_1haxGdVJ2_0),.clk(gclk));
	jdff dff_A_wZD9eGAg9_0(.dout(w_dff_A_Kvt6v9Sw6_0),.din(w_dff_A_wZD9eGAg9_0),.clk(gclk));
	jdff dff_A_Kvt6v9Sw6_0(.dout(w_dff_A_6Glt6atn6_0),.din(w_dff_A_Kvt6v9Sw6_0),.clk(gclk));
	jdff dff_A_6Glt6atn6_0(.dout(w_dff_A_bzvNBOYj0_0),.din(w_dff_A_6Glt6atn6_0),.clk(gclk));
	jdff dff_A_bzvNBOYj0_0(.dout(w_dff_A_6BM5FR752_0),.din(w_dff_A_bzvNBOYj0_0),.clk(gclk));
	jdff dff_A_6BM5FR752_0(.dout(G615),.din(w_dff_A_6BM5FR752_0),.clk(gclk));
	jdff dff_A_VyRNnbsR6_2(.dout(w_dff_A_8v0iwfKN0_0),.din(w_dff_A_VyRNnbsR6_2),.clk(gclk));
	jdff dff_A_8v0iwfKN0_0(.dout(w_dff_A_5c3an98c5_0),.din(w_dff_A_8v0iwfKN0_0),.clk(gclk));
	jdff dff_A_5c3an98c5_0(.dout(w_dff_A_eP0RgtWU9_0),.din(w_dff_A_5c3an98c5_0),.clk(gclk));
	jdff dff_A_eP0RgtWU9_0(.dout(w_dff_A_2lkPwFN80_0),.din(w_dff_A_eP0RgtWU9_0),.clk(gclk));
	jdff dff_A_2lkPwFN80_0(.dout(w_dff_A_ara8B4DS4_0),.din(w_dff_A_2lkPwFN80_0),.clk(gclk));
	jdff dff_A_ara8B4DS4_0(.dout(w_dff_A_JkxiWNce1_0),.din(w_dff_A_ara8B4DS4_0),.clk(gclk));
	jdff dff_A_JkxiWNce1_0(.dout(w_dff_A_yo4P0xeu7_0),.din(w_dff_A_JkxiWNce1_0),.clk(gclk));
	jdff dff_A_yo4P0xeu7_0(.dout(w_dff_A_5BWg8Psx7_0),.din(w_dff_A_yo4P0xeu7_0),.clk(gclk));
	jdff dff_A_5BWg8Psx7_0(.dout(w_dff_A_c08IIq7k5_0),.din(w_dff_A_5BWg8Psx7_0),.clk(gclk));
	jdff dff_A_c08IIq7k5_0(.dout(w_dff_A_vjE7kXum4_0),.din(w_dff_A_c08IIq7k5_0),.clk(gclk));
	jdff dff_A_vjE7kXum4_0(.dout(w_dff_A_OACUKO5e1_0),.din(w_dff_A_vjE7kXum4_0),.clk(gclk));
	jdff dff_A_OACUKO5e1_0(.dout(w_dff_A_EIFAbSCw3_0),.din(w_dff_A_OACUKO5e1_0),.clk(gclk));
	jdff dff_A_EIFAbSCw3_0(.dout(w_dff_A_Uns95WFP8_0),.din(w_dff_A_EIFAbSCw3_0),.clk(gclk));
	jdff dff_A_Uns95WFP8_0(.dout(w_dff_A_ywLwuiAb9_0),.din(w_dff_A_Uns95WFP8_0),.clk(gclk));
	jdff dff_A_ywLwuiAb9_0(.dout(w_dff_A_dQbOsoUn7_0),.din(w_dff_A_ywLwuiAb9_0),.clk(gclk));
	jdff dff_A_dQbOsoUn7_0(.dout(w_dff_A_y1Id65Fp3_0),.din(w_dff_A_dQbOsoUn7_0),.clk(gclk));
	jdff dff_A_y1Id65Fp3_0(.dout(w_dff_A_LwtLdMpv7_0),.din(w_dff_A_y1Id65Fp3_0),.clk(gclk));
	jdff dff_A_LwtLdMpv7_0(.dout(G626),.din(w_dff_A_LwtLdMpv7_0),.clk(gclk));
	jdff dff_A_RZ4RQ0L23_2(.dout(w_dff_A_txr7Wh484_0),.din(w_dff_A_RZ4RQ0L23_2),.clk(gclk));
	jdff dff_A_txr7Wh484_0(.dout(w_dff_A_fn7ZApTB9_0),.din(w_dff_A_txr7Wh484_0),.clk(gclk));
	jdff dff_A_fn7ZApTB9_0(.dout(w_dff_A_iJ58sCCY4_0),.din(w_dff_A_fn7ZApTB9_0),.clk(gclk));
	jdff dff_A_iJ58sCCY4_0(.dout(w_dff_A_mWkPQRQa3_0),.din(w_dff_A_iJ58sCCY4_0),.clk(gclk));
	jdff dff_A_mWkPQRQa3_0(.dout(w_dff_A_WSB7tngo1_0),.din(w_dff_A_mWkPQRQa3_0),.clk(gclk));
	jdff dff_A_WSB7tngo1_0(.dout(w_dff_A_xgaQshQA7_0),.din(w_dff_A_WSB7tngo1_0),.clk(gclk));
	jdff dff_A_xgaQshQA7_0(.dout(w_dff_A_BVDzHZaB2_0),.din(w_dff_A_xgaQshQA7_0),.clk(gclk));
	jdff dff_A_BVDzHZaB2_0(.dout(w_dff_A_O1jl03pm7_0),.din(w_dff_A_BVDzHZaB2_0),.clk(gclk));
	jdff dff_A_O1jl03pm7_0(.dout(w_dff_A_4IB0tKDg2_0),.din(w_dff_A_O1jl03pm7_0),.clk(gclk));
	jdff dff_A_4IB0tKDg2_0(.dout(w_dff_A_iGAv61P90_0),.din(w_dff_A_4IB0tKDg2_0),.clk(gclk));
	jdff dff_A_iGAv61P90_0(.dout(w_dff_A_y24CL9Za1_0),.din(w_dff_A_iGAv61P90_0),.clk(gclk));
	jdff dff_A_y24CL9Za1_0(.dout(w_dff_A_kZduCUAf2_0),.din(w_dff_A_y24CL9Za1_0),.clk(gclk));
	jdff dff_A_kZduCUAf2_0(.dout(w_dff_A_JTr66KAw8_0),.din(w_dff_A_kZduCUAf2_0),.clk(gclk));
	jdff dff_A_JTr66KAw8_0(.dout(w_dff_A_K6d8Q3cU9_0),.din(w_dff_A_JTr66KAw8_0),.clk(gclk));
	jdff dff_A_K6d8Q3cU9_0(.dout(w_dff_A_yoJGiT3X1_0),.din(w_dff_A_K6d8Q3cU9_0),.clk(gclk));
	jdff dff_A_yoJGiT3X1_0(.dout(w_dff_A_BlRKl12i8_0),.din(w_dff_A_yoJGiT3X1_0),.clk(gclk));
	jdff dff_A_BlRKl12i8_0(.dout(G632),.din(w_dff_A_BlRKl12i8_0),.clk(gclk));
	jdff dff_A_lYUtd87F9_1(.dout(w_dff_A_bwbB4dfk5_0),.din(w_dff_A_lYUtd87F9_1),.clk(gclk));
	jdff dff_A_bwbB4dfk5_0(.dout(w_dff_A_8gTHU8iS2_0),.din(w_dff_A_bwbB4dfk5_0),.clk(gclk));
	jdff dff_A_8gTHU8iS2_0(.dout(w_dff_A_BvnYNZOB3_0),.din(w_dff_A_8gTHU8iS2_0),.clk(gclk));
	jdff dff_A_BvnYNZOB3_0(.dout(w_dff_A_QyN45Ac36_0),.din(w_dff_A_BvnYNZOB3_0),.clk(gclk));
	jdff dff_A_QyN45Ac36_0(.dout(w_dff_A_BxAN3miV1_0),.din(w_dff_A_QyN45Ac36_0),.clk(gclk));
	jdff dff_A_BxAN3miV1_0(.dout(w_dff_A_Too8TLhh7_0),.din(w_dff_A_BxAN3miV1_0),.clk(gclk));
	jdff dff_A_Too8TLhh7_0(.dout(w_dff_A_jz0cGITH3_0),.din(w_dff_A_Too8TLhh7_0),.clk(gclk));
	jdff dff_A_jz0cGITH3_0(.dout(w_dff_A_w6kU9sVE5_0),.din(w_dff_A_jz0cGITH3_0),.clk(gclk));
	jdff dff_A_w6kU9sVE5_0(.dout(w_dff_A_QRrpYB9c1_0),.din(w_dff_A_w6kU9sVE5_0),.clk(gclk));
	jdff dff_A_QRrpYB9c1_0(.dout(w_dff_A_FUU9QeKu5_0),.din(w_dff_A_QRrpYB9c1_0),.clk(gclk));
	jdff dff_A_FUU9QeKu5_0(.dout(w_dff_A_TBPKl1lf1_0),.din(w_dff_A_FUU9QeKu5_0),.clk(gclk));
	jdff dff_A_TBPKl1lf1_0(.dout(w_dff_A_UYjP4O1j9_0),.din(w_dff_A_TBPKl1lf1_0),.clk(gclk));
	jdff dff_A_UYjP4O1j9_0(.dout(w_dff_A_AZEwqLtC2_0),.din(w_dff_A_UYjP4O1j9_0),.clk(gclk));
	jdff dff_A_AZEwqLtC2_0(.dout(w_dff_A_wjOrQWWf2_0),.din(w_dff_A_AZEwqLtC2_0),.clk(gclk));
	jdff dff_A_wjOrQWWf2_0(.dout(w_dff_A_rAk1AOeY4_0),.din(w_dff_A_wjOrQWWf2_0),.clk(gclk));
	jdff dff_A_rAk1AOeY4_0(.dout(w_dff_A_sV3M7dZY7_0),.din(w_dff_A_rAk1AOeY4_0),.clk(gclk));
	jdff dff_A_sV3M7dZY7_0(.dout(w_dff_A_mQ3bit1g5_0),.din(w_dff_A_sV3M7dZY7_0),.clk(gclk));
	jdff dff_A_mQ3bit1g5_0(.dout(w_dff_A_KcNSmz6o9_0),.din(w_dff_A_mQ3bit1g5_0),.clk(gclk));
	jdff dff_A_KcNSmz6o9_0(.dout(w_dff_A_hOU7wK100_0),.din(w_dff_A_KcNSmz6o9_0),.clk(gclk));
	jdff dff_A_hOU7wK100_0(.dout(w_dff_A_aHLi1u3A8_0),.din(w_dff_A_hOU7wK100_0),.clk(gclk));
	jdff dff_A_aHLi1u3A8_0(.dout(w_dff_A_DGGQpU6e9_0),.din(w_dff_A_aHLi1u3A8_0),.clk(gclk));
	jdff dff_A_DGGQpU6e9_0(.dout(w_dff_A_GVvo75fl8_0),.din(w_dff_A_DGGQpU6e9_0),.clk(gclk));
	jdff dff_A_GVvo75fl8_0(.dout(G1002),.din(w_dff_A_GVvo75fl8_0),.clk(gclk));
	jdff dff_A_tW43U9KN1_1(.dout(w_dff_A_7s0FSjaT0_0),.din(w_dff_A_tW43U9KN1_1),.clk(gclk));
	jdff dff_A_7s0FSjaT0_0(.dout(w_dff_A_NBBiu6xp2_0),.din(w_dff_A_7s0FSjaT0_0),.clk(gclk));
	jdff dff_A_NBBiu6xp2_0(.dout(w_dff_A_moFeEk9L8_0),.din(w_dff_A_NBBiu6xp2_0),.clk(gclk));
	jdff dff_A_moFeEk9L8_0(.dout(w_dff_A_u35H4Nyf2_0),.din(w_dff_A_moFeEk9L8_0),.clk(gclk));
	jdff dff_A_u35H4Nyf2_0(.dout(w_dff_A_XBD0ESze7_0),.din(w_dff_A_u35H4Nyf2_0),.clk(gclk));
	jdff dff_A_XBD0ESze7_0(.dout(w_dff_A_6PKRrom93_0),.din(w_dff_A_XBD0ESze7_0),.clk(gclk));
	jdff dff_A_6PKRrom93_0(.dout(w_dff_A_jHLZZbYD8_0),.din(w_dff_A_6PKRrom93_0),.clk(gclk));
	jdff dff_A_jHLZZbYD8_0(.dout(w_dff_A_3SyNmhWU4_0),.din(w_dff_A_jHLZZbYD8_0),.clk(gclk));
	jdff dff_A_3SyNmhWU4_0(.dout(w_dff_A_w04x8hvn5_0),.din(w_dff_A_3SyNmhWU4_0),.clk(gclk));
	jdff dff_A_w04x8hvn5_0(.dout(w_dff_A_rQy1K00S9_0),.din(w_dff_A_w04x8hvn5_0),.clk(gclk));
	jdff dff_A_rQy1K00S9_0(.dout(w_dff_A_FTsbSBtP3_0),.din(w_dff_A_rQy1K00S9_0),.clk(gclk));
	jdff dff_A_FTsbSBtP3_0(.dout(w_dff_A_NVQh7i3k5_0),.din(w_dff_A_FTsbSBtP3_0),.clk(gclk));
	jdff dff_A_NVQh7i3k5_0(.dout(w_dff_A_GQzo0G338_0),.din(w_dff_A_NVQh7i3k5_0),.clk(gclk));
	jdff dff_A_GQzo0G338_0(.dout(w_dff_A_fvr5Y7cP2_0),.din(w_dff_A_GQzo0G338_0),.clk(gclk));
	jdff dff_A_fvr5Y7cP2_0(.dout(w_dff_A_rASdqLYY9_0),.din(w_dff_A_fvr5Y7cP2_0),.clk(gclk));
	jdff dff_A_rASdqLYY9_0(.dout(w_dff_A_ZOroC7IB1_0),.din(w_dff_A_rASdqLYY9_0),.clk(gclk));
	jdff dff_A_ZOroC7IB1_0(.dout(w_dff_A_A3B0aA2U6_0),.din(w_dff_A_ZOroC7IB1_0),.clk(gclk));
	jdff dff_A_A3B0aA2U6_0(.dout(w_dff_A_Oo3iQI7s2_0),.din(w_dff_A_A3B0aA2U6_0),.clk(gclk));
	jdff dff_A_Oo3iQI7s2_0(.dout(w_dff_A_vnD58Lnw5_0),.din(w_dff_A_Oo3iQI7s2_0),.clk(gclk));
	jdff dff_A_vnD58Lnw5_0(.dout(w_dff_A_3eEVLCv52_0),.din(w_dff_A_vnD58Lnw5_0),.clk(gclk));
	jdff dff_A_3eEVLCv52_0(.dout(w_dff_A_x4WjN8389_0),.din(w_dff_A_3eEVLCv52_0),.clk(gclk));
	jdff dff_A_x4WjN8389_0(.dout(w_dff_A_DAIpVBCT2_0),.din(w_dff_A_x4WjN8389_0),.clk(gclk));
	jdff dff_A_DAIpVBCT2_0(.dout(G1004),.din(w_dff_A_DAIpVBCT2_0),.clk(gclk));
	jdff dff_A_vKR5DkTS6_2(.dout(w_dff_A_l2Yh8SJN9_0),.din(w_dff_A_vKR5DkTS6_2),.clk(gclk));
	jdff dff_A_l2Yh8SJN9_0(.dout(w_dff_A_hZpNyaxf5_0),.din(w_dff_A_l2Yh8SJN9_0),.clk(gclk));
	jdff dff_A_hZpNyaxf5_0(.dout(w_dff_A_q48AADeD4_0),.din(w_dff_A_hZpNyaxf5_0),.clk(gclk));
	jdff dff_A_q48AADeD4_0(.dout(w_dff_A_KZ6E29cY1_0),.din(w_dff_A_q48AADeD4_0),.clk(gclk));
	jdff dff_A_KZ6E29cY1_0(.dout(w_dff_A_agM5eRlM2_0),.din(w_dff_A_KZ6E29cY1_0),.clk(gclk));
	jdff dff_A_agM5eRlM2_0(.dout(w_dff_A_GTUDroBe6_0),.din(w_dff_A_agM5eRlM2_0),.clk(gclk));
	jdff dff_A_GTUDroBe6_0(.dout(w_dff_A_74FdOBZp5_0),.din(w_dff_A_GTUDroBe6_0),.clk(gclk));
	jdff dff_A_74FdOBZp5_0(.dout(w_dff_A_KQ0wm0q25_0),.din(w_dff_A_74FdOBZp5_0),.clk(gclk));
	jdff dff_A_KQ0wm0q25_0(.dout(w_dff_A_imkArTzf6_0),.din(w_dff_A_KQ0wm0q25_0),.clk(gclk));
	jdff dff_A_imkArTzf6_0(.dout(w_dff_A_ylvXNnnE9_0),.din(w_dff_A_imkArTzf6_0),.clk(gclk));
	jdff dff_A_ylvXNnnE9_0(.dout(w_dff_A_T0qagvLT7_0),.din(w_dff_A_ylvXNnnE9_0),.clk(gclk));
	jdff dff_A_T0qagvLT7_0(.dout(w_dff_A_MFYl9Z271_0),.din(w_dff_A_T0qagvLT7_0),.clk(gclk));
	jdff dff_A_MFYl9Z271_0(.dout(w_dff_A_vaK6s1wt0_0),.din(w_dff_A_MFYl9Z271_0),.clk(gclk));
	jdff dff_A_vaK6s1wt0_0(.dout(G591),.din(w_dff_A_vaK6s1wt0_0),.clk(gclk));
	jdff dff_A_XZnSM4Bv2_2(.dout(w_dff_A_oGdPn1nK8_0),.din(w_dff_A_XZnSM4Bv2_2),.clk(gclk));
	jdff dff_A_oGdPn1nK8_0(.dout(w_dff_A_5Ce3RTXV1_0),.din(w_dff_A_oGdPn1nK8_0),.clk(gclk));
	jdff dff_A_5Ce3RTXV1_0(.dout(w_dff_A_lA1EDnP07_0),.din(w_dff_A_5Ce3RTXV1_0),.clk(gclk));
	jdff dff_A_lA1EDnP07_0(.dout(w_dff_A_PV3IfrPl2_0),.din(w_dff_A_lA1EDnP07_0),.clk(gclk));
	jdff dff_A_PV3IfrPl2_0(.dout(w_dff_A_f1PNTAgp5_0),.din(w_dff_A_PV3IfrPl2_0),.clk(gclk));
	jdff dff_A_f1PNTAgp5_0(.dout(w_dff_A_wHyvzA8D8_0),.din(w_dff_A_f1PNTAgp5_0),.clk(gclk));
	jdff dff_A_wHyvzA8D8_0(.dout(w_dff_A_lo68ThQf3_0),.din(w_dff_A_wHyvzA8D8_0),.clk(gclk));
	jdff dff_A_lo68ThQf3_0(.dout(w_dff_A_ZTqyAL0G6_0),.din(w_dff_A_lo68ThQf3_0),.clk(gclk));
	jdff dff_A_ZTqyAL0G6_0(.dout(w_dff_A_2S9IQ4Vn5_0),.din(w_dff_A_ZTqyAL0G6_0),.clk(gclk));
	jdff dff_A_2S9IQ4Vn5_0(.dout(w_dff_A_2tJdZ4Iw1_0),.din(w_dff_A_2S9IQ4Vn5_0),.clk(gclk));
	jdff dff_A_2tJdZ4Iw1_0(.dout(w_dff_A_3Svn1WWl9_0),.din(w_dff_A_2tJdZ4Iw1_0),.clk(gclk));
	jdff dff_A_3Svn1WWl9_0(.dout(w_dff_A_SgNjeYdC0_0),.din(w_dff_A_3Svn1WWl9_0),.clk(gclk));
	jdff dff_A_SgNjeYdC0_0(.dout(w_dff_A_GqrtkXJw6_0),.din(w_dff_A_SgNjeYdC0_0),.clk(gclk));
	jdff dff_A_GqrtkXJw6_0(.dout(w_dff_A_BxyG4Isx5_0),.din(w_dff_A_GqrtkXJw6_0),.clk(gclk));
	jdff dff_A_BxyG4Isx5_0(.dout(G618),.din(w_dff_A_BxyG4Isx5_0),.clk(gclk));
	jdff dff_A_B0akqYdF7_2(.dout(w_dff_A_qvv5I8vh5_0),.din(w_dff_A_B0akqYdF7_2),.clk(gclk));
	jdff dff_A_qvv5I8vh5_0(.dout(w_dff_A_Rt79gU1P5_0),.din(w_dff_A_qvv5I8vh5_0),.clk(gclk));
	jdff dff_A_Rt79gU1P5_0(.dout(w_dff_A_U7OSUIat9_0),.din(w_dff_A_Rt79gU1P5_0),.clk(gclk));
	jdff dff_A_U7OSUIat9_0(.dout(w_dff_A_BB1WxiYa9_0),.din(w_dff_A_U7OSUIat9_0),.clk(gclk));
	jdff dff_A_BB1WxiYa9_0(.dout(w_dff_A_Tqmo8nN45_0),.din(w_dff_A_BB1WxiYa9_0),.clk(gclk));
	jdff dff_A_Tqmo8nN45_0(.dout(w_dff_A_NrzH5RsR3_0),.din(w_dff_A_Tqmo8nN45_0),.clk(gclk));
	jdff dff_A_NrzH5RsR3_0(.dout(w_dff_A_VMqkaL9U6_0),.din(w_dff_A_NrzH5RsR3_0),.clk(gclk));
	jdff dff_A_VMqkaL9U6_0(.dout(w_dff_A_thk2pDGw4_0),.din(w_dff_A_VMqkaL9U6_0),.clk(gclk));
	jdff dff_A_thk2pDGw4_0(.dout(w_dff_A_TAC9M9JF0_0),.din(w_dff_A_thk2pDGw4_0),.clk(gclk));
	jdff dff_A_TAC9M9JF0_0(.dout(w_dff_A_iksfG1dY1_0),.din(w_dff_A_TAC9M9JF0_0),.clk(gclk));
	jdff dff_A_iksfG1dY1_0(.dout(w_dff_A_UZitD0P75_0),.din(w_dff_A_iksfG1dY1_0),.clk(gclk));
	jdff dff_A_UZitD0P75_0(.dout(w_dff_A_tjDiisG77_0),.din(w_dff_A_UZitD0P75_0),.clk(gclk));
	jdff dff_A_tjDiisG77_0(.dout(w_dff_A_PCsd5L9P9_0),.din(w_dff_A_tjDiisG77_0),.clk(gclk));
	jdff dff_A_PCsd5L9P9_0(.dout(G621),.din(w_dff_A_PCsd5L9P9_0),.clk(gclk));
	jdff dff_A_Znsu090U2_2(.dout(w_dff_A_HUDI3Dhr7_0),.din(w_dff_A_Znsu090U2_2),.clk(gclk));
	jdff dff_A_HUDI3Dhr7_0(.dout(w_dff_A_QhGHobqZ0_0),.din(w_dff_A_HUDI3Dhr7_0),.clk(gclk));
	jdff dff_A_QhGHobqZ0_0(.dout(w_dff_A_c3eQQTJu4_0),.din(w_dff_A_QhGHobqZ0_0),.clk(gclk));
	jdff dff_A_c3eQQTJu4_0(.dout(w_dff_A_hz8SHt0D4_0),.din(w_dff_A_c3eQQTJu4_0),.clk(gclk));
	jdff dff_A_hz8SHt0D4_0(.dout(w_dff_A_sh5jV3hW6_0),.din(w_dff_A_hz8SHt0D4_0),.clk(gclk));
	jdff dff_A_sh5jV3hW6_0(.dout(w_dff_A_1XTfuPD71_0),.din(w_dff_A_sh5jV3hW6_0),.clk(gclk));
	jdff dff_A_1XTfuPD71_0(.dout(w_dff_A_hBPpjwvc4_0),.din(w_dff_A_1XTfuPD71_0),.clk(gclk));
	jdff dff_A_hBPpjwvc4_0(.dout(w_dff_A_TfHZUdBq6_0),.din(w_dff_A_hBPpjwvc4_0),.clk(gclk));
	jdff dff_A_TfHZUdBq6_0(.dout(w_dff_A_wHMlGAhe1_0),.din(w_dff_A_TfHZUdBq6_0),.clk(gclk));
	jdff dff_A_wHMlGAhe1_0(.dout(w_dff_A_Gf2jRHr16_0),.din(w_dff_A_wHMlGAhe1_0),.clk(gclk));
	jdff dff_A_Gf2jRHr16_0(.dout(w_dff_A_sqN5JeLQ7_0),.din(w_dff_A_Gf2jRHr16_0),.clk(gclk));
	jdff dff_A_sqN5JeLQ7_0(.dout(w_dff_A_hxVwygIH9_0),.din(w_dff_A_sqN5JeLQ7_0),.clk(gclk));
	jdff dff_A_hxVwygIH9_0(.dout(w_dff_A_JDnLuERo5_0),.din(w_dff_A_hxVwygIH9_0),.clk(gclk));
	jdff dff_A_JDnLuERo5_0(.dout(w_dff_A_QHnbNUT07_0),.din(w_dff_A_JDnLuERo5_0),.clk(gclk));
	jdff dff_A_QHnbNUT07_0(.dout(G629),.din(w_dff_A_QHnbNUT07_0),.clk(gclk));
	jdff dff_A_hgFfuhYA3_1(.dout(w_dff_A_wAgdn2DK8_0),.din(w_dff_A_hgFfuhYA3_1),.clk(gclk));
	jdff dff_A_wAgdn2DK8_0(.dout(w_dff_A_8EZQGkaj3_0),.din(w_dff_A_wAgdn2DK8_0),.clk(gclk));
	jdff dff_A_8EZQGkaj3_0(.dout(w_dff_A_6HeZkhuj6_0),.din(w_dff_A_8EZQGkaj3_0),.clk(gclk));
	jdff dff_A_6HeZkhuj6_0(.dout(w_dff_A_UWlpq2183_0),.din(w_dff_A_6HeZkhuj6_0),.clk(gclk));
	jdff dff_A_UWlpq2183_0(.dout(w_dff_A_njN7BIqv7_0),.din(w_dff_A_UWlpq2183_0),.clk(gclk));
	jdff dff_A_njN7BIqv7_0(.dout(w_dff_A_3KS7syv66_0),.din(w_dff_A_njN7BIqv7_0),.clk(gclk));
	jdff dff_A_3KS7syv66_0(.dout(w_dff_A_5o9JObNK3_0),.din(w_dff_A_3KS7syv66_0),.clk(gclk));
	jdff dff_A_5o9JObNK3_0(.dout(w_dff_A_6TMyAyPJ9_0),.din(w_dff_A_5o9JObNK3_0),.clk(gclk));
	jdff dff_A_6TMyAyPJ9_0(.dout(w_dff_A_Q196gJ983_0),.din(w_dff_A_6TMyAyPJ9_0),.clk(gclk));
	jdff dff_A_Q196gJ983_0(.dout(w_dff_A_YX4Gu2rD1_0),.din(w_dff_A_Q196gJ983_0),.clk(gclk));
	jdff dff_A_YX4Gu2rD1_0(.dout(w_dff_A_o7Y8otNz4_0),.din(w_dff_A_YX4Gu2rD1_0),.clk(gclk));
	jdff dff_A_o7Y8otNz4_0(.dout(w_dff_A_J3fltsUP7_0),.din(w_dff_A_o7Y8otNz4_0),.clk(gclk));
	jdff dff_A_J3fltsUP7_0(.dout(w_dff_A_XjWylWI51_0),.din(w_dff_A_J3fltsUP7_0),.clk(gclk));
	jdff dff_A_XjWylWI51_0(.dout(w_dff_A_rGc7iKsR2_0),.din(w_dff_A_XjWylWI51_0),.clk(gclk));
	jdff dff_A_rGc7iKsR2_0(.dout(w_dff_A_Wd7ai7VE9_0),.din(w_dff_A_rGc7iKsR2_0),.clk(gclk));
	jdff dff_A_Wd7ai7VE9_0(.dout(w_dff_A_0H6mhUGq6_0),.din(w_dff_A_Wd7ai7VE9_0),.clk(gclk));
	jdff dff_A_0H6mhUGq6_0(.dout(w_dff_A_8TAhpgxJ2_0),.din(w_dff_A_0H6mhUGq6_0),.clk(gclk));
	jdff dff_A_8TAhpgxJ2_0(.dout(w_dff_A_FwMUFPoV6_0),.din(w_dff_A_8TAhpgxJ2_0),.clk(gclk));
	jdff dff_A_FwMUFPoV6_0(.dout(w_dff_A_kKS3FP4J0_0),.din(w_dff_A_FwMUFPoV6_0),.clk(gclk));
	jdff dff_A_kKS3FP4J0_0(.dout(G822),.din(w_dff_A_kKS3FP4J0_0),.clk(gclk));
	jdff dff_A_9ExCEcXI6_1(.dout(w_dff_A_eULcMGbE2_0),.din(w_dff_A_9ExCEcXI6_1),.clk(gclk));
	jdff dff_A_eULcMGbE2_0(.dout(w_dff_A_5WNC0i9U5_0),.din(w_dff_A_eULcMGbE2_0),.clk(gclk));
	jdff dff_A_5WNC0i9U5_0(.dout(w_dff_A_LOuHhHfj4_0),.din(w_dff_A_5WNC0i9U5_0),.clk(gclk));
	jdff dff_A_LOuHhHfj4_0(.dout(w_dff_A_AOIUlj3i0_0),.din(w_dff_A_LOuHhHfj4_0),.clk(gclk));
	jdff dff_A_AOIUlj3i0_0(.dout(w_dff_A_wxpy3BVI8_0),.din(w_dff_A_AOIUlj3i0_0),.clk(gclk));
	jdff dff_A_wxpy3BVI8_0(.dout(w_dff_A_pdWw09zv8_0),.din(w_dff_A_wxpy3BVI8_0),.clk(gclk));
	jdff dff_A_pdWw09zv8_0(.dout(w_dff_A_KQP8SEZB1_0),.din(w_dff_A_pdWw09zv8_0),.clk(gclk));
	jdff dff_A_KQP8SEZB1_0(.dout(w_dff_A_7CfHCbMw1_0),.din(w_dff_A_KQP8SEZB1_0),.clk(gclk));
	jdff dff_A_7CfHCbMw1_0(.dout(w_dff_A_tDp8novG2_0),.din(w_dff_A_7CfHCbMw1_0),.clk(gclk));
	jdff dff_A_tDp8novG2_0(.dout(w_dff_A_rwGFPfjV1_0),.din(w_dff_A_tDp8novG2_0),.clk(gclk));
	jdff dff_A_rwGFPfjV1_0(.dout(w_dff_A_CPYOVB9c5_0),.din(w_dff_A_rwGFPfjV1_0),.clk(gclk));
	jdff dff_A_CPYOVB9c5_0(.dout(w_dff_A_QEwFEsPo3_0),.din(w_dff_A_CPYOVB9c5_0),.clk(gclk));
	jdff dff_A_QEwFEsPo3_0(.dout(w_dff_A_KQ3X0ZOR6_0),.din(w_dff_A_QEwFEsPo3_0),.clk(gclk));
	jdff dff_A_KQ3X0ZOR6_0(.dout(w_dff_A_dv6LnonX7_0),.din(w_dff_A_KQ3X0ZOR6_0),.clk(gclk));
	jdff dff_A_dv6LnonX7_0(.dout(G838),.din(w_dff_A_dv6LnonX7_0),.clk(gclk));
	jdff dff_A_an0UBJ8I1_1(.dout(w_dff_A_gUBJuViZ4_0),.din(w_dff_A_an0UBJ8I1_1),.clk(gclk));
	jdff dff_A_gUBJuViZ4_0(.dout(w_dff_A_EG4FM7dn2_0),.din(w_dff_A_gUBJuViZ4_0),.clk(gclk));
	jdff dff_A_EG4FM7dn2_0(.dout(w_dff_A_hqKisNM08_0),.din(w_dff_A_EG4FM7dn2_0),.clk(gclk));
	jdff dff_A_hqKisNM08_0(.dout(w_dff_A_7m5xpbTN7_0),.din(w_dff_A_hqKisNM08_0),.clk(gclk));
	jdff dff_A_7m5xpbTN7_0(.dout(w_dff_A_jufIAScu7_0),.din(w_dff_A_7m5xpbTN7_0),.clk(gclk));
	jdff dff_A_jufIAScu7_0(.dout(w_dff_A_pAAohuZF1_0),.din(w_dff_A_jufIAScu7_0),.clk(gclk));
	jdff dff_A_pAAohuZF1_0(.dout(w_dff_A_JzpEgPu87_0),.din(w_dff_A_pAAohuZF1_0),.clk(gclk));
	jdff dff_A_JzpEgPu87_0(.dout(w_dff_A_TKvq1jPF5_0),.din(w_dff_A_JzpEgPu87_0),.clk(gclk));
	jdff dff_A_TKvq1jPF5_0(.dout(w_dff_A_CX8VlSlG2_0),.din(w_dff_A_TKvq1jPF5_0),.clk(gclk));
	jdff dff_A_CX8VlSlG2_0(.dout(w_dff_A_0a0JOHZa0_0),.din(w_dff_A_CX8VlSlG2_0),.clk(gclk));
	jdff dff_A_0a0JOHZa0_0(.dout(w_dff_A_QL9xJwti7_0),.din(w_dff_A_0a0JOHZa0_0),.clk(gclk));
	jdff dff_A_QL9xJwti7_0(.dout(w_dff_A_kfqdzEDL3_0),.din(w_dff_A_QL9xJwti7_0),.clk(gclk));
	jdff dff_A_kfqdzEDL3_0(.dout(w_dff_A_2XRKEYz92_0),.din(w_dff_A_kfqdzEDL3_0),.clk(gclk));
	jdff dff_A_2XRKEYz92_0(.dout(w_dff_A_wSJYx65l6_0),.din(w_dff_A_2XRKEYz92_0),.clk(gclk));
	jdff dff_A_wSJYx65l6_0(.dout(w_dff_A_MVi9QUKQ4_0),.din(w_dff_A_wSJYx65l6_0),.clk(gclk));
	jdff dff_A_MVi9QUKQ4_0(.dout(w_dff_A_rbsSBUxY7_0),.din(w_dff_A_MVi9QUKQ4_0),.clk(gclk));
	jdff dff_A_rbsSBUxY7_0(.dout(w_dff_A_6hXiobxC6_0),.din(w_dff_A_rbsSBUxY7_0),.clk(gclk));
	jdff dff_A_6hXiobxC6_0(.dout(G861),.din(w_dff_A_6hXiobxC6_0),.clk(gclk));
	jdff dff_A_J3A90Aak2_1(.dout(w_dff_A_095S7ZBa5_0),.din(w_dff_A_J3A90Aak2_1),.clk(gclk));
	jdff dff_A_095S7ZBa5_0(.dout(w_dff_A_ESVnY7PM7_0),.din(w_dff_A_095S7ZBa5_0),.clk(gclk));
	jdff dff_A_ESVnY7PM7_0(.dout(w_dff_A_GOSnef3m9_0),.din(w_dff_A_ESVnY7PM7_0),.clk(gclk));
	jdff dff_A_GOSnef3m9_0(.dout(w_dff_A_Vbzm2oFo6_0),.din(w_dff_A_GOSnef3m9_0),.clk(gclk));
	jdff dff_A_Vbzm2oFo6_0(.dout(w_dff_A_xxznfzh42_0),.din(w_dff_A_Vbzm2oFo6_0),.clk(gclk));
	jdff dff_A_xxznfzh42_0(.dout(w_dff_A_oK2HLNsr3_0),.din(w_dff_A_xxznfzh42_0),.clk(gclk));
	jdff dff_A_oK2HLNsr3_0(.dout(w_dff_A_WhBfwYZv5_0),.din(w_dff_A_oK2HLNsr3_0),.clk(gclk));
	jdff dff_A_WhBfwYZv5_0(.dout(w_dff_A_rNfutp1c7_0),.din(w_dff_A_WhBfwYZv5_0),.clk(gclk));
	jdff dff_A_rNfutp1c7_0(.dout(w_dff_A_TatpMFv50_0),.din(w_dff_A_rNfutp1c7_0),.clk(gclk));
	jdff dff_A_TatpMFv50_0(.dout(G623),.din(w_dff_A_TatpMFv50_0),.clk(gclk));
	jdff dff_A_PsMfZTAJ4_2(.dout(w_dff_A_AZvzbllH8_0),.din(w_dff_A_PsMfZTAJ4_2),.clk(gclk));
	jdff dff_A_AZvzbllH8_0(.dout(w_dff_A_1LBFoYk27_0),.din(w_dff_A_AZvzbllH8_0),.clk(gclk));
	jdff dff_A_1LBFoYk27_0(.dout(w_dff_A_GvaxARSZ6_0),.din(w_dff_A_1LBFoYk27_0),.clk(gclk));
	jdff dff_A_GvaxARSZ6_0(.dout(w_dff_A_RGKrigig4_0),.din(w_dff_A_GvaxARSZ6_0),.clk(gclk));
	jdff dff_A_RGKrigig4_0(.dout(w_dff_A_22YHxR059_0),.din(w_dff_A_RGKrigig4_0),.clk(gclk));
	jdff dff_A_22YHxR059_0(.dout(w_dff_A_eifgiYac8_0),.din(w_dff_A_22YHxR059_0),.clk(gclk));
	jdff dff_A_eifgiYac8_0(.dout(w_dff_A_RtUT9neU7_0),.din(w_dff_A_eifgiYac8_0),.clk(gclk));
	jdff dff_A_RtUT9neU7_0(.dout(w_dff_A_oSiMinqj7_0),.din(w_dff_A_RtUT9neU7_0),.clk(gclk));
	jdff dff_A_oSiMinqj7_0(.dout(w_dff_A_iKvcm3a23_0),.din(w_dff_A_oSiMinqj7_0),.clk(gclk));
	jdff dff_A_iKvcm3a23_0(.dout(w_dff_A_nZEMvpum1_0),.din(w_dff_A_iKvcm3a23_0),.clk(gclk));
	jdff dff_A_nZEMvpum1_0(.dout(w_dff_A_IxD0SVC77_0),.din(w_dff_A_nZEMvpum1_0),.clk(gclk));
	jdff dff_A_IxD0SVC77_0(.dout(w_dff_A_HVknhIRf2_0),.din(w_dff_A_IxD0SVC77_0),.clk(gclk));
	jdff dff_A_HVknhIRf2_0(.dout(w_dff_A_9n7I7ANS1_0),.din(w_dff_A_HVknhIRf2_0),.clk(gclk));
	jdff dff_A_9n7I7ANS1_0(.dout(G722),.din(w_dff_A_9n7I7ANS1_0),.clk(gclk));
	jdff dff_A_lbSS0iQn2_1(.dout(w_dff_A_sCQVAFv34_0),.din(w_dff_A_lbSS0iQn2_1),.clk(gclk));
	jdff dff_A_sCQVAFv34_0(.dout(w_dff_A_nmGTiiY77_0),.din(w_dff_A_sCQVAFv34_0),.clk(gclk));
	jdff dff_A_nmGTiiY77_0(.dout(w_dff_A_Hq1NbPsd3_0),.din(w_dff_A_nmGTiiY77_0),.clk(gclk));
	jdff dff_A_Hq1NbPsd3_0(.dout(w_dff_A_zMQESlBm2_0),.din(w_dff_A_Hq1NbPsd3_0),.clk(gclk));
	jdff dff_A_zMQESlBm2_0(.dout(w_dff_A_gMPz0CsY7_0),.din(w_dff_A_zMQESlBm2_0),.clk(gclk));
	jdff dff_A_gMPz0CsY7_0(.dout(w_dff_A_brNZPAFR7_0),.din(w_dff_A_gMPz0CsY7_0),.clk(gclk));
	jdff dff_A_brNZPAFR7_0(.dout(w_dff_A_v6oYvakf3_0),.din(w_dff_A_brNZPAFR7_0),.clk(gclk));
	jdff dff_A_v6oYvakf3_0(.dout(w_dff_A_6i2p1qVP1_0),.din(w_dff_A_v6oYvakf3_0),.clk(gclk));
	jdff dff_A_6i2p1qVP1_0(.dout(w_dff_A_uChanSAJ6_0),.din(w_dff_A_6i2p1qVP1_0),.clk(gclk));
	jdff dff_A_uChanSAJ6_0(.dout(w_dff_A_jI2swj6e0_0),.din(w_dff_A_uChanSAJ6_0),.clk(gclk));
	jdff dff_A_jI2swj6e0_0(.dout(w_dff_A_UUzW6DcE1_0),.din(w_dff_A_jI2swj6e0_0),.clk(gclk));
	jdff dff_A_UUzW6DcE1_0(.dout(w_dff_A_3qqKZWbw7_0),.din(w_dff_A_UUzW6DcE1_0),.clk(gclk));
	jdff dff_A_3qqKZWbw7_0(.dout(G832),.din(w_dff_A_3qqKZWbw7_0),.clk(gclk));
	jdff dff_A_D28W5EYA0_1(.dout(w_dff_A_p0u4xb6B4_0),.din(w_dff_A_D28W5EYA0_1),.clk(gclk));
	jdff dff_A_p0u4xb6B4_0(.dout(w_dff_A_eFblj2Xf9_0),.din(w_dff_A_p0u4xb6B4_0),.clk(gclk));
	jdff dff_A_eFblj2Xf9_0(.dout(w_dff_A_quJ1lWA34_0),.din(w_dff_A_eFblj2Xf9_0),.clk(gclk));
	jdff dff_A_quJ1lWA34_0(.dout(w_dff_A_C1xp1yR35_0),.din(w_dff_A_quJ1lWA34_0),.clk(gclk));
	jdff dff_A_C1xp1yR35_0(.dout(w_dff_A_0Lj3NiCX0_0),.din(w_dff_A_C1xp1yR35_0),.clk(gclk));
	jdff dff_A_0Lj3NiCX0_0(.dout(w_dff_A_gTNtLMVa8_0),.din(w_dff_A_0Lj3NiCX0_0),.clk(gclk));
	jdff dff_A_gTNtLMVa8_0(.dout(w_dff_A_SiWz9tmd0_0),.din(w_dff_A_gTNtLMVa8_0),.clk(gclk));
	jdff dff_A_SiWz9tmd0_0(.dout(w_dff_A_3LcXvDW19_0),.din(w_dff_A_SiWz9tmd0_0),.clk(gclk));
	jdff dff_A_3LcXvDW19_0(.dout(w_dff_A_p4evVdpo6_0),.din(w_dff_A_3LcXvDW19_0),.clk(gclk));
	jdff dff_A_p4evVdpo6_0(.dout(w_dff_A_KTLNCtdL9_0),.din(w_dff_A_p4evVdpo6_0),.clk(gclk));
	jdff dff_A_KTLNCtdL9_0(.dout(w_dff_A_zOelNpH78_0),.din(w_dff_A_KTLNCtdL9_0),.clk(gclk));
	jdff dff_A_zOelNpH78_0(.dout(w_dff_A_NzvvGosU3_0),.din(w_dff_A_zOelNpH78_0),.clk(gclk));
	jdff dff_A_NzvvGosU3_0(.dout(w_dff_A_DKQ6jBI75_0),.din(w_dff_A_NzvvGosU3_0),.clk(gclk));
	jdff dff_A_DKQ6jBI75_0(.dout(G834),.din(w_dff_A_DKQ6jBI75_0),.clk(gclk));
	jdff dff_A_4PavxOpF1_1(.dout(w_dff_A_Qv8LXOZe8_0),.din(w_dff_A_4PavxOpF1_1),.clk(gclk));
	jdff dff_A_Qv8LXOZe8_0(.dout(w_dff_A_I4BcIiKF5_0),.din(w_dff_A_Qv8LXOZe8_0),.clk(gclk));
	jdff dff_A_I4BcIiKF5_0(.dout(w_dff_A_HR1U3KUx8_0),.din(w_dff_A_I4BcIiKF5_0),.clk(gclk));
	jdff dff_A_HR1U3KUx8_0(.dout(w_dff_A_anHhA3nr4_0),.din(w_dff_A_HR1U3KUx8_0),.clk(gclk));
	jdff dff_A_anHhA3nr4_0(.dout(w_dff_A_9Aen7PEI7_0),.din(w_dff_A_anHhA3nr4_0),.clk(gclk));
	jdff dff_A_9Aen7PEI7_0(.dout(w_dff_A_J0I4b43A6_0),.din(w_dff_A_9Aen7PEI7_0),.clk(gclk));
	jdff dff_A_J0I4b43A6_0(.dout(w_dff_A_uZTXq8lc1_0),.din(w_dff_A_J0I4b43A6_0),.clk(gclk));
	jdff dff_A_uZTXq8lc1_0(.dout(w_dff_A_iIueJcY23_0),.din(w_dff_A_uZTXq8lc1_0),.clk(gclk));
	jdff dff_A_iIueJcY23_0(.dout(w_dff_A_GoJv94Cg9_0),.din(w_dff_A_iIueJcY23_0),.clk(gclk));
	jdff dff_A_GoJv94Cg9_0(.dout(w_dff_A_TVBGNKJm3_0),.din(w_dff_A_GoJv94Cg9_0),.clk(gclk));
	jdff dff_A_TVBGNKJm3_0(.dout(w_dff_A_z73FdqE16_0),.din(w_dff_A_TVBGNKJm3_0),.clk(gclk));
	jdff dff_A_z73FdqE16_0(.dout(w_dff_A_WbPvDGwR3_0),.din(w_dff_A_z73FdqE16_0),.clk(gclk));
	jdff dff_A_WbPvDGwR3_0(.dout(w_dff_A_7j605oDE4_0),.din(w_dff_A_WbPvDGwR3_0),.clk(gclk));
	jdff dff_A_7j605oDE4_0(.dout(w_dff_A_gfl235sD6_0),.din(w_dff_A_7j605oDE4_0),.clk(gclk));
	jdff dff_A_gfl235sD6_0(.dout(w_dff_A_XbWshpzL5_0),.din(w_dff_A_gfl235sD6_0),.clk(gclk));
	jdff dff_A_XbWshpzL5_0(.dout(G836),.din(w_dff_A_XbWshpzL5_0),.clk(gclk));
	jdff dff_A_uCgvuOjA0_2(.dout(w_dff_A_v0jJKr6S3_0),.din(w_dff_A_uCgvuOjA0_2),.clk(gclk));
	jdff dff_A_v0jJKr6S3_0(.dout(w_dff_A_XrzYRPur9_0),.din(w_dff_A_v0jJKr6S3_0),.clk(gclk));
	jdff dff_A_XrzYRPur9_0(.dout(w_dff_A_wlbXbTYG4_0),.din(w_dff_A_XrzYRPur9_0),.clk(gclk));
	jdff dff_A_wlbXbTYG4_0(.dout(w_dff_A_62uB0t0e8_0),.din(w_dff_A_wlbXbTYG4_0),.clk(gclk));
	jdff dff_A_62uB0t0e8_0(.dout(w_dff_A_CwDC2akM7_0),.din(w_dff_A_62uB0t0e8_0),.clk(gclk));
	jdff dff_A_CwDC2akM7_0(.dout(w_dff_A_tloivukf8_0),.din(w_dff_A_CwDC2akM7_0),.clk(gclk));
	jdff dff_A_tloivukf8_0(.dout(w_dff_A_wPEG65Sn7_0),.din(w_dff_A_tloivukf8_0),.clk(gclk));
	jdff dff_A_wPEG65Sn7_0(.dout(w_dff_A_W9HPife25_0),.din(w_dff_A_wPEG65Sn7_0),.clk(gclk));
	jdff dff_A_W9HPife25_0(.dout(w_dff_A_1ewGm17r1_0),.din(w_dff_A_W9HPife25_0),.clk(gclk));
	jdff dff_A_1ewGm17r1_0(.dout(w_dff_A_hPvTzWf08_0),.din(w_dff_A_1ewGm17r1_0),.clk(gclk));
	jdff dff_A_hPvTzWf08_0(.dout(w_dff_A_8HJp41DM4_0),.din(w_dff_A_hPvTzWf08_0),.clk(gclk));
	jdff dff_A_8HJp41DM4_0(.dout(w_dff_A_xMM7kB9L9_0),.din(w_dff_A_8HJp41DM4_0),.clk(gclk));
	jdff dff_A_xMM7kB9L9_0(.dout(w_dff_A_SkCjaWIe4_0),.din(w_dff_A_xMM7kB9L9_0),.clk(gclk));
	jdff dff_A_SkCjaWIe4_0(.dout(G859),.din(w_dff_A_SkCjaWIe4_0),.clk(gclk));
	jdff dff_A_PwVeE3Jp6_1(.dout(w_dff_A_vvDe9zXd5_0),.din(w_dff_A_PwVeE3Jp6_1),.clk(gclk));
	jdff dff_A_vvDe9zXd5_0(.dout(w_dff_A_D7X7ut397_0),.din(w_dff_A_vvDe9zXd5_0),.clk(gclk));
	jdff dff_A_D7X7ut397_0(.dout(w_dff_A_l8GjwcZV4_0),.din(w_dff_A_D7X7ut397_0),.clk(gclk));
	jdff dff_A_l8GjwcZV4_0(.dout(w_dff_A_3rMJ9UZe3_0),.din(w_dff_A_l8GjwcZV4_0),.clk(gclk));
	jdff dff_A_3rMJ9UZe3_0(.dout(w_dff_A_xgoXUh0e2_0),.din(w_dff_A_3rMJ9UZe3_0),.clk(gclk));
	jdff dff_A_xgoXUh0e2_0(.dout(w_dff_A_7o2950PG1_0),.din(w_dff_A_xgoXUh0e2_0),.clk(gclk));
	jdff dff_A_7o2950PG1_0(.dout(w_dff_A_GQn8F1U73_0),.din(w_dff_A_7o2950PG1_0),.clk(gclk));
	jdff dff_A_GQn8F1U73_0(.dout(w_dff_A_h8qWiK589_0),.din(w_dff_A_GQn8F1U73_0),.clk(gclk));
	jdff dff_A_h8qWiK589_0(.dout(w_dff_A_N75vCvc63_0),.din(w_dff_A_h8qWiK589_0),.clk(gclk));
	jdff dff_A_N75vCvc63_0(.dout(w_dff_A_rZhRhsc42_0),.din(w_dff_A_N75vCvc63_0),.clk(gclk));
	jdff dff_A_rZhRhsc42_0(.dout(w_dff_A_OidMD6HS4_0),.din(w_dff_A_rZhRhsc42_0),.clk(gclk));
	jdff dff_A_OidMD6HS4_0(.dout(w_dff_A_xk218FQj0_0),.din(w_dff_A_OidMD6HS4_0),.clk(gclk));
	jdff dff_A_xk218FQj0_0(.dout(G871),.din(w_dff_A_xk218FQj0_0),.clk(gclk));
	jdff dff_A_ORWvyfmF9_1(.dout(w_dff_A_NTttsbUL7_0),.din(w_dff_A_ORWvyfmF9_1),.clk(gclk));
	jdff dff_A_NTttsbUL7_0(.dout(w_dff_A_OyKzx4fv1_0),.din(w_dff_A_NTttsbUL7_0),.clk(gclk));
	jdff dff_A_OyKzx4fv1_0(.dout(w_dff_A_bMXasXir8_0),.din(w_dff_A_OyKzx4fv1_0),.clk(gclk));
	jdff dff_A_bMXasXir8_0(.dout(w_dff_A_2tKugoVb1_0),.din(w_dff_A_bMXasXir8_0),.clk(gclk));
	jdff dff_A_2tKugoVb1_0(.dout(w_dff_A_RcngK7Hr4_0),.din(w_dff_A_2tKugoVb1_0),.clk(gclk));
	jdff dff_A_RcngK7Hr4_0(.dout(w_dff_A_Qo4FkX5p5_0),.din(w_dff_A_RcngK7Hr4_0),.clk(gclk));
	jdff dff_A_Qo4FkX5p5_0(.dout(w_dff_A_VjyYokhV5_0),.din(w_dff_A_Qo4FkX5p5_0),.clk(gclk));
	jdff dff_A_VjyYokhV5_0(.dout(w_dff_A_52Dt3Y2q1_0),.din(w_dff_A_VjyYokhV5_0),.clk(gclk));
	jdff dff_A_52Dt3Y2q1_0(.dout(w_dff_A_Q1CVm3Fv4_0),.din(w_dff_A_52Dt3Y2q1_0),.clk(gclk));
	jdff dff_A_Q1CVm3Fv4_0(.dout(w_dff_A_O6Qpz3XO9_0),.din(w_dff_A_Q1CVm3Fv4_0),.clk(gclk));
	jdff dff_A_O6Qpz3XO9_0(.dout(w_dff_A_tPCvkRa59_0),.din(w_dff_A_O6Qpz3XO9_0),.clk(gclk));
	jdff dff_A_tPCvkRa59_0(.dout(w_dff_A_EPsyu48S8_0),.din(w_dff_A_tPCvkRa59_0),.clk(gclk));
	jdff dff_A_EPsyu48S8_0(.dout(w_dff_A_jYA1aPvp5_0),.din(w_dff_A_EPsyu48S8_0),.clk(gclk));
	jdff dff_A_jYA1aPvp5_0(.dout(w_dff_A_4MmVsxrl7_0),.din(w_dff_A_jYA1aPvp5_0),.clk(gclk));
	jdff dff_A_4MmVsxrl7_0(.dout(G873),.din(w_dff_A_4MmVsxrl7_0),.clk(gclk));
	jdff dff_A_lkGGGKZR7_1(.dout(w_dff_A_hI1Tcukw9_0),.din(w_dff_A_lkGGGKZR7_1),.clk(gclk));
	jdff dff_A_hI1Tcukw9_0(.dout(w_dff_A_iBqs50su2_0),.din(w_dff_A_hI1Tcukw9_0),.clk(gclk));
	jdff dff_A_iBqs50su2_0(.dout(w_dff_A_nX7Q4mEr4_0),.din(w_dff_A_iBqs50su2_0),.clk(gclk));
	jdff dff_A_nX7Q4mEr4_0(.dout(w_dff_A_dBjPSm9l5_0),.din(w_dff_A_nX7Q4mEr4_0),.clk(gclk));
	jdff dff_A_dBjPSm9l5_0(.dout(w_dff_A_3AnIbj842_0),.din(w_dff_A_dBjPSm9l5_0),.clk(gclk));
	jdff dff_A_3AnIbj842_0(.dout(w_dff_A_eIEMQ4sF1_0),.din(w_dff_A_3AnIbj842_0),.clk(gclk));
	jdff dff_A_eIEMQ4sF1_0(.dout(w_dff_A_qlFVpBF09_0),.din(w_dff_A_eIEMQ4sF1_0),.clk(gclk));
	jdff dff_A_qlFVpBF09_0(.dout(w_dff_A_deqvx5Zb0_0),.din(w_dff_A_qlFVpBF09_0),.clk(gclk));
	jdff dff_A_deqvx5Zb0_0(.dout(w_dff_A_MkKoFrcX8_0),.din(w_dff_A_deqvx5Zb0_0),.clk(gclk));
	jdff dff_A_MkKoFrcX8_0(.dout(w_dff_A_fio9PFVt0_0),.din(w_dff_A_MkKoFrcX8_0),.clk(gclk));
	jdff dff_A_fio9PFVt0_0(.dout(w_dff_A_iAyjbgUq2_0),.din(w_dff_A_fio9PFVt0_0),.clk(gclk));
	jdff dff_A_iAyjbgUq2_0(.dout(w_dff_A_A9GE2VRZ3_0),.din(w_dff_A_iAyjbgUq2_0),.clk(gclk));
	jdff dff_A_A9GE2VRZ3_0(.dout(w_dff_A_WVPwuZV38_0),.din(w_dff_A_A9GE2VRZ3_0),.clk(gclk));
	jdff dff_A_WVPwuZV38_0(.dout(w_dff_A_83uEDLpM4_0),.din(w_dff_A_WVPwuZV38_0),.clk(gclk));
	jdff dff_A_83uEDLpM4_0(.dout(w_dff_A_LYLIQECz2_0),.din(w_dff_A_83uEDLpM4_0),.clk(gclk));
	jdff dff_A_LYLIQECz2_0(.dout(G875),.din(w_dff_A_LYLIQECz2_0),.clk(gclk));
	jdff dff_A_y5o85UER5_1(.dout(w_dff_A_g1MK8hkL5_0),.din(w_dff_A_y5o85UER5_1),.clk(gclk));
	jdff dff_A_g1MK8hkL5_0(.dout(w_dff_A_T9WIBBTr5_0),.din(w_dff_A_g1MK8hkL5_0),.clk(gclk));
	jdff dff_A_T9WIBBTr5_0(.dout(w_dff_A_eSKIkpYy0_0),.din(w_dff_A_T9WIBBTr5_0),.clk(gclk));
	jdff dff_A_eSKIkpYy0_0(.dout(w_dff_A_moeM5zwB5_0),.din(w_dff_A_eSKIkpYy0_0),.clk(gclk));
	jdff dff_A_moeM5zwB5_0(.dout(w_dff_A_kvuU1oFX2_0),.din(w_dff_A_moeM5zwB5_0),.clk(gclk));
	jdff dff_A_kvuU1oFX2_0(.dout(w_dff_A_CFAsKBJq7_0),.din(w_dff_A_kvuU1oFX2_0),.clk(gclk));
	jdff dff_A_CFAsKBJq7_0(.dout(w_dff_A_4EIEZhWY3_0),.din(w_dff_A_CFAsKBJq7_0),.clk(gclk));
	jdff dff_A_4EIEZhWY3_0(.dout(w_dff_A_SWEKU9a34_0),.din(w_dff_A_4EIEZhWY3_0),.clk(gclk));
	jdff dff_A_SWEKU9a34_0(.dout(w_dff_A_Nhj46LBa6_0),.din(w_dff_A_SWEKU9a34_0),.clk(gclk));
	jdff dff_A_Nhj46LBa6_0(.dout(w_dff_A_7hpTfjw56_0),.din(w_dff_A_Nhj46LBa6_0),.clk(gclk));
	jdff dff_A_7hpTfjw56_0(.dout(w_dff_A_o2a6b3xQ4_0),.din(w_dff_A_7hpTfjw56_0),.clk(gclk));
	jdff dff_A_o2a6b3xQ4_0(.dout(w_dff_A_5KMMxAwb2_0),.din(w_dff_A_o2a6b3xQ4_0),.clk(gclk));
	jdff dff_A_5KMMxAwb2_0(.dout(w_dff_A_pqSbxMkD1_0),.din(w_dff_A_5KMMxAwb2_0),.clk(gclk));
	jdff dff_A_pqSbxMkD1_0(.dout(w_dff_A_eEBuOLFI7_0),.din(w_dff_A_pqSbxMkD1_0),.clk(gclk));
	jdff dff_A_eEBuOLFI7_0(.dout(w_dff_A_mR46Ugkq4_0),.din(w_dff_A_eEBuOLFI7_0),.clk(gclk));
	jdff dff_A_mR46Ugkq4_0(.dout(w_dff_A_dCiS2op41_0),.din(w_dff_A_mR46Ugkq4_0),.clk(gclk));
	jdff dff_A_dCiS2op41_0(.dout(G877),.din(w_dff_A_dCiS2op41_0),.clk(gclk));
	jdff dff_A_32pOtW9D1_1(.dout(w_dff_A_XddnKyiD5_0),.din(w_dff_A_32pOtW9D1_1),.clk(gclk));
	jdff dff_A_XddnKyiD5_0(.dout(w_dff_A_OoJRoECC9_0),.din(w_dff_A_XddnKyiD5_0),.clk(gclk));
	jdff dff_A_OoJRoECC9_0(.dout(w_dff_A_nD75eIp11_0),.din(w_dff_A_OoJRoECC9_0),.clk(gclk));
	jdff dff_A_nD75eIp11_0(.dout(w_dff_A_aFRatdU13_0),.din(w_dff_A_nD75eIp11_0),.clk(gclk));
	jdff dff_A_aFRatdU13_0(.dout(w_dff_A_lW3A9Ekv9_0),.din(w_dff_A_aFRatdU13_0),.clk(gclk));
	jdff dff_A_lW3A9Ekv9_0(.dout(w_dff_A_9695fvsc5_0),.din(w_dff_A_lW3A9Ekv9_0),.clk(gclk));
	jdff dff_A_9695fvsc5_0(.dout(w_dff_A_S3U6ijvB5_0),.din(w_dff_A_9695fvsc5_0),.clk(gclk));
	jdff dff_A_S3U6ijvB5_0(.dout(w_dff_A_f70mi43T6_0),.din(w_dff_A_S3U6ijvB5_0),.clk(gclk));
	jdff dff_A_f70mi43T6_0(.dout(w_dff_A_ESCMdPsy2_0),.din(w_dff_A_f70mi43T6_0),.clk(gclk));
	jdff dff_A_ESCMdPsy2_0(.dout(w_dff_A_ES9gYQ6i5_0),.din(w_dff_A_ESCMdPsy2_0),.clk(gclk));
	jdff dff_A_ES9gYQ6i5_0(.dout(w_dff_A_Z7PbR7z03_0),.din(w_dff_A_ES9gYQ6i5_0),.clk(gclk));
	jdff dff_A_Z7PbR7z03_0(.dout(w_dff_A_dpReoaM02_0),.din(w_dff_A_Z7PbR7z03_0),.clk(gclk));
	jdff dff_A_dpReoaM02_0(.dout(w_dff_A_onUMXk6V9_0),.din(w_dff_A_dpReoaM02_0),.clk(gclk));
	jdff dff_A_onUMXk6V9_0(.dout(w_dff_A_Tz4jAXf56_0),.din(w_dff_A_onUMXk6V9_0),.clk(gclk));
	jdff dff_A_Tz4jAXf56_0(.dout(w_dff_A_aIQslsMW3_0),.din(w_dff_A_Tz4jAXf56_0),.clk(gclk));
	jdff dff_A_aIQslsMW3_0(.dout(w_dff_A_xvWGgnOV7_0),.din(w_dff_A_aIQslsMW3_0),.clk(gclk));
	jdff dff_A_xvWGgnOV7_0(.dout(w_dff_A_cLzWTcj00_0),.din(w_dff_A_xvWGgnOV7_0),.clk(gclk));
	jdff dff_A_cLzWTcj00_0(.dout(w_dff_A_csnrMbGv0_0),.din(w_dff_A_cLzWTcj00_0),.clk(gclk));
	jdff dff_A_csnrMbGv0_0(.dout(w_dff_A_cLd5Q0cP9_0),.din(w_dff_A_csnrMbGv0_0),.clk(gclk));
	jdff dff_A_cLd5Q0cP9_0(.dout(G998),.din(w_dff_A_cLd5Q0cP9_0),.clk(gclk));
	jdff dff_A_DX0Mtc6R2_1(.dout(w_dff_A_nTfjI0cF2_0),.din(w_dff_A_DX0Mtc6R2_1),.clk(gclk));
	jdff dff_A_nTfjI0cF2_0(.dout(w_dff_A_ryLxFFBv7_0),.din(w_dff_A_nTfjI0cF2_0),.clk(gclk));
	jdff dff_A_ryLxFFBv7_0(.dout(w_dff_A_7yPlVLkp1_0),.din(w_dff_A_ryLxFFBv7_0),.clk(gclk));
	jdff dff_A_7yPlVLkp1_0(.dout(w_dff_A_ZERoUCzr9_0),.din(w_dff_A_7yPlVLkp1_0),.clk(gclk));
	jdff dff_A_ZERoUCzr9_0(.dout(w_dff_A_JWwDsi4h2_0),.din(w_dff_A_ZERoUCzr9_0),.clk(gclk));
	jdff dff_A_JWwDsi4h2_0(.dout(w_dff_A_6ZUh4y4v1_0),.din(w_dff_A_JWwDsi4h2_0),.clk(gclk));
	jdff dff_A_6ZUh4y4v1_0(.dout(w_dff_A_16vCrZbw8_0),.din(w_dff_A_6ZUh4y4v1_0),.clk(gclk));
	jdff dff_A_16vCrZbw8_0(.dout(w_dff_A_FSZwXZ276_0),.din(w_dff_A_16vCrZbw8_0),.clk(gclk));
	jdff dff_A_FSZwXZ276_0(.dout(w_dff_A_hK9kiUZD7_0),.din(w_dff_A_FSZwXZ276_0),.clk(gclk));
	jdff dff_A_hK9kiUZD7_0(.dout(w_dff_A_wW4156Sl2_0),.din(w_dff_A_hK9kiUZD7_0),.clk(gclk));
	jdff dff_A_wW4156Sl2_0(.dout(w_dff_A_6Opw3FZL5_0),.din(w_dff_A_wW4156Sl2_0),.clk(gclk));
	jdff dff_A_6Opw3FZL5_0(.dout(w_dff_A_fxiYAWL33_0),.din(w_dff_A_6Opw3FZL5_0),.clk(gclk));
	jdff dff_A_fxiYAWL33_0(.dout(w_dff_A_WklZoigz0_0),.din(w_dff_A_fxiYAWL33_0),.clk(gclk));
	jdff dff_A_WklZoigz0_0(.dout(w_dff_A_WQgKZmDb2_0),.din(w_dff_A_WklZoigz0_0),.clk(gclk));
	jdff dff_A_WQgKZmDb2_0(.dout(w_dff_A_mAjVlnfA4_0),.din(w_dff_A_WQgKZmDb2_0),.clk(gclk));
	jdff dff_A_mAjVlnfA4_0(.dout(w_dff_A_Qcn33iHW0_0),.din(w_dff_A_mAjVlnfA4_0),.clk(gclk));
	jdff dff_A_Qcn33iHW0_0(.dout(w_dff_A_6WPFaNR41_0),.din(w_dff_A_Qcn33iHW0_0),.clk(gclk));
	jdff dff_A_6WPFaNR41_0(.dout(w_dff_A_micxCBgF9_0),.din(w_dff_A_6WPFaNR41_0),.clk(gclk));
	jdff dff_A_micxCBgF9_0(.dout(G1000),.din(w_dff_A_micxCBgF9_0),.clk(gclk));
	jdff dff_A_WTTfnauU2_2(.dout(w_dff_A_qiNPFECI1_0),.din(w_dff_A_WTTfnauU2_2),.clk(gclk));
	jdff dff_A_qiNPFECI1_0(.dout(w_dff_A_wUORH9CY2_0),.din(w_dff_A_qiNPFECI1_0),.clk(gclk));
	jdff dff_A_wUORH9CY2_0(.dout(w_dff_A_N39xu8ts0_0),.din(w_dff_A_wUORH9CY2_0),.clk(gclk));
	jdff dff_A_N39xu8ts0_0(.dout(w_dff_A_mIlpv17y8_0),.din(w_dff_A_N39xu8ts0_0),.clk(gclk));
	jdff dff_A_mIlpv17y8_0(.dout(w_dff_A_qm8ipQwt3_0),.din(w_dff_A_mIlpv17y8_0),.clk(gclk));
	jdff dff_A_qm8ipQwt3_0(.dout(w_dff_A_5Wi4odPO4_0),.din(w_dff_A_qm8ipQwt3_0),.clk(gclk));
	jdff dff_A_5Wi4odPO4_0(.dout(w_dff_A_LVK68FTZ8_0),.din(w_dff_A_5Wi4odPO4_0),.clk(gclk));
	jdff dff_A_LVK68FTZ8_0(.dout(G575),.din(w_dff_A_LVK68FTZ8_0),.clk(gclk));
	jdff dff_A_RJ18dgvy4_2(.dout(w_dff_A_ickgKFvR1_0),.din(w_dff_A_RJ18dgvy4_2),.clk(gclk));
	jdff dff_A_ickgKFvR1_0(.dout(w_dff_A_01GTjzFh5_0),.din(w_dff_A_ickgKFvR1_0),.clk(gclk));
	jdff dff_A_01GTjzFh5_0(.dout(w_dff_A_pLEqq7yX9_0),.din(w_dff_A_01GTjzFh5_0),.clk(gclk));
	jdff dff_A_pLEqq7yX9_0(.dout(w_dff_A_26apLcSj0_0),.din(w_dff_A_pLEqq7yX9_0),.clk(gclk));
	jdff dff_A_26apLcSj0_0(.dout(w_dff_A_csXTs7Yw4_0),.din(w_dff_A_26apLcSj0_0),.clk(gclk));
	jdff dff_A_csXTs7Yw4_0(.dout(w_dff_A_pmWRA6JS0_0),.din(w_dff_A_csXTs7Yw4_0),.clk(gclk));
	jdff dff_A_pmWRA6JS0_0(.dout(G585),.din(w_dff_A_pmWRA6JS0_0),.clk(gclk));
	jdff dff_A_cgdxqHwN3_2(.dout(w_dff_A_aoyZcCuj3_0),.din(w_dff_A_cgdxqHwN3_2),.clk(gclk));
	jdff dff_A_aoyZcCuj3_0(.dout(w_dff_A_6ish0ona2_0),.din(w_dff_A_aoyZcCuj3_0),.clk(gclk));
	jdff dff_A_6ish0ona2_0(.dout(w_dff_A_0ZF7D4nz8_0),.din(w_dff_A_6ish0ona2_0),.clk(gclk));
	jdff dff_A_0ZF7D4nz8_0(.dout(w_dff_A_y9XzhXBi3_0),.din(w_dff_A_0ZF7D4nz8_0),.clk(gclk));
	jdff dff_A_y9XzhXBi3_0(.dout(w_dff_A_JIkxsbV44_0),.din(w_dff_A_y9XzhXBi3_0),.clk(gclk));
	jdff dff_A_JIkxsbV44_0(.dout(w_dff_A_NNzvW05A4_0),.din(w_dff_A_JIkxsbV44_0),.clk(gclk));
	jdff dff_A_NNzvW05A4_0(.dout(w_dff_A_ioNsIhzp4_0),.din(w_dff_A_NNzvW05A4_0),.clk(gclk));
	jdff dff_A_ioNsIhzp4_0(.dout(w_dff_A_pekoyJtn2_0),.din(w_dff_A_ioNsIhzp4_0),.clk(gclk));
	jdff dff_A_pekoyJtn2_0(.dout(w_dff_A_0KlY1cIq4_0),.din(w_dff_A_pekoyJtn2_0),.clk(gclk));
	jdff dff_A_0KlY1cIq4_0(.dout(w_dff_A_pSp5ibAu8_0),.din(w_dff_A_0KlY1cIq4_0),.clk(gclk));
	jdff dff_A_pSp5ibAu8_0(.dout(w_dff_A_oMrIBUE60_0),.din(w_dff_A_pSp5ibAu8_0),.clk(gclk));
	jdff dff_A_oMrIBUE60_0(.dout(G661),.din(w_dff_A_oMrIBUE60_0),.clk(gclk));
	jdff dff_A_7W4GWUDP1_2(.dout(w_dff_A_xvOKcKuY6_0),.din(w_dff_A_7W4GWUDP1_2),.clk(gclk));
	jdff dff_A_xvOKcKuY6_0(.dout(w_dff_A_8kfcHEHr0_0),.din(w_dff_A_xvOKcKuY6_0),.clk(gclk));
	jdff dff_A_8kfcHEHr0_0(.dout(w_dff_A_66JR4QGx3_0),.din(w_dff_A_8kfcHEHr0_0),.clk(gclk));
	jdff dff_A_66JR4QGx3_0(.dout(w_dff_A_qbl5jmXt5_0),.din(w_dff_A_66JR4QGx3_0),.clk(gclk));
	jdff dff_A_qbl5jmXt5_0(.dout(w_dff_A_Rjm9jPqe8_0),.din(w_dff_A_qbl5jmXt5_0),.clk(gclk));
	jdff dff_A_Rjm9jPqe8_0(.dout(w_dff_A_IdYvVSNC8_0),.din(w_dff_A_Rjm9jPqe8_0),.clk(gclk));
	jdff dff_A_IdYvVSNC8_0(.dout(w_dff_A_DzCJnUyy5_0),.din(w_dff_A_IdYvVSNC8_0),.clk(gclk));
	jdff dff_A_DzCJnUyy5_0(.dout(w_dff_A_nuMBE6R39_0),.din(w_dff_A_DzCJnUyy5_0),.clk(gclk));
	jdff dff_A_nuMBE6R39_0(.dout(w_dff_A_W8lInqRb8_0),.din(w_dff_A_nuMBE6R39_0),.clk(gclk));
	jdff dff_A_W8lInqRb8_0(.dout(w_dff_A_9U9Fyhuk2_0),.din(w_dff_A_W8lInqRb8_0),.clk(gclk));
	jdff dff_A_9U9Fyhuk2_0(.dout(w_dff_A_iBAJdm7G7_0),.din(w_dff_A_9U9Fyhuk2_0),.clk(gclk));
	jdff dff_A_iBAJdm7G7_0(.dout(G693),.din(w_dff_A_iBAJdm7G7_0),.clk(gclk));
	jdff dff_A_GBVcLEQV9_2(.dout(w_dff_A_DWhri1bT0_0),.din(w_dff_A_GBVcLEQV9_2),.clk(gclk));
	jdff dff_A_DWhri1bT0_0(.dout(w_dff_A_HHLtTfzI9_0),.din(w_dff_A_DWhri1bT0_0),.clk(gclk));
	jdff dff_A_HHLtTfzI9_0(.dout(w_dff_A_EW1wDWNf1_0),.din(w_dff_A_HHLtTfzI9_0),.clk(gclk));
	jdff dff_A_EW1wDWNf1_0(.dout(w_dff_A_ppKmVk3i2_0),.din(w_dff_A_EW1wDWNf1_0),.clk(gclk));
	jdff dff_A_ppKmVk3i2_0(.dout(w_dff_A_h1qgAggJ6_0),.din(w_dff_A_ppKmVk3i2_0),.clk(gclk));
	jdff dff_A_h1qgAggJ6_0(.dout(w_dff_A_kFWA9HyF6_0),.din(w_dff_A_h1qgAggJ6_0),.clk(gclk));
	jdff dff_A_kFWA9HyF6_0(.dout(w_dff_A_chlM9X4k7_0),.din(w_dff_A_kFWA9HyF6_0),.clk(gclk));
	jdff dff_A_chlM9X4k7_0(.dout(G747),.din(w_dff_A_chlM9X4k7_0),.clk(gclk));
	jdff dff_A_nBX0wvip1_2(.dout(w_dff_A_Y6zRAHiT2_0),.din(w_dff_A_nBX0wvip1_2),.clk(gclk));
	jdff dff_A_Y6zRAHiT2_0(.dout(w_dff_A_gsqUxdvN0_0),.din(w_dff_A_Y6zRAHiT2_0),.clk(gclk));
	jdff dff_A_gsqUxdvN0_0(.dout(w_dff_A_LN3kr5iU5_0),.din(w_dff_A_gsqUxdvN0_0),.clk(gclk));
	jdff dff_A_LN3kr5iU5_0(.dout(w_dff_A_hgH6Jr8k8_0),.din(w_dff_A_LN3kr5iU5_0),.clk(gclk));
	jdff dff_A_hgH6Jr8k8_0(.dout(w_dff_A_oa1i2zPk6_0),.din(w_dff_A_hgH6Jr8k8_0),.clk(gclk));
	jdff dff_A_oa1i2zPk6_0(.dout(w_dff_A_alPBq42p3_0),.din(w_dff_A_oa1i2zPk6_0),.clk(gclk));
	jdff dff_A_alPBq42p3_0(.dout(w_dff_A_7d2cgz226_0),.din(w_dff_A_alPBq42p3_0),.clk(gclk));
	jdff dff_A_7d2cgz226_0(.dout(w_dff_A_gvDaQNL11_0),.din(w_dff_A_7d2cgz226_0),.clk(gclk));
	jdff dff_A_gvDaQNL11_0(.dout(G752),.din(w_dff_A_gvDaQNL11_0),.clk(gclk));
	jdff dff_A_7if5Ex0z2_2(.dout(w_dff_A_AiUgCs3j2_0),.din(w_dff_A_7if5Ex0z2_2),.clk(gclk));
	jdff dff_A_AiUgCs3j2_0(.dout(w_dff_A_TwTHJyww3_0),.din(w_dff_A_AiUgCs3j2_0),.clk(gclk));
	jdff dff_A_TwTHJyww3_0(.dout(w_dff_A_IvKZmHXa9_0),.din(w_dff_A_TwTHJyww3_0),.clk(gclk));
	jdff dff_A_IvKZmHXa9_0(.dout(w_dff_A_pxTGSbKb4_0),.din(w_dff_A_IvKZmHXa9_0),.clk(gclk));
	jdff dff_A_pxTGSbKb4_0(.dout(w_dff_A_iB2f7KVS4_0),.din(w_dff_A_pxTGSbKb4_0),.clk(gclk));
	jdff dff_A_iB2f7KVS4_0(.dout(w_dff_A_Evi6oj1V5_0),.din(w_dff_A_iB2f7KVS4_0),.clk(gclk));
	jdff dff_A_Evi6oj1V5_0(.dout(w_dff_A_kB58hnys1_0),.din(w_dff_A_Evi6oj1V5_0),.clk(gclk));
	jdff dff_A_kB58hnys1_0(.dout(w_dff_A_2Rc8y7wi0_0),.din(w_dff_A_kB58hnys1_0),.clk(gclk));
	jdff dff_A_2Rc8y7wi0_0(.dout(w_dff_A_FePXc5eJ4_0),.din(w_dff_A_2Rc8y7wi0_0),.clk(gclk));
	jdff dff_A_FePXc5eJ4_0(.dout(w_dff_A_a8Qk4bxx1_0),.din(w_dff_A_FePXc5eJ4_0),.clk(gclk));
	jdff dff_A_a8Qk4bxx1_0(.dout(G757),.din(w_dff_A_a8Qk4bxx1_0),.clk(gclk));
	jdff dff_A_esKhrEUJ8_2(.dout(w_dff_A_5DTFfIwR9_0),.din(w_dff_A_esKhrEUJ8_2),.clk(gclk));
	jdff dff_A_5DTFfIwR9_0(.dout(w_dff_A_0vWcoYRv3_0),.din(w_dff_A_5DTFfIwR9_0),.clk(gclk));
	jdff dff_A_0vWcoYRv3_0(.dout(w_dff_A_TvWaKho87_0),.din(w_dff_A_0vWcoYRv3_0),.clk(gclk));
	jdff dff_A_TvWaKho87_0(.dout(w_dff_A_SGB4ZzDu8_0),.din(w_dff_A_TvWaKho87_0),.clk(gclk));
	jdff dff_A_SGB4ZzDu8_0(.dout(w_dff_A_wydLsCJt6_0),.din(w_dff_A_SGB4ZzDu8_0),.clk(gclk));
	jdff dff_A_wydLsCJt6_0(.dout(w_dff_A_qg0TwOd41_0),.din(w_dff_A_wydLsCJt6_0),.clk(gclk));
	jdff dff_A_qg0TwOd41_0(.dout(w_dff_A_titBxf2B9_0),.din(w_dff_A_qg0TwOd41_0),.clk(gclk));
	jdff dff_A_titBxf2B9_0(.dout(w_dff_A_kXSjycLt2_0),.din(w_dff_A_titBxf2B9_0),.clk(gclk));
	jdff dff_A_kXSjycLt2_0(.dout(w_dff_A_7YUUNSrQ2_0),.din(w_dff_A_kXSjycLt2_0),.clk(gclk));
	jdff dff_A_7YUUNSrQ2_0(.dout(G762),.din(w_dff_A_7YUUNSrQ2_0),.clk(gclk));
	jdff dff_A_Zo2KDTfC2_2(.dout(w_dff_A_Sz9vAu1E6_0),.din(w_dff_A_Zo2KDTfC2_2),.clk(gclk));
	jdff dff_A_Sz9vAu1E6_0(.dout(w_dff_A_3CMRcvsG8_0),.din(w_dff_A_Sz9vAu1E6_0),.clk(gclk));
	jdff dff_A_3CMRcvsG8_0(.dout(w_dff_A_guSCZ5V70_0),.din(w_dff_A_3CMRcvsG8_0),.clk(gclk));
	jdff dff_A_guSCZ5V70_0(.dout(w_dff_A_utjEpEXv7_0),.din(w_dff_A_guSCZ5V70_0),.clk(gclk));
	jdff dff_A_utjEpEXv7_0(.dout(w_dff_A_07LDldsB9_0),.din(w_dff_A_utjEpEXv7_0),.clk(gclk));
	jdff dff_A_07LDldsB9_0(.dout(w_dff_A_8AryYicP2_0),.din(w_dff_A_07LDldsB9_0),.clk(gclk));
	jdff dff_A_8AryYicP2_0(.dout(w_dff_A_5kDxmMZn0_0),.din(w_dff_A_8AryYicP2_0),.clk(gclk));
	jdff dff_A_5kDxmMZn0_0(.dout(G787),.din(w_dff_A_5kDxmMZn0_0),.clk(gclk));
	jdff dff_A_AdHQiQye7_2(.dout(w_dff_A_AhJMBAbg8_0),.din(w_dff_A_AdHQiQye7_2),.clk(gclk));
	jdff dff_A_AhJMBAbg8_0(.dout(w_dff_A_I6U6F1X47_0),.din(w_dff_A_AhJMBAbg8_0),.clk(gclk));
	jdff dff_A_I6U6F1X47_0(.dout(w_dff_A_WRvWehwM1_0),.din(w_dff_A_I6U6F1X47_0),.clk(gclk));
	jdff dff_A_WRvWehwM1_0(.dout(w_dff_A_FOVkeETD8_0),.din(w_dff_A_WRvWehwM1_0),.clk(gclk));
	jdff dff_A_FOVkeETD8_0(.dout(w_dff_A_8PdqdZtj4_0),.din(w_dff_A_FOVkeETD8_0),.clk(gclk));
	jdff dff_A_8PdqdZtj4_0(.dout(w_dff_A_LBw97b4V0_0),.din(w_dff_A_8PdqdZtj4_0),.clk(gclk));
	jdff dff_A_LBw97b4V0_0(.dout(w_dff_A_XcBEXdFK7_0),.din(w_dff_A_LBw97b4V0_0),.clk(gclk));
	jdff dff_A_XcBEXdFK7_0(.dout(w_dff_A_R7He8G2k5_0),.din(w_dff_A_XcBEXdFK7_0),.clk(gclk));
	jdff dff_A_R7He8G2k5_0(.dout(G792),.din(w_dff_A_R7He8G2k5_0),.clk(gclk));
	jdff dff_A_JuenzXYu0_2(.dout(w_dff_A_M3DLpiA72_0),.din(w_dff_A_JuenzXYu0_2),.clk(gclk));
	jdff dff_A_M3DLpiA72_0(.dout(w_dff_A_PmQtesJW5_0),.din(w_dff_A_M3DLpiA72_0),.clk(gclk));
	jdff dff_A_PmQtesJW5_0(.dout(w_dff_A_uWF7OVIf0_0),.din(w_dff_A_PmQtesJW5_0),.clk(gclk));
	jdff dff_A_uWF7OVIf0_0(.dout(w_dff_A_5orXmOyV5_0),.din(w_dff_A_uWF7OVIf0_0),.clk(gclk));
	jdff dff_A_5orXmOyV5_0(.dout(w_dff_A_IS7AgNOe9_0),.din(w_dff_A_5orXmOyV5_0),.clk(gclk));
	jdff dff_A_IS7AgNOe9_0(.dout(w_dff_A_ylGy2fok4_0),.din(w_dff_A_IS7AgNOe9_0),.clk(gclk));
	jdff dff_A_ylGy2fok4_0(.dout(w_dff_A_eq05BWI14_0),.din(w_dff_A_ylGy2fok4_0),.clk(gclk));
	jdff dff_A_eq05BWI14_0(.dout(w_dff_A_Zr4QqwU15_0),.din(w_dff_A_eq05BWI14_0),.clk(gclk));
	jdff dff_A_Zr4QqwU15_0(.dout(w_dff_A_zrmWGPMr4_0),.din(w_dff_A_Zr4QqwU15_0),.clk(gclk));
	jdff dff_A_zrmWGPMr4_0(.dout(w_dff_A_qu9L4y1s5_0),.din(w_dff_A_zrmWGPMr4_0),.clk(gclk));
	jdff dff_A_qu9L4y1s5_0(.dout(G797),.din(w_dff_A_qu9L4y1s5_0),.clk(gclk));
	jdff dff_A_Oq5Agr8v8_2(.dout(w_dff_A_zfoHNcgE4_0),.din(w_dff_A_Oq5Agr8v8_2),.clk(gclk));
	jdff dff_A_zfoHNcgE4_0(.dout(w_dff_A_LlrZNhX42_0),.din(w_dff_A_zfoHNcgE4_0),.clk(gclk));
	jdff dff_A_LlrZNhX42_0(.dout(w_dff_A_53MU5xUe5_0),.din(w_dff_A_LlrZNhX42_0),.clk(gclk));
	jdff dff_A_53MU5xUe5_0(.dout(w_dff_A_oG3gG4hH5_0),.din(w_dff_A_53MU5xUe5_0),.clk(gclk));
	jdff dff_A_oG3gG4hH5_0(.dout(w_dff_A_H6Wft9bg2_0),.din(w_dff_A_oG3gG4hH5_0),.clk(gclk));
	jdff dff_A_H6Wft9bg2_0(.dout(w_dff_A_CBOLz7UP0_0),.din(w_dff_A_H6Wft9bg2_0),.clk(gclk));
	jdff dff_A_CBOLz7UP0_0(.dout(w_dff_A_atVMBKUE6_0),.din(w_dff_A_CBOLz7UP0_0),.clk(gclk));
	jdff dff_A_atVMBKUE6_0(.dout(w_dff_A_AoKy7gAF3_0),.din(w_dff_A_atVMBKUE6_0),.clk(gclk));
	jdff dff_A_AoKy7gAF3_0(.dout(w_dff_A_QVX67lTB4_0),.din(w_dff_A_AoKy7gAF3_0),.clk(gclk));
	jdff dff_A_QVX67lTB4_0(.dout(G802),.din(w_dff_A_QVX67lTB4_0),.clk(gclk));
	jdff dff_A_oXtvQCRh0_2(.dout(w_dff_A_AFy31fML3_0),.din(w_dff_A_oXtvQCRh0_2),.clk(gclk));
	jdff dff_A_AFy31fML3_0(.dout(w_dff_A_yLTkF0KQ9_0),.din(w_dff_A_AFy31fML3_0),.clk(gclk));
	jdff dff_A_yLTkF0KQ9_0(.dout(w_dff_A_UZ72JWAY2_0),.din(w_dff_A_yLTkF0KQ9_0),.clk(gclk));
	jdff dff_A_UZ72JWAY2_0(.dout(w_dff_A_9pnHBrWs3_0),.din(w_dff_A_UZ72JWAY2_0),.clk(gclk));
	jdff dff_A_9pnHBrWs3_0(.dout(w_dff_A_zry6GCFm8_0),.din(w_dff_A_9pnHBrWs3_0),.clk(gclk));
	jdff dff_A_zry6GCFm8_0(.dout(w_dff_A_h9veY0Y49_0),.din(w_dff_A_zry6GCFm8_0),.clk(gclk));
	jdff dff_A_h9veY0Y49_0(.dout(G642),.din(w_dff_A_h9veY0Y49_0),.clk(gclk));
	jdff dff_A_kmX7ykt16_2(.dout(w_dff_A_8c1TUqnO7_0),.din(w_dff_A_kmX7ykt16_2),.clk(gclk));
	jdff dff_A_8c1TUqnO7_0(.dout(w_dff_A_eKQkdrWr5_0),.din(w_dff_A_8c1TUqnO7_0),.clk(gclk));
	jdff dff_A_eKQkdrWr5_0(.dout(w_dff_A_LYkqClVd5_0),.din(w_dff_A_eKQkdrWr5_0),.clk(gclk));
	jdff dff_A_LYkqClVd5_0(.dout(w_dff_A_5YXDiOFk2_0),.din(w_dff_A_LYkqClVd5_0),.clk(gclk));
	jdff dff_A_5YXDiOFk2_0(.dout(w_dff_A_MjXwIlmF3_0),.din(w_dff_A_5YXDiOFk2_0),.clk(gclk));
	jdff dff_A_MjXwIlmF3_0(.dout(w_dff_A_LoHZeWOW8_0),.din(w_dff_A_MjXwIlmF3_0),.clk(gclk));
	jdff dff_A_LoHZeWOW8_0(.dout(w_dff_A_yyGcsfkC2_0),.din(w_dff_A_LoHZeWOW8_0),.clk(gclk));
	jdff dff_A_yyGcsfkC2_0(.dout(w_dff_A_65IWDiCl7_0),.din(w_dff_A_yyGcsfkC2_0),.clk(gclk));
	jdff dff_A_65IWDiCl7_0(.dout(w_dff_A_cytpHSzO3_0),.din(w_dff_A_65IWDiCl7_0),.clk(gclk));
	jdff dff_A_cytpHSzO3_0(.dout(G664),.din(w_dff_A_cytpHSzO3_0),.clk(gclk));
	jdff dff_A_hZ4sVGkq1_2(.dout(w_dff_A_udKfIzWQ4_0),.din(w_dff_A_hZ4sVGkq1_2),.clk(gclk));
	jdff dff_A_udKfIzWQ4_0(.dout(w_dff_A_vejniamN9_0),.din(w_dff_A_udKfIzWQ4_0),.clk(gclk));
	jdff dff_A_vejniamN9_0(.dout(w_dff_A_neo7xxPE8_0),.din(w_dff_A_vejniamN9_0),.clk(gclk));
	jdff dff_A_neo7xxPE8_0(.dout(w_dff_A_YHclVrpf8_0),.din(w_dff_A_neo7xxPE8_0),.clk(gclk));
	jdff dff_A_YHclVrpf8_0(.dout(w_dff_A_ceJUF5kM6_0),.din(w_dff_A_YHclVrpf8_0),.clk(gclk));
	jdff dff_A_ceJUF5kM6_0(.dout(w_dff_A_bUP0NYwP1_0),.din(w_dff_A_ceJUF5kM6_0),.clk(gclk));
	jdff dff_A_bUP0NYwP1_0(.dout(w_dff_A_ucfcjsAp5_0),.din(w_dff_A_bUP0NYwP1_0),.clk(gclk));
	jdff dff_A_ucfcjsAp5_0(.dout(w_dff_A_TRamPBMB1_0),.din(w_dff_A_ucfcjsAp5_0),.clk(gclk));
	jdff dff_A_TRamPBMB1_0(.dout(w_dff_A_11QVwRVB7_0),.din(w_dff_A_TRamPBMB1_0),.clk(gclk));
	jdff dff_A_11QVwRVB7_0(.dout(G667),.din(w_dff_A_11QVwRVB7_0),.clk(gclk));
	jdff dff_A_IObyZMPk5_2(.dout(w_dff_A_4QyUmgVw0_0),.din(w_dff_A_IObyZMPk5_2),.clk(gclk));
	jdff dff_A_4QyUmgVw0_0(.dout(w_dff_A_StUcGH4c1_0),.din(w_dff_A_4QyUmgVw0_0),.clk(gclk));
	jdff dff_A_StUcGH4c1_0(.dout(w_dff_A_MSnstR2G4_0),.din(w_dff_A_StUcGH4c1_0),.clk(gclk));
	jdff dff_A_MSnstR2G4_0(.dout(w_dff_A_CWFexcX38_0),.din(w_dff_A_MSnstR2G4_0),.clk(gclk));
	jdff dff_A_CWFexcX38_0(.dout(w_dff_A_J7X7YSBc0_0),.din(w_dff_A_CWFexcX38_0),.clk(gclk));
	jdff dff_A_J7X7YSBc0_0(.dout(w_dff_A_lEPF0NfB0_0),.din(w_dff_A_J7X7YSBc0_0),.clk(gclk));
	jdff dff_A_lEPF0NfB0_0(.dout(w_dff_A_T75FYnvw5_0),.din(w_dff_A_lEPF0NfB0_0),.clk(gclk));
	jdff dff_A_T75FYnvw5_0(.dout(w_dff_A_uS2qjpmo0_0),.din(w_dff_A_T75FYnvw5_0),.clk(gclk));
	jdff dff_A_uS2qjpmo0_0(.dout(G670),.din(w_dff_A_uS2qjpmo0_0),.clk(gclk));
	jdff dff_A_GYTpg0iA4_2(.dout(w_dff_A_qr71TKgs6_0),.din(w_dff_A_GYTpg0iA4_2),.clk(gclk));
	jdff dff_A_qr71TKgs6_0(.dout(w_dff_A_fCCOpQyt7_0),.din(w_dff_A_qr71TKgs6_0),.clk(gclk));
	jdff dff_A_fCCOpQyt7_0(.dout(w_dff_A_JvJfqCJj5_0),.din(w_dff_A_fCCOpQyt7_0),.clk(gclk));
	jdff dff_A_JvJfqCJj5_0(.dout(w_dff_A_hYM606gy2_0),.din(w_dff_A_JvJfqCJj5_0),.clk(gclk));
	jdff dff_A_hYM606gy2_0(.dout(w_dff_A_jCghNv7G4_0),.din(w_dff_A_hYM606gy2_0),.clk(gclk));
	jdff dff_A_jCghNv7G4_0(.dout(G676),.din(w_dff_A_jCghNv7G4_0),.clk(gclk));
	jdff dff_A_8eEJ4Fst4_2(.dout(w_dff_A_z29pUF2q2_0),.din(w_dff_A_8eEJ4Fst4_2),.clk(gclk));
	jdff dff_A_z29pUF2q2_0(.dout(w_dff_A_ABvZrmUz6_0),.din(w_dff_A_z29pUF2q2_0),.clk(gclk));
	jdff dff_A_ABvZrmUz6_0(.dout(w_dff_A_9gxXs9RW4_0),.din(w_dff_A_ABvZrmUz6_0),.clk(gclk));
	jdff dff_A_9gxXs9RW4_0(.dout(w_dff_A_ZR5Hs4fi9_0),.din(w_dff_A_9gxXs9RW4_0),.clk(gclk));
	jdff dff_A_ZR5Hs4fi9_0(.dout(w_dff_A_VbV0U5Qh2_0),.din(w_dff_A_ZR5Hs4fi9_0),.clk(gclk));
	jdff dff_A_VbV0U5Qh2_0(.dout(w_dff_A_Otgs3z9w2_0),.din(w_dff_A_VbV0U5Qh2_0),.clk(gclk));
	jdff dff_A_Otgs3z9w2_0(.dout(w_dff_A_OjxKfTJd9_0),.din(w_dff_A_Otgs3z9w2_0),.clk(gclk));
	jdff dff_A_OjxKfTJd9_0(.dout(w_dff_A_3TeE7m7O3_0),.din(w_dff_A_OjxKfTJd9_0),.clk(gclk));
	jdff dff_A_3TeE7m7O3_0(.dout(w_dff_A_P5M5q3K66_0),.din(w_dff_A_3TeE7m7O3_0),.clk(gclk));
	jdff dff_A_P5M5q3K66_0(.dout(G696),.din(w_dff_A_P5M5q3K66_0),.clk(gclk));
	jdff dff_A_2N0KkA108_2(.dout(w_dff_A_DeXEoGm77_0),.din(w_dff_A_2N0KkA108_2),.clk(gclk));
	jdff dff_A_DeXEoGm77_0(.dout(w_dff_A_jRRsxoCY2_0),.din(w_dff_A_DeXEoGm77_0),.clk(gclk));
	jdff dff_A_jRRsxoCY2_0(.dout(w_dff_A_jMVx26Eo7_0),.din(w_dff_A_jRRsxoCY2_0),.clk(gclk));
	jdff dff_A_jMVx26Eo7_0(.dout(w_dff_A_u7lIUA0f9_0),.din(w_dff_A_jMVx26Eo7_0),.clk(gclk));
	jdff dff_A_u7lIUA0f9_0(.dout(w_dff_A_OXHogqZl0_0),.din(w_dff_A_u7lIUA0f9_0),.clk(gclk));
	jdff dff_A_OXHogqZl0_0(.dout(w_dff_A_aFDQzf0f6_0),.din(w_dff_A_OXHogqZl0_0),.clk(gclk));
	jdff dff_A_aFDQzf0f6_0(.dout(w_dff_A_Pe7egUoa6_0),.din(w_dff_A_aFDQzf0f6_0),.clk(gclk));
	jdff dff_A_Pe7egUoa6_0(.dout(w_dff_A_YuQ5v5OO5_0),.din(w_dff_A_Pe7egUoa6_0),.clk(gclk));
	jdff dff_A_YuQ5v5OO5_0(.dout(w_dff_A_CF9Du5FX7_0),.din(w_dff_A_YuQ5v5OO5_0),.clk(gclk));
	jdff dff_A_CF9Du5FX7_0(.dout(G699),.din(w_dff_A_CF9Du5FX7_0),.clk(gclk));
	jdff dff_A_gyEHSMrf9_2(.dout(w_dff_A_nUEvxDSH5_0),.din(w_dff_A_gyEHSMrf9_2),.clk(gclk));
	jdff dff_A_nUEvxDSH5_0(.dout(w_dff_A_6gwONjtW0_0),.din(w_dff_A_nUEvxDSH5_0),.clk(gclk));
	jdff dff_A_6gwONjtW0_0(.dout(w_dff_A_p98PBW9Q3_0),.din(w_dff_A_6gwONjtW0_0),.clk(gclk));
	jdff dff_A_p98PBW9Q3_0(.dout(w_dff_A_MG9fIiLi9_0),.din(w_dff_A_p98PBW9Q3_0),.clk(gclk));
	jdff dff_A_MG9fIiLi9_0(.dout(w_dff_A_xScfjUXN6_0),.din(w_dff_A_MG9fIiLi9_0),.clk(gclk));
	jdff dff_A_xScfjUXN6_0(.dout(w_dff_A_n5ZA8VPH5_0),.din(w_dff_A_xScfjUXN6_0),.clk(gclk));
	jdff dff_A_n5ZA8VPH5_0(.dout(w_dff_A_tuWa77KN8_0),.din(w_dff_A_n5ZA8VPH5_0),.clk(gclk));
	jdff dff_A_tuWa77KN8_0(.dout(w_dff_A_ubA97bsl7_0),.din(w_dff_A_tuWa77KN8_0),.clk(gclk));
	jdff dff_A_ubA97bsl7_0(.dout(G702),.din(w_dff_A_ubA97bsl7_0),.clk(gclk));
	jdff dff_A_6D6rviAx0_2(.dout(w_dff_A_go1YCpUD8_0),.din(w_dff_A_6D6rviAx0_2),.clk(gclk));
	jdff dff_A_go1YCpUD8_0(.dout(w_dff_A_d0mWpsIG6_0),.din(w_dff_A_go1YCpUD8_0),.clk(gclk));
	jdff dff_A_d0mWpsIG6_0(.dout(w_dff_A_d1AauKi04_0),.din(w_dff_A_d0mWpsIG6_0),.clk(gclk));
	jdff dff_A_d1AauKi04_0(.dout(w_dff_A_VnZF5srs2_0),.din(w_dff_A_d1AauKi04_0),.clk(gclk));
	jdff dff_A_VnZF5srs2_0(.dout(w_dff_A_tsj9VRhx1_0),.din(w_dff_A_VnZF5srs2_0),.clk(gclk));
	jdff dff_A_tsj9VRhx1_0(.dout(w_dff_A_8ZQBge4d2_0),.din(w_dff_A_tsj9VRhx1_0),.clk(gclk));
	jdff dff_A_8ZQBge4d2_0(.dout(G818),.din(w_dff_A_8ZQBge4d2_0),.clk(gclk));
	jdff dff_A_yfUFm8z19_2(.dout(w_dff_A_ipkVkOPj4_0),.din(w_dff_A_yfUFm8z19_2),.clk(gclk));
	jdff dff_A_ipkVkOPj4_0(.dout(w_dff_A_nktSdCDh8_0),.din(w_dff_A_ipkVkOPj4_0),.clk(gclk));
	jdff dff_A_nktSdCDh8_0(.dout(w_dff_A_WdVzl2oX6_0),.din(w_dff_A_nktSdCDh8_0),.clk(gclk));
	jdff dff_A_WdVzl2oX6_0(.dout(w_dff_A_DsKGo98l7_0),.din(w_dff_A_WdVzl2oX6_0),.clk(gclk));
	jdff dff_A_DsKGo98l7_0(.dout(w_dff_A_rNDqtyMM3_0),.din(w_dff_A_DsKGo98l7_0),.clk(gclk));
	jdff dff_A_rNDqtyMM3_0(.dout(w_dff_A_ARy93q053_0),.din(w_dff_A_rNDqtyMM3_0),.clk(gclk));
	jdff dff_A_ARy93q053_0(.dout(w_dff_A_pkJbzM3e8_0),.din(w_dff_A_ARy93q053_0),.clk(gclk));
	jdff dff_A_pkJbzM3e8_0(.dout(w_dff_A_61roVGaG6_0),.din(w_dff_A_pkJbzM3e8_0),.clk(gclk));
	jdff dff_A_61roVGaG6_0(.dout(w_dff_A_uaOdc2z75_0),.din(w_dff_A_61roVGaG6_0),.clk(gclk));
	jdff dff_A_uaOdc2z75_0(.dout(G813),.din(w_dff_A_uaOdc2z75_0),.clk(gclk));
	jdff dff_A_JP0ztOG01_1(.dout(w_dff_A_XteXsbNS7_0),.din(w_dff_A_JP0ztOG01_1),.clk(gclk));
	jdff dff_A_XteXsbNS7_0(.dout(w_dff_A_3J3C8zlF7_0),.din(w_dff_A_XteXsbNS7_0),.clk(gclk));
	jdff dff_A_3J3C8zlF7_0(.dout(w_dff_A_IbKSO0nV9_0),.din(w_dff_A_3J3C8zlF7_0),.clk(gclk));
	jdff dff_A_IbKSO0nV9_0(.dout(w_dff_A_0i01aeYu0_0),.din(w_dff_A_IbKSO0nV9_0),.clk(gclk));
	jdff dff_A_0i01aeYu0_0(.dout(w_dff_A_mHR4cvL27_0),.din(w_dff_A_0i01aeYu0_0),.clk(gclk));
	jdff dff_A_mHR4cvL27_0(.dout(w_dff_A_gHpjmiQs1_0),.din(w_dff_A_mHR4cvL27_0),.clk(gclk));
	jdff dff_A_gHpjmiQs1_0(.dout(G824),.din(w_dff_A_gHpjmiQs1_0),.clk(gclk));
	jdff dff_A_BfQNuq0O6_1(.dout(w_dff_A_XBmdcbDl4_0),.din(w_dff_A_BfQNuq0O6_1),.clk(gclk));
	jdff dff_A_XBmdcbDl4_0(.dout(w_dff_A_KFbpGayW2_0),.din(w_dff_A_XBmdcbDl4_0),.clk(gclk));
	jdff dff_A_KFbpGayW2_0(.dout(w_dff_A_K8ITLv3f5_0),.din(w_dff_A_KFbpGayW2_0),.clk(gclk));
	jdff dff_A_K8ITLv3f5_0(.dout(w_dff_A_MqXftXCi9_0),.din(w_dff_A_K8ITLv3f5_0),.clk(gclk));
	jdff dff_A_MqXftXCi9_0(.dout(w_dff_A_QVQFkG3y9_0),.din(w_dff_A_MqXftXCi9_0),.clk(gclk));
	jdff dff_A_QVQFkG3y9_0(.dout(w_dff_A_JlobzhOr4_0),.din(w_dff_A_QVQFkG3y9_0),.clk(gclk));
	jdff dff_A_JlobzhOr4_0(.dout(w_dff_A_U2IuuViG0_0),.din(w_dff_A_JlobzhOr4_0),.clk(gclk));
	jdff dff_A_U2IuuViG0_0(.dout(G826),.din(w_dff_A_U2IuuViG0_0),.clk(gclk));
	jdff dff_A_EMYGxBMS3_1(.dout(w_dff_A_2JoAGth54_0),.din(w_dff_A_EMYGxBMS3_1),.clk(gclk));
	jdff dff_A_2JoAGth54_0(.dout(w_dff_A_U3tmic7N8_0),.din(w_dff_A_2JoAGth54_0),.clk(gclk));
	jdff dff_A_U3tmic7N8_0(.dout(w_dff_A_BP2h6ADM8_0),.din(w_dff_A_U3tmic7N8_0),.clk(gclk));
	jdff dff_A_BP2h6ADM8_0(.dout(w_dff_A_hm9aLquT5_0),.din(w_dff_A_BP2h6ADM8_0),.clk(gclk));
	jdff dff_A_hm9aLquT5_0(.dout(w_dff_A_MdeDkIKL4_0),.din(w_dff_A_hm9aLquT5_0),.clk(gclk));
	jdff dff_A_MdeDkIKL4_0(.dout(w_dff_A_PC2vSuin3_0),.din(w_dff_A_MdeDkIKL4_0),.clk(gclk));
	jdff dff_A_PC2vSuin3_0(.dout(G828),.din(w_dff_A_PC2vSuin3_0),.clk(gclk));
	jdff dff_A_lO1QpRnm5_1(.dout(w_dff_A_gSlZSXwH6_0),.din(w_dff_A_lO1QpRnm5_1),.clk(gclk));
	jdff dff_A_gSlZSXwH6_0(.dout(w_dff_A_4oM9h1By1_0),.din(w_dff_A_gSlZSXwH6_0),.clk(gclk));
	jdff dff_A_4oM9h1By1_0(.dout(w_dff_A_602QKs9Q0_0),.din(w_dff_A_4oM9h1By1_0),.clk(gclk));
	jdff dff_A_602QKs9Q0_0(.dout(w_dff_A_SdQ38IQz7_0),.din(w_dff_A_602QKs9Q0_0),.clk(gclk));
	jdff dff_A_SdQ38IQz7_0(.dout(w_dff_A_HT0lfgmT0_0),.din(w_dff_A_SdQ38IQz7_0),.clk(gclk));
	jdff dff_A_HT0lfgmT0_0(.dout(w_dff_A_sJPm82kd9_0),.din(w_dff_A_HT0lfgmT0_0),.clk(gclk));
	jdff dff_A_sJPm82kd9_0(.dout(w_dff_A_3NYxN2fx2_0),.din(w_dff_A_sJPm82kd9_0),.clk(gclk));
	jdff dff_A_3NYxN2fx2_0(.dout(w_dff_A_rrEDsG667_0),.din(w_dff_A_3NYxN2fx2_0),.clk(gclk));
	jdff dff_A_rrEDsG667_0(.dout(w_dff_A_jRoTd1a24_0),.din(w_dff_A_rrEDsG667_0),.clk(gclk));
	jdff dff_A_jRoTd1a24_0(.dout(w_dff_A_ElkFPYjj3_0),.din(w_dff_A_jRoTd1a24_0),.clk(gclk));
	jdff dff_A_ElkFPYjj3_0(.dout(w_dff_A_bVfZZB9E3_0),.din(w_dff_A_ElkFPYjj3_0),.clk(gclk));
	jdff dff_A_bVfZZB9E3_0(.dout(G830),.din(w_dff_A_bVfZZB9E3_0),.clk(gclk));
	jdff dff_A_895FGv130_2(.dout(w_dff_A_iYY8G84B7_0),.din(w_dff_A_895FGv130_2),.clk(gclk));
	jdff dff_A_iYY8G84B7_0(.dout(w_dff_A_wAm89jr86_0),.din(w_dff_A_iYY8G84B7_0),.clk(gclk));
	jdff dff_A_wAm89jr86_0(.dout(w_dff_A_onCEKMEY6_0),.din(w_dff_A_wAm89jr86_0),.clk(gclk));
	jdff dff_A_onCEKMEY6_0(.dout(w_dff_A_ofDz5DV79_0),.din(w_dff_A_onCEKMEY6_0),.clk(gclk));
	jdff dff_A_ofDz5DV79_0(.dout(w_dff_A_64wp8i3q5_0),.din(w_dff_A_ofDz5DV79_0),.clk(gclk));
	jdff dff_A_64wp8i3q5_0(.dout(w_dff_A_XJybgXKZ4_0),.din(w_dff_A_64wp8i3q5_0),.clk(gclk));
	jdff dff_A_XJybgXKZ4_0(.dout(w_dff_A_8JSSzpdP3_0),.din(w_dff_A_XJybgXKZ4_0),.clk(gclk));
	jdff dff_A_8JSSzpdP3_0(.dout(w_dff_A_NqzCJA5O3_0),.din(w_dff_A_8JSSzpdP3_0),.clk(gclk));
	jdff dff_A_NqzCJA5O3_0(.dout(w_dff_A_K4j0spcf0_0),.din(w_dff_A_NqzCJA5O3_0),.clk(gclk));
	jdff dff_A_K4j0spcf0_0(.dout(w_dff_A_GcND7V5D3_0),.din(w_dff_A_K4j0spcf0_0),.clk(gclk));
	jdff dff_A_GcND7V5D3_0(.dout(w_dff_A_JgKoGoOG6_0),.din(w_dff_A_GcND7V5D3_0),.clk(gclk));
	jdff dff_A_JgKoGoOG6_0(.dout(w_dff_A_0OuHfazO0_0),.din(w_dff_A_JgKoGoOG6_0),.clk(gclk));
	jdff dff_A_0OuHfazO0_0(.dout(w_dff_A_7qxCi5Hh4_0),.din(w_dff_A_0OuHfazO0_0),.clk(gclk));
	jdff dff_A_7qxCi5Hh4_0(.dout(w_dff_A_9g95h1Z50_0),.din(w_dff_A_7qxCi5Hh4_0),.clk(gclk));
	jdff dff_A_9g95h1Z50_0(.dout(w_dff_A_Pop8U8747_0),.din(w_dff_A_9g95h1Z50_0),.clk(gclk));
	jdff dff_A_Pop8U8747_0(.dout(w_dff_A_HT2ozZiF6_0),.din(w_dff_A_Pop8U8747_0),.clk(gclk));
	jdff dff_A_HT2ozZiF6_0(.dout(G854),.din(w_dff_A_HT2ozZiF6_0),.clk(gclk));
	jdff dff_A_6KcRPZEY1_1(.dout(w_dff_A_VL4u1syn8_0),.din(w_dff_A_6KcRPZEY1_1),.clk(gclk));
	jdff dff_A_VL4u1syn8_0(.dout(w_dff_A_qq8TKOja5_0),.din(w_dff_A_VL4u1syn8_0),.clk(gclk));
	jdff dff_A_qq8TKOja5_0(.dout(w_dff_A_ovPhs7Em2_0),.din(w_dff_A_qq8TKOja5_0),.clk(gclk));
	jdff dff_A_ovPhs7Em2_0(.dout(w_dff_A_TZKGaMGi8_0),.din(w_dff_A_ovPhs7Em2_0),.clk(gclk));
	jdff dff_A_TZKGaMGi8_0(.dout(w_dff_A_XuaPGdcM1_0),.din(w_dff_A_TZKGaMGi8_0),.clk(gclk));
	jdff dff_A_XuaPGdcM1_0(.dout(G863),.din(w_dff_A_XuaPGdcM1_0),.clk(gclk));
	jdff dff_A_8HK7cpkl2_1(.dout(w_dff_A_XHwCdkcM9_0),.din(w_dff_A_8HK7cpkl2_1),.clk(gclk));
	jdff dff_A_XHwCdkcM9_0(.dout(w_dff_A_RMCiEWdP1_0),.din(w_dff_A_XHwCdkcM9_0),.clk(gclk));
	jdff dff_A_RMCiEWdP1_0(.dout(w_dff_A_ndgumlmq8_0),.din(w_dff_A_RMCiEWdP1_0),.clk(gclk));
	jdff dff_A_ndgumlmq8_0(.dout(w_dff_A_JKwEgMNF6_0),.din(w_dff_A_ndgumlmq8_0),.clk(gclk));
	jdff dff_A_JKwEgMNF6_0(.dout(w_dff_A_8y39fQ1n8_0),.din(w_dff_A_JKwEgMNF6_0),.clk(gclk));
	jdff dff_A_8y39fQ1n8_0(.dout(w_dff_A_qwXK7NWB1_0),.din(w_dff_A_8y39fQ1n8_0),.clk(gclk));
	jdff dff_A_qwXK7NWB1_0(.dout(w_dff_A_N9gBLWNS1_0),.din(w_dff_A_qwXK7NWB1_0),.clk(gclk));
	jdff dff_A_N9gBLWNS1_0(.dout(w_dff_A_T9EiKK7U8_0),.din(w_dff_A_N9gBLWNS1_0),.clk(gclk));
	jdff dff_A_T9EiKK7U8_0(.dout(G865),.din(w_dff_A_T9EiKK7U8_0),.clk(gclk));
	jdff dff_A_ybOm80nJ7_1(.dout(w_dff_A_pllF5Uob6_0),.din(w_dff_A_ybOm80nJ7_1),.clk(gclk));
	jdff dff_A_pllF5Uob6_0(.dout(w_dff_A_H5JPP1089_0),.din(w_dff_A_pllF5Uob6_0),.clk(gclk));
	jdff dff_A_H5JPP1089_0(.dout(w_dff_A_g4zNuHiz0_0),.din(w_dff_A_H5JPP1089_0),.clk(gclk));
	jdff dff_A_g4zNuHiz0_0(.dout(w_dff_A_tNXXiEgG1_0),.din(w_dff_A_g4zNuHiz0_0),.clk(gclk));
	jdff dff_A_tNXXiEgG1_0(.dout(w_dff_A_NGxlt3pd2_0),.din(w_dff_A_tNXXiEgG1_0),.clk(gclk));
	jdff dff_A_NGxlt3pd2_0(.dout(w_dff_A_N2KlKkZ48_0),.din(w_dff_A_NGxlt3pd2_0),.clk(gclk));
	jdff dff_A_N2KlKkZ48_0(.dout(G867),.din(w_dff_A_N2KlKkZ48_0),.clk(gclk));
	jdff dff_A_YxXv40kT5_1(.dout(w_dff_A_nr5st40n4_0),.din(w_dff_A_YxXv40kT5_1),.clk(gclk));
	jdff dff_A_nr5st40n4_0(.dout(w_dff_A_lEjOuwSH1_0),.din(w_dff_A_nr5st40n4_0),.clk(gclk));
	jdff dff_A_lEjOuwSH1_0(.dout(w_dff_A_eopy3nFu1_0),.din(w_dff_A_lEjOuwSH1_0),.clk(gclk));
	jdff dff_A_eopy3nFu1_0(.dout(w_dff_A_2mUDQUYi4_0),.din(w_dff_A_eopy3nFu1_0),.clk(gclk));
	jdff dff_A_2mUDQUYi4_0(.dout(w_dff_A_eJneS3RH0_0),.din(w_dff_A_2mUDQUYi4_0),.clk(gclk));
	jdff dff_A_eJneS3RH0_0(.dout(w_dff_A_TOixvbg22_0),.din(w_dff_A_eJneS3RH0_0),.clk(gclk));
	jdff dff_A_TOixvbg22_0(.dout(w_dff_A_oERts3xA4_0),.din(w_dff_A_TOixvbg22_0),.clk(gclk));
	jdff dff_A_oERts3xA4_0(.dout(w_dff_A_aSH3WLwF9_0),.din(w_dff_A_oERts3xA4_0),.clk(gclk));
	jdff dff_A_aSH3WLwF9_0(.dout(w_dff_A_UA3c6uSj0_0),.din(w_dff_A_aSH3WLwF9_0),.clk(gclk));
	jdff dff_A_UA3c6uSj0_0(.dout(G869),.din(w_dff_A_UA3c6uSj0_0),.clk(gclk));
	jdff dff_A_9sxuK1rx0_2(.dout(w_dff_A_8Vbysi9b2_0),.din(w_dff_A_9sxuK1rx0_2),.clk(gclk));
	jdff dff_A_8Vbysi9b2_0(.dout(w_dff_A_WpWKO3K38_0),.din(w_dff_A_8Vbysi9b2_0),.clk(gclk));
	jdff dff_A_WpWKO3K38_0(.dout(w_dff_A_0LeTCrT14_0),.din(w_dff_A_WpWKO3K38_0),.clk(gclk));
	jdff dff_A_0LeTCrT14_0(.dout(G712),.din(w_dff_A_0LeTCrT14_0),.clk(gclk));
	jdff dff_A_9ZseDTY54_2(.dout(w_dff_A_HVf0SUn03_0),.din(w_dff_A_9ZseDTY54_2),.clk(gclk));
	jdff dff_A_HVf0SUn03_0(.dout(w_dff_A_dizJkHxB8_0),.din(w_dff_A_HVf0SUn03_0),.clk(gclk));
	jdff dff_A_dizJkHxB8_0(.dout(G727),.din(w_dff_A_dizJkHxB8_0),.clk(gclk));
	jdff dff_A_1o2NTLEO3_2(.dout(w_dff_A_wmaiJ6M16_0),.din(w_dff_A_1o2NTLEO3_2),.clk(gclk));
	jdff dff_A_wmaiJ6M16_0(.dout(w_dff_A_oJAdkQg52_0),.din(w_dff_A_wmaiJ6M16_0),.clk(gclk));
	jdff dff_A_oJAdkQg52_0(.dout(w_dff_A_ejDAC4ma8_0),.din(w_dff_A_oJAdkQg52_0),.clk(gclk));
	jdff dff_A_ejDAC4ma8_0(.dout(G732),.din(w_dff_A_ejDAC4ma8_0),.clk(gclk));
	jdff dff_A_UFCuDxvQ5_2(.dout(w_dff_A_nwSLAHCZ1_0),.din(w_dff_A_UFCuDxvQ5_2),.clk(gclk));
	jdff dff_A_nwSLAHCZ1_0(.dout(w_dff_A_UsCiql2t9_0),.din(w_dff_A_nwSLAHCZ1_0),.clk(gclk));
	jdff dff_A_UsCiql2t9_0(.dout(w_dff_A_cfobi81r2_0),.din(w_dff_A_UsCiql2t9_0),.clk(gclk));
	jdff dff_A_cfobi81r2_0(.dout(G737),.din(w_dff_A_cfobi81r2_0),.clk(gclk));
	jdff dff_A_LJKa69Qm9_2(.dout(w_dff_A_6DDb7pdb3_0),.din(w_dff_A_LJKa69Qm9_2),.clk(gclk));
	jdff dff_A_6DDb7pdb3_0(.dout(w_dff_A_u4CHBI0j2_0),.din(w_dff_A_6DDb7pdb3_0),.clk(gclk));
	jdff dff_A_u4CHBI0j2_0(.dout(w_dff_A_jXQAFSfX9_0),.din(w_dff_A_u4CHBI0j2_0),.clk(gclk));
	jdff dff_A_jXQAFSfX9_0(.dout(w_dff_A_ur4sohGn4_0),.din(w_dff_A_jXQAFSfX9_0),.clk(gclk));
	jdff dff_A_ur4sohGn4_0(.dout(G742),.din(w_dff_A_ur4sohGn4_0),.clk(gclk));
	jdff dff_A_YNkz6Tgg6_2(.dout(w_dff_A_mukuAoNM5_0),.din(w_dff_A_YNkz6Tgg6_2),.clk(gclk));
	jdff dff_A_mukuAoNM5_0(.dout(w_dff_A_pycDjWzk1_0),.din(w_dff_A_mukuAoNM5_0),.clk(gclk));
	jdff dff_A_pycDjWzk1_0(.dout(w_dff_A_6IPccs4l1_0),.din(w_dff_A_pycDjWzk1_0),.clk(gclk));
	jdff dff_A_6IPccs4l1_0(.dout(G772),.din(w_dff_A_6IPccs4l1_0),.clk(gclk));
	jdff dff_A_iVlpqlh74_2(.dout(w_dff_A_c6sjhufo6_0),.din(w_dff_A_iVlpqlh74_2),.clk(gclk));
	jdff dff_A_c6sjhufo6_0(.dout(w_dff_A_elfhUkaj9_0),.din(w_dff_A_c6sjhufo6_0),.clk(gclk));
	jdff dff_A_elfhUkaj9_0(.dout(w_dff_A_lnSRuheC9_0),.din(w_dff_A_elfhUkaj9_0),.clk(gclk));
	jdff dff_A_lnSRuheC9_0(.dout(G777),.din(w_dff_A_lnSRuheC9_0),.clk(gclk));
	jdff dff_A_8lfa568n2_2(.dout(w_dff_A_L4953zrj5_0),.din(w_dff_A_8lfa568n2_2),.clk(gclk));
	jdff dff_A_L4953zrj5_0(.dout(w_dff_A_tvjJ54RO0_0),.din(w_dff_A_L4953zrj5_0),.clk(gclk));
	jdff dff_A_tvjJ54RO0_0(.dout(w_dff_A_p0FFlBzA3_0),.din(w_dff_A_tvjJ54RO0_0),.clk(gclk));
	jdff dff_A_p0FFlBzA3_0(.dout(w_dff_A_xSGnrJLD0_0),.din(w_dff_A_p0FFlBzA3_0),.clk(gclk));
	jdff dff_A_xSGnrJLD0_0(.dout(G782),.din(w_dff_A_xSGnrJLD0_0),.clk(gclk));
	jdff dff_A_iUpifcdH2_2(.dout(w_dff_A_lQAtOq602_0),.din(w_dff_A_iUpifcdH2_2),.clk(gclk));
	jdff dff_A_lQAtOq602_0(.dout(w_dff_A_44bWtlZI3_0),.din(w_dff_A_lQAtOq602_0),.clk(gclk));
	jdff dff_A_44bWtlZI3_0(.dout(w_dff_A_qSB0BDZw9_0),.din(w_dff_A_44bWtlZI3_0),.clk(gclk));
	jdff dff_A_qSB0BDZw9_0(.dout(G645),.din(w_dff_A_qSB0BDZw9_0),.clk(gclk));
	jdff dff_A_2tJJd17T5_2(.dout(w_dff_A_lCoSCkNt9_0),.din(w_dff_A_2tJJd17T5_2),.clk(gclk));
	jdff dff_A_lCoSCkNt9_0(.dout(w_dff_A_xk7Cz47b9_0),.din(w_dff_A_lCoSCkNt9_0),.clk(gclk));
	jdff dff_A_xk7Cz47b9_0(.dout(G648),.din(w_dff_A_xk7Cz47b9_0),.clk(gclk));
	jdff dff_A_8Et3bTWw1_2(.dout(w_dff_A_q80xYIbs9_0),.din(w_dff_A_8Et3bTWw1_2),.clk(gclk));
	jdff dff_A_q80xYIbs9_0(.dout(w_dff_A_hEQsiTAf9_0),.din(w_dff_A_q80xYIbs9_0),.clk(gclk));
	jdff dff_A_hEQsiTAf9_0(.dout(G651),.din(w_dff_A_hEQsiTAf9_0),.clk(gclk));
	jdff dff_A_W8e3w3NF5_2(.dout(w_dff_A_iFsWFNfO5_0),.din(w_dff_A_W8e3w3NF5_2),.clk(gclk));
	jdff dff_A_iFsWFNfO5_0(.dout(G654),.din(w_dff_A_iFsWFNfO5_0),.clk(gclk));
	jdff dff_A_JhrkJhl39_2(.dout(w_dff_A_lkCp01sO9_0),.din(w_dff_A_JhrkJhl39_2),.clk(gclk));
	jdff dff_A_lkCp01sO9_0(.dout(w_dff_A_XYb04rwh0_0),.din(w_dff_A_lkCp01sO9_0),.clk(gclk));
	jdff dff_A_XYb04rwh0_0(.dout(w_dff_A_FsMUJCpF2_0),.din(w_dff_A_XYb04rwh0_0),.clk(gclk));
	jdff dff_A_FsMUJCpF2_0(.dout(G679),.din(w_dff_A_FsMUJCpF2_0),.clk(gclk));
	jdff dff_A_EU9AjEys6_2(.dout(w_dff_A_gBeoBIe98_0),.din(w_dff_A_EU9AjEys6_2),.clk(gclk));
	jdff dff_A_gBeoBIe98_0(.dout(w_dff_A_Agly4Fzj9_0),.din(w_dff_A_gBeoBIe98_0),.clk(gclk));
	jdff dff_A_Agly4Fzj9_0(.dout(G682),.din(w_dff_A_Agly4Fzj9_0),.clk(gclk));
	jdff dff_A_BvotNGEA0_2(.dout(w_dff_A_Kib1mxWx5_0),.din(w_dff_A_BvotNGEA0_2),.clk(gclk));
	jdff dff_A_Kib1mxWx5_0(.dout(w_dff_A_Bbj03Fq73_0),.din(w_dff_A_Kib1mxWx5_0),.clk(gclk));
	jdff dff_A_Bbj03Fq73_0(.dout(G685),.din(w_dff_A_Bbj03Fq73_0),.clk(gclk));
	jdff dff_A_et8vM2y52_2(.dout(w_dff_A_5Kjw3Tkd6_0),.din(w_dff_A_et8vM2y52_2),.clk(gclk));
	jdff dff_A_5Kjw3Tkd6_0(.dout(w_dff_A_LMlsjDrx1_0),.din(w_dff_A_5Kjw3Tkd6_0),.clk(gclk));
	jdff dff_A_LMlsjDrx1_0(.dout(G688),.din(w_dff_A_LMlsjDrx1_0),.clk(gclk));
	jdff dff_A_EMPb80Xy4_2(.dout(w_dff_A_LzkmumMs1_0),.din(w_dff_A_EMPb80Xy4_2),.clk(gclk));
	jdff dff_A_LzkmumMs1_0(.dout(w_dff_A_sTH0gPWI1_0),.din(w_dff_A_LzkmumMs1_0),.clk(gclk));
	jdff dff_A_sTH0gPWI1_0(.dout(w_dff_A_cmeWtwhA1_0),.din(w_dff_A_sTH0gPWI1_0),.clk(gclk));
	jdff dff_A_cmeWtwhA1_0(.dout(w_dff_A_RaE1t2gH7_0),.din(w_dff_A_cmeWtwhA1_0),.clk(gclk));
	jdff dff_A_RaE1t2gH7_0(.dout(w_dff_A_qhYBnWPj1_0),.din(w_dff_A_RaE1t2gH7_0),.clk(gclk));
	jdff dff_A_qhYBnWPj1_0(.dout(G843),.din(w_dff_A_qhYBnWPj1_0),.clk(gclk));
	jdff dff_A_d5yH2TQb2_2(.dout(w_dff_A_0DNiYuTX8_0),.din(w_dff_A_d5yH2TQb2_2),.clk(gclk));
	jdff dff_A_0DNiYuTX8_0(.dout(w_dff_A_z297T3Oe8_0),.din(w_dff_A_0DNiYuTX8_0),.clk(gclk));
	jdff dff_A_z297T3Oe8_0(.dout(w_dff_A_o0pkMQJ63_0),.din(w_dff_A_z297T3Oe8_0),.clk(gclk));
	jdff dff_A_o0pkMQJ63_0(.dout(w_dff_A_KtDh1uLu6_0),.din(w_dff_A_o0pkMQJ63_0),.clk(gclk));
	jdff dff_A_KtDh1uLu6_0(.dout(w_dff_A_Z6lxaLEo3_0),.din(w_dff_A_KtDh1uLu6_0),.clk(gclk));
	jdff dff_A_Z6lxaLEo3_0(.dout(G882),.din(w_dff_A_Z6lxaLEo3_0),.clk(gclk));
	jdff dff_A_uayLeJHg8_2(.dout(G767),.din(w_dff_A_uayLeJHg8_2),.clk(gclk));
	jdff dff_A_Y9j4iuZu8_2(.dout(G807),.din(w_dff_A_Y9j4iuZu8_2),.clk(gclk));
endmodule

