/*

c7552:
	jxor: 228
	jspl: 345
	jspl3: 346
	jnot: 270
	jdff: 2062
	jor: 395
	jand: 513

Summary:
	jxor: 228
	jspl: 345
	jspl3: 346
	jnot: 270
	jdff: 2062
	jor: 395
	jand: 513

The maximum logic level gap of any gate:
	c7552: 21
*/

module rf_c7552(gclk, G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526, G4528, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399);
	input gclk;
	input G1;
	input G5;
	input G9;
	input G12;
	input G15;
	input G18;
	input G23;
	input G26;
	input G29;
	input G32;
	input G35;
	input G38;
	input G41;
	input G44;
	input G47;
	input G50;
	input G53;
	input G54;
	input G55;
	input G56;
	input G57;
	input G58;
	input G59;
	input G60;
	input G61;
	input G62;
	input G63;
	input G64;
	input G65;
	input G66;
	input G69;
	input G70;
	input G73;
	input G74;
	input G75;
	input G76;
	input G77;
	input G78;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G84;
	input G85;
	input G86;
	input G87;
	input G88;
	input G89;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G110;
	input G111;
	input G112;
	input G113;
	input G114;
	input G115;
	input G118;
	input G121;
	input G124;
	input G127;
	input G130;
	input G133;
	input G134;
	input G135;
	input G138;
	input G141;
	input G144;
	input G147;
	input G150;
	input G151;
	input G152;
	input G153;
	input G154;
	input G155;
	input G156;
	input G157;
	input G158;
	input G159;
	input G160;
	input G161;
	input G162;
	input G163;
	input G164;
	input G165;
	input G166;
	input G167;
	input G168;
	input G169;
	input G170;
	input G171;
	input G172;
	input G173;
	input G174;
	input G175;
	input G176;
	input G177;
	input G178;
	input G179;
	input G180;
	input G181;
	input G182;
	input G183;
	input G184;
	input G185;
	input G186;
	input G187;
	input G188;
	input G189;
	input G190;
	input G191;
	input G192;
	input G193;
	input G194;
	input G195;
	input G196;
	input G197;
	input G198;
	input G199;
	input G200;
	input G201;
	input G202;
	input G203;
	input G204;
	input G205;
	input G206;
	input G207;
	input G208;
	input G209;
	input G210;
	input G211;
	input G212;
	input G213;
	input G214;
	input G215;
	input G216;
	input G217;
	input G218;
	input G219;
	input G220;
	input G221;
	input G222;
	input G223;
	input G224;
	input G225;
	input G226;
	input G227;
	input G228;
	input G229;
	input G230;
	input G231;
	input G232;
	input G233;
	input G234;
	input G235;
	input G236;
	input G237;
	input G238;
	input G239;
	input G240;
	input G339;
	input G1197;
	input G1455;
	input G1459;
	input G1462;
	input G1469;
	input G1480;
	input G1486;
	input G1492;
	input G1496;
	input G2204;
	input G2208;
	input G2211;
	input G2218;
	input G2224;
	input G2230;
	input G2236;
	input G2239;
	input G2247;
	input G2253;
	input G2256;
	input G3698;
	input G3701;
	input G3705;
	input G3711;
	input G3717;
	input G3723;
	input G3729;
	input G3737;
	input G3743;
	input G3749;
	input G4393;
	input G4394;
	input G4400;
	input G4405;
	input G4410;
	input G4415;
	input G4420;
	input G4427;
	input G4432;
	input G4437;
	input G4526;
	input G4528;
	output G2;
	output G3;
	output G450;
	output G448;
	output G444;
	output G442;
	output G440;
	output G438;
	output G496;
	output G494;
	output G492;
	output G490;
	output G488;
	output G486;
	output G484;
	output G482;
	output G480;
	output G560;
	output G542;
	output G558;
	output G556;
	output G554;
	output G552;
	output G550;
	output G548;
	output G546;
	output G544;
	output G540;
	output G538;
	output G536;
	output G534;
	output G532;
	output G530;
	output G528;
	output G526;
	output G524;
	output G279;
	output G436;
	output G478;
	output G522;
	output G402;
	output G404;
	output G406;
	output G408;
	output G410;
	output G432;
	output G446;
	output G284;
	output G286;
	output G289;
	output G292;
	output G341;
	output G281;
	output G453;
	output G278;
	output G373;
	output G246;
	output G258;
	output G264;
	output G270;
	output G388;
	output G391;
	output G394;
	output G397;
	output G376;
	output G379;
	output G382;
	output G385;
	output G412;
	output G414;
	output G416;
	output G249;
	output G295;
	output G324;
	output G252;
	output G276;
	output G310;
	output G313;
	output G316;
	output G319;
	output G327;
	output G330;
	output G333;
	output G336;
	output G418;
	output G273;
	output G298;
	output G301;
	output G304;
	output G307;
	output G344;
	output G422;
	output G469;
	output G419;
	output G471;
	output G359;
	output G362;
	output G365;
	output G368;
	output G347;
	output G350;
	output G353;
	output G356;
	output G321;
	output G338;
	output G370;
	output G399;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n347;
	wire n348;
	wire n349;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1134;
	wire n1136;
	wire n1137;
	wire n1139;
	wire n1140;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1146;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1410;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1417;
	wire n1418;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1429;
	wire n1430;
	wire n1432;
	wire n1433;
	wire n1435;
	wire n1436;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1451;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1477;
	wire n1479;
	wire n1480;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1490;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[2:0] w_G5_0;
	wire[2:0] w_G5_1;
	wire[2:0] w_G15_0;
	wire[2:0] w_G18_0;
	wire[2:0] w_G18_1;
	wire[2:0] w_G18_2;
	wire[2:0] w_G18_3;
	wire[2:0] w_G18_4;
	wire[2:0] w_G18_5;
	wire[2:0] w_G18_6;
	wire[2:0] w_G18_7;
	wire[2:0] w_G18_8;
	wire[2:0] w_G18_9;
	wire[2:0] w_G18_10;
	wire[2:0] w_G18_11;
	wire[2:0] w_G18_12;
	wire[2:0] w_G18_13;
	wire[2:0] w_G18_14;
	wire[2:0] w_G18_15;
	wire[2:0] w_G18_16;
	wire[2:0] w_G18_17;
	wire[2:0] w_G18_18;
	wire[2:0] w_G18_19;
	wire[2:0] w_G18_20;
	wire[2:0] w_G18_21;
	wire[2:0] w_G18_22;
	wire[2:0] w_G18_23;
	wire[2:0] w_G18_24;
	wire[2:0] w_G18_25;
	wire[2:0] w_G18_26;
	wire[2:0] w_G18_27;
	wire[2:0] w_G18_28;
	wire[2:0] w_G18_29;
	wire[2:0] w_G18_30;
	wire[2:0] w_G18_31;
	wire[2:0] w_G18_32;
	wire[2:0] w_G18_33;
	wire[2:0] w_G18_34;
	wire[2:0] w_G18_35;
	wire[2:0] w_G18_36;
	wire[2:0] w_G18_37;
	wire[2:0] w_G18_38;
	wire[2:0] w_G18_39;
	wire[2:0] w_G18_40;
	wire[2:0] w_G18_41;
	wire[2:0] w_G18_42;
	wire[2:0] w_G18_43;
	wire[2:0] w_G18_44;
	wire[2:0] w_G18_45;
	wire[2:0] w_G18_46;
	wire[2:0] w_G18_47;
	wire[2:0] w_G18_48;
	wire[2:0] w_G18_49;
	wire[2:0] w_G18_50;
	wire[2:0] w_G18_51;
	wire[2:0] w_G18_52;
	wire[2:0] w_G18_53;
	wire[2:0] w_G18_54;
	wire[2:0] w_G18_55;
	wire[2:0] w_G18_56;
	wire[2:0] w_G18_57;
	wire[2:0] w_G18_58;
	wire[2:0] w_G38_0;
	wire[2:0] w_G38_1;
	wire[2:0] w_G41_0;
	wire[1:0] w_G69_0;
	wire[1:0] w_G70_0;
	wire[2:0] w_G106_0;
	wire[1:0] w_G106_1;
	wire[1:0] w_G229_0;
	wire[2:0] w_G1455_0;
	wire[1:0] w_G1459_0;
	wire[2:0] w_G1462_0;
	wire[2:0] w_G1469_0;
	wire[1:0] w_G1469_1;
	wire[2:0] w_G1480_0;
	wire[2:0] w_G1486_0;
	wire[2:0] w_G1492_0;
	wire[1:0] w_G1492_1;
	wire[2:0] w_G1496_0;
	wire[2:0] w_G2204_0;
	wire[1:0] w_G2208_0;
	wire[2:0] w_G2211_0;
	wire[2:0] w_G2218_0;
	wire[2:0] w_G2224_0;
	wire[1:0] w_G2224_1;
	wire[2:0] w_G2230_0;
	wire[1:0] w_G2230_1;
	wire[2:0] w_G2236_0;
	wire[1:0] w_G2236_1;
	wire[2:0] w_G2239_0;
	wire[2:0] w_G2247_0;
	wire[2:0] w_G2253_0;
	wire[1:0] w_G2253_1;
	wire[2:0] w_G2256_0;
	wire[1:0] w_G2256_1;
	wire[1:0] w_G3698_0;
	wire[2:0] w_G3701_0;
	wire[1:0] w_G3701_1;
	wire[2:0] w_G3705_0;
	wire[2:0] w_G3705_1;
	wire[1:0] w_G3705_2;
	wire[2:0] w_G3711_0;
	wire[1:0] w_G3711_1;
	wire[2:0] w_G3717_0;
	wire[2:0] w_G3717_1;
	wire[1:0] w_G3717_2;
	wire[2:0] w_G3723_0;
	wire[1:0] w_G3723_1;
	wire[2:0] w_G3729_0;
	wire[1:0] w_G3729_1;
	wire[2:0] w_G3737_0;
	wire[1:0] w_G3737_1;
	wire[2:0] w_G3743_0;
	wire[2:0] w_G3743_1;
	wire[2:0] w_G3749_0;
	wire[1:0] w_G3749_1;
	wire[1:0] w_G4393_0;
	wire[2:0] w_G4394_0;
	wire[1:0] w_G4394_1;
	wire[2:0] w_G4400_0;
	wire[2:0] w_G4405_0;
	wire[2:0] w_G4405_1;
	wire[2:0] w_G4410_0;
	wire[1:0] w_G4410_1;
	wire[2:0] w_G4415_0;
	wire[1:0] w_G4415_1;
	wire[2:0] w_G4420_0;
	wire[1:0] w_G4427_0;
	wire[2:0] w_G4432_0;
	wire[1:0] w_G4432_1;
	wire[2:0] w_G4437_0;
	wire[2:0] w_G4526_0;
	wire[1:0] w_G4526_1;
	wire[2:0] w_G4528_0;
	wire w_G404_0;
	wire G404_fa_;
	wire w_G406_0;
	wire G406_fa_;
	wire w_G408_0;
	wire G408_fa_;
	wire w_G410_0;
	wire G410_fa_;
	wire w_G412_0;
	wire G412_fa_;
	wire w_G414_0;
	wire G414_fa_;
	wire w_G416_0;
	wire G416_fa_;
	wire[1:0] w_n345_0;
	wire[1:0] w_n349_0;
	wire[2:0] w_n353_0;
	wire[2:0] w_n354_0;
	wire[2:0] w_n354_1;
	wire[2:0] w_n355_0;
	wire[2:0] w_n355_1;
	wire[2:0] w_n355_2;
	wire[2:0] w_n355_3;
	wire[2:0] w_n355_4;
	wire[2:0] w_n355_5;
	wire[2:0] w_n355_6;
	wire[2:0] w_n355_7;
	wire[2:0] w_n355_8;
	wire[2:0] w_n355_9;
	wire[2:0] w_n355_10;
	wire[2:0] w_n355_11;
	wire[2:0] w_n355_12;
	wire[2:0] w_n355_13;
	wire[2:0] w_n355_14;
	wire[2:0] w_n355_15;
	wire[2:0] w_n355_16;
	wire[2:0] w_n355_17;
	wire[2:0] w_n355_18;
	wire[2:0] w_n355_19;
	wire[2:0] w_n355_20;
	wire[2:0] w_n355_21;
	wire[2:0] w_n355_22;
	wire[2:0] w_n355_23;
	wire[2:0] w_n355_24;
	wire[2:0] w_n355_25;
	wire[1:0] w_n355_26;
	wire[2:0] w_n356_0;
	wire[1:0] w_n358_0;
	wire[1:0] w_n359_0;
	wire[2:0] w_n362_0;
	wire[1:0] w_n364_0;
	wire[1:0] w_n365_0;
	wire[1:0] w_n366_0;
	wire[1:0] w_n370_0;
	wire[2:0] w_n371_0;
	wire[1:0] w_n371_1;
	wire[2:0] w_n372_0;
	wire[2:0] w_n372_1;
	wire[1:0] w_n376_0;
	wire[2:0] w_n377_0;
	wire[2:0] w_n377_1;
	wire[2:0] w_n379_0;
	wire[1:0] w_n379_1;
	wire[2:0] w_n380_0;
	wire[1:0] w_n385_0;
	wire[2:0] w_n386_0;
	wire[2:0] w_n387_0;
	wire[2:0] w_n387_1;
	wire[2:0] w_n388_0;
	wire[1:0] w_n389_0;
	wire[2:0] w_n390_0;
	wire[1:0] w_n390_1;
	wire[2:0] w_n395_0;
	wire[1:0] w_n400_0;
	wire[2:0] w_n401_0;
	wire[2:0] w_n401_1;
	wire[2:0] w_n402_0;
	wire[1:0] w_n402_1;
	wire[1:0] w_n403_0;
	wire[1:0] w_n404_0;
	wire[2:0] w_n405_0;
	wire[2:0] w_n407_0;
	wire[1:0] w_n408_0;
	wire[1:0] w_n410_0;
	wire[2:0] w_n412_0;
	wire[2:0] w_n413_0;
	wire[1:0] w_n413_1;
	wire[2:0] w_n417_0;
	wire[1:0] w_n419_0;
	wire[2:0] w_n422_0;
	wire[2:0] w_n422_1;
	wire[1:0] w_n427_0;
	wire[2:0] w_n428_0;
	wire[2:0] w_n429_0;
	wire[2:0] w_n429_1;
	wire[1:0] w_n429_2;
	wire[1:0] w_n430_0;
	wire[1:0] w_n434_0;
	wire[2:0] w_n435_0;
	wire[1:0] w_n435_1;
	wire[1:0] w_n436_0;
	wire[1:0] w_n437_0;
	wire[1:0] w_n441_0;
	wire[2:0] w_n442_0;
	wire[1:0] w_n443_0;
	wire[1:0] w_n445_0;
	wire[2:0] w_n446_0;
	wire[1:0] w_n446_1;
	wire[1:0] w_n448_0;
	wire[2:0] w_n449_0;
	wire[2:0] w_n450_0;
	wire[1:0] w_n452_0;
	wire[1:0] w_n454_0;
	wire[1:0] w_n455_0;
	wire[2:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[2:0] w_n458_0;
	wire[2:0] w_n460_0;
	wire[1:0] w_n461_0;
	wire[2:0] w_n462_0;
	wire[1:0] w_n464_0;
	wire[2:0] w_n465_0;
	wire[1:0] w_n466_0;
	wire[1:0] w_n468_0;
	wire[2:0] w_n469_0;
	wire[1:0] w_n469_1;
	wire[2:0] w_n470_0;
	wire[2:0] w_n471_0;
	wire[1:0] w_n473_0;
	wire[2:0] w_n474_0;
	wire[1:0] w_n474_1;
	wire[2:0] w_n475_0;
	wire[1:0] w_n475_1;
	wire[1:0] w_n477_0;
	wire[1:0] w_n478_0;
	wire[1:0] w_n479_0;
	wire[2:0] w_n480_0;
	wire[1:0] w_n480_1;
	wire[2:0] w_n481_0;
	wire[1:0] w_n482_0;
	wire[1:0] w_n484_0;
	wire[2:0] w_n485_0;
	wire[2:0] w_n486_0;
	wire[1:0] w_n488_0;
	wire[1:0] w_n489_0;
	wire[2:0] w_n490_0;
	wire[2:0] w_n491_0;
	wire[1:0] w_n491_1;
	wire[1:0] w_n493_0;
	wire[1:0] w_n494_0;
	wire[1:0] w_n502_0;
	wire[1:0] w_n503_0;
	wire[1:0] w_n505_0;
	wire[2:0] w_n507_0;
	wire[2:0] w_n507_1;
	wire[1:0] w_n508_0;
	wire[1:0] w_n509_0;
	wire[1:0] w_n510_0;
	wire[1:0] w_n512_0;
	wire[2:0] w_n514_0;
	wire[2:0] w_n516_0;
	wire[1:0] w_n518_0;
	wire[1:0] w_n519_0;
	wire[2:0] w_n520_0;
	wire[1:0] w_n522_0;
	wire[2:0] w_n523_0;
	wire[2:0] w_n524_0;
	wire[2:0] w_n524_1;
	wire[1:0] w_n524_2;
	wire[2:0] w_n525_0;
	wire[1:0] w_n527_0;
	wire[2:0] w_n528_0;
	wire[1:0] w_n528_1;
	wire[1:0] w_n529_0;
	wire[1:0] w_n530_0;
	wire[2:0] w_n531_0;
	wire[1:0] w_n533_0;
	wire[2:0] w_n534_0;
	wire[1:0] w_n534_1;
	wire[2:0] w_n535_0;
	wire[1:0] w_n535_1;
	wire[1:0] w_n536_0;
	wire[1:0] w_n538_0;
	wire[2:0] w_n539_0;
	wire[1:0] w_n539_1;
	wire[2:0] w_n540_0;
	wire[1:0] w_n542_0;
	wire[1:0] w_n549_0;
	wire[1:0] w_n551_0;
	wire[1:0] w_n552_0;
	wire[1:0] w_n553_0;
	wire[2:0] w_n554_0;
	wire[2:0] w_n556_0;
	wire[1:0] w_n557_0;
	wire[2:0] w_n558_0;
	wire[1:0] w_n560_0;
	wire[2:0] w_n562_0;
	wire[1:0] w_n563_0;
	wire[2:0] w_n564_0;
	wire[2:0] w_n565_0;
	wire[2:0] w_n565_1;
	wire[2:0] w_n565_2;
	wire[2:0] w_n565_3;
	wire[2:0] w_n565_4;
	wire[2:0] w_n565_5;
	wire[2:0] w_n565_6;
	wire[2:0] w_n565_7;
	wire[2:0] w_n565_8;
	wire[2:0] w_n565_9;
	wire[1:0] w_n565_10;
	wire[2:0] w_n567_0;
	wire[1:0] w_n567_1;
	wire[2:0] w_n568_0;
	wire[2:0] w_n569_0;
	wire[1:0] w_n570_0;
	wire[2:0] w_n572_0;
	wire[1:0] w_n572_1;
	wire[2:0] w_n573_0;
	wire[1:0] w_n573_1;
	wire[1:0] w_n574_0;
	wire[1:0] w_n575_0;
	wire[2:0] w_n577_0;
	wire[2:0] w_n578_0;
	wire[1:0] w_n578_1;
	wire[2:0] w_n579_0;
	wire[1:0] w_n580_0;
	wire[1:0] w_n581_0;
	wire[2:0] w_n583_0;
	wire[1:0] w_n583_1;
	wire[2:0] w_n584_0;
	wire[1:0] w_n585_0;
	wire[1:0] w_n586_0;
	wire[2:0] w_n588_0;
	wire[1:0] w_n588_1;
	wire[2:0] w_n589_0;
	wire[1:0] w_n589_1;
	wire[1:0] w_n591_0;
	wire[1:0] w_n592_0;
	wire[1:0] w_n599_0;
	wire[1:0] w_n605_0;
	wire[2:0] w_n606_0;
	wire[2:0] w_n606_1;
	wire[1:0] w_n607_0;
	wire[2:0] w_n608_0;
	wire[1:0] w_n610_0;
	wire[1:0] w_n612_0;
	wire[2:0] w_n613_0;
	wire[2:0] w_n615_0;
	wire[1:0] w_n615_1;
	wire[1:0] w_n617_0;
	wire[2:0] w_n618_0;
	wire[1:0] w_n619_0;
	wire[1:0] w_n620_0;
	wire[2:0] w_n621_0;
	wire[2:0] w_n622_0;
	wire[1:0] w_n622_1;
	wire[2:0] w_n623_0;
	wire[1:0] w_n624_0;
	wire[2:0] w_n625_0;
	wire[1:0] w_n626_0;
	wire[1:0] w_n627_0;
	wire[1:0] w_n628_0;
	wire[1:0] w_n629_0;
	wire[2:0] w_n630_0;
	wire[1:0] w_n631_0;
	wire[1:0] w_n632_0;
	wire[1:0] w_n633_0;
	wire[2:0] w_n634_0;
	wire[2:0] w_n635_0;
	wire[1:0] w_n637_0;
	wire[1:0] w_n642_0;
	wire[1:0] w_n643_0;
	wire[2:0] w_n645_0;
	wire[1:0] w_n647_0;
	wire[2:0] w_n648_0;
	wire[1:0] w_n649_0;
	wire[1:0] w_n650_0;
	wire[1:0] w_n652_0;
	wire[2:0] w_n653_0;
	wire[1:0] w_n653_1;
	wire[1:0] w_n656_0;
	wire[2:0] w_n657_0;
	wire[1:0] w_n657_1;
	wire[2:0] w_n658_0;
	wire[1:0] w_n659_0;
	wire[2:0] w_n660_0;
	wire[1:0] w_n660_1;
	wire[1:0] w_n661_0;
	wire[2:0] w_n662_0;
	wire[1:0] w_n663_0;
	wire[2:0] w_n664_0;
	wire[1:0] w_n664_1;
	wire[2:0] w_n665_0;
	wire[1:0] w_n666_0;
	wire[1:0] w_n667_0;
	wire[2:0] w_n668_0;
	wire[2:0] w_n669_0;
	wire[1:0] w_n671_0;
	wire[1:0] w_n672_0;
	wire[2:0] w_n673_0;
	wire[2:0] w_n674_0;
	wire[1:0] w_n674_1;
	wire[2:0] w_n675_0;
	wire[1:0] w_n676_0;
	wire[2:0] w_n677_0;
	wire[2:0] w_n678_0;
	wire[2:0] w_n679_0;
	wire[1:0] w_n679_1;
	wire[1:0] w_n680_0;
	wire[1:0] w_n683_0;
	wire[1:0] w_n686_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n692_0;
	wire[1:0] w_n693_0;
	wire[2:0] w_n697_0;
	wire[2:0] w_n699_0;
	wire[1:0] w_n699_1;
	wire[2:0] w_n701_0;
	wire[1:0] w_n701_1;
	wire[1:0] w_n703_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n705_0;
	wire[2:0] w_n707_0;
	wire[1:0] w_n708_0;
	wire[2:0] w_n709_0;
	wire[1:0] w_n709_1;
	wire[1:0] w_n710_0;
	wire[1:0] w_n711_0;
	wire[1:0] w_n712_0;
	wire[2:0] w_n713_0;
	wire[1:0] w_n713_1;
	wire[1:0] w_n714_0;
	wire[2:0] w_n715_0;
	wire[2:0] w_n716_0;
	wire[1:0] w_n716_1;
	wire[2:0] w_n720_0;
	wire[1:0] w_n720_1;
	wire[2:0] w_n723_0;
	wire[2:0] w_n727_0;
	wire[1:0] w_n728_0;
	wire[2:0] w_n730_0;
	wire[2:0] w_n734_0;
	wire[1:0] w_n735_0;
	wire[2:0] w_n737_0;
	wire[2:0] w_n741_0;
	wire[1:0] w_n742_0;
	wire[2:0] w_n744_0;
	wire[2:0] w_n748_0;
	wire[1:0] w_n751_0;
	wire[1:0] w_n752_0;
	wire[2:0] w_n754_0;
	wire[2:0] w_n758_0;
	wire[1:0] w_n759_0;
	wire[1:0] w_n764_0;
	wire[1:0] w_n765_0;
	wire[1:0] w_n782_0;
	wire[2:0] w_n784_0;
	wire[2:0] w_n787_0;
	wire[2:0] w_n790_0;
	wire[1:0] w_n790_1;
	wire[2:0] w_n793_0;
	wire[1:0] w_n793_1;
	wire[1:0] w_n795_0;
	wire[2:0] w_n797_0;
	wire[1:0] w_n797_1;
	wire[2:0] w_n801_0;
	wire[1:0] w_n801_1;
	wire[1:0] w_n802_0;
	wire[2:0] w_n804_0;
	wire[2:0] w_n807_0;
	wire[2:0] w_n810_0;
	wire[2:0] w_n812_0;
	wire[2:0] w_n816_0;
	wire[1:0] w_n817_0;
	wire[2:0] w_n819_0;
	wire[2:0] w_n823_0;
	wire[1:0] w_n824_0;
	wire[2:0] w_n827_0;
	wire[2:0] w_n831_0;
	wire[1:0] w_n832_0;
	wire[1:0] w_n834_0;
	wire[1:0] w_n838_0;
	wire[2:0] w_n843_0;
	wire[2:0] w_n847_0;
	wire[1:0] w_n848_0;
	wire[2:0] w_n851_0;
	wire[2:0] w_n855_0;
	wire[1:0] w_n856_0;
	wire[2:0] w_n858_0;
	wire[1:0] w_n859_0;
	wire[1:0] w_n864_0;
	wire[1:0] w_n865_0;
	wire[2:0] w_n869_0;
	wire[2:0] w_n873_0;
	wire[1:0] w_n874_0;
	wire[2:0] w_n878_0;
	wire[2:0] w_n882_0;
	wire[1:0] w_n885_0;
	wire[1:0] w_n887_0;
	wire[1:0] w_n889_0;
	wire[2:0] w_n891_0;
	wire[1:0] w_n891_1;
	wire[2:0] w_n895_0;
	wire[1:0] w_n895_1;
	wire[1:0] w_n896_0;
	wire[2:0] w_n899_0;
	wire[2:0] w_n902_0;
	wire[2:0] w_n905_0;
	wire[2:0] w_n908_0;
	wire[2:0] w_n912_0;
	wire[1:0] w_n913_0;
	wire[2:0] w_n916_0;
	wire[2:0] w_n920_0;
	wire[1:0] w_n921_0;
	wire[1:0] w_n923_0;
	wire[2:0] w_n927_0;
	wire[2:0] w_n931_0;
	wire[1:0] w_n932_0;
	wire[1:0] w_n935_0;
	wire[1:0] w_n937_0;
	wire[1:0] w_n939_0;
	wire[2:0] w_n945_0;
	wire[1:0] w_n945_1;
	wire[2:0] w_n948_0;
	wire[1:0] w_n948_1;
	wire[1:0] w_n950_0;
	wire[1:0] w_n952_0;
	wire[1:0] w_n957_0;
	wire[1:0] w_n972_0;
	wire[1:0] w_n981_0;
	wire[1:0] w_n987_0;
	wire[2:0] w_n988_0;
	wire[2:0] w_n992_0;
	wire[1:0] w_n993_0;
	wire[1:0] w_n994_0;
	wire[2:0] w_n995_0;
	wire[2:0] w_n999_0;
	wire[1:0] w_n1000_0;
	wire[1:0] w_n1003_0;
	wire[1:0] w_n1007_0;
	wire[1:0] w_n1008_0;
	wire[2:0] w_n1009_0;
	wire[1:0] w_n1009_1;
	wire[2:0] w_n1013_0;
	wire[1:0] w_n1013_1;
	wire[1:0] w_n1014_0;
	wire[1:0] w_n1015_0;
	wire[2:0] w_n1016_0;
	wire[2:0] w_n1019_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1044_0;
	wire[2:0] w_n1061_0;
	wire[1:0] w_n1062_0;
	wire[2:0] w_n1066_0;
	wire[1:0] w_n1068_0;
	wire[1:0] w_n1069_0;
	wire[2:0] w_n1073_0;
	wire[1:0] w_n1075_0;
	wire[1:0] w_n1076_0;
	wire[2:0] w_n1077_0;
	wire[2:0] w_n1081_0;
	wire[1:0] w_n1082_0;
	wire[2:0] w_n1086_0;
	wire[1:0] w_n1092_0;
	wire[1:0] w_n1095_0;
	wire[2:0] w_n1096_0;
	wire[2:0] w_n1100_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1104_0;
	wire[1:0] w_n1105_0;
	wire[1:0] w_n1116_0;
	wire[2:0] w_n1122_0;
	wire[2:0] w_n1125_0;
	wire[1:0] w_n1127_0;
	wire[2:0] w_n1128_0;
	wire[1:0] w_n1128_1;
	wire[1:0] w_n1130_0;
	wire[1:0] w_n1136_0;
	wire[1:0] w_n1142_0;
	wire[2:0] w_n1148_0;
	wire[1:0] w_n1156_0;
	wire[1:0] w_n1166_0;
	wire[1:0] w_n1173_0;
	wire[1:0] w_n1189_0;
	wire[1:0] w_n1205_0;
	wire[1:0] w_n1236_0;
	wire[1:0] w_n1244_0;
	wire[1:0] w_n1283_0;
	wire[1:0] w_n1301_0;
	wire[1:0] w_n1309_0;
	wire[1:0] w_n1317_0;
	wire[1:0] w_n1325_0;
	wire[2:0] w_n1359_0;
	wire[2:0] w_n1360_0;
	wire[1:0] w_n1360_1;
	wire[1:0] w_n1361_0;
	wire[1:0] w_n1362_0;
	wire[1:0] w_n1376_0;
	wire[2:0] w_n1380_0;
	wire[1:0] w_n1380_1;
	wire[2:0] w_n1383_0;
	wire[2:0] w_n1383_1;
	wire[2:0] w_n1385_0;
	wire[1:0] w_n1385_1;
	wire[2:0] w_n1389_0;
	wire[1:0] w_n1389_1;
	wire[2:0] w_n1392_0;
	wire[1:0] w_n1392_1;
	wire[1:0] w_n1401_0;
	wire[1:0] w_n1402_0;
	wire[1:0] w_n1403_0;
	wire[1:0] w_n1404_0;
	wire[1:0] w_n1405_0;
	wire[1:0] w_n1406_0;
	wire[1:0] w_n1414_0;
	wire[2:0] w_n1420_0;
	wire[1:0] w_n1421_0;
	wire[1:0] w_n1422_0;
	wire[1:0] w_n1424_0;
	wire[1:0] w_n1425_0;
	wire[2:0] w_n1444_0;
	wire[1:0] w_n1445_0;
	wire[1:0] w_n1447_0;
	wire[1:0] w_n1454_0;
	wire[2:0] w_n1463_0;
	wire[1:0] w_n1464_0;
	wire[1:0] w_n1465_0;
	wire[1:0] w_n1468_0;
	wire[1:0] w_n1469_0;
	wire[1:0] w_n1470_0;
	wire[1:0] w_n1471_0;
	wire[1:0] w_n1472_0;
	wire[1:0] w_n1473_0;
	wire[1:0] w_n1479_0;
	wire[1:0] w_n1482_0;
	wire[1:0] w_n1486_0;
	wire[2:0] w_n1494_0;
	wire[1:0] w_n1501_0;
	wire[1:0] w_n1510_0;
	wire[1:0] w_n1520_0;
	wire[1:0] w_n1536_0;
	wire[1:0] w_n1571_0;
	wire[1:0] w_n1599_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1611_0;
	wire[1:0] w_n1625_0;
	wire[1:0] w_n1642_0;
	wire[1:0] w_n1644_0;
	wire[1:0] w_n1651_0;
	wire[1:0] w_n1654_0;
	wire[1:0] w_n1659_0;
	wire[1:0] w_n1667_0;
	wire[1:0] w_n1670_0;
	wire[1:0] w_n1672_0;
	wire[1:0] w_n1675_0;
	wire[1:0] w_n1680_0;
	wire[1:0] w_n1687_0;
	wire[1:0] w_n1689_0;
	wire[1:0] w_n1699_0;
	wire w_dff_A_9QO5kMsf6_0;
	wire w_dff_A_7yeiBPBK4_0;
	wire w_dff_A_UczSuiSW2_1;
	wire w_dff_A_J3enjoPb9_1;
	wire w_dff_A_nZ0M8cl96_1;
	wire w_dff_A_trt7Zdp61_2;
	wire w_dff_B_FzU78smc9_3;
	wire w_dff_B_QKk2GhSn2_3;
	wire w_dff_B_98XYDJw71_3;
	wire w_dff_B_1hi48cLb9_3;
	wire w_dff_B_0O7tdvpT7_3;
	wire w_dff_B_RlafvuDv0_3;
	wire w_dff_B_c7nUrlS48_3;
	wire w_dff_B_qVGDMjuk5_3;
	wire w_dff_B_l8esVTko5_3;
	wire w_dff_B_gIskj6br3_3;
	wire w_dff_B_HYZgzBaJ0_3;
	wire w_dff_B_Jyrb7Aq96_3;
	wire w_dff_B_7CCFwbtG6_3;
	wire w_dff_B_wwddzhuJ8_3;
	wire w_dff_B_2h7M6AcW9_3;
	wire w_dff_B_9MDYm1pu5_3;
	wire w_dff_B_GEaJHj6j2_0;
	wire w_dff_B_beIsjM3H9_0;
	wire w_dff_B_jYpCtpT52_0;
	wire w_dff_B_3PvZ7pln0_0;
	wire w_dff_B_NzkL4KCy0_0;
	wire w_dff_B_wqq56lm13_0;
	wire w_dff_B_7o9MhInf4_0;
	wire w_dff_A_gWIsP7hv9_0;
	wire w_dff_A_6ENtODDw6_0;
	wire w_dff_A_qE6J2TTm7_0;
	wire w_dff_B_dUmJ2nLu5_3;
	wire w_dff_B_zCbOuQPA0_3;
	wire w_dff_B_ZcdM3jqe8_3;
	wire w_dff_B_FVvdv52x2_3;
	wire w_dff_B_MLds6pbi2_3;
	wire w_dff_B_k3HNFrRD1_3;
	wire w_dff_B_QLKWXMm39_3;
	wire w_dff_B_N6HqhR0y8_3;
	wire w_dff_B_gOHBfbdE9_3;
	wire w_dff_B_yhVRwWBm1_3;
	wire w_dff_B_cxTFjToG5_3;
	wire w_dff_B_qS8OzpVe0_3;
	wire w_dff_B_PoMEaLyb3_3;
	wire w_dff_B_KNTreujU3_3;
	wire w_dff_B_fNpvSgHX4_3;
	wire w_dff_B_p7Uf4fmW9_3;
	wire w_dff_B_ZlWdhG8u9_3;
	wire w_dff_B_WmOCm0RJ3_3;
	wire w_dff_B_805vkh0G7_3;
	wire w_dff_B_t54pZ6mO1_3;
	wire w_dff_B_fBSeNbDi3_3;
	wire w_dff_B_vpIy1vDB9_1;
	wire w_dff_B_1EiMZeuy7_1;
	wire w_dff_B_OCAc2VMT7_1;
	wire w_dff_B_jKZGV9nb8_1;
	wire w_dff_B_D5NeVKLt5_1;
	wire w_dff_B_DbWs0oaN0_1;
	wire w_dff_B_IqtCQLiX5_1;
	wire w_dff_B_IpQODK7f5_1;
	wire w_dff_B_xjehSzm19_1;
	wire w_dff_B_GO6NziZ45_1;
	wire w_dff_B_6CedrUXU4_1;
	wire w_dff_B_HZR9lwyG3_1;
	wire w_dff_B_PqrPMV0z5_1;
	wire w_dff_B_1j8yn1Co1_1;
	wire w_dff_B_fbaVvFO18_1;
	wire w_dff_B_jokLNW1J8_1;
	wire w_dff_B_8iTWyAfu7_1;
	wire w_dff_B_VEBovauy4_1;
	wire w_dff_B_NgxFGKZy6_1;
	wire w_dff_B_yoJOtEfA0_1;
	wire w_dff_B_sa2I5if72_1;
	wire w_dff_B_hWUmrSTw6_1;
	wire w_dff_B_k1hjEaZw6_1;
	wire w_dff_B_kxsOkfov5_1;
	wire w_dff_B_YVoRaUVm1_1;
	wire w_dff_B_unL2ikBW9_1;
	wire w_dff_B_Ul7f0PSX0_1;
	wire w_dff_B_o3urkvCr2_1;
	wire w_dff_B_ZtOmaFTA5_1;
	wire w_dff_B_ZBSCXzLP5_1;
	wire w_dff_B_IcqrIkq40_0;
	wire w_dff_B_Pcx1cnVY3_0;
	wire w_dff_B_mRB84Aq46_0;
	wire w_dff_B_FjQeWa9J1_1;
	wire w_dff_B_4nntlRnQ0_1;
	wire w_dff_B_uf5Db5j67_1;
	wire w_dff_B_wpLSqmpN9_1;
	wire w_dff_B_3YOAXYRg6_1;
	wire w_dff_B_NpqUElue4_1;
	wire w_dff_B_aMRKJmGW8_1;
	wire w_dff_B_4bomZnzS5_1;
	wire w_dff_B_9W3GlZnr3_1;
	wire w_dff_B_bIyzspRH8_1;
	wire w_dff_B_1suRTZFd4_1;
	wire w_dff_B_ixTSlmXd3_1;
	wire w_dff_B_YisDDqVG1_1;
	wire w_dff_B_BfcfbpoJ1_1;
	wire w_dff_B_hedONhuP5_1;
	wire w_dff_B_bEfWGry60_1;
	wire w_dff_B_y7E0SZLh8_1;
	wire w_dff_B_DFsZgEkb6_1;
	wire w_dff_B_r68osuAM6_1;
	wire w_dff_B_PeBK9cnt2_1;
	wire w_dff_B_8PZoI8Si5_1;
	wire w_dff_B_sWOF15J72_1;
	wire w_dff_B_OCC3loJT5_1;
	wire w_dff_B_UuV8fNvE1_1;
	wire w_dff_B_v5I4KI7d8_1;
	wire w_dff_B_vrjz5V6r5_1;
	wire w_dff_B_XHnAdNvx9_1;
	wire w_dff_A_6sApNmgt4_1;
	wire w_dff_A_9ke25cNh8_0;
	wire w_dff_A_LZ0JsTsi0_0;
	wire w_dff_A_2UCs1x1D6_0;
	wire w_dff_A_MC0n00H68_0;
	wire w_dff_A_es7rLjWZ1_0;
	wire w_dff_A_AXC1wYxF0_0;
	wire w_dff_A_3tN9rxVx2_0;
	wire w_dff_A_bR1Dca1U6_0;
	wire w_dff_A_yFlqPns54_0;
	wire w_dff_A_UWLrWuEJ8_0;
	wire w_dff_A_pt1XiaWX8_0;
	wire w_dff_A_mm5g4OxK0_0;
	wire w_dff_A_mlLZNHuO4_0;
	wire w_dff_A_qrcZCWMn1_0;
	wire w_dff_A_2BzIJhw14_0;
	wire w_dff_A_y9h8Fv2q9_0;
	wire w_dff_A_MFr7mmy71_0;
	wire w_dff_A_92nXppBQ8_0;
	wire w_dff_A_Vlr6wKaK1_0;
	wire w_dff_A_QuTrwZn00_0;
	wire w_dff_A_NLUaM75w9_0;
	wire w_dff_A_Tp2fn0a22_0;
	wire w_dff_A_ebvaHMAG2_0;
	wire w_dff_A_iqBvkcJP9_0;
	wire w_dff_A_UjCBY7Yj8_0;
	wire w_dff_A_wiUo5LgO2_0;
	wire w_dff_A_oxIB4Cei6_1;
	wire w_dff_A_KOnG8ukG2_0;
	wire w_dff_A_jh3p7e118_0;
	wire w_dff_A_4lhwOdNW5_0;
	wire w_dff_A_iO6niJPu6_0;
	wire w_dff_A_KnX3nX9b1_0;
	wire w_dff_A_GXzK9WtO3_0;
	wire w_dff_A_WZGcfpE69_0;
	wire w_dff_A_z2YVascr1_0;
	wire w_dff_A_mgsOG2QB8_0;
	wire w_dff_A_jMQ72mdi0_0;
	wire w_dff_A_jbC9VSDC0_0;
	wire w_dff_A_mJAmcchH5_0;
	wire w_dff_A_QHUvUFHM0_0;
	wire w_dff_A_WxDVy1df7_0;
	wire w_dff_A_4YyXivOI6_0;
	wire w_dff_A_hMS5KX0s6_0;
	wire w_dff_A_wasIBB1m9_0;
	wire w_dff_A_AVda3LZ30_0;
	wire w_dff_A_ZAWGvtXM1_0;
	wire w_dff_A_E1S6cTHU0_0;
	wire w_dff_A_PhKk96Qz8_0;
	wire w_dff_A_hQldPRiL2_0;
	wire w_dff_A_5TME2nT46_0;
	wire w_dff_A_PNMpFsm19_0;
	wire w_dff_A_XUoaSZcL4_0;
	wire w_dff_A_5pOQ5Aju4_0;
	wire w_dff_A_10WK5Ss63_1;
	wire w_dff_A_m2OXd8GU0_0;
	wire w_dff_A_RCj1M2n81_0;
	wire w_dff_A_5GzlOVEQ3_0;
	wire w_dff_A_HtgsWHLE0_0;
	wire w_dff_A_wLAdzhAG7_0;
	wire w_dff_A_1FTqlbdL8_0;
	wire w_dff_A_1qKZGVgd2_0;
	wire w_dff_A_mg5a3Dd29_0;
	wire w_dff_A_7xglEOUm7_0;
	wire w_dff_A_IGgBAqn46_0;
	wire w_dff_A_vYWqheHh5_0;
	wire w_dff_A_DdIWD3GI6_0;
	wire w_dff_A_tENZkOfu9_0;
	wire w_dff_A_5rECpUAp8_0;
	wire w_dff_A_ai9ESNxo3_0;
	wire w_dff_A_HPVVcXE57_0;
	wire w_dff_A_2fFXPoYH3_0;
	wire w_dff_A_xs0vf9sa5_0;
	wire w_dff_A_4DCGFR3V4_0;
	wire w_dff_A_1D8OSKsX3_0;
	wire w_dff_A_Wx07uk4D7_0;
	wire w_dff_A_6HNy7nDt6_0;
	wire w_dff_A_rEOCcJTv9_0;
	wire w_dff_A_ocrFkLCU5_0;
	wire w_dff_A_UohQTphH9_0;
	wire w_dff_A_jFIevkki1_0;
	wire w_dff_A_kCaRS6Sy6_1;
	wire w_dff_A_FZW6VcR89_0;
	wire w_dff_A_oVX9haIk8_0;
	wire w_dff_A_rdUe9k8F7_0;
	wire w_dff_A_CAZqmPnc3_0;
	wire w_dff_A_xL6t0IWm9_0;
	wire w_dff_A_JE4n6kCm7_0;
	wire w_dff_A_J9FZsDMu4_0;
	wire w_dff_A_mmmFMqzu3_0;
	wire w_dff_A_NppFIkLE8_0;
	wire w_dff_A_4OarWApE4_0;
	wire w_dff_A_ZuUukkmu1_0;
	wire w_dff_A_QOHK88YV2_0;
	wire w_dff_A_wh25BaB73_0;
	wire w_dff_A_qIvWoEdV6_0;
	wire w_dff_A_TeDyRX4V6_0;
	wire w_dff_A_pEO0k3Wb7_0;
	wire w_dff_A_K2w6pVw00_0;
	wire w_dff_A_cCe9KEAq6_0;
	wire w_dff_A_OgnbogKE4_0;
	wire w_dff_A_z0N22mwn7_0;
	wire w_dff_A_9OXmE5QW8_0;
	wire w_dff_A_tSplufwi4_0;
	wire w_dff_A_jJoz5WTJ6_0;
	wire w_dff_A_WeVAw1Fr1_0;
	wire w_dff_A_xgD2f48o8_0;
	wire w_dff_A_mPJ9Ru6q4_0;
	wire w_dff_A_tz2EUH5g2_1;
	wire w_dff_A_9mG3Lu1n0_0;
	wire w_dff_A_yidHp8eC2_0;
	wire w_dff_A_VzXCQxLY9_0;
	wire w_dff_A_R7HlyTZD5_0;
	wire w_dff_A_nO9k76IR3_0;
	wire w_dff_A_eorpBthw2_0;
	wire w_dff_A_xlEygdER1_0;
	wire w_dff_A_1CxfVFdc6_0;
	wire w_dff_A_Di5cysJZ0_0;
	wire w_dff_A_ks31prln2_0;
	wire w_dff_A_DX9SLhis1_0;
	wire w_dff_A_CY3Dw0K33_0;
	wire w_dff_A_v92hmE3l7_0;
	wire w_dff_A_ew1OSBIm6_0;
	wire w_dff_A_aLXiHK0v8_0;
	wire w_dff_A_GUxv8NP97_0;
	wire w_dff_A_56JtU3Z06_0;
	wire w_dff_A_mEWlNEV93_0;
	wire w_dff_A_uLRusD744_0;
	wire w_dff_A_I9OZLL0H9_0;
	wire w_dff_A_jjejcgTo5_0;
	wire w_dff_A_84PfOtyr1_0;
	wire w_dff_A_vTTYpNhr7_0;
	wire w_dff_A_KdvfegDV5_0;
	wire w_dff_A_iXZXkzMz3_0;
	wire w_dff_A_Ey1u0GRR4_0;
	wire w_dff_A_n6GEbAPE9_1;
	wire w_dff_A_vhSL0ylA8_0;
	wire w_dff_A_vuaj4YVy1_0;
	wire w_dff_A_ouZwcVQa8_0;
	wire w_dff_A_uacfhTVx2_0;
	wire w_dff_A_m98kHR7B0_0;
	wire w_dff_A_scQK8cxc2_0;
	wire w_dff_A_2dNb6GiG8_0;
	wire w_dff_A_kHsCSco35_0;
	wire w_dff_A_gsTwXeFl2_0;
	wire w_dff_A_YgeZsEwQ0_0;
	wire w_dff_A_nKeS3DuD6_0;
	wire w_dff_A_63u1S9YW9_0;
	wire w_dff_A_w9f6qIDK0_0;
	wire w_dff_A_Qk3nP7Dl8_0;
	wire w_dff_A_lRTTKe4K8_0;
	wire w_dff_A_RoPD4Z1f3_0;
	wire w_dff_A_dDsFKOM42_0;
	wire w_dff_A_m2JKHjhT5_0;
	wire w_dff_A_IozIKX6i6_0;
	wire w_dff_A_LnbujqxW7_0;
	wire w_dff_A_OruZdeSh4_0;
	wire w_dff_A_lJltIt2F9_0;
	wire w_dff_A_0J1PsqUz8_0;
	wire w_dff_A_TvVmRDFc7_0;
	wire w_dff_A_M6XVcSha7_0;
	wire w_dff_A_30PmYXmR9_0;
	wire w_dff_A_eZCLFuLa4_1;
	wire w_dff_A_OHMTBp7v4_0;
	wire w_dff_A_2WqyOJTU7_0;
	wire w_dff_A_hV1p6eWM3_0;
	wire w_dff_A_gz2Ewt9K0_0;
	wire w_dff_A_HYR6Vitj0_0;
	wire w_dff_A_lL1Njcps1_0;
	wire w_dff_A_TQQ8cuz43_0;
	wire w_dff_A_xP5lZ3ko5_0;
	wire w_dff_A_GaKABU4J6_0;
	wire w_dff_A_E5uWkL2w0_0;
	wire w_dff_A_QtjBnO1x7_0;
	wire w_dff_A_D3YpL1SM3_0;
	wire w_dff_A_s7s0FuBn6_0;
	wire w_dff_A_olkoY8rg5_0;
	wire w_dff_A_mP9VXzn46_0;
	wire w_dff_A_uUU6biFu6_0;
	wire w_dff_A_AY5aMxLv5_0;
	wire w_dff_A_kcvpou7C5_0;
	wire w_dff_A_sYxXon2S1_0;
	wire w_dff_A_CwLKBqSc5_0;
	wire w_dff_A_8Zpj7t9g1_0;
	wire w_dff_A_rPs7T8ai0_0;
	wire w_dff_A_yZRROB5r1_0;
	wire w_dff_A_hBWYzKIH4_0;
	wire w_dff_A_1fOOLZ0z6_0;
	wire w_dff_A_FVnoGUp58_0;
	wire w_dff_A_7VdHePjq5_1;
	wire w_dff_A_eLwjgnpG0_0;
	wire w_dff_A_NV3ofKnU2_0;
	wire w_dff_A_r6ZTE5W39_0;
	wire w_dff_A_LXc8bHfA0_0;
	wire w_dff_A_2xkbbBgt0_0;
	wire w_dff_A_hW0Jx9WF0_0;
	wire w_dff_A_Y74ITYZM9_0;
	wire w_dff_A_JYT21bjO0_0;
	wire w_dff_A_DByppb385_0;
	wire w_dff_A_oysh2A488_0;
	wire w_dff_A_jgjOjtK23_0;
	wire w_dff_A_3Xy3xQz45_0;
	wire w_dff_A_dtY1ZSAz4_0;
	wire w_dff_A_47B6qsAS5_0;
	wire w_dff_A_dpBByX4E1_0;
	wire w_dff_A_nTUDBs2i7_0;
	wire w_dff_A_sz9DWv3j3_0;
	wire w_dff_A_AbspSUIb2_0;
	wire w_dff_A_funZxtua1_0;
	wire w_dff_A_Z1Fvwk8Q9_0;
	wire w_dff_A_Xi1zp94q0_0;
	wire w_dff_A_m8bmpBbW6_0;
	wire w_dff_A_xSjSqwBd2_0;
	wire w_dff_A_IHoLcdss3_0;
	wire w_dff_A_jz5NWKKy7_0;
	wire w_dff_A_bqWqExrP5_0;
	wire w_dff_A_l63WIzjM6_1;
	wire w_dff_A_erv3MoCl6_0;
	wire w_dff_A_23Nzfjzz4_0;
	wire w_dff_A_hDA8oJ3Z7_0;
	wire w_dff_A_Si5JKb6B2_0;
	wire w_dff_A_1GH6aFFI7_0;
	wire w_dff_A_MRMohy7L5_0;
	wire w_dff_A_XIIBFOiR3_0;
	wire w_dff_A_PSGM1cWS1_0;
	wire w_dff_A_ZQnpKyJs9_0;
	wire w_dff_A_WjTic5P82_0;
	wire w_dff_A_ZkwKTgP03_0;
	wire w_dff_A_akfZ5Bak4_0;
	wire w_dff_A_wFHvd1Lq0_0;
	wire w_dff_A_cpEe7gY65_0;
	wire w_dff_A_tpmFTXUA6_0;
	wire w_dff_A_U2CRmF4K1_0;
	wire w_dff_A_WG28kDGY7_0;
	wire w_dff_A_01xXUPsM1_0;
	wire w_dff_A_TIL8YHkX0_0;
	wire w_dff_A_CU1mMcyK6_0;
	wire w_dff_A_2yxsluPl9_0;
	wire w_dff_A_KtuYRaNB8_0;
	wire w_dff_A_7ddChlGP8_0;
	wire w_dff_A_iTrwKClE9_0;
	wire w_dff_A_hRSgFL8V2_0;
	wire w_dff_A_jAg8ipek3_0;
	wire w_dff_A_38SOXGaA5_1;
	wire w_dff_A_KeiJ0RtT9_0;
	wire w_dff_A_QgRBCdsL6_0;
	wire w_dff_A_VRFKqh112_0;
	wire w_dff_A_3mv3czMj9_0;
	wire w_dff_A_uXxTkFel7_0;
	wire w_dff_A_95MWKwuz3_0;
	wire w_dff_A_NI4HY9Il8_0;
	wire w_dff_A_jcH6biH79_0;
	wire w_dff_A_S9yFVrOo8_0;
	wire w_dff_A_oawsxvSq5_0;
	wire w_dff_A_c60nqKA02_0;
	wire w_dff_A_vh672oYT7_0;
	wire w_dff_A_ubt47kOw0_0;
	wire w_dff_A_QG4AoQJX8_0;
	wire w_dff_A_q4MuepBg4_0;
	wire w_dff_A_trZDxp1t2_0;
	wire w_dff_A_5cCi84ZB8_0;
	wire w_dff_A_N74xfBax7_0;
	wire w_dff_A_e6ywPm164_0;
	wire w_dff_A_fWhcDEEt4_0;
	wire w_dff_A_jHUD2lfR3_0;
	wire w_dff_A_rNKzjgPj4_0;
	wire w_dff_A_WCVQz6gw3_0;
	wire w_dff_A_jhG2YlK52_0;
	wire w_dff_A_yVL49AWJ9_0;
	wire w_dff_A_d1yeIUe78_0;
	wire w_dff_A_SUaMaM1Z9_1;
	wire w_dff_A_RfFlRvc98_0;
	wire w_dff_A_ATamxKvN4_0;
	wire w_dff_A_kG7ZOa896_0;
	wire w_dff_A_eIOSNxwP7_0;
	wire w_dff_A_wkL8Ws237_0;
	wire w_dff_A_VfyBSNvD5_0;
	wire w_dff_A_IPkdxN7Y4_0;
	wire w_dff_A_SipErOe39_0;
	wire w_dff_A_I6XeDiTP7_0;
	wire w_dff_A_UzAQnEMN2_0;
	wire w_dff_A_GVTsDNjh6_0;
	wire w_dff_A_tr5CDcJb0_0;
	wire w_dff_A_56d2YEf73_0;
	wire w_dff_A_0zFHMc236_0;
	wire w_dff_A_2dRy7EHp1_0;
	wire w_dff_A_GLVV54ps2_0;
	wire w_dff_A_jyWGfFm48_0;
	wire w_dff_A_0lk96sWg8_0;
	wire w_dff_A_CySS9Psy9_0;
	wire w_dff_A_v0zKxZPp7_0;
	wire w_dff_A_KZO5bQBU7_0;
	wire w_dff_A_XjBCg3ig5_0;
	wire w_dff_A_NSg3Al6P0_0;
	wire w_dff_A_Adf9uIwU5_0;
	wire w_dff_A_Jjl2wtTR6_0;
	wire w_dff_A_riKnTTVZ4_0;
	wire w_dff_A_3ZgZBMkC9_1;
	wire w_dff_A_IZ5PZk5T1_0;
	wire w_dff_A_KKDlyxGu6_0;
	wire w_dff_A_DUJFvNjE8_0;
	wire w_dff_A_RmTNuhnG8_0;
	wire w_dff_A_SpJoU5tG4_0;
	wire w_dff_A_btUjeE8P2_0;
	wire w_dff_A_iOBp8yYX0_0;
	wire w_dff_A_HGBZ4CNf7_0;
	wire w_dff_A_4UhJp8bi9_0;
	wire w_dff_A_TEl1bOVV8_0;
	wire w_dff_A_Za8Jvuu72_0;
	wire w_dff_A_lhHcrvbB1_0;
	wire w_dff_A_FsEdFg1w7_0;
	wire w_dff_A_B4UEwavN3_0;
	wire w_dff_A_aFdxKZoe1_0;
	wire w_dff_A_FTyiYmxU8_0;
	wire w_dff_A_Rk8kZTiQ8_0;
	wire w_dff_A_OqeN6mxq4_0;
	wire w_dff_A_jctkx6nM4_0;
	wire w_dff_A_RUqYA2zh8_0;
	wire w_dff_A_lqltRERL4_0;
	wire w_dff_A_GLEcxDyd1_0;
	wire w_dff_A_kDxnzNc71_0;
	wire w_dff_A_biqjCc5w0_0;
	wire w_dff_A_Po3bXLZ27_0;
	wire w_dff_A_NP0CdFxh6_0;
	wire w_dff_A_inOpBq5G8_1;
	wire w_dff_A_039U8Q8C1_0;
	wire w_dff_A_PTp0ta9f6_0;
	wire w_dff_A_g708R9XT0_0;
	wire w_dff_A_t3Yp2unN1_0;
	wire w_dff_A_OXpDVo2H8_0;
	wire w_dff_A_sSmWuDKB1_0;
	wire w_dff_A_UKCzLuto4_0;
	wire w_dff_A_NXv5T3ya3_0;
	wire w_dff_A_CAUnL9Al1_0;
	wire w_dff_A_cIcFij5p5_0;
	wire w_dff_A_Ilymf3k60_0;
	wire w_dff_A_8qrfBtfI6_0;
	wire w_dff_A_6SJqKCvb9_0;
	wire w_dff_A_3m0wo6jv8_0;
	wire w_dff_A_yOuD4OE66_0;
	wire w_dff_A_TNs3vqNj5_0;
	wire w_dff_A_LZCfvpDu8_0;
	wire w_dff_A_pSsy8Hzz1_0;
	wire w_dff_A_V89V8Nw91_0;
	wire w_dff_A_zqLwOlIH9_0;
	wire w_dff_A_PXP0deGy6_0;
	wire w_dff_A_yf5cjXBT9_0;
	wire w_dff_A_TLyJCJ7a6_0;
	wire w_dff_A_dMl85Xx90_0;
	wire w_dff_A_8ghSo01x1_0;
	wire w_dff_A_BAVH7tD56_0;
	wire w_dff_A_hlARsFhN7_1;
	wire w_dff_A_SgpPuK3k2_0;
	wire w_dff_A_kIS6r4aZ7_0;
	wire w_dff_A_j1uevwda9_0;
	wire w_dff_A_ulUrA0lV6_0;
	wire w_dff_A_4DfMWjq31_0;
	wire w_dff_A_OuPm1V7O1_0;
	wire w_dff_A_RBfYFazA8_0;
	wire w_dff_A_akxtPTHv4_0;
	wire w_dff_A_m4lMHFXj6_0;
	wire w_dff_A_dmLDFLKy4_0;
	wire w_dff_A_CXZm86Ph2_0;
	wire w_dff_A_wNhqRwne3_0;
	wire w_dff_A_CoksQ7oJ2_0;
	wire w_dff_A_EHcs4mm87_0;
	wire w_dff_A_d0FflE2i1_0;
	wire w_dff_A_osMKI9VY2_0;
	wire w_dff_A_ZsRbECSD5_0;
	wire w_dff_A_srEJcsCX5_0;
	wire w_dff_A_bA9m6G8e2_0;
	wire w_dff_A_3vMVWMoP0_0;
	wire w_dff_A_vU82p77L9_0;
	wire w_dff_A_WY6hktmd5_0;
	wire w_dff_A_LN2CD0su7_0;
	wire w_dff_A_173W7EVh5_0;
	wire w_dff_A_zgz1NpSK5_0;
	wire w_dff_A_zcFDXErM4_0;
	wire w_dff_A_Yw7VDQLa0_1;
	wire w_dff_A_fFw0wmn91_0;
	wire w_dff_A_lJ6ZBqqG7_0;
	wire w_dff_A_kvUmlWvO0_0;
	wire w_dff_A_2hff1qmi7_0;
	wire w_dff_A_xvfhuQGx0_0;
	wire w_dff_A_wIoYfbUU9_0;
	wire w_dff_A_BZdaZaar2_0;
	wire w_dff_A_6EWU5u2h8_0;
	wire w_dff_A_cFMAwVlX6_0;
	wire w_dff_A_kA0hsreO0_0;
	wire w_dff_A_eA4MY8kK1_0;
	wire w_dff_A_sO5rbTRb9_0;
	wire w_dff_A_dciytgMa1_0;
	wire w_dff_A_58Xol0Np8_0;
	wire w_dff_A_NIDDf4Uc5_0;
	wire w_dff_A_arZCFY215_0;
	wire w_dff_A_sOaTfcIY3_0;
	wire w_dff_A_qnPdfFKy6_0;
	wire w_dff_A_xFVdJ6F87_0;
	wire w_dff_A_pAjtyoiV0_0;
	wire w_dff_A_l4uHRBEq2_0;
	wire w_dff_A_eNfHrf2X2_0;
	wire w_dff_A_DAxIzlkR2_0;
	wire w_dff_A_FUjRZ8cJ9_0;
	wire w_dff_A_m8DC2qn42_0;
	wire w_dff_A_z06FxRP62_0;
	wire w_dff_A_iwHRIdkG4_1;
	wire w_dff_A_BGIFbOyj3_0;
	wire w_dff_A_shiOtPBA1_0;
	wire w_dff_A_yQ1frlMq0_0;
	wire w_dff_A_QjrkGQnj0_0;
	wire w_dff_A_VjBlEaz29_0;
	wire w_dff_A_XKRGadRE7_0;
	wire w_dff_A_PuRnX3BE1_0;
	wire w_dff_A_TpKsZdyo3_0;
	wire w_dff_A_hNASR3aM1_0;
	wire w_dff_A_VgJ6n0pj0_0;
	wire w_dff_A_6ho07pFh3_0;
	wire w_dff_A_3jgQ4y4P6_0;
	wire w_dff_A_4yPJU22y0_0;
	wire w_dff_A_tR7DVRlK5_0;
	wire w_dff_A_VCW5Ns853_0;
	wire w_dff_A_z1DAj4V71_0;
	wire w_dff_A_7taAytV31_0;
	wire w_dff_A_SriZSmBP0_0;
	wire w_dff_A_1Jb8n4hz9_0;
	wire w_dff_A_1Xt1UsRl3_0;
	wire w_dff_A_intqS4js7_0;
	wire w_dff_A_k5KwYpQi1_0;
	wire w_dff_A_gmh3UkLG7_0;
	wire w_dff_A_ppx1SayD0_0;
	wire w_dff_A_elGRqeP33_0;
	wire w_dff_A_De9jW90n8_0;
	wire w_dff_A_C0nNn7ci4_1;
	wire w_dff_A_kUPu9xz88_0;
	wire w_dff_A_nTUQs7fh3_0;
	wire w_dff_A_menA27iF4_0;
	wire w_dff_A_Rcnqp6fB2_0;
	wire w_dff_A_ztQaC30v6_0;
	wire w_dff_A_PyRfqxRy5_0;
	wire w_dff_A_Na6L0eqI3_0;
	wire w_dff_A_YUikfB001_0;
	wire w_dff_A_wIpC1jAw5_0;
	wire w_dff_A_iL6rTm147_0;
	wire w_dff_A_RG42v5Fo8_0;
	wire w_dff_A_sPq86jLW4_0;
	wire w_dff_A_YHmzYt8i1_0;
	wire w_dff_A_4OxsawFZ3_0;
	wire w_dff_A_JnSSaOBu9_0;
	wire w_dff_A_kRPMbu3g4_0;
	wire w_dff_A_HUWUs3gN8_0;
	wire w_dff_A_OUZKb1xo5_0;
	wire w_dff_A_9e2NgsCI6_0;
	wire w_dff_A_FsJOpsmq4_0;
	wire w_dff_A_C1xQKPcp3_0;
	wire w_dff_A_SfHDnweU7_0;
	wire w_dff_A_U4Ve1heT3_0;
	wire w_dff_A_Mx8z8elo3_0;
	wire w_dff_A_gUPOrKao8_0;
	wire w_dff_A_Jwe6IFZW0_0;
	wire w_dff_A_d6GEvmtG3_1;
	wire w_dff_A_jatncqTv3_0;
	wire w_dff_A_ZKRR7VyO6_0;
	wire w_dff_A_Dws1yAcj2_0;
	wire w_dff_A_I4b9DIGF2_0;
	wire w_dff_A_Rx6S3XMy1_0;
	wire w_dff_A_4IaJ9Jsx0_0;
	wire w_dff_A_a2yzrX7B0_0;
	wire w_dff_A_MOLNygZT2_0;
	wire w_dff_A_6ruPEoHw7_0;
	wire w_dff_A_74PywZLp3_0;
	wire w_dff_A_cLjHBqcF3_0;
	wire w_dff_A_bvywiqoq9_0;
	wire w_dff_A_lujqbKWz4_0;
	wire w_dff_A_CD3PBN9n0_0;
	wire w_dff_A_7PYJo2uh6_0;
	wire w_dff_A_X0UhJiYk1_0;
	wire w_dff_A_aRRRFv0Y8_0;
	wire w_dff_A_FGG79RbH4_0;
	wire w_dff_A_7YPD08pT7_0;
	wire w_dff_A_YdEAceCT3_0;
	wire w_dff_A_Zuj8yi9w9_0;
	wire w_dff_A_VbVlLpp90_0;
	wire w_dff_A_TSdVQWS17_0;
	wire w_dff_A_RSBOxWA59_0;
	wire w_dff_A_i1Oq1Gay7_0;
	wire w_dff_A_yMBFHVXl3_0;
	wire w_dff_A_0Uka2LbP9_1;
	wire w_dff_A_U360T9CC3_0;
	wire w_dff_A_wPxsm4iK0_0;
	wire w_dff_A_Kg8I0Y0n2_0;
	wire w_dff_A_0j38edxy7_0;
	wire w_dff_A_2Y5icIgb2_0;
	wire w_dff_A_dbHfyyK58_0;
	wire w_dff_A_XZOwo9XQ9_0;
	wire w_dff_A_gLWV1RHN1_0;
	wire w_dff_A_MH5HzhXf2_0;
	wire w_dff_A_PwtvLxwV8_0;
	wire w_dff_A_EzDjUDpC9_0;
	wire w_dff_A_XhltOiFl0_0;
	wire w_dff_A_luhPqDeG9_0;
	wire w_dff_A_LEEInI1R5_0;
	wire w_dff_A_FRn12GRG9_0;
	wire w_dff_A_g0GJsn7h6_0;
	wire w_dff_A_3pNBqtwD8_0;
	wire w_dff_A_zxtyWdo04_0;
	wire w_dff_A_VrctfqQd1_0;
	wire w_dff_A_99TJh3EW7_0;
	wire w_dff_A_JqdtJ06t7_0;
	wire w_dff_A_KtDeLRLl3_0;
	wire w_dff_A_EN5A6FlR1_0;
	wire w_dff_A_ygNdqXwl1_0;
	wire w_dff_A_wMvJbbhA8_0;
	wire w_dff_A_Ttx6l0hr3_0;
	wire w_dff_A_KehafRC34_1;
	wire w_dff_A_RKitj7TC4_0;
	wire w_dff_A_v5Hpp9362_0;
	wire w_dff_A_DHkfGjeT7_0;
	wire w_dff_A_hclh5f0J6_0;
	wire w_dff_A_6b1ZyCH95_0;
	wire w_dff_A_M9861Nx87_0;
	wire w_dff_A_A6i65Hbv0_0;
	wire w_dff_A_26sdpdJF5_0;
	wire w_dff_A_8cjHCRR13_0;
	wire w_dff_A_4JaGGGtg0_0;
	wire w_dff_A_KtwEtyOQ1_0;
	wire w_dff_A_jNqpDRry8_0;
	wire w_dff_A_W14SfSac1_0;
	wire w_dff_A_Hhz4z6hb4_0;
	wire w_dff_A_FSunHFIz8_0;
	wire w_dff_A_6bmdJBYy1_0;
	wire w_dff_A_tL5K89xr9_0;
	wire w_dff_A_m8gXDkFb9_0;
	wire w_dff_A_2cBFxj3S9_0;
	wire w_dff_A_32Jp2cwV4_0;
	wire w_dff_A_Dq4fH5Wd0_0;
	wire w_dff_A_E7cqtWc16_0;
	wire w_dff_A_nNxW80mH2_0;
	wire w_dff_A_9TjaYfXT7_0;
	wire w_dff_A_ML3DyYOs9_0;
	wire w_dff_A_PNfzOgcU1_0;
	wire w_dff_A_jDpzQ2aJ2_1;
	wire w_dff_A_tY6dgRov0_0;
	wire w_dff_A_EHAtL1do0_0;
	wire w_dff_A_i0qYNqRV0_0;
	wire w_dff_A_m6viLzn54_0;
	wire w_dff_A_rw57U0QD9_0;
	wire w_dff_A_gzSKvJmH2_0;
	wire w_dff_A_X6wI6tdu2_0;
	wire w_dff_A_yxJcPIOq2_0;
	wire w_dff_A_6q6pHyw23_0;
	wire w_dff_A_k436aywX5_0;
	wire w_dff_A_LqiquxaA5_0;
	wire w_dff_A_MQPK4MpP8_0;
	wire w_dff_A_diWiusl89_0;
	wire w_dff_A_OFaqqzmH6_0;
	wire w_dff_A_JDeGCL5C5_0;
	wire w_dff_A_6SibfMMf0_0;
	wire w_dff_A_z2Fv1A696_0;
	wire w_dff_A_BVx5WgYL6_0;
	wire w_dff_A_9yBqeMOd0_0;
	wire w_dff_A_CbC1PrI46_0;
	wire w_dff_A_wOYDwEvW2_0;
	wire w_dff_A_wEfDM12M5_0;
	wire w_dff_A_FZBkPWEB6_0;
	wire w_dff_A_IKrTG20f5_0;
	wire w_dff_A_LedmHbcG8_0;
	wire w_dff_A_eUsqHrRl3_0;
	wire w_dff_A_Y9ZWrAog2_1;
	wire w_dff_A_veWLWexF3_0;
	wire w_dff_A_VjLX6Z4I1_0;
	wire w_dff_A_qzyMCrWd1_0;
	wire w_dff_A_eujmvK7H4_0;
	wire w_dff_A_7YKFQXcO3_0;
	wire w_dff_A_12nbvWII9_0;
	wire w_dff_A_2QTP7w2N8_0;
	wire w_dff_A_1PPORM3p0_0;
	wire w_dff_A_leaXiWlx9_0;
	wire w_dff_A_hT6xkbQA0_0;
	wire w_dff_A_psJDiScC5_0;
	wire w_dff_A_1ES4KZKm2_0;
	wire w_dff_A_tTh4NykM4_0;
	wire w_dff_A_3em2Unc16_0;
	wire w_dff_A_ZVgxaHto9_0;
	wire w_dff_A_stIc75sl6_0;
	wire w_dff_A_5r9aLTWK6_0;
	wire w_dff_A_vvVAzQhW6_0;
	wire w_dff_A_A291gemr5_0;
	wire w_dff_A_3J09ytV54_0;
	wire w_dff_A_gVJLw4Hz0_0;
	wire w_dff_A_nTTKElQZ6_0;
	wire w_dff_A_nj8LPSUi8_0;
	wire w_dff_A_TWLlZgxQ6_0;
	wire w_dff_A_ROH6L8Mh1_0;
	wire w_dff_A_gqAy88Wv7_0;
	wire w_dff_A_0ix5qubp0_1;
	wire w_dff_A_60e6HO8E1_0;
	wire w_dff_A_Z2ux1dkz1_0;
	wire w_dff_A_EZ3yinoM9_0;
	wire w_dff_A_QWkUBcJB8_0;
	wire w_dff_A_bGH9w2Qj4_0;
	wire w_dff_A_d0037ciS8_0;
	wire w_dff_A_mY2sA8sQ3_0;
	wire w_dff_A_cOMZIl043_0;
	wire w_dff_A_qFEhImj31_0;
	wire w_dff_A_YbSTgncB9_0;
	wire w_dff_A_ytvceTSx1_0;
	wire w_dff_A_MDckOEme9_0;
	wire w_dff_A_y0MGcsvL5_0;
	wire w_dff_A_dOX4LlK39_0;
	wire w_dff_A_sZLpTzAN4_0;
	wire w_dff_A_Mthay0yB5_0;
	wire w_dff_A_n0OAJnoI5_0;
	wire w_dff_A_YW1X6Ocm5_0;
	wire w_dff_A_xRQAyEz31_0;
	wire w_dff_A_BPAb1zIa4_0;
	wire w_dff_A_EUz3i6PF0_0;
	wire w_dff_A_5PhaOWOG5_0;
	wire w_dff_A_gXxTGb2c8_0;
	wire w_dff_A_Gqzrmer73_0;
	wire w_dff_A_CeobTZQr2_0;
	wire w_dff_A_YbAhygpP0_0;
	wire w_dff_A_wgAbeICk9_1;
	wire w_dff_A_vQ8ykfQd3_0;
	wire w_dff_A_j2h5m3TC8_0;
	wire w_dff_A_Dd33UVEf8_0;
	wire w_dff_A_dzhl3jx75_0;
	wire w_dff_A_meYIlkPJ0_0;
	wire w_dff_A_h8FAtpXP9_0;
	wire w_dff_A_CcuA5gcs9_0;
	wire w_dff_A_kPlsGiaz6_0;
	wire w_dff_A_q47dh4Xv9_0;
	wire w_dff_A_xlbTtHlf3_0;
	wire w_dff_A_uON0jOl05_0;
	wire w_dff_A_qENXP1JA3_0;
	wire w_dff_A_lZXgQIRJ8_0;
	wire w_dff_A_FZ8KGm6o0_0;
	wire w_dff_A_DYVita5t1_0;
	wire w_dff_A_R1FFuPv26_0;
	wire w_dff_A_u3u5S29D7_0;
	wire w_dff_A_Dm5cneEl9_0;
	wire w_dff_A_MBIAjK7l3_0;
	wire w_dff_A_BK3uQb7X5_0;
	wire w_dff_A_DOB6QybZ2_0;
	wire w_dff_A_YgReLinE3_0;
	wire w_dff_A_9rKlEP7H9_0;
	wire w_dff_A_q0Ahveqj8_0;
	wire w_dff_A_LgfPKULk3_0;
	wire w_dff_A_bR8O3B8A6_0;
	wire w_dff_A_CfDvIimZ4_1;
	wire w_dff_A_3SY1fYpy2_0;
	wire w_dff_A_uKP3BkAP2_0;
	wire w_dff_A_O0bRRyHm6_0;
	wire w_dff_A_tG6w6lsh6_0;
	wire w_dff_A_C3h7PFtu4_0;
	wire w_dff_A_l5AKPo0Y7_0;
	wire w_dff_A_AtfozGDW8_0;
	wire w_dff_A_rfKqZ5L64_0;
	wire w_dff_A_1QBmeoPQ4_0;
	wire w_dff_A_8EEFaWvJ3_0;
	wire w_dff_A_SDT7cqFV1_0;
	wire w_dff_A_n6JsGTOj6_0;
	wire w_dff_A_96C6UDXs3_0;
	wire w_dff_A_dXzzdVar1_0;
	wire w_dff_A_7U8X5o2u5_0;
	wire w_dff_A_BEJd0wnq5_0;
	wire w_dff_A_OtxYU6Rj0_0;
	wire w_dff_A_ODJEpXD01_0;
	wire w_dff_A_wDhPmN9S6_0;
	wire w_dff_A_s2FFEnfo6_0;
	wire w_dff_A_8M1x1tpL9_0;
	wire w_dff_A_v6FtbG5R7_0;
	wire w_dff_A_EwTfW2S17_0;
	wire w_dff_A_nwVFLuv12_0;
	wire w_dff_A_clYmrU0C9_0;
	wire w_dff_A_acC3lP8G3_0;
	wire w_dff_A_8brKNuEG7_1;
	wire w_dff_A_aKo1Xqn97_0;
	wire w_dff_A_elwKw87q0_0;
	wire w_dff_A_4fS7H4Po8_0;
	wire w_dff_A_rVUE7aOe2_0;
	wire w_dff_A_t2roooUt4_0;
	wire w_dff_A_95swoQu66_0;
	wire w_dff_A_n6FSe3V11_0;
	wire w_dff_A_XMF7208w7_0;
	wire w_dff_A_9TuXXtwC8_0;
	wire w_dff_A_rEO7qQeb3_0;
	wire w_dff_A_rjuN1Y3Z7_0;
	wire w_dff_A_dVBFye6q9_0;
	wire w_dff_A_JNkmNgcG5_0;
	wire w_dff_A_VbNjRkFM5_0;
	wire w_dff_A_FAQvIRpn3_0;
	wire w_dff_A_VPqPdqFI2_0;
	wire w_dff_A_yJloMtev6_0;
	wire w_dff_A_5X8zdgpV2_0;
	wire w_dff_A_iC4Re1dy6_0;
	wire w_dff_A_Ra8tLkuT0_0;
	wire w_dff_A_gWn9kqhU6_0;
	wire w_dff_A_yh6t0Gq15_0;
	wire w_dff_A_qhpoD1r02_0;
	wire w_dff_A_G2sZBwY77_0;
	wire w_dff_A_2TcBThQC9_0;
	wire w_dff_A_jE64nwd89_0;
	wire w_dff_A_Sld5T4WZ8_1;
	wire w_dff_A_34QmGbZl7_0;
	wire w_dff_A_9KFCa8dQ2_0;
	wire w_dff_A_gote9Jjd3_0;
	wire w_dff_A_YIm6Z9Vd4_0;
	wire w_dff_A_KBMQbzEZ9_0;
	wire w_dff_A_njBJA7ZT7_0;
	wire w_dff_A_B4BINbny2_0;
	wire w_dff_A_xR9vKVC29_0;
	wire w_dff_A_jKxq7Lip5_0;
	wire w_dff_A_dHZk470L8_0;
	wire w_dff_A_TRp6IpqA5_0;
	wire w_dff_A_lmQL2zhz7_0;
	wire w_dff_A_I62zzrR90_0;
	wire w_dff_A_OlGyySJg5_0;
	wire w_dff_A_TDuLjLqF6_0;
	wire w_dff_A_aEu9tbAC6_0;
	wire w_dff_A_BIXzmfRq9_0;
	wire w_dff_A_zRqCkXAm6_0;
	wire w_dff_A_AXlRiLPI0_0;
	wire w_dff_A_yWTt5LKp9_0;
	wire w_dff_A_I6mraCGq5_0;
	wire w_dff_A_KLEEW6wB9_0;
	wire w_dff_A_vJZZpSxL3_0;
	wire w_dff_A_ebtkvx0J8_0;
	wire w_dff_A_0i8fxZ8s6_0;
	wire w_dff_A_p1vOkPhX0_0;
	wire w_dff_A_2zsj2RB06_1;
	wire w_dff_A_4fMokPse6_0;
	wire w_dff_A_tL7I77yW6_0;
	wire w_dff_A_jVhbtRls8_0;
	wire w_dff_A_OwzqNQWn2_0;
	wire w_dff_A_zbNCJ00i7_0;
	wire w_dff_A_GEt8cfV60_0;
	wire w_dff_A_0ed7RTf54_0;
	wire w_dff_A_KDARhFIF8_0;
	wire w_dff_A_S15NTq9M3_0;
	wire w_dff_A_og65d4NS6_0;
	wire w_dff_A_h0OQBv3X3_0;
	wire w_dff_A_2XRTt7va0_0;
	wire w_dff_A_6gimJ83V0_0;
	wire w_dff_A_uNM2lJSj5_0;
	wire w_dff_A_8LKvGAMC6_0;
	wire w_dff_A_WKWR70IY2_0;
	wire w_dff_A_Zr0bAJhg2_0;
	wire w_dff_A_elYa4sC54_0;
	wire w_dff_A_0eIlEFHI3_0;
	wire w_dff_A_GiLMeY3g4_0;
	wire w_dff_A_upXG6BSh9_0;
	wire w_dff_A_8IeNdCz23_0;
	wire w_dff_A_X7apPuCr8_0;
	wire w_dff_A_qTXzhp2l6_0;
	wire w_dff_A_HWXg7uXL3_0;
	wire w_dff_A_9RVvguRJ3_0;
	wire w_dff_A_r0bXZQNs5_1;
	wire w_dff_A_TYUuYlol5_0;
	wire w_dff_A_jJvJxAKt8_0;
	wire w_dff_A_m93Et6xG1_0;
	wire w_dff_A_1kpfSZtl7_0;
	wire w_dff_A_AE3LxU6A4_0;
	wire w_dff_A_OrSPGh5J2_0;
	wire w_dff_A_ZVhf3FjE9_0;
	wire w_dff_A_TWjwJyzN4_0;
	wire w_dff_A_LJxrGtvv2_0;
	wire w_dff_A_XfPcqyW10_0;
	wire w_dff_A_BhqegnN72_0;
	wire w_dff_A_KG2mIWGi2_0;
	wire w_dff_A_ZbKwdjpD8_0;
	wire w_dff_A_3gFPPP905_0;
	wire w_dff_A_R7GQKwCV2_0;
	wire w_dff_A_3WwNRS7P5_0;
	wire w_dff_A_Bbd6QVDF6_0;
	wire w_dff_A_78QWUj3T9_0;
	wire w_dff_A_RqgrTW7a6_0;
	wire w_dff_A_FKCf7JPf3_0;
	wire w_dff_A_lYizDufl3_0;
	wire w_dff_A_dx2puKVE3_0;
	wire w_dff_A_dp9TUOam1_0;
	wire w_dff_A_x89KjzVS8_0;
	wire w_dff_A_5YCHUmkz0_0;
	wire w_dff_A_b8nv0tNG8_0;
	wire w_dff_A_Z2eAlHCZ6_1;
	wire w_dff_A_bcZdGUgK5_0;
	wire w_dff_A_bj7ynTkS4_0;
	wire w_dff_A_nrqFXvBo7_0;
	wire w_dff_A_Uf5PJKEN2_0;
	wire w_dff_A_jFRqfUQs8_0;
	wire w_dff_A_pLS8XMs39_0;
	wire w_dff_A_oeAUcYnB8_0;
	wire w_dff_A_pfw3LPzS8_0;
	wire w_dff_A_kWuZW1Dl3_0;
	wire w_dff_A_bl5dKVag1_0;
	wire w_dff_A_ug0wHStv7_0;
	wire w_dff_A_3fdMy8mA5_0;
	wire w_dff_A_yWHsVoXZ5_0;
	wire w_dff_A_PmVxckrk5_0;
	wire w_dff_A_cRXroEtT6_0;
	wire w_dff_A_3uqfZWDT8_0;
	wire w_dff_A_tTXs6CmS0_0;
	wire w_dff_A_wvKIbn104_0;
	wire w_dff_A_KP4P7DM01_0;
	wire w_dff_A_eq60TIou0_0;
	wire w_dff_A_RWgDBVme1_0;
	wire w_dff_A_ZQVKaTj07_0;
	wire w_dff_A_Zne4Lcdb1_0;
	wire w_dff_A_SIoTOpVS0_0;
	wire w_dff_A_abRDZ85t4_0;
	wire w_dff_A_ffRooCdc0_0;
	wire w_dff_A_iSHkyrCa3_1;
	wire w_dff_A_wldKCeuE7_0;
	wire w_dff_A_x5zorZ2N2_0;
	wire w_dff_A_Kl9a4Opx7_0;
	wire w_dff_A_FPBSg7oK3_0;
	wire w_dff_A_31aDQApI2_0;
	wire w_dff_A_ZLxOp7Wy4_0;
	wire w_dff_A_yeTNJB2x8_0;
	wire w_dff_A_hx8OWPXr2_0;
	wire w_dff_A_p1jZEzf44_0;
	wire w_dff_A_zVRSIu2W3_0;
	wire w_dff_A_rpwQJ1VC3_0;
	wire w_dff_A_fuEY0MX12_0;
	wire w_dff_A_RqQQatKl2_0;
	wire w_dff_A_59zd85SQ5_0;
	wire w_dff_A_87c7SQa24_0;
	wire w_dff_A_Rg5GfciH7_0;
	wire w_dff_A_6Nab88Ga3_0;
	wire w_dff_A_NziXmPSM4_0;
	wire w_dff_A_PvvByTPX0_0;
	wire w_dff_A_YUWj64uu6_0;
	wire w_dff_A_B0mNSMVQ8_0;
	wire w_dff_A_UpxY3T6g7_0;
	wire w_dff_A_1Dxg9UPR4_0;
	wire w_dff_A_uVtiYIfr9_0;
	wire w_dff_A_cF4kbO6V7_0;
	wire w_dff_A_c5Z2LfNb0_0;
	wire w_dff_A_sSU8Nc0v8_1;
	wire w_dff_A_Vd8vT5mw8_0;
	wire w_dff_A_cBRx5XSn9_0;
	wire w_dff_A_FD2JDzAe8_0;
	wire w_dff_A_LXUM44HZ8_0;
	wire w_dff_A_vFSPL2lh6_0;
	wire w_dff_A_L8HFXflp7_0;
	wire w_dff_A_bEWmp0Cu1_0;
	wire w_dff_A_J0Z7YACD8_0;
	wire w_dff_A_M6XJNGtz2_0;
	wire w_dff_A_tSi5QU954_0;
	wire w_dff_A_QgUQ6Eev2_0;
	wire w_dff_A_E8URVVgC8_0;
	wire w_dff_A_8XEOaskD1_0;
	wire w_dff_A_vXyC5kyo2_0;
	wire w_dff_A_6Z2n1XN15_0;
	wire w_dff_A_6Drssuz64_0;
	wire w_dff_A_fJfna1mC2_0;
	wire w_dff_A_AODNTa8Y4_0;
	wire w_dff_A_ohb9x2Yo1_0;
	wire w_dff_A_C0DyVrQP4_0;
	wire w_dff_A_a3lWSis80_0;
	wire w_dff_A_YkBQzBPW6_0;
	wire w_dff_A_6ZTM6K6r9_0;
	wire w_dff_A_S01Z9pJh6_0;
	wire w_dff_A_QvOY3lw56_0;
	wire w_dff_A_CKt7lR0A0_0;
	wire w_dff_A_Of9VtPSQ2_1;
	wire w_dff_A_PaVupGCu8_0;
	wire w_dff_A_XlXcBwfT2_0;
	wire w_dff_A_QFjQFJ8k0_0;
	wire w_dff_A_9q25cNaT0_0;
	wire w_dff_A_1n0AX2pd9_0;
	wire w_dff_A_moSuIVn52_0;
	wire w_dff_A_lppMUx7P5_0;
	wire w_dff_A_iRztI8lv8_0;
	wire w_dff_A_5GR3O3LJ4_0;
	wire w_dff_A_lifUZu2k3_0;
	wire w_dff_A_V0qjYcJ06_0;
	wire w_dff_A_TKBCnWwv2_0;
	wire w_dff_A_JoZRxH766_0;
	wire w_dff_A_csyF3vNs4_0;
	wire w_dff_A_GMMNQUdh9_0;
	wire w_dff_A_DOyVJfzP0_0;
	wire w_dff_A_JVGGwrzx9_0;
	wire w_dff_A_vXnlVzB12_0;
	wire w_dff_A_CpPmcKRx0_0;
	wire w_dff_A_eXqyGPMG6_0;
	wire w_dff_A_k7snMY0i6_0;
	wire w_dff_A_SAhi3Khp4_0;
	wire w_dff_A_78AbOlIQ3_0;
	wire w_dff_A_wpbIjZ4j4_0;
	wire w_dff_A_GbPeiB3i7_0;
	wire w_dff_A_89JoPaTU5_0;
	wire w_dff_A_ztpM8bzy9_1;
	wire w_dff_A_YTA2BZ5I3_0;
	wire w_dff_A_bk2Q4RW43_0;
	wire w_dff_A_gsswx0004_0;
	wire w_dff_A_0xJdXGsN4_0;
	wire w_dff_A_kZcGVlLW3_0;
	wire w_dff_A_Iyd1tB144_0;
	wire w_dff_A_yGTBdxCo1_0;
	wire w_dff_A_peRNmo5t8_0;
	wire w_dff_A_MFlndP3E2_0;
	wire w_dff_A_fBlaoO5U4_0;
	wire w_dff_A_PtxFxaSy4_0;
	wire w_dff_A_BSbI8NYr8_0;
	wire w_dff_A_cavAD3YF0_0;
	wire w_dff_A_2QWqgX0u2_0;
	wire w_dff_A_55crmJhf1_0;
	wire w_dff_A_6cnIPeem5_0;
	wire w_dff_A_iM8ZRctz5_0;
	wire w_dff_A_htYT306Z9_0;
	wire w_dff_A_XOSLuCov6_0;
	wire w_dff_A_UPgu4GZU9_0;
	wire w_dff_A_fwpITZpx7_0;
	wire w_dff_A_SowneOBg8_0;
	wire w_dff_A_sKnAYa0p6_0;
	wire w_dff_A_Qc66GIHC0_0;
	wire w_dff_A_x1lzBeLR7_0;
	wire w_dff_A_1wMcQHme5_0;
	wire w_dff_A_xlD6j1Zi9_1;
	wire w_dff_A_WFX8D3M31_0;
	wire w_dff_A_HTsFE5wa1_0;
	wire w_dff_A_JQvnTFgp9_0;
	wire w_dff_A_QhzKupRl6_0;
	wire w_dff_A_wKWr9rwM1_0;
	wire w_dff_A_r5fBS3tw5_0;
	wire w_dff_A_U1mWXhPx9_0;
	wire w_dff_A_BirBGLRM4_0;
	wire w_dff_A_pqlRep9s4_0;
	wire w_dff_A_n7UdhcRQ5_0;
	wire w_dff_A_VFGVCeBI0_0;
	wire w_dff_A_NTBFRgI07_0;
	wire w_dff_A_z99r3vfj4_0;
	wire w_dff_A_zIxeeIuE7_0;
	wire w_dff_A_uBUobIX13_0;
	wire w_dff_A_BMYthtfc2_0;
	wire w_dff_A_5Z7Y6kIK4_0;
	wire w_dff_A_cJi8gR9v5_0;
	wire w_dff_A_3ls0bRIv3_0;
	wire w_dff_A_VG7KSCzD7_0;
	wire w_dff_A_Ef51zWPW8_0;
	wire w_dff_A_i7bXvKhp7_0;
	wire w_dff_A_oQb5QDZF1_0;
	wire w_dff_A_ae9vdxwT5_0;
	wire w_dff_A_6Ks6GMBT4_0;
	wire w_dff_A_8fgE9Mbg2_0;
	wire w_dff_A_HrHW1qMA5_1;
	wire w_dff_A_EUKT3el10_0;
	wire w_dff_A_am6qkB8O7_0;
	wire w_dff_A_Kwxxnfsg7_0;
	wire w_dff_A_JlJeVVQf2_0;
	wire w_dff_A_hmx2HFlt2_0;
	wire w_dff_A_MCR8gLTZ4_0;
	wire w_dff_A_gGznf6Cf6_0;
	wire w_dff_A_pVYmjbcm9_0;
	wire w_dff_A_l1R2MwS65_0;
	wire w_dff_A_wqHZPVXM5_0;
	wire w_dff_A_VBvUbC149_0;
	wire w_dff_A_LR9doiFJ6_0;
	wire w_dff_A_jykKafmX0_0;
	wire w_dff_A_bB9YN1OB8_0;
	wire w_dff_A_H1cn6M4r3_0;
	wire w_dff_A_sAwmomJL8_0;
	wire w_dff_A_8soKMIOm7_0;
	wire w_dff_A_0Mvz93Qw7_0;
	wire w_dff_A_SajoIkiP4_0;
	wire w_dff_A_Zd97Z9xm1_0;
	wire w_dff_A_c6dqsFPr5_0;
	wire w_dff_A_sTNDFMuf6_0;
	wire w_dff_A_pXsvqIEo4_0;
	wire w_dff_A_Hs586TUD0_0;
	wire w_dff_A_HnFBbxtV7_0;
	wire w_dff_A_TxLtrfLw6_0;
	wire w_dff_A_7HM1DQ839_1;
	wire w_dff_A_slaPthN13_0;
	wire w_dff_A_YGtvSk2a1_0;
	wire w_dff_A_O3mWxzfZ8_0;
	wire w_dff_A_TGV802kf6_0;
	wire w_dff_A_rtzV0jA87_0;
	wire w_dff_A_Z7vxoIqD7_0;
	wire w_dff_A_Gq0fpfWh7_0;
	wire w_dff_A_2ttSukOJ0_0;
	wire w_dff_A_59GyhNNz7_0;
	wire w_dff_A_tcg9Lg7q2_0;
	wire w_dff_A_w6j6igK46_0;
	wire w_dff_A_k7MeAYFZ0_0;
	wire w_dff_A_qoPxUERk8_0;
	wire w_dff_A_L3qDIqAZ0_0;
	wire w_dff_A_dx3MgIUi8_0;
	wire w_dff_A_v0YkqLBK7_0;
	wire w_dff_A_NoRKP3kl9_0;
	wire w_dff_A_XBQlT7uD1_0;
	wire w_dff_A_vxwa7HVZ4_0;
	wire w_dff_A_5iPtCTzu0_0;
	wire w_dff_A_9CM9qpbB9_0;
	wire w_dff_A_NpEibPV07_0;
	wire w_dff_A_e41xzA2k6_0;
	wire w_dff_A_2wodT8tr6_0;
	wire w_dff_A_7gArp3mZ9_0;
	wire w_dff_A_hGOFpqrP7_1;
	wire w_dff_A_dUxLuROW2_0;
	wire w_dff_A_o4lzmtxy2_0;
	wire w_dff_A_hEimCZFb9_0;
	wire w_dff_A_pxTRyZP67_0;
	wire w_dff_A_E8vyQKM88_0;
	wire w_dff_A_mCvSdVtJ6_0;
	wire w_dff_A_LQ4z4i7j8_0;
	wire w_dff_A_KMTyXsnq2_0;
	wire w_dff_A_OVpZpCz27_0;
	wire w_dff_A_qGTsLLm01_0;
	wire w_dff_A_xHqDG8Uq6_0;
	wire w_dff_A_raLbnrIY2_0;
	wire w_dff_A_zwQJNk777_0;
	wire w_dff_A_mbkooX5s5_0;
	wire w_dff_A_IHN0Tpaa5_0;
	wire w_dff_A_Q10zCkCy1_0;
	wire w_dff_A_WMtmX2323_0;
	wire w_dff_A_shvCxdtb1_0;
	wire w_dff_A_ET310NpY6_0;
	wire w_dff_A_xTQCmrBO2_0;
	wire w_dff_A_ZnJv6qjc9_0;
	wire w_dff_A_KbRCv3KB1_0;
	wire w_dff_A_KU2bup1o5_0;
	wire w_dff_A_tapjk4Cf7_0;
	wire w_dff_A_LEd0GuqU0_0;
	wire w_dff_A_FjMIKdmG3_0;
	wire w_dff_A_56ni4neV6_1;
	wire w_dff_A_R5Vj1P5q7_0;
	wire w_dff_A_QWr8flty6_0;
	wire w_dff_A_GtW6k2107_0;
	wire w_dff_A_tDq3HhOq7_0;
	wire w_dff_A_Q4Xugie34_0;
	wire w_dff_A_JC8BfTjG5_0;
	wire w_dff_A_QiqoRcO32_0;
	wire w_dff_A_6AJtieuS4_0;
	wire w_dff_A_XN3Elhhm7_0;
	wire w_dff_A_I4To7Ltp9_0;
	wire w_dff_A_odBDM5Bu5_0;
	wire w_dff_A_lfWSCPaD4_0;
	wire w_dff_A_OS7VMeJR8_0;
	wire w_dff_A_iTc3HYKq6_0;
	wire w_dff_A_gosv3Rzz6_0;
	wire w_dff_A_GNsYfa1T7_0;
	wire w_dff_A_xRDdIrDJ1_0;
	wire w_dff_A_1JdbvD3D8_0;
	wire w_dff_A_kvZw8Kj53_0;
	wire w_dff_A_txsNWER01_0;
	wire w_dff_A_Td4NXJIu5_0;
	wire w_dff_A_z69aD0NZ1_0;
	wire w_dff_A_xbqszPMa7_0;
	wire w_dff_A_UPOudb9i6_0;
	wire w_dff_A_ChtXKLQr0_0;
	wire w_dff_A_I0FN6nyc1_0;
	wire w_dff_A_sAMargQa3_1;
	wire w_dff_A_m2BflVSL6_0;
	wire w_dff_A_fIraQLK07_0;
	wire w_dff_A_A66Nf7J08_0;
	wire w_dff_A_GA9WXupi3_0;
	wire w_dff_A_oOoin8CA8_0;
	wire w_dff_A_ciEf2wi22_0;
	wire w_dff_A_s1gJ98CE2_0;
	wire w_dff_A_ZKWJVfOw4_0;
	wire w_dff_A_PCAAxjED7_0;
	wire w_dff_A_OzdCoDdg1_0;
	wire w_dff_A_zvVnal4D5_0;
	wire w_dff_A_VLfBbvTj2_0;
	wire w_dff_A_LXGn4nOU4_0;
	wire w_dff_A_EgLkMdKR0_0;
	wire w_dff_A_zADllPJ25_0;
	wire w_dff_A_SHtKDGAd4_0;
	wire w_dff_A_QivZwlB87_0;
	wire w_dff_A_awhgtQZa6_0;
	wire w_dff_A_dMILZV8T8_0;
	wire w_dff_A_ISwco8zU4_0;
	wire w_dff_A_cEsRmd8r1_0;
	wire w_dff_A_z3NkZ1Zz8_0;
	wire w_dff_A_nxkUreNI3_0;
	wire w_dff_A_ewcPRaoT8_0;
	wire w_dff_A_hr1ayws02_0;
	wire w_dff_A_oUyfBQsb8_0;
	wire w_dff_A_OZMI4Ga77_2;
	wire w_dff_A_n4ToBhTj3_0;
	wire w_dff_A_Oexla1mg8_0;
	wire w_dff_A_n8YxaAaE9_0;
	wire w_dff_A_GH91YwdK7_0;
	wire w_dff_A_Oslq1ZHc2_0;
	wire w_dff_A_czGeNeLo8_0;
	wire w_dff_A_XpI3nqT53_0;
	wire w_dff_A_axDLYPgR4_0;
	wire w_dff_A_x1gIkGE00_0;
	wire w_dff_A_UY1Vl4A43_0;
	wire w_dff_A_kUuPiZCT1_0;
	wire w_dff_A_LNZgwBAN9_0;
	wire w_dff_A_NcwNWXL39_0;
	wire w_dff_A_UHTWrzuF2_0;
	wire w_dff_A_PEaEW2Jp1_0;
	wire w_dff_A_l6MeY4mM7_0;
	wire w_dff_A_gUTgeiKU5_0;
	wire w_dff_A_xu9AsHLe2_0;
	wire w_dff_A_pSXltQpo6_0;
	wire w_dff_A_5F2korNF4_0;
	wire w_dff_A_6TPs2gno4_0;
	wire w_dff_A_p6bj0BKZ8_0;
	wire w_dff_A_QQO17DdI0_0;
	wire w_dff_A_0Cs0mKtd3_0;
	wire w_dff_A_rJCz512O4_0;
	wire w_dff_A_SGEwqHKw4_1;
	wire w_dff_A_WCjFhd9u8_0;
	wire w_dff_A_ii5WTJeC7_0;
	wire w_dff_A_gTJrP7ff0_0;
	wire w_dff_A_jeZVLKG73_0;
	wire w_dff_A_FZAJqJdk5_0;
	wire w_dff_A_p3KIA5Tw7_0;
	wire w_dff_A_mQUyU7to6_0;
	wire w_dff_A_yVf3E3Uu5_0;
	wire w_dff_A_jl7uMHUv9_0;
	wire w_dff_A_gvJjEoSf3_0;
	wire w_dff_A_EcJpwJNy2_0;
	wire w_dff_A_Bq18wGRS4_0;
	wire w_dff_A_XBwn5tcC5_0;
	wire w_dff_A_qo4tyB984_0;
	wire w_dff_A_LYkosXUf5_0;
	wire w_dff_A_u5We17kT1_0;
	wire w_dff_A_yTQLrgwF3_0;
	wire w_dff_A_M8GcD04g3_0;
	wire w_dff_A_xWHtDopP6_0;
	wire w_dff_A_vxrV3DXv5_0;
	wire w_dff_A_81JwQljV9_0;
	wire w_dff_A_jbDTqvTB5_0;
	wire w_dff_A_sIt0Y2zZ6_0;
	wire w_dff_A_J25vNCWP8_1;
	wire w_dff_A_BkuQIf3C9_0;
	wire w_dff_A_bUcGTBD71_0;
	wire w_dff_A_oH689uGw3_0;
	wire w_dff_A_mwC6lZBd9_0;
	wire w_dff_A_XUmI1UNj4_0;
	wire w_dff_A_cU0zo3iN6_0;
	wire w_dff_A_az6wwGDe5_0;
	wire w_dff_A_zALtfvep0_0;
	wire w_dff_A_PEtQF9Zs2_0;
	wire w_dff_A_h7BfEb0S1_0;
	wire w_dff_A_WCYLutiH9_0;
	wire w_dff_A_PMMcucqa7_0;
	wire w_dff_A_wKNWm0Im7_0;
	wire w_dff_A_drcZnwBR6_0;
	wire w_dff_A_QT2ZJ9WB0_0;
	wire w_dff_A_SlAP4dXO4_0;
	wire w_dff_A_DfKGz3FT7_0;
	wire w_dff_A_2KAjtvHe8_0;
	wire w_dff_A_TEfYyzUs7_0;
	wire w_dff_A_mbFJ79w41_0;
	wire w_dff_A_gs4EZLeV6_0;
	wire w_dff_A_sVf5JINW3_0;
	wire w_dff_A_CAdzPeq91_0;
	wire w_dff_A_6zPirW7D7_1;
	wire w_dff_A_swJY6FON9_0;
	wire w_dff_A_xaDhx7ov5_0;
	wire w_dff_A_UpdGSlPz2_0;
	wire w_dff_A_G6xJVx3O5_0;
	wire w_dff_A_rObM40D18_0;
	wire w_dff_A_Lpa9olqb6_0;
	wire w_dff_A_oQOAjhPd0_0;
	wire w_dff_A_abVQBL915_0;
	wire w_dff_A_pxsPcSCM4_0;
	wire w_dff_A_x2WDlAoM1_0;
	wire w_dff_A_yyUvmJvo3_0;
	wire w_dff_A_z5wRCZwn6_0;
	wire w_dff_A_Ce7shpOP1_0;
	wire w_dff_A_XUqDQT3z8_0;
	wire w_dff_A_pSZMH1zl9_0;
	wire w_dff_A_BmIQnGyM4_0;
	wire w_dff_A_RPpeSkqQ1_0;
	wire w_dff_A_yPmdc3T84_0;
	wire w_dff_A_WIOpWlE71_0;
	wire w_dff_A_7IuK3eYW4_0;
	wire w_dff_A_T6cX8LI91_0;
	wire w_dff_A_vKhBUJMz9_0;
	wire w_dff_A_Wh0cJCrl6_0;
	wire w_dff_A_NzXdC8ZK7_1;
	wire w_dff_A_pn4KMOni0_0;
	wire w_dff_A_QifoiltK8_0;
	wire w_dff_A_aHvpLeWs7_0;
	wire w_dff_A_BRpil0t39_0;
	wire w_dff_A_CVCOIa1X8_0;
	wire w_dff_A_5fxMVuoV7_0;
	wire w_dff_A_O7mUvSFn5_0;
	wire w_dff_A_PLsjc6cc5_0;
	wire w_dff_A_xg6GiZUB3_0;
	wire w_dff_A_VuT2Z1Wn9_0;
	wire w_dff_A_BFwDx8kC1_0;
	wire w_dff_A_TcA86cJC5_0;
	wire w_dff_A_5qZROEJn9_0;
	wire w_dff_A_753z8Nll3_0;
	wire w_dff_A_7quX9Zo90_0;
	wire w_dff_A_kf8qv9KM2_0;
	wire w_dff_A_nQgJ8EyW4_0;
	wire w_dff_A_uCx06Mjp9_0;
	wire w_dff_A_C7IdZ9tA1_0;
	wire w_dff_A_TovBFwZG6_0;
	wire w_dff_A_mKFrwWiS7_0;
	wire w_dff_A_h8GdkFMM1_0;
	wire w_dff_A_9t41dwCj1_0;
	wire w_dff_A_15oUKSIM7_1;
	wire w_dff_A_rV1SaM8m4_0;
	wire w_dff_A_7kl6Y6b35_0;
	wire w_dff_A_OkPxIsGP7_0;
	wire w_dff_A_V7Cwdbaz4_0;
	wire w_dff_A_GQS04JOe1_0;
	wire w_dff_A_D4vzyFZz8_0;
	wire w_dff_A_Elk81OvA1_0;
	wire w_dff_A_ZetmPexk7_0;
	wire w_dff_A_v9me7U372_0;
	wire w_dff_A_z6KKGThk2_0;
	wire w_dff_A_bDpofzk43_0;
	wire w_dff_A_weCviYfJ6_0;
	wire w_dff_A_JFX9dQ9t1_0;
	wire w_dff_A_JWPMpJnY7_0;
	wire w_dff_A_XwDr6baQ2_0;
	wire w_dff_A_xbKGdnls8_0;
	wire w_dff_A_UYM8VOwr7_0;
	wire w_dff_A_025twQV96_0;
	wire w_dff_A_YPyFNXBa0_0;
	wire w_dff_A_sQrSQiKd4_0;
	wire w_dff_A_JV1PFuuH3_0;
	wire w_dff_A_BaP4BC360_0;
	wire w_dff_A_wiyjVIP52_0;
	wire w_dff_A_IVaOQYXD7_0;
	wire w_dff_A_Ld4fhGte8_0;
	wire w_dff_A_V2Sjjcjm2_0;
	wire w_dff_A_FqMa6rxn5_1;
	wire w_dff_A_KxnVtkzY6_0;
	wire w_dff_A_jKIs852d6_0;
	wire w_dff_A_XOUuMD9C8_0;
	wire w_dff_A_ivjdorIe2_0;
	wire w_dff_A_Ge9Q8Dmh1_0;
	wire w_dff_A_Lavmisb85_0;
	wire w_dff_A_dUCZCv3R3_0;
	wire w_dff_A_BKJ67eLy5_0;
	wire w_dff_A_VjEOSWgg9_0;
	wire w_dff_A_9JNxaAIb7_0;
	wire w_dff_A_QrGPKV7s9_0;
	wire w_dff_A_fmQ1iOxl0_0;
	wire w_dff_A_X4n5i12Y8_0;
	wire w_dff_A_MsuKoody8_0;
	wire w_dff_A_YBAXKzI72_0;
	wire w_dff_A_H96RlYwA5_0;
	wire w_dff_A_G1RvKQWe0_0;
	wire w_dff_A_pgDFHFYF3_0;
	wire w_dff_A_023pmYW58_0;
	wire w_dff_A_9ZZai5io4_0;
	wire w_dff_A_UNB6st835_0;
	wire w_dff_A_YZMP34Wf4_0;
	wire w_dff_A_hWw4vhj30_0;
	wire w_dff_A_PFUIfVnV2_0;
	wire w_dff_A_n8HpsUKG8_0;
	wire w_dff_A_mMNe0m2b8_0;
	wire w_dff_A_uzDJ9L3F8_2;
	wire w_dff_A_DFczi5Cy3_0;
	wire w_dff_A_bEg6PutY6_0;
	wire w_dff_A_dXqxX0Ng7_0;
	wire w_dff_A_OaP8C8ge8_0;
	wire w_dff_A_9zm7ukga8_0;
	wire w_dff_A_nqJcaAhV4_0;
	wire w_dff_A_pMluvbk79_0;
	wire w_dff_A_twUM6LXZ7_0;
	wire w_dff_A_9rL0ABE20_0;
	wire w_dff_A_s4WBAphs3_0;
	wire w_dff_A_LS2lmRPx5_0;
	wire w_dff_A_Zk1oiQwt5_0;
	wire w_dff_A_ETPYdynt7_0;
	wire w_dff_A_r7tX8glB7_0;
	wire w_dff_A_WEqtMSzi1_0;
	wire w_dff_A_Llu0yBvG8_0;
	wire w_dff_A_5Lk3h4vZ4_0;
	wire w_dff_A_xUPpYiNs0_0;
	wire w_dff_A_Cl87TgwO7_0;
	wire w_dff_A_u2QYT7gV9_0;
	wire w_dff_A_QtTE4g8n0_0;
	wire w_dff_A_PRGlECK02_0;
	wire w_dff_A_zIwBq5YE5_0;
	wire w_dff_A_S3BlpmZH6_0;
	wire w_dff_A_x6qNQfhM0_1;
	wire w_dff_A_ollMUi7J4_0;
	wire w_dff_A_X0LsElUZ2_0;
	wire w_dff_A_wcaTEiE82_0;
	wire w_dff_A_KqAr2P2W4_0;
	wire w_dff_A_eDd6yCzQ0_0;
	wire w_dff_A_9qFENikU0_0;
	wire w_dff_A_L5KKnOQC6_0;
	wire w_dff_A_aCaHXAuk5_0;
	wire w_dff_A_wqYAbRbZ0_0;
	wire w_dff_A_e9AUNY7E1_0;
	wire w_dff_A_1wqVMcOx7_0;
	wire w_dff_A_BTrkWGRa5_0;
	wire w_dff_A_X2GkVYsK2_0;
	wire w_dff_A_GFRScXE64_0;
	wire w_dff_A_1dymERuQ2_0;
	wire w_dff_A_p9IXDxTq3_0;
	wire w_dff_A_tuNHTqcG6_0;
	wire w_dff_A_3ac1XEpq5_0;
	wire w_dff_A_QZyhMrW18_0;
	wire w_dff_A_IYyvNjoF3_0;
	wire w_dff_A_BRmrOcId6_0;
	wire w_dff_A_8CFnMlOT8_0;
	wire w_dff_A_aDB1Pwe90_0;
	wire w_dff_A_qCtZmxzF6_0;
	wire w_dff_A_DGYT1Nro3_0;
	wire w_dff_A_WJXAWJxz0_2;
	wire w_dff_A_9v7UGhX00_0;
	wire w_dff_A_oxGZTti87_0;
	wire w_dff_A_mCco08TC7_0;
	wire w_dff_A_bKH8u0f57_0;
	wire w_dff_A_jg48mVdB2_0;
	wire w_dff_A_QUDuOjuV3_0;
	wire w_dff_A_nSXQXXB28_0;
	wire w_dff_A_LzFWpX7k9_0;
	wire w_dff_A_ebub0rke1_0;
	wire w_dff_A_6JScAf7E9_0;
	wire w_dff_A_4kH7o5Ex6_0;
	wire w_dff_A_2jrSi9ya2_0;
	wire w_dff_A_GuTi3FQS0_0;
	wire w_dff_A_7y81J92U0_0;
	wire w_dff_A_X7yeDhV98_0;
	wire w_dff_A_csa7LC7O1_0;
	wire w_dff_A_SKKFc0Vi4_0;
	wire w_dff_A_09K4opfR6_0;
	wire w_dff_A_3lBFDCFr9_0;
	wire w_dff_A_Ih72erhV1_0;
	wire w_dff_A_p6Swh93x4_0;
	wire w_dff_A_FN558NaB2_0;
	wire w_dff_A_u6HZNBGs2_0;
	wire w_dff_A_CFzJVzmR7_0;
	wire w_dff_A_1X4oNfns3_2;
	wire w_dff_A_ZhBZZBgd5_0;
	wire w_dff_A_vrlc2RpM8_0;
	wire w_dff_A_FHLtO33B0_0;
	wire w_dff_A_S1NCbxzt8_0;
	wire w_dff_A_4GfGlBmI2_0;
	wire w_dff_A_QsgpELKQ1_0;
	wire w_dff_A_aSXJcHvT5_0;
	wire w_dff_A_vs7GopUV6_0;
	wire w_dff_A_iLrHKmur7_0;
	wire w_dff_A_gLVJe10g9_0;
	wire w_dff_A_jDKNfY3o5_0;
	wire w_dff_A_JPKXI0BP3_0;
	wire w_dff_A_c7dIGHaN4_0;
	wire w_dff_A_CaoHIMYz3_0;
	wire w_dff_A_GfySpbKj7_0;
	wire w_dff_A_pttiFYPI0_0;
	wire w_dff_A_Ihyh8TZa7_0;
	wire w_dff_A_Rw2f9WHk6_0;
	wire w_dff_A_NDiYw3uO0_0;
	wire w_dff_A_0ni8nRFt8_0;
	wire w_dff_A_KYjym8t20_0;
	wire w_dff_A_06FEdL4F2_0;
	wire w_dff_A_u5juNdXE1_0;
	wire w_dff_A_BPLu96TO4_1;
	wire w_dff_A_B2WkPzf57_0;
	wire w_dff_A_LmjfS6Hj3_0;
	wire w_dff_A_IhR9W28s1_0;
	wire w_dff_A_raudKgbW1_0;
	wire w_dff_A_oW8Kzrdr5_0;
	wire w_dff_A_FDFv2MiR7_0;
	wire w_dff_A_PM3C1zbs7_0;
	wire w_dff_A_WZBNOmlY7_0;
	wire w_dff_A_fXJ3jRIS6_0;
	wire w_dff_A_XSXfg8e04_0;
	wire w_dff_A_8nILk8zQ7_0;
	wire w_dff_A_TGsacql63_0;
	wire w_dff_A_0B6ixsIV9_0;
	wire w_dff_A_wG9agYSb6_0;
	wire w_dff_A_cYleF8c42_0;
	wire w_dff_A_P1KVfEbT6_0;
	wire w_dff_A_agUPurLr9_0;
	wire w_dff_A_ZbzVtPQr4_0;
	wire w_dff_A_0OFphQqV0_0;
	wire w_dff_A_MmzAFegM3_0;
	wire w_dff_A_paIQBduA2_0;
	wire w_dff_A_fmRShWyS8_0;
	wire w_dff_A_FntllQ3v5_0;
	wire w_dff_A_rfdWNpQA6_0;
	wire w_dff_A_HTNiFf2C7_0;
	wire w_dff_A_GX6m9gnD6_2;
	wire w_dff_A_Ex4fV9vq1_0;
	wire w_dff_A_WBUNxKt92_0;
	wire w_dff_A_sygmZ1Ir3_0;
	wire w_dff_A_9PWgd9sw8_0;
	wire w_dff_A_IP5rtZp00_0;
	wire w_dff_A_LUsZfq3G6_0;
	wire w_dff_A_Bg0OjLYG3_0;
	wire w_dff_A_lPcWjmYV2_0;
	wire w_dff_A_isYsmanl4_0;
	wire w_dff_A_DMsNzaUo0_0;
	wire w_dff_A_beOfWyyP7_0;
	wire w_dff_A_ry638cHX8_0;
	wire w_dff_A_4Wvqgncc0_0;
	wire w_dff_A_EYJczFbM6_0;
	wire w_dff_A_Xr9txrBs0_0;
	wire w_dff_A_SfdAQZmb0_0;
	wire w_dff_A_98Jc2vF24_0;
	wire w_dff_A_b9r4nJtd6_0;
	wire w_dff_A_RVjpgOoh2_0;
	wire w_dff_A_8FdHHMt39_0;
	wire w_dff_A_hVkwK2D39_0;
	wire w_dff_A_z6N7pVq27_0;
	wire w_dff_A_EXYENh2H3_0;
	wire w_dff_A_Af8wiAcQ9_1;
	wire w_dff_A_aH4naish2_0;
	wire w_dff_A_pashgodO6_0;
	wire w_dff_A_El09sTYD7_0;
	wire w_dff_A_K1aFsXvG3_0;
	wire w_dff_A_jM8U3OSz4_0;
	wire w_dff_A_DbBfKWCV8_0;
	wire w_dff_A_Z6tbIEYD7_0;
	wire w_dff_A_duoFa2TD3_0;
	wire w_dff_A_xdPFVWud3_0;
	wire w_dff_A_amL6RgJj2_0;
	wire w_dff_A_RY2nQBeY6_0;
	wire w_dff_A_y3KRjYep7_0;
	wire w_dff_A_uTB6Ol2B9_0;
	wire w_dff_A_6j4n5Yqy8_0;
	wire w_dff_A_cSUcNv3m2_0;
	wire w_dff_A_JLugpLH33_0;
	wire w_dff_A_geO3nQNh0_0;
	wire w_dff_A_z1lCrkHb7_0;
	wire w_dff_A_YT339kW83_0;
	wire w_dff_A_eTLTVcZb4_0;
	wire w_dff_A_tPE8SIMk4_0;
	wire w_dff_A_25mWouR81_0;
	wire w_dff_A_QcUtAhad9_0;
	wire w_dff_A_2nMDvhkZ0_0;
	wire w_dff_A_vrhFqKrc7_0;
	wire w_dff_A_g4RNV2No7_0;
	wire w_dff_A_0VY9qskf0_2;
	wire w_dff_A_lPgAGG3q1_0;
	wire w_dff_A_APXpKShu5_0;
	wire w_dff_A_gddMmb086_0;
	wire w_dff_A_S9YakP1i6_0;
	wire w_dff_A_M7m6buvZ5_0;
	wire w_dff_A_LUiFWqA37_0;
	wire w_dff_A_ssKtOtWQ2_0;
	wire w_dff_A_UklNp1I48_0;
	wire w_dff_A_GyGplFYw1_0;
	wire w_dff_A_5x6htadB1_0;
	wire w_dff_A_a5CW95X31_0;
	wire w_dff_A_dxGGJhVn3_0;
	wire w_dff_A_t2u1sknl2_0;
	wire w_dff_A_FxF6y2vM8_0;
	wire w_dff_A_7sDV28nT3_0;
	wire w_dff_A_rPiihOKe1_0;
	wire w_dff_A_2SNozCGI0_0;
	wire w_dff_A_4ENMKsBs6_0;
	wire w_dff_A_LUT5gSwh7_0;
	wire w_dff_A_dG3qBhfD4_0;
	wire w_dff_A_fghbiNyz9_0;
	wire w_dff_A_2M9YlSoT1_0;
	wire w_dff_A_9Tb4U9sM0_0;
	wire w_dff_A_7weKCX994_0;
	wire w_dff_A_jkmJ3FGC5_0;
	wire w_dff_A_G6f97vGW1_2;
	wire w_dff_A_s8xf03aG6_0;
	wire w_dff_A_OCU7vohc1_0;
	wire w_dff_A_VrRETt0x9_0;
	wire w_dff_A_nwGFbIDK8_0;
	wire w_dff_A_OmZndJ3G8_0;
	wire w_dff_A_e2Q9b4E56_0;
	wire w_dff_A_FlZOn2Or2_0;
	wire w_dff_A_VocoLcD50_0;
	wire w_dff_A_lcPBdZM54_0;
	wire w_dff_A_hn78JPsk4_0;
	wire w_dff_A_geTMApaP0_0;
	wire w_dff_A_A221yhql8_0;
	wire w_dff_A_3TOpHBz23_0;
	wire w_dff_A_dqX3mFAf6_0;
	wire w_dff_A_GuAxUeW23_0;
	wire w_dff_A_ppNgMf3V4_0;
	wire w_dff_A_bXcR52dd6_0;
	wire w_dff_A_hiw6Tp391_0;
	wire w_dff_A_BqBGIG8B9_0;
	wire w_dff_A_EDqhMU9M5_0;
	wire w_dff_A_tmAqux6d0_2;
	wire w_dff_A_7bncmJrH1_2;
	wire w_dff_A_oxo8IFOF4_0;
	wire w_dff_A_NnB8316l5_0;
	wire w_dff_A_XCkeH2EA7_0;
	wire w_dff_A_Onh8qkL43_0;
	wire w_dff_A_tiBrdGfd2_0;
	wire w_dff_A_yqGXmjzH1_0;
	wire w_dff_A_slq4IEGl3_2;
	wire w_dff_A_49d9nwLz0_0;
	wire w_dff_A_aAWMaHUU6_0;
	wire w_dff_A_TLjT1jhb1_0;
	wire w_dff_A_2fpl2d8b8_0;
	wire w_dff_A_2mIXvj9h8_0;
	wire w_dff_A_P0LTGYCI5_0;
	wire w_dff_A_xynYSXoD0_2;
	wire w_dff_A_7SRXhOvO3_2;
	wire w_dff_A_qCKrcPKM0_0;
	wire w_dff_A_oLHtzAyD0_0;
	wire w_dff_A_y9fU334t0_0;
	wire w_dff_A_iOBIuayx8_0;
	wire w_dff_A_g1FIEsQG9_0;
	wire w_dff_A_QOPMQEOA4_0;
	wire w_dff_A_k6TNAtKY3_0;
	wire w_dff_A_QbskiEbA7_0;
	wire w_dff_A_nHxBmp7f6_0;
	wire w_dff_A_kYpTbEXj1_0;
	wire w_dff_A_djZcg1LF8_0;
	wire w_dff_A_YFqxQxk80_0;
	wire w_dff_A_9djJd31R7_0;
	wire w_dff_A_iLon1dHl7_0;
	wire w_dff_A_ZxG7VkOx2_2;
	wire w_dff_A_buwlAT6j5_0;
	wire w_dff_A_iir7dVLr7_0;
	wire w_dff_A_t99NrWx89_0;
	wire w_dff_A_k2xuEJhq2_0;
	wire w_dff_A_5lcdd36d9_0;
	wire w_dff_A_Jga4aHfz7_0;
	wire w_dff_A_RvlmARqO2_0;
	wire w_dff_A_Ro8C5pz43_0;
	wire w_dff_A_nz3BPLfr4_0;
	wire w_dff_A_TxUb3m2O8_0;
	wire w_dff_A_66DJyi1t6_0;
	wire w_dff_A_SYr65DJ72_0;
	wire w_dff_A_yVq3gOil5_0;
	wire w_dff_A_4yEgPXer3_0;
	wire w_dff_A_2OTiDwfv0_0;
	wire w_dff_A_PUlOZRWD3_0;
	wire w_dff_A_vdMi5oyR9_2;
	wire w_dff_A_7VqXO72Z3_0;
	wire w_dff_A_kHutkUE59_0;
	wire w_dff_A_pMDITxTf6_0;
	wire w_dff_A_r99BU6pK1_0;
	wire w_dff_A_tJLzHwmR6_0;
	wire w_dff_A_cdUZt36Y9_0;
	wire w_dff_A_7DQpceER2_0;
	wire w_dff_A_kJdg2TJO2_0;
	wire w_dff_A_HDjEF4hZ9_0;
	wire w_dff_A_N3DH1ayv2_0;
	wire w_dff_A_ZUqMxNS22_0;
	wire w_dff_A_hlbWUXh28_0;
	wire w_dff_A_pAvAUTJu4_0;
	wire w_dff_A_AYz5eDMm6_0;
	wire w_dff_A_VwaSmJ2w7_0;
	wire w_dff_A_ZKkaejFi5_0;
	wire w_dff_A_kLbTUx1v9_0;
	wire w_dff_A_UGZaqdrl9_2;
	wire w_dff_A_Yc9VjNUH1_0;
	wire w_dff_A_yiTi0O691_0;
	wire w_dff_A_3jugHNN26_0;
	wire w_dff_A_DLBAkYuf0_0;
	wire w_dff_A_fetJtNLW0_0;
	wire w_dff_A_QrLrEXi49_0;
	wire w_dff_A_lcYw7r1L9_0;
	wire w_dff_A_7iTlmmo35_0;
	wire w_dff_A_odoTsM1w6_0;
	wire w_dff_A_OjaMMZRV2_0;
	wire w_dff_A_03qjPbrJ8_0;
	wire w_dff_A_nN49KSXe7_0;
	wire w_dff_A_XCzMfxRA7_0;
	wire w_dff_A_0pppbt6K3_0;
	wire w_dff_A_YQEDeZsF8_0;
	wire w_dff_A_zZCSepld7_0;
	wire w_dff_A_H5ZKYjVU1_0;
	wire w_dff_A_cItHHJ9M8_0;
	wire w_dff_A_Z1rwaf0c9_2;
	wire w_dff_A_lpEtMeBB0_0;
	wire w_dff_A_B7bR7plx4_0;
	wire w_dff_A_YPyXDQlB4_0;
	wire w_dff_A_GzCislSo9_0;
	wire w_dff_A_Pb6qYUgU2_0;
	wire w_dff_A_a0TWqPZN0_0;
	wire w_dff_A_8xeGaHK31_0;
	wire w_dff_A_Nt7mpm9u6_0;
	wire w_dff_A_YSmqPlh66_0;
	wire w_dff_A_8ieq2PLb4_0;
	wire w_dff_A_sIFMCCTq3_0;
	wire w_dff_A_y2NcQUqF0_0;
	wire w_dff_A_6eSmLkqc9_2;
	wire w_dff_A_T7rTPfZH9_0;
	wire w_dff_A_oEjHxI8S8_0;
	wire w_dff_A_6qtVXU9u7_0;
	wire w_dff_A_Dx5l8OnE5_0;
	wire w_dff_A_lFBGzwUw0_0;
	wire w_dff_A_wGNiJXX33_0;
	wire w_dff_A_8NSuVLOE6_0;
	wire w_dff_A_0fddDv9l5_0;
	wire w_dff_A_VWNEkdXj9_0;
	wire w_dff_A_GwCZjVlW8_0;
	wire w_dff_A_NKRZ3IAE1_0;
	wire w_dff_A_IllGmloY9_0;
	wire w_dff_A_m9AUuwwd7_0;
	wire w_dff_A_zlCQ34f47_2;
	wire w_dff_A_TKl59R6U4_0;
	wire w_dff_A_WFvjHIVR2_0;
	wire w_dff_A_9Br4c2dp0_0;
	wire w_dff_A_vWMPW1Se8_0;
	wire w_dff_A_ZFraZAjN7_0;
	wire w_dff_A_7AKyzm9g0_0;
	wire w_dff_A_SS5VBVme5_0;
	wire w_dff_A_4mf447Bi3_0;
	wire w_dff_A_ccXVZmas3_0;
	wire w_dff_A_eqDGjRQR7_0;
	wire w_dff_A_6KGopj4c3_0;
	wire w_dff_A_j3fEP8LP3_0;
	wire w_dff_A_pLJlfSJl1_0;
	wire w_dff_A_zwekv3fv4_2;
	wire w_dff_A_F8BJTSfE3_0;
	wire w_dff_A_U28oKJzG7_0;
	wire w_dff_A_Uk4V7U748_0;
	wire w_dff_A_ttxLDRdL0_0;
	wire w_dff_A_BUxHzEkm9_0;
	wire w_dff_A_P6c34Js75_0;
	wire w_dff_A_CfU4rOil8_0;
	wire w_dff_A_CzMeV7QN3_0;
	wire w_dff_A_p7Ss9eQc5_0;
	wire w_dff_A_F7DMAR7U6_0;
	wire w_dff_A_WNK5iPcp6_0;
	wire w_dff_A_N9fNAT5n7_0;
	wire w_dff_A_zxlsppAi9_0;
	wire w_dff_A_9DBGI9NS8_0;
	wire w_dff_A_QSz4wJVn0_0;
	wire w_dff_A_lCOwNbj03_1;
	wire w_dff_A_OIFj3G9A1_0;
	wire w_dff_A_84NcbFgo0_0;
	wire w_dff_A_JcCbx2fa8_0;
	wire w_dff_A_IM5fMFUJ7_0;
	wire w_dff_A_ZwGittOs1_0;
	wire w_dff_A_lZJniq0H2_0;
	wire w_dff_A_KbWepYJm3_0;
	wire w_dff_A_VkzE3nOL7_0;
	wire w_dff_A_8hSFBnCz5_0;
	wire w_dff_A_OmpXChON8_0;
	wire w_dff_A_dxJhnket5_0;
	wire w_dff_A_58HqTgeW2_0;
	wire w_dff_A_C2XFWLrw2_0;
	wire w_dff_A_IgVUFivB9_0;
	wire w_dff_A_r7VgIBJl5_0;
	wire w_dff_A_sj0YHAtv4_1;
	wire w_dff_A_fswTJykB5_0;
	wire w_dff_A_WgDcwJZP4_0;
	wire w_dff_A_4zcGyYSq2_0;
	wire w_dff_A_z3xdx7EG1_0;
	wire w_dff_A_aIMctxaR4_0;
	wire w_dff_A_XzhAvNwz3_0;
	wire w_dff_A_lgCtd7vg1_0;
	wire w_dff_A_wUbGZ0TX8_0;
	wire w_dff_A_Ff1ch4qe1_0;
	wire w_dff_A_diDwxWGV7_0;
	wire w_dff_A_98STIIH93_0;
	wire w_dff_A_DNtzr0o88_0;
	wire w_dff_A_VdMoBVek6_0;
	wire w_dff_A_0bAyuyYD7_0;
	wire w_dff_A_oYXvcS0d5_0;
	wire w_dff_A_pXJgTd7U2_1;
	wire w_dff_A_0fBnK0dk5_0;
	wire w_dff_A_9H6c9TZi2_0;
	wire w_dff_A_7qN883YS7_0;
	wire w_dff_A_xaVg0qhm5_0;
	wire w_dff_A_UJPSPG4S1_0;
	wire w_dff_A_qQNR8Vp26_0;
	wire w_dff_A_CuYlR7iv7_0;
	wire w_dff_A_ru4lMoYc5_0;
	wire w_dff_A_IwAN1f470_0;
	wire w_dff_A_qVHozKTM8_0;
	wire w_dff_A_wdN7iPWG9_0;
	wire w_dff_A_5GH4LxQw0_0;
	wire w_dff_A_zXAkUw0c5_0;
	wire w_dff_A_uIYyqE1Q1_2;
	wire w_dff_A_7lkjoFMC0_0;
	wire w_dff_A_hG3WFMBp7_0;
	wire w_dff_A_iFfG8cWD7_0;
	wire w_dff_A_PJaBNnYC8_0;
	wire w_dff_A_T2yxENLR8_0;
	wire w_dff_A_BFPRcEdi6_0;
	wire w_dff_A_7i4JzMTm0_2;
	wire w_dff_A_ICTlbeD93_0;
	wire w_dff_A_wNQsUtmF8_0;
	wire w_dff_A_A0q2JVHP4_0;
	wire w_dff_A_iKwEJnzs3_0;
	wire w_dff_A_tmynV1jm6_0;
	wire w_dff_A_BChzxR5r2_0;
	wire w_dff_A_vFD3QYLO8_0;
	wire w_dff_A_l7Tx6VIj5_0;
	wire w_dff_A_A4vaxYBV0_0;
	wire w_dff_A_DICIafTn4_2;
	wire w_dff_A_xKwUIsha4_0;
	wire w_dff_A_u4IoAXrO7_0;
	wire w_dff_A_epYqvhRU1_0;
	wire w_dff_A_6vaKIZ543_0;
	wire w_dff_A_MIboaQFw0_0;
	wire w_dff_A_NQVt2kRm1_2;
	wire w_dff_A_jlQjxoG41_0;
	wire w_dff_A_PmI2oesN5_0;
	wire w_dff_A_4Oh98sEY5_0;
	wire w_dff_A_OkWBMWSE1_0;
	wire w_dff_A_ROJaRKpT5_0;
	wire w_dff_A_lsQP0g3C9_0;
	wire w_dff_A_zAtxwbX66_0;
	wire w_dff_A_MsWlgwaZ9_0;
	wire w_dff_A_ZdlUvHA08_0;
	wire w_dff_A_L1Bufp9g1_2;
	wire w_dff_A_lRTJsLNs9_2;
	wire w_dff_A_9SRkHYKg9_0;
	wire w_dff_A_e3l2gwAl1_0;
	wire w_dff_A_2iq6fmuY0_0;
	wire w_dff_A_neslyGTD7_0;
	wire w_dff_A_lOWCjw8e4_0;
	wire w_dff_A_lnjGnJCt2_2;
	wire w_dff_A_Y5XLu9dj5_0;
	wire w_dff_A_eeanR2vx6_0;
	wire w_dff_A_tYVrD28B9_0;
	wire w_dff_A_1W460Dm57_0;
	wire w_dff_A_BoqqTkn33_0;
	wire w_dff_A_xQQoHkPH4_0;
	wire w_dff_A_8uxDTvgW9_2;
	wire w_dff_A_cPqXYTE18_0;
	wire w_dff_A_voLhiAm82_0;
	wire w_dff_A_YHGunLfs7_0;
	wire w_dff_A_AYxt9uhx6_0;
	wire w_dff_A_JMmm4y7s7_0;
	wire w_dff_A_R9QbWCVT7_0;
	wire w_dff_A_AdMTSGkd2_0;
	wire w_dff_A_msuIofH91_2;
	wire w_dff_A_e7NZZ9Jh9_0;
	wire w_dff_A_WxO82xC60_0;
	wire w_dff_A_Tgt3uhVB7_0;
	wire w_dff_A_3RsOgYAn2_0;
	wire w_dff_A_V2AhAh9a8_0;
	wire w_dff_A_YUlWv93S3_0;
	wire w_dff_A_WPyjfajw6_0;
	wire w_dff_A_6shXyOtb9_2;
	wire w_dff_A_TiDOOqkh8_0;
	wire w_dff_A_YJxM6Mt30_2;
	wire w_dff_A_nsAqMw0Q0_0;
	wire w_dff_A_FTUK2Itj9_0;
	wire w_dff_A_VslLU2ex9_2;
	wire w_dff_A_17APeLJc3_0;
	wire w_dff_A_Gea5GdIC6_0;
	wire w_dff_A_rdoQ9sAy9_0;
	wire w_dff_A_EI1P8NHh9_2;
	wire w_dff_A_iO4BboNG7_0;
	wire w_dff_A_dfsQFtzR5_0;
	wire w_dff_A_vjIvwJmK5_0;
	wire w_dff_A_zFFMkuIJ3_2;
	wire w_dff_A_hl6VS2nb8_0;
	wire w_dff_A_Ti57PiJS2_0;
	wire w_dff_A_iDKQ5rAz6_0;
	wire w_dff_A_ohqNHRVs4_0;
	wire w_dff_A_R3tk25Rf5_0;
	wire w_dff_A_X0BsDltY5_0;
	wire w_dff_A_gT28VCUj6_0;
	wire w_dff_A_T9Mmn4g16_0;
	wire w_dff_A_4O1nbhdD6_0;
	wire w_dff_A_64VC4QjV2_0;
	wire w_dff_A_jsPWeTfS2_0;
	wire w_dff_A_jO93Ve3B1_2;
	wire w_dff_A_OflSHxKU6_2;
	wire w_dff_A_ht6zsPW75_0;
	wire w_dff_A_wCB5TBIl1_0;
	wire w_dff_A_7hPEKW9R3_0;
	wire w_dff_A_dsbSATGu4_2;
	wire w_dff_A_j5V6LuLv2_0;
	wire w_dff_A_OxRSYCGE2_0;
	wire w_dff_A_ZEQWi1pg4_0;
	wire w_dff_A_FvQ315YE3_0;
	wire w_dff_A_ioHSf3dV1_0;
	wire w_dff_A_5LuU9lJA3_2;
	wire w_dff_A_qX5Ij0Hf0_0;
	wire w_dff_A_SnxBONCb1_0;
	wire w_dff_A_Tihw7pkO8_0;
	wire w_dff_A_zi8mZRj11_0;
	wire w_dff_A_J0dSgC1d3_0;
	wire w_dff_A_tQ3YGlOH2_2;
	wire w_dff_A_Wac1H6vR7_0;
	wire w_dff_A_igCfawJ90_0;
	wire w_dff_A_i7PZ4wdJ2_0;
	wire w_dff_A_hiKzcPEr7_0;
	wire w_dff_A_EPOat27B7_0;
	wire w_dff_A_Wc8PTM7X5_0;
	wire w_dff_A_w934NNeU9_0;
	wire w_dff_A_sgRaRusK5_2;
	wire w_dff_A_X25iMPm18_0;
	wire w_dff_A_nw7rdXuS5_0;
	wire w_dff_A_BuVOp8gI7_0;
	wire w_dff_A_scjVvCKs4_0;
	wire w_dff_A_ZhbkMa961_0;
	wire w_dff_A_bu91IbJi1_0;
	wire w_dff_A_9zik9Kzl7_0;
	wire w_dff_A_BoGFj39m3_0;
	wire w_dff_A_OnCKJ4yS2_0;
	wire w_dff_A_ByoYz9dA3_0;
	wire w_dff_A_fuIUMmUJ9_0;
	wire w_dff_A_NUSCYnwC6_0;
	wire w_dff_A_Tf9JfhOZ2_0;
	wire w_dff_A_0s1VMX2B6_2;
	wire w_dff_A_1dn7niiP8_2;
	wire w_dff_A_PDuO5PBw0_2;
	wire w_dff_A_UIpu50357_0;
	wire w_dff_A_a8GoUbFq1_0;
	wire w_dff_A_0X2mtHnC4_0;
	wire w_dff_A_RbZnUKx60_2;
	wire w_dff_A_u16L53ov1_0;
	wire w_dff_A_jJnlQ8lg5_0;
	wire w_dff_A_PKY98M205_0;
	wire w_dff_A_VtwlBwvj4_2;
	wire w_dff_A_MEGQYoZQ8_0;
	wire w_dff_A_e0IBh4tV4_0;
	wire w_dff_A_He7vKV3m7_0;
	wire w_dff_A_0T4TBg678_0;
	wire w_dff_A_xrNjMkcD4_0;
	wire w_dff_A_FgArA67l2_0;
	wire w_dff_A_Ctedzh3r6_0;
	wire w_dff_A_lSAJeN7r2_0;
	wire w_dff_A_LEpBkxa81_0;
	wire w_dff_A_cH5sdleA0_2;
	wire w_dff_A_09nyGtJ86_0;
	wire w_dff_A_8pW9M11I5_0;
	wire w_dff_A_48s4wDcE6_0;
	wire w_dff_A_fGvCaisU3_0;
	wire w_dff_A_BvwSno8Q0_0;
	wire w_dff_A_cZZqkUzd1_0;
	wire w_dff_A_bMJesM9S9_0;
	wire w_dff_A_RKJc31Ei8_0;
	wire w_dff_A_jvOeQbXp8_0;
	wire w_dff_A_j4XNgQ4z2_0;
	wire w_dff_A_lHS6djP02_2;
	wire w_dff_A_mzEkFAxW8_0;
	wire w_dff_A_80KpsHq41_0;
	wire w_dff_A_XU8B1wjo3_0;
	wire w_dff_A_YxbgDcVs8_0;
	wire w_dff_A_GbWXC90o2_0;
	wire w_dff_A_PKh5xbJl3_0;
	wire w_dff_A_YWOxOlqC7_0;
	wire w_dff_A_PgydrYl73_0;
	wire w_dff_A_c2mZSCEB2_0;
	wire w_dff_A_GtHIBI4h7_0;
	wire w_dff_A_qWsczlr09_0;
	wire w_dff_A_2DLI61aZ0_2;
	wire w_dff_A_ZOJQrSh79_0;
	wire w_dff_A_dg8uBm2T5_0;
	wire w_dff_A_itMerj1F4_0;
	wire w_dff_A_fY0orbjl7_0;
	wire w_dff_A_EyeXZHZR0_0;
	wire w_dff_A_XEzsvhyY0_0;
	wire w_dff_A_UpFqKMfv6_0;
	wire w_dff_A_PnLwTg464_0;
	wire w_dff_A_4B8VkiN93_0;
	wire w_dff_A_yxBdb8Hu6_0;
	wire w_dff_A_bYk42HNX2_0;
	wire w_dff_A_1HLKbfCP9_2;
	wire w_dff_A_wgtgLWZW8_0;
	wire w_dff_A_iEf537ix5_0;
	wire w_dff_A_Q5gWqtge2_0;
	wire w_dff_A_JQImtExa2_0;
	wire w_dff_A_NEAW4X7W2_0;
	wire w_dff_A_wfeRvzK13_0;
	wire w_dff_A_NqDqdmRB5_0;
	wire w_dff_A_z5Nuabmv8_0;
	wire w_dff_A_aUo2VDAg5_2;
	wire w_dff_A_TrFPIPHg7_0;
	wire w_dff_A_PcdDueST1_0;
	wire w_dff_A_y0LHmDNq4_0;
	wire w_dff_A_xkssh9pA4_0;
	wire w_dff_A_hYEXsSZI9_0;
	wire w_dff_A_1f6NTWTF5_0;
	wire w_dff_A_GLZYMKPX6_0;
	wire w_dff_A_usVh4LIi3_0;
	wire w_dff_A_6suMEec18_0;
	wire w_dff_A_19A0fWNC1_2;
	wire w_dff_A_zGb8EKUl8_0;
	wire w_dff_A_QsYMua8f1_0;
	wire w_dff_A_ak1EzYwz4_0;
	wire w_dff_A_EersNSW51_0;
	wire w_dff_A_i0DpshIC4_0;
	wire w_dff_A_3aRMGh4s6_0;
	wire w_dff_A_sClgRdwd5_0;
	wire w_dff_A_xEpmNJS08_0;
	wire w_dff_A_e2p8uiMa4_0;
	wire w_dff_A_aevorycp8_2;
	wire w_dff_A_1077YN5D5_0;
	wire w_dff_A_veBJKOnv9_0;
	wire w_dff_A_AShsLy0K8_0;
	wire w_dff_A_fzvrt9aG6_0;
	wire w_dff_A_GOgkxPyM9_0;
	wire w_dff_A_z5vZLAli4_0;
	wire w_dff_A_ojR4bByL9_0;
	wire w_dff_A_Ln9xXAqo0_0;
	wire w_dff_A_bMGOpfbj8_0;
	wire w_dff_A_LwVQP45A9_0;
	wire w_dff_A_BW82lTQW9_0;
	wire w_dff_A_AskpEjKv5_2;
	wire w_dff_A_hUBy5dZx3_0;
	wire w_dff_A_OOgoavvw0_0;
	wire w_dff_A_SIxhEd9F4_0;
	wire w_dff_A_QWCoSs815_0;
	wire w_dff_A_Gw55g2Xc2_2;
	wire w_dff_A_PQd8pTif0_0;
	wire w_dff_A_bDaYB5PH5_0;
	wire w_dff_A_sbLME52K2_0;
	wire w_dff_A_iuBjrNUP2_0;
	wire w_dff_A_RiPI1zBM8_0;
	wire w_dff_A_FwPipHHf7_0;
	wire w_dff_A_ECMPFZkm5_2;
	wire w_dff_A_zT6qpQjp6_0;
	wire w_dff_A_q19Fxxip4_0;
	wire w_dff_A_6gic20X58_0;
	wire w_dff_A_gOEE4jEb7_0;
	jnot g0000(.din(w_G15_0[2]),.dout(w_dff_A_7HM1DQ839_1),.clk(gclk));
	jor g0001(.dina(G57),.dinb(w_G5_1[2]),.dout(w_dff_A_OZMI4Ga77_2),.clk(gclk));
	jnot g0002(.din(G184),.dout(n317),.clk(gclk));
	jnot g0003(.din(G228),.dout(n318),.clk(gclk));
	jor g0004(.dina(n318),.dinb(n317),.dout(n319),.clk(gclk));
	jnot g0005(.din(G150),.dout(n320),.clk(gclk));
	jnot g0006(.din(G240),.dout(n321),.clk(gclk));
	jor g0007(.dina(n321),.dinb(n320),.dout(n322),.clk(gclk));
	jor g0008(.dina(n322),.dinb(n319),.dout(G404_fa_),.clk(gclk));
	jnot g0009(.din(G210),.dout(n324),.clk(gclk));
	jnot g0010(.din(G218),.dout(n325),.clk(gclk));
	jor g0011(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jnot g0012(.din(G152),.dout(n327),.clk(gclk));
	jnot g0013(.din(G230),.dout(n328),.clk(gclk));
	jor g0014(.dina(n328),.dinb(n327),.dout(n329),.clk(gclk));
	jor g0015(.dina(n329),.dinb(n326),.dout(G406_fa_),.clk(gclk));
	jnot g0016(.din(G183),.dout(n331),.clk(gclk));
	jnot g0017(.din(G185),.dout(n332),.clk(gclk));
	jor g0018(.dina(n332),.dinb(n331),.dout(n333),.clk(gclk));
	jnot g0019(.din(G182),.dout(n334),.clk(gclk));
	jnot g0020(.din(G186),.dout(n335),.clk(gclk));
	jor g0021(.dina(n335),.dinb(n334),.dout(n336),.clk(gclk));
	jor g0022(.dina(n336),.dinb(n333),.dout(G408_fa_),.clk(gclk));
	jnot g0023(.din(G172),.dout(n338),.clk(gclk));
	jnot g0024(.din(G188),.dout(n339),.clk(gclk));
	jor g0025(.dina(n339),.dinb(n338),.dout(n340),.clk(gclk));
	jnot g0026(.din(G162),.dout(n341),.clk(gclk));
	jnot g0027(.din(G199),.dout(n342),.clk(gclk));
	jor g0028(.dina(n342),.dinb(n341),.dout(n343),.clk(gclk));
	jor g0029(.dina(n343),.dinb(n340),.dout(G410_fa_),.clk(gclk));
	jnot g0030(.din(G1197),.dout(n345),.clk(gclk));
	jor g0031(.dina(w_n345_0[1]),.dinb(w_G5_1[1]),.dout(w_dff_A_uzDJ9L3F8_2),.clk(gclk));
	jnot g0032(.din(G133),.dout(n347),.clk(gclk));
	jnot g0033(.din(G134),.dout(n348),.clk(gclk));
	jor g0034(.dina(n348),.dinb(n347),.dout(n349),.clk(gclk));
	jor g0035(.dina(w_n349_0[1]),.dinb(w_G5_1[0]),.dout(w_dff_A_1X4oNfns3_2),.clk(gclk));
	jand g0036(.dina(G163),.dinb(w_G1_1[2]),.dout(w_dff_A_0VY9qskf0_2),.clk(gclk));
	jnot g0037(.din(w_G41_0[2]),.dout(n352),.clk(gclk));
	jor g0038(.dina(n352),.dinb(w_G18_58[2]),.dout(n353),.clk(gclk));
	jor g0039(.dina(w_n353_0[2]),.dinb(w_G3701_1[1]),.dout(n354),.clk(gclk));
	jnot g0040(.din(w_G18_58[1]),.dout(n355),.clk(gclk));
	jand g0041(.dina(w_G41_0[1]),.dinb(w_n355_26[1]),.dout(n356),.clk(gclk));
	jand g0042(.dina(w_G229_0[1]),.dinb(w_G18_58[0]),.dout(n357),.clk(gclk));
	jor g0043(.dina(n357),.dinb(w_n356_0[2]),.dout(n358),.clk(gclk));
	jand g0044(.dina(w_G3701_1[0]),.dinb(w_n355_26[0]),.dout(n359),.clk(gclk));
	jnot g0045(.din(w_n359_0[1]),.dout(n360),.clk(gclk));
	jor g0046(.dina(n360),.dinb(w_n358_0[1]),.dout(n361),.clk(gclk));
	jand g0047(.dina(n361),.dinb(w_n354_1[2]),.dout(n362),.clk(gclk));
	jxor g0048(.dina(w_n362_0[2]),.dinb(w_G4526_1[1]),.dout(w_dff_A_G6f97vGW1_2),.clk(gclk));
	jand g0049(.dina(w_G4528_0[2]),.dinb(w_G1496_0[2]),.dout(n364),.clk(gclk));
	jxor g0050(.dina(w_n364_0[1]),.dinb(w_G38_1[2]),.dout(n365),.clk(gclk));
	jnot g0051(.din(w_G3723_1[1]),.dout(n366),.clk(gclk));
	jand g0052(.dina(G235),.dinb(w_G18_57[2]),.dout(n367),.clk(gclk));
	jnot g0053(.din(n367),.dout(n368),.clk(gclk));
	jnot g0054(.din(G103),.dout(n369),.clk(gclk));
	jor g0055(.dina(n369),.dinb(w_G18_57[1]),.dout(n370),.clk(gclk));
	jand g0056(.dina(w_n370_0[1]),.dinb(n368),.dout(n371),.clk(gclk));
	jxor g0057(.dina(w_n371_1[1]),.dinb(w_n366_0[1]),.dout(n372),.clk(gclk));
	jand g0058(.dina(G236),.dinb(w_G18_57[0]),.dout(n373),.clk(gclk));
	jnot g0059(.din(n373),.dout(n374),.clk(gclk));
	jnot g0060(.din(G23),.dout(n375),.clk(gclk));
	jor g0061(.dina(n375),.dinb(w_G18_56[2]),.dout(n376),.clk(gclk));
	jand g0062(.dina(w_n376_0[1]),.dinb(n374),.dout(n377),.clk(gclk));
	jnot g0063(.din(w_n377_1[2]),.dout(n378),.clk(gclk));
	jxor g0064(.dina(n378),.dinb(w_G3717_2[1]),.dout(n379),.clk(gclk));
	jor g0065(.dina(w_n379_1[1]),.dinb(w_n372_1[2]),.dout(n380),.clk(gclk));
	jnot g0066(.din(w_G3711_1[1]),.dout(n381),.clk(gclk));
	jand g0067(.dina(G237),.dinb(w_G18_56[1]),.dout(n382),.clk(gclk));
	jnot g0068(.din(n382),.dout(n383),.clk(gclk));
	jnot g0069(.din(G26),.dout(n384),.clk(gclk));
	jor g0070(.dina(n384),.dinb(w_G18_56[0]),.dout(n385),.clk(gclk));
	jand g0071(.dina(w_n385_0[1]),.dinb(n383),.dout(n386),.clk(gclk));
	jxor g0072(.dina(w_n386_0[2]),.dinb(n381),.dout(n387),.clk(gclk));
	jnot g0073(.din(w_G4526_1[0]),.dout(n388),.clk(gclk));
	jnot g0074(.din(w_G3701_0[2]),.dout(n389),.clk(gclk));
	jand g0075(.dina(w_n356_0[1]),.dinb(w_n389_0[1]),.dout(n390),.clk(gclk));
	jnot g0076(.din(w_G229_0[0]),.dout(n391),.clk(gclk));
	jor g0077(.dina(n391),.dinb(w_n355_25[2]),.dout(n392),.clk(gclk));
	jand g0078(.dina(n392),.dinb(w_n353_0[1]),.dout(n393),.clk(gclk));
	jand g0079(.dina(w_n359_0[0]),.dinb(n393),.dout(n394),.clk(gclk));
	jor g0080(.dina(n394),.dinb(w_n390_1[1]),.dout(n395),.clk(gclk));
	jnot g0081(.din(w_G3705_2[1]),.dout(n396),.clk(gclk));
	jnot g0082(.din(G238),.dout(n397),.clk(gclk));
	jor g0083(.dina(n397),.dinb(w_n355_25[1]),.dout(n398),.clk(gclk));
	jnot g0084(.din(G29),.dout(n399),.clk(gclk));
	jor g0085(.dina(n399),.dinb(w_G18_55[2]),.dout(n400),.clk(gclk));
	jand g0086(.dina(w_n400_0[1]),.dinb(n398),.dout(n401),.clk(gclk));
	jxor g0087(.dina(w_n401_1[2]),.dinb(n396),.dout(n402),.clk(gclk));
	jor g0088(.dina(w_n402_1[1]),.dinb(w_n395_0[2]),.dout(n403),.clk(gclk));
	jor g0089(.dina(w_n403_0[1]),.dinb(w_n388_0[2]),.dout(n404),.clk(gclk));
	jor g0090(.dina(w_n404_0[1]),.dinb(w_n387_1[2]),.dout(n405),.clk(gclk));
	jor g0091(.dina(w_n405_0[2]),.dinb(w_n380_0[2]),.dout(n406),.clk(gclk));
	jor g0092(.dina(w_n386_0[1]),.dinb(w_G3711_1[0]),.dout(n407),.clk(gclk));
	jor g0093(.dina(w_n402_1[0]),.dinb(w_n354_1[1]),.dout(n408),.clk(gclk));
	jor g0094(.dina(w_n408_0[1]),.dinb(w_n387_1[1]),.dout(n409),.clk(gclk));
	jand g0095(.dina(n409),.dinb(w_n407_0[2]),.dout(n410),.clk(gclk));
	jor g0096(.dina(w_n410_0[1]),.dinb(w_n380_0[1]),.dout(n411),.clk(gclk));
	jor g0097(.dina(w_n401_1[1]),.dinb(w_G3705_2[0]),.dout(n412),.clk(gclk));
	jor g0098(.dina(w_n412_0[2]),.dinb(w_n387_1[0]),.dout(n413),.clk(gclk));
	jor g0099(.dina(w_n413_1[1]),.dinb(w_n380_0[0]),.dout(n414),.clk(gclk));
	jor g0100(.dina(w_n371_1[0]),.dinb(w_G3723_1[0]),.dout(n415),.clk(gclk));
	jand g0101(.dina(w_n371_0[2]),.dinb(w_G3723_0[2]),.dout(n416),.clk(gclk));
	jor g0102(.dina(w_n377_1[1]),.dinb(w_G3717_2[0]),.dout(n417),.clk(gclk));
	jor g0103(.dina(w_n417_0[2]),.dinb(n416),.dout(n418),.clk(gclk));
	jand g0104(.dina(n418),.dinb(n415),.dout(n419),.clk(gclk));
	jand g0105(.dina(w_n419_0[1]),.dinb(n414),.dout(n420),.clk(gclk));
	jand g0106(.dina(n420),.dinb(n411),.dout(n421),.clk(gclk));
	jand g0107(.dina(n421),.dinb(n406),.dout(n422),.clk(gclk));
	jnot g0108(.din(w_G3737_1[1]),.dout(n423),.clk(gclk));
	jand g0109(.dina(G233),.dinb(w_G18_55[1]),.dout(n424),.clk(gclk));
	jnot g0110(.din(n424),.dout(n425),.clk(gclk));
	jnot g0111(.din(G127),.dout(n426),.clk(gclk));
	jor g0112(.dina(n426),.dinb(w_G18_55[0]),.dout(n427),.clk(gclk));
	jand g0113(.dina(w_n427_0[1]),.dinb(n425),.dout(n428),.clk(gclk));
	jxor g0114(.dina(w_n428_0[2]),.dinb(n423),.dout(n429),.clk(gclk));
	jnot g0115(.din(w_G3729_1[1]),.dout(n430),.clk(gclk));
	jand g0116(.dina(G234),.dinb(w_G18_54[2]),.dout(n431),.clk(gclk));
	jnot g0117(.din(n431),.dout(n432),.clk(gclk));
	jnot g0118(.din(G130),.dout(n433),.clk(gclk));
	jor g0119(.dina(n433),.dinb(w_G18_54[1]),.dout(n434),.clk(gclk));
	jand g0120(.dina(w_n434_0[1]),.dinb(n432),.dout(n435),.clk(gclk));
	jxor g0121(.dina(w_n435_1[1]),.dinb(w_n430_0[1]),.dout(n436),.clk(gclk));
	jor g0122(.dina(w_n436_0[1]),.dinb(w_n429_2[1]),.dout(n437),.clk(gclk));
	jand g0123(.dina(G231),.dinb(w_G18_54[0]),.dout(n438),.clk(gclk));
	jnot g0124(.din(n438),.dout(n439),.clk(gclk));
	jnot g0125(.din(G100),.dout(n440),.clk(gclk));
	jor g0126(.dina(n440),.dinb(w_G18_53[2]),.dout(n441),.clk(gclk));
	jand g0127(.dina(w_n441_0[1]),.dinb(n439),.dout(n442),.clk(gclk));
	jor g0128(.dina(w_n442_0[2]),.dinb(w_G3749_1[1]),.dout(n443),.clk(gclk));
	jnot g0129(.din(w_n443_0[1]),.dout(n444),.clk(gclk));
	jand g0130(.dina(w_n442_0[1]),.dinb(w_G3749_1[0]),.dout(n445),.clk(gclk));
	jor g0131(.dina(w_n445_0[1]),.dinb(n444),.dout(n446),.clk(gclk));
	jand g0132(.dina(G232),.dinb(w_G18_53[1]),.dout(n447),.clk(gclk));
	jand g0133(.dina(G124),.dinb(w_n355_25[0]),.dout(n448),.clk(gclk));
	jor g0134(.dina(w_n448_0[1]),.dinb(n447),.dout(n449),.clk(gclk));
	jxor g0135(.dina(w_n449_0[2]),.dinb(w_G3743_1[2]),.dout(n450),.clk(gclk));
	jor g0136(.dina(w_n450_0[2]),.dinb(w_n446_1[1]),.dout(n451),.clk(gclk));
	jor g0137(.dina(n451),.dinb(w_n437_0[1]),.dout(n452),.clk(gclk));
	jor g0138(.dina(w_n452_0[1]),.dinb(w_n422_1[2]),.dout(n453),.clk(gclk));
	jnot g0139(.din(w_n449_0[1]),.dout(n454),.clk(gclk));
	jor g0140(.dina(w_n454_0[1]),.dinb(w_G3743_1[1]),.dout(n455),.clk(gclk));
	jand g0141(.dina(w_n454_0[0]),.dinb(w_G3743_1[0]),.dout(n456),.clk(gclk));
	jor g0142(.dina(w_n428_0[1]),.dinb(w_G3737_1[0]),.dout(n457),.clk(gclk));
	jor g0143(.dina(w_n435_1[0]),.dinb(w_G3729_1[0]),.dout(n458),.clk(gclk));
	jor g0144(.dina(w_n458_0[2]),.dinb(w_n429_2[0]),.dout(n459),.clk(gclk));
	jand g0145(.dina(n459),.dinb(w_n457_0[1]),.dout(n460),.clk(gclk));
	jor g0146(.dina(w_n460_0[2]),.dinb(w_n456_0[2]),.dout(n461),.clk(gclk));
	jand g0147(.dina(w_n461_0[1]),.dinb(w_n455_0[1]),.dout(n462),.clk(gclk));
	jand g0148(.dina(w_n462_0[2]),.dinb(w_n443_0[0]),.dout(n463),.clk(gclk));
	jor g0149(.dina(n463),.dinb(w_n445_0[0]),.dout(n464),.clk(gclk));
	jand g0150(.dina(w_n464_0[1]),.dinb(n453),.dout(n465),.clk(gclk));
	jnot g0151(.din(w_G4415_1[1]),.dout(n466),.clk(gclk));
	jand g0152(.dina(G223),.dinb(w_G18_53[0]),.dout(n467),.clk(gclk));
	jand g0153(.dina(G47),.dinb(w_n355_24[2]),.dout(n468),.clk(gclk));
	jor g0154(.dina(w_n468_0[1]),.dinb(n467),.dout(n469),.clk(gclk));
	jxor g0155(.dina(w_n469_1[1]),.dinb(w_n466_0[1]),.dout(n470),.clk(gclk));
	jnot g0156(.din(w_G4400_0[2]),.dout(n471),.clk(gclk));
	jand g0157(.dina(G226),.dinb(w_G18_52[2]),.dout(n472),.clk(gclk));
	jand g0158(.dina(G97),.dinb(w_n355_24[1]),.dout(n473),.clk(gclk));
	jor g0159(.dina(w_n473_0[1]),.dinb(n472),.dout(n474),.clk(gclk));
	jxor g0160(.dina(w_n474_1[1]),.dinb(w_n471_0[2]),.dout(n475),.clk(gclk));
	jand g0161(.dina(G217),.dinb(w_G18_52[1]),.dout(n476),.clk(gclk));
	jand g0162(.dina(G118),.dinb(w_n355_24[0]),.dout(n477),.clk(gclk));
	jor g0163(.dina(w_n477_0[1]),.dinb(n476),.dout(n478),.clk(gclk));
	jnot g0164(.din(w_n478_0[1]),.dout(n479),.clk(gclk));
	jxor g0165(.dina(w_n479_0[1]),.dinb(w_G4394_1[1]),.dout(n480),.clk(gclk));
	jand g0166(.dina(w_n480_1[1]),.dinb(w_n475_1[1]),.dout(n481),.clk(gclk));
	jnot g0167(.din(w_G4410_1[1]),.dout(n482),.clk(gclk));
	jand g0168(.dina(G224),.dinb(w_G18_52[0]),.dout(n483),.clk(gclk));
	jand g0169(.dina(G121),.dinb(w_n355_23[2]),.dout(n484),.clk(gclk));
	jor g0170(.dina(w_n484_0[1]),.dinb(n483),.dout(n485),.clk(gclk));
	jxor g0171(.dina(w_n485_0[2]),.dinb(w_n482_0[1]),.dout(n486),.clk(gclk));
	jand g0172(.dina(G225),.dinb(w_G18_51[2]),.dout(n487),.clk(gclk));
	jand g0173(.dina(G94),.dinb(w_n355_23[1]),.dout(n488),.clk(gclk));
	jor g0174(.dina(w_n488_0[1]),.dinb(n487),.dout(n489),.clk(gclk));
	jnot g0175(.din(w_n489_0[1]),.dout(n490),.clk(gclk));
	jxor g0176(.dina(w_n490_0[2]),.dinb(w_G4405_1[2]),.dout(n491),.clk(gclk));
	jand g0177(.dina(w_n491_1[1]),.dinb(w_n486_0[2]),.dout(n492),.clk(gclk));
	jand g0178(.dina(n492),.dinb(w_n481_0[2]),.dout(n493),.clk(gclk));
	jand g0179(.dina(w_n493_0[1]),.dinb(w_n470_0[2]),.dout(n494),.clk(gclk));
	jnot g0180(.din(w_n494_0[1]),.dout(n495),.clk(gclk));
	jor g0181(.dina(n495),.dinb(w_n465_0[2]),.dout(n496),.clk(gclk));
	jnot g0182(.din(w_n469_1[0]),.dout(n497),.clk(gclk));
	jand g0183(.dina(n497),.dinb(w_G4415_1[0]),.dout(n498),.clk(gclk));
	jand g0184(.dina(w_n469_0[2]),.dinb(w_n466_0[0]),.dout(n499),.clk(gclk));
	jnot g0185(.din(n499),.dout(n500),.clk(gclk));
	jand g0186(.dina(w_n485_0[1]),.dinb(w_n482_0[0]),.dout(n501),.clk(gclk));
	jnot g0187(.din(n501),.dout(n502),.clk(gclk));
	jnot g0188(.din(w_n485_0[0]),.dout(n503),.clk(gclk));
	jand g0189(.dina(w_n503_0[1]),.dinb(w_G4410_1[0]),.dout(n504),.clk(gclk));
	jand g0190(.dina(w_n490_0[1]),.dinb(w_G4405_1[1]),.dout(n505),.clk(gclk));
	jnot g0191(.din(w_n475_1[0]),.dout(n506),.clk(gclk));
	jor g0192(.dina(w_n479_0[0]),.dinb(w_G4394_1[0]),.dout(n507),.clk(gclk));
	jor g0193(.dina(w_n507_1[2]),.dinb(n506),.dout(n508),.clk(gclk));
	jand g0194(.dina(w_n474_1[0]),.dinb(w_n471_0[1]),.dout(n509),.clk(gclk));
	jnot g0195(.din(w_n509_0[1]),.dout(n510),.clk(gclk));
	jor g0196(.dina(w_n490_0[0]),.dinb(w_G4405_1[0]),.dout(n511),.clk(gclk));
	jand g0197(.dina(n511),.dinb(w_n510_0[1]),.dout(n512),.clk(gclk));
	jand g0198(.dina(w_n512_0[1]),.dinb(w_n508_0[1]),.dout(n513),.clk(gclk));
	jor g0199(.dina(n513),.dinb(w_n505_0[1]),.dout(n514),.clk(gclk));
	jor g0200(.dina(w_n514_0[2]),.dinb(n504),.dout(n515),.clk(gclk));
	jand g0201(.dina(n515),.dinb(w_n502_0[1]),.dout(n516),.clk(gclk));
	jand g0202(.dina(w_n516_0[2]),.dinb(n500),.dout(n517),.clk(gclk));
	jor g0203(.dina(n517),.dinb(n498),.dout(n518),.clk(gclk));
	jand g0204(.dina(w_n518_0[1]),.dinb(n496),.dout(n519),.clk(gclk));
	jnot g0205(.din(w_G4427_0[1]),.dout(n520),.clk(gclk));
	jand g0206(.dina(G221),.dinb(w_G18_51[1]),.dout(n521),.clk(gclk));
	jand g0207(.dina(G32),.dinb(w_n355_23[0]),.dout(n522),.clk(gclk));
	jor g0208(.dina(w_n522_0[1]),.dinb(n521),.dout(n523),.clk(gclk));
	jxor g0209(.dina(w_n523_0[2]),.dinb(w_n520_0[2]),.dout(n524),.clk(gclk));
	jnot g0210(.din(w_G4420_0[2]),.dout(n525),.clk(gclk));
	jand g0211(.dina(G222),.dinb(w_G18_51[0]),.dout(n526),.clk(gclk));
	jand g0212(.dina(G35),.dinb(w_n355_22[2]),.dout(n527),.clk(gclk));
	jor g0213(.dina(w_n527_0[1]),.dinb(n526),.dout(n528),.clk(gclk));
	jxor g0214(.dina(w_n528_1[1]),.dinb(w_n525_0[2]),.dout(n529),.clk(gclk));
	jand g0215(.dina(w_n529_0[1]),.dinb(w_n524_2[1]),.dout(n530),.clk(gclk));
	jnot g0216(.din(w_G4437_0[2]),.dout(n531),.clk(gclk));
	jand g0217(.dina(G219),.dinb(w_G18_50[2]),.dout(n532),.clk(gclk));
	jand g0218(.dina(G66),.dinb(w_n355_22[1]),.dout(n533),.clk(gclk));
	jor g0219(.dina(w_n533_0[1]),.dinb(n532),.dout(n534),.clk(gclk));
	jxor g0220(.dina(w_n534_1[1]),.dinb(w_n531_0[2]),.dout(n535),.clk(gclk));
	jnot g0221(.din(w_G4432_1[1]),.dout(n536),.clk(gclk));
	jand g0222(.dina(G220),.dinb(w_G18_50[1]),.dout(n537),.clk(gclk));
	jand g0223(.dina(G50),.dinb(w_n355_22[0]),.dout(n538),.clk(gclk));
	jor g0224(.dina(w_n538_0[1]),.dinb(n537),.dout(n539),.clk(gclk));
	jxor g0225(.dina(w_n539_1[1]),.dinb(w_n536_0[1]),.dout(n540),.clk(gclk));
	jand g0226(.dina(w_n540_0[2]),.dinb(w_n535_1[1]),.dout(n541),.clk(gclk));
	jand g0227(.dina(n541),.dinb(w_n530_0[1]),.dout(n542),.clk(gclk));
	jnot g0228(.din(w_n542_0[1]),.dout(n543),.clk(gclk));
	jor g0229(.dina(n543),.dinb(w_n519_0[1]),.dout(n544),.clk(gclk));
	jnot g0230(.din(w_n534_1[0]),.dout(n545),.clk(gclk));
	jand g0231(.dina(n545),.dinb(w_G4437_0[1]),.dout(n546),.clk(gclk));
	jnot g0232(.din(n546),.dout(n547),.clk(gclk));
	jand g0233(.dina(w_n534_0[2]),.dinb(w_n531_0[1]),.dout(n548),.clk(gclk));
	jand g0234(.dina(w_n539_1[0]),.dinb(w_n536_0[0]),.dout(n549),.clk(gclk));
	jnot g0235(.din(w_n539_0[2]),.dout(n550),.clk(gclk));
	jand g0236(.dina(n550),.dinb(w_G4432_1[0]),.dout(n551),.clk(gclk));
	jnot g0237(.din(w_n551_0[1]),.dout(n552),.clk(gclk));
	jand g0238(.dina(w_n523_0[1]),.dinb(w_n520_0[1]),.dout(n553),.clk(gclk));
	jand g0239(.dina(w_n528_1[0]),.dinb(w_n525_0[1]),.dout(n554),.clk(gclk));
	jand g0240(.dina(w_n554_0[2]),.dinb(w_n524_2[0]),.dout(n555),.clk(gclk));
	jor g0241(.dina(n555),.dinb(w_n553_0[1]),.dout(n556),.clk(gclk));
	jand g0242(.dina(w_n556_0[2]),.dinb(w_n552_0[1]),.dout(n557),.clk(gclk));
	jor g0243(.dina(w_n557_0[1]),.dinb(w_n549_0[1]),.dout(n558),.clk(gclk));
	jor g0244(.dina(w_n558_0[2]),.dinb(n548),.dout(n559),.clk(gclk));
	jand g0245(.dina(n559),.dinb(n547),.dout(n560),.clk(gclk));
	jnot g0246(.din(w_n560_0[1]),.dout(n561),.clk(gclk));
	jand g0247(.dina(n561),.dinb(n544),.dout(n562),.clk(gclk));
	jnot g0248(.din(w_G2236_1[1]),.dout(n563),.clk(gclk));
	jand g0249(.dina(G12),.dinb(G9),.dout(n564),.clk(gclk));
	jnot g0250(.din(w_n564_0[2]),.dout(n565),.clk(gclk));
	jor g0251(.dina(G157),.dinb(w_n355_21[2]),.dout(n566),.clk(gclk));
	jand g0252(.dina(n566),.dinb(w_n565_10[1]),.dout(n567),.clk(gclk));
	jxor g0253(.dina(w_n567_1[1]),.dinb(w_n563_0[1]),.dout(n568),.clk(gclk));
	jnot g0254(.din(w_G2218_0[2]),.dout(n569),.clk(gclk));
	jand g0255(.dina(G138),.dinb(w_n355_21[1]),.dout(n570),.clk(gclk));
	jand g0256(.dina(G160),.dinb(w_G18_50[0]),.dout(n571),.clk(gclk));
	jor g0257(.dina(n571),.dinb(w_n570_0[1]),.dout(n572),.clk(gclk));
	jxor g0258(.dina(w_n572_1[1]),.dinb(w_n569_0[2]),.dout(n573),.clk(gclk));
	jnot g0259(.din(w_G2211_0[2]),.dout(n574),.clk(gclk));
	jand g0260(.dina(G147),.dinb(w_n355_21[0]),.dout(n575),.clk(gclk));
	jand g0261(.dina(G151),.dinb(w_G18_49[2]),.dout(n576),.clk(gclk));
	jor g0262(.dina(n576),.dinb(w_n575_0[1]),.dout(n577),.clk(gclk));
	jxor g0263(.dina(w_n577_0[2]),.dinb(w_n574_0[1]),.dout(n578),.clk(gclk));
	jand g0264(.dina(w_n578_1[1]),.dinb(w_n573_1[1]),.dout(n579),.clk(gclk));
	jnot g0265(.din(w_G2230_1[1]),.dout(n580),.clk(gclk));
	jand g0266(.dina(G135),.dinb(w_n355_20[2]),.dout(n581),.clk(gclk));
	jand g0267(.dina(G158),.dinb(w_G18_49[1]),.dout(n582),.clk(gclk));
	jor g0268(.dina(n582),.dinb(w_n581_0[1]),.dout(n583),.clk(gclk));
	jxor g0269(.dina(w_n583_1[1]),.dinb(w_n580_0[1]),.dout(n584),.clk(gclk));
	jnot g0270(.din(w_G2224_1[1]),.dout(n585),.clk(gclk));
	jand g0271(.dina(G144),.dinb(w_n355_20[1]),.dout(n586),.clk(gclk));
	jand g0272(.dina(G159),.dinb(w_G18_49[0]),.dout(n587),.clk(gclk));
	jor g0273(.dina(n587),.dinb(w_n586_0[1]),.dout(n588),.clk(gclk));
	jxor g0274(.dina(w_n588_1[1]),.dinb(w_n585_0[1]),.dout(n589),.clk(gclk));
	jand g0275(.dina(w_n589_1[1]),.dinb(w_n584_0[2]),.dout(n590),.clk(gclk));
	jand g0276(.dina(n590),.dinb(w_n579_0[2]),.dout(n591),.clk(gclk));
	jand g0277(.dina(w_n591_0[1]),.dinb(w_n568_0[2]),.dout(n592),.clk(gclk));
	jnot g0278(.din(w_n592_0[1]),.dout(n593),.clk(gclk));
	jor g0279(.dina(n593),.dinb(w_n562_0[2]),.dout(n594),.clk(gclk));
	jand g0280(.dina(w_n567_1[0]),.dinb(w_n563_0[0]),.dout(n595),.clk(gclk));
	jnot g0281(.din(n595),.dout(n596),.clk(gclk));
	jnot g0282(.din(w_n567_0[2]),.dout(n597),.clk(gclk));
	jand g0283(.dina(n597),.dinb(w_G2236_1[0]),.dout(n598),.clk(gclk));
	jand g0284(.dina(w_n583_1[0]),.dinb(w_n580_0[0]),.dout(n599),.clk(gclk));
	jnot g0285(.din(w_n599_0[1]),.dout(n600),.clk(gclk));
	jnot g0286(.din(w_n583_0[2]),.dout(n601),.clk(gclk));
	jand g0287(.dina(n601),.dinb(w_G2230_1[0]),.dout(n602),.clk(gclk));
	jnot g0288(.din(w_n588_1[0]),.dout(n603),.clk(gclk));
	jand g0289(.dina(n603),.dinb(w_G2224_1[0]),.dout(n604),.clk(gclk));
	jnot g0290(.din(n604),.dout(n605),.clk(gclk));
	jand g0291(.dina(w_n577_0[1]),.dinb(w_n574_0[0]),.dout(n606),.clk(gclk));
	jand g0292(.dina(w_n606_1[2]),.dinb(w_n573_1[0]),.dout(n607),.clk(gclk));
	jand g0293(.dina(w_n572_1[0]),.dinb(w_n569_0[1]),.dout(n608),.clk(gclk));
	jand g0294(.dina(w_n588_0[2]),.dinb(w_n585_0[0]),.dout(n609),.clk(gclk));
	jor g0295(.dina(n609),.dinb(w_n608_0[2]),.dout(n610),.clk(gclk));
	jor g0296(.dina(w_n610_0[1]),.dinb(w_n607_0[1]),.dout(n611),.clk(gclk));
	jand g0297(.dina(n611),.dinb(w_n605_0[1]),.dout(n612),.clk(gclk));
	jnot g0298(.din(w_n612_0[1]),.dout(n613),.clk(gclk));
	jor g0299(.dina(w_n613_0[2]),.dinb(n602),.dout(n614),.clk(gclk));
	jand g0300(.dina(n614),.dinb(n600),.dout(n615),.clk(gclk));
	jor g0301(.dina(w_n615_1[1]),.dinb(n598),.dout(n616),.clk(gclk));
	jand g0302(.dina(n616),.dinb(n596),.dout(n617),.clk(gclk));
	jand g0303(.dina(w_n617_0[1]),.dinb(n594),.dout(n618),.clk(gclk));
	jnot g0304(.din(w_G2247_0[2]),.dout(n619),.clk(gclk));
	jor g0305(.dina(G155),.dinb(w_n355_20[0]),.dout(n620),.clk(gclk));
	jand g0306(.dina(w_n620_0[1]),.dinb(w_n565_10[0]),.dout(n621),.clk(gclk));
	jxor g0307(.dina(w_n621_0[2]),.dinb(w_n619_0[1]),.dout(n622),.clk(gclk));
	jnot g0308(.din(w_G2239_0[2]),.dout(n623),.clk(gclk));
	jor g0309(.dina(G156),.dinb(w_n355_19[2]),.dout(n624),.clk(gclk));
	jand g0310(.dina(w_n624_0[1]),.dinb(w_n565_9[2]),.dout(n625),.clk(gclk));
	jxor g0311(.dina(w_n625_0[2]),.dinb(w_n623_0[2]),.dout(n626),.clk(gclk));
	jand g0312(.dina(w_n626_0[1]),.dinb(w_n622_1[1]),.dout(n627),.clk(gclk));
	jnot g0313(.din(w_G2256_1[1]),.dout(n628),.clk(gclk));
	jor g0314(.dina(G153),.dinb(w_n355_19[1]),.dout(n629),.clk(gclk));
	jand g0315(.dina(w_n629_0[1]),.dinb(w_n565_9[1]),.dout(n630),.clk(gclk));
	jxor g0316(.dina(w_n630_0[2]),.dinb(w_n628_0[1]),.dout(n631),.clk(gclk));
	jnot g0317(.din(w_G2253_1[1]),.dout(n632),.clk(gclk));
	jor g0318(.dina(G154),.dinb(w_n355_19[0]),.dout(n633),.clk(gclk));
	jand g0319(.dina(w_n633_0[1]),.dinb(w_n565_9[0]),.dout(n634),.clk(gclk));
	jxor g0320(.dina(w_n634_0[2]),.dinb(w_n632_0[1]),.dout(n635),.clk(gclk));
	jand g0321(.dina(w_n635_0[2]),.dinb(w_n631_0[1]),.dout(n636),.clk(gclk));
	jand g0322(.dina(n636),.dinb(w_n627_0[1]),.dout(n637),.clk(gclk));
	jnot g0323(.din(w_n637_0[1]),.dout(n638),.clk(gclk));
	jor g0324(.dina(n638),.dinb(w_n618_0[2]),.dout(n639),.clk(gclk));
	jand g0325(.dina(w_n630_0[1]),.dinb(w_n628_0[0]),.dout(n640),.clk(gclk));
	jnot g0326(.din(n640),.dout(n641),.clk(gclk));
	jand g0327(.dina(w_n634_0[1]),.dinb(w_n632_0[0]),.dout(n642),.clk(gclk));
	jnot g0328(.din(w_n642_0[1]),.dout(n643),.clk(gclk));
	jand g0329(.dina(w_n621_0[1]),.dinb(w_n619_0[0]),.dout(n644),.clk(gclk));
	jand g0330(.dina(w_n625_0[1]),.dinb(w_n623_0[1]),.dout(n645),.clk(gclk));
	jand g0331(.dina(w_n645_0[2]),.dinb(w_n622_1[0]),.dout(n646),.clk(gclk));
	jor g0332(.dina(n646),.dinb(n644),.dout(n647),.clk(gclk));
	jnot g0333(.din(w_n647_0[1]),.dout(n648),.clk(gclk));
	jand g0334(.dina(w_n648_0[2]),.dinb(w_n643_0[1]),.dout(n649),.clk(gclk));
	jnot g0335(.din(w_n630_0[0]),.dout(n650),.clk(gclk));
	jand g0336(.dina(w_n650_0[1]),.dinb(w_G2256_1[0]),.dout(n651),.clk(gclk));
	jnot g0337(.din(w_n634_0[0]),.dout(n652),.clk(gclk));
	jand g0338(.dina(w_n652_0[1]),.dinb(w_G2253_1[0]),.dout(n653),.clk(gclk));
	jor g0339(.dina(w_n653_1[1]),.dinb(n651),.dout(n654),.clk(gclk));
	jor g0340(.dina(n654),.dinb(w_n649_0[1]),.dout(n655),.clk(gclk));
	jand g0341(.dina(n655),.dinb(n641),.dout(n656),.clk(gclk));
	jand g0342(.dina(w_n656_0[1]),.dinb(n639),.dout(n657),.clk(gclk));
	jnot g0343(.din(w_G1486_0[2]),.dout(n658),.clk(gclk));
	jor g0344(.dina(G213),.dinb(w_n355_18[2]),.dout(n659),.clk(gclk));
	jand g0345(.dina(w_n659_0[1]),.dinb(w_n565_8[2]),.dout(n660),.clk(gclk));
	jxor g0346(.dina(w_n660_1[1]),.dinb(w_n658_0[2]),.dout(n661),.clk(gclk));
	jnot g0347(.din(w_G1480_0[2]),.dout(n662),.clk(gclk));
	jor g0348(.dina(G214),.dinb(w_n355_18[1]),.dout(n663),.clk(gclk));
	jand g0349(.dina(w_n663_0[1]),.dinb(w_n565_8[1]),.dout(n664),.clk(gclk));
	jxor g0350(.dina(w_n664_1[1]),.dinb(w_n662_0[2]),.dout(n665),.clk(gclk));
	jnot g0351(.din(w_G106_1[1]),.dout(n666),.clk(gclk));
	jor g0352(.dina(G215),.dinb(w_n355_18[0]),.dout(n667),.clk(gclk));
	jand g0353(.dina(w_n667_0[1]),.dinb(w_n565_8[0]),.dout(n668),.clk(gclk));
	jxor g0354(.dina(w_n668_0[2]),.dinb(w_n666_0[1]),.dout(n669),.clk(gclk));
	jand g0355(.dina(w_n669_0[2]),.dinb(w_n665_0[2]),.dout(n670),.clk(gclk));
	jnot g0356(.din(w_G1469_1[1]),.dout(n671),.clk(gclk));
	jor g0357(.dina(G216),.dinb(w_n355_17[2]),.dout(n672),.clk(gclk));
	jand g0358(.dina(w_n672_0[1]),.dinb(w_n565_7[2]),.dout(n673),.clk(gclk));
	jxor g0359(.dina(w_n673_0[2]),.dinb(w_n671_0[1]),.dout(n674),.clk(gclk));
	jnot g0360(.din(w_G1462_0[2]),.dout(n675),.clk(gclk));
	jor g0361(.dina(G209),.dinb(w_n355_17[1]),.dout(n676),.clk(gclk));
	jand g0362(.dina(w_n676_0[1]),.dinb(w_n565_7[1]),.dout(n677),.clk(gclk));
	jxor g0363(.dina(w_n677_0[2]),.dinb(w_n675_0[2]),.dout(n678),.clk(gclk));
	jand g0364(.dina(w_n678_0[2]),.dinb(w_n674_1[1]),.dout(n679),.clk(gclk));
	jand g0365(.dina(w_n679_1[1]),.dinb(n670),.dout(n680),.clk(gclk));
	jand g0366(.dina(w_n680_0[1]),.dinb(w_n661_0[1]),.dout(n681),.clk(gclk));
	jnot g0367(.din(n681),.dout(n682),.clk(gclk));
	jor g0368(.dina(n682),.dinb(w_n657_1[1]),.dout(n683),.clk(gclk));
	jand g0369(.dina(w_n660_1[0]),.dinb(w_n658_0[1]),.dout(n684),.clk(gclk));
	jor g0370(.dina(w_n660_0[2]),.dinb(w_n658_0[0]),.dout(n685),.clk(gclk));
	jand g0371(.dina(w_n664_1[0]),.dinb(w_n662_0[1]),.dout(n686),.clk(gclk));
	jnot g0372(.din(w_n686_0[1]),.dout(n687),.clk(gclk));
	jor g0373(.dina(w_n664_0[2]),.dinb(w_n662_0[0]),.dout(n688),.clk(gclk));
	jand g0374(.dina(w_n668_0[1]),.dinb(w_n666_0[0]),.dout(n689),.clk(gclk));
	jnot g0375(.din(w_n668_0[0]),.dout(n690),.clk(gclk));
	jand g0376(.dina(w_n690_0[1]),.dinb(w_G106_1[0]),.dout(n691),.clk(gclk));
	jnot g0377(.din(n691),.dout(n692),.clk(gclk));
	jnot g0378(.din(w_n673_0[1]),.dout(n693),.clk(gclk));
	jand g0379(.dina(w_n693_0[1]),.dinb(w_G1469_1[0]),.dout(n694),.clk(gclk));
	jnot g0380(.din(n694),.dout(n695),.clk(gclk));
	jand g0381(.dina(w_n673_0[0]),.dinb(w_n671_0[0]),.dout(n696),.clk(gclk));
	jand g0382(.dina(w_n677_0[1]),.dinb(w_n675_0[1]),.dout(n697),.clk(gclk));
	jor g0383(.dina(w_n697_0[2]),.dinb(n696),.dout(n698),.clk(gclk));
	jand g0384(.dina(n698),.dinb(n695),.dout(n699),.clk(gclk));
	jand g0385(.dina(w_n699_1[1]),.dinb(w_n692_0[1]),.dout(n700),.clk(gclk));
	jor g0386(.dina(n700),.dinb(n689),.dout(n701),.clk(gclk));
	jand g0387(.dina(w_n701_1[1]),.dinb(n688),.dout(n702),.clk(gclk));
	jnot g0388(.din(n702),.dout(n703),.clk(gclk));
	jand g0389(.dina(w_n703_0[1]),.dinb(w_n687_0[1]),.dout(n704),.clk(gclk));
	jnot g0390(.din(w_n704_0[1]),.dout(n705),.clk(gclk));
	jand g0391(.dina(w_n705_0[1]),.dinb(n685),.dout(n706),.clk(gclk));
	jor g0392(.dina(n706),.dinb(n684),.dout(n707),.clk(gclk));
	jnot g0393(.din(w_n707_0[2]),.dout(n708),.clk(gclk));
	jand g0394(.dina(w_n708_0[1]),.dinb(w_n683_0[1]),.dout(n709),.clk(gclk));
	jnot g0395(.din(w_G38_1[1]),.dout(n710),.clk(gclk));
	jand g0396(.dina(w_G4528_0[1]),.dinb(w_G1492_1[1]),.dout(n711),.clk(gclk));
	jxor g0397(.dina(w_n711_0[1]),.dinb(w_n710_0[1]),.dout(n712),.clk(gclk));
	jnot g0398(.din(w_n712_0[1]),.dout(n713),.clk(gclk));
	jor g0399(.dina(w_n713_1[1]),.dinb(w_n709_1[1]),.dout(n714),.clk(gclk));
	jor g0400(.dina(w_n714_0[1]),.dinb(w_n365_0[1]),.dout(n715),.clk(gclk));
	jnot g0401(.din(w_n715_0[2]),.dout(n716),.clk(gclk));
	jnot g0402(.din(w_G1492_1[0]),.dout(n717),.clk(gclk));
	jnot g0403(.din(w_n364_0[0]),.dout(n718),.clk(gclk));
	jor g0404(.dina(n718),.dinb(n717),.dout(n719),.clk(gclk));
	jand g0405(.dina(n719),.dinb(w_G38_1[0]),.dout(n720),.clk(gclk));
	jor g0406(.dina(w_n720_1[1]),.dinb(w_n716_1[1]),.dout(w_dff_A_tmAqux6d0_2),.clk(gclk));
	jor g0407(.dina(G177),.dinb(w_n355_17[0]),.dout(n722),.clk(gclk));
	jand g0408(.dina(n722),.dinb(w_n565_7[0]),.dout(n723),.clk(gclk));
	jand g0409(.dina(w_G2236_0[2]),.dinb(w_G18_48[2]),.dout(n724),.clk(gclk));
	jnot g0410(.din(n724),.dout(n725),.clk(gclk));
	jor g0411(.dina(G64),.dinb(w_G18_48[1]),.dout(n726),.clk(gclk));
	jand g0412(.dina(n726),.dinb(n725),.dout(n727),.clk(gclk));
	jor g0413(.dina(w_n727_0[2]),.dinb(w_n723_0[2]),.dout(n728),.clk(gclk));
	jand g0414(.dina(G178),.dinb(w_G18_48[0]),.dout(n729),.clk(gclk));
	jor g0415(.dina(n729),.dinb(w_n581_0[0]),.dout(n730),.clk(gclk));
	jand g0416(.dina(w_G2230_0[2]),.dinb(w_G18_47[2]),.dout(n731),.clk(gclk));
	jnot g0417(.din(n731),.dout(n732),.clk(gclk));
	jor g0418(.dina(G85),.dinb(w_G18_47[1]),.dout(n733),.clk(gclk));
	jand g0419(.dina(n733),.dinb(n732),.dout(n734),.clk(gclk));
	jor g0420(.dina(w_n734_0[2]),.dinb(w_n730_0[2]),.dout(n735),.clk(gclk));
	jand g0421(.dina(G179),.dinb(w_G18_47[0]),.dout(n736),.clk(gclk));
	jor g0422(.dina(n736),.dinb(w_n586_0[0]),.dout(n737),.clk(gclk));
	jand g0423(.dina(w_G2224_0[2]),.dinb(w_G18_46[2]),.dout(n738),.clk(gclk));
	jnot g0424(.din(n738),.dout(n739),.clk(gclk));
	jor g0425(.dina(G84),.dinb(w_G18_46[1]),.dout(n740),.clk(gclk));
	jand g0426(.dina(n740),.dinb(n739),.dout(n741),.clk(gclk));
	jand g0427(.dina(w_n741_0[2]),.dinb(w_n737_0[2]),.dout(n742),.clk(gclk));
	jand g0428(.dina(G180),.dinb(w_G18_46[0]),.dout(n743),.clk(gclk));
	jor g0429(.dina(n743),.dinb(w_n570_0[0]),.dout(n744),.clk(gclk));
	jand g0430(.dina(w_G2218_0[1]),.dinb(w_G18_45[2]),.dout(n745),.clk(gclk));
	jnot g0431(.din(n745),.dout(n746),.clk(gclk));
	jor g0432(.dina(G83),.dinb(w_G18_45[1]),.dout(n747),.clk(gclk));
	jand g0433(.dina(n747),.dinb(n746),.dout(n748),.clk(gclk));
	jor g0434(.dina(w_n748_0[2]),.dinb(w_n744_0[2]),.dout(n749),.clk(gclk));
	jor g0435(.dina(w_n741_0[1]),.dinb(w_n737_0[1]),.dout(n750),.clk(gclk));
	jand g0436(.dina(n750),.dinb(n749),.dout(n751),.clk(gclk));
	jand g0437(.dina(w_n748_0[1]),.dinb(w_n744_0[1]),.dout(n752),.clk(gclk));
	jand g0438(.dina(G171),.dinb(w_G18_45[0]),.dout(n753),.clk(gclk));
	jor g0439(.dina(n753),.dinb(w_n575_0[0]),.dout(n754),.clk(gclk));
	jand g0440(.dina(w_G2211_0[1]),.dinb(w_G18_44[2]),.dout(n755),.clk(gclk));
	jnot g0441(.din(n755),.dout(n756),.clk(gclk));
	jor g0442(.dina(G65),.dinb(w_G18_44[1]),.dout(n757),.clk(gclk));
	jand g0443(.dina(n757),.dinb(n756),.dout(n758),.clk(gclk));
	jand g0444(.dina(w_n758_0[2]),.dinb(w_n754_0[2]),.dout(n759),.clk(gclk));
	jor g0445(.dina(w_n759_0[1]),.dinb(w_n752_0[1]),.dout(n760),.clk(gclk));
	jand g0446(.dina(n760),.dinb(w_n751_0[1]),.dout(n761),.clk(gclk));
	jor g0447(.dina(n761),.dinb(w_n742_0[1]),.dout(n762),.clk(gclk));
	jand g0448(.dina(n762),.dinb(w_n735_0[1]),.dout(n763),.clk(gclk));
	jand g0449(.dina(w_n734_0[1]),.dinb(w_n730_0[1]),.dout(n764),.clk(gclk));
	jand g0450(.dina(w_n727_0[1]),.dinb(w_n723_0[1]),.dout(n765),.clk(gclk));
	jor g0451(.dina(w_n765_0[1]),.dinb(w_n764_0[1]),.dout(n766),.clk(gclk));
	jor g0452(.dina(n766),.dinb(n763),.dout(n767),.clk(gclk));
	jand g0453(.dina(n767),.dinb(w_n728_0[1]),.dout(n768),.clk(gclk));
	jnot g0454(.din(w_n752_0[0]),.dout(n769),.clk(gclk));
	jand g0455(.dina(n769),.dinb(w_n735_0[0]),.dout(n770),.clk(gclk));
	jnot g0456(.din(w_n742_0[0]),.dout(n771),.clk(gclk));
	jnot g0457(.din(w_n759_0[0]),.dout(n772),.clk(gclk));
	jand g0458(.dina(n772),.dinb(n771),.dout(n773),.clk(gclk));
	jand g0459(.dina(n773),.dinb(n770),.dout(n774),.clk(gclk));
	jnot g0460(.din(w_n765_0[0]),.dout(n775),.clk(gclk));
	jor g0461(.dina(w_n758_0[1]),.dinb(w_n754_0[1]),.dout(n776),.clk(gclk));
	jand g0462(.dina(n776),.dinb(n775),.dout(n777),.clk(gclk));
	jnot g0463(.din(w_n764_0[0]),.dout(n778),.clk(gclk));
	jand g0464(.dina(n778),.dinb(w_n728_0[0]),.dout(n779),.clk(gclk));
	jand g0465(.dina(n779),.dinb(n777),.dout(n780),.clk(gclk));
	jand g0466(.dina(n780),.dinb(w_n751_0[0]),.dout(n781),.clk(gclk));
	jand g0467(.dina(n781),.dinb(n774),.dout(n782),.clk(gclk));
	jand g0468(.dina(G191),.dinb(w_G18_44[0]),.dout(n783),.clk(gclk));
	jor g0469(.dina(n783),.dinb(w_n522_0[0]),.dout(n784),.clk(gclk));
	jor g0470(.dina(G60),.dinb(w_G18_43[2]),.dout(n785),.clk(gclk));
	jor g0471(.dina(w_n520_0[0]),.dinb(w_n355_16[2]),.dout(n786),.clk(gclk));
	jand g0472(.dina(n786),.dinb(n785),.dout(n787),.clk(gclk));
	jxor g0473(.dina(w_n787_0[2]),.dinb(w_n784_0[2]),.dout(n788),.clk(gclk));
	jand g0474(.dina(G189),.dinb(w_G18_43[1]),.dout(n789),.clk(gclk));
	jor g0475(.dina(n789),.dinb(w_n533_0[0]),.dout(n790),.clk(gclk));
	jor g0476(.dina(G62),.dinb(w_G18_43[0]),.dout(n791),.clk(gclk));
	jor g0477(.dina(w_n531_0[0]),.dinb(w_n355_16[1]),.dout(n792),.clk(gclk));
	jand g0478(.dina(n792),.dinb(n791),.dout(n793),.clk(gclk));
	jxor g0479(.dina(w_n793_1[1]),.dinb(w_n790_1[1]),.dout(n794),.clk(gclk));
	jand g0480(.dina(n794),.dinb(n788),.dout(n795),.clk(gclk));
	jand g0481(.dina(G190),.dinb(w_G18_42[2]),.dout(n796),.clk(gclk));
	jor g0482(.dina(n796),.dinb(w_n538_0[0]),.dout(n797),.clk(gclk));
	jor g0483(.dina(G61),.dinb(w_G18_42[1]),.dout(n798),.clk(gclk));
	jand g0484(.dina(w_G4432_0[2]),.dinb(w_G18_42[0]),.dout(n799),.clk(gclk));
	jnot g0485(.din(n799),.dout(n800),.clk(gclk));
	jand g0486(.dina(n800),.dinb(n798),.dout(n801),.clk(gclk));
	jxor g0487(.dina(w_n801_1[1]),.dinb(w_n797_1[1]),.dout(n802),.clk(gclk));
	jand g0488(.dina(G192),.dinb(w_G18_41[2]),.dout(n803),.clk(gclk));
	jor g0489(.dina(n803),.dinb(w_n527_0[0]),.dout(n804),.clk(gclk));
	jor g0490(.dina(G79),.dinb(w_G18_41[1]),.dout(n805),.clk(gclk));
	jor g0491(.dina(w_n525_0[0]),.dinb(w_n355_16[0]),.dout(n806),.clk(gclk));
	jand g0492(.dina(n806),.dinb(n805),.dout(n807),.clk(gclk));
	jxor g0493(.dina(w_n807_0[2]),.dinb(w_n804_0[2]),.dout(n808),.clk(gclk));
	jand g0494(.dina(n808),.dinb(w_n802_0[1]),.dout(n809),.clk(gclk));
	jand g0495(.dina(n809),.dinb(w_n795_0[1]),.dout(n810),.clk(gclk));
	jand g0496(.dina(G196),.dinb(w_G18_41[0]),.dout(n811),.clk(gclk));
	jor g0497(.dina(n811),.dinb(w_n473_0[0]),.dout(n812),.clk(gclk));
	jor g0498(.dina(G78),.dinb(w_G18_40[2]),.dout(n813),.clk(gclk));
	jand g0499(.dina(w_G4400_0[1]),.dinb(w_G18_40[1]),.dout(n814),.clk(gclk));
	jnot g0500(.din(n814),.dout(n815),.clk(gclk));
	jand g0501(.dina(n815),.dinb(n813),.dout(n816),.clk(gclk));
	jor g0502(.dina(w_n816_0[2]),.dinb(w_n812_0[2]),.dout(n817),.clk(gclk));
	jand g0503(.dina(G195),.dinb(w_G18_40[0]),.dout(n818),.clk(gclk));
	jor g0504(.dina(n818),.dinb(w_n488_0[0]),.dout(n819),.clk(gclk));
	jor g0505(.dina(G59),.dinb(w_G18_39[2]),.dout(n820),.clk(gclk));
	jand g0506(.dina(w_G4405_0[2]),.dinb(w_G18_39[1]),.dout(n821),.clk(gclk));
	jnot g0507(.din(n821),.dout(n822),.clk(gclk));
	jand g0508(.dina(n822),.dinb(n820),.dout(n823),.clk(gclk));
	jor g0509(.dina(w_n823_0[2]),.dinb(w_n819_0[2]),.dout(n824),.clk(gclk));
	jand g0510(.dina(w_n824_0[1]),.dinb(w_n817_0[1]),.dout(n825),.clk(gclk));
	jand g0511(.dina(G187),.dinb(w_G18_39[0]),.dout(n826),.clk(gclk));
	jor g0512(.dina(n826),.dinb(w_n477_0[0]),.dout(n827),.clk(gclk));
	jor g0513(.dina(G77),.dinb(w_G18_38[2]),.dout(n828),.clk(gclk));
	jand g0514(.dina(w_G4394_0[2]),.dinb(w_G18_38[1]),.dout(n829),.clk(gclk));
	jnot g0515(.din(n829),.dout(n830),.clk(gclk));
	jand g0516(.dina(n830),.dinb(n828),.dout(n831),.clk(gclk));
	jand g0517(.dina(w_n831_0[2]),.dinb(w_n827_0[2]),.dout(n832),.clk(gclk));
	jnot g0518(.din(w_n832_0[1]),.dout(n833),.clk(gclk));
	jand g0519(.dina(w_n823_0[1]),.dinb(w_n819_0[1]),.dout(n834),.clk(gclk));
	jnot g0520(.din(w_n834_0[1]),.dout(n835),.clk(gclk));
	jand g0521(.dina(n835),.dinb(n833),.dout(n836),.clk(gclk));
	jand g0522(.dina(n836),.dinb(n825),.dout(n837),.clk(gclk));
	jand g0523(.dina(w_n816_0[1]),.dinb(w_n812_0[1]),.dout(n838),.clk(gclk));
	jnot g0524(.din(w_n838_0[1]),.dout(n839),.clk(gclk));
	jor g0525(.dina(w_n831_0[1]),.dinb(w_n827_0[1]),.dout(n840),.clk(gclk));
	jand g0526(.dina(n840),.dinb(n839),.dout(n841),.clk(gclk));
	jand g0527(.dina(G193),.dinb(w_G18_38[0]),.dout(n842),.clk(gclk));
	jor g0528(.dina(n842),.dinb(w_n468_0[0]),.dout(n843),.clk(gclk));
	jor g0529(.dina(G80),.dinb(w_G18_37[2]),.dout(n844),.clk(gclk));
	jand g0530(.dina(w_G4415_0[2]),.dinb(w_G18_37[1]),.dout(n845),.clk(gclk));
	jnot g0531(.din(n845),.dout(n846),.clk(gclk));
	jand g0532(.dina(n846),.dinb(n844),.dout(n847),.clk(gclk));
	jand g0533(.dina(w_n847_0[2]),.dinb(w_n843_0[2]),.dout(n848),.clk(gclk));
	jnot g0534(.din(w_n848_0[1]),.dout(n849),.clk(gclk));
	jand g0535(.dina(G194),.dinb(w_G18_37[0]),.dout(n850),.clk(gclk));
	jor g0536(.dina(n850),.dinb(w_n484_0[0]),.dout(n851),.clk(gclk));
	jor g0537(.dina(G81),.dinb(w_G18_36[2]),.dout(n852),.clk(gclk));
	jand g0538(.dina(w_G4410_0[2]),.dinb(w_G18_36[1]),.dout(n853),.clk(gclk));
	jnot g0539(.din(n853),.dout(n854),.clk(gclk));
	jand g0540(.dina(n854),.dinb(n852),.dout(n855),.clk(gclk));
	jor g0541(.dina(w_n855_0[2]),.dinb(w_n851_0[2]),.dout(n856),.clk(gclk));
	jand g0542(.dina(w_n856_0[1]),.dinb(n849),.dout(n857),.clk(gclk));
	jor g0543(.dina(w_n847_0[1]),.dinb(w_n843_0[1]),.dout(n858),.clk(gclk));
	jand g0544(.dina(w_n855_0[1]),.dinb(w_n851_0[1]),.dout(n859),.clk(gclk));
	jnot g0545(.din(w_n859_0[1]),.dout(n860),.clk(gclk));
	jand g0546(.dina(n860),.dinb(w_n858_0[2]),.dout(n861),.clk(gclk));
	jand g0547(.dina(n861),.dinb(n857),.dout(n862),.clk(gclk));
	jand g0548(.dina(n862),.dinb(n841),.dout(n863),.clk(gclk));
	jand g0549(.dina(n863),.dinb(n837),.dout(n864),.clk(gclk));
	jand g0550(.dina(w_n864_0[1]),.dinb(w_n810_0[2]),.dout(n865),.clk(gclk));
	jand g0551(.dina(G200),.dinb(w_G18_36[0]),.dout(n866),.clk(gclk));
	jnot g0552(.din(n866),.dout(n867),.clk(gclk));
	jand g0553(.dina(n867),.dinb(w_n441_0[0]),.dout(n868),.clk(gclk));
	jnot g0554(.din(n868),.dout(n869),.clk(gclk));
	jor g0555(.dina(G56),.dinb(w_G18_35[2]),.dout(n870),.clk(gclk));
	jand g0556(.dina(w_G3749_0[2]),.dinb(w_G18_35[1]),.dout(n871),.clk(gclk));
	jnot g0557(.din(n871),.dout(n872),.clk(gclk));
	jand g0558(.dina(n872),.dinb(n870),.dout(n873),.clk(gclk));
	jand g0559(.dina(w_n873_0[2]),.dinb(w_n869_0[2]),.dout(n874),.clk(gclk));
	jnot g0560(.din(w_n874_0[1]),.dout(n875),.clk(gclk));
	jnot g0561(.din(w_n427_0[0]),.dout(n876),.clk(gclk));
	jand g0562(.dina(G202),.dinb(w_G18_35[0]),.dout(n877),.clk(gclk));
	jor g0563(.dina(n877),.dinb(n876),.dout(n878),.clk(gclk));
	jor g0564(.dina(G54),.dinb(w_G18_34[2]),.dout(n879),.clk(gclk));
	jand g0565(.dina(w_G3737_0[2]),.dinb(w_G18_34[1]),.dout(n880),.clk(gclk));
	jnot g0566(.din(n880),.dout(n881),.clk(gclk));
	jand g0567(.dina(n881),.dinb(n879),.dout(n882),.clk(gclk));
	jor g0568(.dina(w_n882_0[2]),.dinb(w_n878_0[2]),.dout(n883),.clk(gclk));
	jand g0569(.dina(n883),.dinb(n875),.dout(n884),.clk(gclk));
	jand g0570(.dina(w_n882_0[1]),.dinb(w_n878_0[1]),.dout(n885),.clk(gclk));
	jnot g0571(.din(w_n885_0[1]),.dout(n886),.clk(gclk));
	jor g0572(.dina(w_n873_0[1]),.dinb(w_n869_0[1]),.dout(n887),.clk(gclk));
	jand g0573(.dina(w_n887_0[1]),.dinb(n886),.dout(n888),.clk(gclk));
	jand g0574(.dina(n888),.dinb(n884),.dout(n889),.clk(gclk));
	jand g0575(.dina(G201),.dinb(w_G18_34[0]),.dout(n890),.clk(gclk));
	jor g0576(.dina(n890),.dinb(w_n448_0[0]),.dout(n891),.clk(gclk));
	jor g0577(.dina(G55),.dinb(w_G18_33[2]),.dout(n892),.clk(gclk));
	jand g0578(.dina(w_G3743_0[2]),.dinb(w_G18_33[1]),.dout(n893),.clk(gclk));
	jnot g0579(.din(n893),.dout(n894),.clk(gclk));
	jand g0580(.dina(n894),.dinb(n892),.dout(n895),.clk(gclk));
	jxor g0581(.dina(w_n895_1[1]),.dinb(w_n891_1[1]),.dout(n896),.clk(gclk));
	jnot g0582(.din(w_n434_0[0]),.dout(n897),.clk(gclk));
	jand g0583(.dina(G203),.dinb(w_G18_33[0]),.dout(n898),.clk(gclk));
	jor g0584(.dina(n898),.dinb(n897),.dout(n899),.clk(gclk));
	jor g0585(.dina(G53),.dinb(w_G18_32[2]),.dout(n900),.clk(gclk));
	jor g0586(.dina(w_n430_0[0]),.dinb(w_n355_15[2]),.dout(n901),.clk(gclk));
	jand g0587(.dina(n901),.dinb(n900),.dout(n902),.clk(gclk));
	jxor g0588(.dina(w_n902_0[2]),.dinb(w_n899_0[2]),.dout(n903),.clk(gclk));
	jand g0589(.dina(n903),.dinb(w_n896_0[1]),.dout(n904),.clk(gclk));
	jand g0590(.dina(n904),.dinb(w_n889_0[1]),.dout(n905),.clk(gclk));
	jnot g0591(.din(w_n400_0[0]),.dout(n906),.clk(gclk));
	jand g0592(.dina(G207),.dinb(w_G18_32[1]),.dout(n907),.clk(gclk));
	jor g0593(.dina(n907),.dinb(n906),.dout(n908),.clk(gclk));
	jor g0594(.dina(G74),.dinb(w_G18_32[0]),.dout(n909),.clk(gclk));
	jand g0595(.dina(w_G3705_1[2]),.dinb(w_G18_31[2]),.dout(n910),.clk(gclk));
	jnot g0596(.din(n910),.dout(n911),.clk(gclk));
	jand g0597(.dina(n911),.dinb(n909),.dout(n912),.clk(gclk));
	jor g0598(.dina(w_n912_0[2]),.dinb(w_n908_0[2]),.dout(n913),.clk(gclk));
	jnot g0599(.din(w_n376_0[0]),.dout(n914),.clk(gclk));
	jand g0600(.dina(G205),.dinb(w_G18_31[1]),.dout(n915),.clk(gclk));
	jor g0601(.dina(n915),.dinb(n914),.dout(n916),.clk(gclk));
	jor g0602(.dina(G75),.dinb(w_G18_31[0]),.dout(n917),.clk(gclk));
	jand g0603(.dina(w_G3717_1[2]),.dinb(w_G18_30[2]),.dout(n918),.clk(gclk));
	jnot g0604(.din(n918),.dout(n919),.clk(gclk));
	jand g0605(.dina(n919),.dinb(n917),.dout(n920),.clk(gclk));
	jor g0606(.dina(w_n920_0[2]),.dinb(w_n916_0[2]),.dout(n921),.clk(gclk));
	jand g0607(.dina(w_n921_0[1]),.dinb(w_n913_0[1]),.dout(n922),.clk(gclk));
	jand g0608(.dina(w_n920_0[1]),.dinb(w_n916_0[1]),.dout(n923),.clk(gclk));
	jnot g0609(.din(w_n923_0[1]),.dout(n924),.clk(gclk));
	jnot g0610(.din(w_n385_0[0]),.dout(n925),.clk(gclk));
	jand g0611(.dina(G206),.dinb(w_G18_30[1]),.dout(n926),.clk(gclk));
	jor g0612(.dina(n926),.dinb(n925),.dout(n927),.clk(gclk));
	jor g0613(.dina(G76),.dinb(w_G18_30[0]),.dout(n928),.clk(gclk));
	jand g0614(.dina(w_G3711_0[2]),.dinb(w_G18_29[2]),.dout(n929),.clk(gclk));
	jnot g0615(.din(n929),.dout(n930),.clk(gclk));
	jand g0616(.dina(n930),.dinb(n928),.dout(n931),.clk(gclk));
	jor g0617(.dina(w_n931_0[2]),.dinb(w_n927_0[2]),.dout(n932),.clk(gclk));
	jand g0618(.dina(w_n932_0[1]),.dinb(n924),.dout(n933),.clk(gclk));
	jand g0619(.dina(n933),.dinb(n922),.dout(n934),.clk(gclk));
	jnot g0620(.din(w_G70_0[1]),.dout(n935),.clk(gclk));
	jand g0621(.dina(w_n935_0[1]),.dinb(w_n355_15[1]),.dout(n936),.clk(gclk));
	jnot g0622(.din(n936),.dout(n937),.clk(gclk));
	jor g0623(.dina(w_n937_0[1]),.dinb(w_G41_0[0]),.dout(n938),.clk(gclk));
	jand g0624(.dina(w_n937_0[0]),.dinb(w_n356_0[0]),.dout(n939),.clk(gclk));
	jnot g0625(.din(w_n939_0[1]),.dout(n940),.clk(gclk));
	jand g0626(.dina(n940),.dinb(G89),.dout(n941),.clk(gclk));
	jand g0627(.dina(n941),.dinb(n938),.dout(n942),.clk(gclk));
	jnot g0628(.din(w_n370_0[0]),.dout(n943),.clk(gclk));
	jand g0629(.dina(G204),.dinb(w_G18_29[1]),.dout(n944),.clk(gclk));
	jor g0630(.dina(n944),.dinb(n943),.dout(n945),.clk(gclk));
	jor g0631(.dina(G73),.dinb(w_G18_29[0]),.dout(n946),.clk(gclk));
	jor g0632(.dina(w_n366_0[0]),.dinb(w_n355_15[0]),.dout(n947),.clk(gclk));
	jand g0633(.dina(n947),.dinb(n946),.dout(n948),.clk(gclk));
	jxor g0634(.dina(w_n948_1[1]),.dinb(w_n945_1[1]),.dout(n949),.clk(gclk));
	jand g0635(.dina(w_n912_0[1]),.dinb(w_n908_0[1]),.dout(n950),.clk(gclk));
	jnot g0636(.din(w_n950_0[1]),.dout(n951),.clk(gclk));
	jand g0637(.dina(w_n931_0[1]),.dinb(w_n927_0[1]),.dout(n952),.clk(gclk));
	jnot g0638(.din(w_n952_0[1]),.dout(n953),.clk(gclk));
	jand g0639(.dina(n953),.dinb(n951),.dout(n954),.clk(gclk));
	jand g0640(.dina(n954),.dinb(n949),.dout(n955),.clk(gclk));
	jand g0641(.dina(n955),.dinb(n942),.dout(n956),.clk(gclk));
	jand g0642(.dina(n956),.dinb(n934),.dout(n957),.clk(gclk));
	jand g0643(.dina(w_n957_0[1]),.dinb(w_n905_0[2]),.dout(n958),.clk(gclk));
	jand g0644(.dina(n958),.dinb(w_n865_0[1]),.dout(n959),.clk(gclk));
	jand g0645(.dina(w_n807_0[1]),.dinb(w_n804_0[1]),.dout(n960),.clk(gclk));
	jand g0646(.dina(n960),.dinb(w_n802_0[0]),.dout(n961),.clk(gclk));
	jand g0647(.dina(n961),.dinb(w_n795_0[0]),.dout(n962),.clk(gclk));
	jand g0648(.dina(w_n793_1[0]),.dinb(w_n790_1[0]),.dout(n963),.clk(gclk));
	jand g0649(.dina(w_n787_0[1]),.dinb(w_n784_0[1]),.dout(n964),.clk(gclk));
	jand g0650(.dina(w_n801_1[0]),.dinb(w_n797_1[0]),.dout(n965),.clk(gclk));
	jor g0651(.dina(n965),.dinb(n964),.dout(n966),.clk(gclk));
	jor g0652(.dina(w_n793_0[2]),.dinb(w_n790_0[2]),.dout(n967),.clk(gclk));
	jor g0653(.dina(w_n801_0[2]),.dinb(w_n797_0[2]),.dout(n968),.clk(gclk));
	jand g0654(.dina(n968),.dinb(n967),.dout(n969),.clk(gclk));
	jand g0655(.dina(n969),.dinb(n966),.dout(n970),.clk(gclk));
	jor g0656(.dina(n970),.dinb(n963),.dout(n971),.clk(gclk));
	jor g0657(.dina(n971),.dinb(n962),.dout(n972),.clk(gclk));
	jand g0658(.dina(w_n832_0[0]),.dinb(w_n817_0[0]),.dout(n973),.clk(gclk));
	jor g0659(.dina(w_n838_0[0]),.dinb(w_n834_0[0]),.dout(n974),.clk(gclk));
	jor g0660(.dina(n974),.dinb(n973),.dout(n975),.clk(gclk));
	jand g0661(.dina(w_n858_0[1]),.dinb(w_n856_0[0]),.dout(n976),.clk(gclk));
	jand g0662(.dina(n976),.dinb(w_n824_0[0]),.dout(n977),.clk(gclk));
	jand g0663(.dina(n977),.dinb(n975),.dout(n978),.clk(gclk));
	jand g0664(.dina(w_n859_0[0]),.dinb(w_n858_0[0]),.dout(n979),.clk(gclk));
	jor g0665(.dina(n979),.dinb(w_n848_0[0]),.dout(n980),.clk(gclk));
	jor g0666(.dina(n980),.dinb(n978),.dout(n981),.clk(gclk));
	jand g0667(.dina(w_n981_0[1]),.dinb(w_n810_0[1]),.dout(n982),.clk(gclk));
	jor g0668(.dina(n982),.dinb(w_n972_0[1]),.dout(n983),.clk(gclk));
	jor g0669(.dina(n983),.dinb(n959),.dout(n984),.clk(gclk));
	jand g0670(.dina(n984),.dinb(w_n782_0[1]),.dout(n985),.clk(gclk));
	jor g0671(.dina(n985),.dinb(n768),.dout(n986),.clk(gclk));
	jor g0672(.dina(G173),.dinb(w_n355_14[2]),.dout(n987),.clk(gclk));
	jand g0673(.dina(w_n987_0[1]),.dinb(w_n565_6[2]),.dout(n988),.clk(gclk));
	jand g0674(.dina(w_G2256_0[2]),.dinb(w_G18_28[2]),.dout(n989),.clk(gclk));
	jnot g0675(.din(n989),.dout(n990),.clk(gclk));
	jor g0676(.dina(G110),.dinb(w_G18_28[1]),.dout(n991),.clk(gclk));
	jand g0677(.dina(n991),.dinb(n990),.dout(n992),.clk(gclk));
	jor g0678(.dina(w_n992_0[2]),.dinb(w_n988_0[2]),.dout(n993),.clk(gclk));
	jor g0679(.dina(G175),.dinb(w_n355_14[1]),.dout(n994),.clk(gclk));
	jand g0680(.dina(w_n994_0[1]),.dinb(w_n565_6[1]),.dout(n995),.clk(gclk));
	jand g0681(.dina(w_G2247_0[1]),.dinb(w_G18_28[0]),.dout(n996),.clk(gclk));
	jnot g0682(.din(n996),.dout(n997),.clk(gclk));
	jor g0683(.dina(G86),.dinb(w_G18_27[2]),.dout(n998),.clk(gclk));
	jand g0684(.dina(n998),.dinb(n997),.dout(n999),.clk(gclk));
	jand g0685(.dina(w_n999_0[2]),.dinb(w_n995_0[2]),.dout(n1000),.clk(gclk));
	jnot g0686(.din(w_n1000_0[1]),.dout(n1001),.clk(gclk));
	jand g0687(.dina(n1001),.dinb(w_n993_0[1]),.dout(n1002),.clk(gclk));
	jand g0688(.dina(w_n992_0[1]),.dinb(w_n988_0[1]),.dout(n1003),.clk(gclk));
	jnot g0689(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jor g0690(.dina(w_n999_0[1]),.dinb(w_n995_0[1]),.dout(n1005),.clk(gclk));
	jand g0691(.dina(n1005),.dinb(n1004),.dout(n1006),.clk(gclk));
	jand g0692(.dina(n1006),.dinb(n1002),.dout(n1007),.clk(gclk));
	jor g0693(.dina(G174),.dinb(w_n355_14[0]),.dout(n1008),.clk(gclk));
	jand g0694(.dina(w_n1008_0[1]),.dinb(w_n565_6[0]),.dout(n1009),.clk(gclk));
	jand g0695(.dina(w_G2253_0[2]),.dinb(w_G18_27[1]),.dout(n1010),.clk(gclk));
	jnot g0696(.din(n1010),.dout(n1011),.clk(gclk));
	jor g0697(.dina(G109),.dinb(w_G18_27[0]),.dout(n1012),.clk(gclk));
	jand g0698(.dina(n1012),.dinb(n1011),.dout(n1013),.clk(gclk));
	jxor g0699(.dina(w_n1013_1[1]),.dinb(w_n1009_1[1]),.dout(n1014),.clk(gclk));
	jor g0700(.dina(G176),.dinb(w_n355_13[2]),.dout(n1015),.clk(gclk));
	jand g0701(.dina(w_n1015_0[1]),.dinb(w_n565_5[2]),.dout(n1016),.clk(gclk));
	jor g0702(.dina(w_n623_0[0]),.dinb(w_n355_13[1]),.dout(n1017),.clk(gclk));
	jor g0703(.dina(G63),.dinb(w_G18_26[2]),.dout(n1018),.clk(gclk));
	jand g0704(.dina(n1018),.dinb(n1017),.dout(n1019),.clk(gclk));
	jxor g0705(.dina(w_n1019_0[2]),.dinb(w_n1016_0[2]),.dout(n1020),.clk(gclk));
	jand g0706(.dina(n1020),.dinb(w_n1014_0[1]),.dout(n1021),.clk(gclk));
	jand g0707(.dina(n1021),.dinb(w_n1007_0[1]),.dout(n1022),.clk(gclk));
	jand g0708(.dina(w_n1022_0[1]),.dinb(n986),.dout(n1023),.clk(gclk));
	jand g0709(.dina(w_n948_1[0]),.dinb(w_n945_1[0]),.dout(n1024),.clk(gclk));
	jor g0710(.dina(w_n950_0[0]),.dinb(w_n939_0[0]),.dout(n1025),.clk(gclk));
	jand g0711(.dina(w_n932_0[0]),.dinb(w_n913_0[0]),.dout(n1026),.clk(gclk));
	jand g0712(.dina(n1026),.dinb(n1025),.dout(n1027),.clk(gclk));
	jor g0713(.dina(w_n952_0[0]),.dinb(w_n923_0[0]),.dout(n1028),.clk(gclk));
	jor g0714(.dina(n1028),.dinb(n1027),.dout(n1029),.clk(gclk));
	jor g0715(.dina(w_n948_0[2]),.dinb(w_n945_0[2]),.dout(n1030),.clk(gclk));
	jand g0716(.dina(n1030),.dinb(w_n921_0[0]),.dout(n1031),.clk(gclk));
	jand g0717(.dina(n1031),.dinb(n1029),.dout(n1032),.clk(gclk));
	jor g0718(.dina(n1032),.dinb(n1024),.dout(n1033),.clk(gclk));
	jand g0719(.dina(w_n1033_0[1]),.dinb(w_n905_0[1]),.dout(n1034),.clk(gclk));
	jand g0720(.dina(w_n902_0[1]),.dinb(w_n899_0[1]),.dout(n1035),.clk(gclk));
	jand g0721(.dina(n1035),.dinb(w_n896_0[0]),.dout(n1036),.clk(gclk));
	jand g0722(.dina(n1036),.dinb(w_n889_0[0]),.dout(n1037),.clk(gclk));
	jand g0723(.dina(w_n895_1[0]),.dinb(w_n891_1[0]),.dout(n1038),.clk(gclk));
	jor g0724(.dina(n1038),.dinb(w_n885_0[0]),.dout(n1039),.clk(gclk));
	jor g0725(.dina(w_n895_0[2]),.dinb(w_n891_0[2]),.dout(n1040),.clk(gclk));
	jand g0726(.dina(n1040),.dinb(w_n887_0[0]),.dout(n1041),.clk(gclk));
	jand g0727(.dina(n1041),.dinb(n1039),.dout(n1042),.clk(gclk));
	jor g0728(.dina(n1042),.dinb(w_n874_0[0]),.dout(n1043),.clk(gclk));
	jor g0729(.dina(n1043),.dinb(n1037),.dout(n1044),.clk(gclk));
	jor g0730(.dina(w_n1044_0[1]),.dinb(n1034),.dout(n1045),.clk(gclk));
	jand g0731(.dina(w_n1022_0[0]),.dinb(w_n782_0[0]),.dout(n1046),.clk(gclk));
	jand g0732(.dina(n1046),.dinb(w_n865_0[0]),.dout(n1047),.clk(gclk));
	jand g0733(.dina(n1047),.dinb(n1045),.dout(n1048),.clk(gclk));
	jand g0734(.dina(w_n1019_0[1]),.dinb(w_n1016_0[1]),.dout(n1049),.clk(gclk));
	jand g0735(.dina(n1049),.dinb(w_n1014_0[0]),.dout(n1050),.clk(gclk));
	jand g0736(.dina(n1050),.dinb(w_n1007_0[0]),.dout(n1051),.clk(gclk));
	jand g0737(.dina(w_n1013_1[0]),.dinb(w_n1009_1[0]),.dout(n1052),.clk(gclk));
	jor g0738(.dina(n1052),.dinb(w_n1000_0[0]),.dout(n1053),.clk(gclk));
	jor g0739(.dina(w_n1013_0[2]),.dinb(w_n1009_0[2]),.dout(n1054),.clk(gclk));
	jand g0740(.dina(n1054),.dinb(w_n993_0[0]),.dout(n1055),.clk(gclk));
	jand g0741(.dina(n1055),.dinb(n1053),.dout(n1056),.clk(gclk));
	jor g0742(.dina(n1056),.dinb(w_n1003_0[0]),.dout(n1057),.clk(gclk));
	jor g0743(.dina(n1057),.dinb(n1051),.dout(n1058),.clk(gclk));
	jor g0744(.dina(n1058),.dinb(n1048),.dout(n1059),.clk(gclk));
	jor g0745(.dina(n1059),.dinb(n1023),.dout(n1060),.clk(gclk));
	jor g0746(.dina(G167),.dinb(w_n355_13[0]),.dout(n1061),.clk(gclk));
	jand g0747(.dina(w_n1061_0[2]),.dinb(w_n565_5[1]),.dout(n1062),.clk(gclk));
	jand g0748(.dina(w_G1480_0[1]),.dinb(w_G18_26[1]),.dout(n1063),.clk(gclk));
	jnot g0749(.din(n1063),.dout(n1064),.clk(gclk));
	jor g0750(.dina(G112),.dinb(w_G18_26[0]),.dout(n1065),.clk(gclk));
	jand g0751(.dina(n1065),.dinb(n1064),.dout(n1066),.clk(gclk));
	jor g0752(.dina(w_n1066_0[2]),.dinb(w_n1062_0[1]),.dout(n1067),.clk(gclk));
	jor g0753(.dina(G166),.dinb(w_n355_12[2]),.dout(n1068),.clk(gclk));
	jand g0754(.dina(w_n1068_0[1]),.dinb(w_n565_5[0]),.dout(n1069),.clk(gclk));
	jand g0755(.dina(w_G1486_0[1]),.dinb(w_G18_25[2]),.dout(n1070),.clk(gclk));
	jnot g0756(.din(n1070),.dout(n1071),.clk(gclk));
	jor g0757(.dina(G88),.dinb(w_G18_25[1]),.dout(n1072),.clk(gclk));
	jand g0758(.dina(n1072),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0759(.dina(w_n1073_0[2]),.dinb(w_n1069_0[1]),.dout(n1074),.clk(gclk));
	jand g0760(.dina(n1074),.dinb(n1067),.dout(n1075),.clk(gclk));
	jor g0761(.dina(G169),.dinb(w_n355_12[1]),.dout(n1076),.clk(gclk));
	jand g0762(.dina(w_n1076_0[1]),.dinb(w_n565_4[2]),.dout(n1077),.clk(gclk));
	jand g0763(.dina(w_G1469_0[2]),.dinb(w_G18_25[0]),.dout(n1078),.clk(gclk));
	jnot g0764(.din(n1078),.dout(n1079),.clk(gclk));
	jor g0765(.dina(G111),.dinb(w_G18_24[2]),.dout(n1080),.clk(gclk));
	jand g0766(.dina(n1080),.dinb(n1079),.dout(n1081),.clk(gclk));
	jor g0767(.dina(w_n1081_0[2]),.dinb(w_n1077_0[2]),.dout(n1082),.clk(gclk));
	jand g0768(.dina(w_G1462_0[1]),.dinb(w_G18_24[1]),.dout(n1083),.clk(gclk));
	jnot g0769(.din(n1083),.dout(n1084),.clk(gclk));
	jor g0770(.dina(G113),.dinb(w_G18_24[0]),.dout(n1085),.clk(gclk));
	jand g0771(.dina(n1085),.dinb(n1084),.dout(n1086),.clk(gclk));
	jor g0772(.dina(w_n1086_0[2]),.dinb(w_n565_4[1]),.dout(n1087),.clk(gclk));
	jand g0773(.dina(n1087),.dinb(w_n1082_0[1]),.dout(n1088),.clk(gclk));
	jand g0774(.dina(n1088),.dinb(w_n1075_0[1]),.dout(n1089),.clk(gclk));
	jand g0775(.dina(w_n1081_0[1]),.dinb(w_n1077_0[1]),.dout(n1090),.clk(gclk));
	jand g0776(.dina(w_n1086_0[1]),.dinb(w_n565_4[0]),.dout(n1091),.clk(gclk));
	jor g0777(.dina(n1091),.dinb(n1090),.dout(n1092),.clk(gclk));
	jnot g0778(.din(w_n1092_0[1]),.dout(n1093),.clk(gclk));
	jand g0779(.dina(w_n1066_0[1]),.dinb(w_n1062_0[0]),.dout(n1094),.clk(gclk));
	jor g0780(.dina(G168),.dinb(w_n355_12[0]),.dout(n1095),.clk(gclk));
	jand g0781(.dina(w_n1095_0[1]),.dinb(w_n565_3[2]),.dout(n1096),.clk(gclk));
	jand g0782(.dina(w_G106_0[2]),.dinb(w_G18_23[2]),.dout(n1097),.clk(gclk));
	jnot g0783(.din(n1097),.dout(n1098),.clk(gclk));
	jor g0784(.dina(G87),.dinb(w_G18_23[1]),.dout(n1099),.clk(gclk));
	jand g0785(.dina(n1099),.dinb(n1098),.dout(n1100),.clk(gclk));
	jand g0786(.dina(w_n1100_0[2]),.dinb(w_n1096_0[2]),.dout(n1101),.clk(gclk));
	jor g0787(.dina(n1101),.dinb(n1094),.dout(n1102),.clk(gclk));
	jnot g0788(.din(w_n1102_0[1]),.dout(n1103),.clk(gclk));
	jor g0789(.dina(w_n1100_0[1]),.dinb(w_n1096_0[1]),.dout(n1104),.clk(gclk));
	jand g0790(.dina(w_n1073_0[1]),.dinb(w_n1069_0[0]),.dout(n1105),.clk(gclk));
	jnot g0791(.din(w_n1105_0[1]),.dout(n1106),.clk(gclk));
	jand g0792(.dina(n1106),.dinb(w_n1104_0[1]),.dout(n1107),.clk(gclk));
	jand g0793(.dina(n1107),.dinb(n1103),.dout(n1108),.clk(gclk));
	jand g0794(.dina(n1108),.dinb(n1093),.dout(n1109),.clk(gclk));
	jand g0795(.dina(n1109),.dinb(n1089),.dout(n1110),.clk(gclk));
	jand g0796(.dina(n1110),.dinb(n1060),.dout(n1111),.clk(gclk));
	jand g0797(.dina(w_n1104_0[0]),.dinb(w_n1082_0[0]),.dout(n1112),.clk(gclk));
	jand g0798(.dina(n1112),.dinb(w_n1092_0[0]),.dout(n1113),.clk(gclk));
	jor g0799(.dina(n1113),.dinb(w_n1102_0[0]),.dout(n1114),.clk(gclk));
	jand g0800(.dina(n1114),.dinb(w_n1075_0[0]),.dout(n1115),.clk(gclk));
	jnot g0801(.din(w_G4528_0[0]),.dout(n1116),.clk(gclk));
	jor g0802(.dina(w_G2204_0[2]),.dinb(w_G1455_0[2]),.dout(n1117),.clk(gclk));
	jor g0803(.dina(n1117),.dinb(w_n1116_0[1]),.dout(n1118),.clk(gclk));
	jand g0804(.dina(n1118),.dinb(w_G38_0[2]),.dout(n1119),.clk(gclk));
	jor g0805(.dina(n1119),.dinb(w_n1105_0[0]),.dout(n1120),.clk(gclk));
	jor g0806(.dina(n1120),.dinb(n1115),.dout(n1121),.clk(gclk));
	jor g0807(.dina(n1121),.dinb(n1111),.dout(n1122),.clk(gclk));
	jand g0808(.dina(w_G2204_0[1]),.dinb(w_G1455_0[1]),.dout(n1123),.clk(gclk));
	jor g0809(.dina(w_n1116_0[0]),.dinb(w_G38_0[1]),.dout(n1124),.clk(gclk));
	jor g0810(.dina(n1124),.dinb(n1123),.dout(n1125),.clk(gclk));
	jand g0811(.dina(w_n1125_0[2]),.dinb(w_n1122_0[2]),.dout(w_dff_A_7bncmJrH1_2),.clk(gclk));
	jand g0812(.dina(w_n377_1[0]),.dinb(w_G3717_1[1]),.dout(n1127),.clk(gclk));
	jand g0813(.dina(w_n413_1[0]),.dinb(w_n410_0[0]),.dout(n1128),.clk(gclk));
	jor g0814(.dina(w_n1128_1[1]),.dinb(w_n1127_0[1]),.dout(n1129),.clk(gclk));
	jand g0815(.dina(n1129),.dinb(w_n417_0[1]),.dout(n1130),.clk(gclk));
	jor g0816(.dina(w_n405_0[1]),.dinb(w_n379_1[0]),.dout(n1131),.clk(gclk));
	jand g0817(.dina(n1131),.dinb(w_n1130_0[1]),.dout(n1132),.clk(gclk));
	jxor g0818(.dina(n1132),.dinb(w_n372_1[1]),.dout(w_dff_A_7SRXhOvO3_2),.clk(gclk));
	jand g0819(.dina(w_n1128_1[0]),.dinb(w_n405_0[0]),.dout(n1134),.clk(gclk));
	jxor g0820(.dina(n1134),.dinb(w_n379_0[2]),.dout(w_dff_A_ZxG7VkOx2_2),.clk(gclk));
	jand g0821(.dina(w_n408_0[0]),.dinb(w_n412_0[1]),.dout(n1136),.clk(gclk));
	jand g0822(.dina(w_n1136_0[1]),.dinb(w_n404_0[0]),.dout(n1137),.clk(gclk));
	jxor g0823(.dina(n1137),.dinb(w_n387_0[2]),.dout(w_dff_A_vdMi5oyR9_2),.clk(gclk));
	jor g0824(.dina(w_n395_0[1]),.dinb(w_n388_0[1]),.dout(n1139),.clk(gclk));
	jand g0825(.dina(n1139),.dinb(w_n354_1[0]),.dout(n1140),.clk(gclk));
	jxor g0826(.dina(n1140),.dinb(w_n402_0[2]),.dout(w_dff_A_UGZaqdrl9_2),.clk(gclk));
	jor g0827(.dina(w_n437_0[0]),.dinb(w_n422_1[1]),.dout(n1142),.clk(gclk));
	jor g0828(.dina(w_n1142_0[1]),.dinb(w_n456_0[1]),.dout(n1143),.clk(gclk));
	jand g0829(.dina(n1143),.dinb(w_n462_0[1]),.dout(n1144),.clk(gclk));
	jxor g0830(.dina(n1144),.dinb(w_n446_1[0]),.dout(w_dff_A_Z1rwaf0c9_2),.clk(gclk));
	jand g0831(.dina(w_n1142_0[0]),.dinb(w_n460_0[1]),.dout(n1146),.clk(gclk));
	jxor g0832(.dina(n1146),.dinb(w_n450_0[1]),.dout(w_dff_A_6eSmLkqc9_2),.clk(gclk));
	jand g0833(.dina(w_n435_0[2]),.dinb(w_G3729_0[2]),.dout(n1148),.clk(gclk));
	jor g0834(.dina(w_n1148_0[2]),.dinb(w_n422_1[0]),.dout(n1149),.clk(gclk));
	jand g0835(.dina(n1149),.dinb(w_n458_0[1]),.dout(n1150),.clk(gclk));
	jxor g0836(.dina(n1150),.dinb(w_n429_1[2]),.dout(w_dff_A_zlCQ34f47_2),.clk(gclk));
	jxor g0837(.dina(w_n436_0[0]),.dinb(w_n422_0[2]),.dout(w_dff_A_zwekv3fv4_2),.clk(gclk));
	jxor g0838(.dina(w_n583_0[1]),.dinb(w_n577_0[0]),.dout(n1153),.clk(gclk));
	jxor g0839(.dina(w_n588_0[1]),.dinb(w_n567_0[1]),.dout(n1154),.clk(gclk));
	jxor g0840(.dina(n1154),.dinb(w_n572_0[2]),.dout(n1155),.clk(gclk));
	jnot g0841(.din(w_n625_0[0]),.dout(n1156),.clk(gclk));
	jor g0842(.dina(w_n1156_0[1]),.dinb(w_n620_0[0]),.dout(n1157),.clk(gclk));
	jnot g0843(.din(w_n621_0[0]),.dout(n1158),.clk(gclk));
	jor g0844(.dina(w_n624_0[0]),.dinb(n1158),.dout(n1159),.clk(gclk));
	jand g0845(.dina(n1159),.dinb(n1157),.dout(n1160),.clk(gclk));
	jor g0846(.dina(w_n652_0[0]),.dinb(w_n629_0[0]),.dout(n1161),.clk(gclk));
	jor g0847(.dina(w_n633_0[0]),.dinb(w_n650_0[0]),.dout(n1162),.clk(gclk));
	jand g0848(.dina(n1162),.dinb(n1161),.dout(n1163),.clk(gclk));
	jxor g0849(.dina(n1163),.dinb(n1160),.dout(n1164),.clk(gclk));
	jnot g0850(.din(G141),.dout(n1165),.clk(gclk));
	jor g0851(.dina(n1165),.dinb(w_G18_23[0]),.dout(n1166),.clk(gclk));
	jnot g0852(.din(G161),.dout(n1167),.clk(gclk));
	jor g0853(.dina(n1167),.dinb(w_n355_11[2]),.dout(n1168),.clk(gclk));
	jand g0854(.dina(n1168),.dinb(w_n1166_0[1]),.dout(n1169),.clk(gclk));
	jxor g0855(.dina(n1169),.dinb(n1164),.dout(n1170),.clk(gclk));
	jxor g0856(.dina(n1170),.dinb(n1155),.dout(n1171),.clk(gclk));
	jxor g0857(.dina(n1171),.dinb(n1153),.dout(n1172),.clk(gclk));
	jand g0858(.dina(w_n565_3[1]),.dinb(w_G18_22[2]),.dout(n1173),.clk(gclk));
	jxor g0859(.dina(G212),.dinb(G211),.dout(n1174),.clk(gclk));
	jand g0860(.dina(n1174),.dinb(w_n1173_0[1]),.dout(n1175),.clk(gclk));
	jor g0861(.dina(w_n676_0[0]),.dinb(w_n564_0[1]),.dout(n1176),.clk(gclk));
	jnot g0862(.din(w_n659_0[0]),.dout(n1177),.clk(gclk));
	jand g0863(.dina(w_n664_0[1]),.dinb(n1177),.dout(n1178),.clk(gclk));
	jnot g0864(.din(w_n663_0[0]),.dout(n1179),.clk(gclk));
	jand g0865(.dina(n1179),.dinb(w_n660_0[1]),.dout(n1180),.clk(gclk));
	jor g0866(.dina(n1180),.dinb(n1178),.dout(n1181),.clk(gclk));
	jor g0867(.dina(w_n693_0[0]),.dinb(w_n667_0[0]),.dout(n1182),.clk(gclk));
	jor g0868(.dina(w_n672_0[0]),.dinb(w_n690_0[0]),.dout(n1183),.clk(gclk));
	jand g0869(.dina(n1183),.dinb(n1182),.dout(n1184),.clk(gclk));
	jxor g0870(.dina(n1184),.dinb(n1181),.dout(n1185),.clk(gclk));
	jxor g0871(.dina(n1185),.dinb(n1176),.dout(n1186),.clk(gclk));
	jxor g0872(.dina(n1186),.dinb(n1175),.dout(n1187),.clk(gclk));
	jand g0873(.dina(G239),.dinb(w_G18_22[1]),.dout(n1188),.clk(gclk));
	jand g0874(.dina(G44),.dinb(w_n355_11[1]),.dout(n1189),.clk(gclk));
	jor g0875(.dina(w_n1189_0[1]),.dinb(n1188),.dout(n1190),.clk(gclk));
	jxor g0876(.dina(w_n442_0[0]),.dinb(w_n428_0[0]),.dout(n1191),.clk(gclk));
	jxor g0877(.dina(w_n449_0[0]),.dinb(w_n435_0[1]),.dout(n1192),.clk(gclk));
	jxor g0878(.dina(n1192),.dinb(n1191),.dout(n1193),.clk(gclk));
	jxor g0879(.dina(n1193),.dinb(n1190),.dout(n1194),.clk(gclk));
	jxor g0880(.dina(w_n401_1[0]),.dinb(w_n371_0[1]),.dout(n1195),.clk(gclk));
	jxor g0881(.dina(n1195),.dinb(w_n377_0[2]),.dout(n1196),.clk(gclk));
	jxor g0882(.dina(w_n386_0[0]),.dinb(w_n358_0[0]),.dout(n1197),.clk(gclk));
	jxor g0883(.dina(n1197),.dinb(n1196),.dout(n1198),.clk(gclk));
	jxor g0884(.dina(n1198),.dinb(n1194),.dout(n1199),.clk(gclk));
	jxor g0885(.dina(w_n534_0[1]),.dinb(w_n523_0[0]),.dout(n1200),.clk(gclk));
	jxor g0886(.dina(w_n539_0[1]),.dinb(w_n528_0[2]),.dout(n1201),.clk(gclk));
	jxor g0887(.dina(n1201),.dinb(n1200),.dout(n1202),.clk(gclk));
	jxor g0888(.dina(n1202),.dinb(w_n503_0[0]),.dout(n1203),.clk(gclk));
	jand g0889(.dina(G227),.dinb(w_G18_22[0]),.dout(n1204),.clk(gclk));
	jand g0890(.dina(G115),.dinb(w_n355_11[0]),.dout(n1205),.clk(gclk));
	jor g0891(.dina(w_n1205_0[1]),.dinb(n1204),.dout(n1206),.clk(gclk));
	jxor g0892(.dina(w_n489_0[0]),.dinb(w_n478_0[0]),.dout(n1207),.clk(gclk));
	jxor g0893(.dina(n1207),.dinb(n1206),.dout(n1208),.clk(gclk));
	jxor g0894(.dina(w_n474_0[2]),.dinb(w_n469_0[1]),.dout(n1209),.clk(gclk));
	jxor g0895(.dina(n1209),.dinb(n1208),.dout(n1210),.clk(gclk));
	jxor g0896(.dina(n1210),.dinb(n1203),.dout(n1211),.clk(gclk));
	jor g0897(.dina(n1211),.dinb(n1199),.dout(n1212),.clk(gclk));
	jor g0898(.dina(n1212),.dinb(n1187),.dout(n1213),.clk(gclk));
	jor g0899(.dina(n1213),.dinb(n1172),.dout(G412_fa_),.clk(gclk));
	jxor g0900(.dina(w_n831_0[0]),.dinb(w_n823_0[0]),.dout(n1215),.clk(gclk));
	jxor g0901(.dina(w_n847_0[0]),.dinb(w_n816_0[0]),.dout(n1216),.clk(gclk));
	jxor g0902(.dina(n1216),.dinb(w_n855_0[0]),.dout(n1217),.clk(gclk));
	jxor g0903(.dina(w_n793_0[1]),.dinb(w_n787_0[0]),.dout(n1218),.clk(gclk));
	jxor g0904(.dina(w_n807_0[0]),.dinb(w_n801_0[1]),.dout(n1219),.clk(gclk));
	jxor g0905(.dina(n1219),.dinb(n1218),.dout(n1220),.clk(gclk));
	jor g0906(.dina(w_G4393_0[1]),.dinb(w_n355_10[2]),.dout(n1221),.clk(gclk));
	jnot g0907(.din(G58),.dout(n1222),.clk(gclk));
	jor g0908(.dina(n1222),.dinb(w_G18_21[2]),.dout(n1223),.clk(gclk));
	jand g0909(.dina(n1223),.dinb(n1221),.dout(n1224),.clk(gclk));
	jxor g0910(.dina(n1224),.dinb(n1220),.dout(n1225),.clk(gclk));
	jxor g0911(.dina(n1225),.dinb(n1217),.dout(n1226),.clk(gclk));
	jxor g0912(.dina(n1226),.dinb(n1215),.dout(n1227),.clk(gclk));
	jxor g0913(.dina(w_n389_0[0]),.dinb(w_G3698_0[1]),.dout(n1228),.clk(gclk));
	jor g0914(.dina(n1228),.dinb(w_n355_10[1]),.dout(n1229),.clk(gclk));
	jnot g0915(.din(w_G69_0[1]),.dout(n1230),.clk(gclk));
	jand g0916(.dina(w_n935_0[0]),.dinb(n1230),.dout(n1231),.clk(gclk));
	jand g0917(.dina(w_G70_0[0]),.dinb(w_G69_0[0]),.dout(n1232),.clk(gclk));
	jor g0918(.dina(n1232),.dinb(w_G18_21[1]),.dout(n1233),.clk(gclk));
	jor g0919(.dina(n1233),.dinb(n1231),.dout(n1234),.clk(gclk));
	jand g0920(.dina(n1234),.dinb(n1229),.dout(n1235),.clk(gclk));
	jxor g0921(.dina(n1235),.dinb(w_n912_0[0]),.dout(n1236),.clk(gclk));
	jnot g0922(.din(w_n1236_0[1]),.dout(n1237),.clk(gclk));
	jxor g0923(.dina(w_n948_0[1]),.dinb(w_n931_0[0]),.dout(n1238),.clk(gclk));
	jnot g0924(.din(w_n920_0[0]),.dout(n1239),.clk(gclk));
	jxor g0925(.dina(w_n882_0[0]),.dinb(w_n873_0[0]),.dout(n1240),.clk(gclk));
	jxor g0926(.dina(w_n902_0[0]),.dinb(w_n895_0[1]),.dout(n1241),.clk(gclk));
	jxor g0927(.dina(n1241),.dinb(n1240),.dout(n1242),.clk(gclk));
	jxor g0928(.dina(n1242),.dinb(n1239),.dout(n1243),.clk(gclk));
	jxor g0929(.dina(n1243),.dinb(n1238),.dout(n1244),.clk(gclk));
	jnot g0930(.din(w_n1244_0[1]),.dout(n1245),.clk(gclk));
	jand g0931(.dina(n1245),.dinb(n1237),.dout(n1246),.clk(gclk));
	jand g0932(.dina(w_n1244_0[0]),.dinb(w_n1236_0[0]),.dout(n1247),.clk(gclk));
	jor g0933(.dina(w_G1459_0[1]),.dinb(w_n355_10[0]),.dout(n1248),.clk(gclk));
	jnot g0934(.din(G114),.dout(n1249),.clk(gclk));
	jor g0935(.dina(n1249),.dinb(w_G18_21[0]),.dout(n1250),.clk(gclk));
	jand g0936(.dina(n1250),.dinb(n1248),.dout(n1251),.clk(gclk));
	jxor g0937(.dina(w_n1086_0[0]),.dinb(w_n1081_0[0]),.dout(n1252),.clk(gclk));
	jxor g0938(.dina(n1252),.dinb(n1251),.dout(n1253),.clk(gclk));
	jxor g0939(.dina(w_n1100_0[0]),.dinb(w_n1073_0[0]),.dout(n1254),.clk(gclk));
	jxor g0940(.dina(n1254),.dinb(w_n1066_0[0]),.dout(n1255),.clk(gclk));
	jxor g0941(.dina(w_G1496_0[1]),.dinb(w_G1492_0[2]),.dout(n1256),.clk(gclk));
	jor g0942(.dina(n1256),.dinb(w_n355_9[2]),.dout(n1257),.clk(gclk));
	jxor g0943(.dina(w_G2204_0[0]),.dinb(w_G1455_0[0]),.dout(n1258),.clk(gclk));
	jor g0944(.dina(n1258),.dinb(w_G18_20[2]),.dout(n1259),.clk(gclk));
	jand g0945(.dina(n1259),.dinb(n1257),.dout(n1260),.clk(gclk));
	jxor g0946(.dina(n1260),.dinb(n1255),.dout(n1261),.clk(gclk));
	jxor g0947(.dina(n1261),.dinb(n1253),.dout(n1262),.clk(gclk));
	jxor g0948(.dina(w_n999_0[0]),.dinb(w_n992_0[0]),.dout(n1263),.clk(gclk));
	jxor g0949(.dina(w_n1019_0[0]),.dinb(w_n1013_0[1]),.dout(n1264),.clk(gclk));
	jxor g0950(.dina(n1264),.dinb(n1263),.dout(n1265),.clk(gclk));
	jxor g0951(.dina(n1265),.dinb(w_n727_0[0]),.dout(n1266),.clk(gclk));
	jor g0952(.dina(w_G2208_0[1]),.dinb(w_n355_9[1]),.dout(n1267),.clk(gclk));
	jnot g0953(.din(G82),.dout(n1268),.clk(gclk));
	jor g0954(.dina(n1268),.dinb(w_G18_20[1]),.dout(n1269),.clk(gclk));
	jand g0955(.dina(n1269),.dinb(n1267),.dout(n1270),.clk(gclk));
	jxor g0956(.dina(w_n758_0[0]),.dinb(w_n748_0[0]),.dout(n1271),.clk(gclk));
	jxor g0957(.dina(n1271),.dinb(n1270),.dout(n1272),.clk(gclk));
	jxor g0958(.dina(w_n741_0[0]),.dinb(w_n734_0[0]),.dout(n1273),.clk(gclk));
	jxor g0959(.dina(n1273),.dinb(n1272),.dout(n1274),.clk(gclk));
	jxor g0960(.dina(n1274),.dinb(n1266),.dout(n1275),.clk(gclk));
	jor g0961(.dina(n1275),.dinb(n1262),.dout(n1276),.clk(gclk));
	jor g0962(.dina(n1276),.dinb(n1247),.dout(n1277),.clk(gclk));
	jor g0963(.dina(n1277),.dinb(n1246),.dout(n1278),.clk(gclk));
	jor g0964(.dina(n1278),.dinb(n1227),.dout(G414_fa_),.clk(gclk));
	jnot g0965(.din(w_n1061_0[1]),.dout(n1280),.clk(gclk));
	jnot g0966(.din(G170),.dout(n1281),.clk(gclk));
	jand g0967(.dina(n1281),.dinb(w_G18_20[0]),.dout(n1282),.clk(gclk));
	jxor g0968(.dina(n1282),.dinb(w_n1068_0[0]),.dout(n1283),.clk(gclk));
	jnot g0969(.din(w_n1283_0[1]),.dout(n1284),.clk(gclk));
	jand g0970(.dina(n1284),.dinb(n1280),.dout(n1285),.clk(gclk));
	jand g0971(.dina(w_n1283_0[0]),.dinb(w_n1061_0[0]),.dout(n1286),.clk(gclk));
	jor g0972(.dina(n1286),.dinb(w_n564_0[0]),.dout(n1287),.clk(gclk));
	jor g0973(.dina(n1287),.dinb(n1285),.dout(n1288),.clk(gclk));
	jnot g0974(.din(w_n1077_0[0]),.dout(n1289),.clk(gclk));
	jor g0975(.dina(w_n1095_0[0]),.dinb(n1289),.dout(n1290),.clk(gclk));
	jnot g0976(.din(w_n1096_0[0]),.dout(n1291),.clk(gclk));
	jor g0977(.dina(n1291),.dinb(w_n1076_0[0]),.dout(n1292),.clk(gclk));
	jand g0978(.dina(n1292),.dinb(n1290),.dout(n1293),.clk(gclk));
	jxor g0979(.dina(G165),.dinb(G164),.dout(n1294),.clk(gclk));
	jand g0980(.dina(n1294),.dinb(w_n1173_0[0]),.dout(n1295),.clk(gclk));
	jxor g0981(.dina(n1295),.dinb(n1293),.dout(n1296),.clk(gclk));
	jxor g0982(.dina(n1296),.dinb(n1288),.dout(n1297),.clk(gclk));
	jxor g0983(.dina(w_n790_0[1]),.dinb(w_n784_0[0]),.dout(n1298),.clk(gclk));
	jxor g0984(.dina(w_n804_0[0]),.dinb(w_n797_0[1]),.dout(n1299),.clk(gclk));
	jxor g0985(.dina(n1299),.dinb(n1298),.dout(n1300),.clk(gclk));
	jxor g0986(.dina(n1300),.dinb(w_n851_0[0]),.dout(n1301),.clk(gclk));
	jand g0987(.dina(G197),.dinb(w_G18_19[2]),.dout(n1302),.clk(gclk));
	jor g0988(.dina(n1302),.dinb(w_n1205_0[0]),.dout(n1303),.clk(gclk));
	jnot g0989(.din(n1303),.dout(n1304),.clk(gclk));
	jxor g0990(.dina(w_n827_0[0]),.dinb(w_n819_0[0]),.dout(n1305),.clk(gclk));
	jxor g0991(.dina(n1305),.dinb(n1304),.dout(n1306),.clk(gclk));
	jnot g0992(.din(n1306),.dout(n1307),.clk(gclk));
	jxor g0993(.dina(w_n843_0[0]),.dinb(w_n812_0[0]),.dout(n1308),.clk(gclk));
	jxor g0994(.dina(n1308),.dinb(n1307),.dout(n1309),.clk(gclk));
	jand g0995(.dina(w_n1309_0[1]),.dinb(w_n1301_0[1]),.dout(n1310),.clk(gclk));
	jor g0996(.dina(n1310),.dinb(n1297),.dout(n1311),.clk(gclk));
	jand g0997(.dina(G208),.dinb(w_G18_19[1]),.dout(n1312),.clk(gclk));
	jor g0998(.dina(n1312),.dinb(w_n1189_0[0]),.dout(n1313),.clk(gclk));
	jxor g0999(.dina(w_n878_0[0]),.dinb(w_n869_0[0]),.dout(n1314),.clk(gclk));
	jxor g1000(.dina(w_n899_0[0]),.dinb(w_n891_0[1]),.dout(n1315),.clk(gclk));
	jxor g1001(.dina(n1315),.dinb(n1314),.dout(n1316),.clk(gclk));
	jxor g1002(.dina(n1316),.dinb(n1313),.dout(n1317),.clk(gclk));
	jnot g1003(.din(w_n916_0[0]),.dout(n1318),.clk(gclk));
	jxor g1004(.dina(w_n945_0[1]),.dinb(w_n927_0[0]),.dout(n1319),.clk(gclk));
	jxor g1005(.dina(n1319),.dinb(n1318),.dout(n1320),.clk(gclk));
	jnot g1006(.din(G198),.dout(n1321),.clk(gclk));
	jor g1007(.dina(n1321),.dinb(w_n355_9[0]),.dout(n1322),.clk(gclk));
	jand g1008(.dina(n1322),.dinb(w_n353_0[0]),.dout(n1323),.clk(gclk));
	jxor g1009(.dina(n1323),.dinb(w_n908_0[0]),.dout(n1324),.clk(gclk));
	jxor g1010(.dina(n1324),.dinb(n1320),.dout(n1325),.clk(gclk));
	jand g1011(.dina(w_n1325_0[1]),.dinb(w_n1317_0[1]),.dout(n1326),.clk(gclk));
	jnot g1012(.din(w_n1301_0[0]),.dout(n1327),.clk(gclk));
	jnot g1013(.din(w_n1309_0[0]),.dout(n1328),.clk(gclk));
	jand g1014(.dina(n1328),.dinb(n1327),.dout(n1329),.clk(gclk));
	jnot g1015(.din(w_n1317_0[0]),.dout(n1330),.clk(gclk));
	jnot g1016(.din(w_n1325_0[0]),.dout(n1331),.clk(gclk));
	jand g1017(.dina(n1331),.dinb(n1330),.dout(n1332),.clk(gclk));
	jor g1018(.dina(n1332),.dinb(n1329),.dout(n1333),.clk(gclk));
	jor g1019(.dina(n1333),.dinb(n1326),.dout(n1334),.clk(gclk));
	jor g1020(.dina(n1334),.dinb(n1311),.dout(n1335),.clk(gclk));
	jxor g1021(.dina(w_n744_0[0]),.dinb(w_n730_0[0]),.dout(n1336),.clk(gclk));
	jxor g1022(.dina(n1336),.dinb(w_n737_0[0]),.dout(n1337),.clk(gclk));
	jxor g1023(.dina(w_n754_0[0]),.dinb(w_n723_0[0]),.dout(n1338),.clk(gclk));
	jnot g1024(.din(w_n994_0[0]),.dout(n1339),.clk(gclk));
	jand g1025(.dina(w_n1016_0[0]),.dinb(n1339),.dout(n1340),.clk(gclk));
	jnot g1026(.din(w_n1015_0[0]),.dout(n1341),.clk(gclk));
	jand g1027(.dina(n1341),.dinb(w_n995_0[0]),.dout(n1342),.clk(gclk));
	jor g1028(.dina(n1342),.dinb(n1340),.dout(n1343),.clk(gclk));
	jnot g1029(.din(w_n987_0[0]),.dout(n1344),.clk(gclk));
	jand g1030(.dina(w_n1009_0[1]),.dinb(n1344),.dout(n1345),.clk(gclk));
	jnot g1031(.din(w_n1008_0[0]),.dout(n1346),.clk(gclk));
	jand g1032(.dina(n1346),.dinb(w_n988_0[0]),.dout(n1347),.clk(gclk));
	jor g1033(.dina(n1347),.dinb(n1345),.dout(n1348),.clk(gclk));
	jxor g1034(.dina(n1348),.dinb(n1343),.dout(n1349),.clk(gclk));
	jnot g1035(.din(G181),.dout(n1350),.clk(gclk));
	jor g1036(.dina(n1350),.dinb(w_n355_8[2]),.dout(n1351),.clk(gclk));
	jand g1037(.dina(n1351),.dinb(w_n1166_0[0]),.dout(n1352),.clk(gclk));
	jxor g1038(.dina(n1352),.dinb(n1349),.dout(n1353),.clk(gclk));
	jxor g1039(.dina(n1353),.dinb(n1338),.dout(n1354),.clk(gclk));
	jxor g1040(.dina(n1354),.dinb(n1337),.dout(n1355),.clk(gclk));
	jor g1041(.dina(n1355),.dinb(n1335),.dout(G416_fa_),.clk(gclk));
	jnot g1042(.din(w_n372_1[0]),.dout(n1357),.clk(gclk));
	jxor g1043(.dina(w_n377_0[1]),.dinb(w_G3717_1[0]),.dout(n1358),.clk(gclk));
	jand g1044(.dina(n1358),.dinb(n1357),.dout(n1359),.clk(gclk));
	jnot g1045(.din(w_n387_0[1]),.dout(n1360),.clk(gclk));
	jxor g1046(.dina(w_n401_0[2]),.dinb(w_G3705_1[1]),.dout(n1361),.clk(gclk));
	jand g1047(.dina(w_n1361_0[1]),.dinb(w_n362_0[1]),.dout(n1362),.clk(gclk));
	jand g1048(.dina(w_n1362_0[1]),.dinb(w_G4526_0[2]),.dout(n1363),.clk(gclk));
	jand g1049(.dina(n1363),.dinb(w_n1360_1[1]),.dout(n1364),.clk(gclk));
	jand g1050(.dina(n1364),.dinb(w_n1359_0[2]),.dout(n1365),.clk(gclk));
	jnot g1051(.din(w_n407_0[1]),.dout(n1366),.clk(gclk));
	jand g1052(.dina(w_n1361_0[0]),.dinb(w_n390_1[0]),.dout(n1367),.clk(gclk));
	jand g1053(.dina(n1367),.dinb(w_n1360_1[0]),.dout(n1368),.clk(gclk));
	jor g1054(.dina(n1368),.dinb(n1366),.dout(n1369),.clk(gclk));
	jand g1055(.dina(n1369),.dinb(w_n1359_0[1]),.dout(n1370),.clk(gclk));
	jnot g1056(.din(w_n413_0[2]),.dout(n1371),.clk(gclk));
	jand g1057(.dina(n1371),.dinb(w_n1359_0[0]),.dout(n1372),.clk(gclk));
	jnot g1058(.din(w_n419_0[0]),.dout(n1373),.clk(gclk));
	jor g1059(.dina(n1373),.dinb(n1372),.dout(n1374),.clk(gclk));
	jor g1060(.dina(n1374),.dinb(n1370),.dout(n1375),.clk(gclk));
	jor g1061(.dina(n1375),.dinb(n1365),.dout(n1376),.clk(gclk));
	jnot g1062(.din(w_n452_0[0]),.dout(n1377),.clk(gclk));
	jand g1063(.dina(n1377),.dinb(w_n1376_0[1]),.dout(n1378),.clk(gclk));
	jnot g1064(.din(w_n464_0[0]),.dout(n1379),.clk(gclk));
	jor g1065(.dina(n1379),.dinb(n1378),.dout(n1380),.clk(gclk));
	jand g1066(.dina(w_n494_0[0]),.dinb(w_n1380_1[1]),.dout(n1381),.clk(gclk));
	jnot g1067(.din(w_n518_0[0]),.dout(n1382),.clk(gclk));
	jor g1068(.dina(n1382),.dinb(n1381),.dout(n1383),.clk(gclk));
	jand g1069(.dina(w_n542_0[0]),.dinb(w_n1383_1[2]),.dout(n1384),.clk(gclk));
	jor g1070(.dina(w_n560_0[0]),.dinb(n1384),.dout(n1385),.clk(gclk));
	jxor g1071(.dina(w_n578_1[0]),.dinb(w_n1385_1[1]),.dout(w_dff_A_7i4JzMTm0_2),.clk(gclk));
	jand g1072(.dina(w_n592_0[0]),.dinb(w_n1385_1[0]),.dout(n1387),.clk(gclk));
	jnot g1073(.din(w_n617_0[0]),.dout(n1388),.clk(gclk));
	jor g1074(.dina(n1388),.dinb(n1387),.dout(n1389),.clk(gclk));
	jand g1075(.dina(w_n637_0[0]),.dinb(w_n1389_1[1]),.dout(n1390),.clk(gclk));
	jnot g1076(.din(w_n656_0[0]),.dout(n1391),.clk(gclk));
	jor g1077(.dina(n1391),.dinb(n1390),.dout(n1392),.clk(gclk));
	jxor g1078(.dina(w_n678_0[1]),.dinb(w_n1392_1[1]),.dout(w_dff_A_DICIafTn4_2),.clk(gclk));
	jor g1079(.dina(w_n1033_0[0]),.dinb(w_n957_0[0]),.dout(n1394),.clk(gclk));
	jand g1080(.dina(n1394),.dinb(w_n905_0[0]),.dout(n1395),.clk(gclk));
	jor g1081(.dina(n1395),.dinb(w_n1044_0[0]),.dout(n1396),.clk(gclk));
	jand g1082(.dina(n1396),.dinb(w_n864_0[0]),.dout(n1397),.clk(gclk));
	jor g1083(.dina(n1397),.dinb(w_n981_0[0]),.dout(n1398),.clk(gclk));
	jand g1084(.dina(n1398),.dinb(w_n810_0[0]),.dout(n1399),.clk(gclk));
	jor g1085(.dina(n1399),.dinb(w_n972_0[0]),.dout(w_dff_A_NQVt2kRm1_2),.clk(gclk));
	jnot g1086(.din(w_n568_0[1]),.dout(n1401),.clk(gclk));
	jnot g1087(.din(w_n584_0[1]),.dout(n1402),.clk(gclk));
	jnot g1088(.din(w_n589_1[0]),.dout(n1403),.clk(gclk));
	jnot g1089(.din(w_n579_0[1]),.dout(n1404),.clk(gclk));
	jor g1090(.dina(w_n1404_0[1]),.dinb(w_n562_0[1]),.dout(n1405),.clk(gclk));
	jor g1091(.dina(w_n1405_0[1]),.dinb(w_n1403_0[1]),.dout(n1406),.clk(gclk));
	jor g1092(.dina(w_n1406_0[1]),.dinb(w_n1402_0[1]),.dout(n1407),.clk(gclk));
	jand g1093(.dina(n1407),.dinb(w_n615_1[0]),.dout(n1408),.clk(gclk));
	jxor g1094(.dina(n1408),.dinb(w_n1401_0[1]),.dout(w_dff_A_lRTJsLNs9_2),.clk(gclk));
	jand g1095(.dina(w_n1406_0[0]),.dinb(w_n613_0[1]),.dout(n1410),.clk(gclk));
	jxor g1096(.dina(n1410),.dinb(w_n1402_0[0]),.dout(w_dff_A_lnjGnJCt2_2),.clk(gclk));
	jnot g1097(.din(w_n608_0[1]),.dout(n1412),.clk(gclk));
	jnot g1098(.din(w_n607_0[0]),.dout(n1413),.clk(gclk));
	jand g1099(.dina(n1413),.dinb(n1412),.dout(n1414),.clk(gclk));
	jand g1100(.dina(w_n1414_0[1]),.dinb(w_n1405_0[0]),.dout(n1415),.clk(gclk));
	jxor g1101(.dina(n1415),.dinb(w_n1403_0[0]),.dout(w_dff_A_8uxDTvgW9_2),.clk(gclk));
	jand g1102(.dina(w_n578_0[2]),.dinb(w_n1385_0[2]),.dout(n1417),.clk(gclk));
	jor g1103(.dina(n1417),.dinb(w_n606_1[1]),.dout(n1418),.clk(gclk));
	jxor g1104(.dina(n1418),.dinb(w_n573_0[2]),.dout(w_dff_A_msuIofH91_2),.clk(gclk));
	jnot g1105(.din(w_n661_0[0]),.dout(n1420),.clk(gclk));
	jnot g1106(.din(w_n665_0[1]),.dout(n1421),.clk(gclk));
	jnot g1107(.din(w_n669_0[1]),.dout(n1422),.clk(gclk));
	jnot g1108(.din(w_n679_1[0]),.dout(n1423),.clk(gclk));
	jor g1109(.dina(n1423),.dinb(w_n657_1[0]),.dout(n1424),.clk(gclk));
	jor g1110(.dina(w_n1424_0[1]),.dinb(w_n1422_0[1]),.dout(n1425),.clk(gclk));
	jor g1111(.dina(w_n1425_0[1]),.dinb(w_n1421_0[1]),.dout(n1426),.clk(gclk));
	jand g1112(.dina(n1426),.dinb(w_n704_0[0]),.dout(n1427),.clk(gclk));
	jxor g1113(.dina(n1427),.dinb(w_n1420_0[2]),.dout(w_dff_A_6shXyOtb9_2),.clk(gclk));
	jnot g1114(.din(w_n701_1[0]),.dout(n1429),.clk(gclk));
	jand g1115(.dina(w_n1425_0[0]),.dinb(n1429),.dout(n1430),.clk(gclk));
	jxor g1116(.dina(n1430),.dinb(w_n1421_0[0]),.dout(w_dff_A_YJxM6Mt30_2),.clk(gclk));
	jnot g1117(.din(w_n699_1[0]),.dout(n1432),.clk(gclk));
	jand g1118(.dina(w_n1424_0[0]),.dinb(n1432),.dout(n1433),.clk(gclk));
	jxor g1119(.dina(n1433),.dinb(w_n1422_0[0]),.dout(w_dff_A_VslLU2ex9_2),.clk(gclk));
	jand g1120(.dina(w_n678_0[0]),.dinb(w_n1392_1[0]),.dout(n1435),.clk(gclk));
	jor g1121(.dina(n1435),.dinb(w_n697_0[1]),.dout(n1436),.clk(gclk));
	jxor g1122(.dina(n1436),.dinb(w_n674_1[0]),.dout(w_dff_A_EI1P8NHh9_2),.clk(gclk));
	jor g1123(.dina(w_G408_0),.dinb(w_G404_0),.dout(n1438),.clk(gclk));
	jor g1124(.dina(w_G410_0),.dinb(w_G406_0),.dout(n1439),.clk(gclk));
	jor g1125(.dina(n1439),.dinb(n1438),.dout(n1440),.clk(gclk));
	jor g1126(.dina(w_dff_B_7o9MhInf4_0),.dinb(w_G412_0),.dout(n1441),.clk(gclk));
	jor g1127(.dina(w_dff_B_GEaJHj6j2_0),.dinb(w_G416_0),.dout(n1442),.clk(gclk));
	jor g1128(.dina(n1442),.dinb(w_G414_0),.dout(w_dff_A_zFFMkuIJ3_2),.clk(gclk));
	jnot g1129(.din(w_n631_0[0]),.dout(n1444),.clk(gclk));
	jnot g1130(.din(w_n627_0[0]),.dout(n1445),.clk(gclk));
	jor g1131(.dina(w_n1445_0[1]),.dinb(w_n618_0[1]),.dout(n1446),.clk(gclk));
	jand g1132(.dina(n1446),.dinb(w_n648_0[1]),.dout(n1447),.clk(gclk));
	jor g1133(.dina(w_n1447_0[1]),.dinb(w_n653_1[0]),.dout(n1448),.clk(gclk));
	jand g1134(.dina(n1448),.dinb(w_n643_0[0]),.dout(n1449),.clk(gclk));
	jxor g1135(.dina(n1449),.dinb(w_n1444_0[2]),.dout(w_dff_A_OflSHxKU6_2),.clk(gclk));
	jnot g1136(.din(w_n635_0[1]),.dout(n1451),.clk(gclk));
	jxor g1137(.dina(w_n1447_0[0]),.dinb(w_dff_B_fbaVvFO18_1),.dout(w_dff_A_dsbSATGu4_2),.clk(gclk));
	jand g1138(.dina(w_n1156_0[0]),.dinb(w_G2239_0[1]),.dout(n1453),.clk(gclk));
	jnot g1139(.din(n1453),.dout(n1454),.clk(gclk));
	jand g1140(.dina(w_n1454_0[1]),.dinb(w_n1389_1[0]),.dout(n1455),.clk(gclk));
	jor g1141(.dina(n1455),.dinb(w_n645_0[1]),.dout(n1456),.clk(gclk));
	jxor g1142(.dina(n1456),.dinb(w_n622_0[2]),.dout(w_dff_A_5LuU9lJA3_2),.clk(gclk));
	jxor g1143(.dina(w_n626_0[0]),.dinb(w_n1389_0[2]),.dout(w_dff_A_tQ3YGlOH2_2),.clk(gclk));
	jxor g1144(.dina(w_n480_1[0]),.dinb(w_n1380_1[0]),.dout(w_dff_A_sgRaRusK5_2),.clk(gclk));
	jnot g1145(.din(w_n714_0[0]),.dout(n1460),.clk(gclk));
	jnot g1146(.din(w_n365_0[0]),.dout(n1461),.clk(gclk));
	jor g1147(.dina(w_n711_0[0]),.dinb(w_n710_0[0]),.dout(n1462),.clk(gclk));
	jxor g1148(.dina(n1462),.dinb(n1461),.dout(n1463),.clk(gclk));
	jnot g1149(.din(w_n1463_0[2]),.dout(n1464),.clk(gclk));
	jor g1150(.dina(w_n1464_0[1]),.dinb(n1460),.dout(n1465),.clk(gclk));
	jand g1151(.dina(w_n1465_0[1]),.dinb(w_n715_0[1]),.dout(w_dff_A_0s1VMX2B6_2),.clk(gclk));
	jxor g1152(.dina(w_n713_1[0]),.dinb(w_n709_1[0]),.dout(w_dff_A_PDuO5PBw0_2),.clk(gclk));
	jnot g1153(.din(w_n470_0[1]),.dout(n1468),.clk(gclk));
	jnot g1154(.din(w_n486_0[1]),.dout(n1469),.clk(gclk));
	jnot g1155(.din(w_n491_1[0]),.dout(n1470),.clk(gclk));
	jnot g1156(.din(w_n481_0[1]),.dout(n1471),.clk(gclk));
	jor g1157(.dina(w_n1471_0[1]),.dinb(w_n465_0[1]),.dout(n1472),.clk(gclk));
	jor g1158(.dina(w_n1472_0[1]),.dinb(w_n1470_0[1]),.dout(n1473),.clk(gclk));
	jor g1159(.dina(w_n1473_0[1]),.dinb(w_n1469_0[1]),.dout(n1474),.clk(gclk));
	jand g1160(.dina(n1474),.dinb(w_n516_0[1]),.dout(n1475),.clk(gclk));
	jxor g1161(.dina(n1475),.dinb(w_n1468_0[1]),.dout(w_dff_A_VtwlBwvj4_2),.clk(gclk));
	jand g1162(.dina(w_n1473_0[0]),.dinb(w_n514_0[1]),.dout(n1477),.clk(gclk));
	jxor g1163(.dina(n1477),.dinb(w_n1469_0[0]),.dout(w_dff_A_cH5sdleA0_2),.clk(gclk));
	jand g1164(.dina(w_n508_0[0]),.dinb(w_n510_0[0]),.dout(n1479),.clk(gclk));
	jand g1165(.dina(w_n1479_0[1]),.dinb(w_n1472_0[0]),.dout(n1480),.clk(gclk));
	jxor g1166(.dina(n1480),.dinb(w_n1470_0[0]),.dout(w_dff_A_lHS6djP02_2),.clk(gclk));
	jnot g1167(.din(w_n507_1[1]),.dout(n1482),.clk(gclk));
	jand g1168(.dina(w_n480_0[2]),.dinb(w_n1380_0[2]),.dout(n1483),.clk(gclk));
	jor g1169(.dina(n1483),.dinb(w_n1482_0[1]),.dout(n1484),.clk(gclk));
	jxor g1170(.dina(n1484),.dinb(w_n475_0[2]),.dout(w_dff_A_2DLI61aZ0_2),.clk(gclk));
	jand g1171(.dina(w_n530_0[0]),.dinb(w_n1383_1[1]),.dout(n1486),.clk(gclk));
	jand g1172(.dina(w_n1486_0[1]),.dinb(w_n552_0[0]),.dout(n1487),.clk(gclk));
	jor g1173(.dina(n1487),.dinb(w_n558_0[1]),.dout(n1488),.clk(gclk));
	jxor g1174(.dina(n1488),.dinb(w_n535_1[0]),.dout(w_dff_A_1HLKbfCP9_2),.clk(gclk));
	jor g1175(.dina(w_n1486_0[0]),.dinb(w_n556_0[1]),.dout(n1490),.clk(gclk));
	jxor g1176(.dina(n1490),.dinb(w_n540_0[1]),.dout(w_dff_A_aUo2VDAg5_2),.clk(gclk));
	jnot g1177(.din(w_n528_0[1]),.dout(n1492),.clk(gclk));
	jand g1178(.dina(n1492),.dinb(w_G4420_0[1]),.dout(n1493),.clk(gclk));
	jnot g1179(.din(n1493),.dout(n1494),.clk(gclk));
	jand g1180(.dina(w_n1494_0[2]),.dinb(w_n1383_1[0]),.dout(n1495),.clk(gclk));
	jor g1181(.dina(n1495),.dinb(w_n554_0[1]),.dout(n1496),.clk(gclk));
	jxor g1182(.dina(n1496),.dinb(w_n524_1[2]),.dout(w_dff_A_19A0fWNC1_2),.clk(gclk));
	jxor g1183(.dina(w_n529_0[0]),.dinb(w_n1383_0[2]),.dout(w_dff_A_aevorycp8_2),.clk(gclk));
	jxor g1184(.dina(w_n589_0[2]),.dinb(w_n584_0[0]),.dout(n1499),.clk(gclk));
	jxor g1185(.dina(n1499),.dinb(w_n635_0[0]),.dout(n1500),.clk(gclk));
	jnot g1186(.din(w_n622_0[1]),.dout(n1501),.clk(gclk));
	jnot g1187(.din(w_n653_0[2]),.dout(n1502),.clk(gclk));
	jand g1188(.dina(w_n647_0[0]),.dinb(n1502),.dout(n1503),.clk(gclk));
	jor g1189(.dina(n1503),.dinb(w_n649_0[0]),.dout(n1504),.clk(gclk));
	jxor g1190(.dina(n1504),.dinb(w_n1444_0[1]),.dout(n1505),.clk(gclk));
	jxor g1191(.dina(n1505),.dinb(w_n1501_0[1]),.dout(n1506),.clk(gclk));
	jxor g1192(.dina(n1506),.dinb(w_n1454_0[0]),.dout(n1507),.clk(gclk));
	jand g1193(.dina(n1507),.dinb(w_n618_0[0]),.dout(n1508),.clk(gclk));
	jxor g1194(.dina(w_n645_0[0]),.dinb(w_n1501_0[0]),.dout(n1509),.clk(gclk));
	jand g1195(.dina(w_n648_0[0]),.dinb(w_n1445_0[0]),.dout(n1510),.clk(gclk));
	jnot g1196(.din(w_n1510_0[1]),.dout(n1511),.clk(gclk));
	jor g1197(.dina(n1511),.dinb(w_n642_0[0]),.dout(n1512),.clk(gclk));
	jor g1198(.dina(w_n1510_0[0]),.dinb(w_n653_0[1]),.dout(n1513),.clk(gclk));
	jand g1199(.dina(n1513),.dinb(n1512),.dout(n1514),.clk(gclk));
	jxor g1200(.dina(n1514),.dinb(w_n1444_0[0]),.dout(n1515),.clk(gclk));
	jxor g1201(.dina(n1515),.dinb(n1509),.dout(n1516),.clk(gclk));
	jand g1202(.dina(n1516),.dinb(w_n1389_0[1]),.dout(n1517),.clk(gclk));
	jor g1203(.dina(n1517),.dinb(n1508),.dout(n1518),.clk(gclk));
	jand g1204(.dina(w_n613_0[0]),.dinb(w_n606_1[0]),.dout(n1519),.clk(gclk));
	jnot g1205(.din(w_n606_0[2]),.dout(n1520),.clk(gclk));
	jand g1206(.dina(w_n605_0[0]),.dinb(w_n1520_0[1]),.dout(n1521),.clk(gclk));
	jand g1207(.dina(n1521),.dinb(w_n610_0[0]),.dout(n1522),.clk(gclk));
	jxor g1208(.dina(n1522),.dinb(w_n578_0[1]),.dout(n1523),.clk(gclk));
	jor g1209(.dina(n1523),.dinb(n1519),.dout(n1524),.clk(gclk));
	jor g1210(.dina(w_n572_0[1]),.dinb(w_n569_0[0]),.dout(n1525),.clk(gclk));
	jand g1211(.dina(w_n1520_0[0]),.dinb(n1525),.dout(n1526),.clk(gclk));
	jor g1212(.dina(n1526),.dinb(w_n608_0[0]),.dout(n1527),.clk(gclk));
	jxor g1213(.dina(n1527),.dinb(w_n615_0[2]),.dout(n1528),.clk(gclk));
	jxor g1214(.dina(n1528),.dinb(w_n1401_0[0]),.dout(n1529),.clk(gclk));
	jxor g1215(.dina(n1529),.dinb(n1524),.dout(n1530),.clk(gclk));
	jor g1216(.dina(n1530),.dinb(w_n1385_0[1]),.dout(n1531),.clk(gclk));
	jand g1217(.dina(w_n1414_0[0]),.dinb(w_n1404_0[0]),.dout(n1532),.clk(gclk));
	jxor g1218(.dina(n1532),.dinb(w_n568_0[0]),.dout(n1533),.clk(gclk));
	jxor g1219(.dina(w_n606_0[1]),.dinb(w_n573_0[1]),.dout(n1534),.clk(gclk));
	jand g1220(.dina(w_n589_0[1]),.dinb(w_n579_0[0]),.dout(n1535),.clk(gclk));
	jor g1221(.dina(n1535),.dinb(w_n612_0[0]),.dout(n1536),.clk(gclk));
	jnot g1222(.din(w_n1536_0[1]),.dout(n1537),.clk(gclk));
	jand g1223(.dina(n1537),.dinb(w_n599_0[0]),.dout(n1538),.clk(gclk));
	jnot g1224(.din(w_n591_0[0]),.dout(n1539),.clk(gclk));
	jand g1225(.dina(w_n1536_0[0]),.dinb(n1539),.dout(n1540),.clk(gclk));
	jand g1226(.dina(n1540),.dinb(w_n615_0[1]),.dout(n1541),.clk(gclk));
	jor g1227(.dina(n1541),.dinb(n1538),.dout(n1542),.clk(gclk));
	jxor g1228(.dina(n1542),.dinb(n1534),.dout(n1543),.clk(gclk));
	jxor g1229(.dina(n1543),.dinb(n1533),.dout(n1544),.clk(gclk));
	jor g1230(.dina(n1544),.dinb(w_n562_0[0]),.dout(n1545),.clk(gclk));
	jand g1231(.dina(n1545),.dinb(n1531),.dout(n1546),.clk(gclk));
	jxor g1232(.dina(n1546),.dinb(n1518),.dout(n1547),.clk(gclk));
	jxor g1233(.dina(n1547),.dinb(w_dff_B_ZBSCXzLP5_1),.dout(w_dff_A_AskpEjKv5_2),.clk(gclk));
	jand g1234(.dina(w_n713_0[2]),.dinb(w_n709_0[2]),.dout(n1549),.clk(gclk));
	jor g1235(.dina(n1549),.dinb(w_n1463_0[1]),.dout(n1550),.clk(gclk));
	jnot g1236(.din(w_n683_0[0]),.dout(n1551),.clk(gclk));
	jand g1237(.dina(w_n707_0[1]),.dinb(w_n1392_0[2]),.dout(n1552),.clk(gclk));
	jand g1238(.dina(w_n712_0[0]),.dinb(w_n708_0[0]),.dout(n1553),.clk(gclk));
	jor g1239(.dina(n1553),.dinb(w_n1464_0[0]),.dout(n1554),.clk(gclk));
	jor g1240(.dina(n1554),.dinb(n1552),.dout(n1555),.clk(gclk));
	jor g1241(.dina(n1555),.dinb(n1551),.dout(n1556),.clk(gclk));
	jand g1242(.dina(n1556),.dinb(n1550),.dout(n1557),.clk(gclk));
	jand g1243(.dina(w_n1463_0[0]),.dinb(w_n707_0[0]),.dout(n1558),.clk(gclk));
	jand g1244(.dina(n1558),.dinb(w_n657_0[2]),.dout(n1559),.clk(gclk));
	jor g1245(.dina(n1559),.dinb(n1557),.dout(n1560),.clk(gclk));
	jxor g1246(.dina(w_n669_0[0]),.dinb(w_n665_0[0]),.dout(n1561),.clk(gclk));
	jor g1247(.dina(w_n701_0[2]),.dinb(w_n686_0[0]),.dout(n1562),.clk(gclk));
	jand g1248(.dina(n1562),.dinb(w_n703_0[0]),.dout(n1563),.clk(gclk));
	jxor g1249(.dina(n1563),.dinb(w_n1420_0[1]),.dout(n1564),.clk(gclk));
	jor g1250(.dina(w_n677_0[0]),.dinb(w_n675_0[0]),.dout(n1565),.clk(gclk));
	jxor g1251(.dina(n1565),.dinb(w_n674_0[2]),.dout(n1566),.clk(gclk));
	jxor g1252(.dina(n1566),.dinb(w_n699_0[2]),.dout(n1567),.clk(gclk));
	jxor g1253(.dina(n1567),.dinb(n1564),.dout(n1568),.clk(gclk));
	jand g1254(.dina(n1568),.dinb(w_n657_0[1]),.dout(n1569),.clk(gclk));
	jand g1255(.dina(w_n679_0[2]),.dinb(w_n692_0[0]),.dout(n1570),.clk(gclk));
	jor g1256(.dina(n1570),.dinb(w_n701_0[1]),.dout(n1571),.clk(gclk));
	jor g1257(.dina(w_n1571_0[1]),.dinb(w_n687_0[0]),.dout(n1572),.clk(gclk));
	jnot g1258(.din(w_n1571_0[0]),.dout(n1573),.clk(gclk));
	jor g1259(.dina(n1573),.dinb(w_n680_0[0]),.dout(n1574),.clk(gclk));
	jor g1260(.dina(n1574),.dinb(w_n705_0[0]),.dout(n1575),.clk(gclk));
	jand g1261(.dina(n1575),.dinb(n1572),.dout(n1576),.clk(gclk));
	jor g1262(.dina(w_n699_0[1]),.dinb(w_n679_0[1]),.dout(n1577),.clk(gclk));
	jxor g1263(.dina(n1577),.dinb(w_n1420_0[0]),.dout(n1578),.clk(gclk));
	jxor g1264(.dina(n1578),.dinb(n1576),.dout(n1579),.clk(gclk));
	jxor g1265(.dina(n1579),.dinb(w_n697_0[0]),.dout(n1580),.clk(gclk));
	jxor g1266(.dina(n1580),.dinb(w_n674_0[1]),.dout(n1581),.clk(gclk));
	jand g1267(.dina(n1581),.dinb(w_n1392_0[1]),.dout(n1582),.clk(gclk));
	jor g1268(.dina(n1582),.dinb(n1569),.dout(n1583),.clk(gclk));
	jxor g1269(.dina(n1583),.dinb(n1561),.dout(n1584),.clk(gclk));
	jxor g1270(.dina(w_dff_B_mRB84Aq46_0),.dinb(n1560),.dout(G338),.clk(gclk));
	jxor g1271(.dina(w_n491_0[2]),.dinb(w_n486_0[0]),.dout(n1586),.clk(gclk));
	jxor g1272(.dina(n1586),.dinb(w_n540_0[0]),.dout(n1587),.clk(gclk));
	jnot g1273(.din(w_n535_0[2]),.dout(n1588),.clk(gclk));
	jnot g1274(.din(w_n557_0[0]),.dout(n1589),.clk(gclk));
	jor g1275(.dina(w_n556_0[0]),.dinb(w_n549_0[0]),.dout(n1590),.clk(gclk));
	jand g1276(.dina(n1590),.dinb(n1589),.dout(n1591),.clk(gclk));
	jxor g1277(.dina(n1591),.dinb(n1588),.dout(n1592),.clk(gclk));
	jxor g1278(.dina(w_n1494_0[1]),.dinb(w_n524_1[1]),.dout(n1593),.clk(gclk));
	jxor g1279(.dina(n1593),.dinb(n1592),.dout(n1594),.clk(gclk));
	jand g1280(.dina(n1594),.dinb(w_n519_0[0]),.dout(n1595),.clk(gclk));
	jxor g1281(.dina(w_n554_0[0]),.dinb(w_n524_1[0]),.dout(n1596),.clk(gclk));
	jxor g1282(.dina(n1596),.dinb(w_n535_0[1]),.dout(n1597),.clk(gclk));
	jand g1283(.dina(w_n1494_0[0]),.dinb(w_n524_0[2]),.dout(n1598),.clk(gclk));
	jor g1284(.dina(n1598),.dinb(w_n553_0[0]),.dout(n1599),.clk(gclk));
	jnot g1285(.din(w_n1599_0[1]),.dout(n1600),.clk(gclk));
	jand g1286(.dina(n1600),.dinb(w_n558_0[0]),.dout(n1601),.clk(gclk));
	jand g1287(.dina(w_n1599_0[0]),.dinb(w_n551_0[0]),.dout(n1602),.clk(gclk));
	jor g1288(.dina(n1602),.dinb(n1601),.dout(n1603),.clk(gclk));
	jxor g1289(.dina(n1603),.dinb(n1597),.dout(n1604),.clk(gclk));
	jand g1290(.dina(n1604),.dinb(w_n1383_0[1]),.dout(n1605),.clk(gclk));
	jor g1291(.dina(n1605),.dinb(n1595),.dout(n1606),.clk(gclk));
	jor g1292(.dina(w_n474_0[1]),.dinb(w_n471_0[0]),.dout(n1607),.clk(gclk));
	jand g1293(.dina(w_n507_1[0]),.dinb(n1607),.dout(n1608),.clk(gclk));
	jor g1294(.dina(n1608),.dinb(w_n509_0[0]),.dout(n1609),.clk(gclk));
	jnot g1295(.din(w_n516_0[0]),.dout(n1610),.clk(gclk));
	jnot g1296(.din(w_n514_0[0]),.dout(n1611),.clk(gclk));
	jor g1297(.dina(w_n1611_0[1]),.dinb(w_n507_0[2]),.dout(n1612),.clk(gclk));
	jor g1298(.dina(w_n505_0[0]),.dinb(w_n1482_0[0]),.dout(n1613),.clk(gclk));
	jor g1299(.dina(n1613),.dinb(w_n512_0[0]),.dout(n1614),.clk(gclk));
	jxor g1300(.dina(n1614),.dinb(w_n480_0[1]),.dout(n1615),.clk(gclk));
	jand g1301(.dina(n1615),.dinb(n1612),.dout(n1616),.clk(gclk));
	jxor g1302(.dina(n1616),.dinb(w_n1468_0[0]),.dout(n1617),.clk(gclk));
	jxor g1303(.dina(n1617),.dinb(w_n1610_0[1]),.dout(n1618),.clk(gclk));
	jxor g1304(.dina(n1618),.dinb(n1609),.dout(n1619),.clk(gclk));
	jor g1305(.dina(n1619),.dinb(w_n1380_0[1]),.dout(n1620),.clk(gclk));
	jand g1306(.dina(w_n1479_0[0]),.dinb(w_n1471_0[0]),.dout(n1621),.clk(gclk));
	jxor g1307(.dina(n1621),.dinb(w_n470_0[0]),.dout(n1622),.clk(gclk));
	jxor g1308(.dina(w_n507_0[1]),.dinb(w_n475_0[1]),.dout(n1623),.clk(gclk));
	jand g1309(.dina(w_n491_0[1]),.dinb(w_n481_0[0]),.dout(n1624),.clk(gclk));
	jor g1310(.dina(n1624),.dinb(w_n1611_0[0]),.dout(n1625),.clk(gclk));
	jor g1311(.dina(w_n1625_0[1]),.dinb(w_n502_0[0]),.dout(n1626),.clk(gclk));
	jnot g1312(.din(w_n1625_0[0]),.dout(n1627),.clk(gclk));
	jor g1313(.dina(n1627),.dinb(w_n493_0[0]),.dout(n1628),.clk(gclk));
	jor g1314(.dina(n1628),.dinb(w_n1610_0[0]),.dout(n1629),.clk(gclk));
	jand g1315(.dina(n1629),.dinb(n1626),.dout(n1630),.clk(gclk));
	jxor g1316(.dina(n1630),.dinb(n1623),.dout(n1631),.clk(gclk));
	jxor g1317(.dina(n1631),.dinb(n1622),.dout(n1632),.clk(gclk));
	jor g1318(.dina(n1632),.dinb(w_n465_0[0]),.dout(n1633),.clk(gclk));
	jand g1319(.dina(n1633),.dinb(n1620),.dout(n1634),.clk(gclk));
	jxor g1320(.dina(n1634),.dinb(n1606),.dout(n1635),.clk(gclk));
	jxor g1321(.dina(n1635),.dinb(w_dff_B_ixTSlmXd3_1),.dout(w_dff_A_Gw55g2Xc2_2),.clk(gclk));
	jxor g1322(.dina(w_n450_0[0]),.dinb(w_n1360_0[2]),.dout(n1637),.clk(gclk));
	jnot g1323(.din(w_n455_0[0]),.dout(n1638),.clk(gclk));
	jnot g1324(.din(w_n460_0[0]),.dout(n1639),.clk(gclk));
	jor g1325(.dina(n1639),.dinb(n1638),.dout(n1640),.clk(gclk));
	jand g1326(.dina(n1640),.dinb(w_n461_0[0]),.dout(n1641),.clk(gclk));
	jxor g1327(.dina(n1641),.dinb(w_n446_0[2]),.dout(n1642),.clk(gclk));
	jnot g1328(.din(w_n1642_0[1]),.dout(n1643),.clk(gclk));
	jxor g1329(.dina(w_n1148_0[1]),.dinb(w_n429_1[1]),.dout(n1644),.clk(gclk));
	jnot g1330(.din(w_n1644_0[1]),.dout(n1645),.clk(gclk));
	jor g1331(.dina(n1645),.dinb(n1643),.dout(n1646),.clk(gclk));
	jor g1332(.dina(w_n1644_0[0]),.dinb(w_n1642_0[0]),.dout(n1647),.clk(gclk));
	jand g1333(.dina(n1647),.dinb(w_n422_0[1]),.dout(n1648),.clk(gclk));
	jand g1334(.dina(n1648),.dinb(n1646),.dout(n1649),.clk(gclk));
	jxor g1335(.dina(w_n458_0[0]),.dinb(w_n429_1[0]),.dout(n1650),.clk(gclk));
	jxor g1336(.dina(n1650),.dinb(w_n446_0[1]),.dout(n1651),.clk(gclk));
	jnot g1337(.din(w_n462_0[0]),.dout(n1652),.clk(gclk));
	jor g1338(.dina(w_n1148_0[0]),.dinb(w_n429_0[2]),.dout(n1653),.clk(gclk));
	jand g1339(.dina(n1653),.dinb(w_n457_0[0]),.dout(n1654),.clk(gclk));
	jand g1340(.dina(w_n1654_0[1]),.dinb(n1652),.dout(n1655),.clk(gclk));
	jnot g1341(.din(n1655),.dout(n1656),.clk(gclk));
	jnot g1342(.din(w_n456_0[0]),.dout(n1657),.clk(gclk));
	jor g1343(.dina(w_n1654_0[0]),.dinb(n1657),.dout(n1658),.clk(gclk));
	jand g1344(.dina(n1658),.dinb(n1656),.dout(n1659),.clk(gclk));
	jor g1345(.dina(w_n1659_0[1]),.dinb(w_n1651_0[1]),.dout(n1660),.clk(gclk));
	jnot g1346(.din(w_n1651_0[0]),.dout(n1661),.clk(gclk));
	jnot g1347(.din(w_n1659_0[0]),.dout(n1662),.clk(gclk));
	jor g1348(.dina(n1662),.dinb(n1661),.dout(n1663),.clk(gclk));
	jand g1349(.dina(n1663),.dinb(w_n1376_0[0]),.dout(n1664),.clk(gclk));
	jand g1350(.dina(n1664),.dinb(n1660),.dout(n1665),.clk(gclk));
	jor g1351(.dina(n1665),.dinb(n1649),.dout(n1666),.clk(gclk));
	jand g1352(.dina(w_n1136_0[0]),.dinb(w_n403_0[0]),.dout(n1667),.clk(gclk));
	jnot g1353(.din(w_n1667_0[1]),.dout(n1668),.clk(gclk));
	jor g1354(.dina(n1668),.dinb(w_n1128_0[2]),.dout(n1669),.clk(gclk));
	jnot g1355(.din(w_n1128_0[1]),.dout(n1670),.clk(gclk));
	jand g1356(.dina(w_n1362_0[0]),.dinb(w_n1360_0[1]),.dout(n1671),.clk(gclk));
	jor g1357(.dina(n1671),.dinb(w_n1670_0[1]),.dout(n1672),.clk(gclk));
	jor g1358(.dina(w_n1672_0[1]),.dinb(w_n1667_0[0]),.dout(n1673),.clk(gclk));
	jand g1359(.dina(n1673),.dinb(n1669),.dout(n1674),.clk(gclk));
	jxor g1360(.dina(n1674),.dinb(w_n372_0[2]),.dout(n1675),.clk(gclk));
	jnot g1361(.din(w_n1672_0[0]),.dout(n1676),.clk(gclk));
	jor g1362(.dina(n1676),.dinb(w_n1127_0[0]),.dout(n1677),.clk(gclk));
	jand g1363(.dina(n1677),.dinb(w_n417_0[0]),.dout(n1678),.clk(gclk));
	jxor g1364(.dina(n1678),.dinb(w_n402_0[1]),.dout(n1679),.clk(gclk));
	jxor g1365(.dina(n1679),.dinb(w_n354_0[2]),.dout(n1680),.clk(gclk));
	jnot g1366(.din(w_n1680_0[1]),.dout(n1681),.clk(gclk));
	jand g1367(.dina(n1681),.dinb(w_n1675_0[1]),.dout(n1682),.clk(gclk));
	jnot g1368(.din(w_n1675_0[0]),.dout(n1683),.clk(gclk));
	jand g1369(.dina(w_n1680_0[0]),.dinb(n1683),.dout(n1684),.clk(gclk));
	jor g1370(.dina(n1684),.dinb(w_n388_0[0]),.dout(n1685),.clk(gclk));
	jor g1371(.dina(n1685),.dinb(n1682),.dout(n1686),.clk(gclk));
	jxor g1372(.dina(w_n1130_0[0]),.dinb(w_n372_0[1]),.dout(n1687),.clk(gclk));
	jand g1373(.dina(w_n407_0[0]),.dinb(w_n354_0[1]),.dout(n1688),.clk(gclk));
	jand g1374(.dina(n1688),.dinb(w_n413_0[1]),.dout(n1689),.clk(gclk));
	jand g1375(.dina(w_n1689_0[1]),.dinb(w_n395_0[0]),.dout(n1690),.clk(gclk));
	jnot g1376(.din(w_n1689_0[0]),.dout(n1691),.clk(gclk));
	jand g1377(.dina(w_n1670_0[0]),.dinb(w_n390_0[2]),.dout(n1692),.clk(gclk));
	jor g1378(.dina(n1692),.dinb(w_n362_0[0]),.dout(n1693),.clk(gclk));
	jand g1379(.dina(n1693),.dinb(n1691),.dout(n1694),.clk(gclk));
	jor g1380(.dina(n1694),.dinb(n1690),.dout(n1695),.clk(gclk));
	jand g1381(.dina(w_n401_0[1]),.dinb(w_G3705_1[0]),.dout(n1696),.clk(gclk));
	jor g1382(.dina(n1696),.dinb(w_n390_0[1]),.dout(n1697),.clk(gclk));
	jand g1383(.dina(n1697),.dinb(w_n412_0[0]),.dout(n1698),.clk(gclk));
	jxor g1384(.dina(n1698),.dinb(n1695),.dout(n1699),.clk(gclk));
	jnot g1385(.din(w_n1699_0[1]),.dout(n1700),.clk(gclk));
	jand g1386(.dina(n1700),.dinb(w_n1687_0[1]),.dout(n1701),.clk(gclk));
	jnot g1387(.din(w_n1687_0[0]),.dout(n1702),.clk(gclk));
	jand g1388(.dina(w_n1699_0[0]),.dinb(n1702),.dout(n1703),.clk(gclk));
	jor g1389(.dina(n1703),.dinb(w_G4526_0[1]),.dout(n1704),.clk(gclk));
	jor g1390(.dina(n1704),.dinb(n1701),.dout(n1705),.clk(gclk));
	jand g1391(.dina(n1705),.dinb(n1686),.dout(n1706),.clk(gclk));
	jxor g1392(.dina(n1706),.dinb(w_n379_0[1]),.dout(n1707),.clk(gclk));
	jxor g1393(.dina(n1707),.dinb(n1666),.dout(n1708),.clk(gclk));
	jxor g1394(.dina(n1708),.dinb(w_dff_B_XHnAdNvx9_1),.dout(w_dff_A_ECMPFZkm5_2),.clk(gclk));
	jdff g1395(.din(w_G1_1[1]),.dout(w_dff_A_6sApNmgt4_1));
	jdff g1396(.din(w_G1_1[0]),.dout(w_dff_A_oxIB4Cei6_1));
	jdff g1397(.din(w_G1459_0[0]),.dout(w_dff_A_10WK5Ss63_1));
	jdff g1398(.din(w_G1469_0[1]),.dout(w_dff_A_kCaRS6Sy6_1));
	jdff g1399(.din(w_G1480_0[0]),.dout(w_dff_A_tz2EUH5g2_1));
	jdff g1400(.din(w_G1486_0[0]),.dout(w_dff_A_n6GEbAPE9_1));
	jdff g1401(.din(w_G1492_0[1]),.dout(w_dff_A_eZCLFuLa4_1));
	jdff g1402(.din(w_G1496_0[0]),.dout(w_dff_A_7VdHePjq5_1));
	jdff g1403(.din(w_G2208_0[0]),.dout(w_dff_A_l63WIzjM6_1));
	jdff g1404(.din(w_G2218_0[0]),.dout(w_dff_A_38SOXGaA5_1));
	jdff g1405(.din(w_G2224_0[1]),.dout(w_dff_A_SUaMaM1Z9_1));
	jdff g1406(.din(w_G2230_0[1]),.dout(w_dff_A_3ZgZBMkC9_1));
	jdff g1407(.din(w_G2236_0[1]),.dout(w_dff_A_inOpBq5G8_1));
	jdff g1408(.din(w_G2239_0[0]),.dout(w_dff_A_hlARsFhN7_1));
	jdff g1409(.din(w_G2247_0[0]),.dout(w_dff_A_Yw7VDQLa0_1));
	jdff g1410(.din(w_G2253_0[1]),.dout(w_dff_A_iwHRIdkG4_1));
	jdff g1411(.din(w_G2256_0[1]),.dout(w_dff_A_C0nNn7ci4_1));
	jdff g1412(.din(w_G3698_0[0]),.dout(w_dff_A_d6GEvmtG3_1));
	jdff g1413(.din(w_G3701_0[1]),.dout(w_dff_A_0Uka2LbP9_1));
	jdff g1414(.din(w_G3705_0[2]),.dout(w_dff_A_KehafRC34_1));
	jdff g1415(.din(w_G3711_0[1]),.dout(w_dff_A_jDpzQ2aJ2_1));
	jdff g1416(.din(w_G3717_0[2]),.dout(w_dff_A_Y9ZWrAog2_1));
	jdff g1417(.din(w_G3723_0[1]),.dout(w_dff_A_0ix5qubp0_1));
	jdff g1418(.din(w_G3729_0[1]),.dout(w_dff_A_wgAbeICk9_1));
	jdff g1419(.din(w_G3737_0[1]),.dout(w_dff_A_CfDvIimZ4_1));
	jdff g1420(.din(w_G3743_0[1]),.dout(w_dff_A_8brKNuEG7_1));
	jdff g1421(.din(w_G3749_0[1]),.dout(w_dff_A_Sld5T4WZ8_1));
	jdff g1422(.din(w_G4393_0[0]),.dout(w_dff_A_2zsj2RB06_1));
	jdff g1423(.din(w_G4400_0[0]),.dout(w_dff_A_r0bXZQNs5_1));
	jdff g1424(.din(w_G4405_0[1]),.dout(w_dff_A_Z2eAlHCZ6_1));
	jdff g1425(.din(w_G4410_0[1]),.dout(w_dff_A_iSHkyrCa3_1));
	jdff g1426(.din(w_G4415_0[1]),.dout(w_dff_A_sSU8Nc0v8_1));
	jdff g1427(.din(w_G4420_0[0]),.dout(w_dff_A_Of9VtPSQ2_1));
	jdff g1428(.din(w_G4427_0[0]),.dout(w_dff_A_ztpM8bzy9_1));
	jdff g1429(.din(w_G4432_0[1]),.dout(w_dff_A_xlD6j1Zi9_1));
	jdff g1430(.din(w_G4437_0[0]),.dout(w_dff_A_HrHW1qMA5_1));
	jdff g1431(.din(w_G1462_0[0]),.dout(w_dff_A_hGOFpqrP7_1));
	jdff g1432(.din(w_G2211_0[0]),.dout(w_dff_A_56ni4neV6_1));
	jdff g1433(.din(w_G4394_0[1]),.dout(w_dff_A_sAMargQa3_1));
	jdff g1434(.din(w_G1_0[2]),.dout(w_dff_A_15oUKSIM7_1));
	jdff g1435(.din(w_G106_0[1]),.dout(w_dff_A_FqMa6rxn5_1));
	jnot g1436(.din(w_G15_0[1]),.dout(w_dff_A_x6qNQfhM0_1),.clk(gclk));
	jor g1437(.dina(w_n345_0[0]),.dinb(w_G5_0[2]),.dout(w_dff_A_WJXAWJxz0_2),.clk(gclk));
	jnot g1438(.din(w_G15_0[0]),.dout(w_dff_A_BPLu96TO4_1),.clk(gclk));
	jor g1439(.dina(w_n349_0[0]),.dinb(w_G5_0[1]),.dout(w_dff_A_GX6m9gnD6_2),.clk(gclk));
	jdff g1440(.din(w_G1_0[1]),.dout(w_dff_A_Af8wiAcQ9_1));
	jand g1441(.dina(w_n1125_0[1]),.dinb(w_n1122_0[1]),.dout(w_dff_A_slq4IEGl3_2),.clk(gclk));
	jor g1442(.dina(w_n720_1[0]),.dinb(w_n716_1[0]),.dout(w_dff_A_xynYSXoD0_2),.clk(gclk));
	jand g1443(.dina(w_n1125_0[0]),.dinb(w_n1122_0[0]),.dout(w_dff_A_uIYyqE1Q1_2),.clk(gclk));
	jor g1444(.dina(w_n720_0[2]),.dinb(w_n716_0[2]),.dout(w_dff_A_L1Bufp9g1_2),.clk(gclk));
	jor g1445(.dina(w_n720_0[1]),.dinb(w_n716_0[1]),.dout(w_dff_A_jO93Ve3B1_2),.clk(gclk));
	jand g1446(.dina(w_n1465_0[0]),.dinb(w_n715_0[0]),.dout(w_dff_A_1dn7niiP8_2),.clk(gclk));
	jxor g1447(.dina(w_n713_0[1]),.dinb(w_n709_0[1]),.dout(w_dff_A_RbZnUKx60_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G5_0(.douta(w_G5_0[0]),.doutb(w_dff_A_nZ0M8cl96_1),.doutc(w_dff_A_trt7Zdp61_2),.din(G5));
	jspl3 jspl3_w_G5_1(.douta(w_dff_A_7yeiBPBK4_0),.doutb(w_dff_A_UczSuiSW2_1),.doutc(w_G5_1[2]),.din(w_G5_0[0]));
	jspl3 jspl3_w_G15_0(.douta(w_G15_0[0]),.doutb(w_G15_0[1]),.doutc(w_G15_0[2]),.din(G15));
	jspl3 jspl3_w_G18_0(.douta(w_G18_0[0]),.doutb(w_G18_0[1]),.doutc(w_G18_0[2]),.din(G18));
	jspl3 jspl3_w_G18_1(.douta(w_G18_1[0]),.doutb(w_G18_1[1]),.doutc(w_G18_1[2]),.din(w_G18_0[0]));
	jspl3 jspl3_w_G18_2(.douta(w_G18_2[0]),.doutb(w_G18_2[1]),.doutc(w_G18_2[2]),.din(w_G18_0[1]));
	jspl3 jspl3_w_G18_3(.douta(w_G18_3[0]),.doutb(w_G18_3[1]),.doutc(w_G18_3[2]),.din(w_G18_0[2]));
	jspl3 jspl3_w_G18_4(.douta(w_G18_4[0]),.doutb(w_G18_4[1]),.doutc(w_G18_4[2]),.din(w_G18_1[0]));
	jspl3 jspl3_w_G18_5(.douta(w_G18_5[0]),.doutb(w_G18_5[1]),.doutc(w_G18_5[2]),.din(w_G18_1[1]));
	jspl3 jspl3_w_G18_6(.douta(w_G18_6[0]),.doutb(w_G18_6[1]),.doutc(w_G18_6[2]),.din(w_G18_1[2]));
	jspl3 jspl3_w_G18_7(.douta(w_G18_7[0]),.doutb(w_G18_7[1]),.doutc(w_G18_7[2]),.din(w_G18_2[0]));
	jspl3 jspl3_w_G18_8(.douta(w_G18_8[0]),.doutb(w_G18_8[1]),.doutc(w_G18_8[2]),.din(w_G18_2[1]));
	jspl3 jspl3_w_G18_9(.douta(w_G18_9[0]),.doutb(w_G18_9[1]),.doutc(w_G18_9[2]),.din(w_G18_2[2]));
	jspl3 jspl3_w_G18_10(.douta(w_G18_10[0]),.doutb(w_G18_10[1]),.doutc(w_G18_10[2]),.din(w_G18_3[0]));
	jspl3 jspl3_w_G18_11(.douta(w_G18_11[0]),.doutb(w_G18_11[1]),.doutc(w_G18_11[2]),.din(w_G18_3[1]));
	jspl3 jspl3_w_G18_12(.douta(w_G18_12[0]),.doutb(w_G18_12[1]),.doutc(w_G18_12[2]),.din(w_G18_3[2]));
	jspl3 jspl3_w_G18_13(.douta(w_G18_13[0]),.doutb(w_G18_13[1]),.doutc(w_G18_13[2]),.din(w_G18_4[0]));
	jspl3 jspl3_w_G18_14(.douta(w_G18_14[0]),.doutb(w_G18_14[1]),.doutc(w_G18_14[2]),.din(w_G18_4[1]));
	jspl3 jspl3_w_G18_15(.douta(w_G18_15[0]),.doutb(w_G18_15[1]),.doutc(w_G18_15[2]),.din(w_G18_4[2]));
	jspl3 jspl3_w_G18_16(.douta(w_G18_16[0]),.doutb(w_G18_16[1]),.doutc(w_G18_16[2]),.din(w_G18_5[0]));
	jspl3 jspl3_w_G18_17(.douta(w_G18_17[0]),.doutb(w_G18_17[1]),.doutc(w_G18_17[2]),.din(w_G18_5[1]));
	jspl3 jspl3_w_G18_18(.douta(w_G18_18[0]),.doutb(w_G18_18[1]),.doutc(w_G18_18[2]),.din(w_G18_5[2]));
	jspl3 jspl3_w_G18_19(.douta(w_G18_19[0]),.doutb(w_G18_19[1]),.doutc(w_G18_19[2]),.din(w_G18_6[0]));
	jspl3 jspl3_w_G18_20(.douta(w_G18_20[0]),.doutb(w_G18_20[1]),.doutc(w_G18_20[2]),.din(w_G18_6[1]));
	jspl3 jspl3_w_G18_21(.douta(w_G18_21[0]),.doutb(w_G18_21[1]),.doutc(w_G18_21[2]),.din(w_G18_6[2]));
	jspl3 jspl3_w_G18_22(.douta(w_G18_22[0]),.doutb(w_G18_22[1]),.doutc(w_G18_22[2]),.din(w_G18_7[0]));
	jspl3 jspl3_w_G18_23(.douta(w_G18_23[0]),.doutb(w_G18_23[1]),.doutc(w_G18_23[2]),.din(w_G18_7[1]));
	jspl3 jspl3_w_G18_24(.douta(w_G18_24[0]),.doutb(w_G18_24[1]),.doutc(w_G18_24[2]),.din(w_G18_7[2]));
	jspl3 jspl3_w_G18_25(.douta(w_G18_25[0]),.doutb(w_G18_25[1]),.doutc(w_G18_25[2]),.din(w_G18_8[0]));
	jspl3 jspl3_w_G18_26(.douta(w_G18_26[0]),.doutb(w_G18_26[1]),.doutc(w_G18_26[2]),.din(w_G18_8[1]));
	jspl3 jspl3_w_G18_27(.douta(w_G18_27[0]),.doutb(w_G18_27[1]),.doutc(w_G18_27[2]),.din(w_G18_8[2]));
	jspl3 jspl3_w_G18_28(.douta(w_G18_28[0]),.doutb(w_G18_28[1]),.doutc(w_G18_28[2]),.din(w_G18_9[0]));
	jspl3 jspl3_w_G18_29(.douta(w_G18_29[0]),.doutb(w_G18_29[1]),.doutc(w_G18_29[2]),.din(w_G18_9[1]));
	jspl3 jspl3_w_G18_30(.douta(w_G18_30[0]),.doutb(w_G18_30[1]),.doutc(w_G18_30[2]),.din(w_G18_9[2]));
	jspl3 jspl3_w_G18_31(.douta(w_G18_31[0]),.doutb(w_G18_31[1]),.doutc(w_G18_31[2]),.din(w_G18_10[0]));
	jspl3 jspl3_w_G18_32(.douta(w_G18_32[0]),.doutb(w_G18_32[1]),.doutc(w_G18_32[2]),.din(w_G18_10[1]));
	jspl3 jspl3_w_G18_33(.douta(w_G18_33[0]),.doutb(w_G18_33[1]),.doutc(w_G18_33[2]),.din(w_G18_10[2]));
	jspl3 jspl3_w_G18_34(.douta(w_G18_34[0]),.doutb(w_G18_34[1]),.doutc(w_G18_34[2]),.din(w_G18_11[0]));
	jspl3 jspl3_w_G18_35(.douta(w_G18_35[0]),.doutb(w_G18_35[1]),.doutc(w_G18_35[2]),.din(w_G18_11[1]));
	jspl3 jspl3_w_G18_36(.douta(w_G18_36[0]),.doutb(w_G18_36[1]),.doutc(w_G18_36[2]),.din(w_G18_11[2]));
	jspl3 jspl3_w_G18_37(.douta(w_G18_37[0]),.doutb(w_G18_37[1]),.doutc(w_G18_37[2]),.din(w_G18_12[0]));
	jspl3 jspl3_w_G18_38(.douta(w_G18_38[0]),.doutb(w_G18_38[1]),.doutc(w_G18_38[2]),.din(w_G18_12[1]));
	jspl3 jspl3_w_G18_39(.douta(w_G18_39[0]),.doutb(w_G18_39[1]),.doutc(w_G18_39[2]),.din(w_G18_12[2]));
	jspl3 jspl3_w_G18_40(.douta(w_G18_40[0]),.doutb(w_G18_40[1]),.doutc(w_G18_40[2]),.din(w_G18_13[0]));
	jspl3 jspl3_w_G18_41(.douta(w_G18_41[0]),.doutb(w_G18_41[1]),.doutc(w_G18_41[2]),.din(w_G18_13[1]));
	jspl3 jspl3_w_G18_42(.douta(w_G18_42[0]),.doutb(w_G18_42[1]),.doutc(w_G18_42[2]),.din(w_G18_13[2]));
	jspl3 jspl3_w_G18_43(.douta(w_G18_43[0]),.doutb(w_G18_43[1]),.doutc(w_G18_43[2]),.din(w_G18_14[0]));
	jspl3 jspl3_w_G18_44(.douta(w_G18_44[0]),.doutb(w_G18_44[1]),.doutc(w_G18_44[2]),.din(w_G18_14[1]));
	jspl3 jspl3_w_G18_45(.douta(w_G18_45[0]),.doutb(w_G18_45[1]),.doutc(w_G18_45[2]),.din(w_G18_14[2]));
	jspl3 jspl3_w_G18_46(.douta(w_G18_46[0]),.doutb(w_G18_46[1]),.doutc(w_G18_46[2]),.din(w_G18_15[0]));
	jspl3 jspl3_w_G18_47(.douta(w_G18_47[0]),.doutb(w_G18_47[1]),.doutc(w_G18_47[2]),.din(w_G18_15[1]));
	jspl3 jspl3_w_G18_48(.douta(w_G18_48[0]),.doutb(w_G18_48[1]),.doutc(w_G18_48[2]),.din(w_G18_15[2]));
	jspl3 jspl3_w_G18_49(.douta(w_G18_49[0]),.doutb(w_G18_49[1]),.doutc(w_G18_49[2]),.din(w_G18_16[0]));
	jspl3 jspl3_w_G18_50(.douta(w_G18_50[0]),.doutb(w_G18_50[1]),.doutc(w_G18_50[2]),.din(w_G18_16[1]));
	jspl3 jspl3_w_G18_51(.douta(w_G18_51[0]),.doutb(w_G18_51[1]),.doutc(w_G18_51[2]),.din(w_G18_16[2]));
	jspl3 jspl3_w_G18_52(.douta(w_G18_52[0]),.doutb(w_G18_52[1]),.doutc(w_G18_52[2]),.din(w_G18_17[0]));
	jspl3 jspl3_w_G18_53(.douta(w_G18_53[0]),.doutb(w_G18_53[1]),.doutc(w_G18_53[2]),.din(w_G18_17[1]));
	jspl3 jspl3_w_G18_54(.douta(w_G18_54[0]),.doutb(w_G18_54[1]),.doutc(w_G18_54[2]),.din(w_G18_17[2]));
	jspl3 jspl3_w_G18_55(.douta(w_G18_55[0]),.doutb(w_G18_55[1]),.doutc(w_G18_55[2]),.din(w_G18_18[0]));
	jspl3 jspl3_w_G18_56(.douta(w_G18_56[0]),.doutb(w_G18_56[1]),.doutc(w_G18_56[2]),.din(w_G18_18[1]));
	jspl3 jspl3_w_G18_57(.douta(w_G18_57[0]),.doutb(w_G18_57[1]),.doutc(w_G18_57[2]),.din(w_G18_18[2]));
	jspl3 jspl3_w_G18_58(.douta(w_G18_58[0]),.doutb(w_G18_58[1]),.doutc(w_G18_58[2]),.din(w_G18_19[0]));
	jspl3 jspl3_w_G38_0(.douta(w_G38_0[0]),.doutb(w_G38_0[1]),.doutc(w_G38_0[2]),.din(G38));
	jspl3 jspl3_w_G38_1(.douta(w_G38_1[0]),.doutb(w_G38_1[1]),.doutc(w_G38_1[2]),.din(w_G38_0[0]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_G41_0[1]),.doutc(w_G41_0[2]),.din(G41));
	jspl jspl_w_G69_0(.douta(w_G69_0[0]),.doutb(w_G69_0[1]),.din(G69));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(G70));
	jspl3 jspl3_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.doutc(w_G106_0[2]),.din(G106));
	jspl jspl_w_G106_1(.douta(w_G106_1[0]),.doutb(w_G106_1[1]),.din(w_G106_0[0]));
	jspl jspl_w_G229_0(.douta(w_G229_0[0]),.doutb(w_G229_0[1]),.din(G229));
	jspl3 jspl3_w_G1455_0(.douta(w_G1455_0[0]),.doutb(w_G1455_0[1]),.doutc(w_G1455_0[2]),.din(G1455));
	jspl jspl_w_G1459_0(.douta(w_G1459_0[0]),.doutb(w_G1459_0[1]),.din(G1459));
	jspl3 jspl3_w_G1462_0(.douta(w_G1462_0[0]),.doutb(w_G1462_0[1]),.doutc(w_G1462_0[2]),.din(G1462));
	jspl3 jspl3_w_G1469_0(.douta(w_G1469_0[0]),.doutb(w_G1469_0[1]),.doutc(w_G1469_0[2]),.din(G1469));
	jspl jspl_w_G1469_1(.douta(w_G1469_1[0]),.doutb(w_G1469_1[1]),.din(w_G1469_0[0]));
	jspl3 jspl3_w_G1480_0(.douta(w_G1480_0[0]),.doutb(w_G1480_0[1]),.doutc(w_G1480_0[2]),.din(G1480));
	jspl3 jspl3_w_G1486_0(.douta(w_G1486_0[0]),.doutb(w_G1486_0[1]),.doutc(w_G1486_0[2]),.din(G1486));
	jspl3 jspl3_w_G1492_0(.douta(w_G1492_0[0]),.doutb(w_G1492_0[1]),.doutc(w_G1492_0[2]),.din(G1492));
	jspl jspl_w_G1492_1(.douta(w_G1492_1[0]),.doutb(w_G1492_1[1]),.din(w_G1492_0[0]));
	jspl3 jspl3_w_G1496_0(.douta(w_G1496_0[0]),.doutb(w_G1496_0[1]),.doutc(w_G1496_0[2]),.din(G1496));
	jspl3 jspl3_w_G2204_0(.douta(w_G2204_0[0]),.doutb(w_G2204_0[1]),.doutc(w_G2204_0[2]),.din(G2204));
	jspl jspl_w_G2208_0(.douta(w_G2208_0[0]),.doutb(w_G2208_0[1]),.din(G2208));
	jspl3 jspl3_w_G2211_0(.douta(w_G2211_0[0]),.doutb(w_G2211_0[1]),.doutc(w_G2211_0[2]),.din(G2211));
	jspl3 jspl3_w_G2218_0(.douta(w_G2218_0[0]),.doutb(w_G2218_0[1]),.doutc(w_G2218_0[2]),.din(G2218));
	jspl3 jspl3_w_G2224_0(.douta(w_G2224_0[0]),.doutb(w_G2224_0[1]),.doutc(w_G2224_0[2]),.din(G2224));
	jspl jspl_w_G2224_1(.douta(w_G2224_1[0]),.doutb(w_G2224_1[1]),.din(w_G2224_0[0]));
	jspl3 jspl3_w_G2230_0(.douta(w_G2230_0[0]),.doutb(w_G2230_0[1]),.doutc(w_G2230_0[2]),.din(G2230));
	jspl jspl_w_G2230_1(.douta(w_G2230_1[0]),.doutb(w_G2230_1[1]),.din(w_G2230_0[0]));
	jspl3 jspl3_w_G2236_0(.douta(w_G2236_0[0]),.doutb(w_G2236_0[1]),.doutc(w_G2236_0[2]),.din(G2236));
	jspl jspl_w_G2236_1(.douta(w_G2236_1[0]),.doutb(w_G2236_1[1]),.din(w_G2236_0[0]));
	jspl3 jspl3_w_G2239_0(.douta(w_G2239_0[0]),.doutb(w_G2239_0[1]),.doutc(w_G2239_0[2]),.din(G2239));
	jspl3 jspl3_w_G2247_0(.douta(w_G2247_0[0]),.doutb(w_G2247_0[1]),.doutc(w_G2247_0[2]),.din(G2247));
	jspl3 jspl3_w_G2253_0(.douta(w_G2253_0[0]),.doutb(w_G2253_0[1]),.doutc(w_G2253_0[2]),.din(G2253));
	jspl jspl_w_G2253_1(.douta(w_G2253_1[0]),.doutb(w_G2253_1[1]),.din(w_G2253_0[0]));
	jspl3 jspl3_w_G2256_0(.douta(w_G2256_0[0]),.doutb(w_G2256_0[1]),.doutc(w_G2256_0[2]),.din(G2256));
	jspl jspl_w_G2256_1(.douta(w_G2256_1[0]),.doutb(w_G2256_1[1]),.din(w_G2256_0[0]));
	jspl jspl_w_G3698_0(.douta(w_G3698_0[0]),.doutb(w_G3698_0[1]),.din(G3698));
	jspl3 jspl3_w_G3701_0(.douta(w_G3701_0[0]),.doutb(w_G3701_0[1]),.doutc(w_G3701_0[2]),.din(G3701));
	jspl jspl_w_G3701_1(.douta(w_G3701_1[0]),.doutb(w_G3701_1[1]),.din(w_G3701_0[0]));
	jspl3 jspl3_w_G3705_0(.douta(w_G3705_0[0]),.doutb(w_G3705_0[1]),.doutc(w_G3705_0[2]),.din(G3705));
	jspl3 jspl3_w_G3705_1(.douta(w_G3705_1[0]),.doutb(w_G3705_1[1]),.doutc(w_G3705_1[2]),.din(w_G3705_0[0]));
	jspl jspl_w_G3705_2(.douta(w_G3705_2[0]),.doutb(w_G3705_2[1]),.din(w_G3705_0[1]));
	jspl3 jspl3_w_G3711_0(.douta(w_G3711_0[0]),.doutb(w_G3711_0[1]),.doutc(w_G3711_0[2]),.din(G3711));
	jspl jspl_w_G3711_1(.douta(w_G3711_1[0]),.doutb(w_G3711_1[1]),.din(w_G3711_0[0]));
	jspl3 jspl3_w_G3717_0(.douta(w_G3717_0[0]),.doutb(w_G3717_0[1]),.doutc(w_G3717_0[2]),.din(G3717));
	jspl3 jspl3_w_G3717_1(.douta(w_G3717_1[0]),.doutb(w_G3717_1[1]),.doutc(w_G3717_1[2]),.din(w_G3717_0[0]));
	jspl jspl_w_G3717_2(.douta(w_G3717_2[0]),.doutb(w_G3717_2[1]),.din(w_G3717_0[1]));
	jspl3 jspl3_w_G3723_0(.douta(w_G3723_0[0]),.doutb(w_G3723_0[1]),.doutc(w_G3723_0[2]),.din(G3723));
	jspl jspl_w_G3723_1(.douta(w_G3723_1[0]),.doutb(w_G3723_1[1]),.din(w_G3723_0[0]));
	jspl3 jspl3_w_G3729_0(.douta(w_G3729_0[0]),.doutb(w_G3729_0[1]),.doutc(w_G3729_0[2]),.din(G3729));
	jspl jspl_w_G3729_1(.douta(w_G3729_1[0]),.doutb(w_G3729_1[1]),.din(w_G3729_0[0]));
	jspl3 jspl3_w_G3737_0(.douta(w_G3737_0[0]),.doutb(w_G3737_0[1]),.doutc(w_G3737_0[2]),.din(G3737));
	jspl jspl_w_G3737_1(.douta(w_G3737_1[0]),.doutb(w_G3737_1[1]),.din(w_G3737_0[0]));
	jspl3 jspl3_w_G3743_0(.douta(w_G3743_0[0]),.doutb(w_G3743_0[1]),.doutc(w_G3743_0[2]),.din(G3743));
	jspl3 jspl3_w_G3743_1(.douta(w_G3743_1[0]),.doutb(w_G3743_1[1]),.doutc(w_G3743_1[2]),.din(w_G3743_0[0]));
	jspl3 jspl3_w_G3749_0(.douta(w_G3749_0[0]),.doutb(w_G3749_0[1]),.doutc(w_G3749_0[2]),.din(G3749));
	jspl jspl_w_G3749_1(.douta(w_G3749_1[0]),.doutb(w_G3749_1[1]),.din(w_G3749_0[0]));
	jspl jspl_w_G4393_0(.douta(w_G4393_0[0]),.doutb(w_G4393_0[1]),.din(G4393));
	jspl3 jspl3_w_G4394_0(.douta(w_G4394_0[0]),.doutb(w_G4394_0[1]),.doutc(w_G4394_0[2]),.din(G4394));
	jspl jspl_w_G4394_1(.douta(w_G4394_1[0]),.doutb(w_G4394_1[1]),.din(w_G4394_0[0]));
	jspl3 jspl3_w_G4400_0(.douta(w_G4400_0[0]),.doutb(w_G4400_0[1]),.doutc(w_G4400_0[2]),.din(G4400));
	jspl3 jspl3_w_G4405_0(.douta(w_G4405_0[0]),.doutb(w_G4405_0[1]),.doutc(w_G4405_0[2]),.din(G4405));
	jspl3 jspl3_w_G4405_1(.douta(w_G4405_1[0]),.doutb(w_G4405_1[1]),.doutc(w_G4405_1[2]),.din(w_G4405_0[0]));
	jspl3 jspl3_w_G4410_0(.douta(w_G4410_0[0]),.doutb(w_G4410_0[1]),.doutc(w_G4410_0[2]),.din(G4410));
	jspl jspl_w_G4410_1(.douta(w_G4410_1[0]),.doutb(w_G4410_1[1]),.din(w_G4410_0[0]));
	jspl3 jspl3_w_G4415_0(.douta(w_G4415_0[0]),.doutb(w_G4415_0[1]),.doutc(w_G4415_0[2]),.din(G4415));
	jspl jspl_w_G4415_1(.douta(w_G4415_1[0]),.doutb(w_G4415_1[1]),.din(w_G4415_0[0]));
	jspl3 jspl3_w_G4420_0(.douta(w_G4420_0[0]),.doutb(w_G4420_0[1]),.doutc(w_G4420_0[2]),.din(G4420));
	jspl jspl_w_G4427_0(.douta(w_G4427_0[0]),.doutb(w_G4427_0[1]),.din(G4427));
	jspl3 jspl3_w_G4432_0(.douta(w_G4432_0[0]),.doutb(w_G4432_0[1]),.doutc(w_G4432_0[2]),.din(G4432));
	jspl jspl_w_G4432_1(.douta(w_G4432_1[0]),.doutb(w_G4432_1[1]),.din(w_G4432_0[0]));
	jspl3 jspl3_w_G4437_0(.douta(w_G4437_0[0]),.doutb(w_G4437_0[1]),.doutc(w_G4437_0[2]),.din(G4437));
	jspl3 jspl3_w_G4526_0(.douta(w_G4526_0[0]),.doutb(w_G4526_0[1]),.doutc(w_G4526_0[2]),.din(G4526));
	jspl jspl_w_G4526_1(.douta(w_G4526_1[0]),.doutb(w_G4526_1[1]),.din(w_G4526_0[0]));
	jspl3 jspl3_w_G4528_0(.douta(w_G4528_0[0]),.doutb(w_G4528_0[1]),.doutc(w_G4528_0[2]),.din(G4528));
	jspl jspl_w_G404_0(.douta(w_G404_0),.doutb(w_dff_A_SGEwqHKw4_1),.din(G404_fa_));
	jspl jspl_w_G406_0(.douta(w_G406_0),.doutb(w_dff_A_J25vNCWP8_1),.din(G406_fa_));
	jspl jspl_w_G408_0(.douta(w_G408_0),.doutb(w_dff_A_6zPirW7D7_1),.din(G408_fa_));
	jspl jspl_w_G410_0(.douta(w_G410_0),.doutb(w_dff_A_NzXdC8ZK7_1),.din(G410_fa_));
	jspl jspl_w_G412_0(.douta(w_G412_0),.doutb(w_dff_A_lCOwNbj03_1),.din(G412_fa_));
	jspl jspl_w_G414_0(.douta(w_dff_A_qE6J2TTm7_0),.doutb(w_dff_A_sj0YHAtv4_1),.din(G414_fa_));
	jspl jspl_w_G416_0(.douta(w_G416_0),.doutb(w_dff_A_pXJgTd7U2_1),.din(G416_fa_));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(n345));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl3 jspl3_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.doutc(w_n353_0[2]),.din(n353));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_n354_0[2]),.din(n354));
	jspl3 jspl3_w_n354_1(.douta(w_n354_1[0]),.doutb(w_n354_1[1]),.doutc(w_n354_1[2]),.din(w_n354_0[0]));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl3 jspl3_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.doutc(w_n355_1[2]),.din(w_n355_0[0]));
	jspl3 jspl3_w_n355_2(.douta(w_n355_2[0]),.doutb(w_n355_2[1]),.doutc(w_n355_2[2]),.din(w_n355_0[1]));
	jspl3 jspl3_w_n355_3(.douta(w_n355_3[0]),.doutb(w_n355_3[1]),.doutc(w_n355_3[2]),.din(w_n355_0[2]));
	jspl3 jspl3_w_n355_4(.douta(w_n355_4[0]),.doutb(w_n355_4[1]),.doutc(w_n355_4[2]),.din(w_n355_1[0]));
	jspl3 jspl3_w_n355_5(.douta(w_n355_5[0]),.doutb(w_n355_5[1]),.doutc(w_n355_5[2]),.din(w_n355_1[1]));
	jspl3 jspl3_w_n355_6(.douta(w_n355_6[0]),.doutb(w_n355_6[1]),.doutc(w_n355_6[2]),.din(w_n355_1[2]));
	jspl3 jspl3_w_n355_7(.douta(w_n355_7[0]),.doutb(w_n355_7[1]),.doutc(w_n355_7[2]),.din(w_n355_2[0]));
	jspl3 jspl3_w_n355_8(.douta(w_n355_8[0]),.doutb(w_n355_8[1]),.doutc(w_n355_8[2]),.din(w_n355_2[1]));
	jspl3 jspl3_w_n355_9(.douta(w_n355_9[0]),.doutb(w_n355_9[1]),.doutc(w_n355_9[2]),.din(w_n355_2[2]));
	jspl3 jspl3_w_n355_10(.douta(w_n355_10[0]),.doutb(w_n355_10[1]),.doutc(w_n355_10[2]),.din(w_n355_3[0]));
	jspl3 jspl3_w_n355_11(.douta(w_n355_11[0]),.doutb(w_n355_11[1]),.doutc(w_n355_11[2]),.din(w_n355_3[1]));
	jspl3 jspl3_w_n355_12(.douta(w_n355_12[0]),.doutb(w_n355_12[1]),.doutc(w_n355_12[2]),.din(w_n355_3[2]));
	jspl3 jspl3_w_n355_13(.douta(w_n355_13[0]),.doutb(w_n355_13[1]),.doutc(w_n355_13[2]),.din(w_n355_4[0]));
	jspl3 jspl3_w_n355_14(.douta(w_n355_14[0]),.doutb(w_n355_14[1]),.doutc(w_n355_14[2]),.din(w_n355_4[1]));
	jspl3 jspl3_w_n355_15(.douta(w_n355_15[0]),.doutb(w_n355_15[1]),.doutc(w_n355_15[2]),.din(w_n355_4[2]));
	jspl3 jspl3_w_n355_16(.douta(w_n355_16[0]),.doutb(w_n355_16[1]),.doutc(w_n355_16[2]),.din(w_n355_5[0]));
	jspl3 jspl3_w_n355_17(.douta(w_n355_17[0]),.doutb(w_n355_17[1]),.doutc(w_n355_17[2]),.din(w_n355_5[1]));
	jspl3 jspl3_w_n355_18(.douta(w_n355_18[0]),.doutb(w_n355_18[1]),.doutc(w_n355_18[2]),.din(w_n355_5[2]));
	jspl3 jspl3_w_n355_19(.douta(w_n355_19[0]),.doutb(w_n355_19[1]),.doutc(w_n355_19[2]),.din(w_n355_6[0]));
	jspl3 jspl3_w_n355_20(.douta(w_n355_20[0]),.doutb(w_n355_20[1]),.doutc(w_n355_20[2]),.din(w_n355_6[1]));
	jspl3 jspl3_w_n355_21(.douta(w_n355_21[0]),.doutb(w_n355_21[1]),.doutc(w_n355_21[2]),.din(w_n355_6[2]));
	jspl3 jspl3_w_n355_22(.douta(w_n355_22[0]),.doutb(w_n355_22[1]),.doutc(w_n355_22[2]),.din(w_n355_7[0]));
	jspl3 jspl3_w_n355_23(.douta(w_n355_23[0]),.doutb(w_n355_23[1]),.doutc(w_n355_23[2]),.din(w_n355_7[1]));
	jspl3 jspl3_w_n355_24(.douta(w_n355_24[0]),.doutb(w_n355_24[1]),.doutc(w_n355_24[2]),.din(w_n355_7[2]));
	jspl3 jspl3_w_n355_25(.douta(w_n355_25[0]),.doutb(w_n355_25[1]),.doutc(w_n355_25[2]),.din(w_n355_8[0]));
	jspl jspl_w_n355_26(.douta(w_n355_26[0]),.doutb(w_n355_26[1]),.din(w_n355_8[1]));
	jspl3 jspl3_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.doutc(w_n356_0[2]),.din(n356));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(n358));
	jspl jspl_w_n359_0(.douta(w_n359_0[0]),.doutb(w_n359_0[1]),.din(n359));
	jspl3 jspl3_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.doutc(w_n362_0[2]),.din(n362));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(n366));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(n370));
	jspl3 jspl3_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.doutc(w_n371_0[2]),.din(n371));
	jspl jspl_w_n371_1(.douta(w_n371_1[0]),.doutb(w_n371_1[1]),.din(w_n371_0[0]));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.doutc(w_n372_0[2]),.din(n372));
	jspl3 jspl3_w_n372_1(.douta(w_n372_1[0]),.doutb(w_n372_1[1]),.doutc(w_n372_1[2]),.din(w_n372_0[0]));
	jspl jspl_w_n376_0(.douta(w_n376_0[0]),.doutb(w_n376_0[1]),.din(n376));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_n377_0[2]),.din(n377));
	jspl3 jspl3_w_n377_1(.douta(w_n377_1[0]),.doutb(w_n377_1[1]),.doutc(w_n377_1[2]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n379_0(.douta(w_n379_0[0]),.doutb(w_n379_0[1]),.doutc(w_n379_0[2]),.din(n379));
	jspl jspl_w_n379_1(.douta(w_n379_1[0]),.doutb(w_n379_1[1]),.din(w_n379_0[0]));
	jspl3 jspl3_w_n380_0(.douta(w_n380_0[0]),.doutb(w_n380_0[1]),.doutc(w_n380_0[2]),.din(n380));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl3 jspl3_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.doutc(w_n387_1[2]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_n388_0[2]),.din(n388));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.din(n389));
	jspl3 jspl3_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.doutc(w_n390_0[2]),.din(n390));
	jspl jspl_w_n390_1(.douta(w_n390_1[0]),.doutb(w_n390_1[1]),.din(w_n390_0[0]));
	jspl3 jspl3_w_n395_0(.douta(w_n395_0[0]),.doutb(w_n395_0[1]),.doutc(w_n395_0[2]),.din(n395));
	jspl jspl_w_n400_0(.douta(w_n400_0[0]),.doutb(w_n400_0[1]),.din(n400));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n401_1(.douta(w_n401_1[0]),.doutb(w_n401_1[1]),.doutc(w_n401_1[2]),.din(w_n401_0[0]));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl jspl_w_n402_1(.douta(w_n402_1[0]),.doutb(w_n402_1[1]),.din(w_n402_0[0]));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl jspl_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.din(n404));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl3 jspl3_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.doutc(w_n407_0[2]),.din(n407));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl jspl_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.din(n410));
	jspl3 jspl3_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.doutc(w_n412_0[2]),.din(n412));
	jspl3 jspl3_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.doutc(w_n413_0[2]),.din(n413));
	jspl jspl_w_n413_1(.douta(w_n413_1[0]),.doutb(w_n413_1[1]),.din(w_n413_0[0]));
	jspl3 jspl3_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.doutc(w_n417_0[2]),.din(n417));
	jspl jspl_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.din(n419));
	jspl3 jspl3_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.doutc(w_n422_0[2]),.din(n422));
	jspl3 jspl3_w_n422_1(.douta(w_n422_1[0]),.doutb(w_n422_1[1]),.doutc(w_n422_1[2]),.din(w_n422_0[0]));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(n427));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.doutc(w_n428_0[2]),.din(n428));
	jspl3 jspl3_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.doutc(w_n429_0[2]),.din(n429));
	jspl3 jspl3_w_n429_1(.douta(w_n429_1[0]),.doutb(w_n429_1[1]),.doutc(w_n429_1[2]),.din(w_n429_0[0]));
	jspl jspl_w_n429_2(.douta(w_n429_2[0]),.doutb(w_n429_2[1]),.din(w_n429_0[1]));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl jspl_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.din(w_n435_0[0]));
	jspl jspl_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.din(n436));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl3 jspl3_w_n442_0(.douta(w_n442_0[0]),.doutb(w_n442_0[1]),.doutc(w_n442_0[2]),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.doutc(w_n446_0[2]),.din(n446));
	jspl jspl_w_n446_1(.douta(w_n446_1[0]),.doutb(w_n446_1[1]),.din(w_n446_0[0]));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.din(n448));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n450_0(.douta(w_n450_0[0]),.doutb(w_n450_0[1]),.doutc(w_n450_0[2]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n454_0(.douta(w_n454_0[0]),.doutb(w_n454_0[1]),.din(n454));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.din(n455));
	jspl3 jspl3_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.doutc(w_n456_0[2]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n458_0(.douta(w_n458_0[0]),.doutb(w_n458_0[1]),.doutc(w_n458_0[2]),.din(n458));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl jspl_w_n461_0(.douta(w_n461_0[0]),.doutb(w_n461_0[1]),.din(n461));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(n464));
	jspl3 jspl3_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.doutc(w_n465_0[2]),.din(n465));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(n466));
	jspl jspl_w_n468_0(.douta(w_n468_0[0]),.doutb(w_n468_0[1]),.din(n468));
	jspl3 jspl3_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.doutc(w_n469_0[2]),.din(n469));
	jspl jspl_w_n469_1(.douta(w_n469_1[0]),.doutb(w_n469_1[1]),.din(w_n469_0[0]));
	jspl3 jspl3_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.doutc(w_n470_0[2]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl jspl_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.din(n473));
	jspl3 jspl3_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.doutc(w_n474_0[2]),.din(n474));
	jspl jspl_w_n474_1(.douta(w_n474_1[0]),.doutb(w_n474_1[1]),.din(w_n474_0[0]));
	jspl3 jspl3_w_n475_0(.douta(w_n475_0[0]),.doutb(w_n475_0[1]),.doutc(w_n475_0[2]),.din(n475));
	jspl jspl_w_n475_1(.douta(w_n475_1[0]),.doutb(w_n475_1[1]),.din(w_n475_0[0]));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(n479));
	jspl3 jspl3_w_n480_0(.douta(w_n480_0[0]),.doutb(w_n480_0[1]),.doutc(w_n480_0[2]),.din(n480));
	jspl jspl_w_n480_1(.douta(w_n480_1[0]),.doutb(w_n480_1[1]),.din(w_n480_0[0]));
	jspl3 jspl3_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.doutc(w_n481_0[2]),.din(n481));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl3 jspl3_w_n485_0(.douta(w_n485_0[0]),.doutb(w_n485_0[1]),.doutc(w_n485_0[2]),.din(n485));
	jspl3 jspl3_w_n486_0(.douta(w_n486_0[0]),.doutb(w_n486_0[1]),.doutc(w_n486_0[2]),.din(n486));
	jspl jspl_w_n488_0(.douta(w_n488_0[0]),.doutb(w_n488_0[1]),.din(n488));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(n489));
	jspl3 jspl3_w_n490_0(.douta(w_n490_0[0]),.doutb(w_n490_0[1]),.doutc(w_n490_0[2]),.din(n490));
	jspl3 jspl3_w_n491_0(.douta(w_n491_0[0]),.doutb(w_n491_0[1]),.doutc(w_n491_0[2]),.din(n491));
	jspl jspl_w_n491_1(.douta(w_n491_1[0]),.doutb(w_n491_1[1]),.din(w_n491_0[0]));
	jspl jspl_w_n493_0(.douta(w_n493_0[0]),.doutb(w_n493_0[1]),.din(n493));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl jspl_w_n503_0(.douta(w_n503_0[0]),.doutb(w_n503_0[1]),.din(n503));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(n509));
	jspl jspl_w_n510_0(.douta(w_n510_0[0]),.doutb(w_n510_0[1]),.din(n510));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl3 jspl3_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.doutc(w_n514_0[2]),.din(n514));
	jspl3 jspl3_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.doutc(w_n516_0[2]),.din(n516));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(n519));
	jspl3 jspl3_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.doutc(w_n520_0[2]),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.doutc(w_n523_0[2]),.din(n523));
	jspl3 jspl3_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.doutc(w_n524_0[2]),.din(n524));
	jspl3 jspl3_w_n524_1(.douta(w_n524_1[0]),.doutb(w_n524_1[1]),.doutc(w_n524_1[2]),.din(w_n524_0[0]));
	jspl jspl_w_n524_2(.douta(w_n524_2[0]),.doutb(w_n524_2[1]),.din(w_n524_0[1]));
	jspl3 jspl3_w_n525_0(.douta(w_n525_0[0]),.doutb(w_n525_0[1]),.doutc(w_n525_0[2]),.din(n525));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl3 jspl3_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.doutc(w_n528_0[2]),.din(n528));
	jspl jspl_w_n528_1(.douta(w_n528_1[0]),.doutb(w_n528_1[1]),.din(w_n528_0[0]));
	jspl jspl_w_n529_0(.douta(w_n529_0[0]),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(n530));
	jspl3 jspl3_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.doutc(w_n531_0[2]),.din(n531));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl3 jspl3_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.doutc(w_n534_0[2]),.din(n534));
	jspl jspl_w_n534_1(.douta(w_n534_1[0]),.doutb(w_n534_1[1]),.din(w_n534_0[0]));
	jspl3 jspl3_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.doutc(w_n535_0[2]),.din(n535));
	jspl jspl_w_n535_1(.douta(w_n535_1[0]),.doutb(w_n535_1[1]),.din(w_n535_0[0]));
	jspl jspl_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.din(n536));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl3 jspl3_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.doutc(w_n539_0[2]),.din(n539));
	jspl jspl_w_n539_1(.douta(w_n539_1[0]),.doutb(w_n539_1[1]),.din(w_n539_0[0]));
	jspl3 jspl3_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.doutc(w_n540_0[2]),.din(n540));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n549_0(.douta(w_n549_0[0]),.doutb(w_n549_0[1]),.din(n549));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(n552));
	jspl jspl_w_n553_0(.douta(w_n553_0[0]),.doutb(w_n553_0[1]),.din(n553));
	jspl3 jspl3_w_n554_0(.douta(w_n554_0[0]),.doutb(w_n554_0[1]),.doutc(w_n554_0[2]),.din(n554));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl3 jspl3_w_n558_0(.douta(w_n558_0[0]),.doutb(w_n558_0[1]),.doutc(w_n558_0[2]),.din(n558));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl3 jspl3_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.doutc(w_n562_0[2]),.din(n562));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(n563));
	jspl3 jspl3_w_n564_0(.douta(w_n564_0[0]),.doutb(w_n564_0[1]),.doutc(w_n564_0[2]),.din(n564));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl3 jspl3_w_n565_1(.douta(w_n565_1[0]),.doutb(w_n565_1[1]),.doutc(w_n565_1[2]),.din(w_n565_0[0]));
	jspl3 jspl3_w_n565_2(.douta(w_n565_2[0]),.doutb(w_n565_2[1]),.doutc(w_n565_2[2]),.din(w_n565_0[1]));
	jspl3 jspl3_w_n565_3(.douta(w_n565_3[0]),.doutb(w_n565_3[1]),.doutc(w_n565_3[2]),.din(w_n565_0[2]));
	jspl3 jspl3_w_n565_4(.douta(w_n565_4[0]),.doutb(w_n565_4[1]),.doutc(w_n565_4[2]),.din(w_n565_1[0]));
	jspl3 jspl3_w_n565_5(.douta(w_n565_5[0]),.doutb(w_n565_5[1]),.doutc(w_n565_5[2]),.din(w_n565_1[1]));
	jspl3 jspl3_w_n565_6(.douta(w_n565_6[0]),.doutb(w_n565_6[1]),.doutc(w_n565_6[2]),.din(w_n565_1[2]));
	jspl3 jspl3_w_n565_7(.douta(w_n565_7[0]),.doutb(w_n565_7[1]),.doutc(w_n565_7[2]),.din(w_n565_2[0]));
	jspl3 jspl3_w_n565_8(.douta(w_n565_8[0]),.doutb(w_n565_8[1]),.doutc(w_n565_8[2]),.din(w_n565_2[1]));
	jspl3 jspl3_w_n565_9(.douta(w_n565_9[0]),.doutb(w_n565_9[1]),.doutc(w_n565_9[2]),.din(w_n565_2[2]));
	jspl jspl_w_n565_10(.douta(w_n565_10[0]),.doutb(w_n565_10[1]),.din(w_n565_3[0]));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n567_1(.douta(w_n567_1[0]),.doutb(w_n567_1[1]),.din(w_n567_0[0]));
	jspl3 jspl3_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.doutc(w_n568_0[2]),.din(n568));
	jspl3 jspl3_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.doutc(w_n569_0[2]),.din(n569));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl jspl_w_n572_1(.douta(w_n572_1[0]),.doutb(w_n572_1[1]),.din(w_n572_0[0]));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_n573_0[2]),.din(n573));
	jspl jspl_w_n573_1(.douta(w_n573_1[0]),.doutb(w_n573_1[1]),.din(w_n573_0[0]));
	jspl jspl_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.din(n574));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl3 jspl3_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.doutc(w_n577_0[2]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.doutc(w_n578_0[2]),.din(n578));
	jspl jspl_w_n578_1(.douta(w_n578_1[0]),.doutb(w_n578_1[1]),.din(w_n578_0[0]));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.doutc(w_n579_0[2]),.din(n579));
	jspl jspl_w_n580_0(.douta(w_n580_0[0]),.doutb(w_n580_0[1]),.din(n580));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl3 jspl3_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.doutc(w_n583_0[2]),.din(n583));
	jspl jspl_w_n583_1(.douta(w_n583_1[0]),.doutb(w_n583_1[1]),.din(w_n583_0[0]));
	jspl3 jspl3_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.doutc(w_n584_0[2]),.din(n584));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl jspl_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.din(n586));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n589_0(.douta(w_n589_0[0]),.doutb(w_n589_0[1]),.doutc(w_n589_0[2]),.din(n589));
	jspl jspl_w_n589_1(.douta(w_n589_1[0]),.doutb(w_n589_1[1]),.din(w_n589_0[0]));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(n592));
	jspl jspl_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.din(n599));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl3 jspl3_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.doutc(w_n606_0[2]),.din(n606));
	jspl3 jspl3_w_n606_1(.douta(w_n606_1[0]),.doutb(w_n606_1[1]),.doutc(w_n606_1[2]),.din(w_n606_0[0]));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.doutc(w_n608_0[2]),.din(n608));
	jspl jspl_w_n610_0(.douta(w_n610_0[0]),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.doutc(w_n615_0[2]),.din(n615));
	jspl jspl_w_n615_1(.douta(w_n615_1[0]),.doutb(w_n615_1[1]),.din(w_n615_0[0]));
	jspl jspl_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.din(n617));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.din(n620));
	jspl3 jspl3_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.doutc(w_n621_0[2]),.din(n621));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_n622_0[2]),.din(n622));
	jspl jspl_w_n622_1(.douta(w_n622_1[0]),.doutb(w_n622_1[1]),.din(w_n622_0[0]));
	jspl3 jspl3_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.doutc(w_n623_0[2]),.din(n623));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(n626));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(n628));
	jspl jspl_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.din(n629));
	jspl3 jspl3_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.doutc(w_n630_0[2]),.din(n630));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl jspl_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.din(n633));
	jspl3 jspl3_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.doutc(w_n634_0[2]),.din(n634));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(n637));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl jspl_w_n643_0(.douta(w_n643_0[0]),.doutb(w_n643_0[1]),.din(n643));
	jspl3 jspl3_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.doutc(w_n645_0[2]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(n647));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.doutc(w_n648_0[2]),.din(n648));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl3 jspl3_w_n653_0(.douta(w_n653_0[0]),.doutb(w_n653_0[1]),.doutc(w_n653_0[2]),.din(n653));
	jspl jspl_w_n653_1(.douta(w_n653_1[0]),.doutb(w_n653_1[1]),.din(w_n653_0[0]));
	jspl jspl_w_n656_0(.douta(w_n656_0[0]),.doutb(w_n656_0[1]),.din(n656));
	jspl3 jspl3_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.doutc(w_n657_0[2]),.din(n657));
	jspl jspl_w_n657_1(.douta(w_n657_1[0]),.doutb(w_n657_1[1]),.din(w_n657_0[0]));
	jspl3 jspl3_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.doutc(w_n658_0[2]),.din(n658));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_n660_0[2]),.din(n660));
	jspl jspl_w_n660_1(.douta(w_n660_1[0]),.doutb(w_n660_1[1]),.din(w_n660_0[0]));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl3 jspl3_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.doutc(w_n662_0[2]),.din(n662));
	jspl jspl_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.din(n663));
	jspl3 jspl3_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.doutc(w_n664_0[2]),.din(n664));
	jspl jspl_w_n664_1(.douta(w_n664_1[0]),.doutb(w_n664_1[1]),.din(w_n664_0[0]));
	jspl3 jspl3_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.doutc(w_n665_0[2]),.din(n665));
	jspl jspl_w_n666_0(.douta(w_n666_0[0]),.doutb(w_n666_0[1]),.din(n666));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(n667));
	jspl3 jspl3_w_n668_0(.douta(w_n668_0[0]),.doutb(w_n668_0[1]),.doutc(w_n668_0[2]),.din(n668));
	jspl3 jspl3_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.doutc(w_n669_0[2]),.din(n669));
	jspl jspl_w_n671_0(.douta(w_n671_0[0]),.doutb(w_n671_0[1]),.din(n671));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl3 jspl3_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.doutc(w_n673_0[2]),.din(n673));
	jspl3 jspl3_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.doutc(w_n674_0[2]),.din(n674));
	jspl jspl_w_n674_1(.douta(w_n674_1[0]),.doutb(w_n674_1[1]),.din(w_n674_0[0]));
	jspl3 jspl3_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.doutc(w_n675_0[2]),.din(n675));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl3 jspl3_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.doutc(w_n677_0[2]),.din(n677));
	jspl3 jspl3_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.doutc(w_n678_0[2]),.din(n678));
	jspl3 jspl3_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.doutc(w_n679_0[2]),.din(n679));
	jspl jspl_w_n679_1(.douta(w_n679_1[0]),.doutb(w_n679_1[1]),.din(w_n679_0[0]));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.din(n692));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl3 jspl3_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.doutc(w_n697_0[2]),.din(n697));
	jspl3 jspl3_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.doutc(w_n699_0[2]),.din(n699));
	jspl jspl_w_n699_1(.douta(w_n699_1[0]),.doutb(w_n699_1[1]),.din(w_n699_0[0]));
	jspl3 jspl3_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.doutc(w_n701_0[2]),.din(n701));
	jspl jspl_w_n701_1(.douta(w_n701_1[0]),.doutb(w_n701_1[1]),.din(w_n701_0[0]));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.doutc(w_n707_0[2]),.din(n707));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.din(n708));
	jspl3 jspl3_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.doutc(w_n709_0[2]),.din(n709));
	jspl jspl_w_n709_1(.douta(w_n709_1[0]),.doutb(w_n709_1[1]),.din(w_n709_0[0]));
	jspl jspl_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.din(n712));
	jspl3 jspl3_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.doutc(w_n713_0[2]),.din(n713));
	jspl jspl_w_n713_1(.douta(w_n713_1[0]),.doutb(w_n713_1[1]),.din(w_n713_0[0]));
	jspl jspl_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.din(n714));
	jspl3 jspl3_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.doutc(w_n715_0[2]),.din(n715));
	jspl3 jspl3_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.doutc(w_n716_0[2]),.din(n716));
	jspl jspl_w_n716_1(.douta(w_n716_1[0]),.doutb(w_n716_1[1]),.din(w_n716_0[0]));
	jspl3 jspl3_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.doutc(w_n720_0[2]),.din(w_dff_B_fBSeNbDi3_3));
	jspl jspl_w_n720_1(.douta(w_n720_1[0]),.doutb(w_n720_1[1]),.din(w_n720_0[0]));
	jspl3 jspl3_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.doutc(w_n723_0[2]),.din(n723));
	jspl3 jspl3_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.doutc(w_n727_0[2]),.din(n727));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n730_0(.douta(w_n730_0[0]),.doutb(w_n730_0[1]),.doutc(w_n730_0[2]),.din(n730));
	jspl3 jspl3_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.doutc(w_n734_0[2]),.din(n734));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.din(n735));
	jspl3 jspl3_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_n744_0[2]),.din(n744));
	jspl3 jspl3_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.doutc(w_n748_0[2]),.din(n748));
	jspl jspl_w_n751_0(.douta(w_n751_0[0]),.doutb(w_n751_0[1]),.din(n751));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl3 jspl3_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.doutc(w_n754_0[2]),.din(n754));
	jspl3 jspl3_w_n758_0(.douta(w_n758_0[0]),.doutb(w_n758_0[1]),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(n764));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl3 jspl3_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.doutc(w_n784_0[2]),.din(n784));
	jspl3 jspl3_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.doutc(w_n787_0[2]),.din(n787));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.doutc(w_n790_0[2]),.din(n790));
	jspl jspl_w_n790_1(.douta(w_n790_1[0]),.doutb(w_n790_1[1]),.din(w_n790_0[0]));
	jspl3 jspl3_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.doutc(w_n793_0[2]),.din(n793));
	jspl jspl_w_n793_1(.douta(w_n793_1[0]),.doutb(w_n793_1[1]),.din(w_n793_0[0]));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl jspl_w_n797_1(.douta(w_n797_1[0]),.doutb(w_n797_1[1]),.din(w_n797_0[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl jspl_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.din(w_n801_0[0]));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl3 jspl3_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.doutc(w_n804_0[2]),.din(n804));
	jspl3 jspl3_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.doutc(w_n807_0[2]),.din(n807));
	jspl3 jspl3_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.doutc(w_n810_0[2]),.din(n810));
	jspl3 jspl3_w_n812_0(.douta(w_n812_0[0]),.doutb(w_n812_0[1]),.doutc(w_n812_0[2]),.din(n812));
	jspl3 jspl3_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.doutc(w_n816_0[2]),.din(n816));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(n817));
	jspl3 jspl3_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.doutc(w_n819_0[2]),.din(n819));
	jspl3 jspl3_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.doutc(w_n823_0[2]),.din(n823));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl3 jspl3_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.doutc(w_n827_0[2]),.din(n827));
	jspl3 jspl3_w_n831_0(.douta(w_n831_0[0]),.doutb(w_n831_0[1]),.doutc(w_n831_0[2]),.din(n831));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n838_0(.douta(w_n838_0[0]),.doutb(w_n838_0[1]),.din(n838));
	jspl3 jspl3_w_n843_0(.douta(w_n843_0[0]),.doutb(w_n843_0[1]),.doutc(w_n843_0[2]),.din(n843));
	jspl3 jspl3_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.doutc(w_n847_0[2]),.din(n847));
	jspl jspl_w_n848_0(.douta(w_n848_0[0]),.doutb(w_n848_0[1]),.din(n848));
	jspl3 jspl3_w_n851_0(.douta(w_n851_0[0]),.doutb(w_n851_0[1]),.doutc(w_n851_0[2]),.din(n851));
	jspl3 jspl3_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.doutc(w_n855_0[2]),.din(n855));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl3 jspl3_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.doutc(w_n858_0[2]),.din(n858));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.din(n865));
	jspl3 jspl3_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.doutc(w_n869_0[2]),.din(n869));
	jspl3 jspl3_w_n873_0(.douta(w_n873_0[0]),.doutb(w_n873_0[1]),.doutc(w_n873_0[2]),.din(n873));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(n874));
	jspl3 jspl3_w_n878_0(.douta(w_n878_0[0]),.doutb(w_n878_0[1]),.doutc(w_n878_0[2]),.din(n878));
	jspl3 jspl3_w_n882_0(.douta(w_n882_0[0]),.doutb(w_n882_0[1]),.doutc(w_n882_0[2]),.din(n882));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.din(n887));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl3 jspl3_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.doutc(w_n891_0[2]),.din(n891));
	jspl jspl_w_n891_1(.douta(w_n891_1[0]),.doutb(w_n891_1[1]),.din(w_n891_0[0]));
	jspl3 jspl3_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.doutc(w_n895_0[2]),.din(n895));
	jspl jspl_w_n895_1(.douta(w_n895_1[0]),.doutb(w_n895_1[1]),.din(w_n895_0[0]));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(n896));
	jspl3 jspl3_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.doutc(w_n899_0[2]),.din(n899));
	jspl3 jspl3_w_n902_0(.douta(w_n902_0[0]),.doutb(w_n902_0[1]),.doutc(w_n902_0[2]),.din(n902));
	jspl3 jspl3_w_n905_0(.douta(w_n905_0[0]),.doutb(w_n905_0[1]),.doutc(w_n905_0[2]),.din(n905));
	jspl3 jspl3_w_n908_0(.douta(w_n908_0[0]),.doutb(w_n908_0[1]),.doutc(w_n908_0[2]),.din(n908));
	jspl3 jspl3_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.doutc(w_n912_0[2]),.din(n912));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(n913));
	jspl3 jspl3_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.doutc(w_n916_0[2]),.din(n916));
	jspl3 jspl3_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.doutc(w_n920_0[2]),.din(n920));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(n923));
	jspl3 jspl3_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.doutc(w_n927_0[2]),.din(n927));
	jspl3 jspl3_w_n931_0(.douta(w_n931_0[0]),.doutb(w_n931_0[1]),.doutc(w_n931_0[2]),.din(n931));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n939_0(.douta(w_n939_0[0]),.doutb(w_n939_0[1]),.din(n939));
	jspl3 jspl3_w_n945_0(.douta(w_n945_0[0]),.doutb(w_n945_0[1]),.doutc(w_n945_0[2]),.din(n945));
	jspl jspl_w_n945_1(.douta(w_n945_1[0]),.doutb(w_n945_1[1]),.din(w_n945_0[0]));
	jspl3 jspl3_w_n948_0(.douta(w_n948_0[0]),.doutb(w_n948_0[1]),.doutc(w_n948_0[2]),.din(n948));
	jspl jspl_w_n948_1(.douta(w_n948_1[0]),.doutb(w_n948_1[1]),.din(w_n948_0[0]));
	jspl jspl_w_n950_0(.douta(w_n950_0[0]),.doutb(w_n950_0[1]),.din(n950));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.doutc(w_n988_0[2]),.din(n988));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl3 jspl3_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.doutc(w_n995_0[2]),.din(n995));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.doutc(w_n999_0[2]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.din(n1008));
	jspl3 jspl3_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.doutc(w_n1009_0[2]),.din(n1009));
	jspl jspl_w_n1009_1(.douta(w_n1009_1[0]),.doutb(w_n1009_1[1]),.din(w_n1009_0[0]));
	jspl3 jspl3_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.doutc(w_n1013_0[2]),.din(n1013));
	jspl jspl_w_n1013_1(.douta(w_n1013_1[0]),.doutb(w_n1013_1[1]),.din(w_n1013_0[0]));
	jspl jspl_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.din(n1014));
	jspl jspl_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.din(n1015));
	jspl3 jspl3_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.doutc(w_n1016_0[2]),.din(n1016));
	jspl3 jspl3_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.doutc(w_n1019_0[2]),.din(n1019));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(n1044));
	jspl3 jspl3_w_n1061_0(.douta(w_n1061_0[0]),.doutb(w_n1061_0[1]),.doutc(w_n1061_0[2]),.din(n1061));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.din(n1062));
	jspl3 jspl3_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.doutc(w_n1066_0[2]),.din(n1066));
	jspl jspl_w_n1068_0(.douta(w_n1068_0[0]),.doutb(w_n1068_0[1]),.din(n1068));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(n1069));
	jspl3 jspl3_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.doutc(w_n1073_0[2]),.din(n1073));
	jspl jspl_w_n1075_0(.douta(w_n1075_0[0]),.doutb(w_n1075_0[1]),.din(n1075));
	jspl jspl_w_n1076_0(.douta(w_n1076_0[0]),.doutb(w_n1076_0[1]),.din(n1076));
	jspl3 jspl3_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.doutc(w_n1077_0[2]),.din(n1077));
	jspl3 jspl3_w_n1081_0(.douta(w_n1081_0[0]),.doutb(w_n1081_0[1]),.doutc(w_n1081_0[2]),.din(n1081));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl3 jspl3_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.doutc(w_n1086_0[2]),.din(n1086));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.din(n1095));
	jspl3 jspl3_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.doutc(w_n1096_0[2]),.din(n1096));
	jspl3 jspl3_w_n1100_0(.douta(w_n1100_0[0]),.doutb(w_n1100_0[1]),.doutc(w_n1100_0[2]),.din(n1100));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1104_0(.douta(w_n1104_0[0]),.doutb(w_n1104_0[1]),.din(n1104));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.din(n1105));
	jspl jspl_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.din(n1116));
	jspl3 jspl3_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.doutc(w_n1122_0[2]),.din(n1122));
	jspl3 jspl3_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.doutc(w_n1125_0[2]),.din(w_dff_B_9MDYm1pu5_3));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(n1127));
	jspl3 jspl3_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.doutc(w_n1128_0[2]),.din(n1128));
	jspl jspl_w_n1128_1(.douta(w_n1128_1[0]),.doutb(w_n1128_1[1]),.din(w_n1128_0[0]));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1136_0(.douta(w_n1136_0[0]),.doutb(w_n1136_0[1]),.din(n1136));
	jspl jspl_w_n1142_0(.douta(w_n1142_0[0]),.doutb(w_n1142_0[1]),.din(n1142));
	jspl3 jspl3_w_n1148_0(.douta(w_n1148_0[0]),.doutb(w_n1148_0[1]),.doutc(w_n1148_0[2]),.din(n1148));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(n1156));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(n1173));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(n1283));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl3 jspl3_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.doutc(w_n1359_0[2]),.din(n1359));
	jspl3 jspl3_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.doutc(w_n1360_0[2]),.din(n1360));
	jspl jspl_w_n1360_1(.douta(w_n1360_1[0]),.doutb(w_n1360_1[1]),.din(w_n1360_0[0]));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1362_0(.douta(w_n1362_0[0]),.doutb(w_n1362_0[1]),.din(n1362));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(n1376));
	jspl3 jspl3_w_n1380_0(.douta(w_n1380_0[0]),.doutb(w_n1380_0[1]),.doutc(w_n1380_0[2]),.din(n1380));
	jspl jspl_w_n1380_1(.douta(w_n1380_1[0]),.doutb(w_n1380_1[1]),.din(w_n1380_0[0]));
	jspl3 jspl3_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.doutc(w_n1383_0[2]),.din(n1383));
	jspl3 jspl3_w_n1383_1(.douta(w_n1383_1[0]),.doutb(w_n1383_1[1]),.doutc(w_n1383_1[2]),.din(w_n1383_0[0]));
	jspl3 jspl3_w_n1385_0(.douta(w_n1385_0[0]),.doutb(w_n1385_0[1]),.doutc(w_n1385_0[2]),.din(n1385));
	jspl jspl_w_n1385_1(.douta(w_n1385_1[0]),.doutb(w_n1385_1[1]),.din(w_n1385_0[0]));
	jspl3 jspl3_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.doutc(w_n1389_0[2]),.din(n1389));
	jspl jspl_w_n1389_1(.douta(w_n1389_1[0]),.doutb(w_n1389_1[1]),.din(w_n1389_0[0]));
	jspl3 jspl3_w_n1392_0(.douta(w_n1392_0[0]),.doutb(w_n1392_0[1]),.doutc(w_n1392_0[2]),.din(n1392));
	jspl jspl_w_n1392_1(.douta(w_n1392_1[0]),.doutb(w_n1392_1[1]),.din(w_n1392_0[0]));
	jspl jspl_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_n1401_0[1]),.din(n1401));
	jspl jspl_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_n1402_0[1]),.din(n1402));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_n1404_0[1]),.din(n1404));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl jspl_w_n1406_0(.douta(w_n1406_0[0]),.doutb(w_n1406_0[1]),.din(n1406));
	jspl jspl_w_n1414_0(.douta(w_n1414_0[0]),.doutb(w_n1414_0[1]),.din(n1414));
	jspl3 jspl3_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.doutc(w_n1420_0[2]),.din(n1420));
	jspl jspl_w_n1421_0(.douta(w_n1421_0[0]),.doutb(w_n1421_0[1]),.din(n1421));
	jspl jspl_w_n1422_0(.douta(w_n1422_0[0]),.doutb(w_n1422_0[1]),.din(n1422));
	jspl jspl_w_n1424_0(.douta(w_n1424_0[0]),.doutb(w_n1424_0[1]),.din(n1424));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl3 jspl3_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.doutc(w_n1444_0[2]),.din(n1444));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(n1454));
	jspl3 jspl3_w_n1463_0(.douta(w_n1463_0[0]),.doutb(w_n1463_0[1]),.doutc(w_n1463_0[2]),.din(n1463));
	jspl jspl_w_n1464_0(.douta(w_n1464_0[0]),.doutb(w_n1464_0[1]),.din(n1464));
	jspl jspl_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.din(n1465));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_n1468_0[1]),.din(n1468));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1470_0(.douta(w_n1470_0[0]),.doutb(w_n1470_0[1]),.din(n1470));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(n1471));
	jspl jspl_w_n1472_0(.douta(w_n1472_0[0]),.doutb(w_n1472_0[1]),.din(n1472));
	jspl jspl_w_n1473_0(.douta(w_n1473_0[0]),.doutb(w_n1473_0[1]),.din(n1473));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(n1479));
	jspl jspl_w_n1482_0(.douta(w_n1482_0[0]),.doutb(w_n1482_0[1]),.din(n1482));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(n1486));
	jspl3 jspl3_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.doutc(w_n1494_0[2]),.din(n1494));
	jspl jspl_w_n1501_0(.douta(w_n1501_0[0]),.doutb(w_n1501_0[1]),.din(n1501));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.din(n1520));
	jspl jspl_w_n1536_0(.douta(w_n1536_0[0]),.doutb(w_n1536_0[1]),.din(n1536));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(n1571));
	jspl jspl_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.din(n1611));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl jspl_w_n1642_0(.douta(w_n1642_0[0]),.doutb(w_n1642_0[1]),.din(n1642));
	jspl jspl_w_n1644_0(.douta(w_n1644_0[0]),.doutb(w_n1644_0[1]),.din(n1644));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(n1651));
	jspl jspl_w_n1654_0(.douta(w_n1654_0[0]),.doutb(w_n1654_0[1]),.din(n1654));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1667_0(.douta(w_n1667_0[0]),.doutb(w_n1667_0[1]),.din(n1667));
	jspl jspl_w_n1670_0(.douta(w_n1670_0[0]),.doutb(w_n1670_0[1]),.din(n1670));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(n1672));
	jspl jspl_w_n1675_0(.douta(w_n1675_0[0]),.doutb(w_n1675_0[1]),.din(n1675));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_n1687_0[1]),.din(n1687));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(n1689));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(n1699));
	jdff dff_A_9QO5kMsf6_0(.dout(w_G5_1[0]),.din(w_dff_A_9QO5kMsf6_0),.clk(gclk));
	jdff dff_A_7yeiBPBK4_0(.dout(w_dff_A_9QO5kMsf6_0),.din(w_dff_A_7yeiBPBK4_0),.clk(gclk));
	jdff dff_A_UczSuiSW2_1(.dout(w_G5_1[1]),.din(w_dff_A_UczSuiSW2_1),.clk(gclk));
	jdff dff_A_J3enjoPb9_1(.dout(w_G5_0[1]),.din(w_dff_A_J3enjoPb9_1),.clk(gclk));
	jdff dff_A_nZ0M8cl96_1(.dout(w_dff_A_J3enjoPb9_1),.din(w_dff_A_nZ0M8cl96_1),.clk(gclk));
	jdff dff_A_trt7Zdp61_2(.dout(w_G5_0[2]),.din(w_dff_A_trt7Zdp61_2),.clk(gclk));
	jdff dff_B_FzU78smc9_3(.din(n1125),.dout(w_dff_B_FzU78smc9_3),.clk(gclk));
	jdff dff_B_QKk2GhSn2_3(.din(w_dff_B_FzU78smc9_3),.dout(w_dff_B_QKk2GhSn2_3),.clk(gclk));
	jdff dff_B_98XYDJw71_3(.din(w_dff_B_QKk2GhSn2_3),.dout(w_dff_B_98XYDJw71_3),.clk(gclk));
	jdff dff_B_1hi48cLb9_3(.din(w_dff_B_98XYDJw71_3),.dout(w_dff_B_1hi48cLb9_3),.clk(gclk));
	jdff dff_B_0O7tdvpT7_3(.din(w_dff_B_1hi48cLb9_3),.dout(w_dff_B_0O7tdvpT7_3),.clk(gclk));
	jdff dff_B_RlafvuDv0_3(.din(w_dff_B_0O7tdvpT7_3),.dout(w_dff_B_RlafvuDv0_3),.clk(gclk));
	jdff dff_B_c7nUrlS48_3(.din(w_dff_B_RlafvuDv0_3),.dout(w_dff_B_c7nUrlS48_3),.clk(gclk));
	jdff dff_B_qVGDMjuk5_3(.din(w_dff_B_c7nUrlS48_3),.dout(w_dff_B_qVGDMjuk5_3),.clk(gclk));
	jdff dff_B_l8esVTko5_3(.din(w_dff_B_qVGDMjuk5_3),.dout(w_dff_B_l8esVTko5_3),.clk(gclk));
	jdff dff_B_gIskj6br3_3(.din(w_dff_B_l8esVTko5_3),.dout(w_dff_B_gIskj6br3_3),.clk(gclk));
	jdff dff_B_HYZgzBaJ0_3(.din(w_dff_B_gIskj6br3_3),.dout(w_dff_B_HYZgzBaJ0_3),.clk(gclk));
	jdff dff_B_Jyrb7Aq96_3(.din(w_dff_B_HYZgzBaJ0_3),.dout(w_dff_B_Jyrb7Aq96_3),.clk(gclk));
	jdff dff_B_7CCFwbtG6_3(.din(w_dff_B_Jyrb7Aq96_3),.dout(w_dff_B_7CCFwbtG6_3),.clk(gclk));
	jdff dff_B_wwddzhuJ8_3(.din(w_dff_B_7CCFwbtG6_3),.dout(w_dff_B_wwddzhuJ8_3),.clk(gclk));
	jdff dff_B_2h7M6AcW9_3(.din(w_dff_B_wwddzhuJ8_3),.dout(w_dff_B_2h7M6AcW9_3),.clk(gclk));
	jdff dff_B_9MDYm1pu5_3(.din(w_dff_B_2h7M6AcW9_3),.dout(w_dff_B_9MDYm1pu5_3),.clk(gclk));
	jdff dff_B_GEaJHj6j2_0(.din(n1441),.dout(w_dff_B_GEaJHj6j2_0),.clk(gclk));
	jdff dff_B_beIsjM3H9_0(.din(n1440),.dout(w_dff_B_beIsjM3H9_0),.clk(gclk));
	jdff dff_B_jYpCtpT52_0(.din(w_dff_B_beIsjM3H9_0),.dout(w_dff_B_jYpCtpT52_0),.clk(gclk));
	jdff dff_B_3PvZ7pln0_0(.din(w_dff_B_jYpCtpT52_0),.dout(w_dff_B_3PvZ7pln0_0),.clk(gclk));
	jdff dff_B_NzkL4KCy0_0(.din(w_dff_B_3PvZ7pln0_0),.dout(w_dff_B_NzkL4KCy0_0),.clk(gclk));
	jdff dff_B_wqq56lm13_0(.din(w_dff_B_NzkL4KCy0_0),.dout(w_dff_B_wqq56lm13_0),.clk(gclk));
	jdff dff_B_7o9MhInf4_0(.din(w_dff_B_wqq56lm13_0),.dout(w_dff_B_7o9MhInf4_0),.clk(gclk));
	jdff dff_A_gWIsP7hv9_0(.dout(w_G414_0),.din(w_dff_A_gWIsP7hv9_0),.clk(gclk));
	jdff dff_A_6ENtODDw6_0(.dout(w_dff_A_gWIsP7hv9_0),.din(w_dff_A_6ENtODDw6_0),.clk(gclk));
	jdff dff_A_qE6J2TTm7_0(.dout(w_dff_A_6ENtODDw6_0),.din(w_dff_A_qE6J2TTm7_0),.clk(gclk));
	jdff dff_B_dUmJ2nLu5_3(.din(n720),.dout(w_dff_B_dUmJ2nLu5_3),.clk(gclk));
	jdff dff_B_zCbOuQPA0_3(.din(w_dff_B_dUmJ2nLu5_3),.dout(w_dff_B_zCbOuQPA0_3),.clk(gclk));
	jdff dff_B_ZcdM3jqe8_3(.din(w_dff_B_zCbOuQPA0_3),.dout(w_dff_B_ZcdM3jqe8_3),.clk(gclk));
	jdff dff_B_FVvdv52x2_3(.din(w_dff_B_ZcdM3jqe8_3),.dout(w_dff_B_FVvdv52x2_3),.clk(gclk));
	jdff dff_B_MLds6pbi2_3(.din(w_dff_B_FVvdv52x2_3),.dout(w_dff_B_MLds6pbi2_3),.clk(gclk));
	jdff dff_B_k3HNFrRD1_3(.din(w_dff_B_MLds6pbi2_3),.dout(w_dff_B_k3HNFrRD1_3),.clk(gclk));
	jdff dff_B_QLKWXMm39_3(.din(w_dff_B_k3HNFrRD1_3),.dout(w_dff_B_QLKWXMm39_3),.clk(gclk));
	jdff dff_B_N6HqhR0y8_3(.din(w_dff_B_QLKWXMm39_3),.dout(w_dff_B_N6HqhR0y8_3),.clk(gclk));
	jdff dff_B_gOHBfbdE9_3(.din(w_dff_B_N6HqhR0y8_3),.dout(w_dff_B_gOHBfbdE9_3),.clk(gclk));
	jdff dff_B_yhVRwWBm1_3(.din(w_dff_B_gOHBfbdE9_3),.dout(w_dff_B_yhVRwWBm1_3),.clk(gclk));
	jdff dff_B_cxTFjToG5_3(.din(w_dff_B_yhVRwWBm1_3),.dout(w_dff_B_cxTFjToG5_3),.clk(gclk));
	jdff dff_B_qS8OzpVe0_3(.din(w_dff_B_cxTFjToG5_3),.dout(w_dff_B_qS8OzpVe0_3),.clk(gclk));
	jdff dff_B_PoMEaLyb3_3(.din(w_dff_B_qS8OzpVe0_3),.dout(w_dff_B_PoMEaLyb3_3),.clk(gclk));
	jdff dff_B_KNTreujU3_3(.din(w_dff_B_PoMEaLyb3_3),.dout(w_dff_B_KNTreujU3_3),.clk(gclk));
	jdff dff_B_fNpvSgHX4_3(.din(w_dff_B_KNTreujU3_3),.dout(w_dff_B_fNpvSgHX4_3),.clk(gclk));
	jdff dff_B_p7Uf4fmW9_3(.din(w_dff_B_fNpvSgHX4_3),.dout(w_dff_B_p7Uf4fmW9_3),.clk(gclk));
	jdff dff_B_ZlWdhG8u9_3(.din(w_dff_B_p7Uf4fmW9_3),.dout(w_dff_B_ZlWdhG8u9_3),.clk(gclk));
	jdff dff_B_WmOCm0RJ3_3(.din(w_dff_B_ZlWdhG8u9_3),.dout(w_dff_B_WmOCm0RJ3_3),.clk(gclk));
	jdff dff_B_805vkh0G7_3(.din(w_dff_B_WmOCm0RJ3_3),.dout(w_dff_B_805vkh0G7_3),.clk(gclk));
	jdff dff_B_t54pZ6mO1_3(.din(w_dff_B_805vkh0G7_3),.dout(w_dff_B_t54pZ6mO1_3),.clk(gclk));
	jdff dff_B_fBSeNbDi3_3(.din(w_dff_B_t54pZ6mO1_3),.dout(w_dff_B_fBSeNbDi3_3),.clk(gclk));
	jdff dff_B_vpIy1vDB9_1(.din(n1451),.dout(w_dff_B_vpIy1vDB9_1),.clk(gclk));
	jdff dff_B_1EiMZeuy7_1(.din(w_dff_B_vpIy1vDB9_1),.dout(w_dff_B_1EiMZeuy7_1),.clk(gclk));
	jdff dff_B_OCAc2VMT7_1(.din(w_dff_B_1EiMZeuy7_1),.dout(w_dff_B_OCAc2VMT7_1),.clk(gclk));
	jdff dff_B_jKZGV9nb8_1(.din(w_dff_B_OCAc2VMT7_1),.dout(w_dff_B_jKZGV9nb8_1),.clk(gclk));
	jdff dff_B_D5NeVKLt5_1(.din(w_dff_B_jKZGV9nb8_1),.dout(w_dff_B_D5NeVKLt5_1),.clk(gclk));
	jdff dff_B_DbWs0oaN0_1(.din(w_dff_B_D5NeVKLt5_1),.dout(w_dff_B_DbWs0oaN0_1),.clk(gclk));
	jdff dff_B_IqtCQLiX5_1(.din(w_dff_B_DbWs0oaN0_1),.dout(w_dff_B_IqtCQLiX5_1),.clk(gclk));
	jdff dff_B_IpQODK7f5_1(.din(w_dff_B_IqtCQLiX5_1),.dout(w_dff_B_IpQODK7f5_1),.clk(gclk));
	jdff dff_B_xjehSzm19_1(.din(w_dff_B_IpQODK7f5_1),.dout(w_dff_B_xjehSzm19_1),.clk(gclk));
	jdff dff_B_GO6NziZ45_1(.din(w_dff_B_xjehSzm19_1),.dout(w_dff_B_GO6NziZ45_1),.clk(gclk));
	jdff dff_B_6CedrUXU4_1(.din(w_dff_B_GO6NziZ45_1),.dout(w_dff_B_6CedrUXU4_1),.clk(gclk));
	jdff dff_B_HZR9lwyG3_1(.din(w_dff_B_6CedrUXU4_1),.dout(w_dff_B_HZR9lwyG3_1),.clk(gclk));
	jdff dff_B_PqrPMV0z5_1(.din(w_dff_B_HZR9lwyG3_1),.dout(w_dff_B_PqrPMV0z5_1),.clk(gclk));
	jdff dff_B_1j8yn1Co1_1(.din(w_dff_B_PqrPMV0z5_1),.dout(w_dff_B_1j8yn1Co1_1),.clk(gclk));
	jdff dff_B_fbaVvFO18_1(.din(w_dff_B_1j8yn1Co1_1),.dout(w_dff_B_fbaVvFO18_1),.clk(gclk));
	jdff dff_B_jokLNW1J8_1(.din(n1500),.dout(w_dff_B_jokLNW1J8_1),.clk(gclk));
	jdff dff_B_8iTWyAfu7_1(.din(w_dff_B_jokLNW1J8_1),.dout(w_dff_B_8iTWyAfu7_1),.clk(gclk));
	jdff dff_B_VEBovauy4_1(.din(w_dff_B_8iTWyAfu7_1),.dout(w_dff_B_VEBovauy4_1),.clk(gclk));
	jdff dff_B_NgxFGKZy6_1(.din(w_dff_B_VEBovauy4_1),.dout(w_dff_B_NgxFGKZy6_1),.clk(gclk));
	jdff dff_B_yoJOtEfA0_1(.din(w_dff_B_NgxFGKZy6_1),.dout(w_dff_B_yoJOtEfA0_1),.clk(gclk));
	jdff dff_B_sa2I5if72_1(.din(w_dff_B_yoJOtEfA0_1),.dout(w_dff_B_sa2I5if72_1),.clk(gclk));
	jdff dff_B_hWUmrSTw6_1(.din(w_dff_B_sa2I5if72_1),.dout(w_dff_B_hWUmrSTw6_1),.clk(gclk));
	jdff dff_B_k1hjEaZw6_1(.din(w_dff_B_hWUmrSTw6_1),.dout(w_dff_B_k1hjEaZw6_1),.clk(gclk));
	jdff dff_B_kxsOkfov5_1(.din(w_dff_B_k1hjEaZw6_1),.dout(w_dff_B_kxsOkfov5_1),.clk(gclk));
	jdff dff_B_YVoRaUVm1_1(.din(w_dff_B_kxsOkfov5_1),.dout(w_dff_B_YVoRaUVm1_1),.clk(gclk));
	jdff dff_B_unL2ikBW9_1(.din(w_dff_B_YVoRaUVm1_1),.dout(w_dff_B_unL2ikBW9_1),.clk(gclk));
	jdff dff_B_Ul7f0PSX0_1(.din(w_dff_B_unL2ikBW9_1),.dout(w_dff_B_Ul7f0PSX0_1),.clk(gclk));
	jdff dff_B_o3urkvCr2_1(.din(w_dff_B_Ul7f0PSX0_1),.dout(w_dff_B_o3urkvCr2_1),.clk(gclk));
	jdff dff_B_ZtOmaFTA5_1(.din(w_dff_B_o3urkvCr2_1),.dout(w_dff_B_ZtOmaFTA5_1),.clk(gclk));
	jdff dff_B_ZBSCXzLP5_1(.din(w_dff_B_ZtOmaFTA5_1),.dout(w_dff_B_ZBSCXzLP5_1),.clk(gclk));
	jdff dff_B_IcqrIkq40_0(.din(n1584),.dout(w_dff_B_IcqrIkq40_0),.clk(gclk));
	jdff dff_B_Pcx1cnVY3_0(.din(w_dff_B_IcqrIkq40_0),.dout(w_dff_B_Pcx1cnVY3_0),.clk(gclk));
	jdff dff_B_mRB84Aq46_0(.din(w_dff_B_Pcx1cnVY3_0),.dout(w_dff_B_mRB84Aq46_0),.clk(gclk));
	jdff dff_B_FjQeWa9J1_1(.din(n1587),.dout(w_dff_B_FjQeWa9J1_1),.clk(gclk));
	jdff dff_B_4nntlRnQ0_1(.din(w_dff_B_FjQeWa9J1_1),.dout(w_dff_B_4nntlRnQ0_1),.clk(gclk));
	jdff dff_B_uf5Db5j67_1(.din(w_dff_B_4nntlRnQ0_1),.dout(w_dff_B_uf5Db5j67_1),.clk(gclk));
	jdff dff_B_wpLSqmpN9_1(.din(w_dff_B_uf5Db5j67_1),.dout(w_dff_B_wpLSqmpN9_1),.clk(gclk));
	jdff dff_B_3YOAXYRg6_1(.din(w_dff_B_wpLSqmpN9_1),.dout(w_dff_B_3YOAXYRg6_1),.clk(gclk));
	jdff dff_B_NpqUElue4_1(.din(w_dff_B_3YOAXYRg6_1),.dout(w_dff_B_NpqUElue4_1),.clk(gclk));
	jdff dff_B_aMRKJmGW8_1(.din(w_dff_B_NpqUElue4_1),.dout(w_dff_B_aMRKJmGW8_1),.clk(gclk));
	jdff dff_B_4bomZnzS5_1(.din(w_dff_B_aMRKJmGW8_1),.dout(w_dff_B_4bomZnzS5_1),.clk(gclk));
	jdff dff_B_9W3GlZnr3_1(.din(w_dff_B_4bomZnzS5_1),.dout(w_dff_B_9W3GlZnr3_1),.clk(gclk));
	jdff dff_B_bIyzspRH8_1(.din(w_dff_B_9W3GlZnr3_1),.dout(w_dff_B_bIyzspRH8_1),.clk(gclk));
	jdff dff_B_1suRTZFd4_1(.din(w_dff_B_bIyzspRH8_1),.dout(w_dff_B_1suRTZFd4_1),.clk(gclk));
	jdff dff_B_ixTSlmXd3_1(.din(w_dff_B_1suRTZFd4_1),.dout(w_dff_B_ixTSlmXd3_1),.clk(gclk));
	jdff dff_B_YisDDqVG1_1(.din(n1637),.dout(w_dff_B_YisDDqVG1_1),.clk(gclk));
	jdff dff_B_BfcfbpoJ1_1(.din(w_dff_B_YisDDqVG1_1),.dout(w_dff_B_BfcfbpoJ1_1),.clk(gclk));
	jdff dff_B_hedONhuP5_1(.din(w_dff_B_BfcfbpoJ1_1),.dout(w_dff_B_hedONhuP5_1),.clk(gclk));
	jdff dff_B_bEfWGry60_1(.din(w_dff_B_hedONhuP5_1),.dout(w_dff_B_bEfWGry60_1),.clk(gclk));
	jdff dff_B_y7E0SZLh8_1(.din(w_dff_B_bEfWGry60_1),.dout(w_dff_B_y7E0SZLh8_1),.clk(gclk));
	jdff dff_B_DFsZgEkb6_1(.din(w_dff_B_y7E0SZLh8_1),.dout(w_dff_B_DFsZgEkb6_1),.clk(gclk));
	jdff dff_B_r68osuAM6_1(.din(w_dff_B_DFsZgEkb6_1),.dout(w_dff_B_r68osuAM6_1),.clk(gclk));
	jdff dff_B_PeBK9cnt2_1(.din(w_dff_B_r68osuAM6_1),.dout(w_dff_B_PeBK9cnt2_1),.clk(gclk));
	jdff dff_B_8PZoI8Si5_1(.din(w_dff_B_PeBK9cnt2_1),.dout(w_dff_B_8PZoI8Si5_1),.clk(gclk));
	jdff dff_B_sWOF15J72_1(.din(w_dff_B_8PZoI8Si5_1),.dout(w_dff_B_sWOF15J72_1),.clk(gclk));
	jdff dff_B_OCC3loJT5_1(.din(w_dff_B_sWOF15J72_1),.dout(w_dff_B_OCC3loJT5_1),.clk(gclk));
	jdff dff_B_UuV8fNvE1_1(.din(w_dff_B_OCC3loJT5_1),.dout(w_dff_B_UuV8fNvE1_1),.clk(gclk));
	jdff dff_B_v5I4KI7d8_1(.din(w_dff_B_UuV8fNvE1_1),.dout(w_dff_B_v5I4KI7d8_1),.clk(gclk));
	jdff dff_B_vrjz5V6r5_1(.din(w_dff_B_v5I4KI7d8_1),.dout(w_dff_B_vrjz5V6r5_1),.clk(gclk));
	jdff dff_B_XHnAdNvx9_1(.din(w_dff_B_vrjz5V6r5_1),.dout(w_dff_B_XHnAdNvx9_1),.clk(gclk));
	jdff dff_A_6sApNmgt4_1(.dout(w_dff_A_9ke25cNh8_0),.din(w_dff_A_6sApNmgt4_1),.clk(gclk));
	jdff dff_A_9ke25cNh8_0(.dout(w_dff_A_LZ0JsTsi0_0),.din(w_dff_A_9ke25cNh8_0),.clk(gclk));
	jdff dff_A_LZ0JsTsi0_0(.dout(w_dff_A_2UCs1x1D6_0),.din(w_dff_A_LZ0JsTsi0_0),.clk(gclk));
	jdff dff_A_2UCs1x1D6_0(.dout(w_dff_A_MC0n00H68_0),.din(w_dff_A_2UCs1x1D6_0),.clk(gclk));
	jdff dff_A_MC0n00H68_0(.dout(w_dff_A_es7rLjWZ1_0),.din(w_dff_A_MC0n00H68_0),.clk(gclk));
	jdff dff_A_es7rLjWZ1_0(.dout(w_dff_A_AXC1wYxF0_0),.din(w_dff_A_es7rLjWZ1_0),.clk(gclk));
	jdff dff_A_AXC1wYxF0_0(.dout(w_dff_A_3tN9rxVx2_0),.din(w_dff_A_AXC1wYxF0_0),.clk(gclk));
	jdff dff_A_3tN9rxVx2_0(.dout(w_dff_A_bR1Dca1U6_0),.din(w_dff_A_3tN9rxVx2_0),.clk(gclk));
	jdff dff_A_bR1Dca1U6_0(.dout(w_dff_A_yFlqPns54_0),.din(w_dff_A_bR1Dca1U6_0),.clk(gclk));
	jdff dff_A_yFlqPns54_0(.dout(w_dff_A_UWLrWuEJ8_0),.din(w_dff_A_yFlqPns54_0),.clk(gclk));
	jdff dff_A_UWLrWuEJ8_0(.dout(w_dff_A_pt1XiaWX8_0),.din(w_dff_A_UWLrWuEJ8_0),.clk(gclk));
	jdff dff_A_pt1XiaWX8_0(.dout(w_dff_A_mm5g4OxK0_0),.din(w_dff_A_pt1XiaWX8_0),.clk(gclk));
	jdff dff_A_mm5g4OxK0_0(.dout(w_dff_A_mlLZNHuO4_0),.din(w_dff_A_mm5g4OxK0_0),.clk(gclk));
	jdff dff_A_mlLZNHuO4_0(.dout(w_dff_A_qrcZCWMn1_0),.din(w_dff_A_mlLZNHuO4_0),.clk(gclk));
	jdff dff_A_qrcZCWMn1_0(.dout(w_dff_A_2BzIJhw14_0),.din(w_dff_A_qrcZCWMn1_0),.clk(gclk));
	jdff dff_A_2BzIJhw14_0(.dout(w_dff_A_y9h8Fv2q9_0),.din(w_dff_A_2BzIJhw14_0),.clk(gclk));
	jdff dff_A_y9h8Fv2q9_0(.dout(w_dff_A_MFr7mmy71_0),.din(w_dff_A_y9h8Fv2q9_0),.clk(gclk));
	jdff dff_A_MFr7mmy71_0(.dout(w_dff_A_92nXppBQ8_0),.din(w_dff_A_MFr7mmy71_0),.clk(gclk));
	jdff dff_A_92nXppBQ8_0(.dout(w_dff_A_Vlr6wKaK1_0),.din(w_dff_A_92nXppBQ8_0),.clk(gclk));
	jdff dff_A_Vlr6wKaK1_0(.dout(w_dff_A_QuTrwZn00_0),.din(w_dff_A_Vlr6wKaK1_0),.clk(gclk));
	jdff dff_A_QuTrwZn00_0(.dout(w_dff_A_NLUaM75w9_0),.din(w_dff_A_QuTrwZn00_0),.clk(gclk));
	jdff dff_A_NLUaM75w9_0(.dout(w_dff_A_Tp2fn0a22_0),.din(w_dff_A_NLUaM75w9_0),.clk(gclk));
	jdff dff_A_Tp2fn0a22_0(.dout(w_dff_A_ebvaHMAG2_0),.din(w_dff_A_Tp2fn0a22_0),.clk(gclk));
	jdff dff_A_ebvaHMAG2_0(.dout(w_dff_A_iqBvkcJP9_0),.din(w_dff_A_ebvaHMAG2_0),.clk(gclk));
	jdff dff_A_iqBvkcJP9_0(.dout(w_dff_A_UjCBY7Yj8_0),.din(w_dff_A_iqBvkcJP9_0),.clk(gclk));
	jdff dff_A_UjCBY7Yj8_0(.dout(w_dff_A_wiUo5LgO2_0),.din(w_dff_A_UjCBY7Yj8_0),.clk(gclk));
	jdff dff_A_wiUo5LgO2_0(.dout(G2),.din(w_dff_A_wiUo5LgO2_0),.clk(gclk));
	jdff dff_A_oxIB4Cei6_1(.dout(w_dff_A_KOnG8ukG2_0),.din(w_dff_A_oxIB4Cei6_1),.clk(gclk));
	jdff dff_A_KOnG8ukG2_0(.dout(w_dff_A_jh3p7e118_0),.din(w_dff_A_KOnG8ukG2_0),.clk(gclk));
	jdff dff_A_jh3p7e118_0(.dout(w_dff_A_4lhwOdNW5_0),.din(w_dff_A_jh3p7e118_0),.clk(gclk));
	jdff dff_A_4lhwOdNW5_0(.dout(w_dff_A_iO6niJPu6_0),.din(w_dff_A_4lhwOdNW5_0),.clk(gclk));
	jdff dff_A_iO6niJPu6_0(.dout(w_dff_A_KnX3nX9b1_0),.din(w_dff_A_iO6niJPu6_0),.clk(gclk));
	jdff dff_A_KnX3nX9b1_0(.dout(w_dff_A_GXzK9WtO3_0),.din(w_dff_A_KnX3nX9b1_0),.clk(gclk));
	jdff dff_A_GXzK9WtO3_0(.dout(w_dff_A_WZGcfpE69_0),.din(w_dff_A_GXzK9WtO3_0),.clk(gclk));
	jdff dff_A_WZGcfpE69_0(.dout(w_dff_A_z2YVascr1_0),.din(w_dff_A_WZGcfpE69_0),.clk(gclk));
	jdff dff_A_z2YVascr1_0(.dout(w_dff_A_mgsOG2QB8_0),.din(w_dff_A_z2YVascr1_0),.clk(gclk));
	jdff dff_A_mgsOG2QB8_0(.dout(w_dff_A_jMQ72mdi0_0),.din(w_dff_A_mgsOG2QB8_0),.clk(gclk));
	jdff dff_A_jMQ72mdi0_0(.dout(w_dff_A_jbC9VSDC0_0),.din(w_dff_A_jMQ72mdi0_0),.clk(gclk));
	jdff dff_A_jbC9VSDC0_0(.dout(w_dff_A_mJAmcchH5_0),.din(w_dff_A_jbC9VSDC0_0),.clk(gclk));
	jdff dff_A_mJAmcchH5_0(.dout(w_dff_A_QHUvUFHM0_0),.din(w_dff_A_mJAmcchH5_0),.clk(gclk));
	jdff dff_A_QHUvUFHM0_0(.dout(w_dff_A_WxDVy1df7_0),.din(w_dff_A_QHUvUFHM0_0),.clk(gclk));
	jdff dff_A_WxDVy1df7_0(.dout(w_dff_A_4YyXivOI6_0),.din(w_dff_A_WxDVy1df7_0),.clk(gclk));
	jdff dff_A_4YyXivOI6_0(.dout(w_dff_A_hMS5KX0s6_0),.din(w_dff_A_4YyXivOI6_0),.clk(gclk));
	jdff dff_A_hMS5KX0s6_0(.dout(w_dff_A_wasIBB1m9_0),.din(w_dff_A_hMS5KX0s6_0),.clk(gclk));
	jdff dff_A_wasIBB1m9_0(.dout(w_dff_A_AVda3LZ30_0),.din(w_dff_A_wasIBB1m9_0),.clk(gclk));
	jdff dff_A_AVda3LZ30_0(.dout(w_dff_A_ZAWGvtXM1_0),.din(w_dff_A_AVda3LZ30_0),.clk(gclk));
	jdff dff_A_ZAWGvtXM1_0(.dout(w_dff_A_E1S6cTHU0_0),.din(w_dff_A_ZAWGvtXM1_0),.clk(gclk));
	jdff dff_A_E1S6cTHU0_0(.dout(w_dff_A_PhKk96Qz8_0),.din(w_dff_A_E1S6cTHU0_0),.clk(gclk));
	jdff dff_A_PhKk96Qz8_0(.dout(w_dff_A_hQldPRiL2_0),.din(w_dff_A_PhKk96Qz8_0),.clk(gclk));
	jdff dff_A_hQldPRiL2_0(.dout(w_dff_A_5TME2nT46_0),.din(w_dff_A_hQldPRiL2_0),.clk(gclk));
	jdff dff_A_5TME2nT46_0(.dout(w_dff_A_PNMpFsm19_0),.din(w_dff_A_5TME2nT46_0),.clk(gclk));
	jdff dff_A_PNMpFsm19_0(.dout(w_dff_A_XUoaSZcL4_0),.din(w_dff_A_PNMpFsm19_0),.clk(gclk));
	jdff dff_A_XUoaSZcL4_0(.dout(w_dff_A_5pOQ5Aju4_0),.din(w_dff_A_XUoaSZcL4_0),.clk(gclk));
	jdff dff_A_5pOQ5Aju4_0(.dout(G3),.din(w_dff_A_5pOQ5Aju4_0),.clk(gclk));
	jdff dff_A_10WK5Ss63_1(.dout(w_dff_A_m2OXd8GU0_0),.din(w_dff_A_10WK5Ss63_1),.clk(gclk));
	jdff dff_A_m2OXd8GU0_0(.dout(w_dff_A_RCj1M2n81_0),.din(w_dff_A_m2OXd8GU0_0),.clk(gclk));
	jdff dff_A_RCj1M2n81_0(.dout(w_dff_A_5GzlOVEQ3_0),.din(w_dff_A_RCj1M2n81_0),.clk(gclk));
	jdff dff_A_5GzlOVEQ3_0(.dout(w_dff_A_HtgsWHLE0_0),.din(w_dff_A_5GzlOVEQ3_0),.clk(gclk));
	jdff dff_A_HtgsWHLE0_0(.dout(w_dff_A_wLAdzhAG7_0),.din(w_dff_A_HtgsWHLE0_0),.clk(gclk));
	jdff dff_A_wLAdzhAG7_0(.dout(w_dff_A_1FTqlbdL8_0),.din(w_dff_A_wLAdzhAG7_0),.clk(gclk));
	jdff dff_A_1FTqlbdL8_0(.dout(w_dff_A_1qKZGVgd2_0),.din(w_dff_A_1FTqlbdL8_0),.clk(gclk));
	jdff dff_A_1qKZGVgd2_0(.dout(w_dff_A_mg5a3Dd29_0),.din(w_dff_A_1qKZGVgd2_0),.clk(gclk));
	jdff dff_A_mg5a3Dd29_0(.dout(w_dff_A_7xglEOUm7_0),.din(w_dff_A_mg5a3Dd29_0),.clk(gclk));
	jdff dff_A_7xglEOUm7_0(.dout(w_dff_A_IGgBAqn46_0),.din(w_dff_A_7xglEOUm7_0),.clk(gclk));
	jdff dff_A_IGgBAqn46_0(.dout(w_dff_A_vYWqheHh5_0),.din(w_dff_A_IGgBAqn46_0),.clk(gclk));
	jdff dff_A_vYWqheHh5_0(.dout(w_dff_A_DdIWD3GI6_0),.din(w_dff_A_vYWqheHh5_0),.clk(gclk));
	jdff dff_A_DdIWD3GI6_0(.dout(w_dff_A_tENZkOfu9_0),.din(w_dff_A_DdIWD3GI6_0),.clk(gclk));
	jdff dff_A_tENZkOfu9_0(.dout(w_dff_A_5rECpUAp8_0),.din(w_dff_A_tENZkOfu9_0),.clk(gclk));
	jdff dff_A_5rECpUAp8_0(.dout(w_dff_A_ai9ESNxo3_0),.din(w_dff_A_5rECpUAp8_0),.clk(gclk));
	jdff dff_A_ai9ESNxo3_0(.dout(w_dff_A_HPVVcXE57_0),.din(w_dff_A_ai9ESNxo3_0),.clk(gclk));
	jdff dff_A_HPVVcXE57_0(.dout(w_dff_A_2fFXPoYH3_0),.din(w_dff_A_HPVVcXE57_0),.clk(gclk));
	jdff dff_A_2fFXPoYH3_0(.dout(w_dff_A_xs0vf9sa5_0),.din(w_dff_A_2fFXPoYH3_0),.clk(gclk));
	jdff dff_A_xs0vf9sa5_0(.dout(w_dff_A_4DCGFR3V4_0),.din(w_dff_A_xs0vf9sa5_0),.clk(gclk));
	jdff dff_A_4DCGFR3V4_0(.dout(w_dff_A_1D8OSKsX3_0),.din(w_dff_A_4DCGFR3V4_0),.clk(gclk));
	jdff dff_A_1D8OSKsX3_0(.dout(w_dff_A_Wx07uk4D7_0),.din(w_dff_A_1D8OSKsX3_0),.clk(gclk));
	jdff dff_A_Wx07uk4D7_0(.dout(w_dff_A_6HNy7nDt6_0),.din(w_dff_A_Wx07uk4D7_0),.clk(gclk));
	jdff dff_A_6HNy7nDt6_0(.dout(w_dff_A_rEOCcJTv9_0),.din(w_dff_A_6HNy7nDt6_0),.clk(gclk));
	jdff dff_A_rEOCcJTv9_0(.dout(w_dff_A_ocrFkLCU5_0),.din(w_dff_A_rEOCcJTv9_0),.clk(gclk));
	jdff dff_A_ocrFkLCU5_0(.dout(w_dff_A_UohQTphH9_0),.din(w_dff_A_ocrFkLCU5_0),.clk(gclk));
	jdff dff_A_UohQTphH9_0(.dout(w_dff_A_jFIevkki1_0),.din(w_dff_A_UohQTphH9_0),.clk(gclk));
	jdff dff_A_jFIevkki1_0(.dout(G450),.din(w_dff_A_jFIevkki1_0),.clk(gclk));
	jdff dff_A_kCaRS6Sy6_1(.dout(w_dff_A_FZW6VcR89_0),.din(w_dff_A_kCaRS6Sy6_1),.clk(gclk));
	jdff dff_A_FZW6VcR89_0(.dout(w_dff_A_oVX9haIk8_0),.din(w_dff_A_FZW6VcR89_0),.clk(gclk));
	jdff dff_A_oVX9haIk8_0(.dout(w_dff_A_rdUe9k8F7_0),.din(w_dff_A_oVX9haIk8_0),.clk(gclk));
	jdff dff_A_rdUe9k8F7_0(.dout(w_dff_A_CAZqmPnc3_0),.din(w_dff_A_rdUe9k8F7_0),.clk(gclk));
	jdff dff_A_CAZqmPnc3_0(.dout(w_dff_A_xL6t0IWm9_0),.din(w_dff_A_CAZqmPnc3_0),.clk(gclk));
	jdff dff_A_xL6t0IWm9_0(.dout(w_dff_A_JE4n6kCm7_0),.din(w_dff_A_xL6t0IWm9_0),.clk(gclk));
	jdff dff_A_JE4n6kCm7_0(.dout(w_dff_A_J9FZsDMu4_0),.din(w_dff_A_JE4n6kCm7_0),.clk(gclk));
	jdff dff_A_J9FZsDMu4_0(.dout(w_dff_A_mmmFMqzu3_0),.din(w_dff_A_J9FZsDMu4_0),.clk(gclk));
	jdff dff_A_mmmFMqzu3_0(.dout(w_dff_A_NppFIkLE8_0),.din(w_dff_A_mmmFMqzu3_0),.clk(gclk));
	jdff dff_A_NppFIkLE8_0(.dout(w_dff_A_4OarWApE4_0),.din(w_dff_A_NppFIkLE8_0),.clk(gclk));
	jdff dff_A_4OarWApE4_0(.dout(w_dff_A_ZuUukkmu1_0),.din(w_dff_A_4OarWApE4_0),.clk(gclk));
	jdff dff_A_ZuUukkmu1_0(.dout(w_dff_A_QOHK88YV2_0),.din(w_dff_A_ZuUukkmu1_0),.clk(gclk));
	jdff dff_A_QOHK88YV2_0(.dout(w_dff_A_wh25BaB73_0),.din(w_dff_A_QOHK88YV2_0),.clk(gclk));
	jdff dff_A_wh25BaB73_0(.dout(w_dff_A_qIvWoEdV6_0),.din(w_dff_A_wh25BaB73_0),.clk(gclk));
	jdff dff_A_qIvWoEdV6_0(.dout(w_dff_A_TeDyRX4V6_0),.din(w_dff_A_qIvWoEdV6_0),.clk(gclk));
	jdff dff_A_TeDyRX4V6_0(.dout(w_dff_A_pEO0k3Wb7_0),.din(w_dff_A_TeDyRX4V6_0),.clk(gclk));
	jdff dff_A_pEO0k3Wb7_0(.dout(w_dff_A_K2w6pVw00_0),.din(w_dff_A_pEO0k3Wb7_0),.clk(gclk));
	jdff dff_A_K2w6pVw00_0(.dout(w_dff_A_cCe9KEAq6_0),.din(w_dff_A_K2w6pVw00_0),.clk(gclk));
	jdff dff_A_cCe9KEAq6_0(.dout(w_dff_A_OgnbogKE4_0),.din(w_dff_A_cCe9KEAq6_0),.clk(gclk));
	jdff dff_A_OgnbogKE4_0(.dout(w_dff_A_z0N22mwn7_0),.din(w_dff_A_OgnbogKE4_0),.clk(gclk));
	jdff dff_A_z0N22mwn7_0(.dout(w_dff_A_9OXmE5QW8_0),.din(w_dff_A_z0N22mwn7_0),.clk(gclk));
	jdff dff_A_9OXmE5QW8_0(.dout(w_dff_A_tSplufwi4_0),.din(w_dff_A_9OXmE5QW8_0),.clk(gclk));
	jdff dff_A_tSplufwi4_0(.dout(w_dff_A_jJoz5WTJ6_0),.din(w_dff_A_tSplufwi4_0),.clk(gclk));
	jdff dff_A_jJoz5WTJ6_0(.dout(w_dff_A_WeVAw1Fr1_0),.din(w_dff_A_jJoz5WTJ6_0),.clk(gclk));
	jdff dff_A_WeVAw1Fr1_0(.dout(w_dff_A_xgD2f48o8_0),.din(w_dff_A_WeVAw1Fr1_0),.clk(gclk));
	jdff dff_A_xgD2f48o8_0(.dout(w_dff_A_mPJ9Ru6q4_0),.din(w_dff_A_xgD2f48o8_0),.clk(gclk));
	jdff dff_A_mPJ9Ru6q4_0(.dout(G448),.din(w_dff_A_mPJ9Ru6q4_0),.clk(gclk));
	jdff dff_A_tz2EUH5g2_1(.dout(w_dff_A_9mG3Lu1n0_0),.din(w_dff_A_tz2EUH5g2_1),.clk(gclk));
	jdff dff_A_9mG3Lu1n0_0(.dout(w_dff_A_yidHp8eC2_0),.din(w_dff_A_9mG3Lu1n0_0),.clk(gclk));
	jdff dff_A_yidHp8eC2_0(.dout(w_dff_A_VzXCQxLY9_0),.din(w_dff_A_yidHp8eC2_0),.clk(gclk));
	jdff dff_A_VzXCQxLY9_0(.dout(w_dff_A_R7HlyTZD5_0),.din(w_dff_A_VzXCQxLY9_0),.clk(gclk));
	jdff dff_A_R7HlyTZD5_0(.dout(w_dff_A_nO9k76IR3_0),.din(w_dff_A_R7HlyTZD5_0),.clk(gclk));
	jdff dff_A_nO9k76IR3_0(.dout(w_dff_A_eorpBthw2_0),.din(w_dff_A_nO9k76IR3_0),.clk(gclk));
	jdff dff_A_eorpBthw2_0(.dout(w_dff_A_xlEygdER1_0),.din(w_dff_A_eorpBthw2_0),.clk(gclk));
	jdff dff_A_xlEygdER1_0(.dout(w_dff_A_1CxfVFdc6_0),.din(w_dff_A_xlEygdER1_0),.clk(gclk));
	jdff dff_A_1CxfVFdc6_0(.dout(w_dff_A_Di5cysJZ0_0),.din(w_dff_A_1CxfVFdc6_0),.clk(gclk));
	jdff dff_A_Di5cysJZ0_0(.dout(w_dff_A_ks31prln2_0),.din(w_dff_A_Di5cysJZ0_0),.clk(gclk));
	jdff dff_A_ks31prln2_0(.dout(w_dff_A_DX9SLhis1_0),.din(w_dff_A_ks31prln2_0),.clk(gclk));
	jdff dff_A_DX9SLhis1_0(.dout(w_dff_A_CY3Dw0K33_0),.din(w_dff_A_DX9SLhis1_0),.clk(gclk));
	jdff dff_A_CY3Dw0K33_0(.dout(w_dff_A_v92hmE3l7_0),.din(w_dff_A_CY3Dw0K33_0),.clk(gclk));
	jdff dff_A_v92hmE3l7_0(.dout(w_dff_A_ew1OSBIm6_0),.din(w_dff_A_v92hmE3l7_0),.clk(gclk));
	jdff dff_A_ew1OSBIm6_0(.dout(w_dff_A_aLXiHK0v8_0),.din(w_dff_A_ew1OSBIm6_0),.clk(gclk));
	jdff dff_A_aLXiHK0v8_0(.dout(w_dff_A_GUxv8NP97_0),.din(w_dff_A_aLXiHK0v8_0),.clk(gclk));
	jdff dff_A_GUxv8NP97_0(.dout(w_dff_A_56JtU3Z06_0),.din(w_dff_A_GUxv8NP97_0),.clk(gclk));
	jdff dff_A_56JtU3Z06_0(.dout(w_dff_A_mEWlNEV93_0),.din(w_dff_A_56JtU3Z06_0),.clk(gclk));
	jdff dff_A_mEWlNEV93_0(.dout(w_dff_A_uLRusD744_0),.din(w_dff_A_mEWlNEV93_0),.clk(gclk));
	jdff dff_A_uLRusD744_0(.dout(w_dff_A_I9OZLL0H9_0),.din(w_dff_A_uLRusD744_0),.clk(gclk));
	jdff dff_A_I9OZLL0H9_0(.dout(w_dff_A_jjejcgTo5_0),.din(w_dff_A_I9OZLL0H9_0),.clk(gclk));
	jdff dff_A_jjejcgTo5_0(.dout(w_dff_A_84PfOtyr1_0),.din(w_dff_A_jjejcgTo5_0),.clk(gclk));
	jdff dff_A_84PfOtyr1_0(.dout(w_dff_A_vTTYpNhr7_0),.din(w_dff_A_84PfOtyr1_0),.clk(gclk));
	jdff dff_A_vTTYpNhr7_0(.dout(w_dff_A_KdvfegDV5_0),.din(w_dff_A_vTTYpNhr7_0),.clk(gclk));
	jdff dff_A_KdvfegDV5_0(.dout(w_dff_A_iXZXkzMz3_0),.din(w_dff_A_KdvfegDV5_0),.clk(gclk));
	jdff dff_A_iXZXkzMz3_0(.dout(w_dff_A_Ey1u0GRR4_0),.din(w_dff_A_iXZXkzMz3_0),.clk(gclk));
	jdff dff_A_Ey1u0GRR4_0(.dout(G444),.din(w_dff_A_Ey1u0GRR4_0),.clk(gclk));
	jdff dff_A_n6GEbAPE9_1(.dout(w_dff_A_vhSL0ylA8_0),.din(w_dff_A_n6GEbAPE9_1),.clk(gclk));
	jdff dff_A_vhSL0ylA8_0(.dout(w_dff_A_vuaj4YVy1_0),.din(w_dff_A_vhSL0ylA8_0),.clk(gclk));
	jdff dff_A_vuaj4YVy1_0(.dout(w_dff_A_ouZwcVQa8_0),.din(w_dff_A_vuaj4YVy1_0),.clk(gclk));
	jdff dff_A_ouZwcVQa8_0(.dout(w_dff_A_uacfhTVx2_0),.din(w_dff_A_ouZwcVQa8_0),.clk(gclk));
	jdff dff_A_uacfhTVx2_0(.dout(w_dff_A_m98kHR7B0_0),.din(w_dff_A_uacfhTVx2_0),.clk(gclk));
	jdff dff_A_m98kHR7B0_0(.dout(w_dff_A_scQK8cxc2_0),.din(w_dff_A_m98kHR7B0_0),.clk(gclk));
	jdff dff_A_scQK8cxc2_0(.dout(w_dff_A_2dNb6GiG8_0),.din(w_dff_A_scQK8cxc2_0),.clk(gclk));
	jdff dff_A_2dNb6GiG8_0(.dout(w_dff_A_kHsCSco35_0),.din(w_dff_A_2dNb6GiG8_0),.clk(gclk));
	jdff dff_A_kHsCSco35_0(.dout(w_dff_A_gsTwXeFl2_0),.din(w_dff_A_kHsCSco35_0),.clk(gclk));
	jdff dff_A_gsTwXeFl2_0(.dout(w_dff_A_YgeZsEwQ0_0),.din(w_dff_A_gsTwXeFl2_0),.clk(gclk));
	jdff dff_A_YgeZsEwQ0_0(.dout(w_dff_A_nKeS3DuD6_0),.din(w_dff_A_YgeZsEwQ0_0),.clk(gclk));
	jdff dff_A_nKeS3DuD6_0(.dout(w_dff_A_63u1S9YW9_0),.din(w_dff_A_nKeS3DuD6_0),.clk(gclk));
	jdff dff_A_63u1S9YW9_0(.dout(w_dff_A_w9f6qIDK0_0),.din(w_dff_A_63u1S9YW9_0),.clk(gclk));
	jdff dff_A_w9f6qIDK0_0(.dout(w_dff_A_Qk3nP7Dl8_0),.din(w_dff_A_w9f6qIDK0_0),.clk(gclk));
	jdff dff_A_Qk3nP7Dl8_0(.dout(w_dff_A_lRTTKe4K8_0),.din(w_dff_A_Qk3nP7Dl8_0),.clk(gclk));
	jdff dff_A_lRTTKe4K8_0(.dout(w_dff_A_RoPD4Z1f3_0),.din(w_dff_A_lRTTKe4K8_0),.clk(gclk));
	jdff dff_A_RoPD4Z1f3_0(.dout(w_dff_A_dDsFKOM42_0),.din(w_dff_A_RoPD4Z1f3_0),.clk(gclk));
	jdff dff_A_dDsFKOM42_0(.dout(w_dff_A_m2JKHjhT5_0),.din(w_dff_A_dDsFKOM42_0),.clk(gclk));
	jdff dff_A_m2JKHjhT5_0(.dout(w_dff_A_IozIKX6i6_0),.din(w_dff_A_m2JKHjhT5_0),.clk(gclk));
	jdff dff_A_IozIKX6i6_0(.dout(w_dff_A_LnbujqxW7_0),.din(w_dff_A_IozIKX6i6_0),.clk(gclk));
	jdff dff_A_LnbujqxW7_0(.dout(w_dff_A_OruZdeSh4_0),.din(w_dff_A_LnbujqxW7_0),.clk(gclk));
	jdff dff_A_OruZdeSh4_0(.dout(w_dff_A_lJltIt2F9_0),.din(w_dff_A_OruZdeSh4_0),.clk(gclk));
	jdff dff_A_lJltIt2F9_0(.dout(w_dff_A_0J1PsqUz8_0),.din(w_dff_A_lJltIt2F9_0),.clk(gclk));
	jdff dff_A_0J1PsqUz8_0(.dout(w_dff_A_TvVmRDFc7_0),.din(w_dff_A_0J1PsqUz8_0),.clk(gclk));
	jdff dff_A_TvVmRDFc7_0(.dout(w_dff_A_M6XVcSha7_0),.din(w_dff_A_TvVmRDFc7_0),.clk(gclk));
	jdff dff_A_M6XVcSha7_0(.dout(w_dff_A_30PmYXmR9_0),.din(w_dff_A_M6XVcSha7_0),.clk(gclk));
	jdff dff_A_30PmYXmR9_0(.dout(G442),.din(w_dff_A_30PmYXmR9_0),.clk(gclk));
	jdff dff_A_eZCLFuLa4_1(.dout(w_dff_A_OHMTBp7v4_0),.din(w_dff_A_eZCLFuLa4_1),.clk(gclk));
	jdff dff_A_OHMTBp7v4_0(.dout(w_dff_A_2WqyOJTU7_0),.din(w_dff_A_OHMTBp7v4_0),.clk(gclk));
	jdff dff_A_2WqyOJTU7_0(.dout(w_dff_A_hV1p6eWM3_0),.din(w_dff_A_2WqyOJTU7_0),.clk(gclk));
	jdff dff_A_hV1p6eWM3_0(.dout(w_dff_A_gz2Ewt9K0_0),.din(w_dff_A_hV1p6eWM3_0),.clk(gclk));
	jdff dff_A_gz2Ewt9K0_0(.dout(w_dff_A_HYR6Vitj0_0),.din(w_dff_A_gz2Ewt9K0_0),.clk(gclk));
	jdff dff_A_HYR6Vitj0_0(.dout(w_dff_A_lL1Njcps1_0),.din(w_dff_A_HYR6Vitj0_0),.clk(gclk));
	jdff dff_A_lL1Njcps1_0(.dout(w_dff_A_TQQ8cuz43_0),.din(w_dff_A_lL1Njcps1_0),.clk(gclk));
	jdff dff_A_TQQ8cuz43_0(.dout(w_dff_A_xP5lZ3ko5_0),.din(w_dff_A_TQQ8cuz43_0),.clk(gclk));
	jdff dff_A_xP5lZ3ko5_0(.dout(w_dff_A_GaKABU4J6_0),.din(w_dff_A_xP5lZ3ko5_0),.clk(gclk));
	jdff dff_A_GaKABU4J6_0(.dout(w_dff_A_E5uWkL2w0_0),.din(w_dff_A_GaKABU4J6_0),.clk(gclk));
	jdff dff_A_E5uWkL2w0_0(.dout(w_dff_A_QtjBnO1x7_0),.din(w_dff_A_E5uWkL2w0_0),.clk(gclk));
	jdff dff_A_QtjBnO1x7_0(.dout(w_dff_A_D3YpL1SM3_0),.din(w_dff_A_QtjBnO1x7_0),.clk(gclk));
	jdff dff_A_D3YpL1SM3_0(.dout(w_dff_A_s7s0FuBn6_0),.din(w_dff_A_D3YpL1SM3_0),.clk(gclk));
	jdff dff_A_s7s0FuBn6_0(.dout(w_dff_A_olkoY8rg5_0),.din(w_dff_A_s7s0FuBn6_0),.clk(gclk));
	jdff dff_A_olkoY8rg5_0(.dout(w_dff_A_mP9VXzn46_0),.din(w_dff_A_olkoY8rg5_0),.clk(gclk));
	jdff dff_A_mP9VXzn46_0(.dout(w_dff_A_uUU6biFu6_0),.din(w_dff_A_mP9VXzn46_0),.clk(gclk));
	jdff dff_A_uUU6biFu6_0(.dout(w_dff_A_AY5aMxLv5_0),.din(w_dff_A_uUU6biFu6_0),.clk(gclk));
	jdff dff_A_AY5aMxLv5_0(.dout(w_dff_A_kcvpou7C5_0),.din(w_dff_A_AY5aMxLv5_0),.clk(gclk));
	jdff dff_A_kcvpou7C5_0(.dout(w_dff_A_sYxXon2S1_0),.din(w_dff_A_kcvpou7C5_0),.clk(gclk));
	jdff dff_A_sYxXon2S1_0(.dout(w_dff_A_CwLKBqSc5_0),.din(w_dff_A_sYxXon2S1_0),.clk(gclk));
	jdff dff_A_CwLKBqSc5_0(.dout(w_dff_A_8Zpj7t9g1_0),.din(w_dff_A_CwLKBqSc5_0),.clk(gclk));
	jdff dff_A_8Zpj7t9g1_0(.dout(w_dff_A_rPs7T8ai0_0),.din(w_dff_A_8Zpj7t9g1_0),.clk(gclk));
	jdff dff_A_rPs7T8ai0_0(.dout(w_dff_A_yZRROB5r1_0),.din(w_dff_A_rPs7T8ai0_0),.clk(gclk));
	jdff dff_A_yZRROB5r1_0(.dout(w_dff_A_hBWYzKIH4_0),.din(w_dff_A_yZRROB5r1_0),.clk(gclk));
	jdff dff_A_hBWYzKIH4_0(.dout(w_dff_A_1fOOLZ0z6_0),.din(w_dff_A_hBWYzKIH4_0),.clk(gclk));
	jdff dff_A_1fOOLZ0z6_0(.dout(w_dff_A_FVnoGUp58_0),.din(w_dff_A_1fOOLZ0z6_0),.clk(gclk));
	jdff dff_A_FVnoGUp58_0(.dout(G440),.din(w_dff_A_FVnoGUp58_0),.clk(gclk));
	jdff dff_A_7VdHePjq5_1(.dout(w_dff_A_eLwjgnpG0_0),.din(w_dff_A_7VdHePjq5_1),.clk(gclk));
	jdff dff_A_eLwjgnpG0_0(.dout(w_dff_A_NV3ofKnU2_0),.din(w_dff_A_eLwjgnpG0_0),.clk(gclk));
	jdff dff_A_NV3ofKnU2_0(.dout(w_dff_A_r6ZTE5W39_0),.din(w_dff_A_NV3ofKnU2_0),.clk(gclk));
	jdff dff_A_r6ZTE5W39_0(.dout(w_dff_A_LXc8bHfA0_0),.din(w_dff_A_r6ZTE5W39_0),.clk(gclk));
	jdff dff_A_LXc8bHfA0_0(.dout(w_dff_A_2xkbbBgt0_0),.din(w_dff_A_LXc8bHfA0_0),.clk(gclk));
	jdff dff_A_2xkbbBgt0_0(.dout(w_dff_A_hW0Jx9WF0_0),.din(w_dff_A_2xkbbBgt0_0),.clk(gclk));
	jdff dff_A_hW0Jx9WF0_0(.dout(w_dff_A_Y74ITYZM9_0),.din(w_dff_A_hW0Jx9WF0_0),.clk(gclk));
	jdff dff_A_Y74ITYZM9_0(.dout(w_dff_A_JYT21bjO0_0),.din(w_dff_A_Y74ITYZM9_0),.clk(gclk));
	jdff dff_A_JYT21bjO0_0(.dout(w_dff_A_DByppb385_0),.din(w_dff_A_JYT21bjO0_0),.clk(gclk));
	jdff dff_A_DByppb385_0(.dout(w_dff_A_oysh2A488_0),.din(w_dff_A_DByppb385_0),.clk(gclk));
	jdff dff_A_oysh2A488_0(.dout(w_dff_A_jgjOjtK23_0),.din(w_dff_A_oysh2A488_0),.clk(gclk));
	jdff dff_A_jgjOjtK23_0(.dout(w_dff_A_3Xy3xQz45_0),.din(w_dff_A_jgjOjtK23_0),.clk(gclk));
	jdff dff_A_3Xy3xQz45_0(.dout(w_dff_A_dtY1ZSAz4_0),.din(w_dff_A_3Xy3xQz45_0),.clk(gclk));
	jdff dff_A_dtY1ZSAz4_0(.dout(w_dff_A_47B6qsAS5_0),.din(w_dff_A_dtY1ZSAz4_0),.clk(gclk));
	jdff dff_A_47B6qsAS5_0(.dout(w_dff_A_dpBByX4E1_0),.din(w_dff_A_47B6qsAS5_0),.clk(gclk));
	jdff dff_A_dpBByX4E1_0(.dout(w_dff_A_nTUDBs2i7_0),.din(w_dff_A_dpBByX4E1_0),.clk(gclk));
	jdff dff_A_nTUDBs2i7_0(.dout(w_dff_A_sz9DWv3j3_0),.din(w_dff_A_nTUDBs2i7_0),.clk(gclk));
	jdff dff_A_sz9DWv3j3_0(.dout(w_dff_A_AbspSUIb2_0),.din(w_dff_A_sz9DWv3j3_0),.clk(gclk));
	jdff dff_A_AbspSUIb2_0(.dout(w_dff_A_funZxtua1_0),.din(w_dff_A_AbspSUIb2_0),.clk(gclk));
	jdff dff_A_funZxtua1_0(.dout(w_dff_A_Z1Fvwk8Q9_0),.din(w_dff_A_funZxtua1_0),.clk(gclk));
	jdff dff_A_Z1Fvwk8Q9_0(.dout(w_dff_A_Xi1zp94q0_0),.din(w_dff_A_Z1Fvwk8Q9_0),.clk(gclk));
	jdff dff_A_Xi1zp94q0_0(.dout(w_dff_A_m8bmpBbW6_0),.din(w_dff_A_Xi1zp94q0_0),.clk(gclk));
	jdff dff_A_m8bmpBbW6_0(.dout(w_dff_A_xSjSqwBd2_0),.din(w_dff_A_m8bmpBbW6_0),.clk(gclk));
	jdff dff_A_xSjSqwBd2_0(.dout(w_dff_A_IHoLcdss3_0),.din(w_dff_A_xSjSqwBd2_0),.clk(gclk));
	jdff dff_A_IHoLcdss3_0(.dout(w_dff_A_jz5NWKKy7_0),.din(w_dff_A_IHoLcdss3_0),.clk(gclk));
	jdff dff_A_jz5NWKKy7_0(.dout(w_dff_A_bqWqExrP5_0),.din(w_dff_A_jz5NWKKy7_0),.clk(gclk));
	jdff dff_A_bqWqExrP5_0(.dout(G438),.din(w_dff_A_bqWqExrP5_0),.clk(gclk));
	jdff dff_A_l63WIzjM6_1(.dout(w_dff_A_erv3MoCl6_0),.din(w_dff_A_l63WIzjM6_1),.clk(gclk));
	jdff dff_A_erv3MoCl6_0(.dout(w_dff_A_23Nzfjzz4_0),.din(w_dff_A_erv3MoCl6_0),.clk(gclk));
	jdff dff_A_23Nzfjzz4_0(.dout(w_dff_A_hDA8oJ3Z7_0),.din(w_dff_A_23Nzfjzz4_0),.clk(gclk));
	jdff dff_A_hDA8oJ3Z7_0(.dout(w_dff_A_Si5JKb6B2_0),.din(w_dff_A_hDA8oJ3Z7_0),.clk(gclk));
	jdff dff_A_Si5JKb6B2_0(.dout(w_dff_A_1GH6aFFI7_0),.din(w_dff_A_Si5JKb6B2_0),.clk(gclk));
	jdff dff_A_1GH6aFFI7_0(.dout(w_dff_A_MRMohy7L5_0),.din(w_dff_A_1GH6aFFI7_0),.clk(gclk));
	jdff dff_A_MRMohy7L5_0(.dout(w_dff_A_XIIBFOiR3_0),.din(w_dff_A_MRMohy7L5_0),.clk(gclk));
	jdff dff_A_XIIBFOiR3_0(.dout(w_dff_A_PSGM1cWS1_0),.din(w_dff_A_XIIBFOiR3_0),.clk(gclk));
	jdff dff_A_PSGM1cWS1_0(.dout(w_dff_A_ZQnpKyJs9_0),.din(w_dff_A_PSGM1cWS1_0),.clk(gclk));
	jdff dff_A_ZQnpKyJs9_0(.dout(w_dff_A_WjTic5P82_0),.din(w_dff_A_ZQnpKyJs9_0),.clk(gclk));
	jdff dff_A_WjTic5P82_0(.dout(w_dff_A_ZkwKTgP03_0),.din(w_dff_A_WjTic5P82_0),.clk(gclk));
	jdff dff_A_ZkwKTgP03_0(.dout(w_dff_A_akfZ5Bak4_0),.din(w_dff_A_ZkwKTgP03_0),.clk(gclk));
	jdff dff_A_akfZ5Bak4_0(.dout(w_dff_A_wFHvd1Lq0_0),.din(w_dff_A_akfZ5Bak4_0),.clk(gclk));
	jdff dff_A_wFHvd1Lq0_0(.dout(w_dff_A_cpEe7gY65_0),.din(w_dff_A_wFHvd1Lq0_0),.clk(gclk));
	jdff dff_A_cpEe7gY65_0(.dout(w_dff_A_tpmFTXUA6_0),.din(w_dff_A_cpEe7gY65_0),.clk(gclk));
	jdff dff_A_tpmFTXUA6_0(.dout(w_dff_A_U2CRmF4K1_0),.din(w_dff_A_tpmFTXUA6_0),.clk(gclk));
	jdff dff_A_U2CRmF4K1_0(.dout(w_dff_A_WG28kDGY7_0),.din(w_dff_A_U2CRmF4K1_0),.clk(gclk));
	jdff dff_A_WG28kDGY7_0(.dout(w_dff_A_01xXUPsM1_0),.din(w_dff_A_WG28kDGY7_0),.clk(gclk));
	jdff dff_A_01xXUPsM1_0(.dout(w_dff_A_TIL8YHkX0_0),.din(w_dff_A_01xXUPsM1_0),.clk(gclk));
	jdff dff_A_TIL8YHkX0_0(.dout(w_dff_A_CU1mMcyK6_0),.din(w_dff_A_TIL8YHkX0_0),.clk(gclk));
	jdff dff_A_CU1mMcyK6_0(.dout(w_dff_A_2yxsluPl9_0),.din(w_dff_A_CU1mMcyK6_0),.clk(gclk));
	jdff dff_A_2yxsluPl9_0(.dout(w_dff_A_KtuYRaNB8_0),.din(w_dff_A_2yxsluPl9_0),.clk(gclk));
	jdff dff_A_KtuYRaNB8_0(.dout(w_dff_A_7ddChlGP8_0),.din(w_dff_A_KtuYRaNB8_0),.clk(gclk));
	jdff dff_A_7ddChlGP8_0(.dout(w_dff_A_iTrwKClE9_0),.din(w_dff_A_7ddChlGP8_0),.clk(gclk));
	jdff dff_A_iTrwKClE9_0(.dout(w_dff_A_hRSgFL8V2_0),.din(w_dff_A_iTrwKClE9_0),.clk(gclk));
	jdff dff_A_hRSgFL8V2_0(.dout(w_dff_A_jAg8ipek3_0),.din(w_dff_A_hRSgFL8V2_0),.clk(gclk));
	jdff dff_A_jAg8ipek3_0(.dout(G496),.din(w_dff_A_jAg8ipek3_0),.clk(gclk));
	jdff dff_A_38SOXGaA5_1(.dout(w_dff_A_KeiJ0RtT9_0),.din(w_dff_A_38SOXGaA5_1),.clk(gclk));
	jdff dff_A_KeiJ0RtT9_0(.dout(w_dff_A_QgRBCdsL6_0),.din(w_dff_A_KeiJ0RtT9_0),.clk(gclk));
	jdff dff_A_QgRBCdsL6_0(.dout(w_dff_A_VRFKqh112_0),.din(w_dff_A_QgRBCdsL6_0),.clk(gclk));
	jdff dff_A_VRFKqh112_0(.dout(w_dff_A_3mv3czMj9_0),.din(w_dff_A_VRFKqh112_0),.clk(gclk));
	jdff dff_A_3mv3czMj9_0(.dout(w_dff_A_uXxTkFel7_0),.din(w_dff_A_3mv3czMj9_0),.clk(gclk));
	jdff dff_A_uXxTkFel7_0(.dout(w_dff_A_95MWKwuz3_0),.din(w_dff_A_uXxTkFel7_0),.clk(gclk));
	jdff dff_A_95MWKwuz3_0(.dout(w_dff_A_NI4HY9Il8_0),.din(w_dff_A_95MWKwuz3_0),.clk(gclk));
	jdff dff_A_NI4HY9Il8_0(.dout(w_dff_A_jcH6biH79_0),.din(w_dff_A_NI4HY9Il8_0),.clk(gclk));
	jdff dff_A_jcH6biH79_0(.dout(w_dff_A_S9yFVrOo8_0),.din(w_dff_A_jcH6biH79_0),.clk(gclk));
	jdff dff_A_S9yFVrOo8_0(.dout(w_dff_A_oawsxvSq5_0),.din(w_dff_A_S9yFVrOo8_0),.clk(gclk));
	jdff dff_A_oawsxvSq5_0(.dout(w_dff_A_c60nqKA02_0),.din(w_dff_A_oawsxvSq5_0),.clk(gclk));
	jdff dff_A_c60nqKA02_0(.dout(w_dff_A_vh672oYT7_0),.din(w_dff_A_c60nqKA02_0),.clk(gclk));
	jdff dff_A_vh672oYT7_0(.dout(w_dff_A_ubt47kOw0_0),.din(w_dff_A_vh672oYT7_0),.clk(gclk));
	jdff dff_A_ubt47kOw0_0(.dout(w_dff_A_QG4AoQJX8_0),.din(w_dff_A_ubt47kOw0_0),.clk(gclk));
	jdff dff_A_QG4AoQJX8_0(.dout(w_dff_A_q4MuepBg4_0),.din(w_dff_A_QG4AoQJX8_0),.clk(gclk));
	jdff dff_A_q4MuepBg4_0(.dout(w_dff_A_trZDxp1t2_0),.din(w_dff_A_q4MuepBg4_0),.clk(gclk));
	jdff dff_A_trZDxp1t2_0(.dout(w_dff_A_5cCi84ZB8_0),.din(w_dff_A_trZDxp1t2_0),.clk(gclk));
	jdff dff_A_5cCi84ZB8_0(.dout(w_dff_A_N74xfBax7_0),.din(w_dff_A_5cCi84ZB8_0),.clk(gclk));
	jdff dff_A_N74xfBax7_0(.dout(w_dff_A_e6ywPm164_0),.din(w_dff_A_N74xfBax7_0),.clk(gclk));
	jdff dff_A_e6ywPm164_0(.dout(w_dff_A_fWhcDEEt4_0),.din(w_dff_A_e6ywPm164_0),.clk(gclk));
	jdff dff_A_fWhcDEEt4_0(.dout(w_dff_A_jHUD2lfR3_0),.din(w_dff_A_fWhcDEEt4_0),.clk(gclk));
	jdff dff_A_jHUD2lfR3_0(.dout(w_dff_A_rNKzjgPj4_0),.din(w_dff_A_jHUD2lfR3_0),.clk(gclk));
	jdff dff_A_rNKzjgPj4_0(.dout(w_dff_A_WCVQz6gw3_0),.din(w_dff_A_rNKzjgPj4_0),.clk(gclk));
	jdff dff_A_WCVQz6gw3_0(.dout(w_dff_A_jhG2YlK52_0),.din(w_dff_A_WCVQz6gw3_0),.clk(gclk));
	jdff dff_A_jhG2YlK52_0(.dout(w_dff_A_yVL49AWJ9_0),.din(w_dff_A_jhG2YlK52_0),.clk(gclk));
	jdff dff_A_yVL49AWJ9_0(.dout(w_dff_A_d1yeIUe78_0),.din(w_dff_A_yVL49AWJ9_0),.clk(gclk));
	jdff dff_A_d1yeIUe78_0(.dout(G494),.din(w_dff_A_d1yeIUe78_0),.clk(gclk));
	jdff dff_A_SUaMaM1Z9_1(.dout(w_dff_A_RfFlRvc98_0),.din(w_dff_A_SUaMaM1Z9_1),.clk(gclk));
	jdff dff_A_RfFlRvc98_0(.dout(w_dff_A_ATamxKvN4_0),.din(w_dff_A_RfFlRvc98_0),.clk(gclk));
	jdff dff_A_ATamxKvN4_0(.dout(w_dff_A_kG7ZOa896_0),.din(w_dff_A_ATamxKvN4_0),.clk(gclk));
	jdff dff_A_kG7ZOa896_0(.dout(w_dff_A_eIOSNxwP7_0),.din(w_dff_A_kG7ZOa896_0),.clk(gclk));
	jdff dff_A_eIOSNxwP7_0(.dout(w_dff_A_wkL8Ws237_0),.din(w_dff_A_eIOSNxwP7_0),.clk(gclk));
	jdff dff_A_wkL8Ws237_0(.dout(w_dff_A_VfyBSNvD5_0),.din(w_dff_A_wkL8Ws237_0),.clk(gclk));
	jdff dff_A_VfyBSNvD5_0(.dout(w_dff_A_IPkdxN7Y4_0),.din(w_dff_A_VfyBSNvD5_0),.clk(gclk));
	jdff dff_A_IPkdxN7Y4_0(.dout(w_dff_A_SipErOe39_0),.din(w_dff_A_IPkdxN7Y4_0),.clk(gclk));
	jdff dff_A_SipErOe39_0(.dout(w_dff_A_I6XeDiTP7_0),.din(w_dff_A_SipErOe39_0),.clk(gclk));
	jdff dff_A_I6XeDiTP7_0(.dout(w_dff_A_UzAQnEMN2_0),.din(w_dff_A_I6XeDiTP7_0),.clk(gclk));
	jdff dff_A_UzAQnEMN2_0(.dout(w_dff_A_GVTsDNjh6_0),.din(w_dff_A_UzAQnEMN2_0),.clk(gclk));
	jdff dff_A_GVTsDNjh6_0(.dout(w_dff_A_tr5CDcJb0_0),.din(w_dff_A_GVTsDNjh6_0),.clk(gclk));
	jdff dff_A_tr5CDcJb0_0(.dout(w_dff_A_56d2YEf73_0),.din(w_dff_A_tr5CDcJb0_0),.clk(gclk));
	jdff dff_A_56d2YEf73_0(.dout(w_dff_A_0zFHMc236_0),.din(w_dff_A_56d2YEf73_0),.clk(gclk));
	jdff dff_A_0zFHMc236_0(.dout(w_dff_A_2dRy7EHp1_0),.din(w_dff_A_0zFHMc236_0),.clk(gclk));
	jdff dff_A_2dRy7EHp1_0(.dout(w_dff_A_GLVV54ps2_0),.din(w_dff_A_2dRy7EHp1_0),.clk(gclk));
	jdff dff_A_GLVV54ps2_0(.dout(w_dff_A_jyWGfFm48_0),.din(w_dff_A_GLVV54ps2_0),.clk(gclk));
	jdff dff_A_jyWGfFm48_0(.dout(w_dff_A_0lk96sWg8_0),.din(w_dff_A_jyWGfFm48_0),.clk(gclk));
	jdff dff_A_0lk96sWg8_0(.dout(w_dff_A_CySS9Psy9_0),.din(w_dff_A_0lk96sWg8_0),.clk(gclk));
	jdff dff_A_CySS9Psy9_0(.dout(w_dff_A_v0zKxZPp7_0),.din(w_dff_A_CySS9Psy9_0),.clk(gclk));
	jdff dff_A_v0zKxZPp7_0(.dout(w_dff_A_KZO5bQBU7_0),.din(w_dff_A_v0zKxZPp7_0),.clk(gclk));
	jdff dff_A_KZO5bQBU7_0(.dout(w_dff_A_XjBCg3ig5_0),.din(w_dff_A_KZO5bQBU7_0),.clk(gclk));
	jdff dff_A_XjBCg3ig5_0(.dout(w_dff_A_NSg3Al6P0_0),.din(w_dff_A_XjBCg3ig5_0),.clk(gclk));
	jdff dff_A_NSg3Al6P0_0(.dout(w_dff_A_Adf9uIwU5_0),.din(w_dff_A_NSg3Al6P0_0),.clk(gclk));
	jdff dff_A_Adf9uIwU5_0(.dout(w_dff_A_Jjl2wtTR6_0),.din(w_dff_A_Adf9uIwU5_0),.clk(gclk));
	jdff dff_A_Jjl2wtTR6_0(.dout(w_dff_A_riKnTTVZ4_0),.din(w_dff_A_Jjl2wtTR6_0),.clk(gclk));
	jdff dff_A_riKnTTVZ4_0(.dout(G492),.din(w_dff_A_riKnTTVZ4_0),.clk(gclk));
	jdff dff_A_3ZgZBMkC9_1(.dout(w_dff_A_IZ5PZk5T1_0),.din(w_dff_A_3ZgZBMkC9_1),.clk(gclk));
	jdff dff_A_IZ5PZk5T1_0(.dout(w_dff_A_KKDlyxGu6_0),.din(w_dff_A_IZ5PZk5T1_0),.clk(gclk));
	jdff dff_A_KKDlyxGu6_0(.dout(w_dff_A_DUJFvNjE8_0),.din(w_dff_A_KKDlyxGu6_0),.clk(gclk));
	jdff dff_A_DUJFvNjE8_0(.dout(w_dff_A_RmTNuhnG8_0),.din(w_dff_A_DUJFvNjE8_0),.clk(gclk));
	jdff dff_A_RmTNuhnG8_0(.dout(w_dff_A_SpJoU5tG4_0),.din(w_dff_A_RmTNuhnG8_0),.clk(gclk));
	jdff dff_A_SpJoU5tG4_0(.dout(w_dff_A_btUjeE8P2_0),.din(w_dff_A_SpJoU5tG4_0),.clk(gclk));
	jdff dff_A_btUjeE8P2_0(.dout(w_dff_A_iOBp8yYX0_0),.din(w_dff_A_btUjeE8P2_0),.clk(gclk));
	jdff dff_A_iOBp8yYX0_0(.dout(w_dff_A_HGBZ4CNf7_0),.din(w_dff_A_iOBp8yYX0_0),.clk(gclk));
	jdff dff_A_HGBZ4CNf7_0(.dout(w_dff_A_4UhJp8bi9_0),.din(w_dff_A_HGBZ4CNf7_0),.clk(gclk));
	jdff dff_A_4UhJp8bi9_0(.dout(w_dff_A_TEl1bOVV8_0),.din(w_dff_A_4UhJp8bi9_0),.clk(gclk));
	jdff dff_A_TEl1bOVV8_0(.dout(w_dff_A_Za8Jvuu72_0),.din(w_dff_A_TEl1bOVV8_0),.clk(gclk));
	jdff dff_A_Za8Jvuu72_0(.dout(w_dff_A_lhHcrvbB1_0),.din(w_dff_A_Za8Jvuu72_0),.clk(gclk));
	jdff dff_A_lhHcrvbB1_0(.dout(w_dff_A_FsEdFg1w7_0),.din(w_dff_A_lhHcrvbB1_0),.clk(gclk));
	jdff dff_A_FsEdFg1w7_0(.dout(w_dff_A_B4UEwavN3_0),.din(w_dff_A_FsEdFg1w7_0),.clk(gclk));
	jdff dff_A_B4UEwavN3_0(.dout(w_dff_A_aFdxKZoe1_0),.din(w_dff_A_B4UEwavN3_0),.clk(gclk));
	jdff dff_A_aFdxKZoe1_0(.dout(w_dff_A_FTyiYmxU8_0),.din(w_dff_A_aFdxKZoe1_0),.clk(gclk));
	jdff dff_A_FTyiYmxU8_0(.dout(w_dff_A_Rk8kZTiQ8_0),.din(w_dff_A_FTyiYmxU8_0),.clk(gclk));
	jdff dff_A_Rk8kZTiQ8_0(.dout(w_dff_A_OqeN6mxq4_0),.din(w_dff_A_Rk8kZTiQ8_0),.clk(gclk));
	jdff dff_A_OqeN6mxq4_0(.dout(w_dff_A_jctkx6nM4_0),.din(w_dff_A_OqeN6mxq4_0),.clk(gclk));
	jdff dff_A_jctkx6nM4_0(.dout(w_dff_A_RUqYA2zh8_0),.din(w_dff_A_jctkx6nM4_0),.clk(gclk));
	jdff dff_A_RUqYA2zh8_0(.dout(w_dff_A_lqltRERL4_0),.din(w_dff_A_RUqYA2zh8_0),.clk(gclk));
	jdff dff_A_lqltRERL4_0(.dout(w_dff_A_GLEcxDyd1_0),.din(w_dff_A_lqltRERL4_0),.clk(gclk));
	jdff dff_A_GLEcxDyd1_0(.dout(w_dff_A_kDxnzNc71_0),.din(w_dff_A_GLEcxDyd1_0),.clk(gclk));
	jdff dff_A_kDxnzNc71_0(.dout(w_dff_A_biqjCc5w0_0),.din(w_dff_A_kDxnzNc71_0),.clk(gclk));
	jdff dff_A_biqjCc5w0_0(.dout(w_dff_A_Po3bXLZ27_0),.din(w_dff_A_biqjCc5w0_0),.clk(gclk));
	jdff dff_A_Po3bXLZ27_0(.dout(w_dff_A_NP0CdFxh6_0),.din(w_dff_A_Po3bXLZ27_0),.clk(gclk));
	jdff dff_A_NP0CdFxh6_0(.dout(G490),.din(w_dff_A_NP0CdFxh6_0),.clk(gclk));
	jdff dff_A_inOpBq5G8_1(.dout(w_dff_A_039U8Q8C1_0),.din(w_dff_A_inOpBq5G8_1),.clk(gclk));
	jdff dff_A_039U8Q8C1_0(.dout(w_dff_A_PTp0ta9f6_0),.din(w_dff_A_039U8Q8C1_0),.clk(gclk));
	jdff dff_A_PTp0ta9f6_0(.dout(w_dff_A_g708R9XT0_0),.din(w_dff_A_PTp0ta9f6_0),.clk(gclk));
	jdff dff_A_g708R9XT0_0(.dout(w_dff_A_t3Yp2unN1_0),.din(w_dff_A_g708R9XT0_0),.clk(gclk));
	jdff dff_A_t3Yp2unN1_0(.dout(w_dff_A_OXpDVo2H8_0),.din(w_dff_A_t3Yp2unN1_0),.clk(gclk));
	jdff dff_A_OXpDVo2H8_0(.dout(w_dff_A_sSmWuDKB1_0),.din(w_dff_A_OXpDVo2H8_0),.clk(gclk));
	jdff dff_A_sSmWuDKB1_0(.dout(w_dff_A_UKCzLuto4_0),.din(w_dff_A_sSmWuDKB1_0),.clk(gclk));
	jdff dff_A_UKCzLuto4_0(.dout(w_dff_A_NXv5T3ya3_0),.din(w_dff_A_UKCzLuto4_0),.clk(gclk));
	jdff dff_A_NXv5T3ya3_0(.dout(w_dff_A_CAUnL9Al1_0),.din(w_dff_A_NXv5T3ya3_0),.clk(gclk));
	jdff dff_A_CAUnL9Al1_0(.dout(w_dff_A_cIcFij5p5_0),.din(w_dff_A_CAUnL9Al1_0),.clk(gclk));
	jdff dff_A_cIcFij5p5_0(.dout(w_dff_A_Ilymf3k60_0),.din(w_dff_A_cIcFij5p5_0),.clk(gclk));
	jdff dff_A_Ilymf3k60_0(.dout(w_dff_A_8qrfBtfI6_0),.din(w_dff_A_Ilymf3k60_0),.clk(gclk));
	jdff dff_A_8qrfBtfI6_0(.dout(w_dff_A_6SJqKCvb9_0),.din(w_dff_A_8qrfBtfI6_0),.clk(gclk));
	jdff dff_A_6SJqKCvb9_0(.dout(w_dff_A_3m0wo6jv8_0),.din(w_dff_A_6SJqKCvb9_0),.clk(gclk));
	jdff dff_A_3m0wo6jv8_0(.dout(w_dff_A_yOuD4OE66_0),.din(w_dff_A_3m0wo6jv8_0),.clk(gclk));
	jdff dff_A_yOuD4OE66_0(.dout(w_dff_A_TNs3vqNj5_0),.din(w_dff_A_yOuD4OE66_0),.clk(gclk));
	jdff dff_A_TNs3vqNj5_0(.dout(w_dff_A_LZCfvpDu8_0),.din(w_dff_A_TNs3vqNj5_0),.clk(gclk));
	jdff dff_A_LZCfvpDu8_0(.dout(w_dff_A_pSsy8Hzz1_0),.din(w_dff_A_LZCfvpDu8_0),.clk(gclk));
	jdff dff_A_pSsy8Hzz1_0(.dout(w_dff_A_V89V8Nw91_0),.din(w_dff_A_pSsy8Hzz1_0),.clk(gclk));
	jdff dff_A_V89V8Nw91_0(.dout(w_dff_A_zqLwOlIH9_0),.din(w_dff_A_V89V8Nw91_0),.clk(gclk));
	jdff dff_A_zqLwOlIH9_0(.dout(w_dff_A_PXP0deGy6_0),.din(w_dff_A_zqLwOlIH9_0),.clk(gclk));
	jdff dff_A_PXP0deGy6_0(.dout(w_dff_A_yf5cjXBT9_0),.din(w_dff_A_PXP0deGy6_0),.clk(gclk));
	jdff dff_A_yf5cjXBT9_0(.dout(w_dff_A_TLyJCJ7a6_0),.din(w_dff_A_yf5cjXBT9_0),.clk(gclk));
	jdff dff_A_TLyJCJ7a6_0(.dout(w_dff_A_dMl85Xx90_0),.din(w_dff_A_TLyJCJ7a6_0),.clk(gclk));
	jdff dff_A_dMl85Xx90_0(.dout(w_dff_A_8ghSo01x1_0),.din(w_dff_A_dMl85Xx90_0),.clk(gclk));
	jdff dff_A_8ghSo01x1_0(.dout(w_dff_A_BAVH7tD56_0),.din(w_dff_A_8ghSo01x1_0),.clk(gclk));
	jdff dff_A_BAVH7tD56_0(.dout(G488),.din(w_dff_A_BAVH7tD56_0),.clk(gclk));
	jdff dff_A_hlARsFhN7_1(.dout(w_dff_A_SgpPuK3k2_0),.din(w_dff_A_hlARsFhN7_1),.clk(gclk));
	jdff dff_A_SgpPuK3k2_0(.dout(w_dff_A_kIS6r4aZ7_0),.din(w_dff_A_SgpPuK3k2_0),.clk(gclk));
	jdff dff_A_kIS6r4aZ7_0(.dout(w_dff_A_j1uevwda9_0),.din(w_dff_A_kIS6r4aZ7_0),.clk(gclk));
	jdff dff_A_j1uevwda9_0(.dout(w_dff_A_ulUrA0lV6_0),.din(w_dff_A_j1uevwda9_0),.clk(gclk));
	jdff dff_A_ulUrA0lV6_0(.dout(w_dff_A_4DfMWjq31_0),.din(w_dff_A_ulUrA0lV6_0),.clk(gclk));
	jdff dff_A_4DfMWjq31_0(.dout(w_dff_A_OuPm1V7O1_0),.din(w_dff_A_4DfMWjq31_0),.clk(gclk));
	jdff dff_A_OuPm1V7O1_0(.dout(w_dff_A_RBfYFazA8_0),.din(w_dff_A_OuPm1V7O1_0),.clk(gclk));
	jdff dff_A_RBfYFazA8_0(.dout(w_dff_A_akxtPTHv4_0),.din(w_dff_A_RBfYFazA8_0),.clk(gclk));
	jdff dff_A_akxtPTHv4_0(.dout(w_dff_A_m4lMHFXj6_0),.din(w_dff_A_akxtPTHv4_0),.clk(gclk));
	jdff dff_A_m4lMHFXj6_0(.dout(w_dff_A_dmLDFLKy4_0),.din(w_dff_A_m4lMHFXj6_0),.clk(gclk));
	jdff dff_A_dmLDFLKy4_0(.dout(w_dff_A_CXZm86Ph2_0),.din(w_dff_A_dmLDFLKy4_0),.clk(gclk));
	jdff dff_A_CXZm86Ph2_0(.dout(w_dff_A_wNhqRwne3_0),.din(w_dff_A_CXZm86Ph2_0),.clk(gclk));
	jdff dff_A_wNhqRwne3_0(.dout(w_dff_A_CoksQ7oJ2_0),.din(w_dff_A_wNhqRwne3_0),.clk(gclk));
	jdff dff_A_CoksQ7oJ2_0(.dout(w_dff_A_EHcs4mm87_0),.din(w_dff_A_CoksQ7oJ2_0),.clk(gclk));
	jdff dff_A_EHcs4mm87_0(.dout(w_dff_A_d0FflE2i1_0),.din(w_dff_A_EHcs4mm87_0),.clk(gclk));
	jdff dff_A_d0FflE2i1_0(.dout(w_dff_A_osMKI9VY2_0),.din(w_dff_A_d0FflE2i1_0),.clk(gclk));
	jdff dff_A_osMKI9VY2_0(.dout(w_dff_A_ZsRbECSD5_0),.din(w_dff_A_osMKI9VY2_0),.clk(gclk));
	jdff dff_A_ZsRbECSD5_0(.dout(w_dff_A_srEJcsCX5_0),.din(w_dff_A_ZsRbECSD5_0),.clk(gclk));
	jdff dff_A_srEJcsCX5_0(.dout(w_dff_A_bA9m6G8e2_0),.din(w_dff_A_srEJcsCX5_0),.clk(gclk));
	jdff dff_A_bA9m6G8e2_0(.dout(w_dff_A_3vMVWMoP0_0),.din(w_dff_A_bA9m6G8e2_0),.clk(gclk));
	jdff dff_A_3vMVWMoP0_0(.dout(w_dff_A_vU82p77L9_0),.din(w_dff_A_3vMVWMoP0_0),.clk(gclk));
	jdff dff_A_vU82p77L9_0(.dout(w_dff_A_WY6hktmd5_0),.din(w_dff_A_vU82p77L9_0),.clk(gclk));
	jdff dff_A_WY6hktmd5_0(.dout(w_dff_A_LN2CD0su7_0),.din(w_dff_A_WY6hktmd5_0),.clk(gclk));
	jdff dff_A_LN2CD0su7_0(.dout(w_dff_A_173W7EVh5_0),.din(w_dff_A_LN2CD0su7_0),.clk(gclk));
	jdff dff_A_173W7EVh5_0(.dout(w_dff_A_zgz1NpSK5_0),.din(w_dff_A_173W7EVh5_0),.clk(gclk));
	jdff dff_A_zgz1NpSK5_0(.dout(w_dff_A_zcFDXErM4_0),.din(w_dff_A_zgz1NpSK5_0),.clk(gclk));
	jdff dff_A_zcFDXErM4_0(.dout(G486),.din(w_dff_A_zcFDXErM4_0),.clk(gclk));
	jdff dff_A_Yw7VDQLa0_1(.dout(w_dff_A_fFw0wmn91_0),.din(w_dff_A_Yw7VDQLa0_1),.clk(gclk));
	jdff dff_A_fFw0wmn91_0(.dout(w_dff_A_lJ6ZBqqG7_0),.din(w_dff_A_fFw0wmn91_0),.clk(gclk));
	jdff dff_A_lJ6ZBqqG7_0(.dout(w_dff_A_kvUmlWvO0_0),.din(w_dff_A_lJ6ZBqqG7_0),.clk(gclk));
	jdff dff_A_kvUmlWvO0_0(.dout(w_dff_A_2hff1qmi7_0),.din(w_dff_A_kvUmlWvO0_0),.clk(gclk));
	jdff dff_A_2hff1qmi7_0(.dout(w_dff_A_xvfhuQGx0_0),.din(w_dff_A_2hff1qmi7_0),.clk(gclk));
	jdff dff_A_xvfhuQGx0_0(.dout(w_dff_A_wIoYfbUU9_0),.din(w_dff_A_xvfhuQGx0_0),.clk(gclk));
	jdff dff_A_wIoYfbUU9_0(.dout(w_dff_A_BZdaZaar2_0),.din(w_dff_A_wIoYfbUU9_0),.clk(gclk));
	jdff dff_A_BZdaZaar2_0(.dout(w_dff_A_6EWU5u2h8_0),.din(w_dff_A_BZdaZaar2_0),.clk(gclk));
	jdff dff_A_6EWU5u2h8_0(.dout(w_dff_A_cFMAwVlX6_0),.din(w_dff_A_6EWU5u2h8_0),.clk(gclk));
	jdff dff_A_cFMAwVlX6_0(.dout(w_dff_A_kA0hsreO0_0),.din(w_dff_A_cFMAwVlX6_0),.clk(gclk));
	jdff dff_A_kA0hsreO0_0(.dout(w_dff_A_eA4MY8kK1_0),.din(w_dff_A_kA0hsreO0_0),.clk(gclk));
	jdff dff_A_eA4MY8kK1_0(.dout(w_dff_A_sO5rbTRb9_0),.din(w_dff_A_eA4MY8kK1_0),.clk(gclk));
	jdff dff_A_sO5rbTRb9_0(.dout(w_dff_A_dciytgMa1_0),.din(w_dff_A_sO5rbTRb9_0),.clk(gclk));
	jdff dff_A_dciytgMa1_0(.dout(w_dff_A_58Xol0Np8_0),.din(w_dff_A_dciytgMa1_0),.clk(gclk));
	jdff dff_A_58Xol0Np8_0(.dout(w_dff_A_NIDDf4Uc5_0),.din(w_dff_A_58Xol0Np8_0),.clk(gclk));
	jdff dff_A_NIDDf4Uc5_0(.dout(w_dff_A_arZCFY215_0),.din(w_dff_A_NIDDf4Uc5_0),.clk(gclk));
	jdff dff_A_arZCFY215_0(.dout(w_dff_A_sOaTfcIY3_0),.din(w_dff_A_arZCFY215_0),.clk(gclk));
	jdff dff_A_sOaTfcIY3_0(.dout(w_dff_A_qnPdfFKy6_0),.din(w_dff_A_sOaTfcIY3_0),.clk(gclk));
	jdff dff_A_qnPdfFKy6_0(.dout(w_dff_A_xFVdJ6F87_0),.din(w_dff_A_qnPdfFKy6_0),.clk(gclk));
	jdff dff_A_xFVdJ6F87_0(.dout(w_dff_A_pAjtyoiV0_0),.din(w_dff_A_xFVdJ6F87_0),.clk(gclk));
	jdff dff_A_pAjtyoiV0_0(.dout(w_dff_A_l4uHRBEq2_0),.din(w_dff_A_pAjtyoiV0_0),.clk(gclk));
	jdff dff_A_l4uHRBEq2_0(.dout(w_dff_A_eNfHrf2X2_0),.din(w_dff_A_l4uHRBEq2_0),.clk(gclk));
	jdff dff_A_eNfHrf2X2_0(.dout(w_dff_A_DAxIzlkR2_0),.din(w_dff_A_eNfHrf2X2_0),.clk(gclk));
	jdff dff_A_DAxIzlkR2_0(.dout(w_dff_A_FUjRZ8cJ9_0),.din(w_dff_A_DAxIzlkR2_0),.clk(gclk));
	jdff dff_A_FUjRZ8cJ9_0(.dout(w_dff_A_m8DC2qn42_0),.din(w_dff_A_FUjRZ8cJ9_0),.clk(gclk));
	jdff dff_A_m8DC2qn42_0(.dout(w_dff_A_z06FxRP62_0),.din(w_dff_A_m8DC2qn42_0),.clk(gclk));
	jdff dff_A_z06FxRP62_0(.dout(G484),.din(w_dff_A_z06FxRP62_0),.clk(gclk));
	jdff dff_A_iwHRIdkG4_1(.dout(w_dff_A_BGIFbOyj3_0),.din(w_dff_A_iwHRIdkG4_1),.clk(gclk));
	jdff dff_A_BGIFbOyj3_0(.dout(w_dff_A_shiOtPBA1_0),.din(w_dff_A_BGIFbOyj3_0),.clk(gclk));
	jdff dff_A_shiOtPBA1_0(.dout(w_dff_A_yQ1frlMq0_0),.din(w_dff_A_shiOtPBA1_0),.clk(gclk));
	jdff dff_A_yQ1frlMq0_0(.dout(w_dff_A_QjrkGQnj0_0),.din(w_dff_A_yQ1frlMq0_0),.clk(gclk));
	jdff dff_A_QjrkGQnj0_0(.dout(w_dff_A_VjBlEaz29_0),.din(w_dff_A_QjrkGQnj0_0),.clk(gclk));
	jdff dff_A_VjBlEaz29_0(.dout(w_dff_A_XKRGadRE7_0),.din(w_dff_A_VjBlEaz29_0),.clk(gclk));
	jdff dff_A_XKRGadRE7_0(.dout(w_dff_A_PuRnX3BE1_0),.din(w_dff_A_XKRGadRE7_0),.clk(gclk));
	jdff dff_A_PuRnX3BE1_0(.dout(w_dff_A_TpKsZdyo3_0),.din(w_dff_A_PuRnX3BE1_0),.clk(gclk));
	jdff dff_A_TpKsZdyo3_0(.dout(w_dff_A_hNASR3aM1_0),.din(w_dff_A_TpKsZdyo3_0),.clk(gclk));
	jdff dff_A_hNASR3aM1_0(.dout(w_dff_A_VgJ6n0pj0_0),.din(w_dff_A_hNASR3aM1_0),.clk(gclk));
	jdff dff_A_VgJ6n0pj0_0(.dout(w_dff_A_6ho07pFh3_0),.din(w_dff_A_VgJ6n0pj0_0),.clk(gclk));
	jdff dff_A_6ho07pFh3_0(.dout(w_dff_A_3jgQ4y4P6_0),.din(w_dff_A_6ho07pFh3_0),.clk(gclk));
	jdff dff_A_3jgQ4y4P6_0(.dout(w_dff_A_4yPJU22y0_0),.din(w_dff_A_3jgQ4y4P6_0),.clk(gclk));
	jdff dff_A_4yPJU22y0_0(.dout(w_dff_A_tR7DVRlK5_0),.din(w_dff_A_4yPJU22y0_0),.clk(gclk));
	jdff dff_A_tR7DVRlK5_0(.dout(w_dff_A_VCW5Ns853_0),.din(w_dff_A_tR7DVRlK5_0),.clk(gclk));
	jdff dff_A_VCW5Ns853_0(.dout(w_dff_A_z1DAj4V71_0),.din(w_dff_A_VCW5Ns853_0),.clk(gclk));
	jdff dff_A_z1DAj4V71_0(.dout(w_dff_A_7taAytV31_0),.din(w_dff_A_z1DAj4V71_0),.clk(gclk));
	jdff dff_A_7taAytV31_0(.dout(w_dff_A_SriZSmBP0_0),.din(w_dff_A_7taAytV31_0),.clk(gclk));
	jdff dff_A_SriZSmBP0_0(.dout(w_dff_A_1Jb8n4hz9_0),.din(w_dff_A_SriZSmBP0_0),.clk(gclk));
	jdff dff_A_1Jb8n4hz9_0(.dout(w_dff_A_1Xt1UsRl3_0),.din(w_dff_A_1Jb8n4hz9_0),.clk(gclk));
	jdff dff_A_1Xt1UsRl3_0(.dout(w_dff_A_intqS4js7_0),.din(w_dff_A_1Xt1UsRl3_0),.clk(gclk));
	jdff dff_A_intqS4js7_0(.dout(w_dff_A_k5KwYpQi1_0),.din(w_dff_A_intqS4js7_0),.clk(gclk));
	jdff dff_A_k5KwYpQi1_0(.dout(w_dff_A_gmh3UkLG7_0),.din(w_dff_A_k5KwYpQi1_0),.clk(gclk));
	jdff dff_A_gmh3UkLG7_0(.dout(w_dff_A_ppx1SayD0_0),.din(w_dff_A_gmh3UkLG7_0),.clk(gclk));
	jdff dff_A_ppx1SayD0_0(.dout(w_dff_A_elGRqeP33_0),.din(w_dff_A_ppx1SayD0_0),.clk(gclk));
	jdff dff_A_elGRqeP33_0(.dout(w_dff_A_De9jW90n8_0),.din(w_dff_A_elGRqeP33_0),.clk(gclk));
	jdff dff_A_De9jW90n8_0(.dout(G482),.din(w_dff_A_De9jW90n8_0),.clk(gclk));
	jdff dff_A_C0nNn7ci4_1(.dout(w_dff_A_kUPu9xz88_0),.din(w_dff_A_C0nNn7ci4_1),.clk(gclk));
	jdff dff_A_kUPu9xz88_0(.dout(w_dff_A_nTUQs7fh3_0),.din(w_dff_A_kUPu9xz88_0),.clk(gclk));
	jdff dff_A_nTUQs7fh3_0(.dout(w_dff_A_menA27iF4_0),.din(w_dff_A_nTUQs7fh3_0),.clk(gclk));
	jdff dff_A_menA27iF4_0(.dout(w_dff_A_Rcnqp6fB2_0),.din(w_dff_A_menA27iF4_0),.clk(gclk));
	jdff dff_A_Rcnqp6fB2_0(.dout(w_dff_A_ztQaC30v6_0),.din(w_dff_A_Rcnqp6fB2_0),.clk(gclk));
	jdff dff_A_ztQaC30v6_0(.dout(w_dff_A_PyRfqxRy5_0),.din(w_dff_A_ztQaC30v6_0),.clk(gclk));
	jdff dff_A_PyRfqxRy5_0(.dout(w_dff_A_Na6L0eqI3_0),.din(w_dff_A_PyRfqxRy5_0),.clk(gclk));
	jdff dff_A_Na6L0eqI3_0(.dout(w_dff_A_YUikfB001_0),.din(w_dff_A_Na6L0eqI3_0),.clk(gclk));
	jdff dff_A_YUikfB001_0(.dout(w_dff_A_wIpC1jAw5_0),.din(w_dff_A_YUikfB001_0),.clk(gclk));
	jdff dff_A_wIpC1jAw5_0(.dout(w_dff_A_iL6rTm147_0),.din(w_dff_A_wIpC1jAw5_0),.clk(gclk));
	jdff dff_A_iL6rTm147_0(.dout(w_dff_A_RG42v5Fo8_0),.din(w_dff_A_iL6rTm147_0),.clk(gclk));
	jdff dff_A_RG42v5Fo8_0(.dout(w_dff_A_sPq86jLW4_0),.din(w_dff_A_RG42v5Fo8_0),.clk(gclk));
	jdff dff_A_sPq86jLW4_0(.dout(w_dff_A_YHmzYt8i1_0),.din(w_dff_A_sPq86jLW4_0),.clk(gclk));
	jdff dff_A_YHmzYt8i1_0(.dout(w_dff_A_4OxsawFZ3_0),.din(w_dff_A_YHmzYt8i1_0),.clk(gclk));
	jdff dff_A_4OxsawFZ3_0(.dout(w_dff_A_JnSSaOBu9_0),.din(w_dff_A_4OxsawFZ3_0),.clk(gclk));
	jdff dff_A_JnSSaOBu9_0(.dout(w_dff_A_kRPMbu3g4_0),.din(w_dff_A_JnSSaOBu9_0),.clk(gclk));
	jdff dff_A_kRPMbu3g4_0(.dout(w_dff_A_HUWUs3gN8_0),.din(w_dff_A_kRPMbu3g4_0),.clk(gclk));
	jdff dff_A_HUWUs3gN8_0(.dout(w_dff_A_OUZKb1xo5_0),.din(w_dff_A_HUWUs3gN8_0),.clk(gclk));
	jdff dff_A_OUZKb1xo5_0(.dout(w_dff_A_9e2NgsCI6_0),.din(w_dff_A_OUZKb1xo5_0),.clk(gclk));
	jdff dff_A_9e2NgsCI6_0(.dout(w_dff_A_FsJOpsmq4_0),.din(w_dff_A_9e2NgsCI6_0),.clk(gclk));
	jdff dff_A_FsJOpsmq4_0(.dout(w_dff_A_C1xQKPcp3_0),.din(w_dff_A_FsJOpsmq4_0),.clk(gclk));
	jdff dff_A_C1xQKPcp3_0(.dout(w_dff_A_SfHDnweU7_0),.din(w_dff_A_C1xQKPcp3_0),.clk(gclk));
	jdff dff_A_SfHDnweU7_0(.dout(w_dff_A_U4Ve1heT3_0),.din(w_dff_A_SfHDnweU7_0),.clk(gclk));
	jdff dff_A_U4Ve1heT3_0(.dout(w_dff_A_Mx8z8elo3_0),.din(w_dff_A_U4Ve1heT3_0),.clk(gclk));
	jdff dff_A_Mx8z8elo3_0(.dout(w_dff_A_gUPOrKao8_0),.din(w_dff_A_Mx8z8elo3_0),.clk(gclk));
	jdff dff_A_gUPOrKao8_0(.dout(w_dff_A_Jwe6IFZW0_0),.din(w_dff_A_gUPOrKao8_0),.clk(gclk));
	jdff dff_A_Jwe6IFZW0_0(.dout(G480),.din(w_dff_A_Jwe6IFZW0_0),.clk(gclk));
	jdff dff_A_d6GEvmtG3_1(.dout(w_dff_A_jatncqTv3_0),.din(w_dff_A_d6GEvmtG3_1),.clk(gclk));
	jdff dff_A_jatncqTv3_0(.dout(w_dff_A_ZKRR7VyO6_0),.din(w_dff_A_jatncqTv3_0),.clk(gclk));
	jdff dff_A_ZKRR7VyO6_0(.dout(w_dff_A_Dws1yAcj2_0),.din(w_dff_A_ZKRR7VyO6_0),.clk(gclk));
	jdff dff_A_Dws1yAcj2_0(.dout(w_dff_A_I4b9DIGF2_0),.din(w_dff_A_Dws1yAcj2_0),.clk(gclk));
	jdff dff_A_I4b9DIGF2_0(.dout(w_dff_A_Rx6S3XMy1_0),.din(w_dff_A_I4b9DIGF2_0),.clk(gclk));
	jdff dff_A_Rx6S3XMy1_0(.dout(w_dff_A_4IaJ9Jsx0_0),.din(w_dff_A_Rx6S3XMy1_0),.clk(gclk));
	jdff dff_A_4IaJ9Jsx0_0(.dout(w_dff_A_a2yzrX7B0_0),.din(w_dff_A_4IaJ9Jsx0_0),.clk(gclk));
	jdff dff_A_a2yzrX7B0_0(.dout(w_dff_A_MOLNygZT2_0),.din(w_dff_A_a2yzrX7B0_0),.clk(gclk));
	jdff dff_A_MOLNygZT2_0(.dout(w_dff_A_6ruPEoHw7_0),.din(w_dff_A_MOLNygZT2_0),.clk(gclk));
	jdff dff_A_6ruPEoHw7_0(.dout(w_dff_A_74PywZLp3_0),.din(w_dff_A_6ruPEoHw7_0),.clk(gclk));
	jdff dff_A_74PywZLp3_0(.dout(w_dff_A_cLjHBqcF3_0),.din(w_dff_A_74PywZLp3_0),.clk(gclk));
	jdff dff_A_cLjHBqcF3_0(.dout(w_dff_A_bvywiqoq9_0),.din(w_dff_A_cLjHBqcF3_0),.clk(gclk));
	jdff dff_A_bvywiqoq9_0(.dout(w_dff_A_lujqbKWz4_0),.din(w_dff_A_bvywiqoq9_0),.clk(gclk));
	jdff dff_A_lujqbKWz4_0(.dout(w_dff_A_CD3PBN9n0_0),.din(w_dff_A_lujqbKWz4_0),.clk(gclk));
	jdff dff_A_CD3PBN9n0_0(.dout(w_dff_A_7PYJo2uh6_0),.din(w_dff_A_CD3PBN9n0_0),.clk(gclk));
	jdff dff_A_7PYJo2uh6_0(.dout(w_dff_A_X0UhJiYk1_0),.din(w_dff_A_7PYJo2uh6_0),.clk(gclk));
	jdff dff_A_X0UhJiYk1_0(.dout(w_dff_A_aRRRFv0Y8_0),.din(w_dff_A_X0UhJiYk1_0),.clk(gclk));
	jdff dff_A_aRRRFv0Y8_0(.dout(w_dff_A_FGG79RbH4_0),.din(w_dff_A_aRRRFv0Y8_0),.clk(gclk));
	jdff dff_A_FGG79RbH4_0(.dout(w_dff_A_7YPD08pT7_0),.din(w_dff_A_FGG79RbH4_0),.clk(gclk));
	jdff dff_A_7YPD08pT7_0(.dout(w_dff_A_YdEAceCT3_0),.din(w_dff_A_7YPD08pT7_0),.clk(gclk));
	jdff dff_A_YdEAceCT3_0(.dout(w_dff_A_Zuj8yi9w9_0),.din(w_dff_A_YdEAceCT3_0),.clk(gclk));
	jdff dff_A_Zuj8yi9w9_0(.dout(w_dff_A_VbVlLpp90_0),.din(w_dff_A_Zuj8yi9w9_0),.clk(gclk));
	jdff dff_A_VbVlLpp90_0(.dout(w_dff_A_TSdVQWS17_0),.din(w_dff_A_VbVlLpp90_0),.clk(gclk));
	jdff dff_A_TSdVQWS17_0(.dout(w_dff_A_RSBOxWA59_0),.din(w_dff_A_TSdVQWS17_0),.clk(gclk));
	jdff dff_A_RSBOxWA59_0(.dout(w_dff_A_i1Oq1Gay7_0),.din(w_dff_A_RSBOxWA59_0),.clk(gclk));
	jdff dff_A_i1Oq1Gay7_0(.dout(w_dff_A_yMBFHVXl3_0),.din(w_dff_A_i1Oq1Gay7_0),.clk(gclk));
	jdff dff_A_yMBFHVXl3_0(.dout(G560),.din(w_dff_A_yMBFHVXl3_0),.clk(gclk));
	jdff dff_A_0Uka2LbP9_1(.dout(w_dff_A_U360T9CC3_0),.din(w_dff_A_0Uka2LbP9_1),.clk(gclk));
	jdff dff_A_U360T9CC3_0(.dout(w_dff_A_wPxsm4iK0_0),.din(w_dff_A_U360T9CC3_0),.clk(gclk));
	jdff dff_A_wPxsm4iK0_0(.dout(w_dff_A_Kg8I0Y0n2_0),.din(w_dff_A_wPxsm4iK0_0),.clk(gclk));
	jdff dff_A_Kg8I0Y0n2_0(.dout(w_dff_A_0j38edxy7_0),.din(w_dff_A_Kg8I0Y0n2_0),.clk(gclk));
	jdff dff_A_0j38edxy7_0(.dout(w_dff_A_2Y5icIgb2_0),.din(w_dff_A_0j38edxy7_0),.clk(gclk));
	jdff dff_A_2Y5icIgb2_0(.dout(w_dff_A_dbHfyyK58_0),.din(w_dff_A_2Y5icIgb2_0),.clk(gclk));
	jdff dff_A_dbHfyyK58_0(.dout(w_dff_A_XZOwo9XQ9_0),.din(w_dff_A_dbHfyyK58_0),.clk(gclk));
	jdff dff_A_XZOwo9XQ9_0(.dout(w_dff_A_gLWV1RHN1_0),.din(w_dff_A_XZOwo9XQ9_0),.clk(gclk));
	jdff dff_A_gLWV1RHN1_0(.dout(w_dff_A_MH5HzhXf2_0),.din(w_dff_A_gLWV1RHN1_0),.clk(gclk));
	jdff dff_A_MH5HzhXf2_0(.dout(w_dff_A_PwtvLxwV8_0),.din(w_dff_A_MH5HzhXf2_0),.clk(gclk));
	jdff dff_A_PwtvLxwV8_0(.dout(w_dff_A_EzDjUDpC9_0),.din(w_dff_A_PwtvLxwV8_0),.clk(gclk));
	jdff dff_A_EzDjUDpC9_0(.dout(w_dff_A_XhltOiFl0_0),.din(w_dff_A_EzDjUDpC9_0),.clk(gclk));
	jdff dff_A_XhltOiFl0_0(.dout(w_dff_A_luhPqDeG9_0),.din(w_dff_A_XhltOiFl0_0),.clk(gclk));
	jdff dff_A_luhPqDeG9_0(.dout(w_dff_A_LEEInI1R5_0),.din(w_dff_A_luhPqDeG9_0),.clk(gclk));
	jdff dff_A_LEEInI1R5_0(.dout(w_dff_A_FRn12GRG9_0),.din(w_dff_A_LEEInI1R5_0),.clk(gclk));
	jdff dff_A_FRn12GRG9_0(.dout(w_dff_A_g0GJsn7h6_0),.din(w_dff_A_FRn12GRG9_0),.clk(gclk));
	jdff dff_A_g0GJsn7h6_0(.dout(w_dff_A_3pNBqtwD8_0),.din(w_dff_A_g0GJsn7h6_0),.clk(gclk));
	jdff dff_A_3pNBqtwD8_0(.dout(w_dff_A_zxtyWdo04_0),.din(w_dff_A_3pNBqtwD8_0),.clk(gclk));
	jdff dff_A_zxtyWdo04_0(.dout(w_dff_A_VrctfqQd1_0),.din(w_dff_A_zxtyWdo04_0),.clk(gclk));
	jdff dff_A_VrctfqQd1_0(.dout(w_dff_A_99TJh3EW7_0),.din(w_dff_A_VrctfqQd1_0),.clk(gclk));
	jdff dff_A_99TJh3EW7_0(.dout(w_dff_A_JqdtJ06t7_0),.din(w_dff_A_99TJh3EW7_0),.clk(gclk));
	jdff dff_A_JqdtJ06t7_0(.dout(w_dff_A_KtDeLRLl3_0),.din(w_dff_A_JqdtJ06t7_0),.clk(gclk));
	jdff dff_A_KtDeLRLl3_0(.dout(w_dff_A_EN5A6FlR1_0),.din(w_dff_A_KtDeLRLl3_0),.clk(gclk));
	jdff dff_A_EN5A6FlR1_0(.dout(w_dff_A_ygNdqXwl1_0),.din(w_dff_A_EN5A6FlR1_0),.clk(gclk));
	jdff dff_A_ygNdqXwl1_0(.dout(w_dff_A_wMvJbbhA8_0),.din(w_dff_A_ygNdqXwl1_0),.clk(gclk));
	jdff dff_A_wMvJbbhA8_0(.dout(w_dff_A_Ttx6l0hr3_0),.din(w_dff_A_wMvJbbhA8_0),.clk(gclk));
	jdff dff_A_Ttx6l0hr3_0(.dout(G542),.din(w_dff_A_Ttx6l0hr3_0),.clk(gclk));
	jdff dff_A_KehafRC34_1(.dout(w_dff_A_RKitj7TC4_0),.din(w_dff_A_KehafRC34_1),.clk(gclk));
	jdff dff_A_RKitj7TC4_0(.dout(w_dff_A_v5Hpp9362_0),.din(w_dff_A_RKitj7TC4_0),.clk(gclk));
	jdff dff_A_v5Hpp9362_0(.dout(w_dff_A_DHkfGjeT7_0),.din(w_dff_A_v5Hpp9362_0),.clk(gclk));
	jdff dff_A_DHkfGjeT7_0(.dout(w_dff_A_hclh5f0J6_0),.din(w_dff_A_DHkfGjeT7_0),.clk(gclk));
	jdff dff_A_hclh5f0J6_0(.dout(w_dff_A_6b1ZyCH95_0),.din(w_dff_A_hclh5f0J6_0),.clk(gclk));
	jdff dff_A_6b1ZyCH95_0(.dout(w_dff_A_M9861Nx87_0),.din(w_dff_A_6b1ZyCH95_0),.clk(gclk));
	jdff dff_A_M9861Nx87_0(.dout(w_dff_A_A6i65Hbv0_0),.din(w_dff_A_M9861Nx87_0),.clk(gclk));
	jdff dff_A_A6i65Hbv0_0(.dout(w_dff_A_26sdpdJF5_0),.din(w_dff_A_A6i65Hbv0_0),.clk(gclk));
	jdff dff_A_26sdpdJF5_0(.dout(w_dff_A_8cjHCRR13_0),.din(w_dff_A_26sdpdJF5_0),.clk(gclk));
	jdff dff_A_8cjHCRR13_0(.dout(w_dff_A_4JaGGGtg0_0),.din(w_dff_A_8cjHCRR13_0),.clk(gclk));
	jdff dff_A_4JaGGGtg0_0(.dout(w_dff_A_KtwEtyOQ1_0),.din(w_dff_A_4JaGGGtg0_0),.clk(gclk));
	jdff dff_A_KtwEtyOQ1_0(.dout(w_dff_A_jNqpDRry8_0),.din(w_dff_A_KtwEtyOQ1_0),.clk(gclk));
	jdff dff_A_jNqpDRry8_0(.dout(w_dff_A_W14SfSac1_0),.din(w_dff_A_jNqpDRry8_0),.clk(gclk));
	jdff dff_A_W14SfSac1_0(.dout(w_dff_A_Hhz4z6hb4_0),.din(w_dff_A_W14SfSac1_0),.clk(gclk));
	jdff dff_A_Hhz4z6hb4_0(.dout(w_dff_A_FSunHFIz8_0),.din(w_dff_A_Hhz4z6hb4_0),.clk(gclk));
	jdff dff_A_FSunHFIz8_0(.dout(w_dff_A_6bmdJBYy1_0),.din(w_dff_A_FSunHFIz8_0),.clk(gclk));
	jdff dff_A_6bmdJBYy1_0(.dout(w_dff_A_tL5K89xr9_0),.din(w_dff_A_6bmdJBYy1_0),.clk(gclk));
	jdff dff_A_tL5K89xr9_0(.dout(w_dff_A_m8gXDkFb9_0),.din(w_dff_A_tL5K89xr9_0),.clk(gclk));
	jdff dff_A_m8gXDkFb9_0(.dout(w_dff_A_2cBFxj3S9_0),.din(w_dff_A_m8gXDkFb9_0),.clk(gclk));
	jdff dff_A_2cBFxj3S9_0(.dout(w_dff_A_32Jp2cwV4_0),.din(w_dff_A_2cBFxj3S9_0),.clk(gclk));
	jdff dff_A_32Jp2cwV4_0(.dout(w_dff_A_Dq4fH5Wd0_0),.din(w_dff_A_32Jp2cwV4_0),.clk(gclk));
	jdff dff_A_Dq4fH5Wd0_0(.dout(w_dff_A_E7cqtWc16_0),.din(w_dff_A_Dq4fH5Wd0_0),.clk(gclk));
	jdff dff_A_E7cqtWc16_0(.dout(w_dff_A_nNxW80mH2_0),.din(w_dff_A_E7cqtWc16_0),.clk(gclk));
	jdff dff_A_nNxW80mH2_0(.dout(w_dff_A_9TjaYfXT7_0),.din(w_dff_A_nNxW80mH2_0),.clk(gclk));
	jdff dff_A_9TjaYfXT7_0(.dout(w_dff_A_ML3DyYOs9_0),.din(w_dff_A_9TjaYfXT7_0),.clk(gclk));
	jdff dff_A_ML3DyYOs9_0(.dout(w_dff_A_PNfzOgcU1_0),.din(w_dff_A_ML3DyYOs9_0),.clk(gclk));
	jdff dff_A_PNfzOgcU1_0(.dout(G558),.din(w_dff_A_PNfzOgcU1_0),.clk(gclk));
	jdff dff_A_jDpzQ2aJ2_1(.dout(w_dff_A_tY6dgRov0_0),.din(w_dff_A_jDpzQ2aJ2_1),.clk(gclk));
	jdff dff_A_tY6dgRov0_0(.dout(w_dff_A_EHAtL1do0_0),.din(w_dff_A_tY6dgRov0_0),.clk(gclk));
	jdff dff_A_EHAtL1do0_0(.dout(w_dff_A_i0qYNqRV0_0),.din(w_dff_A_EHAtL1do0_0),.clk(gclk));
	jdff dff_A_i0qYNqRV0_0(.dout(w_dff_A_m6viLzn54_0),.din(w_dff_A_i0qYNqRV0_0),.clk(gclk));
	jdff dff_A_m6viLzn54_0(.dout(w_dff_A_rw57U0QD9_0),.din(w_dff_A_m6viLzn54_0),.clk(gclk));
	jdff dff_A_rw57U0QD9_0(.dout(w_dff_A_gzSKvJmH2_0),.din(w_dff_A_rw57U0QD9_0),.clk(gclk));
	jdff dff_A_gzSKvJmH2_0(.dout(w_dff_A_X6wI6tdu2_0),.din(w_dff_A_gzSKvJmH2_0),.clk(gclk));
	jdff dff_A_X6wI6tdu2_0(.dout(w_dff_A_yxJcPIOq2_0),.din(w_dff_A_X6wI6tdu2_0),.clk(gclk));
	jdff dff_A_yxJcPIOq2_0(.dout(w_dff_A_6q6pHyw23_0),.din(w_dff_A_yxJcPIOq2_0),.clk(gclk));
	jdff dff_A_6q6pHyw23_0(.dout(w_dff_A_k436aywX5_0),.din(w_dff_A_6q6pHyw23_0),.clk(gclk));
	jdff dff_A_k436aywX5_0(.dout(w_dff_A_LqiquxaA5_0),.din(w_dff_A_k436aywX5_0),.clk(gclk));
	jdff dff_A_LqiquxaA5_0(.dout(w_dff_A_MQPK4MpP8_0),.din(w_dff_A_LqiquxaA5_0),.clk(gclk));
	jdff dff_A_MQPK4MpP8_0(.dout(w_dff_A_diWiusl89_0),.din(w_dff_A_MQPK4MpP8_0),.clk(gclk));
	jdff dff_A_diWiusl89_0(.dout(w_dff_A_OFaqqzmH6_0),.din(w_dff_A_diWiusl89_0),.clk(gclk));
	jdff dff_A_OFaqqzmH6_0(.dout(w_dff_A_JDeGCL5C5_0),.din(w_dff_A_OFaqqzmH6_0),.clk(gclk));
	jdff dff_A_JDeGCL5C5_0(.dout(w_dff_A_6SibfMMf0_0),.din(w_dff_A_JDeGCL5C5_0),.clk(gclk));
	jdff dff_A_6SibfMMf0_0(.dout(w_dff_A_z2Fv1A696_0),.din(w_dff_A_6SibfMMf0_0),.clk(gclk));
	jdff dff_A_z2Fv1A696_0(.dout(w_dff_A_BVx5WgYL6_0),.din(w_dff_A_z2Fv1A696_0),.clk(gclk));
	jdff dff_A_BVx5WgYL6_0(.dout(w_dff_A_9yBqeMOd0_0),.din(w_dff_A_BVx5WgYL6_0),.clk(gclk));
	jdff dff_A_9yBqeMOd0_0(.dout(w_dff_A_CbC1PrI46_0),.din(w_dff_A_9yBqeMOd0_0),.clk(gclk));
	jdff dff_A_CbC1PrI46_0(.dout(w_dff_A_wOYDwEvW2_0),.din(w_dff_A_CbC1PrI46_0),.clk(gclk));
	jdff dff_A_wOYDwEvW2_0(.dout(w_dff_A_wEfDM12M5_0),.din(w_dff_A_wOYDwEvW2_0),.clk(gclk));
	jdff dff_A_wEfDM12M5_0(.dout(w_dff_A_FZBkPWEB6_0),.din(w_dff_A_wEfDM12M5_0),.clk(gclk));
	jdff dff_A_FZBkPWEB6_0(.dout(w_dff_A_IKrTG20f5_0),.din(w_dff_A_FZBkPWEB6_0),.clk(gclk));
	jdff dff_A_IKrTG20f5_0(.dout(w_dff_A_LedmHbcG8_0),.din(w_dff_A_IKrTG20f5_0),.clk(gclk));
	jdff dff_A_LedmHbcG8_0(.dout(w_dff_A_eUsqHrRl3_0),.din(w_dff_A_LedmHbcG8_0),.clk(gclk));
	jdff dff_A_eUsqHrRl3_0(.dout(G556),.din(w_dff_A_eUsqHrRl3_0),.clk(gclk));
	jdff dff_A_Y9ZWrAog2_1(.dout(w_dff_A_veWLWexF3_0),.din(w_dff_A_Y9ZWrAog2_1),.clk(gclk));
	jdff dff_A_veWLWexF3_0(.dout(w_dff_A_VjLX6Z4I1_0),.din(w_dff_A_veWLWexF3_0),.clk(gclk));
	jdff dff_A_VjLX6Z4I1_0(.dout(w_dff_A_qzyMCrWd1_0),.din(w_dff_A_VjLX6Z4I1_0),.clk(gclk));
	jdff dff_A_qzyMCrWd1_0(.dout(w_dff_A_eujmvK7H4_0),.din(w_dff_A_qzyMCrWd1_0),.clk(gclk));
	jdff dff_A_eujmvK7H4_0(.dout(w_dff_A_7YKFQXcO3_0),.din(w_dff_A_eujmvK7H4_0),.clk(gclk));
	jdff dff_A_7YKFQXcO3_0(.dout(w_dff_A_12nbvWII9_0),.din(w_dff_A_7YKFQXcO3_0),.clk(gclk));
	jdff dff_A_12nbvWII9_0(.dout(w_dff_A_2QTP7w2N8_0),.din(w_dff_A_12nbvWII9_0),.clk(gclk));
	jdff dff_A_2QTP7w2N8_0(.dout(w_dff_A_1PPORM3p0_0),.din(w_dff_A_2QTP7w2N8_0),.clk(gclk));
	jdff dff_A_1PPORM3p0_0(.dout(w_dff_A_leaXiWlx9_0),.din(w_dff_A_1PPORM3p0_0),.clk(gclk));
	jdff dff_A_leaXiWlx9_0(.dout(w_dff_A_hT6xkbQA0_0),.din(w_dff_A_leaXiWlx9_0),.clk(gclk));
	jdff dff_A_hT6xkbQA0_0(.dout(w_dff_A_psJDiScC5_0),.din(w_dff_A_hT6xkbQA0_0),.clk(gclk));
	jdff dff_A_psJDiScC5_0(.dout(w_dff_A_1ES4KZKm2_0),.din(w_dff_A_psJDiScC5_0),.clk(gclk));
	jdff dff_A_1ES4KZKm2_0(.dout(w_dff_A_tTh4NykM4_0),.din(w_dff_A_1ES4KZKm2_0),.clk(gclk));
	jdff dff_A_tTh4NykM4_0(.dout(w_dff_A_3em2Unc16_0),.din(w_dff_A_tTh4NykM4_0),.clk(gclk));
	jdff dff_A_3em2Unc16_0(.dout(w_dff_A_ZVgxaHto9_0),.din(w_dff_A_3em2Unc16_0),.clk(gclk));
	jdff dff_A_ZVgxaHto9_0(.dout(w_dff_A_stIc75sl6_0),.din(w_dff_A_ZVgxaHto9_0),.clk(gclk));
	jdff dff_A_stIc75sl6_0(.dout(w_dff_A_5r9aLTWK6_0),.din(w_dff_A_stIc75sl6_0),.clk(gclk));
	jdff dff_A_5r9aLTWK6_0(.dout(w_dff_A_vvVAzQhW6_0),.din(w_dff_A_5r9aLTWK6_0),.clk(gclk));
	jdff dff_A_vvVAzQhW6_0(.dout(w_dff_A_A291gemr5_0),.din(w_dff_A_vvVAzQhW6_0),.clk(gclk));
	jdff dff_A_A291gemr5_0(.dout(w_dff_A_3J09ytV54_0),.din(w_dff_A_A291gemr5_0),.clk(gclk));
	jdff dff_A_3J09ytV54_0(.dout(w_dff_A_gVJLw4Hz0_0),.din(w_dff_A_3J09ytV54_0),.clk(gclk));
	jdff dff_A_gVJLw4Hz0_0(.dout(w_dff_A_nTTKElQZ6_0),.din(w_dff_A_gVJLw4Hz0_0),.clk(gclk));
	jdff dff_A_nTTKElQZ6_0(.dout(w_dff_A_nj8LPSUi8_0),.din(w_dff_A_nTTKElQZ6_0),.clk(gclk));
	jdff dff_A_nj8LPSUi8_0(.dout(w_dff_A_TWLlZgxQ6_0),.din(w_dff_A_nj8LPSUi8_0),.clk(gclk));
	jdff dff_A_TWLlZgxQ6_0(.dout(w_dff_A_ROH6L8Mh1_0),.din(w_dff_A_TWLlZgxQ6_0),.clk(gclk));
	jdff dff_A_ROH6L8Mh1_0(.dout(w_dff_A_gqAy88Wv7_0),.din(w_dff_A_ROH6L8Mh1_0),.clk(gclk));
	jdff dff_A_gqAy88Wv7_0(.dout(G554),.din(w_dff_A_gqAy88Wv7_0),.clk(gclk));
	jdff dff_A_0ix5qubp0_1(.dout(w_dff_A_60e6HO8E1_0),.din(w_dff_A_0ix5qubp0_1),.clk(gclk));
	jdff dff_A_60e6HO8E1_0(.dout(w_dff_A_Z2ux1dkz1_0),.din(w_dff_A_60e6HO8E1_0),.clk(gclk));
	jdff dff_A_Z2ux1dkz1_0(.dout(w_dff_A_EZ3yinoM9_0),.din(w_dff_A_Z2ux1dkz1_0),.clk(gclk));
	jdff dff_A_EZ3yinoM9_0(.dout(w_dff_A_QWkUBcJB8_0),.din(w_dff_A_EZ3yinoM9_0),.clk(gclk));
	jdff dff_A_QWkUBcJB8_0(.dout(w_dff_A_bGH9w2Qj4_0),.din(w_dff_A_QWkUBcJB8_0),.clk(gclk));
	jdff dff_A_bGH9w2Qj4_0(.dout(w_dff_A_d0037ciS8_0),.din(w_dff_A_bGH9w2Qj4_0),.clk(gclk));
	jdff dff_A_d0037ciS8_0(.dout(w_dff_A_mY2sA8sQ3_0),.din(w_dff_A_d0037ciS8_0),.clk(gclk));
	jdff dff_A_mY2sA8sQ3_0(.dout(w_dff_A_cOMZIl043_0),.din(w_dff_A_mY2sA8sQ3_0),.clk(gclk));
	jdff dff_A_cOMZIl043_0(.dout(w_dff_A_qFEhImj31_0),.din(w_dff_A_cOMZIl043_0),.clk(gclk));
	jdff dff_A_qFEhImj31_0(.dout(w_dff_A_YbSTgncB9_0),.din(w_dff_A_qFEhImj31_0),.clk(gclk));
	jdff dff_A_YbSTgncB9_0(.dout(w_dff_A_ytvceTSx1_0),.din(w_dff_A_YbSTgncB9_0),.clk(gclk));
	jdff dff_A_ytvceTSx1_0(.dout(w_dff_A_MDckOEme9_0),.din(w_dff_A_ytvceTSx1_0),.clk(gclk));
	jdff dff_A_MDckOEme9_0(.dout(w_dff_A_y0MGcsvL5_0),.din(w_dff_A_MDckOEme9_0),.clk(gclk));
	jdff dff_A_y0MGcsvL5_0(.dout(w_dff_A_dOX4LlK39_0),.din(w_dff_A_y0MGcsvL5_0),.clk(gclk));
	jdff dff_A_dOX4LlK39_0(.dout(w_dff_A_sZLpTzAN4_0),.din(w_dff_A_dOX4LlK39_0),.clk(gclk));
	jdff dff_A_sZLpTzAN4_0(.dout(w_dff_A_Mthay0yB5_0),.din(w_dff_A_sZLpTzAN4_0),.clk(gclk));
	jdff dff_A_Mthay0yB5_0(.dout(w_dff_A_n0OAJnoI5_0),.din(w_dff_A_Mthay0yB5_0),.clk(gclk));
	jdff dff_A_n0OAJnoI5_0(.dout(w_dff_A_YW1X6Ocm5_0),.din(w_dff_A_n0OAJnoI5_0),.clk(gclk));
	jdff dff_A_YW1X6Ocm5_0(.dout(w_dff_A_xRQAyEz31_0),.din(w_dff_A_YW1X6Ocm5_0),.clk(gclk));
	jdff dff_A_xRQAyEz31_0(.dout(w_dff_A_BPAb1zIa4_0),.din(w_dff_A_xRQAyEz31_0),.clk(gclk));
	jdff dff_A_BPAb1zIa4_0(.dout(w_dff_A_EUz3i6PF0_0),.din(w_dff_A_BPAb1zIa4_0),.clk(gclk));
	jdff dff_A_EUz3i6PF0_0(.dout(w_dff_A_5PhaOWOG5_0),.din(w_dff_A_EUz3i6PF0_0),.clk(gclk));
	jdff dff_A_5PhaOWOG5_0(.dout(w_dff_A_gXxTGb2c8_0),.din(w_dff_A_5PhaOWOG5_0),.clk(gclk));
	jdff dff_A_gXxTGb2c8_0(.dout(w_dff_A_Gqzrmer73_0),.din(w_dff_A_gXxTGb2c8_0),.clk(gclk));
	jdff dff_A_Gqzrmer73_0(.dout(w_dff_A_CeobTZQr2_0),.din(w_dff_A_Gqzrmer73_0),.clk(gclk));
	jdff dff_A_CeobTZQr2_0(.dout(w_dff_A_YbAhygpP0_0),.din(w_dff_A_CeobTZQr2_0),.clk(gclk));
	jdff dff_A_YbAhygpP0_0(.dout(G552),.din(w_dff_A_YbAhygpP0_0),.clk(gclk));
	jdff dff_A_wgAbeICk9_1(.dout(w_dff_A_vQ8ykfQd3_0),.din(w_dff_A_wgAbeICk9_1),.clk(gclk));
	jdff dff_A_vQ8ykfQd3_0(.dout(w_dff_A_j2h5m3TC8_0),.din(w_dff_A_vQ8ykfQd3_0),.clk(gclk));
	jdff dff_A_j2h5m3TC8_0(.dout(w_dff_A_Dd33UVEf8_0),.din(w_dff_A_j2h5m3TC8_0),.clk(gclk));
	jdff dff_A_Dd33UVEf8_0(.dout(w_dff_A_dzhl3jx75_0),.din(w_dff_A_Dd33UVEf8_0),.clk(gclk));
	jdff dff_A_dzhl3jx75_0(.dout(w_dff_A_meYIlkPJ0_0),.din(w_dff_A_dzhl3jx75_0),.clk(gclk));
	jdff dff_A_meYIlkPJ0_0(.dout(w_dff_A_h8FAtpXP9_0),.din(w_dff_A_meYIlkPJ0_0),.clk(gclk));
	jdff dff_A_h8FAtpXP9_0(.dout(w_dff_A_CcuA5gcs9_0),.din(w_dff_A_h8FAtpXP9_0),.clk(gclk));
	jdff dff_A_CcuA5gcs9_0(.dout(w_dff_A_kPlsGiaz6_0),.din(w_dff_A_CcuA5gcs9_0),.clk(gclk));
	jdff dff_A_kPlsGiaz6_0(.dout(w_dff_A_q47dh4Xv9_0),.din(w_dff_A_kPlsGiaz6_0),.clk(gclk));
	jdff dff_A_q47dh4Xv9_0(.dout(w_dff_A_xlbTtHlf3_0),.din(w_dff_A_q47dh4Xv9_0),.clk(gclk));
	jdff dff_A_xlbTtHlf3_0(.dout(w_dff_A_uON0jOl05_0),.din(w_dff_A_xlbTtHlf3_0),.clk(gclk));
	jdff dff_A_uON0jOl05_0(.dout(w_dff_A_qENXP1JA3_0),.din(w_dff_A_uON0jOl05_0),.clk(gclk));
	jdff dff_A_qENXP1JA3_0(.dout(w_dff_A_lZXgQIRJ8_0),.din(w_dff_A_qENXP1JA3_0),.clk(gclk));
	jdff dff_A_lZXgQIRJ8_0(.dout(w_dff_A_FZ8KGm6o0_0),.din(w_dff_A_lZXgQIRJ8_0),.clk(gclk));
	jdff dff_A_FZ8KGm6o0_0(.dout(w_dff_A_DYVita5t1_0),.din(w_dff_A_FZ8KGm6o0_0),.clk(gclk));
	jdff dff_A_DYVita5t1_0(.dout(w_dff_A_R1FFuPv26_0),.din(w_dff_A_DYVita5t1_0),.clk(gclk));
	jdff dff_A_R1FFuPv26_0(.dout(w_dff_A_u3u5S29D7_0),.din(w_dff_A_R1FFuPv26_0),.clk(gclk));
	jdff dff_A_u3u5S29D7_0(.dout(w_dff_A_Dm5cneEl9_0),.din(w_dff_A_u3u5S29D7_0),.clk(gclk));
	jdff dff_A_Dm5cneEl9_0(.dout(w_dff_A_MBIAjK7l3_0),.din(w_dff_A_Dm5cneEl9_0),.clk(gclk));
	jdff dff_A_MBIAjK7l3_0(.dout(w_dff_A_BK3uQb7X5_0),.din(w_dff_A_MBIAjK7l3_0),.clk(gclk));
	jdff dff_A_BK3uQb7X5_0(.dout(w_dff_A_DOB6QybZ2_0),.din(w_dff_A_BK3uQb7X5_0),.clk(gclk));
	jdff dff_A_DOB6QybZ2_0(.dout(w_dff_A_YgReLinE3_0),.din(w_dff_A_DOB6QybZ2_0),.clk(gclk));
	jdff dff_A_YgReLinE3_0(.dout(w_dff_A_9rKlEP7H9_0),.din(w_dff_A_YgReLinE3_0),.clk(gclk));
	jdff dff_A_9rKlEP7H9_0(.dout(w_dff_A_q0Ahveqj8_0),.din(w_dff_A_9rKlEP7H9_0),.clk(gclk));
	jdff dff_A_q0Ahveqj8_0(.dout(w_dff_A_LgfPKULk3_0),.din(w_dff_A_q0Ahveqj8_0),.clk(gclk));
	jdff dff_A_LgfPKULk3_0(.dout(w_dff_A_bR8O3B8A6_0),.din(w_dff_A_LgfPKULk3_0),.clk(gclk));
	jdff dff_A_bR8O3B8A6_0(.dout(G550),.din(w_dff_A_bR8O3B8A6_0),.clk(gclk));
	jdff dff_A_CfDvIimZ4_1(.dout(w_dff_A_3SY1fYpy2_0),.din(w_dff_A_CfDvIimZ4_1),.clk(gclk));
	jdff dff_A_3SY1fYpy2_0(.dout(w_dff_A_uKP3BkAP2_0),.din(w_dff_A_3SY1fYpy2_0),.clk(gclk));
	jdff dff_A_uKP3BkAP2_0(.dout(w_dff_A_O0bRRyHm6_0),.din(w_dff_A_uKP3BkAP2_0),.clk(gclk));
	jdff dff_A_O0bRRyHm6_0(.dout(w_dff_A_tG6w6lsh6_0),.din(w_dff_A_O0bRRyHm6_0),.clk(gclk));
	jdff dff_A_tG6w6lsh6_0(.dout(w_dff_A_C3h7PFtu4_0),.din(w_dff_A_tG6w6lsh6_0),.clk(gclk));
	jdff dff_A_C3h7PFtu4_0(.dout(w_dff_A_l5AKPo0Y7_0),.din(w_dff_A_C3h7PFtu4_0),.clk(gclk));
	jdff dff_A_l5AKPo0Y7_0(.dout(w_dff_A_AtfozGDW8_0),.din(w_dff_A_l5AKPo0Y7_0),.clk(gclk));
	jdff dff_A_AtfozGDW8_0(.dout(w_dff_A_rfKqZ5L64_0),.din(w_dff_A_AtfozGDW8_0),.clk(gclk));
	jdff dff_A_rfKqZ5L64_0(.dout(w_dff_A_1QBmeoPQ4_0),.din(w_dff_A_rfKqZ5L64_0),.clk(gclk));
	jdff dff_A_1QBmeoPQ4_0(.dout(w_dff_A_8EEFaWvJ3_0),.din(w_dff_A_1QBmeoPQ4_0),.clk(gclk));
	jdff dff_A_8EEFaWvJ3_0(.dout(w_dff_A_SDT7cqFV1_0),.din(w_dff_A_8EEFaWvJ3_0),.clk(gclk));
	jdff dff_A_SDT7cqFV1_0(.dout(w_dff_A_n6JsGTOj6_0),.din(w_dff_A_SDT7cqFV1_0),.clk(gclk));
	jdff dff_A_n6JsGTOj6_0(.dout(w_dff_A_96C6UDXs3_0),.din(w_dff_A_n6JsGTOj6_0),.clk(gclk));
	jdff dff_A_96C6UDXs3_0(.dout(w_dff_A_dXzzdVar1_0),.din(w_dff_A_96C6UDXs3_0),.clk(gclk));
	jdff dff_A_dXzzdVar1_0(.dout(w_dff_A_7U8X5o2u5_0),.din(w_dff_A_dXzzdVar1_0),.clk(gclk));
	jdff dff_A_7U8X5o2u5_0(.dout(w_dff_A_BEJd0wnq5_0),.din(w_dff_A_7U8X5o2u5_0),.clk(gclk));
	jdff dff_A_BEJd0wnq5_0(.dout(w_dff_A_OtxYU6Rj0_0),.din(w_dff_A_BEJd0wnq5_0),.clk(gclk));
	jdff dff_A_OtxYU6Rj0_0(.dout(w_dff_A_ODJEpXD01_0),.din(w_dff_A_OtxYU6Rj0_0),.clk(gclk));
	jdff dff_A_ODJEpXD01_0(.dout(w_dff_A_wDhPmN9S6_0),.din(w_dff_A_ODJEpXD01_0),.clk(gclk));
	jdff dff_A_wDhPmN9S6_0(.dout(w_dff_A_s2FFEnfo6_0),.din(w_dff_A_wDhPmN9S6_0),.clk(gclk));
	jdff dff_A_s2FFEnfo6_0(.dout(w_dff_A_8M1x1tpL9_0),.din(w_dff_A_s2FFEnfo6_0),.clk(gclk));
	jdff dff_A_8M1x1tpL9_0(.dout(w_dff_A_v6FtbG5R7_0),.din(w_dff_A_8M1x1tpL9_0),.clk(gclk));
	jdff dff_A_v6FtbG5R7_0(.dout(w_dff_A_EwTfW2S17_0),.din(w_dff_A_v6FtbG5R7_0),.clk(gclk));
	jdff dff_A_EwTfW2S17_0(.dout(w_dff_A_nwVFLuv12_0),.din(w_dff_A_EwTfW2S17_0),.clk(gclk));
	jdff dff_A_nwVFLuv12_0(.dout(w_dff_A_clYmrU0C9_0),.din(w_dff_A_nwVFLuv12_0),.clk(gclk));
	jdff dff_A_clYmrU0C9_0(.dout(w_dff_A_acC3lP8G3_0),.din(w_dff_A_clYmrU0C9_0),.clk(gclk));
	jdff dff_A_acC3lP8G3_0(.dout(G548),.din(w_dff_A_acC3lP8G3_0),.clk(gclk));
	jdff dff_A_8brKNuEG7_1(.dout(w_dff_A_aKo1Xqn97_0),.din(w_dff_A_8brKNuEG7_1),.clk(gclk));
	jdff dff_A_aKo1Xqn97_0(.dout(w_dff_A_elwKw87q0_0),.din(w_dff_A_aKo1Xqn97_0),.clk(gclk));
	jdff dff_A_elwKw87q0_0(.dout(w_dff_A_4fS7H4Po8_0),.din(w_dff_A_elwKw87q0_0),.clk(gclk));
	jdff dff_A_4fS7H4Po8_0(.dout(w_dff_A_rVUE7aOe2_0),.din(w_dff_A_4fS7H4Po8_0),.clk(gclk));
	jdff dff_A_rVUE7aOe2_0(.dout(w_dff_A_t2roooUt4_0),.din(w_dff_A_rVUE7aOe2_0),.clk(gclk));
	jdff dff_A_t2roooUt4_0(.dout(w_dff_A_95swoQu66_0),.din(w_dff_A_t2roooUt4_0),.clk(gclk));
	jdff dff_A_95swoQu66_0(.dout(w_dff_A_n6FSe3V11_0),.din(w_dff_A_95swoQu66_0),.clk(gclk));
	jdff dff_A_n6FSe3V11_0(.dout(w_dff_A_XMF7208w7_0),.din(w_dff_A_n6FSe3V11_0),.clk(gclk));
	jdff dff_A_XMF7208w7_0(.dout(w_dff_A_9TuXXtwC8_0),.din(w_dff_A_XMF7208w7_0),.clk(gclk));
	jdff dff_A_9TuXXtwC8_0(.dout(w_dff_A_rEO7qQeb3_0),.din(w_dff_A_9TuXXtwC8_0),.clk(gclk));
	jdff dff_A_rEO7qQeb3_0(.dout(w_dff_A_rjuN1Y3Z7_0),.din(w_dff_A_rEO7qQeb3_0),.clk(gclk));
	jdff dff_A_rjuN1Y3Z7_0(.dout(w_dff_A_dVBFye6q9_0),.din(w_dff_A_rjuN1Y3Z7_0),.clk(gclk));
	jdff dff_A_dVBFye6q9_0(.dout(w_dff_A_JNkmNgcG5_0),.din(w_dff_A_dVBFye6q9_0),.clk(gclk));
	jdff dff_A_JNkmNgcG5_0(.dout(w_dff_A_VbNjRkFM5_0),.din(w_dff_A_JNkmNgcG5_0),.clk(gclk));
	jdff dff_A_VbNjRkFM5_0(.dout(w_dff_A_FAQvIRpn3_0),.din(w_dff_A_VbNjRkFM5_0),.clk(gclk));
	jdff dff_A_FAQvIRpn3_0(.dout(w_dff_A_VPqPdqFI2_0),.din(w_dff_A_FAQvIRpn3_0),.clk(gclk));
	jdff dff_A_VPqPdqFI2_0(.dout(w_dff_A_yJloMtev6_0),.din(w_dff_A_VPqPdqFI2_0),.clk(gclk));
	jdff dff_A_yJloMtev6_0(.dout(w_dff_A_5X8zdgpV2_0),.din(w_dff_A_yJloMtev6_0),.clk(gclk));
	jdff dff_A_5X8zdgpV2_0(.dout(w_dff_A_iC4Re1dy6_0),.din(w_dff_A_5X8zdgpV2_0),.clk(gclk));
	jdff dff_A_iC4Re1dy6_0(.dout(w_dff_A_Ra8tLkuT0_0),.din(w_dff_A_iC4Re1dy6_0),.clk(gclk));
	jdff dff_A_Ra8tLkuT0_0(.dout(w_dff_A_gWn9kqhU6_0),.din(w_dff_A_Ra8tLkuT0_0),.clk(gclk));
	jdff dff_A_gWn9kqhU6_0(.dout(w_dff_A_yh6t0Gq15_0),.din(w_dff_A_gWn9kqhU6_0),.clk(gclk));
	jdff dff_A_yh6t0Gq15_0(.dout(w_dff_A_qhpoD1r02_0),.din(w_dff_A_yh6t0Gq15_0),.clk(gclk));
	jdff dff_A_qhpoD1r02_0(.dout(w_dff_A_G2sZBwY77_0),.din(w_dff_A_qhpoD1r02_0),.clk(gclk));
	jdff dff_A_G2sZBwY77_0(.dout(w_dff_A_2TcBThQC9_0),.din(w_dff_A_G2sZBwY77_0),.clk(gclk));
	jdff dff_A_2TcBThQC9_0(.dout(w_dff_A_jE64nwd89_0),.din(w_dff_A_2TcBThQC9_0),.clk(gclk));
	jdff dff_A_jE64nwd89_0(.dout(G546),.din(w_dff_A_jE64nwd89_0),.clk(gclk));
	jdff dff_A_Sld5T4WZ8_1(.dout(w_dff_A_34QmGbZl7_0),.din(w_dff_A_Sld5T4WZ8_1),.clk(gclk));
	jdff dff_A_34QmGbZl7_0(.dout(w_dff_A_9KFCa8dQ2_0),.din(w_dff_A_34QmGbZl7_0),.clk(gclk));
	jdff dff_A_9KFCa8dQ2_0(.dout(w_dff_A_gote9Jjd3_0),.din(w_dff_A_9KFCa8dQ2_0),.clk(gclk));
	jdff dff_A_gote9Jjd3_0(.dout(w_dff_A_YIm6Z9Vd4_0),.din(w_dff_A_gote9Jjd3_0),.clk(gclk));
	jdff dff_A_YIm6Z9Vd4_0(.dout(w_dff_A_KBMQbzEZ9_0),.din(w_dff_A_YIm6Z9Vd4_0),.clk(gclk));
	jdff dff_A_KBMQbzEZ9_0(.dout(w_dff_A_njBJA7ZT7_0),.din(w_dff_A_KBMQbzEZ9_0),.clk(gclk));
	jdff dff_A_njBJA7ZT7_0(.dout(w_dff_A_B4BINbny2_0),.din(w_dff_A_njBJA7ZT7_0),.clk(gclk));
	jdff dff_A_B4BINbny2_0(.dout(w_dff_A_xR9vKVC29_0),.din(w_dff_A_B4BINbny2_0),.clk(gclk));
	jdff dff_A_xR9vKVC29_0(.dout(w_dff_A_jKxq7Lip5_0),.din(w_dff_A_xR9vKVC29_0),.clk(gclk));
	jdff dff_A_jKxq7Lip5_0(.dout(w_dff_A_dHZk470L8_0),.din(w_dff_A_jKxq7Lip5_0),.clk(gclk));
	jdff dff_A_dHZk470L8_0(.dout(w_dff_A_TRp6IpqA5_0),.din(w_dff_A_dHZk470L8_0),.clk(gclk));
	jdff dff_A_TRp6IpqA5_0(.dout(w_dff_A_lmQL2zhz7_0),.din(w_dff_A_TRp6IpqA5_0),.clk(gclk));
	jdff dff_A_lmQL2zhz7_0(.dout(w_dff_A_I62zzrR90_0),.din(w_dff_A_lmQL2zhz7_0),.clk(gclk));
	jdff dff_A_I62zzrR90_0(.dout(w_dff_A_OlGyySJg5_0),.din(w_dff_A_I62zzrR90_0),.clk(gclk));
	jdff dff_A_OlGyySJg5_0(.dout(w_dff_A_TDuLjLqF6_0),.din(w_dff_A_OlGyySJg5_0),.clk(gclk));
	jdff dff_A_TDuLjLqF6_0(.dout(w_dff_A_aEu9tbAC6_0),.din(w_dff_A_TDuLjLqF6_0),.clk(gclk));
	jdff dff_A_aEu9tbAC6_0(.dout(w_dff_A_BIXzmfRq9_0),.din(w_dff_A_aEu9tbAC6_0),.clk(gclk));
	jdff dff_A_BIXzmfRq9_0(.dout(w_dff_A_zRqCkXAm6_0),.din(w_dff_A_BIXzmfRq9_0),.clk(gclk));
	jdff dff_A_zRqCkXAm6_0(.dout(w_dff_A_AXlRiLPI0_0),.din(w_dff_A_zRqCkXAm6_0),.clk(gclk));
	jdff dff_A_AXlRiLPI0_0(.dout(w_dff_A_yWTt5LKp9_0),.din(w_dff_A_AXlRiLPI0_0),.clk(gclk));
	jdff dff_A_yWTt5LKp9_0(.dout(w_dff_A_I6mraCGq5_0),.din(w_dff_A_yWTt5LKp9_0),.clk(gclk));
	jdff dff_A_I6mraCGq5_0(.dout(w_dff_A_KLEEW6wB9_0),.din(w_dff_A_I6mraCGq5_0),.clk(gclk));
	jdff dff_A_KLEEW6wB9_0(.dout(w_dff_A_vJZZpSxL3_0),.din(w_dff_A_KLEEW6wB9_0),.clk(gclk));
	jdff dff_A_vJZZpSxL3_0(.dout(w_dff_A_ebtkvx0J8_0),.din(w_dff_A_vJZZpSxL3_0),.clk(gclk));
	jdff dff_A_ebtkvx0J8_0(.dout(w_dff_A_0i8fxZ8s6_0),.din(w_dff_A_ebtkvx0J8_0),.clk(gclk));
	jdff dff_A_0i8fxZ8s6_0(.dout(w_dff_A_p1vOkPhX0_0),.din(w_dff_A_0i8fxZ8s6_0),.clk(gclk));
	jdff dff_A_p1vOkPhX0_0(.dout(G544),.din(w_dff_A_p1vOkPhX0_0),.clk(gclk));
	jdff dff_A_2zsj2RB06_1(.dout(w_dff_A_4fMokPse6_0),.din(w_dff_A_2zsj2RB06_1),.clk(gclk));
	jdff dff_A_4fMokPse6_0(.dout(w_dff_A_tL7I77yW6_0),.din(w_dff_A_4fMokPse6_0),.clk(gclk));
	jdff dff_A_tL7I77yW6_0(.dout(w_dff_A_jVhbtRls8_0),.din(w_dff_A_tL7I77yW6_0),.clk(gclk));
	jdff dff_A_jVhbtRls8_0(.dout(w_dff_A_OwzqNQWn2_0),.din(w_dff_A_jVhbtRls8_0),.clk(gclk));
	jdff dff_A_OwzqNQWn2_0(.dout(w_dff_A_zbNCJ00i7_0),.din(w_dff_A_OwzqNQWn2_0),.clk(gclk));
	jdff dff_A_zbNCJ00i7_0(.dout(w_dff_A_GEt8cfV60_0),.din(w_dff_A_zbNCJ00i7_0),.clk(gclk));
	jdff dff_A_GEt8cfV60_0(.dout(w_dff_A_0ed7RTf54_0),.din(w_dff_A_GEt8cfV60_0),.clk(gclk));
	jdff dff_A_0ed7RTf54_0(.dout(w_dff_A_KDARhFIF8_0),.din(w_dff_A_0ed7RTf54_0),.clk(gclk));
	jdff dff_A_KDARhFIF8_0(.dout(w_dff_A_S15NTq9M3_0),.din(w_dff_A_KDARhFIF8_0),.clk(gclk));
	jdff dff_A_S15NTq9M3_0(.dout(w_dff_A_og65d4NS6_0),.din(w_dff_A_S15NTq9M3_0),.clk(gclk));
	jdff dff_A_og65d4NS6_0(.dout(w_dff_A_h0OQBv3X3_0),.din(w_dff_A_og65d4NS6_0),.clk(gclk));
	jdff dff_A_h0OQBv3X3_0(.dout(w_dff_A_2XRTt7va0_0),.din(w_dff_A_h0OQBv3X3_0),.clk(gclk));
	jdff dff_A_2XRTt7va0_0(.dout(w_dff_A_6gimJ83V0_0),.din(w_dff_A_2XRTt7va0_0),.clk(gclk));
	jdff dff_A_6gimJ83V0_0(.dout(w_dff_A_uNM2lJSj5_0),.din(w_dff_A_6gimJ83V0_0),.clk(gclk));
	jdff dff_A_uNM2lJSj5_0(.dout(w_dff_A_8LKvGAMC6_0),.din(w_dff_A_uNM2lJSj5_0),.clk(gclk));
	jdff dff_A_8LKvGAMC6_0(.dout(w_dff_A_WKWR70IY2_0),.din(w_dff_A_8LKvGAMC6_0),.clk(gclk));
	jdff dff_A_WKWR70IY2_0(.dout(w_dff_A_Zr0bAJhg2_0),.din(w_dff_A_WKWR70IY2_0),.clk(gclk));
	jdff dff_A_Zr0bAJhg2_0(.dout(w_dff_A_elYa4sC54_0),.din(w_dff_A_Zr0bAJhg2_0),.clk(gclk));
	jdff dff_A_elYa4sC54_0(.dout(w_dff_A_0eIlEFHI3_0),.din(w_dff_A_elYa4sC54_0),.clk(gclk));
	jdff dff_A_0eIlEFHI3_0(.dout(w_dff_A_GiLMeY3g4_0),.din(w_dff_A_0eIlEFHI3_0),.clk(gclk));
	jdff dff_A_GiLMeY3g4_0(.dout(w_dff_A_upXG6BSh9_0),.din(w_dff_A_GiLMeY3g4_0),.clk(gclk));
	jdff dff_A_upXG6BSh9_0(.dout(w_dff_A_8IeNdCz23_0),.din(w_dff_A_upXG6BSh9_0),.clk(gclk));
	jdff dff_A_8IeNdCz23_0(.dout(w_dff_A_X7apPuCr8_0),.din(w_dff_A_8IeNdCz23_0),.clk(gclk));
	jdff dff_A_X7apPuCr8_0(.dout(w_dff_A_qTXzhp2l6_0),.din(w_dff_A_X7apPuCr8_0),.clk(gclk));
	jdff dff_A_qTXzhp2l6_0(.dout(w_dff_A_HWXg7uXL3_0),.din(w_dff_A_qTXzhp2l6_0),.clk(gclk));
	jdff dff_A_HWXg7uXL3_0(.dout(w_dff_A_9RVvguRJ3_0),.din(w_dff_A_HWXg7uXL3_0),.clk(gclk));
	jdff dff_A_9RVvguRJ3_0(.dout(G540),.din(w_dff_A_9RVvguRJ3_0),.clk(gclk));
	jdff dff_A_r0bXZQNs5_1(.dout(w_dff_A_TYUuYlol5_0),.din(w_dff_A_r0bXZQNs5_1),.clk(gclk));
	jdff dff_A_TYUuYlol5_0(.dout(w_dff_A_jJvJxAKt8_0),.din(w_dff_A_TYUuYlol5_0),.clk(gclk));
	jdff dff_A_jJvJxAKt8_0(.dout(w_dff_A_m93Et6xG1_0),.din(w_dff_A_jJvJxAKt8_0),.clk(gclk));
	jdff dff_A_m93Et6xG1_0(.dout(w_dff_A_1kpfSZtl7_0),.din(w_dff_A_m93Et6xG1_0),.clk(gclk));
	jdff dff_A_1kpfSZtl7_0(.dout(w_dff_A_AE3LxU6A4_0),.din(w_dff_A_1kpfSZtl7_0),.clk(gclk));
	jdff dff_A_AE3LxU6A4_0(.dout(w_dff_A_OrSPGh5J2_0),.din(w_dff_A_AE3LxU6A4_0),.clk(gclk));
	jdff dff_A_OrSPGh5J2_0(.dout(w_dff_A_ZVhf3FjE9_0),.din(w_dff_A_OrSPGh5J2_0),.clk(gclk));
	jdff dff_A_ZVhf3FjE9_0(.dout(w_dff_A_TWjwJyzN4_0),.din(w_dff_A_ZVhf3FjE9_0),.clk(gclk));
	jdff dff_A_TWjwJyzN4_0(.dout(w_dff_A_LJxrGtvv2_0),.din(w_dff_A_TWjwJyzN4_0),.clk(gclk));
	jdff dff_A_LJxrGtvv2_0(.dout(w_dff_A_XfPcqyW10_0),.din(w_dff_A_LJxrGtvv2_0),.clk(gclk));
	jdff dff_A_XfPcqyW10_0(.dout(w_dff_A_BhqegnN72_0),.din(w_dff_A_XfPcqyW10_0),.clk(gclk));
	jdff dff_A_BhqegnN72_0(.dout(w_dff_A_KG2mIWGi2_0),.din(w_dff_A_BhqegnN72_0),.clk(gclk));
	jdff dff_A_KG2mIWGi2_0(.dout(w_dff_A_ZbKwdjpD8_0),.din(w_dff_A_KG2mIWGi2_0),.clk(gclk));
	jdff dff_A_ZbKwdjpD8_0(.dout(w_dff_A_3gFPPP905_0),.din(w_dff_A_ZbKwdjpD8_0),.clk(gclk));
	jdff dff_A_3gFPPP905_0(.dout(w_dff_A_R7GQKwCV2_0),.din(w_dff_A_3gFPPP905_0),.clk(gclk));
	jdff dff_A_R7GQKwCV2_0(.dout(w_dff_A_3WwNRS7P5_0),.din(w_dff_A_R7GQKwCV2_0),.clk(gclk));
	jdff dff_A_3WwNRS7P5_0(.dout(w_dff_A_Bbd6QVDF6_0),.din(w_dff_A_3WwNRS7P5_0),.clk(gclk));
	jdff dff_A_Bbd6QVDF6_0(.dout(w_dff_A_78QWUj3T9_0),.din(w_dff_A_Bbd6QVDF6_0),.clk(gclk));
	jdff dff_A_78QWUj3T9_0(.dout(w_dff_A_RqgrTW7a6_0),.din(w_dff_A_78QWUj3T9_0),.clk(gclk));
	jdff dff_A_RqgrTW7a6_0(.dout(w_dff_A_FKCf7JPf3_0),.din(w_dff_A_RqgrTW7a6_0),.clk(gclk));
	jdff dff_A_FKCf7JPf3_0(.dout(w_dff_A_lYizDufl3_0),.din(w_dff_A_FKCf7JPf3_0),.clk(gclk));
	jdff dff_A_lYizDufl3_0(.dout(w_dff_A_dx2puKVE3_0),.din(w_dff_A_lYizDufl3_0),.clk(gclk));
	jdff dff_A_dx2puKVE3_0(.dout(w_dff_A_dp9TUOam1_0),.din(w_dff_A_dx2puKVE3_0),.clk(gclk));
	jdff dff_A_dp9TUOam1_0(.dout(w_dff_A_x89KjzVS8_0),.din(w_dff_A_dp9TUOam1_0),.clk(gclk));
	jdff dff_A_x89KjzVS8_0(.dout(w_dff_A_5YCHUmkz0_0),.din(w_dff_A_x89KjzVS8_0),.clk(gclk));
	jdff dff_A_5YCHUmkz0_0(.dout(w_dff_A_b8nv0tNG8_0),.din(w_dff_A_5YCHUmkz0_0),.clk(gclk));
	jdff dff_A_b8nv0tNG8_0(.dout(G538),.din(w_dff_A_b8nv0tNG8_0),.clk(gclk));
	jdff dff_A_Z2eAlHCZ6_1(.dout(w_dff_A_bcZdGUgK5_0),.din(w_dff_A_Z2eAlHCZ6_1),.clk(gclk));
	jdff dff_A_bcZdGUgK5_0(.dout(w_dff_A_bj7ynTkS4_0),.din(w_dff_A_bcZdGUgK5_0),.clk(gclk));
	jdff dff_A_bj7ynTkS4_0(.dout(w_dff_A_nrqFXvBo7_0),.din(w_dff_A_bj7ynTkS4_0),.clk(gclk));
	jdff dff_A_nrqFXvBo7_0(.dout(w_dff_A_Uf5PJKEN2_0),.din(w_dff_A_nrqFXvBo7_0),.clk(gclk));
	jdff dff_A_Uf5PJKEN2_0(.dout(w_dff_A_jFRqfUQs8_0),.din(w_dff_A_Uf5PJKEN2_0),.clk(gclk));
	jdff dff_A_jFRqfUQs8_0(.dout(w_dff_A_pLS8XMs39_0),.din(w_dff_A_jFRqfUQs8_0),.clk(gclk));
	jdff dff_A_pLS8XMs39_0(.dout(w_dff_A_oeAUcYnB8_0),.din(w_dff_A_pLS8XMs39_0),.clk(gclk));
	jdff dff_A_oeAUcYnB8_0(.dout(w_dff_A_pfw3LPzS8_0),.din(w_dff_A_oeAUcYnB8_0),.clk(gclk));
	jdff dff_A_pfw3LPzS8_0(.dout(w_dff_A_kWuZW1Dl3_0),.din(w_dff_A_pfw3LPzS8_0),.clk(gclk));
	jdff dff_A_kWuZW1Dl3_0(.dout(w_dff_A_bl5dKVag1_0),.din(w_dff_A_kWuZW1Dl3_0),.clk(gclk));
	jdff dff_A_bl5dKVag1_0(.dout(w_dff_A_ug0wHStv7_0),.din(w_dff_A_bl5dKVag1_0),.clk(gclk));
	jdff dff_A_ug0wHStv7_0(.dout(w_dff_A_3fdMy8mA5_0),.din(w_dff_A_ug0wHStv7_0),.clk(gclk));
	jdff dff_A_3fdMy8mA5_0(.dout(w_dff_A_yWHsVoXZ5_0),.din(w_dff_A_3fdMy8mA5_0),.clk(gclk));
	jdff dff_A_yWHsVoXZ5_0(.dout(w_dff_A_PmVxckrk5_0),.din(w_dff_A_yWHsVoXZ5_0),.clk(gclk));
	jdff dff_A_PmVxckrk5_0(.dout(w_dff_A_cRXroEtT6_0),.din(w_dff_A_PmVxckrk5_0),.clk(gclk));
	jdff dff_A_cRXroEtT6_0(.dout(w_dff_A_3uqfZWDT8_0),.din(w_dff_A_cRXroEtT6_0),.clk(gclk));
	jdff dff_A_3uqfZWDT8_0(.dout(w_dff_A_tTXs6CmS0_0),.din(w_dff_A_3uqfZWDT8_0),.clk(gclk));
	jdff dff_A_tTXs6CmS0_0(.dout(w_dff_A_wvKIbn104_0),.din(w_dff_A_tTXs6CmS0_0),.clk(gclk));
	jdff dff_A_wvKIbn104_0(.dout(w_dff_A_KP4P7DM01_0),.din(w_dff_A_wvKIbn104_0),.clk(gclk));
	jdff dff_A_KP4P7DM01_0(.dout(w_dff_A_eq60TIou0_0),.din(w_dff_A_KP4P7DM01_0),.clk(gclk));
	jdff dff_A_eq60TIou0_0(.dout(w_dff_A_RWgDBVme1_0),.din(w_dff_A_eq60TIou0_0),.clk(gclk));
	jdff dff_A_RWgDBVme1_0(.dout(w_dff_A_ZQVKaTj07_0),.din(w_dff_A_RWgDBVme1_0),.clk(gclk));
	jdff dff_A_ZQVKaTj07_0(.dout(w_dff_A_Zne4Lcdb1_0),.din(w_dff_A_ZQVKaTj07_0),.clk(gclk));
	jdff dff_A_Zne4Lcdb1_0(.dout(w_dff_A_SIoTOpVS0_0),.din(w_dff_A_Zne4Lcdb1_0),.clk(gclk));
	jdff dff_A_SIoTOpVS0_0(.dout(w_dff_A_abRDZ85t4_0),.din(w_dff_A_SIoTOpVS0_0),.clk(gclk));
	jdff dff_A_abRDZ85t4_0(.dout(w_dff_A_ffRooCdc0_0),.din(w_dff_A_abRDZ85t4_0),.clk(gclk));
	jdff dff_A_ffRooCdc0_0(.dout(G536),.din(w_dff_A_ffRooCdc0_0),.clk(gclk));
	jdff dff_A_iSHkyrCa3_1(.dout(w_dff_A_wldKCeuE7_0),.din(w_dff_A_iSHkyrCa3_1),.clk(gclk));
	jdff dff_A_wldKCeuE7_0(.dout(w_dff_A_x5zorZ2N2_0),.din(w_dff_A_wldKCeuE7_0),.clk(gclk));
	jdff dff_A_x5zorZ2N2_0(.dout(w_dff_A_Kl9a4Opx7_0),.din(w_dff_A_x5zorZ2N2_0),.clk(gclk));
	jdff dff_A_Kl9a4Opx7_0(.dout(w_dff_A_FPBSg7oK3_0),.din(w_dff_A_Kl9a4Opx7_0),.clk(gclk));
	jdff dff_A_FPBSg7oK3_0(.dout(w_dff_A_31aDQApI2_0),.din(w_dff_A_FPBSg7oK3_0),.clk(gclk));
	jdff dff_A_31aDQApI2_0(.dout(w_dff_A_ZLxOp7Wy4_0),.din(w_dff_A_31aDQApI2_0),.clk(gclk));
	jdff dff_A_ZLxOp7Wy4_0(.dout(w_dff_A_yeTNJB2x8_0),.din(w_dff_A_ZLxOp7Wy4_0),.clk(gclk));
	jdff dff_A_yeTNJB2x8_0(.dout(w_dff_A_hx8OWPXr2_0),.din(w_dff_A_yeTNJB2x8_0),.clk(gclk));
	jdff dff_A_hx8OWPXr2_0(.dout(w_dff_A_p1jZEzf44_0),.din(w_dff_A_hx8OWPXr2_0),.clk(gclk));
	jdff dff_A_p1jZEzf44_0(.dout(w_dff_A_zVRSIu2W3_0),.din(w_dff_A_p1jZEzf44_0),.clk(gclk));
	jdff dff_A_zVRSIu2W3_0(.dout(w_dff_A_rpwQJ1VC3_0),.din(w_dff_A_zVRSIu2W3_0),.clk(gclk));
	jdff dff_A_rpwQJ1VC3_0(.dout(w_dff_A_fuEY0MX12_0),.din(w_dff_A_rpwQJ1VC3_0),.clk(gclk));
	jdff dff_A_fuEY0MX12_0(.dout(w_dff_A_RqQQatKl2_0),.din(w_dff_A_fuEY0MX12_0),.clk(gclk));
	jdff dff_A_RqQQatKl2_0(.dout(w_dff_A_59zd85SQ5_0),.din(w_dff_A_RqQQatKl2_0),.clk(gclk));
	jdff dff_A_59zd85SQ5_0(.dout(w_dff_A_87c7SQa24_0),.din(w_dff_A_59zd85SQ5_0),.clk(gclk));
	jdff dff_A_87c7SQa24_0(.dout(w_dff_A_Rg5GfciH7_0),.din(w_dff_A_87c7SQa24_0),.clk(gclk));
	jdff dff_A_Rg5GfciH7_0(.dout(w_dff_A_6Nab88Ga3_0),.din(w_dff_A_Rg5GfciH7_0),.clk(gclk));
	jdff dff_A_6Nab88Ga3_0(.dout(w_dff_A_NziXmPSM4_0),.din(w_dff_A_6Nab88Ga3_0),.clk(gclk));
	jdff dff_A_NziXmPSM4_0(.dout(w_dff_A_PvvByTPX0_0),.din(w_dff_A_NziXmPSM4_0),.clk(gclk));
	jdff dff_A_PvvByTPX0_0(.dout(w_dff_A_YUWj64uu6_0),.din(w_dff_A_PvvByTPX0_0),.clk(gclk));
	jdff dff_A_YUWj64uu6_0(.dout(w_dff_A_B0mNSMVQ8_0),.din(w_dff_A_YUWj64uu6_0),.clk(gclk));
	jdff dff_A_B0mNSMVQ8_0(.dout(w_dff_A_UpxY3T6g7_0),.din(w_dff_A_B0mNSMVQ8_0),.clk(gclk));
	jdff dff_A_UpxY3T6g7_0(.dout(w_dff_A_1Dxg9UPR4_0),.din(w_dff_A_UpxY3T6g7_0),.clk(gclk));
	jdff dff_A_1Dxg9UPR4_0(.dout(w_dff_A_uVtiYIfr9_0),.din(w_dff_A_1Dxg9UPR4_0),.clk(gclk));
	jdff dff_A_uVtiYIfr9_0(.dout(w_dff_A_cF4kbO6V7_0),.din(w_dff_A_uVtiYIfr9_0),.clk(gclk));
	jdff dff_A_cF4kbO6V7_0(.dout(w_dff_A_c5Z2LfNb0_0),.din(w_dff_A_cF4kbO6V7_0),.clk(gclk));
	jdff dff_A_c5Z2LfNb0_0(.dout(G534),.din(w_dff_A_c5Z2LfNb0_0),.clk(gclk));
	jdff dff_A_sSU8Nc0v8_1(.dout(w_dff_A_Vd8vT5mw8_0),.din(w_dff_A_sSU8Nc0v8_1),.clk(gclk));
	jdff dff_A_Vd8vT5mw8_0(.dout(w_dff_A_cBRx5XSn9_0),.din(w_dff_A_Vd8vT5mw8_0),.clk(gclk));
	jdff dff_A_cBRx5XSn9_0(.dout(w_dff_A_FD2JDzAe8_0),.din(w_dff_A_cBRx5XSn9_0),.clk(gclk));
	jdff dff_A_FD2JDzAe8_0(.dout(w_dff_A_LXUM44HZ8_0),.din(w_dff_A_FD2JDzAe8_0),.clk(gclk));
	jdff dff_A_LXUM44HZ8_0(.dout(w_dff_A_vFSPL2lh6_0),.din(w_dff_A_LXUM44HZ8_0),.clk(gclk));
	jdff dff_A_vFSPL2lh6_0(.dout(w_dff_A_L8HFXflp7_0),.din(w_dff_A_vFSPL2lh6_0),.clk(gclk));
	jdff dff_A_L8HFXflp7_0(.dout(w_dff_A_bEWmp0Cu1_0),.din(w_dff_A_L8HFXflp7_0),.clk(gclk));
	jdff dff_A_bEWmp0Cu1_0(.dout(w_dff_A_J0Z7YACD8_0),.din(w_dff_A_bEWmp0Cu1_0),.clk(gclk));
	jdff dff_A_J0Z7YACD8_0(.dout(w_dff_A_M6XJNGtz2_0),.din(w_dff_A_J0Z7YACD8_0),.clk(gclk));
	jdff dff_A_M6XJNGtz2_0(.dout(w_dff_A_tSi5QU954_0),.din(w_dff_A_M6XJNGtz2_0),.clk(gclk));
	jdff dff_A_tSi5QU954_0(.dout(w_dff_A_QgUQ6Eev2_0),.din(w_dff_A_tSi5QU954_0),.clk(gclk));
	jdff dff_A_QgUQ6Eev2_0(.dout(w_dff_A_E8URVVgC8_0),.din(w_dff_A_QgUQ6Eev2_0),.clk(gclk));
	jdff dff_A_E8URVVgC8_0(.dout(w_dff_A_8XEOaskD1_0),.din(w_dff_A_E8URVVgC8_0),.clk(gclk));
	jdff dff_A_8XEOaskD1_0(.dout(w_dff_A_vXyC5kyo2_0),.din(w_dff_A_8XEOaskD1_0),.clk(gclk));
	jdff dff_A_vXyC5kyo2_0(.dout(w_dff_A_6Z2n1XN15_0),.din(w_dff_A_vXyC5kyo2_0),.clk(gclk));
	jdff dff_A_6Z2n1XN15_0(.dout(w_dff_A_6Drssuz64_0),.din(w_dff_A_6Z2n1XN15_0),.clk(gclk));
	jdff dff_A_6Drssuz64_0(.dout(w_dff_A_fJfna1mC2_0),.din(w_dff_A_6Drssuz64_0),.clk(gclk));
	jdff dff_A_fJfna1mC2_0(.dout(w_dff_A_AODNTa8Y4_0),.din(w_dff_A_fJfna1mC2_0),.clk(gclk));
	jdff dff_A_AODNTa8Y4_0(.dout(w_dff_A_ohb9x2Yo1_0),.din(w_dff_A_AODNTa8Y4_0),.clk(gclk));
	jdff dff_A_ohb9x2Yo1_0(.dout(w_dff_A_C0DyVrQP4_0),.din(w_dff_A_ohb9x2Yo1_0),.clk(gclk));
	jdff dff_A_C0DyVrQP4_0(.dout(w_dff_A_a3lWSis80_0),.din(w_dff_A_C0DyVrQP4_0),.clk(gclk));
	jdff dff_A_a3lWSis80_0(.dout(w_dff_A_YkBQzBPW6_0),.din(w_dff_A_a3lWSis80_0),.clk(gclk));
	jdff dff_A_YkBQzBPW6_0(.dout(w_dff_A_6ZTM6K6r9_0),.din(w_dff_A_YkBQzBPW6_0),.clk(gclk));
	jdff dff_A_6ZTM6K6r9_0(.dout(w_dff_A_S01Z9pJh6_0),.din(w_dff_A_6ZTM6K6r9_0),.clk(gclk));
	jdff dff_A_S01Z9pJh6_0(.dout(w_dff_A_QvOY3lw56_0),.din(w_dff_A_S01Z9pJh6_0),.clk(gclk));
	jdff dff_A_QvOY3lw56_0(.dout(w_dff_A_CKt7lR0A0_0),.din(w_dff_A_QvOY3lw56_0),.clk(gclk));
	jdff dff_A_CKt7lR0A0_0(.dout(G532),.din(w_dff_A_CKt7lR0A0_0),.clk(gclk));
	jdff dff_A_Of9VtPSQ2_1(.dout(w_dff_A_PaVupGCu8_0),.din(w_dff_A_Of9VtPSQ2_1),.clk(gclk));
	jdff dff_A_PaVupGCu8_0(.dout(w_dff_A_XlXcBwfT2_0),.din(w_dff_A_PaVupGCu8_0),.clk(gclk));
	jdff dff_A_XlXcBwfT2_0(.dout(w_dff_A_QFjQFJ8k0_0),.din(w_dff_A_XlXcBwfT2_0),.clk(gclk));
	jdff dff_A_QFjQFJ8k0_0(.dout(w_dff_A_9q25cNaT0_0),.din(w_dff_A_QFjQFJ8k0_0),.clk(gclk));
	jdff dff_A_9q25cNaT0_0(.dout(w_dff_A_1n0AX2pd9_0),.din(w_dff_A_9q25cNaT0_0),.clk(gclk));
	jdff dff_A_1n0AX2pd9_0(.dout(w_dff_A_moSuIVn52_0),.din(w_dff_A_1n0AX2pd9_0),.clk(gclk));
	jdff dff_A_moSuIVn52_0(.dout(w_dff_A_lppMUx7P5_0),.din(w_dff_A_moSuIVn52_0),.clk(gclk));
	jdff dff_A_lppMUx7P5_0(.dout(w_dff_A_iRztI8lv8_0),.din(w_dff_A_lppMUx7P5_0),.clk(gclk));
	jdff dff_A_iRztI8lv8_0(.dout(w_dff_A_5GR3O3LJ4_0),.din(w_dff_A_iRztI8lv8_0),.clk(gclk));
	jdff dff_A_5GR3O3LJ4_0(.dout(w_dff_A_lifUZu2k3_0),.din(w_dff_A_5GR3O3LJ4_0),.clk(gclk));
	jdff dff_A_lifUZu2k3_0(.dout(w_dff_A_V0qjYcJ06_0),.din(w_dff_A_lifUZu2k3_0),.clk(gclk));
	jdff dff_A_V0qjYcJ06_0(.dout(w_dff_A_TKBCnWwv2_0),.din(w_dff_A_V0qjYcJ06_0),.clk(gclk));
	jdff dff_A_TKBCnWwv2_0(.dout(w_dff_A_JoZRxH766_0),.din(w_dff_A_TKBCnWwv2_0),.clk(gclk));
	jdff dff_A_JoZRxH766_0(.dout(w_dff_A_csyF3vNs4_0),.din(w_dff_A_JoZRxH766_0),.clk(gclk));
	jdff dff_A_csyF3vNs4_0(.dout(w_dff_A_GMMNQUdh9_0),.din(w_dff_A_csyF3vNs4_0),.clk(gclk));
	jdff dff_A_GMMNQUdh9_0(.dout(w_dff_A_DOyVJfzP0_0),.din(w_dff_A_GMMNQUdh9_0),.clk(gclk));
	jdff dff_A_DOyVJfzP0_0(.dout(w_dff_A_JVGGwrzx9_0),.din(w_dff_A_DOyVJfzP0_0),.clk(gclk));
	jdff dff_A_JVGGwrzx9_0(.dout(w_dff_A_vXnlVzB12_0),.din(w_dff_A_JVGGwrzx9_0),.clk(gclk));
	jdff dff_A_vXnlVzB12_0(.dout(w_dff_A_CpPmcKRx0_0),.din(w_dff_A_vXnlVzB12_0),.clk(gclk));
	jdff dff_A_CpPmcKRx0_0(.dout(w_dff_A_eXqyGPMG6_0),.din(w_dff_A_CpPmcKRx0_0),.clk(gclk));
	jdff dff_A_eXqyGPMG6_0(.dout(w_dff_A_k7snMY0i6_0),.din(w_dff_A_eXqyGPMG6_0),.clk(gclk));
	jdff dff_A_k7snMY0i6_0(.dout(w_dff_A_SAhi3Khp4_0),.din(w_dff_A_k7snMY0i6_0),.clk(gclk));
	jdff dff_A_SAhi3Khp4_0(.dout(w_dff_A_78AbOlIQ3_0),.din(w_dff_A_SAhi3Khp4_0),.clk(gclk));
	jdff dff_A_78AbOlIQ3_0(.dout(w_dff_A_wpbIjZ4j4_0),.din(w_dff_A_78AbOlIQ3_0),.clk(gclk));
	jdff dff_A_wpbIjZ4j4_0(.dout(w_dff_A_GbPeiB3i7_0),.din(w_dff_A_wpbIjZ4j4_0),.clk(gclk));
	jdff dff_A_GbPeiB3i7_0(.dout(w_dff_A_89JoPaTU5_0),.din(w_dff_A_GbPeiB3i7_0),.clk(gclk));
	jdff dff_A_89JoPaTU5_0(.dout(G530),.din(w_dff_A_89JoPaTU5_0),.clk(gclk));
	jdff dff_A_ztpM8bzy9_1(.dout(w_dff_A_YTA2BZ5I3_0),.din(w_dff_A_ztpM8bzy9_1),.clk(gclk));
	jdff dff_A_YTA2BZ5I3_0(.dout(w_dff_A_bk2Q4RW43_0),.din(w_dff_A_YTA2BZ5I3_0),.clk(gclk));
	jdff dff_A_bk2Q4RW43_0(.dout(w_dff_A_gsswx0004_0),.din(w_dff_A_bk2Q4RW43_0),.clk(gclk));
	jdff dff_A_gsswx0004_0(.dout(w_dff_A_0xJdXGsN4_0),.din(w_dff_A_gsswx0004_0),.clk(gclk));
	jdff dff_A_0xJdXGsN4_0(.dout(w_dff_A_kZcGVlLW3_0),.din(w_dff_A_0xJdXGsN4_0),.clk(gclk));
	jdff dff_A_kZcGVlLW3_0(.dout(w_dff_A_Iyd1tB144_0),.din(w_dff_A_kZcGVlLW3_0),.clk(gclk));
	jdff dff_A_Iyd1tB144_0(.dout(w_dff_A_yGTBdxCo1_0),.din(w_dff_A_Iyd1tB144_0),.clk(gclk));
	jdff dff_A_yGTBdxCo1_0(.dout(w_dff_A_peRNmo5t8_0),.din(w_dff_A_yGTBdxCo1_0),.clk(gclk));
	jdff dff_A_peRNmo5t8_0(.dout(w_dff_A_MFlndP3E2_0),.din(w_dff_A_peRNmo5t8_0),.clk(gclk));
	jdff dff_A_MFlndP3E2_0(.dout(w_dff_A_fBlaoO5U4_0),.din(w_dff_A_MFlndP3E2_0),.clk(gclk));
	jdff dff_A_fBlaoO5U4_0(.dout(w_dff_A_PtxFxaSy4_0),.din(w_dff_A_fBlaoO5U4_0),.clk(gclk));
	jdff dff_A_PtxFxaSy4_0(.dout(w_dff_A_BSbI8NYr8_0),.din(w_dff_A_PtxFxaSy4_0),.clk(gclk));
	jdff dff_A_BSbI8NYr8_0(.dout(w_dff_A_cavAD3YF0_0),.din(w_dff_A_BSbI8NYr8_0),.clk(gclk));
	jdff dff_A_cavAD3YF0_0(.dout(w_dff_A_2QWqgX0u2_0),.din(w_dff_A_cavAD3YF0_0),.clk(gclk));
	jdff dff_A_2QWqgX0u2_0(.dout(w_dff_A_55crmJhf1_0),.din(w_dff_A_2QWqgX0u2_0),.clk(gclk));
	jdff dff_A_55crmJhf1_0(.dout(w_dff_A_6cnIPeem5_0),.din(w_dff_A_55crmJhf1_0),.clk(gclk));
	jdff dff_A_6cnIPeem5_0(.dout(w_dff_A_iM8ZRctz5_0),.din(w_dff_A_6cnIPeem5_0),.clk(gclk));
	jdff dff_A_iM8ZRctz5_0(.dout(w_dff_A_htYT306Z9_0),.din(w_dff_A_iM8ZRctz5_0),.clk(gclk));
	jdff dff_A_htYT306Z9_0(.dout(w_dff_A_XOSLuCov6_0),.din(w_dff_A_htYT306Z9_0),.clk(gclk));
	jdff dff_A_XOSLuCov6_0(.dout(w_dff_A_UPgu4GZU9_0),.din(w_dff_A_XOSLuCov6_0),.clk(gclk));
	jdff dff_A_UPgu4GZU9_0(.dout(w_dff_A_fwpITZpx7_0),.din(w_dff_A_UPgu4GZU9_0),.clk(gclk));
	jdff dff_A_fwpITZpx7_0(.dout(w_dff_A_SowneOBg8_0),.din(w_dff_A_fwpITZpx7_0),.clk(gclk));
	jdff dff_A_SowneOBg8_0(.dout(w_dff_A_sKnAYa0p6_0),.din(w_dff_A_SowneOBg8_0),.clk(gclk));
	jdff dff_A_sKnAYa0p6_0(.dout(w_dff_A_Qc66GIHC0_0),.din(w_dff_A_sKnAYa0p6_0),.clk(gclk));
	jdff dff_A_Qc66GIHC0_0(.dout(w_dff_A_x1lzBeLR7_0),.din(w_dff_A_Qc66GIHC0_0),.clk(gclk));
	jdff dff_A_x1lzBeLR7_0(.dout(w_dff_A_1wMcQHme5_0),.din(w_dff_A_x1lzBeLR7_0),.clk(gclk));
	jdff dff_A_1wMcQHme5_0(.dout(G528),.din(w_dff_A_1wMcQHme5_0),.clk(gclk));
	jdff dff_A_xlD6j1Zi9_1(.dout(w_dff_A_WFX8D3M31_0),.din(w_dff_A_xlD6j1Zi9_1),.clk(gclk));
	jdff dff_A_WFX8D3M31_0(.dout(w_dff_A_HTsFE5wa1_0),.din(w_dff_A_WFX8D3M31_0),.clk(gclk));
	jdff dff_A_HTsFE5wa1_0(.dout(w_dff_A_JQvnTFgp9_0),.din(w_dff_A_HTsFE5wa1_0),.clk(gclk));
	jdff dff_A_JQvnTFgp9_0(.dout(w_dff_A_QhzKupRl6_0),.din(w_dff_A_JQvnTFgp9_0),.clk(gclk));
	jdff dff_A_QhzKupRl6_0(.dout(w_dff_A_wKWr9rwM1_0),.din(w_dff_A_QhzKupRl6_0),.clk(gclk));
	jdff dff_A_wKWr9rwM1_0(.dout(w_dff_A_r5fBS3tw5_0),.din(w_dff_A_wKWr9rwM1_0),.clk(gclk));
	jdff dff_A_r5fBS3tw5_0(.dout(w_dff_A_U1mWXhPx9_0),.din(w_dff_A_r5fBS3tw5_0),.clk(gclk));
	jdff dff_A_U1mWXhPx9_0(.dout(w_dff_A_BirBGLRM4_0),.din(w_dff_A_U1mWXhPx9_0),.clk(gclk));
	jdff dff_A_BirBGLRM4_0(.dout(w_dff_A_pqlRep9s4_0),.din(w_dff_A_BirBGLRM4_0),.clk(gclk));
	jdff dff_A_pqlRep9s4_0(.dout(w_dff_A_n7UdhcRQ5_0),.din(w_dff_A_pqlRep9s4_0),.clk(gclk));
	jdff dff_A_n7UdhcRQ5_0(.dout(w_dff_A_VFGVCeBI0_0),.din(w_dff_A_n7UdhcRQ5_0),.clk(gclk));
	jdff dff_A_VFGVCeBI0_0(.dout(w_dff_A_NTBFRgI07_0),.din(w_dff_A_VFGVCeBI0_0),.clk(gclk));
	jdff dff_A_NTBFRgI07_0(.dout(w_dff_A_z99r3vfj4_0),.din(w_dff_A_NTBFRgI07_0),.clk(gclk));
	jdff dff_A_z99r3vfj4_0(.dout(w_dff_A_zIxeeIuE7_0),.din(w_dff_A_z99r3vfj4_0),.clk(gclk));
	jdff dff_A_zIxeeIuE7_0(.dout(w_dff_A_uBUobIX13_0),.din(w_dff_A_zIxeeIuE7_0),.clk(gclk));
	jdff dff_A_uBUobIX13_0(.dout(w_dff_A_BMYthtfc2_0),.din(w_dff_A_uBUobIX13_0),.clk(gclk));
	jdff dff_A_BMYthtfc2_0(.dout(w_dff_A_5Z7Y6kIK4_0),.din(w_dff_A_BMYthtfc2_0),.clk(gclk));
	jdff dff_A_5Z7Y6kIK4_0(.dout(w_dff_A_cJi8gR9v5_0),.din(w_dff_A_5Z7Y6kIK4_0),.clk(gclk));
	jdff dff_A_cJi8gR9v5_0(.dout(w_dff_A_3ls0bRIv3_0),.din(w_dff_A_cJi8gR9v5_0),.clk(gclk));
	jdff dff_A_3ls0bRIv3_0(.dout(w_dff_A_VG7KSCzD7_0),.din(w_dff_A_3ls0bRIv3_0),.clk(gclk));
	jdff dff_A_VG7KSCzD7_0(.dout(w_dff_A_Ef51zWPW8_0),.din(w_dff_A_VG7KSCzD7_0),.clk(gclk));
	jdff dff_A_Ef51zWPW8_0(.dout(w_dff_A_i7bXvKhp7_0),.din(w_dff_A_Ef51zWPW8_0),.clk(gclk));
	jdff dff_A_i7bXvKhp7_0(.dout(w_dff_A_oQb5QDZF1_0),.din(w_dff_A_i7bXvKhp7_0),.clk(gclk));
	jdff dff_A_oQb5QDZF1_0(.dout(w_dff_A_ae9vdxwT5_0),.din(w_dff_A_oQb5QDZF1_0),.clk(gclk));
	jdff dff_A_ae9vdxwT5_0(.dout(w_dff_A_6Ks6GMBT4_0),.din(w_dff_A_ae9vdxwT5_0),.clk(gclk));
	jdff dff_A_6Ks6GMBT4_0(.dout(w_dff_A_8fgE9Mbg2_0),.din(w_dff_A_6Ks6GMBT4_0),.clk(gclk));
	jdff dff_A_8fgE9Mbg2_0(.dout(G526),.din(w_dff_A_8fgE9Mbg2_0),.clk(gclk));
	jdff dff_A_HrHW1qMA5_1(.dout(w_dff_A_EUKT3el10_0),.din(w_dff_A_HrHW1qMA5_1),.clk(gclk));
	jdff dff_A_EUKT3el10_0(.dout(w_dff_A_am6qkB8O7_0),.din(w_dff_A_EUKT3el10_0),.clk(gclk));
	jdff dff_A_am6qkB8O7_0(.dout(w_dff_A_Kwxxnfsg7_0),.din(w_dff_A_am6qkB8O7_0),.clk(gclk));
	jdff dff_A_Kwxxnfsg7_0(.dout(w_dff_A_JlJeVVQf2_0),.din(w_dff_A_Kwxxnfsg7_0),.clk(gclk));
	jdff dff_A_JlJeVVQf2_0(.dout(w_dff_A_hmx2HFlt2_0),.din(w_dff_A_JlJeVVQf2_0),.clk(gclk));
	jdff dff_A_hmx2HFlt2_0(.dout(w_dff_A_MCR8gLTZ4_0),.din(w_dff_A_hmx2HFlt2_0),.clk(gclk));
	jdff dff_A_MCR8gLTZ4_0(.dout(w_dff_A_gGznf6Cf6_0),.din(w_dff_A_MCR8gLTZ4_0),.clk(gclk));
	jdff dff_A_gGznf6Cf6_0(.dout(w_dff_A_pVYmjbcm9_0),.din(w_dff_A_gGznf6Cf6_0),.clk(gclk));
	jdff dff_A_pVYmjbcm9_0(.dout(w_dff_A_l1R2MwS65_0),.din(w_dff_A_pVYmjbcm9_0),.clk(gclk));
	jdff dff_A_l1R2MwS65_0(.dout(w_dff_A_wqHZPVXM5_0),.din(w_dff_A_l1R2MwS65_0),.clk(gclk));
	jdff dff_A_wqHZPVXM5_0(.dout(w_dff_A_VBvUbC149_0),.din(w_dff_A_wqHZPVXM5_0),.clk(gclk));
	jdff dff_A_VBvUbC149_0(.dout(w_dff_A_LR9doiFJ6_0),.din(w_dff_A_VBvUbC149_0),.clk(gclk));
	jdff dff_A_LR9doiFJ6_0(.dout(w_dff_A_jykKafmX0_0),.din(w_dff_A_LR9doiFJ6_0),.clk(gclk));
	jdff dff_A_jykKafmX0_0(.dout(w_dff_A_bB9YN1OB8_0),.din(w_dff_A_jykKafmX0_0),.clk(gclk));
	jdff dff_A_bB9YN1OB8_0(.dout(w_dff_A_H1cn6M4r3_0),.din(w_dff_A_bB9YN1OB8_0),.clk(gclk));
	jdff dff_A_H1cn6M4r3_0(.dout(w_dff_A_sAwmomJL8_0),.din(w_dff_A_H1cn6M4r3_0),.clk(gclk));
	jdff dff_A_sAwmomJL8_0(.dout(w_dff_A_8soKMIOm7_0),.din(w_dff_A_sAwmomJL8_0),.clk(gclk));
	jdff dff_A_8soKMIOm7_0(.dout(w_dff_A_0Mvz93Qw7_0),.din(w_dff_A_8soKMIOm7_0),.clk(gclk));
	jdff dff_A_0Mvz93Qw7_0(.dout(w_dff_A_SajoIkiP4_0),.din(w_dff_A_0Mvz93Qw7_0),.clk(gclk));
	jdff dff_A_SajoIkiP4_0(.dout(w_dff_A_Zd97Z9xm1_0),.din(w_dff_A_SajoIkiP4_0),.clk(gclk));
	jdff dff_A_Zd97Z9xm1_0(.dout(w_dff_A_c6dqsFPr5_0),.din(w_dff_A_Zd97Z9xm1_0),.clk(gclk));
	jdff dff_A_c6dqsFPr5_0(.dout(w_dff_A_sTNDFMuf6_0),.din(w_dff_A_c6dqsFPr5_0),.clk(gclk));
	jdff dff_A_sTNDFMuf6_0(.dout(w_dff_A_pXsvqIEo4_0),.din(w_dff_A_sTNDFMuf6_0),.clk(gclk));
	jdff dff_A_pXsvqIEo4_0(.dout(w_dff_A_Hs586TUD0_0),.din(w_dff_A_pXsvqIEo4_0),.clk(gclk));
	jdff dff_A_Hs586TUD0_0(.dout(w_dff_A_HnFBbxtV7_0),.din(w_dff_A_Hs586TUD0_0),.clk(gclk));
	jdff dff_A_HnFBbxtV7_0(.dout(w_dff_A_TxLtrfLw6_0),.din(w_dff_A_HnFBbxtV7_0),.clk(gclk));
	jdff dff_A_TxLtrfLw6_0(.dout(G524),.din(w_dff_A_TxLtrfLw6_0),.clk(gclk));
	jdff dff_A_7HM1DQ839_1(.dout(w_dff_A_slaPthN13_0),.din(w_dff_A_7HM1DQ839_1),.clk(gclk));
	jdff dff_A_slaPthN13_0(.dout(w_dff_A_YGtvSk2a1_0),.din(w_dff_A_slaPthN13_0),.clk(gclk));
	jdff dff_A_YGtvSk2a1_0(.dout(w_dff_A_O3mWxzfZ8_0),.din(w_dff_A_YGtvSk2a1_0),.clk(gclk));
	jdff dff_A_O3mWxzfZ8_0(.dout(w_dff_A_TGV802kf6_0),.din(w_dff_A_O3mWxzfZ8_0),.clk(gclk));
	jdff dff_A_TGV802kf6_0(.dout(w_dff_A_rtzV0jA87_0),.din(w_dff_A_TGV802kf6_0),.clk(gclk));
	jdff dff_A_rtzV0jA87_0(.dout(w_dff_A_Z7vxoIqD7_0),.din(w_dff_A_rtzV0jA87_0),.clk(gclk));
	jdff dff_A_Z7vxoIqD7_0(.dout(w_dff_A_Gq0fpfWh7_0),.din(w_dff_A_Z7vxoIqD7_0),.clk(gclk));
	jdff dff_A_Gq0fpfWh7_0(.dout(w_dff_A_2ttSukOJ0_0),.din(w_dff_A_Gq0fpfWh7_0),.clk(gclk));
	jdff dff_A_2ttSukOJ0_0(.dout(w_dff_A_59GyhNNz7_0),.din(w_dff_A_2ttSukOJ0_0),.clk(gclk));
	jdff dff_A_59GyhNNz7_0(.dout(w_dff_A_tcg9Lg7q2_0),.din(w_dff_A_59GyhNNz7_0),.clk(gclk));
	jdff dff_A_tcg9Lg7q2_0(.dout(w_dff_A_w6j6igK46_0),.din(w_dff_A_tcg9Lg7q2_0),.clk(gclk));
	jdff dff_A_w6j6igK46_0(.dout(w_dff_A_k7MeAYFZ0_0),.din(w_dff_A_w6j6igK46_0),.clk(gclk));
	jdff dff_A_k7MeAYFZ0_0(.dout(w_dff_A_qoPxUERk8_0),.din(w_dff_A_k7MeAYFZ0_0),.clk(gclk));
	jdff dff_A_qoPxUERk8_0(.dout(w_dff_A_L3qDIqAZ0_0),.din(w_dff_A_qoPxUERk8_0),.clk(gclk));
	jdff dff_A_L3qDIqAZ0_0(.dout(w_dff_A_dx3MgIUi8_0),.din(w_dff_A_L3qDIqAZ0_0),.clk(gclk));
	jdff dff_A_dx3MgIUi8_0(.dout(w_dff_A_v0YkqLBK7_0),.din(w_dff_A_dx3MgIUi8_0),.clk(gclk));
	jdff dff_A_v0YkqLBK7_0(.dout(w_dff_A_NoRKP3kl9_0),.din(w_dff_A_v0YkqLBK7_0),.clk(gclk));
	jdff dff_A_NoRKP3kl9_0(.dout(w_dff_A_XBQlT7uD1_0),.din(w_dff_A_NoRKP3kl9_0),.clk(gclk));
	jdff dff_A_XBQlT7uD1_0(.dout(w_dff_A_vxwa7HVZ4_0),.din(w_dff_A_XBQlT7uD1_0),.clk(gclk));
	jdff dff_A_vxwa7HVZ4_0(.dout(w_dff_A_5iPtCTzu0_0),.din(w_dff_A_vxwa7HVZ4_0),.clk(gclk));
	jdff dff_A_5iPtCTzu0_0(.dout(w_dff_A_9CM9qpbB9_0),.din(w_dff_A_5iPtCTzu0_0),.clk(gclk));
	jdff dff_A_9CM9qpbB9_0(.dout(w_dff_A_NpEibPV07_0),.din(w_dff_A_9CM9qpbB9_0),.clk(gclk));
	jdff dff_A_NpEibPV07_0(.dout(w_dff_A_e41xzA2k6_0),.din(w_dff_A_NpEibPV07_0),.clk(gclk));
	jdff dff_A_e41xzA2k6_0(.dout(w_dff_A_2wodT8tr6_0),.din(w_dff_A_e41xzA2k6_0),.clk(gclk));
	jdff dff_A_2wodT8tr6_0(.dout(w_dff_A_7gArp3mZ9_0),.din(w_dff_A_2wodT8tr6_0),.clk(gclk));
	jdff dff_A_7gArp3mZ9_0(.dout(G279),.din(w_dff_A_7gArp3mZ9_0),.clk(gclk));
	jdff dff_A_hGOFpqrP7_1(.dout(w_dff_A_dUxLuROW2_0),.din(w_dff_A_hGOFpqrP7_1),.clk(gclk));
	jdff dff_A_dUxLuROW2_0(.dout(w_dff_A_o4lzmtxy2_0),.din(w_dff_A_dUxLuROW2_0),.clk(gclk));
	jdff dff_A_o4lzmtxy2_0(.dout(w_dff_A_hEimCZFb9_0),.din(w_dff_A_o4lzmtxy2_0),.clk(gclk));
	jdff dff_A_hEimCZFb9_0(.dout(w_dff_A_pxTRyZP67_0),.din(w_dff_A_hEimCZFb9_0),.clk(gclk));
	jdff dff_A_pxTRyZP67_0(.dout(w_dff_A_E8vyQKM88_0),.din(w_dff_A_pxTRyZP67_0),.clk(gclk));
	jdff dff_A_E8vyQKM88_0(.dout(w_dff_A_mCvSdVtJ6_0),.din(w_dff_A_E8vyQKM88_0),.clk(gclk));
	jdff dff_A_mCvSdVtJ6_0(.dout(w_dff_A_LQ4z4i7j8_0),.din(w_dff_A_mCvSdVtJ6_0),.clk(gclk));
	jdff dff_A_LQ4z4i7j8_0(.dout(w_dff_A_KMTyXsnq2_0),.din(w_dff_A_LQ4z4i7j8_0),.clk(gclk));
	jdff dff_A_KMTyXsnq2_0(.dout(w_dff_A_OVpZpCz27_0),.din(w_dff_A_KMTyXsnq2_0),.clk(gclk));
	jdff dff_A_OVpZpCz27_0(.dout(w_dff_A_qGTsLLm01_0),.din(w_dff_A_OVpZpCz27_0),.clk(gclk));
	jdff dff_A_qGTsLLm01_0(.dout(w_dff_A_xHqDG8Uq6_0),.din(w_dff_A_qGTsLLm01_0),.clk(gclk));
	jdff dff_A_xHqDG8Uq6_0(.dout(w_dff_A_raLbnrIY2_0),.din(w_dff_A_xHqDG8Uq6_0),.clk(gclk));
	jdff dff_A_raLbnrIY2_0(.dout(w_dff_A_zwQJNk777_0),.din(w_dff_A_raLbnrIY2_0),.clk(gclk));
	jdff dff_A_zwQJNk777_0(.dout(w_dff_A_mbkooX5s5_0),.din(w_dff_A_zwQJNk777_0),.clk(gclk));
	jdff dff_A_mbkooX5s5_0(.dout(w_dff_A_IHN0Tpaa5_0),.din(w_dff_A_mbkooX5s5_0),.clk(gclk));
	jdff dff_A_IHN0Tpaa5_0(.dout(w_dff_A_Q10zCkCy1_0),.din(w_dff_A_IHN0Tpaa5_0),.clk(gclk));
	jdff dff_A_Q10zCkCy1_0(.dout(w_dff_A_WMtmX2323_0),.din(w_dff_A_Q10zCkCy1_0),.clk(gclk));
	jdff dff_A_WMtmX2323_0(.dout(w_dff_A_shvCxdtb1_0),.din(w_dff_A_WMtmX2323_0),.clk(gclk));
	jdff dff_A_shvCxdtb1_0(.dout(w_dff_A_ET310NpY6_0),.din(w_dff_A_shvCxdtb1_0),.clk(gclk));
	jdff dff_A_ET310NpY6_0(.dout(w_dff_A_xTQCmrBO2_0),.din(w_dff_A_ET310NpY6_0),.clk(gclk));
	jdff dff_A_xTQCmrBO2_0(.dout(w_dff_A_ZnJv6qjc9_0),.din(w_dff_A_xTQCmrBO2_0),.clk(gclk));
	jdff dff_A_ZnJv6qjc9_0(.dout(w_dff_A_KbRCv3KB1_0),.din(w_dff_A_ZnJv6qjc9_0),.clk(gclk));
	jdff dff_A_KbRCv3KB1_0(.dout(w_dff_A_KU2bup1o5_0),.din(w_dff_A_KbRCv3KB1_0),.clk(gclk));
	jdff dff_A_KU2bup1o5_0(.dout(w_dff_A_tapjk4Cf7_0),.din(w_dff_A_KU2bup1o5_0),.clk(gclk));
	jdff dff_A_tapjk4Cf7_0(.dout(w_dff_A_LEd0GuqU0_0),.din(w_dff_A_tapjk4Cf7_0),.clk(gclk));
	jdff dff_A_LEd0GuqU0_0(.dout(w_dff_A_FjMIKdmG3_0),.din(w_dff_A_LEd0GuqU0_0),.clk(gclk));
	jdff dff_A_FjMIKdmG3_0(.dout(G436),.din(w_dff_A_FjMIKdmG3_0),.clk(gclk));
	jdff dff_A_56ni4neV6_1(.dout(w_dff_A_R5Vj1P5q7_0),.din(w_dff_A_56ni4neV6_1),.clk(gclk));
	jdff dff_A_R5Vj1P5q7_0(.dout(w_dff_A_QWr8flty6_0),.din(w_dff_A_R5Vj1P5q7_0),.clk(gclk));
	jdff dff_A_QWr8flty6_0(.dout(w_dff_A_GtW6k2107_0),.din(w_dff_A_QWr8flty6_0),.clk(gclk));
	jdff dff_A_GtW6k2107_0(.dout(w_dff_A_tDq3HhOq7_0),.din(w_dff_A_GtW6k2107_0),.clk(gclk));
	jdff dff_A_tDq3HhOq7_0(.dout(w_dff_A_Q4Xugie34_0),.din(w_dff_A_tDq3HhOq7_0),.clk(gclk));
	jdff dff_A_Q4Xugie34_0(.dout(w_dff_A_JC8BfTjG5_0),.din(w_dff_A_Q4Xugie34_0),.clk(gclk));
	jdff dff_A_JC8BfTjG5_0(.dout(w_dff_A_QiqoRcO32_0),.din(w_dff_A_JC8BfTjG5_0),.clk(gclk));
	jdff dff_A_QiqoRcO32_0(.dout(w_dff_A_6AJtieuS4_0),.din(w_dff_A_QiqoRcO32_0),.clk(gclk));
	jdff dff_A_6AJtieuS4_0(.dout(w_dff_A_XN3Elhhm7_0),.din(w_dff_A_6AJtieuS4_0),.clk(gclk));
	jdff dff_A_XN3Elhhm7_0(.dout(w_dff_A_I4To7Ltp9_0),.din(w_dff_A_XN3Elhhm7_0),.clk(gclk));
	jdff dff_A_I4To7Ltp9_0(.dout(w_dff_A_odBDM5Bu5_0),.din(w_dff_A_I4To7Ltp9_0),.clk(gclk));
	jdff dff_A_odBDM5Bu5_0(.dout(w_dff_A_lfWSCPaD4_0),.din(w_dff_A_odBDM5Bu5_0),.clk(gclk));
	jdff dff_A_lfWSCPaD4_0(.dout(w_dff_A_OS7VMeJR8_0),.din(w_dff_A_lfWSCPaD4_0),.clk(gclk));
	jdff dff_A_OS7VMeJR8_0(.dout(w_dff_A_iTc3HYKq6_0),.din(w_dff_A_OS7VMeJR8_0),.clk(gclk));
	jdff dff_A_iTc3HYKq6_0(.dout(w_dff_A_gosv3Rzz6_0),.din(w_dff_A_iTc3HYKq6_0),.clk(gclk));
	jdff dff_A_gosv3Rzz6_0(.dout(w_dff_A_GNsYfa1T7_0),.din(w_dff_A_gosv3Rzz6_0),.clk(gclk));
	jdff dff_A_GNsYfa1T7_0(.dout(w_dff_A_xRDdIrDJ1_0),.din(w_dff_A_GNsYfa1T7_0),.clk(gclk));
	jdff dff_A_xRDdIrDJ1_0(.dout(w_dff_A_1JdbvD3D8_0),.din(w_dff_A_xRDdIrDJ1_0),.clk(gclk));
	jdff dff_A_1JdbvD3D8_0(.dout(w_dff_A_kvZw8Kj53_0),.din(w_dff_A_1JdbvD3D8_0),.clk(gclk));
	jdff dff_A_kvZw8Kj53_0(.dout(w_dff_A_txsNWER01_0),.din(w_dff_A_kvZw8Kj53_0),.clk(gclk));
	jdff dff_A_txsNWER01_0(.dout(w_dff_A_Td4NXJIu5_0),.din(w_dff_A_txsNWER01_0),.clk(gclk));
	jdff dff_A_Td4NXJIu5_0(.dout(w_dff_A_z69aD0NZ1_0),.din(w_dff_A_Td4NXJIu5_0),.clk(gclk));
	jdff dff_A_z69aD0NZ1_0(.dout(w_dff_A_xbqszPMa7_0),.din(w_dff_A_z69aD0NZ1_0),.clk(gclk));
	jdff dff_A_xbqszPMa7_0(.dout(w_dff_A_UPOudb9i6_0),.din(w_dff_A_xbqszPMa7_0),.clk(gclk));
	jdff dff_A_UPOudb9i6_0(.dout(w_dff_A_ChtXKLQr0_0),.din(w_dff_A_UPOudb9i6_0),.clk(gclk));
	jdff dff_A_ChtXKLQr0_0(.dout(w_dff_A_I0FN6nyc1_0),.din(w_dff_A_ChtXKLQr0_0),.clk(gclk));
	jdff dff_A_I0FN6nyc1_0(.dout(G478),.din(w_dff_A_I0FN6nyc1_0),.clk(gclk));
	jdff dff_A_sAMargQa3_1(.dout(w_dff_A_m2BflVSL6_0),.din(w_dff_A_sAMargQa3_1),.clk(gclk));
	jdff dff_A_m2BflVSL6_0(.dout(w_dff_A_fIraQLK07_0),.din(w_dff_A_m2BflVSL6_0),.clk(gclk));
	jdff dff_A_fIraQLK07_0(.dout(w_dff_A_A66Nf7J08_0),.din(w_dff_A_fIraQLK07_0),.clk(gclk));
	jdff dff_A_A66Nf7J08_0(.dout(w_dff_A_GA9WXupi3_0),.din(w_dff_A_A66Nf7J08_0),.clk(gclk));
	jdff dff_A_GA9WXupi3_0(.dout(w_dff_A_oOoin8CA8_0),.din(w_dff_A_GA9WXupi3_0),.clk(gclk));
	jdff dff_A_oOoin8CA8_0(.dout(w_dff_A_ciEf2wi22_0),.din(w_dff_A_oOoin8CA8_0),.clk(gclk));
	jdff dff_A_ciEf2wi22_0(.dout(w_dff_A_s1gJ98CE2_0),.din(w_dff_A_ciEf2wi22_0),.clk(gclk));
	jdff dff_A_s1gJ98CE2_0(.dout(w_dff_A_ZKWJVfOw4_0),.din(w_dff_A_s1gJ98CE2_0),.clk(gclk));
	jdff dff_A_ZKWJVfOw4_0(.dout(w_dff_A_PCAAxjED7_0),.din(w_dff_A_ZKWJVfOw4_0),.clk(gclk));
	jdff dff_A_PCAAxjED7_0(.dout(w_dff_A_OzdCoDdg1_0),.din(w_dff_A_PCAAxjED7_0),.clk(gclk));
	jdff dff_A_OzdCoDdg1_0(.dout(w_dff_A_zvVnal4D5_0),.din(w_dff_A_OzdCoDdg1_0),.clk(gclk));
	jdff dff_A_zvVnal4D5_0(.dout(w_dff_A_VLfBbvTj2_0),.din(w_dff_A_zvVnal4D5_0),.clk(gclk));
	jdff dff_A_VLfBbvTj2_0(.dout(w_dff_A_LXGn4nOU4_0),.din(w_dff_A_VLfBbvTj2_0),.clk(gclk));
	jdff dff_A_LXGn4nOU4_0(.dout(w_dff_A_EgLkMdKR0_0),.din(w_dff_A_LXGn4nOU4_0),.clk(gclk));
	jdff dff_A_EgLkMdKR0_0(.dout(w_dff_A_zADllPJ25_0),.din(w_dff_A_EgLkMdKR0_0),.clk(gclk));
	jdff dff_A_zADllPJ25_0(.dout(w_dff_A_SHtKDGAd4_0),.din(w_dff_A_zADllPJ25_0),.clk(gclk));
	jdff dff_A_SHtKDGAd4_0(.dout(w_dff_A_QivZwlB87_0),.din(w_dff_A_SHtKDGAd4_0),.clk(gclk));
	jdff dff_A_QivZwlB87_0(.dout(w_dff_A_awhgtQZa6_0),.din(w_dff_A_QivZwlB87_0),.clk(gclk));
	jdff dff_A_awhgtQZa6_0(.dout(w_dff_A_dMILZV8T8_0),.din(w_dff_A_awhgtQZa6_0),.clk(gclk));
	jdff dff_A_dMILZV8T8_0(.dout(w_dff_A_ISwco8zU4_0),.din(w_dff_A_dMILZV8T8_0),.clk(gclk));
	jdff dff_A_ISwco8zU4_0(.dout(w_dff_A_cEsRmd8r1_0),.din(w_dff_A_ISwco8zU4_0),.clk(gclk));
	jdff dff_A_cEsRmd8r1_0(.dout(w_dff_A_z3NkZ1Zz8_0),.din(w_dff_A_cEsRmd8r1_0),.clk(gclk));
	jdff dff_A_z3NkZ1Zz8_0(.dout(w_dff_A_nxkUreNI3_0),.din(w_dff_A_z3NkZ1Zz8_0),.clk(gclk));
	jdff dff_A_nxkUreNI3_0(.dout(w_dff_A_ewcPRaoT8_0),.din(w_dff_A_nxkUreNI3_0),.clk(gclk));
	jdff dff_A_ewcPRaoT8_0(.dout(w_dff_A_hr1ayws02_0),.din(w_dff_A_ewcPRaoT8_0),.clk(gclk));
	jdff dff_A_hr1ayws02_0(.dout(w_dff_A_oUyfBQsb8_0),.din(w_dff_A_hr1ayws02_0),.clk(gclk));
	jdff dff_A_oUyfBQsb8_0(.dout(G522),.din(w_dff_A_oUyfBQsb8_0),.clk(gclk));
	jdff dff_A_OZMI4Ga77_2(.dout(w_dff_A_n4ToBhTj3_0),.din(w_dff_A_OZMI4Ga77_2),.clk(gclk));
	jdff dff_A_n4ToBhTj3_0(.dout(w_dff_A_Oexla1mg8_0),.din(w_dff_A_n4ToBhTj3_0),.clk(gclk));
	jdff dff_A_Oexla1mg8_0(.dout(w_dff_A_n8YxaAaE9_0),.din(w_dff_A_Oexla1mg8_0),.clk(gclk));
	jdff dff_A_n8YxaAaE9_0(.dout(w_dff_A_GH91YwdK7_0),.din(w_dff_A_n8YxaAaE9_0),.clk(gclk));
	jdff dff_A_GH91YwdK7_0(.dout(w_dff_A_Oslq1ZHc2_0),.din(w_dff_A_GH91YwdK7_0),.clk(gclk));
	jdff dff_A_Oslq1ZHc2_0(.dout(w_dff_A_czGeNeLo8_0),.din(w_dff_A_Oslq1ZHc2_0),.clk(gclk));
	jdff dff_A_czGeNeLo8_0(.dout(w_dff_A_XpI3nqT53_0),.din(w_dff_A_czGeNeLo8_0),.clk(gclk));
	jdff dff_A_XpI3nqT53_0(.dout(w_dff_A_axDLYPgR4_0),.din(w_dff_A_XpI3nqT53_0),.clk(gclk));
	jdff dff_A_axDLYPgR4_0(.dout(w_dff_A_x1gIkGE00_0),.din(w_dff_A_axDLYPgR4_0),.clk(gclk));
	jdff dff_A_x1gIkGE00_0(.dout(w_dff_A_UY1Vl4A43_0),.din(w_dff_A_x1gIkGE00_0),.clk(gclk));
	jdff dff_A_UY1Vl4A43_0(.dout(w_dff_A_kUuPiZCT1_0),.din(w_dff_A_UY1Vl4A43_0),.clk(gclk));
	jdff dff_A_kUuPiZCT1_0(.dout(w_dff_A_LNZgwBAN9_0),.din(w_dff_A_kUuPiZCT1_0),.clk(gclk));
	jdff dff_A_LNZgwBAN9_0(.dout(w_dff_A_NcwNWXL39_0),.din(w_dff_A_LNZgwBAN9_0),.clk(gclk));
	jdff dff_A_NcwNWXL39_0(.dout(w_dff_A_UHTWrzuF2_0),.din(w_dff_A_NcwNWXL39_0),.clk(gclk));
	jdff dff_A_UHTWrzuF2_0(.dout(w_dff_A_PEaEW2Jp1_0),.din(w_dff_A_UHTWrzuF2_0),.clk(gclk));
	jdff dff_A_PEaEW2Jp1_0(.dout(w_dff_A_l6MeY4mM7_0),.din(w_dff_A_PEaEW2Jp1_0),.clk(gclk));
	jdff dff_A_l6MeY4mM7_0(.dout(w_dff_A_gUTgeiKU5_0),.din(w_dff_A_l6MeY4mM7_0),.clk(gclk));
	jdff dff_A_gUTgeiKU5_0(.dout(w_dff_A_xu9AsHLe2_0),.din(w_dff_A_gUTgeiKU5_0),.clk(gclk));
	jdff dff_A_xu9AsHLe2_0(.dout(w_dff_A_pSXltQpo6_0),.din(w_dff_A_xu9AsHLe2_0),.clk(gclk));
	jdff dff_A_pSXltQpo6_0(.dout(w_dff_A_5F2korNF4_0),.din(w_dff_A_pSXltQpo6_0),.clk(gclk));
	jdff dff_A_5F2korNF4_0(.dout(w_dff_A_6TPs2gno4_0),.din(w_dff_A_5F2korNF4_0),.clk(gclk));
	jdff dff_A_6TPs2gno4_0(.dout(w_dff_A_p6bj0BKZ8_0),.din(w_dff_A_6TPs2gno4_0),.clk(gclk));
	jdff dff_A_p6bj0BKZ8_0(.dout(w_dff_A_QQO17DdI0_0),.din(w_dff_A_p6bj0BKZ8_0),.clk(gclk));
	jdff dff_A_QQO17DdI0_0(.dout(w_dff_A_0Cs0mKtd3_0),.din(w_dff_A_QQO17DdI0_0),.clk(gclk));
	jdff dff_A_0Cs0mKtd3_0(.dout(w_dff_A_rJCz512O4_0),.din(w_dff_A_0Cs0mKtd3_0),.clk(gclk));
	jdff dff_A_rJCz512O4_0(.dout(G402),.din(w_dff_A_rJCz512O4_0),.clk(gclk));
	jdff dff_A_SGEwqHKw4_1(.dout(w_dff_A_WCjFhd9u8_0),.din(w_dff_A_SGEwqHKw4_1),.clk(gclk));
	jdff dff_A_WCjFhd9u8_0(.dout(w_dff_A_ii5WTJeC7_0),.din(w_dff_A_WCjFhd9u8_0),.clk(gclk));
	jdff dff_A_ii5WTJeC7_0(.dout(w_dff_A_gTJrP7ff0_0),.din(w_dff_A_ii5WTJeC7_0),.clk(gclk));
	jdff dff_A_gTJrP7ff0_0(.dout(w_dff_A_jeZVLKG73_0),.din(w_dff_A_gTJrP7ff0_0),.clk(gclk));
	jdff dff_A_jeZVLKG73_0(.dout(w_dff_A_FZAJqJdk5_0),.din(w_dff_A_jeZVLKG73_0),.clk(gclk));
	jdff dff_A_FZAJqJdk5_0(.dout(w_dff_A_p3KIA5Tw7_0),.din(w_dff_A_FZAJqJdk5_0),.clk(gclk));
	jdff dff_A_p3KIA5Tw7_0(.dout(w_dff_A_mQUyU7to6_0),.din(w_dff_A_p3KIA5Tw7_0),.clk(gclk));
	jdff dff_A_mQUyU7to6_0(.dout(w_dff_A_yVf3E3Uu5_0),.din(w_dff_A_mQUyU7to6_0),.clk(gclk));
	jdff dff_A_yVf3E3Uu5_0(.dout(w_dff_A_jl7uMHUv9_0),.din(w_dff_A_yVf3E3Uu5_0),.clk(gclk));
	jdff dff_A_jl7uMHUv9_0(.dout(w_dff_A_gvJjEoSf3_0),.din(w_dff_A_jl7uMHUv9_0),.clk(gclk));
	jdff dff_A_gvJjEoSf3_0(.dout(w_dff_A_EcJpwJNy2_0),.din(w_dff_A_gvJjEoSf3_0),.clk(gclk));
	jdff dff_A_EcJpwJNy2_0(.dout(w_dff_A_Bq18wGRS4_0),.din(w_dff_A_EcJpwJNy2_0),.clk(gclk));
	jdff dff_A_Bq18wGRS4_0(.dout(w_dff_A_XBwn5tcC5_0),.din(w_dff_A_Bq18wGRS4_0),.clk(gclk));
	jdff dff_A_XBwn5tcC5_0(.dout(w_dff_A_qo4tyB984_0),.din(w_dff_A_XBwn5tcC5_0),.clk(gclk));
	jdff dff_A_qo4tyB984_0(.dout(w_dff_A_LYkosXUf5_0),.din(w_dff_A_qo4tyB984_0),.clk(gclk));
	jdff dff_A_LYkosXUf5_0(.dout(w_dff_A_u5We17kT1_0),.din(w_dff_A_LYkosXUf5_0),.clk(gclk));
	jdff dff_A_u5We17kT1_0(.dout(w_dff_A_yTQLrgwF3_0),.din(w_dff_A_u5We17kT1_0),.clk(gclk));
	jdff dff_A_yTQLrgwF3_0(.dout(w_dff_A_M8GcD04g3_0),.din(w_dff_A_yTQLrgwF3_0),.clk(gclk));
	jdff dff_A_M8GcD04g3_0(.dout(w_dff_A_xWHtDopP6_0),.din(w_dff_A_M8GcD04g3_0),.clk(gclk));
	jdff dff_A_xWHtDopP6_0(.dout(w_dff_A_vxrV3DXv5_0),.din(w_dff_A_xWHtDopP6_0),.clk(gclk));
	jdff dff_A_vxrV3DXv5_0(.dout(w_dff_A_81JwQljV9_0),.din(w_dff_A_vxrV3DXv5_0),.clk(gclk));
	jdff dff_A_81JwQljV9_0(.dout(w_dff_A_jbDTqvTB5_0),.din(w_dff_A_81JwQljV9_0),.clk(gclk));
	jdff dff_A_jbDTqvTB5_0(.dout(w_dff_A_sIt0Y2zZ6_0),.din(w_dff_A_jbDTqvTB5_0),.clk(gclk));
	jdff dff_A_sIt0Y2zZ6_0(.dout(G404),.din(w_dff_A_sIt0Y2zZ6_0),.clk(gclk));
	jdff dff_A_J25vNCWP8_1(.dout(w_dff_A_BkuQIf3C9_0),.din(w_dff_A_J25vNCWP8_1),.clk(gclk));
	jdff dff_A_BkuQIf3C9_0(.dout(w_dff_A_bUcGTBD71_0),.din(w_dff_A_BkuQIf3C9_0),.clk(gclk));
	jdff dff_A_bUcGTBD71_0(.dout(w_dff_A_oH689uGw3_0),.din(w_dff_A_bUcGTBD71_0),.clk(gclk));
	jdff dff_A_oH689uGw3_0(.dout(w_dff_A_mwC6lZBd9_0),.din(w_dff_A_oH689uGw3_0),.clk(gclk));
	jdff dff_A_mwC6lZBd9_0(.dout(w_dff_A_XUmI1UNj4_0),.din(w_dff_A_mwC6lZBd9_0),.clk(gclk));
	jdff dff_A_XUmI1UNj4_0(.dout(w_dff_A_cU0zo3iN6_0),.din(w_dff_A_XUmI1UNj4_0),.clk(gclk));
	jdff dff_A_cU0zo3iN6_0(.dout(w_dff_A_az6wwGDe5_0),.din(w_dff_A_cU0zo3iN6_0),.clk(gclk));
	jdff dff_A_az6wwGDe5_0(.dout(w_dff_A_zALtfvep0_0),.din(w_dff_A_az6wwGDe5_0),.clk(gclk));
	jdff dff_A_zALtfvep0_0(.dout(w_dff_A_PEtQF9Zs2_0),.din(w_dff_A_zALtfvep0_0),.clk(gclk));
	jdff dff_A_PEtQF9Zs2_0(.dout(w_dff_A_h7BfEb0S1_0),.din(w_dff_A_PEtQF9Zs2_0),.clk(gclk));
	jdff dff_A_h7BfEb0S1_0(.dout(w_dff_A_WCYLutiH9_0),.din(w_dff_A_h7BfEb0S1_0),.clk(gclk));
	jdff dff_A_WCYLutiH9_0(.dout(w_dff_A_PMMcucqa7_0),.din(w_dff_A_WCYLutiH9_0),.clk(gclk));
	jdff dff_A_PMMcucqa7_0(.dout(w_dff_A_wKNWm0Im7_0),.din(w_dff_A_PMMcucqa7_0),.clk(gclk));
	jdff dff_A_wKNWm0Im7_0(.dout(w_dff_A_drcZnwBR6_0),.din(w_dff_A_wKNWm0Im7_0),.clk(gclk));
	jdff dff_A_drcZnwBR6_0(.dout(w_dff_A_QT2ZJ9WB0_0),.din(w_dff_A_drcZnwBR6_0),.clk(gclk));
	jdff dff_A_QT2ZJ9WB0_0(.dout(w_dff_A_SlAP4dXO4_0),.din(w_dff_A_QT2ZJ9WB0_0),.clk(gclk));
	jdff dff_A_SlAP4dXO4_0(.dout(w_dff_A_DfKGz3FT7_0),.din(w_dff_A_SlAP4dXO4_0),.clk(gclk));
	jdff dff_A_DfKGz3FT7_0(.dout(w_dff_A_2KAjtvHe8_0),.din(w_dff_A_DfKGz3FT7_0),.clk(gclk));
	jdff dff_A_2KAjtvHe8_0(.dout(w_dff_A_TEfYyzUs7_0),.din(w_dff_A_2KAjtvHe8_0),.clk(gclk));
	jdff dff_A_TEfYyzUs7_0(.dout(w_dff_A_mbFJ79w41_0),.din(w_dff_A_TEfYyzUs7_0),.clk(gclk));
	jdff dff_A_mbFJ79w41_0(.dout(w_dff_A_gs4EZLeV6_0),.din(w_dff_A_mbFJ79w41_0),.clk(gclk));
	jdff dff_A_gs4EZLeV6_0(.dout(w_dff_A_sVf5JINW3_0),.din(w_dff_A_gs4EZLeV6_0),.clk(gclk));
	jdff dff_A_sVf5JINW3_0(.dout(w_dff_A_CAdzPeq91_0),.din(w_dff_A_sVf5JINW3_0),.clk(gclk));
	jdff dff_A_CAdzPeq91_0(.dout(G406),.din(w_dff_A_CAdzPeq91_0),.clk(gclk));
	jdff dff_A_6zPirW7D7_1(.dout(w_dff_A_swJY6FON9_0),.din(w_dff_A_6zPirW7D7_1),.clk(gclk));
	jdff dff_A_swJY6FON9_0(.dout(w_dff_A_xaDhx7ov5_0),.din(w_dff_A_swJY6FON9_0),.clk(gclk));
	jdff dff_A_xaDhx7ov5_0(.dout(w_dff_A_UpdGSlPz2_0),.din(w_dff_A_xaDhx7ov5_0),.clk(gclk));
	jdff dff_A_UpdGSlPz2_0(.dout(w_dff_A_G6xJVx3O5_0),.din(w_dff_A_UpdGSlPz2_0),.clk(gclk));
	jdff dff_A_G6xJVx3O5_0(.dout(w_dff_A_rObM40D18_0),.din(w_dff_A_G6xJVx3O5_0),.clk(gclk));
	jdff dff_A_rObM40D18_0(.dout(w_dff_A_Lpa9olqb6_0),.din(w_dff_A_rObM40D18_0),.clk(gclk));
	jdff dff_A_Lpa9olqb6_0(.dout(w_dff_A_oQOAjhPd0_0),.din(w_dff_A_Lpa9olqb6_0),.clk(gclk));
	jdff dff_A_oQOAjhPd0_0(.dout(w_dff_A_abVQBL915_0),.din(w_dff_A_oQOAjhPd0_0),.clk(gclk));
	jdff dff_A_abVQBL915_0(.dout(w_dff_A_pxsPcSCM4_0),.din(w_dff_A_abVQBL915_0),.clk(gclk));
	jdff dff_A_pxsPcSCM4_0(.dout(w_dff_A_x2WDlAoM1_0),.din(w_dff_A_pxsPcSCM4_0),.clk(gclk));
	jdff dff_A_x2WDlAoM1_0(.dout(w_dff_A_yyUvmJvo3_0),.din(w_dff_A_x2WDlAoM1_0),.clk(gclk));
	jdff dff_A_yyUvmJvo3_0(.dout(w_dff_A_z5wRCZwn6_0),.din(w_dff_A_yyUvmJvo3_0),.clk(gclk));
	jdff dff_A_z5wRCZwn6_0(.dout(w_dff_A_Ce7shpOP1_0),.din(w_dff_A_z5wRCZwn6_0),.clk(gclk));
	jdff dff_A_Ce7shpOP1_0(.dout(w_dff_A_XUqDQT3z8_0),.din(w_dff_A_Ce7shpOP1_0),.clk(gclk));
	jdff dff_A_XUqDQT3z8_0(.dout(w_dff_A_pSZMH1zl9_0),.din(w_dff_A_XUqDQT3z8_0),.clk(gclk));
	jdff dff_A_pSZMH1zl9_0(.dout(w_dff_A_BmIQnGyM4_0),.din(w_dff_A_pSZMH1zl9_0),.clk(gclk));
	jdff dff_A_BmIQnGyM4_0(.dout(w_dff_A_RPpeSkqQ1_0),.din(w_dff_A_BmIQnGyM4_0),.clk(gclk));
	jdff dff_A_RPpeSkqQ1_0(.dout(w_dff_A_yPmdc3T84_0),.din(w_dff_A_RPpeSkqQ1_0),.clk(gclk));
	jdff dff_A_yPmdc3T84_0(.dout(w_dff_A_WIOpWlE71_0),.din(w_dff_A_yPmdc3T84_0),.clk(gclk));
	jdff dff_A_WIOpWlE71_0(.dout(w_dff_A_7IuK3eYW4_0),.din(w_dff_A_WIOpWlE71_0),.clk(gclk));
	jdff dff_A_7IuK3eYW4_0(.dout(w_dff_A_T6cX8LI91_0),.din(w_dff_A_7IuK3eYW4_0),.clk(gclk));
	jdff dff_A_T6cX8LI91_0(.dout(w_dff_A_vKhBUJMz9_0),.din(w_dff_A_T6cX8LI91_0),.clk(gclk));
	jdff dff_A_vKhBUJMz9_0(.dout(w_dff_A_Wh0cJCrl6_0),.din(w_dff_A_vKhBUJMz9_0),.clk(gclk));
	jdff dff_A_Wh0cJCrl6_0(.dout(G408),.din(w_dff_A_Wh0cJCrl6_0),.clk(gclk));
	jdff dff_A_NzXdC8ZK7_1(.dout(w_dff_A_pn4KMOni0_0),.din(w_dff_A_NzXdC8ZK7_1),.clk(gclk));
	jdff dff_A_pn4KMOni0_0(.dout(w_dff_A_QifoiltK8_0),.din(w_dff_A_pn4KMOni0_0),.clk(gclk));
	jdff dff_A_QifoiltK8_0(.dout(w_dff_A_aHvpLeWs7_0),.din(w_dff_A_QifoiltK8_0),.clk(gclk));
	jdff dff_A_aHvpLeWs7_0(.dout(w_dff_A_BRpil0t39_0),.din(w_dff_A_aHvpLeWs7_0),.clk(gclk));
	jdff dff_A_BRpil0t39_0(.dout(w_dff_A_CVCOIa1X8_0),.din(w_dff_A_BRpil0t39_0),.clk(gclk));
	jdff dff_A_CVCOIa1X8_0(.dout(w_dff_A_5fxMVuoV7_0),.din(w_dff_A_CVCOIa1X8_0),.clk(gclk));
	jdff dff_A_5fxMVuoV7_0(.dout(w_dff_A_O7mUvSFn5_0),.din(w_dff_A_5fxMVuoV7_0),.clk(gclk));
	jdff dff_A_O7mUvSFn5_0(.dout(w_dff_A_PLsjc6cc5_0),.din(w_dff_A_O7mUvSFn5_0),.clk(gclk));
	jdff dff_A_PLsjc6cc5_0(.dout(w_dff_A_xg6GiZUB3_0),.din(w_dff_A_PLsjc6cc5_0),.clk(gclk));
	jdff dff_A_xg6GiZUB3_0(.dout(w_dff_A_VuT2Z1Wn9_0),.din(w_dff_A_xg6GiZUB3_0),.clk(gclk));
	jdff dff_A_VuT2Z1Wn9_0(.dout(w_dff_A_BFwDx8kC1_0),.din(w_dff_A_VuT2Z1Wn9_0),.clk(gclk));
	jdff dff_A_BFwDx8kC1_0(.dout(w_dff_A_TcA86cJC5_0),.din(w_dff_A_BFwDx8kC1_0),.clk(gclk));
	jdff dff_A_TcA86cJC5_0(.dout(w_dff_A_5qZROEJn9_0),.din(w_dff_A_TcA86cJC5_0),.clk(gclk));
	jdff dff_A_5qZROEJn9_0(.dout(w_dff_A_753z8Nll3_0),.din(w_dff_A_5qZROEJn9_0),.clk(gclk));
	jdff dff_A_753z8Nll3_0(.dout(w_dff_A_7quX9Zo90_0),.din(w_dff_A_753z8Nll3_0),.clk(gclk));
	jdff dff_A_7quX9Zo90_0(.dout(w_dff_A_kf8qv9KM2_0),.din(w_dff_A_7quX9Zo90_0),.clk(gclk));
	jdff dff_A_kf8qv9KM2_0(.dout(w_dff_A_nQgJ8EyW4_0),.din(w_dff_A_kf8qv9KM2_0),.clk(gclk));
	jdff dff_A_nQgJ8EyW4_0(.dout(w_dff_A_uCx06Mjp9_0),.din(w_dff_A_nQgJ8EyW4_0),.clk(gclk));
	jdff dff_A_uCx06Mjp9_0(.dout(w_dff_A_C7IdZ9tA1_0),.din(w_dff_A_uCx06Mjp9_0),.clk(gclk));
	jdff dff_A_C7IdZ9tA1_0(.dout(w_dff_A_TovBFwZG6_0),.din(w_dff_A_C7IdZ9tA1_0),.clk(gclk));
	jdff dff_A_TovBFwZG6_0(.dout(w_dff_A_mKFrwWiS7_0),.din(w_dff_A_TovBFwZG6_0),.clk(gclk));
	jdff dff_A_mKFrwWiS7_0(.dout(w_dff_A_h8GdkFMM1_0),.din(w_dff_A_mKFrwWiS7_0),.clk(gclk));
	jdff dff_A_h8GdkFMM1_0(.dout(w_dff_A_9t41dwCj1_0),.din(w_dff_A_h8GdkFMM1_0),.clk(gclk));
	jdff dff_A_9t41dwCj1_0(.dout(G410),.din(w_dff_A_9t41dwCj1_0),.clk(gclk));
	jdff dff_A_15oUKSIM7_1(.dout(w_dff_A_rV1SaM8m4_0),.din(w_dff_A_15oUKSIM7_1),.clk(gclk));
	jdff dff_A_rV1SaM8m4_0(.dout(w_dff_A_7kl6Y6b35_0),.din(w_dff_A_rV1SaM8m4_0),.clk(gclk));
	jdff dff_A_7kl6Y6b35_0(.dout(w_dff_A_OkPxIsGP7_0),.din(w_dff_A_7kl6Y6b35_0),.clk(gclk));
	jdff dff_A_OkPxIsGP7_0(.dout(w_dff_A_V7Cwdbaz4_0),.din(w_dff_A_OkPxIsGP7_0),.clk(gclk));
	jdff dff_A_V7Cwdbaz4_0(.dout(w_dff_A_GQS04JOe1_0),.din(w_dff_A_V7Cwdbaz4_0),.clk(gclk));
	jdff dff_A_GQS04JOe1_0(.dout(w_dff_A_D4vzyFZz8_0),.din(w_dff_A_GQS04JOe1_0),.clk(gclk));
	jdff dff_A_D4vzyFZz8_0(.dout(w_dff_A_Elk81OvA1_0),.din(w_dff_A_D4vzyFZz8_0),.clk(gclk));
	jdff dff_A_Elk81OvA1_0(.dout(w_dff_A_ZetmPexk7_0),.din(w_dff_A_Elk81OvA1_0),.clk(gclk));
	jdff dff_A_ZetmPexk7_0(.dout(w_dff_A_v9me7U372_0),.din(w_dff_A_ZetmPexk7_0),.clk(gclk));
	jdff dff_A_v9me7U372_0(.dout(w_dff_A_z6KKGThk2_0),.din(w_dff_A_v9me7U372_0),.clk(gclk));
	jdff dff_A_z6KKGThk2_0(.dout(w_dff_A_bDpofzk43_0),.din(w_dff_A_z6KKGThk2_0),.clk(gclk));
	jdff dff_A_bDpofzk43_0(.dout(w_dff_A_weCviYfJ6_0),.din(w_dff_A_bDpofzk43_0),.clk(gclk));
	jdff dff_A_weCviYfJ6_0(.dout(w_dff_A_JFX9dQ9t1_0),.din(w_dff_A_weCviYfJ6_0),.clk(gclk));
	jdff dff_A_JFX9dQ9t1_0(.dout(w_dff_A_JWPMpJnY7_0),.din(w_dff_A_JFX9dQ9t1_0),.clk(gclk));
	jdff dff_A_JWPMpJnY7_0(.dout(w_dff_A_XwDr6baQ2_0),.din(w_dff_A_JWPMpJnY7_0),.clk(gclk));
	jdff dff_A_XwDr6baQ2_0(.dout(w_dff_A_xbKGdnls8_0),.din(w_dff_A_XwDr6baQ2_0),.clk(gclk));
	jdff dff_A_xbKGdnls8_0(.dout(w_dff_A_UYM8VOwr7_0),.din(w_dff_A_xbKGdnls8_0),.clk(gclk));
	jdff dff_A_UYM8VOwr7_0(.dout(w_dff_A_025twQV96_0),.din(w_dff_A_UYM8VOwr7_0),.clk(gclk));
	jdff dff_A_025twQV96_0(.dout(w_dff_A_YPyFNXBa0_0),.din(w_dff_A_025twQV96_0),.clk(gclk));
	jdff dff_A_YPyFNXBa0_0(.dout(w_dff_A_sQrSQiKd4_0),.din(w_dff_A_YPyFNXBa0_0),.clk(gclk));
	jdff dff_A_sQrSQiKd4_0(.dout(w_dff_A_JV1PFuuH3_0),.din(w_dff_A_sQrSQiKd4_0),.clk(gclk));
	jdff dff_A_JV1PFuuH3_0(.dout(w_dff_A_BaP4BC360_0),.din(w_dff_A_JV1PFuuH3_0),.clk(gclk));
	jdff dff_A_BaP4BC360_0(.dout(w_dff_A_wiyjVIP52_0),.din(w_dff_A_BaP4BC360_0),.clk(gclk));
	jdff dff_A_wiyjVIP52_0(.dout(w_dff_A_IVaOQYXD7_0),.din(w_dff_A_wiyjVIP52_0),.clk(gclk));
	jdff dff_A_IVaOQYXD7_0(.dout(w_dff_A_Ld4fhGte8_0),.din(w_dff_A_IVaOQYXD7_0),.clk(gclk));
	jdff dff_A_Ld4fhGte8_0(.dout(w_dff_A_V2Sjjcjm2_0),.din(w_dff_A_Ld4fhGte8_0),.clk(gclk));
	jdff dff_A_V2Sjjcjm2_0(.dout(G432),.din(w_dff_A_V2Sjjcjm2_0),.clk(gclk));
	jdff dff_A_FqMa6rxn5_1(.dout(w_dff_A_KxnVtkzY6_0),.din(w_dff_A_FqMa6rxn5_1),.clk(gclk));
	jdff dff_A_KxnVtkzY6_0(.dout(w_dff_A_jKIs852d6_0),.din(w_dff_A_KxnVtkzY6_0),.clk(gclk));
	jdff dff_A_jKIs852d6_0(.dout(w_dff_A_XOUuMD9C8_0),.din(w_dff_A_jKIs852d6_0),.clk(gclk));
	jdff dff_A_XOUuMD9C8_0(.dout(w_dff_A_ivjdorIe2_0),.din(w_dff_A_XOUuMD9C8_0),.clk(gclk));
	jdff dff_A_ivjdorIe2_0(.dout(w_dff_A_Ge9Q8Dmh1_0),.din(w_dff_A_ivjdorIe2_0),.clk(gclk));
	jdff dff_A_Ge9Q8Dmh1_0(.dout(w_dff_A_Lavmisb85_0),.din(w_dff_A_Ge9Q8Dmh1_0),.clk(gclk));
	jdff dff_A_Lavmisb85_0(.dout(w_dff_A_dUCZCv3R3_0),.din(w_dff_A_Lavmisb85_0),.clk(gclk));
	jdff dff_A_dUCZCv3R3_0(.dout(w_dff_A_BKJ67eLy5_0),.din(w_dff_A_dUCZCv3R3_0),.clk(gclk));
	jdff dff_A_BKJ67eLy5_0(.dout(w_dff_A_VjEOSWgg9_0),.din(w_dff_A_BKJ67eLy5_0),.clk(gclk));
	jdff dff_A_VjEOSWgg9_0(.dout(w_dff_A_9JNxaAIb7_0),.din(w_dff_A_VjEOSWgg9_0),.clk(gclk));
	jdff dff_A_9JNxaAIb7_0(.dout(w_dff_A_QrGPKV7s9_0),.din(w_dff_A_9JNxaAIb7_0),.clk(gclk));
	jdff dff_A_QrGPKV7s9_0(.dout(w_dff_A_fmQ1iOxl0_0),.din(w_dff_A_QrGPKV7s9_0),.clk(gclk));
	jdff dff_A_fmQ1iOxl0_0(.dout(w_dff_A_X4n5i12Y8_0),.din(w_dff_A_fmQ1iOxl0_0),.clk(gclk));
	jdff dff_A_X4n5i12Y8_0(.dout(w_dff_A_MsuKoody8_0),.din(w_dff_A_X4n5i12Y8_0),.clk(gclk));
	jdff dff_A_MsuKoody8_0(.dout(w_dff_A_YBAXKzI72_0),.din(w_dff_A_MsuKoody8_0),.clk(gclk));
	jdff dff_A_YBAXKzI72_0(.dout(w_dff_A_H96RlYwA5_0),.din(w_dff_A_YBAXKzI72_0),.clk(gclk));
	jdff dff_A_H96RlYwA5_0(.dout(w_dff_A_G1RvKQWe0_0),.din(w_dff_A_H96RlYwA5_0),.clk(gclk));
	jdff dff_A_G1RvKQWe0_0(.dout(w_dff_A_pgDFHFYF3_0),.din(w_dff_A_G1RvKQWe0_0),.clk(gclk));
	jdff dff_A_pgDFHFYF3_0(.dout(w_dff_A_023pmYW58_0),.din(w_dff_A_pgDFHFYF3_0),.clk(gclk));
	jdff dff_A_023pmYW58_0(.dout(w_dff_A_9ZZai5io4_0),.din(w_dff_A_023pmYW58_0),.clk(gclk));
	jdff dff_A_9ZZai5io4_0(.dout(w_dff_A_UNB6st835_0),.din(w_dff_A_9ZZai5io4_0),.clk(gclk));
	jdff dff_A_UNB6st835_0(.dout(w_dff_A_YZMP34Wf4_0),.din(w_dff_A_UNB6st835_0),.clk(gclk));
	jdff dff_A_YZMP34Wf4_0(.dout(w_dff_A_hWw4vhj30_0),.din(w_dff_A_YZMP34Wf4_0),.clk(gclk));
	jdff dff_A_hWw4vhj30_0(.dout(w_dff_A_PFUIfVnV2_0),.din(w_dff_A_hWw4vhj30_0),.clk(gclk));
	jdff dff_A_PFUIfVnV2_0(.dout(w_dff_A_n8HpsUKG8_0),.din(w_dff_A_PFUIfVnV2_0),.clk(gclk));
	jdff dff_A_n8HpsUKG8_0(.dout(w_dff_A_mMNe0m2b8_0),.din(w_dff_A_n8HpsUKG8_0),.clk(gclk));
	jdff dff_A_mMNe0m2b8_0(.dout(G446),.din(w_dff_A_mMNe0m2b8_0),.clk(gclk));
	jdff dff_A_uzDJ9L3F8_2(.dout(w_dff_A_DFczi5Cy3_0),.din(w_dff_A_uzDJ9L3F8_2),.clk(gclk));
	jdff dff_A_DFczi5Cy3_0(.dout(w_dff_A_bEg6PutY6_0),.din(w_dff_A_DFczi5Cy3_0),.clk(gclk));
	jdff dff_A_bEg6PutY6_0(.dout(w_dff_A_dXqxX0Ng7_0),.din(w_dff_A_bEg6PutY6_0),.clk(gclk));
	jdff dff_A_dXqxX0Ng7_0(.dout(w_dff_A_OaP8C8ge8_0),.din(w_dff_A_dXqxX0Ng7_0),.clk(gclk));
	jdff dff_A_OaP8C8ge8_0(.dout(w_dff_A_9zm7ukga8_0),.din(w_dff_A_OaP8C8ge8_0),.clk(gclk));
	jdff dff_A_9zm7ukga8_0(.dout(w_dff_A_nqJcaAhV4_0),.din(w_dff_A_9zm7ukga8_0),.clk(gclk));
	jdff dff_A_nqJcaAhV4_0(.dout(w_dff_A_pMluvbk79_0),.din(w_dff_A_nqJcaAhV4_0),.clk(gclk));
	jdff dff_A_pMluvbk79_0(.dout(w_dff_A_twUM6LXZ7_0),.din(w_dff_A_pMluvbk79_0),.clk(gclk));
	jdff dff_A_twUM6LXZ7_0(.dout(w_dff_A_9rL0ABE20_0),.din(w_dff_A_twUM6LXZ7_0),.clk(gclk));
	jdff dff_A_9rL0ABE20_0(.dout(w_dff_A_s4WBAphs3_0),.din(w_dff_A_9rL0ABE20_0),.clk(gclk));
	jdff dff_A_s4WBAphs3_0(.dout(w_dff_A_LS2lmRPx5_0),.din(w_dff_A_s4WBAphs3_0),.clk(gclk));
	jdff dff_A_LS2lmRPx5_0(.dout(w_dff_A_Zk1oiQwt5_0),.din(w_dff_A_LS2lmRPx5_0),.clk(gclk));
	jdff dff_A_Zk1oiQwt5_0(.dout(w_dff_A_ETPYdynt7_0),.din(w_dff_A_Zk1oiQwt5_0),.clk(gclk));
	jdff dff_A_ETPYdynt7_0(.dout(w_dff_A_r7tX8glB7_0),.din(w_dff_A_ETPYdynt7_0),.clk(gclk));
	jdff dff_A_r7tX8glB7_0(.dout(w_dff_A_WEqtMSzi1_0),.din(w_dff_A_r7tX8glB7_0),.clk(gclk));
	jdff dff_A_WEqtMSzi1_0(.dout(w_dff_A_Llu0yBvG8_0),.din(w_dff_A_WEqtMSzi1_0),.clk(gclk));
	jdff dff_A_Llu0yBvG8_0(.dout(w_dff_A_5Lk3h4vZ4_0),.din(w_dff_A_Llu0yBvG8_0),.clk(gclk));
	jdff dff_A_5Lk3h4vZ4_0(.dout(w_dff_A_xUPpYiNs0_0),.din(w_dff_A_5Lk3h4vZ4_0),.clk(gclk));
	jdff dff_A_xUPpYiNs0_0(.dout(w_dff_A_Cl87TgwO7_0),.din(w_dff_A_xUPpYiNs0_0),.clk(gclk));
	jdff dff_A_Cl87TgwO7_0(.dout(w_dff_A_u2QYT7gV9_0),.din(w_dff_A_Cl87TgwO7_0),.clk(gclk));
	jdff dff_A_u2QYT7gV9_0(.dout(w_dff_A_QtTE4g8n0_0),.din(w_dff_A_u2QYT7gV9_0),.clk(gclk));
	jdff dff_A_QtTE4g8n0_0(.dout(w_dff_A_PRGlECK02_0),.din(w_dff_A_QtTE4g8n0_0),.clk(gclk));
	jdff dff_A_PRGlECK02_0(.dout(w_dff_A_zIwBq5YE5_0),.din(w_dff_A_PRGlECK02_0),.clk(gclk));
	jdff dff_A_zIwBq5YE5_0(.dout(w_dff_A_S3BlpmZH6_0),.din(w_dff_A_zIwBq5YE5_0),.clk(gclk));
	jdff dff_A_S3BlpmZH6_0(.dout(G284),.din(w_dff_A_S3BlpmZH6_0),.clk(gclk));
	jdff dff_A_x6qNQfhM0_1(.dout(w_dff_A_ollMUi7J4_0),.din(w_dff_A_x6qNQfhM0_1),.clk(gclk));
	jdff dff_A_ollMUi7J4_0(.dout(w_dff_A_X0LsElUZ2_0),.din(w_dff_A_ollMUi7J4_0),.clk(gclk));
	jdff dff_A_X0LsElUZ2_0(.dout(w_dff_A_wcaTEiE82_0),.din(w_dff_A_X0LsElUZ2_0),.clk(gclk));
	jdff dff_A_wcaTEiE82_0(.dout(w_dff_A_KqAr2P2W4_0),.din(w_dff_A_wcaTEiE82_0),.clk(gclk));
	jdff dff_A_KqAr2P2W4_0(.dout(w_dff_A_eDd6yCzQ0_0),.din(w_dff_A_KqAr2P2W4_0),.clk(gclk));
	jdff dff_A_eDd6yCzQ0_0(.dout(w_dff_A_9qFENikU0_0),.din(w_dff_A_eDd6yCzQ0_0),.clk(gclk));
	jdff dff_A_9qFENikU0_0(.dout(w_dff_A_L5KKnOQC6_0),.din(w_dff_A_9qFENikU0_0),.clk(gclk));
	jdff dff_A_L5KKnOQC6_0(.dout(w_dff_A_aCaHXAuk5_0),.din(w_dff_A_L5KKnOQC6_0),.clk(gclk));
	jdff dff_A_aCaHXAuk5_0(.dout(w_dff_A_wqYAbRbZ0_0),.din(w_dff_A_aCaHXAuk5_0),.clk(gclk));
	jdff dff_A_wqYAbRbZ0_0(.dout(w_dff_A_e9AUNY7E1_0),.din(w_dff_A_wqYAbRbZ0_0),.clk(gclk));
	jdff dff_A_e9AUNY7E1_0(.dout(w_dff_A_1wqVMcOx7_0),.din(w_dff_A_e9AUNY7E1_0),.clk(gclk));
	jdff dff_A_1wqVMcOx7_0(.dout(w_dff_A_BTrkWGRa5_0),.din(w_dff_A_1wqVMcOx7_0),.clk(gclk));
	jdff dff_A_BTrkWGRa5_0(.dout(w_dff_A_X2GkVYsK2_0),.din(w_dff_A_BTrkWGRa5_0),.clk(gclk));
	jdff dff_A_X2GkVYsK2_0(.dout(w_dff_A_GFRScXE64_0),.din(w_dff_A_X2GkVYsK2_0),.clk(gclk));
	jdff dff_A_GFRScXE64_0(.dout(w_dff_A_1dymERuQ2_0),.din(w_dff_A_GFRScXE64_0),.clk(gclk));
	jdff dff_A_1dymERuQ2_0(.dout(w_dff_A_p9IXDxTq3_0),.din(w_dff_A_1dymERuQ2_0),.clk(gclk));
	jdff dff_A_p9IXDxTq3_0(.dout(w_dff_A_tuNHTqcG6_0),.din(w_dff_A_p9IXDxTq3_0),.clk(gclk));
	jdff dff_A_tuNHTqcG6_0(.dout(w_dff_A_3ac1XEpq5_0),.din(w_dff_A_tuNHTqcG6_0),.clk(gclk));
	jdff dff_A_3ac1XEpq5_0(.dout(w_dff_A_QZyhMrW18_0),.din(w_dff_A_3ac1XEpq5_0),.clk(gclk));
	jdff dff_A_QZyhMrW18_0(.dout(w_dff_A_IYyvNjoF3_0),.din(w_dff_A_QZyhMrW18_0),.clk(gclk));
	jdff dff_A_IYyvNjoF3_0(.dout(w_dff_A_BRmrOcId6_0),.din(w_dff_A_IYyvNjoF3_0),.clk(gclk));
	jdff dff_A_BRmrOcId6_0(.dout(w_dff_A_8CFnMlOT8_0),.din(w_dff_A_BRmrOcId6_0),.clk(gclk));
	jdff dff_A_8CFnMlOT8_0(.dout(w_dff_A_aDB1Pwe90_0),.din(w_dff_A_8CFnMlOT8_0),.clk(gclk));
	jdff dff_A_aDB1Pwe90_0(.dout(w_dff_A_qCtZmxzF6_0),.din(w_dff_A_aDB1Pwe90_0),.clk(gclk));
	jdff dff_A_qCtZmxzF6_0(.dout(w_dff_A_DGYT1Nro3_0),.din(w_dff_A_qCtZmxzF6_0),.clk(gclk));
	jdff dff_A_DGYT1Nro3_0(.dout(G286),.din(w_dff_A_DGYT1Nro3_0),.clk(gclk));
	jdff dff_A_WJXAWJxz0_2(.dout(w_dff_A_9v7UGhX00_0),.din(w_dff_A_WJXAWJxz0_2),.clk(gclk));
	jdff dff_A_9v7UGhX00_0(.dout(w_dff_A_oxGZTti87_0),.din(w_dff_A_9v7UGhX00_0),.clk(gclk));
	jdff dff_A_oxGZTti87_0(.dout(w_dff_A_mCco08TC7_0),.din(w_dff_A_oxGZTti87_0),.clk(gclk));
	jdff dff_A_mCco08TC7_0(.dout(w_dff_A_bKH8u0f57_0),.din(w_dff_A_mCco08TC7_0),.clk(gclk));
	jdff dff_A_bKH8u0f57_0(.dout(w_dff_A_jg48mVdB2_0),.din(w_dff_A_bKH8u0f57_0),.clk(gclk));
	jdff dff_A_jg48mVdB2_0(.dout(w_dff_A_QUDuOjuV3_0),.din(w_dff_A_jg48mVdB2_0),.clk(gclk));
	jdff dff_A_QUDuOjuV3_0(.dout(w_dff_A_nSXQXXB28_0),.din(w_dff_A_QUDuOjuV3_0),.clk(gclk));
	jdff dff_A_nSXQXXB28_0(.dout(w_dff_A_LzFWpX7k9_0),.din(w_dff_A_nSXQXXB28_0),.clk(gclk));
	jdff dff_A_LzFWpX7k9_0(.dout(w_dff_A_ebub0rke1_0),.din(w_dff_A_LzFWpX7k9_0),.clk(gclk));
	jdff dff_A_ebub0rke1_0(.dout(w_dff_A_6JScAf7E9_0),.din(w_dff_A_ebub0rke1_0),.clk(gclk));
	jdff dff_A_6JScAf7E9_0(.dout(w_dff_A_4kH7o5Ex6_0),.din(w_dff_A_6JScAf7E9_0),.clk(gclk));
	jdff dff_A_4kH7o5Ex6_0(.dout(w_dff_A_2jrSi9ya2_0),.din(w_dff_A_4kH7o5Ex6_0),.clk(gclk));
	jdff dff_A_2jrSi9ya2_0(.dout(w_dff_A_GuTi3FQS0_0),.din(w_dff_A_2jrSi9ya2_0),.clk(gclk));
	jdff dff_A_GuTi3FQS0_0(.dout(w_dff_A_7y81J92U0_0),.din(w_dff_A_GuTi3FQS0_0),.clk(gclk));
	jdff dff_A_7y81J92U0_0(.dout(w_dff_A_X7yeDhV98_0),.din(w_dff_A_7y81J92U0_0),.clk(gclk));
	jdff dff_A_X7yeDhV98_0(.dout(w_dff_A_csa7LC7O1_0),.din(w_dff_A_X7yeDhV98_0),.clk(gclk));
	jdff dff_A_csa7LC7O1_0(.dout(w_dff_A_SKKFc0Vi4_0),.din(w_dff_A_csa7LC7O1_0),.clk(gclk));
	jdff dff_A_SKKFc0Vi4_0(.dout(w_dff_A_09K4opfR6_0),.din(w_dff_A_SKKFc0Vi4_0),.clk(gclk));
	jdff dff_A_09K4opfR6_0(.dout(w_dff_A_3lBFDCFr9_0),.din(w_dff_A_09K4opfR6_0),.clk(gclk));
	jdff dff_A_3lBFDCFr9_0(.dout(w_dff_A_Ih72erhV1_0),.din(w_dff_A_3lBFDCFr9_0),.clk(gclk));
	jdff dff_A_Ih72erhV1_0(.dout(w_dff_A_p6Swh93x4_0),.din(w_dff_A_Ih72erhV1_0),.clk(gclk));
	jdff dff_A_p6Swh93x4_0(.dout(w_dff_A_FN558NaB2_0),.din(w_dff_A_p6Swh93x4_0),.clk(gclk));
	jdff dff_A_FN558NaB2_0(.dout(w_dff_A_u6HZNBGs2_0),.din(w_dff_A_FN558NaB2_0),.clk(gclk));
	jdff dff_A_u6HZNBGs2_0(.dout(w_dff_A_CFzJVzmR7_0),.din(w_dff_A_u6HZNBGs2_0),.clk(gclk));
	jdff dff_A_CFzJVzmR7_0(.dout(G289),.din(w_dff_A_CFzJVzmR7_0),.clk(gclk));
	jdff dff_A_1X4oNfns3_2(.dout(w_dff_A_ZhBZZBgd5_0),.din(w_dff_A_1X4oNfns3_2),.clk(gclk));
	jdff dff_A_ZhBZZBgd5_0(.dout(w_dff_A_vrlc2RpM8_0),.din(w_dff_A_ZhBZZBgd5_0),.clk(gclk));
	jdff dff_A_vrlc2RpM8_0(.dout(w_dff_A_FHLtO33B0_0),.din(w_dff_A_vrlc2RpM8_0),.clk(gclk));
	jdff dff_A_FHLtO33B0_0(.dout(w_dff_A_S1NCbxzt8_0),.din(w_dff_A_FHLtO33B0_0),.clk(gclk));
	jdff dff_A_S1NCbxzt8_0(.dout(w_dff_A_4GfGlBmI2_0),.din(w_dff_A_S1NCbxzt8_0),.clk(gclk));
	jdff dff_A_4GfGlBmI2_0(.dout(w_dff_A_QsgpELKQ1_0),.din(w_dff_A_4GfGlBmI2_0),.clk(gclk));
	jdff dff_A_QsgpELKQ1_0(.dout(w_dff_A_aSXJcHvT5_0),.din(w_dff_A_QsgpELKQ1_0),.clk(gclk));
	jdff dff_A_aSXJcHvT5_0(.dout(w_dff_A_vs7GopUV6_0),.din(w_dff_A_aSXJcHvT5_0),.clk(gclk));
	jdff dff_A_vs7GopUV6_0(.dout(w_dff_A_iLrHKmur7_0),.din(w_dff_A_vs7GopUV6_0),.clk(gclk));
	jdff dff_A_iLrHKmur7_0(.dout(w_dff_A_gLVJe10g9_0),.din(w_dff_A_iLrHKmur7_0),.clk(gclk));
	jdff dff_A_gLVJe10g9_0(.dout(w_dff_A_jDKNfY3o5_0),.din(w_dff_A_gLVJe10g9_0),.clk(gclk));
	jdff dff_A_jDKNfY3o5_0(.dout(w_dff_A_JPKXI0BP3_0),.din(w_dff_A_jDKNfY3o5_0),.clk(gclk));
	jdff dff_A_JPKXI0BP3_0(.dout(w_dff_A_c7dIGHaN4_0),.din(w_dff_A_JPKXI0BP3_0),.clk(gclk));
	jdff dff_A_c7dIGHaN4_0(.dout(w_dff_A_CaoHIMYz3_0),.din(w_dff_A_c7dIGHaN4_0),.clk(gclk));
	jdff dff_A_CaoHIMYz3_0(.dout(w_dff_A_GfySpbKj7_0),.din(w_dff_A_CaoHIMYz3_0),.clk(gclk));
	jdff dff_A_GfySpbKj7_0(.dout(w_dff_A_pttiFYPI0_0),.din(w_dff_A_GfySpbKj7_0),.clk(gclk));
	jdff dff_A_pttiFYPI0_0(.dout(w_dff_A_Ihyh8TZa7_0),.din(w_dff_A_pttiFYPI0_0),.clk(gclk));
	jdff dff_A_Ihyh8TZa7_0(.dout(w_dff_A_Rw2f9WHk6_0),.din(w_dff_A_Ihyh8TZa7_0),.clk(gclk));
	jdff dff_A_Rw2f9WHk6_0(.dout(w_dff_A_NDiYw3uO0_0),.din(w_dff_A_Rw2f9WHk6_0),.clk(gclk));
	jdff dff_A_NDiYw3uO0_0(.dout(w_dff_A_0ni8nRFt8_0),.din(w_dff_A_NDiYw3uO0_0),.clk(gclk));
	jdff dff_A_0ni8nRFt8_0(.dout(w_dff_A_KYjym8t20_0),.din(w_dff_A_0ni8nRFt8_0),.clk(gclk));
	jdff dff_A_KYjym8t20_0(.dout(w_dff_A_06FEdL4F2_0),.din(w_dff_A_KYjym8t20_0),.clk(gclk));
	jdff dff_A_06FEdL4F2_0(.dout(w_dff_A_u5juNdXE1_0),.din(w_dff_A_06FEdL4F2_0),.clk(gclk));
	jdff dff_A_u5juNdXE1_0(.dout(G292),.din(w_dff_A_u5juNdXE1_0),.clk(gclk));
	jdff dff_A_BPLu96TO4_1(.dout(w_dff_A_B2WkPzf57_0),.din(w_dff_A_BPLu96TO4_1),.clk(gclk));
	jdff dff_A_B2WkPzf57_0(.dout(w_dff_A_LmjfS6Hj3_0),.din(w_dff_A_B2WkPzf57_0),.clk(gclk));
	jdff dff_A_LmjfS6Hj3_0(.dout(w_dff_A_IhR9W28s1_0),.din(w_dff_A_LmjfS6Hj3_0),.clk(gclk));
	jdff dff_A_IhR9W28s1_0(.dout(w_dff_A_raudKgbW1_0),.din(w_dff_A_IhR9W28s1_0),.clk(gclk));
	jdff dff_A_raudKgbW1_0(.dout(w_dff_A_oW8Kzrdr5_0),.din(w_dff_A_raudKgbW1_0),.clk(gclk));
	jdff dff_A_oW8Kzrdr5_0(.dout(w_dff_A_FDFv2MiR7_0),.din(w_dff_A_oW8Kzrdr5_0),.clk(gclk));
	jdff dff_A_FDFv2MiR7_0(.dout(w_dff_A_PM3C1zbs7_0),.din(w_dff_A_FDFv2MiR7_0),.clk(gclk));
	jdff dff_A_PM3C1zbs7_0(.dout(w_dff_A_WZBNOmlY7_0),.din(w_dff_A_PM3C1zbs7_0),.clk(gclk));
	jdff dff_A_WZBNOmlY7_0(.dout(w_dff_A_fXJ3jRIS6_0),.din(w_dff_A_WZBNOmlY7_0),.clk(gclk));
	jdff dff_A_fXJ3jRIS6_0(.dout(w_dff_A_XSXfg8e04_0),.din(w_dff_A_fXJ3jRIS6_0),.clk(gclk));
	jdff dff_A_XSXfg8e04_0(.dout(w_dff_A_8nILk8zQ7_0),.din(w_dff_A_XSXfg8e04_0),.clk(gclk));
	jdff dff_A_8nILk8zQ7_0(.dout(w_dff_A_TGsacql63_0),.din(w_dff_A_8nILk8zQ7_0),.clk(gclk));
	jdff dff_A_TGsacql63_0(.dout(w_dff_A_0B6ixsIV9_0),.din(w_dff_A_TGsacql63_0),.clk(gclk));
	jdff dff_A_0B6ixsIV9_0(.dout(w_dff_A_wG9agYSb6_0),.din(w_dff_A_0B6ixsIV9_0),.clk(gclk));
	jdff dff_A_wG9agYSb6_0(.dout(w_dff_A_cYleF8c42_0),.din(w_dff_A_wG9agYSb6_0),.clk(gclk));
	jdff dff_A_cYleF8c42_0(.dout(w_dff_A_P1KVfEbT6_0),.din(w_dff_A_cYleF8c42_0),.clk(gclk));
	jdff dff_A_P1KVfEbT6_0(.dout(w_dff_A_agUPurLr9_0),.din(w_dff_A_P1KVfEbT6_0),.clk(gclk));
	jdff dff_A_agUPurLr9_0(.dout(w_dff_A_ZbzVtPQr4_0),.din(w_dff_A_agUPurLr9_0),.clk(gclk));
	jdff dff_A_ZbzVtPQr4_0(.dout(w_dff_A_0OFphQqV0_0),.din(w_dff_A_ZbzVtPQr4_0),.clk(gclk));
	jdff dff_A_0OFphQqV0_0(.dout(w_dff_A_MmzAFegM3_0),.din(w_dff_A_0OFphQqV0_0),.clk(gclk));
	jdff dff_A_MmzAFegM3_0(.dout(w_dff_A_paIQBduA2_0),.din(w_dff_A_MmzAFegM3_0),.clk(gclk));
	jdff dff_A_paIQBduA2_0(.dout(w_dff_A_fmRShWyS8_0),.din(w_dff_A_paIQBduA2_0),.clk(gclk));
	jdff dff_A_fmRShWyS8_0(.dout(w_dff_A_FntllQ3v5_0),.din(w_dff_A_fmRShWyS8_0),.clk(gclk));
	jdff dff_A_FntllQ3v5_0(.dout(w_dff_A_rfdWNpQA6_0),.din(w_dff_A_FntllQ3v5_0),.clk(gclk));
	jdff dff_A_rfdWNpQA6_0(.dout(w_dff_A_HTNiFf2C7_0),.din(w_dff_A_rfdWNpQA6_0),.clk(gclk));
	jdff dff_A_HTNiFf2C7_0(.dout(G341),.din(w_dff_A_HTNiFf2C7_0),.clk(gclk));
	jdff dff_A_GX6m9gnD6_2(.dout(w_dff_A_Ex4fV9vq1_0),.din(w_dff_A_GX6m9gnD6_2),.clk(gclk));
	jdff dff_A_Ex4fV9vq1_0(.dout(w_dff_A_WBUNxKt92_0),.din(w_dff_A_Ex4fV9vq1_0),.clk(gclk));
	jdff dff_A_WBUNxKt92_0(.dout(w_dff_A_sygmZ1Ir3_0),.din(w_dff_A_WBUNxKt92_0),.clk(gclk));
	jdff dff_A_sygmZ1Ir3_0(.dout(w_dff_A_9PWgd9sw8_0),.din(w_dff_A_sygmZ1Ir3_0),.clk(gclk));
	jdff dff_A_9PWgd9sw8_0(.dout(w_dff_A_IP5rtZp00_0),.din(w_dff_A_9PWgd9sw8_0),.clk(gclk));
	jdff dff_A_IP5rtZp00_0(.dout(w_dff_A_LUsZfq3G6_0),.din(w_dff_A_IP5rtZp00_0),.clk(gclk));
	jdff dff_A_LUsZfq3G6_0(.dout(w_dff_A_Bg0OjLYG3_0),.din(w_dff_A_LUsZfq3G6_0),.clk(gclk));
	jdff dff_A_Bg0OjLYG3_0(.dout(w_dff_A_lPcWjmYV2_0),.din(w_dff_A_Bg0OjLYG3_0),.clk(gclk));
	jdff dff_A_lPcWjmYV2_0(.dout(w_dff_A_isYsmanl4_0),.din(w_dff_A_lPcWjmYV2_0),.clk(gclk));
	jdff dff_A_isYsmanl4_0(.dout(w_dff_A_DMsNzaUo0_0),.din(w_dff_A_isYsmanl4_0),.clk(gclk));
	jdff dff_A_DMsNzaUo0_0(.dout(w_dff_A_beOfWyyP7_0),.din(w_dff_A_DMsNzaUo0_0),.clk(gclk));
	jdff dff_A_beOfWyyP7_0(.dout(w_dff_A_ry638cHX8_0),.din(w_dff_A_beOfWyyP7_0),.clk(gclk));
	jdff dff_A_ry638cHX8_0(.dout(w_dff_A_4Wvqgncc0_0),.din(w_dff_A_ry638cHX8_0),.clk(gclk));
	jdff dff_A_4Wvqgncc0_0(.dout(w_dff_A_EYJczFbM6_0),.din(w_dff_A_4Wvqgncc0_0),.clk(gclk));
	jdff dff_A_EYJczFbM6_0(.dout(w_dff_A_Xr9txrBs0_0),.din(w_dff_A_EYJczFbM6_0),.clk(gclk));
	jdff dff_A_Xr9txrBs0_0(.dout(w_dff_A_SfdAQZmb0_0),.din(w_dff_A_Xr9txrBs0_0),.clk(gclk));
	jdff dff_A_SfdAQZmb0_0(.dout(w_dff_A_98Jc2vF24_0),.din(w_dff_A_SfdAQZmb0_0),.clk(gclk));
	jdff dff_A_98Jc2vF24_0(.dout(w_dff_A_b9r4nJtd6_0),.din(w_dff_A_98Jc2vF24_0),.clk(gclk));
	jdff dff_A_b9r4nJtd6_0(.dout(w_dff_A_RVjpgOoh2_0),.din(w_dff_A_b9r4nJtd6_0),.clk(gclk));
	jdff dff_A_RVjpgOoh2_0(.dout(w_dff_A_8FdHHMt39_0),.din(w_dff_A_RVjpgOoh2_0),.clk(gclk));
	jdff dff_A_8FdHHMt39_0(.dout(w_dff_A_hVkwK2D39_0),.din(w_dff_A_8FdHHMt39_0),.clk(gclk));
	jdff dff_A_hVkwK2D39_0(.dout(w_dff_A_z6N7pVq27_0),.din(w_dff_A_hVkwK2D39_0),.clk(gclk));
	jdff dff_A_z6N7pVq27_0(.dout(w_dff_A_EXYENh2H3_0),.din(w_dff_A_z6N7pVq27_0),.clk(gclk));
	jdff dff_A_EXYENh2H3_0(.dout(G281),.din(w_dff_A_EXYENh2H3_0),.clk(gclk));
	jdff dff_A_Af8wiAcQ9_1(.dout(w_dff_A_aH4naish2_0),.din(w_dff_A_Af8wiAcQ9_1),.clk(gclk));
	jdff dff_A_aH4naish2_0(.dout(w_dff_A_pashgodO6_0),.din(w_dff_A_aH4naish2_0),.clk(gclk));
	jdff dff_A_pashgodO6_0(.dout(w_dff_A_El09sTYD7_0),.din(w_dff_A_pashgodO6_0),.clk(gclk));
	jdff dff_A_El09sTYD7_0(.dout(w_dff_A_K1aFsXvG3_0),.din(w_dff_A_El09sTYD7_0),.clk(gclk));
	jdff dff_A_K1aFsXvG3_0(.dout(w_dff_A_jM8U3OSz4_0),.din(w_dff_A_K1aFsXvG3_0),.clk(gclk));
	jdff dff_A_jM8U3OSz4_0(.dout(w_dff_A_DbBfKWCV8_0),.din(w_dff_A_jM8U3OSz4_0),.clk(gclk));
	jdff dff_A_DbBfKWCV8_0(.dout(w_dff_A_Z6tbIEYD7_0),.din(w_dff_A_DbBfKWCV8_0),.clk(gclk));
	jdff dff_A_Z6tbIEYD7_0(.dout(w_dff_A_duoFa2TD3_0),.din(w_dff_A_Z6tbIEYD7_0),.clk(gclk));
	jdff dff_A_duoFa2TD3_0(.dout(w_dff_A_xdPFVWud3_0),.din(w_dff_A_duoFa2TD3_0),.clk(gclk));
	jdff dff_A_xdPFVWud3_0(.dout(w_dff_A_amL6RgJj2_0),.din(w_dff_A_xdPFVWud3_0),.clk(gclk));
	jdff dff_A_amL6RgJj2_0(.dout(w_dff_A_RY2nQBeY6_0),.din(w_dff_A_amL6RgJj2_0),.clk(gclk));
	jdff dff_A_RY2nQBeY6_0(.dout(w_dff_A_y3KRjYep7_0),.din(w_dff_A_RY2nQBeY6_0),.clk(gclk));
	jdff dff_A_y3KRjYep7_0(.dout(w_dff_A_uTB6Ol2B9_0),.din(w_dff_A_y3KRjYep7_0),.clk(gclk));
	jdff dff_A_uTB6Ol2B9_0(.dout(w_dff_A_6j4n5Yqy8_0),.din(w_dff_A_uTB6Ol2B9_0),.clk(gclk));
	jdff dff_A_6j4n5Yqy8_0(.dout(w_dff_A_cSUcNv3m2_0),.din(w_dff_A_6j4n5Yqy8_0),.clk(gclk));
	jdff dff_A_cSUcNv3m2_0(.dout(w_dff_A_JLugpLH33_0),.din(w_dff_A_cSUcNv3m2_0),.clk(gclk));
	jdff dff_A_JLugpLH33_0(.dout(w_dff_A_geO3nQNh0_0),.din(w_dff_A_JLugpLH33_0),.clk(gclk));
	jdff dff_A_geO3nQNh0_0(.dout(w_dff_A_z1lCrkHb7_0),.din(w_dff_A_geO3nQNh0_0),.clk(gclk));
	jdff dff_A_z1lCrkHb7_0(.dout(w_dff_A_YT339kW83_0),.din(w_dff_A_z1lCrkHb7_0),.clk(gclk));
	jdff dff_A_YT339kW83_0(.dout(w_dff_A_eTLTVcZb4_0),.din(w_dff_A_YT339kW83_0),.clk(gclk));
	jdff dff_A_eTLTVcZb4_0(.dout(w_dff_A_tPE8SIMk4_0),.din(w_dff_A_eTLTVcZb4_0),.clk(gclk));
	jdff dff_A_tPE8SIMk4_0(.dout(w_dff_A_25mWouR81_0),.din(w_dff_A_tPE8SIMk4_0),.clk(gclk));
	jdff dff_A_25mWouR81_0(.dout(w_dff_A_QcUtAhad9_0),.din(w_dff_A_25mWouR81_0),.clk(gclk));
	jdff dff_A_QcUtAhad9_0(.dout(w_dff_A_2nMDvhkZ0_0),.din(w_dff_A_QcUtAhad9_0),.clk(gclk));
	jdff dff_A_2nMDvhkZ0_0(.dout(w_dff_A_vrhFqKrc7_0),.din(w_dff_A_2nMDvhkZ0_0),.clk(gclk));
	jdff dff_A_vrhFqKrc7_0(.dout(w_dff_A_g4RNV2No7_0),.din(w_dff_A_vrhFqKrc7_0),.clk(gclk));
	jdff dff_A_g4RNV2No7_0(.dout(G453),.din(w_dff_A_g4RNV2No7_0),.clk(gclk));
	jdff dff_A_0VY9qskf0_2(.dout(w_dff_A_lPgAGG3q1_0),.din(w_dff_A_0VY9qskf0_2),.clk(gclk));
	jdff dff_A_lPgAGG3q1_0(.dout(w_dff_A_APXpKShu5_0),.din(w_dff_A_lPgAGG3q1_0),.clk(gclk));
	jdff dff_A_APXpKShu5_0(.dout(w_dff_A_gddMmb086_0),.din(w_dff_A_APXpKShu5_0),.clk(gclk));
	jdff dff_A_gddMmb086_0(.dout(w_dff_A_S9YakP1i6_0),.din(w_dff_A_gddMmb086_0),.clk(gclk));
	jdff dff_A_S9YakP1i6_0(.dout(w_dff_A_M7m6buvZ5_0),.din(w_dff_A_S9YakP1i6_0),.clk(gclk));
	jdff dff_A_M7m6buvZ5_0(.dout(w_dff_A_LUiFWqA37_0),.din(w_dff_A_M7m6buvZ5_0),.clk(gclk));
	jdff dff_A_LUiFWqA37_0(.dout(w_dff_A_ssKtOtWQ2_0),.din(w_dff_A_LUiFWqA37_0),.clk(gclk));
	jdff dff_A_ssKtOtWQ2_0(.dout(w_dff_A_UklNp1I48_0),.din(w_dff_A_ssKtOtWQ2_0),.clk(gclk));
	jdff dff_A_UklNp1I48_0(.dout(w_dff_A_GyGplFYw1_0),.din(w_dff_A_UklNp1I48_0),.clk(gclk));
	jdff dff_A_GyGplFYw1_0(.dout(w_dff_A_5x6htadB1_0),.din(w_dff_A_GyGplFYw1_0),.clk(gclk));
	jdff dff_A_5x6htadB1_0(.dout(w_dff_A_a5CW95X31_0),.din(w_dff_A_5x6htadB1_0),.clk(gclk));
	jdff dff_A_a5CW95X31_0(.dout(w_dff_A_dxGGJhVn3_0),.din(w_dff_A_a5CW95X31_0),.clk(gclk));
	jdff dff_A_dxGGJhVn3_0(.dout(w_dff_A_t2u1sknl2_0),.din(w_dff_A_dxGGJhVn3_0),.clk(gclk));
	jdff dff_A_t2u1sknl2_0(.dout(w_dff_A_FxF6y2vM8_0),.din(w_dff_A_t2u1sknl2_0),.clk(gclk));
	jdff dff_A_FxF6y2vM8_0(.dout(w_dff_A_7sDV28nT3_0),.din(w_dff_A_FxF6y2vM8_0),.clk(gclk));
	jdff dff_A_7sDV28nT3_0(.dout(w_dff_A_rPiihOKe1_0),.din(w_dff_A_7sDV28nT3_0),.clk(gclk));
	jdff dff_A_rPiihOKe1_0(.dout(w_dff_A_2SNozCGI0_0),.din(w_dff_A_rPiihOKe1_0),.clk(gclk));
	jdff dff_A_2SNozCGI0_0(.dout(w_dff_A_4ENMKsBs6_0),.din(w_dff_A_2SNozCGI0_0),.clk(gclk));
	jdff dff_A_4ENMKsBs6_0(.dout(w_dff_A_LUT5gSwh7_0),.din(w_dff_A_4ENMKsBs6_0),.clk(gclk));
	jdff dff_A_LUT5gSwh7_0(.dout(w_dff_A_dG3qBhfD4_0),.din(w_dff_A_LUT5gSwh7_0),.clk(gclk));
	jdff dff_A_dG3qBhfD4_0(.dout(w_dff_A_fghbiNyz9_0),.din(w_dff_A_dG3qBhfD4_0),.clk(gclk));
	jdff dff_A_fghbiNyz9_0(.dout(w_dff_A_2M9YlSoT1_0),.din(w_dff_A_fghbiNyz9_0),.clk(gclk));
	jdff dff_A_2M9YlSoT1_0(.dout(w_dff_A_9Tb4U9sM0_0),.din(w_dff_A_2M9YlSoT1_0),.clk(gclk));
	jdff dff_A_9Tb4U9sM0_0(.dout(w_dff_A_7weKCX994_0),.din(w_dff_A_9Tb4U9sM0_0),.clk(gclk));
	jdff dff_A_7weKCX994_0(.dout(w_dff_A_jkmJ3FGC5_0),.din(w_dff_A_7weKCX994_0),.clk(gclk));
	jdff dff_A_jkmJ3FGC5_0(.dout(G278),.din(w_dff_A_jkmJ3FGC5_0),.clk(gclk));
	jdff dff_A_G6f97vGW1_2(.dout(w_dff_A_s8xf03aG6_0),.din(w_dff_A_G6f97vGW1_2),.clk(gclk));
	jdff dff_A_s8xf03aG6_0(.dout(w_dff_A_OCU7vohc1_0),.din(w_dff_A_s8xf03aG6_0),.clk(gclk));
	jdff dff_A_OCU7vohc1_0(.dout(w_dff_A_VrRETt0x9_0),.din(w_dff_A_OCU7vohc1_0),.clk(gclk));
	jdff dff_A_VrRETt0x9_0(.dout(w_dff_A_nwGFbIDK8_0),.din(w_dff_A_VrRETt0x9_0),.clk(gclk));
	jdff dff_A_nwGFbIDK8_0(.dout(w_dff_A_OmZndJ3G8_0),.din(w_dff_A_nwGFbIDK8_0),.clk(gclk));
	jdff dff_A_OmZndJ3G8_0(.dout(w_dff_A_e2Q9b4E56_0),.din(w_dff_A_OmZndJ3G8_0),.clk(gclk));
	jdff dff_A_e2Q9b4E56_0(.dout(w_dff_A_FlZOn2Or2_0),.din(w_dff_A_e2Q9b4E56_0),.clk(gclk));
	jdff dff_A_FlZOn2Or2_0(.dout(w_dff_A_VocoLcD50_0),.din(w_dff_A_FlZOn2Or2_0),.clk(gclk));
	jdff dff_A_VocoLcD50_0(.dout(w_dff_A_lcPBdZM54_0),.din(w_dff_A_VocoLcD50_0),.clk(gclk));
	jdff dff_A_lcPBdZM54_0(.dout(w_dff_A_hn78JPsk4_0),.din(w_dff_A_lcPBdZM54_0),.clk(gclk));
	jdff dff_A_hn78JPsk4_0(.dout(w_dff_A_geTMApaP0_0),.din(w_dff_A_hn78JPsk4_0),.clk(gclk));
	jdff dff_A_geTMApaP0_0(.dout(w_dff_A_A221yhql8_0),.din(w_dff_A_geTMApaP0_0),.clk(gclk));
	jdff dff_A_A221yhql8_0(.dout(w_dff_A_3TOpHBz23_0),.din(w_dff_A_A221yhql8_0),.clk(gclk));
	jdff dff_A_3TOpHBz23_0(.dout(w_dff_A_dqX3mFAf6_0),.din(w_dff_A_3TOpHBz23_0),.clk(gclk));
	jdff dff_A_dqX3mFAf6_0(.dout(w_dff_A_GuAxUeW23_0),.din(w_dff_A_dqX3mFAf6_0),.clk(gclk));
	jdff dff_A_GuAxUeW23_0(.dout(w_dff_A_ppNgMf3V4_0),.din(w_dff_A_GuAxUeW23_0),.clk(gclk));
	jdff dff_A_ppNgMf3V4_0(.dout(w_dff_A_bXcR52dd6_0),.din(w_dff_A_ppNgMf3V4_0),.clk(gclk));
	jdff dff_A_bXcR52dd6_0(.dout(w_dff_A_hiw6Tp391_0),.din(w_dff_A_bXcR52dd6_0),.clk(gclk));
	jdff dff_A_hiw6Tp391_0(.dout(w_dff_A_BqBGIG8B9_0),.din(w_dff_A_hiw6Tp391_0),.clk(gclk));
	jdff dff_A_BqBGIG8B9_0(.dout(w_dff_A_EDqhMU9M5_0),.din(w_dff_A_BqBGIG8B9_0),.clk(gclk));
	jdff dff_A_EDqhMU9M5_0(.dout(G373),.din(w_dff_A_EDqhMU9M5_0),.clk(gclk));
	jdff dff_A_tmAqux6d0_2(.dout(G246),.din(w_dff_A_tmAqux6d0_2),.clk(gclk));
	jdff dff_A_7bncmJrH1_2(.dout(w_dff_A_oxo8IFOF4_0),.din(w_dff_A_7bncmJrH1_2),.clk(gclk));
	jdff dff_A_oxo8IFOF4_0(.dout(w_dff_A_NnB8316l5_0),.din(w_dff_A_oxo8IFOF4_0),.clk(gclk));
	jdff dff_A_NnB8316l5_0(.dout(w_dff_A_XCkeH2EA7_0),.din(w_dff_A_NnB8316l5_0),.clk(gclk));
	jdff dff_A_XCkeH2EA7_0(.dout(w_dff_A_Onh8qkL43_0),.din(w_dff_A_XCkeH2EA7_0),.clk(gclk));
	jdff dff_A_Onh8qkL43_0(.dout(w_dff_A_tiBrdGfd2_0),.din(w_dff_A_Onh8qkL43_0),.clk(gclk));
	jdff dff_A_tiBrdGfd2_0(.dout(w_dff_A_yqGXmjzH1_0),.din(w_dff_A_tiBrdGfd2_0),.clk(gclk));
	jdff dff_A_yqGXmjzH1_0(.dout(G258),.din(w_dff_A_yqGXmjzH1_0),.clk(gclk));
	jdff dff_A_slq4IEGl3_2(.dout(w_dff_A_49d9nwLz0_0),.din(w_dff_A_slq4IEGl3_2),.clk(gclk));
	jdff dff_A_49d9nwLz0_0(.dout(w_dff_A_aAWMaHUU6_0),.din(w_dff_A_49d9nwLz0_0),.clk(gclk));
	jdff dff_A_aAWMaHUU6_0(.dout(w_dff_A_TLjT1jhb1_0),.din(w_dff_A_aAWMaHUU6_0),.clk(gclk));
	jdff dff_A_TLjT1jhb1_0(.dout(w_dff_A_2fpl2d8b8_0),.din(w_dff_A_TLjT1jhb1_0),.clk(gclk));
	jdff dff_A_2fpl2d8b8_0(.dout(w_dff_A_2mIXvj9h8_0),.din(w_dff_A_2fpl2d8b8_0),.clk(gclk));
	jdff dff_A_2mIXvj9h8_0(.dout(w_dff_A_P0LTGYCI5_0),.din(w_dff_A_2mIXvj9h8_0),.clk(gclk));
	jdff dff_A_P0LTGYCI5_0(.dout(G264),.din(w_dff_A_P0LTGYCI5_0),.clk(gclk));
	jdff dff_A_xynYSXoD0_2(.dout(G270),.din(w_dff_A_xynYSXoD0_2),.clk(gclk));
	jdff dff_A_7SRXhOvO3_2(.dout(w_dff_A_qCKrcPKM0_0),.din(w_dff_A_7SRXhOvO3_2),.clk(gclk));
	jdff dff_A_qCKrcPKM0_0(.dout(w_dff_A_oLHtzAyD0_0),.din(w_dff_A_qCKrcPKM0_0),.clk(gclk));
	jdff dff_A_oLHtzAyD0_0(.dout(w_dff_A_y9fU334t0_0),.din(w_dff_A_oLHtzAyD0_0),.clk(gclk));
	jdff dff_A_y9fU334t0_0(.dout(w_dff_A_iOBIuayx8_0),.din(w_dff_A_y9fU334t0_0),.clk(gclk));
	jdff dff_A_iOBIuayx8_0(.dout(w_dff_A_g1FIEsQG9_0),.din(w_dff_A_iOBIuayx8_0),.clk(gclk));
	jdff dff_A_g1FIEsQG9_0(.dout(w_dff_A_QOPMQEOA4_0),.din(w_dff_A_g1FIEsQG9_0),.clk(gclk));
	jdff dff_A_QOPMQEOA4_0(.dout(w_dff_A_k6TNAtKY3_0),.din(w_dff_A_QOPMQEOA4_0),.clk(gclk));
	jdff dff_A_k6TNAtKY3_0(.dout(w_dff_A_QbskiEbA7_0),.din(w_dff_A_k6TNAtKY3_0),.clk(gclk));
	jdff dff_A_QbskiEbA7_0(.dout(w_dff_A_nHxBmp7f6_0),.din(w_dff_A_QbskiEbA7_0),.clk(gclk));
	jdff dff_A_nHxBmp7f6_0(.dout(w_dff_A_kYpTbEXj1_0),.din(w_dff_A_nHxBmp7f6_0),.clk(gclk));
	jdff dff_A_kYpTbEXj1_0(.dout(w_dff_A_djZcg1LF8_0),.din(w_dff_A_kYpTbEXj1_0),.clk(gclk));
	jdff dff_A_djZcg1LF8_0(.dout(w_dff_A_YFqxQxk80_0),.din(w_dff_A_djZcg1LF8_0),.clk(gclk));
	jdff dff_A_YFqxQxk80_0(.dout(w_dff_A_9djJd31R7_0),.din(w_dff_A_YFqxQxk80_0),.clk(gclk));
	jdff dff_A_9djJd31R7_0(.dout(w_dff_A_iLon1dHl7_0),.din(w_dff_A_9djJd31R7_0),.clk(gclk));
	jdff dff_A_iLon1dHl7_0(.dout(G388),.din(w_dff_A_iLon1dHl7_0),.clk(gclk));
	jdff dff_A_ZxG7VkOx2_2(.dout(w_dff_A_buwlAT6j5_0),.din(w_dff_A_ZxG7VkOx2_2),.clk(gclk));
	jdff dff_A_buwlAT6j5_0(.dout(w_dff_A_iir7dVLr7_0),.din(w_dff_A_buwlAT6j5_0),.clk(gclk));
	jdff dff_A_iir7dVLr7_0(.dout(w_dff_A_t99NrWx89_0),.din(w_dff_A_iir7dVLr7_0),.clk(gclk));
	jdff dff_A_t99NrWx89_0(.dout(w_dff_A_k2xuEJhq2_0),.din(w_dff_A_t99NrWx89_0),.clk(gclk));
	jdff dff_A_k2xuEJhq2_0(.dout(w_dff_A_5lcdd36d9_0),.din(w_dff_A_k2xuEJhq2_0),.clk(gclk));
	jdff dff_A_5lcdd36d9_0(.dout(w_dff_A_Jga4aHfz7_0),.din(w_dff_A_5lcdd36d9_0),.clk(gclk));
	jdff dff_A_Jga4aHfz7_0(.dout(w_dff_A_RvlmARqO2_0),.din(w_dff_A_Jga4aHfz7_0),.clk(gclk));
	jdff dff_A_RvlmARqO2_0(.dout(w_dff_A_Ro8C5pz43_0),.din(w_dff_A_RvlmARqO2_0),.clk(gclk));
	jdff dff_A_Ro8C5pz43_0(.dout(w_dff_A_nz3BPLfr4_0),.din(w_dff_A_Ro8C5pz43_0),.clk(gclk));
	jdff dff_A_nz3BPLfr4_0(.dout(w_dff_A_TxUb3m2O8_0),.din(w_dff_A_nz3BPLfr4_0),.clk(gclk));
	jdff dff_A_TxUb3m2O8_0(.dout(w_dff_A_66DJyi1t6_0),.din(w_dff_A_TxUb3m2O8_0),.clk(gclk));
	jdff dff_A_66DJyi1t6_0(.dout(w_dff_A_SYr65DJ72_0),.din(w_dff_A_66DJyi1t6_0),.clk(gclk));
	jdff dff_A_SYr65DJ72_0(.dout(w_dff_A_yVq3gOil5_0),.din(w_dff_A_SYr65DJ72_0),.clk(gclk));
	jdff dff_A_yVq3gOil5_0(.dout(w_dff_A_4yEgPXer3_0),.din(w_dff_A_yVq3gOil5_0),.clk(gclk));
	jdff dff_A_4yEgPXer3_0(.dout(w_dff_A_2OTiDwfv0_0),.din(w_dff_A_4yEgPXer3_0),.clk(gclk));
	jdff dff_A_2OTiDwfv0_0(.dout(w_dff_A_PUlOZRWD3_0),.din(w_dff_A_2OTiDwfv0_0),.clk(gclk));
	jdff dff_A_PUlOZRWD3_0(.dout(G391),.din(w_dff_A_PUlOZRWD3_0),.clk(gclk));
	jdff dff_A_vdMi5oyR9_2(.dout(w_dff_A_7VqXO72Z3_0),.din(w_dff_A_vdMi5oyR9_2),.clk(gclk));
	jdff dff_A_7VqXO72Z3_0(.dout(w_dff_A_kHutkUE59_0),.din(w_dff_A_7VqXO72Z3_0),.clk(gclk));
	jdff dff_A_kHutkUE59_0(.dout(w_dff_A_pMDITxTf6_0),.din(w_dff_A_kHutkUE59_0),.clk(gclk));
	jdff dff_A_pMDITxTf6_0(.dout(w_dff_A_r99BU6pK1_0),.din(w_dff_A_pMDITxTf6_0),.clk(gclk));
	jdff dff_A_r99BU6pK1_0(.dout(w_dff_A_tJLzHwmR6_0),.din(w_dff_A_r99BU6pK1_0),.clk(gclk));
	jdff dff_A_tJLzHwmR6_0(.dout(w_dff_A_cdUZt36Y9_0),.din(w_dff_A_tJLzHwmR6_0),.clk(gclk));
	jdff dff_A_cdUZt36Y9_0(.dout(w_dff_A_7DQpceER2_0),.din(w_dff_A_cdUZt36Y9_0),.clk(gclk));
	jdff dff_A_7DQpceER2_0(.dout(w_dff_A_kJdg2TJO2_0),.din(w_dff_A_7DQpceER2_0),.clk(gclk));
	jdff dff_A_kJdg2TJO2_0(.dout(w_dff_A_HDjEF4hZ9_0),.din(w_dff_A_kJdg2TJO2_0),.clk(gclk));
	jdff dff_A_HDjEF4hZ9_0(.dout(w_dff_A_N3DH1ayv2_0),.din(w_dff_A_HDjEF4hZ9_0),.clk(gclk));
	jdff dff_A_N3DH1ayv2_0(.dout(w_dff_A_ZUqMxNS22_0),.din(w_dff_A_N3DH1ayv2_0),.clk(gclk));
	jdff dff_A_ZUqMxNS22_0(.dout(w_dff_A_hlbWUXh28_0),.din(w_dff_A_ZUqMxNS22_0),.clk(gclk));
	jdff dff_A_hlbWUXh28_0(.dout(w_dff_A_pAvAUTJu4_0),.din(w_dff_A_hlbWUXh28_0),.clk(gclk));
	jdff dff_A_pAvAUTJu4_0(.dout(w_dff_A_AYz5eDMm6_0),.din(w_dff_A_pAvAUTJu4_0),.clk(gclk));
	jdff dff_A_AYz5eDMm6_0(.dout(w_dff_A_VwaSmJ2w7_0),.din(w_dff_A_AYz5eDMm6_0),.clk(gclk));
	jdff dff_A_VwaSmJ2w7_0(.dout(w_dff_A_ZKkaejFi5_0),.din(w_dff_A_VwaSmJ2w7_0),.clk(gclk));
	jdff dff_A_ZKkaejFi5_0(.dout(w_dff_A_kLbTUx1v9_0),.din(w_dff_A_ZKkaejFi5_0),.clk(gclk));
	jdff dff_A_kLbTUx1v9_0(.dout(G394),.din(w_dff_A_kLbTUx1v9_0),.clk(gclk));
	jdff dff_A_UGZaqdrl9_2(.dout(w_dff_A_Yc9VjNUH1_0),.din(w_dff_A_UGZaqdrl9_2),.clk(gclk));
	jdff dff_A_Yc9VjNUH1_0(.dout(w_dff_A_yiTi0O691_0),.din(w_dff_A_Yc9VjNUH1_0),.clk(gclk));
	jdff dff_A_yiTi0O691_0(.dout(w_dff_A_3jugHNN26_0),.din(w_dff_A_yiTi0O691_0),.clk(gclk));
	jdff dff_A_3jugHNN26_0(.dout(w_dff_A_DLBAkYuf0_0),.din(w_dff_A_3jugHNN26_0),.clk(gclk));
	jdff dff_A_DLBAkYuf0_0(.dout(w_dff_A_fetJtNLW0_0),.din(w_dff_A_DLBAkYuf0_0),.clk(gclk));
	jdff dff_A_fetJtNLW0_0(.dout(w_dff_A_QrLrEXi49_0),.din(w_dff_A_fetJtNLW0_0),.clk(gclk));
	jdff dff_A_QrLrEXi49_0(.dout(w_dff_A_lcYw7r1L9_0),.din(w_dff_A_QrLrEXi49_0),.clk(gclk));
	jdff dff_A_lcYw7r1L9_0(.dout(w_dff_A_7iTlmmo35_0),.din(w_dff_A_lcYw7r1L9_0),.clk(gclk));
	jdff dff_A_7iTlmmo35_0(.dout(w_dff_A_odoTsM1w6_0),.din(w_dff_A_7iTlmmo35_0),.clk(gclk));
	jdff dff_A_odoTsM1w6_0(.dout(w_dff_A_OjaMMZRV2_0),.din(w_dff_A_odoTsM1w6_0),.clk(gclk));
	jdff dff_A_OjaMMZRV2_0(.dout(w_dff_A_03qjPbrJ8_0),.din(w_dff_A_OjaMMZRV2_0),.clk(gclk));
	jdff dff_A_03qjPbrJ8_0(.dout(w_dff_A_nN49KSXe7_0),.din(w_dff_A_03qjPbrJ8_0),.clk(gclk));
	jdff dff_A_nN49KSXe7_0(.dout(w_dff_A_XCzMfxRA7_0),.din(w_dff_A_nN49KSXe7_0),.clk(gclk));
	jdff dff_A_XCzMfxRA7_0(.dout(w_dff_A_0pppbt6K3_0),.din(w_dff_A_XCzMfxRA7_0),.clk(gclk));
	jdff dff_A_0pppbt6K3_0(.dout(w_dff_A_YQEDeZsF8_0),.din(w_dff_A_0pppbt6K3_0),.clk(gclk));
	jdff dff_A_YQEDeZsF8_0(.dout(w_dff_A_zZCSepld7_0),.din(w_dff_A_YQEDeZsF8_0),.clk(gclk));
	jdff dff_A_zZCSepld7_0(.dout(w_dff_A_H5ZKYjVU1_0),.din(w_dff_A_zZCSepld7_0),.clk(gclk));
	jdff dff_A_H5ZKYjVU1_0(.dout(w_dff_A_cItHHJ9M8_0),.din(w_dff_A_H5ZKYjVU1_0),.clk(gclk));
	jdff dff_A_cItHHJ9M8_0(.dout(G397),.din(w_dff_A_cItHHJ9M8_0),.clk(gclk));
	jdff dff_A_Z1rwaf0c9_2(.dout(w_dff_A_lpEtMeBB0_0),.din(w_dff_A_Z1rwaf0c9_2),.clk(gclk));
	jdff dff_A_lpEtMeBB0_0(.dout(w_dff_A_B7bR7plx4_0),.din(w_dff_A_lpEtMeBB0_0),.clk(gclk));
	jdff dff_A_B7bR7plx4_0(.dout(w_dff_A_YPyXDQlB4_0),.din(w_dff_A_B7bR7plx4_0),.clk(gclk));
	jdff dff_A_YPyXDQlB4_0(.dout(w_dff_A_GzCislSo9_0),.din(w_dff_A_YPyXDQlB4_0),.clk(gclk));
	jdff dff_A_GzCislSo9_0(.dout(w_dff_A_Pb6qYUgU2_0),.din(w_dff_A_GzCislSo9_0),.clk(gclk));
	jdff dff_A_Pb6qYUgU2_0(.dout(w_dff_A_a0TWqPZN0_0),.din(w_dff_A_Pb6qYUgU2_0),.clk(gclk));
	jdff dff_A_a0TWqPZN0_0(.dout(w_dff_A_8xeGaHK31_0),.din(w_dff_A_a0TWqPZN0_0),.clk(gclk));
	jdff dff_A_8xeGaHK31_0(.dout(w_dff_A_Nt7mpm9u6_0),.din(w_dff_A_8xeGaHK31_0),.clk(gclk));
	jdff dff_A_Nt7mpm9u6_0(.dout(w_dff_A_YSmqPlh66_0),.din(w_dff_A_Nt7mpm9u6_0),.clk(gclk));
	jdff dff_A_YSmqPlh66_0(.dout(w_dff_A_8ieq2PLb4_0),.din(w_dff_A_YSmqPlh66_0),.clk(gclk));
	jdff dff_A_8ieq2PLb4_0(.dout(w_dff_A_sIFMCCTq3_0),.din(w_dff_A_8ieq2PLb4_0),.clk(gclk));
	jdff dff_A_sIFMCCTq3_0(.dout(w_dff_A_y2NcQUqF0_0),.din(w_dff_A_sIFMCCTq3_0),.clk(gclk));
	jdff dff_A_y2NcQUqF0_0(.dout(G376),.din(w_dff_A_y2NcQUqF0_0),.clk(gclk));
	jdff dff_A_6eSmLkqc9_2(.dout(w_dff_A_T7rTPfZH9_0),.din(w_dff_A_6eSmLkqc9_2),.clk(gclk));
	jdff dff_A_T7rTPfZH9_0(.dout(w_dff_A_oEjHxI8S8_0),.din(w_dff_A_T7rTPfZH9_0),.clk(gclk));
	jdff dff_A_oEjHxI8S8_0(.dout(w_dff_A_6qtVXU9u7_0),.din(w_dff_A_oEjHxI8S8_0),.clk(gclk));
	jdff dff_A_6qtVXU9u7_0(.dout(w_dff_A_Dx5l8OnE5_0),.din(w_dff_A_6qtVXU9u7_0),.clk(gclk));
	jdff dff_A_Dx5l8OnE5_0(.dout(w_dff_A_lFBGzwUw0_0),.din(w_dff_A_Dx5l8OnE5_0),.clk(gclk));
	jdff dff_A_lFBGzwUw0_0(.dout(w_dff_A_wGNiJXX33_0),.din(w_dff_A_lFBGzwUw0_0),.clk(gclk));
	jdff dff_A_wGNiJXX33_0(.dout(w_dff_A_8NSuVLOE6_0),.din(w_dff_A_wGNiJXX33_0),.clk(gclk));
	jdff dff_A_8NSuVLOE6_0(.dout(w_dff_A_0fddDv9l5_0),.din(w_dff_A_8NSuVLOE6_0),.clk(gclk));
	jdff dff_A_0fddDv9l5_0(.dout(w_dff_A_VWNEkdXj9_0),.din(w_dff_A_0fddDv9l5_0),.clk(gclk));
	jdff dff_A_VWNEkdXj9_0(.dout(w_dff_A_GwCZjVlW8_0),.din(w_dff_A_VWNEkdXj9_0),.clk(gclk));
	jdff dff_A_GwCZjVlW8_0(.dout(w_dff_A_NKRZ3IAE1_0),.din(w_dff_A_GwCZjVlW8_0),.clk(gclk));
	jdff dff_A_NKRZ3IAE1_0(.dout(w_dff_A_IllGmloY9_0),.din(w_dff_A_NKRZ3IAE1_0),.clk(gclk));
	jdff dff_A_IllGmloY9_0(.dout(w_dff_A_m9AUuwwd7_0),.din(w_dff_A_IllGmloY9_0),.clk(gclk));
	jdff dff_A_m9AUuwwd7_0(.dout(G379),.din(w_dff_A_m9AUuwwd7_0),.clk(gclk));
	jdff dff_A_zlCQ34f47_2(.dout(w_dff_A_TKl59R6U4_0),.din(w_dff_A_zlCQ34f47_2),.clk(gclk));
	jdff dff_A_TKl59R6U4_0(.dout(w_dff_A_WFvjHIVR2_0),.din(w_dff_A_TKl59R6U4_0),.clk(gclk));
	jdff dff_A_WFvjHIVR2_0(.dout(w_dff_A_9Br4c2dp0_0),.din(w_dff_A_WFvjHIVR2_0),.clk(gclk));
	jdff dff_A_9Br4c2dp0_0(.dout(w_dff_A_vWMPW1Se8_0),.din(w_dff_A_9Br4c2dp0_0),.clk(gclk));
	jdff dff_A_vWMPW1Se8_0(.dout(w_dff_A_ZFraZAjN7_0),.din(w_dff_A_vWMPW1Se8_0),.clk(gclk));
	jdff dff_A_ZFraZAjN7_0(.dout(w_dff_A_7AKyzm9g0_0),.din(w_dff_A_ZFraZAjN7_0),.clk(gclk));
	jdff dff_A_7AKyzm9g0_0(.dout(w_dff_A_SS5VBVme5_0),.din(w_dff_A_7AKyzm9g0_0),.clk(gclk));
	jdff dff_A_SS5VBVme5_0(.dout(w_dff_A_4mf447Bi3_0),.din(w_dff_A_SS5VBVme5_0),.clk(gclk));
	jdff dff_A_4mf447Bi3_0(.dout(w_dff_A_ccXVZmas3_0),.din(w_dff_A_4mf447Bi3_0),.clk(gclk));
	jdff dff_A_ccXVZmas3_0(.dout(w_dff_A_eqDGjRQR7_0),.din(w_dff_A_ccXVZmas3_0),.clk(gclk));
	jdff dff_A_eqDGjRQR7_0(.dout(w_dff_A_6KGopj4c3_0),.din(w_dff_A_eqDGjRQR7_0),.clk(gclk));
	jdff dff_A_6KGopj4c3_0(.dout(w_dff_A_j3fEP8LP3_0),.din(w_dff_A_6KGopj4c3_0),.clk(gclk));
	jdff dff_A_j3fEP8LP3_0(.dout(w_dff_A_pLJlfSJl1_0),.din(w_dff_A_j3fEP8LP3_0),.clk(gclk));
	jdff dff_A_pLJlfSJl1_0(.dout(G382),.din(w_dff_A_pLJlfSJl1_0),.clk(gclk));
	jdff dff_A_zwekv3fv4_2(.dout(w_dff_A_F8BJTSfE3_0),.din(w_dff_A_zwekv3fv4_2),.clk(gclk));
	jdff dff_A_F8BJTSfE3_0(.dout(w_dff_A_U28oKJzG7_0),.din(w_dff_A_F8BJTSfE3_0),.clk(gclk));
	jdff dff_A_U28oKJzG7_0(.dout(w_dff_A_Uk4V7U748_0),.din(w_dff_A_U28oKJzG7_0),.clk(gclk));
	jdff dff_A_Uk4V7U748_0(.dout(w_dff_A_ttxLDRdL0_0),.din(w_dff_A_Uk4V7U748_0),.clk(gclk));
	jdff dff_A_ttxLDRdL0_0(.dout(w_dff_A_BUxHzEkm9_0),.din(w_dff_A_ttxLDRdL0_0),.clk(gclk));
	jdff dff_A_BUxHzEkm9_0(.dout(w_dff_A_P6c34Js75_0),.din(w_dff_A_BUxHzEkm9_0),.clk(gclk));
	jdff dff_A_P6c34Js75_0(.dout(w_dff_A_CfU4rOil8_0),.din(w_dff_A_P6c34Js75_0),.clk(gclk));
	jdff dff_A_CfU4rOil8_0(.dout(w_dff_A_CzMeV7QN3_0),.din(w_dff_A_CfU4rOil8_0),.clk(gclk));
	jdff dff_A_CzMeV7QN3_0(.dout(w_dff_A_p7Ss9eQc5_0),.din(w_dff_A_CzMeV7QN3_0),.clk(gclk));
	jdff dff_A_p7Ss9eQc5_0(.dout(w_dff_A_F7DMAR7U6_0),.din(w_dff_A_p7Ss9eQc5_0),.clk(gclk));
	jdff dff_A_F7DMAR7U6_0(.dout(w_dff_A_WNK5iPcp6_0),.din(w_dff_A_F7DMAR7U6_0),.clk(gclk));
	jdff dff_A_WNK5iPcp6_0(.dout(w_dff_A_N9fNAT5n7_0),.din(w_dff_A_WNK5iPcp6_0),.clk(gclk));
	jdff dff_A_N9fNAT5n7_0(.dout(w_dff_A_zxlsppAi9_0),.din(w_dff_A_N9fNAT5n7_0),.clk(gclk));
	jdff dff_A_zxlsppAi9_0(.dout(w_dff_A_9DBGI9NS8_0),.din(w_dff_A_zxlsppAi9_0),.clk(gclk));
	jdff dff_A_9DBGI9NS8_0(.dout(w_dff_A_QSz4wJVn0_0),.din(w_dff_A_9DBGI9NS8_0),.clk(gclk));
	jdff dff_A_QSz4wJVn0_0(.dout(G385),.din(w_dff_A_QSz4wJVn0_0),.clk(gclk));
	jdff dff_A_lCOwNbj03_1(.dout(w_dff_A_OIFj3G9A1_0),.din(w_dff_A_lCOwNbj03_1),.clk(gclk));
	jdff dff_A_OIFj3G9A1_0(.dout(w_dff_A_84NcbFgo0_0),.din(w_dff_A_OIFj3G9A1_0),.clk(gclk));
	jdff dff_A_84NcbFgo0_0(.dout(w_dff_A_JcCbx2fa8_0),.din(w_dff_A_84NcbFgo0_0),.clk(gclk));
	jdff dff_A_JcCbx2fa8_0(.dout(w_dff_A_IM5fMFUJ7_0),.din(w_dff_A_JcCbx2fa8_0),.clk(gclk));
	jdff dff_A_IM5fMFUJ7_0(.dout(w_dff_A_ZwGittOs1_0),.din(w_dff_A_IM5fMFUJ7_0),.clk(gclk));
	jdff dff_A_ZwGittOs1_0(.dout(w_dff_A_lZJniq0H2_0),.din(w_dff_A_ZwGittOs1_0),.clk(gclk));
	jdff dff_A_lZJniq0H2_0(.dout(w_dff_A_KbWepYJm3_0),.din(w_dff_A_lZJniq0H2_0),.clk(gclk));
	jdff dff_A_KbWepYJm3_0(.dout(w_dff_A_VkzE3nOL7_0),.din(w_dff_A_KbWepYJm3_0),.clk(gclk));
	jdff dff_A_VkzE3nOL7_0(.dout(w_dff_A_8hSFBnCz5_0),.din(w_dff_A_VkzE3nOL7_0),.clk(gclk));
	jdff dff_A_8hSFBnCz5_0(.dout(w_dff_A_OmpXChON8_0),.din(w_dff_A_8hSFBnCz5_0),.clk(gclk));
	jdff dff_A_OmpXChON8_0(.dout(w_dff_A_dxJhnket5_0),.din(w_dff_A_OmpXChON8_0),.clk(gclk));
	jdff dff_A_dxJhnket5_0(.dout(w_dff_A_58HqTgeW2_0),.din(w_dff_A_dxJhnket5_0),.clk(gclk));
	jdff dff_A_58HqTgeW2_0(.dout(w_dff_A_C2XFWLrw2_0),.din(w_dff_A_58HqTgeW2_0),.clk(gclk));
	jdff dff_A_C2XFWLrw2_0(.dout(w_dff_A_IgVUFivB9_0),.din(w_dff_A_C2XFWLrw2_0),.clk(gclk));
	jdff dff_A_IgVUFivB9_0(.dout(w_dff_A_r7VgIBJl5_0),.din(w_dff_A_IgVUFivB9_0),.clk(gclk));
	jdff dff_A_r7VgIBJl5_0(.dout(G412),.din(w_dff_A_r7VgIBJl5_0),.clk(gclk));
	jdff dff_A_sj0YHAtv4_1(.dout(w_dff_A_fswTJykB5_0),.din(w_dff_A_sj0YHAtv4_1),.clk(gclk));
	jdff dff_A_fswTJykB5_0(.dout(w_dff_A_WgDcwJZP4_0),.din(w_dff_A_fswTJykB5_0),.clk(gclk));
	jdff dff_A_WgDcwJZP4_0(.dout(w_dff_A_4zcGyYSq2_0),.din(w_dff_A_WgDcwJZP4_0),.clk(gclk));
	jdff dff_A_4zcGyYSq2_0(.dout(w_dff_A_z3xdx7EG1_0),.din(w_dff_A_4zcGyYSq2_0),.clk(gclk));
	jdff dff_A_z3xdx7EG1_0(.dout(w_dff_A_aIMctxaR4_0),.din(w_dff_A_z3xdx7EG1_0),.clk(gclk));
	jdff dff_A_aIMctxaR4_0(.dout(w_dff_A_XzhAvNwz3_0),.din(w_dff_A_aIMctxaR4_0),.clk(gclk));
	jdff dff_A_XzhAvNwz3_0(.dout(w_dff_A_lgCtd7vg1_0),.din(w_dff_A_XzhAvNwz3_0),.clk(gclk));
	jdff dff_A_lgCtd7vg1_0(.dout(w_dff_A_wUbGZ0TX8_0),.din(w_dff_A_lgCtd7vg1_0),.clk(gclk));
	jdff dff_A_wUbGZ0TX8_0(.dout(w_dff_A_Ff1ch4qe1_0),.din(w_dff_A_wUbGZ0TX8_0),.clk(gclk));
	jdff dff_A_Ff1ch4qe1_0(.dout(w_dff_A_diDwxWGV7_0),.din(w_dff_A_Ff1ch4qe1_0),.clk(gclk));
	jdff dff_A_diDwxWGV7_0(.dout(w_dff_A_98STIIH93_0),.din(w_dff_A_diDwxWGV7_0),.clk(gclk));
	jdff dff_A_98STIIH93_0(.dout(w_dff_A_DNtzr0o88_0),.din(w_dff_A_98STIIH93_0),.clk(gclk));
	jdff dff_A_DNtzr0o88_0(.dout(w_dff_A_VdMoBVek6_0),.din(w_dff_A_DNtzr0o88_0),.clk(gclk));
	jdff dff_A_VdMoBVek6_0(.dout(w_dff_A_0bAyuyYD7_0),.din(w_dff_A_VdMoBVek6_0),.clk(gclk));
	jdff dff_A_0bAyuyYD7_0(.dout(w_dff_A_oYXvcS0d5_0),.din(w_dff_A_0bAyuyYD7_0),.clk(gclk));
	jdff dff_A_oYXvcS0d5_0(.dout(G414),.din(w_dff_A_oYXvcS0d5_0),.clk(gclk));
	jdff dff_A_pXJgTd7U2_1(.dout(w_dff_A_0fBnK0dk5_0),.din(w_dff_A_pXJgTd7U2_1),.clk(gclk));
	jdff dff_A_0fBnK0dk5_0(.dout(w_dff_A_9H6c9TZi2_0),.din(w_dff_A_0fBnK0dk5_0),.clk(gclk));
	jdff dff_A_9H6c9TZi2_0(.dout(w_dff_A_7qN883YS7_0),.din(w_dff_A_9H6c9TZi2_0),.clk(gclk));
	jdff dff_A_7qN883YS7_0(.dout(w_dff_A_xaVg0qhm5_0),.din(w_dff_A_7qN883YS7_0),.clk(gclk));
	jdff dff_A_xaVg0qhm5_0(.dout(w_dff_A_UJPSPG4S1_0),.din(w_dff_A_xaVg0qhm5_0),.clk(gclk));
	jdff dff_A_UJPSPG4S1_0(.dout(w_dff_A_qQNR8Vp26_0),.din(w_dff_A_UJPSPG4S1_0),.clk(gclk));
	jdff dff_A_qQNR8Vp26_0(.dout(w_dff_A_CuYlR7iv7_0),.din(w_dff_A_qQNR8Vp26_0),.clk(gclk));
	jdff dff_A_CuYlR7iv7_0(.dout(w_dff_A_ru4lMoYc5_0),.din(w_dff_A_CuYlR7iv7_0),.clk(gclk));
	jdff dff_A_ru4lMoYc5_0(.dout(w_dff_A_IwAN1f470_0),.din(w_dff_A_ru4lMoYc5_0),.clk(gclk));
	jdff dff_A_IwAN1f470_0(.dout(w_dff_A_qVHozKTM8_0),.din(w_dff_A_IwAN1f470_0),.clk(gclk));
	jdff dff_A_qVHozKTM8_0(.dout(w_dff_A_wdN7iPWG9_0),.din(w_dff_A_qVHozKTM8_0),.clk(gclk));
	jdff dff_A_wdN7iPWG9_0(.dout(w_dff_A_5GH4LxQw0_0),.din(w_dff_A_wdN7iPWG9_0),.clk(gclk));
	jdff dff_A_5GH4LxQw0_0(.dout(w_dff_A_zXAkUw0c5_0),.din(w_dff_A_5GH4LxQw0_0),.clk(gclk));
	jdff dff_A_zXAkUw0c5_0(.dout(G416),.din(w_dff_A_zXAkUw0c5_0),.clk(gclk));
	jdff dff_A_uIYyqE1Q1_2(.dout(w_dff_A_7lkjoFMC0_0),.din(w_dff_A_uIYyqE1Q1_2),.clk(gclk));
	jdff dff_A_7lkjoFMC0_0(.dout(w_dff_A_hG3WFMBp7_0),.din(w_dff_A_7lkjoFMC0_0),.clk(gclk));
	jdff dff_A_hG3WFMBp7_0(.dout(w_dff_A_iFfG8cWD7_0),.din(w_dff_A_hG3WFMBp7_0),.clk(gclk));
	jdff dff_A_iFfG8cWD7_0(.dout(w_dff_A_PJaBNnYC8_0),.din(w_dff_A_iFfG8cWD7_0),.clk(gclk));
	jdff dff_A_PJaBNnYC8_0(.dout(w_dff_A_T2yxENLR8_0),.din(w_dff_A_PJaBNnYC8_0),.clk(gclk));
	jdff dff_A_T2yxENLR8_0(.dout(w_dff_A_BFPRcEdi6_0),.din(w_dff_A_T2yxENLR8_0),.clk(gclk));
	jdff dff_A_BFPRcEdi6_0(.dout(G249),.din(w_dff_A_BFPRcEdi6_0),.clk(gclk));
	jdff dff_A_7i4JzMTm0_2(.dout(w_dff_A_ICTlbeD93_0),.din(w_dff_A_7i4JzMTm0_2),.clk(gclk));
	jdff dff_A_ICTlbeD93_0(.dout(w_dff_A_wNQsUtmF8_0),.din(w_dff_A_ICTlbeD93_0),.clk(gclk));
	jdff dff_A_wNQsUtmF8_0(.dout(w_dff_A_A0q2JVHP4_0),.din(w_dff_A_wNQsUtmF8_0),.clk(gclk));
	jdff dff_A_A0q2JVHP4_0(.dout(w_dff_A_iKwEJnzs3_0),.din(w_dff_A_A0q2JVHP4_0),.clk(gclk));
	jdff dff_A_iKwEJnzs3_0(.dout(w_dff_A_tmynV1jm6_0),.din(w_dff_A_iKwEJnzs3_0),.clk(gclk));
	jdff dff_A_tmynV1jm6_0(.dout(w_dff_A_BChzxR5r2_0),.din(w_dff_A_tmynV1jm6_0),.clk(gclk));
	jdff dff_A_BChzxR5r2_0(.dout(w_dff_A_vFD3QYLO8_0),.din(w_dff_A_BChzxR5r2_0),.clk(gclk));
	jdff dff_A_vFD3QYLO8_0(.dout(w_dff_A_l7Tx6VIj5_0),.din(w_dff_A_vFD3QYLO8_0),.clk(gclk));
	jdff dff_A_l7Tx6VIj5_0(.dout(w_dff_A_A4vaxYBV0_0),.din(w_dff_A_l7Tx6VIj5_0),.clk(gclk));
	jdff dff_A_A4vaxYBV0_0(.dout(G295),.din(w_dff_A_A4vaxYBV0_0),.clk(gclk));
	jdff dff_A_DICIafTn4_2(.dout(w_dff_A_xKwUIsha4_0),.din(w_dff_A_DICIafTn4_2),.clk(gclk));
	jdff dff_A_xKwUIsha4_0(.dout(w_dff_A_u4IoAXrO7_0),.din(w_dff_A_xKwUIsha4_0),.clk(gclk));
	jdff dff_A_u4IoAXrO7_0(.dout(w_dff_A_epYqvhRU1_0),.din(w_dff_A_u4IoAXrO7_0),.clk(gclk));
	jdff dff_A_epYqvhRU1_0(.dout(w_dff_A_6vaKIZ543_0),.din(w_dff_A_epYqvhRU1_0),.clk(gclk));
	jdff dff_A_6vaKIZ543_0(.dout(w_dff_A_MIboaQFw0_0),.din(w_dff_A_6vaKIZ543_0),.clk(gclk));
	jdff dff_A_MIboaQFw0_0(.dout(G324),.din(w_dff_A_MIboaQFw0_0),.clk(gclk));
	jdff dff_A_NQVt2kRm1_2(.dout(w_dff_A_jlQjxoG41_0),.din(w_dff_A_NQVt2kRm1_2),.clk(gclk));
	jdff dff_A_jlQjxoG41_0(.dout(w_dff_A_PmI2oesN5_0),.din(w_dff_A_jlQjxoG41_0),.clk(gclk));
	jdff dff_A_PmI2oesN5_0(.dout(w_dff_A_4Oh98sEY5_0),.din(w_dff_A_PmI2oesN5_0),.clk(gclk));
	jdff dff_A_4Oh98sEY5_0(.dout(w_dff_A_OkWBMWSE1_0),.din(w_dff_A_4Oh98sEY5_0),.clk(gclk));
	jdff dff_A_OkWBMWSE1_0(.dout(w_dff_A_ROJaRKpT5_0),.din(w_dff_A_OkWBMWSE1_0),.clk(gclk));
	jdff dff_A_ROJaRKpT5_0(.dout(w_dff_A_lsQP0g3C9_0),.din(w_dff_A_ROJaRKpT5_0),.clk(gclk));
	jdff dff_A_lsQP0g3C9_0(.dout(w_dff_A_zAtxwbX66_0),.din(w_dff_A_lsQP0g3C9_0),.clk(gclk));
	jdff dff_A_zAtxwbX66_0(.dout(w_dff_A_MsWlgwaZ9_0),.din(w_dff_A_zAtxwbX66_0),.clk(gclk));
	jdff dff_A_MsWlgwaZ9_0(.dout(w_dff_A_ZdlUvHA08_0),.din(w_dff_A_MsWlgwaZ9_0),.clk(gclk));
	jdff dff_A_ZdlUvHA08_0(.dout(G252),.din(w_dff_A_ZdlUvHA08_0),.clk(gclk));
	jdff dff_A_L1Bufp9g1_2(.dout(G276),.din(w_dff_A_L1Bufp9g1_2),.clk(gclk));
	jdff dff_A_lRTJsLNs9_2(.dout(w_dff_A_9SRkHYKg9_0),.din(w_dff_A_lRTJsLNs9_2),.clk(gclk));
	jdff dff_A_9SRkHYKg9_0(.dout(w_dff_A_e3l2gwAl1_0),.din(w_dff_A_9SRkHYKg9_0),.clk(gclk));
	jdff dff_A_e3l2gwAl1_0(.dout(w_dff_A_2iq6fmuY0_0),.din(w_dff_A_e3l2gwAl1_0),.clk(gclk));
	jdff dff_A_2iq6fmuY0_0(.dout(w_dff_A_neslyGTD7_0),.din(w_dff_A_2iq6fmuY0_0),.clk(gclk));
	jdff dff_A_neslyGTD7_0(.dout(w_dff_A_lOWCjw8e4_0),.din(w_dff_A_neslyGTD7_0),.clk(gclk));
	jdff dff_A_lOWCjw8e4_0(.dout(G310),.din(w_dff_A_lOWCjw8e4_0),.clk(gclk));
	jdff dff_A_lnjGnJCt2_2(.dout(w_dff_A_Y5XLu9dj5_0),.din(w_dff_A_lnjGnJCt2_2),.clk(gclk));
	jdff dff_A_Y5XLu9dj5_0(.dout(w_dff_A_eeanR2vx6_0),.din(w_dff_A_Y5XLu9dj5_0),.clk(gclk));
	jdff dff_A_eeanR2vx6_0(.dout(w_dff_A_tYVrD28B9_0),.din(w_dff_A_eeanR2vx6_0),.clk(gclk));
	jdff dff_A_tYVrD28B9_0(.dout(w_dff_A_1W460Dm57_0),.din(w_dff_A_tYVrD28B9_0),.clk(gclk));
	jdff dff_A_1W460Dm57_0(.dout(w_dff_A_BoqqTkn33_0),.din(w_dff_A_1W460Dm57_0),.clk(gclk));
	jdff dff_A_BoqqTkn33_0(.dout(w_dff_A_xQQoHkPH4_0),.din(w_dff_A_BoqqTkn33_0),.clk(gclk));
	jdff dff_A_xQQoHkPH4_0(.dout(G313),.din(w_dff_A_xQQoHkPH4_0),.clk(gclk));
	jdff dff_A_8uxDTvgW9_2(.dout(w_dff_A_cPqXYTE18_0),.din(w_dff_A_8uxDTvgW9_2),.clk(gclk));
	jdff dff_A_cPqXYTE18_0(.dout(w_dff_A_voLhiAm82_0),.din(w_dff_A_cPqXYTE18_0),.clk(gclk));
	jdff dff_A_voLhiAm82_0(.dout(w_dff_A_YHGunLfs7_0),.din(w_dff_A_voLhiAm82_0),.clk(gclk));
	jdff dff_A_YHGunLfs7_0(.dout(w_dff_A_AYxt9uhx6_0),.din(w_dff_A_YHGunLfs7_0),.clk(gclk));
	jdff dff_A_AYxt9uhx6_0(.dout(w_dff_A_JMmm4y7s7_0),.din(w_dff_A_AYxt9uhx6_0),.clk(gclk));
	jdff dff_A_JMmm4y7s7_0(.dout(w_dff_A_R9QbWCVT7_0),.din(w_dff_A_JMmm4y7s7_0),.clk(gclk));
	jdff dff_A_R9QbWCVT7_0(.dout(w_dff_A_AdMTSGkd2_0),.din(w_dff_A_R9QbWCVT7_0),.clk(gclk));
	jdff dff_A_AdMTSGkd2_0(.dout(G316),.din(w_dff_A_AdMTSGkd2_0),.clk(gclk));
	jdff dff_A_msuIofH91_2(.dout(w_dff_A_e7NZZ9Jh9_0),.din(w_dff_A_msuIofH91_2),.clk(gclk));
	jdff dff_A_e7NZZ9Jh9_0(.dout(w_dff_A_WxO82xC60_0),.din(w_dff_A_e7NZZ9Jh9_0),.clk(gclk));
	jdff dff_A_WxO82xC60_0(.dout(w_dff_A_Tgt3uhVB7_0),.din(w_dff_A_WxO82xC60_0),.clk(gclk));
	jdff dff_A_Tgt3uhVB7_0(.dout(w_dff_A_3RsOgYAn2_0),.din(w_dff_A_Tgt3uhVB7_0),.clk(gclk));
	jdff dff_A_3RsOgYAn2_0(.dout(w_dff_A_V2AhAh9a8_0),.din(w_dff_A_3RsOgYAn2_0),.clk(gclk));
	jdff dff_A_V2AhAh9a8_0(.dout(w_dff_A_YUlWv93S3_0),.din(w_dff_A_V2AhAh9a8_0),.clk(gclk));
	jdff dff_A_YUlWv93S3_0(.dout(w_dff_A_WPyjfajw6_0),.din(w_dff_A_YUlWv93S3_0),.clk(gclk));
	jdff dff_A_WPyjfajw6_0(.dout(G319),.din(w_dff_A_WPyjfajw6_0),.clk(gclk));
	jdff dff_A_6shXyOtb9_2(.dout(w_dff_A_TiDOOqkh8_0),.din(w_dff_A_6shXyOtb9_2),.clk(gclk));
	jdff dff_A_TiDOOqkh8_0(.dout(G327),.din(w_dff_A_TiDOOqkh8_0),.clk(gclk));
	jdff dff_A_YJxM6Mt30_2(.dout(w_dff_A_nsAqMw0Q0_0),.din(w_dff_A_YJxM6Mt30_2),.clk(gclk));
	jdff dff_A_nsAqMw0Q0_0(.dout(w_dff_A_FTUK2Itj9_0),.din(w_dff_A_nsAqMw0Q0_0),.clk(gclk));
	jdff dff_A_FTUK2Itj9_0(.dout(G330),.din(w_dff_A_FTUK2Itj9_0),.clk(gclk));
	jdff dff_A_VslLU2ex9_2(.dout(w_dff_A_17APeLJc3_0),.din(w_dff_A_VslLU2ex9_2),.clk(gclk));
	jdff dff_A_17APeLJc3_0(.dout(w_dff_A_Gea5GdIC6_0),.din(w_dff_A_17APeLJc3_0),.clk(gclk));
	jdff dff_A_Gea5GdIC6_0(.dout(w_dff_A_rdoQ9sAy9_0),.din(w_dff_A_Gea5GdIC6_0),.clk(gclk));
	jdff dff_A_rdoQ9sAy9_0(.dout(G333),.din(w_dff_A_rdoQ9sAy9_0),.clk(gclk));
	jdff dff_A_EI1P8NHh9_2(.dout(w_dff_A_iO4BboNG7_0),.din(w_dff_A_EI1P8NHh9_2),.clk(gclk));
	jdff dff_A_iO4BboNG7_0(.dout(w_dff_A_dfsQFtzR5_0),.din(w_dff_A_iO4BboNG7_0),.clk(gclk));
	jdff dff_A_dfsQFtzR5_0(.dout(w_dff_A_vjIvwJmK5_0),.din(w_dff_A_dfsQFtzR5_0),.clk(gclk));
	jdff dff_A_vjIvwJmK5_0(.dout(G336),.din(w_dff_A_vjIvwJmK5_0),.clk(gclk));
	jdff dff_A_zFFMkuIJ3_2(.dout(w_dff_A_hl6VS2nb8_0),.din(w_dff_A_zFFMkuIJ3_2),.clk(gclk));
	jdff dff_A_hl6VS2nb8_0(.dout(w_dff_A_Ti57PiJS2_0),.din(w_dff_A_hl6VS2nb8_0),.clk(gclk));
	jdff dff_A_Ti57PiJS2_0(.dout(w_dff_A_iDKQ5rAz6_0),.din(w_dff_A_Ti57PiJS2_0),.clk(gclk));
	jdff dff_A_iDKQ5rAz6_0(.dout(w_dff_A_ohqNHRVs4_0),.din(w_dff_A_iDKQ5rAz6_0),.clk(gclk));
	jdff dff_A_ohqNHRVs4_0(.dout(w_dff_A_R3tk25Rf5_0),.din(w_dff_A_ohqNHRVs4_0),.clk(gclk));
	jdff dff_A_R3tk25Rf5_0(.dout(w_dff_A_X0BsDltY5_0),.din(w_dff_A_R3tk25Rf5_0),.clk(gclk));
	jdff dff_A_X0BsDltY5_0(.dout(w_dff_A_gT28VCUj6_0),.din(w_dff_A_X0BsDltY5_0),.clk(gclk));
	jdff dff_A_gT28VCUj6_0(.dout(w_dff_A_T9Mmn4g16_0),.din(w_dff_A_gT28VCUj6_0),.clk(gclk));
	jdff dff_A_T9Mmn4g16_0(.dout(w_dff_A_4O1nbhdD6_0),.din(w_dff_A_T9Mmn4g16_0),.clk(gclk));
	jdff dff_A_4O1nbhdD6_0(.dout(w_dff_A_64VC4QjV2_0),.din(w_dff_A_4O1nbhdD6_0),.clk(gclk));
	jdff dff_A_64VC4QjV2_0(.dout(w_dff_A_jsPWeTfS2_0),.din(w_dff_A_64VC4QjV2_0),.clk(gclk));
	jdff dff_A_jsPWeTfS2_0(.dout(G418),.din(w_dff_A_jsPWeTfS2_0),.clk(gclk));
	jdff dff_A_jO93Ve3B1_2(.dout(G273),.din(w_dff_A_jO93Ve3B1_2),.clk(gclk));
	jdff dff_A_OflSHxKU6_2(.dout(w_dff_A_ht6zsPW75_0),.din(w_dff_A_OflSHxKU6_2),.clk(gclk));
	jdff dff_A_ht6zsPW75_0(.dout(w_dff_A_wCB5TBIl1_0),.din(w_dff_A_ht6zsPW75_0),.clk(gclk));
	jdff dff_A_wCB5TBIl1_0(.dout(w_dff_A_7hPEKW9R3_0),.din(w_dff_A_wCB5TBIl1_0),.clk(gclk));
	jdff dff_A_7hPEKW9R3_0(.dout(G298),.din(w_dff_A_7hPEKW9R3_0),.clk(gclk));
	jdff dff_A_dsbSATGu4_2(.dout(w_dff_A_j5V6LuLv2_0),.din(w_dff_A_dsbSATGu4_2),.clk(gclk));
	jdff dff_A_j5V6LuLv2_0(.dout(w_dff_A_OxRSYCGE2_0),.din(w_dff_A_j5V6LuLv2_0),.clk(gclk));
	jdff dff_A_OxRSYCGE2_0(.dout(w_dff_A_ZEQWi1pg4_0),.din(w_dff_A_OxRSYCGE2_0),.clk(gclk));
	jdff dff_A_ZEQWi1pg4_0(.dout(w_dff_A_FvQ315YE3_0),.din(w_dff_A_ZEQWi1pg4_0),.clk(gclk));
	jdff dff_A_FvQ315YE3_0(.dout(w_dff_A_ioHSf3dV1_0),.din(w_dff_A_FvQ315YE3_0),.clk(gclk));
	jdff dff_A_ioHSf3dV1_0(.dout(G301),.din(w_dff_A_ioHSf3dV1_0),.clk(gclk));
	jdff dff_A_5LuU9lJA3_2(.dout(w_dff_A_qX5Ij0Hf0_0),.din(w_dff_A_5LuU9lJA3_2),.clk(gclk));
	jdff dff_A_qX5Ij0Hf0_0(.dout(w_dff_A_SnxBONCb1_0),.din(w_dff_A_qX5Ij0Hf0_0),.clk(gclk));
	jdff dff_A_SnxBONCb1_0(.dout(w_dff_A_Tihw7pkO8_0),.din(w_dff_A_SnxBONCb1_0),.clk(gclk));
	jdff dff_A_Tihw7pkO8_0(.dout(w_dff_A_zi8mZRj11_0),.din(w_dff_A_Tihw7pkO8_0),.clk(gclk));
	jdff dff_A_zi8mZRj11_0(.dout(w_dff_A_J0dSgC1d3_0),.din(w_dff_A_zi8mZRj11_0),.clk(gclk));
	jdff dff_A_J0dSgC1d3_0(.dout(G304),.din(w_dff_A_J0dSgC1d3_0),.clk(gclk));
	jdff dff_A_tQ3YGlOH2_2(.dout(w_dff_A_Wac1H6vR7_0),.din(w_dff_A_tQ3YGlOH2_2),.clk(gclk));
	jdff dff_A_Wac1H6vR7_0(.dout(w_dff_A_igCfawJ90_0),.din(w_dff_A_Wac1H6vR7_0),.clk(gclk));
	jdff dff_A_igCfawJ90_0(.dout(w_dff_A_i7PZ4wdJ2_0),.din(w_dff_A_igCfawJ90_0),.clk(gclk));
	jdff dff_A_i7PZ4wdJ2_0(.dout(w_dff_A_hiKzcPEr7_0),.din(w_dff_A_i7PZ4wdJ2_0),.clk(gclk));
	jdff dff_A_hiKzcPEr7_0(.dout(w_dff_A_EPOat27B7_0),.din(w_dff_A_hiKzcPEr7_0),.clk(gclk));
	jdff dff_A_EPOat27B7_0(.dout(w_dff_A_Wc8PTM7X5_0),.din(w_dff_A_EPOat27B7_0),.clk(gclk));
	jdff dff_A_Wc8PTM7X5_0(.dout(w_dff_A_w934NNeU9_0),.din(w_dff_A_Wc8PTM7X5_0),.clk(gclk));
	jdff dff_A_w934NNeU9_0(.dout(G307),.din(w_dff_A_w934NNeU9_0),.clk(gclk));
	jdff dff_A_sgRaRusK5_2(.dout(w_dff_A_X25iMPm18_0),.din(w_dff_A_sgRaRusK5_2),.clk(gclk));
	jdff dff_A_X25iMPm18_0(.dout(w_dff_A_nw7rdXuS5_0),.din(w_dff_A_X25iMPm18_0),.clk(gclk));
	jdff dff_A_nw7rdXuS5_0(.dout(w_dff_A_BuVOp8gI7_0),.din(w_dff_A_nw7rdXuS5_0),.clk(gclk));
	jdff dff_A_BuVOp8gI7_0(.dout(w_dff_A_scjVvCKs4_0),.din(w_dff_A_BuVOp8gI7_0),.clk(gclk));
	jdff dff_A_scjVvCKs4_0(.dout(w_dff_A_ZhbkMa961_0),.din(w_dff_A_scjVvCKs4_0),.clk(gclk));
	jdff dff_A_ZhbkMa961_0(.dout(w_dff_A_bu91IbJi1_0),.din(w_dff_A_ZhbkMa961_0),.clk(gclk));
	jdff dff_A_bu91IbJi1_0(.dout(w_dff_A_9zik9Kzl7_0),.din(w_dff_A_bu91IbJi1_0),.clk(gclk));
	jdff dff_A_9zik9Kzl7_0(.dout(w_dff_A_BoGFj39m3_0),.din(w_dff_A_9zik9Kzl7_0),.clk(gclk));
	jdff dff_A_BoGFj39m3_0(.dout(w_dff_A_OnCKJ4yS2_0),.din(w_dff_A_BoGFj39m3_0),.clk(gclk));
	jdff dff_A_OnCKJ4yS2_0(.dout(w_dff_A_ByoYz9dA3_0),.din(w_dff_A_OnCKJ4yS2_0),.clk(gclk));
	jdff dff_A_ByoYz9dA3_0(.dout(w_dff_A_fuIUMmUJ9_0),.din(w_dff_A_ByoYz9dA3_0),.clk(gclk));
	jdff dff_A_fuIUMmUJ9_0(.dout(w_dff_A_NUSCYnwC6_0),.din(w_dff_A_fuIUMmUJ9_0),.clk(gclk));
	jdff dff_A_NUSCYnwC6_0(.dout(w_dff_A_Tf9JfhOZ2_0),.din(w_dff_A_NUSCYnwC6_0),.clk(gclk));
	jdff dff_A_Tf9JfhOZ2_0(.dout(G344),.din(w_dff_A_Tf9JfhOZ2_0),.clk(gclk));
	jdff dff_A_0s1VMX2B6_2(.dout(G422),.din(w_dff_A_0s1VMX2B6_2),.clk(gclk));
	jdff dff_A_1dn7niiP8_2(.dout(G469),.din(w_dff_A_1dn7niiP8_2),.clk(gclk));
	jdff dff_A_PDuO5PBw0_2(.dout(w_dff_A_UIpu50357_0),.din(w_dff_A_PDuO5PBw0_2),.clk(gclk));
	jdff dff_A_UIpu50357_0(.dout(w_dff_A_a8GoUbFq1_0),.din(w_dff_A_UIpu50357_0),.clk(gclk));
	jdff dff_A_a8GoUbFq1_0(.dout(w_dff_A_0X2mtHnC4_0),.din(w_dff_A_a8GoUbFq1_0),.clk(gclk));
	jdff dff_A_0X2mtHnC4_0(.dout(G419),.din(w_dff_A_0X2mtHnC4_0),.clk(gclk));
	jdff dff_A_RbZnUKx60_2(.dout(w_dff_A_u16L53ov1_0),.din(w_dff_A_RbZnUKx60_2),.clk(gclk));
	jdff dff_A_u16L53ov1_0(.dout(w_dff_A_jJnlQ8lg5_0),.din(w_dff_A_u16L53ov1_0),.clk(gclk));
	jdff dff_A_jJnlQ8lg5_0(.dout(w_dff_A_PKY98M205_0),.din(w_dff_A_jJnlQ8lg5_0),.clk(gclk));
	jdff dff_A_PKY98M205_0(.dout(G471),.din(w_dff_A_PKY98M205_0),.clk(gclk));
	jdff dff_A_VtwlBwvj4_2(.dout(w_dff_A_MEGQYoZQ8_0),.din(w_dff_A_VtwlBwvj4_2),.clk(gclk));
	jdff dff_A_MEGQYoZQ8_0(.dout(w_dff_A_e0IBh4tV4_0),.din(w_dff_A_MEGQYoZQ8_0),.clk(gclk));
	jdff dff_A_e0IBh4tV4_0(.dout(w_dff_A_He7vKV3m7_0),.din(w_dff_A_e0IBh4tV4_0),.clk(gclk));
	jdff dff_A_He7vKV3m7_0(.dout(w_dff_A_0T4TBg678_0),.din(w_dff_A_He7vKV3m7_0),.clk(gclk));
	jdff dff_A_0T4TBg678_0(.dout(w_dff_A_xrNjMkcD4_0),.din(w_dff_A_0T4TBg678_0),.clk(gclk));
	jdff dff_A_xrNjMkcD4_0(.dout(w_dff_A_FgArA67l2_0),.din(w_dff_A_xrNjMkcD4_0),.clk(gclk));
	jdff dff_A_FgArA67l2_0(.dout(w_dff_A_Ctedzh3r6_0),.din(w_dff_A_FgArA67l2_0),.clk(gclk));
	jdff dff_A_Ctedzh3r6_0(.dout(w_dff_A_lSAJeN7r2_0),.din(w_dff_A_Ctedzh3r6_0),.clk(gclk));
	jdff dff_A_lSAJeN7r2_0(.dout(w_dff_A_LEpBkxa81_0),.din(w_dff_A_lSAJeN7r2_0),.clk(gclk));
	jdff dff_A_LEpBkxa81_0(.dout(G359),.din(w_dff_A_LEpBkxa81_0),.clk(gclk));
	jdff dff_A_cH5sdleA0_2(.dout(w_dff_A_09nyGtJ86_0),.din(w_dff_A_cH5sdleA0_2),.clk(gclk));
	jdff dff_A_09nyGtJ86_0(.dout(w_dff_A_8pW9M11I5_0),.din(w_dff_A_09nyGtJ86_0),.clk(gclk));
	jdff dff_A_8pW9M11I5_0(.dout(w_dff_A_48s4wDcE6_0),.din(w_dff_A_8pW9M11I5_0),.clk(gclk));
	jdff dff_A_48s4wDcE6_0(.dout(w_dff_A_fGvCaisU3_0),.din(w_dff_A_48s4wDcE6_0),.clk(gclk));
	jdff dff_A_fGvCaisU3_0(.dout(w_dff_A_BvwSno8Q0_0),.din(w_dff_A_fGvCaisU3_0),.clk(gclk));
	jdff dff_A_BvwSno8Q0_0(.dout(w_dff_A_cZZqkUzd1_0),.din(w_dff_A_BvwSno8Q0_0),.clk(gclk));
	jdff dff_A_cZZqkUzd1_0(.dout(w_dff_A_bMJesM9S9_0),.din(w_dff_A_cZZqkUzd1_0),.clk(gclk));
	jdff dff_A_bMJesM9S9_0(.dout(w_dff_A_RKJc31Ei8_0),.din(w_dff_A_bMJesM9S9_0),.clk(gclk));
	jdff dff_A_RKJc31Ei8_0(.dout(w_dff_A_jvOeQbXp8_0),.din(w_dff_A_RKJc31Ei8_0),.clk(gclk));
	jdff dff_A_jvOeQbXp8_0(.dout(w_dff_A_j4XNgQ4z2_0),.din(w_dff_A_jvOeQbXp8_0),.clk(gclk));
	jdff dff_A_j4XNgQ4z2_0(.dout(G362),.din(w_dff_A_j4XNgQ4z2_0),.clk(gclk));
	jdff dff_A_lHS6djP02_2(.dout(w_dff_A_mzEkFAxW8_0),.din(w_dff_A_lHS6djP02_2),.clk(gclk));
	jdff dff_A_mzEkFAxW8_0(.dout(w_dff_A_80KpsHq41_0),.din(w_dff_A_mzEkFAxW8_0),.clk(gclk));
	jdff dff_A_80KpsHq41_0(.dout(w_dff_A_XU8B1wjo3_0),.din(w_dff_A_80KpsHq41_0),.clk(gclk));
	jdff dff_A_XU8B1wjo3_0(.dout(w_dff_A_YxbgDcVs8_0),.din(w_dff_A_XU8B1wjo3_0),.clk(gclk));
	jdff dff_A_YxbgDcVs8_0(.dout(w_dff_A_GbWXC90o2_0),.din(w_dff_A_YxbgDcVs8_0),.clk(gclk));
	jdff dff_A_GbWXC90o2_0(.dout(w_dff_A_PKh5xbJl3_0),.din(w_dff_A_GbWXC90o2_0),.clk(gclk));
	jdff dff_A_PKh5xbJl3_0(.dout(w_dff_A_YWOxOlqC7_0),.din(w_dff_A_PKh5xbJl3_0),.clk(gclk));
	jdff dff_A_YWOxOlqC7_0(.dout(w_dff_A_PgydrYl73_0),.din(w_dff_A_YWOxOlqC7_0),.clk(gclk));
	jdff dff_A_PgydrYl73_0(.dout(w_dff_A_c2mZSCEB2_0),.din(w_dff_A_PgydrYl73_0),.clk(gclk));
	jdff dff_A_c2mZSCEB2_0(.dout(w_dff_A_GtHIBI4h7_0),.din(w_dff_A_c2mZSCEB2_0),.clk(gclk));
	jdff dff_A_GtHIBI4h7_0(.dout(w_dff_A_qWsczlr09_0),.din(w_dff_A_GtHIBI4h7_0),.clk(gclk));
	jdff dff_A_qWsczlr09_0(.dout(G365),.din(w_dff_A_qWsczlr09_0),.clk(gclk));
	jdff dff_A_2DLI61aZ0_2(.dout(w_dff_A_ZOJQrSh79_0),.din(w_dff_A_2DLI61aZ0_2),.clk(gclk));
	jdff dff_A_ZOJQrSh79_0(.dout(w_dff_A_dg8uBm2T5_0),.din(w_dff_A_ZOJQrSh79_0),.clk(gclk));
	jdff dff_A_dg8uBm2T5_0(.dout(w_dff_A_itMerj1F4_0),.din(w_dff_A_dg8uBm2T5_0),.clk(gclk));
	jdff dff_A_itMerj1F4_0(.dout(w_dff_A_fY0orbjl7_0),.din(w_dff_A_itMerj1F4_0),.clk(gclk));
	jdff dff_A_fY0orbjl7_0(.dout(w_dff_A_EyeXZHZR0_0),.din(w_dff_A_fY0orbjl7_0),.clk(gclk));
	jdff dff_A_EyeXZHZR0_0(.dout(w_dff_A_XEzsvhyY0_0),.din(w_dff_A_EyeXZHZR0_0),.clk(gclk));
	jdff dff_A_XEzsvhyY0_0(.dout(w_dff_A_UpFqKMfv6_0),.din(w_dff_A_XEzsvhyY0_0),.clk(gclk));
	jdff dff_A_UpFqKMfv6_0(.dout(w_dff_A_PnLwTg464_0),.din(w_dff_A_UpFqKMfv6_0),.clk(gclk));
	jdff dff_A_PnLwTg464_0(.dout(w_dff_A_4B8VkiN93_0),.din(w_dff_A_PnLwTg464_0),.clk(gclk));
	jdff dff_A_4B8VkiN93_0(.dout(w_dff_A_yxBdb8Hu6_0),.din(w_dff_A_4B8VkiN93_0),.clk(gclk));
	jdff dff_A_yxBdb8Hu6_0(.dout(w_dff_A_bYk42HNX2_0),.din(w_dff_A_yxBdb8Hu6_0),.clk(gclk));
	jdff dff_A_bYk42HNX2_0(.dout(G368),.din(w_dff_A_bYk42HNX2_0),.clk(gclk));
	jdff dff_A_1HLKbfCP9_2(.dout(w_dff_A_wgtgLWZW8_0),.din(w_dff_A_1HLKbfCP9_2),.clk(gclk));
	jdff dff_A_wgtgLWZW8_0(.dout(w_dff_A_iEf537ix5_0),.din(w_dff_A_wgtgLWZW8_0),.clk(gclk));
	jdff dff_A_iEf537ix5_0(.dout(w_dff_A_Q5gWqtge2_0),.din(w_dff_A_iEf537ix5_0),.clk(gclk));
	jdff dff_A_Q5gWqtge2_0(.dout(w_dff_A_JQImtExa2_0),.din(w_dff_A_Q5gWqtge2_0),.clk(gclk));
	jdff dff_A_JQImtExa2_0(.dout(w_dff_A_NEAW4X7W2_0),.din(w_dff_A_JQImtExa2_0),.clk(gclk));
	jdff dff_A_NEAW4X7W2_0(.dout(w_dff_A_wfeRvzK13_0),.din(w_dff_A_NEAW4X7W2_0),.clk(gclk));
	jdff dff_A_wfeRvzK13_0(.dout(w_dff_A_NqDqdmRB5_0),.din(w_dff_A_wfeRvzK13_0),.clk(gclk));
	jdff dff_A_NqDqdmRB5_0(.dout(w_dff_A_z5Nuabmv8_0),.din(w_dff_A_NqDqdmRB5_0),.clk(gclk));
	jdff dff_A_z5Nuabmv8_0(.dout(G347),.din(w_dff_A_z5Nuabmv8_0),.clk(gclk));
	jdff dff_A_aUo2VDAg5_2(.dout(w_dff_A_TrFPIPHg7_0),.din(w_dff_A_aUo2VDAg5_2),.clk(gclk));
	jdff dff_A_TrFPIPHg7_0(.dout(w_dff_A_PcdDueST1_0),.din(w_dff_A_TrFPIPHg7_0),.clk(gclk));
	jdff dff_A_PcdDueST1_0(.dout(w_dff_A_y0LHmDNq4_0),.din(w_dff_A_PcdDueST1_0),.clk(gclk));
	jdff dff_A_y0LHmDNq4_0(.dout(w_dff_A_xkssh9pA4_0),.din(w_dff_A_y0LHmDNq4_0),.clk(gclk));
	jdff dff_A_xkssh9pA4_0(.dout(w_dff_A_hYEXsSZI9_0),.din(w_dff_A_xkssh9pA4_0),.clk(gclk));
	jdff dff_A_hYEXsSZI9_0(.dout(w_dff_A_1f6NTWTF5_0),.din(w_dff_A_hYEXsSZI9_0),.clk(gclk));
	jdff dff_A_1f6NTWTF5_0(.dout(w_dff_A_GLZYMKPX6_0),.din(w_dff_A_1f6NTWTF5_0),.clk(gclk));
	jdff dff_A_GLZYMKPX6_0(.dout(w_dff_A_usVh4LIi3_0),.din(w_dff_A_GLZYMKPX6_0),.clk(gclk));
	jdff dff_A_usVh4LIi3_0(.dout(w_dff_A_6suMEec18_0),.din(w_dff_A_usVh4LIi3_0),.clk(gclk));
	jdff dff_A_6suMEec18_0(.dout(G350),.din(w_dff_A_6suMEec18_0),.clk(gclk));
	jdff dff_A_19A0fWNC1_2(.dout(w_dff_A_zGb8EKUl8_0),.din(w_dff_A_19A0fWNC1_2),.clk(gclk));
	jdff dff_A_zGb8EKUl8_0(.dout(w_dff_A_QsYMua8f1_0),.din(w_dff_A_zGb8EKUl8_0),.clk(gclk));
	jdff dff_A_QsYMua8f1_0(.dout(w_dff_A_ak1EzYwz4_0),.din(w_dff_A_QsYMua8f1_0),.clk(gclk));
	jdff dff_A_ak1EzYwz4_0(.dout(w_dff_A_EersNSW51_0),.din(w_dff_A_ak1EzYwz4_0),.clk(gclk));
	jdff dff_A_EersNSW51_0(.dout(w_dff_A_i0DpshIC4_0),.din(w_dff_A_EersNSW51_0),.clk(gclk));
	jdff dff_A_i0DpshIC4_0(.dout(w_dff_A_3aRMGh4s6_0),.din(w_dff_A_i0DpshIC4_0),.clk(gclk));
	jdff dff_A_3aRMGh4s6_0(.dout(w_dff_A_sClgRdwd5_0),.din(w_dff_A_3aRMGh4s6_0),.clk(gclk));
	jdff dff_A_sClgRdwd5_0(.dout(w_dff_A_xEpmNJS08_0),.din(w_dff_A_sClgRdwd5_0),.clk(gclk));
	jdff dff_A_xEpmNJS08_0(.dout(w_dff_A_e2p8uiMa4_0),.din(w_dff_A_xEpmNJS08_0),.clk(gclk));
	jdff dff_A_e2p8uiMa4_0(.dout(G353),.din(w_dff_A_e2p8uiMa4_0),.clk(gclk));
	jdff dff_A_aevorycp8_2(.dout(w_dff_A_1077YN5D5_0),.din(w_dff_A_aevorycp8_2),.clk(gclk));
	jdff dff_A_1077YN5D5_0(.dout(w_dff_A_veBJKOnv9_0),.din(w_dff_A_1077YN5D5_0),.clk(gclk));
	jdff dff_A_veBJKOnv9_0(.dout(w_dff_A_AShsLy0K8_0),.din(w_dff_A_veBJKOnv9_0),.clk(gclk));
	jdff dff_A_AShsLy0K8_0(.dout(w_dff_A_fzvrt9aG6_0),.din(w_dff_A_AShsLy0K8_0),.clk(gclk));
	jdff dff_A_fzvrt9aG6_0(.dout(w_dff_A_GOgkxPyM9_0),.din(w_dff_A_fzvrt9aG6_0),.clk(gclk));
	jdff dff_A_GOgkxPyM9_0(.dout(w_dff_A_z5vZLAli4_0),.din(w_dff_A_GOgkxPyM9_0),.clk(gclk));
	jdff dff_A_z5vZLAli4_0(.dout(w_dff_A_ojR4bByL9_0),.din(w_dff_A_z5vZLAli4_0),.clk(gclk));
	jdff dff_A_ojR4bByL9_0(.dout(w_dff_A_Ln9xXAqo0_0),.din(w_dff_A_ojR4bByL9_0),.clk(gclk));
	jdff dff_A_Ln9xXAqo0_0(.dout(w_dff_A_bMGOpfbj8_0),.din(w_dff_A_Ln9xXAqo0_0),.clk(gclk));
	jdff dff_A_bMGOpfbj8_0(.dout(w_dff_A_LwVQP45A9_0),.din(w_dff_A_bMGOpfbj8_0),.clk(gclk));
	jdff dff_A_LwVQP45A9_0(.dout(w_dff_A_BW82lTQW9_0),.din(w_dff_A_LwVQP45A9_0),.clk(gclk));
	jdff dff_A_BW82lTQW9_0(.dout(G356),.din(w_dff_A_BW82lTQW9_0),.clk(gclk));
	jdff dff_A_AskpEjKv5_2(.dout(w_dff_A_hUBy5dZx3_0),.din(w_dff_A_AskpEjKv5_2),.clk(gclk));
	jdff dff_A_hUBy5dZx3_0(.dout(w_dff_A_OOgoavvw0_0),.din(w_dff_A_hUBy5dZx3_0),.clk(gclk));
	jdff dff_A_OOgoavvw0_0(.dout(w_dff_A_SIxhEd9F4_0),.din(w_dff_A_OOgoavvw0_0),.clk(gclk));
	jdff dff_A_SIxhEd9F4_0(.dout(w_dff_A_QWCoSs815_0),.din(w_dff_A_SIxhEd9F4_0),.clk(gclk));
	jdff dff_A_QWCoSs815_0(.dout(G321),.din(w_dff_A_QWCoSs815_0),.clk(gclk));
	jdff dff_A_Gw55g2Xc2_2(.dout(w_dff_A_PQd8pTif0_0),.din(w_dff_A_Gw55g2Xc2_2),.clk(gclk));
	jdff dff_A_PQd8pTif0_0(.dout(w_dff_A_bDaYB5PH5_0),.din(w_dff_A_PQd8pTif0_0),.clk(gclk));
	jdff dff_A_bDaYB5PH5_0(.dout(w_dff_A_sbLME52K2_0),.din(w_dff_A_bDaYB5PH5_0),.clk(gclk));
	jdff dff_A_sbLME52K2_0(.dout(w_dff_A_iuBjrNUP2_0),.din(w_dff_A_sbLME52K2_0),.clk(gclk));
	jdff dff_A_iuBjrNUP2_0(.dout(w_dff_A_RiPI1zBM8_0),.din(w_dff_A_iuBjrNUP2_0),.clk(gclk));
	jdff dff_A_RiPI1zBM8_0(.dout(w_dff_A_FwPipHHf7_0),.din(w_dff_A_RiPI1zBM8_0),.clk(gclk));
	jdff dff_A_FwPipHHf7_0(.dout(G370),.din(w_dff_A_FwPipHHf7_0),.clk(gclk));
	jdff dff_A_ECMPFZkm5_2(.dout(w_dff_A_zT6qpQjp6_0),.din(w_dff_A_ECMPFZkm5_2),.clk(gclk));
	jdff dff_A_zT6qpQjp6_0(.dout(w_dff_A_q19Fxxip4_0),.din(w_dff_A_zT6qpQjp6_0),.clk(gclk));
	jdff dff_A_q19Fxxip4_0(.dout(w_dff_A_6gic20X58_0),.din(w_dff_A_q19Fxxip4_0),.clk(gclk));
	jdff dff_A_6gic20X58_0(.dout(w_dff_A_gOEE4jEb7_0),.din(w_dff_A_6gic20X58_0),.clk(gclk));
	jdff dff_A_gOEE4jEb7_0(.dout(G399),.din(w_dff_A_gOEE4jEb7_0),.clk(gclk));
endmodule

