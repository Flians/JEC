/*

c6288:
	jxor: 446
	jspl: 940
	jspl3: 260
	jnot: 330
	jdff: 1618
	jand: 683
	jor: 331

Summary:
	jxor: 446
	jspl: 940
	jspl3: 260
	jnot: 330
	jdff: 1618
	jand: 683
	jor: 331

The maximum logic level gap of any gate:
	c6288: 60
*/

module rf_c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G1gat_1;
	wire[2:0] w_G1gat_2;
	wire[2:0] w_G1gat_3;
	wire[2:0] w_G1gat_4;
	wire[2:0] w_G1gat_5;
	wire[2:0] w_G1gat_6;
	wire[1:0] w_G1gat_7;
	wire[2:0] w_G18gat_0;
	wire[2:0] w_G18gat_1;
	wire[2:0] w_G18gat_2;
	wire[2:0] w_G18gat_3;
	wire[2:0] w_G18gat_4;
	wire[2:0] w_G18gat_5;
	wire[2:0] w_G18gat_6;
	wire[2:0] w_G18gat_7;
	wire[2:0] w_G35gat_0;
	wire[2:0] w_G35gat_1;
	wire[2:0] w_G35gat_2;
	wire[2:0] w_G35gat_3;
	wire[2:0] w_G35gat_4;
	wire[2:0] w_G35gat_5;
	wire[2:0] w_G35gat_6;
	wire[2:0] w_G35gat_7;
	wire[2:0] w_G52gat_0;
	wire[2:0] w_G52gat_1;
	wire[2:0] w_G52gat_2;
	wire[2:0] w_G52gat_3;
	wire[2:0] w_G52gat_4;
	wire[2:0] w_G52gat_5;
	wire[2:0] w_G52gat_6;
	wire[2:0] w_G52gat_7;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G69gat_1;
	wire[2:0] w_G69gat_2;
	wire[2:0] w_G69gat_3;
	wire[2:0] w_G69gat_4;
	wire[2:0] w_G69gat_5;
	wire[2:0] w_G69gat_6;
	wire[1:0] w_G69gat_7;
	wire[2:0] w_G86gat_0;
	wire[2:0] w_G86gat_1;
	wire[2:0] w_G86gat_2;
	wire[2:0] w_G86gat_3;
	wire[2:0] w_G86gat_4;
	wire[2:0] w_G86gat_5;
	wire[2:0] w_G86gat_6;
	wire[1:0] w_G86gat_7;
	wire[2:0] w_G103gat_0;
	wire[2:0] w_G103gat_1;
	wire[2:0] w_G103gat_2;
	wire[2:0] w_G103gat_3;
	wire[2:0] w_G103gat_4;
	wire[2:0] w_G103gat_5;
	wire[2:0] w_G103gat_6;
	wire[1:0] w_G103gat_7;
	wire[2:0] w_G120gat_0;
	wire[2:0] w_G120gat_1;
	wire[2:0] w_G120gat_2;
	wire[2:0] w_G120gat_3;
	wire[2:0] w_G120gat_4;
	wire[2:0] w_G120gat_5;
	wire[2:0] w_G120gat_6;
	wire[1:0] w_G120gat_7;
	wire[2:0] w_G137gat_0;
	wire[2:0] w_G137gat_1;
	wire[2:0] w_G137gat_2;
	wire[2:0] w_G137gat_3;
	wire[2:0] w_G137gat_4;
	wire[2:0] w_G137gat_5;
	wire[2:0] w_G137gat_6;
	wire[1:0] w_G137gat_7;
	wire[2:0] w_G154gat_0;
	wire[2:0] w_G154gat_1;
	wire[2:0] w_G154gat_2;
	wire[2:0] w_G154gat_3;
	wire[2:0] w_G154gat_4;
	wire[2:0] w_G154gat_5;
	wire[2:0] w_G154gat_6;
	wire[1:0] w_G154gat_7;
	wire[2:0] w_G171gat_0;
	wire[2:0] w_G171gat_1;
	wire[2:0] w_G171gat_2;
	wire[2:0] w_G171gat_3;
	wire[2:0] w_G171gat_4;
	wire[2:0] w_G171gat_5;
	wire[2:0] w_G171gat_6;
	wire[1:0] w_G171gat_7;
	wire[2:0] w_G188gat_0;
	wire[2:0] w_G188gat_1;
	wire[2:0] w_G188gat_2;
	wire[2:0] w_G188gat_3;
	wire[2:0] w_G188gat_4;
	wire[2:0] w_G188gat_5;
	wire[2:0] w_G188gat_6;
	wire[1:0] w_G188gat_7;
	wire[2:0] w_G205gat_0;
	wire[2:0] w_G205gat_1;
	wire[2:0] w_G205gat_2;
	wire[2:0] w_G205gat_3;
	wire[2:0] w_G205gat_4;
	wire[2:0] w_G205gat_5;
	wire[2:0] w_G205gat_6;
	wire[1:0] w_G205gat_7;
	wire[2:0] w_G222gat_0;
	wire[2:0] w_G222gat_1;
	wire[2:0] w_G222gat_2;
	wire[2:0] w_G222gat_3;
	wire[2:0] w_G222gat_4;
	wire[2:0] w_G222gat_5;
	wire[2:0] w_G222gat_6;
	wire[1:0] w_G222gat_7;
	wire[2:0] w_G239gat_0;
	wire[2:0] w_G239gat_1;
	wire[2:0] w_G239gat_2;
	wire[2:0] w_G239gat_3;
	wire[2:0] w_G239gat_4;
	wire[2:0] w_G239gat_5;
	wire[2:0] w_G239gat_6;
	wire[1:0] w_G239gat_7;
	wire[2:0] w_G256gat_0;
	wire[2:0] w_G256gat_1;
	wire[2:0] w_G256gat_2;
	wire[2:0] w_G256gat_3;
	wire[2:0] w_G256gat_4;
	wire[2:0] w_G256gat_5;
	wire[2:0] w_G256gat_6;
	wire[1:0] w_G256gat_7;
	wire[2:0] w_G273gat_0;
	wire[2:0] w_G273gat_1;
	wire[2:0] w_G273gat_2;
	wire[2:0] w_G273gat_3;
	wire[2:0] w_G273gat_4;
	wire[2:0] w_G273gat_5;
	wire[2:0] w_G273gat_6;
	wire[2:0] w_G273gat_7;
	wire[2:0] w_G290gat_0;
	wire[2:0] w_G290gat_1;
	wire[2:0] w_G290gat_2;
	wire[2:0] w_G290gat_3;
	wire[2:0] w_G290gat_4;
	wire[2:0] w_G290gat_5;
	wire[2:0] w_G290gat_6;
	wire[2:0] w_G290gat_7;
	wire[2:0] w_G307gat_0;
	wire[2:0] w_G307gat_1;
	wire[2:0] w_G307gat_2;
	wire[2:0] w_G307gat_3;
	wire[2:0] w_G307gat_4;
	wire[2:0] w_G307gat_5;
	wire[2:0] w_G307gat_6;
	wire[2:0] w_G307gat_7;
	wire[2:0] w_G324gat_0;
	wire[2:0] w_G324gat_1;
	wire[2:0] w_G324gat_2;
	wire[2:0] w_G324gat_3;
	wire[2:0] w_G324gat_4;
	wire[2:0] w_G324gat_5;
	wire[2:0] w_G324gat_6;
	wire[1:0] w_G324gat_7;
	wire[2:0] w_G341gat_0;
	wire[2:0] w_G341gat_1;
	wire[2:0] w_G341gat_2;
	wire[2:0] w_G341gat_3;
	wire[2:0] w_G341gat_4;
	wire[2:0] w_G341gat_5;
	wire[2:0] w_G341gat_6;
	wire[1:0] w_G341gat_7;
	wire[2:0] w_G358gat_0;
	wire[2:0] w_G358gat_1;
	wire[2:0] w_G358gat_2;
	wire[2:0] w_G358gat_3;
	wire[2:0] w_G358gat_4;
	wire[2:0] w_G358gat_5;
	wire[2:0] w_G358gat_6;
	wire[1:0] w_G358gat_7;
	wire[2:0] w_G375gat_0;
	wire[2:0] w_G375gat_1;
	wire[2:0] w_G375gat_2;
	wire[2:0] w_G375gat_3;
	wire[2:0] w_G375gat_4;
	wire[2:0] w_G375gat_5;
	wire[2:0] w_G375gat_6;
	wire[1:0] w_G375gat_7;
	wire[2:0] w_G392gat_0;
	wire[2:0] w_G392gat_1;
	wire[2:0] w_G392gat_2;
	wire[2:0] w_G392gat_3;
	wire[2:0] w_G392gat_4;
	wire[2:0] w_G392gat_5;
	wire[2:0] w_G392gat_6;
	wire[1:0] w_G392gat_7;
	wire[2:0] w_G409gat_0;
	wire[2:0] w_G409gat_1;
	wire[2:0] w_G409gat_2;
	wire[2:0] w_G409gat_3;
	wire[2:0] w_G409gat_4;
	wire[2:0] w_G409gat_5;
	wire[2:0] w_G409gat_6;
	wire[1:0] w_G409gat_7;
	wire[2:0] w_G426gat_0;
	wire[2:0] w_G426gat_1;
	wire[2:0] w_G426gat_2;
	wire[2:0] w_G426gat_3;
	wire[2:0] w_G426gat_4;
	wire[2:0] w_G426gat_5;
	wire[2:0] w_G426gat_6;
	wire[1:0] w_G426gat_7;
	wire[2:0] w_G443gat_0;
	wire[2:0] w_G443gat_1;
	wire[2:0] w_G443gat_2;
	wire[2:0] w_G443gat_3;
	wire[2:0] w_G443gat_4;
	wire[2:0] w_G443gat_5;
	wire[2:0] w_G443gat_6;
	wire[1:0] w_G443gat_7;
	wire[2:0] w_G460gat_0;
	wire[2:0] w_G460gat_1;
	wire[2:0] w_G460gat_2;
	wire[2:0] w_G460gat_3;
	wire[2:0] w_G460gat_4;
	wire[2:0] w_G460gat_5;
	wire[2:0] w_G460gat_6;
	wire[1:0] w_G460gat_7;
	wire[2:0] w_G477gat_0;
	wire[2:0] w_G477gat_1;
	wire[2:0] w_G477gat_2;
	wire[2:0] w_G477gat_3;
	wire[2:0] w_G477gat_4;
	wire[2:0] w_G477gat_5;
	wire[2:0] w_G477gat_6;
	wire[1:0] w_G477gat_7;
	wire[2:0] w_G494gat_0;
	wire[2:0] w_G494gat_1;
	wire[2:0] w_G494gat_2;
	wire[2:0] w_G494gat_3;
	wire[2:0] w_G494gat_4;
	wire[2:0] w_G494gat_5;
	wire[2:0] w_G494gat_6;
	wire[1:0] w_G494gat_7;
	wire[2:0] w_G511gat_0;
	wire[2:0] w_G511gat_1;
	wire[2:0] w_G511gat_2;
	wire[2:0] w_G511gat_3;
	wire[2:0] w_G511gat_4;
	wire[2:0] w_G511gat_5;
	wire[2:0] w_G511gat_6;
	wire[1:0] w_G511gat_7;
	wire[2:0] w_G528gat_0;
	wire[2:0] w_G528gat_1;
	wire[2:0] w_G528gat_2;
	wire[2:0] w_G528gat_3;
	wire[2:0] w_G528gat_4;
	wire[2:0] w_G528gat_5;
	wire[2:0] w_G528gat_6;
	wire[1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire[1:0] w_n65_0;
	wire[1:0] w_n69_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n72_0;
	wire[1:0] w_n75_0;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[1:0] w_n81_0;
	wire[2:0] w_n82_0;
	wire[1:0] w_n82_1;
	wire[1:0] w_n84_0;
	wire[1:0] w_n85_0;
	wire[1:0] w_n87_0;
	wire[1:0] w_n89_0;
	wire[1:0] w_n93_0;
	wire[1:0] w_n94_0;
	wire[1:0] w_n96_0;
	wire[1:0] w_n99_0;
	wire[2:0] w_n100_0;
	wire[1:0] w_n100_1;
	wire[2:0] w_n101_0;
	wire[1:0] w_n103_0;
	wire[1:0] w_n104_0;
	wire[1:0] w_n107_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n110_0;
	wire[1:0] w_n115_0;
	wire[1:0] w_n116_0;
	wire[2:0] w_n126_0;
	wire[1:0] w_n128_0;
	wire[1:0] w_n129_0;
	wire[1:0] w_n130_0;
	wire[1:0] w_n131_0;
	wire[2:0] w_n132_0;
	wire[2:0] w_n133_0;
	wire[1:0] w_n138_0;
	wire[1:0] w_n139_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n142_0;
	wire[1:0] w_n143_0;
	wire[1:0] w_n145_0;
	wire[1:0] w_n150_0;
	wire[1:0] w_n151_0;
	wire[2:0] w_n156_0;
	wire[1:0] w_n158_0;
	wire[1:0] w_n163_0;
	wire[1:0] w_n165_0;
	wire[1:0] w_n166_0;
	wire[1:0] w_n168_0;
	wire[2:0] w_n169_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n172_0;
	wire[1:0] w_n174_0;
	wire[1:0] w_n175_0;
	wire[1:0] w_n176_0;
	wire[1:0] w_n177_0;
	wire[1:0] w_n178_0;
	wire[1:0] w_n180_0;
	wire[1:0] w_n181_0;
	wire[1:0] w_n183_0;
	wire[1:0] w_n188_0;
	wire[1:0] w_n189_0;
	wire[2:0] w_n194_0;
	wire[1:0] w_n196_0;
	wire[1:0] w_n199_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n207_0;
	wire[1:0] w_n209_0;
	wire[2:0] w_n210_0;
	wire[1:0] w_n210_1;
	wire[1:0] w_n213_0;
	wire[1:0] w_n215_0;
	wire[1:0] w_n216_0;
	wire[1:0] w_n217_0;
	wire[1:0] w_n218_0;
	wire[1:0] w_n219_0;
	wire[1:0] w_n220_0;
	wire[1:0] w_n221_0;
	wire[1:0] w_n223_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n226_0;
	wire[1:0] w_n231_0;
	wire[1:0] w_n232_0;
	wire[2:0] w_n237_0;
	wire[1:0] w_n239_0;
	wire[1:0] w_n242_0;
	wire[1:0] w_n244_0;
	wire[1:0] w_n247_0;
	wire[1:0] w_n249_0;
	wire[1:0] w_n252_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n255_0;
	wire[1:0] w_n257_0;
	wire[2:0] w_n258_0;
	wire[1:0] w_n259_0;
	wire[1:0] w_n261_0;
	wire[1:0] w_n264_0;
	wire[1:0] w_n265_0;
	wire[1:0] w_n266_0;
	wire[1:0] w_n267_0;
	wire[1:0] w_n268_0;
	wire[1:0] w_n269_0;
	wire[1:0] w_n270_0;
	wire[1:0] w_n271_0;
	wire[1:0] w_n272_0;
	wire[1:0] w_n274_0;
	wire[1:0] w_n275_0;
	wire[1:0] w_n277_0;
	wire[1:0] w_n282_0;
	wire[1:0] w_n283_0;
	wire[2:0] w_n288_0;
	wire[1:0] w_n290_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n295_0;
	wire[1:0] w_n298_0;
	wire[1:0] w_n300_0;
	wire[1:0] w_n303_0;
	wire[1:0] w_n305_0;
	wire[1:0] w_n308_0;
	wire[1:0] w_n310_0;
	wire[1:0] w_n311_0;
	wire[1:0] w_n313_0;
	wire[2:0] w_n314_0;
	wire[1:0] w_n315_0;
	wire[1:0] w_n317_0;
	wire[1:0] w_n320_0;
	wire[1:0] w_n321_0;
	wire[1:0] w_n322_0;
	wire[1:0] w_n323_0;
	wire[1:0] w_n324_0;
	wire[1:0] w_n325_0;
	wire[1:0] w_n326_0;
	wire[1:0] w_n327_0;
	wire[1:0] w_n328_0;
	wire[1:0] w_n329_0;
	wire[1:0] w_n330_0;
	wire[1:0] w_n332_0;
	wire[1:0] w_n333_0;
	wire[1:0] w_n335_0;
	wire[1:0] w_n340_0;
	wire[1:0] w_n341_0;
	wire[2:0] w_n346_0;
	wire[1:0] w_n348_0;
	wire[1:0] w_n351_0;
	wire[1:0] w_n353_0;
	wire[1:0] w_n356_0;
	wire[1:0] w_n358_0;
	wire[1:0] w_n361_0;
	wire[1:0] w_n363_0;
	wire[1:0] w_n366_0;
	wire[1:0] w_n368_0;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n373_0;
	wire[1:0] w_n375_0;
	wire[2:0] w_n376_0;
	wire[1:0] w_n377_0;
	wire[1:0] w_n380_0;
	wire[1:0] w_n382_0;
	wire[1:0] w_n383_0;
	wire[1:0] w_n384_0;
	wire[1:0] w_n385_0;
	wire[1:0] w_n386_0;
	wire[1:0] w_n387_0;
	wire[1:0] w_n388_0;
	wire[1:0] w_n389_0;
	wire[1:0] w_n390_0;
	wire[1:0] w_n391_0;
	wire[1:0] w_n392_0;
	wire[1:0] w_n393_0;
	wire[1:0] w_n394_0;
	wire[1:0] w_n396_0;
	wire[1:0] w_n397_0;
	wire[1:0] w_n399_0;
	wire[1:0] w_n404_0;
	wire[1:0] w_n405_0;
	wire[2:0] w_n410_0;
	wire[1:0] w_n412_0;
	wire[1:0] w_n415_0;
	wire[1:0] w_n417_0;
	wire[1:0] w_n420_0;
	wire[1:0] w_n422_0;
	wire[1:0] w_n425_0;
	wire[1:0] w_n427_0;
	wire[1:0] w_n430_0;
	wire[1:0] w_n432_0;
	wire[1:0] w_n435_0;
	wire[1:0] w_n437_0;
	wire[1:0] w_n441_0;
	wire[1:0] w_n442_0;
	wire[1:0] w_n443_0;
	wire[1:0] w_n445_0;
	wire[2:0] w_n446_0;
	wire[1:0] w_n447_0;
	wire[1:0] w_n450_0;
	wire[1:0] w_n452_0;
	wire[1:0] w_n453_0;
	wire[1:0] w_n454_0;
	wire[1:0] w_n455_0;
	wire[1:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[1:0] w_n458_0;
	wire[1:0] w_n459_0;
	wire[1:0] w_n460_0;
	wire[1:0] w_n461_0;
	wire[1:0] w_n462_0;
	wire[1:0] w_n463_0;
	wire[1:0] w_n464_0;
	wire[1:0] w_n465_0;
	wire[1:0] w_n466_0;
	wire[1:0] w_n468_0;
	wire[1:0] w_n469_0;
	wire[1:0] w_n471_0;
	wire[1:0] w_n476_0;
	wire[1:0] w_n477_0;
	wire[2:0] w_n482_0;
	wire[1:0] w_n484_0;
	wire[1:0] w_n487_0;
	wire[1:0] w_n489_0;
	wire[1:0] w_n492_0;
	wire[1:0] w_n494_0;
	wire[1:0] w_n497_0;
	wire[1:0] w_n499_0;
	wire[1:0] w_n502_0;
	wire[1:0] w_n504_0;
	wire[1:0] w_n507_0;
	wire[1:0] w_n509_0;
	wire[1:0] w_n512_0;
	wire[1:0] w_n514_0;
	wire[1:0] w_n518_0;
	wire[1:0] w_n519_0;
	wire[1:0] w_n520_0;
	wire[1:0] w_n522_0;
	wire[2:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n527_0;
	wire[1:0] w_n529_0;
	wire[1:0] w_n530_0;
	wire[1:0] w_n531_0;
	wire[1:0] w_n532_0;
	wire[1:0] w_n533_0;
	wire[1:0] w_n534_0;
	wire[1:0] w_n535_0;
	wire[1:0] w_n536_0;
	wire[1:0] w_n537_0;
	wire[1:0] w_n538_0;
	wire[1:0] w_n539_0;
	wire[1:0] w_n540_0;
	wire[1:0] w_n541_0;
	wire[1:0] w_n542_0;
	wire[1:0] w_n543_0;
	wire[1:0] w_n544_0;
	wire[1:0] w_n545_0;
	wire[1:0] w_n547_0;
	wire[1:0] w_n548_0;
	wire[1:0] w_n550_0;
	wire[1:0] w_n555_0;
	wire[1:0] w_n556_0;
	wire[2:0] w_n561_0;
	wire[1:0] w_n563_0;
	wire[1:0] w_n566_0;
	wire[1:0] w_n568_0;
	wire[1:0] w_n571_0;
	wire[1:0] w_n573_0;
	wire[1:0] w_n576_0;
	wire[1:0] w_n578_0;
	wire[1:0] w_n581_0;
	wire[1:0] w_n583_0;
	wire[1:0] w_n586_0;
	wire[1:0] w_n588_0;
	wire[1:0] w_n591_0;
	wire[1:0] w_n593_0;
	wire[1:0] w_n596_0;
	wire[1:0] w_n598_0;
	wire[1:0] w_n602_0;
	wire[1:0] w_n603_0;
	wire[1:0] w_n604_0;
	wire[1:0] w_n606_0;
	wire[2:0] w_n607_0;
	wire[1:0] w_n608_0;
	wire[1:0] w_n611_0;
	wire[1:0] w_n613_0;
	wire[1:0] w_n614_0;
	wire[1:0] w_n615_0;
	wire[1:0] w_n616_0;
	wire[1:0] w_n617_0;
	wire[1:0] w_n618_0;
	wire[1:0] w_n619_0;
	wire[1:0] w_n620_0;
	wire[1:0] w_n621_0;
	wire[1:0] w_n622_0;
	wire[1:0] w_n623_0;
	wire[1:0] w_n624_0;
	wire[1:0] w_n625_0;
	wire[1:0] w_n626_0;
	wire[1:0] w_n627_0;
	wire[1:0] w_n628_0;
	wire[1:0] w_n629_0;
	wire[1:0] w_n630_0;
	wire[1:0] w_n631_0;
	wire[1:0] w_n633_0;
	wire[1:0] w_n634_0;
	wire[1:0] w_n636_0;
	wire[1:0] w_n641_0;
	wire[1:0] w_n642_0;
	wire[2:0] w_n647_0;
	wire[1:0] w_n649_0;
	wire[1:0] w_n652_0;
	wire[1:0] w_n654_0;
	wire[1:0] w_n657_0;
	wire[1:0] w_n659_0;
	wire[1:0] w_n662_0;
	wire[1:0] w_n664_0;
	wire[1:0] w_n667_0;
	wire[1:0] w_n669_0;
	wire[1:0] w_n672_0;
	wire[1:0] w_n674_0;
	wire[1:0] w_n677_0;
	wire[1:0] w_n679_0;
	wire[1:0] w_n682_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n693_0;
	wire[1:0] w_n694_0;
	wire[2:0] w_n695_0;
	wire[1:0] w_n697_0;
	wire[2:0] w_n698_0;
	wire[1:0] w_n699_0;
	wire[1:0] w_n702_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n705_0;
	wire[1:0] w_n706_0;
	wire[1:0] w_n707_0;
	wire[1:0] w_n708_0;
	wire[1:0] w_n709_0;
	wire[1:0] w_n710_0;
	wire[1:0] w_n711_0;
	wire[1:0] w_n712_0;
	wire[1:0] w_n713_0;
	wire[1:0] w_n714_0;
	wire[1:0] w_n715_0;
	wire[1:0] w_n716_0;
	wire[1:0] w_n717_0;
	wire[1:0] w_n718_0;
	wire[1:0] w_n719_0;
	wire[1:0] w_n720_0;
	wire[1:0] w_n721_0;
	wire[1:0] w_n722_0;
	wire[1:0] w_n723_0;
	wire[1:0] w_n724_0;
	wire[1:0] w_n726_0;
	wire[1:0] w_n727_0;
	wire[1:0] w_n729_0;
	wire[1:0] w_n734_0;
	wire[1:0] w_n735_0;
	wire[2:0] w_n740_0;
	wire[1:0] w_n742_0;
	wire[1:0] w_n745_0;
	wire[1:0] w_n747_0;
	wire[1:0] w_n750_0;
	wire[1:0] w_n752_0;
	wire[1:0] w_n755_0;
	wire[1:0] w_n757_0;
	wire[1:0] w_n760_0;
	wire[1:0] w_n762_0;
	wire[1:0] w_n765_0;
	wire[1:0] w_n767_0;
	wire[1:0] w_n770_0;
	wire[1:0] w_n772_0;
	wire[1:0] w_n775_0;
	wire[1:0] w_n777_0;
	wire[1:0] w_n780_0;
	wire[1:0] w_n782_0;
	wire[1:0] w_n785_0;
	wire[1:0] w_n787_0;
	wire[1:0] w_n791_0;
	wire[1:0] w_n792_0;
	wire[1:0] w_n793_0;
	wire[1:0] w_n795_0;
	wire[2:0] w_n797_0;
	wire[1:0] w_n800_0;
	wire[1:0] w_n802_0;
	wire[1:0] w_n803_0;
	wire[1:0] w_n804_0;
	wire[1:0] w_n805_0;
	wire[1:0] w_n806_0;
	wire[1:0] w_n807_0;
	wire[1:0] w_n808_0;
	wire[1:0] w_n809_0;
	wire[1:0] w_n810_0;
	wire[1:0] w_n811_0;
	wire[1:0] w_n812_0;
	wire[1:0] w_n813_0;
	wire[1:0] w_n814_0;
	wire[1:0] w_n815_0;
	wire[1:0] w_n816_0;
	wire[1:0] w_n817_0;
	wire[1:0] w_n818_0;
	wire[1:0] w_n819_0;
	wire[1:0] w_n820_0;
	wire[1:0] w_n821_0;
	wire[1:0] w_n822_0;
	wire[1:0] w_n823_0;
	wire[1:0] w_n824_0;
	wire[1:0] w_n826_0;
	wire[1:0] w_n827_0;
	wire[1:0] w_n829_0;
	wire[1:0] w_n834_0;
	wire[1:0] w_n835_0;
	wire[1:0] w_n839_0;
	wire[1:0] w_n840_0;
	wire[2:0] w_n844_0;
	wire[1:0] w_n846_0;
	wire[1:0] w_n849_0;
	wire[1:0] w_n851_0;
	wire[1:0] w_n854_0;
	wire[1:0] w_n856_0;
	wire[1:0] w_n859_0;
	wire[1:0] w_n861_0;
	wire[1:0] w_n864_0;
	wire[1:0] w_n866_0;
	wire[1:0] w_n869_0;
	wire[1:0] w_n871_0;
	wire[1:0] w_n874_0;
	wire[1:0] w_n876_0;
	wire[1:0] w_n879_0;
	wire[1:0] w_n881_0;
	wire[1:0] w_n884_0;
	wire[1:0] w_n886_0;
	wire[1:0] w_n889_0;
	wire[1:0] w_n891_0;
	wire[1:0] w_n895_0;
	wire[1:0] w_n896_0;
	wire[1:0] w_n897_0;
	wire[1:0] w_n898_0;
	wire[1:0] w_n901_0;
	wire[1:0] w_n903_0;
	wire[1:0] w_n906_0;
	wire[1:0] w_n907_0;
	wire[1:0] w_n908_0;
	wire[1:0] w_n909_0;
	wire[1:0] w_n910_0;
	wire[1:0] w_n911_0;
	wire[1:0] w_n912_0;
	wire[1:0] w_n913_0;
	wire[1:0] w_n914_0;
	wire[1:0] w_n915_0;
	wire[1:0] w_n916_0;
	wire[1:0] w_n917_0;
	wire[1:0] w_n918_0;
	wire[1:0] w_n919_0;
	wire[1:0] w_n920_0;
	wire[1:0] w_n921_0;
	wire[1:0] w_n922_0;
	wire[1:0] w_n923_0;
	wire[1:0] w_n924_0;
	wire[1:0] w_n925_0;
	wire[1:0] w_n926_0;
	wire[2:0] w_n927_0;
	wire[1:0] w_n929_0;
	wire[1:0] w_n930_0;
	wire[1:0] w_n931_0;
	wire[1:0] w_n932_0;
	wire[1:0] w_n937_0;
	wire[1:0] w_n938_0;
	wire[2:0] w_n942_0;
	wire[1:0] w_n943_0;
	wire[1:0] w_n949_0;
	wire[1:0] w_n951_0;
	wire[1:0] w_n954_0;
	wire[1:0] w_n956_0;
	wire[1:0] w_n959_0;
	wire[1:0] w_n961_0;
	wire[1:0] w_n964_0;
	wire[1:0] w_n966_0;
	wire[1:0] w_n969_0;
	wire[1:0] w_n971_0;
	wire[1:0] w_n974_0;
	wire[1:0] w_n976_0;
	wire[1:0] w_n979_0;
	wire[1:0] w_n981_0;
	wire[1:0] w_n984_0;
	wire[1:0] w_n986_0;
	wire[1:0] w_n989_0;
	wire[1:0] w_n991_0;
	wire[1:0] w_n994_0;
	wire[1:0] w_n996_0;
	wire[1:0] w_n999_0;
	wire[1:0] w_n1001_0;
	wire[1:0] w_n1005_0;
	wire[1:0] w_n1006_0;
	wire[1:0] w_n1008_0;
	wire[1:0] w_n1009_0;
	wire[1:0] w_n1010_0;
	wire[1:0] w_n1011_0;
	wire[1:0] w_n1012_0;
	wire[1:0] w_n1013_0;
	wire[1:0] w_n1014_0;
	wire[1:0] w_n1015_0;
	wire[1:0] w_n1016_0;
	wire[1:0] w_n1017_0;
	wire[1:0] w_n1018_0;
	wire[1:0] w_n1019_0;
	wire[1:0] w_n1020_0;
	wire[1:0] w_n1021_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1023_0;
	wire[1:0] w_n1024_0;
	wire[1:0] w_n1025_0;
	wire[1:0] w_n1026_0;
	wire[1:0] w_n1027_0;
	wire[1:0] w_n1028_0;
	wire[1:0] w_n1029_0;
	wire[1:0] w_n1030_0;
	wire[1:0] w_n1031_0;
	wire[1:0] w_n1032_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1034_0;
	wire[1:0] w_n1035_0;
	wire[1:0] w_n1037_0;
	wire[1:0] w_n1039_0;
	wire[1:0] w_n1043_0;
	wire[1:0] w_n1044_0;
	wire[1:0] w_n1048_0;
	wire[1:0] w_n1049_0;
	wire[1:0] w_n1052_0;
	wire[1:0] w_n1054_0;
	wire[1:0] w_n1057_0;
	wire[1:0] w_n1059_0;
	wire[1:0] w_n1062_0;
	wire[1:0] w_n1064_0;
	wire[1:0] w_n1067_0;
	wire[1:0] w_n1069_0;
	wire[1:0] w_n1072_0;
	wire[1:0] w_n1074_0;
	wire[1:0] w_n1077_0;
	wire[1:0] w_n1079_0;
	wire[1:0] w_n1082_0;
	wire[1:0] w_n1084_0;
	wire[1:0] w_n1087_0;
	wire[1:0] w_n1089_0;
	wire[1:0] w_n1092_0;
	wire[1:0] w_n1094_0;
	wire[1:0] w_n1097_0;
	wire[1:0] w_n1099_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1103_0;
	wire[1:0] w_n1109_0;
	wire[1:0] w_n1110_0;
	wire[1:0] w_n1114_0;
	wire[1:0] w_n1115_0;
	wire[1:0] w_n1116_0;
	wire[1:0] w_n1117_0;
	wire[1:0] w_n1118_0;
	wire[1:0] w_n1119_0;
	wire[1:0] w_n1120_0;
	wire[1:0] w_n1121_0;
	wire[1:0] w_n1122_0;
	wire[1:0] w_n1123_0;
	wire[1:0] w_n1124_0;
	wire[1:0] w_n1125_0;
	wire[1:0] w_n1126_0;
	wire[1:0] w_n1127_0;
	wire[1:0] w_n1128_0;
	wire[1:0] w_n1129_0;
	wire[1:0] w_n1130_0;
	wire[1:0] w_n1131_0;
	wire[1:0] w_n1132_0;
	wire[1:0] w_n1133_0;
	wire[1:0] w_n1134_0;
	wire[1:0] w_n1135_0;
	wire[1:0] w_n1137_0;
	wire[1:0] w_n1138_0;
	wire[1:0] w_n1139_0;
	wire[1:0] w_n1140_0;
	wire[1:0] w_n1141_0;
	wire[1:0] w_n1147_0;
	wire[1:0] w_n1151_0;
	wire[1:0] w_n1152_0;
	wire[1:0] w_n1156_0;
	wire[1:0] w_n1158_0;
	wire[1:0] w_n1161_0;
	wire[1:0] w_n1163_0;
	wire[1:0] w_n1166_0;
	wire[1:0] w_n1168_0;
	wire[1:0] w_n1171_0;
	wire[1:0] w_n1173_0;
	wire[1:0] w_n1176_0;
	wire[1:0] w_n1178_0;
	wire[1:0] w_n1181_0;
	wire[1:0] w_n1183_0;
	wire[1:0] w_n1186_0;
	wire[1:0] w_n1188_0;
	wire[1:0] w_n1191_0;
	wire[1:0] w_n1193_0;
	wire[1:0] w_n1196_0;
	wire[1:0] w_n1198_0;
	wire[1:0] w_n1201_0;
	wire[1:0] w_n1203_0;
	wire[1:0] w_n1206_0;
	wire[1:0] w_n1207_0;
	wire[1:0] w_n1208_0;
	wire[1:0] w_n1210_0;
	wire[1:0] w_n1212_0;
	wire[1:0] w_n1213_0;
	wire[1:0] w_n1214_0;
	wire[1:0] w_n1215_0;
	wire[1:0] w_n1216_0;
	wire[1:0] w_n1217_0;
	wire[1:0] w_n1218_0;
	wire[1:0] w_n1219_0;
	wire[1:0] w_n1220_0;
	wire[1:0] w_n1221_0;
	wire[1:0] w_n1222_0;
	wire[1:0] w_n1223_0;
	wire[1:0] w_n1224_0;
	wire[1:0] w_n1225_0;
	wire[1:0] w_n1226_0;
	wire[1:0] w_n1227_0;
	wire[1:0] w_n1228_0;
	wire[1:0] w_n1229_0;
	wire[1:0] w_n1230_0;
	wire[1:0] w_n1231_0;
	wire[1:0] w_n1232_0;
	wire[1:0] w_n1234_0;
	wire[1:0] w_n1236_0;
	wire[1:0] w_n1237_0;
	wire[1:0] w_n1238_0;
	wire[1:0] w_n1244_0;
	wire[1:0] w_n1247_0;
	wire[1:0] w_n1248_0;
	wire[1:0] w_n1251_0;
	wire[1:0] w_n1253_0;
	wire[1:0] w_n1256_0;
	wire[1:0] w_n1258_0;
	wire[1:0] w_n1261_0;
	wire[1:0] w_n1263_0;
	wire[1:0] w_n1266_0;
	wire[1:0] w_n1268_0;
	wire[1:0] w_n1271_0;
	wire[1:0] w_n1273_0;
	wire[1:0] w_n1276_0;
	wire[1:0] w_n1278_0;
	wire[1:0] w_n1281_0;
	wire[1:0] w_n1283_0;
	wire[1:0] w_n1286_0;
	wire[1:0] w_n1288_0;
	wire[1:0] w_n1291_0;
	wire[1:0] w_n1293_0;
	wire[1:0] w_n1296_0;
	wire[1:0] w_n1297_0;
	wire[1:0] w_n1298_0;
	wire[1:0] w_n1301_0;
	wire[1:0] w_n1303_0;
	wire[1:0] w_n1304_0;
	wire[1:0] w_n1305_0;
	wire[1:0] w_n1306_0;
	wire[1:0] w_n1307_0;
	wire[1:0] w_n1308_0;
	wire[1:0] w_n1309_0;
	wire[1:0] w_n1310_0;
	wire[1:0] w_n1311_0;
	wire[1:0] w_n1312_0;
	wire[1:0] w_n1313_0;
	wire[1:0] w_n1314_0;
	wire[1:0] w_n1315_0;
	wire[1:0] w_n1316_0;
	wire[1:0] w_n1317_0;
	wire[1:0] w_n1318_0;
	wire[1:0] w_n1319_0;
	wire[1:0] w_n1320_0;
	wire[1:0] w_n1321_0;
	wire[1:0] w_n1322_0;
	wire[1:0] w_n1324_0;
	wire[1:0] w_n1325_0;
	wire[1:0] w_n1326_0;
	wire[1:0] w_n1332_0;
	wire[1:0] w_n1337_0;
	wire[1:0] w_n1338_0;
	wire[1:0] w_n1341_0;
	wire[1:0] w_n1343_0;
	wire[1:0] w_n1346_0;
	wire[1:0] w_n1348_0;
	wire[1:0] w_n1351_0;
	wire[1:0] w_n1353_0;
	wire[1:0] w_n1356_0;
	wire[1:0] w_n1358_0;
	wire[1:0] w_n1361_0;
	wire[1:0] w_n1363_0;
	wire[1:0] w_n1366_0;
	wire[1:0] w_n1368_0;
	wire[1:0] w_n1371_0;
	wire[1:0] w_n1373_0;
	wire[1:0] w_n1376_0;
	wire[1:0] w_n1378_0;
	wire[1:0] w_n1381_0;
	wire[1:0] w_n1382_0;
	wire[1:0] w_n1383_0;
	wire[1:0] w_n1386_0;
	wire[1:0] w_n1388_0;
	wire[1:0] w_n1389_0;
	wire[1:0] w_n1390_0;
	wire[1:0] w_n1391_0;
	wire[1:0] w_n1392_0;
	wire[1:0] w_n1393_0;
	wire[1:0] w_n1394_0;
	wire[1:0] w_n1395_0;
	wire[1:0] w_n1396_0;
	wire[1:0] w_n1397_0;
	wire[1:0] w_n1398_0;
	wire[1:0] w_n1399_0;
	wire[1:0] w_n1400_0;
	wire[1:0] w_n1401_0;
	wire[1:0] w_n1402_0;
	wire[1:0] w_n1403_0;
	wire[1:0] w_n1404_0;
	wire[1:0] w_n1405_0;
	wire[1:0] w_n1407_0;
	wire[1:0] w_n1409_0;
	wire[1:0] w_n1410_0;
	wire[1:0] w_n1415_0;
	wire[1:0] w_n1420_0;
	wire[1:0] w_n1421_0;
	wire[1:0] w_n1424_0;
	wire[1:0] w_n1426_0;
	wire[1:0] w_n1429_0;
	wire[1:0] w_n1431_0;
	wire[1:0] w_n1434_0;
	wire[1:0] w_n1436_0;
	wire[1:0] w_n1439_0;
	wire[1:0] w_n1441_0;
	wire[1:0] w_n1444_0;
	wire[1:0] w_n1446_0;
	wire[1:0] w_n1449_0;
	wire[1:0] w_n1451_0;
	wire[1:0] w_n1454_0;
	wire[1:0] w_n1456_0;
	wire[1:0] w_n1459_0;
	wire[1:0] w_n1460_0;
	wire[1:0] w_n1461_0;
	wire[1:0] w_n1464_0;
	wire[1:0] w_n1466_0;
	wire[1:0] w_n1467_0;
	wire[1:0] w_n1468_0;
	wire[1:0] w_n1469_0;
	wire[1:0] w_n1470_0;
	wire[1:0] w_n1471_0;
	wire[1:0] w_n1472_0;
	wire[1:0] w_n1473_0;
	wire[1:0] w_n1474_0;
	wire[1:0] w_n1475_0;
	wire[1:0] w_n1476_0;
	wire[1:0] w_n1477_0;
	wire[1:0] w_n1478_0;
	wire[1:0] w_n1479_0;
	wire[1:0] w_n1480_0;
	wire[1:0] w_n1481_0;
	wire[1:0] w_n1483_0;
	wire[1:0] w_n1485_0;
	wire[1:0] w_n1486_0;
	wire[1:0] w_n1491_0;
	wire[1:0] w_n1496_0;
	wire[1:0] w_n1497_0;
	wire[1:0] w_n1500_0;
	wire[1:0] w_n1502_0;
	wire[1:0] w_n1505_0;
	wire[1:0] w_n1507_0;
	wire[1:0] w_n1510_0;
	wire[1:0] w_n1512_0;
	wire[1:0] w_n1515_0;
	wire[1:0] w_n1517_0;
	wire[1:0] w_n1520_0;
	wire[1:0] w_n1522_0;
	wire[1:0] w_n1525_0;
	wire[1:0] w_n1527_0;
	wire[1:0] w_n1530_0;
	wire[1:0] w_n1531_0;
	wire[1:0] w_n1532_0;
	wire[1:0] w_n1535_0;
	wire[1:0] w_n1537_0;
	wire[1:0] w_n1538_0;
	wire[1:0] w_n1539_0;
	wire[1:0] w_n1540_0;
	wire[1:0] w_n1541_0;
	wire[1:0] w_n1542_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1544_0;
	wire[1:0] w_n1545_0;
	wire[1:0] w_n1546_0;
	wire[1:0] w_n1547_0;
	wire[1:0] w_n1548_0;
	wire[1:0] w_n1549_0;
	wire[1:0] w_n1550_0;
	wire[1:0] w_n1552_0;
	wire[1:0] w_n1554_0;
	wire[1:0] w_n1555_0;
	wire[1:0] w_n1560_0;
	wire[1:0] w_n1565_0;
	wire[1:0] w_n1566_0;
	wire[1:0] w_n1569_0;
	wire[1:0] w_n1571_0;
	wire[1:0] w_n1574_0;
	wire[1:0] w_n1576_0;
	wire[1:0] w_n1579_0;
	wire[1:0] w_n1581_0;
	wire[1:0] w_n1584_0;
	wire[1:0] w_n1586_0;
	wire[1:0] w_n1589_0;
	wire[1:0] w_n1591_0;
	wire[1:0] w_n1594_0;
	wire[1:0] w_n1595_0;
	wire[1:0] w_n1596_0;
	wire[1:0] w_n1599_0;
	wire[1:0] w_n1601_0;
	wire[1:0] w_n1602_0;
	wire[1:0] w_n1603_0;
	wire[1:0] w_n1604_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1606_0;
	wire[1:0] w_n1607_0;
	wire[1:0] w_n1608_0;
	wire[1:0] w_n1609_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1611_0;
	wire[1:0] w_n1612_0;
	wire[1:0] w_n1614_0;
	wire[1:0] w_n1616_0;
	wire[1:0] w_n1617_0;
	wire[1:0] w_n1622_0;
	wire[1:0] w_n1627_0;
	wire[1:0] w_n1628_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1633_0;
	wire[1:0] w_n1636_0;
	wire[1:0] w_n1638_0;
	wire[1:0] w_n1641_0;
	wire[1:0] w_n1643_0;
	wire[1:0] w_n1646_0;
	wire[1:0] w_n1648_0;
	wire[1:0] w_n1651_0;
	wire[1:0] w_n1652_0;
	wire[1:0] w_n1653_0;
	wire[1:0] w_n1656_0;
	wire[1:0] w_n1658_0;
	wire[1:0] w_n1659_0;
	wire[1:0] w_n1660_0;
	wire[1:0] w_n1661_0;
	wire[1:0] w_n1662_0;
	wire[1:0] w_n1663_0;
	wire[1:0] w_n1664_0;
	wire[1:0] w_n1665_0;
	wire[1:0] w_n1666_0;
	wire[1:0] w_n1667_0;
	wire[1:0] w_n1669_0;
	wire[1:0] w_n1671_0;
	wire[1:0] w_n1672_0;
	wire[1:0] w_n1677_0;
	wire[1:0] w_n1682_0;
	wire[1:0] w_n1684_0;
	wire[1:0] w_n1687_0;
	wire[1:0] w_n1689_0;
	wire[1:0] w_n1692_0;
	wire[1:0] w_n1694_0;
	wire[1:0] w_n1697_0;
	wire[1:0] w_n1699_0;
	wire[1:0] w_n1702_0;
	wire[1:0] w_n1703_0;
	wire[1:0] w_n1704_0;
	wire[1:0] w_n1707_0;
	wire[1:0] w_n1709_0;
	wire[1:0] w_n1710_0;
	wire[1:0] w_n1711_0;
	wire[1:0] w_n1712_0;
	wire[1:0] w_n1713_0;
	wire[1:0] w_n1714_0;
	wire[1:0] w_n1715_0;
	wire[1:0] w_n1716_0;
	wire[1:0] w_n1717_0;
	wire[1:0] w_n1719_0;
	wire[1:0] w_n1720_0;
	wire[1:0] w_n1725_0;
	wire[1:0] w_n1728_0;
	wire[1:0] w_n1730_0;
	wire[1:0] w_n1733_0;
	wire[1:0] w_n1735_0;
	wire[1:0] w_n1738_0;
	wire[1:0] w_n1740_0;
	wire[1:0] w_n1743_0;
	wire[1:0] w_n1744_0;
	wire[1:0] w_n1745_0;
	wire[1:0] w_n1748_0;
	wire[1:0] w_n1750_0;
	wire[1:0] w_n1751_0;
	wire[1:0] w_n1752_0;
	wire[1:0] w_n1753_0;
	wire[1:0] w_n1754_0;
	wire[1:0] w_n1755_0;
	wire[1:0] w_n1756_0;
	wire[1:0] w_n1757_0;
	wire[1:0] w_n1758_0;
	wire[1:0] w_n1765_0;
	wire[1:0] w_n1768_0;
	wire[1:0] w_n1770_0;
	wire[1:0] w_n1773_0;
	wire[1:0] w_n1775_0;
	wire[1:0] w_n1778_0;
	wire[1:0] w_n1779_0;
	wire[1:0] w_n1780_0;
	wire[1:0] w_n1783_0;
	wire[1:0] w_n1785_0;
	wire[1:0] w_n1786_0;
	wire[1:0] w_n1787_0;
	wire[1:0] w_n1788_0;
	wire[1:0] w_n1789_0;
	wire[1:0] w_n1790_0;
	wire[1:0] w_n1791_0;
	wire[1:0] w_n1798_0;
	wire[1:0] w_n1801_0;
	wire[1:0] w_n1803_0;
	wire[1:0] w_n1806_0;
	wire[1:0] w_n1807_0;
	wire[1:0] w_n1808_0;
	wire[1:0] w_n1811_0;
	wire[1:0] w_n1813_0;
	wire[1:0] w_n1814_0;
	wire[1:0] w_n1815_0;
	wire[1:0] w_n1816_0;
	wire[1:0] w_n1817_0;
	wire[1:0] w_n1824_0;
	wire[1:0] w_n1827_0;
	wire[1:0] w_n1828_0;
	wire[1:0] w_n1829_0;
	wire[1:0] w_n1832_0;
	wire[1:0] w_n1834_0;
	wire[1:0] w_n1835_0;
	wire[1:0] w_n1836_0;
	wire[1:0] w_n1838_0;
	wire[1:0] w_n1841_0;
	wire[1:0] w_n1848_0;
	wire[1:0] w_n1849_0;
	wire w_dff_B_bbppiPhb7_1;
	wire w_dff_B_AvIxvPmF5_1;
	wire w_dff_B_jTjV4pz17_1;
	wire w_dff_B_0LjNHhat3_1;
	wire w_dff_B_FZ3q2YcR3_1;
	wire w_dff_B_qcojHCOn8_1;
	wire w_dff_B_bDc5GmoL9_1;
	wire w_dff_B_5ukqYSMc0_1;
	wire w_dff_B_migKC2OD1_1;
	wire w_dff_B_U7JZyBM13_1;
	wire w_dff_B_Y2Q3omrR4_1;
	wire w_dff_B_PgYh4dwy6_1;
	wire w_dff_B_v0ge0q491_1;
	wire w_dff_B_hAehoMhR4_1;
	wire w_dff_B_p9QM19To9_1;
	wire w_dff_B_UJv3YTAA8_1;
	wire w_dff_B_rggcB22Q3_1;
	wire w_dff_B_6N3bllvZ7_1;
	wire w_dff_B_5rTwhrzE4_1;
	wire w_dff_B_tOmEsRbI4_1;
	wire w_dff_B_JhvV744d7_1;
	wire w_dff_B_yn8sG5gV0_1;
	wire w_dff_B_rTAhQaIy5_1;
	wire w_dff_B_CmYDUPhJ4_1;
	wire w_dff_B_Upm07QLC4_1;
	wire w_dff_B_proUJcUP0_1;
	wire w_dff_B_aOGmcA4y5_1;
	wire w_dff_B_YcYBpuWM3_1;
	wire w_dff_B_XRvb5gxl5_1;
	wire w_dff_B_fwhTfTdf5_1;
	wire w_dff_B_u4htHALd8_1;
	wire w_dff_B_aFy0JXQc9_1;
	wire w_dff_B_gW3FhgDb6_1;
	wire w_dff_B_0aYWqcgP5_1;
	wire w_dff_B_mpRUR74K0_1;
	wire w_dff_B_c68VdqjT0_1;
	wire w_dff_B_HnOS8sg78_1;
	wire w_dff_B_87qx4Hrz1_1;
	wire w_dff_B_6cDtbgj96_1;
	wire w_dff_B_30443sQP7_1;
	wire w_dff_B_hYOv1wcl4_1;
	wire w_dff_B_5y8ARYGA0_1;
	wire w_dff_B_kxKSSoxD1_1;
	wire w_dff_B_E57Rn5bm7_1;
	wire w_dff_B_TyH78zMm2_1;
	wire w_dff_B_KNzEJ7Tm8_1;
	wire w_dff_B_iK6D8GFi2_1;
	wire w_dff_B_kIZuIE5P6_1;
	wire w_dff_B_6CwcnaX19_1;
	wire w_dff_B_qN1tNO329_1;
	wire w_dff_B_6oZvyY0P2_1;
	wire w_dff_B_OxDLKM6A4_1;
	wire w_dff_B_oxBe3N5y3_1;
	wire w_dff_B_SjcxDkzW4_1;
	wire w_dff_B_eoiU48Fu6_1;
	wire w_dff_B_dyi3x6cZ1_1;
	wire w_dff_B_MkWRSGne5_1;
	wire w_dff_B_4nkAMVf06_1;
	wire w_dff_B_g9msoVzN5_1;
	wire w_dff_B_s1gSvCsW5_1;
	wire w_dff_B_Q4crtiAT9_1;
	wire w_dff_B_xzZGX8Mf4_1;
	wire w_dff_B_8DqYEO6r5_1;
	wire w_dff_B_fY2PG9Q50_1;
	wire w_dff_B_WEE1FcfJ1_1;
	wire w_dff_B_3sZshMf70_1;
	wire w_dff_B_ltcvYspb2_1;
	wire w_dff_B_ZWVFB0pd8_1;
	wire w_dff_B_2MNp1Nwe7_1;
	wire w_dff_B_4L0Rtspp9_1;
	wire w_dff_B_qR4ebJi07_1;
	wire w_dff_B_V0FnKv5p0_1;
	wire w_dff_B_0JgJWV5x0_1;
	wire w_dff_B_fddkuUJa3_1;
	wire w_dff_B_Xpk1Nv1t8_1;
	wire w_dff_B_GhC6Xt7D1_1;
	wire w_dff_B_sLNvUs3e8_1;
	wire w_dff_B_GJA0rymt0_1;
	wire w_dff_B_tQMba3r72_1;
	wire w_dff_B_yXcJsc5P4_1;
	wire w_dff_B_shhv4Tye1_1;
	wire w_dff_B_XbVzYS2p8_1;
	wire w_dff_B_37AB7eTi2_1;
	wire w_dff_B_QouHpRJl8_1;
	wire w_dff_B_WBt48WoY6_1;
	wire w_dff_B_TgCdYDGj2_1;
	wire w_dff_B_5yhAp5iP6_1;
	wire w_dff_B_dcbNGr257_1;
	wire w_dff_B_C4gKgDTb4_1;
	wire w_dff_B_t9FLso1H6_1;
	wire w_dff_B_qUc528Iy9_1;
	wire w_dff_B_kbrQWFFZ8_1;
	wire w_dff_B_Yo3uftzK8_1;
	wire w_dff_B_DoPaIDCY3_1;
	wire w_dff_B_q0g7copr0_1;
	wire w_dff_B_r2JZQDKa6_1;
	wire w_dff_B_dXVPzbuD2_1;
	wire w_dff_B_l6ibNJLf0_1;
	wire w_dff_B_naw2xN6C7_1;
	wire w_dff_B_Nksj6Jr94_1;
	wire w_dff_B_ugtd4XIZ5_1;
	wire w_dff_B_FDdO9CcS1_1;
	wire w_dff_B_S9iSXbef9_1;
	wire w_dff_B_1dURD0NL3_1;
	wire w_dff_B_ICEp6Czp6_1;
	wire w_dff_B_P02rJtwH9_1;
	wire w_dff_B_YDKnW1wb3_1;
	wire w_dff_B_xJZCAaJe5_1;
	wire w_dff_B_3chGe1H86_1;
	wire w_dff_B_toAbKKVg2_1;
	wire w_dff_B_cSgI2MDr0_1;
	wire w_dff_B_oyzKLNjM5_1;
	wire w_dff_B_9RlXIP708_1;
	wire w_dff_B_aFmFTcfr2_1;
	wire w_dff_B_A60PPsHR6_1;
	wire w_dff_B_9GIUgHZk6_1;
	wire w_dff_B_ij0Oc1JR6_1;
	wire w_dff_B_S9Jtk2y21_1;
	wire w_dff_B_dCUpUq7u1_1;
	wire w_dff_B_UK7e50Xv1_1;
	wire w_dff_B_P2Tdt8LC4_1;
	wire w_dff_B_9otp8oGy8_1;
	wire w_dff_B_QqXGKpnH8_1;
	wire w_dff_B_HhtfZ3Z65_1;
	wire w_dff_B_CZorwbve9_1;
	wire w_dff_B_0xT7CAzJ5_1;
	wire w_dff_B_ZKuaVAcV6_1;
	wire w_dff_B_7FgAbger1_1;
	wire w_dff_B_Mzox2m156_1;
	wire w_dff_B_R6CM2PpY5_1;
	wire w_dff_B_Q2Jfq5qy7_1;
	wire w_dff_B_BCMy1xRw9_1;
	wire w_dff_B_uYwllOdJ1_1;
	wire w_dff_B_0HJtWpZl3_1;
	wire w_dff_B_7mwDdNrj3_1;
	wire w_dff_B_tgQZfhrL0_1;
	wire w_dff_B_Ff3fkwRn6_1;
	wire w_dff_B_C1KqM5Zq9_1;
	wire w_dff_B_SjOWITER0_1;
	wire w_dff_B_tTrZGqmv4_1;
	wire w_dff_B_ld6u9pkR6_1;
	wire w_dff_B_PWPgwCeY7_1;
	wire w_dff_B_RWF06jY82_1;
	wire w_dff_B_Mcjq08GE7_1;
	wire w_dff_B_igGtsUuN6_1;
	wire w_dff_B_eRqVPqVl8_1;
	wire w_dff_B_F8tX5Snw8_1;
	wire w_dff_B_d2JEphAb6_1;
	wire w_dff_B_xKaeNnVZ8_1;
	wire w_dff_B_QHvZffoJ2_1;
	wire w_dff_B_49orrsqK4_1;
	wire w_dff_B_a80AzxBE0_1;
	wire w_dff_B_U6pCYpOd8_1;
	wire w_dff_B_JgoRaaFd2_1;
	wire w_dff_B_ROjjjfPG1_1;
	wire w_dff_B_KBNO8qCX6_1;
	wire w_dff_B_eiIrvGNx6_1;
	wire w_dff_B_eKxwp02R0_1;
	wire w_dff_B_j0ZXAfue4_1;
	wire w_dff_B_q4SCnHRo3_1;
	wire w_dff_B_yqUuNiF27_1;
	wire w_dff_B_6gAHwBbU4_1;
	wire w_dff_B_9uRagnYN2_1;
	wire w_dff_B_yvbGykZv8_1;
	wire w_dff_B_Rf84pPBc9_1;
	wire w_dff_B_UaYS03Sm0_1;
	wire w_dff_B_Lv8aYlRS2_1;
	wire w_dff_B_nKxXnrAS9_1;
	wire w_dff_B_RI7p9Pgb4_1;
	wire w_dff_B_MjVwJuex5_1;
	wire w_dff_B_IeQ4Mc0m0_1;
	wire w_dff_B_gagweyfX1_1;
	wire w_dff_B_vImXVMkq9_1;
	wire w_dff_B_Fy0Ny00m6_1;
	wire w_dff_B_m2D6RYDR1_1;
	wire w_dff_B_pkyARCTV1_1;
	wire w_dff_B_wCo3a4uh3_1;
	wire w_dff_B_adX6pACi2_1;
	wire w_dff_B_nmUoOWI66_1;
	wire w_dff_B_SEGCZxaa1_1;
	wire w_dff_B_TSwSvq6g1_1;
	wire w_dff_B_1mC62K1r5_1;
	wire w_dff_B_mJvpMM5J6_1;
	wire w_dff_B_7g41H3jB4_1;
	wire w_dff_B_SMAtpfSw4_1;
	wire w_dff_B_R6hwYzDj5_1;
	wire w_dff_B_3bWrEArN2_1;
	wire w_dff_B_vYwylIjI8_1;
	wire w_dff_B_p6j5WuPh1_1;
	wire w_dff_B_LM4YDIdJ9_1;
	wire w_dff_B_rYnpfGur9_1;
	wire w_dff_B_WjD0aMZd3_1;
	wire w_dff_B_QPjPjBpq5_1;
	wire w_dff_B_aDRMe4PM0_1;
	wire w_dff_B_e4yJMXLs2_1;
	wire w_dff_B_FbGaAzP94_1;
	wire w_dff_B_kRlxDcRM9_1;
	wire w_dff_B_K1GLlw1c3_1;
	wire w_dff_B_tpgJ8gqe1_1;
	wire w_dff_B_Xe6Nxzol9_1;
	wire w_dff_B_Ba2xc9xv1_1;
	wire w_dff_B_9H4eVJqS1_1;
	wire w_dff_B_QxYkCHCB4_1;
	wire w_dff_B_9DOl2dlq1_1;
	wire w_dff_B_TLypH8Ai2_1;
	wire w_dff_B_kCdFSZW74_1;
	wire w_dff_B_7uOlee4C1_1;
	wire w_dff_B_EnuMKhEj9_1;
	wire w_dff_B_s0KFe9fj8_1;
	wire w_dff_B_TVXLodJF2_1;
	wire w_dff_B_KSR3uyc06_1;
	wire w_dff_B_chq6mbe15_1;
	wire w_dff_B_mRhf5AEx1_1;
	wire w_dff_B_WB3M9t5M1_1;
	wire w_dff_B_eVZxnaxN8_1;
	wire w_dff_B_DdqK9DK56_1;
	wire w_dff_B_3fbI7QoG4_1;
	wire w_dff_B_hD5JL3X31_1;
	wire w_dff_B_T0axEqJp4_1;
	wire w_dff_B_1b3jWi2f0_1;
	wire w_dff_B_2WwhoMh78_1;
	wire w_dff_B_wdK9Ir0v9_1;
	wire w_dff_B_y3iiGRBm9_1;
	wire w_dff_B_HdQzN8y37_1;
	wire w_dff_B_cK9Wfv0w3_1;
	wire w_dff_B_3DTy8LOv2_1;
	wire w_dff_B_tLOrQI8M4_1;
	wire w_dff_B_rKWA5vRt1_1;
	wire w_dff_B_o87l8aUU6_1;
	wire w_dff_B_LJrdZcoV6_1;
	wire w_dff_B_3iq7gh183_1;
	wire w_dff_B_eOcfunNn6_1;
	wire w_dff_B_M44iwoup2_1;
	wire w_dff_B_NZWnolkN1_1;
	wire w_dff_B_HRJjBXxx8_1;
	wire w_dff_B_iOqjcP361_1;
	wire w_dff_B_pZsGzh8i1_1;
	wire w_dff_B_HiqvZNM75_1;
	wire w_dff_B_58S1dTmc4_1;
	wire w_dff_B_AIeOHJQc4_1;
	wire w_dff_B_y7GOh2GO1_1;
	wire w_dff_B_1GvLUgkk3_1;
	wire w_dff_B_VKTN7njI5_1;
	wire w_dff_B_ENsKRcJM1_1;
	wire w_dff_B_nLYm0xp18_1;
	wire w_dff_B_nm5uEQUF1_1;
	wire w_dff_B_leim9mt08_1;
	wire w_dff_B_4OcNLf0j8_1;
	wire w_dff_B_yT9SxfeR2_1;
	wire w_dff_B_Gpk7ezK60_1;
	wire w_dff_B_GV3mzXQq6_1;
	wire w_dff_B_eRvdZ90j5_1;
	wire w_dff_B_FaZyKaHO6_1;
	wire w_dff_B_Q1e6kKlY1_1;
	wire w_dff_B_HjgawN2L4_1;
	wire w_dff_B_Fwoz4kiq8_1;
	wire w_dff_B_m5fpVlLg8_1;
	wire w_dff_B_vzpSX2mR4_1;
	wire w_dff_B_GWrfhdjj7_1;
	wire w_dff_B_azPfQlIz8_1;
	wire w_dff_B_RojonLnm3_1;
	wire w_dff_B_0svLXzdR2_1;
	wire w_dff_B_6HtfvSOS6_1;
	wire w_dff_B_4X46y0Zx8_1;
	wire w_dff_B_9XwRkT5m5_1;
	wire w_dff_B_JDgGXXA50_1;
	wire w_dff_B_bJFpnRci9_1;
	wire w_dff_B_XbohPpsD3_1;
	wire w_dff_B_N8lpKHza2_1;
	wire w_dff_B_dvW6l90d8_1;
	wire w_dff_B_d6sjpxFq3_1;
	wire w_dff_B_gdriOl6g3_1;
	wire w_dff_B_fo7zCS5x4_1;
	wire w_dff_B_7bwNHSSY3_1;
	wire w_dff_B_hrismID71_1;
	wire w_dff_B_XrvHtSpy0_1;
	wire w_dff_B_qP46jQbq7_1;
	wire w_dff_B_Lp0w4pKz5_1;
	wire w_dff_B_JaaTS2r72_1;
	wire w_dff_B_xVwlfayq0_1;
	wire w_dff_B_FPu8Wwva5_1;
	wire w_dff_B_1oXggIs45_1;
	wire w_dff_B_KPVkZZ1V2_1;
	wire w_dff_B_WDY1Kifv8_1;
	wire w_dff_B_7kyrPZGY8_1;
	wire w_dff_B_lFBVzJRX8_1;
	wire w_dff_B_j0VSIXt63_1;
	wire w_dff_B_xPBzHC7Q5_1;
	wire w_dff_B_hONsmt908_1;
	wire w_dff_B_FVWJcb5u2_1;
	wire w_dff_B_3SjG0wVu9_1;
	wire w_dff_B_A1I68soy3_1;
	wire w_dff_B_8JRnPKiX5_1;
	wire w_dff_B_tDYKRwZI0_1;
	wire w_dff_B_hBPbpSF41_1;
	wire w_dff_B_kihbHujo9_1;
	wire w_dff_B_G1s9zMRU0_1;
	wire w_dff_B_hcVLaKD18_1;
	wire w_dff_B_tril6glz3_1;
	wire w_dff_B_f9GTB9Qv4_1;
	wire w_dff_B_5nRltPhm2_1;
	wire w_dff_B_TTlbWxqY0_1;
	wire w_dff_B_6A8co7Y52_1;
	wire w_dff_B_CrUABUte0_1;
	wire w_dff_B_r7vsu1Nx8_1;
	wire w_dff_B_1VqjD5nW2_1;
	wire w_dff_B_J5Fk6Dix5_1;
	wire w_dff_B_IIvwCoP80_1;
	wire w_dff_B_hnLLpKD29_1;
	wire w_dff_B_n8LY6GXK0_1;
	wire w_dff_B_VqgwCVqI3_1;
	wire w_dff_B_5l941F006_1;
	wire w_dff_B_ukXY0LS96_1;
	wire w_dff_B_DvN4zRQK4_1;
	wire w_dff_B_bNcWidkD1_1;
	wire w_dff_B_e8CpMAeq7_1;
	wire w_dff_B_GLpHVpJ71_1;
	wire w_dff_B_w224alA12_1;
	wire w_dff_B_lX1idXQ92_1;
	wire w_dff_B_X10zzGzj2_1;
	wire w_dff_B_omWaHplO9_1;
	wire w_dff_B_Y6maJJWP2_1;
	wire w_dff_B_LMy4L1Qn7_1;
	wire w_dff_B_ls9Yo28U4_1;
	wire w_dff_B_vrSgv7pe0_1;
	wire w_dff_B_Z4eQIBYN1_1;
	wire w_dff_B_uZtKOEGq0_1;
	wire w_dff_B_xiNNoxFZ7_1;
	wire w_dff_B_w2Kbh6uf6_1;
	wire w_dff_B_fP7WTlcY5_1;
	wire w_dff_B_lQr3XVAK2_0;
	wire w_dff_B_jaXDnHrE5_1;
	wire w_dff_B_9wBv86Ac4_1;
	wire w_dff_B_fvAVpMFh9_1;
	wire w_dff_B_vJGQTYef9_1;
	wire w_dff_B_tkLLvKi47_1;
	wire w_dff_B_u5sNaIjK6_1;
	wire w_dff_B_nPcle7br3_1;
	wire w_dff_B_yBkNdTAm7_1;
	wire w_dff_B_aBIokkte6_1;
	wire w_dff_B_tCAIVqgo6_1;
	wire w_dff_B_kiUSm16c5_1;
	wire w_dff_B_HxyBNYEG0_1;
	wire w_dff_B_dZMtG6911_1;
	wire w_dff_B_hzE7q2Sk5_0;
	wire w_dff_B_M75Ir0bP4_0;
	wire w_dff_B_uR6tgjXS1_0;
	wire w_dff_B_o6DSENKN7_0;
	wire w_dff_B_1VrmdnFO5_0;
	wire w_dff_B_wBAEPCUH7_0;
	wire w_dff_B_XMCAzU8D6_0;
	wire w_dff_B_TvpWawKz1_0;
	wire w_dff_B_wkIjs8mN0_0;
	wire w_dff_B_xwv9vb1o5_0;
	wire w_dff_B_r6oV5yp74_0;
	wire w_dff_B_rGI5WH8Q5_1;
	wire w_dff_B_KOkLL7AE8_1;
	wire w_dff_B_ePLJXcwg3_1;
	wire w_dff_B_hUuTLsCD0_1;
	wire w_dff_B_S0A38z4p1_1;
	wire w_dff_B_EGWBvchY7_1;
	wire w_dff_B_xNPsICqc2_1;
	wire w_dff_B_ATuq1jgw3_1;
	wire w_dff_B_9yHiEcDe7_1;
	wire w_dff_B_AIQlOzkn9_1;
	wire w_dff_B_qcB4i5Lp4_1;
	wire w_dff_B_iWYRQ4ys9_0;
	wire w_dff_B_9V90CMJQ5_0;
	wire w_dff_B_ILgibT5O4_0;
	wire w_dff_B_j6mQpogF4_0;
	wire w_dff_B_M99bmLne9_0;
	wire w_dff_B_0JsVgMXC5_0;
	wire w_dff_B_qXfIvdzc3_0;
	wire w_dff_B_vlFBUAih6_0;
	wire w_dff_B_Fso2apb72_0;
	wire w_dff_B_Mr2wOWV55_0;
	wire w_dff_B_EnAgxTet0_1;
	wire w_dff_B_7uuecxy63_1;
	wire w_dff_B_Nve3TPCf6_1;
	wire w_dff_B_dVl77WSQ0_1;
	wire w_dff_B_UgyF34N34_1;
	wire w_dff_B_vuOcyOYu8_1;
	wire w_dff_B_dW6bcvXe1_1;
	wire w_dff_B_fFrwz9Kn1_1;
	wire w_dff_B_3aU9GhEG7_1;
	wire w_dff_B_oepmN3JF2_1;
	wire w_dff_B_j2KrgK254_1;
	wire w_dff_B_dA0HCEG48_0;
	wire w_dff_B_FrlL5QKw2_0;
	wire w_dff_B_IJ6pwduu0_0;
	wire w_dff_B_T53wAaOn3_0;
	wire w_dff_B_tdxjmLkO7_0;
	wire w_dff_B_SkyAzguN9_0;
	wire w_dff_B_LpsxhZDt1_0;
	wire w_dff_B_GuIOCIJb2_0;
	wire w_dff_B_KkbU6eaE5_0;
	wire w_dff_B_S11eF9xM5_0;
	wire w_dff_B_wMnVA5vf0_1;
	wire w_dff_B_YRmfgDlQ7_1;
	wire w_dff_B_pqd1WIft9_1;
	wire w_dff_B_kiTDo6Kq4_1;
	wire w_dff_B_YX0j1f3L9_1;
	wire w_dff_B_29pD1IvM8_1;
	wire w_dff_B_3g9DAuUi8_1;
	wire w_dff_B_U9vd2RPF0_1;
	wire w_dff_B_CVMHTWgo6_1;
	wire w_dff_B_ZL5KMlUy4_1;
	wire w_dff_B_IOofLOGl5_1;
	wire w_dff_B_jd8bIYSw8_0;
	wire w_dff_B_KPUmYetE3_0;
	wire w_dff_B_VMl6ZMXJ6_0;
	wire w_dff_B_fqJm61u26_0;
	wire w_dff_B_V9aPycDz6_0;
	wire w_dff_B_I7mBGZew2_0;
	wire w_dff_B_OEd8LnQS6_0;
	wire w_dff_B_ss3azBuR8_0;
	wire w_dff_B_bZAGdl4l4_0;
	wire w_dff_B_BE1ml2kz8_0;
	wire w_dff_B_hYszWuVb0_1;
	wire w_dff_B_e55ES3g08_1;
	wire w_dff_B_qY7AI4fe1_1;
	wire w_dff_B_YByykTAO4_1;
	wire w_dff_B_pOUOZQxt6_1;
	wire w_dff_B_pWBfprob9_1;
	wire w_dff_B_dJN2MV1C9_1;
	wire w_dff_B_VGF49Dzw2_1;
	wire w_dff_B_aAjyqMuW4_1;
	wire w_dff_B_C10XhRCQ3_1;
	wire w_dff_B_kjNYoeB98_1;
	wire w_dff_B_I9vmdZhI1_0;
	wire w_dff_B_9Thgu8DF7_0;
	wire w_dff_B_qODYfE2y9_0;
	wire w_dff_B_9f9ANNgz1_0;
	wire w_dff_B_AYakFLww5_0;
	wire w_dff_B_eCcqk5O08_0;
	wire w_dff_B_grq4Gk7X6_0;
	wire w_dff_B_XJeiFyyT6_0;
	wire w_dff_B_V3IDgEqV0_0;
	wire w_dff_B_EOQdpHEL7_0;
	wire w_dff_B_lnKr4Z7M8_1;
	wire w_dff_B_8ryk7nNh3_1;
	wire w_dff_B_xT2rPhOl3_1;
	wire w_dff_B_cyBPuupf1_1;
	wire w_dff_B_RtfzpUNm3_1;
	wire w_dff_B_5IUnnD3o3_1;
	wire w_dff_B_cInorMwj2_1;
	wire w_dff_B_xnrt3JKO3_1;
	wire w_dff_B_566lHE4j0_1;
	wire w_dff_B_Rt7hsOhw1_1;
	wire w_dff_B_E0Q23Cbc3_1;
	wire w_dff_B_Te4K5kvL8_0;
	wire w_dff_B_HrG0XZDw7_0;
	wire w_dff_B_5V2AectB7_0;
	wire w_dff_B_vyjlDjqI7_0;
	wire w_dff_B_37Ud5FH85_0;
	wire w_dff_B_2VjCm8n39_0;
	wire w_dff_B_Xsyp27mk8_0;
	wire w_dff_B_9EHMQM611_0;
	wire w_dff_B_JgvJPJc61_0;
	wire w_dff_B_UVLAc0EO0_1;
	wire w_dff_B_ldjYnZOI1_1;
	wire w_dff_B_8qoqtQM48_1;
	wire w_dff_B_a3dab27L0_1;
	wire w_dff_B_zJk2ODOZ0_1;
	wire w_dff_B_gh0oauVX4_1;
	wire w_dff_B_Zy8hjRZX6_1;
	wire w_dff_B_yrkT1iFw0_1;
	wire w_dff_B_recaVOal6_1;
	wire w_dff_B_mdApH64o0_1;
	wire w_dff_B_ZACUQHss7_0;
	wire w_dff_B_b66iRCz56_0;
	wire w_dff_B_C0krQAGI3_0;
	wire w_dff_B_lZH28Lpf5_0;
	wire w_dff_B_0PpXJGId1_0;
	wire w_dff_B_I3gLJUfE5_0;
	wire w_dff_B_lJpb3XBs9_0;
	wire w_dff_B_L0Rmnoh95_0;
	wire w_dff_B_NtB9GY9u5_1;
	wire w_dff_B_kc2SXV4C9_1;
	wire w_dff_B_lIn9U0oC5_1;
	wire w_dff_B_vMqNVLf12_1;
	wire w_dff_B_eK3ZCjBO5_1;
	wire w_dff_B_ZLlHNbcU6_1;
	wire w_dff_B_4HoTxXe18_1;
	wire w_dff_B_vK72Semg3_1;
	wire w_dff_B_hSZeGp3d4_1;
	wire w_dff_B_mlg2U20o0_1;
	wire w_dff_B_lK74pQE89_0;
	wire w_dff_B_M2oIsJN86_0;
	wire w_dff_B_qero6xuu1_0;
	wire w_dff_B_9ZpKI2PX1_0;
	wire w_dff_B_nH3r2rMY5_0;
	wire w_dff_B_eMl8xzca9_0;
	wire w_dff_B_C1LZVcf42_0;
	wire w_dff_B_KPH1H2a54_0;
	wire w_dff_B_SkgusjyV0_1;
	wire w_dff_B_xg0A5I4d9_1;
	wire w_dff_B_5i3qlVWW0_1;
	wire w_dff_B_B4WHnUco5_1;
	wire w_dff_B_ealkyqLW8_1;
	wire w_dff_B_RwCo48J74_1;
	wire w_dff_B_Gby1XeE97_1;
	wire w_dff_B_ykjfpplL7_1;
	wire w_dff_B_PRkjS5AF3_0;
	wire w_dff_B_zJBKnvHv2_0;
	wire w_dff_B_ORoFsjNZ9_0;
	wire w_dff_B_dN8MtqrG4_0;
	wire w_dff_B_mMBcqcDb9_0;
	wire w_dff_B_GiR5nEIQ5_0;
	wire w_dff_B_nptbMNFz7_1;
	wire w_dff_B_ybqZzHbw3_1;
	wire w_dff_B_lyZevIjg9_1;
	wire w_dff_B_0dddYj4P1_1;
	wire w_dff_B_vvQWjoHL8_1;
	wire w_dff_B_FY27eXD76_1;
	wire w_dff_B_nLY9nNaa0_1;
	wire w_dff_B_4sthuPwJ9_0;
	wire w_dff_B_00MQZg730_0;
	wire w_dff_B_RFCXNyKI4_0;
	wire w_dff_B_ur5vXtRu1_0;
	wire w_dff_B_6uiefIB11_0;
	wire w_dff_B_I9SQWbCD5_1;
	wire w_dff_B_71iVHwuC6_1;
	wire w_dff_B_SUufHxY01_1;
	wire w_dff_B_tkTdiyXq4_1;
	wire w_dff_B_1GNZutHk9_1;
	wire w_dff_B_lqat5rQz4_1;
	wire w_dff_B_TqqQ4Yxt6_0;
	wire w_dff_B_JkGMiJWi8_0;
	wire w_dff_B_3E5T5ux09_0;
	wire w_dff_B_FsUF8c9E3_0;
	wire w_dff_B_NR9urmj73_1;
	wire w_dff_B_vpyJeysS8_1;
	wire w_dff_B_AURzPvBv7_1;
	wire w_dff_B_nG2AdicV6_1;
	wire w_dff_B_avGxlZft2_1;
	wire w_dff_A_7UVDgp5P2_1;
	wire w_dff_B_wDX4iwEr7_2;
	wire w_dff_B_39iS0oOH0_1;
	wire w_dff_B_Vw5ca9Im3_1;
	wire w_dff_B_2un0XYhY5_1;
	wire w_dff_B_PH0q2cYe9_1;
	wire w_dff_B_oci1c3qe0_1;
	wire w_dff_B_GX6DC5BQ6_1;
	wire w_dff_B_APQpbtXG4_1;
	wire w_dff_B_mzf3UAuW1_1;
	wire w_dff_B_44uZDAnU6_1;
	wire w_dff_B_JW3HweTE7_1;
	wire w_dff_B_rPUbm3kx1_1;
	wire w_dff_B_Qkzi8O9h3_1;
	wire w_dff_B_pS4HvURR3_1;
	wire w_dff_B_hckTMUBH6_1;
	wire w_dff_B_MoKKPG2t4_0;
	wire w_dff_A_DmL1QnrY4_0;
	wire w_dff_A_er5FX7J50_0;
	wire w_dff_A_bTCAl6WQ9_1;
	wire w_dff_A_0ScrAvYA0_0;
	wire w_dff_A_qLQNHc772_0;
	wire w_dff_A_sQAbRgXs7_0;
	wire w_dff_A_vSrC9zRj6_0;
	wire w_dff_A_TpQrlgLG0_0;
	wire w_dff_A_gMDywc4O0_0;
	wire w_dff_A_tBK1z3xF2_0;
	wire w_dff_A_uUoxld6q6_0;
	wire w_dff_A_TSALyH9y1_0;
	wire w_dff_A_8ps0W6gc6_0;
	wire w_dff_A_SfDcYrZF8_0;
	wire w_dff_A_r7UZrAKR5_0;
	wire w_dff_A_5wePWLCf3_0;
	wire w_dff_A_c6DtyH4Z5_0;
	wire w_dff_A_yUtL0ibs1_0;
	wire w_dff_A_w9w5rUgd2_0;
	wire w_dff_A_k6MJjzzb4_0;
	wire w_dff_A_oFhV9Yys2_0;
	wire w_dff_A_JySU2AdA9_0;
	wire w_dff_A_KL1R5lLa0_0;
	wire w_dff_A_QlsXtofC7_0;
	wire w_dff_A_Ml9p01M16_0;
	wire w_dff_A_hgOBoV5l6_0;
	wire w_dff_A_wZoIVWxZ6_0;
	wire w_dff_A_Hus5icBz9_0;
	wire w_dff_A_b67jr6Eg0_0;
	wire w_dff_A_ykMKu8d73_0;
	wire w_dff_A_V9d7Aimv6_0;
	wire w_dff_A_7JUV1yZB5_0;
	wire w_dff_A_LULJGEXV8_0;
	wire w_dff_A_uLmT33eu7_0;
	wire w_dff_A_CDSpkiVt9_0;
	wire w_dff_A_czkmhjny3_0;
	wire w_dff_A_k853RhGH4_0;
	wire w_dff_A_aj8YeYcW4_0;
	wire w_dff_A_Nfl5jsIK7_0;
	wire w_dff_A_9TjwUSOj3_0;
	wire w_dff_A_WJ4WcMJ96_0;
	wire w_dff_A_eAcLipFN6_0;
	wire w_dff_A_CjbjKJoK4_0;
	wire w_dff_A_xsCKGOOr4_0;
	wire w_dff_A_kfiwen4i4_0;
	wire w_dff_A_EhPrHA807_0;
	wire w_dff_A_PStkDCsD2_0;
	wire w_dff_A_PqZ9lHp65_0;
	wire w_dff_A_N5TV2sMd6_0;
	wire w_dff_A_1HmaeqVb3_0;
	wire w_dff_A_yHb2qhDd5_0;
	wire w_dff_A_SRkecX2R9_0;
	wire w_dff_A_TMtIDAje4_0;
	wire w_dff_A_hsT0ClWq5_0;
	wire w_dff_A_jvqCnlvm2_0;
	wire w_dff_A_KLP8Ccrj8_0;
	wire w_dff_A_HMvn4lKJ5_0;
	wire w_dff_A_g1u098Kg4_0;
	wire w_dff_A_qD6Vc4tY9_0;
	wire w_dff_A_nwd66FEe1_0;
	wire w_dff_A_djA9kIsB9_0;
	wire w_dff_A_cVpNKl5A7_0;
	wire w_dff_A_JccXoHeQ7_0;
	wire w_dff_A_UdverVv39_0;
	wire w_dff_A_d1Vwirj30_0;
	wire w_dff_A_3DOedldN8_0;
	wire w_dff_A_aVw6sbrF0_0;
	wire w_dff_A_7PPz50Jf7_0;
	wire w_dff_A_bjUMuoak4_0;
	wire w_dff_A_5CgO0BtO3_0;
	wire w_dff_A_4BrFiUsN2_0;
	wire w_dff_A_YHZsrDRc7_0;
	wire w_dff_A_CFwdSuc96_0;
	wire w_dff_A_mKQsCMmW1_0;
	wire w_dff_A_CaANVt3b2_0;
	wire w_dff_A_i7WgIhzW9_0;
	wire w_dff_A_Ylhs6zuk8_0;
	wire w_dff_A_PCFOBIdG2_2;
	wire w_dff_A_2Mzr1ECC3_0;
	wire w_dff_A_6QKawOoD4_0;
	wire w_dff_A_qtsaskvR9_0;
	wire w_dff_A_Sfvt9r7P4_0;
	wire w_dff_A_q7zQL3ts8_0;
	wire w_dff_A_fIX6F0zj0_0;
	wire w_dff_A_vYgo1J5r7_0;
	wire w_dff_A_kruFvQBM7_0;
	wire w_dff_A_IV5qeMYJ4_0;
	wire w_dff_A_HfrdipqK3_0;
	wire w_dff_A_KzklCMRf5_0;
	wire w_dff_A_TOlj5WV82_0;
	wire w_dff_A_20sgbXbq4_0;
	wire w_dff_A_TcYi2j4C9_0;
	wire w_dff_A_AANIZtXG9_0;
	wire w_dff_A_0MjJmIVK0_0;
	wire w_dff_A_o8qRoWCs1_0;
	wire w_dff_A_xRSwZSJU0_0;
	wire w_dff_A_fuC9qxw03_0;
	wire w_dff_A_yOpVah1B5_0;
	wire w_dff_A_L9WocArF1_0;
	wire w_dff_A_40Vxe5di2_0;
	wire w_dff_A_W9DxnpiI7_0;
	wire w_dff_A_YHCbXd5w3_0;
	wire w_dff_A_Re9knHc57_0;
	wire w_dff_A_XOXyhfpa9_0;
	wire w_dff_A_LsnChDDU8_0;
	wire w_dff_A_ZmF08uMv9_0;
	wire w_dff_A_bYxj8sBs4_0;
	wire w_dff_A_iiqDTF3D9_0;
	wire w_dff_A_K79vuuDa3_0;
	wire w_dff_A_f7m85JD31_0;
	wire w_dff_A_BbEZIhoi3_0;
	wire w_dff_A_BfSG9JWu2_0;
	wire w_dff_A_sC9H0qdR7_0;
	wire w_dff_A_GnSGWHR24_0;
	wire w_dff_A_9uD8Bf8N0_0;
	wire w_dff_A_z35CjSuA4_0;
	wire w_dff_A_PBj5hJAw0_0;
	wire w_dff_A_BhJGv6NN6_0;
	wire w_dff_A_p09tgYgj6_0;
	wire w_dff_A_79XkmjZf6_0;
	wire w_dff_A_fInH4XCV8_0;
	wire w_dff_A_SHtWT2Ly0_0;
	wire w_dff_A_KT4lCMgo8_0;
	wire w_dff_A_dWzDn9il4_0;
	wire w_dff_A_cUp3s2dx7_0;
	wire w_dff_A_xij6pl4g4_0;
	wire w_dff_A_TqnhkYWe8_0;
	wire w_dff_A_4k5xBdMV0_0;
	wire w_dff_A_WkaFB5Xi3_0;
	wire w_dff_A_aMyXT85o1_0;
	wire w_dff_A_kEIejvSk1_0;
	wire w_dff_A_pmcdxPhG1_0;
	wire w_dff_A_spjh1imy7_0;
	wire w_dff_A_5Otg00Ik3_0;
	wire w_dff_A_tezjCjUI0_0;
	wire w_dff_A_urczoHXB2_0;
	wire w_dff_A_MXXMO5ot8_0;
	wire w_dff_A_uGgSWvGW4_0;
	wire w_dff_A_M4EEyhLj5_0;
	wire w_dff_A_BoXyyHj22_0;
	wire w_dff_A_KXOUefs93_0;
	wire w_dff_A_9WUW8n335_0;
	wire w_dff_A_A8KvOhOl2_0;
	wire w_dff_A_7h32TuHA1_0;
	wire w_dff_A_ZHltzi1X1_0;
	wire w_dff_A_3wjTuG9P9_0;
	wire w_dff_A_xfIO8r2W7_0;
	wire w_dff_A_a0upQTJm5_0;
	wire w_dff_A_yRiCeCrV9_0;
	wire w_dff_A_gydU51Oe5_2;
	wire w_dff_A_f0BGSe2f5_0;
	wire w_dff_A_Z82EQlDJ0_0;
	wire w_dff_A_8FEFZ3Sz6_0;
	wire w_dff_A_YKmMqeaU2_0;
	wire w_dff_A_Nlbuindq6_0;
	wire w_dff_A_aooHxRTH7_0;
	wire w_dff_A_02m7LUoB2_0;
	wire w_dff_A_Ey6ruAB05_0;
	wire w_dff_A_y3NXqFwT3_0;
	wire w_dff_A_NKMh9XOT2_0;
	wire w_dff_A_sODMZWVr2_0;
	wire w_dff_A_EmYJyEwV8_0;
	wire w_dff_A_jpwXQkDx7_0;
	wire w_dff_A_e7PbWgvi1_0;
	wire w_dff_A_CmrDmMdF6_0;
	wire w_dff_A_fYsxbyRn4_0;
	wire w_dff_A_kJxXDTez0_0;
	wire w_dff_A_2msFmwVe4_0;
	wire w_dff_A_Y1vpadBU8_0;
	wire w_dff_A_IR9ELOl26_0;
	wire w_dff_A_LbQzRoPG2_0;
	wire w_dff_A_PbrkiFNE5_0;
	wire w_dff_A_PsTxWtSE7_0;
	wire w_dff_A_o7jEZkWX4_0;
	wire w_dff_A_7t3XfWNz9_0;
	wire w_dff_A_XgoMQO123_0;
	wire w_dff_A_wG1z2PhT4_0;
	wire w_dff_A_QuhbicoL8_0;
	wire w_dff_A_pYRUjwUH3_0;
	wire w_dff_A_6lbBUaA12_0;
	wire w_dff_A_02XnWht50_0;
	wire w_dff_A_yZOGwDdy5_0;
	wire w_dff_A_fXIKyH653_0;
	wire w_dff_A_cfc6UD1e7_0;
	wire w_dff_A_NMSQm9MR7_0;
	wire w_dff_A_5u7OaqjL0_0;
	wire w_dff_A_kK3LOHlJ4_0;
	wire w_dff_A_4rjhZXYO1_0;
	wire w_dff_A_PrmI54Ub1_0;
	wire w_dff_A_IUVx0WOO6_0;
	wire w_dff_A_x7acFD1t4_0;
	wire w_dff_A_EXnmhxjQ7_0;
	wire w_dff_A_SV20HDXb9_0;
	wire w_dff_A_S1NUcAYo4_0;
	wire w_dff_A_KjQWqlTc9_0;
	wire w_dff_A_W7rxWAuA6_0;
	wire w_dff_A_gGrn6bqt5_0;
	wire w_dff_A_tvdmtwT72_0;
	wire w_dff_A_g3iGdPqK3_0;
	wire w_dff_A_nb6Nw2eq1_0;
	wire w_dff_A_KDkDbngu1_0;
	wire w_dff_A_halcnJiQ9_0;
	wire w_dff_A_8uHcXYeR0_0;
	wire w_dff_A_gC3Qiwfd9_0;
	wire w_dff_A_o0s4HBiH8_0;
	wire w_dff_A_npWGeNy41_0;
	wire w_dff_A_7cSNeZNJ3_0;
	wire w_dff_A_MEfw7ESU9_0;
	wire w_dff_A_Aj5JIvaH9_0;
	wire w_dff_A_DcTs0AJE7_0;
	wire w_dff_A_xyrkQMju2_0;
	wire w_dff_A_VhTIUq7m4_0;
	wire w_dff_A_tmLdcmJc5_0;
	wire w_dff_A_XJUDcSpe1_0;
	wire w_dff_A_q39y2On41_0;
	wire w_dff_A_lOleXO5M1_0;
	wire w_dff_A_jGqRSgYq8_0;
	wire w_dff_A_1EyJbabK4_0;
	wire w_dff_A_prb6lJFG0_2;
	wire w_dff_A_OxDidKSP6_0;
	wire w_dff_A_nhZic5li8_0;
	wire w_dff_A_qVQCv1YV5_0;
	wire w_dff_A_uOX3vY8y9_0;
	wire w_dff_A_jiOCJq2f3_0;
	wire w_dff_A_GViBomQK2_0;
	wire w_dff_A_BPR3l0ig8_0;
	wire w_dff_A_BVTRRFdk0_0;
	wire w_dff_A_sHcPSkRH4_0;
	wire w_dff_A_BaoC3HYn5_0;
	wire w_dff_A_vtT2dp4p0_0;
	wire w_dff_A_v1QtNPQd3_0;
	wire w_dff_A_N14FrFCB5_0;
	wire w_dff_A_tDFYfXtJ0_0;
	wire w_dff_A_NWvUz3em2_0;
	wire w_dff_A_xgo9767D0_0;
	wire w_dff_A_1dlcXUkU6_0;
	wire w_dff_A_tK44xAL30_0;
	wire w_dff_A_XSa6KXDS5_0;
	wire w_dff_A_i5QkZB390_0;
	wire w_dff_A_KRykysKq3_0;
	wire w_dff_A_dJJBCedG5_0;
	wire w_dff_A_gKHGj8eP3_0;
	wire w_dff_A_EN3SHpej0_0;
	wire w_dff_A_visgnOOx6_0;
	wire w_dff_A_BaUCnUCu8_0;
	wire w_dff_A_868bPX6R5_0;
	wire w_dff_A_djX1Utye9_0;
	wire w_dff_A_L5yEuaN89_0;
	wire w_dff_A_FtbR5yr94_0;
	wire w_dff_A_7OJ4VoAa6_0;
	wire w_dff_A_fgphuv9K2_0;
	wire w_dff_A_98YRb6NB4_0;
	wire w_dff_A_Nd46zg6l7_0;
	wire w_dff_A_8ZNJjnBP0_0;
	wire w_dff_A_smKaSlsP2_0;
	wire w_dff_A_xGrdbFud0_0;
	wire w_dff_A_qInHphzq1_0;
	wire w_dff_A_O9y1Lb8v6_0;
	wire w_dff_A_VhWduckN3_0;
	wire w_dff_A_xsRKr0yu5_0;
	wire w_dff_A_40cJkeo17_0;
	wire w_dff_A_18VOsNQB2_0;
	wire w_dff_A_9sdn0RMT2_0;
	wire w_dff_A_98yKo7043_0;
	wire w_dff_A_uhu3chIJ6_0;
	wire w_dff_A_W66ZXEkR4_0;
	wire w_dff_A_Z4KDpIEW7_0;
	wire w_dff_A_RbhZD9fC4_0;
	wire w_dff_A_W8eiWEpY2_0;
	wire w_dff_A_fh2Rwq3V3_0;
	wire w_dff_A_dX8P4xxg6_0;
	wire w_dff_A_7fRx0Mrl3_0;
	wire w_dff_A_auYM8PUv0_0;
	wire w_dff_A_hLHArS1K8_0;
	wire w_dff_A_qWyZckTx6_0;
	wire w_dff_A_TXm0458n1_0;
	wire w_dff_A_o8ZbXhrK7_0;
	wire w_dff_A_ycn3xqJR2_0;
	wire w_dff_A_Ljgp1K857_0;
	wire w_dff_A_WVhfadmC6_0;
	wire w_dff_A_YMi4KCxM8_0;
	wire w_dff_A_B2GAhc2t0_0;
	wire w_dff_A_KptnlIbk0_0;
	wire w_dff_A_usnr3rUr2_0;
	wire w_dff_A_wOXl4S3M1_2;
	wire w_dff_A_7hy5QJns0_0;
	wire w_dff_A_9hqhv14t9_0;
	wire w_dff_A_Eg2t6DAC9_0;
	wire w_dff_A_Ucnyg9uT8_0;
	wire w_dff_A_HFgQc5mW3_0;
	wire w_dff_A_m2Fx4NjN1_0;
	wire w_dff_A_cNwbseb57_0;
	wire w_dff_A_8434XY279_0;
	wire w_dff_A_JxH1Zs8H1_0;
	wire w_dff_A_J77lj9Wa2_0;
	wire w_dff_A_TxcUI6uj4_0;
	wire w_dff_A_EwTEVRUW8_0;
	wire w_dff_A_0EUdAcGq7_0;
	wire w_dff_A_trISoiH85_0;
	wire w_dff_A_GSLkOisb4_0;
	wire w_dff_A_6xvPxCsa1_0;
	wire w_dff_A_1uvFQFdB0_0;
	wire w_dff_A_bcgkZdub8_0;
	wire w_dff_A_XauOiins2_0;
	wire w_dff_A_vABrxvFW2_0;
	wire w_dff_A_NpsOMvbQ7_0;
	wire w_dff_A_7ONuRJUz4_0;
	wire w_dff_A_qnQvu6wG7_0;
	wire w_dff_A_yHLzZtqQ6_0;
	wire w_dff_A_S3XagoCB4_0;
	wire w_dff_A_qJZC3b2K1_0;
	wire w_dff_A_h7xJIght0_0;
	wire w_dff_A_pA7sS7h18_0;
	wire w_dff_A_uPneUDtG5_0;
	wire w_dff_A_pGczmvaZ8_0;
	wire w_dff_A_mQKarlVz4_0;
	wire w_dff_A_2ghvIAro6_0;
	wire w_dff_A_pEinz4bu7_0;
	wire w_dff_A_kIk9LCbv3_0;
	wire w_dff_A_UE3MjOxz0_0;
	wire w_dff_A_zyUsQLb01_0;
	wire w_dff_A_ZInLNyof0_0;
	wire w_dff_A_xXkyusC57_0;
	wire w_dff_A_jCgXjnTd6_0;
	wire w_dff_A_Zz3Cu5Ob4_0;
	wire w_dff_A_hTm1wQGb2_0;
	wire w_dff_A_3tHjbWCs9_0;
	wire w_dff_A_SNvfIzRR2_0;
	wire w_dff_A_FCM4mrq16_0;
	wire w_dff_A_YKJtArdH0_0;
	wire w_dff_A_CeUtBCTm7_0;
	wire w_dff_A_8KD9NmQT3_0;
	wire w_dff_A_Mbfv8Efu0_0;
	wire w_dff_A_OjDTsPix5_0;
	wire w_dff_A_sbFXTfGl4_0;
	wire w_dff_A_kJXpJdIh5_0;
	wire w_dff_A_7nFt87XP2_0;
	wire w_dff_A_hhzOfGZQ0_0;
	wire w_dff_A_uQ4sCpKG5_0;
	wire w_dff_A_nnY1DhGg0_0;
	wire w_dff_A_40tFfYE27_0;
	wire w_dff_A_rLL3qYXL8_0;
	wire w_dff_A_y6YoDGeR0_0;
	wire w_dff_A_Xi7DDEN93_0;
	wire w_dff_A_FS9LwAhT9_0;
	wire w_dff_A_DWaR64Ip1_0;
	wire w_dff_A_ZLjqwxAp1_0;
	wire w_dff_A_SMosFExk3_2;
	wire w_dff_A_2rCC6sEb4_0;
	wire w_dff_A_vqOlRl3Q0_0;
	wire w_dff_A_UJhNnV2O6_0;
	wire w_dff_A_Mr6dVPRD9_0;
	wire w_dff_A_2ayOVf0n1_0;
	wire w_dff_A_wPTN0wP55_0;
	wire w_dff_A_ACi7K8od9_0;
	wire w_dff_A_44a2eiLU9_0;
	wire w_dff_A_23gJRQ5g7_0;
	wire w_dff_A_EhztXqOr7_0;
	wire w_dff_A_ihWLOVIY5_0;
	wire w_dff_A_eld0vHKq7_0;
	wire w_dff_A_et9QRQjx2_0;
	wire w_dff_A_bq4bkuOx6_0;
	wire w_dff_A_uAHb1l8Y4_0;
	wire w_dff_A_xT3nxTPf5_0;
	wire w_dff_A_7CDVaAUy7_0;
	wire w_dff_A_osUikJmw5_0;
	wire w_dff_A_I2bKiwRX6_0;
	wire w_dff_A_X3JIcfeP8_0;
	wire w_dff_A_yXilKSbz2_0;
	wire w_dff_A_7BArrZLc7_0;
	wire w_dff_A_k9e5vIjO4_0;
	wire w_dff_A_KPYifWeK0_0;
	wire w_dff_A_gI5v4pFM6_0;
	wire w_dff_A_NR8ptgg72_0;
	wire w_dff_A_gh4Usdza2_0;
	wire w_dff_A_Y3nZJsFV5_0;
	wire w_dff_A_uAOadEvp4_0;
	wire w_dff_A_K3I5LBL13_0;
	wire w_dff_A_cnLgQGrX1_0;
	wire w_dff_A_Lb5zGbly4_0;
	wire w_dff_A_iqgWX9BT3_0;
	wire w_dff_A_jzmE2qCb1_0;
	wire w_dff_A_sq9MCJmi6_0;
	wire w_dff_A_pT415re51_0;
	wire w_dff_A_5iaHRD7b2_0;
	wire w_dff_A_38zF5tBq1_0;
	wire w_dff_A_2sRk0kPJ0_0;
	wire w_dff_A_ltnelA0H8_0;
	wire w_dff_A_7Pslk3Ky0_0;
	wire w_dff_A_C910CYpl6_0;
	wire w_dff_A_3zgdTU2Q9_0;
	wire w_dff_A_er3PfDBR0_0;
	wire w_dff_A_skDCO7qN4_0;
	wire w_dff_A_YhshNMAx9_0;
	wire w_dff_A_NPpsaEtJ7_0;
	wire w_dff_A_jo3nTC6z3_0;
	wire w_dff_A_sl9S4LCA8_0;
	wire w_dff_A_0z457G1N3_0;
	wire w_dff_A_MLvBmDwZ0_0;
	wire w_dff_A_eESDDvKH1_0;
	wire w_dff_A_lYy1cg6K2_0;
	wire w_dff_A_GndAPpUj6_0;
	wire w_dff_A_O1F8qIlQ6_0;
	wire w_dff_A_elzVeDOa0_0;
	wire w_dff_A_BWlKDNSe1_0;
	wire w_dff_A_lIGMU9qz9_0;
	wire w_dff_A_zKZSf5z96_0;
	wire w_dff_A_6toCtfid3_2;
	wire w_dff_A_1A78CLq23_0;
	wire w_dff_A_DT8YxD0y7_0;
	wire w_dff_A_4W3S1Zbk1_0;
	wire w_dff_A_uwhYlclb7_0;
	wire w_dff_A_FpsAau1M8_0;
	wire w_dff_A_SpVZiSAV6_0;
	wire w_dff_A_EwKqoT1F5_0;
	wire w_dff_A_rPgrdZFb1_0;
	wire w_dff_A_SomvLv1L6_0;
	wire w_dff_A_9cUXX2Kj1_0;
	wire w_dff_A_q9RO1Lzg6_0;
	wire w_dff_A_Kk4RyuDK6_0;
	wire w_dff_A_P2tdFThs6_0;
	wire w_dff_A_7O78XgBo2_0;
	wire w_dff_A_rXPTY3mI5_0;
	wire w_dff_A_muS7FTk72_0;
	wire w_dff_A_6ys0O7wf0_0;
	wire w_dff_A_BexIlYpB4_0;
	wire w_dff_A_xhkygyeT1_0;
	wire w_dff_A_yg0mGmLT6_0;
	wire w_dff_A_lApmStI82_0;
	wire w_dff_A_r1any91t6_0;
	wire w_dff_A_TgB9vsIv2_0;
	wire w_dff_A_1MSyKHFW4_0;
	wire w_dff_A_6OgsMwFq5_0;
	wire w_dff_A_Syyluhm85_0;
	wire w_dff_A_b4VCfP1L0_0;
	wire w_dff_A_JCARhnNj2_0;
	wire w_dff_A_w5pCZ8tj4_0;
	wire w_dff_A_5kMaIGTd8_0;
	wire w_dff_A_SYbL35Ts2_0;
	wire w_dff_A_rpveoWhk8_0;
	wire w_dff_A_LUS4asnZ0_0;
	wire w_dff_A_utui7ytj2_0;
	wire w_dff_A_Kcypql472_0;
	wire w_dff_A_BA1l9tEx7_0;
	wire w_dff_A_bVNmCXeP0_0;
	wire w_dff_A_eShxbMli4_0;
	wire w_dff_A_gx5S1IAV7_0;
	wire w_dff_A_sn3BQ7i11_0;
	wire w_dff_A_KqcQUQlx2_0;
	wire w_dff_A_OJdOHBX93_0;
	wire w_dff_A_PPTuMW0k7_0;
	wire w_dff_A_mtgH9WXw2_0;
	wire w_dff_A_jCkkOiMF2_0;
	wire w_dff_A_UNBsOa8C7_0;
	wire w_dff_A_S8XShES05_0;
	wire w_dff_A_aYJ2pzRp7_0;
	wire w_dff_A_YxHxLVnZ8_0;
	wire w_dff_A_9ctmFtp53_0;
	wire w_dff_A_zIiicibX8_0;
	wire w_dff_A_JgzCnWIR8_0;
	wire w_dff_A_tuDxqGzk5_0;
	wire w_dff_A_0Ucy4uLc4_0;
	wire w_dff_A_50w7r7GH6_0;
	wire w_dff_A_unRZLVOU2_0;
	wire w_dff_A_oHiEz1mj9_2;
	wire w_dff_A_WWEIev9b4_0;
	wire w_dff_A_uA6SoFcj8_0;
	wire w_dff_A_Im5bakEX7_0;
	wire w_dff_A_wwh3wwVl4_0;
	wire w_dff_A_pCktsyqg6_0;
	wire w_dff_A_XarRVOir2_0;
	wire w_dff_A_ICpnhRlR4_0;
	wire w_dff_A_ElF2a2Pl4_0;
	wire w_dff_A_dmInaRWU6_0;
	wire w_dff_A_8chgmXkn3_0;
	wire w_dff_A_aIfZjx4G2_0;
	wire w_dff_A_czBZEWN88_0;
	wire w_dff_A_YpT2eter7_0;
	wire w_dff_A_GRhhVCMk5_0;
	wire w_dff_A_26MYKpXU1_0;
	wire w_dff_A_7M7Y0dV11_0;
	wire w_dff_A_8plRAxtm9_0;
	wire w_dff_A_dSTa3YCe5_0;
	wire w_dff_A_8ryPOv5L2_0;
	wire w_dff_A_0vaBFGXN1_0;
	wire w_dff_A_QMaXO7Iw3_0;
	wire w_dff_A_HocgjUo00_0;
	wire w_dff_A_SLpt4ERs3_0;
	wire w_dff_A_qyeJ6crN4_0;
	wire w_dff_A_WJ0JzlSi6_0;
	wire w_dff_A_hHFyBcm03_0;
	wire w_dff_A_J2WU4fNO3_0;
	wire w_dff_A_jIC19Oib5_0;
	wire w_dff_A_4towJrA42_0;
	wire w_dff_A_W70XScJL3_0;
	wire w_dff_A_su1sO7qz0_0;
	wire w_dff_A_Nb2pKhfa6_0;
	wire w_dff_A_eBsCWehA7_0;
	wire w_dff_A_wn4ZLpoS3_0;
	wire w_dff_A_alTNogDg2_0;
	wire w_dff_A_tdBlQ9uE9_0;
	wire w_dff_A_PVQwOhb35_0;
	wire w_dff_A_qkcyUDQB5_0;
	wire w_dff_A_9uT8iI8J1_0;
	wire w_dff_A_KIEFJ4uB8_0;
	wire w_dff_A_SshSlihQ9_0;
	wire w_dff_A_2DiWrGUt5_0;
	wire w_dff_A_KCmVgIDG9_0;
	wire w_dff_A_KGvGrEZY2_0;
	wire w_dff_A_c4XxgjSx9_0;
	wire w_dff_A_eR3kaN9e3_0;
	wire w_dff_A_wVtDgxO92_0;
	wire w_dff_A_vS3u9BTU9_0;
	wire w_dff_A_71hOUxa46_0;
	wire w_dff_A_wCDoon3U0_0;
	wire w_dff_A_VRpSlWHe7_0;
	wire w_dff_A_mO9XADgl5_0;
	wire w_dff_A_mAXKtItz3_0;
	wire w_dff_A_Rbm3HLMi5_2;
	wire w_dff_A_171O33842_0;
	wire w_dff_A_DgfunnHf5_0;
	wire w_dff_A_1XEqnQNl3_0;
	wire w_dff_A_Itlvq3gT1_0;
	wire w_dff_A_AQvVTgB18_0;
	wire w_dff_A_rt7aZmnp6_0;
	wire w_dff_A_rYS2JgCZ8_0;
	wire w_dff_A_n08vK04M5_0;
	wire w_dff_A_A9qrLozT8_0;
	wire w_dff_A_STfqNvTT5_0;
	wire w_dff_A_DLGn9dEN8_0;
	wire w_dff_A_q4Bm408v2_0;
	wire w_dff_A_xtWdB1hM3_0;
	wire w_dff_A_rdPXo40U9_0;
	wire w_dff_A_0EUS7Gy69_0;
	wire w_dff_A_m60602m17_0;
	wire w_dff_A_UsNhS3ZC6_0;
	wire w_dff_A_JUsV8DUM7_0;
	wire w_dff_A_PprRIjDj7_0;
	wire w_dff_A_VG0Dc0401_0;
	wire w_dff_A_w6xc5oFK2_0;
	wire w_dff_A_DAZddbCR9_0;
	wire w_dff_A_e4Zjc54A7_0;
	wire w_dff_A_IvS6FEvt9_0;
	wire w_dff_A_N0mB9gaT8_0;
	wire w_dff_A_S3Cycj0C1_0;
	wire w_dff_A_vIrNo3oQ7_0;
	wire w_dff_A_Qt9cfgkr9_0;
	wire w_dff_A_dtsgTO692_0;
	wire w_dff_A_xXp27jWL2_0;
	wire w_dff_A_oaq6qhw19_0;
	wire w_dff_A_sPKFS5bJ4_0;
	wire w_dff_A_H3oeM2KD5_0;
	wire w_dff_A_EdoQ8exD1_0;
	wire w_dff_A_oz8yjHUa0_0;
	wire w_dff_A_wxH53mKv5_0;
	wire w_dff_A_UXx9YtCx2_0;
	wire w_dff_A_Fs05k84w1_0;
	wire w_dff_A_ukihaXIE7_0;
	wire w_dff_A_LsGwcZjm2_0;
	wire w_dff_A_CilGgzuw8_0;
	wire w_dff_A_cmY3SbYL4_0;
	wire w_dff_A_vGdK8Ez57_0;
	wire w_dff_A_efN5jWQA2_0;
	wire w_dff_A_N5qTMZjD4_0;
	wire w_dff_A_qi3aoIvW9_0;
	wire w_dff_A_VLbPaEW49_0;
	wire w_dff_A_lHUTu3Ql0_0;
	wire w_dff_A_lcM46GUp5_0;
	wire w_dff_A_3EWNILvx8_0;
	wire w_dff_A_nwOyaoey4_2;
	wire w_dff_A_X9oxnlGG7_0;
	wire w_dff_A_MdrQzZCY2_0;
	wire w_dff_A_VplQJjIg6_0;
	wire w_dff_A_Jk7DRYxx6_0;
	wire w_dff_A_xGAsp6qN3_0;
	wire w_dff_A_EMZY7AgU3_0;
	wire w_dff_A_tmHqdvq06_0;
	wire w_dff_A_SdTKA03y4_0;
	wire w_dff_A_dCdlsUtN6_0;
	wire w_dff_A_Rh70a2QI7_0;
	wire w_dff_A_NYsT8Ru43_0;
	wire w_dff_A_hz06ag0v6_0;
	wire w_dff_A_z7HCUJXW2_0;
	wire w_dff_A_htzWotAw5_0;
	wire w_dff_A_bDjX3uyT9_0;
	wire w_dff_A_8JbD8Mhb1_0;
	wire w_dff_A_lmeM88u52_0;
	wire w_dff_A_cDuUjgib5_0;
	wire w_dff_A_hAmdzvUy5_0;
	wire w_dff_A_tBiijj7F5_0;
	wire w_dff_A_iCFNLp680_0;
	wire w_dff_A_FfWlSijm1_0;
	wire w_dff_A_oI5hKF827_0;
	wire w_dff_A_eL1AppEj4_0;
	wire w_dff_A_o8ntKq7g2_0;
	wire w_dff_A_xxlrpDic0_0;
	wire w_dff_A_bryDQU6H2_0;
	wire w_dff_A_OnUyEe4a4_0;
	wire w_dff_A_b1OGVNak8_0;
	wire w_dff_A_pdhXn80u2_0;
	wire w_dff_A_mJ2pnWn60_0;
	wire w_dff_A_UhzvvQa80_0;
	wire w_dff_A_E0O0qPjW6_0;
	wire w_dff_A_3f0HYPBW2_0;
	wire w_dff_A_VnIb08re1_0;
	wire w_dff_A_4ELMRuYw3_0;
	wire w_dff_A_iTXTK2Dw1_0;
	wire w_dff_A_pPoAfbmZ8_0;
	wire w_dff_A_P4bBWatu1_0;
	wire w_dff_A_5uOQzi5I1_0;
	wire w_dff_A_W1c0Qucw6_0;
	wire w_dff_A_XMNoKD2T4_0;
	wire w_dff_A_Ob7pC4jD4_0;
	wire w_dff_A_Fa1pGlJZ8_0;
	wire w_dff_A_KAdki1ij5_0;
	wire w_dff_A_Wja5gqcN2_0;
	wire w_dff_A_YIEnXGgf1_0;
	wire w_dff_A_Vd7i4kR94_2;
	wire w_dff_A_Pu9Wjaa81_0;
	wire w_dff_A_y832RBgu8_0;
	wire w_dff_A_2HY3uVQV7_0;
	wire w_dff_A_Eh1vioIX1_0;
	wire w_dff_A_U6Jo0qeT7_0;
	wire w_dff_A_qrJIZ9aJ4_0;
	wire w_dff_A_QOg5krL15_0;
	wire w_dff_A_PeBKsD8r3_0;
	wire w_dff_A_ruFNp6fX8_0;
	wire w_dff_A_voWj35FN8_0;
	wire w_dff_A_sXUZFv1v8_0;
	wire w_dff_A_rVMVXYnb2_0;
	wire w_dff_A_ngOg0wGB5_0;
	wire w_dff_A_YbGuxqbD1_0;
	wire w_dff_A_ibqyDZsC2_0;
	wire w_dff_A_mEkAvLwo5_0;
	wire w_dff_A_9JRzzrQQ1_0;
	wire w_dff_A_PfmQXbOq6_0;
	wire w_dff_A_5iqj2tZi3_0;
	wire w_dff_A_lB2yMDCX9_0;
	wire w_dff_A_f3F18Xvh9_0;
	wire w_dff_A_CAV4BSWD0_0;
	wire w_dff_A_K8iX0db10_0;
	wire w_dff_A_Z8TAfvkZ8_0;
	wire w_dff_A_3YbNqBzd0_0;
	wire w_dff_A_BrkJvYdD8_0;
	wire w_dff_A_DhkUnXQC1_0;
	wire w_dff_A_nd5FsRW52_0;
	wire w_dff_A_nBhH7AQT1_0;
	wire w_dff_A_MwUq6KdQ6_0;
	wire w_dff_A_Bp9tMnD25_0;
	wire w_dff_A_n2iIoE575_0;
	wire w_dff_A_HNyFd3XT2_0;
	wire w_dff_A_f0fxSfn54_0;
	wire w_dff_A_bI00JPe37_0;
	wire w_dff_A_0sIfIjAV3_0;
	wire w_dff_A_CKX7qzNz6_0;
	wire w_dff_A_g7OldxJj7_0;
	wire w_dff_A_1dQWdZgN8_0;
	wire w_dff_A_PbxyKYi87_0;
	wire w_dff_A_2KYOE4Va3_0;
	wire w_dff_A_escM5kvZ4_0;
	wire w_dff_A_NlBn5b4h2_0;
	wire w_dff_A_XNdtygn63_0;
	wire w_dff_A_guWKCtIU7_2;
	wire w_dff_A_lZJWPPFQ8_0;
	wire w_dff_A_SRBWEpiC6_0;
	wire w_dff_A_JN3xHNET9_0;
	wire w_dff_A_7iVXD8Sp4_0;
	wire w_dff_A_OUTL29Vo9_0;
	wire w_dff_A_eXcYIxyU9_0;
	wire w_dff_A_fuT2LR7C2_0;
	wire w_dff_A_bibjArTY6_0;
	wire w_dff_A_aEm5TNCV5_0;
	wire w_dff_A_6X0Hkh105_0;
	wire w_dff_A_LxsGgTfI2_0;
	wire w_dff_A_RUjfs1g04_0;
	wire w_dff_A_5frHibc22_0;
	wire w_dff_A_Lx6Rpnzz6_0;
	wire w_dff_A_j8yhVrs60_0;
	wire w_dff_A_FBuJaati5_0;
	wire w_dff_A_0njTq2o26_0;
	wire w_dff_A_0k8lcele9_0;
	wire w_dff_A_I2mqRNHs6_0;
	wire w_dff_A_cM7FXky90_0;
	wire w_dff_A_ndKk4ywE9_0;
	wire w_dff_A_rFyx1reS0_0;
	wire w_dff_A_N3nbda6R0_0;
	wire w_dff_A_BwdpbHXw3_0;
	wire w_dff_A_GIkqeymX2_0;
	wire w_dff_A_GC9J6uZz8_0;
	wire w_dff_A_ZVpwNGuK0_0;
	wire w_dff_A_MFiTvBbX4_0;
	wire w_dff_A_MaHDXhzZ9_0;
	wire w_dff_A_sDLdcoCN1_0;
	wire w_dff_A_dOPFCIKj0_0;
	wire w_dff_A_dngdOybR0_0;
	wire w_dff_A_HYouyW4f7_0;
	wire w_dff_A_P4px86Pf8_0;
	wire w_dff_A_6Gs0xb4l6_0;
	wire w_dff_A_fxvU3Dhu5_0;
	wire w_dff_A_0mg0BSQh3_0;
	wire w_dff_A_QzLDgINi9_0;
	wire w_dff_A_Zf4DBYiT4_0;
	wire w_dff_A_TsWhlDO92_0;
	wire w_dff_A_6nk7GkCt1_0;
	wire w_dff_A_8K6sinQo2_2;
	wire w_dff_A_GfPQn7GX3_0;
	wire w_dff_A_JNnXggAV3_0;
	wire w_dff_A_RXF1Y7ws6_0;
	wire w_dff_A_ofXrKFV59_0;
	wire w_dff_A_f4fQlerU7_0;
	wire w_dff_A_1fN5ouJP5_0;
	wire w_dff_A_zU7Jeund6_0;
	wire w_dff_A_DdzN2HBs7_0;
	wire w_dff_A_M7zlZhe93_0;
	wire w_dff_A_yssQJ5ap2_0;
	wire w_dff_A_A7J1Gk0G7_0;
	wire w_dff_A_Dw9LjXUF7_0;
	wire w_dff_A_lyw1ITQV8_0;
	wire w_dff_A_kWwfDxtK4_0;
	wire w_dff_A_cCr8Tswj7_0;
	wire w_dff_A_nFgjYuYT0_0;
	wire w_dff_A_plHmViy87_0;
	wire w_dff_A_BR26NNCS8_0;
	wire w_dff_A_7gPHeTGa1_0;
	wire w_dff_A_WiaY6IOK6_0;
	wire w_dff_A_Vo80r9JR8_0;
	wire w_dff_A_SpoRhbOs9_0;
	wire w_dff_A_sgO7idng4_0;
	wire w_dff_A_SMpKunVy7_0;
	wire w_dff_A_JurrIsLZ7_0;
	wire w_dff_A_jYyqzmar3_0;
	wire w_dff_A_jqO2OKA84_0;
	wire w_dff_A_XL3D0XrL0_0;
	wire w_dff_A_mzN4nRDF2_0;
	wire w_dff_A_EQUZUBrn5_0;
	wire w_dff_A_tYOakAXO1_0;
	wire w_dff_A_KCFnn8lv5_0;
	wire w_dff_A_YGZhVVr04_0;
	wire w_dff_A_jtk7yuY95_0;
	wire w_dff_A_R3asqZOm8_0;
	wire w_dff_A_KAtYWEx24_0;
	wire w_dff_A_xAs5my3L6_0;
	wire w_dff_A_TkAKGVbx0_0;
	wire w_dff_A_bgSyLykw2_2;
	wire w_dff_A_ntCRt9Xm2_0;
	wire w_dff_A_Sgrhl8zQ8_0;
	wire w_dff_A_ZePkzJr66_0;
	wire w_dff_A_dhwgM6kh5_0;
	wire w_dff_A_BoEvaWQw6_0;
	wire w_dff_A_pGVXO9u82_0;
	wire w_dff_A_VJPXJRPA5_0;
	wire w_dff_A_7kCwRQcM5_0;
	wire w_dff_A_Kxs5Dtx22_0;
	wire w_dff_A_6aNgm7qc6_0;
	wire w_dff_A_1my3cUMa0_0;
	wire w_dff_A_iVHRFBGG3_0;
	wire w_dff_A_rU7hAwhA0_0;
	wire w_dff_A_me30UN9W4_0;
	wire w_dff_A_ShzFT1zM2_0;
	wire w_dff_A_ZTjzSqwx2_0;
	wire w_dff_A_3U7yrEdy9_0;
	wire w_dff_A_0ATY7b6R9_0;
	wire w_dff_A_WwRyUwzb2_0;
	wire w_dff_A_hYAG7MK33_0;
	wire w_dff_A_SDJMsobg9_0;
	wire w_dff_A_fSOs6jWy6_0;
	wire w_dff_A_DczPKTpz3_0;
	wire w_dff_A_kCL466yC7_0;
	wire w_dff_A_H7OGRi6A5_0;
	wire w_dff_A_bnWgRYoh5_0;
	wire w_dff_A_YS7a8fLk6_0;
	wire w_dff_A_LmWMfktV1_0;
	wire w_dff_A_lwv9BZYb9_0;
	wire w_dff_A_tSjzfsgx4_0;
	wire w_dff_A_u8VmXTca9_0;
	wire w_dff_A_oojI1ZYQ6_0;
	wire w_dff_A_oIIRsrEb9_0;
	wire w_dff_A_OpzbgR6U0_0;
	wire w_dff_A_XgOMPC0j8_0;
	wire w_dff_A_HUPrWpUI2_2;
	wire w_dff_A_64QSWXVK6_0;
	wire w_dff_A_PFHLJvTo9_0;
	wire w_dff_A_pZdJIG9B4_0;
	wire w_dff_A_9LDmQsRC7_0;
	wire w_dff_A_bWPyAhAK8_0;
	wire w_dff_A_CEfgBgMP8_0;
	wire w_dff_A_HaxRrwB50_0;
	wire w_dff_A_WYz39Sl44_0;
	wire w_dff_A_Ju5LJsON5_0;
	wire w_dff_A_5IYbzKHa0_0;
	wire w_dff_A_FhudYR129_0;
	wire w_dff_A_WQMPsREa2_0;
	wire w_dff_A_DcRdYJQx1_0;
	wire w_dff_A_3NVsXQ8R2_0;
	wire w_dff_A_I8O7RJY53_0;
	wire w_dff_A_gEj68g6m7_0;
	wire w_dff_A_Rj970DGQ4_0;
	wire w_dff_A_JXVDUVx24_0;
	wire w_dff_A_ub5KuGH98_0;
	wire w_dff_A_PXFymSUC6_0;
	wire w_dff_A_9AAylEAF5_0;
	wire w_dff_A_bKlsDN5c9_0;
	wire w_dff_A_tkELLfEE5_0;
	wire w_dff_A_FuWYUGHm4_0;
	wire w_dff_A_EgKCktUe0_0;
	wire w_dff_A_HOOPbwb98_0;
	wire w_dff_A_KuElOmoQ7_0;
	wire w_dff_A_Eb4f4YI32_0;
	wire w_dff_A_Y9VpNMDr4_0;
	wire w_dff_A_Az6wZtah5_0;
	wire w_dff_A_DseTCSk85_0;
	wire w_dff_A_CC5pY0xT4_0;
	wire w_dff_A_dkRXDqWE6_2;
	wire w_dff_A_yiZ3IYnb0_0;
	wire w_dff_A_GRbEqwlc5_0;
	wire w_dff_A_yNueZH6b5_0;
	wire w_dff_A_9aGsA8D06_0;
	wire w_dff_A_G5bZRDvy3_0;
	wire w_dff_A_SW2Ij6fh7_0;
	wire w_dff_A_Wqyn8iDX4_0;
	wire w_dff_A_A9O1UhMb5_0;
	wire w_dff_A_jgzE7U3v1_0;
	wire w_dff_A_RRDgoQ4P2_0;
	wire w_dff_A_JO6bXnkI9_0;
	wire w_dff_A_4qBoBvWY9_0;
	wire w_dff_A_mOp6pj7s1_0;
	wire w_dff_A_DFjpI4MN9_0;
	wire w_dff_A_H81wNIv47_0;
	wire w_dff_A_cRG8EHzL2_0;
	wire w_dff_A_QTKL9rY99_0;
	wire w_dff_A_adSknmPh5_0;
	wire w_dff_A_Hzp84igx3_0;
	wire w_dff_A_TQiCZPPG1_0;
	wire w_dff_A_7CdSWMpS2_0;
	wire w_dff_A_nMYswItO5_0;
	wire w_dff_A_kDn3tEb55_0;
	wire w_dff_A_hIceY3HB1_0;
	wire w_dff_A_Bt7icd6K9_0;
	wire w_dff_A_K8uXSM0B5_0;
	wire w_dff_A_R5A5ubKE6_0;
	wire w_dff_A_rIj6fq011_0;
	wire w_dff_A_ukbNP34h2_0;
	wire w_dff_A_XP7KI9S09_2;
	wire w_dff_A_QYT2rliR4_0;
	wire w_dff_A_N9SMenpp5_0;
	wire w_dff_A_UgK9U5FT0_0;
	wire w_dff_A_7PBadlrA1_0;
	wire w_dff_A_y2udl6fQ1_0;
	wire w_dff_A_oVl7XIuV5_0;
	wire w_dff_A_7ZQ1NyRU9_0;
	wire w_dff_A_HoujgT4A7_0;
	wire w_dff_A_mIL9qtZM0_0;
	wire w_dff_A_SxwH9dxH1_0;
	wire w_dff_A_35805j6E7_0;
	wire w_dff_A_6aAhYsJY9_0;
	wire w_dff_A_LVMOG8c84_0;
	wire w_dff_A_asFbVqi07_0;
	wire w_dff_A_OwHt3ajN5_0;
	wire w_dff_A_8bxLa27V0_0;
	wire w_dff_A_0w5p6SzL5_0;
	wire w_dff_A_G2RhsFcW6_0;
	wire w_dff_A_h6gZP8qM5_0;
	wire w_dff_A_UtcDfwkz2_0;
	wire w_dff_A_SKWDjgK36_0;
	wire w_dff_A_lsoqaHTn7_0;
	wire w_dff_A_n4q0mMOi0_0;
	wire w_dff_A_quTNwDxI6_0;
	wire w_dff_A_rZolB5tP1_0;
	wire w_dff_A_5z3SpYsC8_0;
	wire w_dff_A_L2Nd2Iat2_0;
	wire w_dff_A_muYCmXs49_2;
	wire w_dff_A_RhmMgHzJ2_0;
	wire w_dff_A_Y1oVLQD46_0;
	wire w_dff_A_xdwiQXY37_0;
	wire w_dff_A_PkRSJyfj3_0;
	wire w_dff_A_4gLnuB6Z8_0;
	wire w_dff_A_asP64sgb1_0;
	wire w_dff_A_dByGgPP52_0;
	wire w_dff_A_jDheKlDP8_0;
	wire w_dff_A_pWlC6zdb2_0;
	wire w_dff_A_uehCxuEK1_0;
	wire w_dff_A_DYt4QheT0_0;
	wire w_dff_A_aGaicp3P0_0;
	wire w_dff_A_1i05DgVs6_0;
	wire w_dff_A_2stMxxT16_0;
	wire w_dff_A_5YBeaBvd9_0;
	wire w_dff_A_KDw3NH4l1_0;
	wire w_dff_A_lEuD209Z0_0;
	wire w_dff_A_mir0XGtj0_0;
	wire w_dff_A_Jj3fJt1g0_0;
	wire w_dff_A_kpQ2LYBI7_0;
	wire w_dff_A_agb1MY1J7_0;
	wire w_dff_A_yQbmpn760_0;
	wire w_dff_A_l8Ot5fQK3_0;
	wire w_dff_A_NSXzSIEr5_0;
	wire w_dff_A_smKVEayf3_0;
	wire w_dff_A_MsaMqHPq5_2;
	wire w_dff_A_EWidRBpa7_0;
	wire w_dff_A_J3bF2UZ40_0;
	wire w_dff_A_NU4fQv7S1_0;
	wire w_dff_A_e6F23xlq3_0;
	wire w_dff_A_MR7cQP7V6_0;
	wire w_dff_A_jurMbIww6_0;
	wire w_dff_A_RLAmi19d0_0;
	wire w_dff_A_cY6jLVdC3_0;
	wire w_dff_A_8lanbtLS9_0;
	wire w_dff_A_akO7jPOA8_0;
	wire w_dff_A_llQc2Dv85_0;
	wire w_dff_A_oLB8ljKD0_0;
	wire w_dff_A_okEQeA9W3_0;
	wire w_dff_A_exmAmJc02_0;
	wire w_dff_A_NhFTfx3R2_0;
	wire w_dff_A_OZiNN5vz2_0;
	wire w_dff_A_oZf1kPbn0_0;
	wire w_dff_A_iZqQD9uf0_0;
	wire w_dff_A_gFb0YsbJ8_0;
	wire w_dff_A_EYGGr5a33_0;
	wire w_dff_A_XyirquLk5_0;
	wire w_dff_A_4aciwrKU0_0;
	wire w_dff_A_2xQ6EuHI9_0;
	wire w_dff_A_1vLH8UxP8_0;
	wire w_dff_A_2H3dPpHv5_2;
	wire w_dff_A_zGqYnJ693_0;
	wire w_dff_A_SINlhkzL7_0;
	wire w_dff_A_Bc6xhLxp3_0;
	wire w_dff_A_XyAd7eVI4_0;
	wire w_dff_A_PZ2v6xN74_0;
	wire w_dff_A_bw8PlNid0_0;
	wire w_dff_A_xtiPKrGv5_0;
	wire w_dff_A_eLofanXw5_0;
	wire w_dff_A_PKXkb4Os1_0;
	wire w_dff_A_SRpbTUPX1_0;
	wire w_dff_A_0XXQL3WG8_0;
	wire w_dff_A_TGwhWh9a2_0;
	wire w_dff_A_0TEZQyNz2_0;
	wire w_dff_A_jG0KZhr14_0;
	wire w_dff_A_V4sVFDLJ3_0;
	wire w_dff_A_g5ZRMeTb6_0;
	wire w_dff_A_fewmH9SB0_0;
	wire w_dff_A_MS0plOq66_0;
	wire w_dff_A_DHiYfBnH8_0;
	wire w_dff_A_Sil1Kgkq5_0;
	wire w_dff_A_cy4DZ6lv3_0;
	wire w_dff_A_csOQGDMp5_0;
	wire w_dff_A_nFZwUN7m5_2;
	wire w_dff_A_wCP1GDwg3_0;
	wire w_dff_A_TuJYL9Bw9_0;
	wire w_dff_A_bQHtmJrg1_0;
	wire w_dff_A_EHh4ViMa5_0;
	wire w_dff_A_v1wTa9oT6_0;
	wire w_dff_A_0BRWUEF80_0;
	wire w_dff_A_ZHZDjXgd2_0;
	wire w_dff_A_cDq0aF7i9_0;
	wire w_dff_A_k3rsHM7N8_0;
	wire w_dff_A_kta9keZ81_0;
	wire w_dff_A_JckzmQxj7_0;
	wire w_dff_A_DjcrbS1d8_0;
	wire w_dff_A_lcs140vB1_0;
	wire w_dff_A_rgnMc04L7_0;
	wire w_dff_A_rcswlGYS6_0;
	wire w_dff_A_Nvj4k6Rj6_0;
	wire w_dff_A_n7maCWAC0_0;
	wire w_dff_A_wcRGgzfw3_0;
	wire w_dff_A_p0dNXKDc3_0;
	wire w_dff_A_7A6bt52y7_0;
	wire w_dff_A_BTnUMnAU7_2;
	wire w_dff_A_yDpE8sMw3_0;
	wire w_dff_A_zAbpuylL6_0;
	wire w_dff_A_Jniz9VPd4_0;
	wire w_dff_A_ynRMVfXO9_0;
	wire w_dff_A_CyTXiea32_0;
	wire w_dff_A_cfWCba7g3_0;
	wire w_dff_A_rL3YDsfb0_0;
	wire w_dff_A_5eiugd7Z3_0;
	wire w_dff_A_DzHrCLbt5_0;
	wire w_dff_A_FI9jyE854_0;
	wire w_dff_A_H3LZ7MPh8_0;
	wire w_dff_A_sCCm3opL9_0;
	wire w_dff_A_dYeziSMj6_0;
	wire w_dff_A_vmKejPkQ0_0;
	wire w_dff_A_CJtxRjim8_0;
	wire w_dff_A_1ctpGbgg5_0;
	wire w_dff_A_JKXbp7w75_0;
	wire w_dff_A_LRHSc0ac9_0;
	wire w_dff_A_96BrlB423_2;
	wire w_dff_A_6L2TBEwC3_0;
	wire w_dff_A_ECb3B5yj2_0;
	wire w_dff_A_N9Ade0XG7_0;
	wire w_dff_A_HVjBrLV06_0;
	wire w_dff_A_LMhO7NQ81_0;
	wire w_dff_A_XQ8lBCio4_0;
	wire w_dff_A_EQFvMxPh9_0;
	wire w_dff_A_4RSN6NPj4_0;
	wire w_dff_A_Ge9Wk7tA2_0;
	wire w_dff_A_GPo7kuIa4_0;
	wire w_dff_A_VXvFFCb12_0;
	wire w_dff_A_KZLK5GGh2_0;
	wire w_dff_A_rG1oGnWq8_0;
	wire w_dff_A_BazaDLNT9_0;
	wire w_dff_A_UJbvnSdq0_0;
	wire w_dff_A_Eh2gmav45_0;
	wire w_dff_A_oWs98O0Y7_2;
	wire w_dff_A_YbnRnyt18_0;
	wire w_dff_A_DYu5ZkHt0_0;
	wire w_dff_A_pkr6GAxp8_0;
	wire w_dff_A_3C4cP3FN5_0;
	wire w_dff_A_WxBtqsJX7_0;
	wire w_dff_A_rPkki8Nx6_0;
	wire w_dff_A_AXNVxNfd5_0;
	wire w_dff_A_UcjgaseF0_0;
	wire w_dff_A_rvDdg6zP3_0;
	wire w_dff_A_2U5jOXBD8_0;
	wire w_dff_A_FIRCRgyq9_0;
	wire w_dff_A_PMzcuCJm9_0;
	wire w_dff_A_Qm1n0uAa5_0;
	wire w_dff_A_PRGfI1FU0_0;
	wire w_dff_A_IFaEiPVG2_2;
	wire w_dff_A_g1szHesY8_0;
	wire w_dff_A_TBgoZo4N9_0;
	wire w_dff_A_baN9XbAo0_0;
	wire w_dff_A_RlyKUGeq5_0;
	wire w_dff_A_Sq8ptWYj3_0;
	wire w_dff_A_3t4g6c3I0_0;
	wire w_dff_A_7eom11wB9_0;
	wire w_dff_A_2x5unCXl3_0;
	wire w_dff_A_RJKDsMbD7_0;
	wire w_dff_A_Re64RGVU3_0;
	wire w_dff_A_bFU1C6921_0;
	wire w_dff_A_H4DQHubn4_0;
	wire w_dff_A_iPM9LwlQ1_2;
	wire w_dff_A_BSFUGiiD3_0;
	wire w_dff_A_U6tWwpAv3_0;
	wire w_dff_A_60EC0Zj36_0;
	wire w_dff_A_Ui8GvQhv0_0;
	wire w_dff_A_MtvFY0gW8_0;
	wire w_dff_A_5vIlxAwr8_0;
	wire w_dff_A_ukTT6Mmc0_0;
	wire w_dff_A_e7uD8wLC2_0;
	wire w_dff_A_CmzlbS8M7_0;
	wire w_dff_A_hVZ4EwjM5_0;
	wire w_dff_A_4ZSUinxL1_2;
	wire w_dff_A_8vznccM88_0;
	wire w_dff_A_4EbhWlwH9_0;
	wire w_dff_A_0FB3gmKz9_0;
	wire w_dff_A_I3FHZ6Ns0_0;
	wire w_dff_A_L0s8w6739_0;
	wire w_dff_A_DbJuQ1rh1_0;
	wire w_dff_A_jMcL0vjA6_0;
	wire w_dff_A_Ip7LTZOl9_0;
	wire w_dff_A_jerCFLUD1_2;
	wire w_dff_A_OzM6UivC1_0;
	wire w_dff_A_UwqzvO0V4_0;
	wire w_dff_A_7qdSojmy8_0;
	wire w_dff_A_UFwoG57b5_0;
	wire w_dff_A_NcaGpnbc9_0;
	wire w_dff_A_WS5t0grE8_0;
	wire w_dff_A_AZmphtiy6_2;
	wire w_dff_A_ro53mV445_0;
	wire w_dff_A_yYNv67ns6_0;
	wire w_dff_A_k7BRES2e4_0;
	wire w_dff_A_ihGoirPu7_0;
	wire w_dff_A_VrGQGW8r1_2;
	wire w_dff_A_TSBcsTUK5_0;
	wire w_dff_A_2SWcjTOU1_0;
	wire w_dff_A_JNspNrBf3_2;
	jand g0000(.dina(w_G273gat_7[2]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G273gat_7[1]),.dinb(w_G18gat_7[2]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_G290gat_7[2]),.dinb(w_G1gat_7[0]),.dout(n66),.clk(gclk));
	jor g0003(.dina(n66),.dinb(w_n65_0[1]),.dout(n67),.clk(gclk));
	jand g0004(.dina(w_G290gat_7[1]),.dinb(w_G18gat_7[1]),.dout(n68),.clk(gclk));
	jand g0005(.dina(n68),.dinb(w_G545gat_0),.dout(n69),.clk(gclk));
	jnot g0006(.din(w_n69_0[1]),.dout(n70),.clk(gclk));
	jand g0007(.dina(w_n70_0[1]),.dinb(w_dff_B_bbppiPhb7_1),.dout(w_dff_A_PCFOBIdG2_2),.clk(gclk));
	jand g0008(.dina(w_G307gat_7[2]),.dinb(w_G1gat_6[2]),.dout(n72),.clk(gclk));
	jnot g0009(.din(w_n72_0[1]),.dout(n73),.clk(gclk));
	jnot g0010(.din(w_G18gat_7[0]),.dout(n74),.clk(gclk));
	jnot g0011(.din(w_G290gat_7[0]),.dout(n75),.clk(gclk));
	jor g0012(.dina(w_n75_0[1]),.dinb(n74),.dout(n76),.clk(gclk));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G273gat_7[0]),.dout(n78),.clk(gclk));
	jor g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79),.clk(gclk));
	jand g0016(.dina(n79),.dinb(n76),.dout(n80),.clk(gclk));
	jand g0017(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jand g0018(.dina(w_n81_0[1]),.dinb(w_n65_0[0]),.dout(n82),.clk(gclk));
	jor g0019(.dina(w_n82_1[1]),.dinb(n80),.dout(n83),.clk(gclk));
	jand g0020(.dina(n83),.dinb(w_n70_0[0]),.dout(n84),.clk(gclk));
	jnot g0021(.din(w_n82_1[0]),.dout(n85),.clk(gclk));
	jand g0022(.dina(w_n85_0[1]),.dinb(w_n69_0[0]),.dout(n86),.clk(gclk));
	jor g0023(.dina(w_dff_B_MoKKPG2t4_0),.dinb(w_n84_0[1]),.dout(n87),.clk(gclk));
	jxor g0024(.dina(w_n87_0[1]),.dinb(w_dff_B_FZ3q2YcR3_1),.dout(w_dff_A_gydU51Oe5_2),.clk(gclk));
	jand g0025(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n89),.clk(gclk));
	jnot g0026(.din(w_n89_0[1]),.dout(n90),.clk(gclk));
	jnot g0027(.din(w_n84_0[0]),.dout(n91),.clk(gclk));
	jor g0028(.dina(w_n87_0[0]),.dinb(w_n72_0[0]),.dout(n92),.clk(gclk));
	jand g0029(.dina(n92),.dinb(w_dff_B_hckTMUBH6_1),.dout(n93),.clk(gclk));
	jand g0030(.dina(w_G307gat_7[1]),.dinb(w_G18gat_6[2]),.dout(n94),.clk(gclk));
	jnot g0031(.din(w_n94_0[1]),.dout(n95),.clk(gclk));
	jand g0032(.dina(w_G273gat_6[2]),.dinb(w_G52gat_7[2]),.dout(n96),.clk(gclk));
	jor g0033(.dina(w_n96_0[1]),.dinb(w_n81_0[0]),.dout(n97),.clk(gclk));
	jand g0034(.dina(w_G273gat_6[1]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G290gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jand g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100),.clk(gclk));
	jnot g0037(.din(w_n100_1[1]),.dout(n101),.clk(gclk));
	jand g0038(.dina(w_n101_0[2]),.dinb(n97),.dout(n102),.clk(gclk));
	jor g0039(.dina(n102),.dinb(w_n82_0[2]),.dout(n103),.clk(gclk));
	jand g0040(.dina(w_n101_0[1]),.dinb(w_n82_0[1]),.dout(n104),.clk(gclk));
	jnot g0041(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jand g0042(.dina(n105),.dinb(w_n103_0[1]),.dout(n106),.clk(gclk));
	jxor g0043(.dina(n106),.dinb(n95),.dout(n107),.clk(gclk));
	jxor g0044(.dina(w_n107_0[1]),.dinb(w_n93_0[1]),.dout(n108),.clk(gclk));
	jxor g0045(.dina(w_n108_0[1]),.dinb(w_dff_B_PgYh4dwy6_1),.dout(w_dff_A_prb6lJFG0_2),.clk(gclk));
	jand g0046(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n110),.clk(gclk));
	jnot g0047(.din(w_n110_0[1]),.dout(n111),.clk(gclk));
	jnot g0048(.din(w_n107_0[0]),.dout(n112),.clk(gclk));
	jor g0049(.dina(n112),.dinb(w_n93_0[0]),.dout(n113),.clk(gclk));
	jor g0050(.dina(w_n108_0[0]),.dinb(w_n89_0[0]),.dout(n114),.clk(gclk));
	jand g0051(.dina(n114),.dinb(w_dff_B_pS4HvURR3_1),.dout(n115),.clk(gclk));
	jand g0052(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n116),.clk(gclk));
	jnot g0053(.din(w_n116_0[1]),.dout(n117),.clk(gclk));
	jor g0054(.dina(w_n75_0[0]),.dinb(w_n77_0[0]),.dout(n118),.clk(gclk));
	jnot g0055(.din(w_G52gat_7[0]),.dout(n119),.clk(gclk));
	jor g0056(.dina(w_n78_0[0]),.dinb(n119),.dout(n120),.clk(gclk));
	jand g0057(.dina(n120),.dinb(n118),.dout(n121),.clk(gclk));
	jor g0058(.dina(w_n100_1[0]),.dinb(n121),.dout(n122),.clk(gclk));
	jand g0059(.dina(n122),.dinb(w_n85_0[0]),.dout(n123),.clk(gclk));
	jor g0060(.dina(w_n104_0[0]),.dinb(n123),.dout(n124),.clk(gclk));
	jor g0061(.dina(n124),.dinb(w_n94_0[0]),.dout(n125),.clk(gclk));
	jand g0062(.dina(n125),.dinb(w_n103_0[0]),.dout(n126),.clk(gclk));
	jand g0063(.dina(w_G307gat_7[0]),.dinb(w_G35gat_6[2]),.dout(n127),.clk(gclk));
	jnot g0064(.din(n127),.dout(n128),.clk(gclk));
	jand g0065(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[1]),.dout(n129),.clk(gclk));
	jor g0066(.dina(w_n129_0[1]),.dinb(w_n99_0[0]),.dout(n130),.clk(gclk));
	jand g0067(.dina(w_G290gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n131),.clk(gclk));
	jand g0068(.dina(w_n131_0[1]),.dinb(w_n96_0[0]),.dout(n132),.clk(gclk));
	jnot g0069(.din(w_n132_0[2]),.dout(n133),.clk(gclk));
	jand g0070(.dina(w_n133_0[2]),.dinb(w_n130_0[1]),.dout(n134),.clk(gclk));
	jor g0071(.dina(n134),.dinb(w_n100_0[2]),.dout(n135),.clk(gclk));
	jand g0072(.dina(w_n133_0[1]),.dinb(w_n100_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(n136),.dout(n137),.clk(gclk));
	jand g0074(.dina(n137),.dinb(n135),.dout(n138),.clk(gclk));
	jxor g0075(.dina(w_n138_0[1]),.dinb(w_n128_0[1]),.dout(n139),.clk(gclk));
	jnot g0076(.din(w_n139_0[1]),.dout(n140),.clk(gclk));
	jxor g0077(.dina(w_n140_0[1]),.dinb(w_n126_0[2]),.dout(n141),.clk(gclk));
	jxor g0078(.dina(n141),.dinb(n117),.dout(n142),.clk(gclk));
	jxor g0079(.dina(w_n142_0[1]),.dinb(w_n115_0[1]),.dout(n143),.clk(gclk));
	jxor g0080(.dina(w_n143_0[1]),.dinb(w_dff_B_yn8sG5gV0_1),.dout(w_dff_A_wOXl4S3M1_2),.clk(gclk));
	jand g0081(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n145),.clk(gclk));
	jnot g0082(.din(w_n145_0[1]),.dout(n146),.clk(gclk));
	jnot g0083(.din(w_n142_0[0]),.dout(n147),.clk(gclk));
	jor g0084(.dina(n147),.dinb(w_n115_0[0]),.dout(n148),.clk(gclk));
	jor g0085(.dina(w_n143_0[0]),.dinb(w_n110_0[0]),.dout(n149),.clk(gclk));
	jand g0086(.dina(n149),.dinb(w_dff_B_Qkzi8O9h3_1),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n151),.clk(gclk));
	jnot g0088(.din(w_n151_0[1]),.dout(n152),.clk(gclk));
	jor g0089(.dina(w_n140_0[0]),.dinb(w_n126_0[1]),.dout(n153),.clk(gclk));
	jxor g0090(.dina(w_n139_0[0]),.dinb(w_n126_0[0]),.dout(n154),.clk(gclk));
	jor g0091(.dina(n154),.dinb(w_n116_0[0]),.dout(n155),.clk(gclk));
	jand g0092(.dina(n155),.dinb(n153),.dout(n156),.clk(gclk));
	jand g0093(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n157),.clk(gclk));
	jnot g0094(.din(n157),.dout(n158),.clk(gclk));
	jnot g0095(.din(w_n130_0[0]),.dout(n159),.clk(gclk));
	jor g0096(.dina(w_n132_0[1]),.dinb(n159),.dout(n160),.clk(gclk));
	jand g0097(.dina(n160),.dinb(w_n101_0[0]),.dout(n161),.clk(gclk));
	jand g0098(.dina(w_n138_0[0]),.dinb(w_n128_0[0]),.dout(n162),.clk(gclk));
	jor g0099(.dina(n162),.dinb(n161),.dout(n163),.clk(gclk));
	jand g0100(.dina(w_G307gat_6[2]),.dinb(w_G52gat_6[2]),.dout(n164),.clk(gclk));
	jnot g0101(.din(n164),.dout(n165),.clk(gclk));
	jand g0102(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n166),.clk(gclk));
	jor g0103(.dina(w_n166_0[1]),.dinb(w_n131_0[0]),.dout(n167),.clk(gclk));
	jand g0104(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n168),.clk(gclk));
	jand g0105(.dina(w_n168_0[1]),.dinb(w_n129_0[0]),.dout(n169),.clk(gclk));
	jnot g0106(.din(w_n169_0[2]),.dout(n170),.clk(gclk));
	jand g0107(.dina(w_n170_0[1]),.dinb(n167),.dout(n171),.clk(gclk));
	jor g0108(.dina(n171),.dinb(w_n132_0[0]),.dout(n172),.clk(gclk));
	jor g0109(.dina(w_n169_0[1]),.dinb(w_n133_0[0]),.dout(n173),.clk(gclk));
	jand g0110(.dina(n173),.dinb(w_n172_0[1]),.dout(n174),.clk(gclk));
	jxor g0111(.dina(w_n174_0[1]),.dinb(w_n165_0[1]),.dout(n175),.clk(gclk));
	jxor g0112(.dina(w_n175_0[1]),.dinb(w_n163_0[1]),.dout(n176),.clk(gclk));
	jxor g0113(.dina(w_n176_0[1]),.dinb(w_n158_0[1]),.dout(n177),.clk(gclk));
	jnot g0114(.din(w_n177_0[1]),.dout(n178),.clk(gclk));
	jxor g0115(.dina(w_n178_0[1]),.dinb(w_n156_0[2]),.dout(n179),.clk(gclk));
	jxor g0116(.dina(n179),.dinb(n152),.dout(n180),.clk(gclk));
	jxor g0117(.dina(w_n180_0[1]),.dinb(w_n150_0[1]),.dout(n181),.clk(gclk));
	jxor g0118(.dina(w_n181_0[1]),.dinb(w_dff_B_mpRUR74K0_1),.dout(w_dff_A_SMosFExk3_2),.clk(gclk));
	jand g0119(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n183),.clk(gclk));
	jnot g0120(.din(w_n183_0[1]),.dout(n184),.clk(gclk));
	jnot g0121(.din(w_n180_0[0]),.dout(n185),.clk(gclk));
	jor g0122(.dina(n185),.dinb(w_n150_0[0]),.dout(n186),.clk(gclk));
	jor g0123(.dina(w_n181_0[0]),.dinb(w_n145_0[0]),.dout(n187),.clk(gclk));
	jand g0124(.dina(n187),.dinb(w_dff_B_rPUbm3kx1_1),.dout(n188),.clk(gclk));
	jand g0125(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n189),.clk(gclk));
	jnot g0126(.din(w_n189_0[1]),.dout(n190),.clk(gclk));
	jor g0127(.dina(w_n178_0[0]),.dinb(w_n156_0[1]),.dout(n191),.clk(gclk));
	jxor g0128(.dina(w_n177_0[0]),.dinb(w_n156_0[0]),.dout(n192),.clk(gclk));
	jor g0129(.dina(n192),.dinb(w_n151_0[0]),.dout(n193),.clk(gclk));
	jand g0130(.dina(n193),.dinb(n191),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n195),.clk(gclk));
	jnot g0132(.din(n195),.dout(n196),.clk(gclk));
	jand g0133(.dina(w_n175_0[0]),.dinb(w_n163_0[0]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_n176_0[0]),.dinb(w_n158_0[0]),.dout(n198),.clk(gclk));
	jor g0135(.dina(n198),.dinb(n197),.dout(n199),.clk(gclk));
	jand g0136(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n200),.clk(gclk));
	jnot g0137(.din(n200),.dout(n201),.clk(gclk));
	jnot g0138(.din(w_n172_0[0]),.dout(n202),.clk(gclk));
	jand g0139(.dina(w_n174_0[0]),.dinb(w_n165_0[0]),.dout(n203),.clk(gclk));
	jor g0140(.dina(n203),.dinb(n202),.dout(n204),.clk(gclk));
	jand g0141(.dina(w_G307gat_6[1]),.dinb(w_G69gat_6[2]),.dout(n205),.clk(gclk));
	jnot g0142(.din(n205),.dout(n206),.clk(gclk));
	jand g0143(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n207),.clk(gclk));
	jor g0144(.dina(w_n207_0[1]),.dinb(w_n168_0[0]),.dout(n208),.clk(gclk));
	jand g0145(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n209),.clk(gclk));
	jand g0146(.dina(w_n209_0[1]),.dinb(w_n166_0[0]),.dout(n210),.clk(gclk));
	jnot g0147(.din(w_n210_1[1]),.dout(n211),.clk(gclk));
	jand g0148(.dina(n211),.dinb(n208),.dout(n212),.clk(gclk));
	jor g0149(.dina(n212),.dinb(w_n169_0[0]),.dout(n213),.clk(gclk));
	jor g0150(.dina(w_n210_1[0]),.dinb(w_n170_0[0]),.dout(n214),.clk(gclk));
	jand g0151(.dina(n214),.dinb(w_n213_0[1]),.dout(n215),.clk(gclk));
	jxor g0152(.dina(w_n215_0[1]),.dinb(w_n206_0[1]),.dout(n216),.clk(gclk));
	jxor g0153(.dina(w_n216_0[1]),.dinb(w_n204_0[1]),.dout(n217),.clk(gclk));
	jxor g0154(.dina(w_n217_0[1]),.dinb(w_n201_0[1]),.dout(n218),.clk(gclk));
	jxor g0155(.dina(w_n218_0[1]),.dinb(w_n199_0[1]),.dout(n219),.clk(gclk));
	jxor g0156(.dina(w_n219_0[1]),.dinb(w_n196_0[1]),.dout(n220),.clk(gclk));
	jnot g0157(.din(w_n220_0[1]),.dout(n221),.clk(gclk));
	jxor g0158(.dina(w_n221_0[1]),.dinb(w_n194_0[2]),.dout(n222),.clk(gclk));
	jxor g0159(.dina(n222),.dinb(n190),.dout(n223),.clk(gclk));
	jxor g0160(.dina(w_n223_0[1]),.dinb(w_n188_0[1]),.dout(n224),.clk(gclk));
	jxor g0161(.dina(w_n224_0[1]),.dinb(w_dff_B_6oZvyY0P2_1),.dout(w_dff_A_6toCtfid3_2),.clk(gclk));
	jand g0162(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n226),.clk(gclk));
	jnot g0163(.din(w_n226_0[1]),.dout(n227),.clk(gclk));
	jnot g0164(.din(w_n223_0[0]),.dout(n228),.clk(gclk));
	jor g0165(.dina(n228),.dinb(w_n188_0[0]),.dout(n229),.clk(gclk));
	jor g0166(.dina(w_n224_0[0]),.dinb(w_n183_0[0]),.dout(n230),.clk(gclk));
	jand g0167(.dina(n230),.dinb(w_dff_B_JW3HweTE7_1),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n232),.clk(gclk));
	jnot g0169(.din(w_n232_0[1]),.dout(n233),.clk(gclk));
	jor g0170(.dina(w_n221_0[0]),.dinb(w_n194_0[1]),.dout(n234),.clk(gclk));
	jxor g0171(.dina(w_n220_0[0]),.dinb(w_n194_0[0]),.dout(n235),.clk(gclk));
	jor g0172(.dina(n235),.dinb(w_n189_0[0]),.dout(n236),.clk(gclk));
	jand g0173(.dina(n236),.dinb(n234),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n238),.clk(gclk));
	jnot g0175(.din(n238),.dout(n239),.clk(gclk));
	jand g0176(.dina(w_n218_0[0]),.dinb(w_n199_0[0]),.dout(n240),.clk(gclk));
	jand g0177(.dina(w_n219_0[0]),.dinb(w_n196_0[0]),.dout(n241),.clk(gclk));
	jor g0178(.dina(n241),.dinb(n240),.dout(n242),.clk(gclk));
	jand g0179(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(n243),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_n216_0[0]),.dinb(w_n204_0[0]),.dout(n245),.clk(gclk));
	jand g0182(.dina(w_n217_0[0]),.dinb(w_n201_0[0]),.dout(n246),.clk(gclk));
	jor g0183(.dina(n246),.dinb(n245),.dout(n247),.clk(gclk));
	jand g0184(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n248),.clk(gclk));
	jnot g0185(.din(n248),.dout(n249),.clk(gclk));
	jnot g0186(.din(w_n213_0[0]),.dout(n250),.clk(gclk));
	jand g0187(.dina(w_n215_0[0]),.dinb(w_n206_0[0]),.dout(n251),.clk(gclk));
	jor g0188(.dina(n251),.dinb(n250),.dout(n252),.clk(gclk));
	jand g0189(.dina(w_G307gat_6[0]),.dinb(w_G86gat_6[2]),.dout(n253),.clk(gclk));
	jnot g0190(.din(n253),.dout(n254),.clk(gclk));
	jand g0191(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n255),.clk(gclk));
	jor g0192(.dina(w_n255_0[1]),.dinb(w_n209_0[0]),.dout(n256),.clk(gclk));
	jand g0193(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n257),.clk(gclk));
	jand g0194(.dina(w_n257_0[1]),.dinb(w_n207_0[0]),.dout(n258),.clk(gclk));
	jnot g0195(.din(w_n258_0[2]),.dout(n259),.clk(gclk));
	jand g0196(.dina(w_n259_0[1]),.dinb(n256),.dout(n260),.clk(gclk));
	jor g0197(.dina(n260),.dinb(w_n210_0[2]),.dout(n261),.clk(gclk));
	jand g0198(.dina(w_n259_0[0]),.dinb(w_n210_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(n262),.dout(n263),.clk(gclk));
	jand g0200(.dina(n263),.dinb(w_n261_0[1]),.dout(n264),.clk(gclk));
	jxor g0201(.dina(w_n264_0[1]),.dinb(w_n254_0[1]),.dout(n265),.clk(gclk));
	jxor g0202(.dina(w_n265_0[1]),.dinb(w_n252_0[1]),.dout(n266),.clk(gclk));
	jxor g0203(.dina(w_n266_0[1]),.dinb(w_n249_0[1]),.dout(n267),.clk(gclk));
	jxor g0204(.dina(w_n267_0[1]),.dinb(w_n247_0[1]),.dout(n268),.clk(gclk));
	jxor g0205(.dina(w_n268_0[1]),.dinb(w_n244_0[1]),.dout(n269),.clk(gclk));
	jxor g0206(.dina(w_n269_0[1]),.dinb(w_n242_0[1]),.dout(n270),.clk(gclk));
	jxor g0207(.dina(w_n270_0[1]),.dinb(w_n239_0[1]),.dout(n271),.clk(gclk));
	jnot g0208(.din(w_n271_0[1]),.dout(n272),.clk(gclk));
	jxor g0209(.dina(w_n272_0[1]),.dinb(w_n237_0[2]),.dout(n273),.clk(gclk));
	jxor g0210(.dina(n273),.dinb(n233),.dout(n274),.clk(gclk));
	jxor g0211(.dina(w_n274_0[1]),.dinb(w_n231_0[1]),.dout(n275),.clk(gclk));
	jxor g0212(.dina(w_n275_0[1]),.dinb(w_dff_B_4L0Rtspp9_1),.dout(w_dff_A_oHiEz1mj9_2),.clk(gclk));
	jand g0213(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n277),.clk(gclk));
	jnot g0214(.din(w_n277_0[1]),.dout(n278),.clk(gclk));
	jnot g0215(.din(w_n274_0[0]),.dout(n279),.clk(gclk));
	jor g0216(.dina(n279),.dinb(w_n231_0[0]),.dout(n280),.clk(gclk));
	jor g0217(.dina(w_n275_0[0]),.dinb(w_n226_0[0]),.dout(n281),.clk(gclk));
	jand g0218(.dina(n281),.dinb(w_dff_B_44uZDAnU6_1),.dout(n282),.clk(gclk));
	jand g0219(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(w_n283_0[1]),.dout(n284),.clk(gclk));
	jor g0221(.dina(w_n272_0[0]),.dinb(w_n237_0[1]),.dout(n285),.clk(gclk));
	jxor g0222(.dina(w_n271_0[0]),.dinb(w_n237_0[0]),.dout(n286),.clk(gclk));
	jor g0223(.dina(n286),.dinb(w_n232_0[0]),.dout(n287),.clk(gclk));
	jand g0224(.dina(n287),.dinb(n285),.dout(n288),.clk(gclk));
	jand g0225(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n289),.clk(gclk));
	jnot g0226(.din(n289),.dout(n290),.clk(gclk));
	jand g0227(.dina(w_n269_0[0]),.dinb(w_n242_0[0]),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n270_0[0]),.dinb(w_n239_0[0]),.dout(n292),.clk(gclk));
	jor g0229(.dina(n292),.dinb(n291),.dout(n293),.clk(gclk));
	jand g0230(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_n267_0[0]),.dinb(w_n247_0[0]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n268_0[0]),.dinb(w_n244_0[0]),.dout(n297),.clk(gclk));
	jor g0234(.dina(n297),.dinb(n296),.dout(n298),.clk(gclk));
	jand g0235(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n299),.clk(gclk));
	jnot g0236(.din(n299),.dout(n300),.clk(gclk));
	jand g0237(.dina(w_n265_0[0]),.dinb(w_n252_0[0]),.dout(n301),.clk(gclk));
	jand g0238(.dina(w_n266_0[0]),.dinb(w_n249_0[0]),.dout(n302),.clk(gclk));
	jor g0239(.dina(n302),.dinb(n301),.dout(n303),.clk(gclk));
	jand g0240(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n304),.clk(gclk));
	jnot g0241(.din(n304),.dout(n305),.clk(gclk));
	jnot g0242(.din(w_n261_0[0]),.dout(n306),.clk(gclk));
	jand g0243(.dina(w_n264_0[0]),.dinb(w_n254_0[0]),.dout(n307),.clk(gclk));
	jor g0244(.dina(n307),.dinb(n306),.dout(n308),.clk(gclk));
	jand g0245(.dina(w_G307gat_5[2]),.dinb(w_G103gat_6[2]),.dout(n309),.clk(gclk));
	jnot g0246(.din(n309),.dout(n310),.clk(gclk));
	jand g0247(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n311),.clk(gclk));
	jor g0248(.dina(w_n311_0[1]),.dinb(w_n257_0[0]),.dout(n312),.clk(gclk));
	jand g0249(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n313),.clk(gclk));
	jand g0250(.dina(w_n313_0[1]),.dinb(w_n255_0[0]),.dout(n314),.clk(gclk));
	jnot g0251(.din(w_n314_0[2]),.dout(n315),.clk(gclk));
	jand g0252(.dina(w_n315_0[1]),.dinb(n312),.dout(n316),.clk(gclk));
	jor g0253(.dina(n316),.dinb(w_n258_0[1]),.dout(n317),.clk(gclk));
	jand g0254(.dina(w_n315_0[0]),.dinb(w_n258_0[0]),.dout(n318),.clk(gclk));
	jnot g0255(.din(n318),.dout(n319),.clk(gclk));
	jand g0256(.dina(n319),.dinb(w_n317_0[1]),.dout(n320),.clk(gclk));
	jxor g0257(.dina(w_n320_0[1]),.dinb(w_n310_0[1]),.dout(n321),.clk(gclk));
	jxor g0258(.dina(w_n321_0[1]),.dinb(w_n308_0[1]),.dout(n322),.clk(gclk));
	jxor g0259(.dina(w_n322_0[1]),.dinb(w_n305_0[1]),.dout(n323),.clk(gclk));
	jxor g0260(.dina(w_n323_0[1]),.dinb(w_n303_0[1]),.dout(n324),.clk(gclk));
	jxor g0261(.dina(w_n324_0[1]),.dinb(w_n300_0[1]),.dout(n325),.clk(gclk));
	jxor g0262(.dina(w_n325_0[1]),.dinb(w_n298_0[1]),.dout(n326),.clk(gclk));
	jxor g0263(.dina(w_n326_0[1]),.dinb(w_n295_0[1]),.dout(n327),.clk(gclk));
	jxor g0264(.dina(w_n327_0[1]),.dinb(w_n293_0[1]),.dout(n328),.clk(gclk));
	jxor g0265(.dina(w_n328_0[1]),.dinb(w_n290_0[1]),.dout(n329),.clk(gclk));
	jnot g0266(.din(w_n329_0[1]),.dout(n330),.clk(gclk));
	jxor g0267(.dina(w_n330_0[1]),.dinb(w_n288_0[2]),.dout(n331),.clk(gclk));
	jxor g0268(.dina(n331),.dinb(n284),.dout(n332),.clk(gclk));
	jxor g0269(.dina(w_n332_0[1]),.dinb(w_n282_0[1]),.dout(n333),.clk(gclk));
	jxor g0270(.dina(w_n333_0[1]),.dinb(w_dff_B_kbrQWFFZ8_1),.dout(w_dff_A_Rbm3HLMi5_2),.clk(gclk));
	jand g0271(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n335),.clk(gclk));
	jnot g0272(.din(w_n335_0[1]),.dout(n336),.clk(gclk));
	jnot g0273(.din(w_n332_0[0]),.dout(n337),.clk(gclk));
	jor g0274(.dina(n337),.dinb(w_n282_0[0]),.dout(n338),.clk(gclk));
	jor g0275(.dina(w_n333_0[0]),.dinb(w_n277_0[0]),.dout(n339),.clk(gclk));
	jand g0276(.dina(n339),.dinb(w_dff_B_mzf3UAuW1_1),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n341),.clk(gclk));
	jnot g0278(.din(w_n341_0[1]),.dout(n342),.clk(gclk));
	jor g0279(.dina(w_n330_0[0]),.dinb(w_n288_0[1]),.dout(n343),.clk(gclk));
	jxor g0280(.dina(w_n329_0[0]),.dinb(w_n288_0[0]),.dout(n344),.clk(gclk));
	jor g0281(.dina(n344),.dinb(w_n283_0[0]),.dout(n345),.clk(gclk));
	jand g0282(.dina(n345),.dinb(n343),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n347),.clk(gclk));
	jnot g0284(.din(n347),.dout(n348),.clk(gclk));
	jand g0285(.dina(w_n327_0[0]),.dinb(w_n293_0[0]),.dout(n349),.clk(gclk));
	jand g0286(.dina(w_n328_0[0]),.dinb(w_n290_0[0]),.dout(n350),.clk(gclk));
	jor g0287(.dina(n350),.dinb(n349),.dout(n351),.clk(gclk));
	jand g0288(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n352),.clk(gclk));
	jnot g0289(.din(n352),.dout(n353),.clk(gclk));
	jand g0290(.dina(w_n325_0[0]),.dinb(w_n298_0[0]),.dout(n354),.clk(gclk));
	jand g0291(.dina(w_n326_0[0]),.dinb(w_n295_0[0]),.dout(n355),.clk(gclk));
	jor g0292(.dina(n355),.dinb(n354),.dout(n356),.clk(gclk));
	jand g0293(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n357),.clk(gclk));
	jnot g0294(.din(n357),.dout(n358),.clk(gclk));
	jand g0295(.dina(w_n323_0[0]),.dinb(w_n303_0[0]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_n324_0[0]),.dinb(w_n300_0[0]),.dout(n360),.clk(gclk));
	jor g0297(.dina(n360),.dinb(n359),.dout(n361),.clk(gclk));
	jand g0298(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n362),.clk(gclk));
	jnot g0299(.din(n362),.dout(n363),.clk(gclk));
	jand g0300(.dina(w_n321_0[0]),.dinb(w_n308_0[0]),.dout(n364),.clk(gclk));
	jand g0301(.dina(w_n322_0[0]),.dinb(w_n305_0[0]),.dout(n365),.clk(gclk));
	jor g0302(.dina(n365),.dinb(n364),.dout(n366),.clk(gclk));
	jand g0303(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n367),.clk(gclk));
	jnot g0304(.din(n367),.dout(n368),.clk(gclk));
	jnot g0305(.din(w_n317_0[0]),.dout(n369),.clk(gclk));
	jand g0306(.dina(w_n320_0[0]),.dinb(w_n310_0[0]),.dout(n370),.clk(gclk));
	jor g0307(.dina(n370),.dinb(n369),.dout(n371),.clk(gclk));
	jand g0308(.dina(w_G307gat_5[1]),.dinb(w_G120gat_6[2]),.dout(n372),.clk(gclk));
	jand g0309(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n373),.clk(gclk));
	jor g0310(.dina(w_n373_0[1]),.dinb(w_n313_0[0]),.dout(n374),.clk(gclk));
	jand g0311(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n375),.clk(gclk));
	jand g0312(.dina(w_n375_0[1]),.dinb(w_n311_0[0]),.dout(n376),.clk(gclk));
	jnot g0313(.din(w_n376_0[2]),.dout(n377),.clk(gclk));
	jand g0314(.dina(w_n377_0[1]),.dinb(n374),.dout(n378),.clk(gclk));
	jor g0315(.dina(n378),.dinb(w_n314_0[1]),.dout(n379),.clk(gclk));
	jnot g0316(.din(n379),.dout(n380),.clk(gclk));
	jand g0317(.dina(w_n377_0[0]),.dinb(w_n314_0[0]),.dout(n381),.clk(gclk));
	jor g0318(.dina(n381),.dinb(w_n380_0[1]),.dout(n382),.clk(gclk));
	jxor g0319(.dina(w_n382_0[1]),.dinb(w_n372_0[1]),.dout(n383),.clk(gclk));
	jxor g0320(.dina(w_n383_0[1]),.dinb(w_n371_0[1]),.dout(n384),.clk(gclk));
	jxor g0321(.dina(w_n384_0[1]),.dinb(w_n368_0[1]),.dout(n385),.clk(gclk));
	jxor g0322(.dina(w_n385_0[1]),.dinb(w_n366_0[1]),.dout(n386),.clk(gclk));
	jxor g0323(.dina(w_n386_0[1]),.dinb(w_n363_0[1]),.dout(n387),.clk(gclk));
	jxor g0324(.dina(w_n387_0[1]),.dinb(w_n361_0[1]),.dout(n388),.clk(gclk));
	jxor g0325(.dina(w_n388_0[1]),.dinb(w_n358_0[1]),.dout(n389),.clk(gclk));
	jxor g0326(.dina(w_n389_0[1]),.dinb(w_n356_0[1]),.dout(n390),.clk(gclk));
	jxor g0327(.dina(w_n390_0[1]),.dinb(w_n353_0[1]),.dout(n391),.clk(gclk));
	jxor g0328(.dina(w_n391_0[1]),.dinb(w_n351_0[1]),.dout(n392),.clk(gclk));
	jxor g0329(.dina(w_n392_0[1]),.dinb(w_n348_0[1]),.dout(n393),.clk(gclk));
	jnot g0330(.din(w_n393_0[1]),.dout(n394),.clk(gclk));
	jxor g0331(.dina(w_n394_0[1]),.dinb(w_n346_0[2]),.dout(n395),.clk(gclk));
	jxor g0332(.dina(n395),.dinb(n342),.dout(n396),.clk(gclk));
	jxor g0333(.dina(w_n396_0[1]),.dinb(w_n340_0[1]),.dout(n397),.clk(gclk));
	jxor g0334(.dina(w_n397_0[1]),.dinb(w_dff_B_ij0Oc1JR6_1),.dout(w_dff_A_nwOyaoey4_2),.clk(gclk));
	jand g0335(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n399),.clk(gclk));
	jnot g0336(.din(w_n399_0[1]),.dout(n400),.clk(gclk));
	jnot g0337(.din(w_n396_0[0]),.dout(n401),.clk(gclk));
	jor g0338(.dina(n401),.dinb(w_n340_0[0]),.dout(n402),.clk(gclk));
	jor g0339(.dina(w_n397_0[0]),.dinb(w_n335_0[0]),.dout(n403),.clk(gclk));
	jand g0340(.dina(n403),.dinb(w_dff_B_APQpbtXG4_1),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n405),.clk(gclk));
	jnot g0342(.din(w_n405_0[1]),.dout(n406),.clk(gclk));
	jor g0343(.dina(w_n394_0[0]),.dinb(w_n346_0[1]),.dout(n407),.clk(gclk));
	jxor g0344(.dina(w_n393_0[0]),.dinb(w_n346_0[0]),.dout(n408),.clk(gclk));
	jor g0345(.dina(n408),.dinb(w_n341_0[0]),.dout(n409),.clk(gclk));
	jand g0346(.dina(n409),.dinb(n407),.dout(n410),.clk(gclk));
	jand g0347(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n411),.clk(gclk));
	jnot g0348(.din(n411),.dout(n412),.clk(gclk));
	jand g0349(.dina(w_n391_0[0]),.dinb(w_n351_0[0]),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n392_0[0]),.dinb(w_n348_0[0]),.dout(n414),.clk(gclk));
	jor g0351(.dina(n414),.dinb(n413),.dout(n415),.clk(gclk));
	jand g0352(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n416),.clk(gclk));
	jnot g0353(.din(n416),.dout(n417),.clk(gclk));
	jand g0354(.dina(w_n389_0[0]),.dinb(w_n356_0[0]),.dout(n418),.clk(gclk));
	jand g0355(.dina(w_n390_0[0]),.dinb(w_n353_0[0]),.dout(n419),.clk(gclk));
	jor g0356(.dina(n419),.dinb(n418),.dout(n420),.clk(gclk));
	jand g0357(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n421),.clk(gclk));
	jnot g0358(.din(n421),.dout(n422),.clk(gclk));
	jand g0359(.dina(w_n387_0[0]),.dinb(w_n361_0[0]),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_n388_0[0]),.dinb(w_n358_0[0]),.dout(n424),.clk(gclk));
	jor g0361(.dina(n424),.dinb(n423),.dout(n425),.clk(gclk));
	jand g0362(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n426),.clk(gclk));
	jnot g0363(.din(n426),.dout(n427),.clk(gclk));
	jand g0364(.dina(w_n385_0[0]),.dinb(w_n366_0[0]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_n386_0[0]),.dinb(w_n363_0[0]),.dout(n429),.clk(gclk));
	jor g0366(.dina(n429),.dinb(n428),.dout(n430),.clk(gclk));
	jand g0367(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n431),.clk(gclk));
	jnot g0368(.din(n431),.dout(n432),.clk(gclk));
	jand g0369(.dina(w_n383_0[0]),.dinb(w_n371_0[0]),.dout(n433),.clk(gclk));
	jand g0370(.dina(w_n384_0[0]),.dinb(w_n368_0[0]),.dout(n434),.clk(gclk));
	jor g0371(.dina(n434),.dinb(n433),.dout(n435),.clk(gclk));
	jand g0372(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n436),.clk(gclk));
	jnot g0373(.din(n436),.dout(n437),.clk(gclk));
	jnot g0374(.din(w_n372_0[0]),.dout(n438),.clk(gclk));
	jnot g0375(.din(w_n382_0[0]),.dout(n439),.clk(gclk));
	jand g0376(.dina(n439),.dinb(n438),.dout(n440),.clk(gclk));
	jor g0377(.dina(n440),.dinb(w_n380_0[0]),.dout(n441),.clk(gclk));
	jand g0378(.dina(w_G307gat_5[0]),.dinb(w_G137gat_6[2]),.dout(n442),.clk(gclk));
	jand g0379(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n443),.clk(gclk));
	jor g0380(.dina(w_n443_0[1]),.dinb(w_n375_0[0]),.dout(n444),.clk(gclk));
	jand g0381(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n445),.clk(gclk));
	jand g0382(.dina(w_n445_0[1]),.dinb(w_n373_0[0]),.dout(n446),.clk(gclk));
	jnot g0383(.din(w_n446_0[2]),.dout(n447),.clk(gclk));
	jand g0384(.dina(w_n447_0[1]),.dinb(n444),.dout(n448),.clk(gclk));
	jor g0385(.dina(n448),.dinb(w_n376_0[1]),.dout(n449),.clk(gclk));
	jnot g0386(.din(n449),.dout(n450),.clk(gclk));
	jand g0387(.dina(w_n447_0[0]),.dinb(w_n376_0[0]),.dout(n451),.clk(gclk));
	jor g0388(.dina(n451),.dinb(w_n450_0[1]),.dout(n452),.clk(gclk));
	jxor g0389(.dina(w_n452_0[1]),.dinb(w_n442_0[1]),.dout(n453),.clk(gclk));
	jxor g0390(.dina(w_n453_0[1]),.dinb(w_n441_0[1]),.dout(n454),.clk(gclk));
	jxor g0391(.dina(w_n454_0[1]),.dinb(w_n437_0[1]),.dout(n455),.clk(gclk));
	jxor g0392(.dina(w_n455_0[1]),.dinb(w_n435_0[1]),.dout(n456),.clk(gclk));
	jxor g0393(.dina(w_n456_0[1]),.dinb(w_n432_0[1]),.dout(n457),.clk(gclk));
	jxor g0394(.dina(w_n457_0[1]),.dinb(w_n430_0[1]),.dout(n458),.clk(gclk));
	jxor g0395(.dina(w_n458_0[1]),.dinb(w_n427_0[1]),.dout(n459),.clk(gclk));
	jxor g0396(.dina(w_n459_0[1]),.dinb(w_n425_0[1]),.dout(n460),.clk(gclk));
	jxor g0397(.dina(w_n460_0[1]),.dinb(w_n422_0[1]),.dout(n461),.clk(gclk));
	jxor g0398(.dina(w_n461_0[1]),.dinb(w_n420_0[1]),.dout(n462),.clk(gclk));
	jxor g0399(.dina(w_n462_0[1]),.dinb(w_n417_0[1]),.dout(n463),.clk(gclk));
	jxor g0400(.dina(w_n463_0[1]),.dinb(w_n415_0[1]),.dout(n464),.clk(gclk));
	jxor g0401(.dina(w_n464_0[1]),.dinb(w_n412_0[1]),.dout(n465),.clk(gclk));
	jnot g0402(.din(w_n465_0[1]),.dout(n466),.clk(gclk));
	jxor g0403(.dina(w_n466_0[1]),.dinb(w_n410_0[2]),.dout(n467),.clk(gclk));
	jxor g0404(.dina(n467),.dinb(n406),.dout(n468),.clk(gclk));
	jxor g0405(.dina(w_n468_0[1]),.dinb(w_n404_0[1]),.dout(n469),.clk(gclk));
	jxor g0406(.dina(w_n469_0[1]),.dinb(w_dff_B_igGtsUuN6_1),.dout(w_dff_A_Vd7i4kR94_2),.clk(gclk));
	jand g0407(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n471),.clk(gclk));
	jnot g0408(.din(w_n471_0[1]),.dout(n472),.clk(gclk));
	jnot g0409(.din(w_n468_0[0]),.dout(n473),.clk(gclk));
	jor g0410(.dina(n473),.dinb(w_n404_0[0]),.dout(n474),.clk(gclk));
	jor g0411(.dina(w_n469_0[0]),.dinb(w_n399_0[0]),.dout(n475),.clk(gclk));
	jand g0412(.dina(n475),.dinb(w_dff_B_GX6DC5BQ6_1),.dout(n476),.clk(gclk));
	jand g0413(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n477),.clk(gclk));
	jnot g0414(.din(w_n477_0[1]),.dout(n478),.clk(gclk));
	jor g0415(.dina(w_n466_0[0]),.dinb(w_n410_0[1]),.dout(n479),.clk(gclk));
	jxor g0416(.dina(w_n465_0[0]),.dinb(w_n410_0[0]),.dout(n480),.clk(gclk));
	jor g0417(.dina(n480),.dinb(w_n405_0[0]),.dout(n481),.clk(gclk));
	jand g0418(.dina(n481),.dinb(n479),.dout(n482),.clk(gclk));
	jand g0419(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n463_0[0]),.dinb(w_n415_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n464_0[0]),.dinb(w_n412_0[0]),.dout(n486),.clk(gclk));
	jor g0423(.dina(n486),.dinb(n485),.dout(n487),.clk(gclk));
	jand g0424(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n461_0[0]),.dinb(w_n420_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n462_0[0]),.dinb(w_n417_0[0]),.dout(n491),.clk(gclk));
	jor g0428(.dina(n491),.dinb(n490),.dout(n492),.clk(gclk));
	jand g0429(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jand g0431(.dina(w_n459_0[0]),.dinb(w_n425_0[0]),.dout(n495),.clk(gclk));
	jand g0432(.dina(w_n460_0[0]),.dinb(w_n422_0[0]),.dout(n496),.clk(gclk));
	jor g0433(.dina(n496),.dinb(n495),.dout(n497),.clk(gclk));
	jand g0434(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_n457_0[0]),.dinb(w_n430_0[0]),.dout(n500),.clk(gclk));
	jand g0437(.dina(w_n458_0[0]),.dinb(w_n427_0[0]),.dout(n501),.clk(gclk));
	jor g0438(.dina(n501),.dinb(n500),.dout(n502),.clk(gclk));
	jand g0439(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n503),.clk(gclk));
	jnot g0440(.din(n503),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_n455_0[0]),.dinb(w_n435_0[0]),.dout(n505),.clk(gclk));
	jand g0442(.dina(w_n456_0[0]),.dinb(w_n432_0[0]),.dout(n506),.clk(gclk));
	jor g0443(.dina(n506),.dinb(n505),.dout(n507),.clk(gclk));
	jand g0444(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n508),.clk(gclk));
	jnot g0445(.din(n508),.dout(n509),.clk(gclk));
	jand g0446(.dina(w_n453_0[0]),.dinb(w_n441_0[0]),.dout(n510),.clk(gclk));
	jand g0447(.dina(w_n454_0[0]),.dinb(w_n437_0[0]),.dout(n511),.clk(gclk));
	jor g0448(.dina(n511),.dinb(n510),.dout(n512),.clk(gclk));
	jand g0449(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n513),.clk(gclk));
	jnot g0450(.din(n513),.dout(n514),.clk(gclk));
	jnot g0451(.din(w_n442_0[0]),.dout(n515),.clk(gclk));
	jnot g0452(.din(w_n452_0[0]),.dout(n516),.clk(gclk));
	jand g0453(.dina(n516),.dinb(n515),.dout(n517),.clk(gclk));
	jor g0454(.dina(n517),.dinb(w_n450_0[0]),.dout(n518),.clk(gclk));
	jand g0455(.dina(w_G307gat_4[2]),.dinb(w_G154gat_6[2]),.dout(n519),.clk(gclk));
	jand g0456(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n520),.clk(gclk));
	jor g0457(.dina(w_n520_0[1]),.dinb(w_n445_0[0]),.dout(n521),.clk(gclk));
	jand g0458(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n522),.clk(gclk));
	jand g0459(.dina(w_n522_0[1]),.dinb(w_n443_0[0]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[2]),.dout(n524),.clk(gclk));
	jand g0461(.dina(w_n524_0[1]),.dinb(n521),.dout(n525),.clk(gclk));
	jor g0462(.dina(n525),.dinb(w_n446_0[1]),.dout(n526),.clk(gclk));
	jnot g0463(.din(n526),.dout(n527),.clk(gclk));
	jand g0464(.dina(w_n524_0[0]),.dinb(w_n446_0[0]),.dout(n528),.clk(gclk));
	jor g0465(.dina(n528),.dinb(w_n527_0[1]),.dout(n529),.clk(gclk));
	jxor g0466(.dina(w_n529_0[1]),.dinb(w_n519_0[1]),.dout(n530),.clk(gclk));
	jxor g0467(.dina(w_n530_0[1]),.dinb(w_n518_0[1]),.dout(n531),.clk(gclk));
	jxor g0468(.dina(w_n531_0[1]),.dinb(w_n514_0[1]),.dout(n532),.clk(gclk));
	jxor g0469(.dina(w_n532_0[1]),.dinb(w_n512_0[1]),.dout(n533),.clk(gclk));
	jxor g0470(.dina(w_n533_0[1]),.dinb(w_n509_0[1]),.dout(n534),.clk(gclk));
	jxor g0471(.dina(w_n534_0[1]),.dinb(w_n507_0[1]),.dout(n535),.clk(gclk));
	jxor g0472(.dina(w_n535_0[1]),.dinb(w_n504_0[1]),.dout(n536),.clk(gclk));
	jxor g0473(.dina(w_n536_0[1]),.dinb(w_n502_0[1]),.dout(n537),.clk(gclk));
	jxor g0474(.dina(w_n537_0[1]),.dinb(w_n499_0[1]),.dout(n538),.clk(gclk));
	jxor g0475(.dina(w_n538_0[1]),.dinb(w_n497_0[1]),.dout(n539),.clk(gclk));
	jxor g0476(.dina(w_n539_0[1]),.dinb(w_n494_0[1]),.dout(n540),.clk(gclk));
	jxor g0477(.dina(w_n540_0[1]),.dinb(w_n492_0[1]),.dout(n541),.clk(gclk));
	jxor g0478(.dina(w_n541_0[1]),.dinb(w_n489_0[1]),.dout(n542),.clk(gclk));
	jxor g0479(.dina(w_n542_0[1]),.dinb(w_n487_0[1]),.dout(n543),.clk(gclk));
	jxor g0480(.dina(w_n543_0[1]),.dinb(w_n484_0[1]),.dout(n544),.clk(gclk));
	jnot g0481(.din(w_n544_0[1]),.dout(n545),.clk(gclk));
	jxor g0482(.dina(w_n545_0[1]),.dinb(w_n482_0[2]),.dout(n546),.clk(gclk));
	jxor g0483(.dina(n546),.dinb(n478),.dout(n547),.clk(gclk));
	jxor g0484(.dina(w_n547_0[1]),.dinb(w_n476_0[1]),.dout(n548),.clk(gclk));
	jxor g0485(.dina(w_n548_0[1]),.dinb(w_dff_B_pkyARCTV1_1),.dout(w_dff_A_guWKCtIU7_2),.clk(gclk));
	jand g0486(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n550),.clk(gclk));
	jnot g0487(.din(w_n550_0[1]),.dout(n551),.clk(gclk));
	jnot g0488(.din(w_n547_0[0]),.dout(n552),.clk(gclk));
	jor g0489(.dina(n552),.dinb(w_n476_0[0]),.dout(n553),.clk(gclk));
	jor g0490(.dina(w_n548_0[0]),.dinb(w_n471_0[0]),.dout(n554),.clk(gclk));
	jand g0491(.dina(n554),.dinb(w_dff_B_oci1c3qe0_1),.dout(n555),.clk(gclk));
	jand g0492(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n556),.clk(gclk));
	jnot g0493(.din(w_n556_0[1]),.dout(n557),.clk(gclk));
	jor g0494(.dina(w_n545_0[0]),.dinb(w_n482_0[1]),.dout(n558),.clk(gclk));
	jxor g0495(.dina(w_n544_0[0]),.dinb(w_n482_0[0]),.dout(n559),.clk(gclk));
	jor g0496(.dina(n559),.dinb(w_n477_0[0]),.dout(n560),.clk(gclk));
	jand g0497(.dina(n560),.dinb(n558),.dout(n561),.clk(gclk));
	jand g0498(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n562),.clk(gclk));
	jnot g0499(.din(n562),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n542_0[0]),.dinb(w_n487_0[0]),.dout(n564),.clk(gclk));
	jand g0501(.dina(w_n543_0[0]),.dinb(w_n484_0[0]),.dout(n565),.clk(gclk));
	jor g0502(.dina(n565),.dinb(n564),.dout(n566),.clk(gclk));
	jand g0503(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n567),.clk(gclk));
	jnot g0504(.din(n567),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n540_0[0]),.dinb(w_n492_0[0]),.dout(n569),.clk(gclk));
	jand g0506(.dina(w_n541_0[0]),.dinb(w_n489_0[0]),.dout(n570),.clk(gclk));
	jor g0507(.dina(n570),.dinb(n569),.dout(n571),.clk(gclk));
	jand g0508(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n572),.clk(gclk));
	jnot g0509(.din(n572),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n538_0[0]),.dinb(w_n497_0[0]),.dout(n574),.clk(gclk));
	jand g0511(.dina(w_n539_0[0]),.dinb(w_n494_0[0]),.dout(n575),.clk(gclk));
	jor g0512(.dina(n575),.dinb(n574),.dout(n576),.clk(gclk));
	jand g0513(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n577),.clk(gclk));
	jnot g0514(.din(n577),.dout(n578),.clk(gclk));
	jand g0515(.dina(w_n536_0[0]),.dinb(w_n502_0[0]),.dout(n579),.clk(gclk));
	jand g0516(.dina(w_n537_0[0]),.dinb(w_n499_0[0]),.dout(n580),.clk(gclk));
	jor g0517(.dina(n580),.dinb(n579),.dout(n581),.clk(gclk));
	jand g0518(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n582),.clk(gclk));
	jnot g0519(.din(n582),.dout(n583),.clk(gclk));
	jand g0520(.dina(w_n534_0[0]),.dinb(w_n507_0[0]),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_n535_0[0]),.dinb(w_n504_0[0]),.dout(n585),.clk(gclk));
	jor g0522(.dina(n585),.dinb(n584),.dout(n586),.clk(gclk));
	jand g0523(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n587),.clk(gclk));
	jnot g0524(.din(n587),.dout(n588),.clk(gclk));
	jand g0525(.dina(w_n532_0[0]),.dinb(w_n512_0[0]),.dout(n589),.clk(gclk));
	jand g0526(.dina(w_n533_0[0]),.dinb(w_n509_0[0]),.dout(n590),.clk(gclk));
	jor g0527(.dina(n590),.dinb(n589),.dout(n591),.clk(gclk));
	jand g0528(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n592),.clk(gclk));
	jnot g0529(.din(n592),.dout(n593),.clk(gclk));
	jand g0530(.dina(w_n530_0[0]),.dinb(w_n518_0[0]),.dout(n594),.clk(gclk));
	jand g0531(.dina(w_n531_0[0]),.dinb(w_n514_0[0]),.dout(n595),.clk(gclk));
	jor g0532(.dina(n595),.dinb(n594),.dout(n596),.clk(gclk));
	jand g0533(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n597),.clk(gclk));
	jnot g0534(.din(n597),.dout(n598),.clk(gclk));
	jnot g0535(.din(w_n519_0[0]),.dout(n599),.clk(gclk));
	jnot g0536(.din(w_n529_0[0]),.dout(n600),.clk(gclk));
	jand g0537(.dina(n600),.dinb(n599),.dout(n601),.clk(gclk));
	jor g0538(.dina(n601),.dinb(w_n527_0[0]),.dout(n602),.clk(gclk));
	jand g0539(.dina(w_G307gat_4[1]),.dinb(w_G171gat_6[2]),.dout(n603),.clk(gclk));
	jand g0540(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n604),.clk(gclk));
	jor g0541(.dina(w_n604_0[1]),.dinb(w_n522_0[0]),.dout(n605),.clk(gclk));
	jand g0542(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n606),.clk(gclk));
	jand g0543(.dina(w_n606_0[1]),.dinb(w_n520_0[0]),.dout(n607),.clk(gclk));
	jnot g0544(.din(w_n607_0[2]),.dout(n608),.clk(gclk));
	jand g0545(.dina(w_n608_0[1]),.dinb(n605),.dout(n609),.clk(gclk));
	jor g0546(.dina(n609),.dinb(w_n523_0[1]),.dout(n610),.clk(gclk));
	jnot g0547(.din(n610),.dout(n611),.clk(gclk));
	jand g0548(.dina(w_n608_0[0]),.dinb(w_n523_0[0]),.dout(n612),.clk(gclk));
	jor g0549(.dina(n612),.dinb(w_n611_0[1]),.dout(n613),.clk(gclk));
	jxor g0550(.dina(w_n613_0[1]),.dinb(w_n603_0[1]),.dout(n614),.clk(gclk));
	jxor g0551(.dina(w_n614_0[1]),.dinb(w_n602_0[1]),.dout(n615),.clk(gclk));
	jxor g0552(.dina(w_n615_0[1]),.dinb(w_n598_0[1]),.dout(n616),.clk(gclk));
	jxor g0553(.dina(w_n616_0[1]),.dinb(w_n596_0[1]),.dout(n617),.clk(gclk));
	jxor g0554(.dina(w_n617_0[1]),.dinb(w_n593_0[1]),.dout(n618),.clk(gclk));
	jxor g0555(.dina(w_n618_0[1]),.dinb(w_n591_0[1]),.dout(n619),.clk(gclk));
	jxor g0556(.dina(w_n619_0[1]),.dinb(w_n588_0[1]),.dout(n620),.clk(gclk));
	jxor g0557(.dina(w_n620_0[1]),.dinb(w_n586_0[1]),.dout(n621),.clk(gclk));
	jxor g0558(.dina(w_n621_0[1]),.dinb(w_n583_0[1]),.dout(n622),.clk(gclk));
	jxor g0559(.dina(w_n622_0[1]),.dinb(w_n581_0[1]),.dout(n623),.clk(gclk));
	jxor g0560(.dina(w_n623_0[1]),.dinb(w_n578_0[1]),.dout(n624),.clk(gclk));
	jxor g0561(.dina(w_n624_0[1]),.dinb(w_n576_0[1]),.dout(n625),.clk(gclk));
	jxor g0562(.dina(w_n625_0[1]),.dinb(w_n573_0[1]),.dout(n626),.clk(gclk));
	jxor g0563(.dina(w_n626_0[1]),.dinb(w_n571_0[1]),.dout(n627),.clk(gclk));
	jxor g0564(.dina(w_n627_0[1]),.dinb(w_n568_0[1]),.dout(n628),.clk(gclk));
	jxor g0565(.dina(w_n628_0[1]),.dinb(w_n566_0[1]),.dout(n629),.clk(gclk));
	jxor g0566(.dina(w_n629_0[1]),.dinb(w_n563_0[1]),.dout(n630),.clk(gclk));
	jnot g0567(.din(w_n630_0[1]),.dout(n631),.clk(gclk));
	jxor g0568(.dina(w_n631_0[1]),.dinb(w_n561_0[2]),.dout(n632),.clk(gclk));
	jxor g0569(.dina(n632),.dinb(n557),.dout(n633),.clk(gclk));
	jxor g0570(.dina(w_n633_0[1]),.dinb(w_n555_0[1]),.dout(n634),.clk(gclk));
	jxor g0571(.dina(w_n634_0[1]),.dinb(w_dff_B_TVXLodJF2_1),.dout(w_dff_A_8K6sinQo2_2),.clk(gclk));
	jand g0572(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n636),.clk(gclk));
	jnot g0573(.din(w_n636_0[1]),.dout(n637),.clk(gclk));
	jnot g0574(.din(w_n633_0[0]),.dout(n638),.clk(gclk));
	jor g0575(.dina(n638),.dinb(w_n555_0[0]),.dout(n639),.clk(gclk));
	jor g0576(.dina(w_n634_0[0]),.dinb(w_n550_0[0]),.dout(n640),.clk(gclk));
	jand g0577(.dina(n640),.dinb(w_dff_B_PH0q2cYe9_1),.dout(n641),.clk(gclk));
	jand g0578(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n642),.clk(gclk));
	jnot g0579(.din(w_n642_0[1]),.dout(n643),.clk(gclk));
	jor g0580(.dina(w_n631_0[0]),.dinb(w_n561_0[1]),.dout(n644),.clk(gclk));
	jxor g0581(.dina(w_n630_0[0]),.dinb(w_n561_0[0]),.dout(n645),.clk(gclk));
	jor g0582(.dina(n645),.dinb(w_n556_0[0]),.dout(n646),.clk(gclk));
	jand g0583(.dina(n646),.dinb(n644),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n648),.clk(gclk));
	jnot g0585(.din(n648),.dout(n649),.clk(gclk));
	jand g0586(.dina(w_n628_0[0]),.dinb(w_n566_0[0]),.dout(n650),.clk(gclk));
	jand g0587(.dina(w_n629_0[0]),.dinb(w_n563_0[0]),.dout(n651),.clk(gclk));
	jor g0588(.dina(n651),.dinb(n650),.dout(n652),.clk(gclk));
	jand g0589(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n653),.clk(gclk));
	jnot g0590(.din(n653),.dout(n654),.clk(gclk));
	jand g0591(.dina(w_n626_0[0]),.dinb(w_n571_0[0]),.dout(n655),.clk(gclk));
	jand g0592(.dina(w_n627_0[0]),.dinb(w_n568_0[0]),.dout(n656),.clk(gclk));
	jor g0593(.dina(n656),.dinb(n655),.dout(n657),.clk(gclk));
	jand g0594(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n658),.clk(gclk));
	jnot g0595(.din(n658),.dout(n659),.clk(gclk));
	jand g0596(.dina(w_n624_0[0]),.dinb(w_n576_0[0]),.dout(n660),.clk(gclk));
	jand g0597(.dina(w_n625_0[0]),.dinb(w_n573_0[0]),.dout(n661),.clk(gclk));
	jor g0598(.dina(n661),.dinb(n660),.dout(n662),.clk(gclk));
	jand g0599(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n663),.clk(gclk));
	jnot g0600(.din(n663),.dout(n664),.clk(gclk));
	jand g0601(.dina(w_n622_0[0]),.dinb(w_n581_0[0]),.dout(n665),.clk(gclk));
	jand g0602(.dina(w_n623_0[0]),.dinb(w_n578_0[0]),.dout(n666),.clk(gclk));
	jor g0603(.dina(n666),.dinb(n665),.dout(n667),.clk(gclk));
	jand g0604(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n668),.clk(gclk));
	jnot g0605(.din(n668),.dout(n669),.clk(gclk));
	jand g0606(.dina(w_n620_0[0]),.dinb(w_n586_0[0]),.dout(n670),.clk(gclk));
	jand g0607(.dina(w_n621_0[0]),.dinb(w_n583_0[0]),.dout(n671),.clk(gclk));
	jor g0608(.dina(n671),.dinb(n670),.dout(n672),.clk(gclk));
	jand g0609(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_n618_0[0]),.dinb(w_n591_0[0]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n619_0[0]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jor g0613(.dina(n676),.dinb(n675),.dout(n677),.clk(gclk));
	jand g0614(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n678),.clk(gclk));
	jnot g0615(.din(n678),.dout(n679),.clk(gclk));
	jand g0616(.dina(w_n616_0[0]),.dinb(w_n596_0[0]),.dout(n680),.clk(gclk));
	jand g0617(.dina(w_n617_0[0]),.dinb(w_n593_0[0]),.dout(n681),.clk(gclk));
	jor g0618(.dina(n681),.dinb(n680),.dout(n682),.clk(gclk));
	jand g0619(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n683),.clk(gclk));
	jnot g0620(.din(n683),.dout(n684),.clk(gclk));
	jand g0621(.dina(w_n614_0[0]),.dinb(w_n602_0[0]),.dout(n685),.clk(gclk));
	jand g0622(.dina(w_n615_0[0]),.dinb(w_n598_0[0]),.dout(n686),.clk(gclk));
	jor g0623(.dina(n686),.dinb(n685),.dout(n687),.clk(gclk));
	jand g0624(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n688),.clk(gclk));
	jnot g0625(.din(n688),.dout(n689),.clk(gclk));
	jnot g0626(.din(w_n603_0[0]),.dout(n690),.clk(gclk));
	jnot g0627(.din(w_n613_0[0]),.dout(n691),.clk(gclk));
	jand g0628(.dina(n691),.dinb(n690),.dout(n692),.clk(gclk));
	jor g0629(.dina(n692),.dinb(w_n611_0[0]),.dout(n693),.clk(gclk));
	jand g0630(.dina(w_G307gat_4[0]),.dinb(w_G188gat_6[2]),.dout(n694),.clk(gclk));
	jand g0631(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n695),.clk(gclk));
	jor g0632(.dina(w_n695_0[2]),.dinb(w_n606_0[0]),.dout(n696),.clk(gclk));
	jand g0633(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n697),.clk(gclk));
	jand g0634(.dina(w_n697_0[1]),.dinb(w_n604_0[0]),.dout(n698),.clk(gclk));
	jnot g0635(.din(w_n698_0[2]),.dout(n699),.clk(gclk));
	jand g0636(.dina(w_n699_0[1]),.dinb(n696),.dout(n700),.clk(gclk));
	jor g0637(.dina(n700),.dinb(w_n607_0[1]),.dout(n701),.clk(gclk));
	jnot g0638(.din(n701),.dout(n702),.clk(gclk));
	jand g0639(.dina(w_n699_0[0]),.dinb(w_n607_0[0]),.dout(n703),.clk(gclk));
	jor g0640(.dina(n703),.dinb(w_n702_0[1]),.dout(n704),.clk(gclk));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_n694_0[1]),.dout(n705),.clk(gclk));
	jxor g0642(.dina(w_n705_0[1]),.dinb(w_n693_0[1]),.dout(n706),.clk(gclk));
	jxor g0643(.dina(w_n706_0[1]),.dinb(w_n689_0[1]),.dout(n707),.clk(gclk));
	jxor g0644(.dina(w_n707_0[1]),.dinb(w_n687_0[1]),.dout(n708),.clk(gclk));
	jxor g0645(.dina(w_n708_0[1]),.dinb(w_n684_0[1]),.dout(n709),.clk(gclk));
	jxor g0646(.dina(w_n709_0[1]),.dinb(w_n682_0[1]),.dout(n710),.clk(gclk));
	jxor g0647(.dina(w_n710_0[1]),.dinb(w_n679_0[1]),.dout(n711),.clk(gclk));
	jxor g0648(.dina(w_n711_0[1]),.dinb(w_n677_0[1]),.dout(n712),.clk(gclk));
	jxor g0649(.dina(w_n712_0[1]),.dinb(w_n674_0[1]),.dout(n713),.clk(gclk));
	jxor g0650(.dina(w_n713_0[1]),.dinb(w_n672_0[1]),.dout(n714),.clk(gclk));
	jxor g0651(.dina(w_n714_0[1]),.dinb(w_n669_0[1]),.dout(n715),.clk(gclk));
	jxor g0652(.dina(w_n715_0[1]),.dinb(w_n667_0[1]),.dout(n716),.clk(gclk));
	jxor g0653(.dina(w_n716_0[1]),.dinb(w_n664_0[1]),.dout(n717),.clk(gclk));
	jxor g0654(.dina(w_n717_0[1]),.dinb(w_n662_0[1]),.dout(n718),.clk(gclk));
	jxor g0655(.dina(w_n718_0[1]),.dinb(w_n659_0[1]),.dout(n719),.clk(gclk));
	jxor g0656(.dina(w_n719_0[1]),.dinb(w_n657_0[1]),.dout(n720),.clk(gclk));
	jxor g0657(.dina(w_n720_0[1]),.dinb(w_n654_0[1]),.dout(n721),.clk(gclk));
	jxor g0658(.dina(w_n721_0[1]),.dinb(w_n652_0[1]),.dout(n722),.clk(gclk));
	jxor g0659(.dina(w_n722_0[1]),.dinb(w_n649_0[1]),.dout(n723),.clk(gclk));
	jnot g0660(.din(w_n723_0[1]),.dout(n724),.clk(gclk));
	jxor g0661(.dina(w_n724_0[1]),.dinb(w_n647_0[2]),.dout(n725),.clk(gclk));
	jxor g0662(.dina(n725),.dinb(n643),.dout(n726),.clk(gclk));
	jxor g0663(.dina(w_n726_0[1]),.dinb(w_n641_0[1]),.dout(n727),.clk(gclk));
	jxor g0664(.dina(w_n727_0[1]),.dinb(w_dff_B_leim9mt08_1),.dout(w_dff_A_bgSyLykw2_2),.clk(gclk));
	jand g0665(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n729),.clk(gclk));
	jnot g0666(.din(w_n729_0[1]),.dout(n730),.clk(gclk));
	jnot g0667(.din(w_n726_0[0]),.dout(n731),.clk(gclk));
	jor g0668(.dina(n731),.dinb(w_n641_0[0]),.dout(n732),.clk(gclk));
	jor g0669(.dina(w_n727_0[0]),.dinb(w_n636_0[0]),.dout(n733),.clk(gclk));
	jand g0670(.dina(n733),.dinb(w_dff_B_2un0XYhY5_1),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n735),.clk(gclk));
	jnot g0672(.din(w_n735_0[1]),.dout(n736),.clk(gclk));
	jor g0673(.dina(w_n724_0[0]),.dinb(w_n647_0[1]),.dout(n737),.clk(gclk));
	jxor g0674(.dina(w_n723_0[0]),.dinb(w_n647_0[0]),.dout(n738),.clk(gclk));
	jor g0675(.dina(n738),.dinb(w_n642_0[0]),.dout(n739),.clk(gclk));
	jand g0676(.dina(n739),.dinb(n737),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n741),.clk(gclk));
	jnot g0678(.din(n741),.dout(n742),.clk(gclk));
	jand g0679(.dina(w_n721_0[0]),.dinb(w_n652_0[0]),.dout(n743),.clk(gclk));
	jand g0680(.dina(w_n722_0[0]),.dinb(w_n649_0[0]),.dout(n744),.clk(gclk));
	jor g0681(.dina(n744),.dinb(n743),.dout(n745),.clk(gclk));
	jand g0682(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n746),.clk(gclk));
	jnot g0683(.din(n746),.dout(n747),.clk(gclk));
	jand g0684(.dina(w_n719_0[0]),.dinb(w_n657_0[0]),.dout(n748),.clk(gclk));
	jand g0685(.dina(w_n720_0[0]),.dinb(w_n654_0[0]),.dout(n749),.clk(gclk));
	jor g0686(.dina(n749),.dinb(n748),.dout(n750),.clk(gclk));
	jand g0687(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n751),.clk(gclk));
	jnot g0688(.din(n751),.dout(n752),.clk(gclk));
	jand g0689(.dina(w_n717_0[0]),.dinb(w_n662_0[0]),.dout(n753),.clk(gclk));
	jand g0690(.dina(w_n718_0[0]),.dinb(w_n659_0[0]),.dout(n754),.clk(gclk));
	jor g0691(.dina(n754),.dinb(n753),.dout(n755),.clk(gclk));
	jand g0692(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n756),.clk(gclk));
	jnot g0693(.din(n756),.dout(n757),.clk(gclk));
	jand g0694(.dina(w_n715_0[0]),.dinb(w_n667_0[0]),.dout(n758),.clk(gclk));
	jand g0695(.dina(w_n716_0[0]),.dinb(w_n664_0[0]),.dout(n759),.clk(gclk));
	jor g0696(.dina(n759),.dinb(n758),.dout(n760),.clk(gclk));
	jand g0697(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n761),.clk(gclk));
	jnot g0698(.din(n761),.dout(n762),.clk(gclk));
	jand g0699(.dina(w_n713_0[0]),.dinb(w_n672_0[0]),.dout(n763),.clk(gclk));
	jand g0700(.dina(w_n714_0[0]),.dinb(w_n669_0[0]),.dout(n764),.clk(gclk));
	jor g0701(.dina(n764),.dinb(n763),.dout(n765),.clk(gclk));
	jand g0702(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(w_n711_0[0]),.dinb(w_n677_0[0]),.dout(n768),.clk(gclk));
	jand g0705(.dina(w_n712_0[0]),.dinb(w_n674_0[0]),.dout(n769),.clk(gclk));
	jor g0706(.dina(n769),.dinb(n768),.dout(n770),.clk(gclk));
	jand g0707(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n771),.clk(gclk));
	jnot g0708(.din(n771),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n709_0[0]),.dinb(w_n682_0[0]),.dout(n773),.clk(gclk));
	jand g0710(.dina(w_n710_0[0]),.dinb(w_n679_0[0]),.dout(n774),.clk(gclk));
	jor g0711(.dina(n774),.dinb(n773),.dout(n775),.clk(gclk));
	jand g0712(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n776),.clk(gclk));
	jnot g0713(.din(n776),.dout(n777),.clk(gclk));
	jand g0714(.dina(w_n707_0[0]),.dinb(w_n687_0[0]),.dout(n778),.clk(gclk));
	jand g0715(.dina(w_n708_0[0]),.dinb(w_n684_0[0]),.dout(n779),.clk(gclk));
	jor g0716(.dina(n779),.dinb(n778),.dout(n780),.clk(gclk));
	jand g0717(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n781),.clk(gclk));
	jnot g0718(.din(n781),.dout(n782),.clk(gclk));
	jand g0719(.dina(w_n705_0[0]),.dinb(w_n693_0[0]),.dout(n783),.clk(gclk));
	jand g0720(.dina(w_n706_0[0]),.dinb(w_n689_0[0]),.dout(n784),.clk(gclk));
	jor g0721(.dina(n784),.dinb(n783),.dout(n785),.clk(gclk));
	jand g0722(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n786),.clk(gclk));
	jnot g0723(.din(n786),.dout(n787),.clk(gclk));
	jnot g0724(.din(w_n694_0[0]),.dout(n788),.clk(gclk));
	jnot g0725(.din(w_n704_0[0]),.dout(n789),.clk(gclk));
	jand g0726(.dina(n789),.dinb(n788),.dout(n790),.clk(gclk));
	jor g0727(.dina(n790),.dinb(w_n702_0[0]),.dout(n791),.clk(gclk));
	jand g0728(.dina(w_G307gat_3[2]),.dinb(w_G205gat_6[2]),.dout(n792),.clk(gclk));
	jand g0729(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n793),.clk(gclk));
	jor g0730(.dina(w_n793_0[1]),.dinb(w_n697_0[0]),.dout(n794),.clk(gclk));
	jand g0731(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n795),.clk(gclk));
	jand g0732(.dina(w_n795_0[1]),.dinb(w_n695_0[1]),.dout(n796),.clk(gclk));
	jnot g0733(.din(n796),.dout(n797),.clk(gclk));
	jand g0734(.dina(w_n797_0[2]),.dinb(n794),.dout(n798),.clk(gclk));
	jor g0735(.dina(n798),.dinb(w_n698_0[1]),.dout(n799),.clk(gclk));
	jnot g0736(.din(n799),.dout(n800),.clk(gclk));
	jand g0737(.dina(w_n797_0[1]),.dinb(w_n698_0[0]),.dout(n801),.clk(gclk));
	jor g0738(.dina(n801),.dinb(w_n800_0[1]),.dout(n802),.clk(gclk));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n792_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_n791_0[1]),.dout(n804),.clk(gclk));
	jxor g0741(.dina(w_n804_0[1]),.dinb(w_n787_0[1]),.dout(n805),.clk(gclk));
	jxor g0742(.dina(w_n805_0[1]),.dinb(w_n785_0[1]),.dout(n806),.clk(gclk));
	jxor g0743(.dina(w_n806_0[1]),.dinb(w_n782_0[1]),.dout(n807),.clk(gclk));
	jxor g0744(.dina(w_n807_0[1]),.dinb(w_n780_0[1]),.dout(n808),.clk(gclk));
	jxor g0745(.dina(w_n808_0[1]),.dinb(w_n777_0[1]),.dout(n809),.clk(gclk));
	jxor g0746(.dina(w_n809_0[1]),.dinb(w_n775_0[1]),.dout(n810),.clk(gclk));
	jxor g0747(.dina(w_n810_0[1]),.dinb(w_n772_0[1]),.dout(n811),.clk(gclk));
	jxor g0748(.dina(w_n811_0[1]),.dinb(w_n770_0[1]),.dout(n812),.clk(gclk));
	jxor g0749(.dina(w_n812_0[1]),.dinb(w_n767_0[1]),.dout(n813),.clk(gclk));
	jxor g0750(.dina(w_n813_0[1]),.dinb(w_n765_0[1]),.dout(n814),.clk(gclk));
	jxor g0751(.dina(w_n814_0[1]),.dinb(w_n762_0[1]),.dout(n815),.clk(gclk));
	jxor g0752(.dina(w_n815_0[1]),.dinb(w_n760_0[1]),.dout(n816),.clk(gclk));
	jxor g0753(.dina(w_n816_0[1]),.dinb(w_n757_0[1]),.dout(n817),.clk(gclk));
	jxor g0754(.dina(w_n817_0[1]),.dinb(w_n755_0[1]),.dout(n818),.clk(gclk));
	jxor g0755(.dina(w_n818_0[1]),.dinb(w_n752_0[1]),.dout(n819),.clk(gclk));
	jxor g0756(.dina(w_n819_0[1]),.dinb(w_n750_0[1]),.dout(n820),.clk(gclk));
	jxor g0757(.dina(w_n820_0[1]),.dinb(w_n747_0[1]),.dout(n821),.clk(gclk));
	jxor g0758(.dina(w_n821_0[1]),.dinb(w_n745_0[1]),.dout(n822),.clk(gclk));
	jxor g0759(.dina(w_n822_0[1]),.dinb(w_n742_0[1]),.dout(n823),.clk(gclk));
	jnot g0760(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jxor g0761(.dina(w_n824_0[1]),.dinb(w_n740_0[2]),.dout(n825),.clk(gclk));
	jxor g0762(.dina(n825),.dinb(n736),.dout(n826),.clk(gclk));
	jxor g0763(.dina(w_n826_0[1]),.dinb(w_n734_0[1]),.dout(n827),.clk(gclk));
	jxor g0764(.dina(w_n827_0[1]),.dinb(w_dff_B_j0VSIXt63_1),.dout(w_dff_A_HUPrWpUI2_2),.clk(gclk));
	jand g0765(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n829),.clk(gclk));
	jnot g0766(.din(w_n829_0[1]),.dout(n830),.clk(gclk));
	jnot g0767(.din(w_n826_0[0]),.dout(n831),.clk(gclk));
	jor g0768(.dina(n831),.dinb(w_n734_0[0]),.dout(n832),.clk(gclk));
	jor g0769(.dina(w_n827_0[0]),.dinb(w_n729_0[0]),.dout(n833),.clk(gclk));
	jand g0770(.dina(n833),.dinb(w_dff_B_Vw5ca9Im3_1),.dout(n834),.clk(gclk));
	jand g0771(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n835),.clk(gclk));
	jor g0772(.dina(w_n824_0[0]),.dinb(w_n740_0[1]),.dout(n836),.clk(gclk));
	jxor g0773(.dina(w_n823_0[0]),.dinb(w_n740_0[0]),.dout(n837),.clk(gclk));
	jor g0774(.dina(n837),.dinb(w_n735_0[0]),.dout(n838),.clk(gclk));
	jand g0775(.dina(n838),.dinb(n836),.dout(n839),.clk(gclk));
	jand g0776(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n840),.clk(gclk));
	jnot g0777(.din(w_n840_0[1]),.dout(n841),.clk(gclk));
	jand g0778(.dina(w_n821_0[0]),.dinb(w_n745_0[0]),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n822_0[0]),.dinb(w_n742_0[0]),.dout(n843),.clk(gclk));
	jor g0780(.dina(n843),.dinb(n842),.dout(n844),.clk(gclk));
	jand g0781(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n845),.clk(gclk));
	jnot g0782(.din(n845),.dout(n846),.clk(gclk));
	jand g0783(.dina(w_n819_0[0]),.dinb(w_n750_0[0]),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n820_0[0]),.dinb(w_n747_0[0]),.dout(n848),.clk(gclk));
	jor g0785(.dina(n848),.dinb(n847),.dout(n849),.clk(gclk));
	jand g0786(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n850),.clk(gclk));
	jnot g0787(.din(n850),.dout(n851),.clk(gclk));
	jand g0788(.dina(w_n817_0[0]),.dinb(w_n755_0[0]),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n818_0[0]),.dinb(w_n752_0[0]),.dout(n853),.clk(gclk));
	jor g0790(.dina(n853),.dinb(n852),.dout(n854),.clk(gclk));
	jand g0791(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n855),.clk(gclk));
	jnot g0792(.din(n855),.dout(n856),.clk(gclk));
	jand g0793(.dina(w_n815_0[0]),.dinb(w_n760_0[0]),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n816_0[0]),.dinb(w_n757_0[0]),.dout(n858),.clk(gclk));
	jor g0795(.dina(n858),.dinb(n857),.dout(n859),.clk(gclk));
	jand g0796(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n860),.clk(gclk));
	jnot g0797(.din(n860),.dout(n861),.clk(gclk));
	jand g0798(.dina(w_n813_0[0]),.dinb(w_n765_0[0]),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n814_0[0]),.dinb(w_n762_0[0]),.dout(n863),.clk(gclk));
	jor g0800(.dina(n863),.dinb(n862),.dout(n864),.clk(gclk));
	jand g0801(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n865),.clk(gclk));
	jnot g0802(.din(n865),.dout(n866),.clk(gclk));
	jand g0803(.dina(w_n811_0[0]),.dinb(w_n770_0[0]),.dout(n867),.clk(gclk));
	jand g0804(.dina(w_n812_0[0]),.dinb(w_n767_0[0]),.dout(n868),.clk(gclk));
	jor g0805(.dina(n868),.dinb(n867),.dout(n869),.clk(gclk));
	jand g0806(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n870),.clk(gclk));
	jnot g0807(.din(n870),.dout(n871),.clk(gclk));
	jand g0808(.dina(w_n809_0[0]),.dinb(w_n775_0[0]),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_n810_0[0]),.dinb(w_n772_0[0]),.dout(n873),.clk(gclk));
	jor g0810(.dina(n873),.dinb(n872),.dout(n874),.clk(gclk));
	jand g0811(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n875),.clk(gclk));
	jnot g0812(.din(n875),.dout(n876),.clk(gclk));
	jand g0813(.dina(w_n807_0[0]),.dinb(w_n780_0[0]),.dout(n877),.clk(gclk));
	jand g0814(.dina(w_n808_0[0]),.dinb(w_n777_0[0]),.dout(n878),.clk(gclk));
	jor g0815(.dina(n878),.dinb(n877),.dout(n879),.clk(gclk));
	jand g0816(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n880),.clk(gclk));
	jnot g0817(.din(n880),.dout(n881),.clk(gclk));
	jand g0818(.dina(w_n805_0[0]),.dinb(w_n785_0[0]),.dout(n882),.clk(gclk));
	jand g0819(.dina(w_n806_0[0]),.dinb(w_n782_0[0]),.dout(n883),.clk(gclk));
	jor g0820(.dina(n883),.dinb(n882),.dout(n884),.clk(gclk));
	jand g0821(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n885),.clk(gclk));
	jnot g0822(.din(n885),.dout(n886),.clk(gclk));
	jand g0823(.dina(w_n803_0[0]),.dinb(w_n791_0[0]),.dout(n887),.clk(gclk));
	jand g0824(.dina(w_n804_0[0]),.dinb(w_n787_0[0]),.dout(n888),.clk(gclk));
	jor g0825(.dina(n888),.dinb(n887),.dout(n889),.clk(gclk));
	jand g0826(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n890),.clk(gclk));
	jnot g0827(.din(n890),.dout(n891),.clk(gclk));
	jnot g0828(.din(w_n792_0[0]),.dout(n892),.clk(gclk));
	jnot g0829(.din(w_n802_0[0]),.dout(n893),.clk(gclk));
	jand g0830(.dina(n893),.dinb(n892),.dout(n894),.clk(gclk));
	jor g0831(.dina(n894),.dinb(w_n800_0[0]),.dout(n895),.clk(gclk));
	jand g0832(.dina(w_G307gat_3[1]),.dinb(w_G222gat_6[2]),.dout(n896),.clk(gclk));
	jnot g0833(.din(w_n795_0[0]),.dout(n897),.clk(gclk));
	jand g0834(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n898),.clk(gclk));
	jand g0835(.dina(w_n898_0[1]),.dinb(w_n897_0[1]),.dout(n899),.clk(gclk));
	jnot g0836(.din(n899),.dout(n900),.clk(gclk));
	jor g0837(.dina(w_n898_0[0]),.dinb(w_n897_0[0]),.dout(n901),.clk(gclk));
	jand g0838(.dina(w_n901_0[1]),.dinb(w_n797_0[0]),.dout(n902),.clk(gclk));
	jand g0839(.dina(n902),.dinb(n900),.dout(n903),.clk(gclk));
	jnot g0840(.din(w_n901_0[0]),.dout(n904),.clk(gclk));
	jand g0841(.dina(n904),.dinb(w_n695_0[0]),.dout(n905),.clk(gclk));
	jor g0842(.dina(n905),.dinb(w_n903_0[1]),.dout(n906),.clk(gclk));
	jxor g0843(.dina(w_n906_0[1]),.dinb(w_n896_0[1]),.dout(n907),.clk(gclk));
	jxor g0844(.dina(w_n907_0[1]),.dinb(w_n895_0[1]),.dout(n908),.clk(gclk));
	jxor g0845(.dina(w_n908_0[1]),.dinb(w_n891_0[1]),.dout(n909),.clk(gclk));
	jxor g0846(.dina(w_n909_0[1]),.dinb(w_n889_0[1]),.dout(n910),.clk(gclk));
	jxor g0847(.dina(w_n910_0[1]),.dinb(w_n886_0[1]),.dout(n911),.clk(gclk));
	jxor g0848(.dina(w_n911_0[1]),.dinb(w_n884_0[1]),.dout(n912),.clk(gclk));
	jxor g0849(.dina(w_n912_0[1]),.dinb(w_n881_0[1]),.dout(n913),.clk(gclk));
	jxor g0850(.dina(w_n913_0[1]),.dinb(w_n879_0[1]),.dout(n914),.clk(gclk));
	jxor g0851(.dina(w_n914_0[1]),.dinb(w_n876_0[1]),.dout(n915),.clk(gclk));
	jxor g0852(.dina(w_n915_0[1]),.dinb(w_n874_0[1]),.dout(n916),.clk(gclk));
	jxor g0853(.dina(w_n916_0[1]),.dinb(w_n871_0[1]),.dout(n917),.clk(gclk));
	jxor g0854(.dina(w_n917_0[1]),.dinb(w_n869_0[1]),.dout(n918),.clk(gclk));
	jxor g0855(.dina(w_n918_0[1]),.dinb(w_n866_0[1]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(w_n919_0[1]),.dinb(w_n864_0[1]),.dout(n920),.clk(gclk));
	jxor g0857(.dina(w_n920_0[1]),.dinb(w_n861_0[1]),.dout(n921),.clk(gclk));
	jxor g0858(.dina(w_n921_0[1]),.dinb(w_n859_0[1]),.dout(n922),.clk(gclk));
	jxor g0859(.dina(w_n922_0[1]),.dinb(w_n856_0[1]),.dout(n923),.clk(gclk));
	jxor g0860(.dina(w_n923_0[1]),.dinb(w_n854_0[1]),.dout(n924),.clk(gclk));
	jxor g0861(.dina(w_n924_0[1]),.dinb(w_n851_0[1]),.dout(n925),.clk(gclk));
	jxor g0862(.dina(w_n925_0[1]),.dinb(w_n849_0[1]),.dout(n926),.clk(gclk));
	jxor g0863(.dina(w_n926_0[1]),.dinb(w_n846_0[1]),.dout(n927),.clk(gclk));
	jxor g0864(.dina(w_n927_0[2]),.dinb(w_n844_0[2]),.dout(n928),.clk(gclk));
	jxor g0865(.dina(n928),.dinb(n841),.dout(n929),.clk(gclk));
	jxor g0866(.dina(w_n929_0[1]),.dinb(w_n839_0[1]),.dout(n930),.clk(gclk));
	jxor g0867(.dina(w_n930_0[1]),.dinb(w_n835_0[1]),.dout(n931),.clk(gclk));
	jxor g0868(.dina(w_n931_0[1]),.dinb(w_n834_0[1]),.dout(n932),.clk(gclk));
	jxor g0869(.dina(w_n932_0[1]),.dinb(w_dff_B_fP7WTlcY5_1),.dout(w_dff_A_dkRXDqWE6_2),.clk(gclk));
	jnot g0870(.din(w_n931_0[0]),.dout(n934),.clk(gclk));
	jor g0871(.dina(n934),.dinb(w_n834_0[0]),.dout(n935),.clk(gclk));
	jor g0872(.dina(w_n932_0[0]),.dinb(w_n829_0[0]),.dout(n936),.clk(gclk));
	jand g0873(.dina(n936),.dinb(w_dff_B_39iS0oOH0_1),.dout(n937),.clk(gclk));
	jand g0874(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n938),.clk(gclk));
	jnot g0875(.din(w_n929_0[0]),.dout(n939),.clk(gclk));
	jor g0876(.dina(n939),.dinb(w_n839_0[0]),.dout(n940),.clk(gclk));
	jor g0877(.dina(w_n930_0[0]),.dinb(w_n835_0[0]),.dout(n941),.clk(gclk));
	jand g0878(.dina(n941),.dinb(n940),.dout(n942),.clk(gclk));
	jand g0879(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n943),.clk(gclk));
	jand g0880(.dina(w_n927_0[1]),.dinb(w_n844_0[1]),.dout(n944),.clk(gclk));
	jnot g0881(.din(n944),.dout(n945),.clk(gclk));
	jnot g0882(.din(w_n927_0[0]),.dout(n946),.clk(gclk));
	jxor g0883(.dina(n946),.dinb(w_n844_0[0]),.dout(n947),.clk(gclk));
	jor g0884(.dina(n947),.dinb(w_n840_0[0]),.dout(n948),.clk(gclk));
	jand g0885(.dina(n948),.dinb(n945),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n950),.clk(gclk));
	jnot g0887(.din(n950),.dout(n951),.clk(gclk));
	jand g0888(.dina(w_n925_0[0]),.dinb(w_n849_0[0]),.dout(n952),.clk(gclk));
	jand g0889(.dina(w_n926_0[0]),.dinb(w_n846_0[0]),.dout(n953),.clk(gclk));
	jor g0890(.dina(n953),.dinb(n952),.dout(n954),.clk(gclk));
	jand g0891(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n955),.clk(gclk));
	jnot g0892(.din(n955),.dout(n956),.clk(gclk));
	jand g0893(.dina(w_n923_0[0]),.dinb(w_n854_0[0]),.dout(n957),.clk(gclk));
	jand g0894(.dina(w_n924_0[0]),.dinb(w_n851_0[0]),.dout(n958),.clk(gclk));
	jor g0895(.dina(n958),.dinb(n957),.dout(n959),.clk(gclk));
	jand g0896(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n960),.clk(gclk));
	jnot g0897(.din(n960),.dout(n961),.clk(gclk));
	jand g0898(.dina(w_n921_0[0]),.dinb(w_n859_0[0]),.dout(n962),.clk(gclk));
	jand g0899(.dina(w_n922_0[0]),.dinb(w_n856_0[0]),.dout(n963),.clk(gclk));
	jor g0900(.dina(n963),.dinb(n962),.dout(n964),.clk(gclk));
	jand g0901(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n965),.clk(gclk));
	jnot g0902(.din(n965),.dout(n966),.clk(gclk));
	jand g0903(.dina(w_n919_0[0]),.dinb(w_n864_0[0]),.dout(n967),.clk(gclk));
	jand g0904(.dina(w_n920_0[0]),.dinb(w_n861_0[0]),.dout(n968),.clk(gclk));
	jor g0905(.dina(n968),.dinb(n967),.dout(n969),.clk(gclk));
	jand g0906(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n970),.clk(gclk));
	jnot g0907(.din(n970),.dout(n971),.clk(gclk));
	jand g0908(.dina(w_n917_0[0]),.dinb(w_n869_0[0]),.dout(n972),.clk(gclk));
	jand g0909(.dina(w_n918_0[0]),.dinb(w_n866_0[0]),.dout(n973),.clk(gclk));
	jor g0910(.dina(n973),.dinb(n972),.dout(n974),.clk(gclk));
	jand g0911(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(w_n915_0[0]),.dinb(w_n874_0[0]),.dout(n977),.clk(gclk));
	jand g0914(.dina(w_n916_0[0]),.dinb(w_n871_0[0]),.dout(n978),.clk(gclk));
	jor g0915(.dina(n978),.dinb(n977),.dout(n979),.clk(gclk));
	jand g0916(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n980),.clk(gclk));
	jnot g0917(.din(n980),.dout(n981),.clk(gclk));
	jand g0918(.dina(w_n913_0[0]),.dinb(w_n879_0[0]),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_n914_0[0]),.dinb(w_n876_0[0]),.dout(n983),.clk(gclk));
	jor g0920(.dina(n983),.dinb(n982),.dout(n984),.clk(gclk));
	jand g0921(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n985),.clk(gclk));
	jnot g0922(.din(n985),.dout(n986),.clk(gclk));
	jand g0923(.dina(w_n911_0[0]),.dinb(w_n884_0[0]),.dout(n987),.clk(gclk));
	jand g0924(.dina(w_n912_0[0]),.dinb(w_n881_0[0]),.dout(n988),.clk(gclk));
	jor g0925(.dina(n988),.dinb(n987),.dout(n989),.clk(gclk));
	jand g0926(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n990),.clk(gclk));
	jnot g0927(.din(n990),.dout(n991),.clk(gclk));
	jand g0928(.dina(w_n909_0[0]),.dinb(w_n889_0[0]),.dout(n992),.clk(gclk));
	jand g0929(.dina(w_n910_0[0]),.dinb(w_n886_0[0]),.dout(n993),.clk(gclk));
	jor g0930(.dina(n993),.dinb(n992),.dout(n994),.clk(gclk));
	jand g0931(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n995),.clk(gclk));
	jnot g0932(.din(n995),.dout(n996),.clk(gclk));
	jand g0933(.dina(w_n907_0[0]),.dinb(w_n895_0[0]),.dout(n997),.clk(gclk));
	jand g0934(.dina(w_n908_0[0]),.dinb(w_n891_0[0]),.dout(n998),.clk(gclk));
	jor g0935(.dina(n998),.dinb(n997),.dout(n999),.clk(gclk));
	jand g0936(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n1000),.clk(gclk));
	jnot g0937(.din(n1000),.dout(n1001),.clk(gclk));
	jnot g0938(.din(w_n896_0[0]),.dout(n1002),.clk(gclk));
	jnot g0939(.din(w_n906_0[0]),.dout(n1003),.clk(gclk));
	jand g0940(.dina(n1003),.dinb(n1002),.dout(n1004),.clk(gclk));
	jor g0941(.dina(n1004),.dinb(w_n903_0[0]),.dout(n1005),.clk(gclk));
	jand g0942(.dina(w_G307gat_3[0]),.dinb(w_G239gat_6[2]),.dout(n1006),.clk(gclk));
	jand g0943(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n1007),.clk(gclk));
	jnot g0944(.din(n1007),.dout(n1008),.clk(gclk));
	jor g0945(.dina(w_n1008_0[1]),.dinb(w_n793_0[0]),.dout(n1009),.clk(gclk));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n1006_0[1]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(w_n1010_0[1]),.dinb(w_n1005_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n1001_0[1]),.dout(n1012),.clk(gclk));
	jxor g0949(.dina(w_n1012_0[1]),.dinb(w_n999_0[1]),.dout(n1013),.clk(gclk));
	jxor g0950(.dina(w_n1013_0[1]),.dinb(w_n996_0[1]),.dout(n1014),.clk(gclk));
	jxor g0951(.dina(w_n1014_0[1]),.dinb(w_n994_0[1]),.dout(n1015),.clk(gclk));
	jxor g0952(.dina(w_n1015_0[1]),.dinb(w_n991_0[1]),.dout(n1016),.clk(gclk));
	jxor g0953(.dina(w_n1016_0[1]),.dinb(w_n989_0[1]),.dout(n1017),.clk(gclk));
	jxor g0954(.dina(w_n1017_0[1]),.dinb(w_n986_0[1]),.dout(n1018),.clk(gclk));
	jxor g0955(.dina(w_n1018_0[1]),.dinb(w_n984_0[1]),.dout(n1019),.clk(gclk));
	jxor g0956(.dina(w_n1019_0[1]),.dinb(w_n981_0[1]),.dout(n1020),.clk(gclk));
	jxor g0957(.dina(w_n1020_0[1]),.dinb(w_n979_0[1]),.dout(n1021),.clk(gclk));
	jxor g0958(.dina(w_n1021_0[1]),.dinb(w_n976_0[1]),.dout(n1022),.clk(gclk));
	jxor g0959(.dina(w_n1022_0[1]),.dinb(w_n974_0[1]),.dout(n1023),.clk(gclk));
	jxor g0960(.dina(w_n1023_0[1]),.dinb(w_n971_0[1]),.dout(n1024),.clk(gclk));
	jxor g0961(.dina(w_n1024_0[1]),.dinb(w_n969_0[1]),.dout(n1025),.clk(gclk));
	jxor g0962(.dina(w_n1025_0[1]),.dinb(w_n966_0[1]),.dout(n1026),.clk(gclk));
	jxor g0963(.dina(w_n1026_0[1]),.dinb(w_n964_0[1]),.dout(n1027),.clk(gclk));
	jxor g0964(.dina(w_n1027_0[1]),.dinb(w_n961_0[1]),.dout(n1028),.clk(gclk));
	jxor g0965(.dina(w_n1028_0[1]),.dinb(w_n959_0[1]),.dout(n1029),.clk(gclk));
	jxor g0966(.dina(w_n1029_0[1]),.dinb(w_n956_0[1]),.dout(n1030),.clk(gclk));
	jxor g0967(.dina(w_n1030_0[1]),.dinb(w_n954_0[1]),.dout(n1031),.clk(gclk));
	jxor g0968(.dina(w_n1031_0[1]),.dinb(w_n951_0[1]),.dout(n1032),.clk(gclk));
	jxor g0969(.dina(w_n1032_0[1]),.dinb(w_n949_0[1]),.dout(n1033),.clk(gclk));
	jxor g0970(.dina(w_n1033_0[1]),.dinb(w_n943_0[1]),.dout(n1034),.clk(gclk));
	jnot g0971(.din(w_n1034_0[1]),.dout(n1035),.clk(gclk));
	jxor g0972(.dina(w_n1035_0[1]),.dinb(w_n942_0[2]),.dout(n1036),.clk(gclk));
	jxor g0973(.dina(n1036),.dinb(w_n938_0[1]),.dout(n1037),.clk(gclk));
	jxor g0974(.dina(w_n1037_0[1]),.dinb(w_n937_0[1]),.dout(w_dff_A_XP7KI9S09_2),.clk(gclk));
	jand g0975(.dina(w_n1037_0[0]),.dinb(w_n937_0[0]),.dout(n1039),.clk(gclk));
	jor g0976(.dina(w_n1035_0[0]),.dinb(w_n942_0[1]),.dout(n1040),.clk(gclk));
	jxor g0977(.dina(w_n1034_0[0]),.dinb(w_n942_0[0]),.dout(n1041),.clk(gclk));
	jor g0978(.dina(n1041),.dinb(w_n938_0[0]),.dout(n1042),.clk(gclk));
	jand g0979(.dina(n1042),.dinb(n1040),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1044),.clk(gclk));
	jnot g0981(.din(w_n1032_0[0]),.dout(n1045),.clk(gclk));
	jor g0982(.dina(n1045),.dinb(w_n949_0[0]),.dout(n1046),.clk(gclk));
	jor g0983(.dina(w_n1033_0[0]),.dinb(w_n943_0[0]),.dout(n1047),.clk(gclk));
	jand g0984(.dina(n1047),.dinb(n1046),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n1030_0[0]),.dinb(w_n954_0[0]),.dout(n1050),.clk(gclk));
	jand g0987(.dina(w_n1031_0[0]),.dinb(w_n951_0[0]),.dout(n1051),.clk(gclk));
	jor g0988(.dina(n1051),.dinb(n1050),.dout(n1052),.clk(gclk));
	jand g0989(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1053),.clk(gclk));
	jnot g0990(.din(n1053),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n1028_0[0]),.dinb(w_n959_0[0]),.dout(n1055),.clk(gclk));
	jand g0992(.dina(w_n1029_0[0]),.dinb(w_n956_0[0]),.dout(n1056),.clk(gclk));
	jor g0993(.dina(n1056),.dinb(n1055),.dout(n1057),.clk(gclk));
	jand g0994(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1058),.clk(gclk));
	jnot g0995(.din(n1058),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n1026_0[0]),.dinb(w_n964_0[0]),.dout(n1060),.clk(gclk));
	jand g0997(.dina(w_n1027_0[0]),.dinb(w_n961_0[0]),.dout(n1061),.clk(gclk));
	jor g0998(.dina(n1061),.dinb(n1060),.dout(n1062),.clk(gclk));
	jand g0999(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1063),.clk(gclk));
	jnot g1000(.din(n1063),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n1024_0[0]),.dinb(w_n969_0[0]),.dout(n1065),.clk(gclk));
	jand g1002(.dina(w_n1025_0[0]),.dinb(w_n966_0[0]),.dout(n1066),.clk(gclk));
	jor g1003(.dina(n1066),.dinb(n1065),.dout(n1067),.clk(gclk));
	jand g1004(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1068),.clk(gclk));
	jnot g1005(.din(n1068),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n1022_0[0]),.dinb(w_n974_0[0]),.dout(n1070),.clk(gclk));
	jand g1007(.dina(w_n1023_0[0]),.dinb(w_n971_0[0]),.dout(n1071),.clk(gclk));
	jor g1008(.dina(n1071),.dinb(n1070),.dout(n1072),.clk(gclk));
	jand g1009(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1073),.clk(gclk));
	jnot g1010(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n1020_0[0]),.dinb(w_n979_0[0]),.dout(n1075),.clk(gclk));
	jand g1012(.dina(w_n1021_0[0]),.dinb(w_n976_0[0]),.dout(n1076),.clk(gclk));
	jor g1013(.dina(n1076),.dinb(n1075),.dout(n1077),.clk(gclk));
	jand g1014(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1078),.clk(gclk));
	jnot g1015(.din(n1078),.dout(n1079),.clk(gclk));
	jand g1016(.dina(w_n1018_0[0]),.dinb(w_n984_0[0]),.dout(n1080),.clk(gclk));
	jand g1017(.dina(w_n1019_0[0]),.dinb(w_n981_0[0]),.dout(n1081),.clk(gclk));
	jor g1018(.dina(n1081),.dinb(n1080),.dout(n1082),.clk(gclk));
	jand g1019(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1083),.clk(gclk));
	jnot g1020(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1021(.dina(w_n1016_0[0]),.dinb(w_n989_0[0]),.dout(n1085),.clk(gclk));
	jand g1022(.dina(w_n1017_0[0]),.dinb(w_n986_0[0]),.dout(n1086),.clk(gclk));
	jor g1023(.dina(n1086),.dinb(n1085),.dout(n1087),.clk(gclk));
	jand g1024(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1088),.clk(gclk));
	jnot g1025(.din(n1088),.dout(n1089),.clk(gclk));
	jand g1026(.dina(w_n1014_0[0]),.dinb(w_n994_0[0]),.dout(n1090),.clk(gclk));
	jand g1027(.dina(w_n1015_0[0]),.dinb(w_n991_0[0]),.dout(n1091),.clk(gclk));
	jor g1028(.dina(n1091),.dinb(n1090),.dout(n1092),.clk(gclk));
	jand g1029(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1093),.clk(gclk));
	jnot g1030(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1031(.dina(w_n1012_0[0]),.dinb(w_n999_0[0]),.dout(n1095),.clk(gclk));
	jand g1032(.dina(w_n1013_0[0]),.dinb(w_n996_0[0]),.dout(n1096),.clk(gclk));
	jor g1033(.dina(n1096),.dinb(n1095),.dout(n1097),.clk(gclk));
	jand g1034(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1098),.clk(gclk));
	jnot g1035(.din(n1098),.dout(n1099),.clk(gclk));
	jand g1036(.dina(w_n1010_0[0]),.dinb(w_n1005_0[0]),.dout(n1100),.clk(gclk));
	jand g1037(.dina(w_n1011_0[0]),.dinb(w_n1001_0[0]),.dout(n1101),.clk(gclk));
	jor g1038(.dina(n1101),.dinb(n1100),.dout(n1102),.clk(gclk));
	jand g1039(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1103),.clk(gclk));
	jand g1040(.dina(w_G307gat_2[2]),.dinb(w_G256gat_6[2]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(w_n1006_0[0]),.dout(n1105),.clk(gclk));
	jnot g1042(.din(w_n1009_0[0]),.dout(n1106),.clk(gclk));
	jand g1043(.dina(n1106),.dinb(n1105),.dout(n1107),.clk(gclk));
	jor g1044(.dina(n1107),.dinb(w_n1008_0[0]),.dout(n1108),.clk(gclk));
	jnot g1045(.din(n1108),.dout(n1109),.clk(gclk));
	jor g1046(.dina(w_n1109_0[1]),.dinb(n1104),.dout(n1110),.clk(gclk));
	jand g1047(.dina(w_n1109_0[0]),.dinb(w_G307gat_2[1]),.dout(n1111),.clk(gclk));
	jnot g1048(.din(n1111),.dout(n1112),.clk(gclk));
	jand g1049(.dina(n1112),.dinb(w_n1110_0[1]),.dout(n1113),.clk(gclk));
	jnot g1050(.din(n1113),.dout(n1114),.clk(gclk));
	jxor g1051(.dina(w_n1114_0[1]),.dinb(w_n1103_0[1]),.dout(n1115),.clk(gclk));
	jxor g1052(.dina(w_n1115_0[1]),.dinb(w_n1102_0[1]),.dout(n1116),.clk(gclk));
	jxor g1053(.dina(w_n1116_0[1]),.dinb(w_n1099_0[1]),.dout(n1117),.clk(gclk));
	jxor g1054(.dina(w_n1117_0[1]),.dinb(w_n1097_0[1]),.dout(n1118),.clk(gclk));
	jxor g1055(.dina(w_n1118_0[1]),.dinb(w_n1094_0[1]),.dout(n1119),.clk(gclk));
	jxor g1056(.dina(w_n1119_0[1]),.dinb(w_n1092_0[1]),.dout(n1120),.clk(gclk));
	jxor g1057(.dina(w_n1120_0[1]),.dinb(w_n1089_0[1]),.dout(n1121),.clk(gclk));
	jxor g1058(.dina(w_n1121_0[1]),.dinb(w_n1087_0[1]),.dout(n1122),.clk(gclk));
	jxor g1059(.dina(w_n1122_0[1]),.dinb(w_n1084_0[1]),.dout(n1123),.clk(gclk));
	jxor g1060(.dina(w_n1123_0[1]),.dinb(w_n1082_0[1]),.dout(n1124),.clk(gclk));
	jxor g1061(.dina(w_n1124_0[1]),.dinb(w_n1079_0[1]),.dout(n1125),.clk(gclk));
	jxor g1062(.dina(w_n1125_0[1]),.dinb(w_n1077_0[1]),.dout(n1126),.clk(gclk));
	jxor g1063(.dina(w_n1126_0[1]),.dinb(w_n1074_0[1]),.dout(n1127),.clk(gclk));
	jxor g1064(.dina(w_n1127_0[1]),.dinb(w_n1072_0[1]),.dout(n1128),.clk(gclk));
	jxor g1065(.dina(w_n1128_0[1]),.dinb(w_n1069_0[1]),.dout(n1129),.clk(gclk));
	jxor g1066(.dina(w_n1129_0[1]),.dinb(w_n1067_0[1]),.dout(n1130),.clk(gclk));
	jxor g1067(.dina(w_n1130_0[1]),.dinb(w_n1064_0[1]),.dout(n1131),.clk(gclk));
	jxor g1068(.dina(w_n1131_0[1]),.dinb(w_n1062_0[1]),.dout(n1132),.clk(gclk));
	jxor g1069(.dina(w_n1132_0[1]),.dinb(w_n1059_0[1]),.dout(n1133),.clk(gclk));
	jxor g1070(.dina(w_n1133_0[1]),.dinb(w_n1057_0[1]),.dout(n1134),.clk(gclk));
	jxor g1071(.dina(w_n1134_0[1]),.dinb(w_n1054_0[1]),.dout(n1135),.clk(gclk));
	jxor g1072(.dina(w_n1135_0[1]),.dinb(w_n1052_0[1]),.dout(n1136),.clk(gclk));
	jnot g1073(.din(n1136),.dout(n1137),.clk(gclk));
	jxor g1074(.dina(w_n1137_0[1]),.dinb(w_n1049_0[1]),.dout(n1138),.clk(gclk));
	jxor g1075(.dina(w_n1138_0[1]),.dinb(w_n1048_0[1]),.dout(n1139),.clk(gclk));
	jxor g1076(.dina(w_n1139_0[1]),.dinb(w_n1044_0[1]),.dout(n1140),.clk(gclk));
	jxor g1077(.dina(w_n1140_0[1]),.dinb(w_n1043_0[1]),.dout(n1141),.clk(gclk));
	jnot g1078(.din(w_n1141_0[1]),.dout(n1142),.clk(gclk));
	jxor g1079(.dina(n1142),.dinb(w_n1039_0[1]),.dout(w_dff_A_muYCmXs49_2),.clk(gclk));
	jnot g1080(.din(w_n1140_0[0]),.dout(n1144),.clk(gclk));
	jor g1081(.dina(n1144),.dinb(w_n1043_0[0]),.dout(n1145),.clk(gclk));
	jor g1082(.dina(w_n1141_0[0]),.dinb(w_n1039_0[0]),.dout(n1146),.clk(gclk));
	jand g1083(.dina(n1146),.dinb(w_dff_B_avGxlZft2_1),.dout(n1147),.clk(gclk));
	jnot g1084(.din(w_n1138_0[0]),.dout(n1148),.clk(gclk));
	jor g1085(.dina(n1148),.dinb(w_n1048_0[0]),.dout(n1149),.clk(gclk));
	jor g1086(.dina(w_n1139_0[0]),.dinb(w_n1044_0[0]),.dout(n1150),.clk(gclk));
	jand g1087(.dina(n1150),.dinb(n1149),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1135_0[0]),.dinb(w_n1052_0[0]),.dout(n1153),.clk(gclk));
	jnot g1090(.din(n1153),.dout(n1154),.clk(gclk));
	jor g1091(.dina(w_n1137_0[0]),.dinb(w_n1049_0[0]),.dout(n1155),.clk(gclk));
	jand g1092(.dina(n1155),.dinb(n1154),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1157),.clk(gclk));
	jnot g1094(.din(n1157),.dout(n1158),.clk(gclk));
	jand g1095(.dina(w_n1133_0[0]),.dinb(w_n1057_0[0]),.dout(n1159),.clk(gclk));
	jand g1096(.dina(w_n1134_0[0]),.dinb(w_n1054_0[0]),.dout(n1160),.clk(gclk));
	jor g1097(.dina(n1160),.dinb(n1159),.dout(n1161),.clk(gclk));
	jand g1098(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1162),.clk(gclk));
	jnot g1099(.din(n1162),.dout(n1163),.clk(gclk));
	jand g1100(.dina(w_n1131_0[0]),.dinb(w_n1062_0[0]),.dout(n1164),.clk(gclk));
	jand g1101(.dina(w_n1132_0[0]),.dinb(w_n1059_0[0]),.dout(n1165),.clk(gclk));
	jor g1102(.dina(n1165),.dinb(n1164),.dout(n1166),.clk(gclk));
	jand g1103(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1167),.clk(gclk));
	jnot g1104(.din(n1167),.dout(n1168),.clk(gclk));
	jand g1105(.dina(w_n1129_0[0]),.dinb(w_n1067_0[0]),.dout(n1169),.clk(gclk));
	jand g1106(.dina(w_n1130_0[0]),.dinb(w_n1064_0[0]),.dout(n1170),.clk(gclk));
	jor g1107(.dina(n1170),.dinb(n1169),.dout(n1171),.clk(gclk));
	jand g1108(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1172),.clk(gclk));
	jnot g1109(.din(n1172),.dout(n1173),.clk(gclk));
	jand g1110(.dina(w_n1127_0[0]),.dinb(w_n1072_0[0]),.dout(n1174),.clk(gclk));
	jand g1111(.dina(w_n1128_0[0]),.dinb(w_n1069_0[0]),.dout(n1175),.clk(gclk));
	jor g1112(.dina(n1175),.dinb(n1174),.dout(n1176),.clk(gclk));
	jand g1113(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1177),.clk(gclk));
	jnot g1114(.din(n1177),.dout(n1178),.clk(gclk));
	jand g1115(.dina(w_n1125_0[0]),.dinb(w_n1077_0[0]),.dout(n1179),.clk(gclk));
	jand g1116(.dina(w_n1126_0[0]),.dinb(w_n1074_0[0]),.dout(n1180),.clk(gclk));
	jor g1117(.dina(n1180),.dinb(n1179),.dout(n1181),.clk(gclk));
	jand g1118(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1182),.clk(gclk));
	jnot g1119(.din(n1182),.dout(n1183),.clk(gclk));
	jand g1120(.dina(w_n1123_0[0]),.dinb(w_n1082_0[0]),.dout(n1184),.clk(gclk));
	jand g1121(.dina(w_n1124_0[0]),.dinb(w_n1079_0[0]),.dout(n1185),.clk(gclk));
	jor g1122(.dina(n1185),.dinb(n1184),.dout(n1186),.clk(gclk));
	jand g1123(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1187),.clk(gclk));
	jnot g1124(.din(n1187),.dout(n1188),.clk(gclk));
	jand g1125(.dina(w_n1121_0[0]),.dinb(w_n1087_0[0]),.dout(n1189),.clk(gclk));
	jand g1126(.dina(w_n1122_0[0]),.dinb(w_n1084_0[0]),.dout(n1190),.clk(gclk));
	jor g1127(.dina(n1190),.dinb(n1189),.dout(n1191),.clk(gclk));
	jand g1128(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1192),.clk(gclk));
	jnot g1129(.din(n1192),.dout(n1193),.clk(gclk));
	jand g1130(.dina(w_n1119_0[0]),.dinb(w_n1092_0[0]),.dout(n1194),.clk(gclk));
	jand g1131(.dina(w_n1120_0[0]),.dinb(w_n1089_0[0]),.dout(n1195),.clk(gclk));
	jor g1132(.dina(n1195),.dinb(n1194),.dout(n1196),.clk(gclk));
	jand g1133(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1197),.clk(gclk));
	jnot g1134(.din(n1197),.dout(n1198),.clk(gclk));
	jand g1135(.dina(w_n1117_0[0]),.dinb(w_n1097_0[0]),.dout(n1199),.clk(gclk));
	jand g1136(.dina(w_n1118_0[0]),.dinb(w_n1094_0[0]),.dout(n1200),.clk(gclk));
	jor g1137(.dina(n1200),.dinb(n1199),.dout(n1201),.clk(gclk));
	jand g1138(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jand g1140(.dina(w_n1115_0[0]),.dinb(w_n1102_0[0]),.dout(n1204),.clk(gclk));
	jand g1141(.dina(w_n1116_0[0]),.dinb(w_n1099_0[0]),.dout(n1205),.clk(gclk));
	jor g1142(.dina(n1205),.dinb(n1204),.dout(n1206),.clk(gclk));
	jand g1143(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1207),.clk(gclk));
	jand g1144(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1208),.clk(gclk));
	jor g1145(.dina(w_n1114_0[0]),.dinb(w_n1103_0[0]),.dout(n1209),.clk(gclk));
	jand g1146(.dina(n1209),.dinb(w_n1110_0[0]),.dout(n1210),.clk(gclk));
	jxor g1147(.dina(w_n1210_0[1]),.dinb(w_n1208_0[1]),.dout(n1211),.clk(gclk));
	jnot g1148(.din(n1211),.dout(n1212),.clk(gclk));
	jxor g1149(.dina(w_n1212_0[1]),.dinb(w_n1207_0[1]),.dout(n1213),.clk(gclk));
	jxor g1150(.dina(w_n1213_0[1]),.dinb(w_n1206_0[1]),.dout(n1214),.clk(gclk));
	jxor g1151(.dina(w_n1214_0[1]),.dinb(w_n1203_0[1]),.dout(n1215),.clk(gclk));
	jxor g1152(.dina(w_n1215_0[1]),.dinb(w_n1201_0[1]),.dout(n1216),.clk(gclk));
	jxor g1153(.dina(w_n1216_0[1]),.dinb(w_n1198_0[1]),.dout(n1217),.clk(gclk));
	jxor g1154(.dina(w_n1217_0[1]),.dinb(w_n1196_0[1]),.dout(n1218),.clk(gclk));
	jxor g1155(.dina(w_n1218_0[1]),.dinb(w_n1193_0[1]),.dout(n1219),.clk(gclk));
	jxor g1156(.dina(w_n1219_0[1]),.dinb(w_n1191_0[1]),.dout(n1220),.clk(gclk));
	jxor g1157(.dina(w_n1220_0[1]),.dinb(w_n1188_0[1]),.dout(n1221),.clk(gclk));
	jxor g1158(.dina(w_n1221_0[1]),.dinb(w_n1186_0[1]),.dout(n1222),.clk(gclk));
	jxor g1159(.dina(w_n1222_0[1]),.dinb(w_n1183_0[1]),.dout(n1223),.clk(gclk));
	jxor g1160(.dina(w_n1223_0[1]),.dinb(w_n1181_0[1]),.dout(n1224),.clk(gclk));
	jxor g1161(.dina(w_n1224_0[1]),.dinb(w_n1178_0[1]),.dout(n1225),.clk(gclk));
	jxor g1162(.dina(w_n1225_0[1]),.dinb(w_n1176_0[1]),.dout(n1226),.clk(gclk));
	jxor g1163(.dina(w_n1226_0[1]),.dinb(w_n1173_0[1]),.dout(n1227),.clk(gclk));
	jxor g1164(.dina(w_n1227_0[1]),.dinb(w_n1171_0[1]),.dout(n1228),.clk(gclk));
	jxor g1165(.dina(w_n1228_0[1]),.dinb(w_n1168_0[1]),.dout(n1229),.clk(gclk));
	jxor g1166(.dina(w_n1229_0[1]),.dinb(w_n1166_0[1]),.dout(n1230),.clk(gclk));
	jxor g1167(.dina(w_n1230_0[1]),.dinb(w_n1163_0[1]),.dout(n1231),.clk(gclk));
	jxor g1168(.dina(w_n1231_0[1]),.dinb(w_n1161_0[1]),.dout(n1232),.clk(gclk));
	jxor g1169(.dina(w_n1232_0[1]),.dinb(w_n1158_0[1]),.dout(n1233),.clk(gclk));
	jnot g1170(.din(n1233),.dout(n1234),.clk(gclk));
	jxor g1171(.dina(w_n1234_0[1]),.dinb(w_n1156_0[1]),.dout(n1235),.clk(gclk));
	jnot g1172(.din(n1235),.dout(n1236),.clk(gclk));
	jxor g1173(.dina(w_n1236_0[1]),.dinb(w_n1152_0[1]),.dout(n1237),.clk(gclk));
	jxor g1174(.dina(w_n1237_0[1]),.dinb(w_n1151_0[1]),.dout(n1238),.clk(gclk));
	jnot g1175(.din(w_n1238_0[1]),.dout(n1239),.clk(gclk));
	jxor g1176(.dina(n1239),.dinb(w_n1147_0[1]),.dout(w_dff_A_MsaMqHPq5_2),.clk(gclk));
	jnot g1177(.din(w_n1237_0[0]),.dout(n1241),.clk(gclk));
	jor g1178(.dina(n1241),.dinb(w_n1151_0[0]),.dout(n1242),.clk(gclk));
	jor g1179(.dina(w_n1238_0[0]),.dinb(w_n1147_0[0]),.dout(n1243),.clk(gclk));
	jand g1180(.dina(n1243),.dinb(w_dff_B_nG2AdicV6_1),.dout(n1244),.clk(gclk));
	jor g1181(.dina(w_n1234_0[0]),.dinb(w_n1156_0[0]),.dout(n1245),.clk(gclk));
	jor g1182(.dina(w_n1236_0[0]),.dinb(w_n1152_0[0]),.dout(n1246),.clk(gclk));
	jand g1183(.dina(n1246),.dinb(n1245),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1231_0[0]),.dinb(w_n1161_0[0]),.dout(n1249),.clk(gclk));
	jand g1186(.dina(w_n1232_0[0]),.dinb(w_n1158_0[0]),.dout(n1250),.clk(gclk));
	jor g1187(.dina(n1250),.dinb(n1249),.dout(n1251),.clk(gclk));
	jand g1188(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1252),.clk(gclk));
	jnot g1189(.din(n1252),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1229_0[0]),.dinb(w_n1166_0[0]),.dout(n1254),.clk(gclk));
	jand g1191(.dina(w_n1230_0[0]),.dinb(w_n1163_0[0]),.dout(n1255),.clk(gclk));
	jor g1192(.dina(n1255),.dinb(n1254),.dout(n1256),.clk(gclk));
	jand g1193(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1257),.clk(gclk));
	jnot g1194(.din(n1257),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1227_0[0]),.dinb(w_n1171_0[0]),.dout(n1259),.clk(gclk));
	jand g1196(.dina(w_n1228_0[0]),.dinb(w_n1168_0[0]),.dout(n1260),.clk(gclk));
	jor g1197(.dina(n1260),.dinb(n1259),.dout(n1261),.clk(gclk));
	jand g1198(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1262),.clk(gclk));
	jnot g1199(.din(n1262),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1225_0[0]),.dinb(w_n1176_0[0]),.dout(n1264),.clk(gclk));
	jand g1201(.dina(w_n1226_0[0]),.dinb(w_n1173_0[0]),.dout(n1265),.clk(gclk));
	jor g1202(.dina(n1265),.dinb(n1264),.dout(n1266),.clk(gclk));
	jand g1203(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1267),.clk(gclk));
	jnot g1204(.din(n1267),.dout(n1268),.clk(gclk));
	jand g1205(.dina(w_n1223_0[0]),.dinb(w_n1181_0[0]),.dout(n1269),.clk(gclk));
	jand g1206(.dina(w_n1224_0[0]),.dinb(w_n1178_0[0]),.dout(n1270),.clk(gclk));
	jor g1207(.dina(n1270),.dinb(n1269),.dout(n1271),.clk(gclk));
	jand g1208(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1272),.clk(gclk));
	jnot g1209(.din(n1272),.dout(n1273),.clk(gclk));
	jand g1210(.dina(w_n1221_0[0]),.dinb(w_n1186_0[0]),.dout(n1274),.clk(gclk));
	jand g1211(.dina(w_n1222_0[0]),.dinb(w_n1183_0[0]),.dout(n1275),.clk(gclk));
	jor g1212(.dina(n1275),.dinb(n1274),.dout(n1276),.clk(gclk));
	jand g1213(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1277),.clk(gclk));
	jnot g1214(.din(n1277),.dout(n1278),.clk(gclk));
	jand g1215(.dina(w_n1219_0[0]),.dinb(w_n1191_0[0]),.dout(n1279),.clk(gclk));
	jand g1216(.dina(w_n1220_0[0]),.dinb(w_n1188_0[0]),.dout(n1280),.clk(gclk));
	jor g1217(.dina(n1280),.dinb(n1279),.dout(n1281),.clk(gclk));
	jand g1218(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1282),.clk(gclk));
	jnot g1219(.din(n1282),.dout(n1283),.clk(gclk));
	jand g1220(.dina(w_n1217_0[0]),.dinb(w_n1196_0[0]),.dout(n1284),.clk(gclk));
	jand g1221(.dina(w_n1218_0[0]),.dinb(w_n1193_0[0]),.dout(n1285),.clk(gclk));
	jor g1222(.dina(n1285),.dinb(n1284),.dout(n1286),.clk(gclk));
	jand g1223(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1287),.clk(gclk));
	jnot g1224(.din(n1287),.dout(n1288),.clk(gclk));
	jand g1225(.dina(w_n1215_0[0]),.dinb(w_n1201_0[0]),.dout(n1289),.clk(gclk));
	jand g1226(.dina(w_n1216_0[0]),.dinb(w_n1198_0[0]),.dout(n1290),.clk(gclk));
	jor g1227(.dina(n1290),.dinb(n1289),.dout(n1291),.clk(gclk));
	jand g1228(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jand g1230(.dina(w_n1213_0[0]),.dinb(w_n1206_0[0]),.dout(n1294),.clk(gclk));
	jand g1231(.dina(w_n1214_0[0]),.dinb(w_n1203_0[0]),.dout(n1295),.clk(gclk));
	jor g1232(.dina(n1295),.dinb(n1294),.dout(n1296),.clk(gclk));
	jand g1233(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1297),.clk(gclk));
	jand g1234(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1298),.clk(gclk));
	jor g1235(.dina(w_n1210_0[0]),.dinb(w_n1208_0[0]),.dout(n1299),.clk(gclk));
	jor g1236(.dina(w_n1212_0[0]),.dinb(w_n1207_0[0]),.dout(n1300),.clk(gclk));
	jand g1237(.dina(n1300),.dinb(n1299),.dout(n1301),.clk(gclk));
	jxor g1238(.dina(w_n1301_0[1]),.dinb(w_n1298_0[1]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(n1302),.dout(n1303),.clk(gclk));
	jxor g1240(.dina(w_n1303_0[1]),.dinb(w_n1297_0[1]),.dout(n1304),.clk(gclk));
	jxor g1241(.dina(w_n1304_0[1]),.dinb(w_n1296_0[1]),.dout(n1305),.clk(gclk));
	jxor g1242(.dina(w_n1305_0[1]),.dinb(w_n1293_0[1]),.dout(n1306),.clk(gclk));
	jxor g1243(.dina(w_n1306_0[1]),.dinb(w_n1291_0[1]),.dout(n1307),.clk(gclk));
	jxor g1244(.dina(w_n1307_0[1]),.dinb(w_n1288_0[1]),.dout(n1308),.clk(gclk));
	jxor g1245(.dina(w_n1308_0[1]),.dinb(w_n1286_0[1]),.dout(n1309),.clk(gclk));
	jxor g1246(.dina(w_n1309_0[1]),.dinb(w_n1283_0[1]),.dout(n1310),.clk(gclk));
	jxor g1247(.dina(w_n1310_0[1]),.dinb(w_n1281_0[1]),.dout(n1311),.clk(gclk));
	jxor g1248(.dina(w_n1311_0[1]),.dinb(w_n1278_0[1]),.dout(n1312),.clk(gclk));
	jxor g1249(.dina(w_n1312_0[1]),.dinb(w_n1276_0[1]),.dout(n1313),.clk(gclk));
	jxor g1250(.dina(w_n1313_0[1]),.dinb(w_n1273_0[1]),.dout(n1314),.clk(gclk));
	jxor g1251(.dina(w_n1314_0[1]),.dinb(w_n1271_0[1]),.dout(n1315),.clk(gclk));
	jxor g1252(.dina(w_n1315_0[1]),.dinb(w_n1268_0[1]),.dout(n1316),.clk(gclk));
	jxor g1253(.dina(w_n1316_0[1]),.dinb(w_n1266_0[1]),.dout(n1317),.clk(gclk));
	jxor g1254(.dina(w_n1317_0[1]),.dinb(w_n1263_0[1]),.dout(n1318),.clk(gclk));
	jxor g1255(.dina(w_n1318_0[1]),.dinb(w_n1261_0[1]),.dout(n1319),.clk(gclk));
	jxor g1256(.dina(w_n1319_0[1]),.dinb(w_n1258_0[1]),.dout(n1320),.clk(gclk));
	jxor g1257(.dina(w_n1320_0[1]),.dinb(w_n1256_0[1]),.dout(n1321),.clk(gclk));
	jxor g1258(.dina(w_n1321_0[1]),.dinb(w_n1253_0[1]),.dout(n1322),.clk(gclk));
	jxor g1259(.dina(w_n1322_0[1]),.dinb(w_n1251_0[1]),.dout(n1323),.clk(gclk));
	jnot g1260(.din(n1323),.dout(n1324),.clk(gclk));
	jxor g1261(.dina(w_n1324_0[1]),.dinb(w_n1248_0[1]),.dout(n1325),.clk(gclk));
	jxor g1262(.dina(w_n1325_0[1]),.dinb(w_n1247_0[1]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(w_n1326_0[1]),.dout(n1327),.clk(gclk));
	jxor g1264(.dina(w_dff_B_lQr3XVAK2_0),.dinb(w_n1244_0[1]),.dout(w_dff_A_2H3dPpHv5_2),.clk(gclk));
	jnot g1265(.din(w_n1325_0[0]),.dout(n1329),.clk(gclk));
	jor g1266(.dina(n1329),.dinb(w_n1247_0[0]),.dout(n1330),.clk(gclk));
	jor g1267(.dina(w_n1326_0[0]),.dinb(w_n1244_0[0]),.dout(n1331),.clk(gclk));
	jand g1268(.dina(n1331),.dinb(w_dff_B_AURzPvBv7_1),.dout(n1332),.clk(gclk));
	jnot g1269(.din(w_n1251_0[0]),.dout(n1333),.clk(gclk));
	jnot g1270(.din(w_n1322_0[0]),.dout(n1334),.clk(gclk));
	jor g1271(.dina(n1334),.dinb(n1333),.dout(n1335),.clk(gclk));
	jor g1272(.dina(w_n1324_0[0]),.dinb(w_n1248_0[0]),.dout(n1336),.clk(gclk));
	jand g1273(.dina(n1336),.dinb(n1335),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1320_0[0]),.dinb(w_n1256_0[0]),.dout(n1339),.clk(gclk));
	jand g1276(.dina(w_n1321_0[0]),.dinb(w_n1253_0[0]),.dout(n1340),.clk(gclk));
	jor g1277(.dina(n1340),.dinb(n1339),.dout(n1341),.clk(gclk));
	jand g1278(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1342),.clk(gclk));
	jnot g1279(.din(n1342),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1318_0[0]),.dinb(w_n1261_0[0]),.dout(n1344),.clk(gclk));
	jand g1281(.dina(w_n1319_0[0]),.dinb(w_n1258_0[0]),.dout(n1345),.clk(gclk));
	jor g1282(.dina(n1345),.dinb(n1344),.dout(n1346),.clk(gclk));
	jand g1283(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1347),.clk(gclk));
	jnot g1284(.din(n1347),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1316_0[0]),.dinb(w_n1266_0[0]),.dout(n1349),.clk(gclk));
	jand g1286(.dina(w_n1317_0[0]),.dinb(w_n1263_0[0]),.dout(n1350),.clk(gclk));
	jor g1287(.dina(n1350),.dinb(n1349),.dout(n1351),.clk(gclk));
	jand g1288(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1352),.clk(gclk));
	jnot g1289(.din(n1352),.dout(n1353),.clk(gclk));
	jand g1290(.dina(w_n1314_0[0]),.dinb(w_n1271_0[0]),.dout(n1354),.clk(gclk));
	jand g1291(.dina(w_n1315_0[0]),.dinb(w_n1268_0[0]),.dout(n1355),.clk(gclk));
	jor g1292(.dina(n1355),.dinb(n1354),.dout(n1356),.clk(gclk));
	jand g1293(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1357),.clk(gclk));
	jnot g1294(.din(n1357),.dout(n1358),.clk(gclk));
	jand g1295(.dina(w_n1312_0[0]),.dinb(w_n1276_0[0]),.dout(n1359),.clk(gclk));
	jand g1296(.dina(w_n1313_0[0]),.dinb(w_n1273_0[0]),.dout(n1360),.clk(gclk));
	jor g1297(.dina(n1360),.dinb(n1359),.dout(n1361),.clk(gclk));
	jand g1298(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1362),.clk(gclk));
	jnot g1299(.din(n1362),.dout(n1363),.clk(gclk));
	jand g1300(.dina(w_n1310_0[0]),.dinb(w_n1281_0[0]),.dout(n1364),.clk(gclk));
	jand g1301(.dina(w_n1311_0[0]),.dinb(w_n1278_0[0]),.dout(n1365),.clk(gclk));
	jor g1302(.dina(n1365),.dinb(n1364),.dout(n1366),.clk(gclk));
	jand g1303(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1367),.clk(gclk));
	jnot g1304(.din(n1367),.dout(n1368),.clk(gclk));
	jand g1305(.dina(w_n1308_0[0]),.dinb(w_n1286_0[0]),.dout(n1369),.clk(gclk));
	jand g1306(.dina(w_n1309_0[0]),.dinb(w_n1283_0[0]),.dout(n1370),.clk(gclk));
	jor g1307(.dina(n1370),.dinb(n1369),.dout(n1371),.clk(gclk));
	jand g1308(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1372),.clk(gclk));
	jnot g1309(.din(n1372),.dout(n1373),.clk(gclk));
	jand g1310(.dina(w_n1306_0[0]),.dinb(w_n1291_0[0]),.dout(n1374),.clk(gclk));
	jand g1311(.dina(w_n1307_0[0]),.dinb(w_n1288_0[0]),.dout(n1375),.clk(gclk));
	jor g1312(.dina(n1375),.dinb(n1374),.dout(n1376),.clk(gclk));
	jand g1313(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jand g1315(.dina(w_n1304_0[0]),.dinb(w_n1296_0[0]),.dout(n1379),.clk(gclk));
	jand g1316(.dina(w_n1305_0[0]),.dinb(w_n1293_0[0]),.dout(n1380),.clk(gclk));
	jor g1317(.dina(n1380),.dinb(n1379),.dout(n1381),.clk(gclk));
	jand g1318(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1382),.clk(gclk));
	jand g1319(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1383),.clk(gclk));
	jor g1320(.dina(w_n1301_0[0]),.dinb(w_n1298_0[0]),.dout(n1384),.clk(gclk));
	jor g1321(.dina(w_n1303_0[0]),.dinb(w_n1297_0[0]),.dout(n1385),.clk(gclk));
	jand g1322(.dina(n1385),.dinb(n1384),.dout(n1386),.clk(gclk));
	jxor g1323(.dina(w_n1386_0[1]),.dinb(w_n1383_0[1]),.dout(n1387),.clk(gclk));
	jnot g1324(.din(n1387),.dout(n1388),.clk(gclk));
	jxor g1325(.dina(w_n1388_0[1]),.dinb(w_n1382_0[1]),.dout(n1389),.clk(gclk));
	jxor g1326(.dina(w_n1389_0[1]),.dinb(w_n1381_0[1]),.dout(n1390),.clk(gclk));
	jxor g1327(.dina(w_n1390_0[1]),.dinb(w_n1378_0[1]),.dout(n1391),.clk(gclk));
	jxor g1328(.dina(w_n1391_0[1]),.dinb(w_n1376_0[1]),.dout(n1392),.clk(gclk));
	jxor g1329(.dina(w_n1392_0[1]),.dinb(w_n1373_0[1]),.dout(n1393),.clk(gclk));
	jxor g1330(.dina(w_n1393_0[1]),.dinb(w_n1371_0[1]),.dout(n1394),.clk(gclk));
	jxor g1331(.dina(w_n1394_0[1]),.dinb(w_n1368_0[1]),.dout(n1395),.clk(gclk));
	jxor g1332(.dina(w_n1395_0[1]),.dinb(w_n1366_0[1]),.dout(n1396),.clk(gclk));
	jxor g1333(.dina(w_n1396_0[1]),.dinb(w_n1363_0[1]),.dout(n1397),.clk(gclk));
	jxor g1334(.dina(w_n1397_0[1]),.dinb(w_n1361_0[1]),.dout(n1398),.clk(gclk));
	jxor g1335(.dina(w_n1398_0[1]),.dinb(w_n1358_0[1]),.dout(n1399),.clk(gclk));
	jxor g1336(.dina(w_n1399_0[1]),.dinb(w_n1356_0[1]),.dout(n1400),.clk(gclk));
	jxor g1337(.dina(w_n1400_0[1]),.dinb(w_n1353_0[1]),.dout(n1401),.clk(gclk));
	jxor g1338(.dina(w_n1401_0[1]),.dinb(w_n1351_0[1]),.dout(n1402),.clk(gclk));
	jxor g1339(.dina(w_n1402_0[1]),.dinb(w_n1348_0[1]),.dout(n1403),.clk(gclk));
	jxor g1340(.dina(w_n1403_0[1]),.dinb(w_n1346_0[1]),.dout(n1404),.clk(gclk));
	jxor g1341(.dina(w_n1404_0[1]),.dinb(w_n1343_0[1]),.dout(n1405),.clk(gclk));
	jxor g1342(.dina(w_n1405_0[1]),.dinb(w_n1341_0[1]),.dout(n1406),.clk(gclk));
	jnot g1343(.din(n1406),.dout(n1407),.clk(gclk));
	jxor g1344(.dina(w_n1407_0[1]),.dinb(w_n1338_0[1]),.dout(n1408),.clk(gclk));
	jnot g1345(.din(n1408),.dout(n1409),.clk(gclk));
	jxor g1346(.dina(w_n1409_0[1]),.dinb(w_n1337_0[1]),.dout(n1410),.clk(gclk));
	jxor g1347(.dina(w_n1410_0[1]),.dinb(w_n1332_0[1]),.dout(w_dff_A_nFZwUN7m5_2),.clk(gclk));
	jor g1348(.dina(w_n1409_0[0]),.dinb(w_n1337_0[0]),.dout(n1412),.clk(gclk));
	jnot g1349(.din(w_n1410_0[0]),.dout(n1413),.clk(gclk));
	jor g1350(.dina(w_dff_B_FsUF8c9E3_0),.dinb(w_n1332_0[0]),.dout(n1414),.clk(gclk));
	jand g1351(.dina(n1414),.dinb(w_dff_B_lqat5rQz4_1),.dout(n1415),.clk(gclk));
	jnot g1352(.din(w_n1341_0[0]),.dout(n1416),.clk(gclk));
	jnot g1353(.din(w_n1405_0[0]),.dout(n1417),.clk(gclk));
	jor g1354(.dina(n1417),.dinb(n1416),.dout(n1418),.clk(gclk));
	jor g1355(.dina(w_n1407_0[0]),.dinb(w_n1338_0[0]),.dout(n1419),.clk(gclk));
	jand g1356(.dina(n1419),.dinb(n1418),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1403_0[0]),.dinb(w_n1346_0[0]),.dout(n1422),.clk(gclk));
	jand g1359(.dina(w_n1404_0[0]),.dinb(w_n1343_0[0]),.dout(n1423),.clk(gclk));
	jor g1360(.dina(n1423),.dinb(n1422),.dout(n1424),.clk(gclk));
	jand g1361(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1425),.clk(gclk));
	jnot g1362(.din(n1425),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1401_0[0]),.dinb(w_n1351_0[0]),.dout(n1427),.clk(gclk));
	jand g1364(.dina(w_n1402_0[0]),.dinb(w_n1348_0[0]),.dout(n1428),.clk(gclk));
	jor g1365(.dina(n1428),.dinb(n1427),.dout(n1429),.clk(gclk));
	jand g1366(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1430),.clk(gclk));
	jnot g1367(.din(n1430),.dout(n1431),.clk(gclk));
	jand g1368(.dina(w_n1399_0[0]),.dinb(w_n1356_0[0]),.dout(n1432),.clk(gclk));
	jand g1369(.dina(w_n1400_0[0]),.dinb(w_n1353_0[0]),.dout(n1433),.clk(gclk));
	jor g1370(.dina(n1433),.dinb(n1432),.dout(n1434),.clk(gclk));
	jand g1371(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1435),.clk(gclk));
	jnot g1372(.din(n1435),.dout(n1436),.clk(gclk));
	jand g1373(.dina(w_n1397_0[0]),.dinb(w_n1361_0[0]),.dout(n1437),.clk(gclk));
	jand g1374(.dina(w_n1398_0[0]),.dinb(w_n1358_0[0]),.dout(n1438),.clk(gclk));
	jor g1375(.dina(n1438),.dinb(n1437),.dout(n1439),.clk(gclk));
	jand g1376(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1440),.clk(gclk));
	jnot g1377(.din(n1440),.dout(n1441),.clk(gclk));
	jand g1378(.dina(w_n1395_0[0]),.dinb(w_n1366_0[0]),.dout(n1442),.clk(gclk));
	jand g1379(.dina(w_n1396_0[0]),.dinb(w_n1363_0[0]),.dout(n1443),.clk(gclk));
	jor g1380(.dina(n1443),.dinb(n1442),.dout(n1444),.clk(gclk));
	jand g1381(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1445),.clk(gclk));
	jnot g1382(.din(n1445),.dout(n1446),.clk(gclk));
	jand g1383(.dina(w_n1393_0[0]),.dinb(w_n1371_0[0]),.dout(n1447),.clk(gclk));
	jand g1384(.dina(w_n1394_0[0]),.dinb(w_n1368_0[0]),.dout(n1448),.clk(gclk));
	jor g1385(.dina(n1448),.dinb(n1447),.dout(n1449),.clk(gclk));
	jand g1386(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1450),.clk(gclk));
	jnot g1387(.din(n1450),.dout(n1451),.clk(gclk));
	jand g1388(.dina(w_n1391_0[0]),.dinb(w_n1376_0[0]),.dout(n1452),.clk(gclk));
	jand g1389(.dina(w_n1392_0[0]),.dinb(w_n1373_0[0]),.dout(n1453),.clk(gclk));
	jor g1390(.dina(n1453),.dinb(n1452),.dout(n1454),.clk(gclk));
	jand g1391(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1455),.clk(gclk));
	jnot g1392(.din(n1455),.dout(n1456),.clk(gclk));
	jand g1393(.dina(w_n1389_0[0]),.dinb(w_n1381_0[0]),.dout(n1457),.clk(gclk));
	jand g1394(.dina(w_n1390_0[0]),.dinb(w_n1378_0[0]),.dout(n1458),.clk(gclk));
	jor g1395(.dina(n1458),.dinb(n1457),.dout(n1459),.clk(gclk));
	jand g1396(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1460),.clk(gclk));
	jand g1397(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1461),.clk(gclk));
	jor g1398(.dina(w_n1386_0[0]),.dinb(w_n1383_0[0]),.dout(n1462),.clk(gclk));
	jor g1399(.dina(w_n1388_0[0]),.dinb(w_n1382_0[0]),.dout(n1463),.clk(gclk));
	jand g1400(.dina(n1463),.dinb(n1462),.dout(n1464),.clk(gclk));
	jxor g1401(.dina(w_n1464_0[1]),.dinb(w_n1461_0[1]),.dout(n1465),.clk(gclk));
	jnot g1402(.din(n1465),.dout(n1466),.clk(gclk));
	jxor g1403(.dina(w_n1466_0[1]),.dinb(w_n1460_0[1]),.dout(n1467),.clk(gclk));
	jxor g1404(.dina(w_n1467_0[1]),.dinb(w_n1459_0[1]),.dout(n1468),.clk(gclk));
	jxor g1405(.dina(w_n1468_0[1]),.dinb(w_n1456_0[1]),.dout(n1469),.clk(gclk));
	jxor g1406(.dina(w_n1469_0[1]),.dinb(w_n1454_0[1]),.dout(n1470),.clk(gclk));
	jxor g1407(.dina(w_n1470_0[1]),.dinb(w_n1451_0[1]),.dout(n1471),.clk(gclk));
	jxor g1408(.dina(w_n1471_0[1]),.dinb(w_n1449_0[1]),.dout(n1472),.clk(gclk));
	jxor g1409(.dina(w_n1472_0[1]),.dinb(w_n1446_0[1]),.dout(n1473),.clk(gclk));
	jxor g1410(.dina(w_n1473_0[1]),.dinb(w_n1444_0[1]),.dout(n1474),.clk(gclk));
	jxor g1411(.dina(w_n1474_0[1]),.dinb(w_n1441_0[1]),.dout(n1475),.clk(gclk));
	jxor g1412(.dina(w_n1475_0[1]),.dinb(w_n1439_0[1]),.dout(n1476),.clk(gclk));
	jxor g1413(.dina(w_n1476_0[1]),.dinb(w_n1436_0[1]),.dout(n1477),.clk(gclk));
	jxor g1414(.dina(w_n1477_0[1]),.dinb(w_n1434_0[1]),.dout(n1478),.clk(gclk));
	jxor g1415(.dina(w_n1478_0[1]),.dinb(w_n1431_0[1]),.dout(n1479),.clk(gclk));
	jxor g1416(.dina(w_n1479_0[1]),.dinb(w_n1429_0[1]),.dout(n1480),.clk(gclk));
	jxor g1417(.dina(w_n1480_0[1]),.dinb(w_n1426_0[1]),.dout(n1481),.clk(gclk));
	jxor g1418(.dina(w_n1481_0[1]),.dinb(w_n1424_0[1]),.dout(n1482),.clk(gclk));
	jnot g1419(.din(n1482),.dout(n1483),.clk(gclk));
	jxor g1420(.dina(w_n1483_0[1]),.dinb(w_n1421_0[1]),.dout(n1484),.clk(gclk));
	jnot g1421(.din(n1484),.dout(n1485),.clk(gclk));
	jxor g1422(.dina(w_n1485_0[1]),.dinb(w_n1420_0[1]),.dout(n1486),.clk(gclk));
	jxor g1423(.dina(w_n1486_0[1]),.dinb(w_n1415_0[1]),.dout(w_dff_A_BTnUMnAU7_2),.clk(gclk));
	jor g1424(.dina(w_n1485_0[0]),.dinb(w_n1420_0[0]),.dout(n1488),.clk(gclk));
	jnot g1425(.din(w_n1486_0[0]),.dout(n1489),.clk(gclk));
	jor g1426(.dina(w_dff_B_6uiefIB11_0),.dinb(w_n1415_0[0]),.dout(n1490),.clk(gclk));
	jand g1427(.dina(n1490),.dinb(w_dff_B_nLY9nNaa0_1),.dout(n1491),.clk(gclk));
	jnot g1428(.din(w_n1424_0[0]),.dout(n1492),.clk(gclk));
	jnot g1429(.din(w_n1481_0[0]),.dout(n1493),.clk(gclk));
	jor g1430(.dina(n1493),.dinb(n1492),.dout(n1494),.clk(gclk));
	jor g1431(.dina(w_n1483_0[0]),.dinb(w_n1421_0[0]),.dout(n1495),.clk(gclk));
	jand g1432(.dina(n1495),.dinb(n1494),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1479_0[0]),.dinb(w_n1429_0[0]),.dout(n1498),.clk(gclk));
	jand g1435(.dina(w_n1480_0[0]),.dinb(w_n1426_0[0]),.dout(n1499),.clk(gclk));
	jor g1436(.dina(n1499),.dinb(n1498),.dout(n1500),.clk(gclk));
	jand g1437(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1501),.clk(gclk));
	jnot g1438(.din(n1501),.dout(n1502),.clk(gclk));
	jand g1439(.dina(w_n1477_0[0]),.dinb(w_n1434_0[0]),.dout(n1503),.clk(gclk));
	jand g1440(.dina(w_n1478_0[0]),.dinb(w_n1431_0[0]),.dout(n1504),.clk(gclk));
	jor g1441(.dina(n1504),.dinb(n1503),.dout(n1505),.clk(gclk));
	jand g1442(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1506),.clk(gclk));
	jnot g1443(.din(n1506),.dout(n1507),.clk(gclk));
	jand g1444(.dina(w_n1475_0[0]),.dinb(w_n1439_0[0]),.dout(n1508),.clk(gclk));
	jand g1445(.dina(w_n1476_0[0]),.dinb(w_n1436_0[0]),.dout(n1509),.clk(gclk));
	jor g1446(.dina(n1509),.dinb(n1508),.dout(n1510),.clk(gclk));
	jand g1447(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1511),.clk(gclk));
	jnot g1448(.din(n1511),.dout(n1512),.clk(gclk));
	jand g1449(.dina(w_n1473_0[0]),.dinb(w_n1444_0[0]),.dout(n1513),.clk(gclk));
	jand g1450(.dina(w_n1474_0[0]),.dinb(w_n1441_0[0]),.dout(n1514),.clk(gclk));
	jor g1451(.dina(n1514),.dinb(n1513),.dout(n1515),.clk(gclk));
	jand g1452(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1516),.clk(gclk));
	jnot g1453(.din(n1516),.dout(n1517),.clk(gclk));
	jand g1454(.dina(w_n1471_0[0]),.dinb(w_n1449_0[0]),.dout(n1518),.clk(gclk));
	jand g1455(.dina(w_n1472_0[0]),.dinb(w_n1446_0[0]),.dout(n1519),.clk(gclk));
	jor g1456(.dina(n1519),.dinb(n1518),.dout(n1520),.clk(gclk));
	jand g1457(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1521),.clk(gclk));
	jnot g1458(.din(n1521),.dout(n1522),.clk(gclk));
	jand g1459(.dina(w_n1469_0[0]),.dinb(w_n1454_0[0]),.dout(n1523),.clk(gclk));
	jand g1460(.dina(w_n1470_0[0]),.dinb(w_n1451_0[0]),.dout(n1524),.clk(gclk));
	jor g1461(.dina(n1524),.dinb(n1523),.dout(n1525),.clk(gclk));
	jand g1462(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1526),.clk(gclk));
	jnot g1463(.din(n1526),.dout(n1527),.clk(gclk));
	jand g1464(.dina(w_n1467_0[0]),.dinb(w_n1459_0[0]),.dout(n1528),.clk(gclk));
	jand g1465(.dina(w_n1468_0[0]),.dinb(w_n1456_0[0]),.dout(n1529),.clk(gclk));
	jor g1466(.dina(n1529),.dinb(n1528),.dout(n1530),.clk(gclk));
	jand g1467(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1531),.clk(gclk));
	jand g1468(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1532),.clk(gclk));
	jor g1469(.dina(w_n1464_0[0]),.dinb(w_n1461_0[0]),.dout(n1533),.clk(gclk));
	jor g1470(.dina(w_n1466_0[0]),.dinb(w_n1460_0[0]),.dout(n1534),.clk(gclk));
	jand g1471(.dina(n1534),.dinb(n1533),.dout(n1535),.clk(gclk));
	jxor g1472(.dina(w_n1535_0[1]),.dinb(w_n1532_0[1]),.dout(n1536),.clk(gclk));
	jnot g1473(.din(n1536),.dout(n1537),.clk(gclk));
	jxor g1474(.dina(w_n1537_0[1]),.dinb(w_n1531_0[1]),.dout(n1538),.clk(gclk));
	jxor g1475(.dina(w_n1538_0[1]),.dinb(w_n1530_0[1]),.dout(n1539),.clk(gclk));
	jxor g1476(.dina(w_n1539_0[1]),.dinb(w_n1527_0[1]),.dout(n1540),.clk(gclk));
	jxor g1477(.dina(w_n1540_0[1]),.dinb(w_n1525_0[1]),.dout(n1541),.clk(gclk));
	jxor g1478(.dina(w_n1541_0[1]),.dinb(w_n1522_0[1]),.dout(n1542),.clk(gclk));
	jxor g1479(.dina(w_n1542_0[1]),.dinb(w_n1520_0[1]),.dout(n1543),.clk(gclk));
	jxor g1480(.dina(w_n1543_0[1]),.dinb(w_n1517_0[1]),.dout(n1544),.clk(gclk));
	jxor g1481(.dina(w_n1544_0[1]),.dinb(w_n1515_0[1]),.dout(n1545),.clk(gclk));
	jxor g1482(.dina(w_n1545_0[1]),.dinb(w_n1512_0[1]),.dout(n1546),.clk(gclk));
	jxor g1483(.dina(w_n1546_0[1]),.dinb(w_n1510_0[1]),.dout(n1547),.clk(gclk));
	jxor g1484(.dina(w_n1547_0[1]),.dinb(w_n1507_0[1]),.dout(n1548),.clk(gclk));
	jxor g1485(.dina(w_n1548_0[1]),.dinb(w_n1505_0[1]),.dout(n1549),.clk(gclk));
	jxor g1486(.dina(w_n1549_0[1]),.dinb(w_n1502_0[1]),.dout(n1550),.clk(gclk));
	jxor g1487(.dina(w_n1550_0[1]),.dinb(w_n1500_0[1]),.dout(n1551),.clk(gclk));
	jnot g1488(.din(n1551),.dout(n1552),.clk(gclk));
	jxor g1489(.dina(w_n1552_0[1]),.dinb(w_n1497_0[1]),.dout(n1553),.clk(gclk));
	jnot g1490(.din(n1553),.dout(n1554),.clk(gclk));
	jxor g1491(.dina(w_n1554_0[1]),.dinb(w_n1496_0[1]),.dout(n1555),.clk(gclk));
	jxor g1492(.dina(w_n1555_0[1]),.dinb(w_n1491_0[1]),.dout(w_dff_A_96BrlB423_2),.clk(gclk));
	jor g1493(.dina(w_n1554_0[0]),.dinb(w_n1496_0[0]),.dout(n1557),.clk(gclk));
	jnot g1494(.din(w_n1555_0[0]),.dout(n1558),.clk(gclk));
	jor g1495(.dina(w_dff_B_GiR5nEIQ5_0),.dinb(w_n1491_0[0]),.dout(n1559),.clk(gclk));
	jand g1496(.dina(n1559),.dinb(w_dff_B_ykjfpplL7_1),.dout(n1560),.clk(gclk));
	jnot g1497(.din(w_n1500_0[0]),.dout(n1561),.clk(gclk));
	jnot g1498(.din(w_n1550_0[0]),.dout(n1562),.clk(gclk));
	jor g1499(.dina(n1562),.dinb(n1561),.dout(n1563),.clk(gclk));
	jor g1500(.dina(w_n1552_0[0]),.dinb(w_n1497_0[0]),.dout(n1564),.clk(gclk));
	jand g1501(.dina(n1564),.dinb(n1563),.dout(n1565),.clk(gclk));
	jand g1502(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1566),.clk(gclk));
	jand g1503(.dina(w_n1548_0[0]),.dinb(w_n1505_0[0]),.dout(n1567),.clk(gclk));
	jand g1504(.dina(w_n1549_0[0]),.dinb(w_n1502_0[0]),.dout(n1568),.clk(gclk));
	jor g1505(.dina(n1568),.dinb(n1567),.dout(n1569),.clk(gclk));
	jand g1506(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1570),.clk(gclk));
	jnot g1507(.din(n1570),.dout(n1571),.clk(gclk));
	jand g1508(.dina(w_n1546_0[0]),.dinb(w_n1510_0[0]),.dout(n1572),.clk(gclk));
	jand g1509(.dina(w_n1547_0[0]),.dinb(w_n1507_0[0]),.dout(n1573),.clk(gclk));
	jor g1510(.dina(n1573),.dinb(n1572),.dout(n1574),.clk(gclk));
	jand g1511(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1575),.clk(gclk));
	jnot g1512(.din(n1575),.dout(n1576),.clk(gclk));
	jand g1513(.dina(w_n1544_0[0]),.dinb(w_n1515_0[0]),.dout(n1577),.clk(gclk));
	jand g1514(.dina(w_n1545_0[0]),.dinb(w_n1512_0[0]),.dout(n1578),.clk(gclk));
	jor g1515(.dina(n1578),.dinb(n1577),.dout(n1579),.clk(gclk));
	jand g1516(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1580),.clk(gclk));
	jnot g1517(.din(n1580),.dout(n1581),.clk(gclk));
	jand g1518(.dina(w_n1542_0[0]),.dinb(w_n1520_0[0]),.dout(n1582),.clk(gclk));
	jand g1519(.dina(w_n1543_0[0]),.dinb(w_n1517_0[0]),.dout(n1583),.clk(gclk));
	jor g1520(.dina(n1583),.dinb(n1582),.dout(n1584),.clk(gclk));
	jand g1521(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1585),.clk(gclk));
	jnot g1522(.din(n1585),.dout(n1586),.clk(gclk));
	jand g1523(.dina(w_n1540_0[0]),.dinb(w_n1525_0[0]),.dout(n1587),.clk(gclk));
	jand g1524(.dina(w_n1541_0[0]),.dinb(w_n1522_0[0]),.dout(n1588),.clk(gclk));
	jor g1525(.dina(n1588),.dinb(n1587),.dout(n1589),.clk(gclk));
	jand g1526(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1590),.clk(gclk));
	jnot g1527(.din(n1590),.dout(n1591),.clk(gclk));
	jand g1528(.dina(w_n1538_0[0]),.dinb(w_n1530_0[0]),.dout(n1592),.clk(gclk));
	jand g1529(.dina(w_n1539_0[0]),.dinb(w_n1527_0[0]),.dout(n1593),.clk(gclk));
	jor g1530(.dina(n1593),.dinb(n1592),.dout(n1594),.clk(gclk));
	jand g1531(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1595),.clk(gclk));
	jand g1532(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1596),.clk(gclk));
	jor g1533(.dina(w_n1535_0[0]),.dinb(w_n1532_0[0]),.dout(n1597),.clk(gclk));
	jor g1534(.dina(w_n1537_0[0]),.dinb(w_n1531_0[0]),.dout(n1598),.clk(gclk));
	jand g1535(.dina(n1598),.dinb(n1597),.dout(n1599),.clk(gclk));
	jxor g1536(.dina(w_n1599_0[1]),.dinb(w_n1596_0[1]),.dout(n1600),.clk(gclk));
	jnot g1537(.din(n1600),.dout(n1601),.clk(gclk));
	jxor g1538(.dina(w_n1601_0[1]),.dinb(w_n1595_0[1]),.dout(n1602),.clk(gclk));
	jxor g1539(.dina(w_n1602_0[1]),.dinb(w_n1594_0[1]),.dout(n1603),.clk(gclk));
	jxor g1540(.dina(w_n1603_0[1]),.dinb(w_n1591_0[1]),.dout(n1604),.clk(gclk));
	jxor g1541(.dina(w_n1604_0[1]),.dinb(w_n1589_0[1]),.dout(n1605),.clk(gclk));
	jxor g1542(.dina(w_n1605_0[1]),.dinb(w_n1586_0[1]),.dout(n1606),.clk(gclk));
	jxor g1543(.dina(w_n1606_0[1]),.dinb(w_n1584_0[1]),.dout(n1607),.clk(gclk));
	jxor g1544(.dina(w_n1607_0[1]),.dinb(w_n1581_0[1]),.dout(n1608),.clk(gclk));
	jxor g1545(.dina(w_n1608_0[1]),.dinb(w_n1579_0[1]),.dout(n1609),.clk(gclk));
	jxor g1546(.dina(w_n1609_0[1]),.dinb(w_n1576_0[1]),.dout(n1610),.clk(gclk));
	jxor g1547(.dina(w_n1610_0[1]),.dinb(w_n1574_0[1]),.dout(n1611),.clk(gclk));
	jxor g1548(.dina(w_n1611_0[1]),.dinb(w_n1571_0[1]),.dout(n1612),.clk(gclk));
	jxor g1549(.dina(w_n1612_0[1]),.dinb(w_n1569_0[1]),.dout(n1613),.clk(gclk));
	jnot g1550(.din(n1613),.dout(n1614),.clk(gclk));
	jxor g1551(.dina(w_n1614_0[1]),.dinb(w_n1566_0[1]),.dout(n1615),.clk(gclk));
	jnot g1552(.din(n1615),.dout(n1616),.clk(gclk));
	jxor g1553(.dina(w_n1616_0[1]),.dinb(w_n1565_0[1]),.dout(n1617),.clk(gclk));
	jxor g1554(.dina(w_n1617_0[1]),.dinb(w_n1560_0[1]),.dout(w_dff_A_oWs98O0Y7_2),.clk(gclk));
	jor g1555(.dina(w_n1616_0[0]),.dinb(w_n1565_0[0]),.dout(n1619),.clk(gclk));
	jnot g1556(.din(w_n1617_0[0]),.dout(n1620),.clk(gclk));
	jor g1557(.dina(w_dff_B_KPH1H2a54_0),.dinb(w_n1560_0[0]),.dout(n1621),.clk(gclk));
	jand g1558(.dina(n1621),.dinb(w_dff_B_mlg2U20o0_1),.dout(n1622),.clk(gclk));
	jnot g1559(.din(w_n1569_0[0]),.dout(n1623),.clk(gclk));
	jnot g1560(.din(w_n1612_0[0]),.dout(n1624),.clk(gclk));
	jor g1561(.dina(n1624),.dinb(n1623),.dout(n1625),.clk(gclk));
	jor g1562(.dina(w_n1614_0[0]),.dinb(w_n1566_0[0]),.dout(n1626),.clk(gclk));
	jand g1563(.dina(n1626),.dinb(n1625),.dout(n1627),.clk(gclk));
	jand g1564(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1628),.clk(gclk));
	jand g1565(.dina(w_n1610_0[0]),.dinb(w_n1574_0[0]),.dout(n1629),.clk(gclk));
	jand g1566(.dina(w_n1611_0[0]),.dinb(w_n1571_0[0]),.dout(n1630),.clk(gclk));
	jor g1567(.dina(n1630),.dinb(n1629),.dout(n1631),.clk(gclk));
	jand g1568(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1632),.clk(gclk));
	jnot g1569(.din(n1632),.dout(n1633),.clk(gclk));
	jand g1570(.dina(w_n1608_0[0]),.dinb(w_n1579_0[0]),.dout(n1634),.clk(gclk));
	jand g1571(.dina(w_n1609_0[0]),.dinb(w_n1576_0[0]),.dout(n1635),.clk(gclk));
	jor g1572(.dina(n1635),.dinb(n1634),.dout(n1636),.clk(gclk));
	jand g1573(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jand g1575(.dina(w_n1606_0[0]),.dinb(w_n1584_0[0]),.dout(n1639),.clk(gclk));
	jand g1576(.dina(w_n1607_0[0]),.dinb(w_n1581_0[0]),.dout(n1640),.clk(gclk));
	jor g1577(.dina(n1640),.dinb(n1639),.dout(n1641),.clk(gclk));
	jand g1578(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1642),.clk(gclk));
	jnot g1579(.din(n1642),.dout(n1643),.clk(gclk));
	jand g1580(.dina(w_n1604_0[0]),.dinb(w_n1589_0[0]),.dout(n1644),.clk(gclk));
	jand g1581(.dina(w_n1605_0[0]),.dinb(w_n1586_0[0]),.dout(n1645),.clk(gclk));
	jor g1582(.dina(n1645),.dinb(n1644),.dout(n1646),.clk(gclk));
	jand g1583(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(n1647),.dout(n1648),.clk(gclk));
	jand g1585(.dina(w_n1602_0[0]),.dinb(w_n1594_0[0]),.dout(n1649),.clk(gclk));
	jand g1586(.dina(w_n1603_0[0]),.dinb(w_n1591_0[0]),.dout(n1650),.clk(gclk));
	jor g1587(.dina(n1650),.dinb(n1649),.dout(n1651),.clk(gclk));
	jand g1588(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1652),.clk(gclk));
	jand g1589(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1653),.clk(gclk));
	jor g1590(.dina(w_n1599_0[0]),.dinb(w_n1596_0[0]),.dout(n1654),.clk(gclk));
	jor g1591(.dina(w_n1601_0[0]),.dinb(w_n1595_0[0]),.dout(n1655),.clk(gclk));
	jand g1592(.dina(n1655),.dinb(n1654),.dout(n1656),.clk(gclk));
	jxor g1593(.dina(w_n1656_0[1]),.dinb(w_n1653_0[1]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jxor g1595(.dina(w_n1658_0[1]),.dinb(w_n1652_0[1]),.dout(n1659),.clk(gclk));
	jxor g1596(.dina(w_n1659_0[1]),.dinb(w_n1651_0[1]),.dout(n1660),.clk(gclk));
	jxor g1597(.dina(w_n1660_0[1]),.dinb(w_n1648_0[1]),.dout(n1661),.clk(gclk));
	jxor g1598(.dina(w_n1661_0[1]),.dinb(w_n1646_0[1]),.dout(n1662),.clk(gclk));
	jxor g1599(.dina(w_n1662_0[1]),.dinb(w_n1643_0[1]),.dout(n1663),.clk(gclk));
	jxor g1600(.dina(w_n1663_0[1]),.dinb(w_n1641_0[1]),.dout(n1664),.clk(gclk));
	jxor g1601(.dina(w_n1664_0[1]),.dinb(w_n1638_0[1]),.dout(n1665),.clk(gclk));
	jxor g1602(.dina(w_n1665_0[1]),.dinb(w_n1636_0[1]),.dout(n1666),.clk(gclk));
	jxor g1603(.dina(w_n1666_0[1]),.dinb(w_n1633_0[1]),.dout(n1667),.clk(gclk));
	jxor g1604(.dina(w_n1667_0[1]),.dinb(w_n1631_0[1]),.dout(n1668),.clk(gclk));
	jnot g1605(.din(n1668),.dout(n1669),.clk(gclk));
	jxor g1606(.dina(w_n1669_0[1]),.dinb(w_n1628_0[1]),.dout(n1670),.clk(gclk));
	jnot g1607(.din(n1670),.dout(n1671),.clk(gclk));
	jxor g1608(.dina(w_n1671_0[1]),.dinb(w_n1627_0[1]),.dout(n1672),.clk(gclk));
	jxor g1609(.dina(w_n1672_0[1]),.dinb(w_n1622_0[1]),.dout(w_dff_A_IFaEiPVG2_2),.clk(gclk));
	jor g1610(.dina(w_n1671_0[0]),.dinb(w_n1627_0[0]),.dout(n1674),.clk(gclk));
	jnot g1611(.din(w_n1672_0[0]),.dout(n1675),.clk(gclk));
	jor g1612(.dina(w_dff_B_L0Rmnoh95_0),.dinb(w_n1622_0[0]),.dout(n1676),.clk(gclk));
	jand g1613(.dina(n1676),.dinb(w_dff_B_mdApH64o0_1),.dout(n1677),.clk(gclk));
	jnot g1614(.din(w_n1631_0[0]),.dout(n1678),.clk(gclk));
	jnot g1615(.din(w_n1667_0[0]),.dout(n1679),.clk(gclk));
	jor g1616(.dina(n1679),.dinb(n1678),.dout(n1680),.clk(gclk));
	jor g1617(.dina(w_n1669_0[0]),.dinb(w_n1628_0[0]),.dout(n1681),.clk(gclk));
	jand g1618(.dina(n1681),.dinb(n1680),.dout(n1682),.clk(gclk));
	jand g1619(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1683),.clk(gclk));
	jnot g1620(.din(n1683),.dout(n1684),.clk(gclk));
	jand g1621(.dina(w_n1665_0[0]),.dinb(w_n1636_0[0]),.dout(n1685),.clk(gclk));
	jand g1622(.dina(w_n1666_0[0]),.dinb(w_n1633_0[0]),.dout(n1686),.clk(gclk));
	jor g1623(.dina(n1686),.dinb(n1685),.dout(n1687),.clk(gclk));
	jand g1624(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1688),.clk(gclk));
	jnot g1625(.din(n1688),.dout(n1689),.clk(gclk));
	jand g1626(.dina(w_n1663_0[0]),.dinb(w_n1641_0[0]),.dout(n1690),.clk(gclk));
	jand g1627(.dina(w_n1664_0[0]),.dinb(w_n1638_0[0]),.dout(n1691),.clk(gclk));
	jor g1628(.dina(n1691),.dinb(n1690),.dout(n1692),.clk(gclk));
	jand g1629(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1693),.clk(gclk));
	jnot g1630(.din(n1693),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1661_0[0]),.dinb(w_n1646_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1662_0[0]),.dinb(w_n1643_0[0]),.dout(n1696),.clk(gclk));
	jor g1633(.dina(n1696),.dinb(n1695),.dout(n1697),.clk(gclk));
	jand g1634(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1659_0[0]),.dinb(w_n1651_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1660_0[0]),.dinb(w_n1648_0[0]),.dout(n1701),.clk(gclk));
	jor g1638(.dina(n1701),.dinb(n1700),.dout(n1702),.clk(gclk));
	jand g1639(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1703),.clk(gclk));
	jand g1640(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1704),.clk(gclk));
	jor g1641(.dina(w_n1656_0[0]),.dinb(w_n1653_0[0]),.dout(n1705),.clk(gclk));
	jor g1642(.dina(w_n1658_0[0]),.dinb(w_n1652_0[0]),.dout(n1706),.clk(gclk));
	jand g1643(.dina(n1706),.dinb(n1705),.dout(n1707),.clk(gclk));
	jxor g1644(.dina(w_n1707_0[1]),.dinb(w_n1704_0[1]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jxor g1646(.dina(w_n1709_0[1]),.dinb(w_n1703_0[1]),.dout(n1710),.clk(gclk));
	jxor g1647(.dina(w_n1710_0[1]),.dinb(w_n1702_0[1]),.dout(n1711),.clk(gclk));
	jxor g1648(.dina(w_n1711_0[1]),.dinb(w_n1699_0[1]),.dout(n1712),.clk(gclk));
	jxor g1649(.dina(w_n1712_0[1]),.dinb(w_n1697_0[1]),.dout(n1713),.clk(gclk));
	jxor g1650(.dina(w_n1713_0[1]),.dinb(w_n1694_0[1]),.dout(n1714),.clk(gclk));
	jxor g1651(.dina(w_n1714_0[1]),.dinb(w_n1692_0[1]),.dout(n1715),.clk(gclk));
	jxor g1652(.dina(w_n1715_0[1]),.dinb(w_n1689_0[1]),.dout(n1716),.clk(gclk));
	jxor g1653(.dina(w_n1716_0[1]),.dinb(w_n1687_0[1]),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1684_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1682_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1677_0[1]),.dout(w_dff_A_iPM9LwlQ1_2),.clk(gclk));
	jor g1658(.dina(w_n1719_0[0]),.dinb(w_n1682_0[0]),.dout(n1722),.clk(gclk));
	jnot g1659(.din(w_n1720_0[0]),.dout(n1723),.clk(gclk));
	jor g1660(.dina(w_dff_B_JgvJPJc61_0),.dinb(w_n1677_0[0]),.dout(n1724),.clk(gclk));
	jand g1661(.dina(n1724),.dinb(w_dff_B_E0Q23Cbc3_1),.dout(n1725),.clk(gclk));
	jand g1662(.dina(w_n1716_0[0]),.dinb(w_n1687_0[0]),.dout(n1726),.clk(gclk));
	jand g1663(.dina(w_n1717_0[0]),.dinb(w_n1684_0[0]),.dout(n1727),.clk(gclk));
	jor g1664(.dina(n1727),.dinb(n1726),.dout(n1728),.clk(gclk));
	jand g1665(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(n1729),.dout(n1730),.clk(gclk));
	jand g1667(.dina(w_n1714_0[0]),.dinb(w_n1692_0[0]),.dout(n1731),.clk(gclk));
	jand g1668(.dina(w_n1715_0[0]),.dinb(w_n1689_0[0]),.dout(n1732),.clk(gclk));
	jor g1669(.dina(n1732),.dinb(n1731),.dout(n1733),.clk(gclk));
	jand g1670(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1734),.clk(gclk));
	jnot g1671(.din(n1734),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1712_0[0]),.dinb(w_n1697_0[0]),.dout(n1736),.clk(gclk));
	jand g1673(.dina(w_n1713_0[0]),.dinb(w_n1694_0[0]),.dout(n1737),.clk(gclk));
	jor g1674(.dina(n1737),.dinb(n1736),.dout(n1738),.clk(gclk));
	jand g1675(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1739),.clk(gclk));
	jnot g1676(.din(n1739),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1710_0[0]),.dinb(w_n1702_0[0]),.dout(n1741),.clk(gclk));
	jand g1678(.dina(w_n1711_0[0]),.dinb(w_n1699_0[0]),.dout(n1742),.clk(gclk));
	jor g1679(.dina(n1742),.dinb(n1741),.dout(n1743),.clk(gclk));
	jand g1680(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1745),.clk(gclk));
	jor g1682(.dina(w_n1707_0[0]),.dinb(w_n1704_0[0]),.dout(n1746),.clk(gclk));
	jor g1683(.dina(w_n1709_0[0]),.dinb(w_n1703_0[0]),.dout(n1747),.clk(gclk));
	jand g1684(.dina(n1747),.dinb(n1746),.dout(n1748),.clk(gclk));
	jxor g1685(.dina(w_n1748_0[1]),.dinb(w_n1745_0[1]),.dout(n1749),.clk(gclk));
	jnot g1686(.din(n1749),.dout(n1750),.clk(gclk));
	jxor g1687(.dina(w_n1750_0[1]),.dinb(w_n1744_0[1]),.dout(n1751),.clk(gclk));
	jxor g1688(.dina(w_n1751_0[1]),.dinb(w_n1743_0[1]),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1740_0[1]),.dout(n1753),.clk(gclk));
	jxor g1690(.dina(w_n1753_0[1]),.dinb(w_n1738_0[1]),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1735_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1733_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1730_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1728_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1725_0[1]),.dout(w_dff_A_4ZSUinxL1_2),.clk(gclk));
	jnot g1696(.din(w_n1728_0[0]),.dout(n1760),.clk(gclk));
	jnot g1697(.din(w_n1757_0[0]),.dout(n1761),.clk(gclk));
	jor g1698(.dina(n1761),.dinb(n1760),.dout(n1762),.clk(gclk));
	jnot g1699(.din(w_n1758_0[0]),.dout(n1763),.clk(gclk));
	jor g1700(.dina(w_dff_B_EOQdpHEL7_0),.dinb(w_n1725_0[0]),.dout(n1764),.clk(gclk));
	jand g1701(.dina(n1764),.dinb(w_dff_B_kjNYoeB98_1),.dout(n1765),.clk(gclk));
	jand g1702(.dina(w_n1755_0[0]),.dinb(w_n1733_0[0]),.dout(n1766),.clk(gclk));
	jand g1703(.dina(w_n1756_0[0]),.dinb(w_n1730_0[0]),.dout(n1767),.clk(gclk));
	jor g1704(.dina(n1767),.dinb(n1766),.dout(n1768),.clk(gclk));
	jand g1705(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1769),.clk(gclk));
	jnot g1706(.din(n1769),.dout(n1770),.clk(gclk));
	jand g1707(.dina(w_n1753_0[0]),.dinb(w_n1738_0[0]),.dout(n1771),.clk(gclk));
	jand g1708(.dina(w_n1754_0[0]),.dinb(w_n1735_0[0]),.dout(n1772),.clk(gclk));
	jor g1709(.dina(n1772),.dinb(n1771),.dout(n1773),.clk(gclk));
	jand g1710(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1774),.clk(gclk));
	jnot g1711(.din(n1774),.dout(n1775),.clk(gclk));
	jand g1712(.dina(w_n1751_0[0]),.dinb(w_n1743_0[0]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_n1752_0[0]),.dinb(w_n1740_0[0]),.dout(n1777),.clk(gclk));
	jor g1714(.dina(n1777),.dinb(n1776),.dout(n1778),.clk(gclk));
	jand g1715(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1779),.clk(gclk));
	jand g1716(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1780),.clk(gclk));
	jor g1717(.dina(w_n1748_0[0]),.dinb(w_n1745_0[0]),.dout(n1781),.clk(gclk));
	jor g1718(.dina(w_n1750_0[0]),.dinb(w_n1744_0[0]),.dout(n1782),.clk(gclk));
	jand g1719(.dina(n1782),.dinb(n1781),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1780_0[1]),.dout(n1784),.clk(gclk));
	jnot g1721(.din(n1784),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1779_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1778_0[1]),.dout(n1787),.clk(gclk));
	jxor g1724(.dina(w_n1787_0[1]),.dinb(w_n1775_0[1]),.dout(n1788),.clk(gclk));
	jxor g1725(.dina(w_n1788_0[1]),.dinb(w_n1773_0[1]),.dout(n1789),.clk(gclk));
	jxor g1726(.dina(w_n1789_0[1]),.dinb(w_n1770_0[1]),.dout(n1790),.clk(gclk));
	jxor g1727(.dina(w_n1790_0[1]),.dinb(w_n1768_0[1]),.dout(n1791),.clk(gclk));
	jxor g1728(.dina(w_n1791_0[1]),.dinb(w_n1765_0[1]),.dout(w_dff_A_jerCFLUD1_2),.clk(gclk));
	jnot g1729(.din(w_n1768_0[0]),.dout(n1793),.clk(gclk));
	jnot g1730(.din(w_n1790_0[0]),.dout(n1794),.clk(gclk));
	jor g1731(.dina(n1794),.dinb(n1793),.dout(n1795),.clk(gclk));
	jnot g1732(.din(w_n1791_0[0]),.dout(n1796),.clk(gclk));
	jor g1733(.dina(w_dff_B_BE1ml2kz8_0),.dinb(w_n1765_0[0]),.dout(n1797),.clk(gclk));
	jand g1734(.dina(n1797),.dinb(w_dff_B_IOofLOGl5_1),.dout(n1798),.clk(gclk));
	jand g1735(.dina(w_n1788_0[0]),.dinb(w_n1773_0[0]),.dout(n1799),.clk(gclk));
	jand g1736(.dina(w_n1789_0[0]),.dinb(w_n1770_0[0]),.dout(n1800),.clk(gclk));
	jor g1737(.dina(n1800),.dinb(n1799),.dout(n1801),.clk(gclk));
	jand g1738(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jand g1740(.dina(w_n1786_0[0]),.dinb(w_n1778_0[0]),.dout(n1804),.clk(gclk));
	jand g1741(.dina(w_n1787_0[0]),.dinb(w_n1775_0[0]),.dout(n1805),.clk(gclk));
	jor g1742(.dina(n1805),.dinb(n1804),.dout(n1806),.clk(gclk));
	jand g1743(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1807),.clk(gclk));
	jand g1744(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1808),.clk(gclk));
	jor g1745(.dina(w_n1783_0[0]),.dinb(w_n1780_0[0]),.dout(n1809),.clk(gclk));
	jor g1746(.dina(w_n1785_0[0]),.dinb(w_n1779_0[0]),.dout(n1810),.clk(gclk));
	jand g1747(.dina(n1810),.dinb(n1809),.dout(n1811),.clk(gclk));
	jxor g1748(.dina(w_n1811_0[1]),.dinb(w_n1808_0[1]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(n1812),.dout(n1813),.clk(gclk));
	jxor g1750(.dina(w_n1813_0[1]),.dinb(w_n1807_0[1]),.dout(n1814),.clk(gclk));
	jxor g1751(.dina(w_n1814_0[1]),.dinb(w_n1806_0[1]),.dout(n1815),.clk(gclk));
	jxor g1752(.dina(w_n1815_0[1]),.dinb(w_n1803_0[1]),.dout(n1816),.clk(gclk));
	jxor g1753(.dina(w_n1816_0[1]),.dinb(w_n1801_0[1]),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1817_0[1]),.dinb(w_n1798_0[1]),.dout(w_dff_A_AZmphtiy6_2),.clk(gclk));
	jnot g1755(.din(w_n1801_0[0]),.dout(n1819),.clk(gclk));
	jnot g1756(.din(w_n1816_0[0]),.dout(n1820),.clk(gclk));
	jor g1757(.dina(n1820),.dinb(n1819),.dout(n1821),.clk(gclk));
	jnot g1758(.din(w_n1817_0[0]),.dout(n1822),.clk(gclk));
	jor g1759(.dina(w_dff_B_S11eF9xM5_0),.dinb(w_n1798_0[0]),.dout(n1823),.clk(gclk));
	jand g1760(.dina(n1823),.dinb(w_dff_B_j2KrgK254_1),.dout(n1824),.clk(gclk));
	jand g1761(.dina(w_n1814_0[0]),.dinb(w_n1806_0[0]),.dout(n1825),.clk(gclk));
	jand g1762(.dina(w_n1815_0[0]),.dinb(w_n1803_0[0]),.dout(n1826),.clk(gclk));
	jor g1763(.dina(n1826),.dinb(n1825),.dout(n1827),.clk(gclk));
	jand g1764(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1828),.clk(gclk));
	jand g1765(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1829),.clk(gclk));
	jor g1766(.dina(w_n1811_0[0]),.dinb(w_n1808_0[0]),.dout(n1830),.clk(gclk));
	jor g1767(.dina(w_n1813_0[0]),.dinb(w_n1807_0[0]),.dout(n1831),.clk(gclk));
	jand g1768(.dina(n1831),.dinb(n1830),.dout(n1832),.clk(gclk));
	jxor g1769(.dina(w_n1832_0[1]),.dinb(w_n1829_0[1]),.dout(n1833),.clk(gclk));
	jnot g1770(.din(n1833),.dout(n1834),.clk(gclk));
	jxor g1771(.dina(w_n1834_0[1]),.dinb(w_n1828_0[1]),.dout(n1835),.clk(gclk));
	jxor g1772(.dina(w_n1835_0[1]),.dinb(w_n1827_0[1]),.dout(n1836),.clk(gclk));
	jxor g1773(.dina(w_n1836_0[1]),.dinb(w_n1824_0[1]),.dout(w_dff_A_VrGQGW8r1_2),.clk(gclk));
	jand g1774(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1838),.clk(gclk));
	jor g1775(.dina(w_n1832_0[0]),.dinb(w_n1829_0[0]),.dout(n1839),.clk(gclk));
	jor g1776(.dina(w_n1834_0[0]),.dinb(w_n1828_0[0]),.dout(n1840),.clk(gclk));
	jand g1777(.dina(n1840),.dinb(n1839),.dout(n1841),.clk(gclk));
	jor g1778(.dina(w_n1841_0[1]),.dinb(w_n1838_0[1]),.dout(n1842),.clk(gclk));
	jnot g1779(.din(w_n1827_0[0]),.dout(n1843),.clk(gclk));
	jnot g1780(.din(w_n1835_0[0]),.dout(n1844),.clk(gclk));
	jor g1781(.dina(n1844),.dinb(n1843),.dout(n1845),.clk(gclk));
	jnot g1782(.din(w_n1836_0[0]),.dout(n1846),.clk(gclk));
	jor g1783(.dina(w_dff_B_Mr2wOWV55_0),.dinb(w_n1824_0[0]),.dout(n1847),.clk(gclk));
	jand g1784(.dina(n1847),.dinb(w_dff_B_qcB4i5Lp4_1),.dout(n1848),.clk(gclk));
	jxor g1785(.dina(w_n1841_0[0]),.dinb(w_n1838_0[0]),.dout(n1849),.clk(gclk));
	jnot g1786(.din(w_n1849_0[1]),.dout(n1850),.clk(gclk));
	jor g1787(.dina(w_dff_B_r6oV5yp74_0),.dinb(w_n1848_0[1]),.dout(n1851),.clk(gclk));
	jand g1788(.dina(n1851),.dinb(w_dff_B_dZMtG6911_1),.dout(G6287gat),.clk(gclk));
	jxor g1789(.dina(w_n1849_0[0]),.dinb(w_n1848_0[0]),.dout(w_dff_A_JNspNrBf3_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl3 jspl3_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.doutc(w_G18gat_7[2]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl3 jspl3_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.doutc(w_G273gat_7[2]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_G307gat_2[1]),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl3 jspl3_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.doutc(w_G307gat_7[2]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(w_dff_A_bTCAl6WQ9_1),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n69_0(.douta(w_dff_A_er5FX7J50_0),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_dff_A_DmL1QnrY4_0),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n72_0(.douta(w_n72_0[0]),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.din(n81));
	jspl3 jspl3_w_n82_0(.douta(w_n82_0[0]),.doutb(w_n82_0[1]),.doutc(w_n82_0[2]),.din(n82));
	jspl jspl_w_n82_1(.douta(w_n82_1[0]),.doutb(w_n82_1[1]),.din(w_n82_0[0]));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl jspl_w_n87_0(.douta(w_n87_0[0]),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_n89_0[0]),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl jspl_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n100_0(.douta(w_n100_0[0]),.doutb(w_n100_0[1]),.doutc(w_n100_0[2]),.din(n100));
	jspl jspl_w_n100_1(.douta(w_n100_1[0]),.doutb(w_n100_1[1]),.din(w_n100_0[0]));
	jspl3 jspl3_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.din(n103));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.din(n110));
	jspl jspl_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.din(n115));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.din(n116));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n129_0(.douta(w_n129_0[0]),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.doutc(w_n133_0[2]),.din(n133));
	jspl jspl_w_n138_0(.douta(w_n138_0[0]),.doutb(w_n138_0[1]),.din(n138));
	jspl jspl_w_n139_0(.douta(w_n139_0[0]),.doutb(w_n139_0[1]),.din(n139));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n150_0(.douta(w_n150_0[0]),.doutb(w_n150_0[1]),.din(n150));
	jspl jspl_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.din(n151));
	jspl3 jspl3_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.doutc(w_n156_0[2]),.din(n156));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(n158));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(n165));
	jspl jspl_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.din(n166));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.doutc(w_n169_0[2]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl jspl_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.din(n177));
	jspl jspl_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.din(n178));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl jspl_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.din(n181));
	jspl jspl_w_n183_0(.douta(w_n183_0[0]),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.doutc(w_n194_0[2]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.din(n196));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.din(n209));
	jspl3 jspl3_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.doutc(w_n210_0[2]),.din(n210));
	jspl jspl_w_n210_1(.douta(w_n210_1[0]),.doutb(w_n210_1[1]),.din(w_n210_0[0]));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl jspl_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.din(n215));
	jspl jspl_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.din(n216));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.din(n221));
	jspl jspl_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.din(n223));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.din(n231));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n237_0(.douta(w_n237_0[0]),.doutb(w_n237_0[1]),.doutc(w_n237_0[2]),.din(n237));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(n239));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.din(n244));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_n257_0[1]),.din(n257));
	jspl3 jspl3_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.doutc(w_n258_0[2]),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(n265));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(n267));
	jspl jspl_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.din(n268));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.din(n269));
	jspl jspl_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.din(n270));
	jspl jspl_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.din(n283));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(n290));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(n295));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_n300_0[1]),.din(n300));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(n305));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(n310));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.doutc(w_n314_0[2]),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.din(n317));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.din(n321));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(n323));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.din(n326));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(n327));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(n330));
	jspl jspl_w_n332_0(.douta(w_n332_0[0]),.doutb(w_n332_0[1]),.din(n332));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.din(n335));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl jspl_w_n341_0(.douta(w_n341_0[0]),.doutb(w_n341_0[1]),.din(n341));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n351_0(.douta(w_n351_0[0]),.doutb(w_n351_0[1]),.din(n351));
	jspl jspl_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.din(n353));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(n356));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(n358));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(n363));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(n366));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(n368));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl3 jspl3_w_n376_0(.douta(w_n376_0[0]),.doutb(w_n376_0[1]),.doutc(w_n376_0[2]),.din(n376));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.din(n377));
	jspl jspl_w_n380_0(.douta(w_n380_0[0]),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.din(n382));
	jspl jspl_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.din(n383));
	jspl jspl_w_n384_0(.douta(w_n384_0[0]),.doutb(w_n384_0[1]),.din(n384));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl jspl_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.din(n387));
	jspl jspl_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.din(n388));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.din(n389));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(n390));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(n391));
	jspl jspl_w_n392_0(.douta(w_n392_0[0]),.doutb(w_n392_0[1]),.din(n392));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.din(n396));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n399_0(.douta(w_n399_0[0]),.doutb(w_n399_0[1]),.din(n399));
	jspl jspl_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_n410_0[2]),.din(n410));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(n412));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl jspl_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.din(n417));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.din(n420));
	jspl jspl_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.din(n422));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(n427));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(n432));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_n442_0[1]),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.doutc(w_n446_0[2]),.din(n446));
	jspl jspl_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.din(n447));
	jspl jspl_w_n450_0(.douta(w_n450_0[0]),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.din(n453));
	jspl jspl_w_n454_0(.douta(w_n454_0[0]),.doutb(w_n454_0[1]),.din(n454));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.din(n455));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl jspl_w_n458_0(.douta(w_n458_0[0]),.doutb(w_n458_0[1]),.din(n458));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(n459));
	jspl jspl_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.din(n460));
	jspl jspl_w_n461_0(.douta(w_n461_0[0]),.doutb(w_n461_0[1]),.din(n461));
	jspl jspl_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.din(n462));
	jspl jspl_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.din(n463));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(n464));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(n466));
	jspl jspl_w_n468_0(.douta(w_n468_0[0]),.doutb(w_n468_0[1]),.din(n468));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(n469));
	jspl jspl_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.din(n471));
	jspl jspl_w_n476_0(.douta(w_n476_0[0]),.doutb(w_n476_0[1]),.din(n476));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl3 jspl3_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.doutc(w_n482_0[2]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(n489));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl jspl_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.din(n497));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(n499));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(n509));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(n519));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.doutc(w_n523_0[2]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_n529_0[0]),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(n530));
	jspl jspl_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.din(n531));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(n532));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.din(n535));
	jspl jspl_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.din(n536));
	jspl jspl_w_n537_0(.douta(w_n537_0[0]),.doutb(w_n537_0[1]),.din(n537));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(n547));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.din(n556));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(n563));
	jspl jspl_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.din(n566));
	jspl jspl_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.din(n568));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.din(n571));
	jspl jspl_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.din(n573));
	jspl jspl_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.din(n576));
	jspl jspl_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.din(n578));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl jspl_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.din(n583));
	jspl jspl_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(n588));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(n596));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(n606));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n611_0(.douta(w_n611_0[0]),.doutb(w_n611_0[1]),.din(n611));
	jspl jspl_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.din(n613));
	jspl jspl_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.din(n614));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl jspl_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.din(n617));
	jspl jspl_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.din(n618));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.din(n620));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.din(n621));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.din(n625));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(n626));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(n628));
	jspl jspl_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.din(n629));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.din(n633));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl jspl_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.din(n636));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.doutc(w_n647_0[2]),.din(n647));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(n654));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(n662));
	jspl jspl_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.din(n664));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(n667));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(n669));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(n674));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.din(n679));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.doutc(w_n695_0[2]),.din(n695));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl3 jspl3_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.doutc(w_n698_0[2]),.din(n698));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n702_0(.douta(w_n702_0[0]),.doutb(w_n702_0[1]),.din(n702));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.din(n707));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.din(n708));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(n709));
	jspl jspl_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl jspl_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.din(n714));
	jspl jspl_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.din(n715));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl jspl_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.din(n718));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(n719));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(n721));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(n724));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.din(n729));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(n734));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.din(n735));
	jspl3 jspl3_w_n740_0(.douta(w_n740_0[0]),.doutb(w_n740_0[1]),.doutc(w_n740_0[2]),.din(n740));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(n747));
	jspl jspl_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl jspl_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.din(n755));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(n762));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl jspl_w_n770_0(.douta(w_n770_0[0]),.doutb(w_n770_0[1]),.din(n770));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(n772));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(n787));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl jspl_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.din(n793));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl jspl_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(n803));
	jspl jspl_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.din(n804));
	jspl jspl_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.din(n806));
	jspl jspl_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.din(n807));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.din(n808));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(n811));
	jspl jspl_w_n812_0(.douta(w_n812_0[0]),.doutb(w_n812_0[1]),.din(n812));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl jspl_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.din(n814));
	jspl jspl_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(n817));
	jspl jspl_w_n818_0(.douta(w_n818_0[0]),.doutb(w_n818_0[1]),.din(n818));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(n819));
	jspl jspl_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.din(n820));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(n821));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(n822));
	jspl jspl_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n826_0(.douta(w_n826_0[0]),.doutb(w_n826_0[1]),.din(n826));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n829_0(.douta(w_n829_0[0]),.doutb(w_n829_0[1]),.din(n829));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl jspl_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.din(n840));
	jspl3 jspl3_w_n844_0(.douta(w_n844_0[0]),.doutb(w_n844_0[1]),.doutc(w_n844_0[2]),.din(n844));
	jspl jspl_w_n846_0(.douta(w_n846_0[0]),.doutb(w_n846_0[1]),.din(n846));
	jspl jspl_w_n849_0(.douta(w_n849_0[0]),.doutb(w_n849_0[1]),.din(n849));
	jspl jspl_w_n851_0(.douta(w_n851_0[0]),.doutb(w_n851_0[1]),.din(n851));
	jspl jspl_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.din(n854));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(n861));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(n866));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(n874));
	jspl jspl_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.din(n876));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(n886));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(n891));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(n896));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(n898));
	jspl jspl_w_n901_0(.douta(w_n901_0[0]),.doutb(w_n901_0[1]),.din(n901));
	jspl jspl_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n906_0(.douta(w_n906_0[0]),.doutb(w_n906_0[1]),.din(n906));
	jspl jspl_w_n907_0(.douta(w_n907_0[0]),.doutb(w_n907_0[1]),.din(n907));
	jspl jspl_w_n908_0(.douta(w_n908_0[0]),.doutb(w_n908_0[1]),.din(n908));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(n910));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(n911));
	jspl jspl_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.din(n912));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(n913));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.din(n915));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(n916));
	jspl jspl_w_n917_0(.douta(w_n917_0[0]),.doutb(w_n917_0[1]),.din(n917));
	jspl jspl_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.din(n918));
	jspl jspl_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.din(n919));
	jspl jspl_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.din(n920));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(n923));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(n924));
	jspl jspl_w_n925_0(.douta(w_n925_0[0]),.doutb(w_n925_0[1]),.din(n925));
	jspl jspl_w_n926_0(.douta(w_n926_0[0]),.doutb(w_n926_0[1]),.din(n926));
	jspl3 jspl3_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.doutc(w_n927_0[2]),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(n929));
	jspl jspl_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.din(n930));
	jspl jspl_w_n931_0(.douta(w_n931_0[0]),.doutb(w_n931_0[1]),.din(n931));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(n938));
	jspl3 jspl3_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.doutc(w_n942_0[2]),.din(n942));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_n943_0[1]),.din(n943));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(n949));
	jspl jspl_w_n951_0(.douta(w_n951_0[0]),.doutb(w_n951_0[1]),.din(n951));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n956_0(.douta(w_n956_0[0]),.doutb(w_n956_0[1]),.din(n956));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(n959));
	jspl jspl_w_n961_0(.douta(w_n961_0[0]),.doutb(w_n961_0[1]),.din(n961));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.din(n966));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_n971_0[1]),.din(n971));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n976_0(.douta(w_n976_0[0]),.doutb(w_n976_0[1]),.din(n976));
	jspl jspl_w_n979_0(.douta(w_n979_0[0]),.doutb(w_n979_0[1]),.din(n979));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(n991));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(n996));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.din(n1006));
	jspl jspl_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1010_0(.douta(w_n1010_0[0]),.doutb(w_n1010_0[1]),.din(n1010));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.din(n1012));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl jspl_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.din(n1014));
	jspl jspl_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.din(n1015));
	jspl jspl_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.din(n1016));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(n1018));
	jspl jspl_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.din(n1019));
	jspl jspl_w_n1020_0(.douta(w_n1020_0[0]),.doutb(w_n1020_0[1]),.din(n1020));
	jspl jspl_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.din(n1021));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(n1023));
	jspl jspl_w_n1024_0(.douta(w_n1024_0[0]),.doutb(w_n1024_0[1]),.din(n1024));
	jspl jspl_w_n1025_0(.douta(w_n1025_0[0]),.doutb(w_n1025_0[1]),.din(n1025));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1027_0(.douta(w_n1027_0[0]),.doutb(w_n1027_0[1]),.din(n1027));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(n1028));
	jspl jspl_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.din(n1029));
	jspl jspl_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.din(n1030));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.din(n1032));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1034_0(.douta(w_n1034_0[0]),.doutb(w_n1034_0[1]),.din(n1034));
	jspl jspl_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.din(n1035));
	jspl jspl_w_n1037_0(.douta(w_n1037_0[0]),.doutb(w_n1037_0[1]),.din(w_dff_B_wDX4iwEr7_2));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_dff_A_7UVDgp5P2_1),.din(n1039));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(n1043));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(n1044));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(n1048));
	jspl jspl_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.din(n1049));
	jspl jspl_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.din(n1054));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.din(n1057));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(n1059));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.din(n1062));
	jspl jspl_w_n1064_0(.douta(w_n1064_0[0]),.doutb(w_n1064_0[1]),.din(n1064));
	jspl jspl_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.din(n1067));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(n1069));
	jspl jspl_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.din(n1072));
	jspl jspl_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.din(n1074));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(n1077));
	jspl jspl_w_n1079_0(.douta(w_n1079_0[0]),.doutb(w_n1079_0[1]),.din(n1079));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(n1084));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(n1087));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(n1089));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(n1094));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(n1103));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1110_0(.douta(w_n1110_0[0]),.doutb(w_n1110_0[1]),.din(n1110));
	jspl jspl_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.din(n1114));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.din(n1116));
	jspl jspl_w_n1117_0(.douta(w_n1117_0[0]),.doutb(w_n1117_0[1]),.din(n1117));
	jspl jspl_w_n1118_0(.douta(w_n1118_0[0]),.doutb(w_n1118_0[1]),.din(n1118));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(n1119));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl jspl_w_n1121_0(.douta(w_n1121_0[0]),.doutb(w_n1121_0[1]),.din(n1121));
	jspl jspl_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.din(n1122));
	jspl jspl_w_n1123_0(.douta(w_n1123_0[0]),.doutb(w_n1123_0[1]),.din(n1123));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.din(n1125));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(n1126));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(n1127));
	jspl jspl_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.din(n1128));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(n1131));
	jspl jspl_w_n1132_0(.douta(w_n1132_0[0]),.doutb(w_n1132_0[1]),.din(n1132));
	jspl jspl_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.din(n1133));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1135_0(.douta(w_n1135_0[0]),.doutb(w_n1135_0[1]),.din(n1135));
	jspl jspl_w_n1137_0(.douta(w_n1137_0[0]),.doutb(w_n1137_0[1]),.din(n1137));
	jspl jspl_w_n1138_0(.douta(w_n1138_0[0]),.doutb(w_n1138_0[1]),.din(n1138));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1140_0(.douta(w_n1140_0[0]),.doutb(w_n1140_0[1]),.din(n1140));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(n1141));
	jspl jspl_w_n1147_0(.douta(w_n1147_0[0]),.doutb(w_n1147_0[1]),.din(n1147));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(n1151));
	jspl jspl_w_n1152_0(.douta(w_n1152_0[0]),.doutb(w_n1152_0[1]),.din(n1152));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(n1156));
	jspl jspl_w_n1158_0(.douta(w_n1158_0[0]),.doutb(w_n1158_0[1]),.din(n1158));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(n1161));
	jspl jspl_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.din(n1163));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl jspl_w_n1168_0(.douta(w_n1168_0[0]),.doutb(w_n1168_0[1]),.din(n1168));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(n1171));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(n1173));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(n1176));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.din(n1178));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(n1183));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(n1186));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(n1188));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(n1191));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(n1193));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(n1198));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(n1203));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(n1206));
	jspl jspl_w_n1207_0(.douta(w_n1207_0[0]),.doutb(w_n1207_0[1]),.din(n1207));
	jspl jspl_w_n1208_0(.douta(w_n1208_0[0]),.doutb(w_n1208_0[1]),.din(n1208));
	jspl jspl_w_n1210_0(.douta(w_n1210_0[0]),.doutb(w_n1210_0[1]),.din(n1210));
	jspl jspl_w_n1212_0(.douta(w_n1212_0[0]),.doutb(w_n1212_0[1]),.din(n1212));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1214_0(.douta(w_n1214_0[0]),.doutb(w_n1214_0[1]),.din(n1214));
	jspl jspl_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.din(n1215));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(n1217));
	jspl jspl_w_n1218_0(.douta(w_n1218_0[0]),.doutb(w_n1218_0[1]),.din(n1218));
	jspl jspl_w_n1219_0(.douta(w_n1219_0[0]),.doutb(w_n1219_0[1]),.din(n1219));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1221_0(.douta(w_n1221_0[0]),.doutb(w_n1221_0[1]),.din(n1221));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(n1222));
	jspl jspl_w_n1223_0(.douta(w_n1223_0[0]),.doutb(w_n1223_0[1]),.din(n1223));
	jspl jspl_w_n1224_0(.douta(w_n1224_0[0]),.doutb(w_n1224_0[1]),.din(n1224));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(n1225));
	jspl jspl_w_n1226_0(.douta(w_n1226_0[0]),.doutb(w_n1226_0[1]),.din(n1226));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(n1227));
	jspl jspl_w_n1228_0(.douta(w_n1228_0[0]),.doutb(w_n1228_0[1]),.din(n1228));
	jspl jspl_w_n1229_0(.douta(w_n1229_0[0]),.doutb(w_n1229_0[1]),.din(n1229));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1231_0(.douta(w_n1231_0[0]),.doutb(w_n1231_0[1]),.din(n1231));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(n1232));
	jspl jspl_w_n1234_0(.douta(w_n1234_0[0]),.doutb(w_n1234_0[1]),.din(n1234));
	jspl jspl_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(n1237));
	jspl jspl_w_n1238_0(.douta(w_n1238_0[0]),.doutb(w_n1238_0[1]),.din(n1238));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(n1247));
	jspl jspl_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.din(n1248));
	jspl jspl_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.din(n1251));
	jspl jspl_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.din(n1253));
	jspl jspl_w_n1256_0(.douta(w_n1256_0[0]),.doutb(w_n1256_0[1]),.din(n1256));
	jspl jspl_w_n1258_0(.douta(w_n1258_0[0]),.doutb(w_n1258_0[1]),.din(n1258));
	jspl jspl_w_n1261_0(.douta(w_n1261_0[0]),.doutb(w_n1261_0[1]),.din(n1261));
	jspl jspl_w_n1263_0(.douta(w_n1263_0[0]),.doutb(w_n1263_0[1]),.din(n1263));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(n1266));
	jspl jspl_w_n1268_0(.douta(w_n1268_0[0]),.doutb(w_n1268_0[1]),.din(n1268));
	jspl jspl_w_n1271_0(.douta(w_n1271_0[0]),.doutb(w_n1271_0[1]),.din(n1271));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(n1273));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(n1276));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(n1278));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(n1281));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(n1283));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(n1286));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(n1288));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_n1291_0[1]),.din(n1291));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(n1293));
	jspl jspl_w_n1296_0(.douta(w_n1296_0[0]),.doutb(w_n1296_0[1]),.din(n1296));
	jspl jspl_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.din(n1297));
	jspl jspl_w_n1298_0(.douta(w_n1298_0[0]),.doutb(w_n1298_0[1]),.din(n1298));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1303_0(.douta(w_n1303_0[0]),.doutb(w_n1303_0[1]),.din(n1303));
	jspl jspl_w_n1304_0(.douta(w_n1304_0[0]),.doutb(w_n1304_0[1]),.din(n1304));
	jspl jspl_w_n1305_0(.douta(w_n1305_0[0]),.doutb(w_n1305_0[1]),.din(n1305));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(n1307));
	jspl jspl_w_n1308_0(.douta(w_n1308_0[0]),.doutb(w_n1308_0[1]),.din(n1308));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl jspl_w_n1311_0(.douta(w_n1311_0[0]),.doutb(w_n1311_0[1]),.din(n1311));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(n1312));
	jspl jspl_w_n1313_0(.douta(w_n1313_0[0]),.doutb(w_n1313_0[1]),.din(n1313));
	jspl jspl_w_n1314_0(.douta(w_n1314_0[0]),.doutb(w_n1314_0[1]),.din(n1314));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.din(n1316));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1318_0(.douta(w_n1318_0[0]),.doutb(w_n1318_0[1]),.din(n1318));
	jspl jspl_w_n1319_0(.douta(w_n1319_0[0]),.doutb(w_n1319_0[1]),.din(n1319));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.din(n1321));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.din(n1322));
	jspl jspl_w_n1324_0(.douta(w_n1324_0[0]),.doutb(w_n1324_0[1]),.din(n1324));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl jspl_w_n1326_0(.douta(w_n1326_0[0]),.doutb(w_n1326_0[1]),.din(n1326));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(n1332));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(n1337));
	jspl jspl_w_n1338_0(.douta(w_n1338_0[0]),.doutb(w_n1338_0[1]),.din(n1338));
	jspl jspl_w_n1341_0(.douta(w_n1341_0[0]),.doutb(w_n1341_0[1]),.din(n1341));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(n1343));
	jspl jspl_w_n1346_0(.douta(w_n1346_0[0]),.doutb(w_n1346_0[1]),.din(n1346));
	jspl jspl_w_n1348_0(.douta(w_n1348_0[0]),.doutb(w_n1348_0[1]),.din(n1348));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(n1351));
	jspl jspl_w_n1353_0(.douta(w_n1353_0[0]),.doutb(w_n1353_0[1]),.din(n1353));
	jspl jspl_w_n1356_0(.douta(w_n1356_0[0]),.doutb(w_n1356_0[1]),.din(n1356));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(n1363));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(n1366));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(n1368));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(n1373));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(n1376));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(n1378));
	jspl jspl_w_n1381_0(.douta(w_n1381_0[0]),.doutb(w_n1381_0[1]),.din(n1381));
	jspl jspl_w_n1382_0(.douta(w_n1382_0[0]),.doutb(w_n1382_0[1]),.din(n1382));
	jspl jspl_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.din(n1383));
	jspl jspl_w_n1386_0(.douta(w_n1386_0[0]),.doutb(w_n1386_0[1]),.din(n1386));
	jspl jspl_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_n1388_0[1]),.din(n1388));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(n1389));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(n1390));
	jspl jspl_w_n1391_0(.douta(w_n1391_0[0]),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1392_0(.douta(w_n1392_0[0]),.doutb(w_n1392_0[1]),.din(n1392));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(n1395));
	jspl jspl_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.din(n1396));
	jspl jspl_w_n1397_0(.douta(w_n1397_0[0]),.doutb(w_n1397_0[1]),.din(n1397));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(n1399));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(n1400));
	jspl jspl_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_n1401_0[1]),.din(n1401));
	jspl jspl_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_n1402_0[1]),.din(n1402));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_n1404_0[1]),.din(n1404));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl jspl_w_n1407_0(.douta(w_n1407_0[0]),.doutb(w_n1407_0[1]),.din(n1407));
	jspl jspl_w_n1409_0(.douta(w_n1409_0[0]),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(n1410));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(n1415));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(n1420));
	jspl jspl_w_n1421_0(.douta(w_n1421_0[0]),.doutb(w_n1421_0[1]),.din(n1421));
	jspl jspl_w_n1424_0(.douta(w_n1424_0[0]),.doutb(w_n1424_0[1]),.din(n1424));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(n1426));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(n1431));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(n1436));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(n1444));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(n1449));
	jspl jspl_w_n1451_0(.douta(w_n1451_0[0]),.doutb(w_n1451_0[1]),.din(n1451));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(n1454));
	jspl jspl_w_n1456_0(.douta(w_n1456_0[0]),.doutb(w_n1456_0[1]),.din(n1456));
	jspl jspl_w_n1459_0(.douta(w_n1459_0[0]),.doutb(w_n1459_0[1]),.din(n1459));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(n1460));
	jspl jspl_w_n1461_0(.douta(w_n1461_0[0]),.doutb(w_n1461_0[1]),.din(n1461));
	jspl jspl_w_n1464_0(.douta(w_n1464_0[0]),.doutb(w_n1464_0[1]),.din(n1464));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(n1466));
	jspl jspl_w_n1467_0(.douta(w_n1467_0[0]),.doutb(w_n1467_0[1]),.din(n1467));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_n1468_0[1]),.din(n1468));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1470_0(.douta(w_n1470_0[0]),.doutb(w_n1470_0[1]),.din(n1470));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(n1471));
	jspl jspl_w_n1472_0(.douta(w_n1472_0[0]),.doutb(w_n1472_0[1]),.din(n1472));
	jspl jspl_w_n1473_0(.douta(w_n1473_0[0]),.doutb(w_n1473_0[1]),.din(n1473));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(n1474));
	jspl jspl_w_n1475_0(.douta(w_n1475_0[0]),.doutb(w_n1475_0[1]),.din(n1475));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(n1476));
	jspl jspl_w_n1477_0(.douta(w_n1477_0[0]),.doutb(w_n1477_0[1]),.din(n1477));
	jspl jspl_w_n1478_0(.douta(w_n1478_0[0]),.doutb(w_n1478_0[1]),.din(n1478));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(n1479));
	jspl jspl_w_n1480_0(.douta(w_n1480_0[0]),.doutb(w_n1480_0[1]),.din(n1480));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(n1481));
	jspl jspl_w_n1483_0(.douta(w_n1483_0[0]),.doutb(w_n1483_0[1]),.din(n1483));
	jspl jspl_w_n1485_0(.douta(w_n1485_0[0]),.doutb(w_n1485_0[1]),.din(n1485));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(n1486));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(n1491));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(n1496));
	jspl jspl_w_n1497_0(.douta(w_n1497_0[0]),.doutb(w_n1497_0[1]),.din(n1497));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(n1500));
	jspl jspl_w_n1502_0(.douta(w_n1502_0[0]),.doutb(w_n1502_0[1]),.din(n1502));
	jspl jspl_w_n1505_0(.douta(w_n1505_0[0]),.doutb(w_n1505_0[1]),.din(n1505));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(n1507));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(n1512));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(n1515));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(n1517));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.din(n1520));
	jspl jspl_w_n1522_0(.douta(w_n1522_0[0]),.doutb(w_n1522_0[1]),.din(n1522));
	jspl jspl_w_n1525_0(.douta(w_n1525_0[0]),.doutb(w_n1525_0[1]),.din(n1525));
	jspl jspl_w_n1527_0(.douta(w_n1527_0[0]),.doutb(w_n1527_0[1]),.din(n1527));
	jspl jspl_w_n1530_0(.douta(w_n1530_0[0]),.doutb(w_n1530_0[1]),.din(n1530));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(n1531));
	jspl jspl_w_n1532_0(.douta(w_n1532_0[0]),.doutb(w_n1532_0[1]),.din(n1532));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(n1535));
	jspl jspl_w_n1537_0(.douta(w_n1537_0[0]),.doutb(w_n1537_0[1]),.din(n1537));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.din(n1539));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(n1540));
	jspl jspl_w_n1541_0(.douta(w_n1541_0[0]),.doutb(w_n1541_0[1]),.din(n1541));
	jspl jspl_w_n1542_0(.douta(w_n1542_0[0]),.doutb(w_n1542_0[1]),.din(n1542));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1544_0(.douta(w_n1544_0[0]),.doutb(w_n1544_0[1]),.din(n1544));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1546_0(.douta(w_n1546_0[0]),.doutb(w_n1546_0[1]),.din(n1546));
	jspl jspl_w_n1547_0(.douta(w_n1547_0[0]),.doutb(w_n1547_0[1]),.din(n1547));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(n1548));
	jspl jspl_w_n1549_0(.douta(w_n1549_0[0]),.doutb(w_n1549_0[1]),.din(n1549));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_n1550_0[1]),.din(n1550));
	jspl jspl_w_n1552_0(.douta(w_n1552_0[0]),.doutb(w_n1552_0[1]),.din(n1552));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(n1565));
	jspl jspl_w_n1566_0(.douta(w_n1566_0[0]),.doutb(w_n1566_0[1]),.din(n1566));
	jspl jspl_w_n1569_0(.douta(w_n1569_0[0]),.doutb(w_n1569_0[1]),.din(n1569));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(n1571));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(n1574));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(n1576));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(n1579));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_n1581_0[1]),.din(n1581));
	jspl jspl_w_n1584_0(.douta(w_n1584_0[0]),.doutb(w_n1584_0[1]),.din(n1584));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.din(n1586));
	jspl jspl_w_n1589_0(.douta(w_n1589_0[0]),.doutb(w_n1589_0[1]),.din(n1589));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1594_0(.douta(w_n1594_0[0]),.doutb(w_n1594_0[1]),.din(n1594));
	jspl jspl_w_n1595_0(.douta(w_n1595_0[0]),.doutb(w_n1595_0[1]),.din(n1595));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_n1603_0[1]),.din(n1603));
	jspl jspl_w_n1604_0(.douta(w_n1604_0[0]),.doutb(w_n1604_0[1]),.din(n1604));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1606_0(.douta(w_n1606_0[0]),.doutb(w_n1606_0[1]),.din(n1606));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1608_0(.douta(w_n1608_0[0]),.doutb(w_n1608_0[1]),.din(n1608));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.din(n1611));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(n1612));
	jspl jspl_w_n1614_0(.douta(w_n1614_0[0]),.doutb(w_n1614_0[1]),.din(n1614));
	jspl jspl_w_n1616_0(.douta(w_n1616_0[0]),.doutb(w_n1616_0[1]),.din(n1616));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_n1617_0[1]),.din(n1617));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(n1622));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(n1628));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(n1631));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(n1633));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(n1636));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(n1638));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_n1641_0[1]),.din(n1641));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(n1643));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(n1646));
	jspl jspl_w_n1648_0(.douta(w_n1648_0[0]),.doutb(w_n1648_0[1]),.din(n1648));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(n1651));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_n1652_0[1]),.din(n1652));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(n1653));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(n1656));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(n1658));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1660_0(.douta(w_n1660_0[0]),.doutb(w_n1660_0[1]),.din(n1660));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(n1661));
	jspl jspl_w_n1662_0(.douta(w_n1662_0[0]),.doutb(w_n1662_0[1]),.din(n1662));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(n1663));
	jspl jspl_w_n1664_0(.douta(w_n1664_0[0]),.doutb(w_n1664_0[1]),.din(n1664));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(n1666));
	jspl jspl_w_n1667_0(.douta(w_n1667_0[0]),.doutb(w_n1667_0[1]),.din(n1667));
	jspl jspl_w_n1669_0(.douta(w_n1669_0[0]),.doutb(w_n1669_0[1]),.din(n1669));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(n1671));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(n1672));
	jspl jspl_w_n1677_0(.douta(w_n1677_0[0]),.doutb(w_n1677_0[1]),.din(n1677));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(n1682));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(n1684));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_n1687_0[1]),.din(n1687));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(n1689));
	jspl jspl_w_n1692_0(.douta(w_n1692_0[0]),.doutb(w_n1692_0[1]),.din(n1692));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(n1694));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_n1697_0[1]),.din(n1697));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(n1699));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(n1702));
	jspl jspl_w_n1703_0(.douta(w_n1703_0[0]),.doutb(w_n1703_0[1]),.din(n1703));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(n1704));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(n1707));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(n1709));
	jspl jspl_w_n1710_0(.douta(w_n1710_0[0]),.doutb(w_n1710_0[1]),.din(n1710));
	jspl jspl_w_n1711_0(.douta(w_n1711_0[0]),.doutb(w_n1711_0[1]),.din(n1711));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(n1712));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(n1713));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(n1714));
	jspl jspl_w_n1715_0(.douta(w_n1715_0[0]),.doutb(w_n1715_0[1]),.din(n1715));
	jspl jspl_w_n1716_0(.douta(w_n1716_0[0]),.doutb(w_n1716_0[1]),.din(n1716));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_n1720_0[1]),.din(n1720));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1728_0(.douta(w_n1728_0[0]),.doutb(w_n1728_0[1]),.din(n1728));
	jspl jspl_w_n1730_0(.douta(w_n1730_0[0]),.doutb(w_n1730_0[1]),.din(n1730));
	jspl jspl_w_n1733_0(.douta(w_n1733_0[0]),.doutb(w_n1733_0[1]),.din(n1733));
	jspl jspl_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.din(n1735));
	jspl jspl_w_n1738_0(.douta(w_n1738_0[0]),.doutb(w_n1738_0[1]),.din(n1738));
	jspl jspl_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.din(n1740));
	jspl jspl_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.din(n1743));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(n1744));
	jspl jspl_w_n1745_0(.douta(w_n1745_0[0]),.doutb(w_n1745_0[1]),.din(n1745));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(n1748));
	jspl jspl_w_n1750_0(.douta(w_n1750_0[0]),.doutb(w_n1750_0[1]),.din(n1750));
	jspl jspl_w_n1751_0(.douta(w_n1751_0[0]),.doutb(w_n1751_0[1]),.din(n1751));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1753_0(.douta(w_n1753_0[0]),.doutb(w_n1753_0[1]),.din(n1753));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_n1758_0[1]),.din(n1758));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl jspl_w_n1768_0(.douta(w_n1768_0[0]),.doutb(w_n1768_0[1]),.din(n1768));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(n1770));
	jspl jspl_w_n1773_0(.douta(w_n1773_0[0]),.doutb(w_n1773_0[1]),.din(n1773));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(n1775));
	jspl jspl_w_n1778_0(.douta(w_n1778_0[0]),.doutb(w_n1778_0[1]),.din(n1778));
	jspl jspl_w_n1779_0(.douta(w_n1779_0[0]),.doutb(w_n1779_0[1]),.din(n1779));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(n1780));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_n1786_0[1]),.din(n1786));
	jspl jspl_w_n1787_0(.douta(w_n1787_0[0]),.doutb(w_n1787_0[1]),.din(n1787));
	jspl jspl_w_n1788_0(.douta(w_n1788_0[0]),.doutb(w_n1788_0[1]),.din(n1788));
	jspl jspl_w_n1789_0(.douta(w_n1789_0[0]),.doutb(w_n1789_0[1]),.din(n1789));
	jspl jspl_w_n1790_0(.douta(w_n1790_0[0]),.doutb(w_n1790_0[1]),.din(n1790));
	jspl jspl_w_n1791_0(.douta(w_n1791_0[0]),.doutb(w_n1791_0[1]),.din(n1791));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(n1798));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_n1801_0[1]),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(n1803));
	jspl jspl_w_n1806_0(.douta(w_n1806_0[0]),.doutb(w_n1806_0[1]),.din(n1806));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(n1807));
	jspl jspl_w_n1808_0(.douta(w_n1808_0[0]),.doutb(w_n1808_0[1]),.din(n1808));
	jspl jspl_w_n1811_0(.douta(w_n1811_0[0]),.doutb(w_n1811_0[1]),.din(n1811));
	jspl jspl_w_n1813_0(.douta(w_n1813_0[0]),.doutb(w_n1813_0[1]),.din(n1813));
	jspl jspl_w_n1814_0(.douta(w_n1814_0[0]),.doutb(w_n1814_0[1]),.din(n1814));
	jspl jspl_w_n1815_0(.douta(w_n1815_0[0]),.doutb(w_n1815_0[1]),.din(n1815));
	jspl jspl_w_n1816_0(.douta(w_n1816_0[0]),.doutb(w_n1816_0[1]),.din(n1816));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_n1817_0[1]),.din(n1817));
	jspl jspl_w_n1824_0(.douta(w_n1824_0[0]),.doutb(w_n1824_0[1]),.din(n1824));
	jspl jspl_w_n1827_0(.douta(w_n1827_0[0]),.doutb(w_n1827_0[1]),.din(n1827));
	jspl jspl_w_n1828_0(.douta(w_n1828_0[0]),.doutb(w_n1828_0[1]),.din(n1828));
	jspl jspl_w_n1829_0(.douta(w_n1829_0[0]),.doutb(w_n1829_0[1]),.din(n1829));
	jspl jspl_w_n1832_0(.douta(w_n1832_0[0]),.doutb(w_n1832_0[1]),.din(n1832));
	jspl jspl_w_n1834_0(.douta(w_n1834_0[0]),.doutb(w_n1834_0[1]),.din(n1834));
	jspl jspl_w_n1835_0(.douta(w_n1835_0[0]),.doutb(w_n1835_0[1]),.din(n1835));
	jspl jspl_w_n1836_0(.douta(w_n1836_0[0]),.doutb(w_n1836_0[1]),.din(n1836));
	jspl jspl_w_n1838_0(.douta(w_n1838_0[0]),.doutb(w_n1838_0[1]),.din(n1838));
	jspl jspl_w_n1841_0(.douta(w_n1841_0[0]),.doutb(w_n1841_0[1]),.din(n1841));
	jspl jspl_w_n1848_0(.douta(w_n1848_0[0]),.doutb(w_n1848_0[1]),.din(n1848));
	jspl jspl_w_n1849_0(.douta(w_n1849_0[0]),.doutb(w_n1849_0[1]),.din(n1849));
	jdff dff_B_bbppiPhb7_1(.din(n67),.dout(w_dff_B_bbppiPhb7_1),.clk(gclk));
	jdff dff_B_AvIxvPmF5_1(.din(n73),.dout(w_dff_B_AvIxvPmF5_1),.clk(gclk));
	jdff dff_B_jTjV4pz17_1(.din(w_dff_B_AvIxvPmF5_1),.dout(w_dff_B_jTjV4pz17_1),.clk(gclk));
	jdff dff_B_0LjNHhat3_1(.din(w_dff_B_jTjV4pz17_1),.dout(w_dff_B_0LjNHhat3_1),.clk(gclk));
	jdff dff_B_FZ3q2YcR3_1(.din(w_dff_B_0LjNHhat3_1),.dout(w_dff_B_FZ3q2YcR3_1),.clk(gclk));
	jdff dff_B_qcojHCOn8_1(.din(n90),.dout(w_dff_B_qcojHCOn8_1),.clk(gclk));
	jdff dff_B_bDc5GmoL9_1(.din(w_dff_B_qcojHCOn8_1),.dout(w_dff_B_bDc5GmoL9_1),.clk(gclk));
	jdff dff_B_5ukqYSMc0_1(.din(w_dff_B_bDc5GmoL9_1),.dout(w_dff_B_5ukqYSMc0_1),.clk(gclk));
	jdff dff_B_migKC2OD1_1(.din(w_dff_B_5ukqYSMc0_1),.dout(w_dff_B_migKC2OD1_1),.clk(gclk));
	jdff dff_B_U7JZyBM13_1(.din(w_dff_B_migKC2OD1_1),.dout(w_dff_B_U7JZyBM13_1),.clk(gclk));
	jdff dff_B_Y2Q3omrR4_1(.din(w_dff_B_U7JZyBM13_1),.dout(w_dff_B_Y2Q3omrR4_1),.clk(gclk));
	jdff dff_B_PgYh4dwy6_1(.din(w_dff_B_Y2Q3omrR4_1),.dout(w_dff_B_PgYh4dwy6_1),.clk(gclk));
	jdff dff_B_v0ge0q491_1(.din(n111),.dout(w_dff_B_v0ge0q491_1),.clk(gclk));
	jdff dff_B_hAehoMhR4_1(.din(w_dff_B_v0ge0q491_1),.dout(w_dff_B_hAehoMhR4_1),.clk(gclk));
	jdff dff_B_p9QM19To9_1(.din(w_dff_B_hAehoMhR4_1),.dout(w_dff_B_p9QM19To9_1),.clk(gclk));
	jdff dff_B_UJv3YTAA8_1(.din(w_dff_B_p9QM19To9_1),.dout(w_dff_B_UJv3YTAA8_1),.clk(gclk));
	jdff dff_B_rggcB22Q3_1(.din(w_dff_B_UJv3YTAA8_1),.dout(w_dff_B_rggcB22Q3_1),.clk(gclk));
	jdff dff_B_6N3bllvZ7_1(.din(w_dff_B_rggcB22Q3_1),.dout(w_dff_B_6N3bllvZ7_1),.clk(gclk));
	jdff dff_B_5rTwhrzE4_1(.din(w_dff_B_6N3bllvZ7_1),.dout(w_dff_B_5rTwhrzE4_1),.clk(gclk));
	jdff dff_B_tOmEsRbI4_1(.din(w_dff_B_5rTwhrzE4_1),.dout(w_dff_B_tOmEsRbI4_1),.clk(gclk));
	jdff dff_B_JhvV744d7_1(.din(w_dff_B_tOmEsRbI4_1),.dout(w_dff_B_JhvV744d7_1),.clk(gclk));
	jdff dff_B_yn8sG5gV0_1(.din(w_dff_B_JhvV744d7_1),.dout(w_dff_B_yn8sG5gV0_1),.clk(gclk));
	jdff dff_B_rTAhQaIy5_1(.din(n146),.dout(w_dff_B_rTAhQaIy5_1),.clk(gclk));
	jdff dff_B_CmYDUPhJ4_1(.din(w_dff_B_rTAhQaIy5_1),.dout(w_dff_B_CmYDUPhJ4_1),.clk(gclk));
	jdff dff_B_Upm07QLC4_1(.din(w_dff_B_CmYDUPhJ4_1),.dout(w_dff_B_Upm07QLC4_1),.clk(gclk));
	jdff dff_B_proUJcUP0_1(.din(w_dff_B_Upm07QLC4_1),.dout(w_dff_B_proUJcUP0_1),.clk(gclk));
	jdff dff_B_aOGmcA4y5_1(.din(w_dff_B_proUJcUP0_1),.dout(w_dff_B_aOGmcA4y5_1),.clk(gclk));
	jdff dff_B_YcYBpuWM3_1(.din(w_dff_B_aOGmcA4y5_1),.dout(w_dff_B_YcYBpuWM3_1),.clk(gclk));
	jdff dff_B_XRvb5gxl5_1(.din(w_dff_B_YcYBpuWM3_1),.dout(w_dff_B_XRvb5gxl5_1),.clk(gclk));
	jdff dff_B_fwhTfTdf5_1(.din(w_dff_B_XRvb5gxl5_1),.dout(w_dff_B_fwhTfTdf5_1),.clk(gclk));
	jdff dff_B_u4htHALd8_1(.din(w_dff_B_fwhTfTdf5_1),.dout(w_dff_B_u4htHALd8_1),.clk(gclk));
	jdff dff_B_aFy0JXQc9_1(.din(w_dff_B_u4htHALd8_1),.dout(w_dff_B_aFy0JXQc9_1),.clk(gclk));
	jdff dff_B_gW3FhgDb6_1(.din(w_dff_B_aFy0JXQc9_1),.dout(w_dff_B_gW3FhgDb6_1),.clk(gclk));
	jdff dff_B_0aYWqcgP5_1(.din(w_dff_B_gW3FhgDb6_1),.dout(w_dff_B_0aYWqcgP5_1),.clk(gclk));
	jdff dff_B_mpRUR74K0_1(.din(w_dff_B_0aYWqcgP5_1),.dout(w_dff_B_mpRUR74K0_1),.clk(gclk));
	jdff dff_B_c68VdqjT0_1(.din(n184),.dout(w_dff_B_c68VdqjT0_1),.clk(gclk));
	jdff dff_B_HnOS8sg78_1(.din(w_dff_B_c68VdqjT0_1),.dout(w_dff_B_HnOS8sg78_1),.clk(gclk));
	jdff dff_B_87qx4Hrz1_1(.din(w_dff_B_HnOS8sg78_1),.dout(w_dff_B_87qx4Hrz1_1),.clk(gclk));
	jdff dff_B_6cDtbgj96_1(.din(w_dff_B_87qx4Hrz1_1),.dout(w_dff_B_6cDtbgj96_1),.clk(gclk));
	jdff dff_B_30443sQP7_1(.din(w_dff_B_6cDtbgj96_1),.dout(w_dff_B_30443sQP7_1),.clk(gclk));
	jdff dff_B_hYOv1wcl4_1(.din(w_dff_B_30443sQP7_1),.dout(w_dff_B_hYOv1wcl4_1),.clk(gclk));
	jdff dff_B_5y8ARYGA0_1(.din(w_dff_B_hYOv1wcl4_1),.dout(w_dff_B_5y8ARYGA0_1),.clk(gclk));
	jdff dff_B_kxKSSoxD1_1(.din(w_dff_B_5y8ARYGA0_1),.dout(w_dff_B_kxKSSoxD1_1),.clk(gclk));
	jdff dff_B_E57Rn5bm7_1(.din(w_dff_B_kxKSSoxD1_1),.dout(w_dff_B_E57Rn5bm7_1),.clk(gclk));
	jdff dff_B_TyH78zMm2_1(.din(w_dff_B_E57Rn5bm7_1),.dout(w_dff_B_TyH78zMm2_1),.clk(gclk));
	jdff dff_B_KNzEJ7Tm8_1(.din(w_dff_B_TyH78zMm2_1),.dout(w_dff_B_KNzEJ7Tm8_1),.clk(gclk));
	jdff dff_B_iK6D8GFi2_1(.din(w_dff_B_KNzEJ7Tm8_1),.dout(w_dff_B_iK6D8GFi2_1),.clk(gclk));
	jdff dff_B_kIZuIE5P6_1(.din(w_dff_B_iK6D8GFi2_1),.dout(w_dff_B_kIZuIE5P6_1),.clk(gclk));
	jdff dff_B_6CwcnaX19_1(.din(w_dff_B_kIZuIE5P6_1),.dout(w_dff_B_6CwcnaX19_1),.clk(gclk));
	jdff dff_B_qN1tNO329_1(.din(w_dff_B_6CwcnaX19_1),.dout(w_dff_B_qN1tNO329_1),.clk(gclk));
	jdff dff_B_6oZvyY0P2_1(.din(w_dff_B_qN1tNO329_1),.dout(w_dff_B_6oZvyY0P2_1),.clk(gclk));
	jdff dff_B_OxDLKM6A4_1(.din(n227),.dout(w_dff_B_OxDLKM6A4_1),.clk(gclk));
	jdff dff_B_oxBe3N5y3_1(.din(w_dff_B_OxDLKM6A4_1),.dout(w_dff_B_oxBe3N5y3_1),.clk(gclk));
	jdff dff_B_SjcxDkzW4_1(.din(w_dff_B_oxBe3N5y3_1),.dout(w_dff_B_SjcxDkzW4_1),.clk(gclk));
	jdff dff_B_eoiU48Fu6_1(.din(w_dff_B_SjcxDkzW4_1),.dout(w_dff_B_eoiU48Fu6_1),.clk(gclk));
	jdff dff_B_dyi3x6cZ1_1(.din(w_dff_B_eoiU48Fu6_1),.dout(w_dff_B_dyi3x6cZ1_1),.clk(gclk));
	jdff dff_B_MkWRSGne5_1(.din(w_dff_B_dyi3x6cZ1_1),.dout(w_dff_B_MkWRSGne5_1),.clk(gclk));
	jdff dff_B_4nkAMVf06_1(.din(w_dff_B_MkWRSGne5_1),.dout(w_dff_B_4nkAMVf06_1),.clk(gclk));
	jdff dff_B_g9msoVzN5_1(.din(w_dff_B_4nkAMVf06_1),.dout(w_dff_B_g9msoVzN5_1),.clk(gclk));
	jdff dff_B_s1gSvCsW5_1(.din(w_dff_B_g9msoVzN5_1),.dout(w_dff_B_s1gSvCsW5_1),.clk(gclk));
	jdff dff_B_Q4crtiAT9_1(.din(w_dff_B_s1gSvCsW5_1),.dout(w_dff_B_Q4crtiAT9_1),.clk(gclk));
	jdff dff_B_xzZGX8Mf4_1(.din(w_dff_B_Q4crtiAT9_1),.dout(w_dff_B_xzZGX8Mf4_1),.clk(gclk));
	jdff dff_B_8DqYEO6r5_1(.din(w_dff_B_xzZGX8Mf4_1),.dout(w_dff_B_8DqYEO6r5_1),.clk(gclk));
	jdff dff_B_fY2PG9Q50_1(.din(w_dff_B_8DqYEO6r5_1),.dout(w_dff_B_fY2PG9Q50_1),.clk(gclk));
	jdff dff_B_WEE1FcfJ1_1(.din(w_dff_B_fY2PG9Q50_1),.dout(w_dff_B_WEE1FcfJ1_1),.clk(gclk));
	jdff dff_B_3sZshMf70_1(.din(w_dff_B_WEE1FcfJ1_1),.dout(w_dff_B_3sZshMf70_1),.clk(gclk));
	jdff dff_B_ltcvYspb2_1(.din(w_dff_B_3sZshMf70_1),.dout(w_dff_B_ltcvYspb2_1),.clk(gclk));
	jdff dff_B_ZWVFB0pd8_1(.din(w_dff_B_ltcvYspb2_1),.dout(w_dff_B_ZWVFB0pd8_1),.clk(gclk));
	jdff dff_B_2MNp1Nwe7_1(.din(w_dff_B_ZWVFB0pd8_1),.dout(w_dff_B_2MNp1Nwe7_1),.clk(gclk));
	jdff dff_B_4L0Rtspp9_1(.din(w_dff_B_2MNp1Nwe7_1),.dout(w_dff_B_4L0Rtspp9_1),.clk(gclk));
	jdff dff_B_qR4ebJi07_1(.din(n278),.dout(w_dff_B_qR4ebJi07_1),.clk(gclk));
	jdff dff_B_V0FnKv5p0_1(.din(w_dff_B_qR4ebJi07_1),.dout(w_dff_B_V0FnKv5p0_1),.clk(gclk));
	jdff dff_B_0JgJWV5x0_1(.din(w_dff_B_V0FnKv5p0_1),.dout(w_dff_B_0JgJWV5x0_1),.clk(gclk));
	jdff dff_B_fddkuUJa3_1(.din(w_dff_B_0JgJWV5x0_1),.dout(w_dff_B_fddkuUJa3_1),.clk(gclk));
	jdff dff_B_Xpk1Nv1t8_1(.din(w_dff_B_fddkuUJa3_1),.dout(w_dff_B_Xpk1Nv1t8_1),.clk(gclk));
	jdff dff_B_GhC6Xt7D1_1(.din(w_dff_B_Xpk1Nv1t8_1),.dout(w_dff_B_GhC6Xt7D1_1),.clk(gclk));
	jdff dff_B_sLNvUs3e8_1(.din(w_dff_B_GhC6Xt7D1_1),.dout(w_dff_B_sLNvUs3e8_1),.clk(gclk));
	jdff dff_B_GJA0rymt0_1(.din(w_dff_B_sLNvUs3e8_1),.dout(w_dff_B_GJA0rymt0_1),.clk(gclk));
	jdff dff_B_tQMba3r72_1(.din(w_dff_B_GJA0rymt0_1),.dout(w_dff_B_tQMba3r72_1),.clk(gclk));
	jdff dff_B_yXcJsc5P4_1(.din(w_dff_B_tQMba3r72_1),.dout(w_dff_B_yXcJsc5P4_1),.clk(gclk));
	jdff dff_B_shhv4Tye1_1(.din(w_dff_B_yXcJsc5P4_1),.dout(w_dff_B_shhv4Tye1_1),.clk(gclk));
	jdff dff_B_XbVzYS2p8_1(.din(w_dff_B_shhv4Tye1_1),.dout(w_dff_B_XbVzYS2p8_1),.clk(gclk));
	jdff dff_B_37AB7eTi2_1(.din(w_dff_B_XbVzYS2p8_1),.dout(w_dff_B_37AB7eTi2_1),.clk(gclk));
	jdff dff_B_QouHpRJl8_1(.din(w_dff_B_37AB7eTi2_1),.dout(w_dff_B_QouHpRJl8_1),.clk(gclk));
	jdff dff_B_WBt48WoY6_1(.din(w_dff_B_QouHpRJl8_1),.dout(w_dff_B_WBt48WoY6_1),.clk(gclk));
	jdff dff_B_TgCdYDGj2_1(.din(w_dff_B_WBt48WoY6_1),.dout(w_dff_B_TgCdYDGj2_1),.clk(gclk));
	jdff dff_B_5yhAp5iP6_1(.din(w_dff_B_TgCdYDGj2_1),.dout(w_dff_B_5yhAp5iP6_1),.clk(gclk));
	jdff dff_B_dcbNGr257_1(.din(w_dff_B_5yhAp5iP6_1),.dout(w_dff_B_dcbNGr257_1),.clk(gclk));
	jdff dff_B_C4gKgDTb4_1(.din(w_dff_B_dcbNGr257_1),.dout(w_dff_B_C4gKgDTb4_1),.clk(gclk));
	jdff dff_B_t9FLso1H6_1(.din(w_dff_B_C4gKgDTb4_1),.dout(w_dff_B_t9FLso1H6_1),.clk(gclk));
	jdff dff_B_qUc528Iy9_1(.din(w_dff_B_t9FLso1H6_1),.dout(w_dff_B_qUc528Iy9_1),.clk(gclk));
	jdff dff_B_kbrQWFFZ8_1(.din(w_dff_B_qUc528Iy9_1),.dout(w_dff_B_kbrQWFFZ8_1),.clk(gclk));
	jdff dff_B_Yo3uftzK8_1(.din(n336),.dout(w_dff_B_Yo3uftzK8_1),.clk(gclk));
	jdff dff_B_DoPaIDCY3_1(.din(w_dff_B_Yo3uftzK8_1),.dout(w_dff_B_DoPaIDCY3_1),.clk(gclk));
	jdff dff_B_q0g7copr0_1(.din(w_dff_B_DoPaIDCY3_1),.dout(w_dff_B_q0g7copr0_1),.clk(gclk));
	jdff dff_B_r2JZQDKa6_1(.din(w_dff_B_q0g7copr0_1),.dout(w_dff_B_r2JZQDKa6_1),.clk(gclk));
	jdff dff_B_dXVPzbuD2_1(.din(w_dff_B_r2JZQDKa6_1),.dout(w_dff_B_dXVPzbuD2_1),.clk(gclk));
	jdff dff_B_l6ibNJLf0_1(.din(w_dff_B_dXVPzbuD2_1),.dout(w_dff_B_l6ibNJLf0_1),.clk(gclk));
	jdff dff_B_naw2xN6C7_1(.din(w_dff_B_l6ibNJLf0_1),.dout(w_dff_B_naw2xN6C7_1),.clk(gclk));
	jdff dff_B_Nksj6Jr94_1(.din(w_dff_B_naw2xN6C7_1),.dout(w_dff_B_Nksj6Jr94_1),.clk(gclk));
	jdff dff_B_ugtd4XIZ5_1(.din(w_dff_B_Nksj6Jr94_1),.dout(w_dff_B_ugtd4XIZ5_1),.clk(gclk));
	jdff dff_B_FDdO9CcS1_1(.din(w_dff_B_ugtd4XIZ5_1),.dout(w_dff_B_FDdO9CcS1_1),.clk(gclk));
	jdff dff_B_S9iSXbef9_1(.din(w_dff_B_FDdO9CcS1_1),.dout(w_dff_B_S9iSXbef9_1),.clk(gclk));
	jdff dff_B_1dURD0NL3_1(.din(w_dff_B_S9iSXbef9_1),.dout(w_dff_B_1dURD0NL3_1),.clk(gclk));
	jdff dff_B_ICEp6Czp6_1(.din(w_dff_B_1dURD0NL3_1),.dout(w_dff_B_ICEp6Czp6_1),.clk(gclk));
	jdff dff_B_P02rJtwH9_1(.din(w_dff_B_ICEp6Czp6_1),.dout(w_dff_B_P02rJtwH9_1),.clk(gclk));
	jdff dff_B_YDKnW1wb3_1(.din(w_dff_B_P02rJtwH9_1),.dout(w_dff_B_YDKnW1wb3_1),.clk(gclk));
	jdff dff_B_xJZCAaJe5_1(.din(w_dff_B_YDKnW1wb3_1),.dout(w_dff_B_xJZCAaJe5_1),.clk(gclk));
	jdff dff_B_3chGe1H86_1(.din(w_dff_B_xJZCAaJe5_1),.dout(w_dff_B_3chGe1H86_1),.clk(gclk));
	jdff dff_B_toAbKKVg2_1(.din(w_dff_B_3chGe1H86_1),.dout(w_dff_B_toAbKKVg2_1),.clk(gclk));
	jdff dff_B_cSgI2MDr0_1(.din(w_dff_B_toAbKKVg2_1),.dout(w_dff_B_cSgI2MDr0_1),.clk(gclk));
	jdff dff_B_oyzKLNjM5_1(.din(w_dff_B_cSgI2MDr0_1),.dout(w_dff_B_oyzKLNjM5_1),.clk(gclk));
	jdff dff_B_9RlXIP708_1(.din(w_dff_B_oyzKLNjM5_1),.dout(w_dff_B_9RlXIP708_1),.clk(gclk));
	jdff dff_B_aFmFTcfr2_1(.din(w_dff_B_9RlXIP708_1),.dout(w_dff_B_aFmFTcfr2_1),.clk(gclk));
	jdff dff_B_A60PPsHR6_1(.din(w_dff_B_aFmFTcfr2_1),.dout(w_dff_B_A60PPsHR6_1),.clk(gclk));
	jdff dff_B_9GIUgHZk6_1(.din(w_dff_B_A60PPsHR6_1),.dout(w_dff_B_9GIUgHZk6_1),.clk(gclk));
	jdff dff_B_ij0Oc1JR6_1(.din(w_dff_B_9GIUgHZk6_1),.dout(w_dff_B_ij0Oc1JR6_1),.clk(gclk));
	jdff dff_B_S9Jtk2y21_1(.din(n400),.dout(w_dff_B_S9Jtk2y21_1),.clk(gclk));
	jdff dff_B_dCUpUq7u1_1(.din(w_dff_B_S9Jtk2y21_1),.dout(w_dff_B_dCUpUq7u1_1),.clk(gclk));
	jdff dff_B_UK7e50Xv1_1(.din(w_dff_B_dCUpUq7u1_1),.dout(w_dff_B_UK7e50Xv1_1),.clk(gclk));
	jdff dff_B_P2Tdt8LC4_1(.din(w_dff_B_UK7e50Xv1_1),.dout(w_dff_B_P2Tdt8LC4_1),.clk(gclk));
	jdff dff_B_9otp8oGy8_1(.din(w_dff_B_P2Tdt8LC4_1),.dout(w_dff_B_9otp8oGy8_1),.clk(gclk));
	jdff dff_B_QqXGKpnH8_1(.din(w_dff_B_9otp8oGy8_1),.dout(w_dff_B_QqXGKpnH8_1),.clk(gclk));
	jdff dff_B_HhtfZ3Z65_1(.din(w_dff_B_QqXGKpnH8_1),.dout(w_dff_B_HhtfZ3Z65_1),.clk(gclk));
	jdff dff_B_CZorwbve9_1(.din(w_dff_B_HhtfZ3Z65_1),.dout(w_dff_B_CZorwbve9_1),.clk(gclk));
	jdff dff_B_0xT7CAzJ5_1(.din(w_dff_B_CZorwbve9_1),.dout(w_dff_B_0xT7CAzJ5_1),.clk(gclk));
	jdff dff_B_ZKuaVAcV6_1(.din(w_dff_B_0xT7CAzJ5_1),.dout(w_dff_B_ZKuaVAcV6_1),.clk(gclk));
	jdff dff_B_7FgAbger1_1(.din(w_dff_B_ZKuaVAcV6_1),.dout(w_dff_B_7FgAbger1_1),.clk(gclk));
	jdff dff_B_Mzox2m156_1(.din(w_dff_B_7FgAbger1_1),.dout(w_dff_B_Mzox2m156_1),.clk(gclk));
	jdff dff_B_R6CM2PpY5_1(.din(w_dff_B_Mzox2m156_1),.dout(w_dff_B_R6CM2PpY5_1),.clk(gclk));
	jdff dff_B_Q2Jfq5qy7_1(.din(w_dff_B_R6CM2PpY5_1),.dout(w_dff_B_Q2Jfq5qy7_1),.clk(gclk));
	jdff dff_B_BCMy1xRw9_1(.din(w_dff_B_Q2Jfq5qy7_1),.dout(w_dff_B_BCMy1xRw9_1),.clk(gclk));
	jdff dff_B_uYwllOdJ1_1(.din(w_dff_B_BCMy1xRw9_1),.dout(w_dff_B_uYwllOdJ1_1),.clk(gclk));
	jdff dff_B_0HJtWpZl3_1(.din(w_dff_B_uYwllOdJ1_1),.dout(w_dff_B_0HJtWpZl3_1),.clk(gclk));
	jdff dff_B_7mwDdNrj3_1(.din(w_dff_B_0HJtWpZl3_1),.dout(w_dff_B_7mwDdNrj3_1),.clk(gclk));
	jdff dff_B_tgQZfhrL0_1(.din(w_dff_B_7mwDdNrj3_1),.dout(w_dff_B_tgQZfhrL0_1),.clk(gclk));
	jdff dff_B_Ff3fkwRn6_1(.din(w_dff_B_tgQZfhrL0_1),.dout(w_dff_B_Ff3fkwRn6_1),.clk(gclk));
	jdff dff_B_C1KqM5Zq9_1(.din(w_dff_B_Ff3fkwRn6_1),.dout(w_dff_B_C1KqM5Zq9_1),.clk(gclk));
	jdff dff_B_SjOWITER0_1(.din(w_dff_B_C1KqM5Zq9_1),.dout(w_dff_B_SjOWITER0_1),.clk(gclk));
	jdff dff_B_tTrZGqmv4_1(.din(w_dff_B_SjOWITER0_1),.dout(w_dff_B_tTrZGqmv4_1),.clk(gclk));
	jdff dff_B_ld6u9pkR6_1(.din(w_dff_B_tTrZGqmv4_1),.dout(w_dff_B_ld6u9pkR6_1),.clk(gclk));
	jdff dff_B_PWPgwCeY7_1(.din(w_dff_B_ld6u9pkR6_1),.dout(w_dff_B_PWPgwCeY7_1),.clk(gclk));
	jdff dff_B_RWF06jY82_1(.din(w_dff_B_PWPgwCeY7_1),.dout(w_dff_B_RWF06jY82_1),.clk(gclk));
	jdff dff_B_Mcjq08GE7_1(.din(w_dff_B_RWF06jY82_1),.dout(w_dff_B_Mcjq08GE7_1),.clk(gclk));
	jdff dff_B_igGtsUuN6_1(.din(w_dff_B_Mcjq08GE7_1),.dout(w_dff_B_igGtsUuN6_1),.clk(gclk));
	jdff dff_B_eRqVPqVl8_1(.din(n472),.dout(w_dff_B_eRqVPqVl8_1),.clk(gclk));
	jdff dff_B_F8tX5Snw8_1(.din(w_dff_B_eRqVPqVl8_1),.dout(w_dff_B_F8tX5Snw8_1),.clk(gclk));
	jdff dff_B_d2JEphAb6_1(.din(w_dff_B_F8tX5Snw8_1),.dout(w_dff_B_d2JEphAb6_1),.clk(gclk));
	jdff dff_B_xKaeNnVZ8_1(.din(w_dff_B_d2JEphAb6_1),.dout(w_dff_B_xKaeNnVZ8_1),.clk(gclk));
	jdff dff_B_QHvZffoJ2_1(.din(w_dff_B_xKaeNnVZ8_1),.dout(w_dff_B_QHvZffoJ2_1),.clk(gclk));
	jdff dff_B_49orrsqK4_1(.din(w_dff_B_QHvZffoJ2_1),.dout(w_dff_B_49orrsqK4_1),.clk(gclk));
	jdff dff_B_a80AzxBE0_1(.din(w_dff_B_49orrsqK4_1),.dout(w_dff_B_a80AzxBE0_1),.clk(gclk));
	jdff dff_B_U6pCYpOd8_1(.din(w_dff_B_a80AzxBE0_1),.dout(w_dff_B_U6pCYpOd8_1),.clk(gclk));
	jdff dff_B_JgoRaaFd2_1(.din(w_dff_B_U6pCYpOd8_1),.dout(w_dff_B_JgoRaaFd2_1),.clk(gclk));
	jdff dff_B_ROjjjfPG1_1(.din(w_dff_B_JgoRaaFd2_1),.dout(w_dff_B_ROjjjfPG1_1),.clk(gclk));
	jdff dff_B_KBNO8qCX6_1(.din(w_dff_B_ROjjjfPG1_1),.dout(w_dff_B_KBNO8qCX6_1),.clk(gclk));
	jdff dff_B_eiIrvGNx6_1(.din(w_dff_B_KBNO8qCX6_1),.dout(w_dff_B_eiIrvGNx6_1),.clk(gclk));
	jdff dff_B_eKxwp02R0_1(.din(w_dff_B_eiIrvGNx6_1),.dout(w_dff_B_eKxwp02R0_1),.clk(gclk));
	jdff dff_B_j0ZXAfue4_1(.din(w_dff_B_eKxwp02R0_1),.dout(w_dff_B_j0ZXAfue4_1),.clk(gclk));
	jdff dff_B_q4SCnHRo3_1(.din(w_dff_B_j0ZXAfue4_1),.dout(w_dff_B_q4SCnHRo3_1),.clk(gclk));
	jdff dff_B_yqUuNiF27_1(.din(w_dff_B_q4SCnHRo3_1),.dout(w_dff_B_yqUuNiF27_1),.clk(gclk));
	jdff dff_B_6gAHwBbU4_1(.din(w_dff_B_yqUuNiF27_1),.dout(w_dff_B_6gAHwBbU4_1),.clk(gclk));
	jdff dff_B_9uRagnYN2_1(.din(w_dff_B_6gAHwBbU4_1),.dout(w_dff_B_9uRagnYN2_1),.clk(gclk));
	jdff dff_B_yvbGykZv8_1(.din(w_dff_B_9uRagnYN2_1),.dout(w_dff_B_yvbGykZv8_1),.clk(gclk));
	jdff dff_B_Rf84pPBc9_1(.din(w_dff_B_yvbGykZv8_1),.dout(w_dff_B_Rf84pPBc9_1),.clk(gclk));
	jdff dff_B_UaYS03Sm0_1(.din(w_dff_B_Rf84pPBc9_1),.dout(w_dff_B_UaYS03Sm0_1),.clk(gclk));
	jdff dff_B_Lv8aYlRS2_1(.din(w_dff_B_UaYS03Sm0_1),.dout(w_dff_B_Lv8aYlRS2_1),.clk(gclk));
	jdff dff_B_nKxXnrAS9_1(.din(w_dff_B_Lv8aYlRS2_1),.dout(w_dff_B_nKxXnrAS9_1),.clk(gclk));
	jdff dff_B_RI7p9Pgb4_1(.din(w_dff_B_nKxXnrAS9_1),.dout(w_dff_B_RI7p9Pgb4_1),.clk(gclk));
	jdff dff_B_MjVwJuex5_1(.din(w_dff_B_RI7p9Pgb4_1),.dout(w_dff_B_MjVwJuex5_1),.clk(gclk));
	jdff dff_B_IeQ4Mc0m0_1(.din(w_dff_B_MjVwJuex5_1),.dout(w_dff_B_IeQ4Mc0m0_1),.clk(gclk));
	jdff dff_B_gagweyfX1_1(.din(w_dff_B_IeQ4Mc0m0_1),.dout(w_dff_B_gagweyfX1_1),.clk(gclk));
	jdff dff_B_vImXVMkq9_1(.din(w_dff_B_gagweyfX1_1),.dout(w_dff_B_vImXVMkq9_1),.clk(gclk));
	jdff dff_B_Fy0Ny00m6_1(.din(w_dff_B_vImXVMkq9_1),.dout(w_dff_B_Fy0Ny00m6_1),.clk(gclk));
	jdff dff_B_m2D6RYDR1_1(.din(w_dff_B_Fy0Ny00m6_1),.dout(w_dff_B_m2D6RYDR1_1),.clk(gclk));
	jdff dff_B_pkyARCTV1_1(.din(w_dff_B_m2D6RYDR1_1),.dout(w_dff_B_pkyARCTV1_1),.clk(gclk));
	jdff dff_B_wCo3a4uh3_1(.din(n551),.dout(w_dff_B_wCo3a4uh3_1),.clk(gclk));
	jdff dff_B_adX6pACi2_1(.din(w_dff_B_wCo3a4uh3_1),.dout(w_dff_B_adX6pACi2_1),.clk(gclk));
	jdff dff_B_nmUoOWI66_1(.din(w_dff_B_adX6pACi2_1),.dout(w_dff_B_nmUoOWI66_1),.clk(gclk));
	jdff dff_B_SEGCZxaa1_1(.din(w_dff_B_nmUoOWI66_1),.dout(w_dff_B_SEGCZxaa1_1),.clk(gclk));
	jdff dff_B_TSwSvq6g1_1(.din(w_dff_B_SEGCZxaa1_1),.dout(w_dff_B_TSwSvq6g1_1),.clk(gclk));
	jdff dff_B_1mC62K1r5_1(.din(w_dff_B_TSwSvq6g1_1),.dout(w_dff_B_1mC62K1r5_1),.clk(gclk));
	jdff dff_B_mJvpMM5J6_1(.din(w_dff_B_1mC62K1r5_1),.dout(w_dff_B_mJvpMM5J6_1),.clk(gclk));
	jdff dff_B_7g41H3jB4_1(.din(w_dff_B_mJvpMM5J6_1),.dout(w_dff_B_7g41H3jB4_1),.clk(gclk));
	jdff dff_B_SMAtpfSw4_1(.din(w_dff_B_7g41H3jB4_1),.dout(w_dff_B_SMAtpfSw4_1),.clk(gclk));
	jdff dff_B_R6hwYzDj5_1(.din(w_dff_B_SMAtpfSw4_1),.dout(w_dff_B_R6hwYzDj5_1),.clk(gclk));
	jdff dff_B_3bWrEArN2_1(.din(w_dff_B_R6hwYzDj5_1),.dout(w_dff_B_3bWrEArN2_1),.clk(gclk));
	jdff dff_B_vYwylIjI8_1(.din(w_dff_B_3bWrEArN2_1),.dout(w_dff_B_vYwylIjI8_1),.clk(gclk));
	jdff dff_B_p6j5WuPh1_1(.din(w_dff_B_vYwylIjI8_1),.dout(w_dff_B_p6j5WuPh1_1),.clk(gclk));
	jdff dff_B_LM4YDIdJ9_1(.din(w_dff_B_p6j5WuPh1_1),.dout(w_dff_B_LM4YDIdJ9_1),.clk(gclk));
	jdff dff_B_rYnpfGur9_1(.din(w_dff_B_LM4YDIdJ9_1),.dout(w_dff_B_rYnpfGur9_1),.clk(gclk));
	jdff dff_B_WjD0aMZd3_1(.din(w_dff_B_rYnpfGur9_1),.dout(w_dff_B_WjD0aMZd3_1),.clk(gclk));
	jdff dff_B_QPjPjBpq5_1(.din(w_dff_B_WjD0aMZd3_1),.dout(w_dff_B_QPjPjBpq5_1),.clk(gclk));
	jdff dff_B_aDRMe4PM0_1(.din(w_dff_B_QPjPjBpq5_1),.dout(w_dff_B_aDRMe4PM0_1),.clk(gclk));
	jdff dff_B_e4yJMXLs2_1(.din(w_dff_B_aDRMe4PM0_1),.dout(w_dff_B_e4yJMXLs2_1),.clk(gclk));
	jdff dff_B_FbGaAzP94_1(.din(w_dff_B_e4yJMXLs2_1),.dout(w_dff_B_FbGaAzP94_1),.clk(gclk));
	jdff dff_B_kRlxDcRM9_1(.din(w_dff_B_FbGaAzP94_1),.dout(w_dff_B_kRlxDcRM9_1),.clk(gclk));
	jdff dff_B_K1GLlw1c3_1(.din(w_dff_B_kRlxDcRM9_1),.dout(w_dff_B_K1GLlw1c3_1),.clk(gclk));
	jdff dff_B_tpgJ8gqe1_1(.din(w_dff_B_K1GLlw1c3_1),.dout(w_dff_B_tpgJ8gqe1_1),.clk(gclk));
	jdff dff_B_Xe6Nxzol9_1(.din(w_dff_B_tpgJ8gqe1_1),.dout(w_dff_B_Xe6Nxzol9_1),.clk(gclk));
	jdff dff_B_Ba2xc9xv1_1(.din(w_dff_B_Xe6Nxzol9_1),.dout(w_dff_B_Ba2xc9xv1_1),.clk(gclk));
	jdff dff_B_9H4eVJqS1_1(.din(w_dff_B_Ba2xc9xv1_1),.dout(w_dff_B_9H4eVJqS1_1),.clk(gclk));
	jdff dff_B_QxYkCHCB4_1(.din(w_dff_B_9H4eVJqS1_1),.dout(w_dff_B_QxYkCHCB4_1),.clk(gclk));
	jdff dff_B_9DOl2dlq1_1(.din(w_dff_B_QxYkCHCB4_1),.dout(w_dff_B_9DOl2dlq1_1),.clk(gclk));
	jdff dff_B_TLypH8Ai2_1(.din(w_dff_B_9DOl2dlq1_1),.dout(w_dff_B_TLypH8Ai2_1),.clk(gclk));
	jdff dff_B_kCdFSZW74_1(.din(w_dff_B_TLypH8Ai2_1),.dout(w_dff_B_kCdFSZW74_1),.clk(gclk));
	jdff dff_B_7uOlee4C1_1(.din(w_dff_B_kCdFSZW74_1),.dout(w_dff_B_7uOlee4C1_1),.clk(gclk));
	jdff dff_B_EnuMKhEj9_1(.din(w_dff_B_7uOlee4C1_1),.dout(w_dff_B_EnuMKhEj9_1),.clk(gclk));
	jdff dff_B_s0KFe9fj8_1(.din(w_dff_B_EnuMKhEj9_1),.dout(w_dff_B_s0KFe9fj8_1),.clk(gclk));
	jdff dff_B_TVXLodJF2_1(.din(w_dff_B_s0KFe9fj8_1),.dout(w_dff_B_TVXLodJF2_1),.clk(gclk));
	jdff dff_B_KSR3uyc06_1(.din(n637),.dout(w_dff_B_KSR3uyc06_1),.clk(gclk));
	jdff dff_B_chq6mbe15_1(.din(w_dff_B_KSR3uyc06_1),.dout(w_dff_B_chq6mbe15_1),.clk(gclk));
	jdff dff_B_mRhf5AEx1_1(.din(w_dff_B_chq6mbe15_1),.dout(w_dff_B_mRhf5AEx1_1),.clk(gclk));
	jdff dff_B_WB3M9t5M1_1(.din(w_dff_B_mRhf5AEx1_1),.dout(w_dff_B_WB3M9t5M1_1),.clk(gclk));
	jdff dff_B_eVZxnaxN8_1(.din(w_dff_B_WB3M9t5M1_1),.dout(w_dff_B_eVZxnaxN8_1),.clk(gclk));
	jdff dff_B_DdqK9DK56_1(.din(w_dff_B_eVZxnaxN8_1),.dout(w_dff_B_DdqK9DK56_1),.clk(gclk));
	jdff dff_B_3fbI7QoG4_1(.din(w_dff_B_DdqK9DK56_1),.dout(w_dff_B_3fbI7QoG4_1),.clk(gclk));
	jdff dff_B_hD5JL3X31_1(.din(w_dff_B_3fbI7QoG4_1),.dout(w_dff_B_hD5JL3X31_1),.clk(gclk));
	jdff dff_B_T0axEqJp4_1(.din(w_dff_B_hD5JL3X31_1),.dout(w_dff_B_T0axEqJp4_1),.clk(gclk));
	jdff dff_B_1b3jWi2f0_1(.din(w_dff_B_T0axEqJp4_1),.dout(w_dff_B_1b3jWi2f0_1),.clk(gclk));
	jdff dff_B_2WwhoMh78_1(.din(w_dff_B_1b3jWi2f0_1),.dout(w_dff_B_2WwhoMh78_1),.clk(gclk));
	jdff dff_B_wdK9Ir0v9_1(.din(w_dff_B_2WwhoMh78_1),.dout(w_dff_B_wdK9Ir0v9_1),.clk(gclk));
	jdff dff_B_y3iiGRBm9_1(.din(w_dff_B_wdK9Ir0v9_1),.dout(w_dff_B_y3iiGRBm9_1),.clk(gclk));
	jdff dff_B_HdQzN8y37_1(.din(w_dff_B_y3iiGRBm9_1),.dout(w_dff_B_HdQzN8y37_1),.clk(gclk));
	jdff dff_B_cK9Wfv0w3_1(.din(w_dff_B_HdQzN8y37_1),.dout(w_dff_B_cK9Wfv0w3_1),.clk(gclk));
	jdff dff_B_3DTy8LOv2_1(.din(w_dff_B_cK9Wfv0w3_1),.dout(w_dff_B_3DTy8LOv2_1),.clk(gclk));
	jdff dff_B_tLOrQI8M4_1(.din(w_dff_B_3DTy8LOv2_1),.dout(w_dff_B_tLOrQI8M4_1),.clk(gclk));
	jdff dff_B_rKWA5vRt1_1(.din(w_dff_B_tLOrQI8M4_1),.dout(w_dff_B_rKWA5vRt1_1),.clk(gclk));
	jdff dff_B_o87l8aUU6_1(.din(w_dff_B_rKWA5vRt1_1),.dout(w_dff_B_o87l8aUU6_1),.clk(gclk));
	jdff dff_B_LJrdZcoV6_1(.din(w_dff_B_o87l8aUU6_1),.dout(w_dff_B_LJrdZcoV6_1),.clk(gclk));
	jdff dff_B_3iq7gh183_1(.din(w_dff_B_LJrdZcoV6_1),.dout(w_dff_B_3iq7gh183_1),.clk(gclk));
	jdff dff_B_eOcfunNn6_1(.din(w_dff_B_3iq7gh183_1),.dout(w_dff_B_eOcfunNn6_1),.clk(gclk));
	jdff dff_B_M44iwoup2_1(.din(w_dff_B_eOcfunNn6_1),.dout(w_dff_B_M44iwoup2_1),.clk(gclk));
	jdff dff_B_NZWnolkN1_1(.din(w_dff_B_M44iwoup2_1),.dout(w_dff_B_NZWnolkN1_1),.clk(gclk));
	jdff dff_B_HRJjBXxx8_1(.din(w_dff_B_NZWnolkN1_1),.dout(w_dff_B_HRJjBXxx8_1),.clk(gclk));
	jdff dff_B_iOqjcP361_1(.din(w_dff_B_HRJjBXxx8_1),.dout(w_dff_B_iOqjcP361_1),.clk(gclk));
	jdff dff_B_pZsGzh8i1_1(.din(w_dff_B_iOqjcP361_1),.dout(w_dff_B_pZsGzh8i1_1),.clk(gclk));
	jdff dff_B_HiqvZNM75_1(.din(w_dff_B_pZsGzh8i1_1),.dout(w_dff_B_HiqvZNM75_1),.clk(gclk));
	jdff dff_B_58S1dTmc4_1(.din(w_dff_B_HiqvZNM75_1),.dout(w_dff_B_58S1dTmc4_1),.clk(gclk));
	jdff dff_B_AIeOHJQc4_1(.din(w_dff_B_58S1dTmc4_1),.dout(w_dff_B_AIeOHJQc4_1),.clk(gclk));
	jdff dff_B_y7GOh2GO1_1(.din(w_dff_B_AIeOHJQc4_1),.dout(w_dff_B_y7GOh2GO1_1),.clk(gclk));
	jdff dff_B_1GvLUgkk3_1(.din(w_dff_B_y7GOh2GO1_1),.dout(w_dff_B_1GvLUgkk3_1),.clk(gclk));
	jdff dff_B_VKTN7njI5_1(.din(w_dff_B_1GvLUgkk3_1),.dout(w_dff_B_VKTN7njI5_1),.clk(gclk));
	jdff dff_B_ENsKRcJM1_1(.din(w_dff_B_VKTN7njI5_1),.dout(w_dff_B_ENsKRcJM1_1),.clk(gclk));
	jdff dff_B_nLYm0xp18_1(.din(w_dff_B_ENsKRcJM1_1),.dout(w_dff_B_nLYm0xp18_1),.clk(gclk));
	jdff dff_B_nm5uEQUF1_1(.din(w_dff_B_nLYm0xp18_1),.dout(w_dff_B_nm5uEQUF1_1),.clk(gclk));
	jdff dff_B_leim9mt08_1(.din(w_dff_B_nm5uEQUF1_1),.dout(w_dff_B_leim9mt08_1),.clk(gclk));
	jdff dff_B_4OcNLf0j8_1(.din(n730),.dout(w_dff_B_4OcNLf0j8_1),.clk(gclk));
	jdff dff_B_yT9SxfeR2_1(.din(w_dff_B_4OcNLf0j8_1),.dout(w_dff_B_yT9SxfeR2_1),.clk(gclk));
	jdff dff_B_Gpk7ezK60_1(.din(w_dff_B_yT9SxfeR2_1),.dout(w_dff_B_Gpk7ezK60_1),.clk(gclk));
	jdff dff_B_GV3mzXQq6_1(.din(w_dff_B_Gpk7ezK60_1),.dout(w_dff_B_GV3mzXQq6_1),.clk(gclk));
	jdff dff_B_eRvdZ90j5_1(.din(w_dff_B_GV3mzXQq6_1),.dout(w_dff_B_eRvdZ90j5_1),.clk(gclk));
	jdff dff_B_FaZyKaHO6_1(.din(w_dff_B_eRvdZ90j5_1),.dout(w_dff_B_FaZyKaHO6_1),.clk(gclk));
	jdff dff_B_Q1e6kKlY1_1(.din(w_dff_B_FaZyKaHO6_1),.dout(w_dff_B_Q1e6kKlY1_1),.clk(gclk));
	jdff dff_B_HjgawN2L4_1(.din(w_dff_B_Q1e6kKlY1_1),.dout(w_dff_B_HjgawN2L4_1),.clk(gclk));
	jdff dff_B_Fwoz4kiq8_1(.din(w_dff_B_HjgawN2L4_1),.dout(w_dff_B_Fwoz4kiq8_1),.clk(gclk));
	jdff dff_B_m5fpVlLg8_1(.din(w_dff_B_Fwoz4kiq8_1),.dout(w_dff_B_m5fpVlLg8_1),.clk(gclk));
	jdff dff_B_vzpSX2mR4_1(.din(w_dff_B_m5fpVlLg8_1),.dout(w_dff_B_vzpSX2mR4_1),.clk(gclk));
	jdff dff_B_GWrfhdjj7_1(.din(w_dff_B_vzpSX2mR4_1),.dout(w_dff_B_GWrfhdjj7_1),.clk(gclk));
	jdff dff_B_azPfQlIz8_1(.din(w_dff_B_GWrfhdjj7_1),.dout(w_dff_B_azPfQlIz8_1),.clk(gclk));
	jdff dff_B_RojonLnm3_1(.din(w_dff_B_azPfQlIz8_1),.dout(w_dff_B_RojonLnm3_1),.clk(gclk));
	jdff dff_B_0svLXzdR2_1(.din(w_dff_B_RojonLnm3_1),.dout(w_dff_B_0svLXzdR2_1),.clk(gclk));
	jdff dff_B_6HtfvSOS6_1(.din(w_dff_B_0svLXzdR2_1),.dout(w_dff_B_6HtfvSOS6_1),.clk(gclk));
	jdff dff_B_4X46y0Zx8_1(.din(w_dff_B_6HtfvSOS6_1),.dout(w_dff_B_4X46y0Zx8_1),.clk(gclk));
	jdff dff_B_9XwRkT5m5_1(.din(w_dff_B_4X46y0Zx8_1),.dout(w_dff_B_9XwRkT5m5_1),.clk(gclk));
	jdff dff_B_JDgGXXA50_1(.din(w_dff_B_9XwRkT5m5_1),.dout(w_dff_B_JDgGXXA50_1),.clk(gclk));
	jdff dff_B_bJFpnRci9_1(.din(w_dff_B_JDgGXXA50_1),.dout(w_dff_B_bJFpnRci9_1),.clk(gclk));
	jdff dff_B_XbohPpsD3_1(.din(w_dff_B_bJFpnRci9_1),.dout(w_dff_B_XbohPpsD3_1),.clk(gclk));
	jdff dff_B_N8lpKHza2_1(.din(w_dff_B_XbohPpsD3_1),.dout(w_dff_B_N8lpKHza2_1),.clk(gclk));
	jdff dff_B_dvW6l90d8_1(.din(w_dff_B_N8lpKHza2_1),.dout(w_dff_B_dvW6l90d8_1),.clk(gclk));
	jdff dff_B_d6sjpxFq3_1(.din(w_dff_B_dvW6l90d8_1),.dout(w_dff_B_d6sjpxFq3_1),.clk(gclk));
	jdff dff_B_gdriOl6g3_1(.din(w_dff_B_d6sjpxFq3_1),.dout(w_dff_B_gdriOl6g3_1),.clk(gclk));
	jdff dff_B_fo7zCS5x4_1(.din(w_dff_B_gdriOl6g3_1),.dout(w_dff_B_fo7zCS5x4_1),.clk(gclk));
	jdff dff_B_7bwNHSSY3_1(.din(w_dff_B_fo7zCS5x4_1),.dout(w_dff_B_7bwNHSSY3_1),.clk(gclk));
	jdff dff_B_hrismID71_1(.din(w_dff_B_7bwNHSSY3_1),.dout(w_dff_B_hrismID71_1),.clk(gclk));
	jdff dff_B_XrvHtSpy0_1(.din(w_dff_B_hrismID71_1),.dout(w_dff_B_XrvHtSpy0_1),.clk(gclk));
	jdff dff_B_qP46jQbq7_1(.din(w_dff_B_XrvHtSpy0_1),.dout(w_dff_B_qP46jQbq7_1),.clk(gclk));
	jdff dff_B_Lp0w4pKz5_1(.din(w_dff_B_qP46jQbq7_1),.dout(w_dff_B_Lp0w4pKz5_1),.clk(gclk));
	jdff dff_B_JaaTS2r72_1(.din(w_dff_B_Lp0w4pKz5_1),.dout(w_dff_B_JaaTS2r72_1),.clk(gclk));
	jdff dff_B_xVwlfayq0_1(.din(w_dff_B_JaaTS2r72_1),.dout(w_dff_B_xVwlfayq0_1),.clk(gclk));
	jdff dff_B_FPu8Wwva5_1(.din(w_dff_B_xVwlfayq0_1),.dout(w_dff_B_FPu8Wwva5_1),.clk(gclk));
	jdff dff_B_1oXggIs45_1(.din(w_dff_B_FPu8Wwva5_1),.dout(w_dff_B_1oXggIs45_1),.clk(gclk));
	jdff dff_B_KPVkZZ1V2_1(.din(w_dff_B_1oXggIs45_1),.dout(w_dff_B_KPVkZZ1V2_1),.clk(gclk));
	jdff dff_B_WDY1Kifv8_1(.din(w_dff_B_KPVkZZ1V2_1),.dout(w_dff_B_WDY1Kifv8_1),.clk(gclk));
	jdff dff_B_7kyrPZGY8_1(.din(w_dff_B_WDY1Kifv8_1),.dout(w_dff_B_7kyrPZGY8_1),.clk(gclk));
	jdff dff_B_lFBVzJRX8_1(.din(w_dff_B_7kyrPZGY8_1),.dout(w_dff_B_lFBVzJRX8_1),.clk(gclk));
	jdff dff_B_j0VSIXt63_1(.din(w_dff_B_lFBVzJRX8_1),.dout(w_dff_B_j0VSIXt63_1),.clk(gclk));
	jdff dff_B_xPBzHC7Q5_1(.din(n830),.dout(w_dff_B_xPBzHC7Q5_1),.clk(gclk));
	jdff dff_B_hONsmt908_1(.din(w_dff_B_xPBzHC7Q5_1),.dout(w_dff_B_hONsmt908_1),.clk(gclk));
	jdff dff_B_FVWJcb5u2_1(.din(w_dff_B_hONsmt908_1),.dout(w_dff_B_FVWJcb5u2_1),.clk(gclk));
	jdff dff_B_3SjG0wVu9_1(.din(w_dff_B_FVWJcb5u2_1),.dout(w_dff_B_3SjG0wVu9_1),.clk(gclk));
	jdff dff_B_A1I68soy3_1(.din(w_dff_B_3SjG0wVu9_1),.dout(w_dff_B_A1I68soy3_1),.clk(gclk));
	jdff dff_B_8JRnPKiX5_1(.din(w_dff_B_A1I68soy3_1),.dout(w_dff_B_8JRnPKiX5_1),.clk(gclk));
	jdff dff_B_tDYKRwZI0_1(.din(w_dff_B_8JRnPKiX5_1),.dout(w_dff_B_tDYKRwZI0_1),.clk(gclk));
	jdff dff_B_hBPbpSF41_1(.din(w_dff_B_tDYKRwZI0_1),.dout(w_dff_B_hBPbpSF41_1),.clk(gclk));
	jdff dff_B_kihbHujo9_1(.din(w_dff_B_hBPbpSF41_1),.dout(w_dff_B_kihbHujo9_1),.clk(gclk));
	jdff dff_B_G1s9zMRU0_1(.din(w_dff_B_kihbHujo9_1),.dout(w_dff_B_G1s9zMRU0_1),.clk(gclk));
	jdff dff_B_hcVLaKD18_1(.din(w_dff_B_G1s9zMRU0_1),.dout(w_dff_B_hcVLaKD18_1),.clk(gclk));
	jdff dff_B_tril6glz3_1(.din(w_dff_B_hcVLaKD18_1),.dout(w_dff_B_tril6glz3_1),.clk(gclk));
	jdff dff_B_f9GTB9Qv4_1(.din(w_dff_B_tril6glz3_1),.dout(w_dff_B_f9GTB9Qv4_1),.clk(gclk));
	jdff dff_B_5nRltPhm2_1(.din(w_dff_B_f9GTB9Qv4_1),.dout(w_dff_B_5nRltPhm2_1),.clk(gclk));
	jdff dff_B_TTlbWxqY0_1(.din(w_dff_B_5nRltPhm2_1),.dout(w_dff_B_TTlbWxqY0_1),.clk(gclk));
	jdff dff_B_6A8co7Y52_1(.din(w_dff_B_TTlbWxqY0_1),.dout(w_dff_B_6A8co7Y52_1),.clk(gclk));
	jdff dff_B_CrUABUte0_1(.din(w_dff_B_6A8co7Y52_1),.dout(w_dff_B_CrUABUte0_1),.clk(gclk));
	jdff dff_B_r7vsu1Nx8_1(.din(w_dff_B_CrUABUte0_1),.dout(w_dff_B_r7vsu1Nx8_1),.clk(gclk));
	jdff dff_B_1VqjD5nW2_1(.din(w_dff_B_r7vsu1Nx8_1),.dout(w_dff_B_1VqjD5nW2_1),.clk(gclk));
	jdff dff_B_J5Fk6Dix5_1(.din(w_dff_B_1VqjD5nW2_1),.dout(w_dff_B_J5Fk6Dix5_1),.clk(gclk));
	jdff dff_B_IIvwCoP80_1(.din(w_dff_B_J5Fk6Dix5_1),.dout(w_dff_B_IIvwCoP80_1),.clk(gclk));
	jdff dff_B_hnLLpKD29_1(.din(w_dff_B_IIvwCoP80_1),.dout(w_dff_B_hnLLpKD29_1),.clk(gclk));
	jdff dff_B_n8LY6GXK0_1(.din(w_dff_B_hnLLpKD29_1),.dout(w_dff_B_n8LY6GXK0_1),.clk(gclk));
	jdff dff_B_VqgwCVqI3_1(.din(w_dff_B_n8LY6GXK0_1),.dout(w_dff_B_VqgwCVqI3_1),.clk(gclk));
	jdff dff_B_5l941F006_1(.din(w_dff_B_VqgwCVqI3_1),.dout(w_dff_B_5l941F006_1),.clk(gclk));
	jdff dff_B_ukXY0LS96_1(.din(w_dff_B_5l941F006_1),.dout(w_dff_B_ukXY0LS96_1),.clk(gclk));
	jdff dff_B_DvN4zRQK4_1(.din(w_dff_B_ukXY0LS96_1),.dout(w_dff_B_DvN4zRQK4_1),.clk(gclk));
	jdff dff_B_bNcWidkD1_1(.din(w_dff_B_DvN4zRQK4_1),.dout(w_dff_B_bNcWidkD1_1),.clk(gclk));
	jdff dff_B_e8CpMAeq7_1(.din(w_dff_B_bNcWidkD1_1),.dout(w_dff_B_e8CpMAeq7_1),.clk(gclk));
	jdff dff_B_GLpHVpJ71_1(.din(w_dff_B_e8CpMAeq7_1),.dout(w_dff_B_GLpHVpJ71_1),.clk(gclk));
	jdff dff_B_w224alA12_1(.din(w_dff_B_GLpHVpJ71_1),.dout(w_dff_B_w224alA12_1),.clk(gclk));
	jdff dff_B_lX1idXQ92_1(.din(w_dff_B_w224alA12_1),.dout(w_dff_B_lX1idXQ92_1),.clk(gclk));
	jdff dff_B_X10zzGzj2_1(.din(w_dff_B_lX1idXQ92_1),.dout(w_dff_B_X10zzGzj2_1),.clk(gclk));
	jdff dff_B_omWaHplO9_1(.din(w_dff_B_X10zzGzj2_1),.dout(w_dff_B_omWaHplO9_1),.clk(gclk));
	jdff dff_B_Y6maJJWP2_1(.din(w_dff_B_omWaHplO9_1),.dout(w_dff_B_Y6maJJWP2_1),.clk(gclk));
	jdff dff_B_LMy4L1Qn7_1(.din(w_dff_B_Y6maJJWP2_1),.dout(w_dff_B_LMy4L1Qn7_1),.clk(gclk));
	jdff dff_B_ls9Yo28U4_1(.din(w_dff_B_LMy4L1Qn7_1),.dout(w_dff_B_ls9Yo28U4_1),.clk(gclk));
	jdff dff_B_vrSgv7pe0_1(.din(w_dff_B_ls9Yo28U4_1),.dout(w_dff_B_vrSgv7pe0_1),.clk(gclk));
	jdff dff_B_Z4eQIBYN1_1(.din(w_dff_B_vrSgv7pe0_1),.dout(w_dff_B_Z4eQIBYN1_1),.clk(gclk));
	jdff dff_B_uZtKOEGq0_1(.din(w_dff_B_Z4eQIBYN1_1),.dout(w_dff_B_uZtKOEGq0_1),.clk(gclk));
	jdff dff_B_xiNNoxFZ7_1(.din(w_dff_B_uZtKOEGq0_1),.dout(w_dff_B_xiNNoxFZ7_1),.clk(gclk));
	jdff dff_B_w2Kbh6uf6_1(.din(w_dff_B_xiNNoxFZ7_1),.dout(w_dff_B_w2Kbh6uf6_1),.clk(gclk));
	jdff dff_B_fP7WTlcY5_1(.din(w_dff_B_w2Kbh6uf6_1),.dout(w_dff_B_fP7WTlcY5_1),.clk(gclk));
	jdff dff_B_lQr3XVAK2_0(.din(n1327),.dout(w_dff_B_lQr3XVAK2_0),.clk(gclk));
	jdff dff_B_jaXDnHrE5_1(.din(n1842),.dout(w_dff_B_jaXDnHrE5_1),.clk(gclk));
	jdff dff_B_9wBv86Ac4_1(.din(w_dff_B_jaXDnHrE5_1),.dout(w_dff_B_9wBv86Ac4_1),.clk(gclk));
	jdff dff_B_fvAVpMFh9_1(.din(w_dff_B_9wBv86Ac4_1),.dout(w_dff_B_fvAVpMFh9_1),.clk(gclk));
	jdff dff_B_vJGQTYef9_1(.din(w_dff_B_fvAVpMFh9_1),.dout(w_dff_B_vJGQTYef9_1),.clk(gclk));
	jdff dff_B_tkLLvKi47_1(.din(w_dff_B_vJGQTYef9_1),.dout(w_dff_B_tkLLvKi47_1),.clk(gclk));
	jdff dff_B_u5sNaIjK6_1(.din(w_dff_B_tkLLvKi47_1),.dout(w_dff_B_u5sNaIjK6_1),.clk(gclk));
	jdff dff_B_nPcle7br3_1(.din(w_dff_B_u5sNaIjK6_1),.dout(w_dff_B_nPcle7br3_1),.clk(gclk));
	jdff dff_B_yBkNdTAm7_1(.din(w_dff_B_nPcle7br3_1),.dout(w_dff_B_yBkNdTAm7_1),.clk(gclk));
	jdff dff_B_aBIokkte6_1(.din(w_dff_B_yBkNdTAm7_1),.dout(w_dff_B_aBIokkte6_1),.clk(gclk));
	jdff dff_B_tCAIVqgo6_1(.din(w_dff_B_aBIokkte6_1),.dout(w_dff_B_tCAIVqgo6_1),.clk(gclk));
	jdff dff_B_kiUSm16c5_1(.din(w_dff_B_tCAIVqgo6_1),.dout(w_dff_B_kiUSm16c5_1),.clk(gclk));
	jdff dff_B_HxyBNYEG0_1(.din(w_dff_B_kiUSm16c5_1),.dout(w_dff_B_HxyBNYEG0_1),.clk(gclk));
	jdff dff_B_dZMtG6911_1(.din(w_dff_B_HxyBNYEG0_1),.dout(w_dff_B_dZMtG6911_1),.clk(gclk));
	jdff dff_B_hzE7q2Sk5_0(.din(n1850),.dout(w_dff_B_hzE7q2Sk5_0),.clk(gclk));
	jdff dff_B_M75Ir0bP4_0(.din(w_dff_B_hzE7q2Sk5_0),.dout(w_dff_B_M75Ir0bP4_0),.clk(gclk));
	jdff dff_B_uR6tgjXS1_0(.din(w_dff_B_M75Ir0bP4_0),.dout(w_dff_B_uR6tgjXS1_0),.clk(gclk));
	jdff dff_B_o6DSENKN7_0(.din(w_dff_B_uR6tgjXS1_0),.dout(w_dff_B_o6DSENKN7_0),.clk(gclk));
	jdff dff_B_1VrmdnFO5_0(.din(w_dff_B_o6DSENKN7_0),.dout(w_dff_B_1VrmdnFO5_0),.clk(gclk));
	jdff dff_B_wBAEPCUH7_0(.din(w_dff_B_1VrmdnFO5_0),.dout(w_dff_B_wBAEPCUH7_0),.clk(gclk));
	jdff dff_B_XMCAzU8D6_0(.din(w_dff_B_wBAEPCUH7_0),.dout(w_dff_B_XMCAzU8D6_0),.clk(gclk));
	jdff dff_B_TvpWawKz1_0(.din(w_dff_B_XMCAzU8D6_0),.dout(w_dff_B_TvpWawKz1_0),.clk(gclk));
	jdff dff_B_wkIjs8mN0_0(.din(w_dff_B_TvpWawKz1_0),.dout(w_dff_B_wkIjs8mN0_0),.clk(gclk));
	jdff dff_B_xwv9vb1o5_0(.din(w_dff_B_wkIjs8mN0_0),.dout(w_dff_B_xwv9vb1o5_0),.clk(gclk));
	jdff dff_B_r6oV5yp74_0(.din(w_dff_B_xwv9vb1o5_0),.dout(w_dff_B_r6oV5yp74_0),.clk(gclk));
	jdff dff_B_rGI5WH8Q5_1(.din(n1845),.dout(w_dff_B_rGI5WH8Q5_1),.clk(gclk));
	jdff dff_B_KOkLL7AE8_1(.din(w_dff_B_rGI5WH8Q5_1),.dout(w_dff_B_KOkLL7AE8_1),.clk(gclk));
	jdff dff_B_ePLJXcwg3_1(.din(w_dff_B_KOkLL7AE8_1),.dout(w_dff_B_ePLJXcwg3_1),.clk(gclk));
	jdff dff_B_hUuTLsCD0_1(.din(w_dff_B_ePLJXcwg3_1),.dout(w_dff_B_hUuTLsCD0_1),.clk(gclk));
	jdff dff_B_S0A38z4p1_1(.din(w_dff_B_hUuTLsCD0_1),.dout(w_dff_B_S0A38z4p1_1),.clk(gclk));
	jdff dff_B_EGWBvchY7_1(.din(w_dff_B_S0A38z4p1_1),.dout(w_dff_B_EGWBvchY7_1),.clk(gclk));
	jdff dff_B_xNPsICqc2_1(.din(w_dff_B_EGWBvchY7_1),.dout(w_dff_B_xNPsICqc2_1),.clk(gclk));
	jdff dff_B_ATuq1jgw3_1(.din(w_dff_B_xNPsICqc2_1),.dout(w_dff_B_ATuq1jgw3_1),.clk(gclk));
	jdff dff_B_9yHiEcDe7_1(.din(w_dff_B_ATuq1jgw3_1),.dout(w_dff_B_9yHiEcDe7_1),.clk(gclk));
	jdff dff_B_AIQlOzkn9_1(.din(w_dff_B_9yHiEcDe7_1),.dout(w_dff_B_AIQlOzkn9_1),.clk(gclk));
	jdff dff_B_qcB4i5Lp4_1(.din(w_dff_B_AIQlOzkn9_1),.dout(w_dff_B_qcB4i5Lp4_1),.clk(gclk));
	jdff dff_B_iWYRQ4ys9_0(.din(n1846),.dout(w_dff_B_iWYRQ4ys9_0),.clk(gclk));
	jdff dff_B_9V90CMJQ5_0(.din(w_dff_B_iWYRQ4ys9_0),.dout(w_dff_B_9V90CMJQ5_0),.clk(gclk));
	jdff dff_B_ILgibT5O4_0(.din(w_dff_B_9V90CMJQ5_0),.dout(w_dff_B_ILgibT5O4_0),.clk(gclk));
	jdff dff_B_j6mQpogF4_0(.din(w_dff_B_ILgibT5O4_0),.dout(w_dff_B_j6mQpogF4_0),.clk(gclk));
	jdff dff_B_M99bmLne9_0(.din(w_dff_B_j6mQpogF4_0),.dout(w_dff_B_M99bmLne9_0),.clk(gclk));
	jdff dff_B_0JsVgMXC5_0(.din(w_dff_B_M99bmLne9_0),.dout(w_dff_B_0JsVgMXC5_0),.clk(gclk));
	jdff dff_B_qXfIvdzc3_0(.din(w_dff_B_0JsVgMXC5_0),.dout(w_dff_B_qXfIvdzc3_0),.clk(gclk));
	jdff dff_B_vlFBUAih6_0(.din(w_dff_B_qXfIvdzc3_0),.dout(w_dff_B_vlFBUAih6_0),.clk(gclk));
	jdff dff_B_Fso2apb72_0(.din(w_dff_B_vlFBUAih6_0),.dout(w_dff_B_Fso2apb72_0),.clk(gclk));
	jdff dff_B_Mr2wOWV55_0(.din(w_dff_B_Fso2apb72_0),.dout(w_dff_B_Mr2wOWV55_0),.clk(gclk));
	jdff dff_B_EnAgxTet0_1(.din(n1821),.dout(w_dff_B_EnAgxTet0_1),.clk(gclk));
	jdff dff_B_7uuecxy63_1(.din(w_dff_B_EnAgxTet0_1),.dout(w_dff_B_7uuecxy63_1),.clk(gclk));
	jdff dff_B_Nve3TPCf6_1(.din(w_dff_B_7uuecxy63_1),.dout(w_dff_B_Nve3TPCf6_1),.clk(gclk));
	jdff dff_B_dVl77WSQ0_1(.din(w_dff_B_Nve3TPCf6_1),.dout(w_dff_B_dVl77WSQ0_1),.clk(gclk));
	jdff dff_B_UgyF34N34_1(.din(w_dff_B_dVl77WSQ0_1),.dout(w_dff_B_UgyF34N34_1),.clk(gclk));
	jdff dff_B_vuOcyOYu8_1(.din(w_dff_B_UgyF34N34_1),.dout(w_dff_B_vuOcyOYu8_1),.clk(gclk));
	jdff dff_B_dW6bcvXe1_1(.din(w_dff_B_vuOcyOYu8_1),.dout(w_dff_B_dW6bcvXe1_1),.clk(gclk));
	jdff dff_B_fFrwz9Kn1_1(.din(w_dff_B_dW6bcvXe1_1),.dout(w_dff_B_fFrwz9Kn1_1),.clk(gclk));
	jdff dff_B_3aU9GhEG7_1(.din(w_dff_B_fFrwz9Kn1_1),.dout(w_dff_B_3aU9GhEG7_1),.clk(gclk));
	jdff dff_B_oepmN3JF2_1(.din(w_dff_B_3aU9GhEG7_1),.dout(w_dff_B_oepmN3JF2_1),.clk(gclk));
	jdff dff_B_j2KrgK254_1(.din(w_dff_B_oepmN3JF2_1),.dout(w_dff_B_j2KrgK254_1),.clk(gclk));
	jdff dff_B_dA0HCEG48_0(.din(n1822),.dout(w_dff_B_dA0HCEG48_0),.clk(gclk));
	jdff dff_B_FrlL5QKw2_0(.din(w_dff_B_dA0HCEG48_0),.dout(w_dff_B_FrlL5QKw2_0),.clk(gclk));
	jdff dff_B_IJ6pwduu0_0(.din(w_dff_B_FrlL5QKw2_0),.dout(w_dff_B_IJ6pwduu0_0),.clk(gclk));
	jdff dff_B_T53wAaOn3_0(.din(w_dff_B_IJ6pwduu0_0),.dout(w_dff_B_T53wAaOn3_0),.clk(gclk));
	jdff dff_B_tdxjmLkO7_0(.din(w_dff_B_T53wAaOn3_0),.dout(w_dff_B_tdxjmLkO7_0),.clk(gclk));
	jdff dff_B_SkyAzguN9_0(.din(w_dff_B_tdxjmLkO7_0),.dout(w_dff_B_SkyAzguN9_0),.clk(gclk));
	jdff dff_B_LpsxhZDt1_0(.din(w_dff_B_SkyAzguN9_0),.dout(w_dff_B_LpsxhZDt1_0),.clk(gclk));
	jdff dff_B_GuIOCIJb2_0(.din(w_dff_B_LpsxhZDt1_0),.dout(w_dff_B_GuIOCIJb2_0),.clk(gclk));
	jdff dff_B_KkbU6eaE5_0(.din(w_dff_B_GuIOCIJb2_0),.dout(w_dff_B_KkbU6eaE5_0),.clk(gclk));
	jdff dff_B_S11eF9xM5_0(.din(w_dff_B_KkbU6eaE5_0),.dout(w_dff_B_S11eF9xM5_0),.clk(gclk));
	jdff dff_B_wMnVA5vf0_1(.din(n1795),.dout(w_dff_B_wMnVA5vf0_1),.clk(gclk));
	jdff dff_B_YRmfgDlQ7_1(.din(w_dff_B_wMnVA5vf0_1),.dout(w_dff_B_YRmfgDlQ7_1),.clk(gclk));
	jdff dff_B_pqd1WIft9_1(.din(w_dff_B_YRmfgDlQ7_1),.dout(w_dff_B_pqd1WIft9_1),.clk(gclk));
	jdff dff_B_kiTDo6Kq4_1(.din(w_dff_B_pqd1WIft9_1),.dout(w_dff_B_kiTDo6Kq4_1),.clk(gclk));
	jdff dff_B_YX0j1f3L9_1(.din(w_dff_B_kiTDo6Kq4_1),.dout(w_dff_B_YX0j1f3L9_1),.clk(gclk));
	jdff dff_B_29pD1IvM8_1(.din(w_dff_B_YX0j1f3L9_1),.dout(w_dff_B_29pD1IvM8_1),.clk(gclk));
	jdff dff_B_3g9DAuUi8_1(.din(w_dff_B_29pD1IvM8_1),.dout(w_dff_B_3g9DAuUi8_1),.clk(gclk));
	jdff dff_B_U9vd2RPF0_1(.din(w_dff_B_3g9DAuUi8_1),.dout(w_dff_B_U9vd2RPF0_1),.clk(gclk));
	jdff dff_B_CVMHTWgo6_1(.din(w_dff_B_U9vd2RPF0_1),.dout(w_dff_B_CVMHTWgo6_1),.clk(gclk));
	jdff dff_B_ZL5KMlUy4_1(.din(w_dff_B_CVMHTWgo6_1),.dout(w_dff_B_ZL5KMlUy4_1),.clk(gclk));
	jdff dff_B_IOofLOGl5_1(.din(w_dff_B_ZL5KMlUy4_1),.dout(w_dff_B_IOofLOGl5_1),.clk(gclk));
	jdff dff_B_jd8bIYSw8_0(.din(n1796),.dout(w_dff_B_jd8bIYSw8_0),.clk(gclk));
	jdff dff_B_KPUmYetE3_0(.din(w_dff_B_jd8bIYSw8_0),.dout(w_dff_B_KPUmYetE3_0),.clk(gclk));
	jdff dff_B_VMl6ZMXJ6_0(.din(w_dff_B_KPUmYetE3_0),.dout(w_dff_B_VMl6ZMXJ6_0),.clk(gclk));
	jdff dff_B_fqJm61u26_0(.din(w_dff_B_VMl6ZMXJ6_0),.dout(w_dff_B_fqJm61u26_0),.clk(gclk));
	jdff dff_B_V9aPycDz6_0(.din(w_dff_B_fqJm61u26_0),.dout(w_dff_B_V9aPycDz6_0),.clk(gclk));
	jdff dff_B_I7mBGZew2_0(.din(w_dff_B_V9aPycDz6_0),.dout(w_dff_B_I7mBGZew2_0),.clk(gclk));
	jdff dff_B_OEd8LnQS6_0(.din(w_dff_B_I7mBGZew2_0),.dout(w_dff_B_OEd8LnQS6_0),.clk(gclk));
	jdff dff_B_ss3azBuR8_0(.din(w_dff_B_OEd8LnQS6_0),.dout(w_dff_B_ss3azBuR8_0),.clk(gclk));
	jdff dff_B_bZAGdl4l4_0(.din(w_dff_B_ss3azBuR8_0),.dout(w_dff_B_bZAGdl4l4_0),.clk(gclk));
	jdff dff_B_BE1ml2kz8_0(.din(w_dff_B_bZAGdl4l4_0),.dout(w_dff_B_BE1ml2kz8_0),.clk(gclk));
	jdff dff_B_hYszWuVb0_1(.din(n1762),.dout(w_dff_B_hYszWuVb0_1),.clk(gclk));
	jdff dff_B_e55ES3g08_1(.din(w_dff_B_hYszWuVb0_1),.dout(w_dff_B_e55ES3g08_1),.clk(gclk));
	jdff dff_B_qY7AI4fe1_1(.din(w_dff_B_e55ES3g08_1),.dout(w_dff_B_qY7AI4fe1_1),.clk(gclk));
	jdff dff_B_YByykTAO4_1(.din(w_dff_B_qY7AI4fe1_1),.dout(w_dff_B_YByykTAO4_1),.clk(gclk));
	jdff dff_B_pOUOZQxt6_1(.din(w_dff_B_YByykTAO4_1),.dout(w_dff_B_pOUOZQxt6_1),.clk(gclk));
	jdff dff_B_pWBfprob9_1(.din(w_dff_B_pOUOZQxt6_1),.dout(w_dff_B_pWBfprob9_1),.clk(gclk));
	jdff dff_B_dJN2MV1C9_1(.din(w_dff_B_pWBfprob9_1),.dout(w_dff_B_dJN2MV1C9_1),.clk(gclk));
	jdff dff_B_VGF49Dzw2_1(.din(w_dff_B_dJN2MV1C9_1),.dout(w_dff_B_VGF49Dzw2_1),.clk(gclk));
	jdff dff_B_aAjyqMuW4_1(.din(w_dff_B_VGF49Dzw2_1),.dout(w_dff_B_aAjyqMuW4_1),.clk(gclk));
	jdff dff_B_C10XhRCQ3_1(.din(w_dff_B_aAjyqMuW4_1),.dout(w_dff_B_C10XhRCQ3_1),.clk(gclk));
	jdff dff_B_kjNYoeB98_1(.din(w_dff_B_C10XhRCQ3_1),.dout(w_dff_B_kjNYoeB98_1),.clk(gclk));
	jdff dff_B_I9vmdZhI1_0(.din(n1763),.dout(w_dff_B_I9vmdZhI1_0),.clk(gclk));
	jdff dff_B_9Thgu8DF7_0(.din(w_dff_B_I9vmdZhI1_0),.dout(w_dff_B_9Thgu8DF7_0),.clk(gclk));
	jdff dff_B_qODYfE2y9_0(.din(w_dff_B_9Thgu8DF7_0),.dout(w_dff_B_qODYfE2y9_0),.clk(gclk));
	jdff dff_B_9f9ANNgz1_0(.din(w_dff_B_qODYfE2y9_0),.dout(w_dff_B_9f9ANNgz1_0),.clk(gclk));
	jdff dff_B_AYakFLww5_0(.din(w_dff_B_9f9ANNgz1_0),.dout(w_dff_B_AYakFLww5_0),.clk(gclk));
	jdff dff_B_eCcqk5O08_0(.din(w_dff_B_AYakFLww5_0),.dout(w_dff_B_eCcqk5O08_0),.clk(gclk));
	jdff dff_B_grq4Gk7X6_0(.din(w_dff_B_eCcqk5O08_0),.dout(w_dff_B_grq4Gk7X6_0),.clk(gclk));
	jdff dff_B_XJeiFyyT6_0(.din(w_dff_B_grq4Gk7X6_0),.dout(w_dff_B_XJeiFyyT6_0),.clk(gclk));
	jdff dff_B_V3IDgEqV0_0(.din(w_dff_B_XJeiFyyT6_0),.dout(w_dff_B_V3IDgEqV0_0),.clk(gclk));
	jdff dff_B_EOQdpHEL7_0(.din(w_dff_B_V3IDgEqV0_0),.dout(w_dff_B_EOQdpHEL7_0),.clk(gclk));
	jdff dff_B_lnKr4Z7M8_1(.din(n1722),.dout(w_dff_B_lnKr4Z7M8_1),.clk(gclk));
	jdff dff_B_8ryk7nNh3_1(.din(w_dff_B_lnKr4Z7M8_1),.dout(w_dff_B_8ryk7nNh3_1),.clk(gclk));
	jdff dff_B_xT2rPhOl3_1(.din(w_dff_B_8ryk7nNh3_1),.dout(w_dff_B_xT2rPhOl3_1),.clk(gclk));
	jdff dff_B_cyBPuupf1_1(.din(w_dff_B_xT2rPhOl3_1),.dout(w_dff_B_cyBPuupf1_1),.clk(gclk));
	jdff dff_B_RtfzpUNm3_1(.din(w_dff_B_cyBPuupf1_1),.dout(w_dff_B_RtfzpUNm3_1),.clk(gclk));
	jdff dff_B_5IUnnD3o3_1(.din(w_dff_B_RtfzpUNm3_1),.dout(w_dff_B_5IUnnD3o3_1),.clk(gclk));
	jdff dff_B_cInorMwj2_1(.din(w_dff_B_5IUnnD3o3_1),.dout(w_dff_B_cInorMwj2_1),.clk(gclk));
	jdff dff_B_xnrt3JKO3_1(.din(w_dff_B_cInorMwj2_1),.dout(w_dff_B_xnrt3JKO3_1),.clk(gclk));
	jdff dff_B_566lHE4j0_1(.din(w_dff_B_xnrt3JKO3_1),.dout(w_dff_B_566lHE4j0_1),.clk(gclk));
	jdff dff_B_Rt7hsOhw1_1(.din(w_dff_B_566lHE4j0_1),.dout(w_dff_B_Rt7hsOhw1_1),.clk(gclk));
	jdff dff_B_E0Q23Cbc3_1(.din(w_dff_B_Rt7hsOhw1_1),.dout(w_dff_B_E0Q23Cbc3_1),.clk(gclk));
	jdff dff_B_Te4K5kvL8_0(.din(n1723),.dout(w_dff_B_Te4K5kvL8_0),.clk(gclk));
	jdff dff_B_HrG0XZDw7_0(.din(w_dff_B_Te4K5kvL8_0),.dout(w_dff_B_HrG0XZDw7_0),.clk(gclk));
	jdff dff_B_5V2AectB7_0(.din(w_dff_B_HrG0XZDw7_0),.dout(w_dff_B_5V2AectB7_0),.clk(gclk));
	jdff dff_B_vyjlDjqI7_0(.din(w_dff_B_5V2AectB7_0),.dout(w_dff_B_vyjlDjqI7_0),.clk(gclk));
	jdff dff_B_37Ud5FH85_0(.din(w_dff_B_vyjlDjqI7_0),.dout(w_dff_B_37Ud5FH85_0),.clk(gclk));
	jdff dff_B_2VjCm8n39_0(.din(w_dff_B_37Ud5FH85_0),.dout(w_dff_B_2VjCm8n39_0),.clk(gclk));
	jdff dff_B_Xsyp27mk8_0(.din(w_dff_B_2VjCm8n39_0),.dout(w_dff_B_Xsyp27mk8_0),.clk(gclk));
	jdff dff_B_9EHMQM611_0(.din(w_dff_B_Xsyp27mk8_0),.dout(w_dff_B_9EHMQM611_0),.clk(gclk));
	jdff dff_B_JgvJPJc61_0(.din(w_dff_B_9EHMQM611_0),.dout(w_dff_B_JgvJPJc61_0),.clk(gclk));
	jdff dff_B_UVLAc0EO0_1(.din(n1674),.dout(w_dff_B_UVLAc0EO0_1),.clk(gclk));
	jdff dff_B_ldjYnZOI1_1(.din(w_dff_B_UVLAc0EO0_1),.dout(w_dff_B_ldjYnZOI1_1),.clk(gclk));
	jdff dff_B_8qoqtQM48_1(.din(w_dff_B_ldjYnZOI1_1),.dout(w_dff_B_8qoqtQM48_1),.clk(gclk));
	jdff dff_B_a3dab27L0_1(.din(w_dff_B_8qoqtQM48_1),.dout(w_dff_B_a3dab27L0_1),.clk(gclk));
	jdff dff_B_zJk2ODOZ0_1(.din(w_dff_B_a3dab27L0_1),.dout(w_dff_B_zJk2ODOZ0_1),.clk(gclk));
	jdff dff_B_gh0oauVX4_1(.din(w_dff_B_zJk2ODOZ0_1),.dout(w_dff_B_gh0oauVX4_1),.clk(gclk));
	jdff dff_B_Zy8hjRZX6_1(.din(w_dff_B_gh0oauVX4_1),.dout(w_dff_B_Zy8hjRZX6_1),.clk(gclk));
	jdff dff_B_yrkT1iFw0_1(.din(w_dff_B_Zy8hjRZX6_1),.dout(w_dff_B_yrkT1iFw0_1),.clk(gclk));
	jdff dff_B_recaVOal6_1(.din(w_dff_B_yrkT1iFw0_1),.dout(w_dff_B_recaVOal6_1),.clk(gclk));
	jdff dff_B_mdApH64o0_1(.din(w_dff_B_recaVOal6_1),.dout(w_dff_B_mdApH64o0_1),.clk(gclk));
	jdff dff_B_ZACUQHss7_0(.din(n1675),.dout(w_dff_B_ZACUQHss7_0),.clk(gclk));
	jdff dff_B_b66iRCz56_0(.din(w_dff_B_ZACUQHss7_0),.dout(w_dff_B_b66iRCz56_0),.clk(gclk));
	jdff dff_B_C0krQAGI3_0(.din(w_dff_B_b66iRCz56_0),.dout(w_dff_B_C0krQAGI3_0),.clk(gclk));
	jdff dff_B_lZH28Lpf5_0(.din(w_dff_B_C0krQAGI3_0),.dout(w_dff_B_lZH28Lpf5_0),.clk(gclk));
	jdff dff_B_0PpXJGId1_0(.din(w_dff_B_lZH28Lpf5_0),.dout(w_dff_B_0PpXJGId1_0),.clk(gclk));
	jdff dff_B_I3gLJUfE5_0(.din(w_dff_B_0PpXJGId1_0),.dout(w_dff_B_I3gLJUfE5_0),.clk(gclk));
	jdff dff_B_lJpb3XBs9_0(.din(w_dff_B_I3gLJUfE5_0),.dout(w_dff_B_lJpb3XBs9_0),.clk(gclk));
	jdff dff_B_L0Rmnoh95_0(.din(w_dff_B_lJpb3XBs9_0),.dout(w_dff_B_L0Rmnoh95_0),.clk(gclk));
	jdff dff_B_NtB9GY9u5_1(.din(n1619),.dout(w_dff_B_NtB9GY9u5_1),.clk(gclk));
	jdff dff_B_kc2SXV4C9_1(.din(w_dff_B_NtB9GY9u5_1),.dout(w_dff_B_kc2SXV4C9_1),.clk(gclk));
	jdff dff_B_lIn9U0oC5_1(.din(w_dff_B_kc2SXV4C9_1),.dout(w_dff_B_lIn9U0oC5_1),.clk(gclk));
	jdff dff_B_vMqNVLf12_1(.din(w_dff_B_lIn9U0oC5_1),.dout(w_dff_B_vMqNVLf12_1),.clk(gclk));
	jdff dff_B_eK3ZCjBO5_1(.din(w_dff_B_vMqNVLf12_1),.dout(w_dff_B_eK3ZCjBO5_1),.clk(gclk));
	jdff dff_B_ZLlHNbcU6_1(.din(w_dff_B_eK3ZCjBO5_1),.dout(w_dff_B_ZLlHNbcU6_1),.clk(gclk));
	jdff dff_B_4HoTxXe18_1(.din(w_dff_B_ZLlHNbcU6_1),.dout(w_dff_B_4HoTxXe18_1),.clk(gclk));
	jdff dff_B_vK72Semg3_1(.din(w_dff_B_4HoTxXe18_1),.dout(w_dff_B_vK72Semg3_1),.clk(gclk));
	jdff dff_B_hSZeGp3d4_1(.din(w_dff_B_vK72Semg3_1),.dout(w_dff_B_hSZeGp3d4_1),.clk(gclk));
	jdff dff_B_mlg2U20o0_1(.din(w_dff_B_hSZeGp3d4_1),.dout(w_dff_B_mlg2U20o0_1),.clk(gclk));
	jdff dff_B_lK74pQE89_0(.din(n1620),.dout(w_dff_B_lK74pQE89_0),.clk(gclk));
	jdff dff_B_M2oIsJN86_0(.din(w_dff_B_lK74pQE89_0),.dout(w_dff_B_M2oIsJN86_0),.clk(gclk));
	jdff dff_B_qero6xuu1_0(.din(w_dff_B_M2oIsJN86_0),.dout(w_dff_B_qero6xuu1_0),.clk(gclk));
	jdff dff_B_9ZpKI2PX1_0(.din(w_dff_B_qero6xuu1_0),.dout(w_dff_B_9ZpKI2PX1_0),.clk(gclk));
	jdff dff_B_nH3r2rMY5_0(.din(w_dff_B_9ZpKI2PX1_0),.dout(w_dff_B_nH3r2rMY5_0),.clk(gclk));
	jdff dff_B_eMl8xzca9_0(.din(w_dff_B_nH3r2rMY5_0),.dout(w_dff_B_eMl8xzca9_0),.clk(gclk));
	jdff dff_B_C1LZVcf42_0(.din(w_dff_B_eMl8xzca9_0),.dout(w_dff_B_C1LZVcf42_0),.clk(gclk));
	jdff dff_B_KPH1H2a54_0(.din(w_dff_B_C1LZVcf42_0),.dout(w_dff_B_KPH1H2a54_0),.clk(gclk));
	jdff dff_B_SkgusjyV0_1(.din(n1557),.dout(w_dff_B_SkgusjyV0_1),.clk(gclk));
	jdff dff_B_xg0A5I4d9_1(.din(w_dff_B_SkgusjyV0_1),.dout(w_dff_B_xg0A5I4d9_1),.clk(gclk));
	jdff dff_B_5i3qlVWW0_1(.din(w_dff_B_xg0A5I4d9_1),.dout(w_dff_B_5i3qlVWW0_1),.clk(gclk));
	jdff dff_B_B4WHnUco5_1(.din(w_dff_B_5i3qlVWW0_1),.dout(w_dff_B_B4WHnUco5_1),.clk(gclk));
	jdff dff_B_ealkyqLW8_1(.din(w_dff_B_B4WHnUco5_1),.dout(w_dff_B_ealkyqLW8_1),.clk(gclk));
	jdff dff_B_RwCo48J74_1(.din(w_dff_B_ealkyqLW8_1),.dout(w_dff_B_RwCo48J74_1),.clk(gclk));
	jdff dff_B_Gby1XeE97_1(.din(w_dff_B_RwCo48J74_1),.dout(w_dff_B_Gby1XeE97_1),.clk(gclk));
	jdff dff_B_ykjfpplL7_1(.din(w_dff_B_Gby1XeE97_1),.dout(w_dff_B_ykjfpplL7_1),.clk(gclk));
	jdff dff_B_PRkjS5AF3_0(.din(n1558),.dout(w_dff_B_PRkjS5AF3_0),.clk(gclk));
	jdff dff_B_zJBKnvHv2_0(.din(w_dff_B_PRkjS5AF3_0),.dout(w_dff_B_zJBKnvHv2_0),.clk(gclk));
	jdff dff_B_ORoFsjNZ9_0(.din(w_dff_B_zJBKnvHv2_0),.dout(w_dff_B_ORoFsjNZ9_0),.clk(gclk));
	jdff dff_B_dN8MtqrG4_0(.din(w_dff_B_ORoFsjNZ9_0),.dout(w_dff_B_dN8MtqrG4_0),.clk(gclk));
	jdff dff_B_mMBcqcDb9_0(.din(w_dff_B_dN8MtqrG4_0),.dout(w_dff_B_mMBcqcDb9_0),.clk(gclk));
	jdff dff_B_GiR5nEIQ5_0(.din(w_dff_B_mMBcqcDb9_0),.dout(w_dff_B_GiR5nEIQ5_0),.clk(gclk));
	jdff dff_B_nptbMNFz7_1(.din(n1488),.dout(w_dff_B_nptbMNFz7_1),.clk(gclk));
	jdff dff_B_ybqZzHbw3_1(.din(w_dff_B_nptbMNFz7_1),.dout(w_dff_B_ybqZzHbw3_1),.clk(gclk));
	jdff dff_B_lyZevIjg9_1(.din(w_dff_B_ybqZzHbw3_1),.dout(w_dff_B_lyZevIjg9_1),.clk(gclk));
	jdff dff_B_0dddYj4P1_1(.din(w_dff_B_lyZevIjg9_1),.dout(w_dff_B_0dddYj4P1_1),.clk(gclk));
	jdff dff_B_vvQWjoHL8_1(.din(w_dff_B_0dddYj4P1_1),.dout(w_dff_B_vvQWjoHL8_1),.clk(gclk));
	jdff dff_B_FY27eXD76_1(.din(w_dff_B_vvQWjoHL8_1),.dout(w_dff_B_FY27eXD76_1),.clk(gclk));
	jdff dff_B_nLY9nNaa0_1(.din(w_dff_B_FY27eXD76_1),.dout(w_dff_B_nLY9nNaa0_1),.clk(gclk));
	jdff dff_B_4sthuPwJ9_0(.din(n1489),.dout(w_dff_B_4sthuPwJ9_0),.clk(gclk));
	jdff dff_B_00MQZg730_0(.din(w_dff_B_4sthuPwJ9_0),.dout(w_dff_B_00MQZg730_0),.clk(gclk));
	jdff dff_B_RFCXNyKI4_0(.din(w_dff_B_00MQZg730_0),.dout(w_dff_B_RFCXNyKI4_0),.clk(gclk));
	jdff dff_B_ur5vXtRu1_0(.din(w_dff_B_RFCXNyKI4_0),.dout(w_dff_B_ur5vXtRu1_0),.clk(gclk));
	jdff dff_B_6uiefIB11_0(.din(w_dff_B_ur5vXtRu1_0),.dout(w_dff_B_6uiefIB11_0),.clk(gclk));
	jdff dff_B_I9SQWbCD5_1(.din(n1412),.dout(w_dff_B_I9SQWbCD5_1),.clk(gclk));
	jdff dff_B_71iVHwuC6_1(.din(w_dff_B_I9SQWbCD5_1),.dout(w_dff_B_71iVHwuC6_1),.clk(gclk));
	jdff dff_B_SUufHxY01_1(.din(w_dff_B_71iVHwuC6_1),.dout(w_dff_B_SUufHxY01_1),.clk(gclk));
	jdff dff_B_tkTdiyXq4_1(.din(w_dff_B_SUufHxY01_1),.dout(w_dff_B_tkTdiyXq4_1),.clk(gclk));
	jdff dff_B_1GNZutHk9_1(.din(w_dff_B_tkTdiyXq4_1),.dout(w_dff_B_1GNZutHk9_1),.clk(gclk));
	jdff dff_B_lqat5rQz4_1(.din(w_dff_B_1GNZutHk9_1),.dout(w_dff_B_lqat5rQz4_1),.clk(gclk));
	jdff dff_B_TqqQ4Yxt6_0(.din(n1413),.dout(w_dff_B_TqqQ4Yxt6_0),.clk(gclk));
	jdff dff_B_JkGMiJWi8_0(.din(w_dff_B_TqqQ4Yxt6_0),.dout(w_dff_B_JkGMiJWi8_0),.clk(gclk));
	jdff dff_B_3E5T5ux09_0(.din(w_dff_B_JkGMiJWi8_0),.dout(w_dff_B_3E5T5ux09_0),.clk(gclk));
	jdff dff_B_FsUF8c9E3_0(.din(w_dff_B_3E5T5ux09_0),.dout(w_dff_B_FsUF8c9E3_0),.clk(gclk));
	jdff dff_B_NR9urmj73_1(.din(n1330),.dout(w_dff_B_NR9urmj73_1),.clk(gclk));
	jdff dff_B_vpyJeysS8_1(.din(w_dff_B_NR9urmj73_1),.dout(w_dff_B_vpyJeysS8_1),.clk(gclk));
	jdff dff_B_AURzPvBv7_1(.din(w_dff_B_vpyJeysS8_1),.dout(w_dff_B_AURzPvBv7_1),.clk(gclk));
	jdff dff_B_nG2AdicV6_1(.din(n1242),.dout(w_dff_B_nG2AdicV6_1),.clk(gclk));
	jdff dff_B_avGxlZft2_1(.din(n1145),.dout(w_dff_B_avGxlZft2_1),.clk(gclk));
	jdff dff_A_7UVDgp5P2_1(.dout(w_n1039_0[1]),.din(w_dff_A_7UVDgp5P2_1),.clk(gclk));
	jdff dff_B_wDX4iwEr7_2(.din(n1037),.dout(w_dff_B_wDX4iwEr7_2),.clk(gclk));
	jdff dff_B_39iS0oOH0_1(.din(n935),.dout(w_dff_B_39iS0oOH0_1),.clk(gclk));
	jdff dff_B_Vw5ca9Im3_1(.din(n832),.dout(w_dff_B_Vw5ca9Im3_1),.clk(gclk));
	jdff dff_B_2un0XYhY5_1(.din(n732),.dout(w_dff_B_2un0XYhY5_1),.clk(gclk));
	jdff dff_B_PH0q2cYe9_1(.din(n639),.dout(w_dff_B_PH0q2cYe9_1),.clk(gclk));
	jdff dff_B_oci1c3qe0_1(.din(n553),.dout(w_dff_B_oci1c3qe0_1),.clk(gclk));
	jdff dff_B_GX6DC5BQ6_1(.din(n474),.dout(w_dff_B_GX6DC5BQ6_1),.clk(gclk));
	jdff dff_B_APQpbtXG4_1(.din(n402),.dout(w_dff_B_APQpbtXG4_1),.clk(gclk));
	jdff dff_B_mzf3UAuW1_1(.din(n338),.dout(w_dff_B_mzf3UAuW1_1),.clk(gclk));
	jdff dff_B_44uZDAnU6_1(.din(n280),.dout(w_dff_B_44uZDAnU6_1),.clk(gclk));
	jdff dff_B_JW3HweTE7_1(.din(n229),.dout(w_dff_B_JW3HweTE7_1),.clk(gclk));
	jdff dff_B_rPUbm3kx1_1(.din(n186),.dout(w_dff_B_rPUbm3kx1_1),.clk(gclk));
	jdff dff_B_Qkzi8O9h3_1(.din(n148),.dout(w_dff_B_Qkzi8O9h3_1),.clk(gclk));
	jdff dff_B_pS4HvURR3_1(.din(n113),.dout(w_dff_B_pS4HvURR3_1),.clk(gclk));
	jdff dff_B_hckTMUBH6_1(.din(n91),.dout(w_dff_B_hckTMUBH6_1),.clk(gclk));
	jdff dff_B_MoKKPG2t4_0(.din(n86),.dout(w_dff_B_MoKKPG2t4_0),.clk(gclk));
	jdff dff_A_DmL1QnrY4_0(.dout(w_n70_0[0]),.din(w_dff_A_DmL1QnrY4_0),.clk(gclk));
	jdff dff_A_er5FX7J50_0(.dout(w_n69_0[0]),.din(w_dff_A_er5FX7J50_0),.clk(gclk));
	jdff dff_A_bTCAl6WQ9_1(.dout(w_dff_A_0ScrAvYA0_0),.din(w_dff_A_bTCAl6WQ9_1),.clk(gclk));
	jdff dff_A_0ScrAvYA0_0(.dout(w_dff_A_qLQNHc772_0),.din(w_dff_A_0ScrAvYA0_0),.clk(gclk));
	jdff dff_A_qLQNHc772_0(.dout(w_dff_A_sQAbRgXs7_0),.din(w_dff_A_qLQNHc772_0),.clk(gclk));
	jdff dff_A_sQAbRgXs7_0(.dout(w_dff_A_vSrC9zRj6_0),.din(w_dff_A_sQAbRgXs7_0),.clk(gclk));
	jdff dff_A_vSrC9zRj6_0(.dout(w_dff_A_TpQrlgLG0_0),.din(w_dff_A_vSrC9zRj6_0),.clk(gclk));
	jdff dff_A_TpQrlgLG0_0(.dout(w_dff_A_gMDywc4O0_0),.din(w_dff_A_TpQrlgLG0_0),.clk(gclk));
	jdff dff_A_gMDywc4O0_0(.dout(w_dff_A_tBK1z3xF2_0),.din(w_dff_A_gMDywc4O0_0),.clk(gclk));
	jdff dff_A_tBK1z3xF2_0(.dout(w_dff_A_uUoxld6q6_0),.din(w_dff_A_tBK1z3xF2_0),.clk(gclk));
	jdff dff_A_uUoxld6q6_0(.dout(w_dff_A_TSALyH9y1_0),.din(w_dff_A_uUoxld6q6_0),.clk(gclk));
	jdff dff_A_TSALyH9y1_0(.dout(w_dff_A_8ps0W6gc6_0),.din(w_dff_A_TSALyH9y1_0),.clk(gclk));
	jdff dff_A_8ps0W6gc6_0(.dout(w_dff_A_SfDcYrZF8_0),.din(w_dff_A_8ps0W6gc6_0),.clk(gclk));
	jdff dff_A_SfDcYrZF8_0(.dout(w_dff_A_r7UZrAKR5_0),.din(w_dff_A_SfDcYrZF8_0),.clk(gclk));
	jdff dff_A_r7UZrAKR5_0(.dout(w_dff_A_5wePWLCf3_0),.din(w_dff_A_r7UZrAKR5_0),.clk(gclk));
	jdff dff_A_5wePWLCf3_0(.dout(w_dff_A_c6DtyH4Z5_0),.din(w_dff_A_5wePWLCf3_0),.clk(gclk));
	jdff dff_A_c6DtyH4Z5_0(.dout(w_dff_A_yUtL0ibs1_0),.din(w_dff_A_c6DtyH4Z5_0),.clk(gclk));
	jdff dff_A_yUtL0ibs1_0(.dout(w_dff_A_w9w5rUgd2_0),.din(w_dff_A_yUtL0ibs1_0),.clk(gclk));
	jdff dff_A_w9w5rUgd2_0(.dout(w_dff_A_k6MJjzzb4_0),.din(w_dff_A_w9w5rUgd2_0),.clk(gclk));
	jdff dff_A_k6MJjzzb4_0(.dout(w_dff_A_oFhV9Yys2_0),.din(w_dff_A_k6MJjzzb4_0),.clk(gclk));
	jdff dff_A_oFhV9Yys2_0(.dout(w_dff_A_JySU2AdA9_0),.din(w_dff_A_oFhV9Yys2_0),.clk(gclk));
	jdff dff_A_JySU2AdA9_0(.dout(w_dff_A_KL1R5lLa0_0),.din(w_dff_A_JySU2AdA9_0),.clk(gclk));
	jdff dff_A_KL1R5lLa0_0(.dout(w_dff_A_QlsXtofC7_0),.din(w_dff_A_KL1R5lLa0_0),.clk(gclk));
	jdff dff_A_QlsXtofC7_0(.dout(w_dff_A_Ml9p01M16_0),.din(w_dff_A_QlsXtofC7_0),.clk(gclk));
	jdff dff_A_Ml9p01M16_0(.dout(w_dff_A_hgOBoV5l6_0),.din(w_dff_A_Ml9p01M16_0),.clk(gclk));
	jdff dff_A_hgOBoV5l6_0(.dout(w_dff_A_wZoIVWxZ6_0),.din(w_dff_A_hgOBoV5l6_0),.clk(gclk));
	jdff dff_A_wZoIVWxZ6_0(.dout(w_dff_A_Hus5icBz9_0),.din(w_dff_A_wZoIVWxZ6_0),.clk(gclk));
	jdff dff_A_Hus5icBz9_0(.dout(w_dff_A_b67jr6Eg0_0),.din(w_dff_A_Hus5icBz9_0),.clk(gclk));
	jdff dff_A_b67jr6Eg0_0(.dout(w_dff_A_ykMKu8d73_0),.din(w_dff_A_b67jr6Eg0_0),.clk(gclk));
	jdff dff_A_ykMKu8d73_0(.dout(w_dff_A_V9d7Aimv6_0),.din(w_dff_A_ykMKu8d73_0),.clk(gclk));
	jdff dff_A_V9d7Aimv6_0(.dout(w_dff_A_7JUV1yZB5_0),.din(w_dff_A_V9d7Aimv6_0),.clk(gclk));
	jdff dff_A_7JUV1yZB5_0(.dout(w_dff_A_LULJGEXV8_0),.din(w_dff_A_7JUV1yZB5_0),.clk(gclk));
	jdff dff_A_LULJGEXV8_0(.dout(w_dff_A_uLmT33eu7_0),.din(w_dff_A_LULJGEXV8_0),.clk(gclk));
	jdff dff_A_uLmT33eu7_0(.dout(w_dff_A_CDSpkiVt9_0),.din(w_dff_A_uLmT33eu7_0),.clk(gclk));
	jdff dff_A_CDSpkiVt9_0(.dout(w_dff_A_czkmhjny3_0),.din(w_dff_A_CDSpkiVt9_0),.clk(gclk));
	jdff dff_A_czkmhjny3_0(.dout(w_dff_A_k853RhGH4_0),.din(w_dff_A_czkmhjny3_0),.clk(gclk));
	jdff dff_A_k853RhGH4_0(.dout(w_dff_A_aj8YeYcW4_0),.din(w_dff_A_k853RhGH4_0),.clk(gclk));
	jdff dff_A_aj8YeYcW4_0(.dout(w_dff_A_Nfl5jsIK7_0),.din(w_dff_A_aj8YeYcW4_0),.clk(gclk));
	jdff dff_A_Nfl5jsIK7_0(.dout(w_dff_A_9TjwUSOj3_0),.din(w_dff_A_Nfl5jsIK7_0),.clk(gclk));
	jdff dff_A_9TjwUSOj3_0(.dout(w_dff_A_WJ4WcMJ96_0),.din(w_dff_A_9TjwUSOj3_0),.clk(gclk));
	jdff dff_A_WJ4WcMJ96_0(.dout(w_dff_A_eAcLipFN6_0),.din(w_dff_A_WJ4WcMJ96_0),.clk(gclk));
	jdff dff_A_eAcLipFN6_0(.dout(w_dff_A_CjbjKJoK4_0),.din(w_dff_A_eAcLipFN6_0),.clk(gclk));
	jdff dff_A_CjbjKJoK4_0(.dout(w_dff_A_xsCKGOOr4_0),.din(w_dff_A_CjbjKJoK4_0),.clk(gclk));
	jdff dff_A_xsCKGOOr4_0(.dout(w_dff_A_kfiwen4i4_0),.din(w_dff_A_xsCKGOOr4_0),.clk(gclk));
	jdff dff_A_kfiwen4i4_0(.dout(w_dff_A_EhPrHA807_0),.din(w_dff_A_kfiwen4i4_0),.clk(gclk));
	jdff dff_A_EhPrHA807_0(.dout(w_dff_A_PStkDCsD2_0),.din(w_dff_A_EhPrHA807_0),.clk(gclk));
	jdff dff_A_PStkDCsD2_0(.dout(w_dff_A_PqZ9lHp65_0),.din(w_dff_A_PStkDCsD2_0),.clk(gclk));
	jdff dff_A_PqZ9lHp65_0(.dout(w_dff_A_N5TV2sMd6_0),.din(w_dff_A_PqZ9lHp65_0),.clk(gclk));
	jdff dff_A_N5TV2sMd6_0(.dout(w_dff_A_1HmaeqVb3_0),.din(w_dff_A_N5TV2sMd6_0),.clk(gclk));
	jdff dff_A_1HmaeqVb3_0(.dout(w_dff_A_yHb2qhDd5_0),.din(w_dff_A_1HmaeqVb3_0),.clk(gclk));
	jdff dff_A_yHb2qhDd5_0(.dout(w_dff_A_SRkecX2R9_0),.din(w_dff_A_yHb2qhDd5_0),.clk(gclk));
	jdff dff_A_SRkecX2R9_0(.dout(w_dff_A_TMtIDAje4_0),.din(w_dff_A_SRkecX2R9_0),.clk(gclk));
	jdff dff_A_TMtIDAje4_0(.dout(w_dff_A_hsT0ClWq5_0),.din(w_dff_A_TMtIDAje4_0),.clk(gclk));
	jdff dff_A_hsT0ClWq5_0(.dout(w_dff_A_jvqCnlvm2_0),.din(w_dff_A_hsT0ClWq5_0),.clk(gclk));
	jdff dff_A_jvqCnlvm2_0(.dout(w_dff_A_KLP8Ccrj8_0),.din(w_dff_A_jvqCnlvm2_0),.clk(gclk));
	jdff dff_A_KLP8Ccrj8_0(.dout(w_dff_A_HMvn4lKJ5_0),.din(w_dff_A_KLP8Ccrj8_0),.clk(gclk));
	jdff dff_A_HMvn4lKJ5_0(.dout(w_dff_A_g1u098Kg4_0),.din(w_dff_A_HMvn4lKJ5_0),.clk(gclk));
	jdff dff_A_g1u098Kg4_0(.dout(w_dff_A_qD6Vc4tY9_0),.din(w_dff_A_g1u098Kg4_0),.clk(gclk));
	jdff dff_A_qD6Vc4tY9_0(.dout(w_dff_A_nwd66FEe1_0),.din(w_dff_A_qD6Vc4tY9_0),.clk(gclk));
	jdff dff_A_nwd66FEe1_0(.dout(w_dff_A_djA9kIsB9_0),.din(w_dff_A_nwd66FEe1_0),.clk(gclk));
	jdff dff_A_djA9kIsB9_0(.dout(w_dff_A_cVpNKl5A7_0),.din(w_dff_A_djA9kIsB9_0),.clk(gclk));
	jdff dff_A_cVpNKl5A7_0(.dout(w_dff_A_JccXoHeQ7_0),.din(w_dff_A_cVpNKl5A7_0),.clk(gclk));
	jdff dff_A_JccXoHeQ7_0(.dout(w_dff_A_UdverVv39_0),.din(w_dff_A_JccXoHeQ7_0),.clk(gclk));
	jdff dff_A_UdverVv39_0(.dout(w_dff_A_d1Vwirj30_0),.din(w_dff_A_UdverVv39_0),.clk(gclk));
	jdff dff_A_d1Vwirj30_0(.dout(w_dff_A_3DOedldN8_0),.din(w_dff_A_d1Vwirj30_0),.clk(gclk));
	jdff dff_A_3DOedldN8_0(.dout(w_dff_A_aVw6sbrF0_0),.din(w_dff_A_3DOedldN8_0),.clk(gclk));
	jdff dff_A_aVw6sbrF0_0(.dout(w_dff_A_7PPz50Jf7_0),.din(w_dff_A_aVw6sbrF0_0),.clk(gclk));
	jdff dff_A_7PPz50Jf7_0(.dout(w_dff_A_bjUMuoak4_0),.din(w_dff_A_7PPz50Jf7_0),.clk(gclk));
	jdff dff_A_bjUMuoak4_0(.dout(w_dff_A_5CgO0BtO3_0),.din(w_dff_A_bjUMuoak4_0),.clk(gclk));
	jdff dff_A_5CgO0BtO3_0(.dout(w_dff_A_4BrFiUsN2_0),.din(w_dff_A_5CgO0BtO3_0),.clk(gclk));
	jdff dff_A_4BrFiUsN2_0(.dout(w_dff_A_YHZsrDRc7_0),.din(w_dff_A_4BrFiUsN2_0),.clk(gclk));
	jdff dff_A_YHZsrDRc7_0(.dout(w_dff_A_CFwdSuc96_0),.din(w_dff_A_YHZsrDRc7_0),.clk(gclk));
	jdff dff_A_CFwdSuc96_0(.dout(w_dff_A_mKQsCMmW1_0),.din(w_dff_A_CFwdSuc96_0),.clk(gclk));
	jdff dff_A_mKQsCMmW1_0(.dout(w_dff_A_CaANVt3b2_0),.din(w_dff_A_mKQsCMmW1_0),.clk(gclk));
	jdff dff_A_CaANVt3b2_0(.dout(w_dff_A_i7WgIhzW9_0),.din(w_dff_A_CaANVt3b2_0),.clk(gclk));
	jdff dff_A_i7WgIhzW9_0(.dout(w_dff_A_Ylhs6zuk8_0),.din(w_dff_A_i7WgIhzW9_0),.clk(gclk));
	jdff dff_A_Ylhs6zuk8_0(.dout(G545gat),.din(w_dff_A_Ylhs6zuk8_0),.clk(gclk));
	jdff dff_A_PCFOBIdG2_2(.dout(w_dff_A_2Mzr1ECC3_0),.din(w_dff_A_PCFOBIdG2_2),.clk(gclk));
	jdff dff_A_2Mzr1ECC3_0(.dout(w_dff_A_6QKawOoD4_0),.din(w_dff_A_2Mzr1ECC3_0),.clk(gclk));
	jdff dff_A_6QKawOoD4_0(.dout(w_dff_A_qtsaskvR9_0),.din(w_dff_A_6QKawOoD4_0),.clk(gclk));
	jdff dff_A_qtsaskvR9_0(.dout(w_dff_A_Sfvt9r7P4_0),.din(w_dff_A_qtsaskvR9_0),.clk(gclk));
	jdff dff_A_Sfvt9r7P4_0(.dout(w_dff_A_q7zQL3ts8_0),.din(w_dff_A_Sfvt9r7P4_0),.clk(gclk));
	jdff dff_A_q7zQL3ts8_0(.dout(w_dff_A_fIX6F0zj0_0),.din(w_dff_A_q7zQL3ts8_0),.clk(gclk));
	jdff dff_A_fIX6F0zj0_0(.dout(w_dff_A_vYgo1J5r7_0),.din(w_dff_A_fIX6F0zj0_0),.clk(gclk));
	jdff dff_A_vYgo1J5r7_0(.dout(w_dff_A_kruFvQBM7_0),.din(w_dff_A_vYgo1J5r7_0),.clk(gclk));
	jdff dff_A_kruFvQBM7_0(.dout(w_dff_A_IV5qeMYJ4_0),.din(w_dff_A_kruFvQBM7_0),.clk(gclk));
	jdff dff_A_IV5qeMYJ4_0(.dout(w_dff_A_HfrdipqK3_0),.din(w_dff_A_IV5qeMYJ4_0),.clk(gclk));
	jdff dff_A_HfrdipqK3_0(.dout(w_dff_A_KzklCMRf5_0),.din(w_dff_A_HfrdipqK3_0),.clk(gclk));
	jdff dff_A_KzklCMRf5_0(.dout(w_dff_A_TOlj5WV82_0),.din(w_dff_A_KzklCMRf5_0),.clk(gclk));
	jdff dff_A_TOlj5WV82_0(.dout(w_dff_A_20sgbXbq4_0),.din(w_dff_A_TOlj5WV82_0),.clk(gclk));
	jdff dff_A_20sgbXbq4_0(.dout(w_dff_A_TcYi2j4C9_0),.din(w_dff_A_20sgbXbq4_0),.clk(gclk));
	jdff dff_A_TcYi2j4C9_0(.dout(w_dff_A_AANIZtXG9_0),.din(w_dff_A_TcYi2j4C9_0),.clk(gclk));
	jdff dff_A_AANIZtXG9_0(.dout(w_dff_A_0MjJmIVK0_0),.din(w_dff_A_AANIZtXG9_0),.clk(gclk));
	jdff dff_A_0MjJmIVK0_0(.dout(w_dff_A_o8qRoWCs1_0),.din(w_dff_A_0MjJmIVK0_0),.clk(gclk));
	jdff dff_A_o8qRoWCs1_0(.dout(w_dff_A_xRSwZSJU0_0),.din(w_dff_A_o8qRoWCs1_0),.clk(gclk));
	jdff dff_A_xRSwZSJU0_0(.dout(w_dff_A_fuC9qxw03_0),.din(w_dff_A_xRSwZSJU0_0),.clk(gclk));
	jdff dff_A_fuC9qxw03_0(.dout(w_dff_A_yOpVah1B5_0),.din(w_dff_A_fuC9qxw03_0),.clk(gclk));
	jdff dff_A_yOpVah1B5_0(.dout(w_dff_A_L9WocArF1_0),.din(w_dff_A_yOpVah1B5_0),.clk(gclk));
	jdff dff_A_L9WocArF1_0(.dout(w_dff_A_40Vxe5di2_0),.din(w_dff_A_L9WocArF1_0),.clk(gclk));
	jdff dff_A_40Vxe5di2_0(.dout(w_dff_A_W9DxnpiI7_0),.din(w_dff_A_40Vxe5di2_0),.clk(gclk));
	jdff dff_A_W9DxnpiI7_0(.dout(w_dff_A_YHCbXd5w3_0),.din(w_dff_A_W9DxnpiI7_0),.clk(gclk));
	jdff dff_A_YHCbXd5w3_0(.dout(w_dff_A_Re9knHc57_0),.din(w_dff_A_YHCbXd5w3_0),.clk(gclk));
	jdff dff_A_Re9knHc57_0(.dout(w_dff_A_XOXyhfpa9_0),.din(w_dff_A_Re9knHc57_0),.clk(gclk));
	jdff dff_A_XOXyhfpa9_0(.dout(w_dff_A_LsnChDDU8_0),.din(w_dff_A_XOXyhfpa9_0),.clk(gclk));
	jdff dff_A_LsnChDDU8_0(.dout(w_dff_A_ZmF08uMv9_0),.din(w_dff_A_LsnChDDU8_0),.clk(gclk));
	jdff dff_A_ZmF08uMv9_0(.dout(w_dff_A_bYxj8sBs4_0),.din(w_dff_A_ZmF08uMv9_0),.clk(gclk));
	jdff dff_A_bYxj8sBs4_0(.dout(w_dff_A_iiqDTF3D9_0),.din(w_dff_A_bYxj8sBs4_0),.clk(gclk));
	jdff dff_A_iiqDTF3D9_0(.dout(w_dff_A_K79vuuDa3_0),.din(w_dff_A_iiqDTF3D9_0),.clk(gclk));
	jdff dff_A_K79vuuDa3_0(.dout(w_dff_A_f7m85JD31_0),.din(w_dff_A_K79vuuDa3_0),.clk(gclk));
	jdff dff_A_f7m85JD31_0(.dout(w_dff_A_BbEZIhoi3_0),.din(w_dff_A_f7m85JD31_0),.clk(gclk));
	jdff dff_A_BbEZIhoi3_0(.dout(w_dff_A_BfSG9JWu2_0),.din(w_dff_A_BbEZIhoi3_0),.clk(gclk));
	jdff dff_A_BfSG9JWu2_0(.dout(w_dff_A_sC9H0qdR7_0),.din(w_dff_A_BfSG9JWu2_0),.clk(gclk));
	jdff dff_A_sC9H0qdR7_0(.dout(w_dff_A_GnSGWHR24_0),.din(w_dff_A_sC9H0qdR7_0),.clk(gclk));
	jdff dff_A_GnSGWHR24_0(.dout(w_dff_A_9uD8Bf8N0_0),.din(w_dff_A_GnSGWHR24_0),.clk(gclk));
	jdff dff_A_9uD8Bf8N0_0(.dout(w_dff_A_z35CjSuA4_0),.din(w_dff_A_9uD8Bf8N0_0),.clk(gclk));
	jdff dff_A_z35CjSuA4_0(.dout(w_dff_A_PBj5hJAw0_0),.din(w_dff_A_z35CjSuA4_0),.clk(gclk));
	jdff dff_A_PBj5hJAw0_0(.dout(w_dff_A_BhJGv6NN6_0),.din(w_dff_A_PBj5hJAw0_0),.clk(gclk));
	jdff dff_A_BhJGv6NN6_0(.dout(w_dff_A_p09tgYgj6_0),.din(w_dff_A_BhJGv6NN6_0),.clk(gclk));
	jdff dff_A_p09tgYgj6_0(.dout(w_dff_A_79XkmjZf6_0),.din(w_dff_A_p09tgYgj6_0),.clk(gclk));
	jdff dff_A_79XkmjZf6_0(.dout(w_dff_A_fInH4XCV8_0),.din(w_dff_A_79XkmjZf6_0),.clk(gclk));
	jdff dff_A_fInH4XCV8_0(.dout(w_dff_A_SHtWT2Ly0_0),.din(w_dff_A_fInH4XCV8_0),.clk(gclk));
	jdff dff_A_SHtWT2Ly0_0(.dout(w_dff_A_KT4lCMgo8_0),.din(w_dff_A_SHtWT2Ly0_0),.clk(gclk));
	jdff dff_A_KT4lCMgo8_0(.dout(w_dff_A_dWzDn9il4_0),.din(w_dff_A_KT4lCMgo8_0),.clk(gclk));
	jdff dff_A_dWzDn9il4_0(.dout(w_dff_A_cUp3s2dx7_0),.din(w_dff_A_dWzDn9il4_0),.clk(gclk));
	jdff dff_A_cUp3s2dx7_0(.dout(w_dff_A_xij6pl4g4_0),.din(w_dff_A_cUp3s2dx7_0),.clk(gclk));
	jdff dff_A_xij6pl4g4_0(.dout(w_dff_A_TqnhkYWe8_0),.din(w_dff_A_xij6pl4g4_0),.clk(gclk));
	jdff dff_A_TqnhkYWe8_0(.dout(w_dff_A_4k5xBdMV0_0),.din(w_dff_A_TqnhkYWe8_0),.clk(gclk));
	jdff dff_A_4k5xBdMV0_0(.dout(w_dff_A_WkaFB5Xi3_0),.din(w_dff_A_4k5xBdMV0_0),.clk(gclk));
	jdff dff_A_WkaFB5Xi3_0(.dout(w_dff_A_aMyXT85o1_0),.din(w_dff_A_WkaFB5Xi3_0),.clk(gclk));
	jdff dff_A_aMyXT85o1_0(.dout(w_dff_A_kEIejvSk1_0),.din(w_dff_A_aMyXT85o1_0),.clk(gclk));
	jdff dff_A_kEIejvSk1_0(.dout(w_dff_A_pmcdxPhG1_0),.din(w_dff_A_kEIejvSk1_0),.clk(gclk));
	jdff dff_A_pmcdxPhG1_0(.dout(w_dff_A_spjh1imy7_0),.din(w_dff_A_pmcdxPhG1_0),.clk(gclk));
	jdff dff_A_spjh1imy7_0(.dout(w_dff_A_5Otg00Ik3_0),.din(w_dff_A_spjh1imy7_0),.clk(gclk));
	jdff dff_A_5Otg00Ik3_0(.dout(w_dff_A_tezjCjUI0_0),.din(w_dff_A_5Otg00Ik3_0),.clk(gclk));
	jdff dff_A_tezjCjUI0_0(.dout(w_dff_A_urczoHXB2_0),.din(w_dff_A_tezjCjUI0_0),.clk(gclk));
	jdff dff_A_urczoHXB2_0(.dout(w_dff_A_MXXMO5ot8_0),.din(w_dff_A_urczoHXB2_0),.clk(gclk));
	jdff dff_A_MXXMO5ot8_0(.dout(w_dff_A_uGgSWvGW4_0),.din(w_dff_A_MXXMO5ot8_0),.clk(gclk));
	jdff dff_A_uGgSWvGW4_0(.dout(w_dff_A_M4EEyhLj5_0),.din(w_dff_A_uGgSWvGW4_0),.clk(gclk));
	jdff dff_A_M4EEyhLj5_0(.dout(w_dff_A_BoXyyHj22_0),.din(w_dff_A_M4EEyhLj5_0),.clk(gclk));
	jdff dff_A_BoXyyHj22_0(.dout(w_dff_A_KXOUefs93_0),.din(w_dff_A_BoXyyHj22_0),.clk(gclk));
	jdff dff_A_KXOUefs93_0(.dout(w_dff_A_9WUW8n335_0),.din(w_dff_A_KXOUefs93_0),.clk(gclk));
	jdff dff_A_9WUW8n335_0(.dout(w_dff_A_A8KvOhOl2_0),.din(w_dff_A_9WUW8n335_0),.clk(gclk));
	jdff dff_A_A8KvOhOl2_0(.dout(w_dff_A_7h32TuHA1_0),.din(w_dff_A_A8KvOhOl2_0),.clk(gclk));
	jdff dff_A_7h32TuHA1_0(.dout(w_dff_A_ZHltzi1X1_0),.din(w_dff_A_7h32TuHA1_0),.clk(gclk));
	jdff dff_A_ZHltzi1X1_0(.dout(w_dff_A_3wjTuG9P9_0),.din(w_dff_A_ZHltzi1X1_0),.clk(gclk));
	jdff dff_A_3wjTuG9P9_0(.dout(w_dff_A_xfIO8r2W7_0),.din(w_dff_A_3wjTuG9P9_0),.clk(gclk));
	jdff dff_A_xfIO8r2W7_0(.dout(w_dff_A_a0upQTJm5_0),.din(w_dff_A_xfIO8r2W7_0),.clk(gclk));
	jdff dff_A_a0upQTJm5_0(.dout(w_dff_A_yRiCeCrV9_0),.din(w_dff_A_a0upQTJm5_0),.clk(gclk));
	jdff dff_A_yRiCeCrV9_0(.dout(G1581gat),.din(w_dff_A_yRiCeCrV9_0),.clk(gclk));
	jdff dff_A_gydU51Oe5_2(.dout(w_dff_A_f0BGSe2f5_0),.din(w_dff_A_gydU51Oe5_2),.clk(gclk));
	jdff dff_A_f0BGSe2f5_0(.dout(w_dff_A_Z82EQlDJ0_0),.din(w_dff_A_f0BGSe2f5_0),.clk(gclk));
	jdff dff_A_Z82EQlDJ0_0(.dout(w_dff_A_8FEFZ3Sz6_0),.din(w_dff_A_Z82EQlDJ0_0),.clk(gclk));
	jdff dff_A_8FEFZ3Sz6_0(.dout(w_dff_A_YKmMqeaU2_0),.din(w_dff_A_8FEFZ3Sz6_0),.clk(gclk));
	jdff dff_A_YKmMqeaU2_0(.dout(w_dff_A_Nlbuindq6_0),.din(w_dff_A_YKmMqeaU2_0),.clk(gclk));
	jdff dff_A_Nlbuindq6_0(.dout(w_dff_A_aooHxRTH7_0),.din(w_dff_A_Nlbuindq6_0),.clk(gclk));
	jdff dff_A_aooHxRTH7_0(.dout(w_dff_A_02m7LUoB2_0),.din(w_dff_A_aooHxRTH7_0),.clk(gclk));
	jdff dff_A_02m7LUoB2_0(.dout(w_dff_A_Ey6ruAB05_0),.din(w_dff_A_02m7LUoB2_0),.clk(gclk));
	jdff dff_A_Ey6ruAB05_0(.dout(w_dff_A_y3NXqFwT3_0),.din(w_dff_A_Ey6ruAB05_0),.clk(gclk));
	jdff dff_A_y3NXqFwT3_0(.dout(w_dff_A_NKMh9XOT2_0),.din(w_dff_A_y3NXqFwT3_0),.clk(gclk));
	jdff dff_A_NKMh9XOT2_0(.dout(w_dff_A_sODMZWVr2_0),.din(w_dff_A_NKMh9XOT2_0),.clk(gclk));
	jdff dff_A_sODMZWVr2_0(.dout(w_dff_A_EmYJyEwV8_0),.din(w_dff_A_sODMZWVr2_0),.clk(gclk));
	jdff dff_A_EmYJyEwV8_0(.dout(w_dff_A_jpwXQkDx7_0),.din(w_dff_A_EmYJyEwV8_0),.clk(gclk));
	jdff dff_A_jpwXQkDx7_0(.dout(w_dff_A_e7PbWgvi1_0),.din(w_dff_A_jpwXQkDx7_0),.clk(gclk));
	jdff dff_A_e7PbWgvi1_0(.dout(w_dff_A_CmrDmMdF6_0),.din(w_dff_A_e7PbWgvi1_0),.clk(gclk));
	jdff dff_A_CmrDmMdF6_0(.dout(w_dff_A_fYsxbyRn4_0),.din(w_dff_A_CmrDmMdF6_0),.clk(gclk));
	jdff dff_A_fYsxbyRn4_0(.dout(w_dff_A_kJxXDTez0_0),.din(w_dff_A_fYsxbyRn4_0),.clk(gclk));
	jdff dff_A_kJxXDTez0_0(.dout(w_dff_A_2msFmwVe4_0),.din(w_dff_A_kJxXDTez0_0),.clk(gclk));
	jdff dff_A_2msFmwVe4_0(.dout(w_dff_A_Y1vpadBU8_0),.din(w_dff_A_2msFmwVe4_0),.clk(gclk));
	jdff dff_A_Y1vpadBU8_0(.dout(w_dff_A_IR9ELOl26_0),.din(w_dff_A_Y1vpadBU8_0),.clk(gclk));
	jdff dff_A_IR9ELOl26_0(.dout(w_dff_A_LbQzRoPG2_0),.din(w_dff_A_IR9ELOl26_0),.clk(gclk));
	jdff dff_A_LbQzRoPG2_0(.dout(w_dff_A_PbrkiFNE5_0),.din(w_dff_A_LbQzRoPG2_0),.clk(gclk));
	jdff dff_A_PbrkiFNE5_0(.dout(w_dff_A_PsTxWtSE7_0),.din(w_dff_A_PbrkiFNE5_0),.clk(gclk));
	jdff dff_A_PsTxWtSE7_0(.dout(w_dff_A_o7jEZkWX4_0),.din(w_dff_A_PsTxWtSE7_0),.clk(gclk));
	jdff dff_A_o7jEZkWX4_0(.dout(w_dff_A_7t3XfWNz9_0),.din(w_dff_A_o7jEZkWX4_0),.clk(gclk));
	jdff dff_A_7t3XfWNz9_0(.dout(w_dff_A_XgoMQO123_0),.din(w_dff_A_7t3XfWNz9_0),.clk(gclk));
	jdff dff_A_XgoMQO123_0(.dout(w_dff_A_wG1z2PhT4_0),.din(w_dff_A_XgoMQO123_0),.clk(gclk));
	jdff dff_A_wG1z2PhT4_0(.dout(w_dff_A_QuhbicoL8_0),.din(w_dff_A_wG1z2PhT4_0),.clk(gclk));
	jdff dff_A_QuhbicoL8_0(.dout(w_dff_A_pYRUjwUH3_0),.din(w_dff_A_QuhbicoL8_0),.clk(gclk));
	jdff dff_A_pYRUjwUH3_0(.dout(w_dff_A_6lbBUaA12_0),.din(w_dff_A_pYRUjwUH3_0),.clk(gclk));
	jdff dff_A_6lbBUaA12_0(.dout(w_dff_A_02XnWht50_0),.din(w_dff_A_6lbBUaA12_0),.clk(gclk));
	jdff dff_A_02XnWht50_0(.dout(w_dff_A_yZOGwDdy5_0),.din(w_dff_A_02XnWht50_0),.clk(gclk));
	jdff dff_A_yZOGwDdy5_0(.dout(w_dff_A_fXIKyH653_0),.din(w_dff_A_yZOGwDdy5_0),.clk(gclk));
	jdff dff_A_fXIKyH653_0(.dout(w_dff_A_cfc6UD1e7_0),.din(w_dff_A_fXIKyH653_0),.clk(gclk));
	jdff dff_A_cfc6UD1e7_0(.dout(w_dff_A_NMSQm9MR7_0),.din(w_dff_A_cfc6UD1e7_0),.clk(gclk));
	jdff dff_A_NMSQm9MR7_0(.dout(w_dff_A_5u7OaqjL0_0),.din(w_dff_A_NMSQm9MR7_0),.clk(gclk));
	jdff dff_A_5u7OaqjL0_0(.dout(w_dff_A_kK3LOHlJ4_0),.din(w_dff_A_5u7OaqjL0_0),.clk(gclk));
	jdff dff_A_kK3LOHlJ4_0(.dout(w_dff_A_4rjhZXYO1_0),.din(w_dff_A_kK3LOHlJ4_0),.clk(gclk));
	jdff dff_A_4rjhZXYO1_0(.dout(w_dff_A_PrmI54Ub1_0),.din(w_dff_A_4rjhZXYO1_0),.clk(gclk));
	jdff dff_A_PrmI54Ub1_0(.dout(w_dff_A_IUVx0WOO6_0),.din(w_dff_A_PrmI54Ub1_0),.clk(gclk));
	jdff dff_A_IUVx0WOO6_0(.dout(w_dff_A_x7acFD1t4_0),.din(w_dff_A_IUVx0WOO6_0),.clk(gclk));
	jdff dff_A_x7acFD1t4_0(.dout(w_dff_A_EXnmhxjQ7_0),.din(w_dff_A_x7acFD1t4_0),.clk(gclk));
	jdff dff_A_EXnmhxjQ7_0(.dout(w_dff_A_SV20HDXb9_0),.din(w_dff_A_EXnmhxjQ7_0),.clk(gclk));
	jdff dff_A_SV20HDXb9_0(.dout(w_dff_A_S1NUcAYo4_0),.din(w_dff_A_SV20HDXb9_0),.clk(gclk));
	jdff dff_A_S1NUcAYo4_0(.dout(w_dff_A_KjQWqlTc9_0),.din(w_dff_A_S1NUcAYo4_0),.clk(gclk));
	jdff dff_A_KjQWqlTc9_0(.dout(w_dff_A_W7rxWAuA6_0),.din(w_dff_A_KjQWqlTc9_0),.clk(gclk));
	jdff dff_A_W7rxWAuA6_0(.dout(w_dff_A_gGrn6bqt5_0),.din(w_dff_A_W7rxWAuA6_0),.clk(gclk));
	jdff dff_A_gGrn6bqt5_0(.dout(w_dff_A_tvdmtwT72_0),.din(w_dff_A_gGrn6bqt5_0),.clk(gclk));
	jdff dff_A_tvdmtwT72_0(.dout(w_dff_A_g3iGdPqK3_0),.din(w_dff_A_tvdmtwT72_0),.clk(gclk));
	jdff dff_A_g3iGdPqK3_0(.dout(w_dff_A_nb6Nw2eq1_0),.din(w_dff_A_g3iGdPqK3_0),.clk(gclk));
	jdff dff_A_nb6Nw2eq1_0(.dout(w_dff_A_KDkDbngu1_0),.din(w_dff_A_nb6Nw2eq1_0),.clk(gclk));
	jdff dff_A_KDkDbngu1_0(.dout(w_dff_A_halcnJiQ9_0),.din(w_dff_A_KDkDbngu1_0),.clk(gclk));
	jdff dff_A_halcnJiQ9_0(.dout(w_dff_A_8uHcXYeR0_0),.din(w_dff_A_halcnJiQ9_0),.clk(gclk));
	jdff dff_A_8uHcXYeR0_0(.dout(w_dff_A_gC3Qiwfd9_0),.din(w_dff_A_8uHcXYeR0_0),.clk(gclk));
	jdff dff_A_gC3Qiwfd9_0(.dout(w_dff_A_o0s4HBiH8_0),.din(w_dff_A_gC3Qiwfd9_0),.clk(gclk));
	jdff dff_A_o0s4HBiH8_0(.dout(w_dff_A_npWGeNy41_0),.din(w_dff_A_o0s4HBiH8_0),.clk(gclk));
	jdff dff_A_npWGeNy41_0(.dout(w_dff_A_7cSNeZNJ3_0),.din(w_dff_A_npWGeNy41_0),.clk(gclk));
	jdff dff_A_7cSNeZNJ3_0(.dout(w_dff_A_MEfw7ESU9_0),.din(w_dff_A_7cSNeZNJ3_0),.clk(gclk));
	jdff dff_A_MEfw7ESU9_0(.dout(w_dff_A_Aj5JIvaH9_0),.din(w_dff_A_MEfw7ESU9_0),.clk(gclk));
	jdff dff_A_Aj5JIvaH9_0(.dout(w_dff_A_DcTs0AJE7_0),.din(w_dff_A_Aj5JIvaH9_0),.clk(gclk));
	jdff dff_A_DcTs0AJE7_0(.dout(w_dff_A_xyrkQMju2_0),.din(w_dff_A_DcTs0AJE7_0),.clk(gclk));
	jdff dff_A_xyrkQMju2_0(.dout(w_dff_A_VhTIUq7m4_0),.din(w_dff_A_xyrkQMju2_0),.clk(gclk));
	jdff dff_A_VhTIUq7m4_0(.dout(w_dff_A_tmLdcmJc5_0),.din(w_dff_A_VhTIUq7m4_0),.clk(gclk));
	jdff dff_A_tmLdcmJc5_0(.dout(w_dff_A_XJUDcSpe1_0),.din(w_dff_A_tmLdcmJc5_0),.clk(gclk));
	jdff dff_A_XJUDcSpe1_0(.dout(w_dff_A_q39y2On41_0),.din(w_dff_A_XJUDcSpe1_0),.clk(gclk));
	jdff dff_A_q39y2On41_0(.dout(w_dff_A_lOleXO5M1_0),.din(w_dff_A_q39y2On41_0),.clk(gclk));
	jdff dff_A_lOleXO5M1_0(.dout(w_dff_A_jGqRSgYq8_0),.din(w_dff_A_lOleXO5M1_0),.clk(gclk));
	jdff dff_A_jGqRSgYq8_0(.dout(w_dff_A_1EyJbabK4_0),.din(w_dff_A_jGqRSgYq8_0),.clk(gclk));
	jdff dff_A_1EyJbabK4_0(.dout(G1901gat),.din(w_dff_A_1EyJbabK4_0),.clk(gclk));
	jdff dff_A_prb6lJFG0_2(.dout(w_dff_A_OxDidKSP6_0),.din(w_dff_A_prb6lJFG0_2),.clk(gclk));
	jdff dff_A_OxDidKSP6_0(.dout(w_dff_A_nhZic5li8_0),.din(w_dff_A_OxDidKSP6_0),.clk(gclk));
	jdff dff_A_nhZic5li8_0(.dout(w_dff_A_qVQCv1YV5_0),.din(w_dff_A_nhZic5li8_0),.clk(gclk));
	jdff dff_A_qVQCv1YV5_0(.dout(w_dff_A_uOX3vY8y9_0),.din(w_dff_A_qVQCv1YV5_0),.clk(gclk));
	jdff dff_A_uOX3vY8y9_0(.dout(w_dff_A_jiOCJq2f3_0),.din(w_dff_A_uOX3vY8y9_0),.clk(gclk));
	jdff dff_A_jiOCJq2f3_0(.dout(w_dff_A_GViBomQK2_0),.din(w_dff_A_jiOCJq2f3_0),.clk(gclk));
	jdff dff_A_GViBomQK2_0(.dout(w_dff_A_BPR3l0ig8_0),.din(w_dff_A_GViBomQK2_0),.clk(gclk));
	jdff dff_A_BPR3l0ig8_0(.dout(w_dff_A_BVTRRFdk0_0),.din(w_dff_A_BPR3l0ig8_0),.clk(gclk));
	jdff dff_A_BVTRRFdk0_0(.dout(w_dff_A_sHcPSkRH4_0),.din(w_dff_A_BVTRRFdk0_0),.clk(gclk));
	jdff dff_A_sHcPSkRH4_0(.dout(w_dff_A_BaoC3HYn5_0),.din(w_dff_A_sHcPSkRH4_0),.clk(gclk));
	jdff dff_A_BaoC3HYn5_0(.dout(w_dff_A_vtT2dp4p0_0),.din(w_dff_A_BaoC3HYn5_0),.clk(gclk));
	jdff dff_A_vtT2dp4p0_0(.dout(w_dff_A_v1QtNPQd3_0),.din(w_dff_A_vtT2dp4p0_0),.clk(gclk));
	jdff dff_A_v1QtNPQd3_0(.dout(w_dff_A_N14FrFCB5_0),.din(w_dff_A_v1QtNPQd3_0),.clk(gclk));
	jdff dff_A_N14FrFCB5_0(.dout(w_dff_A_tDFYfXtJ0_0),.din(w_dff_A_N14FrFCB5_0),.clk(gclk));
	jdff dff_A_tDFYfXtJ0_0(.dout(w_dff_A_NWvUz3em2_0),.din(w_dff_A_tDFYfXtJ0_0),.clk(gclk));
	jdff dff_A_NWvUz3em2_0(.dout(w_dff_A_xgo9767D0_0),.din(w_dff_A_NWvUz3em2_0),.clk(gclk));
	jdff dff_A_xgo9767D0_0(.dout(w_dff_A_1dlcXUkU6_0),.din(w_dff_A_xgo9767D0_0),.clk(gclk));
	jdff dff_A_1dlcXUkU6_0(.dout(w_dff_A_tK44xAL30_0),.din(w_dff_A_1dlcXUkU6_0),.clk(gclk));
	jdff dff_A_tK44xAL30_0(.dout(w_dff_A_XSa6KXDS5_0),.din(w_dff_A_tK44xAL30_0),.clk(gclk));
	jdff dff_A_XSa6KXDS5_0(.dout(w_dff_A_i5QkZB390_0),.din(w_dff_A_XSa6KXDS5_0),.clk(gclk));
	jdff dff_A_i5QkZB390_0(.dout(w_dff_A_KRykysKq3_0),.din(w_dff_A_i5QkZB390_0),.clk(gclk));
	jdff dff_A_KRykysKq3_0(.dout(w_dff_A_dJJBCedG5_0),.din(w_dff_A_KRykysKq3_0),.clk(gclk));
	jdff dff_A_dJJBCedG5_0(.dout(w_dff_A_gKHGj8eP3_0),.din(w_dff_A_dJJBCedG5_0),.clk(gclk));
	jdff dff_A_gKHGj8eP3_0(.dout(w_dff_A_EN3SHpej0_0),.din(w_dff_A_gKHGj8eP3_0),.clk(gclk));
	jdff dff_A_EN3SHpej0_0(.dout(w_dff_A_visgnOOx6_0),.din(w_dff_A_EN3SHpej0_0),.clk(gclk));
	jdff dff_A_visgnOOx6_0(.dout(w_dff_A_BaUCnUCu8_0),.din(w_dff_A_visgnOOx6_0),.clk(gclk));
	jdff dff_A_BaUCnUCu8_0(.dout(w_dff_A_868bPX6R5_0),.din(w_dff_A_BaUCnUCu8_0),.clk(gclk));
	jdff dff_A_868bPX6R5_0(.dout(w_dff_A_djX1Utye9_0),.din(w_dff_A_868bPX6R5_0),.clk(gclk));
	jdff dff_A_djX1Utye9_0(.dout(w_dff_A_L5yEuaN89_0),.din(w_dff_A_djX1Utye9_0),.clk(gclk));
	jdff dff_A_L5yEuaN89_0(.dout(w_dff_A_FtbR5yr94_0),.din(w_dff_A_L5yEuaN89_0),.clk(gclk));
	jdff dff_A_FtbR5yr94_0(.dout(w_dff_A_7OJ4VoAa6_0),.din(w_dff_A_FtbR5yr94_0),.clk(gclk));
	jdff dff_A_7OJ4VoAa6_0(.dout(w_dff_A_fgphuv9K2_0),.din(w_dff_A_7OJ4VoAa6_0),.clk(gclk));
	jdff dff_A_fgphuv9K2_0(.dout(w_dff_A_98YRb6NB4_0),.din(w_dff_A_fgphuv9K2_0),.clk(gclk));
	jdff dff_A_98YRb6NB4_0(.dout(w_dff_A_Nd46zg6l7_0),.din(w_dff_A_98YRb6NB4_0),.clk(gclk));
	jdff dff_A_Nd46zg6l7_0(.dout(w_dff_A_8ZNJjnBP0_0),.din(w_dff_A_Nd46zg6l7_0),.clk(gclk));
	jdff dff_A_8ZNJjnBP0_0(.dout(w_dff_A_smKaSlsP2_0),.din(w_dff_A_8ZNJjnBP0_0),.clk(gclk));
	jdff dff_A_smKaSlsP2_0(.dout(w_dff_A_xGrdbFud0_0),.din(w_dff_A_smKaSlsP2_0),.clk(gclk));
	jdff dff_A_xGrdbFud0_0(.dout(w_dff_A_qInHphzq1_0),.din(w_dff_A_xGrdbFud0_0),.clk(gclk));
	jdff dff_A_qInHphzq1_0(.dout(w_dff_A_O9y1Lb8v6_0),.din(w_dff_A_qInHphzq1_0),.clk(gclk));
	jdff dff_A_O9y1Lb8v6_0(.dout(w_dff_A_VhWduckN3_0),.din(w_dff_A_O9y1Lb8v6_0),.clk(gclk));
	jdff dff_A_VhWduckN3_0(.dout(w_dff_A_xsRKr0yu5_0),.din(w_dff_A_VhWduckN3_0),.clk(gclk));
	jdff dff_A_xsRKr0yu5_0(.dout(w_dff_A_40cJkeo17_0),.din(w_dff_A_xsRKr0yu5_0),.clk(gclk));
	jdff dff_A_40cJkeo17_0(.dout(w_dff_A_18VOsNQB2_0),.din(w_dff_A_40cJkeo17_0),.clk(gclk));
	jdff dff_A_18VOsNQB2_0(.dout(w_dff_A_9sdn0RMT2_0),.din(w_dff_A_18VOsNQB2_0),.clk(gclk));
	jdff dff_A_9sdn0RMT2_0(.dout(w_dff_A_98yKo7043_0),.din(w_dff_A_9sdn0RMT2_0),.clk(gclk));
	jdff dff_A_98yKo7043_0(.dout(w_dff_A_uhu3chIJ6_0),.din(w_dff_A_98yKo7043_0),.clk(gclk));
	jdff dff_A_uhu3chIJ6_0(.dout(w_dff_A_W66ZXEkR4_0),.din(w_dff_A_uhu3chIJ6_0),.clk(gclk));
	jdff dff_A_W66ZXEkR4_0(.dout(w_dff_A_Z4KDpIEW7_0),.din(w_dff_A_W66ZXEkR4_0),.clk(gclk));
	jdff dff_A_Z4KDpIEW7_0(.dout(w_dff_A_RbhZD9fC4_0),.din(w_dff_A_Z4KDpIEW7_0),.clk(gclk));
	jdff dff_A_RbhZD9fC4_0(.dout(w_dff_A_W8eiWEpY2_0),.din(w_dff_A_RbhZD9fC4_0),.clk(gclk));
	jdff dff_A_W8eiWEpY2_0(.dout(w_dff_A_fh2Rwq3V3_0),.din(w_dff_A_W8eiWEpY2_0),.clk(gclk));
	jdff dff_A_fh2Rwq3V3_0(.dout(w_dff_A_dX8P4xxg6_0),.din(w_dff_A_fh2Rwq3V3_0),.clk(gclk));
	jdff dff_A_dX8P4xxg6_0(.dout(w_dff_A_7fRx0Mrl3_0),.din(w_dff_A_dX8P4xxg6_0),.clk(gclk));
	jdff dff_A_7fRx0Mrl3_0(.dout(w_dff_A_auYM8PUv0_0),.din(w_dff_A_7fRx0Mrl3_0),.clk(gclk));
	jdff dff_A_auYM8PUv0_0(.dout(w_dff_A_hLHArS1K8_0),.din(w_dff_A_auYM8PUv0_0),.clk(gclk));
	jdff dff_A_hLHArS1K8_0(.dout(w_dff_A_qWyZckTx6_0),.din(w_dff_A_hLHArS1K8_0),.clk(gclk));
	jdff dff_A_qWyZckTx6_0(.dout(w_dff_A_TXm0458n1_0),.din(w_dff_A_qWyZckTx6_0),.clk(gclk));
	jdff dff_A_TXm0458n1_0(.dout(w_dff_A_o8ZbXhrK7_0),.din(w_dff_A_TXm0458n1_0),.clk(gclk));
	jdff dff_A_o8ZbXhrK7_0(.dout(w_dff_A_ycn3xqJR2_0),.din(w_dff_A_o8ZbXhrK7_0),.clk(gclk));
	jdff dff_A_ycn3xqJR2_0(.dout(w_dff_A_Ljgp1K857_0),.din(w_dff_A_ycn3xqJR2_0),.clk(gclk));
	jdff dff_A_Ljgp1K857_0(.dout(w_dff_A_WVhfadmC6_0),.din(w_dff_A_Ljgp1K857_0),.clk(gclk));
	jdff dff_A_WVhfadmC6_0(.dout(w_dff_A_YMi4KCxM8_0),.din(w_dff_A_WVhfadmC6_0),.clk(gclk));
	jdff dff_A_YMi4KCxM8_0(.dout(w_dff_A_B2GAhc2t0_0),.din(w_dff_A_YMi4KCxM8_0),.clk(gclk));
	jdff dff_A_B2GAhc2t0_0(.dout(w_dff_A_KptnlIbk0_0),.din(w_dff_A_B2GAhc2t0_0),.clk(gclk));
	jdff dff_A_KptnlIbk0_0(.dout(w_dff_A_usnr3rUr2_0),.din(w_dff_A_KptnlIbk0_0),.clk(gclk));
	jdff dff_A_usnr3rUr2_0(.dout(G2223gat),.din(w_dff_A_usnr3rUr2_0),.clk(gclk));
	jdff dff_A_wOXl4S3M1_2(.dout(w_dff_A_7hy5QJns0_0),.din(w_dff_A_wOXl4S3M1_2),.clk(gclk));
	jdff dff_A_7hy5QJns0_0(.dout(w_dff_A_9hqhv14t9_0),.din(w_dff_A_7hy5QJns0_0),.clk(gclk));
	jdff dff_A_9hqhv14t9_0(.dout(w_dff_A_Eg2t6DAC9_0),.din(w_dff_A_9hqhv14t9_0),.clk(gclk));
	jdff dff_A_Eg2t6DAC9_0(.dout(w_dff_A_Ucnyg9uT8_0),.din(w_dff_A_Eg2t6DAC9_0),.clk(gclk));
	jdff dff_A_Ucnyg9uT8_0(.dout(w_dff_A_HFgQc5mW3_0),.din(w_dff_A_Ucnyg9uT8_0),.clk(gclk));
	jdff dff_A_HFgQc5mW3_0(.dout(w_dff_A_m2Fx4NjN1_0),.din(w_dff_A_HFgQc5mW3_0),.clk(gclk));
	jdff dff_A_m2Fx4NjN1_0(.dout(w_dff_A_cNwbseb57_0),.din(w_dff_A_m2Fx4NjN1_0),.clk(gclk));
	jdff dff_A_cNwbseb57_0(.dout(w_dff_A_8434XY279_0),.din(w_dff_A_cNwbseb57_0),.clk(gclk));
	jdff dff_A_8434XY279_0(.dout(w_dff_A_JxH1Zs8H1_0),.din(w_dff_A_8434XY279_0),.clk(gclk));
	jdff dff_A_JxH1Zs8H1_0(.dout(w_dff_A_J77lj9Wa2_0),.din(w_dff_A_JxH1Zs8H1_0),.clk(gclk));
	jdff dff_A_J77lj9Wa2_0(.dout(w_dff_A_TxcUI6uj4_0),.din(w_dff_A_J77lj9Wa2_0),.clk(gclk));
	jdff dff_A_TxcUI6uj4_0(.dout(w_dff_A_EwTEVRUW8_0),.din(w_dff_A_TxcUI6uj4_0),.clk(gclk));
	jdff dff_A_EwTEVRUW8_0(.dout(w_dff_A_0EUdAcGq7_0),.din(w_dff_A_EwTEVRUW8_0),.clk(gclk));
	jdff dff_A_0EUdAcGq7_0(.dout(w_dff_A_trISoiH85_0),.din(w_dff_A_0EUdAcGq7_0),.clk(gclk));
	jdff dff_A_trISoiH85_0(.dout(w_dff_A_GSLkOisb4_0),.din(w_dff_A_trISoiH85_0),.clk(gclk));
	jdff dff_A_GSLkOisb4_0(.dout(w_dff_A_6xvPxCsa1_0),.din(w_dff_A_GSLkOisb4_0),.clk(gclk));
	jdff dff_A_6xvPxCsa1_0(.dout(w_dff_A_1uvFQFdB0_0),.din(w_dff_A_6xvPxCsa1_0),.clk(gclk));
	jdff dff_A_1uvFQFdB0_0(.dout(w_dff_A_bcgkZdub8_0),.din(w_dff_A_1uvFQFdB0_0),.clk(gclk));
	jdff dff_A_bcgkZdub8_0(.dout(w_dff_A_XauOiins2_0),.din(w_dff_A_bcgkZdub8_0),.clk(gclk));
	jdff dff_A_XauOiins2_0(.dout(w_dff_A_vABrxvFW2_0),.din(w_dff_A_XauOiins2_0),.clk(gclk));
	jdff dff_A_vABrxvFW2_0(.dout(w_dff_A_NpsOMvbQ7_0),.din(w_dff_A_vABrxvFW2_0),.clk(gclk));
	jdff dff_A_NpsOMvbQ7_0(.dout(w_dff_A_7ONuRJUz4_0),.din(w_dff_A_NpsOMvbQ7_0),.clk(gclk));
	jdff dff_A_7ONuRJUz4_0(.dout(w_dff_A_qnQvu6wG7_0),.din(w_dff_A_7ONuRJUz4_0),.clk(gclk));
	jdff dff_A_qnQvu6wG7_0(.dout(w_dff_A_yHLzZtqQ6_0),.din(w_dff_A_qnQvu6wG7_0),.clk(gclk));
	jdff dff_A_yHLzZtqQ6_0(.dout(w_dff_A_S3XagoCB4_0),.din(w_dff_A_yHLzZtqQ6_0),.clk(gclk));
	jdff dff_A_S3XagoCB4_0(.dout(w_dff_A_qJZC3b2K1_0),.din(w_dff_A_S3XagoCB4_0),.clk(gclk));
	jdff dff_A_qJZC3b2K1_0(.dout(w_dff_A_h7xJIght0_0),.din(w_dff_A_qJZC3b2K1_0),.clk(gclk));
	jdff dff_A_h7xJIght0_0(.dout(w_dff_A_pA7sS7h18_0),.din(w_dff_A_h7xJIght0_0),.clk(gclk));
	jdff dff_A_pA7sS7h18_0(.dout(w_dff_A_uPneUDtG5_0),.din(w_dff_A_pA7sS7h18_0),.clk(gclk));
	jdff dff_A_uPneUDtG5_0(.dout(w_dff_A_pGczmvaZ8_0),.din(w_dff_A_uPneUDtG5_0),.clk(gclk));
	jdff dff_A_pGczmvaZ8_0(.dout(w_dff_A_mQKarlVz4_0),.din(w_dff_A_pGczmvaZ8_0),.clk(gclk));
	jdff dff_A_mQKarlVz4_0(.dout(w_dff_A_2ghvIAro6_0),.din(w_dff_A_mQKarlVz4_0),.clk(gclk));
	jdff dff_A_2ghvIAro6_0(.dout(w_dff_A_pEinz4bu7_0),.din(w_dff_A_2ghvIAro6_0),.clk(gclk));
	jdff dff_A_pEinz4bu7_0(.dout(w_dff_A_kIk9LCbv3_0),.din(w_dff_A_pEinz4bu7_0),.clk(gclk));
	jdff dff_A_kIk9LCbv3_0(.dout(w_dff_A_UE3MjOxz0_0),.din(w_dff_A_kIk9LCbv3_0),.clk(gclk));
	jdff dff_A_UE3MjOxz0_0(.dout(w_dff_A_zyUsQLb01_0),.din(w_dff_A_UE3MjOxz0_0),.clk(gclk));
	jdff dff_A_zyUsQLb01_0(.dout(w_dff_A_ZInLNyof0_0),.din(w_dff_A_zyUsQLb01_0),.clk(gclk));
	jdff dff_A_ZInLNyof0_0(.dout(w_dff_A_xXkyusC57_0),.din(w_dff_A_ZInLNyof0_0),.clk(gclk));
	jdff dff_A_xXkyusC57_0(.dout(w_dff_A_jCgXjnTd6_0),.din(w_dff_A_xXkyusC57_0),.clk(gclk));
	jdff dff_A_jCgXjnTd6_0(.dout(w_dff_A_Zz3Cu5Ob4_0),.din(w_dff_A_jCgXjnTd6_0),.clk(gclk));
	jdff dff_A_Zz3Cu5Ob4_0(.dout(w_dff_A_hTm1wQGb2_0),.din(w_dff_A_Zz3Cu5Ob4_0),.clk(gclk));
	jdff dff_A_hTm1wQGb2_0(.dout(w_dff_A_3tHjbWCs9_0),.din(w_dff_A_hTm1wQGb2_0),.clk(gclk));
	jdff dff_A_3tHjbWCs9_0(.dout(w_dff_A_SNvfIzRR2_0),.din(w_dff_A_3tHjbWCs9_0),.clk(gclk));
	jdff dff_A_SNvfIzRR2_0(.dout(w_dff_A_FCM4mrq16_0),.din(w_dff_A_SNvfIzRR2_0),.clk(gclk));
	jdff dff_A_FCM4mrq16_0(.dout(w_dff_A_YKJtArdH0_0),.din(w_dff_A_FCM4mrq16_0),.clk(gclk));
	jdff dff_A_YKJtArdH0_0(.dout(w_dff_A_CeUtBCTm7_0),.din(w_dff_A_YKJtArdH0_0),.clk(gclk));
	jdff dff_A_CeUtBCTm7_0(.dout(w_dff_A_8KD9NmQT3_0),.din(w_dff_A_CeUtBCTm7_0),.clk(gclk));
	jdff dff_A_8KD9NmQT3_0(.dout(w_dff_A_Mbfv8Efu0_0),.din(w_dff_A_8KD9NmQT3_0),.clk(gclk));
	jdff dff_A_Mbfv8Efu0_0(.dout(w_dff_A_OjDTsPix5_0),.din(w_dff_A_Mbfv8Efu0_0),.clk(gclk));
	jdff dff_A_OjDTsPix5_0(.dout(w_dff_A_sbFXTfGl4_0),.din(w_dff_A_OjDTsPix5_0),.clk(gclk));
	jdff dff_A_sbFXTfGl4_0(.dout(w_dff_A_kJXpJdIh5_0),.din(w_dff_A_sbFXTfGl4_0),.clk(gclk));
	jdff dff_A_kJXpJdIh5_0(.dout(w_dff_A_7nFt87XP2_0),.din(w_dff_A_kJXpJdIh5_0),.clk(gclk));
	jdff dff_A_7nFt87XP2_0(.dout(w_dff_A_hhzOfGZQ0_0),.din(w_dff_A_7nFt87XP2_0),.clk(gclk));
	jdff dff_A_hhzOfGZQ0_0(.dout(w_dff_A_uQ4sCpKG5_0),.din(w_dff_A_hhzOfGZQ0_0),.clk(gclk));
	jdff dff_A_uQ4sCpKG5_0(.dout(w_dff_A_nnY1DhGg0_0),.din(w_dff_A_uQ4sCpKG5_0),.clk(gclk));
	jdff dff_A_nnY1DhGg0_0(.dout(w_dff_A_40tFfYE27_0),.din(w_dff_A_nnY1DhGg0_0),.clk(gclk));
	jdff dff_A_40tFfYE27_0(.dout(w_dff_A_rLL3qYXL8_0),.din(w_dff_A_40tFfYE27_0),.clk(gclk));
	jdff dff_A_rLL3qYXL8_0(.dout(w_dff_A_y6YoDGeR0_0),.din(w_dff_A_rLL3qYXL8_0),.clk(gclk));
	jdff dff_A_y6YoDGeR0_0(.dout(w_dff_A_Xi7DDEN93_0),.din(w_dff_A_y6YoDGeR0_0),.clk(gclk));
	jdff dff_A_Xi7DDEN93_0(.dout(w_dff_A_FS9LwAhT9_0),.din(w_dff_A_Xi7DDEN93_0),.clk(gclk));
	jdff dff_A_FS9LwAhT9_0(.dout(w_dff_A_DWaR64Ip1_0),.din(w_dff_A_FS9LwAhT9_0),.clk(gclk));
	jdff dff_A_DWaR64Ip1_0(.dout(w_dff_A_ZLjqwxAp1_0),.din(w_dff_A_DWaR64Ip1_0),.clk(gclk));
	jdff dff_A_ZLjqwxAp1_0(.dout(G2548gat),.din(w_dff_A_ZLjqwxAp1_0),.clk(gclk));
	jdff dff_A_SMosFExk3_2(.dout(w_dff_A_2rCC6sEb4_0),.din(w_dff_A_SMosFExk3_2),.clk(gclk));
	jdff dff_A_2rCC6sEb4_0(.dout(w_dff_A_vqOlRl3Q0_0),.din(w_dff_A_2rCC6sEb4_0),.clk(gclk));
	jdff dff_A_vqOlRl3Q0_0(.dout(w_dff_A_UJhNnV2O6_0),.din(w_dff_A_vqOlRl3Q0_0),.clk(gclk));
	jdff dff_A_UJhNnV2O6_0(.dout(w_dff_A_Mr6dVPRD9_0),.din(w_dff_A_UJhNnV2O6_0),.clk(gclk));
	jdff dff_A_Mr6dVPRD9_0(.dout(w_dff_A_2ayOVf0n1_0),.din(w_dff_A_Mr6dVPRD9_0),.clk(gclk));
	jdff dff_A_2ayOVf0n1_0(.dout(w_dff_A_wPTN0wP55_0),.din(w_dff_A_2ayOVf0n1_0),.clk(gclk));
	jdff dff_A_wPTN0wP55_0(.dout(w_dff_A_ACi7K8od9_0),.din(w_dff_A_wPTN0wP55_0),.clk(gclk));
	jdff dff_A_ACi7K8od9_0(.dout(w_dff_A_44a2eiLU9_0),.din(w_dff_A_ACi7K8od9_0),.clk(gclk));
	jdff dff_A_44a2eiLU9_0(.dout(w_dff_A_23gJRQ5g7_0),.din(w_dff_A_44a2eiLU9_0),.clk(gclk));
	jdff dff_A_23gJRQ5g7_0(.dout(w_dff_A_EhztXqOr7_0),.din(w_dff_A_23gJRQ5g7_0),.clk(gclk));
	jdff dff_A_EhztXqOr7_0(.dout(w_dff_A_ihWLOVIY5_0),.din(w_dff_A_EhztXqOr7_0),.clk(gclk));
	jdff dff_A_ihWLOVIY5_0(.dout(w_dff_A_eld0vHKq7_0),.din(w_dff_A_ihWLOVIY5_0),.clk(gclk));
	jdff dff_A_eld0vHKq7_0(.dout(w_dff_A_et9QRQjx2_0),.din(w_dff_A_eld0vHKq7_0),.clk(gclk));
	jdff dff_A_et9QRQjx2_0(.dout(w_dff_A_bq4bkuOx6_0),.din(w_dff_A_et9QRQjx2_0),.clk(gclk));
	jdff dff_A_bq4bkuOx6_0(.dout(w_dff_A_uAHb1l8Y4_0),.din(w_dff_A_bq4bkuOx6_0),.clk(gclk));
	jdff dff_A_uAHb1l8Y4_0(.dout(w_dff_A_xT3nxTPf5_0),.din(w_dff_A_uAHb1l8Y4_0),.clk(gclk));
	jdff dff_A_xT3nxTPf5_0(.dout(w_dff_A_7CDVaAUy7_0),.din(w_dff_A_xT3nxTPf5_0),.clk(gclk));
	jdff dff_A_7CDVaAUy7_0(.dout(w_dff_A_osUikJmw5_0),.din(w_dff_A_7CDVaAUy7_0),.clk(gclk));
	jdff dff_A_osUikJmw5_0(.dout(w_dff_A_I2bKiwRX6_0),.din(w_dff_A_osUikJmw5_0),.clk(gclk));
	jdff dff_A_I2bKiwRX6_0(.dout(w_dff_A_X3JIcfeP8_0),.din(w_dff_A_I2bKiwRX6_0),.clk(gclk));
	jdff dff_A_X3JIcfeP8_0(.dout(w_dff_A_yXilKSbz2_0),.din(w_dff_A_X3JIcfeP8_0),.clk(gclk));
	jdff dff_A_yXilKSbz2_0(.dout(w_dff_A_7BArrZLc7_0),.din(w_dff_A_yXilKSbz2_0),.clk(gclk));
	jdff dff_A_7BArrZLc7_0(.dout(w_dff_A_k9e5vIjO4_0),.din(w_dff_A_7BArrZLc7_0),.clk(gclk));
	jdff dff_A_k9e5vIjO4_0(.dout(w_dff_A_KPYifWeK0_0),.din(w_dff_A_k9e5vIjO4_0),.clk(gclk));
	jdff dff_A_KPYifWeK0_0(.dout(w_dff_A_gI5v4pFM6_0),.din(w_dff_A_KPYifWeK0_0),.clk(gclk));
	jdff dff_A_gI5v4pFM6_0(.dout(w_dff_A_NR8ptgg72_0),.din(w_dff_A_gI5v4pFM6_0),.clk(gclk));
	jdff dff_A_NR8ptgg72_0(.dout(w_dff_A_gh4Usdza2_0),.din(w_dff_A_NR8ptgg72_0),.clk(gclk));
	jdff dff_A_gh4Usdza2_0(.dout(w_dff_A_Y3nZJsFV5_0),.din(w_dff_A_gh4Usdza2_0),.clk(gclk));
	jdff dff_A_Y3nZJsFV5_0(.dout(w_dff_A_uAOadEvp4_0),.din(w_dff_A_Y3nZJsFV5_0),.clk(gclk));
	jdff dff_A_uAOadEvp4_0(.dout(w_dff_A_K3I5LBL13_0),.din(w_dff_A_uAOadEvp4_0),.clk(gclk));
	jdff dff_A_K3I5LBL13_0(.dout(w_dff_A_cnLgQGrX1_0),.din(w_dff_A_K3I5LBL13_0),.clk(gclk));
	jdff dff_A_cnLgQGrX1_0(.dout(w_dff_A_Lb5zGbly4_0),.din(w_dff_A_cnLgQGrX1_0),.clk(gclk));
	jdff dff_A_Lb5zGbly4_0(.dout(w_dff_A_iqgWX9BT3_0),.din(w_dff_A_Lb5zGbly4_0),.clk(gclk));
	jdff dff_A_iqgWX9BT3_0(.dout(w_dff_A_jzmE2qCb1_0),.din(w_dff_A_iqgWX9BT3_0),.clk(gclk));
	jdff dff_A_jzmE2qCb1_0(.dout(w_dff_A_sq9MCJmi6_0),.din(w_dff_A_jzmE2qCb1_0),.clk(gclk));
	jdff dff_A_sq9MCJmi6_0(.dout(w_dff_A_pT415re51_0),.din(w_dff_A_sq9MCJmi6_0),.clk(gclk));
	jdff dff_A_pT415re51_0(.dout(w_dff_A_5iaHRD7b2_0),.din(w_dff_A_pT415re51_0),.clk(gclk));
	jdff dff_A_5iaHRD7b2_0(.dout(w_dff_A_38zF5tBq1_0),.din(w_dff_A_5iaHRD7b2_0),.clk(gclk));
	jdff dff_A_38zF5tBq1_0(.dout(w_dff_A_2sRk0kPJ0_0),.din(w_dff_A_38zF5tBq1_0),.clk(gclk));
	jdff dff_A_2sRk0kPJ0_0(.dout(w_dff_A_ltnelA0H8_0),.din(w_dff_A_2sRk0kPJ0_0),.clk(gclk));
	jdff dff_A_ltnelA0H8_0(.dout(w_dff_A_7Pslk3Ky0_0),.din(w_dff_A_ltnelA0H8_0),.clk(gclk));
	jdff dff_A_7Pslk3Ky0_0(.dout(w_dff_A_C910CYpl6_0),.din(w_dff_A_7Pslk3Ky0_0),.clk(gclk));
	jdff dff_A_C910CYpl6_0(.dout(w_dff_A_3zgdTU2Q9_0),.din(w_dff_A_C910CYpl6_0),.clk(gclk));
	jdff dff_A_3zgdTU2Q9_0(.dout(w_dff_A_er3PfDBR0_0),.din(w_dff_A_3zgdTU2Q9_0),.clk(gclk));
	jdff dff_A_er3PfDBR0_0(.dout(w_dff_A_skDCO7qN4_0),.din(w_dff_A_er3PfDBR0_0),.clk(gclk));
	jdff dff_A_skDCO7qN4_0(.dout(w_dff_A_YhshNMAx9_0),.din(w_dff_A_skDCO7qN4_0),.clk(gclk));
	jdff dff_A_YhshNMAx9_0(.dout(w_dff_A_NPpsaEtJ7_0),.din(w_dff_A_YhshNMAx9_0),.clk(gclk));
	jdff dff_A_NPpsaEtJ7_0(.dout(w_dff_A_jo3nTC6z3_0),.din(w_dff_A_NPpsaEtJ7_0),.clk(gclk));
	jdff dff_A_jo3nTC6z3_0(.dout(w_dff_A_sl9S4LCA8_0),.din(w_dff_A_jo3nTC6z3_0),.clk(gclk));
	jdff dff_A_sl9S4LCA8_0(.dout(w_dff_A_0z457G1N3_0),.din(w_dff_A_sl9S4LCA8_0),.clk(gclk));
	jdff dff_A_0z457G1N3_0(.dout(w_dff_A_MLvBmDwZ0_0),.din(w_dff_A_0z457G1N3_0),.clk(gclk));
	jdff dff_A_MLvBmDwZ0_0(.dout(w_dff_A_eESDDvKH1_0),.din(w_dff_A_MLvBmDwZ0_0),.clk(gclk));
	jdff dff_A_eESDDvKH1_0(.dout(w_dff_A_lYy1cg6K2_0),.din(w_dff_A_eESDDvKH1_0),.clk(gclk));
	jdff dff_A_lYy1cg6K2_0(.dout(w_dff_A_GndAPpUj6_0),.din(w_dff_A_lYy1cg6K2_0),.clk(gclk));
	jdff dff_A_GndAPpUj6_0(.dout(w_dff_A_O1F8qIlQ6_0),.din(w_dff_A_GndAPpUj6_0),.clk(gclk));
	jdff dff_A_O1F8qIlQ6_0(.dout(w_dff_A_elzVeDOa0_0),.din(w_dff_A_O1F8qIlQ6_0),.clk(gclk));
	jdff dff_A_elzVeDOa0_0(.dout(w_dff_A_BWlKDNSe1_0),.din(w_dff_A_elzVeDOa0_0),.clk(gclk));
	jdff dff_A_BWlKDNSe1_0(.dout(w_dff_A_lIGMU9qz9_0),.din(w_dff_A_BWlKDNSe1_0),.clk(gclk));
	jdff dff_A_lIGMU9qz9_0(.dout(w_dff_A_zKZSf5z96_0),.din(w_dff_A_lIGMU9qz9_0),.clk(gclk));
	jdff dff_A_zKZSf5z96_0(.dout(G2877gat),.din(w_dff_A_zKZSf5z96_0),.clk(gclk));
	jdff dff_A_6toCtfid3_2(.dout(w_dff_A_1A78CLq23_0),.din(w_dff_A_6toCtfid3_2),.clk(gclk));
	jdff dff_A_1A78CLq23_0(.dout(w_dff_A_DT8YxD0y7_0),.din(w_dff_A_1A78CLq23_0),.clk(gclk));
	jdff dff_A_DT8YxD0y7_0(.dout(w_dff_A_4W3S1Zbk1_0),.din(w_dff_A_DT8YxD0y7_0),.clk(gclk));
	jdff dff_A_4W3S1Zbk1_0(.dout(w_dff_A_uwhYlclb7_0),.din(w_dff_A_4W3S1Zbk1_0),.clk(gclk));
	jdff dff_A_uwhYlclb7_0(.dout(w_dff_A_FpsAau1M8_0),.din(w_dff_A_uwhYlclb7_0),.clk(gclk));
	jdff dff_A_FpsAau1M8_0(.dout(w_dff_A_SpVZiSAV6_0),.din(w_dff_A_FpsAau1M8_0),.clk(gclk));
	jdff dff_A_SpVZiSAV6_0(.dout(w_dff_A_EwKqoT1F5_0),.din(w_dff_A_SpVZiSAV6_0),.clk(gclk));
	jdff dff_A_EwKqoT1F5_0(.dout(w_dff_A_rPgrdZFb1_0),.din(w_dff_A_EwKqoT1F5_0),.clk(gclk));
	jdff dff_A_rPgrdZFb1_0(.dout(w_dff_A_SomvLv1L6_0),.din(w_dff_A_rPgrdZFb1_0),.clk(gclk));
	jdff dff_A_SomvLv1L6_0(.dout(w_dff_A_9cUXX2Kj1_0),.din(w_dff_A_SomvLv1L6_0),.clk(gclk));
	jdff dff_A_9cUXX2Kj1_0(.dout(w_dff_A_q9RO1Lzg6_0),.din(w_dff_A_9cUXX2Kj1_0),.clk(gclk));
	jdff dff_A_q9RO1Lzg6_0(.dout(w_dff_A_Kk4RyuDK6_0),.din(w_dff_A_q9RO1Lzg6_0),.clk(gclk));
	jdff dff_A_Kk4RyuDK6_0(.dout(w_dff_A_P2tdFThs6_0),.din(w_dff_A_Kk4RyuDK6_0),.clk(gclk));
	jdff dff_A_P2tdFThs6_0(.dout(w_dff_A_7O78XgBo2_0),.din(w_dff_A_P2tdFThs6_0),.clk(gclk));
	jdff dff_A_7O78XgBo2_0(.dout(w_dff_A_rXPTY3mI5_0),.din(w_dff_A_7O78XgBo2_0),.clk(gclk));
	jdff dff_A_rXPTY3mI5_0(.dout(w_dff_A_muS7FTk72_0),.din(w_dff_A_rXPTY3mI5_0),.clk(gclk));
	jdff dff_A_muS7FTk72_0(.dout(w_dff_A_6ys0O7wf0_0),.din(w_dff_A_muS7FTk72_0),.clk(gclk));
	jdff dff_A_6ys0O7wf0_0(.dout(w_dff_A_BexIlYpB4_0),.din(w_dff_A_6ys0O7wf0_0),.clk(gclk));
	jdff dff_A_BexIlYpB4_0(.dout(w_dff_A_xhkygyeT1_0),.din(w_dff_A_BexIlYpB4_0),.clk(gclk));
	jdff dff_A_xhkygyeT1_0(.dout(w_dff_A_yg0mGmLT6_0),.din(w_dff_A_xhkygyeT1_0),.clk(gclk));
	jdff dff_A_yg0mGmLT6_0(.dout(w_dff_A_lApmStI82_0),.din(w_dff_A_yg0mGmLT6_0),.clk(gclk));
	jdff dff_A_lApmStI82_0(.dout(w_dff_A_r1any91t6_0),.din(w_dff_A_lApmStI82_0),.clk(gclk));
	jdff dff_A_r1any91t6_0(.dout(w_dff_A_TgB9vsIv2_0),.din(w_dff_A_r1any91t6_0),.clk(gclk));
	jdff dff_A_TgB9vsIv2_0(.dout(w_dff_A_1MSyKHFW4_0),.din(w_dff_A_TgB9vsIv2_0),.clk(gclk));
	jdff dff_A_1MSyKHFW4_0(.dout(w_dff_A_6OgsMwFq5_0),.din(w_dff_A_1MSyKHFW4_0),.clk(gclk));
	jdff dff_A_6OgsMwFq5_0(.dout(w_dff_A_Syyluhm85_0),.din(w_dff_A_6OgsMwFq5_0),.clk(gclk));
	jdff dff_A_Syyluhm85_0(.dout(w_dff_A_b4VCfP1L0_0),.din(w_dff_A_Syyluhm85_0),.clk(gclk));
	jdff dff_A_b4VCfP1L0_0(.dout(w_dff_A_JCARhnNj2_0),.din(w_dff_A_b4VCfP1L0_0),.clk(gclk));
	jdff dff_A_JCARhnNj2_0(.dout(w_dff_A_w5pCZ8tj4_0),.din(w_dff_A_JCARhnNj2_0),.clk(gclk));
	jdff dff_A_w5pCZ8tj4_0(.dout(w_dff_A_5kMaIGTd8_0),.din(w_dff_A_w5pCZ8tj4_0),.clk(gclk));
	jdff dff_A_5kMaIGTd8_0(.dout(w_dff_A_SYbL35Ts2_0),.din(w_dff_A_5kMaIGTd8_0),.clk(gclk));
	jdff dff_A_SYbL35Ts2_0(.dout(w_dff_A_rpveoWhk8_0),.din(w_dff_A_SYbL35Ts2_0),.clk(gclk));
	jdff dff_A_rpveoWhk8_0(.dout(w_dff_A_LUS4asnZ0_0),.din(w_dff_A_rpveoWhk8_0),.clk(gclk));
	jdff dff_A_LUS4asnZ0_0(.dout(w_dff_A_utui7ytj2_0),.din(w_dff_A_LUS4asnZ0_0),.clk(gclk));
	jdff dff_A_utui7ytj2_0(.dout(w_dff_A_Kcypql472_0),.din(w_dff_A_utui7ytj2_0),.clk(gclk));
	jdff dff_A_Kcypql472_0(.dout(w_dff_A_BA1l9tEx7_0),.din(w_dff_A_Kcypql472_0),.clk(gclk));
	jdff dff_A_BA1l9tEx7_0(.dout(w_dff_A_bVNmCXeP0_0),.din(w_dff_A_BA1l9tEx7_0),.clk(gclk));
	jdff dff_A_bVNmCXeP0_0(.dout(w_dff_A_eShxbMli4_0),.din(w_dff_A_bVNmCXeP0_0),.clk(gclk));
	jdff dff_A_eShxbMli4_0(.dout(w_dff_A_gx5S1IAV7_0),.din(w_dff_A_eShxbMli4_0),.clk(gclk));
	jdff dff_A_gx5S1IAV7_0(.dout(w_dff_A_sn3BQ7i11_0),.din(w_dff_A_gx5S1IAV7_0),.clk(gclk));
	jdff dff_A_sn3BQ7i11_0(.dout(w_dff_A_KqcQUQlx2_0),.din(w_dff_A_sn3BQ7i11_0),.clk(gclk));
	jdff dff_A_KqcQUQlx2_0(.dout(w_dff_A_OJdOHBX93_0),.din(w_dff_A_KqcQUQlx2_0),.clk(gclk));
	jdff dff_A_OJdOHBX93_0(.dout(w_dff_A_PPTuMW0k7_0),.din(w_dff_A_OJdOHBX93_0),.clk(gclk));
	jdff dff_A_PPTuMW0k7_0(.dout(w_dff_A_mtgH9WXw2_0),.din(w_dff_A_PPTuMW0k7_0),.clk(gclk));
	jdff dff_A_mtgH9WXw2_0(.dout(w_dff_A_jCkkOiMF2_0),.din(w_dff_A_mtgH9WXw2_0),.clk(gclk));
	jdff dff_A_jCkkOiMF2_0(.dout(w_dff_A_UNBsOa8C7_0),.din(w_dff_A_jCkkOiMF2_0),.clk(gclk));
	jdff dff_A_UNBsOa8C7_0(.dout(w_dff_A_S8XShES05_0),.din(w_dff_A_UNBsOa8C7_0),.clk(gclk));
	jdff dff_A_S8XShES05_0(.dout(w_dff_A_aYJ2pzRp7_0),.din(w_dff_A_S8XShES05_0),.clk(gclk));
	jdff dff_A_aYJ2pzRp7_0(.dout(w_dff_A_YxHxLVnZ8_0),.din(w_dff_A_aYJ2pzRp7_0),.clk(gclk));
	jdff dff_A_YxHxLVnZ8_0(.dout(w_dff_A_9ctmFtp53_0),.din(w_dff_A_YxHxLVnZ8_0),.clk(gclk));
	jdff dff_A_9ctmFtp53_0(.dout(w_dff_A_zIiicibX8_0),.din(w_dff_A_9ctmFtp53_0),.clk(gclk));
	jdff dff_A_zIiicibX8_0(.dout(w_dff_A_JgzCnWIR8_0),.din(w_dff_A_zIiicibX8_0),.clk(gclk));
	jdff dff_A_JgzCnWIR8_0(.dout(w_dff_A_tuDxqGzk5_0),.din(w_dff_A_JgzCnWIR8_0),.clk(gclk));
	jdff dff_A_tuDxqGzk5_0(.dout(w_dff_A_0Ucy4uLc4_0),.din(w_dff_A_tuDxqGzk5_0),.clk(gclk));
	jdff dff_A_0Ucy4uLc4_0(.dout(w_dff_A_50w7r7GH6_0),.din(w_dff_A_0Ucy4uLc4_0),.clk(gclk));
	jdff dff_A_50w7r7GH6_0(.dout(w_dff_A_unRZLVOU2_0),.din(w_dff_A_50w7r7GH6_0),.clk(gclk));
	jdff dff_A_unRZLVOU2_0(.dout(G3211gat),.din(w_dff_A_unRZLVOU2_0),.clk(gclk));
	jdff dff_A_oHiEz1mj9_2(.dout(w_dff_A_WWEIev9b4_0),.din(w_dff_A_oHiEz1mj9_2),.clk(gclk));
	jdff dff_A_WWEIev9b4_0(.dout(w_dff_A_uA6SoFcj8_0),.din(w_dff_A_WWEIev9b4_0),.clk(gclk));
	jdff dff_A_uA6SoFcj8_0(.dout(w_dff_A_Im5bakEX7_0),.din(w_dff_A_uA6SoFcj8_0),.clk(gclk));
	jdff dff_A_Im5bakEX7_0(.dout(w_dff_A_wwh3wwVl4_0),.din(w_dff_A_Im5bakEX7_0),.clk(gclk));
	jdff dff_A_wwh3wwVl4_0(.dout(w_dff_A_pCktsyqg6_0),.din(w_dff_A_wwh3wwVl4_0),.clk(gclk));
	jdff dff_A_pCktsyqg6_0(.dout(w_dff_A_XarRVOir2_0),.din(w_dff_A_pCktsyqg6_0),.clk(gclk));
	jdff dff_A_XarRVOir2_0(.dout(w_dff_A_ICpnhRlR4_0),.din(w_dff_A_XarRVOir2_0),.clk(gclk));
	jdff dff_A_ICpnhRlR4_0(.dout(w_dff_A_ElF2a2Pl4_0),.din(w_dff_A_ICpnhRlR4_0),.clk(gclk));
	jdff dff_A_ElF2a2Pl4_0(.dout(w_dff_A_dmInaRWU6_0),.din(w_dff_A_ElF2a2Pl4_0),.clk(gclk));
	jdff dff_A_dmInaRWU6_0(.dout(w_dff_A_8chgmXkn3_0),.din(w_dff_A_dmInaRWU6_0),.clk(gclk));
	jdff dff_A_8chgmXkn3_0(.dout(w_dff_A_aIfZjx4G2_0),.din(w_dff_A_8chgmXkn3_0),.clk(gclk));
	jdff dff_A_aIfZjx4G2_0(.dout(w_dff_A_czBZEWN88_0),.din(w_dff_A_aIfZjx4G2_0),.clk(gclk));
	jdff dff_A_czBZEWN88_0(.dout(w_dff_A_YpT2eter7_0),.din(w_dff_A_czBZEWN88_0),.clk(gclk));
	jdff dff_A_YpT2eter7_0(.dout(w_dff_A_GRhhVCMk5_0),.din(w_dff_A_YpT2eter7_0),.clk(gclk));
	jdff dff_A_GRhhVCMk5_0(.dout(w_dff_A_26MYKpXU1_0),.din(w_dff_A_GRhhVCMk5_0),.clk(gclk));
	jdff dff_A_26MYKpXU1_0(.dout(w_dff_A_7M7Y0dV11_0),.din(w_dff_A_26MYKpXU1_0),.clk(gclk));
	jdff dff_A_7M7Y0dV11_0(.dout(w_dff_A_8plRAxtm9_0),.din(w_dff_A_7M7Y0dV11_0),.clk(gclk));
	jdff dff_A_8plRAxtm9_0(.dout(w_dff_A_dSTa3YCe5_0),.din(w_dff_A_8plRAxtm9_0),.clk(gclk));
	jdff dff_A_dSTa3YCe5_0(.dout(w_dff_A_8ryPOv5L2_0),.din(w_dff_A_dSTa3YCe5_0),.clk(gclk));
	jdff dff_A_8ryPOv5L2_0(.dout(w_dff_A_0vaBFGXN1_0),.din(w_dff_A_8ryPOv5L2_0),.clk(gclk));
	jdff dff_A_0vaBFGXN1_0(.dout(w_dff_A_QMaXO7Iw3_0),.din(w_dff_A_0vaBFGXN1_0),.clk(gclk));
	jdff dff_A_QMaXO7Iw3_0(.dout(w_dff_A_HocgjUo00_0),.din(w_dff_A_QMaXO7Iw3_0),.clk(gclk));
	jdff dff_A_HocgjUo00_0(.dout(w_dff_A_SLpt4ERs3_0),.din(w_dff_A_HocgjUo00_0),.clk(gclk));
	jdff dff_A_SLpt4ERs3_0(.dout(w_dff_A_qyeJ6crN4_0),.din(w_dff_A_SLpt4ERs3_0),.clk(gclk));
	jdff dff_A_qyeJ6crN4_0(.dout(w_dff_A_WJ0JzlSi6_0),.din(w_dff_A_qyeJ6crN4_0),.clk(gclk));
	jdff dff_A_WJ0JzlSi6_0(.dout(w_dff_A_hHFyBcm03_0),.din(w_dff_A_WJ0JzlSi6_0),.clk(gclk));
	jdff dff_A_hHFyBcm03_0(.dout(w_dff_A_J2WU4fNO3_0),.din(w_dff_A_hHFyBcm03_0),.clk(gclk));
	jdff dff_A_J2WU4fNO3_0(.dout(w_dff_A_jIC19Oib5_0),.din(w_dff_A_J2WU4fNO3_0),.clk(gclk));
	jdff dff_A_jIC19Oib5_0(.dout(w_dff_A_4towJrA42_0),.din(w_dff_A_jIC19Oib5_0),.clk(gclk));
	jdff dff_A_4towJrA42_0(.dout(w_dff_A_W70XScJL3_0),.din(w_dff_A_4towJrA42_0),.clk(gclk));
	jdff dff_A_W70XScJL3_0(.dout(w_dff_A_su1sO7qz0_0),.din(w_dff_A_W70XScJL3_0),.clk(gclk));
	jdff dff_A_su1sO7qz0_0(.dout(w_dff_A_Nb2pKhfa6_0),.din(w_dff_A_su1sO7qz0_0),.clk(gclk));
	jdff dff_A_Nb2pKhfa6_0(.dout(w_dff_A_eBsCWehA7_0),.din(w_dff_A_Nb2pKhfa6_0),.clk(gclk));
	jdff dff_A_eBsCWehA7_0(.dout(w_dff_A_wn4ZLpoS3_0),.din(w_dff_A_eBsCWehA7_0),.clk(gclk));
	jdff dff_A_wn4ZLpoS3_0(.dout(w_dff_A_alTNogDg2_0),.din(w_dff_A_wn4ZLpoS3_0),.clk(gclk));
	jdff dff_A_alTNogDg2_0(.dout(w_dff_A_tdBlQ9uE9_0),.din(w_dff_A_alTNogDg2_0),.clk(gclk));
	jdff dff_A_tdBlQ9uE9_0(.dout(w_dff_A_PVQwOhb35_0),.din(w_dff_A_tdBlQ9uE9_0),.clk(gclk));
	jdff dff_A_PVQwOhb35_0(.dout(w_dff_A_qkcyUDQB5_0),.din(w_dff_A_PVQwOhb35_0),.clk(gclk));
	jdff dff_A_qkcyUDQB5_0(.dout(w_dff_A_9uT8iI8J1_0),.din(w_dff_A_qkcyUDQB5_0),.clk(gclk));
	jdff dff_A_9uT8iI8J1_0(.dout(w_dff_A_KIEFJ4uB8_0),.din(w_dff_A_9uT8iI8J1_0),.clk(gclk));
	jdff dff_A_KIEFJ4uB8_0(.dout(w_dff_A_SshSlihQ9_0),.din(w_dff_A_KIEFJ4uB8_0),.clk(gclk));
	jdff dff_A_SshSlihQ9_0(.dout(w_dff_A_2DiWrGUt5_0),.din(w_dff_A_SshSlihQ9_0),.clk(gclk));
	jdff dff_A_2DiWrGUt5_0(.dout(w_dff_A_KCmVgIDG9_0),.din(w_dff_A_2DiWrGUt5_0),.clk(gclk));
	jdff dff_A_KCmVgIDG9_0(.dout(w_dff_A_KGvGrEZY2_0),.din(w_dff_A_KCmVgIDG9_0),.clk(gclk));
	jdff dff_A_KGvGrEZY2_0(.dout(w_dff_A_c4XxgjSx9_0),.din(w_dff_A_KGvGrEZY2_0),.clk(gclk));
	jdff dff_A_c4XxgjSx9_0(.dout(w_dff_A_eR3kaN9e3_0),.din(w_dff_A_c4XxgjSx9_0),.clk(gclk));
	jdff dff_A_eR3kaN9e3_0(.dout(w_dff_A_wVtDgxO92_0),.din(w_dff_A_eR3kaN9e3_0),.clk(gclk));
	jdff dff_A_wVtDgxO92_0(.dout(w_dff_A_vS3u9BTU9_0),.din(w_dff_A_wVtDgxO92_0),.clk(gclk));
	jdff dff_A_vS3u9BTU9_0(.dout(w_dff_A_71hOUxa46_0),.din(w_dff_A_vS3u9BTU9_0),.clk(gclk));
	jdff dff_A_71hOUxa46_0(.dout(w_dff_A_wCDoon3U0_0),.din(w_dff_A_71hOUxa46_0),.clk(gclk));
	jdff dff_A_wCDoon3U0_0(.dout(w_dff_A_VRpSlWHe7_0),.din(w_dff_A_wCDoon3U0_0),.clk(gclk));
	jdff dff_A_VRpSlWHe7_0(.dout(w_dff_A_mO9XADgl5_0),.din(w_dff_A_VRpSlWHe7_0),.clk(gclk));
	jdff dff_A_mO9XADgl5_0(.dout(w_dff_A_mAXKtItz3_0),.din(w_dff_A_mO9XADgl5_0),.clk(gclk));
	jdff dff_A_mAXKtItz3_0(.dout(G3552gat),.din(w_dff_A_mAXKtItz3_0),.clk(gclk));
	jdff dff_A_Rbm3HLMi5_2(.dout(w_dff_A_171O33842_0),.din(w_dff_A_Rbm3HLMi5_2),.clk(gclk));
	jdff dff_A_171O33842_0(.dout(w_dff_A_DgfunnHf5_0),.din(w_dff_A_171O33842_0),.clk(gclk));
	jdff dff_A_DgfunnHf5_0(.dout(w_dff_A_1XEqnQNl3_0),.din(w_dff_A_DgfunnHf5_0),.clk(gclk));
	jdff dff_A_1XEqnQNl3_0(.dout(w_dff_A_Itlvq3gT1_0),.din(w_dff_A_1XEqnQNl3_0),.clk(gclk));
	jdff dff_A_Itlvq3gT1_0(.dout(w_dff_A_AQvVTgB18_0),.din(w_dff_A_Itlvq3gT1_0),.clk(gclk));
	jdff dff_A_AQvVTgB18_0(.dout(w_dff_A_rt7aZmnp6_0),.din(w_dff_A_AQvVTgB18_0),.clk(gclk));
	jdff dff_A_rt7aZmnp6_0(.dout(w_dff_A_rYS2JgCZ8_0),.din(w_dff_A_rt7aZmnp6_0),.clk(gclk));
	jdff dff_A_rYS2JgCZ8_0(.dout(w_dff_A_n08vK04M5_0),.din(w_dff_A_rYS2JgCZ8_0),.clk(gclk));
	jdff dff_A_n08vK04M5_0(.dout(w_dff_A_A9qrLozT8_0),.din(w_dff_A_n08vK04M5_0),.clk(gclk));
	jdff dff_A_A9qrLozT8_0(.dout(w_dff_A_STfqNvTT5_0),.din(w_dff_A_A9qrLozT8_0),.clk(gclk));
	jdff dff_A_STfqNvTT5_0(.dout(w_dff_A_DLGn9dEN8_0),.din(w_dff_A_STfqNvTT5_0),.clk(gclk));
	jdff dff_A_DLGn9dEN8_0(.dout(w_dff_A_q4Bm408v2_0),.din(w_dff_A_DLGn9dEN8_0),.clk(gclk));
	jdff dff_A_q4Bm408v2_0(.dout(w_dff_A_xtWdB1hM3_0),.din(w_dff_A_q4Bm408v2_0),.clk(gclk));
	jdff dff_A_xtWdB1hM3_0(.dout(w_dff_A_rdPXo40U9_0),.din(w_dff_A_xtWdB1hM3_0),.clk(gclk));
	jdff dff_A_rdPXo40U9_0(.dout(w_dff_A_0EUS7Gy69_0),.din(w_dff_A_rdPXo40U9_0),.clk(gclk));
	jdff dff_A_0EUS7Gy69_0(.dout(w_dff_A_m60602m17_0),.din(w_dff_A_0EUS7Gy69_0),.clk(gclk));
	jdff dff_A_m60602m17_0(.dout(w_dff_A_UsNhS3ZC6_0),.din(w_dff_A_m60602m17_0),.clk(gclk));
	jdff dff_A_UsNhS3ZC6_0(.dout(w_dff_A_JUsV8DUM7_0),.din(w_dff_A_UsNhS3ZC6_0),.clk(gclk));
	jdff dff_A_JUsV8DUM7_0(.dout(w_dff_A_PprRIjDj7_0),.din(w_dff_A_JUsV8DUM7_0),.clk(gclk));
	jdff dff_A_PprRIjDj7_0(.dout(w_dff_A_VG0Dc0401_0),.din(w_dff_A_PprRIjDj7_0),.clk(gclk));
	jdff dff_A_VG0Dc0401_0(.dout(w_dff_A_w6xc5oFK2_0),.din(w_dff_A_VG0Dc0401_0),.clk(gclk));
	jdff dff_A_w6xc5oFK2_0(.dout(w_dff_A_DAZddbCR9_0),.din(w_dff_A_w6xc5oFK2_0),.clk(gclk));
	jdff dff_A_DAZddbCR9_0(.dout(w_dff_A_e4Zjc54A7_0),.din(w_dff_A_DAZddbCR9_0),.clk(gclk));
	jdff dff_A_e4Zjc54A7_0(.dout(w_dff_A_IvS6FEvt9_0),.din(w_dff_A_e4Zjc54A7_0),.clk(gclk));
	jdff dff_A_IvS6FEvt9_0(.dout(w_dff_A_N0mB9gaT8_0),.din(w_dff_A_IvS6FEvt9_0),.clk(gclk));
	jdff dff_A_N0mB9gaT8_0(.dout(w_dff_A_S3Cycj0C1_0),.din(w_dff_A_N0mB9gaT8_0),.clk(gclk));
	jdff dff_A_S3Cycj0C1_0(.dout(w_dff_A_vIrNo3oQ7_0),.din(w_dff_A_S3Cycj0C1_0),.clk(gclk));
	jdff dff_A_vIrNo3oQ7_0(.dout(w_dff_A_Qt9cfgkr9_0),.din(w_dff_A_vIrNo3oQ7_0),.clk(gclk));
	jdff dff_A_Qt9cfgkr9_0(.dout(w_dff_A_dtsgTO692_0),.din(w_dff_A_Qt9cfgkr9_0),.clk(gclk));
	jdff dff_A_dtsgTO692_0(.dout(w_dff_A_xXp27jWL2_0),.din(w_dff_A_dtsgTO692_0),.clk(gclk));
	jdff dff_A_xXp27jWL2_0(.dout(w_dff_A_oaq6qhw19_0),.din(w_dff_A_xXp27jWL2_0),.clk(gclk));
	jdff dff_A_oaq6qhw19_0(.dout(w_dff_A_sPKFS5bJ4_0),.din(w_dff_A_oaq6qhw19_0),.clk(gclk));
	jdff dff_A_sPKFS5bJ4_0(.dout(w_dff_A_H3oeM2KD5_0),.din(w_dff_A_sPKFS5bJ4_0),.clk(gclk));
	jdff dff_A_H3oeM2KD5_0(.dout(w_dff_A_EdoQ8exD1_0),.din(w_dff_A_H3oeM2KD5_0),.clk(gclk));
	jdff dff_A_EdoQ8exD1_0(.dout(w_dff_A_oz8yjHUa0_0),.din(w_dff_A_EdoQ8exD1_0),.clk(gclk));
	jdff dff_A_oz8yjHUa0_0(.dout(w_dff_A_wxH53mKv5_0),.din(w_dff_A_oz8yjHUa0_0),.clk(gclk));
	jdff dff_A_wxH53mKv5_0(.dout(w_dff_A_UXx9YtCx2_0),.din(w_dff_A_wxH53mKv5_0),.clk(gclk));
	jdff dff_A_UXx9YtCx2_0(.dout(w_dff_A_Fs05k84w1_0),.din(w_dff_A_UXx9YtCx2_0),.clk(gclk));
	jdff dff_A_Fs05k84w1_0(.dout(w_dff_A_ukihaXIE7_0),.din(w_dff_A_Fs05k84w1_0),.clk(gclk));
	jdff dff_A_ukihaXIE7_0(.dout(w_dff_A_LsGwcZjm2_0),.din(w_dff_A_ukihaXIE7_0),.clk(gclk));
	jdff dff_A_LsGwcZjm2_0(.dout(w_dff_A_CilGgzuw8_0),.din(w_dff_A_LsGwcZjm2_0),.clk(gclk));
	jdff dff_A_CilGgzuw8_0(.dout(w_dff_A_cmY3SbYL4_0),.din(w_dff_A_CilGgzuw8_0),.clk(gclk));
	jdff dff_A_cmY3SbYL4_0(.dout(w_dff_A_vGdK8Ez57_0),.din(w_dff_A_cmY3SbYL4_0),.clk(gclk));
	jdff dff_A_vGdK8Ez57_0(.dout(w_dff_A_efN5jWQA2_0),.din(w_dff_A_vGdK8Ez57_0),.clk(gclk));
	jdff dff_A_efN5jWQA2_0(.dout(w_dff_A_N5qTMZjD4_0),.din(w_dff_A_efN5jWQA2_0),.clk(gclk));
	jdff dff_A_N5qTMZjD4_0(.dout(w_dff_A_qi3aoIvW9_0),.din(w_dff_A_N5qTMZjD4_0),.clk(gclk));
	jdff dff_A_qi3aoIvW9_0(.dout(w_dff_A_VLbPaEW49_0),.din(w_dff_A_qi3aoIvW9_0),.clk(gclk));
	jdff dff_A_VLbPaEW49_0(.dout(w_dff_A_lHUTu3Ql0_0),.din(w_dff_A_VLbPaEW49_0),.clk(gclk));
	jdff dff_A_lHUTu3Ql0_0(.dout(w_dff_A_lcM46GUp5_0),.din(w_dff_A_lHUTu3Ql0_0),.clk(gclk));
	jdff dff_A_lcM46GUp5_0(.dout(w_dff_A_3EWNILvx8_0),.din(w_dff_A_lcM46GUp5_0),.clk(gclk));
	jdff dff_A_3EWNILvx8_0(.dout(G3895gat),.din(w_dff_A_3EWNILvx8_0),.clk(gclk));
	jdff dff_A_nwOyaoey4_2(.dout(w_dff_A_X9oxnlGG7_0),.din(w_dff_A_nwOyaoey4_2),.clk(gclk));
	jdff dff_A_X9oxnlGG7_0(.dout(w_dff_A_MdrQzZCY2_0),.din(w_dff_A_X9oxnlGG7_0),.clk(gclk));
	jdff dff_A_MdrQzZCY2_0(.dout(w_dff_A_VplQJjIg6_0),.din(w_dff_A_MdrQzZCY2_0),.clk(gclk));
	jdff dff_A_VplQJjIg6_0(.dout(w_dff_A_Jk7DRYxx6_0),.din(w_dff_A_VplQJjIg6_0),.clk(gclk));
	jdff dff_A_Jk7DRYxx6_0(.dout(w_dff_A_xGAsp6qN3_0),.din(w_dff_A_Jk7DRYxx6_0),.clk(gclk));
	jdff dff_A_xGAsp6qN3_0(.dout(w_dff_A_EMZY7AgU3_0),.din(w_dff_A_xGAsp6qN3_0),.clk(gclk));
	jdff dff_A_EMZY7AgU3_0(.dout(w_dff_A_tmHqdvq06_0),.din(w_dff_A_EMZY7AgU3_0),.clk(gclk));
	jdff dff_A_tmHqdvq06_0(.dout(w_dff_A_SdTKA03y4_0),.din(w_dff_A_tmHqdvq06_0),.clk(gclk));
	jdff dff_A_SdTKA03y4_0(.dout(w_dff_A_dCdlsUtN6_0),.din(w_dff_A_SdTKA03y4_0),.clk(gclk));
	jdff dff_A_dCdlsUtN6_0(.dout(w_dff_A_Rh70a2QI7_0),.din(w_dff_A_dCdlsUtN6_0),.clk(gclk));
	jdff dff_A_Rh70a2QI7_0(.dout(w_dff_A_NYsT8Ru43_0),.din(w_dff_A_Rh70a2QI7_0),.clk(gclk));
	jdff dff_A_NYsT8Ru43_0(.dout(w_dff_A_hz06ag0v6_0),.din(w_dff_A_NYsT8Ru43_0),.clk(gclk));
	jdff dff_A_hz06ag0v6_0(.dout(w_dff_A_z7HCUJXW2_0),.din(w_dff_A_hz06ag0v6_0),.clk(gclk));
	jdff dff_A_z7HCUJXW2_0(.dout(w_dff_A_htzWotAw5_0),.din(w_dff_A_z7HCUJXW2_0),.clk(gclk));
	jdff dff_A_htzWotAw5_0(.dout(w_dff_A_bDjX3uyT9_0),.din(w_dff_A_htzWotAw5_0),.clk(gclk));
	jdff dff_A_bDjX3uyT9_0(.dout(w_dff_A_8JbD8Mhb1_0),.din(w_dff_A_bDjX3uyT9_0),.clk(gclk));
	jdff dff_A_8JbD8Mhb1_0(.dout(w_dff_A_lmeM88u52_0),.din(w_dff_A_8JbD8Mhb1_0),.clk(gclk));
	jdff dff_A_lmeM88u52_0(.dout(w_dff_A_cDuUjgib5_0),.din(w_dff_A_lmeM88u52_0),.clk(gclk));
	jdff dff_A_cDuUjgib5_0(.dout(w_dff_A_hAmdzvUy5_0),.din(w_dff_A_cDuUjgib5_0),.clk(gclk));
	jdff dff_A_hAmdzvUy5_0(.dout(w_dff_A_tBiijj7F5_0),.din(w_dff_A_hAmdzvUy5_0),.clk(gclk));
	jdff dff_A_tBiijj7F5_0(.dout(w_dff_A_iCFNLp680_0),.din(w_dff_A_tBiijj7F5_0),.clk(gclk));
	jdff dff_A_iCFNLp680_0(.dout(w_dff_A_FfWlSijm1_0),.din(w_dff_A_iCFNLp680_0),.clk(gclk));
	jdff dff_A_FfWlSijm1_0(.dout(w_dff_A_oI5hKF827_0),.din(w_dff_A_FfWlSijm1_0),.clk(gclk));
	jdff dff_A_oI5hKF827_0(.dout(w_dff_A_eL1AppEj4_0),.din(w_dff_A_oI5hKF827_0),.clk(gclk));
	jdff dff_A_eL1AppEj4_0(.dout(w_dff_A_o8ntKq7g2_0),.din(w_dff_A_eL1AppEj4_0),.clk(gclk));
	jdff dff_A_o8ntKq7g2_0(.dout(w_dff_A_xxlrpDic0_0),.din(w_dff_A_o8ntKq7g2_0),.clk(gclk));
	jdff dff_A_xxlrpDic0_0(.dout(w_dff_A_bryDQU6H2_0),.din(w_dff_A_xxlrpDic0_0),.clk(gclk));
	jdff dff_A_bryDQU6H2_0(.dout(w_dff_A_OnUyEe4a4_0),.din(w_dff_A_bryDQU6H2_0),.clk(gclk));
	jdff dff_A_OnUyEe4a4_0(.dout(w_dff_A_b1OGVNak8_0),.din(w_dff_A_OnUyEe4a4_0),.clk(gclk));
	jdff dff_A_b1OGVNak8_0(.dout(w_dff_A_pdhXn80u2_0),.din(w_dff_A_b1OGVNak8_0),.clk(gclk));
	jdff dff_A_pdhXn80u2_0(.dout(w_dff_A_mJ2pnWn60_0),.din(w_dff_A_pdhXn80u2_0),.clk(gclk));
	jdff dff_A_mJ2pnWn60_0(.dout(w_dff_A_UhzvvQa80_0),.din(w_dff_A_mJ2pnWn60_0),.clk(gclk));
	jdff dff_A_UhzvvQa80_0(.dout(w_dff_A_E0O0qPjW6_0),.din(w_dff_A_UhzvvQa80_0),.clk(gclk));
	jdff dff_A_E0O0qPjW6_0(.dout(w_dff_A_3f0HYPBW2_0),.din(w_dff_A_E0O0qPjW6_0),.clk(gclk));
	jdff dff_A_3f0HYPBW2_0(.dout(w_dff_A_VnIb08re1_0),.din(w_dff_A_3f0HYPBW2_0),.clk(gclk));
	jdff dff_A_VnIb08re1_0(.dout(w_dff_A_4ELMRuYw3_0),.din(w_dff_A_VnIb08re1_0),.clk(gclk));
	jdff dff_A_4ELMRuYw3_0(.dout(w_dff_A_iTXTK2Dw1_0),.din(w_dff_A_4ELMRuYw3_0),.clk(gclk));
	jdff dff_A_iTXTK2Dw1_0(.dout(w_dff_A_pPoAfbmZ8_0),.din(w_dff_A_iTXTK2Dw1_0),.clk(gclk));
	jdff dff_A_pPoAfbmZ8_0(.dout(w_dff_A_P4bBWatu1_0),.din(w_dff_A_pPoAfbmZ8_0),.clk(gclk));
	jdff dff_A_P4bBWatu1_0(.dout(w_dff_A_5uOQzi5I1_0),.din(w_dff_A_P4bBWatu1_0),.clk(gclk));
	jdff dff_A_5uOQzi5I1_0(.dout(w_dff_A_W1c0Qucw6_0),.din(w_dff_A_5uOQzi5I1_0),.clk(gclk));
	jdff dff_A_W1c0Qucw6_0(.dout(w_dff_A_XMNoKD2T4_0),.din(w_dff_A_W1c0Qucw6_0),.clk(gclk));
	jdff dff_A_XMNoKD2T4_0(.dout(w_dff_A_Ob7pC4jD4_0),.din(w_dff_A_XMNoKD2T4_0),.clk(gclk));
	jdff dff_A_Ob7pC4jD4_0(.dout(w_dff_A_Fa1pGlJZ8_0),.din(w_dff_A_Ob7pC4jD4_0),.clk(gclk));
	jdff dff_A_Fa1pGlJZ8_0(.dout(w_dff_A_KAdki1ij5_0),.din(w_dff_A_Fa1pGlJZ8_0),.clk(gclk));
	jdff dff_A_KAdki1ij5_0(.dout(w_dff_A_Wja5gqcN2_0),.din(w_dff_A_KAdki1ij5_0),.clk(gclk));
	jdff dff_A_Wja5gqcN2_0(.dout(w_dff_A_YIEnXGgf1_0),.din(w_dff_A_Wja5gqcN2_0),.clk(gclk));
	jdff dff_A_YIEnXGgf1_0(.dout(G4241gat),.din(w_dff_A_YIEnXGgf1_0),.clk(gclk));
	jdff dff_A_Vd7i4kR94_2(.dout(w_dff_A_Pu9Wjaa81_0),.din(w_dff_A_Vd7i4kR94_2),.clk(gclk));
	jdff dff_A_Pu9Wjaa81_0(.dout(w_dff_A_y832RBgu8_0),.din(w_dff_A_Pu9Wjaa81_0),.clk(gclk));
	jdff dff_A_y832RBgu8_0(.dout(w_dff_A_2HY3uVQV7_0),.din(w_dff_A_y832RBgu8_0),.clk(gclk));
	jdff dff_A_2HY3uVQV7_0(.dout(w_dff_A_Eh1vioIX1_0),.din(w_dff_A_2HY3uVQV7_0),.clk(gclk));
	jdff dff_A_Eh1vioIX1_0(.dout(w_dff_A_U6Jo0qeT7_0),.din(w_dff_A_Eh1vioIX1_0),.clk(gclk));
	jdff dff_A_U6Jo0qeT7_0(.dout(w_dff_A_qrJIZ9aJ4_0),.din(w_dff_A_U6Jo0qeT7_0),.clk(gclk));
	jdff dff_A_qrJIZ9aJ4_0(.dout(w_dff_A_QOg5krL15_0),.din(w_dff_A_qrJIZ9aJ4_0),.clk(gclk));
	jdff dff_A_QOg5krL15_0(.dout(w_dff_A_PeBKsD8r3_0),.din(w_dff_A_QOg5krL15_0),.clk(gclk));
	jdff dff_A_PeBKsD8r3_0(.dout(w_dff_A_ruFNp6fX8_0),.din(w_dff_A_PeBKsD8r3_0),.clk(gclk));
	jdff dff_A_ruFNp6fX8_0(.dout(w_dff_A_voWj35FN8_0),.din(w_dff_A_ruFNp6fX8_0),.clk(gclk));
	jdff dff_A_voWj35FN8_0(.dout(w_dff_A_sXUZFv1v8_0),.din(w_dff_A_voWj35FN8_0),.clk(gclk));
	jdff dff_A_sXUZFv1v8_0(.dout(w_dff_A_rVMVXYnb2_0),.din(w_dff_A_sXUZFv1v8_0),.clk(gclk));
	jdff dff_A_rVMVXYnb2_0(.dout(w_dff_A_ngOg0wGB5_0),.din(w_dff_A_rVMVXYnb2_0),.clk(gclk));
	jdff dff_A_ngOg0wGB5_0(.dout(w_dff_A_YbGuxqbD1_0),.din(w_dff_A_ngOg0wGB5_0),.clk(gclk));
	jdff dff_A_YbGuxqbD1_0(.dout(w_dff_A_ibqyDZsC2_0),.din(w_dff_A_YbGuxqbD1_0),.clk(gclk));
	jdff dff_A_ibqyDZsC2_0(.dout(w_dff_A_mEkAvLwo5_0),.din(w_dff_A_ibqyDZsC2_0),.clk(gclk));
	jdff dff_A_mEkAvLwo5_0(.dout(w_dff_A_9JRzzrQQ1_0),.din(w_dff_A_mEkAvLwo5_0),.clk(gclk));
	jdff dff_A_9JRzzrQQ1_0(.dout(w_dff_A_PfmQXbOq6_0),.din(w_dff_A_9JRzzrQQ1_0),.clk(gclk));
	jdff dff_A_PfmQXbOq6_0(.dout(w_dff_A_5iqj2tZi3_0),.din(w_dff_A_PfmQXbOq6_0),.clk(gclk));
	jdff dff_A_5iqj2tZi3_0(.dout(w_dff_A_lB2yMDCX9_0),.din(w_dff_A_5iqj2tZi3_0),.clk(gclk));
	jdff dff_A_lB2yMDCX9_0(.dout(w_dff_A_f3F18Xvh9_0),.din(w_dff_A_lB2yMDCX9_0),.clk(gclk));
	jdff dff_A_f3F18Xvh9_0(.dout(w_dff_A_CAV4BSWD0_0),.din(w_dff_A_f3F18Xvh9_0),.clk(gclk));
	jdff dff_A_CAV4BSWD0_0(.dout(w_dff_A_K8iX0db10_0),.din(w_dff_A_CAV4BSWD0_0),.clk(gclk));
	jdff dff_A_K8iX0db10_0(.dout(w_dff_A_Z8TAfvkZ8_0),.din(w_dff_A_K8iX0db10_0),.clk(gclk));
	jdff dff_A_Z8TAfvkZ8_0(.dout(w_dff_A_3YbNqBzd0_0),.din(w_dff_A_Z8TAfvkZ8_0),.clk(gclk));
	jdff dff_A_3YbNqBzd0_0(.dout(w_dff_A_BrkJvYdD8_0),.din(w_dff_A_3YbNqBzd0_0),.clk(gclk));
	jdff dff_A_BrkJvYdD8_0(.dout(w_dff_A_DhkUnXQC1_0),.din(w_dff_A_BrkJvYdD8_0),.clk(gclk));
	jdff dff_A_DhkUnXQC1_0(.dout(w_dff_A_nd5FsRW52_0),.din(w_dff_A_DhkUnXQC1_0),.clk(gclk));
	jdff dff_A_nd5FsRW52_0(.dout(w_dff_A_nBhH7AQT1_0),.din(w_dff_A_nd5FsRW52_0),.clk(gclk));
	jdff dff_A_nBhH7AQT1_0(.dout(w_dff_A_MwUq6KdQ6_0),.din(w_dff_A_nBhH7AQT1_0),.clk(gclk));
	jdff dff_A_MwUq6KdQ6_0(.dout(w_dff_A_Bp9tMnD25_0),.din(w_dff_A_MwUq6KdQ6_0),.clk(gclk));
	jdff dff_A_Bp9tMnD25_0(.dout(w_dff_A_n2iIoE575_0),.din(w_dff_A_Bp9tMnD25_0),.clk(gclk));
	jdff dff_A_n2iIoE575_0(.dout(w_dff_A_HNyFd3XT2_0),.din(w_dff_A_n2iIoE575_0),.clk(gclk));
	jdff dff_A_HNyFd3XT2_0(.dout(w_dff_A_f0fxSfn54_0),.din(w_dff_A_HNyFd3XT2_0),.clk(gclk));
	jdff dff_A_f0fxSfn54_0(.dout(w_dff_A_bI00JPe37_0),.din(w_dff_A_f0fxSfn54_0),.clk(gclk));
	jdff dff_A_bI00JPe37_0(.dout(w_dff_A_0sIfIjAV3_0),.din(w_dff_A_bI00JPe37_0),.clk(gclk));
	jdff dff_A_0sIfIjAV3_0(.dout(w_dff_A_CKX7qzNz6_0),.din(w_dff_A_0sIfIjAV3_0),.clk(gclk));
	jdff dff_A_CKX7qzNz6_0(.dout(w_dff_A_g7OldxJj7_0),.din(w_dff_A_CKX7qzNz6_0),.clk(gclk));
	jdff dff_A_g7OldxJj7_0(.dout(w_dff_A_1dQWdZgN8_0),.din(w_dff_A_g7OldxJj7_0),.clk(gclk));
	jdff dff_A_1dQWdZgN8_0(.dout(w_dff_A_PbxyKYi87_0),.din(w_dff_A_1dQWdZgN8_0),.clk(gclk));
	jdff dff_A_PbxyKYi87_0(.dout(w_dff_A_2KYOE4Va3_0),.din(w_dff_A_PbxyKYi87_0),.clk(gclk));
	jdff dff_A_2KYOE4Va3_0(.dout(w_dff_A_escM5kvZ4_0),.din(w_dff_A_2KYOE4Va3_0),.clk(gclk));
	jdff dff_A_escM5kvZ4_0(.dout(w_dff_A_NlBn5b4h2_0),.din(w_dff_A_escM5kvZ4_0),.clk(gclk));
	jdff dff_A_NlBn5b4h2_0(.dout(w_dff_A_XNdtygn63_0),.din(w_dff_A_NlBn5b4h2_0),.clk(gclk));
	jdff dff_A_XNdtygn63_0(.dout(G4591gat),.din(w_dff_A_XNdtygn63_0),.clk(gclk));
	jdff dff_A_guWKCtIU7_2(.dout(w_dff_A_lZJWPPFQ8_0),.din(w_dff_A_guWKCtIU7_2),.clk(gclk));
	jdff dff_A_lZJWPPFQ8_0(.dout(w_dff_A_SRBWEpiC6_0),.din(w_dff_A_lZJWPPFQ8_0),.clk(gclk));
	jdff dff_A_SRBWEpiC6_0(.dout(w_dff_A_JN3xHNET9_0),.din(w_dff_A_SRBWEpiC6_0),.clk(gclk));
	jdff dff_A_JN3xHNET9_0(.dout(w_dff_A_7iVXD8Sp4_0),.din(w_dff_A_JN3xHNET9_0),.clk(gclk));
	jdff dff_A_7iVXD8Sp4_0(.dout(w_dff_A_OUTL29Vo9_0),.din(w_dff_A_7iVXD8Sp4_0),.clk(gclk));
	jdff dff_A_OUTL29Vo9_0(.dout(w_dff_A_eXcYIxyU9_0),.din(w_dff_A_OUTL29Vo9_0),.clk(gclk));
	jdff dff_A_eXcYIxyU9_0(.dout(w_dff_A_fuT2LR7C2_0),.din(w_dff_A_eXcYIxyU9_0),.clk(gclk));
	jdff dff_A_fuT2LR7C2_0(.dout(w_dff_A_bibjArTY6_0),.din(w_dff_A_fuT2LR7C2_0),.clk(gclk));
	jdff dff_A_bibjArTY6_0(.dout(w_dff_A_aEm5TNCV5_0),.din(w_dff_A_bibjArTY6_0),.clk(gclk));
	jdff dff_A_aEm5TNCV5_0(.dout(w_dff_A_6X0Hkh105_0),.din(w_dff_A_aEm5TNCV5_0),.clk(gclk));
	jdff dff_A_6X0Hkh105_0(.dout(w_dff_A_LxsGgTfI2_0),.din(w_dff_A_6X0Hkh105_0),.clk(gclk));
	jdff dff_A_LxsGgTfI2_0(.dout(w_dff_A_RUjfs1g04_0),.din(w_dff_A_LxsGgTfI2_0),.clk(gclk));
	jdff dff_A_RUjfs1g04_0(.dout(w_dff_A_5frHibc22_0),.din(w_dff_A_RUjfs1g04_0),.clk(gclk));
	jdff dff_A_5frHibc22_0(.dout(w_dff_A_Lx6Rpnzz6_0),.din(w_dff_A_5frHibc22_0),.clk(gclk));
	jdff dff_A_Lx6Rpnzz6_0(.dout(w_dff_A_j8yhVrs60_0),.din(w_dff_A_Lx6Rpnzz6_0),.clk(gclk));
	jdff dff_A_j8yhVrs60_0(.dout(w_dff_A_FBuJaati5_0),.din(w_dff_A_j8yhVrs60_0),.clk(gclk));
	jdff dff_A_FBuJaati5_0(.dout(w_dff_A_0njTq2o26_0),.din(w_dff_A_FBuJaati5_0),.clk(gclk));
	jdff dff_A_0njTq2o26_0(.dout(w_dff_A_0k8lcele9_0),.din(w_dff_A_0njTq2o26_0),.clk(gclk));
	jdff dff_A_0k8lcele9_0(.dout(w_dff_A_I2mqRNHs6_0),.din(w_dff_A_0k8lcele9_0),.clk(gclk));
	jdff dff_A_I2mqRNHs6_0(.dout(w_dff_A_cM7FXky90_0),.din(w_dff_A_I2mqRNHs6_0),.clk(gclk));
	jdff dff_A_cM7FXky90_0(.dout(w_dff_A_ndKk4ywE9_0),.din(w_dff_A_cM7FXky90_0),.clk(gclk));
	jdff dff_A_ndKk4ywE9_0(.dout(w_dff_A_rFyx1reS0_0),.din(w_dff_A_ndKk4ywE9_0),.clk(gclk));
	jdff dff_A_rFyx1reS0_0(.dout(w_dff_A_N3nbda6R0_0),.din(w_dff_A_rFyx1reS0_0),.clk(gclk));
	jdff dff_A_N3nbda6R0_0(.dout(w_dff_A_BwdpbHXw3_0),.din(w_dff_A_N3nbda6R0_0),.clk(gclk));
	jdff dff_A_BwdpbHXw3_0(.dout(w_dff_A_GIkqeymX2_0),.din(w_dff_A_BwdpbHXw3_0),.clk(gclk));
	jdff dff_A_GIkqeymX2_0(.dout(w_dff_A_GC9J6uZz8_0),.din(w_dff_A_GIkqeymX2_0),.clk(gclk));
	jdff dff_A_GC9J6uZz8_0(.dout(w_dff_A_ZVpwNGuK0_0),.din(w_dff_A_GC9J6uZz8_0),.clk(gclk));
	jdff dff_A_ZVpwNGuK0_0(.dout(w_dff_A_MFiTvBbX4_0),.din(w_dff_A_ZVpwNGuK0_0),.clk(gclk));
	jdff dff_A_MFiTvBbX4_0(.dout(w_dff_A_MaHDXhzZ9_0),.din(w_dff_A_MFiTvBbX4_0),.clk(gclk));
	jdff dff_A_MaHDXhzZ9_0(.dout(w_dff_A_sDLdcoCN1_0),.din(w_dff_A_MaHDXhzZ9_0),.clk(gclk));
	jdff dff_A_sDLdcoCN1_0(.dout(w_dff_A_dOPFCIKj0_0),.din(w_dff_A_sDLdcoCN1_0),.clk(gclk));
	jdff dff_A_dOPFCIKj0_0(.dout(w_dff_A_dngdOybR0_0),.din(w_dff_A_dOPFCIKj0_0),.clk(gclk));
	jdff dff_A_dngdOybR0_0(.dout(w_dff_A_HYouyW4f7_0),.din(w_dff_A_dngdOybR0_0),.clk(gclk));
	jdff dff_A_HYouyW4f7_0(.dout(w_dff_A_P4px86Pf8_0),.din(w_dff_A_HYouyW4f7_0),.clk(gclk));
	jdff dff_A_P4px86Pf8_0(.dout(w_dff_A_6Gs0xb4l6_0),.din(w_dff_A_P4px86Pf8_0),.clk(gclk));
	jdff dff_A_6Gs0xb4l6_0(.dout(w_dff_A_fxvU3Dhu5_0),.din(w_dff_A_6Gs0xb4l6_0),.clk(gclk));
	jdff dff_A_fxvU3Dhu5_0(.dout(w_dff_A_0mg0BSQh3_0),.din(w_dff_A_fxvU3Dhu5_0),.clk(gclk));
	jdff dff_A_0mg0BSQh3_0(.dout(w_dff_A_QzLDgINi9_0),.din(w_dff_A_0mg0BSQh3_0),.clk(gclk));
	jdff dff_A_QzLDgINi9_0(.dout(w_dff_A_Zf4DBYiT4_0),.din(w_dff_A_QzLDgINi9_0),.clk(gclk));
	jdff dff_A_Zf4DBYiT4_0(.dout(w_dff_A_TsWhlDO92_0),.din(w_dff_A_Zf4DBYiT4_0),.clk(gclk));
	jdff dff_A_TsWhlDO92_0(.dout(w_dff_A_6nk7GkCt1_0),.din(w_dff_A_TsWhlDO92_0),.clk(gclk));
	jdff dff_A_6nk7GkCt1_0(.dout(G4946gat),.din(w_dff_A_6nk7GkCt1_0),.clk(gclk));
	jdff dff_A_8K6sinQo2_2(.dout(w_dff_A_GfPQn7GX3_0),.din(w_dff_A_8K6sinQo2_2),.clk(gclk));
	jdff dff_A_GfPQn7GX3_0(.dout(w_dff_A_JNnXggAV3_0),.din(w_dff_A_GfPQn7GX3_0),.clk(gclk));
	jdff dff_A_JNnXggAV3_0(.dout(w_dff_A_RXF1Y7ws6_0),.din(w_dff_A_JNnXggAV3_0),.clk(gclk));
	jdff dff_A_RXF1Y7ws6_0(.dout(w_dff_A_ofXrKFV59_0),.din(w_dff_A_RXF1Y7ws6_0),.clk(gclk));
	jdff dff_A_ofXrKFV59_0(.dout(w_dff_A_f4fQlerU7_0),.din(w_dff_A_ofXrKFV59_0),.clk(gclk));
	jdff dff_A_f4fQlerU7_0(.dout(w_dff_A_1fN5ouJP5_0),.din(w_dff_A_f4fQlerU7_0),.clk(gclk));
	jdff dff_A_1fN5ouJP5_0(.dout(w_dff_A_zU7Jeund6_0),.din(w_dff_A_1fN5ouJP5_0),.clk(gclk));
	jdff dff_A_zU7Jeund6_0(.dout(w_dff_A_DdzN2HBs7_0),.din(w_dff_A_zU7Jeund6_0),.clk(gclk));
	jdff dff_A_DdzN2HBs7_0(.dout(w_dff_A_M7zlZhe93_0),.din(w_dff_A_DdzN2HBs7_0),.clk(gclk));
	jdff dff_A_M7zlZhe93_0(.dout(w_dff_A_yssQJ5ap2_0),.din(w_dff_A_M7zlZhe93_0),.clk(gclk));
	jdff dff_A_yssQJ5ap2_0(.dout(w_dff_A_A7J1Gk0G7_0),.din(w_dff_A_yssQJ5ap2_0),.clk(gclk));
	jdff dff_A_A7J1Gk0G7_0(.dout(w_dff_A_Dw9LjXUF7_0),.din(w_dff_A_A7J1Gk0G7_0),.clk(gclk));
	jdff dff_A_Dw9LjXUF7_0(.dout(w_dff_A_lyw1ITQV8_0),.din(w_dff_A_Dw9LjXUF7_0),.clk(gclk));
	jdff dff_A_lyw1ITQV8_0(.dout(w_dff_A_kWwfDxtK4_0),.din(w_dff_A_lyw1ITQV8_0),.clk(gclk));
	jdff dff_A_kWwfDxtK4_0(.dout(w_dff_A_cCr8Tswj7_0),.din(w_dff_A_kWwfDxtK4_0),.clk(gclk));
	jdff dff_A_cCr8Tswj7_0(.dout(w_dff_A_nFgjYuYT0_0),.din(w_dff_A_cCr8Tswj7_0),.clk(gclk));
	jdff dff_A_nFgjYuYT0_0(.dout(w_dff_A_plHmViy87_0),.din(w_dff_A_nFgjYuYT0_0),.clk(gclk));
	jdff dff_A_plHmViy87_0(.dout(w_dff_A_BR26NNCS8_0),.din(w_dff_A_plHmViy87_0),.clk(gclk));
	jdff dff_A_BR26NNCS8_0(.dout(w_dff_A_7gPHeTGa1_0),.din(w_dff_A_BR26NNCS8_0),.clk(gclk));
	jdff dff_A_7gPHeTGa1_0(.dout(w_dff_A_WiaY6IOK6_0),.din(w_dff_A_7gPHeTGa1_0),.clk(gclk));
	jdff dff_A_WiaY6IOK6_0(.dout(w_dff_A_Vo80r9JR8_0),.din(w_dff_A_WiaY6IOK6_0),.clk(gclk));
	jdff dff_A_Vo80r9JR8_0(.dout(w_dff_A_SpoRhbOs9_0),.din(w_dff_A_Vo80r9JR8_0),.clk(gclk));
	jdff dff_A_SpoRhbOs9_0(.dout(w_dff_A_sgO7idng4_0),.din(w_dff_A_SpoRhbOs9_0),.clk(gclk));
	jdff dff_A_sgO7idng4_0(.dout(w_dff_A_SMpKunVy7_0),.din(w_dff_A_sgO7idng4_0),.clk(gclk));
	jdff dff_A_SMpKunVy7_0(.dout(w_dff_A_JurrIsLZ7_0),.din(w_dff_A_SMpKunVy7_0),.clk(gclk));
	jdff dff_A_JurrIsLZ7_0(.dout(w_dff_A_jYyqzmar3_0),.din(w_dff_A_JurrIsLZ7_0),.clk(gclk));
	jdff dff_A_jYyqzmar3_0(.dout(w_dff_A_jqO2OKA84_0),.din(w_dff_A_jYyqzmar3_0),.clk(gclk));
	jdff dff_A_jqO2OKA84_0(.dout(w_dff_A_XL3D0XrL0_0),.din(w_dff_A_jqO2OKA84_0),.clk(gclk));
	jdff dff_A_XL3D0XrL0_0(.dout(w_dff_A_mzN4nRDF2_0),.din(w_dff_A_XL3D0XrL0_0),.clk(gclk));
	jdff dff_A_mzN4nRDF2_0(.dout(w_dff_A_EQUZUBrn5_0),.din(w_dff_A_mzN4nRDF2_0),.clk(gclk));
	jdff dff_A_EQUZUBrn5_0(.dout(w_dff_A_tYOakAXO1_0),.din(w_dff_A_EQUZUBrn5_0),.clk(gclk));
	jdff dff_A_tYOakAXO1_0(.dout(w_dff_A_KCFnn8lv5_0),.din(w_dff_A_tYOakAXO1_0),.clk(gclk));
	jdff dff_A_KCFnn8lv5_0(.dout(w_dff_A_YGZhVVr04_0),.din(w_dff_A_KCFnn8lv5_0),.clk(gclk));
	jdff dff_A_YGZhVVr04_0(.dout(w_dff_A_jtk7yuY95_0),.din(w_dff_A_YGZhVVr04_0),.clk(gclk));
	jdff dff_A_jtk7yuY95_0(.dout(w_dff_A_R3asqZOm8_0),.din(w_dff_A_jtk7yuY95_0),.clk(gclk));
	jdff dff_A_R3asqZOm8_0(.dout(w_dff_A_KAtYWEx24_0),.din(w_dff_A_R3asqZOm8_0),.clk(gclk));
	jdff dff_A_KAtYWEx24_0(.dout(w_dff_A_xAs5my3L6_0),.din(w_dff_A_KAtYWEx24_0),.clk(gclk));
	jdff dff_A_xAs5my3L6_0(.dout(w_dff_A_TkAKGVbx0_0),.din(w_dff_A_xAs5my3L6_0),.clk(gclk));
	jdff dff_A_TkAKGVbx0_0(.dout(G5308gat),.din(w_dff_A_TkAKGVbx0_0),.clk(gclk));
	jdff dff_A_bgSyLykw2_2(.dout(w_dff_A_ntCRt9Xm2_0),.din(w_dff_A_bgSyLykw2_2),.clk(gclk));
	jdff dff_A_ntCRt9Xm2_0(.dout(w_dff_A_Sgrhl8zQ8_0),.din(w_dff_A_ntCRt9Xm2_0),.clk(gclk));
	jdff dff_A_Sgrhl8zQ8_0(.dout(w_dff_A_ZePkzJr66_0),.din(w_dff_A_Sgrhl8zQ8_0),.clk(gclk));
	jdff dff_A_ZePkzJr66_0(.dout(w_dff_A_dhwgM6kh5_0),.din(w_dff_A_ZePkzJr66_0),.clk(gclk));
	jdff dff_A_dhwgM6kh5_0(.dout(w_dff_A_BoEvaWQw6_0),.din(w_dff_A_dhwgM6kh5_0),.clk(gclk));
	jdff dff_A_BoEvaWQw6_0(.dout(w_dff_A_pGVXO9u82_0),.din(w_dff_A_BoEvaWQw6_0),.clk(gclk));
	jdff dff_A_pGVXO9u82_0(.dout(w_dff_A_VJPXJRPA5_0),.din(w_dff_A_pGVXO9u82_0),.clk(gclk));
	jdff dff_A_VJPXJRPA5_0(.dout(w_dff_A_7kCwRQcM5_0),.din(w_dff_A_VJPXJRPA5_0),.clk(gclk));
	jdff dff_A_7kCwRQcM5_0(.dout(w_dff_A_Kxs5Dtx22_0),.din(w_dff_A_7kCwRQcM5_0),.clk(gclk));
	jdff dff_A_Kxs5Dtx22_0(.dout(w_dff_A_6aNgm7qc6_0),.din(w_dff_A_Kxs5Dtx22_0),.clk(gclk));
	jdff dff_A_6aNgm7qc6_0(.dout(w_dff_A_1my3cUMa0_0),.din(w_dff_A_6aNgm7qc6_0),.clk(gclk));
	jdff dff_A_1my3cUMa0_0(.dout(w_dff_A_iVHRFBGG3_0),.din(w_dff_A_1my3cUMa0_0),.clk(gclk));
	jdff dff_A_iVHRFBGG3_0(.dout(w_dff_A_rU7hAwhA0_0),.din(w_dff_A_iVHRFBGG3_0),.clk(gclk));
	jdff dff_A_rU7hAwhA0_0(.dout(w_dff_A_me30UN9W4_0),.din(w_dff_A_rU7hAwhA0_0),.clk(gclk));
	jdff dff_A_me30UN9W4_0(.dout(w_dff_A_ShzFT1zM2_0),.din(w_dff_A_me30UN9W4_0),.clk(gclk));
	jdff dff_A_ShzFT1zM2_0(.dout(w_dff_A_ZTjzSqwx2_0),.din(w_dff_A_ShzFT1zM2_0),.clk(gclk));
	jdff dff_A_ZTjzSqwx2_0(.dout(w_dff_A_3U7yrEdy9_0),.din(w_dff_A_ZTjzSqwx2_0),.clk(gclk));
	jdff dff_A_3U7yrEdy9_0(.dout(w_dff_A_0ATY7b6R9_0),.din(w_dff_A_3U7yrEdy9_0),.clk(gclk));
	jdff dff_A_0ATY7b6R9_0(.dout(w_dff_A_WwRyUwzb2_0),.din(w_dff_A_0ATY7b6R9_0),.clk(gclk));
	jdff dff_A_WwRyUwzb2_0(.dout(w_dff_A_hYAG7MK33_0),.din(w_dff_A_WwRyUwzb2_0),.clk(gclk));
	jdff dff_A_hYAG7MK33_0(.dout(w_dff_A_SDJMsobg9_0),.din(w_dff_A_hYAG7MK33_0),.clk(gclk));
	jdff dff_A_SDJMsobg9_0(.dout(w_dff_A_fSOs6jWy6_0),.din(w_dff_A_SDJMsobg9_0),.clk(gclk));
	jdff dff_A_fSOs6jWy6_0(.dout(w_dff_A_DczPKTpz3_0),.din(w_dff_A_fSOs6jWy6_0),.clk(gclk));
	jdff dff_A_DczPKTpz3_0(.dout(w_dff_A_kCL466yC7_0),.din(w_dff_A_DczPKTpz3_0),.clk(gclk));
	jdff dff_A_kCL466yC7_0(.dout(w_dff_A_H7OGRi6A5_0),.din(w_dff_A_kCL466yC7_0),.clk(gclk));
	jdff dff_A_H7OGRi6A5_0(.dout(w_dff_A_bnWgRYoh5_0),.din(w_dff_A_H7OGRi6A5_0),.clk(gclk));
	jdff dff_A_bnWgRYoh5_0(.dout(w_dff_A_YS7a8fLk6_0),.din(w_dff_A_bnWgRYoh5_0),.clk(gclk));
	jdff dff_A_YS7a8fLk6_0(.dout(w_dff_A_LmWMfktV1_0),.din(w_dff_A_YS7a8fLk6_0),.clk(gclk));
	jdff dff_A_LmWMfktV1_0(.dout(w_dff_A_lwv9BZYb9_0),.din(w_dff_A_LmWMfktV1_0),.clk(gclk));
	jdff dff_A_lwv9BZYb9_0(.dout(w_dff_A_tSjzfsgx4_0),.din(w_dff_A_lwv9BZYb9_0),.clk(gclk));
	jdff dff_A_tSjzfsgx4_0(.dout(w_dff_A_u8VmXTca9_0),.din(w_dff_A_tSjzfsgx4_0),.clk(gclk));
	jdff dff_A_u8VmXTca9_0(.dout(w_dff_A_oojI1ZYQ6_0),.din(w_dff_A_u8VmXTca9_0),.clk(gclk));
	jdff dff_A_oojI1ZYQ6_0(.dout(w_dff_A_oIIRsrEb9_0),.din(w_dff_A_oojI1ZYQ6_0),.clk(gclk));
	jdff dff_A_oIIRsrEb9_0(.dout(w_dff_A_OpzbgR6U0_0),.din(w_dff_A_oIIRsrEb9_0),.clk(gclk));
	jdff dff_A_OpzbgR6U0_0(.dout(w_dff_A_XgOMPC0j8_0),.din(w_dff_A_OpzbgR6U0_0),.clk(gclk));
	jdff dff_A_XgOMPC0j8_0(.dout(G5672gat),.din(w_dff_A_XgOMPC0j8_0),.clk(gclk));
	jdff dff_A_HUPrWpUI2_2(.dout(w_dff_A_64QSWXVK6_0),.din(w_dff_A_HUPrWpUI2_2),.clk(gclk));
	jdff dff_A_64QSWXVK6_0(.dout(w_dff_A_PFHLJvTo9_0),.din(w_dff_A_64QSWXVK6_0),.clk(gclk));
	jdff dff_A_PFHLJvTo9_0(.dout(w_dff_A_pZdJIG9B4_0),.din(w_dff_A_PFHLJvTo9_0),.clk(gclk));
	jdff dff_A_pZdJIG9B4_0(.dout(w_dff_A_9LDmQsRC7_0),.din(w_dff_A_pZdJIG9B4_0),.clk(gclk));
	jdff dff_A_9LDmQsRC7_0(.dout(w_dff_A_bWPyAhAK8_0),.din(w_dff_A_9LDmQsRC7_0),.clk(gclk));
	jdff dff_A_bWPyAhAK8_0(.dout(w_dff_A_CEfgBgMP8_0),.din(w_dff_A_bWPyAhAK8_0),.clk(gclk));
	jdff dff_A_CEfgBgMP8_0(.dout(w_dff_A_HaxRrwB50_0),.din(w_dff_A_CEfgBgMP8_0),.clk(gclk));
	jdff dff_A_HaxRrwB50_0(.dout(w_dff_A_WYz39Sl44_0),.din(w_dff_A_HaxRrwB50_0),.clk(gclk));
	jdff dff_A_WYz39Sl44_0(.dout(w_dff_A_Ju5LJsON5_0),.din(w_dff_A_WYz39Sl44_0),.clk(gclk));
	jdff dff_A_Ju5LJsON5_0(.dout(w_dff_A_5IYbzKHa0_0),.din(w_dff_A_Ju5LJsON5_0),.clk(gclk));
	jdff dff_A_5IYbzKHa0_0(.dout(w_dff_A_FhudYR129_0),.din(w_dff_A_5IYbzKHa0_0),.clk(gclk));
	jdff dff_A_FhudYR129_0(.dout(w_dff_A_WQMPsREa2_0),.din(w_dff_A_FhudYR129_0),.clk(gclk));
	jdff dff_A_WQMPsREa2_0(.dout(w_dff_A_DcRdYJQx1_0),.din(w_dff_A_WQMPsREa2_0),.clk(gclk));
	jdff dff_A_DcRdYJQx1_0(.dout(w_dff_A_3NVsXQ8R2_0),.din(w_dff_A_DcRdYJQx1_0),.clk(gclk));
	jdff dff_A_3NVsXQ8R2_0(.dout(w_dff_A_I8O7RJY53_0),.din(w_dff_A_3NVsXQ8R2_0),.clk(gclk));
	jdff dff_A_I8O7RJY53_0(.dout(w_dff_A_gEj68g6m7_0),.din(w_dff_A_I8O7RJY53_0),.clk(gclk));
	jdff dff_A_gEj68g6m7_0(.dout(w_dff_A_Rj970DGQ4_0),.din(w_dff_A_gEj68g6m7_0),.clk(gclk));
	jdff dff_A_Rj970DGQ4_0(.dout(w_dff_A_JXVDUVx24_0),.din(w_dff_A_Rj970DGQ4_0),.clk(gclk));
	jdff dff_A_JXVDUVx24_0(.dout(w_dff_A_ub5KuGH98_0),.din(w_dff_A_JXVDUVx24_0),.clk(gclk));
	jdff dff_A_ub5KuGH98_0(.dout(w_dff_A_PXFymSUC6_0),.din(w_dff_A_ub5KuGH98_0),.clk(gclk));
	jdff dff_A_PXFymSUC6_0(.dout(w_dff_A_9AAylEAF5_0),.din(w_dff_A_PXFymSUC6_0),.clk(gclk));
	jdff dff_A_9AAylEAF5_0(.dout(w_dff_A_bKlsDN5c9_0),.din(w_dff_A_9AAylEAF5_0),.clk(gclk));
	jdff dff_A_bKlsDN5c9_0(.dout(w_dff_A_tkELLfEE5_0),.din(w_dff_A_bKlsDN5c9_0),.clk(gclk));
	jdff dff_A_tkELLfEE5_0(.dout(w_dff_A_FuWYUGHm4_0),.din(w_dff_A_tkELLfEE5_0),.clk(gclk));
	jdff dff_A_FuWYUGHm4_0(.dout(w_dff_A_EgKCktUe0_0),.din(w_dff_A_FuWYUGHm4_0),.clk(gclk));
	jdff dff_A_EgKCktUe0_0(.dout(w_dff_A_HOOPbwb98_0),.din(w_dff_A_EgKCktUe0_0),.clk(gclk));
	jdff dff_A_HOOPbwb98_0(.dout(w_dff_A_KuElOmoQ7_0),.din(w_dff_A_HOOPbwb98_0),.clk(gclk));
	jdff dff_A_KuElOmoQ7_0(.dout(w_dff_A_Eb4f4YI32_0),.din(w_dff_A_KuElOmoQ7_0),.clk(gclk));
	jdff dff_A_Eb4f4YI32_0(.dout(w_dff_A_Y9VpNMDr4_0),.din(w_dff_A_Eb4f4YI32_0),.clk(gclk));
	jdff dff_A_Y9VpNMDr4_0(.dout(w_dff_A_Az6wZtah5_0),.din(w_dff_A_Y9VpNMDr4_0),.clk(gclk));
	jdff dff_A_Az6wZtah5_0(.dout(w_dff_A_DseTCSk85_0),.din(w_dff_A_Az6wZtah5_0),.clk(gclk));
	jdff dff_A_DseTCSk85_0(.dout(w_dff_A_CC5pY0xT4_0),.din(w_dff_A_DseTCSk85_0),.clk(gclk));
	jdff dff_A_CC5pY0xT4_0(.dout(G5971gat),.din(w_dff_A_CC5pY0xT4_0),.clk(gclk));
	jdff dff_A_dkRXDqWE6_2(.dout(w_dff_A_yiZ3IYnb0_0),.din(w_dff_A_dkRXDqWE6_2),.clk(gclk));
	jdff dff_A_yiZ3IYnb0_0(.dout(w_dff_A_GRbEqwlc5_0),.din(w_dff_A_yiZ3IYnb0_0),.clk(gclk));
	jdff dff_A_GRbEqwlc5_0(.dout(w_dff_A_yNueZH6b5_0),.din(w_dff_A_GRbEqwlc5_0),.clk(gclk));
	jdff dff_A_yNueZH6b5_0(.dout(w_dff_A_9aGsA8D06_0),.din(w_dff_A_yNueZH6b5_0),.clk(gclk));
	jdff dff_A_9aGsA8D06_0(.dout(w_dff_A_G5bZRDvy3_0),.din(w_dff_A_9aGsA8D06_0),.clk(gclk));
	jdff dff_A_G5bZRDvy3_0(.dout(w_dff_A_SW2Ij6fh7_0),.din(w_dff_A_G5bZRDvy3_0),.clk(gclk));
	jdff dff_A_SW2Ij6fh7_0(.dout(w_dff_A_Wqyn8iDX4_0),.din(w_dff_A_SW2Ij6fh7_0),.clk(gclk));
	jdff dff_A_Wqyn8iDX4_0(.dout(w_dff_A_A9O1UhMb5_0),.din(w_dff_A_Wqyn8iDX4_0),.clk(gclk));
	jdff dff_A_A9O1UhMb5_0(.dout(w_dff_A_jgzE7U3v1_0),.din(w_dff_A_A9O1UhMb5_0),.clk(gclk));
	jdff dff_A_jgzE7U3v1_0(.dout(w_dff_A_RRDgoQ4P2_0),.din(w_dff_A_jgzE7U3v1_0),.clk(gclk));
	jdff dff_A_RRDgoQ4P2_0(.dout(w_dff_A_JO6bXnkI9_0),.din(w_dff_A_RRDgoQ4P2_0),.clk(gclk));
	jdff dff_A_JO6bXnkI9_0(.dout(w_dff_A_4qBoBvWY9_0),.din(w_dff_A_JO6bXnkI9_0),.clk(gclk));
	jdff dff_A_4qBoBvWY9_0(.dout(w_dff_A_mOp6pj7s1_0),.din(w_dff_A_4qBoBvWY9_0),.clk(gclk));
	jdff dff_A_mOp6pj7s1_0(.dout(w_dff_A_DFjpI4MN9_0),.din(w_dff_A_mOp6pj7s1_0),.clk(gclk));
	jdff dff_A_DFjpI4MN9_0(.dout(w_dff_A_H81wNIv47_0),.din(w_dff_A_DFjpI4MN9_0),.clk(gclk));
	jdff dff_A_H81wNIv47_0(.dout(w_dff_A_cRG8EHzL2_0),.din(w_dff_A_H81wNIv47_0),.clk(gclk));
	jdff dff_A_cRG8EHzL2_0(.dout(w_dff_A_QTKL9rY99_0),.din(w_dff_A_cRG8EHzL2_0),.clk(gclk));
	jdff dff_A_QTKL9rY99_0(.dout(w_dff_A_adSknmPh5_0),.din(w_dff_A_QTKL9rY99_0),.clk(gclk));
	jdff dff_A_adSknmPh5_0(.dout(w_dff_A_Hzp84igx3_0),.din(w_dff_A_adSknmPh5_0),.clk(gclk));
	jdff dff_A_Hzp84igx3_0(.dout(w_dff_A_TQiCZPPG1_0),.din(w_dff_A_Hzp84igx3_0),.clk(gclk));
	jdff dff_A_TQiCZPPG1_0(.dout(w_dff_A_7CdSWMpS2_0),.din(w_dff_A_TQiCZPPG1_0),.clk(gclk));
	jdff dff_A_7CdSWMpS2_0(.dout(w_dff_A_nMYswItO5_0),.din(w_dff_A_7CdSWMpS2_0),.clk(gclk));
	jdff dff_A_nMYswItO5_0(.dout(w_dff_A_kDn3tEb55_0),.din(w_dff_A_nMYswItO5_0),.clk(gclk));
	jdff dff_A_kDn3tEb55_0(.dout(w_dff_A_hIceY3HB1_0),.din(w_dff_A_kDn3tEb55_0),.clk(gclk));
	jdff dff_A_hIceY3HB1_0(.dout(w_dff_A_Bt7icd6K9_0),.din(w_dff_A_hIceY3HB1_0),.clk(gclk));
	jdff dff_A_Bt7icd6K9_0(.dout(w_dff_A_K8uXSM0B5_0),.din(w_dff_A_Bt7icd6K9_0),.clk(gclk));
	jdff dff_A_K8uXSM0B5_0(.dout(w_dff_A_R5A5ubKE6_0),.din(w_dff_A_K8uXSM0B5_0),.clk(gclk));
	jdff dff_A_R5A5ubKE6_0(.dout(w_dff_A_rIj6fq011_0),.din(w_dff_A_R5A5ubKE6_0),.clk(gclk));
	jdff dff_A_rIj6fq011_0(.dout(w_dff_A_ukbNP34h2_0),.din(w_dff_A_rIj6fq011_0),.clk(gclk));
	jdff dff_A_ukbNP34h2_0(.dout(G6123gat),.din(w_dff_A_ukbNP34h2_0),.clk(gclk));
	jdff dff_A_XP7KI9S09_2(.dout(w_dff_A_QYT2rliR4_0),.din(w_dff_A_XP7KI9S09_2),.clk(gclk));
	jdff dff_A_QYT2rliR4_0(.dout(w_dff_A_N9SMenpp5_0),.din(w_dff_A_QYT2rliR4_0),.clk(gclk));
	jdff dff_A_N9SMenpp5_0(.dout(w_dff_A_UgK9U5FT0_0),.din(w_dff_A_N9SMenpp5_0),.clk(gclk));
	jdff dff_A_UgK9U5FT0_0(.dout(w_dff_A_7PBadlrA1_0),.din(w_dff_A_UgK9U5FT0_0),.clk(gclk));
	jdff dff_A_7PBadlrA1_0(.dout(w_dff_A_y2udl6fQ1_0),.din(w_dff_A_7PBadlrA1_0),.clk(gclk));
	jdff dff_A_y2udl6fQ1_0(.dout(w_dff_A_oVl7XIuV5_0),.din(w_dff_A_y2udl6fQ1_0),.clk(gclk));
	jdff dff_A_oVl7XIuV5_0(.dout(w_dff_A_7ZQ1NyRU9_0),.din(w_dff_A_oVl7XIuV5_0),.clk(gclk));
	jdff dff_A_7ZQ1NyRU9_0(.dout(w_dff_A_HoujgT4A7_0),.din(w_dff_A_7ZQ1NyRU9_0),.clk(gclk));
	jdff dff_A_HoujgT4A7_0(.dout(w_dff_A_mIL9qtZM0_0),.din(w_dff_A_HoujgT4A7_0),.clk(gclk));
	jdff dff_A_mIL9qtZM0_0(.dout(w_dff_A_SxwH9dxH1_0),.din(w_dff_A_mIL9qtZM0_0),.clk(gclk));
	jdff dff_A_SxwH9dxH1_0(.dout(w_dff_A_35805j6E7_0),.din(w_dff_A_SxwH9dxH1_0),.clk(gclk));
	jdff dff_A_35805j6E7_0(.dout(w_dff_A_6aAhYsJY9_0),.din(w_dff_A_35805j6E7_0),.clk(gclk));
	jdff dff_A_6aAhYsJY9_0(.dout(w_dff_A_LVMOG8c84_0),.din(w_dff_A_6aAhYsJY9_0),.clk(gclk));
	jdff dff_A_LVMOG8c84_0(.dout(w_dff_A_asFbVqi07_0),.din(w_dff_A_LVMOG8c84_0),.clk(gclk));
	jdff dff_A_asFbVqi07_0(.dout(w_dff_A_OwHt3ajN5_0),.din(w_dff_A_asFbVqi07_0),.clk(gclk));
	jdff dff_A_OwHt3ajN5_0(.dout(w_dff_A_8bxLa27V0_0),.din(w_dff_A_OwHt3ajN5_0),.clk(gclk));
	jdff dff_A_8bxLa27V0_0(.dout(w_dff_A_0w5p6SzL5_0),.din(w_dff_A_8bxLa27V0_0),.clk(gclk));
	jdff dff_A_0w5p6SzL5_0(.dout(w_dff_A_G2RhsFcW6_0),.din(w_dff_A_0w5p6SzL5_0),.clk(gclk));
	jdff dff_A_G2RhsFcW6_0(.dout(w_dff_A_h6gZP8qM5_0),.din(w_dff_A_G2RhsFcW6_0),.clk(gclk));
	jdff dff_A_h6gZP8qM5_0(.dout(w_dff_A_UtcDfwkz2_0),.din(w_dff_A_h6gZP8qM5_0),.clk(gclk));
	jdff dff_A_UtcDfwkz2_0(.dout(w_dff_A_SKWDjgK36_0),.din(w_dff_A_UtcDfwkz2_0),.clk(gclk));
	jdff dff_A_SKWDjgK36_0(.dout(w_dff_A_lsoqaHTn7_0),.din(w_dff_A_SKWDjgK36_0),.clk(gclk));
	jdff dff_A_lsoqaHTn7_0(.dout(w_dff_A_n4q0mMOi0_0),.din(w_dff_A_lsoqaHTn7_0),.clk(gclk));
	jdff dff_A_n4q0mMOi0_0(.dout(w_dff_A_quTNwDxI6_0),.din(w_dff_A_n4q0mMOi0_0),.clk(gclk));
	jdff dff_A_quTNwDxI6_0(.dout(w_dff_A_rZolB5tP1_0),.din(w_dff_A_quTNwDxI6_0),.clk(gclk));
	jdff dff_A_rZolB5tP1_0(.dout(w_dff_A_5z3SpYsC8_0),.din(w_dff_A_rZolB5tP1_0),.clk(gclk));
	jdff dff_A_5z3SpYsC8_0(.dout(w_dff_A_L2Nd2Iat2_0),.din(w_dff_A_5z3SpYsC8_0),.clk(gclk));
	jdff dff_A_L2Nd2Iat2_0(.dout(G6150gat),.din(w_dff_A_L2Nd2Iat2_0),.clk(gclk));
	jdff dff_A_muYCmXs49_2(.dout(w_dff_A_RhmMgHzJ2_0),.din(w_dff_A_muYCmXs49_2),.clk(gclk));
	jdff dff_A_RhmMgHzJ2_0(.dout(w_dff_A_Y1oVLQD46_0),.din(w_dff_A_RhmMgHzJ2_0),.clk(gclk));
	jdff dff_A_Y1oVLQD46_0(.dout(w_dff_A_xdwiQXY37_0),.din(w_dff_A_Y1oVLQD46_0),.clk(gclk));
	jdff dff_A_xdwiQXY37_0(.dout(w_dff_A_PkRSJyfj3_0),.din(w_dff_A_xdwiQXY37_0),.clk(gclk));
	jdff dff_A_PkRSJyfj3_0(.dout(w_dff_A_4gLnuB6Z8_0),.din(w_dff_A_PkRSJyfj3_0),.clk(gclk));
	jdff dff_A_4gLnuB6Z8_0(.dout(w_dff_A_asP64sgb1_0),.din(w_dff_A_4gLnuB6Z8_0),.clk(gclk));
	jdff dff_A_asP64sgb1_0(.dout(w_dff_A_dByGgPP52_0),.din(w_dff_A_asP64sgb1_0),.clk(gclk));
	jdff dff_A_dByGgPP52_0(.dout(w_dff_A_jDheKlDP8_0),.din(w_dff_A_dByGgPP52_0),.clk(gclk));
	jdff dff_A_jDheKlDP8_0(.dout(w_dff_A_pWlC6zdb2_0),.din(w_dff_A_jDheKlDP8_0),.clk(gclk));
	jdff dff_A_pWlC6zdb2_0(.dout(w_dff_A_uehCxuEK1_0),.din(w_dff_A_pWlC6zdb2_0),.clk(gclk));
	jdff dff_A_uehCxuEK1_0(.dout(w_dff_A_DYt4QheT0_0),.din(w_dff_A_uehCxuEK1_0),.clk(gclk));
	jdff dff_A_DYt4QheT0_0(.dout(w_dff_A_aGaicp3P0_0),.din(w_dff_A_DYt4QheT0_0),.clk(gclk));
	jdff dff_A_aGaicp3P0_0(.dout(w_dff_A_1i05DgVs6_0),.din(w_dff_A_aGaicp3P0_0),.clk(gclk));
	jdff dff_A_1i05DgVs6_0(.dout(w_dff_A_2stMxxT16_0),.din(w_dff_A_1i05DgVs6_0),.clk(gclk));
	jdff dff_A_2stMxxT16_0(.dout(w_dff_A_5YBeaBvd9_0),.din(w_dff_A_2stMxxT16_0),.clk(gclk));
	jdff dff_A_5YBeaBvd9_0(.dout(w_dff_A_KDw3NH4l1_0),.din(w_dff_A_5YBeaBvd9_0),.clk(gclk));
	jdff dff_A_KDw3NH4l1_0(.dout(w_dff_A_lEuD209Z0_0),.din(w_dff_A_KDw3NH4l1_0),.clk(gclk));
	jdff dff_A_lEuD209Z0_0(.dout(w_dff_A_mir0XGtj0_0),.din(w_dff_A_lEuD209Z0_0),.clk(gclk));
	jdff dff_A_mir0XGtj0_0(.dout(w_dff_A_Jj3fJt1g0_0),.din(w_dff_A_mir0XGtj0_0),.clk(gclk));
	jdff dff_A_Jj3fJt1g0_0(.dout(w_dff_A_kpQ2LYBI7_0),.din(w_dff_A_Jj3fJt1g0_0),.clk(gclk));
	jdff dff_A_kpQ2LYBI7_0(.dout(w_dff_A_agb1MY1J7_0),.din(w_dff_A_kpQ2LYBI7_0),.clk(gclk));
	jdff dff_A_agb1MY1J7_0(.dout(w_dff_A_yQbmpn760_0),.din(w_dff_A_agb1MY1J7_0),.clk(gclk));
	jdff dff_A_yQbmpn760_0(.dout(w_dff_A_l8Ot5fQK3_0),.din(w_dff_A_yQbmpn760_0),.clk(gclk));
	jdff dff_A_l8Ot5fQK3_0(.dout(w_dff_A_NSXzSIEr5_0),.din(w_dff_A_l8Ot5fQK3_0),.clk(gclk));
	jdff dff_A_NSXzSIEr5_0(.dout(w_dff_A_smKVEayf3_0),.din(w_dff_A_NSXzSIEr5_0),.clk(gclk));
	jdff dff_A_smKVEayf3_0(.dout(G6160gat),.din(w_dff_A_smKVEayf3_0),.clk(gclk));
	jdff dff_A_MsaMqHPq5_2(.dout(w_dff_A_EWidRBpa7_0),.din(w_dff_A_MsaMqHPq5_2),.clk(gclk));
	jdff dff_A_EWidRBpa7_0(.dout(w_dff_A_J3bF2UZ40_0),.din(w_dff_A_EWidRBpa7_0),.clk(gclk));
	jdff dff_A_J3bF2UZ40_0(.dout(w_dff_A_NU4fQv7S1_0),.din(w_dff_A_J3bF2UZ40_0),.clk(gclk));
	jdff dff_A_NU4fQv7S1_0(.dout(w_dff_A_e6F23xlq3_0),.din(w_dff_A_NU4fQv7S1_0),.clk(gclk));
	jdff dff_A_e6F23xlq3_0(.dout(w_dff_A_MR7cQP7V6_0),.din(w_dff_A_e6F23xlq3_0),.clk(gclk));
	jdff dff_A_MR7cQP7V6_0(.dout(w_dff_A_jurMbIww6_0),.din(w_dff_A_MR7cQP7V6_0),.clk(gclk));
	jdff dff_A_jurMbIww6_0(.dout(w_dff_A_RLAmi19d0_0),.din(w_dff_A_jurMbIww6_0),.clk(gclk));
	jdff dff_A_RLAmi19d0_0(.dout(w_dff_A_cY6jLVdC3_0),.din(w_dff_A_RLAmi19d0_0),.clk(gclk));
	jdff dff_A_cY6jLVdC3_0(.dout(w_dff_A_8lanbtLS9_0),.din(w_dff_A_cY6jLVdC3_0),.clk(gclk));
	jdff dff_A_8lanbtLS9_0(.dout(w_dff_A_akO7jPOA8_0),.din(w_dff_A_8lanbtLS9_0),.clk(gclk));
	jdff dff_A_akO7jPOA8_0(.dout(w_dff_A_llQc2Dv85_0),.din(w_dff_A_akO7jPOA8_0),.clk(gclk));
	jdff dff_A_llQc2Dv85_0(.dout(w_dff_A_oLB8ljKD0_0),.din(w_dff_A_llQc2Dv85_0),.clk(gclk));
	jdff dff_A_oLB8ljKD0_0(.dout(w_dff_A_okEQeA9W3_0),.din(w_dff_A_oLB8ljKD0_0),.clk(gclk));
	jdff dff_A_okEQeA9W3_0(.dout(w_dff_A_exmAmJc02_0),.din(w_dff_A_okEQeA9W3_0),.clk(gclk));
	jdff dff_A_exmAmJc02_0(.dout(w_dff_A_NhFTfx3R2_0),.din(w_dff_A_exmAmJc02_0),.clk(gclk));
	jdff dff_A_NhFTfx3R2_0(.dout(w_dff_A_OZiNN5vz2_0),.din(w_dff_A_NhFTfx3R2_0),.clk(gclk));
	jdff dff_A_OZiNN5vz2_0(.dout(w_dff_A_oZf1kPbn0_0),.din(w_dff_A_OZiNN5vz2_0),.clk(gclk));
	jdff dff_A_oZf1kPbn0_0(.dout(w_dff_A_iZqQD9uf0_0),.din(w_dff_A_oZf1kPbn0_0),.clk(gclk));
	jdff dff_A_iZqQD9uf0_0(.dout(w_dff_A_gFb0YsbJ8_0),.din(w_dff_A_iZqQD9uf0_0),.clk(gclk));
	jdff dff_A_gFb0YsbJ8_0(.dout(w_dff_A_EYGGr5a33_0),.din(w_dff_A_gFb0YsbJ8_0),.clk(gclk));
	jdff dff_A_EYGGr5a33_0(.dout(w_dff_A_XyirquLk5_0),.din(w_dff_A_EYGGr5a33_0),.clk(gclk));
	jdff dff_A_XyirquLk5_0(.dout(w_dff_A_4aciwrKU0_0),.din(w_dff_A_XyirquLk5_0),.clk(gclk));
	jdff dff_A_4aciwrKU0_0(.dout(w_dff_A_2xQ6EuHI9_0),.din(w_dff_A_4aciwrKU0_0),.clk(gclk));
	jdff dff_A_2xQ6EuHI9_0(.dout(w_dff_A_1vLH8UxP8_0),.din(w_dff_A_2xQ6EuHI9_0),.clk(gclk));
	jdff dff_A_1vLH8UxP8_0(.dout(G6170gat),.din(w_dff_A_1vLH8UxP8_0),.clk(gclk));
	jdff dff_A_2H3dPpHv5_2(.dout(w_dff_A_zGqYnJ693_0),.din(w_dff_A_2H3dPpHv5_2),.clk(gclk));
	jdff dff_A_zGqYnJ693_0(.dout(w_dff_A_SINlhkzL7_0),.din(w_dff_A_zGqYnJ693_0),.clk(gclk));
	jdff dff_A_SINlhkzL7_0(.dout(w_dff_A_Bc6xhLxp3_0),.din(w_dff_A_SINlhkzL7_0),.clk(gclk));
	jdff dff_A_Bc6xhLxp3_0(.dout(w_dff_A_XyAd7eVI4_0),.din(w_dff_A_Bc6xhLxp3_0),.clk(gclk));
	jdff dff_A_XyAd7eVI4_0(.dout(w_dff_A_PZ2v6xN74_0),.din(w_dff_A_XyAd7eVI4_0),.clk(gclk));
	jdff dff_A_PZ2v6xN74_0(.dout(w_dff_A_bw8PlNid0_0),.din(w_dff_A_PZ2v6xN74_0),.clk(gclk));
	jdff dff_A_bw8PlNid0_0(.dout(w_dff_A_xtiPKrGv5_0),.din(w_dff_A_bw8PlNid0_0),.clk(gclk));
	jdff dff_A_xtiPKrGv5_0(.dout(w_dff_A_eLofanXw5_0),.din(w_dff_A_xtiPKrGv5_0),.clk(gclk));
	jdff dff_A_eLofanXw5_0(.dout(w_dff_A_PKXkb4Os1_0),.din(w_dff_A_eLofanXw5_0),.clk(gclk));
	jdff dff_A_PKXkb4Os1_0(.dout(w_dff_A_SRpbTUPX1_0),.din(w_dff_A_PKXkb4Os1_0),.clk(gclk));
	jdff dff_A_SRpbTUPX1_0(.dout(w_dff_A_0XXQL3WG8_0),.din(w_dff_A_SRpbTUPX1_0),.clk(gclk));
	jdff dff_A_0XXQL3WG8_0(.dout(w_dff_A_TGwhWh9a2_0),.din(w_dff_A_0XXQL3WG8_0),.clk(gclk));
	jdff dff_A_TGwhWh9a2_0(.dout(w_dff_A_0TEZQyNz2_0),.din(w_dff_A_TGwhWh9a2_0),.clk(gclk));
	jdff dff_A_0TEZQyNz2_0(.dout(w_dff_A_jG0KZhr14_0),.din(w_dff_A_0TEZQyNz2_0),.clk(gclk));
	jdff dff_A_jG0KZhr14_0(.dout(w_dff_A_V4sVFDLJ3_0),.din(w_dff_A_jG0KZhr14_0),.clk(gclk));
	jdff dff_A_V4sVFDLJ3_0(.dout(w_dff_A_g5ZRMeTb6_0),.din(w_dff_A_V4sVFDLJ3_0),.clk(gclk));
	jdff dff_A_g5ZRMeTb6_0(.dout(w_dff_A_fewmH9SB0_0),.din(w_dff_A_g5ZRMeTb6_0),.clk(gclk));
	jdff dff_A_fewmH9SB0_0(.dout(w_dff_A_MS0plOq66_0),.din(w_dff_A_fewmH9SB0_0),.clk(gclk));
	jdff dff_A_MS0plOq66_0(.dout(w_dff_A_DHiYfBnH8_0),.din(w_dff_A_MS0plOq66_0),.clk(gclk));
	jdff dff_A_DHiYfBnH8_0(.dout(w_dff_A_Sil1Kgkq5_0),.din(w_dff_A_DHiYfBnH8_0),.clk(gclk));
	jdff dff_A_Sil1Kgkq5_0(.dout(w_dff_A_cy4DZ6lv3_0),.din(w_dff_A_Sil1Kgkq5_0),.clk(gclk));
	jdff dff_A_cy4DZ6lv3_0(.dout(w_dff_A_csOQGDMp5_0),.din(w_dff_A_cy4DZ6lv3_0),.clk(gclk));
	jdff dff_A_csOQGDMp5_0(.dout(G6180gat),.din(w_dff_A_csOQGDMp5_0),.clk(gclk));
	jdff dff_A_nFZwUN7m5_2(.dout(w_dff_A_wCP1GDwg3_0),.din(w_dff_A_nFZwUN7m5_2),.clk(gclk));
	jdff dff_A_wCP1GDwg3_0(.dout(w_dff_A_TuJYL9Bw9_0),.din(w_dff_A_wCP1GDwg3_0),.clk(gclk));
	jdff dff_A_TuJYL9Bw9_0(.dout(w_dff_A_bQHtmJrg1_0),.din(w_dff_A_TuJYL9Bw9_0),.clk(gclk));
	jdff dff_A_bQHtmJrg1_0(.dout(w_dff_A_EHh4ViMa5_0),.din(w_dff_A_bQHtmJrg1_0),.clk(gclk));
	jdff dff_A_EHh4ViMa5_0(.dout(w_dff_A_v1wTa9oT6_0),.din(w_dff_A_EHh4ViMa5_0),.clk(gclk));
	jdff dff_A_v1wTa9oT6_0(.dout(w_dff_A_0BRWUEF80_0),.din(w_dff_A_v1wTa9oT6_0),.clk(gclk));
	jdff dff_A_0BRWUEF80_0(.dout(w_dff_A_ZHZDjXgd2_0),.din(w_dff_A_0BRWUEF80_0),.clk(gclk));
	jdff dff_A_ZHZDjXgd2_0(.dout(w_dff_A_cDq0aF7i9_0),.din(w_dff_A_ZHZDjXgd2_0),.clk(gclk));
	jdff dff_A_cDq0aF7i9_0(.dout(w_dff_A_k3rsHM7N8_0),.din(w_dff_A_cDq0aF7i9_0),.clk(gclk));
	jdff dff_A_k3rsHM7N8_0(.dout(w_dff_A_kta9keZ81_0),.din(w_dff_A_k3rsHM7N8_0),.clk(gclk));
	jdff dff_A_kta9keZ81_0(.dout(w_dff_A_JckzmQxj7_0),.din(w_dff_A_kta9keZ81_0),.clk(gclk));
	jdff dff_A_JckzmQxj7_0(.dout(w_dff_A_DjcrbS1d8_0),.din(w_dff_A_JckzmQxj7_0),.clk(gclk));
	jdff dff_A_DjcrbS1d8_0(.dout(w_dff_A_lcs140vB1_0),.din(w_dff_A_DjcrbS1d8_0),.clk(gclk));
	jdff dff_A_lcs140vB1_0(.dout(w_dff_A_rgnMc04L7_0),.din(w_dff_A_lcs140vB1_0),.clk(gclk));
	jdff dff_A_rgnMc04L7_0(.dout(w_dff_A_rcswlGYS6_0),.din(w_dff_A_rgnMc04L7_0),.clk(gclk));
	jdff dff_A_rcswlGYS6_0(.dout(w_dff_A_Nvj4k6Rj6_0),.din(w_dff_A_rcswlGYS6_0),.clk(gclk));
	jdff dff_A_Nvj4k6Rj6_0(.dout(w_dff_A_n7maCWAC0_0),.din(w_dff_A_Nvj4k6Rj6_0),.clk(gclk));
	jdff dff_A_n7maCWAC0_0(.dout(w_dff_A_wcRGgzfw3_0),.din(w_dff_A_n7maCWAC0_0),.clk(gclk));
	jdff dff_A_wcRGgzfw3_0(.dout(w_dff_A_p0dNXKDc3_0),.din(w_dff_A_wcRGgzfw3_0),.clk(gclk));
	jdff dff_A_p0dNXKDc3_0(.dout(w_dff_A_7A6bt52y7_0),.din(w_dff_A_p0dNXKDc3_0),.clk(gclk));
	jdff dff_A_7A6bt52y7_0(.dout(G6190gat),.din(w_dff_A_7A6bt52y7_0),.clk(gclk));
	jdff dff_A_BTnUMnAU7_2(.dout(w_dff_A_yDpE8sMw3_0),.din(w_dff_A_BTnUMnAU7_2),.clk(gclk));
	jdff dff_A_yDpE8sMw3_0(.dout(w_dff_A_zAbpuylL6_0),.din(w_dff_A_yDpE8sMw3_0),.clk(gclk));
	jdff dff_A_zAbpuylL6_0(.dout(w_dff_A_Jniz9VPd4_0),.din(w_dff_A_zAbpuylL6_0),.clk(gclk));
	jdff dff_A_Jniz9VPd4_0(.dout(w_dff_A_ynRMVfXO9_0),.din(w_dff_A_Jniz9VPd4_0),.clk(gclk));
	jdff dff_A_ynRMVfXO9_0(.dout(w_dff_A_CyTXiea32_0),.din(w_dff_A_ynRMVfXO9_0),.clk(gclk));
	jdff dff_A_CyTXiea32_0(.dout(w_dff_A_cfWCba7g3_0),.din(w_dff_A_CyTXiea32_0),.clk(gclk));
	jdff dff_A_cfWCba7g3_0(.dout(w_dff_A_rL3YDsfb0_0),.din(w_dff_A_cfWCba7g3_0),.clk(gclk));
	jdff dff_A_rL3YDsfb0_0(.dout(w_dff_A_5eiugd7Z3_0),.din(w_dff_A_rL3YDsfb0_0),.clk(gclk));
	jdff dff_A_5eiugd7Z3_0(.dout(w_dff_A_DzHrCLbt5_0),.din(w_dff_A_5eiugd7Z3_0),.clk(gclk));
	jdff dff_A_DzHrCLbt5_0(.dout(w_dff_A_FI9jyE854_0),.din(w_dff_A_DzHrCLbt5_0),.clk(gclk));
	jdff dff_A_FI9jyE854_0(.dout(w_dff_A_H3LZ7MPh8_0),.din(w_dff_A_FI9jyE854_0),.clk(gclk));
	jdff dff_A_H3LZ7MPh8_0(.dout(w_dff_A_sCCm3opL9_0),.din(w_dff_A_H3LZ7MPh8_0),.clk(gclk));
	jdff dff_A_sCCm3opL9_0(.dout(w_dff_A_dYeziSMj6_0),.din(w_dff_A_sCCm3opL9_0),.clk(gclk));
	jdff dff_A_dYeziSMj6_0(.dout(w_dff_A_vmKejPkQ0_0),.din(w_dff_A_dYeziSMj6_0),.clk(gclk));
	jdff dff_A_vmKejPkQ0_0(.dout(w_dff_A_CJtxRjim8_0),.din(w_dff_A_vmKejPkQ0_0),.clk(gclk));
	jdff dff_A_CJtxRjim8_0(.dout(w_dff_A_1ctpGbgg5_0),.din(w_dff_A_CJtxRjim8_0),.clk(gclk));
	jdff dff_A_1ctpGbgg5_0(.dout(w_dff_A_JKXbp7w75_0),.din(w_dff_A_1ctpGbgg5_0),.clk(gclk));
	jdff dff_A_JKXbp7w75_0(.dout(w_dff_A_LRHSc0ac9_0),.din(w_dff_A_JKXbp7w75_0),.clk(gclk));
	jdff dff_A_LRHSc0ac9_0(.dout(G6200gat),.din(w_dff_A_LRHSc0ac9_0),.clk(gclk));
	jdff dff_A_96BrlB423_2(.dout(w_dff_A_6L2TBEwC3_0),.din(w_dff_A_96BrlB423_2),.clk(gclk));
	jdff dff_A_6L2TBEwC3_0(.dout(w_dff_A_ECb3B5yj2_0),.din(w_dff_A_6L2TBEwC3_0),.clk(gclk));
	jdff dff_A_ECb3B5yj2_0(.dout(w_dff_A_N9Ade0XG7_0),.din(w_dff_A_ECb3B5yj2_0),.clk(gclk));
	jdff dff_A_N9Ade0XG7_0(.dout(w_dff_A_HVjBrLV06_0),.din(w_dff_A_N9Ade0XG7_0),.clk(gclk));
	jdff dff_A_HVjBrLV06_0(.dout(w_dff_A_LMhO7NQ81_0),.din(w_dff_A_HVjBrLV06_0),.clk(gclk));
	jdff dff_A_LMhO7NQ81_0(.dout(w_dff_A_XQ8lBCio4_0),.din(w_dff_A_LMhO7NQ81_0),.clk(gclk));
	jdff dff_A_XQ8lBCio4_0(.dout(w_dff_A_EQFvMxPh9_0),.din(w_dff_A_XQ8lBCio4_0),.clk(gclk));
	jdff dff_A_EQFvMxPh9_0(.dout(w_dff_A_4RSN6NPj4_0),.din(w_dff_A_EQFvMxPh9_0),.clk(gclk));
	jdff dff_A_4RSN6NPj4_0(.dout(w_dff_A_Ge9Wk7tA2_0),.din(w_dff_A_4RSN6NPj4_0),.clk(gclk));
	jdff dff_A_Ge9Wk7tA2_0(.dout(w_dff_A_GPo7kuIa4_0),.din(w_dff_A_Ge9Wk7tA2_0),.clk(gclk));
	jdff dff_A_GPo7kuIa4_0(.dout(w_dff_A_VXvFFCb12_0),.din(w_dff_A_GPo7kuIa4_0),.clk(gclk));
	jdff dff_A_VXvFFCb12_0(.dout(w_dff_A_KZLK5GGh2_0),.din(w_dff_A_VXvFFCb12_0),.clk(gclk));
	jdff dff_A_KZLK5GGh2_0(.dout(w_dff_A_rG1oGnWq8_0),.din(w_dff_A_KZLK5GGh2_0),.clk(gclk));
	jdff dff_A_rG1oGnWq8_0(.dout(w_dff_A_BazaDLNT9_0),.din(w_dff_A_rG1oGnWq8_0),.clk(gclk));
	jdff dff_A_BazaDLNT9_0(.dout(w_dff_A_UJbvnSdq0_0),.din(w_dff_A_BazaDLNT9_0),.clk(gclk));
	jdff dff_A_UJbvnSdq0_0(.dout(w_dff_A_Eh2gmav45_0),.din(w_dff_A_UJbvnSdq0_0),.clk(gclk));
	jdff dff_A_Eh2gmav45_0(.dout(G6210gat),.din(w_dff_A_Eh2gmav45_0),.clk(gclk));
	jdff dff_A_oWs98O0Y7_2(.dout(w_dff_A_YbnRnyt18_0),.din(w_dff_A_oWs98O0Y7_2),.clk(gclk));
	jdff dff_A_YbnRnyt18_0(.dout(w_dff_A_DYu5ZkHt0_0),.din(w_dff_A_YbnRnyt18_0),.clk(gclk));
	jdff dff_A_DYu5ZkHt0_0(.dout(w_dff_A_pkr6GAxp8_0),.din(w_dff_A_DYu5ZkHt0_0),.clk(gclk));
	jdff dff_A_pkr6GAxp8_0(.dout(w_dff_A_3C4cP3FN5_0),.din(w_dff_A_pkr6GAxp8_0),.clk(gclk));
	jdff dff_A_3C4cP3FN5_0(.dout(w_dff_A_WxBtqsJX7_0),.din(w_dff_A_3C4cP3FN5_0),.clk(gclk));
	jdff dff_A_WxBtqsJX7_0(.dout(w_dff_A_rPkki8Nx6_0),.din(w_dff_A_WxBtqsJX7_0),.clk(gclk));
	jdff dff_A_rPkki8Nx6_0(.dout(w_dff_A_AXNVxNfd5_0),.din(w_dff_A_rPkki8Nx6_0),.clk(gclk));
	jdff dff_A_AXNVxNfd5_0(.dout(w_dff_A_UcjgaseF0_0),.din(w_dff_A_AXNVxNfd5_0),.clk(gclk));
	jdff dff_A_UcjgaseF0_0(.dout(w_dff_A_rvDdg6zP3_0),.din(w_dff_A_UcjgaseF0_0),.clk(gclk));
	jdff dff_A_rvDdg6zP3_0(.dout(w_dff_A_2U5jOXBD8_0),.din(w_dff_A_rvDdg6zP3_0),.clk(gclk));
	jdff dff_A_2U5jOXBD8_0(.dout(w_dff_A_FIRCRgyq9_0),.din(w_dff_A_2U5jOXBD8_0),.clk(gclk));
	jdff dff_A_FIRCRgyq9_0(.dout(w_dff_A_PMzcuCJm9_0),.din(w_dff_A_FIRCRgyq9_0),.clk(gclk));
	jdff dff_A_PMzcuCJm9_0(.dout(w_dff_A_Qm1n0uAa5_0),.din(w_dff_A_PMzcuCJm9_0),.clk(gclk));
	jdff dff_A_Qm1n0uAa5_0(.dout(w_dff_A_PRGfI1FU0_0),.din(w_dff_A_Qm1n0uAa5_0),.clk(gclk));
	jdff dff_A_PRGfI1FU0_0(.dout(G6220gat),.din(w_dff_A_PRGfI1FU0_0),.clk(gclk));
	jdff dff_A_IFaEiPVG2_2(.dout(w_dff_A_g1szHesY8_0),.din(w_dff_A_IFaEiPVG2_2),.clk(gclk));
	jdff dff_A_g1szHesY8_0(.dout(w_dff_A_TBgoZo4N9_0),.din(w_dff_A_g1szHesY8_0),.clk(gclk));
	jdff dff_A_TBgoZo4N9_0(.dout(w_dff_A_baN9XbAo0_0),.din(w_dff_A_TBgoZo4N9_0),.clk(gclk));
	jdff dff_A_baN9XbAo0_0(.dout(w_dff_A_RlyKUGeq5_0),.din(w_dff_A_baN9XbAo0_0),.clk(gclk));
	jdff dff_A_RlyKUGeq5_0(.dout(w_dff_A_Sq8ptWYj3_0),.din(w_dff_A_RlyKUGeq5_0),.clk(gclk));
	jdff dff_A_Sq8ptWYj3_0(.dout(w_dff_A_3t4g6c3I0_0),.din(w_dff_A_Sq8ptWYj3_0),.clk(gclk));
	jdff dff_A_3t4g6c3I0_0(.dout(w_dff_A_7eom11wB9_0),.din(w_dff_A_3t4g6c3I0_0),.clk(gclk));
	jdff dff_A_7eom11wB9_0(.dout(w_dff_A_2x5unCXl3_0),.din(w_dff_A_7eom11wB9_0),.clk(gclk));
	jdff dff_A_2x5unCXl3_0(.dout(w_dff_A_RJKDsMbD7_0),.din(w_dff_A_2x5unCXl3_0),.clk(gclk));
	jdff dff_A_RJKDsMbD7_0(.dout(w_dff_A_Re64RGVU3_0),.din(w_dff_A_RJKDsMbD7_0),.clk(gclk));
	jdff dff_A_Re64RGVU3_0(.dout(w_dff_A_bFU1C6921_0),.din(w_dff_A_Re64RGVU3_0),.clk(gclk));
	jdff dff_A_bFU1C6921_0(.dout(w_dff_A_H4DQHubn4_0),.din(w_dff_A_bFU1C6921_0),.clk(gclk));
	jdff dff_A_H4DQHubn4_0(.dout(G6230gat),.din(w_dff_A_H4DQHubn4_0),.clk(gclk));
	jdff dff_A_iPM9LwlQ1_2(.dout(w_dff_A_BSFUGiiD3_0),.din(w_dff_A_iPM9LwlQ1_2),.clk(gclk));
	jdff dff_A_BSFUGiiD3_0(.dout(w_dff_A_U6tWwpAv3_0),.din(w_dff_A_BSFUGiiD3_0),.clk(gclk));
	jdff dff_A_U6tWwpAv3_0(.dout(w_dff_A_60EC0Zj36_0),.din(w_dff_A_U6tWwpAv3_0),.clk(gclk));
	jdff dff_A_60EC0Zj36_0(.dout(w_dff_A_Ui8GvQhv0_0),.din(w_dff_A_60EC0Zj36_0),.clk(gclk));
	jdff dff_A_Ui8GvQhv0_0(.dout(w_dff_A_MtvFY0gW8_0),.din(w_dff_A_Ui8GvQhv0_0),.clk(gclk));
	jdff dff_A_MtvFY0gW8_0(.dout(w_dff_A_5vIlxAwr8_0),.din(w_dff_A_MtvFY0gW8_0),.clk(gclk));
	jdff dff_A_5vIlxAwr8_0(.dout(w_dff_A_ukTT6Mmc0_0),.din(w_dff_A_5vIlxAwr8_0),.clk(gclk));
	jdff dff_A_ukTT6Mmc0_0(.dout(w_dff_A_e7uD8wLC2_0),.din(w_dff_A_ukTT6Mmc0_0),.clk(gclk));
	jdff dff_A_e7uD8wLC2_0(.dout(w_dff_A_CmzlbS8M7_0),.din(w_dff_A_e7uD8wLC2_0),.clk(gclk));
	jdff dff_A_CmzlbS8M7_0(.dout(w_dff_A_hVZ4EwjM5_0),.din(w_dff_A_CmzlbS8M7_0),.clk(gclk));
	jdff dff_A_hVZ4EwjM5_0(.dout(G6240gat),.din(w_dff_A_hVZ4EwjM5_0),.clk(gclk));
	jdff dff_A_4ZSUinxL1_2(.dout(w_dff_A_8vznccM88_0),.din(w_dff_A_4ZSUinxL1_2),.clk(gclk));
	jdff dff_A_8vznccM88_0(.dout(w_dff_A_4EbhWlwH9_0),.din(w_dff_A_8vznccM88_0),.clk(gclk));
	jdff dff_A_4EbhWlwH9_0(.dout(w_dff_A_0FB3gmKz9_0),.din(w_dff_A_4EbhWlwH9_0),.clk(gclk));
	jdff dff_A_0FB3gmKz9_0(.dout(w_dff_A_I3FHZ6Ns0_0),.din(w_dff_A_0FB3gmKz9_0),.clk(gclk));
	jdff dff_A_I3FHZ6Ns0_0(.dout(w_dff_A_L0s8w6739_0),.din(w_dff_A_I3FHZ6Ns0_0),.clk(gclk));
	jdff dff_A_L0s8w6739_0(.dout(w_dff_A_DbJuQ1rh1_0),.din(w_dff_A_L0s8w6739_0),.clk(gclk));
	jdff dff_A_DbJuQ1rh1_0(.dout(w_dff_A_jMcL0vjA6_0),.din(w_dff_A_DbJuQ1rh1_0),.clk(gclk));
	jdff dff_A_jMcL0vjA6_0(.dout(w_dff_A_Ip7LTZOl9_0),.din(w_dff_A_jMcL0vjA6_0),.clk(gclk));
	jdff dff_A_Ip7LTZOl9_0(.dout(G6250gat),.din(w_dff_A_Ip7LTZOl9_0),.clk(gclk));
	jdff dff_A_jerCFLUD1_2(.dout(w_dff_A_OzM6UivC1_0),.din(w_dff_A_jerCFLUD1_2),.clk(gclk));
	jdff dff_A_OzM6UivC1_0(.dout(w_dff_A_UwqzvO0V4_0),.din(w_dff_A_OzM6UivC1_0),.clk(gclk));
	jdff dff_A_UwqzvO0V4_0(.dout(w_dff_A_7qdSojmy8_0),.din(w_dff_A_UwqzvO0V4_0),.clk(gclk));
	jdff dff_A_7qdSojmy8_0(.dout(w_dff_A_UFwoG57b5_0),.din(w_dff_A_7qdSojmy8_0),.clk(gclk));
	jdff dff_A_UFwoG57b5_0(.dout(w_dff_A_NcaGpnbc9_0),.din(w_dff_A_UFwoG57b5_0),.clk(gclk));
	jdff dff_A_NcaGpnbc9_0(.dout(w_dff_A_WS5t0grE8_0),.din(w_dff_A_NcaGpnbc9_0),.clk(gclk));
	jdff dff_A_WS5t0grE8_0(.dout(G6260gat),.din(w_dff_A_WS5t0grE8_0),.clk(gclk));
	jdff dff_A_AZmphtiy6_2(.dout(w_dff_A_ro53mV445_0),.din(w_dff_A_AZmphtiy6_2),.clk(gclk));
	jdff dff_A_ro53mV445_0(.dout(w_dff_A_yYNv67ns6_0),.din(w_dff_A_ro53mV445_0),.clk(gclk));
	jdff dff_A_yYNv67ns6_0(.dout(w_dff_A_k7BRES2e4_0),.din(w_dff_A_yYNv67ns6_0),.clk(gclk));
	jdff dff_A_k7BRES2e4_0(.dout(w_dff_A_ihGoirPu7_0),.din(w_dff_A_k7BRES2e4_0),.clk(gclk));
	jdff dff_A_ihGoirPu7_0(.dout(G6270gat),.din(w_dff_A_ihGoirPu7_0),.clk(gclk));
	jdff dff_A_VrGQGW8r1_2(.dout(w_dff_A_TSBcsTUK5_0),.din(w_dff_A_VrGQGW8r1_2),.clk(gclk));
	jdff dff_A_TSBcsTUK5_0(.dout(w_dff_A_2SWcjTOU1_0),.din(w_dff_A_TSBcsTUK5_0),.clk(gclk));
	jdff dff_A_2SWcjTOU1_0(.dout(G6280gat),.din(w_dff_A_2SWcjTOU1_0),.clk(gclk));
	jdff dff_A_JNspNrBf3_2(.dout(G6288gat),.din(w_dff_A_JNspNrBf3_2),.clk(gclk));
endmodule

