/*

c432:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jcb: 110
	jdff: 752
	jand: 111

Summary:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jcb: 110
	jdff: 752
	jand: 111
*/

module c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n43;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n150;
	wire n151;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n217;
	wire n218;
	wire n219;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n235;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n244;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n262;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G4gat_0;
	wire [2:0] w_G8gat_0;
	wire [2:0] w_G11gat_0;
	wire [2:0] w_G14gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G21gat_0;
	wire [1:0] w_G21gat_1;
	wire [1:0] w_G24gat_0;
	wire [1:0] w_G27gat_0;
	wire [1:0] w_G30gat_0;
	wire [2:0] w_G34gat_0;
	wire [2:0] w_G37gat_0;
	wire [1:0] w_G40gat_0;
	wire [2:0] w_G43gat_0;
	wire [1:0] w_G43gat_1;
	wire [1:0] w_G47gat_0;
	wire [2:0] w_G50gat_0;
	wire [1:0] w_G53gat_0;
	wire [2:0] w_G56gat_0;
	wire [2:0] w_G60gat_0;
	wire [2:0] w_G63gat_0;
	wire [1:0] w_G66gat_0;
	wire [2:0] w_G69gat_0;
	wire [2:0] w_G73gat_0;
	wire [1:0] w_G76gat_0;
	wire [1:0] w_G79gat_0;
	wire [2:0] w_G82gat_0;
	wire [2:0] w_G86gat_0;
	wire [1:0] w_G86gat_1;
	wire [2:0] w_G89gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G95gat_0;
	wire [2:0] w_G99gat_0;
	wire [2:0] w_G102gat_0;
	wire [1:0] w_G105gat_0;
	wire [2:0] w_G108gat_0;
	wire [2:0] w_G112gat_0;
	wire [1:0] w_G115gat_0;
	wire [2:0] w_G223gat_0;
	wire [2:0] w_G223gat_1;
	wire [2:0] w_G223gat_2;
	wire [1:0] w_G223gat_3;
	wire G223gat_fa_;
	wire [2:0] w_G329gat_0;
	wire [2:0] w_G329gat_1;
	wire [2:0] w_G329gat_2;
	wire [2:0] w_G329gat_3;
	wire [2:0] w_G329gat_4;
	wire [2:0] w_G329gat_5;
	wire w_G329gat_6;
	wire G329gat_fa_;
	wire [2:0] w_G370gat_0;
	wire [2:0] w_G370gat_1;
	wire w_G370gat_2;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire [1:0] w_n43_0;
	wire [1:0] w_n44_0;
	wire [1:0] w_n47_0;
	wire [1:0] w_n52_0;
	wire [1:0] w_n53_0;
	wire [1:0] w_n56_0;
	wire [1:0] w_n58_0;
	wire [1:0] w_n61_0;
	wire [1:0] w_n63_0;
	wire [1:0] w_n69_0;
	wire [1:0] w_n71_0;
	wire [1:0] w_n72_0;
	wire [1:0] w_n73_0;
	wire [1:0] w_n77_0;
	wire [1:0] w_n78_0;
	wire [1:0] w_n79_0;
	wire [1:0] w_n82_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n87_0;
	wire [1:0] w_n89_0;
	wire [2:0] w_n94_0;
	wire [2:0] w_n94_1;
	wire [2:0] w_n94_2;
	wire [2:0] w_n94_3;
	wire [1:0] w_n94_4;
	wire [1:0] w_n96_0;
	wire [1:0] w_n98_0;
	wire [1:0] w_n100_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n109_0;
	wire [2:0] w_n114_0;
	wire [1:0] w_n115_0;
	wire [1:0] w_n119_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n123_0;
	wire [2:0] w_n126_0;
	wire [1:0] w_n128_0;
	wire [2:0] w_n130_0;
	wire [1:0] w_n132_0;
	wire [1:0] w_n139_0;
	wire [1:0] w_n141_0;
	wire [1:0] w_n142_0;
	wire [1:0] w_n145_0;
	wire [1:0] w_n146_0;
	wire [1:0] w_n147_0;
	wire [1:0] w_n150_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n154_0;
	wire [1:0] w_n156_0;
	wire [1:0] w_n159_0;
	wire [1:0] w_n164_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n174_0;
	wire [1:0] w_n177_0;
	wire [2:0] w_n182_0;
	wire [2:0] w_n182_1;
	wire [2:0] w_n182_2;
	wire [1:0] w_n182_3;
	wire [1:0] w_n184_0;
	wire [1:0] w_n188_0;
	wire [1:0] w_n191_0;
	wire [1:0] w_n193_0;
	wire [1:0] w_n197_0;
	wire [1:0] w_n198_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n217_0;
	wire [1:0] w_n219_0;
	wire [1:0] w_n222_0;
	wire [1:0] w_n224_0;
	wire [1:0] w_n231_0;
	wire [1:0] w_n254_0;
	wire [1:0] w_n260_0;
	wire [2:0] w_n271_0;
	wire [2:0] w_n271_1;
	wire [2:0] w_n271_2;
	wire [1:0] w_n271_3;
	wire [1:0] w_n274_0;
	wire [1:0] w_n281_0;
	wire [1:0] w_n283_0;
	wire [1:0] w_n286_0;
	wire [1:0] w_n290_0;
	wire [1:0] w_n293_0;
	wire [1:0] w_n296_0;
	wire [1:0] w_n303_0;
	wire [1:0] w_n305_0;
	wire [1:0] w_n313_0;
	wire [1:0] w_n314_0;
	wire [2:0] w_n317_0;
	wire [1:0] w_n319_0;
	wire w_dff_B_NNAzo5ez5_1;
	wire w_dff_B_LjWFwRck8_1;
	wire w_dff_B_KumAQcfB7_1;
	wire w_dff_B_re7nzJSS3_0;
	wire w_dff_B_7RirBMnF4_0;
	wire w_dff_B_DlRgxCvk4_0;
	wire w_dff_B_cqLXRr0u4_0;
	wire w_dff_B_eX5WKZFn6_0;
	wire w_dff_B_XTwMCCN78_0;
	wire w_dff_B_DT7GTFZ78_1;
	wire w_dff_A_VbrR3Svo9_0;
	wire w_dff_A_57a6Uuz23_0;
	wire w_dff_B_4CsutdP87_0;
	wire w_dff_B_rSWyHv3o3_0;
	wire w_dff_B_QTBEKGTI2_0;
	wire w_dff_B_BRRmZ4vR4_0;
	wire w_dff_B_kRRpcpBl2_0;
	wire w_dff_B_H7dSlUJY2_0;
	wire w_dff_B_wi0W0TXf6_0;
	wire w_dff_B_5VZfKCJ99_0;
	wire w_dff_B_aBdLMG4F6_0;
	wire w_dff_B_gyyUuk2t2_0;
	wire w_dff_B_1NKPMYqv0_0;
	wire w_dff_B_ykPddIkY9_0;
	wire w_dff_B_huyq7yRr4_0;
	wire w_dff_A_l8TA9xag9_0;
	wire w_dff_A_lC6q45058_0;
	wire w_dff_B_qacHT2eE3_2;
	wire w_dff_B_pDlUUxKz7_2;
	wire w_dff_A_QzSmpVMj2_0;
	wire w_dff_A_ajmtU2Kc5_0;
	wire w_dff_A_AUtTnTtB4_0;
	wire w_dff_A_YxinQqic0_0;
	wire w_dff_A_jLUDdNHJ6_0;
	wire w_dff_B_kx9oFqVr3_0;
	wire w_dff_B_sTlSopjC5_0;
	wire w_dff_B_0jpW6hqj9_0;
	wire w_dff_A_y4kzilGs0_0;
	wire w_dff_A_2gWDS8Pv5_0;
	wire w_dff_A_CESwO5LL4_0;
	wire w_dff_A_aghYQyFm5_0;
	wire w_dff_A_nCOlxojz0_0;
	wire w_dff_B_MKx9TkqZ7_0;
	wire w_dff_B_1WgPJZoq7_0;
	wire w_dff_B_hlTOnxwO7_0;
	wire w_dff_B_STSxD65J2_0;
	wire w_dff_B_WZY9NVfD0_0;
	wire w_dff_B_pMmHWCzx8_1;
	wire w_dff_B_SuetQrwe0_1;
	wire w_dff_B_kJU5ADqp7_1;
	wire w_dff_B_PbAjnpRW2_1;
	wire w_dff_B_tYvIWOvL3_1;
	wire w_dff_B_pOpfgyo86_1;
	wire w_dff_B_WXG14XJK5_1;
	wire w_dff_B_6COZDPs56_1;
	wire w_dff_B_iLSo7CQV5_1;
	wire w_dff_B_5aytIf7K8_1;
	wire w_dff_B_LGlF82Bj9_1;
	wire w_dff_B_WxnLOgQu4_1;
	wire w_dff_B_CbHy5VSx4_1;
	wire w_dff_B_AsHoFPKM0_1;
	wire w_dff_B_usN9BBhI1_1;
	wire w_dff_B_XdWY8pKv6_1;
	wire w_dff_B_fFN1zz8A3_1;
	wire w_dff_B_QzanNSGG8_1;
	wire w_dff_B_MCw2aYup6_1;
	wire w_dff_B_G9r9K1T88_1;
	wire w_dff_B_nDzhsVir4_1;
	wire w_dff_B_9LZIO7vR5_1;
	wire w_dff_B_zI66Mbb68_1;
	wire w_dff_B_BlhSNEHh9_1;
	wire w_dff_B_nKBhQB1W6_1;
	wire w_dff_B_mtQiiog55_0;
	wire w_dff_B_q1ZvadfE8_0;
	wire w_dff_B_RuLZw8Ua2_0;
	wire w_dff_B_VDGaAm5s7_0;
	wire w_dff_B_FzdHCtZe2_0;
	wire w_dff_B_dBUvcGT71_0;
	wire w_dff_A_IbpRZwoY1_1;
	wire w_dff_A_6SQvWR6o7_1;
	wire w_dff_A_nSldGmhS8_1;
	wire w_dff_A_ER1SrXHP2_1;
	wire w_dff_A_tPfc51Xj1_1;
	wire w_dff_A_5PS2gS7j8_0;
	wire w_dff_A_YDJ1gxww5_0;
	wire w_dff_B_qCFSnN2y9_2;
	wire w_dff_B_vHMFABkU9_2;
	wire w_dff_B_cw23lUTm5_2;
	wire w_dff_B_k1nrhP409_1;
	wire w_dff_B_kBUEQRTF0_1;
	wire w_dff_B_63L91ISR7_1;
	wire w_dff_B_ADThpRlJ6_1;
	wire w_dff_B_UEHS9Rue4_1;
	wire w_dff_B_cx9NWvkF0_1;
	wire w_dff_B_0ez9y9bH3_3;
	wire w_dff_B_BhTVwoiE5_3;
	wire w_dff_B_hXQrdu6m1_3;
	wire w_dff_A_fJ3BgBZi1_0;
	wire w_dff_A_bwjzrf8s6_0;
	wire w_dff_A_E2ysPMuG0_0;
	wire w_dff_A_rtfRFXE34_0;
	wire w_dff_A_twwzGNpN2_0;
	wire w_dff_A_hueS9QO64_1;
	wire w_dff_B_NfZgjlwf5_1;
	wire w_dff_A_NT74VLku4_0;
	wire w_dff_A_cE2g9gf94_0;
	wire w_dff_A_W0FYNaVC8_0;
	wire w_dff_A_wO3lTOII3_0;
	wire w_dff_A_PRB0O4F03_0;
	wire w_dff_A_NFUlC0aO7_0;
	wire w_dff_A_RLmbjydG7_0;
	wire w_dff_A_jUKicEId0_0;
	wire w_dff_B_QPu4F5w71_2;
	wire w_dff_B_74pYg0I73_2;
	wire w_dff_B_kMHmiD887_2;
	wire w_dff_B_4d9Ks3Kf6_2;
	wire w_dff_B_2QA2Dpgb7_2;
	wire w_dff_B_m7tctwbd5_2;
	wire w_dff_B_13boSzhX0_2;
	wire w_dff_B_LhaKIiE29_2;
	wire w_dff_B_4wcdZRlD8_2;
	wire w_dff_B_dAgSW9SZ3_2;
	wire w_dff_A_IYR4xoeH0_0;
	wire w_dff_A_xZN92ch06_0;
	wire w_dff_A_E8iWS6TP6_0;
	wire w_dff_A_c3fldacj6_0;
	wire w_dff_A_p5dQdp7B1_0;
	wire w_dff_A_bDMsQRBX9_0;
	wire w_dff_A_4EA5zdRI4_0;
	wire w_dff_A_jovG9FKY9_0;
	wire w_dff_A_UBfoKA1H8_1;
	wire w_dff_A_Kz7b49HT1_1;
	wire w_dff_A_TRga1sTf0_0;
	wire w_dff_A_5jgl3oVI5_0;
	wire w_dff_A_ydR0BTVG5_0;
	wire w_dff_A_ZYiiNVLQ6_0;
	wire w_dff_A_x99nVF944_0;
	wire w_dff_A_kpfsJ6rd1_0;
	wire w_dff_A_uG6fHCXf6_0;
	wire w_dff_A_fH58VTXp6_0;
	wire w_dff_B_klVZumzE8_2;
	wire w_dff_B_uUPXFwHZ8_2;
	wire w_dff_B_qNaHHyIp1_2;
	wire w_dff_B_ZdyRjlON2_2;
	wire w_dff_B_xww0tWIQ3_2;
	wire w_dff_B_p270DQTj0_2;
	wire w_dff_A_xj2sYUjV9_0;
	wire w_dff_A_R0QeNTxd5_0;
	wire w_dff_A_DgzJYiL52_0;
	wire w_dff_A_ydn6721I3_0;
	wire w_dff_A_gl96Tb8m4_0;
	wire w_dff_A_SxYdW0EY2_0;
	wire w_dff_A_iz3CEMhh3_0;
	wire w_dff_A_sOYWmSRN7_0;
	wire w_dff_A_OdLRWxCG1_0;
	wire w_dff_A_lQ80jKB65_0;
	wire w_dff_A_Jn7ijbyN7_0;
	wire w_dff_A_BdJINvIe4_0;
	wire w_dff_B_aUb5jDP07_1;
	wire w_dff_B_7h3X1Cgb7_1;
	wire w_dff_B_lutzR7G29_1;
	wire w_dff_B_IttGQTE16_1;
	wire w_dff_B_lq9qRrrh7_1;
	wire w_dff_B_r4DKtmoG9_1;
	wire w_dff_B_mgImKyoN3_1;
	wire w_dff_B_dg3ww7RA6_1;
	wire w_dff_B_VCU9QS1w1_1;
	wire w_dff_B_RTlDi3Jd6_1;
	wire w_dff_B_wOlzNPsq8_1;
	wire w_dff_B_wjvURLz65_1;
	wire w_dff_B_p18gYLXB7_1;
	wire w_dff_B_hhYWuN8p8_1;
	wire w_dff_B_jRmp4DZU2_1;
	wire w_dff_B_WB9UUlEd5_1;
	wire w_dff_B_oq4HkBVB6_1;
	wire w_dff_B_nzZemYMx0_1;
	wire w_dff_B_SLm6IIqn0_1;
	wire w_dff_A_s7LV3qY29_0;
	wire w_dff_A_zLyxdrxy5_0;
	wire w_dff_A_qiqysHQD8_0;
	wire w_dff_A_amCkDlQG0_0;
	wire w_dff_A_unzlrDbQ0_0;
	wire w_dff_A_DLenJcZs5_0;
	wire w_dff_A_33WDRoqx6_0;
	wire w_dff_A_n6XHEdUj8_0;
	wire w_dff_A_aoPBYSjc7_1;
	wire w_dff_A_GVLtgWZY8_1;
	wire w_dff_A_ONnW7Y279_1;
	wire w_dff_A_TjsBU9JQ2_1;
	wire w_dff_A_Gd3cNstL9_1;
	wire w_dff_A_xsQPmKib1_1;
	wire w_dff_A_P8Drobbj0_1;
	wire w_dff_A_d13K1z2Z8_1;
	wire w_dff_A_7CHHER2a3_1;
	wire w_dff_A_fIl2YIaC5_1;
	wire w_dff_A_xUkjWZZx2_1;
	wire w_dff_A_UQ0gZUMf1_1;
	wire w_dff_B_0Fm7J8cP5_0;
	wire w_dff_B_NB6VqPUe9_0;
	wire w_dff_B_OX8CYYjJ6_0;
	wire w_dff_A_EZ66K8I56_0;
	wire w_dff_A_QIXAY9WK7_0;
	wire w_dff_A_uC5b3hSA3_0;
	wire w_dff_A_h4em9AGo8_0;
	wire w_dff_A_tIGfwHGg2_0;
	wire w_dff_A_J8QPLg9J7_0;
	wire w_dff_A_MFJeeaF62_0;
	wire w_dff_A_1sgwg0GZ7_0;
	wire w_dff_B_j6icMxLW8_2;
	wire w_dff_B_ViB2Df705_2;
	wire w_dff_B_X6v2frNB4_2;
	wire w_dff_B_GhwuFCdQ1_2;
	wire w_dff_B_mQ6TBImH6_2;
	wire w_dff_B_T1KCYwbu9_2;
	wire w_dff_A_ZQM77ijN8_0;
	wire w_dff_A_gLHxr5VE8_0;
	wire w_dff_A_UH5r1ecC3_0;
	wire w_dff_A_i1NsmZSa3_0;
	wire w_dff_A_kUCTXTQI4_0;
	wire w_dff_A_w64DdZxZ0_0;
	wire w_dff_A_h2w8RUEb4_0;
	wire w_dff_A_ZW076xdY9_0;
	wire w_dff_A_7p5qUIwD9_0;
	wire w_dff_A_4DZfS5Xn2_0;
	wire w_dff_A_sHGoiaU70_0;
	wire w_dff_A_T3NsGRQx8_0;
	wire w_dff_A_hMVbeRty0_1;
	wire w_dff_A_i0yxT9Qv6_1;
	wire w_dff_A_Hw8MJEYn1_1;
	wire w_dff_A_yYO2Wevq8_1;
	wire w_dff_A_X7C3Aba86_1;
	wire w_dff_A_etXGr1iD5_1;
	wire w_dff_A_ct50e6pk0_1;
	wire w_dff_A_bVOGG39t0_1;
	wire w_dff_A_iYtOsyqy6_1;
	wire w_dff_A_YSMFNW3H9_1;
	wire w_dff_A_F9SGUW079_1;
	wire w_dff_A_9bFtK4IS8_0;
	wire w_dff_A_OIwkqYyV4_0;
	wire w_dff_A_ZUT9YEWU6_0;
	wire w_dff_A_ZXqWWYqh1_0;
	wire w_dff_B_yha5fpCJ9_1;
	wire w_dff_B_JanIzsh28_1;
	wire w_dff_B_YM6zdRQQ9_0;
	wire w_dff_B_lk5jbvF57_0;
	wire w_dff_B_RJacCCyX8_0;
	wire w_dff_A_otWel9Ab8_0;
	wire w_dff_A_4bvWgYgg2_0;
	wire w_dff_A_vwNK0Yky6_0;
	wire w_dff_A_jS1q47vm7_0;
	wire w_dff_A_dYdWcGhN9_0;
	wire w_dff_A_Cwm2wRgm1_0;
	wire w_dff_A_LjWVac3z9_0;
	wire w_dff_A_lvyuG3S28_0;
	wire w_dff_B_hCMkpj2D8_2;
	wire w_dff_B_lMUpE1dq4_2;
	wire w_dff_B_ApHbSPsA1_2;
	wire w_dff_B_80e3dtk22_2;
	wire w_dff_B_8KIQ7lgq9_2;
	wire w_dff_B_gn2lZ5EV5_2;
	wire w_dff_A_yTMzwNf05_0;
	wire w_dff_A_8uQ57ghq4_0;
	wire w_dff_A_cqIW7l3Z6_0;
	wire w_dff_A_i7h7aHMk0_0;
	wire w_dff_A_OXIsrcsI1_0;
	wire w_dff_A_Pwv98ANR5_0;
	wire w_dff_A_8V1RKfWy8_0;
	wire w_dff_A_pGQcxazk7_0;
	wire w_dff_A_qttq73nH6_0;
	wire w_dff_A_7MLCmt1f9_0;
	wire w_dff_A_A3IUWPZP3_0;
	wire w_dff_A_flv45uwV2_0;
	wire w_dff_A_8hk90B1W0_0;
	wire w_dff_A_lTONVAEu1_0;
	wire w_dff_A_BNcYI1jW3_0;
	wire w_dff_A_CTsZFhOj0_1;
	wire w_dff_A_aZStHclE5_1;
	wire w_dff_B_94FtYurF3_0;
	wire w_dff_B_dPRfy0Oi2_0;
	wire w_dff_B_s94aZ1uZ9_0;
	wire w_dff_B_e0UwjMc36_0;
	wire w_dff_A_euxpM8qG3_0;
	wire w_dff_A_uDc6K0OK8_0;
	wire w_dff_A_Xpzl2Exo1_0;
	wire w_dff_A_XEUslydH8_0;
	wire w_dff_A_zAmybL963_0;
	wire w_dff_A_WaC0xmkI5_0;
	wire w_dff_A_lZKOxCBE9_0;
	wire w_dff_A_Co4vapyC6_0;
	wire w_dff_A_U5NXQK7T8_0;
	wire w_dff_A_wl7cV57o1_0;
	wire w_dff_A_F2ypEOLn8_0;
	wire w_dff_A_vjRiOPuB4_0;
	wire w_dff_A_oAQZktvN8_0;
	wire w_dff_A_4hKiCFt56_0;
	wire w_dff_A_Tkq26vvM1_0;
	wire w_dff_A_NM4lVzEs6_0;
	wire w_dff_A_y0w11bp89_0;
	wire w_dff_A_o1lx5Zeh3_0;
	wire w_dff_A_FwWBv6J41_0;
	wire w_dff_A_PRHZWjfF4_0;
	wire w_dff_A_Og0IvzaN0_0;
	wire w_dff_A_CVbHa7rN5_0;
	wire w_dff_A_kje4BfZV4_0;
	wire w_dff_A_JlmQPkRc7_0;
	wire w_dff_A_7Z8y3gVK5_0;
	wire w_dff_A_Azx8s1LO1_0;
	wire w_dff_B_RoMW8FnH0_1;
	wire w_dff_B_HtIDmsE94_1;
	wire w_dff_B_tAdIrQVR3_1;
	wire w_dff_B_CUo1k0AK5_1;
	wire w_dff_B_4wmQmU9N4_1;
	wire w_dff_A_N9RnvfVd9_0;
	wire w_dff_A_v5evyWm53_0;
	wire w_dff_A_OLtuKuaT3_0;
	wire w_dff_A_yjadT7ge8_0;
	wire w_dff_B_BfUpeLkb6_1;
	wire w_dff_B_bDjw6hKi6_1;
	wire w_dff_B_PRYKRpCi3_1;
	wire w_dff_B_LcjHbqcO6_1;
	wire w_dff_B_ahmtxd9L6_0;
	wire w_dff_B_UUwDZErp8_0;
	wire w_dff_B_kYUNMXF78_0;
	wire w_dff_A_qedJcAie1_0;
	wire w_dff_A_5xI6FYCb3_0;
	wire w_dff_A_kCt4opwe3_0;
	wire w_dff_A_7hBtspxo9_0;
	wire w_dff_A_PK1iZVts9_0;
	wire w_dff_A_WKMAoyGh9_0;
	wire w_dff_A_GEBICV0d9_0;
	wire w_dff_A_xxkv2tFz2_0;
	wire w_dff_A_OcNDm2Cr7_0;
	wire w_dff_A_amCOZp3N3_0;
	wire w_dff_B_kmbGbOWT9_1;
	wire w_dff_B_xONieWA89_1;
	wire w_dff_A_45LdLgW39_0;
	wire w_dff_B_16gvVIQX6_0;
	wire w_dff_B_dqwQiNEy2_0;
	wire w_dff_B_4tnmKcOD0_0;
	wire w_dff_A_51j4moIv4_0;
	wire w_dff_A_IGXwJl4N5_0;
	wire w_dff_A_BjmicdfJ7_0;
	wire w_dff_A_SXsHS5Nr3_0;
	wire w_dff_A_Im4Zx6Q98_0;
	wire w_dff_A_pcrO7N6p0_0;
	wire w_dff_A_Kp35cWIA9_0;
	wire w_dff_A_rzK6xVI06_0;
	wire w_dff_A_HijxTHh74_0;
	wire w_dff_A_pqUeLYjz8_0;
	wire w_dff_A_rj2cDQlh2_0;
	wire w_dff_A_gspv3eSZ3_0;
	wire w_dff_A_OEAQYrDn7_0;
	wire w_dff_A_kNaO7n3e3_0;
	wire w_dff_A_sO1JVLwy0_0;
	wire w_dff_A_BCX9q4bR9_0;
	wire w_dff_A_qru0Po659_0;
	wire w_dff_A_JrGztQ1P5_0;
	wire w_dff_A_ygsYRx3b7_0;
	wire w_dff_B_mMGdF3hJ9_2;
	wire w_dff_B_j8uXlFgC4_2;
	wire w_dff_B_ElnPzp5u5_2;
	wire w_dff_B_sXxwHUdg3_2;
	wire w_dff_B_ZzIRq4707_2;
	wire w_dff_B_xxngIuti1_2;
	wire w_dff_B_y1WVhjcL2_2;
	wire w_dff_B_y6fsy1og2_2;
	wire w_dff_B_tCHJSG9R8_2;
	wire w_dff_B_vPY4wFJg5_2;
	wire w_dff_A_9ctAOboP5_0;
	wire w_dff_A_Sgezy1ZD9_0;
	wire w_dff_A_wNHs7BF89_0;
	wire w_dff_A_K7qbLHhz0_0;
	wire w_dff_A_JwycmPio6_0;
	wire w_dff_A_NjnZNVek5_0;
	wire w_dff_A_N7OVrmsV2_0;
	wire w_dff_A_6ukVAaVQ2_0;
	wire w_dff_A_fMMmZkVI5_1;
	wire w_dff_A_ErzZilkO7_1;
	wire w_dff_A_7HH9ZPhQ7_0;
	wire w_dff_A_G7dKXof11_0;
	wire w_dff_A_zN5Gn6sK1_0;
	wire w_dff_A_H3mov8WQ6_0;
	wire w_dff_A_4B4Ax9XZ3_0;
	wire w_dff_A_3igUQjgO4_0;
	wire w_dff_A_u46OFi9Y9_0;
	wire w_dff_A_5SMsCezM6_0;
	wire w_dff_A_gmRkcWga9_0;
	wire w_dff_B_0cKDbo398_2;
	wire w_dff_B_hK7q5ME77_2;
	wire w_dff_B_V9hL6yDC8_2;
	wire w_dff_B_Hr3aWMtA7_2;
	wire w_dff_B_2xp4turu3_2;
	wire w_dff_A_IemfyM1A4_0;
	wire w_dff_A_h0YWiSR97_0;
	wire w_dff_A_TRtyb1yV4_0;
	wire w_dff_A_D9worTUj9_0;
	wire w_dff_A_Ha33DfY80_0;
	wire w_dff_A_Ss42PQcG9_0;
	wire w_dff_A_PRuzpXi84_0;
	wire w_dff_A_NxZ1ansZ3_0;
	wire w_dff_A_YO0lsnOw4_0;
	wire w_dff_A_Mij1yVR26_0;
	wire w_dff_A_YrPtC6Qu3_0;
	wire w_dff_A_98gxp4xM3_0;
	wire w_dff_A_ThHCmN9U9_1;
	wire w_dff_B_PfcDVYKc0_2;
	wire w_dff_B_ngZQ1Hzr1_2;
	wire w_dff_B_AvNIJiip3_2;
	wire w_dff_A_gRzdTXiH8_0;
	wire w_dff_A_60aJI0iE4_0;
	wire w_dff_A_slz6LnE38_0;
	wire w_dff_A_y5QS8XdQ4_0;
	wire w_dff_A_rkrCP9Nh7_0;
	wire w_dff_A_DBLhnoT00_0;
	wire w_dff_A_687nKNvu5_0;
	wire w_dff_A_Dv6BYRCd0_0;
	wire w_dff_A_eS3giYuP3_0;
	wire w_dff_A_qZrV8PM09_0;
	wire w_dff_A_F46ApbvD1_0;
	wire w_dff_A_6uo0edn53_0;
	wire w_dff_A_hCQ3erfp1_0;
	wire w_dff_A_OqN5NvHD9_0;
	wire w_dff_A_01WeINRc4_1;
	wire w_dff_A_0zNXGn6v8_1;
	wire w_dff_A_FY84Pajv3_1;
	wire w_dff_A_PIFyp6Mc1_1;
	wire w_dff_B_dh5i1UYv0_3;
	wire w_dff_B_Mvf6uajc4_3;
	wire w_dff_B_LLA56UmP6_3;
	wire w_dff_B_Dq1UPj7x4_3;
	wire w_dff_B_2zO58puS2_3;
	wire w_dff_A_stysf4x63_0;
	wire w_dff_A_ZzbkiKXP8_0;
	wire w_dff_A_qDqggfUI9_0;
	wire w_dff_A_RgXeAOyg4_1;
	wire w_dff_A_gjPjgQxL4_1;
	wire w_dff_A_e5jZYph45_1;
	wire w_dff_A_5T9DzNF45_1;
	wire w_dff_A_E9EqQVzh5_1;
	wire w_dff_A_Xg4AYU0B8_1;
	wire w_dff_A_lB43AEcG3_1;
	wire w_dff_A_HLQlrUyS4_2;
	wire w_dff_A_VRX6WUSF8_2;
	wire w_dff_A_I4sHbNO93_2;
	wire w_dff_A_ae1AmbqQ3_2;
	wire w_dff_A_1dAyMAjO7_2;
	wire w_dff_A_0SmGn8rt8_2;
	wire w_dff_A_Ys6RiXrh8_2;
	wire w_dff_A_N5aIXP5K9_0;
	wire w_dff_A_QfhYA8MQ7_0;
	wire w_dff_A_TADIeDG23_0;
	wire w_dff_A_GS2qVlTL6_0;
	wire w_dff_A_Esef1Cy66_0;
	wire w_dff_A_qNSIVEWK5_0;
	wire w_dff_A_NQYZ3OtY0_0;
	wire w_dff_A_AuCjO2Rd0_0;
	wire w_dff_A_rzcpK0X44_1;
	wire w_dff_A_RveaSCQI7_1;
	wire w_dff_A_lcaJCISS7_1;
	wire w_dff_A_Q5I9TeQr4_1;
	wire w_dff_B_iHX2EVeZ1_3;
	wire w_dff_B_mrxKIk5a2_3;
	wire w_dff_B_diEUpV051_3;
	wire w_dff_B_WzroyfKe4_3;
	wire w_dff_B_2BcIh0H47_3;
	wire w_dff_A_KCWSiRUj0_0;
	wire w_dff_A_jdfQKXCQ2_0;
	wire w_dff_A_K5bHggug5_0;
	wire w_dff_A_BSIq8CKJ4_1;
	wire w_dff_A_1LQ596uY6_1;
	wire w_dff_A_74lpbGHW9_1;
	wire w_dff_A_lzaRgxEL0_1;
	wire w_dff_A_LmwynoSP5_1;
	wire w_dff_A_PARIs3hI1_1;
	wire w_dff_A_6CSFh7d00_1;
	wire w_dff_A_TOho2NGc7_2;
	wire w_dff_A_0Hj1w6ek6_2;
	wire w_dff_A_HyRLz8mU1_2;
	wire w_dff_A_QV749GuN9_2;
	wire w_dff_A_wEc8Mubu0_2;
	wire w_dff_A_7xqCXz1e3_2;
	wire w_dff_A_KwcRjYcX8_2;
	wire w_dff_A_saQb2HaH3_1;
	wire w_dff_A_XvdXSowH1_1;
	wire w_dff_A_KKGaIIYi5_1;
	wire w_dff_A_w7DTeoif4_1;
	wire w_dff_A_klqXxfI94_0;
	wire w_dff_A_t254wNan5_0;
	wire w_dff_A_SsooMSsU0_0;
	wire w_dff_A_k4Q3J28A3_0;
	wire w_dff_A_Zie9ZKbO8_0;
	wire w_dff_A_uKQ7X8Ye8_0;
	wire w_dff_A_QBSlD7Dg1_0;
	wire w_dff_B_wT6b7cE44_1;
	wire w_dff_B_9j3xKf2N8_1;
	wire w_dff_B_z3JBK7ly4_1;
	wire w_dff_B_Prui9E6n3_1;
	wire w_dff_B_m8JfDSuB2_1;
	wire w_dff_A_1ux9T1S57_0;
	wire w_dff_A_qPJ96Qa95_0;
	wire w_dff_A_HTvPTl7u9_0;
	wire w_dff_A_ILbgMFZF7_0;
	wire w_dff_A_bvwyD8wS4_0;
	wire w_dff_A_nc9zCKgV8_0;
	wire w_dff_A_DqS6Uenx5_0;
	wire w_dff_A_nCUDPzqM2_1;
	wire w_dff_A_etTlYGfi6_1;
	wire w_dff_A_EYMhh2NP2_1;
	wire w_dff_A_2AgsyYxV7_0;
	wire w_dff_A_UYDvcHSI1_0;
	wire w_dff_A_LXsqiYb71_0;
	wire w_dff_A_K5gZdYiz0_0;
	wire w_dff_A_o1CtH3px7_0;
	wire w_dff_A_6GEmcsxw8_0;
	wire w_dff_A_rPGBybKv5_0;
	wire w_dff_A_wqcMWBRI4_0;
	wire w_dff_A_3KiuoKLP4_0;
	wire w_dff_A_PeqWGNTD6_0;
	wire w_dff_A_F8LbHkJN7_0;
	wire w_dff_A_0HDFWRb66_2;
	wire w_dff_A_fppVYlUd0_2;
	wire w_dff_A_9REwY6lZ9_2;
	wire w_dff_A_kShLKGpb9_2;
	wire w_dff_A_7uBotQ7w8_2;
	wire w_dff_A_ZMC09e0a7_2;
	wire w_dff_A_GrXrPVvO1_0;
	wire w_dff_A_zXE8161e9_0;
	wire w_dff_A_kcZW8rLt0_0;
	wire w_dff_A_Zypb9wwg6_0;
	wire w_dff_A_Pm7bGHyd0_0;
	wire w_dff_A_fdhJtzY19_0;
	wire w_dff_A_oXRlq6rw9_0;
	wire w_dff_A_CDO7FLDy4_0;
	wire w_dff_B_9AEKi8Wd3_2;
	wire w_dff_B_n9yB6g0j6_2;
	wire w_dff_B_sc1awKeY9_2;
	wire w_dff_B_i7erxtH59_2;
	wire w_dff_B_Vyv08kLF5_2;
	wire w_dff_A_VSbvciKf9_0;
	wire w_dff_A_FaB9VHLX3_0;
	wire w_dff_A_Ygu4L3Fl5_0;
	wire w_dff_A_upJ1DuWE0_0;
	wire w_dff_A_uADjZGxX3_0;
	wire w_dff_A_EkgfeO7E3_0;
	wire w_dff_A_B9xrlfVz5_0;
	wire w_dff_A_nsrhvbI39_1;
	wire w_dff_A_QoTXlDAs2_1;
	wire w_dff_A_R0XfIb7R3_1;
	wire w_dff_B_WrgAAFQT6_1;
	wire w_dff_B_L4gTz73F1_1;
	wire w_dff_B_KmI86kS49_1;
	wire w_dff_B_8FQ5nRby9_1;
	wire w_dff_B_SxfERUy20_1;
	wire w_dff_A_LmBsVYOJ1_0;
	wire w_dff_A_vdXwpCaN8_0;
	wire w_dff_A_YjA6dPWN9_0;
	wire w_dff_A_Q7oYwNKj6_1;
	wire w_dff_A_nqjCgffJ3_1;
	wire w_dff_A_ldZQdspU7_1;
	wire w_dff_A_MJd0lSQh5_1;
	wire w_dff_A_u5QpBoZE8_1;
	wire w_dff_A_PFOYwTxd2_1;
	wire w_dff_A_sIDebUwH7_1;
	wire w_dff_A_BnZ8GJYy9_0;
	wire w_dff_A_SPrxYeus6_0;
	wire w_dff_A_tJ2kkDH47_0;
	wire w_dff_A_Ka4lySTd9_0;
	wire w_dff_A_KxULQEaE2_0;
	wire w_dff_A_Px12xE5V5_0;
	wire w_dff_A_pFsUduFA4_0;
	wire w_dff_A_PUtd6XR36_0;
	wire w_dff_B_INznXfhf6_2;
	wire w_dff_B_MiTTpgiV0_2;
	wire w_dff_B_7f13l2KJ8_2;
	wire w_dff_B_2AkHVdqx1_2;
	wire w_dff_B_tHKxWh0D8_2;
	wire w_dff_A_TvXMT8YZ3_0;
	wire w_dff_A_zezalJ4X7_0;
	wire w_dff_A_goJCiRP38_0;
	wire w_dff_A_Tt5DhScb6_0;
	wire w_dff_A_os6HbrYI5_0;
	wire w_dff_A_6WhEq6Vx3_0;
	wire w_dff_A_KxQ4NtnU9_0;
	wire w_dff_A_WOWvNLkQ1_1;
	wire w_dff_A_KZWlUtOU4_1;
	wire w_dff_A_kYYK6bRS4_1;
	wire w_dff_A_MyYSfVuL7_0;
	wire w_dff_A_kqsKzx969_0;
	wire w_dff_A_PtH4u72W1_0;
	wire w_dff_A_zBbLDxvQ0_0;
	wire w_dff_B_LNRer4O56_1;
	wire w_dff_A_bG27XOGL8_0;
	wire w_dff_A_v4vcAIMn0_0;
	wire w_dff_A_WlB0py4B6_0;
	wire w_dff_A_SAaoQR5h7_0;
	wire w_dff_A_fjnOabEE3_0;
	wire w_dff_A_4RWu16j10_0;
	wire w_dff_A_EV2sJo6k3_0;
	wire w_dff_A_gaki3A8c6_0;
	wire w_dff_A_7D03RUXx3_0;
	wire w_dff_A_xsn42MhW1_0;
	wire w_dff_A_bZ6zyFUp1_0;
	wire w_dff_A_YTuRB6Gf8_0;
	wire w_dff_A_JUJu95Zx7_0;
	wire w_dff_A_LR7YmvsM5_0;
	wire w_dff_B_A8pZF0mD5_0;
	wire w_dff_A_QNhJK7rH4_0;
	wire w_dff_A_jNCouyL34_0;
	wire w_dff_A_H3BVJhYs1_0;
	wire w_dff_A_xGrMqJsJ5_0;
	wire w_dff_A_Xagkc7CY7_0;
	wire w_dff_A_Ta83EDWr3_0;
	wire w_dff_A_vJO7fpZQ4_0;
	wire w_dff_A_IlkKZJFh0_0;
	wire w_dff_A_AXMTzXvf2_0;
	wire w_dff_A_EtBe2ehS1_0;
	wire w_dff_A_AtdiSjA13_0;
	wire w_dff_A_A2XPuU905_0;
	wire w_dff_A_hSCnyLzu4_0;
	wire w_dff_A_JceNb8cT8_0;
	wire w_dff_A_0K2V6HLY3_0;
	wire w_dff_B_ctJnivF36_2;
	wire w_dff_B_rHP0cAYc5_2;
	wire w_dff_B_JCPlyy7P0_2;
	wire w_dff_B_xpLdf9kD2_2;
	wire w_dff_B_qb1tUmSa4_2;
	wire w_dff_A_ciQpGTVL6_0;
	wire w_dff_A_9bMwNqAm2_0;
	wire w_dff_A_GK8arUIn6_0;
	wire w_dff_A_VSeaxf1k8_0;
	wire w_dff_A_dcHtOUie7_0;
	wire w_dff_A_QVr0zDOh5_0;
	wire w_dff_A_oxSmCrPp1_0;
	wire w_dff_A_EK9hzRGP0_1;
	wire w_dff_A_WTrN4iro9_1;
	wire w_dff_A_r9UuOjSk8_1;
	wire w_dff_A_N7fbQPkr9_1;
	wire w_dff_A_aTbF4cHM8_1;
	wire w_dff_A_FWcx9C3Y3_1;
	wire w_dff_A_1ipRx2DE7_1;
	wire w_dff_A_LnOkSJ5j2_1;
	wire w_dff_A_BxmwBAfp9_0;
	wire w_dff_A_AwL1qWK18_0;
	wire w_dff_A_otO67G9I2_0;
	wire w_dff_A_mpTh07YM3_0;
	wire w_dff_A_QeiAwPo49_0;
	wire w_dff_A_ackFX2VS9_2;
	wire w_dff_A_7tHy1G102_0;
	wire w_dff_A_qVT9keJC1_0;
	wire w_dff_A_yODH62IO5_0;
	wire w_dff_A_cXNwIErP0_0;
	wire w_dff_A_3nvwjmDD0_0;
	wire w_dff_A_8Q9aDmsZ4_0;
	wire w_dff_A_S9cH5ASg8_1;
	wire w_dff_A_APOtbspc7_0;
	wire w_dff_A_f3Xi4Qwd0_0;
	wire w_dff_A_aVFwHXl16_0;
	wire w_dff_A_Gis9XQrO3_0;
	wire w_dff_A_v7VY6Ps68_0;
	wire w_dff_A_mK9E1x6N7_0;
	wire w_dff_A_spUQlFXn1_1;
	wire w_dff_A_EHE0HbeY6_0;
	wire w_dff_A_ykbCGbil4_0;
	wire w_dff_A_HcPEVzBh4_0;
	wire w_dff_A_qQqlwDc46_0;
	wire w_dff_A_ykuSPxPC3_0;
	wire w_dff_A_yhPEyTC79_2;
	wire w_dff_A_S9UKB6UZ7_0;
	wire w_dff_A_Ve4z2LmU5_0;
	wire w_dff_A_VTN8bKRk0_0;
	wire w_dff_A_Gos5lcXw0_0;
	wire w_dff_A_qQ3Kzdjq6_0;
	wire w_dff_A_fFAyDfkg4_0;
	wire w_dff_A_ccVj2SPm1_1;
	wire w_dff_A_gr0LHtEM7_0;
	wire w_dff_A_jlg59BuU9_0;
	wire w_dff_A_AV8qV57X8_0;
	wire w_dff_A_iS2sVosO3_0;
	wire w_dff_A_EIPkYlR64_0;
	wire w_dff_A_x97kb6s77_2;
	wire w_dff_A_HH5XMtOD5_0;
	wire w_dff_A_mt9U9CVX7_0;
	wire w_dff_A_cxvNp9Vi8_0;
	wire w_dff_A_yHbq8kSS5_0;
	wire w_dff_A_ZHctAwEN9_0;
	wire w_dff_A_iwJkMMKv3_0;
	wire w_dff_A_bZE7w3OJ6_1;
	wire w_dff_A_KWD4Dwzu7_0;
	wire w_dff_A_6iCdptVu6_0;
	wire w_dff_A_2Ov9wwNx0_0;
	wire w_dff_A_3WsiLQ5r3_0;
	wire w_dff_A_cSh138lx0_0;
	wire w_dff_A_mNTfqqc63_2;
	wire w_dff_A_I73cHgpi9_0;
	wire w_dff_A_fHB4XJih3_0;
	wire w_dff_A_KbVKz9Mn1_0;
	wire w_dff_A_EuZn7Eiy6_0;
	wire w_dff_A_8WY9Fg2k9_0;
	wire w_dff_A_hJhMiXj88_0;
	wire w_dff_A_kRPglyTL6_1;
	wire w_dff_A_WyQy5OLV6_0;
	wire w_dff_A_7ewoJsAz5_0;
	wire w_dff_A_pv6JlPPU4_0;
	wire w_dff_A_bjbEQ63G7_1;
	wire w_dff_A_4XfPiDUQ5_1;
	wire w_dff_A_KwYcxXwP8_2;
	wire w_dff_A_UyYShGjK6_0;
	wire w_dff_A_pq1DDwcH6_0;
	wire w_dff_A_Q2VAeA2m4_1;
	wire w_dff_A_XMo7uwTd9_0;
	wire w_dff_A_AsJ4Gvp40_0;
	wire w_dff_A_p1w3Gei79_0;
	wire w_dff_A_syGEktSd7_0;
	wire w_dff_A_tQeqhSFR8_0;
	wire w_dff_A_RuHE0NNv0_2;
	wire w_dff_A_xc9obCm23_0;
	wire w_dff_A_813ZqyV73_0;
	wire w_dff_A_j4wWfytA0_0;
	wire w_dff_A_9GXswcgi6_0;
	wire w_dff_A_0Vl9meXi0_0;
	wire w_dff_A_Ds2KCWjB4_0;
	wire w_dff_A_zx77paec5_1;
	wire w_dff_A_4SCBLVVK6_1;
	wire w_dff_A_tH6gJrwO5_0;
	wire w_dff_A_fgwqndJK0_1;
	wire w_dff_A_S0Zpzih35_1;
	wire w_dff_A_NTnB0OF15_1;
	wire w_dff_A_Nj3ox54D2_1;
	wire w_dff_A_68cmWWIi9_1;
	wire w_dff_A_xeQ0w4hR0_2;
	wire w_dff_A_jXWkyhs01_0;
	wire w_dff_A_SPilwwnD3_0;
	wire w_dff_A_u7R7yUNg8_0;
	wire w_dff_A_PDTzFAbJ0_0;
	wire w_dff_A_KKzrVnWZ8_0;
	wire w_dff_A_V77Qgtx09_0;
	wire w_dff_A_1TIcpTGE4_0;
	wire w_dff_A_ofGCrke68_0;
	wire w_dff_A_cs9ejUyk0_0;
	wire w_dff_A_mGFoBZuA1_0;
	wire w_dff_A_eO7y5zfd3_0;
	wire w_dff_A_nJ8mA2cN9_0;
	wire w_dff_A_UAZ4UGCm2_0;
	wire w_dff_A_dZ1WiuOi5_2;
	wire w_dff_A_BZGd1Zbo3_1;
	wire w_dff_A_2lFAT6Du2_1;
	wire w_dff_A_HcHjp5KW6_1;
	wire w_dff_A_kLajnnKD6_1;
	wire w_dff_A_DMqNZfW33_1;
	wire w_dff_A_HVDqM4J37_1;
	wire w_dff_A_ITHjWEV05_1;
	wire w_dff_A_ByEd35Mx2_1;
	jnot g000(.din(w_G76gat_0[1]),.dout(n43),.clk(gclk));
	jand g001(.dina(w_G82gat_0[2]),.dinb(w_n43_0[1]),.dout(n44),.clk(gclk));
	jnot g002(.din(w_G24gat_0[1]),.dout(n45),.clk(gclk));
	jand g003(.dina(w_G30gat_0[1]),.dinb(n45),.dout(n46),.clk(gclk));
	jnot g004(.din(w_G11gat_0[2]),.dout(n47),.clk(gclk));
	jand g005(.dina(w_G17gat_0[2]),.dinb(w_n47_0[1]),.dout(n48),.clk(gclk));
	jcb g006(.dina(n48),.dinb(n46),.dout(n49));
	jcb g007(.dina(n49),.dinb(w_n44_0[1]),.dout(n50));
	jnot g008(.din(w_G37gat_0[2]),.dout(n51),.clk(gclk));
	jand g009(.dina(w_G43gat_1[1]),.dinb(n51),.dout(n52),.clk(gclk));
	jnot g010(.din(w_G63gat_0[2]),.dout(n53),.clk(gclk));
	jand g011(.dina(w_G69gat_0[2]),.dinb(w_n53_0[1]),.dout(n54),.clk(gclk));
	jcb g012(.dina(n54),.dinb(w_n52_0[1]),.dout(n55));
	jnot g013(.din(w_G102gat_0[2]),.dout(n56),.clk(gclk));
	jand g014(.dina(w_G108gat_0[2]),.dinb(w_n56_0[1]),.dout(n57),.clk(gclk));
	jnot g015(.din(w_G50gat_0[2]),.dout(n58),.clk(gclk));
	jand g016(.dina(w_G56gat_0[2]),.dinb(w_n58_0[1]),.dout(n59),.clk(gclk));
	jcb g017(.dina(n59),.dinb(n57),.dout(n60));
	jnot g018(.din(w_G89gat_0[2]),.dout(n61),.clk(gclk));
	jand g019(.dina(w_G95gat_0[2]),.dinb(w_n61_0[1]),.dout(n62),.clk(gclk));
	jnot g020(.din(w_G1gat_0[2]),.dout(n63),.clk(gclk));
	jand g021(.dina(w_G4gat_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jcb g022(.dina(n64),.dinb(n62),.dout(n65));
	jcb g023(.dina(n65),.dinb(n60),.dout(n66));
	jcb g024(.dina(n66),.dinb(n55),.dout(n67));
	jcb g025(.dina(n67),.dinb(n50),.dout(G223gat_fa_));
	jnot g026(.din(w_G112gat_0[2]),.dout(n69),.clk(gclk));
	jnot g027(.din(w_n44_0[0]),.dout(n70),.clk(gclk));
	jnot g028(.din(w_G30gat_0[0]),.dout(n71),.clk(gclk));
	jcb g029(.dina(w_n71_0[1]),.dinb(w_G24gat_0[0]),.dout(n72));
	jnot g030(.din(w_G17gat_0[1]),.dout(n73),.clk(gclk));
	jcb g031(.dina(w_n73_0[1]),.dinb(w_G11gat_0[1]),.dout(n74));
	jand g032(.dina(n74),.dinb(w_n72_0[1]),.dout(n75),.clk(gclk));
	jand g033(.dina(w_dff_B_A8pZF0mD5_0),.dinb(n70),.dout(n76),.clk(gclk));
	jnot g034(.din(w_G43gat_1[0]),.dout(n77),.clk(gclk));
	jcb g035(.dina(w_n77_0[1]),.dinb(w_G37gat_0[1]),.dout(n78));
	jnot g036(.din(w_G69gat_0[1]),.dout(n79),.clk(gclk));
	jcb g037(.dina(w_n79_0[1]),.dinb(w_G63gat_0[1]),.dout(n80));
	jand g038(.dina(n80),.dinb(w_n78_0[1]),.dout(n81),.clk(gclk));
	jnot g039(.din(w_G108gat_0[1]),.dout(n82),.clk(gclk));
	jcb g040(.dina(w_n82_0[1]),.dinb(w_G102gat_0[1]),.dout(n83));
	jnot g041(.din(w_G56gat_0[1]),.dout(n84),.clk(gclk));
	jcb g042(.dina(w_n84_0[1]),.dinb(w_G50gat_0[1]),.dout(n85));
	jand g043(.dina(n85),.dinb(n83),.dout(n86),.clk(gclk));
	jnot g044(.din(w_G95gat_0[1]),.dout(n87),.clk(gclk));
	jcb g045(.dina(w_n87_0[1]),.dinb(w_G89gat_0[1]),.dout(n88));
	jnot g046(.din(w_G4gat_0[1]),.dout(n89),.clk(gclk));
	jcb g047(.dina(w_n89_0[1]),.dinb(w_G1gat_0[1]),.dout(n90));
	jand g048(.dina(n90),.dinb(n88),.dout(n91),.clk(gclk));
	jand g049(.dina(n91),.dinb(n86),.dout(n92),.clk(gclk));
	jand g050(.dina(n92),.dinb(w_dff_B_LNRer4O56_1),.dout(n93),.clk(gclk));
	jand g051(.dina(n93),.dinb(n76),.dout(n94),.clk(gclk));
	jcb g052(.dina(w_n94_4[1]),.dinb(w_n56_0[0]),.dout(n95));
	jand g053(.dina(n95),.dinb(w_G108gat_0[0]),.dout(n96),.clk(gclk));
	jand g054(.dina(w_n96_0[1]),.dinb(w_n69_0[1]),.dout(n97),.clk(gclk));
	jnot g055(.din(w_G8gat_0[2]),.dout(n98),.clk(gclk));
	jcb g056(.dina(w_n94_4[0]),.dinb(w_n63_0[0]),.dout(n99));
	jand g057(.dina(n99),.dinb(w_G4gat_0[0]),.dout(n100),.clk(gclk));
	jand g058(.dina(w_n100_0[1]),.dinb(w_n98_0[1]),.dout(n101),.clk(gclk));
	jcb g059(.dina(n101),.dinb(n97),.dout(n102));
	jnot g060(.din(w_G99gat_0[2]),.dout(n103),.clk(gclk));
	jcb g061(.dina(w_n94_3[2]),.dinb(w_n61_0[0]),.dout(n104));
	jand g062(.dina(n104),.dinb(w_G95gat_0[0]),.dout(n105),.clk(gclk));
	jand g063(.dina(n105),.dinb(w_dff_B_SxfERUy20_1),.dout(n106),.clk(gclk));
	jnot g064(.din(w_G73gat_0[2]),.dout(n107),.clk(gclk));
	jcb g065(.dina(w_n94_3[1]),.dinb(w_n53_0[0]),.dout(n108));
	jand g066(.dina(n108),.dinb(w_G69gat_0[0]),.dout(n109),.clk(gclk));
	jand g067(.dina(w_n109_0[1]),.dinb(w_n107_0[1]),.dout(n110),.clk(gclk));
	jcb g068(.dina(n110),.dinb(n106),.dout(n111));
	jcb g069(.dina(n111),.dinb(n102),.dout(n112));
	jxor g070(.dina(w_n94_3[0]),.dinb(w_n72_0[0]),.dout(n113),.clk(gclk));
	jcb g071(.dina(n113),.dinb(w_n71_0[0]),.dout(n114));
	jcb g072(.dina(w_n114_0[2]),.dinb(w_G34gat_0[2]),.dout(n115));
	jnot g073(.din(w_n115_0[1]),.dout(n116),.clk(gclk));
	jnot g074(.din(w_G60gat_0[2]),.dout(n117),.clk(gclk));
	jcb g075(.dina(w_n94_2[2]),.dinb(w_n58_0[0]),.dout(n118));
	jand g076(.dina(n118),.dinb(w_G56gat_0[0]),.dout(n119),.clk(gclk));
	jand g077(.dina(w_n119_0[1]),.dinb(w_dff_B_m8JfDSuB2_1),.dout(n120),.clk(gclk));
	jxor g078(.dina(w_n94_2[1]),.dinb(w_n52_0[0]),.dout(n121),.clk(gclk));
	jnot g079(.din(w_G47gat_0[1]),.dout(n122),.clk(gclk));
	jand g080(.dina(n122),.dinb(w_G43gat_0[2]),.dout(n123),.clk(gclk));
	jand g081(.dina(w_n123_0[1]),.dinb(w_n121_0[1]),.dout(n124),.clk(gclk));
	jcb g082(.dina(n124),.dinb(n120),.dout(n125));
	jnot g083(.din(w_G86gat_1[1]),.dout(n126),.clk(gclk));
	jcb g084(.dina(w_n94_2[0]),.dinb(w_n43_0[0]),.dout(n127));
	jand g085(.dina(n127),.dinb(w_G82gat_0[1]),.dout(n128),.clk(gclk));
	jand g086(.dina(w_n128_0[1]),.dinb(w_n126_0[2]),.dout(n129),.clk(gclk));
	jnot g087(.din(w_G21gat_1[1]),.dout(n130),.clk(gclk));
	jcb g088(.dina(w_n94_1[2]),.dinb(w_n47_0[0]),.dout(n131));
	jand g089(.dina(n131),.dinb(w_G17gat_0[0]),.dout(n132),.clk(gclk));
	jand g090(.dina(w_n132_0[1]),.dinb(w_n130_0[2]),.dout(n133),.clk(gclk));
	jcb g091(.dina(n133),.dinb(n129),.dout(n134));
	jcb g092(.dina(n134),.dinb(n125),.dout(n135));
	jcb g093(.dina(n135),.dinb(n116),.dout(n136));
	jcb g094(.dina(n136),.dinb(n112),.dout(G329gat_fa_));
	jand g095(.dina(w_G223gat_3[1]),.dinb(w_G89gat_0[0]),.dout(n138),.clk(gclk));
	jcb g096(.dina(n138),.dinb(w_n87_0[0]),.dout(n139));
	jand g097(.dina(w_G329gat_6),.dinb(w_G99gat_0[1]),.dout(n140),.clk(gclk));
	jcb g098(.dina(n140),.dinb(w_n139_0[1]),.dout(n141));
	jcb g099(.dina(w_n141_0[1]),.dinb(w_G105gat_0[1]),.dout(n142));
	jnot g100(.din(w_n142_0[1]),.dout(n143),.clk(gclk));
	jand g101(.dina(w_G223gat_3[0]),.dinb(w_G50gat_0[0]),.dout(n144),.clk(gclk));
	jcb g102(.dina(n144),.dinb(w_n84_0[0]),.dout(n145));
	jcb g103(.dina(w_n145_0[1]),.dinb(w_G60gat_0[1]),.dout(n146));
	jand g104(.dina(w_G329gat_5[2]),.dinb(w_n146_0[1]),.dout(n147),.clk(gclk));
	jnot g105(.din(w_n147_0[1]),.dout(n148),.clk(gclk));
	jnot g106(.din(w_G66gat_0[1]),.dout(n150),.clk(gclk));
	jand g107(.dina(w_n119_0[0]),.dinb(w_n150_0[1]),.dout(n151),.clk(gclk));
	jand g108(.dina(w_n151_0[1]),.dinb(n148),.dout(n153),.clk(gclk));
	jnot g109(.din(w_G79gat_0[1]),.dout(n154),.clk(gclk));
	jand g110(.dina(w_G223gat_2[2]),.dinb(w_G102gat_0[0]),.dout(n155),.clk(gclk));
	jcb g111(.dina(n155),.dinb(w_n82_0[0]),.dout(n156));
	jcb g112(.dina(w_n156_0[1]),.dinb(w_G112gat_0[1]),.dout(n157));
	jand g113(.dina(w_G223gat_2[1]),.dinb(w_G1gat_0[0]),.dout(n158),.clk(gclk));
	jcb g114(.dina(n158),.dinb(w_n89_0[0]),.dout(n159));
	jcb g115(.dina(w_n159_0[1]),.dinb(w_G8gat_0[1]),.dout(n160));
	jand g116(.dina(n160),.dinb(n157),.dout(n161),.clk(gclk));
	jcb g117(.dina(w_n139_0[0]),.dinb(w_G99gat_0[0]),.dout(n162));
	jand g118(.dina(w_G223gat_2[0]),.dinb(w_G63gat_0[0]),.dout(n163),.clk(gclk));
	jcb g119(.dina(n163),.dinb(w_n79_0[0]),.dout(n164));
	jcb g120(.dina(w_n164_0[1]),.dinb(w_G73gat_0[1]),.dout(n165));
	jand g121(.dina(n165),.dinb(n162),.dout(n166),.clk(gclk));
	jand g122(.dina(n166),.dinb(n161),.dout(n167),.clk(gclk));
	jxor g123(.dina(w_n94_1[1]),.dinb(w_n78_0[0]),.dout(n168),.clk(gclk));
	jnot g124(.din(w_n123_0[0]),.dout(n169),.clk(gclk));
	jcb g125(.dina(w_dff_B_4tnmKcOD0_0),.dinb(n168),.dout(n170));
	jand g126(.dina(w_n170_0[1]),.dinb(w_n146_0[0]),.dout(n171),.clk(gclk));
	jnot g127(.din(w_G82gat_0[0]),.dout(n172),.clk(gclk));
	jand g128(.dina(w_G223gat_1[2]),.dinb(w_G76gat_0[0]),.dout(n173),.clk(gclk));
	jcb g129(.dina(n173),.dinb(w_dff_B_xONieWA89_1),.dout(n174));
	jcb g130(.dina(w_n174_0[1]),.dinb(w_G86gat_1[0]),.dout(n175));
	jand g131(.dina(w_G223gat_1[1]),.dinb(w_G11gat_0[0]),.dout(n176),.clk(gclk));
	jcb g132(.dina(n176),.dinb(w_n73_0[0]),.dout(n177));
	jcb g133(.dina(w_n177_0[1]),.dinb(w_G21gat_1[0]),.dout(n178));
	jand g134(.dina(n178),.dinb(n175),.dout(n179),.clk(gclk));
	jand g135(.dina(w_dff_B_kYUNMXF78_0),.dinb(n171),.dout(n180),.clk(gclk));
	jand g136(.dina(n180),.dinb(w_n115_0[0]),.dout(n181),.clk(gclk));
	jand g137(.dina(n181),.dinb(w_dff_B_LcjHbqcO6_1),.dout(n182),.clk(gclk));
	jcb g138(.dina(w_n182_3[1]),.dinb(w_n107_0[0]),.dout(n183));
	jand g139(.dina(n183),.dinb(w_n109_0[0]),.dout(n184),.clk(gclk));
	jand g140(.dina(w_n184_0[1]),.dinb(w_n154_0[1]),.dout(n185),.clk(gclk));
	jcb g141(.dina(n185),.dinb(w_dff_B_4wmQmU9N4_1),.dout(n186));
	jcb g142(.dina(n186),.dinb(w_dff_B_tAdIrQVR3_1),.dout(n187));
	jand g143(.dina(w_G329gat_5[1]),.dinb(w_n170_0[0]),.dout(n188),.clk(gclk));
	jnot g144(.din(w_n188_0[1]),.dout(n189),.clk(gclk));
	jnot g145(.din(w_G53gat_0[1]),.dout(n191),.clk(gclk));
	jand g146(.dina(w_n191_0[1]),.dinb(w_G43gat_0[1]),.dout(n192),.clk(gclk));
	jand g147(.dina(w_dff_B_e0UwjMc36_0),.dinb(w_n121_0[0]),.dout(n193),.clk(gclk));
	jand g148(.dina(w_n193_0[1]),.dinb(n189),.dout(n195),.clk(gclk));
	jcb g149(.dina(w_n182_3[0]),.dinb(w_n130_0[1]),.dout(n196));
	jand g150(.dina(n196),.dinb(w_n132_0[0]),.dout(n197),.clk(gclk));
	jnot g151(.din(w_G27gat_0[1]),.dout(n198),.clk(gclk));
	jcb g152(.dina(w_G329gat_5[0]),.dinb(w_G21gat_0[2]),.dout(n199));
	jand g153(.dina(n199),.dinb(w_n198_0[1]),.dout(n200),.clk(gclk));
	jand g154(.dina(w_dff_B_RJacCCyX8_0),.dinb(w_n197_0[1]),.dout(n201),.clk(gclk));
	jcb g155(.dina(n201),.dinb(w_dff_B_JanIzsh28_1),.dout(n202));
	jcb g156(.dina(w_n182_2[2]),.dinb(w_n126_0[1]),.dout(n203));
	jand g157(.dina(n203),.dinb(w_n128_0[0]),.dout(n204),.clk(gclk));
	jnot g158(.din(w_G92gat_0[2]),.dout(n205),.clk(gclk));
	jcb g159(.dina(w_G329gat_4[2]),.dinb(w_G86gat_0[2]),.dout(n206));
	jand g160(.dina(n206),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jand g161(.dina(w_dff_B_OX8CYYjJ6_0),.dinb(w_n204_0[1]),.dout(n208),.clk(gclk));
	jnot g162(.din(w_G14gat_0[2]),.dout(n209),.clk(gclk));
	jcb g163(.dina(w_n182_2[1]),.dinb(w_n98_0[0]),.dout(n210));
	jand g164(.dina(n210),.dinb(w_n100_0[0]),.dout(n211),.clk(gclk));
	jand g165(.dina(n211),.dinb(w_dff_B_SLm6IIqn0_1),.dout(n212),.clk(gclk));
	jcb g166(.dina(n212),.dinb(n208),.dout(n213));
	jnot g167(.din(w_G34gat_0[1]),.dout(n214),.clk(gclk));
	jcb g168(.dina(w_n182_2[0]),.dinb(w_dff_B_VCU9QS1w1_1),.dout(n215));
	jnot g169(.din(w_G40gat_0[1]),.dout(n217),.clk(gclk));
	jnot g170(.din(w_n114_0[1]),.dout(n218),.clk(gclk));
	jand g171(.dina(n218),.dinb(w_n217_0[1]),.dout(n219),.clk(gclk));
	jand g172(.dina(w_n219_0[1]),.dinb(n215),.dout(n221),.clk(gclk));
	jnot g173(.din(w_G115gat_0[1]),.dout(n222),.clk(gclk));
	jcb g174(.dina(w_n182_1[2]),.dinb(w_n69_0[0]),.dout(n223));
	jand g175(.dina(n223),.dinb(w_n96_0[0]),.dout(n224),.clk(gclk));
	jand g176(.dina(w_n224_0[1]),.dinb(w_n222_0[1]),.dout(n225),.clk(gclk));
	jcb g177(.dina(n225),.dinb(w_dff_B_NfZgjlwf5_1),.dout(n226));
	jcb g178(.dina(n226),.dinb(n213),.dout(n227));
	jcb g179(.dina(n227),.dinb(n202),.dout(n228));
	jcb g180(.dina(n228),.dinb(n187),.dout(G370gat_fa_));
	jand g181(.dina(w_G329gat_4[1]),.dinb(w_G8gat_0[0]),.dout(n230),.clk(gclk));
	jcb g182(.dina(n230),.dinb(w_n159_0[0]),.dout(n231));
	jand g183(.dina(w_G370gat_2),.dinb(w_G14gat_0[1]),.dout(n232),.clk(gclk));
	jcb g184(.dina(n232),.dinb(w_n231_0[1]),.dout(n233));
	jnot g185(.din(w_n151_0[0]),.dout(n235),.clk(gclk));
	jcb g186(.dina(n235),.dinb(w_n147_0[0]),.dout(n237));
	jand g187(.dina(w_G329gat_4[0]),.dinb(w_G73gat_0[0]),.dout(n238),.clk(gclk));
	jcb g188(.dina(n238),.dinb(w_n164_0[0]),.dout(n239));
	jcb g189(.dina(n239),.dinb(w_G79gat_0[0]),.dout(n240));
	jand g190(.dina(n240),.dinb(n237),.dout(n241),.clk(gclk));
	jand g191(.dina(n241),.dinb(w_n142_0[0]),.dout(n242),.clk(gclk));
	jnot g192(.din(w_n193_0[0]),.dout(n244),.clk(gclk));
	jcb g193(.dina(n244),.dinb(w_n188_0[0]),.dout(n246));
	jand g194(.dina(w_G329gat_3[2]),.dinb(w_G21gat_0[1]),.dout(n247),.clk(gclk));
	jcb g195(.dina(n247),.dinb(w_n177_0[0]),.dout(n248));
	jand g196(.dina(w_n182_1[1]),.dinb(w_n130_0[0]),.dout(n249),.clk(gclk));
	jcb g197(.dina(n249),.dinb(w_G27gat_0[0]),.dout(n250));
	jcb g198(.dina(n250),.dinb(w_dff_B_cx9NWvkF0_1),.dout(n251));
	jand g199(.dina(n251),.dinb(w_dff_B_63L91ISR7_1),.dout(n252),.clk(gclk));
	jand g200(.dina(w_G329gat_3[1]),.dinb(w_G86gat_0[1]),.dout(n253),.clk(gclk));
	jcb g201(.dina(n253),.dinb(w_n174_0[0]),.dout(n254));
	jand g202(.dina(w_n182_1[0]),.dinb(w_n126_0[0]),.dout(n255),.clk(gclk));
	jcb g203(.dina(n255),.dinb(w_G92gat_0[1]),.dout(n256));
	jcb g204(.dina(n256),.dinb(w_n254_0[1]),.dout(n257));
	jcb g205(.dina(w_n231_0[0]),.dinb(w_G14gat_0[0]),.dout(n258));
	jand g206(.dina(w_dff_B_dBUvcGT71_0),.dinb(n257),.dout(n259),.clk(gclk));
	jand g207(.dina(w_G329gat_3[0]),.dinb(w_G34gat_0[0]),.dout(n260),.clk(gclk));
	jnot g208(.din(w_n219_0[0]),.dout(n262),.clk(gclk));
	jcb g209(.dina(n262),.dinb(w_n260_0[1]),.dout(n264));
	jand g210(.dina(w_G329gat_2[2]),.dinb(w_G112gat_0[0]),.dout(n265),.clk(gclk));
	jcb g211(.dina(n265),.dinb(w_n156_0[0]),.dout(n266));
	jcb g212(.dina(n266),.dinb(w_G115gat_0[0]),.dout(n267));
	jand g213(.dina(w_dff_B_RuLZw8Ua2_0),.dinb(n264),.dout(n268),.clk(gclk));
	jand g214(.dina(w_dff_B_q1ZvadfE8_0),.dinb(n259),.dout(n269),.clk(gclk));
	jand g215(.dina(n269),.dinb(w_dff_B_nKBhQB1W6_1),.dout(n270),.clk(gclk));
	jand g216(.dina(n270),.dinb(w_dff_B_BlhSNEHh9_1),.dout(n271),.clk(gclk));
	jcb g217(.dina(w_n271_3[1]),.dinb(w_n150_0[0]),.dout(n272));
	jand g218(.dina(w_G329gat_2[1]),.dinb(w_G60gat_0[0]),.dout(n273),.clk(gclk));
	jcb g219(.dina(n273),.dinb(w_n145_0[0]),.dout(n274));
	jnot g220(.din(w_n274_0[1]),.dout(n275),.clk(gclk));
	jand g221(.dina(w_dff_B_XTwMCCN78_0),.dinb(n272),.dout(n276),.clk(gclk));
	jcb g222(.dina(w_n271_3[0]),.dinb(w_n191_0[0]),.dout(n277));
	jand g223(.dina(w_G329gat_2[0]),.dinb(w_G47gat_0[0]),.dout(n278),.clk(gclk));
	jand g224(.dina(w_G223gat_1[0]),.dinb(w_G37gat_0[0]),.dout(n279),.clk(gclk));
	jcb g225(.dina(n279),.dinb(w_n77_0[0]),.dout(n280));
	jcb g226(.dina(w_dff_B_WZY9NVfD0_0),.dinb(n278),.dout(n281));
	jnot g227(.din(w_n281_0[1]),.dout(n282),.clk(gclk));
	jand g228(.dina(w_dff_B_huyq7yRr4_0),.dinb(n277),.dout(n283),.clk(gclk));
	jcb g229(.dina(w_n283_0[1]),.dinb(n276),.dout(n284));
	jcb g230(.dina(w_n271_2[2]),.dinb(w_n198_0[0]),.dout(n285));
	jand g231(.dina(n285),.dinb(w_n197_0[0]),.dout(n286),.clk(gclk));
	jcb g232(.dina(w_n271_2[1]),.dinb(w_n217_0[0]),.dout(n287));
	jcb g233(.dina(w_n114_0[0]),.dinb(w_n260_0[0]),.dout(n290));
	jnot g234(.din(w_n290_0[1]),.dout(n291),.clk(gclk));
	jand g235(.dina(w_dff_B_H7dSlUJY2_0),.dinb(n287),.dout(n292),.clk(gclk));
	jcb g236(.dina(n292),.dinb(w_n286_0[1]),.dout(n293));
	jcb g237(.dina(w_n293_0[1]),.dinb(n284),.dout(G430gat_fa_));
	jcb g238(.dina(w_n271_2[0]),.dinb(w_n205_0[0]),.dout(n295));
	jand g239(.dina(n295),.dinb(w_n204_0[0]),.dout(n296),.clk(gclk));
	jcb g240(.dina(w_n271_1[2]),.dinb(w_n222_0[0]),.dout(n297));
	jand g241(.dina(n297),.dinb(w_n224_0[0]),.dout(n298),.clk(gclk));
	jcb g242(.dina(n298),.dinb(w_n296_0[1]),.dout(n299));
	jnot g243(.din(w_n141_0[0]),.dout(n300),.clk(gclk));
	jnot g244(.din(w_G105gat_0[0]),.dout(n301),.clk(gclk));
	jcb g245(.dina(w_n271_1[1]),.dinb(w_dff_B_G9r9K1T88_1),.dout(n302));
	jand g246(.dina(n302),.dinb(w_dff_B_pOpfgyo86_1),.dout(n303),.clk(gclk));
	jcb g247(.dina(w_n271_1[0]),.dinb(w_n154_0[0]),.dout(n304));
	jand g248(.dina(n304),.dinb(w_n184_0[0]),.dout(n305),.clk(gclk));
	jcb g249(.dina(w_n305_0[1]),.dinb(w_n303_0[1]),.dout(n306));
	jcb g250(.dina(n306),.dinb(n299),.dout(n307));
	jcb g251(.dina(n307),.dinb(w_G430gat_0),.dout(n308));
	jand g252(.dina(n308),.dinb(w_dff_B_KumAQcfB7_1),.dout(G421gat),.clk(gclk));
	jand g253(.dina(w_G370gat_1[2]),.dinb(w_G66gat_0[0]),.dout(n310),.clk(gclk));
	jcb g254(.dina(w_n274_0[0]),.dinb(n310),.dout(n311));
	jand g255(.dina(w_G370gat_1[1]),.dinb(w_G53gat_0[0]),.dout(n312),.clk(gclk));
	jcb g256(.dina(w_n281_0[0]),.dinb(n312),.dout(n313));
	jand g257(.dina(w_n313_0[1]),.dinb(n311),.dout(n314),.clk(gclk));
	jand g258(.dina(w_n296_0[0]),.dinb(w_n314_0[1]),.dout(n315),.clk(gclk));
	jand g259(.dina(w_G370gat_1[0]),.dinb(w_G40gat_0[0]),.dout(n316),.clk(gclk));
	jcb g260(.dina(w_n290_0[0]),.dinb(n316),.dout(n317));
	jand g261(.dina(w_n305_0[0]),.dinb(w_n317_0[2]),.dout(n318),.clk(gclk));
	jand g262(.dina(n318),.dinb(w_n314_0[0]),.dout(n319),.clk(gclk));
	jcb g263(.dina(w_n319_0[1]),.dinb(w_n293_0[0]),.dout(n320));
	jcb g264(.dina(n320),.dinb(w_dff_B_DT7GTFZ78_1),.dout(G431gat));
	jand g265(.dina(w_n303_0[0]),.dinb(w_n317_0[1]),.dout(n322),.clk(gclk));
	jand g266(.dina(w_G370gat_0[2]),.dinb(w_G92gat_0[0]),.dout(n323),.clk(gclk));
	jcb g267(.dina(n323),.dinb(w_n254_0[0]),.dout(n324));
	jand g268(.dina(n324),.dinb(w_n313_0[0]),.dout(n325),.clk(gclk));
	jand g269(.dina(w_dff_B_0jpW6hqj9_0),.dinb(n322),.dout(n326),.clk(gclk));
	jand g270(.dina(w_n317_0[0]),.dinb(w_n283_0[0]),.dout(n327),.clk(gclk));
	jcb g271(.dina(n327),.dinb(w_n286_0[0]),.dout(n328));
	jcb g272(.dina(w_dff_B_wi0W0TXf6_0),.dinb(w_n319_0[0]),.dout(n329));
	jcb g273(.dina(n329),.dinb(n326),.dout(G432gat));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_8Q9aDmsZ4_0),.doutb(w_dff_A_S9cH5ASg8_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_dff_A_QeiAwPo49_0),.doutb(w_G4gat_0[1]),.doutc(w_dff_A_ackFX2VS9_2),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_KxQ4NtnU9_0),.doutb(w_dff_A_kYYK6bRS4_1),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G11gat_0(.douta(w_dff_A_Ds2KCWjB4_0),.doutb(w_dff_A_zx77paec5_1),.doutc(w_G11gat_0[2]),.din(G11gat));
	jspl3 jspl3_w_G14gat_0(.douta(w_dff_A_n6XHEdUj8_0),.doutb(w_dff_A_UQ0gZUMf1_1),.doutc(w_G14gat_0[2]),.din(G14gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_dff_A_tQeqhSFR8_0),.doutb(w_G17gat_0[1]),.doutc(w_dff_A_RuHE0NNv0_2),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_G21gat_0[0]),.doutb(w_dff_A_lB43AEcG3_1),.doutc(w_dff_A_Ys6RiXrh8_2),.din(G21gat));
	jspl jspl_w_G21gat_1(.douta(w_dff_A_qDqggfUI9_0),.doutb(w_G21gat_1[1]),.din(w_G21gat_0[0]));
	jspl jspl_w_G24gat_0(.douta(w_dff_A_tH6gJrwO5_0),.doutb(w_G24gat_0[1]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_dff_A_A3IUWPZP3_0),.doutb(w_G27gat_0[1]),.din(G27gat));
	jspl jspl_w_G30gat_0(.douta(w_G30gat_0[0]),.doutb(w_dff_A_4SCBLVVK6_1),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_dff_A_F8LbHkJN7_0),.doutb(w_G34gat_0[1]),.doutc(w_dff_A_ZMC09e0a7_2),.din(G34gat));
	jspl3 jspl3_w_G37gat_0(.douta(w_dff_A_pq1DDwcH6_0),.doutb(w_dff_A_Q2VAeA2m4_1),.doutc(w_G37gat_0[2]),.din(G37gat));
	jspl jspl_w_G40gat_0(.douta(w_dff_A_BdJINvIe4_0),.doutb(w_G40gat_0[1]),.din(G40gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_G43gat_0[0]),.doutb(w_dff_A_4XfPiDUQ5_1),.doutc(w_dff_A_KwYcxXwP8_2),.din(G43gat));
	jspl jspl_w_G43gat_1(.douta(w_G43gat_1[0]),.doutb(w_dff_A_bjbEQ63G7_1),.din(w_G43gat_0[0]));
	jspl jspl_w_G47gat_0(.douta(w_dff_A_QBSlD7Dg1_0),.doutb(w_G47gat_0[1]),.din(G47gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_dff_A_fFAyDfkg4_0),.doutb(w_dff_A_ccVj2SPm1_1),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_dff_A_Azx8s1LO1_0),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_dff_A_ykuSPxPC3_0),.doutb(w_G56gat_0[1]),.doutc(w_dff_A_yhPEyTC79_2),.din(G56gat));
	jspl3 jspl3_w_G60gat_0(.douta(w_dff_A_DqS6Uenx5_0),.doutb(w_dff_A_EYMhh2NP2_1),.doutc(w_G60gat_0[2]),.din(G60gat));
	jspl3 jspl3_w_G63gat_0(.douta(w_dff_A_hJhMiXj88_0),.doutb(w_dff_A_kRPglyTL6_1),.doutc(w_G63gat_0[2]),.din(G63gat));
	jspl jspl_w_G66gat_0(.douta(w_dff_A_98gxp4xM3_0),.doutb(w_G66gat_0[1]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_dff_A_cSh138lx0_0),.doutb(w_G69gat_0[1]),.doutc(w_dff_A_mNTfqqc63_2),.din(G69gat));
	jspl3 jspl3_w_G73gat_0(.douta(w_dff_A_B9xrlfVz5_0),.doutb(w_dff_A_R0XfIb7R3_1),.doutc(w_G73gat_0[2]),.din(G73gat));
	jspl jspl_w_G76gat_0(.douta(w_dff_A_V77Qgtx09_0),.doutb(w_G76gat_0[1]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_dff_A_6ukVAaVQ2_0),.doutb(w_G79gat_0[1]),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_G82gat_0[0]),.doutb(w_dff_A_68cmWWIi9_1),.doutc(w_dff_A_xeQ0w4hR0_2),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_dff_A_6CSFh7d00_1),.doutc(w_dff_A_KwcRjYcX8_2),.din(G86gat));
	jspl jspl_w_G86gat_1(.douta(w_dff_A_K5bHggug5_0),.doutb(w_G86gat_1[1]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G89gat_0(.douta(w_dff_A_mK9E1x6N7_0),.doutb(w_dff_A_spUQlFXn1_1),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_T3NsGRQx8_0),.doutb(w_dff_A_F9SGUW079_1),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_dff_A_UAZ4UGCm2_0),.doutb(w_G95gat_0[1]),.doutc(w_dff_A_dZ1WiuOi5_2),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_YjA6dPWN9_0),.doutb(w_dff_A_sIDebUwH7_1),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl3 jspl3_w_G102gat_0(.douta(w_dff_A_iwJkMMKv3_0),.doutb(w_dff_A_bZE7w3OJ6_1),.doutc(w_G102gat_0[2]),.din(G102gat));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_dff_A_ByEd35Mx2_1),.din(G105gat));
	jspl3 jspl3_w_G108gat_0(.douta(w_dff_A_EIPkYlR64_0),.doutb(w_G108gat_0[1]),.doutc(w_dff_A_x97kb6s77_2),.din(G108gat));
	jspl3 jspl3_w_G112gat_0(.douta(w_dff_A_oxSmCrPp1_0),.doutb(w_dff_A_r9UuOjSk8_1),.doutc(w_G112gat_0[2]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_dff_A_jovG9FKY9_0),.doutb(w_G115gat_0[1]),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(G223gat),.din(w_G223gat_0[2]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl3 jspl3_w_G329gat_4(.douta(w_G329gat_4[0]),.doutb(w_G329gat_4[1]),.doutc(w_G329gat_4[2]),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G329gat_5(.douta(w_G329gat_5[0]),.doutb(w_G329gat_5[1]),.doutc(w_G329gat_5[2]),.din(w_G329gat_1[1]));
	jspl jspl_w_G329gat_6(.douta(w_G329gat_6),.doutb(G329gat),.din(w_G329gat_1[2]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_G370gat_1[2]),.din(w_G370gat_0[0]));
	jspl jspl_w_G370gat_2(.douta(w_G370gat_2),.doutb(G370gat),.din(w_G370gat_0[1]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(G430gat),.din(G430gat_fa_));
	jspl jspl_w_n43_0(.douta(w_dff_A_PDTzFAbJ0_0),.doutb(w_n43_0[1]),.din(n43));
	jspl jspl_w_n44_0(.douta(w_n44_0[0]),.doutb(w_n44_0[1]),.din(n44));
	jspl jspl_w_n47_0(.douta(w_dff_A_9GXswcgi6_0),.doutb(w_n47_0[1]),.din(n47));
	jspl jspl_w_n52_0(.douta(w_dff_A_pv6JlPPU4_0),.doutb(w_n52_0[1]),.din(n52));
	jspl jspl_w_n53_0(.douta(w_dff_A_EuZn7Eiy6_0),.doutb(w_n53_0[1]),.din(n53));
	jspl jspl_w_n56_0(.douta(w_dff_A_yHbq8kSS5_0),.doutb(w_n56_0[1]),.din(n56));
	jspl jspl_w_n58_0(.douta(w_dff_A_Gos5lcXw0_0),.doutb(w_n58_0[1]),.din(n58));
	jspl jspl_w_n61_0(.douta(w_dff_A_Gis9XQrO3_0),.doutb(w_n61_0[1]),.din(n61));
	jspl jspl_w_n63_0(.douta(w_dff_A_cXNwIErP0_0),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n69_0(.douta(w_dff_A_0K2V6HLY3_0),.doutb(w_n69_0[1]),.din(w_dff_B_qb1tUmSa4_2));
	jspl jspl_w_n71_0(.douta(w_dff_A_AtdiSjA13_0),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n72_0(.douta(w_dff_A_Ta83EDWr3_0),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n73_0(.douta(w_dff_A_jNCouyL34_0),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n77_0(.douta(w_dff_A_LR7YmvsM5_0),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_dff_A_YTuRB6Gf8_0),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n79_0(.douta(w_dff_A_gaki3A8c6_0),.doutb(w_n79_0[1]),.din(n79));
	jspl jspl_w_n82_0(.douta(w_dff_A_4RWu16j10_0),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_dff_A_SAaoQR5h7_0),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n87_0(.douta(w_dff_A_ofGCrke68_0),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_dff_A_v4vcAIMn0_0),.doutb(w_n89_0[1]),.din(n89));
	jspl3 jspl3_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl3 jspl3_w_n94_1(.douta(w_n94_1[0]),.doutb(w_n94_1[1]),.doutc(w_n94_1[2]),.din(w_n94_0[0]));
	jspl3 jspl3_w_n94_2(.douta(w_n94_2[0]),.doutb(w_n94_2[1]),.doutc(w_n94_2[2]),.din(w_n94_0[1]));
	jspl3 jspl3_w_n94_3(.douta(w_n94_3[0]),.doutb(w_n94_3[1]),.doutc(w_n94_3[2]),.din(w_n94_0[2]));
	jspl jspl_w_n94_4(.douta(w_n94_4[0]),.doutb(w_n94_4[1]),.din(w_n94_1[0]));
	jspl jspl_w_n96_0(.douta(w_dff_A_zBbLDxvQ0_0),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_dff_A_PUtd6XR36_0),.doutb(w_n98_0[1]),.din(w_dff_B_tHKxWh0D8_2));
	jspl jspl_w_n100_0(.douta(w_dff_A_Ka4lySTd9_0),.doutb(w_n100_0[1]),.din(n100));
	jspl jspl_w_n107_0(.douta(w_dff_A_CDO7FLDy4_0),.doutb(w_n107_0[1]),.din(w_dff_B_Vyv08kLF5_2));
	jspl jspl_w_n109_0(.douta(w_dff_A_Zypb9wwg6_0),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n114_0(.douta(w_dff_A_K5gZdYiz0_0),.doutb(w_n114_0[1]),.doutc(w_n114_0[2]),.din(n114));
	jspl jspl_w_n115_0(.douta(w_dff_A_UYDvcHSI1_0),.doutb(w_n115_0[1]),.din(n115));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n123_0(.douta(w_n123_0[0]),.doutb(w_dff_A_w7DTeoif4_1),.din(n123));
	jspl3 jspl3_w_n126_0(.douta(w_dff_A_AuCjO2Rd0_0),.doutb(w_dff_A_Q5I9TeQr4_1),.doutc(w_n126_0[2]),.din(w_dff_B_2BcIh0H47_3));
	jspl jspl_w_n128_0(.douta(w_dff_A_GS2qVlTL6_0),.doutb(w_n128_0[1]),.din(n128));
	jspl3 jspl3_w_n130_0(.douta(w_dff_A_OqN5NvHD9_0),.doutb(w_dff_A_PIFyp6Mc1_1),.doutc(w_n130_0[2]),.din(w_dff_B_2zO58puS2_3));
	jspl jspl_w_n132_0(.douta(w_dff_A_qZrV8PM09_0),.doutb(w_n132_0[1]),.din(n132));
	jspl jspl_w_n139_0(.douta(w_n139_0[0]),.doutb(w_dff_A_LnOkSJ5j2_1),.din(n139));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_dff_A_DBLhnoT00_0),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n145_0(.douta(w_dff_A_rkrCP9Nh7_0),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_ThHCmN9U9_1),.din(w_dff_B_AvNIJiip3_2));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl jspl_w_n150_0(.douta(w_dff_A_gmRkcWga9_0),.doutb(w_n150_0[1]),.din(w_dff_B_2xp4turu3_2));
	jspl jspl_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_ErzZilkO7_1),.din(n151));
	jspl jspl_w_n154_0(.douta(w_dff_A_ygsYRx3b7_0),.doutb(w_n154_0[1]),.din(w_dff_B_vPY4wFJg5_2));
	jspl jspl_w_n156_0(.douta(w_dff_A_sO1JVLwy0_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n159_0(.douta(w_dff_A_pqUeLYjz8_0),.doutb(w_n159_0[1]),.din(n159));
	jspl jspl_w_n164_0(.douta(w_dff_A_Im4Zx6Q98_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n170_0(.douta(w_dff_A_45LdLgW39_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n174_0(.douta(w_dff_A_amCOZp3N3_0),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n177_0(.douta(w_dff_A_PK1iZVts9_0),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n182_2(.douta(w_n182_2[0]),.doutb(w_n182_2[1]),.doutc(w_n182_2[2]),.din(w_n182_0[1]));
	jspl jspl_w_n182_3(.douta(w_n182_3[0]),.doutb(w_n182_3[1]),.din(w_n182_0[2]));
	jspl jspl_w_n184_0(.douta(w_dff_A_yjadT7ge8_0),.doutb(w_n184_0[1]),.din(n184));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n191_0(.douta(w_dff_A_4hKiCFt56_0),.doutb(w_n191_0[1]),.din(n191));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_dff_A_aZStHclE5_1),.din(n193));
	jspl jspl_w_n197_0(.douta(w_dff_A_BNcYI1jW3_0),.doutb(w_n197_0[1]),.din(n197));
	jspl jspl_w_n198_0(.douta(w_dff_A_lvyuG3S28_0),.doutb(w_n198_0[1]),.din(w_dff_B_gn2lZ5EV5_2));
	jspl jspl_w_n204_0(.douta(w_dff_A_ZXqWWYqh1_0),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n205_0(.douta(w_dff_A_1sgwg0GZ7_0),.doutb(w_n205_0[1]),.din(w_dff_B_T1KCYwbu9_2));
	jspl jspl_w_n217_0(.douta(w_dff_A_fH58VTXp6_0),.doutb(w_n217_0[1]),.din(w_dff_B_p270DQTj0_2));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_dff_A_Kz7b49HT1_1),.din(n219));
	jspl jspl_w_n222_0(.douta(w_dff_A_jUKicEId0_0),.doutb(w_n222_0[1]),.din(w_dff_B_dAgSW9SZ3_2));
	jspl jspl_w_n224_0(.douta(w_dff_A_wO3lTOII3_0),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_dff_A_tPfc51Xj1_1),.din(n231));
	jspl jspl_w_n254_0(.douta(w_dff_A_YDJ1gxww5_0),.doutb(w_n254_0[1]),.din(w_dff_B_cw23lUTm5_2));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_dff_A_hueS9QO64_1),.din(n260));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_n271_1[0]),.doutb(w_n271_1[1]),.doutc(w_n271_1[2]),.din(w_n271_0[0]));
	jspl3 jspl3_w_n271_2(.douta(w_n271_2[0]),.doutb(w_n271_2[1]),.doutc(w_n271_2[2]),.din(w_n271_0[1]));
	jspl jspl_w_n271_3(.douta(w_n271_3[0]),.doutb(w_n271_3[1]),.din(w_n271_0[2]));
	jspl jspl_w_n274_0(.douta(w_dff_A_jLUDdNHJ6_0),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n281_0(.douta(w_dff_A_nCOlxojz0_0),.doutb(w_n281_0[1]),.din(n281));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.din(n283));
	jspl jspl_w_n286_0(.douta(w_dff_A_l8TA9xag9_0),.doutb(w_n286_0[1]),.din(n286));
	jspl jspl_w_n290_0(.douta(w_dff_A_twwzGNpN2_0),.doutb(w_n290_0[1]),.din(n290));
	jspl jspl_w_n293_0(.douta(w_dff_A_57a6Uuz23_0),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(n305));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl jspl_w_n314_0(.douta(w_dff_A_lC6q45058_0),.doutb(w_n314_0[1]),.din(w_dff_B_pDlUUxKz7_2));
	jspl3 jspl3_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.doutc(w_n317_0[2]),.din(w_dff_B_hXQrdu6m1_3));
	jspl jspl_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.din(n319));
	jdff dff_B_NNAzo5ez5_1(.din(n233),.dout(w_dff_B_NNAzo5ez5_1),.clk(gclk));
	jdff dff_B_LjWFwRck8_1(.din(w_dff_B_NNAzo5ez5_1),.dout(w_dff_B_LjWFwRck8_1),.clk(gclk));
	jdff dff_B_KumAQcfB7_1(.din(w_dff_B_LjWFwRck8_1),.dout(w_dff_B_KumAQcfB7_1),.clk(gclk));
	jdff dff_B_re7nzJSS3_0(.din(n275),.dout(w_dff_B_re7nzJSS3_0),.clk(gclk));
	jdff dff_B_7RirBMnF4_0(.din(w_dff_B_re7nzJSS3_0),.dout(w_dff_B_7RirBMnF4_0),.clk(gclk));
	jdff dff_B_DlRgxCvk4_0(.din(w_dff_B_7RirBMnF4_0),.dout(w_dff_B_DlRgxCvk4_0),.clk(gclk));
	jdff dff_B_cqLXRr0u4_0(.din(w_dff_B_DlRgxCvk4_0),.dout(w_dff_B_cqLXRr0u4_0),.clk(gclk));
	jdff dff_B_eX5WKZFn6_0(.din(w_dff_B_cqLXRr0u4_0),.dout(w_dff_B_eX5WKZFn6_0),.clk(gclk));
	jdff dff_B_XTwMCCN78_0(.din(w_dff_B_eX5WKZFn6_0),.dout(w_dff_B_XTwMCCN78_0),.clk(gclk));
	jdff dff_B_DT7GTFZ78_1(.din(n315),.dout(w_dff_B_DT7GTFZ78_1),.clk(gclk));
	jdff dff_A_VbrR3Svo9_0(.dout(w_n293_0[0]),.din(w_dff_A_VbrR3Svo9_0),.clk(gclk));
	jdff dff_A_57a6Uuz23_0(.dout(w_dff_A_VbrR3Svo9_0),.din(w_dff_A_57a6Uuz23_0),.clk(gclk));
	jdff dff_B_4CsutdP87_0(.din(n291),.dout(w_dff_B_4CsutdP87_0),.clk(gclk));
	jdff dff_B_rSWyHv3o3_0(.din(w_dff_B_4CsutdP87_0),.dout(w_dff_B_rSWyHv3o3_0),.clk(gclk));
	jdff dff_B_QTBEKGTI2_0(.din(w_dff_B_rSWyHv3o3_0),.dout(w_dff_B_QTBEKGTI2_0),.clk(gclk));
	jdff dff_B_BRRmZ4vR4_0(.din(w_dff_B_QTBEKGTI2_0),.dout(w_dff_B_BRRmZ4vR4_0),.clk(gclk));
	jdff dff_B_kRRpcpBl2_0(.din(w_dff_B_BRRmZ4vR4_0),.dout(w_dff_B_kRRpcpBl2_0),.clk(gclk));
	jdff dff_B_H7dSlUJY2_0(.din(w_dff_B_kRRpcpBl2_0),.dout(w_dff_B_H7dSlUJY2_0),.clk(gclk));
	jdff dff_B_wi0W0TXf6_0(.din(n328),.dout(w_dff_B_wi0W0TXf6_0),.clk(gclk));
	jdff dff_B_5VZfKCJ99_0(.din(n282),.dout(w_dff_B_5VZfKCJ99_0),.clk(gclk));
	jdff dff_B_aBdLMG4F6_0(.din(w_dff_B_5VZfKCJ99_0),.dout(w_dff_B_aBdLMG4F6_0),.clk(gclk));
	jdff dff_B_gyyUuk2t2_0(.din(w_dff_B_aBdLMG4F6_0),.dout(w_dff_B_gyyUuk2t2_0),.clk(gclk));
	jdff dff_B_1NKPMYqv0_0(.din(w_dff_B_gyyUuk2t2_0),.dout(w_dff_B_1NKPMYqv0_0),.clk(gclk));
	jdff dff_B_ykPddIkY9_0(.din(w_dff_B_1NKPMYqv0_0),.dout(w_dff_B_ykPddIkY9_0),.clk(gclk));
	jdff dff_B_huyq7yRr4_0(.din(w_dff_B_ykPddIkY9_0),.dout(w_dff_B_huyq7yRr4_0),.clk(gclk));
	jdff dff_A_l8TA9xag9_0(.dout(w_n286_0[0]),.din(w_dff_A_l8TA9xag9_0),.clk(gclk));
	jdff dff_A_lC6q45058_0(.dout(w_n314_0[0]),.din(w_dff_A_lC6q45058_0),.clk(gclk));
	jdff dff_B_qacHT2eE3_2(.din(n314),.dout(w_dff_B_qacHT2eE3_2),.clk(gclk));
	jdff dff_B_pDlUUxKz7_2(.din(w_dff_B_qacHT2eE3_2),.dout(w_dff_B_pDlUUxKz7_2),.clk(gclk));
	jdff dff_A_QzSmpVMj2_0(.dout(w_n274_0[0]),.din(w_dff_A_QzSmpVMj2_0),.clk(gclk));
	jdff dff_A_ajmtU2Kc5_0(.dout(w_dff_A_QzSmpVMj2_0),.din(w_dff_A_ajmtU2Kc5_0),.clk(gclk));
	jdff dff_A_AUtTnTtB4_0(.dout(w_dff_A_ajmtU2Kc5_0),.din(w_dff_A_AUtTnTtB4_0),.clk(gclk));
	jdff dff_A_YxinQqic0_0(.dout(w_dff_A_AUtTnTtB4_0),.din(w_dff_A_YxinQqic0_0),.clk(gclk));
	jdff dff_A_jLUDdNHJ6_0(.dout(w_dff_A_YxinQqic0_0),.din(w_dff_A_jLUDdNHJ6_0),.clk(gclk));
	jdff dff_B_kx9oFqVr3_0(.din(n325),.dout(w_dff_B_kx9oFqVr3_0),.clk(gclk));
	jdff dff_B_sTlSopjC5_0(.din(w_dff_B_kx9oFqVr3_0),.dout(w_dff_B_sTlSopjC5_0),.clk(gclk));
	jdff dff_B_0jpW6hqj9_0(.din(w_dff_B_sTlSopjC5_0),.dout(w_dff_B_0jpW6hqj9_0),.clk(gclk));
	jdff dff_A_y4kzilGs0_0(.dout(w_n281_0[0]),.din(w_dff_A_y4kzilGs0_0),.clk(gclk));
	jdff dff_A_2gWDS8Pv5_0(.dout(w_dff_A_y4kzilGs0_0),.din(w_dff_A_2gWDS8Pv5_0),.clk(gclk));
	jdff dff_A_CESwO5LL4_0(.dout(w_dff_A_2gWDS8Pv5_0),.din(w_dff_A_CESwO5LL4_0),.clk(gclk));
	jdff dff_A_aghYQyFm5_0(.dout(w_dff_A_CESwO5LL4_0),.din(w_dff_A_aghYQyFm5_0),.clk(gclk));
	jdff dff_A_nCOlxojz0_0(.dout(w_dff_A_aghYQyFm5_0),.din(w_dff_A_nCOlxojz0_0),.clk(gclk));
	jdff dff_B_MKx9TkqZ7_0(.din(n280),.dout(w_dff_B_MKx9TkqZ7_0),.clk(gclk));
	jdff dff_B_1WgPJZoq7_0(.din(w_dff_B_MKx9TkqZ7_0),.dout(w_dff_B_1WgPJZoq7_0),.clk(gclk));
	jdff dff_B_hlTOnxwO7_0(.din(w_dff_B_1WgPJZoq7_0),.dout(w_dff_B_hlTOnxwO7_0),.clk(gclk));
	jdff dff_B_STSxD65J2_0(.din(w_dff_B_hlTOnxwO7_0),.dout(w_dff_B_STSxD65J2_0),.clk(gclk));
	jdff dff_B_WZY9NVfD0_0(.din(w_dff_B_STSxD65J2_0),.dout(w_dff_B_WZY9NVfD0_0),.clk(gclk));
	jdff dff_B_pMmHWCzx8_1(.din(n300),.dout(w_dff_B_pMmHWCzx8_1),.clk(gclk));
	jdff dff_B_SuetQrwe0_1(.din(w_dff_B_pMmHWCzx8_1),.dout(w_dff_B_SuetQrwe0_1),.clk(gclk));
	jdff dff_B_kJU5ADqp7_1(.din(w_dff_B_SuetQrwe0_1),.dout(w_dff_B_kJU5ADqp7_1),.clk(gclk));
	jdff dff_B_PbAjnpRW2_1(.din(w_dff_B_kJU5ADqp7_1),.dout(w_dff_B_PbAjnpRW2_1),.clk(gclk));
	jdff dff_B_tYvIWOvL3_1(.din(w_dff_B_PbAjnpRW2_1),.dout(w_dff_B_tYvIWOvL3_1),.clk(gclk));
	jdff dff_B_pOpfgyo86_1(.din(w_dff_B_tYvIWOvL3_1),.dout(w_dff_B_pOpfgyo86_1),.clk(gclk));
	jdff dff_B_WXG14XJK5_1(.din(n301),.dout(w_dff_B_WXG14XJK5_1),.clk(gclk));
	jdff dff_B_6COZDPs56_1(.din(w_dff_B_WXG14XJK5_1),.dout(w_dff_B_6COZDPs56_1),.clk(gclk));
	jdff dff_B_iLSo7CQV5_1(.din(w_dff_B_6COZDPs56_1),.dout(w_dff_B_iLSo7CQV5_1),.clk(gclk));
	jdff dff_B_5aytIf7K8_1(.din(w_dff_B_iLSo7CQV5_1),.dout(w_dff_B_5aytIf7K8_1),.clk(gclk));
	jdff dff_B_LGlF82Bj9_1(.din(w_dff_B_5aytIf7K8_1),.dout(w_dff_B_LGlF82Bj9_1),.clk(gclk));
	jdff dff_B_WxnLOgQu4_1(.din(w_dff_B_LGlF82Bj9_1),.dout(w_dff_B_WxnLOgQu4_1),.clk(gclk));
	jdff dff_B_CbHy5VSx4_1(.din(w_dff_B_WxnLOgQu4_1),.dout(w_dff_B_CbHy5VSx4_1),.clk(gclk));
	jdff dff_B_AsHoFPKM0_1(.din(w_dff_B_CbHy5VSx4_1),.dout(w_dff_B_AsHoFPKM0_1),.clk(gclk));
	jdff dff_B_usN9BBhI1_1(.din(w_dff_B_AsHoFPKM0_1),.dout(w_dff_B_usN9BBhI1_1),.clk(gclk));
	jdff dff_B_XdWY8pKv6_1(.din(w_dff_B_usN9BBhI1_1),.dout(w_dff_B_XdWY8pKv6_1),.clk(gclk));
	jdff dff_B_fFN1zz8A3_1(.din(w_dff_B_XdWY8pKv6_1),.dout(w_dff_B_fFN1zz8A3_1),.clk(gclk));
	jdff dff_B_QzanNSGG8_1(.din(w_dff_B_fFN1zz8A3_1),.dout(w_dff_B_QzanNSGG8_1),.clk(gclk));
	jdff dff_B_MCw2aYup6_1(.din(w_dff_B_QzanNSGG8_1),.dout(w_dff_B_MCw2aYup6_1),.clk(gclk));
	jdff dff_B_G9r9K1T88_1(.din(w_dff_B_MCw2aYup6_1),.dout(w_dff_B_G9r9K1T88_1),.clk(gclk));
	jdff dff_B_nDzhsVir4_1(.din(n242),.dout(w_dff_B_nDzhsVir4_1),.clk(gclk));
	jdff dff_B_9LZIO7vR5_1(.din(w_dff_B_nDzhsVir4_1),.dout(w_dff_B_9LZIO7vR5_1),.clk(gclk));
	jdff dff_B_zI66Mbb68_1(.din(w_dff_B_9LZIO7vR5_1),.dout(w_dff_B_zI66Mbb68_1),.clk(gclk));
	jdff dff_B_BlhSNEHh9_1(.din(w_dff_B_zI66Mbb68_1),.dout(w_dff_B_BlhSNEHh9_1),.clk(gclk));
	jdff dff_B_nKBhQB1W6_1(.din(n252),.dout(w_dff_B_nKBhQB1W6_1),.clk(gclk));
	jdff dff_B_mtQiiog55_0(.din(n268),.dout(w_dff_B_mtQiiog55_0),.clk(gclk));
	jdff dff_B_q1ZvadfE8_0(.din(w_dff_B_mtQiiog55_0),.dout(w_dff_B_q1ZvadfE8_0),.clk(gclk));
	jdff dff_B_RuLZw8Ua2_0(.din(n267),.dout(w_dff_B_RuLZw8Ua2_0),.clk(gclk));
	jdff dff_B_VDGaAm5s7_0(.din(n258),.dout(w_dff_B_VDGaAm5s7_0),.clk(gclk));
	jdff dff_B_FzdHCtZe2_0(.din(w_dff_B_VDGaAm5s7_0),.dout(w_dff_B_FzdHCtZe2_0),.clk(gclk));
	jdff dff_B_dBUvcGT71_0(.din(w_dff_B_FzdHCtZe2_0),.dout(w_dff_B_dBUvcGT71_0),.clk(gclk));
	jdff dff_A_IbpRZwoY1_1(.dout(w_n231_0[1]),.din(w_dff_A_IbpRZwoY1_1),.clk(gclk));
	jdff dff_A_6SQvWR6o7_1(.dout(w_dff_A_IbpRZwoY1_1),.din(w_dff_A_6SQvWR6o7_1),.clk(gclk));
	jdff dff_A_nSldGmhS8_1(.dout(w_dff_A_6SQvWR6o7_1),.din(w_dff_A_nSldGmhS8_1),.clk(gclk));
	jdff dff_A_ER1SrXHP2_1(.dout(w_dff_A_nSldGmhS8_1),.din(w_dff_A_ER1SrXHP2_1),.clk(gclk));
	jdff dff_A_tPfc51Xj1_1(.dout(w_dff_A_ER1SrXHP2_1),.din(w_dff_A_tPfc51Xj1_1),.clk(gclk));
	jdff dff_A_5PS2gS7j8_0(.dout(w_n254_0[0]),.din(w_dff_A_5PS2gS7j8_0),.clk(gclk));
	jdff dff_A_YDJ1gxww5_0(.dout(w_dff_A_5PS2gS7j8_0),.din(w_dff_A_YDJ1gxww5_0),.clk(gclk));
	jdff dff_B_qCFSnN2y9_2(.din(n254),.dout(w_dff_B_qCFSnN2y9_2),.clk(gclk));
	jdff dff_B_vHMFABkU9_2(.din(w_dff_B_qCFSnN2y9_2),.dout(w_dff_B_vHMFABkU9_2),.clk(gclk));
	jdff dff_B_cw23lUTm5_2(.din(w_dff_B_vHMFABkU9_2),.dout(w_dff_B_cw23lUTm5_2),.clk(gclk));
	jdff dff_B_k1nrhP409_1(.din(n246),.dout(w_dff_B_k1nrhP409_1),.clk(gclk));
	jdff dff_B_kBUEQRTF0_1(.din(w_dff_B_k1nrhP409_1),.dout(w_dff_B_kBUEQRTF0_1),.clk(gclk));
	jdff dff_B_63L91ISR7_1(.din(w_dff_B_kBUEQRTF0_1),.dout(w_dff_B_63L91ISR7_1),.clk(gclk));
	jdff dff_B_ADThpRlJ6_1(.din(n248),.dout(w_dff_B_ADThpRlJ6_1),.clk(gclk));
	jdff dff_B_UEHS9Rue4_1(.din(w_dff_B_ADThpRlJ6_1),.dout(w_dff_B_UEHS9Rue4_1),.clk(gclk));
	jdff dff_B_cx9NWvkF0_1(.din(w_dff_B_UEHS9Rue4_1),.dout(w_dff_B_cx9NWvkF0_1),.clk(gclk));
	jdff dff_B_0ez9y9bH3_3(.din(n317),.dout(w_dff_B_0ez9y9bH3_3),.clk(gclk));
	jdff dff_B_BhTVwoiE5_3(.din(w_dff_B_0ez9y9bH3_3),.dout(w_dff_B_BhTVwoiE5_3),.clk(gclk));
	jdff dff_B_hXQrdu6m1_3(.din(w_dff_B_BhTVwoiE5_3),.dout(w_dff_B_hXQrdu6m1_3),.clk(gclk));
	jdff dff_A_fJ3BgBZi1_0(.dout(w_n290_0[0]),.din(w_dff_A_fJ3BgBZi1_0),.clk(gclk));
	jdff dff_A_bwjzrf8s6_0(.dout(w_dff_A_fJ3BgBZi1_0),.din(w_dff_A_bwjzrf8s6_0),.clk(gclk));
	jdff dff_A_E2ysPMuG0_0(.dout(w_dff_A_bwjzrf8s6_0),.din(w_dff_A_E2ysPMuG0_0),.clk(gclk));
	jdff dff_A_rtfRFXE34_0(.dout(w_dff_A_E2ysPMuG0_0),.din(w_dff_A_rtfRFXE34_0),.clk(gclk));
	jdff dff_A_twwzGNpN2_0(.dout(w_dff_A_rtfRFXE34_0),.din(w_dff_A_twwzGNpN2_0),.clk(gclk));
	jdff dff_A_hueS9QO64_1(.dout(w_n260_0[1]),.din(w_dff_A_hueS9QO64_1),.clk(gclk));
	jdff dff_B_NfZgjlwf5_1(.din(n221),.dout(w_dff_B_NfZgjlwf5_1),.clk(gclk));
	jdff dff_A_NT74VLku4_0(.dout(w_n224_0[0]),.din(w_dff_A_NT74VLku4_0),.clk(gclk));
	jdff dff_A_cE2g9gf94_0(.dout(w_dff_A_NT74VLku4_0),.din(w_dff_A_cE2g9gf94_0),.clk(gclk));
	jdff dff_A_W0FYNaVC8_0(.dout(w_dff_A_cE2g9gf94_0),.din(w_dff_A_W0FYNaVC8_0),.clk(gclk));
	jdff dff_A_wO3lTOII3_0(.dout(w_dff_A_W0FYNaVC8_0),.din(w_dff_A_wO3lTOII3_0),.clk(gclk));
	jdff dff_A_PRB0O4F03_0(.dout(w_n222_0[0]),.din(w_dff_A_PRB0O4F03_0),.clk(gclk));
	jdff dff_A_NFUlC0aO7_0(.dout(w_dff_A_PRB0O4F03_0),.din(w_dff_A_NFUlC0aO7_0),.clk(gclk));
	jdff dff_A_RLmbjydG7_0(.dout(w_dff_A_NFUlC0aO7_0),.din(w_dff_A_RLmbjydG7_0),.clk(gclk));
	jdff dff_A_jUKicEId0_0(.dout(w_dff_A_RLmbjydG7_0),.din(w_dff_A_jUKicEId0_0),.clk(gclk));
	jdff dff_B_QPu4F5w71_2(.din(n222),.dout(w_dff_B_QPu4F5w71_2),.clk(gclk));
	jdff dff_B_74pYg0I73_2(.din(w_dff_B_QPu4F5w71_2),.dout(w_dff_B_74pYg0I73_2),.clk(gclk));
	jdff dff_B_kMHmiD887_2(.din(w_dff_B_74pYg0I73_2),.dout(w_dff_B_kMHmiD887_2),.clk(gclk));
	jdff dff_B_4d9Ks3Kf6_2(.din(w_dff_B_kMHmiD887_2),.dout(w_dff_B_4d9Ks3Kf6_2),.clk(gclk));
	jdff dff_B_2QA2Dpgb7_2(.din(w_dff_B_4d9Ks3Kf6_2),.dout(w_dff_B_2QA2Dpgb7_2),.clk(gclk));
	jdff dff_B_m7tctwbd5_2(.din(w_dff_B_2QA2Dpgb7_2),.dout(w_dff_B_m7tctwbd5_2),.clk(gclk));
	jdff dff_B_13boSzhX0_2(.din(w_dff_B_m7tctwbd5_2),.dout(w_dff_B_13boSzhX0_2),.clk(gclk));
	jdff dff_B_LhaKIiE29_2(.din(w_dff_B_13boSzhX0_2),.dout(w_dff_B_LhaKIiE29_2),.clk(gclk));
	jdff dff_B_4wcdZRlD8_2(.din(w_dff_B_LhaKIiE29_2),.dout(w_dff_B_4wcdZRlD8_2),.clk(gclk));
	jdff dff_B_dAgSW9SZ3_2(.din(w_dff_B_4wcdZRlD8_2),.dout(w_dff_B_dAgSW9SZ3_2),.clk(gclk));
	jdff dff_A_IYR4xoeH0_0(.dout(w_G115gat_0[0]),.din(w_dff_A_IYR4xoeH0_0),.clk(gclk));
	jdff dff_A_xZN92ch06_0(.dout(w_dff_A_IYR4xoeH0_0),.din(w_dff_A_xZN92ch06_0),.clk(gclk));
	jdff dff_A_E8iWS6TP6_0(.dout(w_dff_A_xZN92ch06_0),.din(w_dff_A_E8iWS6TP6_0),.clk(gclk));
	jdff dff_A_c3fldacj6_0(.dout(w_dff_A_E8iWS6TP6_0),.din(w_dff_A_c3fldacj6_0),.clk(gclk));
	jdff dff_A_p5dQdp7B1_0(.dout(w_dff_A_c3fldacj6_0),.din(w_dff_A_p5dQdp7B1_0),.clk(gclk));
	jdff dff_A_bDMsQRBX9_0(.dout(w_dff_A_p5dQdp7B1_0),.din(w_dff_A_bDMsQRBX9_0),.clk(gclk));
	jdff dff_A_4EA5zdRI4_0(.dout(w_dff_A_bDMsQRBX9_0),.din(w_dff_A_4EA5zdRI4_0),.clk(gclk));
	jdff dff_A_jovG9FKY9_0(.dout(w_dff_A_4EA5zdRI4_0),.din(w_dff_A_jovG9FKY9_0),.clk(gclk));
	jdff dff_A_UBfoKA1H8_1(.dout(w_n219_0[1]),.din(w_dff_A_UBfoKA1H8_1),.clk(gclk));
	jdff dff_A_Kz7b49HT1_1(.dout(w_dff_A_UBfoKA1H8_1),.din(w_dff_A_Kz7b49HT1_1),.clk(gclk));
	jdff dff_A_TRga1sTf0_0(.dout(w_n217_0[0]),.din(w_dff_A_TRga1sTf0_0),.clk(gclk));
	jdff dff_A_5jgl3oVI5_0(.dout(w_dff_A_TRga1sTf0_0),.din(w_dff_A_5jgl3oVI5_0),.clk(gclk));
	jdff dff_A_ydR0BTVG5_0(.dout(w_dff_A_5jgl3oVI5_0),.din(w_dff_A_ydR0BTVG5_0),.clk(gclk));
	jdff dff_A_ZYiiNVLQ6_0(.dout(w_dff_A_ydR0BTVG5_0),.din(w_dff_A_ZYiiNVLQ6_0),.clk(gclk));
	jdff dff_A_x99nVF944_0(.dout(w_dff_A_ZYiiNVLQ6_0),.din(w_dff_A_x99nVF944_0),.clk(gclk));
	jdff dff_A_kpfsJ6rd1_0(.dout(w_dff_A_x99nVF944_0),.din(w_dff_A_kpfsJ6rd1_0),.clk(gclk));
	jdff dff_A_uG6fHCXf6_0(.dout(w_dff_A_kpfsJ6rd1_0),.din(w_dff_A_uG6fHCXf6_0),.clk(gclk));
	jdff dff_A_fH58VTXp6_0(.dout(w_dff_A_uG6fHCXf6_0),.din(w_dff_A_fH58VTXp6_0),.clk(gclk));
	jdff dff_B_klVZumzE8_2(.din(n217),.dout(w_dff_B_klVZumzE8_2),.clk(gclk));
	jdff dff_B_uUPXFwHZ8_2(.din(w_dff_B_klVZumzE8_2),.dout(w_dff_B_uUPXFwHZ8_2),.clk(gclk));
	jdff dff_B_qNaHHyIp1_2(.din(w_dff_B_uUPXFwHZ8_2),.dout(w_dff_B_qNaHHyIp1_2),.clk(gclk));
	jdff dff_B_ZdyRjlON2_2(.din(w_dff_B_qNaHHyIp1_2),.dout(w_dff_B_ZdyRjlON2_2),.clk(gclk));
	jdff dff_B_xww0tWIQ3_2(.din(w_dff_B_ZdyRjlON2_2),.dout(w_dff_B_xww0tWIQ3_2),.clk(gclk));
	jdff dff_B_p270DQTj0_2(.din(w_dff_B_xww0tWIQ3_2),.dout(w_dff_B_p270DQTj0_2),.clk(gclk));
	jdff dff_A_xj2sYUjV9_0(.dout(w_G40gat_0[0]),.din(w_dff_A_xj2sYUjV9_0),.clk(gclk));
	jdff dff_A_R0QeNTxd5_0(.dout(w_dff_A_xj2sYUjV9_0),.din(w_dff_A_R0QeNTxd5_0),.clk(gclk));
	jdff dff_A_DgzJYiL52_0(.dout(w_dff_A_R0QeNTxd5_0),.din(w_dff_A_DgzJYiL52_0),.clk(gclk));
	jdff dff_A_ydn6721I3_0(.dout(w_dff_A_DgzJYiL52_0),.din(w_dff_A_ydn6721I3_0),.clk(gclk));
	jdff dff_A_gl96Tb8m4_0(.dout(w_dff_A_ydn6721I3_0),.din(w_dff_A_gl96Tb8m4_0),.clk(gclk));
	jdff dff_A_SxYdW0EY2_0(.dout(w_dff_A_gl96Tb8m4_0),.din(w_dff_A_SxYdW0EY2_0),.clk(gclk));
	jdff dff_A_iz3CEMhh3_0(.dout(w_dff_A_SxYdW0EY2_0),.din(w_dff_A_iz3CEMhh3_0),.clk(gclk));
	jdff dff_A_sOYWmSRN7_0(.dout(w_dff_A_iz3CEMhh3_0),.din(w_dff_A_sOYWmSRN7_0),.clk(gclk));
	jdff dff_A_OdLRWxCG1_0(.dout(w_dff_A_sOYWmSRN7_0),.din(w_dff_A_OdLRWxCG1_0),.clk(gclk));
	jdff dff_A_lQ80jKB65_0(.dout(w_dff_A_OdLRWxCG1_0),.din(w_dff_A_lQ80jKB65_0),.clk(gclk));
	jdff dff_A_Jn7ijbyN7_0(.dout(w_dff_A_lQ80jKB65_0),.din(w_dff_A_Jn7ijbyN7_0),.clk(gclk));
	jdff dff_A_BdJINvIe4_0(.dout(w_dff_A_Jn7ijbyN7_0),.din(w_dff_A_BdJINvIe4_0),.clk(gclk));
	jdff dff_B_aUb5jDP07_1(.din(n214),.dout(w_dff_B_aUb5jDP07_1),.clk(gclk));
	jdff dff_B_7h3X1Cgb7_1(.din(w_dff_B_aUb5jDP07_1),.dout(w_dff_B_7h3X1Cgb7_1),.clk(gclk));
	jdff dff_B_lutzR7G29_1(.din(w_dff_B_7h3X1Cgb7_1),.dout(w_dff_B_lutzR7G29_1),.clk(gclk));
	jdff dff_B_IttGQTE16_1(.din(w_dff_B_lutzR7G29_1),.dout(w_dff_B_IttGQTE16_1),.clk(gclk));
	jdff dff_B_lq9qRrrh7_1(.din(w_dff_B_IttGQTE16_1),.dout(w_dff_B_lq9qRrrh7_1),.clk(gclk));
	jdff dff_B_r4DKtmoG9_1(.din(w_dff_B_lq9qRrrh7_1),.dout(w_dff_B_r4DKtmoG9_1),.clk(gclk));
	jdff dff_B_mgImKyoN3_1(.din(w_dff_B_r4DKtmoG9_1),.dout(w_dff_B_mgImKyoN3_1),.clk(gclk));
	jdff dff_B_dg3ww7RA6_1(.din(w_dff_B_mgImKyoN3_1),.dout(w_dff_B_dg3ww7RA6_1),.clk(gclk));
	jdff dff_B_VCU9QS1w1_1(.din(w_dff_B_dg3ww7RA6_1),.dout(w_dff_B_VCU9QS1w1_1),.clk(gclk));
	jdff dff_B_RTlDi3Jd6_1(.din(n209),.dout(w_dff_B_RTlDi3Jd6_1),.clk(gclk));
	jdff dff_B_wOlzNPsq8_1(.din(w_dff_B_RTlDi3Jd6_1),.dout(w_dff_B_wOlzNPsq8_1),.clk(gclk));
	jdff dff_B_wjvURLz65_1(.din(w_dff_B_wOlzNPsq8_1),.dout(w_dff_B_wjvURLz65_1),.clk(gclk));
	jdff dff_B_p18gYLXB7_1(.din(w_dff_B_wjvURLz65_1),.dout(w_dff_B_p18gYLXB7_1),.clk(gclk));
	jdff dff_B_hhYWuN8p8_1(.din(w_dff_B_p18gYLXB7_1),.dout(w_dff_B_hhYWuN8p8_1),.clk(gclk));
	jdff dff_B_jRmp4DZU2_1(.din(w_dff_B_hhYWuN8p8_1),.dout(w_dff_B_jRmp4DZU2_1),.clk(gclk));
	jdff dff_B_WB9UUlEd5_1(.din(w_dff_B_jRmp4DZU2_1),.dout(w_dff_B_WB9UUlEd5_1),.clk(gclk));
	jdff dff_B_oq4HkBVB6_1(.din(w_dff_B_WB9UUlEd5_1),.dout(w_dff_B_oq4HkBVB6_1),.clk(gclk));
	jdff dff_B_nzZemYMx0_1(.din(w_dff_B_oq4HkBVB6_1),.dout(w_dff_B_nzZemYMx0_1),.clk(gclk));
	jdff dff_B_SLm6IIqn0_1(.din(w_dff_B_nzZemYMx0_1),.dout(w_dff_B_SLm6IIqn0_1),.clk(gclk));
	jdff dff_A_s7LV3qY29_0(.dout(w_G14gat_0[0]),.din(w_dff_A_s7LV3qY29_0),.clk(gclk));
	jdff dff_A_zLyxdrxy5_0(.dout(w_dff_A_s7LV3qY29_0),.din(w_dff_A_zLyxdrxy5_0),.clk(gclk));
	jdff dff_A_qiqysHQD8_0(.dout(w_dff_A_zLyxdrxy5_0),.din(w_dff_A_qiqysHQD8_0),.clk(gclk));
	jdff dff_A_amCkDlQG0_0(.dout(w_dff_A_qiqysHQD8_0),.din(w_dff_A_amCkDlQG0_0),.clk(gclk));
	jdff dff_A_unzlrDbQ0_0(.dout(w_dff_A_amCkDlQG0_0),.din(w_dff_A_unzlrDbQ0_0),.clk(gclk));
	jdff dff_A_DLenJcZs5_0(.dout(w_dff_A_unzlrDbQ0_0),.din(w_dff_A_DLenJcZs5_0),.clk(gclk));
	jdff dff_A_33WDRoqx6_0(.dout(w_dff_A_DLenJcZs5_0),.din(w_dff_A_33WDRoqx6_0),.clk(gclk));
	jdff dff_A_n6XHEdUj8_0(.dout(w_dff_A_33WDRoqx6_0),.din(w_dff_A_n6XHEdUj8_0),.clk(gclk));
	jdff dff_A_aoPBYSjc7_1(.dout(w_G14gat_0[1]),.din(w_dff_A_aoPBYSjc7_1),.clk(gclk));
	jdff dff_A_GVLtgWZY8_1(.dout(w_dff_A_aoPBYSjc7_1),.din(w_dff_A_GVLtgWZY8_1),.clk(gclk));
	jdff dff_A_ONnW7Y279_1(.dout(w_dff_A_GVLtgWZY8_1),.din(w_dff_A_ONnW7Y279_1),.clk(gclk));
	jdff dff_A_TjsBU9JQ2_1(.dout(w_dff_A_ONnW7Y279_1),.din(w_dff_A_TjsBU9JQ2_1),.clk(gclk));
	jdff dff_A_Gd3cNstL9_1(.dout(w_dff_A_TjsBU9JQ2_1),.din(w_dff_A_Gd3cNstL9_1),.clk(gclk));
	jdff dff_A_xsQPmKib1_1(.dout(w_dff_A_Gd3cNstL9_1),.din(w_dff_A_xsQPmKib1_1),.clk(gclk));
	jdff dff_A_P8Drobbj0_1(.dout(w_dff_A_xsQPmKib1_1),.din(w_dff_A_P8Drobbj0_1),.clk(gclk));
	jdff dff_A_d13K1z2Z8_1(.dout(w_dff_A_P8Drobbj0_1),.din(w_dff_A_d13K1z2Z8_1),.clk(gclk));
	jdff dff_A_7CHHER2a3_1(.dout(w_dff_A_d13K1z2Z8_1),.din(w_dff_A_7CHHER2a3_1),.clk(gclk));
	jdff dff_A_fIl2YIaC5_1(.dout(w_dff_A_7CHHER2a3_1),.din(w_dff_A_fIl2YIaC5_1),.clk(gclk));
	jdff dff_A_xUkjWZZx2_1(.dout(w_dff_A_fIl2YIaC5_1),.din(w_dff_A_xUkjWZZx2_1),.clk(gclk));
	jdff dff_A_UQ0gZUMf1_1(.dout(w_dff_A_xUkjWZZx2_1),.din(w_dff_A_UQ0gZUMf1_1),.clk(gclk));
	jdff dff_B_0Fm7J8cP5_0(.din(n207),.dout(w_dff_B_0Fm7J8cP5_0),.clk(gclk));
	jdff dff_B_NB6VqPUe9_0(.din(w_dff_B_0Fm7J8cP5_0),.dout(w_dff_B_NB6VqPUe9_0),.clk(gclk));
	jdff dff_B_OX8CYYjJ6_0(.din(w_dff_B_NB6VqPUe9_0),.dout(w_dff_B_OX8CYYjJ6_0),.clk(gclk));
	jdff dff_A_EZ66K8I56_0(.dout(w_n205_0[0]),.din(w_dff_A_EZ66K8I56_0),.clk(gclk));
	jdff dff_A_QIXAY9WK7_0(.dout(w_dff_A_EZ66K8I56_0),.din(w_dff_A_QIXAY9WK7_0),.clk(gclk));
	jdff dff_A_uC5b3hSA3_0(.dout(w_dff_A_QIXAY9WK7_0),.din(w_dff_A_uC5b3hSA3_0),.clk(gclk));
	jdff dff_A_h4em9AGo8_0(.dout(w_dff_A_uC5b3hSA3_0),.din(w_dff_A_h4em9AGo8_0),.clk(gclk));
	jdff dff_A_tIGfwHGg2_0(.dout(w_dff_A_h4em9AGo8_0),.din(w_dff_A_tIGfwHGg2_0),.clk(gclk));
	jdff dff_A_J8QPLg9J7_0(.dout(w_dff_A_tIGfwHGg2_0),.din(w_dff_A_J8QPLg9J7_0),.clk(gclk));
	jdff dff_A_MFJeeaF62_0(.dout(w_dff_A_J8QPLg9J7_0),.din(w_dff_A_MFJeeaF62_0),.clk(gclk));
	jdff dff_A_1sgwg0GZ7_0(.dout(w_dff_A_MFJeeaF62_0),.din(w_dff_A_1sgwg0GZ7_0),.clk(gclk));
	jdff dff_B_j6icMxLW8_2(.din(n205),.dout(w_dff_B_j6icMxLW8_2),.clk(gclk));
	jdff dff_B_ViB2Df705_2(.din(w_dff_B_j6icMxLW8_2),.dout(w_dff_B_ViB2Df705_2),.clk(gclk));
	jdff dff_B_X6v2frNB4_2(.din(w_dff_B_ViB2Df705_2),.dout(w_dff_B_X6v2frNB4_2),.clk(gclk));
	jdff dff_B_GhwuFCdQ1_2(.din(w_dff_B_X6v2frNB4_2),.dout(w_dff_B_GhwuFCdQ1_2),.clk(gclk));
	jdff dff_B_mQ6TBImH6_2(.din(w_dff_B_GhwuFCdQ1_2),.dout(w_dff_B_mQ6TBImH6_2),.clk(gclk));
	jdff dff_B_T1KCYwbu9_2(.din(w_dff_B_mQ6TBImH6_2),.dout(w_dff_B_T1KCYwbu9_2),.clk(gclk));
	jdff dff_A_ZQM77ijN8_0(.dout(w_G92gat_0[0]),.din(w_dff_A_ZQM77ijN8_0),.clk(gclk));
	jdff dff_A_gLHxr5VE8_0(.dout(w_dff_A_ZQM77ijN8_0),.din(w_dff_A_gLHxr5VE8_0),.clk(gclk));
	jdff dff_A_UH5r1ecC3_0(.dout(w_dff_A_gLHxr5VE8_0),.din(w_dff_A_UH5r1ecC3_0),.clk(gclk));
	jdff dff_A_i1NsmZSa3_0(.dout(w_dff_A_UH5r1ecC3_0),.din(w_dff_A_i1NsmZSa3_0),.clk(gclk));
	jdff dff_A_kUCTXTQI4_0(.dout(w_dff_A_i1NsmZSa3_0),.din(w_dff_A_kUCTXTQI4_0),.clk(gclk));
	jdff dff_A_w64DdZxZ0_0(.dout(w_dff_A_kUCTXTQI4_0),.din(w_dff_A_w64DdZxZ0_0),.clk(gclk));
	jdff dff_A_h2w8RUEb4_0(.dout(w_dff_A_w64DdZxZ0_0),.din(w_dff_A_h2w8RUEb4_0),.clk(gclk));
	jdff dff_A_ZW076xdY9_0(.dout(w_dff_A_h2w8RUEb4_0),.din(w_dff_A_ZW076xdY9_0),.clk(gclk));
	jdff dff_A_7p5qUIwD9_0(.dout(w_dff_A_ZW076xdY9_0),.din(w_dff_A_7p5qUIwD9_0),.clk(gclk));
	jdff dff_A_4DZfS5Xn2_0(.dout(w_dff_A_7p5qUIwD9_0),.din(w_dff_A_4DZfS5Xn2_0),.clk(gclk));
	jdff dff_A_sHGoiaU70_0(.dout(w_dff_A_4DZfS5Xn2_0),.din(w_dff_A_sHGoiaU70_0),.clk(gclk));
	jdff dff_A_T3NsGRQx8_0(.dout(w_dff_A_sHGoiaU70_0),.din(w_dff_A_T3NsGRQx8_0),.clk(gclk));
	jdff dff_A_hMVbeRty0_1(.dout(w_G92gat_0[1]),.din(w_dff_A_hMVbeRty0_1),.clk(gclk));
	jdff dff_A_i0yxT9Qv6_1(.dout(w_dff_A_hMVbeRty0_1),.din(w_dff_A_i0yxT9Qv6_1),.clk(gclk));
	jdff dff_A_Hw8MJEYn1_1(.dout(w_dff_A_i0yxT9Qv6_1),.din(w_dff_A_Hw8MJEYn1_1),.clk(gclk));
	jdff dff_A_yYO2Wevq8_1(.dout(w_dff_A_Hw8MJEYn1_1),.din(w_dff_A_yYO2Wevq8_1),.clk(gclk));
	jdff dff_A_X7C3Aba86_1(.dout(w_dff_A_yYO2Wevq8_1),.din(w_dff_A_X7C3Aba86_1),.clk(gclk));
	jdff dff_A_etXGr1iD5_1(.dout(w_dff_A_X7C3Aba86_1),.din(w_dff_A_etXGr1iD5_1),.clk(gclk));
	jdff dff_A_ct50e6pk0_1(.dout(w_dff_A_etXGr1iD5_1),.din(w_dff_A_ct50e6pk0_1),.clk(gclk));
	jdff dff_A_bVOGG39t0_1(.dout(w_dff_A_ct50e6pk0_1),.din(w_dff_A_bVOGG39t0_1),.clk(gclk));
	jdff dff_A_iYtOsyqy6_1(.dout(w_dff_A_bVOGG39t0_1),.din(w_dff_A_iYtOsyqy6_1),.clk(gclk));
	jdff dff_A_YSMFNW3H9_1(.dout(w_dff_A_iYtOsyqy6_1),.din(w_dff_A_YSMFNW3H9_1),.clk(gclk));
	jdff dff_A_F9SGUW079_1(.dout(w_dff_A_YSMFNW3H9_1),.din(w_dff_A_F9SGUW079_1),.clk(gclk));
	jdff dff_A_9bFtK4IS8_0(.dout(w_n204_0[0]),.din(w_dff_A_9bFtK4IS8_0),.clk(gclk));
	jdff dff_A_OIwkqYyV4_0(.dout(w_dff_A_9bFtK4IS8_0),.din(w_dff_A_OIwkqYyV4_0),.clk(gclk));
	jdff dff_A_ZUT9YEWU6_0(.dout(w_dff_A_OIwkqYyV4_0),.din(w_dff_A_ZUT9YEWU6_0),.clk(gclk));
	jdff dff_A_ZXqWWYqh1_0(.dout(w_dff_A_ZUT9YEWU6_0),.din(w_dff_A_ZXqWWYqh1_0),.clk(gclk));
	jdff dff_B_yha5fpCJ9_1(.din(n195),.dout(w_dff_B_yha5fpCJ9_1),.clk(gclk));
	jdff dff_B_JanIzsh28_1(.din(w_dff_B_yha5fpCJ9_1),.dout(w_dff_B_JanIzsh28_1),.clk(gclk));
	jdff dff_B_YM6zdRQQ9_0(.din(n200),.dout(w_dff_B_YM6zdRQQ9_0),.clk(gclk));
	jdff dff_B_lk5jbvF57_0(.din(w_dff_B_YM6zdRQQ9_0),.dout(w_dff_B_lk5jbvF57_0),.clk(gclk));
	jdff dff_B_RJacCCyX8_0(.din(w_dff_B_lk5jbvF57_0),.dout(w_dff_B_RJacCCyX8_0),.clk(gclk));
	jdff dff_A_otWel9Ab8_0(.dout(w_n198_0[0]),.din(w_dff_A_otWel9Ab8_0),.clk(gclk));
	jdff dff_A_4bvWgYgg2_0(.dout(w_dff_A_otWel9Ab8_0),.din(w_dff_A_4bvWgYgg2_0),.clk(gclk));
	jdff dff_A_vwNK0Yky6_0(.dout(w_dff_A_4bvWgYgg2_0),.din(w_dff_A_vwNK0Yky6_0),.clk(gclk));
	jdff dff_A_jS1q47vm7_0(.dout(w_dff_A_vwNK0Yky6_0),.din(w_dff_A_jS1q47vm7_0),.clk(gclk));
	jdff dff_A_dYdWcGhN9_0(.dout(w_dff_A_jS1q47vm7_0),.din(w_dff_A_dYdWcGhN9_0),.clk(gclk));
	jdff dff_A_Cwm2wRgm1_0(.dout(w_dff_A_dYdWcGhN9_0),.din(w_dff_A_Cwm2wRgm1_0),.clk(gclk));
	jdff dff_A_LjWVac3z9_0(.dout(w_dff_A_Cwm2wRgm1_0),.din(w_dff_A_LjWVac3z9_0),.clk(gclk));
	jdff dff_A_lvyuG3S28_0(.dout(w_dff_A_LjWVac3z9_0),.din(w_dff_A_lvyuG3S28_0),.clk(gclk));
	jdff dff_B_hCMkpj2D8_2(.din(n198),.dout(w_dff_B_hCMkpj2D8_2),.clk(gclk));
	jdff dff_B_lMUpE1dq4_2(.din(w_dff_B_hCMkpj2D8_2),.dout(w_dff_B_lMUpE1dq4_2),.clk(gclk));
	jdff dff_B_ApHbSPsA1_2(.din(w_dff_B_lMUpE1dq4_2),.dout(w_dff_B_ApHbSPsA1_2),.clk(gclk));
	jdff dff_B_80e3dtk22_2(.din(w_dff_B_ApHbSPsA1_2),.dout(w_dff_B_80e3dtk22_2),.clk(gclk));
	jdff dff_B_8KIQ7lgq9_2(.din(w_dff_B_80e3dtk22_2),.dout(w_dff_B_8KIQ7lgq9_2),.clk(gclk));
	jdff dff_B_gn2lZ5EV5_2(.din(w_dff_B_8KIQ7lgq9_2),.dout(w_dff_B_gn2lZ5EV5_2),.clk(gclk));
	jdff dff_A_yTMzwNf05_0(.dout(w_G27gat_0[0]),.din(w_dff_A_yTMzwNf05_0),.clk(gclk));
	jdff dff_A_8uQ57ghq4_0(.dout(w_dff_A_yTMzwNf05_0),.din(w_dff_A_8uQ57ghq4_0),.clk(gclk));
	jdff dff_A_cqIW7l3Z6_0(.dout(w_dff_A_8uQ57ghq4_0),.din(w_dff_A_cqIW7l3Z6_0),.clk(gclk));
	jdff dff_A_i7h7aHMk0_0(.dout(w_dff_A_cqIW7l3Z6_0),.din(w_dff_A_i7h7aHMk0_0),.clk(gclk));
	jdff dff_A_OXIsrcsI1_0(.dout(w_dff_A_i7h7aHMk0_0),.din(w_dff_A_OXIsrcsI1_0),.clk(gclk));
	jdff dff_A_Pwv98ANR5_0(.dout(w_dff_A_OXIsrcsI1_0),.din(w_dff_A_Pwv98ANR5_0),.clk(gclk));
	jdff dff_A_8V1RKfWy8_0(.dout(w_dff_A_Pwv98ANR5_0),.din(w_dff_A_8V1RKfWy8_0),.clk(gclk));
	jdff dff_A_pGQcxazk7_0(.dout(w_dff_A_8V1RKfWy8_0),.din(w_dff_A_pGQcxazk7_0),.clk(gclk));
	jdff dff_A_qttq73nH6_0(.dout(w_dff_A_pGQcxazk7_0),.din(w_dff_A_qttq73nH6_0),.clk(gclk));
	jdff dff_A_7MLCmt1f9_0(.dout(w_dff_A_qttq73nH6_0),.din(w_dff_A_7MLCmt1f9_0),.clk(gclk));
	jdff dff_A_A3IUWPZP3_0(.dout(w_dff_A_7MLCmt1f9_0),.din(w_dff_A_A3IUWPZP3_0),.clk(gclk));
	jdff dff_A_flv45uwV2_0(.dout(w_n197_0[0]),.din(w_dff_A_flv45uwV2_0),.clk(gclk));
	jdff dff_A_8hk90B1W0_0(.dout(w_dff_A_flv45uwV2_0),.din(w_dff_A_8hk90B1W0_0),.clk(gclk));
	jdff dff_A_lTONVAEu1_0(.dout(w_dff_A_8hk90B1W0_0),.din(w_dff_A_lTONVAEu1_0),.clk(gclk));
	jdff dff_A_BNcYI1jW3_0(.dout(w_dff_A_lTONVAEu1_0),.din(w_dff_A_BNcYI1jW3_0),.clk(gclk));
	jdff dff_A_CTsZFhOj0_1(.dout(w_n193_0[1]),.din(w_dff_A_CTsZFhOj0_1),.clk(gclk));
	jdff dff_A_aZStHclE5_1(.dout(w_dff_A_CTsZFhOj0_1),.din(w_dff_A_aZStHclE5_1),.clk(gclk));
	jdff dff_B_94FtYurF3_0(.din(n192),.dout(w_dff_B_94FtYurF3_0),.clk(gclk));
	jdff dff_B_dPRfy0Oi2_0(.din(w_dff_B_94FtYurF3_0),.dout(w_dff_B_dPRfy0Oi2_0),.clk(gclk));
	jdff dff_B_s94aZ1uZ9_0(.din(w_dff_B_dPRfy0Oi2_0),.dout(w_dff_B_s94aZ1uZ9_0),.clk(gclk));
	jdff dff_B_e0UwjMc36_0(.din(w_dff_B_s94aZ1uZ9_0),.dout(w_dff_B_e0UwjMc36_0),.clk(gclk));
	jdff dff_A_euxpM8qG3_0(.dout(w_n191_0[0]),.din(w_dff_A_euxpM8qG3_0),.clk(gclk));
	jdff dff_A_uDc6K0OK8_0(.dout(w_dff_A_euxpM8qG3_0),.din(w_dff_A_uDc6K0OK8_0),.clk(gclk));
	jdff dff_A_Xpzl2Exo1_0(.dout(w_dff_A_uDc6K0OK8_0),.din(w_dff_A_Xpzl2Exo1_0),.clk(gclk));
	jdff dff_A_XEUslydH8_0(.dout(w_dff_A_Xpzl2Exo1_0),.din(w_dff_A_XEUslydH8_0),.clk(gclk));
	jdff dff_A_zAmybL963_0(.dout(w_dff_A_XEUslydH8_0),.din(w_dff_A_zAmybL963_0),.clk(gclk));
	jdff dff_A_WaC0xmkI5_0(.dout(w_dff_A_zAmybL963_0),.din(w_dff_A_WaC0xmkI5_0),.clk(gclk));
	jdff dff_A_lZKOxCBE9_0(.dout(w_dff_A_WaC0xmkI5_0),.din(w_dff_A_lZKOxCBE9_0),.clk(gclk));
	jdff dff_A_Co4vapyC6_0(.dout(w_dff_A_lZKOxCBE9_0),.din(w_dff_A_Co4vapyC6_0),.clk(gclk));
	jdff dff_A_U5NXQK7T8_0(.dout(w_dff_A_Co4vapyC6_0),.din(w_dff_A_U5NXQK7T8_0),.clk(gclk));
	jdff dff_A_wl7cV57o1_0(.dout(w_dff_A_U5NXQK7T8_0),.din(w_dff_A_wl7cV57o1_0),.clk(gclk));
	jdff dff_A_F2ypEOLn8_0(.dout(w_dff_A_wl7cV57o1_0),.din(w_dff_A_F2ypEOLn8_0),.clk(gclk));
	jdff dff_A_vjRiOPuB4_0(.dout(w_dff_A_F2ypEOLn8_0),.din(w_dff_A_vjRiOPuB4_0),.clk(gclk));
	jdff dff_A_oAQZktvN8_0(.dout(w_dff_A_vjRiOPuB4_0),.din(w_dff_A_oAQZktvN8_0),.clk(gclk));
	jdff dff_A_4hKiCFt56_0(.dout(w_dff_A_oAQZktvN8_0),.din(w_dff_A_4hKiCFt56_0),.clk(gclk));
	jdff dff_A_Tkq26vvM1_0(.dout(w_G53gat_0[0]),.din(w_dff_A_Tkq26vvM1_0),.clk(gclk));
	jdff dff_A_NM4lVzEs6_0(.dout(w_dff_A_Tkq26vvM1_0),.din(w_dff_A_NM4lVzEs6_0),.clk(gclk));
	jdff dff_A_y0w11bp89_0(.dout(w_dff_A_NM4lVzEs6_0),.din(w_dff_A_y0w11bp89_0),.clk(gclk));
	jdff dff_A_o1lx5Zeh3_0(.dout(w_dff_A_y0w11bp89_0),.din(w_dff_A_o1lx5Zeh3_0),.clk(gclk));
	jdff dff_A_FwWBv6J41_0(.dout(w_dff_A_o1lx5Zeh3_0),.din(w_dff_A_FwWBv6J41_0),.clk(gclk));
	jdff dff_A_PRHZWjfF4_0(.dout(w_dff_A_FwWBv6J41_0),.din(w_dff_A_PRHZWjfF4_0),.clk(gclk));
	jdff dff_A_Og0IvzaN0_0(.dout(w_dff_A_PRHZWjfF4_0),.din(w_dff_A_Og0IvzaN0_0),.clk(gclk));
	jdff dff_A_CVbHa7rN5_0(.dout(w_dff_A_Og0IvzaN0_0),.din(w_dff_A_CVbHa7rN5_0),.clk(gclk));
	jdff dff_A_kje4BfZV4_0(.dout(w_dff_A_CVbHa7rN5_0),.din(w_dff_A_kje4BfZV4_0),.clk(gclk));
	jdff dff_A_JlmQPkRc7_0(.dout(w_dff_A_kje4BfZV4_0),.din(w_dff_A_JlmQPkRc7_0),.clk(gclk));
	jdff dff_A_7Z8y3gVK5_0(.dout(w_dff_A_JlmQPkRc7_0),.din(w_dff_A_7Z8y3gVK5_0),.clk(gclk));
	jdff dff_A_Azx8s1LO1_0(.dout(w_dff_A_7Z8y3gVK5_0),.din(w_dff_A_Azx8s1LO1_0),.clk(gclk));
	jdff dff_B_RoMW8FnH0_1(.din(n143),.dout(w_dff_B_RoMW8FnH0_1),.clk(gclk));
	jdff dff_B_HtIDmsE94_1(.din(w_dff_B_RoMW8FnH0_1),.dout(w_dff_B_HtIDmsE94_1),.clk(gclk));
	jdff dff_B_tAdIrQVR3_1(.din(w_dff_B_HtIDmsE94_1),.dout(w_dff_B_tAdIrQVR3_1),.clk(gclk));
	jdff dff_B_CUo1k0AK5_1(.din(n153),.dout(w_dff_B_CUo1k0AK5_1),.clk(gclk));
	jdff dff_B_4wmQmU9N4_1(.din(w_dff_B_CUo1k0AK5_1),.dout(w_dff_B_4wmQmU9N4_1),.clk(gclk));
	jdff dff_A_N9RnvfVd9_0(.dout(w_n184_0[0]),.din(w_dff_A_N9RnvfVd9_0),.clk(gclk));
	jdff dff_A_v5evyWm53_0(.dout(w_dff_A_N9RnvfVd9_0),.din(w_dff_A_v5evyWm53_0),.clk(gclk));
	jdff dff_A_OLtuKuaT3_0(.dout(w_dff_A_v5evyWm53_0),.din(w_dff_A_OLtuKuaT3_0),.clk(gclk));
	jdff dff_A_yjadT7ge8_0(.dout(w_dff_A_OLtuKuaT3_0),.din(w_dff_A_yjadT7ge8_0),.clk(gclk));
	jdff dff_B_BfUpeLkb6_1(.din(n167),.dout(w_dff_B_BfUpeLkb6_1),.clk(gclk));
	jdff dff_B_bDjw6hKi6_1(.din(w_dff_B_BfUpeLkb6_1),.dout(w_dff_B_bDjw6hKi6_1),.clk(gclk));
	jdff dff_B_PRYKRpCi3_1(.din(w_dff_B_bDjw6hKi6_1),.dout(w_dff_B_PRYKRpCi3_1),.clk(gclk));
	jdff dff_B_LcjHbqcO6_1(.din(w_dff_B_PRYKRpCi3_1),.dout(w_dff_B_LcjHbqcO6_1),.clk(gclk));
	jdff dff_B_ahmtxd9L6_0(.din(n179),.dout(w_dff_B_ahmtxd9L6_0),.clk(gclk));
	jdff dff_B_UUwDZErp8_0(.din(w_dff_B_ahmtxd9L6_0),.dout(w_dff_B_UUwDZErp8_0),.clk(gclk));
	jdff dff_B_kYUNMXF78_0(.din(w_dff_B_UUwDZErp8_0),.dout(w_dff_B_kYUNMXF78_0),.clk(gclk));
	jdff dff_A_qedJcAie1_0(.dout(w_n177_0[0]),.din(w_dff_A_qedJcAie1_0),.clk(gclk));
	jdff dff_A_5xI6FYCb3_0(.dout(w_dff_A_qedJcAie1_0),.din(w_dff_A_5xI6FYCb3_0),.clk(gclk));
	jdff dff_A_kCt4opwe3_0(.dout(w_dff_A_5xI6FYCb3_0),.din(w_dff_A_kCt4opwe3_0),.clk(gclk));
	jdff dff_A_7hBtspxo9_0(.dout(w_dff_A_kCt4opwe3_0),.din(w_dff_A_7hBtspxo9_0),.clk(gclk));
	jdff dff_A_PK1iZVts9_0(.dout(w_dff_A_7hBtspxo9_0),.din(w_dff_A_PK1iZVts9_0),.clk(gclk));
	jdff dff_A_WKMAoyGh9_0(.dout(w_n174_0[0]),.din(w_dff_A_WKMAoyGh9_0),.clk(gclk));
	jdff dff_A_GEBICV0d9_0(.dout(w_dff_A_WKMAoyGh9_0),.din(w_dff_A_GEBICV0d9_0),.clk(gclk));
	jdff dff_A_xxkv2tFz2_0(.dout(w_dff_A_GEBICV0d9_0),.din(w_dff_A_xxkv2tFz2_0),.clk(gclk));
	jdff dff_A_OcNDm2Cr7_0(.dout(w_dff_A_xxkv2tFz2_0),.din(w_dff_A_OcNDm2Cr7_0),.clk(gclk));
	jdff dff_A_amCOZp3N3_0(.dout(w_dff_A_OcNDm2Cr7_0),.din(w_dff_A_amCOZp3N3_0),.clk(gclk));
	jdff dff_B_kmbGbOWT9_1(.din(n172),.dout(w_dff_B_kmbGbOWT9_1),.clk(gclk));
	jdff dff_B_xONieWA89_1(.din(w_dff_B_kmbGbOWT9_1),.dout(w_dff_B_xONieWA89_1),.clk(gclk));
	jdff dff_A_45LdLgW39_0(.dout(w_n170_0[0]),.din(w_dff_A_45LdLgW39_0),.clk(gclk));
	jdff dff_B_16gvVIQX6_0(.din(n169),.dout(w_dff_B_16gvVIQX6_0),.clk(gclk));
	jdff dff_B_dqwQiNEy2_0(.din(w_dff_B_16gvVIQX6_0),.dout(w_dff_B_dqwQiNEy2_0),.clk(gclk));
	jdff dff_B_4tnmKcOD0_0(.din(w_dff_B_dqwQiNEy2_0),.dout(w_dff_B_4tnmKcOD0_0),.clk(gclk));
	jdff dff_A_51j4moIv4_0(.dout(w_n164_0[0]),.din(w_dff_A_51j4moIv4_0),.clk(gclk));
	jdff dff_A_IGXwJl4N5_0(.dout(w_dff_A_51j4moIv4_0),.din(w_dff_A_IGXwJl4N5_0),.clk(gclk));
	jdff dff_A_BjmicdfJ7_0(.dout(w_dff_A_IGXwJl4N5_0),.din(w_dff_A_BjmicdfJ7_0),.clk(gclk));
	jdff dff_A_SXsHS5Nr3_0(.dout(w_dff_A_BjmicdfJ7_0),.din(w_dff_A_SXsHS5Nr3_0),.clk(gclk));
	jdff dff_A_Im4Zx6Q98_0(.dout(w_dff_A_SXsHS5Nr3_0),.din(w_dff_A_Im4Zx6Q98_0),.clk(gclk));
	jdff dff_A_pcrO7N6p0_0(.dout(w_n159_0[0]),.din(w_dff_A_pcrO7N6p0_0),.clk(gclk));
	jdff dff_A_Kp35cWIA9_0(.dout(w_dff_A_pcrO7N6p0_0),.din(w_dff_A_Kp35cWIA9_0),.clk(gclk));
	jdff dff_A_rzK6xVI06_0(.dout(w_dff_A_Kp35cWIA9_0),.din(w_dff_A_rzK6xVI06_0),.clk(gclk));
	jdff dff_A_HijxTHh74_0(.dout(w_dff_A_rzK6xVI06_0),.din(w_dff_A_HijxTHh74_0),.clk(gclk));
	jdff dff_A_pqUeLYjz8_0(.dout(w_dff_A_HijxTHh74_0),.din(w_dff_A_pqUeLYjz8_0),.clk(gclk));
	jdff dff_A_rj2cDQlh2_0(.dout(w_n156_0[0]),.din(w_dff_A_rj2cDQlh2_0),.clk(gclk));
	jdff dff_A_gspv3eSZ3_0(.dout(w_dff_A_rj2cDQlh2_0),.din(w_dff_A_gspv3eSZ3_0),.clk(gclk));
	jdff dff_A_OEAQYrDn7_0(.dout(w_dff_A_gspv3eSZ3_0),.din(w_dff_A_OEAQYrDn7_0),.clk(gclk));
	jdff dff_A_kNaO7n3e3_0(.dout(w_dff_A_OEAQYrDn7_0),.din(w_dff_A_kNaO7n3e3_0),.clk(gclk));
	jdff dff_A_sO1JVLwy0_0(.dout(w_dff_A_kNaO7n3e3_0),.din(w_dff_A_sO1JVLwy0_0),.clk(gclk));
	jdff dff_A_BCX9q4bR9_0(.dout(w_n154_0[0]),.din(w_dff_A_BCX9q4bR9_0),.clk(gclk));
	jdff dff_A_qru0Po659_0(.dout(w_dff_A_BCX9q4bR9_0),.din(w_dff_A_qru0Po659_0),.clk(gclk));
	jdff dff_A_JrGztQ1P5_0(.dout(w_dff_A_qru0Po659_0),.din(w_dff_A_JrGztQ1P5_0),.clk(gclk));
	jdff dff_A_ygsYRx3b7_0(.dout(w_dff_A_JrGztQ1P5_0),.din(w_dff_A_ygsYRx3b7_0),.clk(gclk));
	jdff dff_B_mMGdF3hJ9_2(.din(n154),.dout(w_dff_B_mMGdF3hJ9_2),.clk(gclk));
	jdff dff_B_j8uXlFgC4_2(.din(w_dff_B_mMGdF3hJ9_2),.dout(w_dff_B_j8uXlFgC4_2),.clk(gclk));
	jdff dff_B_ElnPzp5u5_2(.din(w_dff_B_j8uXlFgC4_2),.dout(w_dff_B_ElnPzp5u5_2),.clk(gclk));
	jdff dff_B_sXxwHUdg3_2(.din(w_dff_B_ElnPzp5u5_2),.dout(w_dff_B_sXxwHUdg3_2),.clk(gclk));
	jdff dff_B_ZzIRq4707_2(.din(w_dff_B_sXxwHUdg3_2),.dout(w_dff_B_ZzIRq4707_2),.clk(gclk));
	jdff dff_B_xxngIuti1_2(.din(w_dff_B_ZzIRq4707_2),.dout(w_dff_B_xxngIuti1_2),.clk(gclk));
	jdff dff_B_y1WVhjcL2_2(.din(w_dff_B_xxngIuti1_2),.dout(w_dff_B_y1WVhjcL2_2),.clk(gclk));
	jdff dff_B_y6fsy1og2_2(.din(w_dff_B_y1WVhjcL2_2),.dout(w_dff_B_y6fsy1og2_2),.clk(gclk));
	jdff dff_B_tCHJSG9R8_2(.din(w_dff_B_y6fsy1og2_2),.dout(w_dff_B_tCHJSG9R8_2),.clk(gclk));
	jdff dff_B_vPY4wFJg5_2(.din(w_dff_B_tCHJSG9R8_2),.dout(w_dff_B_vPY4wFJg5_2),.clk(gclk));
	jdff dff_A_9ctAOboP5_0(.dout(w_G79gat_0[0]),.din(w_dff_A_9ctAOboP5_0),.clk(gclk));
	jdff dff_A_Sgezy1ZD9_0(.dout(w_dff_A_9ctAOboP5_0),.din(w_dff_A_Sgezy1ZD9_0),.clk(gclk));
	jdff dff_A_wNHs7BF89_0(.dout(w_dff_A_Sgezy1ZD9_0),.din(w_dff_A_wNHs7BF89_0),.clk(gclk));
	jdff dff_A_K7qbLHhz0_0(.dout(w_dff_A_wNHs7BF89_0),.din(w_dff_A_K7qbLHhz0_0),.clk(gclk));
	jdff dff_A_JwycmPio6_0(.dout(w_dff_A_K7qbLHhz0_0),.din(w_dff_A_JwycmPio6_0),.clk(gclk));
	jdff dff_A_NjnZNVek5_0(.dout(w_dff_A_JwycmPio6_0),.din(w_dff_A_NjnZNVek5_0),.clk(gclk));
	jdff dff_A_N7OVrmsV2_0(.dout(w_dff_A_NjnZNVek5_0),.din(w_dff_A_N7OVrmsV2_0),.clk(gclk));
	jdff dff_A_6ukVAaVQ2_0(.dout(w_dff_A_N7OVrmsV2_0),.din(w_dff_A_6ukVAaVQ2_0),.clk(gclk));
	jdff dff_A_fMMmZkVI5_1(.dout(w_n151_0[1]),.din(w_dff_A_fMMmZkVI5_1),.clk(gclk));
	jdff dff_A_ErzZilkO7_1(.dout(w_dff_A_fMMmZkVI5_1),.din(w_dff_A_ErzZilkO7_1),.clk(gclk));
	jdff dff_A_7HH9ZPhQ7_0(.dout(w_n150_0[0]),.din(w_dff_A_7HH9ZPhQ7_0),.clk(gclk));
	jdff dff_A_G7dKXof11_0(.dout(w_dff_A_7HH9ZPhQ7_0),.din(w_dff_A_G7dKXof11_0),.clk(gclk));
	jdff dff_A_zN5Gn6sK1_0(.dout(w_dff_A_G7dKXof11_0),.din(w_dff_A_zN5Gn6sK1_0),.clk(gclk));
	jdff dff_A_H3mov8WQ6_0(.dout(w_dff_A_zN5Gn6sK1_0),.din(w_dff_A_H3mov8WQ6_0),.clk(gclk));
	jdff dff_A_4B4Ax9XZ3_0(.dout(w_dff_A_H3mov8WQ6_0),.din(w_dff_A_4B4Ax9XZ3_0),.clk(gclk));
	jdff dff_A_3igUQjgO4_0(.dout(w_dff_A_4B4Ax9XZ3_0),.din(w_dff_A_3igUQjgO4_0),.clk(gclk));
	jdff dff_A_u46OFi9Y9_0(.dout(w_dff_A_3igUQjgO4_0),.din(w_dff_A_u46OFi9Y9_0),.clk(gclk));
	jdff dff_A_5SMsCezM6_0(.dout(w_dff_A_u46OFi9Y9_0),.din(w_dff_A_5SMsCezM6_0),.clk(gclk));
	jdff dff_A_gmRkcWga9_0(.dout(w_dff_A_5SMsCezM6_0),.din(w_dff_A_gmRkcWga9_0),.clk(gclk));
	jdff dff_B_0cKDbo398_2(.din(n150),.dout(w_dff_B_0cKDbo398_2),.clk(gclk));
	jdff dff_B_hK7q5ME77_2(.din(w_dff_B_0cKDbo398_2),.dout(w_dff_B_hK7q5ME77_2),.clk(gclk));
	jdff dff_B_V9hL6yDC8_2(.din(w_dff_B_hK7q5ME77_2),.dout(w_dff_B_V9hL6yDC8_2),.clk(gclk));
	jdff dff_B_Hr3aWMtA7_2(.din(w_dff_B_V9hL6yDC8_2),.dout(w_dff_B_Hr3aWMtA7_2),.clk(gclk));
	jdff dff_B_2xp4turu3_2(.din(w_dff_B_Hr3aWMtA7_2),.dout(w_dff_B_2xp4turu3_2),.clk(gclk));
	jdff dff_A_IemfyM1A4_0(.dout(w_G66gat_0[0]),.din(w_dff_A_IemfyM1A4_0),.clk(gclk));
	jdff dff_A_h0YWiSR97_0(.dout(w_dff_A_IemfyM1A4_0),.din(w_dff_A_h0YWiSR97_0),.clk(gclk));
	jdff dff_A_TRtyb1yV4_0(.dout(w_dff_A_h0YWiSR97_0),.din(w_dff_A_TRtyb1yV4_0),.clk(gclk));
	jdff dff_A_D9worTUj9_0(.dout(w_dff_A_TRtyb1yV4_0),.din(w_dff_A_D9worTUj9_0),.clk(gclk));
	jdff dff_A_Ha33DfY80_0(.dout(w_dff_A_D9worTUj9_0),.din(w_dff_A_Ha33DfY80_0),.clk(gclk));
	jdff dff_A_Ss42PQcG9_0(.dout(w_dff_A_Ha33DfY80_0),.din(w_dff_A_Ss42PQcG9_0),.clk(gclk));
	jdff dff_A_PRuzpXi84_0(.dout(w_dff_A_Ss42PQcG9_0),.din(w_dff_A_PRuzpXi84_0),.clk(gclk));
	jdff dff_A_NxZ1ansZ3_0(.dout(w_dff_A_PRuzpXi84_0),.din(w_dff_A_NxZ1ansZ3_0),.clk(gclk));
	jdff dff_A_YO0lsnOw4_0(.dout(w_dff_A_NxZ1ansZ3_0),.din(w_dff_A_YO0lsnOw4_0),.clk(gclk));
	jdff dff_A_Mij1yVR26_0(.dout(w_dff_A_YO0lsnOw4_0),.din(w_dff_A_Mij1yVR26_0),.clk(gclk));
	jdff dff_A_YrPtC6Qu3_0(.dout(w_dff_A_Mij1yVR26_0),.din(w_dff_A_YrPtC6Qu3_0),.clk(gclk));
	jdff dff_A_98gxp4xM3_0(.dout(w_dff_A_YrPtC6Qu3_0),.din(w_dff_A_98gxp4xM3_0),.clk(gclk));
	jdff dff_A_ThHCmN9U9_1(.dout(w_n146_0[1]),.din(w_dff_A_ThHCmN9U9_1),.clk(gclk));
	jdff dff_B_PfcDVYKc0_2(.din(n146),.dout(w_dff_B_PfcDVYKc0_2),.clk(gclk));
	jdff dff_B_ngZQ1Hzr1_2(.din(w_dff_B_PfcDVYKc0_2),.dout(w_dff_B_ngZQ1Hzr1_2),.clk(gclk));
	jdff dff_B_AvNIJiip3_2(.din(w_dff_B_ngZQ1Hzr1_2),.dout(w_dff_B_AvNIJiip3_2),.clk(gclk));
	jdff dff_A_gRzdTXiH8_0(.dout(w_n145_0[0]),.din(w_dff_A_gRzdTXiH8_0),.clk(gclk));
	jdff dff_A_60aJI0iE4_0(.dout(w_dff_A_gRzdTXiH8_0),.din(w_dff_A_60aJI0iE4_0),.clk(gclk));
	jdff dff_A_slz6LnE38_0(.dout(w_dff_A_60aJI0iE4_0),.din(w_dff_A_slz6LnE38_0),.clk(gclk));
	jdff dff_A_y5QS8XdQ4_0(.dout(w_dff_A_slz6LnE38_0),.din(w_dff_A_y5QS8XdQ4_0),.clk(gclk));
	jdff dff_A_rkrCP9Nh7_0(.dout(w_dff_A_y5QS8XdQ4_0),.din(w_dff_A_rkrCP9Nh7_0),.clk(gclk));
	jdff dff_A_DBLhnoT00_0(.dout(w_n142_0[0]),.din(w_dff_A_DBLhnoT00_0),.clk(gclk));
	jdff dff_A_687nKNvu5_0(.dout(w_n132_0[0]),.din(w_dff_A_687nKNvu5_0),.clk(gclk));
	jdff dff_A_Dv6BYRCd0_0(.dout(w_dff_A_687nKNvu5_0),.din(w_dff_A_Dv6BYRCd0_0),.clk(gclk));
	jdff dff_A_eS3giYuP3_0(.dout(w_dff_A_Dv6BYRCd0_0),.din(w_dff_A_eS3giYuP3_0),.clk(gclk));
	jdff dff_A_qZrV8PM09_0(.dout(w_dff_A_eS3giYuP3_0),.din(w_dff_A_qZrV8PM09_0),.clk(gclk));
	jdff dff_A_F46ApbvD1_0(.dout(w_n130_0[0]),.din(w_dff_A_F46ApbvD1_0),.clk(gclk));
	jdff dff_A_6uo0edn53_0(.dout(w_dff_A_F46ApbvD1_0),.din(w_dff_A_6uo0edn53_0),.clk(gclk));
	jdff dff_A_hCQ3erfp1_0(.dout(w_dff_A_6uo0edn53_0),.din(w_dff_A_hCQ3erfp1_0),.clk(gclk));
	jdff dff_A_OqN5NvHD9_0(.dout(w_dff_A_hCQ3erfp1_0),.din(w_dff_A_OqN5NvHD9_0),.clk(gclk));
	jdff dff_A_01WeINRc4_1(.dout(w_n130_0[1]),.din(w_dff_A_01WeINRc4_1),.clk(gclk));
	jdff dff_A_0zNXGn6v8_1(.dout(w_dff_A_01WeINRc4_1),.din(w_dff_A_0zNXGn6v8_1),.clk(gclk));
	jdff dff_A_FY84Pajv3_1(.dout(w_dff_A_0zNXGn6v8_1),.din(w_dff_A_FY84Pajv3_1),.clk(gclk));
	jdff dff_A_PIFyp6Mc1_1(.dout(w_dff_A_FY84Pajv3_1),.din(w_dff_A_PIFyp6Mc1_1),.clk(gclk));
	jdff dff_B_dh5i1UYv0_3(.din(n130),.dout(w_dff_B_dh5i1UYv0_3),.clk(gclk));
	jdff dff_B_Mvf6uajc4_3(.din(w_dff_B_dh5i1UYv0_3),.dout(w_dff_B_Mvf6uajc4_3),.clk(gclk));
	jdff dff_B_LLA56UmP6_3(.din(w_dff_B_Mvf6uajc4_3),.dout(w_dff_B_LLA56UmP6_3),.clk(gclk));
	jdff dff_B_Dq1UPj7x4_3(.din(w_dff_B_LLA56UmP6_3),.dout(w_dff_B_Dq1UPj7x4_3),.clk(gclk));
	jdff dff_B_2zO58puS2_3(.din(w_dff_B_Dq1UPj7x4_3),.dout(w_dff_B_2zO58puS2_3),.clk(gclk));
	jdff dff_A_stysf4x63_0(.dout(w_G21gat_1[0]),.din(w_dff_A_stysf4x63_0),.clk(gclk));
	jdff dff_A_ZzbkiKXP8_0(.dout(w_dff_A_stysf4x63_0),.din(w_dff_A_ZzbkiKXP8_0),.clk(gclk));
	jdff dff_A_qDqggfUI9_0(.dout(w_dff_A_ZzbkiKXP8_0),.din(w_dff_A_qDqggfUI9_0),.clk(gclk));
	jdff dff_A_RgXeAOyg4_1(.dout(w_G21gat_0[1]),.din(w_dff_A_RgXeAOyg4_1),.clk(gclk));
	jdff dff_A_gjPjgQxL4_1(.dout(w_dff_A_RgXeAOyg4_1),.din(w_dff_A_gjPjgQxL4_1),.clk(gclk));
	jdff dff_A_e5jZYph45_1(.dout(w_dff_A_gjPjgQxL4_1),.din(w_dff_A_e5jZYph45_1),.clk(gclk));
	jdff dff_A_5T9DzNF45_1(.dout(w_dff_A_e5jZYph45_1),.din(w_dff_A_5T9DzNF45_1),.clk(gclk));
	jdff dff_A_E9EqQVzh5_1(.dout(w_dff_A_5T9DzNF45_1),.din(w_dff_A_E9EqQVzh5_1),.clk(gclk));
	jdff dff_A_Xg4AYU0B8_1(.dout(w_dff_A_E9EqQVzh5_1),.din(w_dff_A_Xg4AYU0B8_1),.clk(gclk));
	jdff dff_A_lB43AEcG3_1(.dout(w_dff_A_Xg4AYU0B8_1),.din(w_dff_A_lB43AEcG3_1),.clk(gclk));
	jdff dff_A_HLQlrUyS4_2(.dout(w_G21gat_0[2]),.din(w_dff_A_HLQlrUyS4_2),.clk(gclk));
	jdff dff_A_VRX6WUSF8_2(.dout(w_dff_A_HLQlrUyS4_2),.din(w_dff_A_VRX6WUSF8_2),.clk(gclk));
	jdff dff_A_I4sHbNO93_2(.dout(w_dff_A_VRX6WUSF8_2),.din(w_dff_A_I4sHbNO93_2),.clk(gclk));
	jdff dff_A_ae1AmbqQ3_2(.dout(w_dff_A_I4sHbNO93_2),.din(w_dff_A_ae1AmbqQ3_2),.clk(gclk));
	jdff dff_A_1dAyMAjO7_2(.dout(w_dff_A_ae1AmbqQ3_2),.din(w_dff_A_1dAyMAjO7_2),.clk(gclk));
	jdff dff_A_0SmGn8rt8_2(.dout(w_dff_A_1dAyMAjO7_2),.din(w_dff_A_0SmGn8rt8_2),.clk(gclk));
	jdff dff_A_Ys6RiXrh8_2(.dout(w_dff_A_0SmGn8rt8_2),.din(w_dff_A_Ys6RiXrh8_2),.clk(gclk));
	jdff dff_A_N5aIXP5K9_0(.dout(w_n128_0[0]),.din(w_dff_A_N5aIXP5K9_0),.clk(gclk));
	jdff dff_A_QfhYA8MQ7_0(.dout(w_dff_A_N5aIXP5K9_0),.din(w_dff_A_QfhYA8MQ7_0),.clk(gclk));
	jdff dff_A_TADIeDG23_0(.dout(w_dff_A_QfhYA8MQ7_0),.din(w_dff_A_TADIeDG23_0),.clk(gclk));
	jdff dff_A_GS2qVlTL6_0(.dout(w_dff_A_TADIeDG23_0),.din(w_dff_A_GS2qVlTL6_0),.clk(gclk));
	jdff dff_A_Esef1Cy66_0(.dout(w_n126_0[0]),.din(w_dff_A_Esef1Cy66_0),.clk(gclk));
	jdff dff_A_qNSIVEWK5_0(.dout(w_dff_A_Esef1Cy66_0),.din(w_dff_A_qNSIVEWK5_0),.clk(gclk));
	jdff dff_A_NQYZ3OtY0_0(.dout(w_dff_A_qNSIVEWK5_0),.din(w_dff_A_NQYZ3OtY0_0),.clk(gclk));
	jdff dff_A_AuCjO2Rd0_0(.dout(w_dff_A_NQYZ3OtY0_0),.din(w_dff_A_AuCjO2Rd0_0),.clk(gclk));
	jdff dff_A_rzcpK0X44_1(.dout(w_n126_0[1]),.din(w_dff_A_rzcpK0X44_1),.clk(gclk));
	jdff dff_A_RveaSCQI7_1(.dout(w_dff_A_rzcpK0X44_1),.din(w_dff_A_RveaSCQI7_1),.clk(gclk));
	jdff dff_A_lcaJCISS7_1(.dout(w_dff_A_RveaSCQI7_1),.din(w_dff_A_lcaJCISS7_1),.clk(gclk));
	jdff dff_A_Q5I9TeQr4_1(.dout(w_dff_A_lcaJCISS7_1),.din(w_dff_A_Q5I9TeQr4_1),.clk(gclk));
	jdff dff_B_iHX2EVeZ1_3(.din(n126),.dout(w_dff_B_iHX2EVeZ1_3),.clk(gclk));
	jdff dff_B_mrxKIk5a2_3(.din(w_dff_B_iHX2EVeZ1_3),.dout(w_dff_B_mrxKIk5a2_3),.clk(gclk));
	jdff dff_B_diEUpV051_3(.din(w_dff_B_mrxKIk5a2_3),.dout(w_dff_B_diEUpV051_3),.clk(gclk));
	jdff dff_B_WzroyfKe4_3(.din(w_dff_B_diEUpV051_3),.dout(w_dff_B_WzroyfKe4_3),.clk(gclk));
	jdff dff_B_2BcIh0H47_3(.din(w_dff_B_WzroyfKe4_3),.dout(w_dff_B_2BcIh0H47_3),.clk(gclk));
	jdff dff_A_KCWSiRUj0_0(.dout(w_G86gat_1[0]),.din(w_dff_A_KCWSiRUj0_0),.clk(gclk));
	jdff dff_A_jdfQKXCQ2_0(.dout(w_dff_A_KCWSiRUj0_0),.din(w_dff_A_jdfQKXCQ2_0),.clk(gclk));
	jdff dff_A_K5bHggug5_0(.dout(w_dff_A_jdfQKXCQ2_0),.din(w_dff_A_K5bHggug5_0),.clk(gclk));
	jdff dff_A_BSIq8CKJ4_1(.dout(w_G86gat_0[1]),.din(w_dff_A_BSIq8CKJ4_1),.clk(gclk));
	jdff dff_A_1LQ596uY6_1(.dout(w_dff_A_BSIq8CKJ4_1),.din(w_dff_A_1LQ596uY6_1),.clk(gclk));
	jdff dff_A_74lpbGHW9_1(.dout(w_dff_A_1LQ596uY6_1),.din(w_dff_A_74lpbGHW9_1),.clk(gclk));
	jdff dff_A_lzaRgxEL0_1(.dout(w_dff_A_74lpbGHW9_1),.din(w_dff_A_lzaRgxEL0_1),.clk(gclk));
	jdff dff_A_LmwynoSP5_1(.dout(w_dff_A_lzaRgxEL0_1),.din(w_dff_A_LmwynoSP5_1),.clk(gclk));
	jdff dff_A_PARIs3hI1_1(.dout(w_dff_A_LmwynoSP5_1),.din(w_dff_A_PARIs3hI1_1),.clk(gclk));
	jdff dff_A_6CSFh7d00_1(.dout(w_dff_A_PARIs3hI1_1),.din(w_dff_A_6CSFh7d00_1),.clk(gclk));
	jdff dff_A_TOho2NGc7_2(.dout(w_G86gat_0[2]),.din(w_dff_A_TOho2NGc7_2),.clk(gclk));
	jdff dff_A_0Hj1w6ek6_2(.dout(w_dff_A_TOho2NGc7_2),.din(w_dff_A_0Hj1w6ek6_2),.clk(gclk));
	jdff dff_A_HyRLz8mU1_2(.dout(w_dff_A_0Hj1w6ek6_2),.din(w_dff_A_HyRLz8mU1_2),.clk(gclk));
	jdff dff_A_QV749GuN9_2(.dout(w_dff_A_HyRLz8mU1_2),.din(w_dff_A_QV749GuN9_2),.clk(gclk));
	jdff dff_A_wEc8Mubu0_2(.dout(w_dff_A_QV749GuN9_2),.din(w_dff_A_wEc8Mubu0_2),.clk(gclk));
	jdff dff_A_7xqCXz1e3_2(.dout(w_dff_A_wEc8Mubu0_2),.din(w_dff_A_7xqCXz1e3_2),.clk(gclk));
	jdff dff_A_KwcRjYcX8_2(.dout(w_dff_A_7xqCXz1e3_2),.din(w_dff_A_KwcRjYcX8_2),.clk(gclk));
	jdff dff_A_saQb2HaH3_1(.dout(w_n123_0[1]),.din(w_dff_A_saQb2HaH3_1),.clk(gclk));
	jdff dff_A_XvdXSowH1_1(.dout(w_dff_A_saQb2HaH3_1),.din(w_dff_A_XvdXSowH1_1),.clk(gclk));
	jdff dff_A_KKGaIIYi5_1(.dout(w_dff_A_XvdXSowH1_1),.din(w_dff_A_KKGaIIYi5_1),.clk(gclk));
	jdff dff_A_w7DTeoif4_1(.dout(w_dff_A_KKGaIIYi5_1),.din(w_dff_A_w7DTeoif4_1),.clk(gclk));
	jdff dff_A_klqXxfI94_0(.dout(w_G47gat_0[0]),.din(w_dff_A_klqXxfI94_0),.clk(gclk));
	jdff dff_A_t254wNan5_0(.dout(w_dff_A_klqXxfI94_0),.din(w_dff_A_t254wNan5_0),.clk(gclk));
	jdff dff_A_SsooMSsU0_0(.dout(w_dff_A_t254wNan5_0),.din(w_dff_A_SsooMSsU0_0),.clk(gclk));
	jdff dff_A_k4Q3J28A3_0(.dout(w_dff_A_SsooMSsU0_0),.din(w_dff_A_k4Q3J28A3_0),.clk(gclk));
	jdff dff_A_Zie9ZKbO8_0(.dout(w_dff_A_k4Q3J28A3_0),.din(w_dff_A_Zie9ZKbO8_0),.clk(gclk));
	jdff dff_A_uKQ7X8Ye8_0(.dout(w_dff_A_Zie9ZKbO8_0),.din(w_dff_A_uKQ7X8Ye8_0),.clk(gclk));
	jdff dff_A_QBSlD7Dg1_0(.dout(w_dff_A_uKQ7X8Ye8_0),.din(w_dff_A_QBSlD7Dg1_0),.clk(gclk));
	jdff dff_B_wT6b7cE44_1(.din(n117),.dout(w_dff_B_wT6b7cE44_1),.clk(gclk));
	jdff dff_B_9j3xKf2N8_1(.din(w_dff_B_wT6b7cE44_1),.dout(w_dff_B_9j3xKf2N8_1),.clk(gclk));
	jdff dff_B_z3JBK7ly4_1(.din(w_dff_B_9j3xKf2N8_1),.dout(w_dff_B_z3JBK7ly4_1),.clk(gclk));
	jdff dff_B_Prui9E6n3_1(.din(w_dff_B_z3JBK7ly4_1),.dout(w_dff_B_Prui9E6n3_1),.clk(gclk));
	jdff dff_B_m8JfDSuB2_1(.din(w_dff_B_Prui9E6n3_1),.dout(w_dff_B_m8JfDSuB2_1),.clk(gclk));
	jdff dff_A_1ux9T1S57_0(.dout(w_G60gat_0[0]),.din(w_dff_A_1ux9T1S57_0),.clk(gclk));
	jdff dff_A_qPJ96Qa95_0(.dout(w_dff_A_1ux9T1S57_0),.din(w_dff_A_qPJ96Qa95_0),.clk(gclk));
	jdff dff_A_HTvPTl7u9_0(.dout(w_dff_A_qPJ96Qa95_0),.din(w_dff_A_HTvPTl7u9_0),.clk(gclk));
	jdff dff_A_ILbgMFZF7_0(.dout(w_dff_A_HTvPTl7u9_0),.din(w_dff_A_ILbgMFZF7_0),.clk(gclk));
	jdff dff_A_bvwyD8wS4_0(.dout(w_dff_A_ILbgMFZF7_0),.din(w_dff_A_bvwyD8wS4_0),.clk(gclk));
	jdff dff_A_nc9zCKgV8_0(.dout(w_dff_A_bvwyD8wS4_0),.din(w_dff_A_nc9zCKgV8_0),.clk(gclk));
	jdff dff_A_DqS6Uenx5_0(.dout(w_dff_A_nc9zCKgV8_0),.din(w_dff_A_DqS6Uenx5_0),.clk(gclk));
	jdff dff_A_nCUDPzqM2_1(.dout(w_G60gat_0[1]),.din(w_dff_A_nCUDPzqM2_1),.clk(gclk));
	jdff dff_A_etTlYGfi6_1(.dout(w_dff_A_nCUDPzqM2_1),.din(w_dff_A_etTlYGfi6_1),.clk(gclk));
	jdff dff_A_EYMhh2NP2_1(.dout(w_dff_A_etTlYGfi6_1),.din(w_dff_A_EYMhh2NP2_1),.clk(gclk));
	jdff dff_A_2AgsyYxV7_0(.dout(w_n115_0[0]),.din(w_dff_A_2AgsyYxV7_0),.clk(gclk));
	jdff dff_A_UYDvcHSI1_0(.dout(w_dff_A_2AgsyYxV7_0),.din(w_dff_A_UYDvcHSI1_0),.clk(gclk));
	jdff dff_A_LXsqiYb71_0(.dout(w_n114_0[0]),.din(w_dff_A_LXsqiYb71_0),.clk(gclk));
	jdff dff_A_K5gZdYiz0_0(.dout(w_dff_A_LXsqiYb71_0),.din(w_dff_A_K5gZdYiz0_0),.clk(gclk));
	jdff dff_A_o1CtH3px7_0(.dout(w_G34gat_0[0]),.din(w_dff_A_o1CtH3px7_0),.clk(gclk));
	jdff dff_A_6GEmcsxw8_0(.dout(w_dff_A_o1CtH3px7_0),.din(w_dff_A_6GEmcsxw8_0),.clk(gclk));
	jdff dff_A_rPGBybKv5_0(.dout(w_dff_A_6GEmcsxw8_0),.din(w_dff_A_rPGBybKv5_0),.clk(gclk));
	jdff dff_A_wqcMWBRI4_0(.dout(w_dff_A_rPGBybKv5_0),.din(w_dff_A_wqcMWBRI4_0),.clk(gclk));
	jdff dff_A_3KiuoKLP4_0(.dout(w_dff_A_wqcMWBRI4_0),.din(w_dff_A_3KiuoKLP4_0),.clk(gclk));
	jdff dff_A_PeqWGNTD6_0(.dout(w_dff_A_3KiuoKLP4_0),.din(w_dff_A_PeqWGNTD6_0),.clk(gclk));
	jdff dff_A_F8LbHkJN7_0(.dout(w_dff_A_PeqWGNTD6_0),.din(w_dff_A_F8LbHkJN7_0),.clk(gclk));
	jdff dff_A_0HDFWRb66_2(.dout(w_G34gat_0[2]),.din(w_dff_A_0HDFWRb66_2),.clk(gclk));
	jdff dff_A_fppVYlUd0_2(.dout(w_dff_A_0HDFWRb66_2),.din(w_dff_A_fppVYlUd0_2),.clk(gclk));
	jdff dff_A_9REwY6lZ9_2(.dout(w_dff_A_fppVYlUd0_2),.din(w_dff_A_9REwY6lZ9_2),.clk(gclk));
	jdff dff_A_kShLKGpb9_2(.dout(w_dff_A_9REwY6lZ9_2),.din(w_dff_A_kShLKGpb9_2),.clk(gclk));
	jdff dff_A_7uBotQ7w8_2(.dout(w_dff_A_kShLKGpb9_2),.din(w_dff_A_7uBotQ7w8_2),.clk(gclk));
	jdff dff_A_ZMC09e0a7_2(.dout(w_dff_A_7uBotQ7w8_2),.din(w_dff_A_ZMC09e0a7_2),.clk(gclk));
	jdff dff_A_GrXrPVvO1_0(.dout(w_n109_0[0]),.din(w_dff_A_GrXrPVvO1_0),.clk(gclk));
	jdff dff_A_zXE8161e9_0(.dout(w_dff_A_GrXrPVvO1_0),.din(w_dff_A_zXE8161e9_0),.clk(gclk));
	jdff dff_A_kcZW8rLt0_0(.dout(w_dff_A_zXE8161e9_0),.din(w_dff_A_kcZW8rLt0_0),.clk(gclk));
	jdff dff_A_Zypb9wwg6_0(.dout(w_dff_A_kcZW8rLt0_0),.din(w_dff_A_Zypb9wwg6_0),.clk(gclk));
	jdff dff_A_Pm7bGHyd0_0(.dout(w_n107_0[0]),.din(w_dff_A_Pm7bGHyd0_0),.clk(gclk));
	jdff dff_A_fdhJtzY19_0(.dout(w_dff_A_Pm7bGHyd0_0),.din(w_dff_A_fdhJtzY19_0),.clk(gclk));
	jdff dff_A_oXRlq6rw9_0(.dout(w_dff_A_fdhJtzY19_0),.din(w_dff_A_oXRlq6rw9_0),.clk(gclk));
	jdff dff_A_CDO7FLDy4_0(.dout(w_dff_A_oXRlq6rw9_0),.din(w_dff_A_CDO7FLDy4_0),.clk(gclk));
	jdff dff_B_9AEKi8Wd3_2(.din(n107),.dout(w_dff_B_9AEKi8Wd3_2),.clk(gclk));
	jdff dff_B_n9yB6g0j6_2(.din(w_dff_B_9AEKi8Wd3_2),.dout(w_dff_B_n9yB6g0j6_2),.clk(gclk));
	jdff dff_B_sc1awKeY9_2(.din(w_dff_B_n9yB6g0j6_2),.dout(w_dff_B_sc1awKeY9_2),.clk(gclk));
	jdff dff_B_i7erxtH59_2(.din(w_dff_B_sc1awKeY9_2),.dout(w_dff_B_i7erxtH59_2),.clk(gclk));
	jdff dff_B_Vyv08kLF5_2(.din(w_dff_B_i7erxtH59_2),.dout(w_dff_B_Vyv08kLF5_2),.clk(gclk));
	jdff dff_A_VSbvciKf9_0(.dout(w_G73gat_0[0]),.din(w_dff_A_VSbvciKf9_0),.clk(gclk));
	jdff dff_A_FaB9VHLX3_0(.dout(w_dff_A_VSbvciKf9_0),.din(w_dff_A_FaB9VHLX3_0),.clk(gclk));
	jdff dff_A_Ygu4L3Fl5_0(.dout(w_dff_A_FaB9VHLX3_0),.din(w_dff_A_Ygu4L3Fl5_0),.clk(gclk));
	jdff dff_A_upJ1DuWE0_0(.dout(w_dff_A_Ygu4L3Fl5_0),.din(w_dff_A_upJ1DuWE0_0),.clk(gclk));
	jdff dff_A_uADjZGxX3_0(.dout(w_dff_A_upJ1DuWE0_0),.din(w_dff_A_uADjZGxX3_0),.clk(gclk));
	jdff dff_A_EkgfeO7E3_0(.dout(w_dff_A_uADjZGxX3_0),.din(w_dff_A_EkgfeO7E3_0),.clk(gclk));
	jdff dff_A_B9xrlfVz5_0(.dout(w_dff_A_EkgfeO7E3_0),.din(w_dff_A_B9xrlfVz5_0),.clk(gclk));
	jdff dff_A_nsrhvbI39_1(.dout(w_G73gat_0[1]),.din(w_dff_A_nsrhvbI39_1),.clk(gclk));
	jdff dff_A_QoTXlDAs2_1(.dout(w_dff_A_nsrhvbI39_1),.din(w_dff_A_QoTXlDAs2_1),.clk(gclk));
	jdff dff_A_R0XfIb7R3_1(.dout(w_dff_A_QoTXlDAs2_1),.din(w_dff_A_R0XfIb7R3_1),.clk(gclk));
	jdff dff_B_WrgAAFQT6_1(.din(n103),.dout(w_dff_B_WrgAAFQT6_1),.clk(gclk));
	jdff dff_B_L4gTz73F1_1(.din(w_dff_B_WrgAAFQT6_1),.dout(w_dff_B_L4gTz73F1_1),.clk(gclk));
	jdff dff_B_KmI86kS49_1(.din(w_dff_B_L4gTz73F1_1),.dout(w_dff_B_KmI86kS49_1),.clk(gclk));
	jdff dff_B_8FQ5nRby9_1(.din(w_dff_B_KmI86kS49_1),.dout(w_dff_B_8FQ5nRby9_1),.clk(gclk));
	jdff dff_B_SxfERUy20_1(.din(w_dff_B_8FQ5nRby9_1),.dout(w_dff_B_SxfERUy20_1),.clk(gclk));
	jdff dff_A_LmBsVYOJ1_0(.dout(w_G99gat_0[0]),.din(w_dff_A_LmBsVYOJ1_0),.clk(gclk));
	jdff dff_A_vdXwpCaN8_0(.dout(w_dff_A_LmBsVYOJ1_0),.din(w_dff_A_vdXwpCaN8_0),.clk(gclk));
	jdff dff_A_YjA6dPWN9_0(.dout(w_dff_A_vdXwpCaN8_0),.din(w_dff_A_YjA6dPWN9_0),.clk(gclk));
	jdff dff_A_Q7oYwNKj6_1(.dout(w_G99gat_0[1]),.din(w_dff_A_Q7oYwNKj6_1),.clk(gclk));
	jdff dff_A_nqjCgffJ3_1(.dout(w_dff_A_Q7oYwNKj6_1),.din(w_dff_A_nqjCgffJ3_1),.clk(gclk));
	jdff dff_A_ldZQdspU7_1(.dout(w_dff_A_nqjCgffJ3_1),.din(w_dff_A_ldZQdspU7_1),.clk(gclk));
	jdff dff_A_MJd0lSQh5_1(.dout(w_dff_A_ldZQdspU7_1),.din(w_dff_A_MJd0lSQh5_1),.clk(gclk));
	jdff dff_A_u5QpBoZE8_1(.dout(w_dff_A_MJd0lSQh5_1),.din(w_dff_A_u5QpBoZE8_1),.clk(gclk));
	jdff dff_A_PFOYwTxd2_1(.dout(w_dff_A_u5QpBoZE8_1),.din(w_dff_A_PFOYwTxd2_1),.clk(gclk));
	jdff dff_A_sIDebUwH7_1(.dout(w_dff_A_PFOYwTxd2_1),.din(w_dff_A_sIDebUwH7_1),.clk(gclk));
	jdff dff_A_BnZ8GJYy9_0(.dout(w_n100_0[0]),.din(w_dff_A_BnZ8GJYy9_0),.clk(gclk));
	jdff dff_A_SPrxYeus6_0(.dout(w_dff_A_BnZ8GJYy9_0),.din(w_dff_A_SPrxYeus6_0),.clk(gclk));
	jdff dff_A_tJ2kkDH47_0(.dout(w_dff_A_SPrxYeus6_0),.din(w_dff_A_tJ2kkDH47_0),.clk(gclk));
	jdff dff_A_Ka4lySTd9_0(.dout(w_dff_A_tJ2kkDH47_0),.din(w_dff_A_Ka4lySTd9_0),.clk(gclk));
	jdff dff_A_KxULQEaE2_0(.dout(w_n98_0[0]),.din(w_dff_A_KxULQEaE2_0),.clk(gclk));
	jdff dff_A_Px12xE5V5_0(.dout(w_dff_A_KxULQEaE2_0),.din(w_dff_A_Px12xE5V5_0),.clk(gclk));
	jdff dff_A_pFsUduFA4_0(.dout(w_dff_A_Px12xE5V5_0),.din(w_dff_A_pFsUduFA4_0),.clk(gclk));
	jdff dff_A_PUtd6XR36_0(.dout(w_dff_A_pFsUduFA4_0),.din(w_dff_A_PUtd6XR36_0),.clk(gclk));
	jdff dff_B_INznXfhf6_2(.din(n98),.dout(w_dff_B_INznXfhf6_2),.clk(gclk));
	jdff dff_B_MiTTpgiV0_2(.din(w_dff_B_INznXfhf6_2),.dout(w_dff_B_MiTTpgiV0_2),.clk(gclk));
	jdff dff_B_7f13l2KJ8_2(.din(w_dff_B_MiTTpgiV0_2),.dout(w_dff_B_7f13l2KJ8_2),.clk(gclk));
	jdff dff_B_2AkHVdqx1_2(.din(w_dff_B_7f13l2KJ8_2),.dout(w_dff_B_2AkHVdqx1_2),.clk(gclk));
	jdff dff_B_tHKxWh0D8_2(.din(w_dff_B_2AkHVdqx1_2),.dout(w_dff_B_tHKxWh0D8_2),.clk(gclk));
	jdff dff_A_TvXMT8YZ3_0(.dout(w_G8gat_0[0]),.din(w_dff_A_TvXMT8YZ3_0),.clk(gclk));
	jdff dff_A_zezalJ4X7_0(.dout(w_dff_A_TvXMT8YZ3_0),.din(w_dff_A_zezalJ4X7_0),.clk(gclk));
	jdff dff_A_goJCiRP38_0(.dout(w_dff_A_zezalJ4X7_0),.din(w_dff_A_goJCiRP38_0),.clk(gclk));
	jdff dff_A_Tt5DhScb6_0(.dout(w_dff_A_goJCiRP38_0),.din(w_dff_A_Tt5DhScb6_0),.clk(gclk));
	jdff dff_A_os6HbrYI5_0(.dout(w_dff_A_Tt5DhScb6_0),.din(w_dff_A_os6HbrYI5_0),.clk(gclk));
	jdff dff_A_6WhEq6Vx3_0(.dout(w_dff_A_os6HbrYI5_0),.din(w_dff_A_6WhEq6Vx3_0),.clk(gclk));
	jdff dff_A_KxQ4NtnU9_0(.dout(w_dff_A_6WhEq6Vx3_0),.din(w_dff_A_KxQ4NtnU9_0),.clk(gclk));
	jdff dff_A_WOWvNLkQ1_1(.dout(w_G8gat_0[1]),.din(w_dff_A_WOWvNLkQ1_1),.clk(gclk));
	jdff dff_A_KZWlUtOU4_1(.dout(w_dff_A_WOWvNLkQ1_1),.din(w_dff_A_KZWlUtOU4_1),.clk(gclk));
	jdff dff_A_kYYK6bRS4_1(.dout(w_dff_A_KZWlUtOU4_1),.din(w_dff_A_kYYK6bRS4_1),.clk(gclk));
	jdff dff_A_MyYSfVuL7_0(.dout(w_n96_0[0]),.din(w_dff_A_MyYSfVuL7_0),.clk(gclk));
	jdff dff_A_kqsKzx969_0(.dout(w_dff_A_MyYSfVuL7_0),.din(w_dff_A_kqsKzx969_0),.clk(gclk));
	jdff dff_A_PtH4u72W1_0(.dout(w_dff_A_kqsKzx969_0),.din(w_dff_A_PtH4u72W1_0),.clk(gclk));
	jdff dff_A_zBbLDxvQ0_0(.dout(w_dff_A_PtH4u72W1_0),.din(w_dff_A_zBbLDxvQ0_0),.clk(gclk));
	jdff dff_B_LNRer4O56_1(.din(n81),.dout(w_dff_B_LNRer4O56_1),.clk(gclk));
	jdff dff_A_bG27XOGL8_0(.dout(w_n89_0[0]),.din(w_dff_A_bG27XOGL8_0),.clk(gclk));
	jdff dff_A_v4vcAIMn0_0(.dout(w_dff_A_bG27XOGL8_0),.din(w_dff_A_v4vcAIMn0_0),.clk(gclk));
	jdff dff_A_WlB0py4B6_0(.dout(w_n84_0[0]),.din(w_dff_A_WlB0py4B6_0),.clk(gclk));
	jdff dff_A_SAaoQR5h7_0(.dout(w_dff_A_WlB0py4B6_0),.din(w_dff_A_SAaoQR5h7_0),.clk(gclk));
	jdff dff_A_fjnOabEE3_0(.dout(w_n82_0[0]),.din(w_dff_A_fjnOabEE3_0),.clk(gclk));
	jdff dff_A_4RWu16j10_0(.dout(w_dff_A_fjnOabEE3_0),.din(w_dff_A_4RWu16j10_0),.clk(gclk));
	jdff dff_A_EV2sJo6k3_0(.dout(w_n79_0[0]),.din(w_dff_A_EV2sJo6k3_0),.clk(gclk));
	jdff dff_A_gaki3A8c6_0(.dout(w_dff_A_EV2sJo6k3_0),.din(w_dff_A_gaki3A8c6_0),.clk(gclk));
	jdff dff_A_7D03RUXx3_0(.dout(w_n78_0[0]),.din(w_dff_A_7D03RUXx3_0),.clk(gclk));
	jdff dff_A_xsn42MhW1_0(.dout(w_dff_A_7D03RUXx3_0),.din(w_dff_A_xsn42MhW1_0),.clk(gclk));
	jdff dff_A_bZ6zyFUp1_0(.dout(w_dff_A_xsn42MhW1_0),.din(w_dff_A_bZ6zyFUp1_0),.clk(gclk));
	jdff dff_A_YTuRB6Gf8_0(.dout(w_dff_A_bZ6zyFUp1_0),.din(w_dff_A_YTuRB6Gf8_0),.clk(gclk));
	jdff dff_A_JUJu95Zx7_0(.dout(w_n77_0[0]),.din(w_dff_A_JUJu95Zx7_0),.clk(gclk));
	jdff dff_A_LR7YmvsM5_0(.dout(w_dff_A_JUJu95Zx7_0),.din(w_dff_A_LR7YmvsM5_0),.clk(gclk));
	jdff dff_B_A8pZF0mD5_0(.din(n75),.dout(w_dff_B_A8pZF0mD5_0),.clk(gclk));
	jdff dff_A_QNhJK7rH4_0(.dout(w_n73_0[0]),.din(w_dff_A_QNhJK7rH4_0),.clk(gclk));
	jdff dff_A_jNCouyL34_0(.dout(w_dff_A_QNhJK7rH4_0),.din(w_dff_A_jNCouyL34_0),.clk(gclk));
	jdff dff_A_H3BVJhYs1_0(.dout(w_n72_0[0]),.din(w_dff_A_H3BVJhYs1_0),.clk(gclk));
	jdff dff_A_xGrMqJsJ5_0(.dout(w_dff_A_H3BVJhYs1_0),.din(w_dff_A_xGrMqJsJ5_0),.clk(gclk));
	jdff dff_A_Xagkc7CY7_0(.dout(w_dff_A_xGrMqJsJ5_0),.din(w_dff_A_Xagkc7CY7_0),.clk(gclk));
	jdff dff_A_Ta83EDWr3_0(.dout(w_dff_A_Xagkc7CY7_0),.din(w_dff_A_Ta83EDWr3_0),.clk(gclk));
	jdff dff_A_vJO7fpZQ4_0(.dout(w_n71_0[0]),.din(w_dff_A_vJO7fpZQ4_0),.clk(gclk));
	jdff dff_A_IlkKZJFh0_0(.dout(w_dff_A_vJO7fpZQ4_0),.din(w_dff_A_IlkKZJFh0_0),.clk(gclk));
	jdff dff_A_AXMTzXvf2_0(.dout(w_dff_A_IlkKZJFh0_0),.din(w_dff_A_AXMTzXvf2_0),.clk(gclk));
	jdff dff_A_EtBe2ehS1_0(.dout(w_dff_A_AXMTzXvf2_0),.din(w_dff_A_EtBe2ehS1_0),.clk(gclk));
	jdff dff_A_AtdiSjA13_0(.dout(w_dff_A_EtBe2ehS1_0),.din(w_dff_A_AtdiSjA13_0),.clk(gclk));
	jdff dff_A_A2XPuU905_0(.dout(w_n69_0[0]),.din(w_dff_A_A2XPuU905_0),.clk(gclk));
	jdff dff_A_hSCnyLzu4_0(.dout(w_dff_A_A2XPuU905_0),.din(w_dff_A_hSCnyLzu4_0),.clk(gclk));
	jdff dff_A_JceNb8cT8_0(.dout(w_dff_A_hSCnyLzu4_0),.din(w_dff_A_JceNb8cT8_0),.clk(gclk));
	jdff dff_A_0K2V6HLY3_0(.dout(w_dff_A_JceNb8cT8_0),.din(w_dff_A_0K2V6HLY3_0),.clk(gclk));
	jdff dff_B_ctJnivF36_2(.din(n69),.dout(w_dff_B_ctJnivF36_2),.clk(gclk));
	jdff dff_B_rHP0cAYc5_2(.din(w_dff_B_ctJnivF36_2),.dout(w_dff_B_rHP0cAYc5_2),.clk(gclk));
	jdff dff_B_JCPlyy7P0_2(.din(w_dff_B_rHP0cAYc5_2),.dout(w_dff_B_JCPlyy7P0_2),.clk(gclk));
	jdff dff_B_xpLdf9kD2_2(.din(w_dff_B_JCPlyy7P0_2),.dout(w_dff_B_xpLdf9kD2_2),.clk(gclk));
	jdff dff_B_qb1tUmSa4_2(.din(w_dff_B_xpLdf9kD2_2),.dout(w_dff_B_qb1tUmSa4_2),.clk(gclk));
	jdff dff_A_ciQpGTVL6_0(.dout(w_G112gat_0[0]),.din(w_dff_A_ciQpGTVL6_0),.clk(gclk));
	jdff dff_A_9bMwNqAm2_0(.dout(w_dff_A_ciQpGTVL6_0),.din(w_dff_A_9bMwNqAm2_0),.clk(gclk));
	jdff dff_A_GK8arUIn6_0(.dout(w_dff_A_9bMwNqAm2_0),.din(w_dff_A_GK8arUIn6_0),.clk(gclk));
	jdff dff_A_VSeaxf1k8_0(.dout(w_dff_A_GK8arUIn6_0),.din(w_dff_A_VSeaxf1k8_0),.clk(gclk));
	jdff dff_A_dcHtOUie7_0(.dout(w_dff_A_VSeaxf1k8_0),.din(w_dff_A_dcHtOUie7_0),.clk(gclk));
	jdff dff_A_QVr0zDOh5_0(.dout(w_dff_A_dcHtOUie7_0),.din(w_dff_A_QVr0zDOh5_0),.clk(gclk));
	jdff dff_A_oxSmCrPp1_0(.dout(w_dff_A_QVr0zDOh5_0),.din(w_dff_A_oxSmCrPp1_0),.clk(gclk));
	jdff dff_A_EK9hzRGP0_1(.dout(w_G112gat_0[1]),.din(w_dff_A_EK9hzRGP0_1),.clk(gclk));
	jdff dff_A_WTrN4iro9_1(.dout(w_dff_A_EK9hzRGP0_1),.din(w_dff_A_WTrN4iro9_1),.clk(gclk));
	jdff dff_A_r9UuOjSk8_1(.dout(w_dff_A_WTrN4iro9_1),.din(w_dff_A_r9UuOjSk8_1),.clk(gclk));
	jdff dff_A_N7fbQPkr9_1(.dout(w_n139_0[1]),.din(w_dff_A_N7fbQPkr9_1),.clk(gclk));
	jdff dff_A_aTbF4cHM8_1(.dout(w_dff_A_N7fbQPkr9_1),.din(w_dff_A_aTbF4cHM8_1),.clk(gclk));
	jdff dff_A_FWcx9C3Y3_1(.dout(w_dff_A_aTbF4cHM8_1),.din(w_dff_A_FWcx9C3Y3_1),.clk(gclk));
	jdff dff_A_1ipRx2DE7_1(.dout(w_dff_A_FWcx9C3Y3_1),.din(w_dff_A_1ipRx2DE7_1),.clk(gclk));
	jdff dff_A_LnOkSJ5j2_1(.dout(w_dff_A_1ipRx2DE7_1),.din(w_dff_A_LnOkSJ5j2_1),.clk(gclk));
	jdff dff_A_BxmwBAfp9_0(.dout(w_G4gat_0[0]),.din(w_dff_A_BxmwBAfp9_0),.clk(gclk));
	jdff dff_A_AwL1qWK18_0(.dout(w_dff_A_BxmwBAfp9_0),.din(w_dff_A_AwL1qWK18_0),.clk(gclk));
	jdff dff_A_otO67G9I2_0(.dout(w_dff_A_AwL1qWK18_0),.din(w_dff_A_otO67G9I2_0),.clk(gclk));
	jdff dff_A_mpTh07YM3_0(.dout(w_dff_A_otO67G9I2_0),.din(w_dff_A_mpTh07YM3_0),.clk(gclk));
	jdff dff_A_QeiAwPo49_0(.dout(w_dff_A_mpTh07YM3_0),.din(w_dff_A_QeiAwPo49_0),.clk(gclk));
	jdff dff_A_ackFX2VS9_2(.dout(w_G4gat_0[2]),.din(w_dff_A_ackFX2VS9_2),.clk(gclk));
	jdff dff_A_7tHy1G102_0(.dout(w_n63_0[0]),.din(w_dff_A_7tHy1G102_0),.clk(gclk));
	jdff dff_A_qVT9keJC1_0(.dout(w_dff_A_7tHy1G102_0),.din(w_dff_A_qVT9keJC1_0),.clk(gclk));
	jdff dff_A_yODH62IO5_0(.dout(w_dff_A_qVT9keJC1_0),.din(w_dff_A_yODH62IO5_0),.clk(gclk));
	jdff dff_A_cXNwIErP0_0(.dout(w_dff_A_yODH62IO5_0),.din(w_dff_A_cXNwIErP0_0),.clk(gclk));
	jdff dff_A_3nvwjmDD0_0(.dout(w_G1gat_0[0]),.din(w_dff_A_3nvwjmDD0_0),.clk(gclk));
	jdff dff_A_8Q9aDmsZ4_0(.dout(w_dff_A_3nvwjmDD0_0),.din(w_dff_A_8Q9aDmsZ4_0),.clk(gclk));
	jdff dff_A_S9cH5ASg8_1(.dout(w_G1gat_0[1]),.din(w_dff_A_S9cH5ASg8_1),.clk(gclk));
	jdff dff_A_APOtbspc7_0(.dout(w_n61_0[0]),.din(w_dff_A_APOtbspc7_0),.clk(gclk));
	jdff dff_A_f3Xi4Qwd0_0(.dout(w_dff_A_APOtbspc7_0),.din(w_dff_A_f3Xi4Qwd0_0),.clk(gclk));
	jdff dff_A_aVFwHXl16_0(.dout(w_dff_A_f3Xi4Qwd0_0),.din(w_dff_A_aVFwHXl16_0),.clk(gclk));
	jdff dff_A_Gis9XQrO3_0(.dout(w_dff_A_aVFwHXl16_0),.din(w_dff_A_Gis9XQrO3_0),.clk(gclk));
	jdff dff_A_v7VY6Ps68_0(.dout(w_G89gat_0[0]),.din(w_dff_A_v7VY6Ps68_0),.clk(gclk));
	jdff dff_A_mK9E1x6N7_0(.dout(w_dff_A_v7VY6Ps68_0),.din(w_dff_A_mK9E1x6N7_0),.clk(gclk));
	jdff dff_A_spUQlFXn1_1(.dout(w_G89gat_0[1]),.din(w_dff_A_spUQlFXn1_1),.clk(gclk));
	jdff dff_A_EHE0HbeY6_0(.dout(w_G56gat_0[0]),.din(w_dff_A_EHE0HbeY6_0),.clk(gclk));
	jdff dff_A_ykbCGbil4_0(.dout(w_dff_A_EHE0HbeY6_0),.din(w_dff_A_ykbCGbil4_0),.clk(gclk));
	jdff dff_A_HcPEVzBh4_0(.dout(w_dff_A_ykbCGbil4_0),.din(w_dff_A_HcPEVzBh4_0),.clk(gclk));
	jdff dff_A_qQqlwDc46_0(.dout(w_dff_A_HcPEVzBh4_0),.din(w_dff_A_qQqlwDc46_0),.clk(gclk));
	jdff dff_A_ykuSPxPC3_0(.dout(w_dff_A_qQqlwDc46_0),.din(w_dff_A_ykuSPxPC3_0),.clk(gclk));
	jdff dff_A_yhPEyTC79_2(.dout(w_G56gat_0[2]),.din(w_dff_A_yhPEyTC79_2),.clk(gclk));
	jdff dff_A_S9UKB6UZ7_0(.dout(w_n58_0[0]),.din(w_dff_A_S9UKB6UZ7_0),.clk(gclk));
	jdff dff_A_Ve4z2LmU5_0(.dout(w_dff_A_S9UKB6UZ7_0),.din(w_dff_A_Ve4z2LmU5_0),.clk(gclk));
	jdff dff_A_VTN8bKRk0_0(.dout(w_dff_A_Ve4z2LmU5_0),.din(w_dff_A_VTN8bKRk0_0),.clk(gclk));
	jdff dff_A_Gos5lcXw0_0(.dout(w_dff_A_VTN8bKRk0_0),.din(w_dff_A_Gos5lcXw0_0),.clk(gclk));
	jdff dff_A_qQ3Kzdjq6_0(.dout(w_G50gat_0[0]),.din(w_dff_A_qQ3Kzdjq6_0),.clk(gclk));
	jdff dff_A_fFAyDfkg4_0(.dout(w_dff_A_qQ3Kzdjq6_0),.din(w_dff_A_fFAyDfkg4_0),.clk(gclk));
	jdff dff_A_ccVj2SPm1_1(.dout(w_G50gat_0[1]),.din(w_dff_A_ccVj2SPm1_1),.clk(gclk));
	jdff dff_A_gr0LHtEM7_0(.dout(w_G108gat_0[0]),.din(w_dff_A_gr0LHtEM7_0),.clk(gclk));
	jdff dff_A_jlg59BuU9_0(.dout(w_dff_A_gr0LHtEM7_0),.din(w_dff_A_jlg59BuU9_0),.clk(gclk));
	jdff dff_A_AV8qV57X8_0(.dout(w_dff_A_jlg59BuU9_0),.din(w_dff_A_AV8qV57X8_0),.clk(gclk));
	jdff dff_A_iS2sVosO3_0(.dout(w_dff_A_AV8qV57X8_0),.din(w_dff_A_iS2sVosO3_0),.clk(gclk));
	jdff dff_A_EIPkYlR64_0(.dout(w_dff_A_iS2sVosO3_0),.din(w_dff_A_EIPkYlR64_0),.clk(gclk));
	jdff dff_A_x97kb6s77_2(.dout(w_G108gat_0[2]),.din(w_dff_A_x97kb6s77_2),.clk(gclk));
	jdff dff_A_HH5XMtOD5_0(.dout(w_n56_0[0]),.din(w_dff_A_HH5XMtOD5_0),.clk(gclk));
	jdff dff_A_mt9U9CVX7_0(.dout(w_dff_A_HH5XMtOD5_0),.din(w_dff_A_mt9U9CVX7_0),.clk(gclk));
	jdff dff_A_cxvNp9Vi8_0(.dout(w_dff_A_mt9U9CVX7_0),.din(w_dff_A_cxvNp9Vi8_0),.clk(gclk));
	jdff dff_A_yHbq8kSS5_0(.dout(w_dff_A_cxvNp9Vi8_0),.din(w_dff_A_yHbq8kSS5_0),.clk(gclk));
	jdff dff_A_ZHctAwEN9_0(.dout(w_G102gat_0[0]),.din(w_dff_A_ZHctAwEN9_0),.clk(gclk));
	jdff dff_A_iwJkMMKv3_0(.dout(w_dff_A_ZHctAwEN9_0),.din(w_dff_A_iwJkMMKv3_0),.clk(gclk));
	jdff dff_A_bZE7w3OJ6_1(.dout(w_G102gat_0[1]),.din(w_dff_A_bZE7w3OJ6_1),.clk(gclk));
	jdff dff_A_KWD4Dwzu7_0(.dout(w_G69gat_0[0]),.din(w_dff_A_KWD4Dwzu7_0),.clk(gclk));
	jdff dff_A_6iCdptVu6_0(.dout(w_dff_A_KWD4Dwzu7_0),.din(w_dff_A_6iCdptVu6_0),.clk(gclk));
	jdff dff_A_2Ov9wwNx0_0(.dout(w_dff_A_6iCdptVu6_0),.din(w_dff_A_2Ov9wwNx0_0),.clk(gclk));
	jdff dff_A_3WsiLQ5r3_0(.dout(w_dff_A_2Ov9wwNx0_0),.din(w_dff_A_3WsiLQ5r3_0),.clk(gclk));
	jdff dff_A_cSh138lx0_0(.dout(w_dff_A_3WsiLQ5r3_0),.din(w_dff_A_cSh138lx0_0),.clk(gclk));
	jdff dff_A_mNTfqqc63_2(.dout(w_G69gat_0[2]),.din(w_dff_A_mNTfqqc63_2),.clk(gclk));
	jdff dff_A_I73cHgpi9_0(.dout(w_n53_0[0]),.din(w_dff_A_I73cHgpi9_0),.clk(gclk));
	jdff dff_A_fHB4XJih3_0(.dout(w_dff_A_I73cHgpi9_0),.din(w_dff_A_fHB4XJih3_0),.clk(gclk));
	jdff dff_A_KbVKz9Mn1_0(.dout(w_dff_A_fHB4XJih3_0),.din(w_dff_A_KbVKz9Mn1_0),.clk(gclk));
	jdff dff_A_EuZn7Eiy6_0(.dout(w_dff_A_KbVKz9Mn1_0),.din(w_dff_A_EuZn7Eiy6_0),.clk(gclk));
	jdff dff_A_8WY9Fg2k9_0(.dout(w_G63gat_0[0]),.din(w_dff_A_8WY9Fg2k9_0),.clk(gclk));
	jdff dff_A_hJhMiXj88_0(.dout(w_dff_A_8WY9Fg2k9_0),.din(w_dff_A_hJhMiXj88_0),.clk(gclk));
	jdff dff_A_kRPglyTL6_1(.dout(w_G63gat_0[1]),.din(w_dff_A_kRPglyTL6_1),.clk(gclk));
	jdff dff_A_WyQy5OLV6_0(.dout(w_n52_0[0]),.din(w_dff_A_WyQy5OLV6_0),.clk(gclk));
	jdff dff_A_7ewoJsAz5_0(.dout(w_dff_A_WyQy5OLV6_0),.din(w_dff_A_7ewoJsAz5_0),.clk(gclk));
	jdff dff_A_pv6JlPPU4_0(.dout(w_dff_A_7ewoJsAz5_0),.din(w_dff_A_pv6JlPPU4_0),.clk(gclk));
	jdff dff_A_bjbEQ63G7_1(.dout(w_G43gat_1[1]),.din(w_dff_A_bjbEQ63G7_1),.clk(gclk));
	jdff dff_A_4XfPiDUQ5_1(.dout(w_G43gat_0[1]),.din(w_dff_A_4XfPiDUQ5_1),.clk(gclk));
	jdff dff_A_KwYcxXwP8_2(.dout(w_G43gat_0[2]),.din(w_dff_A_KwYcxXwP8_2),.clk(gclk));
	jdff dff_A_UyYShGjK6_0(.dout(w_G37gat_0[0]),.din(w_dff_A_UyYShGjK6_0),.clk(gclk));
	jdff dff_A_pq1DDwcH6_0(.dout(w_dff_A_UyYShGjK6_0),.din(w_dff_A_pq1DDwcH6_0),.clk(gclk));
	jdff dff_A_Q2VAeA2m4_1(.dout(w_G37gat_0[1]),.din(w_dff_A_Q2VAeA2m4_1),.clk(gclk));
	jdff dff_A_XMo7uwTd9_0(.dout(w_G17gat_0[0]),.din(w_dff_A_XMo7uwTd9_0),.clk(gclk));
	jdff dff_A_AsJ4Gvp40_0(.dout(w_dff_A_XMo7uwTd9_0),.din(w_dff_A_AsJ4Gvp40_0),.clk(gclk));
	jdff dff_A_p1w3Gei79_0(.dout(w_dff_A_AsJ4Gvp40_0),.din(w_dff_A_p1w3Gei79_0),.clk(gclk));
	jdff dff_A_syGEktSd7_0(.dout(w_dff_A_p1w3Gei79_0),.din(w_dff_A_syGEktSd7_0),.clk(gclk));
	jdff dff_A_tQeqhSFR8_0(.dout(w_dff_A_syGEktSd7_0),.din(w_dff_A_tQeqhSFR8_0),.clk(gclk));
	jdff dff_A_RuHE0NNv0_2(.dout(w_G17gat_0[2]),.din(w_dff_A_RuHE0NNv0_2),.clk(gclk));
	jdff dff_A_xc9obCm23_0(.dout(w_n47_0[0]),.din(w_dff_A_xc9obCm23_0),.clk(gclk));
	jdff dff_A_813ZqyV73_0(.dout(w_dff_A_xc9obCm23_0),.din(w_dff_A_813ZqyV73_0),.clk(gclk));
	jdff dff_A_j4wWfytA0_0(.dout(w_dff_A_813ZqyV73_0),.din(w_dff_A_j4wWfytA0_0),.clk(gclk));
	jdff dff_A_9GXswcgi6_0(.dout(w_dff_A_j4wWfytA0_0),.din(w_dff_A_9GXswcgi6_0),.clk(gclk));
	jdff dff_A_0Vl9meXi0_0(.dout(w_G11gat_0[0]),.din(w_dff_A_0Vl9meXi0_0),.clk(gclk));
	jdff dff_A_Ds2KCWjB4_0(.dout(w_dff_A_0Vl9meXi0_0),.din(w_dff_A_Ds2KCWjB4_0),.clk(gclk));
	jdff dff_A_zx77paec5_1(.dout(w_G11gat_0[1]),.din(w_dff_A_zx77paec5_1),.clk(gclk));
	jdff dff_A_4SCBLVVK6_1(.dout(w_G30gat_0[1]),.din(w_dff_A_4SCBLVVK6_1),.clk(gclk));
	jdff dff_A_tH6gJrwO5_0(.dout(w_G24gat_0[0]),.din(w_dff_A_tH6gJrwO5_0),.clk(gclk));
	jdff dff_A_fgwqndJK0_1(.dout(w_G82gat_0[1]),.din(w_dff_A_fgwqndJK0_1),.clk(gclk));
	jdff dff_A_S0Zpzih35_1(.dout(w_dff_A_fgwqndJK0_1),.din(w_dff_A_S0Zpzih35_1),.clk(gclk));
	jdff dff_A_NTnB0OF15_1(.dout(w_dff_A_S0Zpzih35_1),.din(w_dff_A_NTnB0OF15_1),.clk(gclk));
	jdff dff_A_Nj3ox54D2_1(.dout(w_dff_A_NTnB0OF15_1),.din(w_dff_A_Nj3ox54D2_1),.clk(gclk));
	jdff dff_A_68cmWWIi9_1(.dout(w_dff_A_Nj3ox54D2_1),.din(w_dff_A_68cmWWIi9_1),.clk(gclk));
	jdff dff_A_xeQ0w4hR0_2(.dout(w_G82gat_0[2]),.din(w_dff_A_xeQ0w4hR0_2),.clk(gclk));
	jdff dff_A_jXWkyhs01_0(.dout(w_n43_0[0]),.din(w_dff_A_jXWkyhs01_0),.clk(gclk));
	jdff dff_A_SPilwwnD3_0(.dout(w_dff_A_jXWkyhs01_0),.din(w_dff_A_SPilwwnD3_0),.clk(gclk));
	jdff dff_A_u7R7yUNg8_0(.dout(w_dff_A_SPilwwnD3_0),.din(w_dff_A_u7R7yUNg8_0),.clk(gclk));
	jdff dff_A_PDTzFAbJ0_0(.dout(w_dff_A_u7R7yUNg8_0),.din(w_dff_A_PDTzFAbJ0_0),.clk(gclk));
	jdff dff_A_KKzrVnWZ8_0(.dout(w_G76gat_0[0]),.din(w_dff_A_KKzrVnWZ8_0),.clk(gclk));
	jdff dff_A_V77Qgtx09_0(.dout(w_dff_A_KKzrVnWZ8_0),.din(w_dff_A_V77Qgtx09_0),.clk(gclk));
	jdff dff_A_1TIcpTGE4_0(.dout(w_n87_0[0]),.din(w_dff_A_1TIcpTGE4_0),.clk(gclk));
	jdff dff_A_ofGCrke68_0(.dout(w_dff_A_1TIcpTGE4_0),.din(w_dff_A_ofGCrke68_0),.clk(gclk));
	jdff dff_A_cs9ejUyk0_0(.dout(w_G95gat_0[0]),.din(w_dff_A_cs9ejUyk0_0),.clk(gclk));
	jdff dff_A_mGFoBZuA1_0(.dout(w_dff_A_cs9ejUyk0_0),.din(w_dff_A_mGFoBZuA1_0),.clk(gclk));
	jdff dff_A_eO7y5zfd3_0(.dout(w_dff_A_mGFoBZuA1_0),.din(w_dff_A_eO7y5zfd3_0),.clk(gclk));
	jdff dff_A_nJ8mA2cN9_0(.dout(w_dff_A_eO7y5zfd3_0),.din(w_dff_A_nJ8mA2cN9_0),.clk(gclk));
	jdff dff_A_UAZ4UGCm2_0(.dout(w_dff_A_nJ8mA2cN9_0),.din(w_dff_A_UAZ4UGCm2_0),.clk(gclk));
	jdff dff_A_dZ1WiuOi5_2(.dout(w_G95gat_0[2]),.din(w_dff_A_dZ1WiuOi5_2),.clk(gclk));
	jdff dff_A_BZGd1Zbo3_1(.dout(w_G105gat_0[1]),.din(w_dff_A_BZGd1Zbo3_1),.clk(gclk));
	jdff dff_A_2lFAT6Du2_1(.dout(w_dff_A_BZGd1Zbo3_1),.din(w_dff_A_2lFAT6Du2_1),.clk(gclk));
	jdff dff_A_HcHjp5KW6_1(.dout(w_dff_A_2lFAT6Du2_1),.din(w_dff_A_HcHjp5KW6_1),.clk(gclk));
	jdff dff_A_kLajnnKD6_1(.dout(w_dff_A_HcHjp5KW6_1),.din(w_dff_A_kLajnnKD6_1),.clk(gclk));
	jdff dff_A_DMqNZfW33_1(.dout(w_dff_A_kLajnnKD6_1),.din(w_dff_A_DMqNZfW33_1),.clk(gclk));
	jdff dff_A_HVDqM4J37_1(.dout(w_dff_A_DMqNZfW33_1),.din(w_dff_A_HVDqM4J37_1),.clk(gclk));
	jdff dff_A_ITHjWEV05_1(.dout(w_dff_A_HVDqM4J37_1),.din(w_dff_A_ITHjWEV05_1),.clk(gclk));
	jdff dff_A_ByEd35Mx2_1(.dout(w_dff_A_ITHjWEV05_1),.din(w_dff_A_ByEd35Mx2_1),.clk(gclk));
endmodule

