/*
gf_c432:
	jxor: 1
	jspl: 84
	jspl3: 48
	jnot: 47
	jdff: 1154
	jand: 104
	jor: 104

Summary:
	jxor: 1
	jspl: 84
	jspl3: 48
	jnot: 47
	jdff: 1154
	jand: 104
	jor: 104

The maximum logic level gap of any gate:
	gf_c432: 7
*/

module gf_c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n43;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G4gat_0;
	wire [2:0] w_G8gat_0;
	wire [2:0] w_G11gat_0;
	wire [2:0] w_G14gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G21gat_0;
	wire [2:0] w_G24gat_0;
	wire [1:0] w_G27gat_0;
	wire [2:0] w_G30gat_0;
	wire [2:0] w_G34gat_0;
	wire [1:0] w_G40gat_0;
	wire [1:0] w_G43gat_0;
	wire [2:0] w_G47gat_0;
	wire [1:0] w_G50gat_0;
	wire [1:0] w_G53gat_0;
	wire [2:0] w_G56gat_0;
	wire [1:0] w_G56gat_1;
	wire [1:0] w_G60gat_0;
	wire [2:0] w_G63gat_0;
	wire [2:0] w_G66gat_0;
	wire [2:0] w_G69gat_0;
	wire [2:0] w_G73gat_0;
	wire [2:0] w_G76gat_0;
	wire [1:0] w_G79gat_0;
	wire [2:0] w_G82gat_0;
	wire [2:0] w_G86gat_0;
	wire [2:0] w_G89gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G95gat_0;
	wire [2:0] w_G99gat_0;
	wire [1:0] w_G102gat_0;
	wire [1:0] w_G105gat_0;
	wire [2:0] w_G108gat_0;
	wire [2:0] w_G112gat_0;
	wire [1:0] w_G115gat_0;
	wire [2:0] w_G223gat_0;
	wire [2:0] w_G223gat_1;
	wire [2:0] w_G223gat_2;
	wire [2:0] w_G223gat_3;
	wire w_G223gat_4;
	wire G223gat_fa_;
	wire [2:0] w_G329gat_0;
	wire [2:0] w_G329gat_1;
	wire [2:0] w_G329gat_2;
	wire [2:0] w_G329gat_3;
	wire w_G329gat_4;
	wire G329gat_fa_;
	wire [2:0] w_G370gat_0;
	wire [1:0] w_G370gat_1;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire [1:0] w_n43_0;
	wire [1:0] w_n44_0;
	wire [1:0] w_n45_0;
	wire [2:0] w_n46_0;
	wire [1:0] w_n47_0;
	wire [1:0] w_n49_0;
	wire [1:0] w_n51_0;
	wire [1:0] w_n54_0;
	wire [1:0] w_n57_0;
	wire [1:0] w_n60_0;
	wire [1:0] w_n62_0;
	wire [1:0] w_n64_0;
	wire [1:0] w_n70_0;
	wire [1:0] w_n73_0;
	wire [1:0] w_n75_0;
	wire [1:0] w_n78_0;
	wire [1:0] w_n80_0;
	wire [1:0] w_n81_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n86_0;
	wire [1:0] w_n88_0;
	wire [2:0] w_n93_0;
	wire [2:0] w_n93_1;
	wire [2:0] w_n93_2;
	wire [2:0] w_n93_3;
	wire [1:0] w_n95_0;
	wire [1:0] w_n102_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n106_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n111_0;
	wire [1:0] w_n113_0;
	wire [1:0] w_n117_0;
	wire [2:0] w_n119_0;
	wire [1:0] w_n120_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n123_0;
	wire [1:0] w_n125_0;
	wire [1:0] w_n127_0;
	wire [2:0] w_n131_0;
	wire [1:0] w_n138_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n141_0;
	wire [1:0] w_n144_0;
	wire [1:0] w_n145_0;
	wire [1:0] w_n147_0;
	wire [1:0] w_n149_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n156_0;
	wire [1:0] w_n159_0;
	wire [1:0] w_n164_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n173_0;
	wire [2:0] w_n181_0;
	wire [2:0] w_n181_1;
	wire [2:0] w_n181_2;
	wire [1:0] w_n183_0;
	wire [1:0] w_n185_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n202_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n206_0;
	wire [1:0] w_n209_0;
	wire [1:0] w_n211_0;
	wire [1:0] w_n222_0;
	wire [1:0] w_n227_0;
	wire [1:0] w_n230_0;
	wire [2:0] w_n246_0;
	wire [2:0] w_n246_1;
	wire [2:0] w_n246_2;
	wire [1:0] w_n248_0;
	wire [1:0] w_n250_0;
	wire [1:0] w_n251_0;
	wire [1:0] w_n253_0;
	wire [1:0] w_n254_0;
	wire [1:0] w_n257_0;
	wire [1:0] w_n264_0;
	wire [1:0] w_n265_0;
	wire [1:0] w_n269_0;
	wire [1:0] w_n271_0;
	wire [1:0] w_n281_0;
	wire [1:0] w_n288_0;
	wire [1:0] w_n290_0;
	wire w_dff_B_vwebLdyM5_0;
	wire w_dff_B_oLBFTUv28_0;
	wire w_dff_B_SoG1fvF07_0;
	wire w_dff_B_79cmHCEP3_0;
	wire w_dff_B_wCIJXmYt4_0;
	wire w_dff_B_qxQuhH704_0;
	wire w_dff_B_gUf4KBF24_0;
	wire w_dff_B_3oNaz6UP6_0;
	wire w_dff_B_8uzFWmwk8_0;
	wire w_dff_B_r4O0bDM98_2;
	wire w_dff_A_ePfqqCRY9_0;
	wire w_dff_B_RfiQmJcF3_2;
	wire w_dff_A_V53s9Bud7_1;
	wire w_dff_B_43yBtcuU3_1;
	wire w_dff_B_KVHQTPUU2_1;
	wire w_dff_B_tOvj13OK4_1;
	wire w_dff_B_qrDAUZOZ2_1;
	wire w_dff_B_FgqCtSzS2_1;
	wire w_dff_B_KOSLGNRT6_1;
	wire w_dff_B_LmmiM9Xv9_1;
	wire w_dff_B_LfGHjFt56_1;
	wire w_dff_B_CPy1CaQU2_1;
	wire w_dff_B_25uQAo1M0_1;
	wire w_dff_B_hSBrOcX19_1;
	wire w_dff_B_E0fz8Fo44_1;
	wire w_dff_B_cMRFAcil9_1;
	wire w_dff_B_WnVUmdgl8_1;
	wire w_dff_B_wwQQdLiQ3_1;
	wire w_dff_B_yN1SrVII7_1;
	wire w_dff_B_O01IHSQm2_1;
	wire w_dff_B_szApWXCv5_1;
	wire w_dff_B_pOZNkinj4_1;
	wire w_dff_B_zQrb1Bal0_1;
	wire w_dff_B_ODz5wPXy6_1;
	wire w_dff_B_4KOH86ug3_1;
	wire w_dff_B_CN6R47Uy5_1;
	wire w_dff_B_HKO3SEqS9_1;
	wire w_dff_B_uui4NYYm0_2;
	wire w_dff_A_XDeI3lnr5_0;
	wire w_dff_A_e9DjkIqI4_0;
	wire w_dff_A_svtpdesh5_0;
	wire w_dff_B_eJEne66E0_1;
	wire w_dff_A_GZGs2fVn7_0;
	wire w_dff_A_6UT3alEb7_0;
	wire w_dff_A_ssRhug4y7_0;
	wire w_dff_A_2GaXWSBg2_0;
	wire w_dff_A_cVOe3GPp0_0;
	wire w_dff_A_cQsYk8by8_0;
	wire w_dff_B_d4byrfUW0_1;
	wire w_dff_B_38Cgd16t7_1;
	wire w_dff_B_JDh6NcOG2_1;
	wire w_dff_B_PCjPAHOB3_1;
	wire w_dff_B_PLk0RNOm6_1;
	wire w_dff_B_6Urc5rC95_1;
	wire w_dff_B_3iyEOD4r6_1;
	wire w_dff_B_E92dO7Rk5_0;
	wire w_dff_B_iO0msDPq8_0;
	wire w_dff_B_vuu4jUCe9_0;
	wire w_dff_B_iwDUkmAt4_0;
	wire w_dff_A_bwA1ag0Z4_1;
	wire w_dff_A_KlHbBqMD0_1;
	wire w_dff_A_OITiqYk01_1;
	wire w_dff_A_75VzJehO6_1;
	wire w_dff_A_e9JMKHNp3_1;
	wire w_dff_B_K8XvReoO8_1;
	wire w_dff_B_esJ086AR6_0;
	wire w_dff_A_IOZJOknJ8_0;
	wire w_dff_A_8aKTlphy4_0;
	wire w_dff_A_3fXteCz35_0;
	wire w_dff_A_DR3j0Nzw8_0;
	wire w_dff_A_ZNZawBni9_0;
	wire w_dff_A_MtDsypUi6_0;
	wire w_dff_A_ISmlcl4W5_0;
	wire w_dff_A_QEWSt3uY8_0;
	wire w_dff_A_emJaql312_0;
	wire w_dff_A_tpC5tqD67_0;
	wire w_dff_A_qGfc80q32_0;
	wire w_dff_B_7WqDrcLp1_2;
	wire w_dff_B_9ID2y5OB1_2;
	wire w_dff_B_yfSETw2Y7_2;
	wire w_dff_B_z9yi05R28_2;
	wire w_dff_B_fFJEMfJy2_2;
	wire w_dff_B_Ri7WhaH01_2;
	wire w_dff_B_RGAJpQ5v8_2;
	wire w_dff_B_PJRQGn585_2;
	wire w_dff_B_88KCtT4B9_2;
	wire w_dff_B_KXRq1A8e9_2;
	wire w_dff_B_w7y06zHV5_2;
	wire w_dff_B_BsuvV6W49_2;
	wire w_dff_B_ks6N9hNk0_2;
	wire w_dff_B_bgzYbinz7_2;
	wire w_dff_A_olLEk2cE6_0;
	wire w_dff_A_UbvmZKng4_0;
	wire w_dff_A_VRvNWvrO0_0;
	wire w_dff_A_4fTmYll73_0;
	wire w_dff_A_OWTt24nJ5_0;
	wire w_dff_A_dbQqSDnz1_0;
	wire w_dff_A_RhOqGTS71_0;
	wire w_dff_A_Q5X4imaJ6_0;
	wire w_dff_A_kavg2DEy0_0;
	wire w_dff_A_0searHjC4_0;
	wire w_dff_A_seRwWBH32_0;
	wire w_dff_B_ZgxHQ6Hk4_2;
	wire w_dff_B_bzAcanZg5_2;
	wire w_dff_B_PA8Pnz9I4_2;
	wire w_dff_B_OGPoxPg14_2;
	wire w_dff_B_t73EmK7g8_2;
	wire w_dff_B_eg2rpMol3_2;
	wire w_dff_B_RYjBlcNS3_2;
	wire w_dff_B_0GnCNoDc7_2;
	wire w_dff_B_xvkXV2VS7_2;
	wire w_dff_B_nFb1iLfC0_2;
	wire w_dff_B_JKd3r0gC1_2;
	wire w_dff_B_17S53n1d3_2;
	wire w_dff_B_IwNFJkjs7_2;
	wire w_dff_B_JHCPCgkZ6_2;
	wire w_dff_B_GDaQqjpP7_1;
	wire w_dff_B_f2VOUnh55_1;
	wire w_dff_B_LUQePqha0_1;
	wire w_dff_B_SAF5a7wU9_1;
	wire w_dff_B_yKHAQ7bZ8_1;
	wire w_dff_B_X07PlIy63_1;
	wire w_dff_B_m65lksJo0_1;
	wire w_dff_B_0erNJKzh6_1;
	wire w_dff_B_iZMOoaEc6_1;
	wire w_dff_B_R9RicJHW6_1;
	wire w_dff_B_aDb6Ttog1_1;
	wire w_dff_B_m0F1ncWq9_1;
	wire w_dff_B_bw5EIPSK4_1;
	wire w_dff_B_XRoBwbH59_1;
	wire w_dff_B_bwo9Ndcl8_1;
	wire w_dff_B_O2ProZuN1_1;
	wire w_dff_B_tDQLSqeZ0_1;
	wire w_dff_B_rnxsM0XU5_1;
	wire w_dff_B_hikrsU7Z5_1;
	wire w_dff_B_8IOPiCWU6_1;
	wire w_dff_B_4MbmWuke4_1;
	wire w_dff_B_KTg1yAft1_1;
	wire w_dff_B_XEkyDelF6_1;
	wire w_dff_B_9z3QR0bs6_1;
	wire w_dff_B_AftZ3Wo78_1;
	wire w_dff_B_7nSYDCnB8_1;
	wire w_dff_B_GotyeNsY1_1;
	wire w_dff_B_PlDjCZY22_1;
	wire w_dff_A_PiFD3WSk3_0;
	wire w_dff_A_OMLjdNpq0_0;
	wire w_dff_A_eBwg2Bxj9_0;
	wire w_dff_A_TLy8opGb5_0;
	wire w_dff_A_zvdmaR5U2_0;
	wire w_dff_B_QQbq5IlY3_2;
	wire w_dff_B_OZd97weI4_2;
	wire w_dff_B_P5IQ1JFW2_2;
	wire w_dff_B_iunqsuTI3_2;
	wire w_dff_B_gtk4BpM27_2;
	wire w_dff_B_AOsJNhcZ1_2;
	wire w_dff_B_pzAcnuhG5_2;
	wire w_dff_B_Dbx0aZZD7_2;
	wire w_dff_B_MnC1J1qK4_2;
	wire w_dff_B_dcRO4kWi7_2;
	wire w_dff_B_cjtuyWXx7_2;
	wire w_dff_B_iyYNJnsV9_2;
	wire w_dff_B_1JorpXEE6_2;
	wire w_dff_B_y54Z7sHy7_2;
	wire w_dff_B_oiWBOB7h9_2;
	wire w_dff_A_DgN3MSVq3_0;
	wire w_dff_A_82TKdms76_0;
	wire w_dff_A_3SzNbMJf1_0;
	wire w_dff_A_jeePaV4h6_0;
	wire w_dff_A_xnsN78VT8_0;
	wire w_dff_B_GIyhLYus5_2;
	wire w_dff_B_PwQ2kG6V7_2;
	wire w_dff_B_ZbC8dhtR8_2;
	wire w_dff_B_2SXjRmGM2_2;
	wire w_dff_B_LvX2UqvK5_2;
	wire w_dff_B_BKDMNEAh6_2;
	wire w_dff_B_O2oHx9JX0_2;
	wire w_dff_B_3IVECn2B0_2;
	wire w_dff_B_B5gS4YMs9_2;
	wire w_dff_B_Laq60N2c5_2;
	wire w_dff_B_TO6m9H4P8_2;
	wire w_dff_B_R8eM2w5n0_2;
	wire w_dff_B_cEebf5uW0_2;
	wire w_dff_B_jl8Wcy995_2;
	wire w_dff_A_RM1anhUw6_0;
	wire w_dff_A_sKthbOZ28_0;
	wire w_dff_A_ZcZgjok87_0;
	wire w_dff_A_D2pY2psu8_0;
	wire w_dff_A_fMuf9xEt9_0;
	wire w_dff_A_8Dmcj8nY2_0;
	wire w_dff_A_UtKslg8F9_0;
	wire w_dff_A_1hTnlo0v1_0;
	wire w_dff_A_frZW8Ixb0_0;
	wire w_dff_B_ZhxoKhHD8_1;
	wire w_dff_B_zJt6HAym3_0;
	wire w_dff_A_WPTe1u9q5_0;
	wire w_dff_A_GSNYGnTk2_0;
	wire w_dff_A_kqEjlvSJ1_0;
	wire w_dff_A_VCL4iba75_0;
	wire w_dff_A_1w8blDM99_0;
	wire w_dff_A_qWk2rJrB6_0;
	wire w_dff_A_DzX34acp6_0;
	wire w_dff_A_aCCqTrBc7_0;
	wire w_dff_A_SWPagyCX3_0;
	wire w_dff_A_QTPwGdp08_0;
	wire w_dff_A_Rq4e2tBh2_0;
	wire w_dff_A_NxpvU0VK7_0;
	wire w_dff_A_wgEUhDkE2_0;
	wire w_dff_A_arkkcmbz7_0;
	wire w_dff_A_mAgQsyME8_0;
	wire w_dff_A_kNAQRqxn5_0;
	wire w_dff_A_vY8QnSd14_0;
	wire w_dff_A_zzuNB8Ds1_0;
	wire w_dff_A_FAluccEs6_0;
	wire w_dff_A_1gshwirA9_0;
	wire w_dff_A_dxkrPtun8_0;
	wire w_dff_A_u6BXhCcu8_0;
	wire w_dff_A_bsEdBsHB3_0;
	wire w_dff_A_UOSQooNn3_0;
	wire w_dff_A_1B5QYVXI4_0;
	wire w_dff_A_XJLVieiL0_0;
	wire w_dff_A_jFB0XQEE4_0;
	wire w_dff_A_UP0ZRpiA9_0;
	wire w_dff_A_iuNc7Xhb9_0;
	wire w_dff_A_HRDrLIPA2_0;
	wire w_dff_A_yzk0Ipx60_0;
	wire w_dff_A_RAmVZyC48_0;
	wire w_dff_A_n93NZ9wV0_0;
	wire w_dff_A_ITq3EleO6_0;
	wire w_dff_A_mCrN3Lj91_0;
	wire w_dff_A_4hKeouNQ8_0;
	wire w_dff_A_CQcrHCBb6_0;
	wire w_dff_A_C1l3zL6B5_0;
	wire w_dff_A_YD7hr8tY0_0;
	wire w_dff_A_i0KCF6q20_0;
	wire w_dff_A_4dtMxGzU6_0;
	wire w_dff_A_z1qq2N689_0;
	wire w_dff_A_cDTPGoMq9_0;
	wire w_dff_A_ieM7F0Qu8_0;
	wire w_dff_A_z9Dm9cNI4_0;
	wire w_dff_A_bNf7nTdS6_0;
	wire w_dff_A_67IY7bF71_0;
	wire w_dff_A_KCe3CFxT9_0;
	wire w_dff_A_V9xet9mD8_0;
	wire w_dff_A_Ce1tMWSv9_0;
	wire w_dff_A_lorB278v7_0;
	wire w_dff_A_8sSn4NmT8_0;
	wire w_dff_A_TPK5Ey768_0;
	wire w_dff_A_1LZv9Un12_0;
	wire w_dff_A_loKggvBq6_0;
	wire w_dff_A_FEf1B7nZ7_0;
	wire w_dff_A_2uLs2c3S9_1;
	wire w_dff_A_AhuKunsi1_1;
	wire w_dff_A_pcFbUBcz9_1;
	wire w_dff_A_s3eF31HN8_1;
	wire w_dff_A_MsmPoJDb8_1;
	wire w_dff_A_Xfxgwyf14_1;
	wire w_dff_A_FFB9MV8l1_1;
	wire w_dff_A_LVJrnfm42_1;
	wire w_dff_A_14DWDvVg9_1;
	wire w_dff_A_3upgWeKT5_1;
	wire w_dff_A_kTp2LQFU5_1;
	wire w_dff_A_b2buw0UU4_1;
	wire w_dff_A_OGEALcHA6_1;
	wire w_dff_A_MxjzSkw00_1;
	wire w_dff_A_PWYb19Y21_1;
	wire w_dff_A_f59jYA8P5_0;
	wire w_dff_A_pRmMQpeE8_0;
	wire w_dff_A_QIn5Lzi67_0;
	wire w_dff_A_AjrOsry46_0;
	wire w_dff_A_Qx88tkmG9_0;
	wire w_dff_A_l6vhJiZM3_0;
	wire w_dff_A_isqtWgis2_0;
	wire w_dff_A_ITwmwsQp0_0;
	wire w_dff_A_wBFge4ko1_0;
	wire w_dff_A_ZxDfTi8f3_0;
	wire w_dff_A_wwlGmWnf0_0;
	wire w_dff_A_yTO17ioo5_0;
	wire w_dff_A_Cw8fn0Qz3_0;
	wire w_dff_A_Dgi3RNPu2_0;
	wire w_dff_A_tOFYThyM9_0;
	wire w_dff_A_AUmjnKpy6_0;
	wire w_dff_A_kz696BsN3_0;
	wire w_dff_A_PsC3Z56w8_0;
	wire w_dff_A_32rDj0y51_0;
	wire w_dff_A_awSD8oBC8_0;
	wire w_dff_A_bMTPEd8B3_0;
	wire w_dff_A_KgaLiSJk5_0;
	wire w_dff_A_SifZUAWh9_0;
	wire w_dff_A_WB3qmmwu6_0;
	wire w_dff_A_1mWI1GVB8_0;
	wire w_dff_A_X7CJlDZg1_0;
	wire w_dff_A_HjH7T54d8_1;
	wire w_dff_A_Jjd5WVeh4_1;
	wire w_dff_A_vzidcSnN8_1;
	wire w_dff_A_0BDYz8ZI6_1;
	wire w_dff_A_dSPJwEna1_1;
	wire w_dff_A_wA5Uq0Mn6_1;
	wire w_dff_A_CmdJG8Ph9_1;
	wire w_dff_A_CzKBE1lf3_1;
	wire w_dff_A_J9fnEt7q1_1;
	wire w_dff_A_s4X9JNUG4_1;
	wire w_dff_A_6TGauh890_1;
	wire w_dff_A_4bV3bnYD5_1;
	wire w_dff_A_eSG4JE0Y4_1;
	wire w_dff_A_cyGpAo5m7_1;
	wire w_dff_A_zfRanZFb5_1;
	wire w_dff_B_Vv1U1Xsw1_1;
	wire w_dff_B_8QAkKt3M0_1;
	wire w_dff_B_355MOtrO4_1;
	wire w_dff_B_it2znLd43_1;
	wire w_dff_B_NyDAsDHa5_1;
	wire w_dff_A_ly6rZopT4_0;
	wire w_dff_A_gyXE4MHt9_0;
	wire w_dff_A_iWtpklWD3_0;
	wire w_dff_A_ukOAbM1O3_0;
	wire w_dff_A_KHlim5GW8_0;
	wire w_dff_A_o4Gn8Rp16_0;
	wire w_dff_A_htKJlJg06_0;
	wire w_dff_A_iyv5sVN33_0;
	wire w_dff_A_jUuZdhSc6_0;
	wire w_dff_A_qUxF57Qh6_0;
	wire w_dff_A_Q9c17TY98_0;
	wire w_dff_A_xKPOWsTF8_0;
	wire w_dff_A_C3dt0v0v1_0;
	wire w_dff_A_FZnNBvdh3_0;
	wire w_dff_A_xWYS2Qnl3_0;
	wire w_dff_A_WUcUq3Y59_0;
	wire w_dff_A_8TKz3JAl9_0;
	wire w_dff_A_hMc6BZEG9_0;
	wire w_dff_A_Qp1Rk47H9_0;
	wire w_dff_A_pw1kHjUz2_0;
	wire w_dff_A_6mPWo1Ja7_1;
	wire w_dff_A_b0eEEZzx3_1;
	wire w_dff_A_RChVbdHd9_1;
	wire w_dff_A_Ug4oAg0y9_1;
	wire w_dff_A_CpzthAVL9_1;
	wire w_dff_A_r3ILZe7g6_1;
	wire w_dff_A_jco5sZSn2_1;
	wire w_dff_A_tBcWuE1L0_1;
	wire w_dff_A_f9fvTdNm4_1;
	wire w_dff_A_RzDsK4NF5_1;
	wire w_dff_A_ymJMnyH77_1;
	wire w_dff_A_8JAKO9mK3_1;
	wire w_dff_A_JpuSwqI38_1;
	wire w_dff_A_TlcIV72U0_1;
	wire w_dff_A_EGfukxDR9_1;
	wire w_dff_A_IYKTXbQ26_0;
	wire w_dff_A_3MUahvAy4_0;
	wire w_dff_A_YYeBLsx88_0;
	wire w_dff_A_VYWMwE812_0;
	wire w_dff_A_CmjLWyko3_0;
	wire w_dff_A_9zRzmdzM7_0;
	wire w_dff_A_SyYmKoxZ3_0;
	wire w_dff_A_cU0uybh90_0;
	wire w_dff_A_FClwhfiw9_0;
	wire w_dff_A_gUxxbEq39_0;
	wire w_dff_A_Ee5Gfiu55_0;
	wire w_dff_A_MFKm1KjX7_0;
	wire w_dff_A_1MGRnFlX9_0;
	wire w_dff_A_rBTwsf5d4_0;
	wire w_dff_A_KwV5G41l5_0;
	wire w_dff_A_XQDfzSS13_1;
	wire w_dff_B_fpzEPT5I7_0;
	wire w_dff_B_m25x534I1_0;
	wire w_dff_B_7DzAXQHl2_0;
	wire w_dff_B_LUBtFMM42_0;
	wire w_dff_B_JCNH5Y7g8_0;
	wire w_dff_B_VFPT1eVQ5_0;
	wire w_dff_A_cAgb6sJp5_0;
	wire w_dff_A_UwRY90fB9_0;
	wire w_dff_A_oy9L780f9_0;
	wire w_dff_A_YZGk8nx20_0;
	wire w_dff_A_XGUntYs56_0;
	wire w_dff_A_83uB0iM15_0;
	wire w_dff_A_HlQglHUY2_0;
	wire w_dff_A_bF9J1icF2_0;
	wire w_dff_A_vDrPrNMf5_0;
	wire w_dff_A_zbeykTCV7_0;
	wire w_dff_A_AsDAUV2P7_0;
	wire w_dff_A_MDnOkpYB1_0;
	wire w_dff_B_A5e2h8VR1_2;
	wire w_dff_B_YI0AwNSz6_2;
	wire w_dff_B_2X8y0zbI3_2;
	wire w_dff_B_3tLIWoyx4_2;
	wire w_dff_B_ygig0ASU9_2;
	wire w_dff_B_VUJKNZ2w6_2;
	wire w_dff_B_1M8i8mw79_2;
	wire w_dff_A_TehYMzBl8_0;
	wire w_dff_A_Fn7Iv4Cx7_0;
	wire w_dff_A_HE2idggS8_0;
	wire w_dff_A_yrQ2Xsar7_0;
	wire w_dff_A_2vSLHRkS3_0;
	wire w_dff_A_2iqLDpq24_0;
	wire w_dff_A_OsNwv2H67_0;
	wire w_dff_A_KBGWrlXH4_0;
	wire w_dff_A_2c9lvAsF9_0;
	wire w_dff_A_4C9omT440_0;
	wire w_dff_A_9n1BOoKH9_0;
	wire w_dff_A_HDcVbxuz4_0;
	wire w_dff_A_3z2JhcZs3_0;
	wire w_dff_A_FMq6roSG4_0;
	wire w_dff_A_7U1ypy1a6_0;
	wire w_dff_A_WpQyq9FU3_0;
	wire w_dff_A_0X4VuQBb3_0;
	wire w_dff_A_4KdI0J6J9_0;
	wire w_dff_A_NXAvvox10_0;
	wire w_dff_A_rA6U099P1_0;
	wire w_dff_A_iZIDpyIr3_0;
	wire w_dff_B_NqK5r0uJ8_1;
	wire w_dff_B_KqJio3Rg4_1;
	wire w_dff_B_pYwWI0Mm8_1;
	wire w_dff_B_ka8Zgljp4_1;
	wire w_dff_B_Fyq44NgT7_1;
	wire w_dff_B_ZdKfvdf30_1;
	wire w_dff_B_447HS49Y5_1;
	wire w_dff_B_vJDXMRpC0_1;
	wire w_dff_A_ukWOq8tP3_0;
	wire w_dff_A_YYqfWhRq9_0;
	wire w_dff_A_CXIqUqbt1_0;
	wire w_dff_A_Rmm5znAV3_0;
	wire w_dff_A_iLzFQlOm1_0;
	wire w_dff_A_o9WJ33q89_0;
	wire w_dff_A_fnI5mclx4_0;
	wire w_dff_A_DcKErPU78_0;
	wire w_dff_A_oBfutAC63_0;
	wire w_dff_A_BVrgXk641_0;
	wire w_dff_A_GtwakSja0_0;
	wire w_dff_A_8y8N3Guq4_0;
	wire w_dff_A_j1MTcUuX6_0;
	wire w_dff_A_BTCMwIhv4_0;
	wire w_dff_A_0vTTxGiD2_0;
	wire w_dff_A_YR1Vi4Ty3_0;
	wire w_dff_A_uIcAZ2sq8_0;
	wire w_dff_A_sOSeQPg69_0;
	wire w_dff_B_ppkxjZnz4_2;
	wire w_dff_B_MvqA1pyZ4_2;
	wire w_dff_B_nYPoKPki5_2;
	wire w_dff_B_Z878v3sO5_2;
	wire w_dff_B_bzuIyA295_2;
	wire w_dff_B_NgIky2cZ8_2;
	wire w_dff_B_jlkyKIwC3_2;
	wire w_dff_A_t0fwS1Fi4_0;
	wire w_dff_A_eBAMU7Fu8_0;
	wire w_dff_A_qiARuj7l3_0;
	wire w_dff_A_Fx7tNW6C3_0;
	wire w_dff_A_KQeLt5oc7_0;
	wire w_dff_A_yXhG2H8g8_0;
	wire w_dff_A_PNEJJfWC8_0;
	wire w_dff_A_iXm02h9u9_0;
	wire w_dff_A_ZJXP5Yfj7_0;
	wire w_dff_A_UGzvVhbG3_0;
	wire w_dff_A_TNwq3u6B6_0;
	wire w_dff_B_IOWr197e6_2;
	wire w_dff_B_OkO0mU4i5_2;
	wire w_dff_B_JbGIOMH40_2;
	wire w_dff_B_L9v1PK3V0_2;
	wire w_dff_B_uW5GfRcs4_2;
	wire w_dff_B_s9Nl5gDw7_2;
	wire w_dff_B_aWMZslLJ7_2;
	wire w_dff_B_tFxJeg604_1;
	wire w_dff_B_kNpHvdbT1_0;
	wire w_dff_A_wK59n6K32_0;
	wire w_dff_A_Fot6INnu1_0;
	wire w_dff_A_m4w3asQE4_0;
	wire w_dff_A_ep4zO53T7_0;
	wire w_dff_A_jNCJ47D70_0;
	wire w_dff_A_jvJV2ZFZ2_0;
	wire w_dff_A_q0VOqsmD5_0;
	wire w_dff_A_oYvf3OG94_0;
	wire w_dff_A_qPPMUy726_0;
	wire w_dff_A_7Lu1vTHu9_0;
	wire w_dff_A_mLXAvt4n0_0;
	wire w_dff_B_b4dbHZai5_2;
	wire w_dff_B_eurmNImh1_2;
	wire w_dff_B_Yp7sK7kU0_2;
	wire w_dff_B_FEn4Q8Yo7_2;
	wire w_dff_B_TVEWEfFY6_2;
	wire w_dff_B_MJmaSI9H1_2;
	wire w_dff_B_kRvHPEm09_2;
	wire w_dff_A_iJzAqBOW0_0;
	wire w_dff_A_UBAr06oW3_0;
	wire w_dff_A_zLWEIj8B8_0;
	wire w_dff_A_19qyuNKG3_0;
	wire w_dff_A_eMNfuXmO1_0;
	wire w_dff_A_XMNTUH095_0;
	wire w_dff_A_hB2DIHX84_0;
	wire w_dff_A_tUk0OBpo4_0;
	wire w_dff_A_QdaKPHcP5_0;
	wire w_dff_A_Wkzy1KtS0_0;
	wire w_dff_A_V88cwFC23_0;
	wire w_dff_B_dA3SBpJ68_2;
	wire w_dff_B_G1ZeSt958_2;
	wire w_dff_B_3aBa0O241_2;
	wire w_dff_B_Wus2GaKB4_2;
	wire w_dff_B_5oAjXXeq8_2;
	wire w_dff_B_U9Vb01T34_2;
	wire w_dff_B_93DoIoKW3_2;
	wire w_dff_B_4Hy0jiv52_1;
	wire w_dff_B_ecmWlFWi7_1;
	wire w_dff_B_hhc665Rx5_1;
	wire w_dff_B_AnQhNxo99_1;
	wire w_dff_B_DQXU00sF7_1;
	wire w_dff_B_djL2IWfi4_1;
	wire w_dff_B_awY5TtCk8_1;
	wire w_dff_A_0gGFO1si5_0;
	wire w_dff_A_w5VXco6n2_0;
	wire w_dff_A_O5BubKlF6_0;
	wire w_dff_A_uvZBCxhN2_0;
	wire w_dff_A_IbJJYA8K7_0;
	wire w_dff_A_cRMZYc3B1_0;
	wire w_dff_A_dAdDwizU1_0;
	wire w_dff_A_cIgXDEL30_0;
	wire w_dff_A_1e8abMSn7_0;
	wire w_dff_A_yCXfxgGn8_0;
	wire w_dff_A_dM4HeqPw5_0;
	wire w_dff_B_7S11WjdZ4_2;
	wire w_dff_B_CXrh2OYW4_2;
	wire w_dff_B_6Cbbxs066_2;
	wire w_dff_B_nZFvdqNt7_2;
	wire w_dff_B_ubgIpsNP6_2;
	wire w_dff_B_WMzIhlvR0_2;
	wire w_dff_B_du5n4KHy9_2;
	wire w_dff_A_HsvVj9Sr9_1;
	wire w_dff_A_GfVaUSdR8_1;
	wire w_dff_A_TazNC8XV7_1;
	wire w_dff_A_QCoJQIcB1_1;
	wire w_dff_A_efO9Ivv29_1;
	wire w_dff_A_TLOHSE780_1;
	wire w_dff_A_gevF5jCx6_1;
	wire w_dff_A_W2xbkyoo0_1;
	wire w_dff_A_kPjP12Jp9_1;
	wire w_dff_A_DrfipQrw9_1;
	wire w_dff_A_KAZwzF9R4_1;
	wire w_dff_A_qrbowgNY3_1;
	wire w_dff_A_RC5qWVzk6_1;
	wire w_dff_A_SbUyfcqN9_1;
	wire w_dff_A_UzWk0GRm9_1;
	wire w_dff_A_rN8koomI5_0;
	wire w_dff_A_PzEU658U9_0;
	wire w_dff_A_mOfbwand3_0;
	wire w_dff_A_AkUplPZz5_0;
	wire w_dff_A_UkbINEYs0_0;
	wire w_dff_B_i0JwDmKu3_2;
	wire w_dff_B_nkkH4yCR3_2;
	wire w_dff_B_4zpay2Qy5_2;
	wire w_dff_B_1gHkALnk9_2;
	wire w_dff_B_cqrnNfOR2_2;
	wire w_dff_B_P2897u1Q3_2;
	wire w_dff_B_IaRzRIba6_2;
	wire w_dff_B_Q13EOOKL1_2;
	wire w_dff_B_1GMVD8i19_2;
	wire w_dff_B_J8W4Nmss9_2;
	wire w_dff_B_hbK7XanY0_2;
	wire w_dff_B_180tNT1g1_2;
	wire w_dff_B_KfyEUUMm8_2;
	wire w_dff_B_jWf3GUkZ9_2;
	wire w_dff_A_QD8Sn8xn6_0;
	wire w_dff_A_hnXEFaRo3_0;
	wire w_dff_A_ubLSppHX7_0;
	wire w_dff_A_fChuHLr85_0;
	wire w_dff_A_p5a7Vwgh8_0;
	wire w_dff_A_gj7DxBKd2_0;
	wire w_dff_A_xuEWtplg7_0;
	wire w_dff_A_gHCh00wX9_0;
	wire w_dff_A_56IQBdFD6_0;
	wire w_dff_A_Ntc4VIEX7_0;
	wire w_dff_A_UCyxuw599_0;
	wire w_dff_A_sPIJUNzg2_0;
	wire w_dff_A_fwbZKcqG5_0;
	wire w_dff_A_5Rzh4lej4_0;
	wire w_dff_A_PkvW4NuJ6_0;
	wire w_dff_A_IQsc8pdn6_0;
	wire w_dff_A_qx6bSRxL0_0;
	wire w_dff_A_1ZnpfZau8_0;
	wire w_dff_A_eYlnGbmT1_0;
	wire w_dff_A_YZFvLYFV8_0;
	wire w_dff_A_4ovGi05V3_0;
	wire w_dff_B_NQ6qWZcn7_1;
	wire w_dff_B_MGjLvvx48_1;
	wire w_dff_A_azkryNac6_0;
	wire w_dff_A_NU4en6Er5_0;
	wire w_dff_A_4Obfc4wf3_0;
	wire w_dff_A_TwTZHlF69_0;
	wire w_dff_A_jyiK3bZm1_0;
	wire w_dff_A_hGZTRHHC4_0;
	wire w_dff_A_CphBLeP64_0;
	wire w_dff_A_6LwEWqdP7_0;
	wire w_dff_A_d3psj1Pa9_1;
	wire w_dff_A_jn0pbfpr1_1;
	wire w_dff_A_G66HetqF0_1;
	wire w_dff_A_2DcnsPvc6_1;
	wire w_dff_A_LL1Dh6kU8_1;
	wire w_dff_A_my1kK3pL0_1;
	wire w_dff_A_ofCS9CID6_1;
	wire w_dff_A_T6pXnsGV7_1;
	wire w_dff_A_AH4PL5i43_1;
	wire w_dff_A_i4JLvFh20_1;
	wire w_dff_A_m22eKOdL3_1;
	wire w_dff_A_ETi4jrU66_1;
	wire w_dff_A_JLloTRJ83_1;
	wire w_dff_A_gnRA4fNu1_0;
	wire w_dff_A_7cwWfYfj1_0;
	wire w_dff_A_tF4grip08_0;
	wire w_dff_A_yEMOP4rc7_0;
	wire w_dff_A_7o0mONMx5_0;
	wire w_dff_A_Z6xDi7py5_0;
	wire w_dff_A_keSjFFSW4_0;
	wire w_dff_A_FmMZyJLw4_0;
	wire w_dff_A_GQSUqkXk1_0;
	wire w_dff_A_0GQ949Hm5_0;
	wire w_dff_A_5LXmG0EF7_0;
	wire w_dff_A_OkcAVjAQ3_0;
	wire w_dff_A_7ZIDyrBl4_0;
	wire w_dff_A_tJnszgV80_0;
	wire w_dff_A_5K6pCmpL2_0;
	wire w_dff_A_e9MGPYqX1_0;
	wire w_dff_A_MP349w4b3_0;
	wire w_dff_A_F67Yb6UX5_0;
	wire w_dff_A_Le75QP4r4_0;
	wire w_dff_A_d0c6zVx68_1;
	wire w_dff_A_7n9lGIWn3_1;
	wire w_dff_A_fBde5rFb6_1;
	wire w_dff_A_I8xSQwyx5_1;
	wire w_dff_A_sDy1bD010_1;
	wire w_dff_A_8JQYqsyZ2_1;
	wire w_dff_A_zm39boY64_1;
	wire w_dff_A_tttNuUrm6_1;
	wire w_dff_A_Bn1RDwuN2_0;
	wire w_dff_A_0hA8ov3Z6_0;
	wire w_dff_A_4UeZc7LN8_0;
	wire w_dff_A_1XKNu4IG7_0;
	wire w_dff_A_KphDdd8P5_0;
	wire w_dff_A_HOZpH2xk1_0;
	wire w_dff_A_wj4A0kFJ0_0;
	wire w_dff_A_lTb9FXNb9_0;
	wire w_dff_A_yzggL9pr8_0;
	wire w_dff_A_zhixABwN9_0;
	wire w_dff_A_8r4FoLHq8_0;
	wire w_dff_A_HTtol3Ui3_0;
	wire w_dff_A_Fw3USXt87_0;
	wire w_dff_A_oYqhOt2F2_0;
	wire w_dff_A_H7KaN3Pn9_0;
	wire w_dff_A_G3oHU4zl8_0;
	wire w_dff_A_xGqxvpuB2_0;
	wire w_dff_A_YPeFjJbQ3_0;
	wire w_dff_A_8NTOvryK9_0;
	wire w_dff_A_Wj9TiAki9_1;
	wire w_dff_A_IxTDQcvy2_1;
	wire w_dff_A_0R3kRCOl1_1;
	wire w_dff_A_h5QL0kCJ5_1;
	wire w_dff_A_LYIfWeTe0_1;
	wire w_dff_A_ox9oGVPL0_1;
	wire w_dff_A_n0dbXPoS4_1;
	wire w_dff_A_4RTxeQTv8_1;
	wire w_dff_A_CMuI8L6j7_1;
	wire w_dff_A_G9lrbznW0_1;
	wire w_dff_A_KeFNm4pW6_1;
	wire w_dff_A_kC62ZcDW3_1;
	wire w_dff_A_jcY5vvGb8_1;
	wire w_dff_A_wRopOt5L7_1;
	wire w_dff_A_22tN93cK1_1;
	wire w_dff_A_us47lpq66_1;
	wire w_dff_A_AC2CS2hU4_0;
	wire w_dff_A_shvZ5KCl4_0;
	wire w_dff_A_yPTK2SJA6_0;
	wire w_dff_A_BUk5ewy63_0;
	wire w_dff_A_i5tkwe6P9_0;
	wire w_dff_B_iEHWkATf7_2;
	wire w_dff_B_eWavxSBs5_2;
	wire w_dff_B_GVnRsVxf0_2;
	wire w_dff_B_flLocZ0f0_2;
	wire w_dff_B_8H0gQXti6_2;
	wire w_dff_B_4MgC1ltu4_2;
	wire w_dff_B_A00qhiij1_2;
	wire w_dff_A_lolXuHU57_0;
	wire w_dff_A_druw62o49_0;
	wire w_dff_A_EWhHvAiG8_0;
	wire w_dff_A_Vjp4mi7i3_0;
	wire w_dff_A_uHBZwbJl4_0;
	wire w_dff_A_7h7Fu2Q37_0;
	wire w_dff_A_aBwOw3bx5_0;
	wire w_dff_A_L8UYUXoS7_0;
	wire w_dff_A_wOe423ER8_0;
	wire w_dff_A_VvECfKTc5_0;
	wire w_dff_A_Ca2DWTUk9_0;
	wire w_dff_A_WYBF2niX3_0;
	wire w_dff_A_Eb5WXesu6_0;
	wire w_dff_B_NkP5lfii7_1;
	wire w_dff_B_rpyFMvjf6_0;
	wire w_dff_A_AV111u4x0_0;
	wire w_dff_A_wo8KVVH63_0;
	wire w_dff_A_ccHW2PQS0_0;
	wire w_dff_A_Xhx1JmBs3_0;
	wire w_dff_A_XsWQRDXO9_0;
	wire w_dff_A_4GiB9DAe3_0;
	wire w_dff_B_ceKxluQL1_1;
	wire w_dff_B_ixQvM5mF6_1;
	wire w_dff_B_rwvNWt2F9_1;
	wire w_dff_B_DThuhYie8_1;
	wire w_dff_B_rOFVomLb6_1;
	wire w_dff_B_KXeC1Orn6_1;
	wire w_dff_A_k3fKdYD15_0;
	wire w_dff_A_whBlaFGt4_0;
	wire w_dff_A_CuHV83vG7_0;
	wire w_dff_A_HSg7n5MY5_0;
	wire w_dff_A_cIuwW6t58_0;
	wire w_dff_A_D1ma7eyi6_0;
	wire w_dff_A_EdJiK31x6_0;
	wire w_dff_A_r3BlC9AS4_0;
	wire w_dff_A_Dsjj1ZWE9_0;
	wire w_dff_A_yUVK0bzL0_0;
	wire w_dff_A_bUhEWbP29_0;
	wire w_dff_A_07xr8NJQ7_0;
	wire w_dff_A_IGg9SyEP8_0;
	wire w_dff_A_A4cTJAJG0_1;
	wire w_dff_A_VelxpJ7w3_1;
	wire w_dff_A_pbbzKgfQ3_1;
	wire w_dff_A_CrRJtig80_1;
	wire w_dff_A_16ISkeaI6_1;
	wire w_dff_A_9HJ1m68B0_1;
	wire w_dff_A_MRcXXCTX4_1;
	wire w_dff_A_Go6c1lDV5_1;
	wire w_dff_A_8zIyKzcm6_0;
	wire w_dff_A_BXapyMDz5_0;
	wire w_dff_A_FBcAiRaI0_0;
	wire w_dff_A_jyNHHBvE5_0;
	wire w_dff_A_t01SNbxc5_0;
	wire w_dff_A_LLFs3lMj2_0;
	wire w_dff_A_O0hk1lCZ9_0;
	wire w_dff_A_iy7XwnFi0_0;
	wire w_dff_A_9ClCkjFc1_0;
	wire w_dff_A_nDCd2ZVJ3_0;
	wire w_dff_A_PV5SEcjm8_0;
	wire w_dff_A_TfER06w00_0;
	wire w_dff_A_azgze0TS8_0;
	wire w_dff_A_4T1XvxtM9_0;
	wire w_dff_A_syqbI9W44_0;
	wire w_dff_A_NlPQNhwO8_0;
	wire w_dff_A_Cd7ZuZQ00_0;
	wire w_dff_A_ZMqb7ndf1_0;
	wire w_dff_A_qZdLlFXE3_0;
	wire w_dff_A_6QRAG9CT9_1;
	wire w_dff_A_AcLiwcxi2_1;
	wire w_dff_A_qcwqUm645_1;
	wire w_dff_A_dYv6qkAD3_1;
	wire w_dff_A_dVLWKPsM2_1;
	wire w_dff_A_aGjZh8xo6_1;
	wire w_dff_A_uxhi2cct6_1;
	wire w_dff_A_z7fBMfWI3_1;
	wire w_dff_A_2oNqJcOO7_0;
	wire w_dff_A_HRjeNp6v5_0;
	wire w_dff_A_aQ800rtG2_0;
	wire w_dff_A_2zq3WU0W6_0;
	wire w_dff_A_uV1tepnh5_0;
	wire w_dff_A_sKncualL7_0;
	wire w_dff_A_5RRJF1ak2_1;
	wire w_dff_A_L1yUcqb50_1;
	wire w_dff_A_dkLUS4L14_1;
	wire w_dff_A_2m4pnNzZ3_1;
	wire w_dff_A_euCG29MY4_1;
	wire w_dff_A_GzJpBzPy9_1;
	wire w_dff_A_TQUWBhtX2_0;
	wire w_dff_A_vJIq0LWk4_0;
	wire w_dff_A_NYzJIYwp2_0;
	wire w_dff_A_duF1Fab66_0;
	wire w_dff_A_HqieGEOn9_0;
	wire w_dff_A_STDLK6Qv8_0;
	wire w_dff_A_nZgFW8Dk0_0;
	wire w_dff_A_EV2WFCl09_0;
	wire w_dff_A_MvLqRxip3_1;
	wire w_dff_A_wLWdPZcw9_1;
	wire w_dff_A_bLQHGVVf3_1;
	wire w_dff_A_VFNv39zM4_1;
	wire w_dff_A_bvzu4eKc1_1;
	wire w_dff_A_O7QdYVcU6_1;
	wire w_dff_A_NazXc7KQ6_1;
	wire w_dff_A_7yy3x1e71_1;
	wire w_dff_A_xPBJ9FAM0_1;
	wire w_dff_A_fQLewJoZ8_1;
	wire w_dff_A_9vng2tpv8_1;
	wire w_dff_A_chPBt41z6_1;
	wire w_dff_A_xwKVzm7V8_1;
	wire w_dff_A_BRBQYKct3_0;
	wire w_dff_A_7nwawlw80_0;
	wire w_dff_A_IOns0ZG35_0;
	wire w_dff_A_0UIFhdOv2_0;
	wire w_dff_A_DZmf4tuv4_0;
	wire w_dff_A_YjxOWqGe8_0;
	wire w_dff_B_YwTz4Rdk3_1;
	wire w_dff_B_13jNcIH78_1;
	wire w_dff_A_JInPuuqa8_0;
	wire w_dff_A_G1Aw1gSS7_0;
	wire w_dff_A_aNspGlsp1_0;
	wire w_dff_A_GDQYNaQN9_0;
	wire w_dff_A_kSn583jH5_0;
	wire w_dff_A_TBubJOYM9_0;
	wire w_dff_A_8WMfvOJY9_0;
	wire w_dff_A_B6ddvVpF3_0;
	wire w_dff_A_IaUakkkr1_0;
	wire w_dff_A_fk6MrzLy9_0;
	wire w_dff_A_UMoQmOdK2_0;
	wire w_dff_A_qqnjVmhM7_0;
	wire w_dff_A_hrgFTxrx9_0;
	wire w_dff_A_7AlZQU0f4_0;
	wire w_dff_A_9mFFV7fQ3_0;
	wire w_dff_A_XFRjWb0e7_0;
	wire w_dff_A_AB5AJAx93_0;
	wire w_dff_A_7sx2afBE9_0;
	wire w_dff_A_rlN0UfkF4_0;
	wire w_dff_A_ZeyIuTAQ0_0;
	wire w_dff_A_XfAAkZ0G4_0;
	wire w_dff_A_s1kCKJxT9_0;
	wire w_dff_A_JwZoJf724_0;
	wire w_dff_A_2sB8qnBj9_0;
	wire w_dff_A_dmo9lwF68_0;
	wire w_dff_A_cN0njtaj5_0;
	wire w_dff_A_uwlUsmnk9_0;
	wire w_dff_A_CNqPklHs0_0;
	wire w_dff_A_EODEH6fW7_0;
	wire w_dff_A_GjiScDiW3_0;
	wire w_dff_A_R73CpPBc0_0;
	wire w_dff_A_nhp2kmJQ0_0;
	wire w_dff_A_X3q7bKiM4_0;
	wire w_dff_A_RNTOFx799_0;
	wire w_dff_A_SN7SJ5w29_0;
	wire w_dff_A_Y8ekKrsm4_0;
	wire w_dff_A_IqGY3AHw1_0;
	wire w_dff_A_bSHxnqms8_0;
	wire w_dff_A_anc3jKno6_0;
	wire w_dff_A_AOrQJtKy9_0;
	wire w_dff_A_YHIgEvW72_0;
	wire w_dff_A_M8ITuz5Y3_0;
	wire w_dff_A_hXIi3Tfy1_0;
	wire w_dff_A_ReeXbjtY2_0;
	wire w_dff_A_9ygUFtzK9_0;
	wire w_dff_A_cGZvoynY1_1;
	wire w_dff_A_TPD2k8Xz9_1;
	wire w_dff_A_TqNdzYTj2_1;
	wire w_dff_A_ETYGaLcs1_1;
	wire w_dff_A_kkX8SL0T2_1;
	wire w_dff_A_1J93v6sV9_1;
	wire w_dff_A_uMKEEnY32_1;
	wire w_dff_A_2UsyUsik1_1;
	wire w_dff_A_XHwaf2sQ1_0;
	wire w_dff_A_9NlhitPg0_0;
	wire w_dff_A_omjH5Oei0_0;
	wire w_dff_A_nhH959ff2_0;
	wire w_dff_A_xQEWaPFd4_0;
	wire w_dff_B_ixIUlemi6_2;
	wire w_dff_B_oN58kuea0_2;
	wire w_dff_B_Q9b2boXO0_2;
	wire w_dff_B_vHmKgquF2_2;
	wire w_dff_B_t6OXCiwM1_2;
	wire w_dff_B_yn1gTL1Z5_2;
	wire w_dff_B_IF04gzgP6_2;
	wire w_dff_A_bU10WHIn3_0;
	wire w_dff_A_hvrbYllE2_0;
	wire w_dff_A_TxrgJKPe2_0;
	wire w_dff_A_3UCTd4K72_0;
	wire w_dff_A_QMSVHAYt5_0;
	wire w_dff_A_hyeI8XLQ6_0;
	wire w_dff_A_Cz0JYlKT3_0;
	wire w_dff_A_h8TvgjHo5_0;
	wire w_dff_A_GwkEOQSb7_0;
	wire w_dff_A_HivPc0ry6_0;
	wire w_dff_A_NSJpxvh96_0;
	wire w_dff_A_PjSU1GIe5_0;
	wire w_dff_A_YZreO8RO2_0;
	wire w_dff_A_HUmFkQhw3_1;
	wire w_dff_A_EKVT5ugf1_1;
	wire w_dff_A_AZ5gkIHl5_1;
	wire w_dff_A_mj4enfqA6_1;
	wire w_dff_A_b3uE29Xi6_1;
	wire w_dff_A_SfkfkjLP5_1;
	wire w_dff_A_ilKvU5Xf7_1;
	wire w_dff_A_EE1vAm416_1;
	wire w_dff_A_U9Sinh8X8_0;
	wire w_dff_A_1CKWLqAN1_0;
	wire w_dff_A_1jdCjZXD7_0;
	wire w_dff_A_ScTkoQ8O2_0;
	wire w_dff_A_4sJ3XD5G4_0;
	wire w_dff_A_zUsGRMpU8_0;
	wire w_dff_B_iVWKt9F30_1;
	wire w_dff_B_7OeTX8tP1_1;
	wire w_dff_A_cLYJzDLR9_0;
	wire w_dff_A_9d8Zy8bX8_0;
	wire w_dff_A_I8zY70O09_0;
	wire w_dff_A_nKaof8P33_0;
	wire w_dff_A_AsYHRkx51_0;
	wire w_dff_A_kwJpDK9d3_0;
	wire w_dff_A_pJCoHLR02_0;
	wire w_dff_A_SeAMmSL87_0;
	wire w_dff_A_qakHzVMB1_0;
	wire w_dff_A_NZCBwXPu8_0;
	wire w_dff_A_8Ff8nEbI3_0;
	wire w_dff_A_6gIMxOOk2_0;
	wire w_dff_A_NE6oXFhM3_0;
	wire w_dff_A_jCLSgv0p3_2;
	wire w_dff_A_pRmSFdzO9_0;
	wire w_dff_A_tW2aJNWD6_0;
	wire w_dff_A_eTIT3P1E9_0;
	wire w_dff_A_lbMIEfNe9_0;
	wire w_dff_A_iOnzaU6I2_0;
	wire w_dff_A_9dUrKNKd3_0;
	wire w_dff_A_0ivgQ7UW7_1;
	wire w_dff_A_sQG3aNIQ2_0;
	wire w_dff_A_NSLkkRcy3_0;
	wire w_dff_A_NZvhiyj07_0;
	wire w_dff_A_TtnypJFA6_0;
	wire w_dff_A_JuVeqah71_0;
	wire w_dff_A_VfX4Xf9w3_0;
	wire w_dff_A_9RG3yveU9_0;
	wire w_dff_A_27ER9Jzv1_0;
	wire w_dff_A_tSk2aKxK9_0;
	wire w_dff_A_R0n8zemA2_0;
	wire w_dff_A_wyeJougk1_0;
	wire w_dff_A_rq5gl4iL9_0;
	wire w_dff_A_1s5F0kqf1_0;
	wire w_dff_A_m3tq5pOZ7_2;
	wire w_dff_A_bc99Wd5Z3_0;
	wire w_dff_A_vtgvAEaQ7_0;
	wire w_dff_A_jei1LsGN8_0;
	wire w_dff_A_sOO6HaqA6_0;
	wire w_dff_A_d2JnQgsp2_0;
	wire w_dff_A_lKn6yJlJ6_0;
	wire w_dff_A_TRRJesDS2_1;
	wire w_dff_A_xVmFd9Dm5_0;
	wire w_dff_A_uMGYBVYl1_0;
	wire w_dff_A_EiSnpKIJ6_0;
	wire w_dff_A_T7qDgt7E6_0;
	wire w_dff_A_dOTcBzwc9_0;
	wire w_dff_A_gGNBgYqU5_0;
	wire w_dff_A_pcgnEsJ98_0;
	wire w_dff_A_GmnGWvfI8_0;
	wire w_dff_A_VHqVsIXk3_0;
	wire w_dff_A_2D6P5aMx2_0;
	wire w_dff_A_WiWzKvF72_0;
	wire w_dff_A_S1nC82Tx3_0;
	wire w_dff_A_u2Wkcub51_0;
	wire w_dff_A_CPVaA3YE2_2;
	wire w_dff_A_hl3QBdk34_0;
	wire w_dff_A_M4NHu0WP6_0;
	wire w_dff_A_2GBha37m9_0;
	wire w_dff_A_dTgi6XPn2_0;
	wire w_dff_A_7fGXVDn78_0;
	wire w_dff_A_9feHHqEP9_0;
	wire w_dff_A_ZUmlp4ih2_1;
	wire w_dff_A_893RPwEf4_0;
	wire w_dff_A_luoqwI3p0_0;
	wire w_dff_A_dZEkaBhF4_0;
	wire w_dff_A_QWq5YH7x7_0;
	wire w_dff_A_s3FmS4px5_0;
	wire w_dff_A_2z1I5Puz3_0;
	wire w_dff_A_ULD4DwGY1_0;
	wire w_dff_A_VeGUxuiq8_0;
	wire w_dff_A_ZKU1lP1t1_0;
	wire w_dff_A_NMfp3Yml3_0;
	wire w_dff_A_5iMHirOA5_0;
	wire w_dff_A_2jtw5R4j9_0;
	wire w_dff_A_EcgTezgs3_0;
	wire w_dff_A_wfQ7uCxp3_0;
	wire w_dff_A_GiJdxXtb8_0;
	wire w_dff_A_bgcdtyLP4_0;
	wire w_dff_A_0bQ4fxyL7_0;
	wire w_dff_A_eSJpdP357_0;
	wire w_dff_A_C69Ak8SM2_0;
	wire w_dff_A_m4p2c9nk5_0;
	wire w_dff_A_A1f7VNc53_0;
	wire w_dff_A_xY1SuJ7Y7_0;
	wire w_dff_A_INVL3gxL2_0;
	wire w_dff_A_mziMIdWz5_0;
	wire w_dff_A_KULj1DkY4_0;
	wire w_dff_A_dZOlZMLW4_1;
	wire w_dff_A_LVGuxcLB1_1;
	wire w_dff_A_wmTR8ict7_1;
	wire w_dff_A_yFShnhJM9_1;
	wire w_dff_A_ZMA7FEMY9_1;
	wire w_dff_A_qhPKt9yi6_1;
	wire w_dff_A_ySmVm7jB4_1;
	wire w_dff_A_oiBtZd8U0_1;
	wire w_dff_A_FBpKnxet5_1;
	wire w_dff_A_fYIfsCf14_1;
	wire w_dff_A_xozF5Ach0_1;
	wire w_dff_A_pdTn0NBz5_1;
	wire w_dff_A_UrBp0ROh1_1;
	wire w_dff_A_SbqqBJrZ8_1;
	wire w_dff_A_PcM4HkA08_1;
	wire w_dff_A_Ht3awnJL8_1;
	wire w_dff_A_2ixDfRJv6_1;
	wire w_dff_A_j3CELniN6_1;
	wire w_dff_A_p3oH2QIB6_1;
	wire w_dff_A_c91kfoCy9_1;
	wire w_dff_A_x2trJ02B9_1;
	wire w_dff_A_KLpJZTcl2_1;
	wire w_dff_A_t52nroUK4_1;
	wire w_dff_A_68hQuQow0_2;
	wire w_dff_A_UAyRo1Zw5_2;
	wire w_dff_A_cZX06fTd3_2;
	wire w_dff_A_rhNdrFvP2_2;
	wire w_dff_A_84alNLuP1_2;
	wire w_dff_A_3RBbZaOv7_2;
	wire w_dff_A_HM7Xt9M00_2;
	wire w_dff_A_sns6gJAF5_0;
	wire w_dff_A_ygNnZWiE9_0;
	wire w_dff_A_UYxhPOTK9_0;
	wire w_dff_A_OstBHuum1_0;
	wire w_dff_A_LXonWnii7_0;
	wire w_dff_A_ReADckMX0_0;
	wire w_dff_A_4tjV6s9y4_0;
	wire w_dff_A_44Q1Hx1w5_0;
	wire w_dff_A_ErKFxt4K2_0;
	wire w_dff_A_l0mWy9y61_0;
	wire w_dff_A_QmPZJawy2_0;
	wire w_dff_A_mVgvovWA6_0;
	wire w_dff_A_s7Pv9KOO4_0;
	wire w_dff_A_TclB1t9Z4_0;
	wire w_dff_A_GkEWWy088_2;
	wire w_dff_A_VhMnQ70e8_0;
	wire w_dff_A_RbLgk9ah9_0;
	wire w_dff_A_NcyuVqO52_0;
	wire w_dff_A_FKAcYUAm7_0;
	wire w_dff_A_cLWxCmsI0_0;
	wire w_dff_A_w7lt1dcp9_0;
	wire w_dff_A_AuOKD7660_1;
	wire w_dff_A_LaLU8o9Q5_0;
	wire w_dff_A_CCVTszga5_0;
	wire w_dff_A_52ov8LUL3_0;
	wire w_dff_A_tN7AdNdI6_0;
	wire w_dff_A_HE4889sh5_0;
	wire w_dff_A_jCXMQBrh3_0;
	wire w_dff_A_1r8vJFC17_0;
	wire w_dff_A_5hpQmw7i6_0;
	wire w_dff_A_Y53OLZNa4_0;
	wire w_dff_A_VqdGLU0k9_0;
	wire w_dff_A_VUb1qwie9_0;
	wire w_dff_A_i1HZzGEE2_0;
	wire w_dff_A_KATBrZG45_0;
	wire w_dff_A_2GQp74W96_2;
	wire w_dff_A_oZF4Mh1o2_0;
	wire w_dff_A_DC01FJdH6_0;
	wire w_dff_A_2N3DnU7i7_0;
	wire w_dff_A_gyI1bUZ51_0;
	wire w_dff_A_e7Fk9voQ8_0;
	wire w_dff_A_X0lqFf1U5_0;
	wire w_dff_A_asY2EJUK6_1;
	wire w_dff_A_iICP0BMf4_0;
	wire w_dff_A_5Q2BFT2c6_0;
	wire w_dff_A_cSSoVR0x0_0;
	wire w_dff_A_tH7PkBp22_0;
	wire w_dff_A_BvclH8Jb5_0;
	wire w_dff_A_DfSg4lqe1_0;
	wire w_dff_A_pOArUeeG7_0;
	wire w_dff_A_kAOLIRaY0_0;
	wire w_dff_A_A8Ooo5bE8_0;
	wire w_dff_A_hKHameyp3_0;
	wire w_dff_A_Jtk8u1bt3_0;
	wire w_dff_A_UnP2Bxod0_0;
	wire w_dff_A_7wRvwOcp8_0;
	wire w_dff_A_CDaLzzUH4_2;
	wire w_dff_A_EMEt9F877_0;
	wire w_dff_A_vP4Y4k477_0;
	wire w_dff_A_ZQ72B3iZ6_0;
	wire w_dff_A_B7Epgujb4_0;
	wire w_dff_A_ywAkzHm66_1;
	wire w_dff_B_Ml2pD0BU8_1;
	wire w_dff_A_Gv5iyWLq3_0;
	wire w_dff_A_OQjvPBdC0_0;
	wire w_dff_A_FDkYign09_0;
	wire w_dff_A_Q0N3R1ey1_0;
	wire w_dff_A_sOhfZZak9_0;
	wire w_dff_A_q6JCB2dB3_0;
	wire w_dff_A_XNVAdMtj9_0;
	wire w_dff_A_GRRshK6s2_0;
	wire w_dff_A_gyc3Z5Gb4_0;
	wire w_dff_A_PXIAEZS05_0;
	wire w_dff_A_qgQcvee10_0;
	wire w_dff_A_wbdwtidA6_0;
	wire w_dff_A_MieW2VVm4_0;
	wire w_dff_A_ebpXr9Hh7_1;
	wire w_dff_A_NucbvHI39_1;
	wire w_dff_A_iWOI8SEZ1_1;
	wire w_dff_A_MbjdOFz08_1;
	wire w_dff_A_gvY4XCXn2_1;
	wire w_dff_A_SH013tnM8_1;
	wire w_dff_A_IAtl95gj8_1;
	wire w_dff_A_W3svUPV46_1;
	wire w_dff_A_4i46PGmI0_2;
	wire w_dff_A_xAe2rTE61_0;
	wire w_dff_A_2znjptDJ4_0;
	wire w_dff_A_UfIjYvQB1_0;
	wire w_dff_A_TNcbctzq1_0;
	wire w_dff_A_YwwioSY85_0;
	wire w_dff_A_N65usaMv8_0;
	wire w_dff_A_45DDNgtQ3_0;
	wire w_dff_A_o6ixDT2s2_0;
	wire w_dff_A_pz45IahK8_0;
	wire w_dff_A_JaxLAtvC3_0;
	wire w_dff_A_70y3XZk07_0;
	wire w_dff_A_WfdLipTW7_0;
	wire w_dff_A_cnpsrrmk0_0;
	wire w_dff_A_mWIZI3vw2_0;
	wire w_dff_A_9vXIbKq39_0;
	wire w_dff_A_zUzEfCVk4_0;
	wire w_dff_A_81gjaSbA7_0;
	wire w_dff_A_ojfR0qZ85_0;
	wire w_dff_A_bgSF60ae4_0;
	wire w_dff_A_7z1ywyqd3_0;
	wire w_dff_A_ObiHwby38_0;
	wire w_dff_A_usOypx327_0;
	wire w_dff_A_zdoTkP3m3_1;
	wire w_dff_A_SEMGl6Zg8_1;
	wire w_dff_A_FgI7NOuD4_0;
	wire w_dff_A_W85J9Emz9_0;
	wire w_dff_A_6RXb5wTr2_0;
	wire w_dff_A_yAs7j40J5_0;
	wire w_dff_A_nxGMixCD4_0;
	wire w_dff_A_iBZzaS8T9_0;
	wire w_dff_A_fo5d3vHc4_0;
	wire w_dff_A_cxMmrtHl2_0;
	wire w_dff_A_jEd241Z64_0;
	wire w_dff_A_uHCETZMJ0_0;
	wire w_dff_A_mIpwl0R25_0;
	wire w_dff_A_KSXBSmRr2_0;
	wire w_dff_A_HrY8qfug8_0;
	wire w_dff_A_F6lggsDY0_0;
	wire w_dff_A_5ANkbwFV0_0;
	wire w_dff_A_bl0NvcbN2_0;
	wire w_dff_A_fU2MW94j0_0;
	wire w_dff_A_N81KYzpx5_0;
	wire w_dff_A_8gq10dYw0_0;
	wire w_dff_A_7QgaQTST6_0;
	wire w_dff_A_n8EDLT5F7_1;
	wire w_dff_A_g5CDUu0d0_0;
	wire w_dff_A_QGRhmXyi2_0;
	wire w_dff_A_046ZAo3f0_0;
	wire w_dff_A_p08ej82O1_0;
	wire w_dff_A_CSDyzqPJ5_0;
	wire w_dff_A_NrCqfr6e4_0;
	wire w_dff_A_yhzrV6pF0_0;
	wire w_dff_A_lrl24h1E3_0;
	wire w_dff_A_43gH8nQM2_0;
	wire w_dff_A_qXojXBgN6_0;
	wire w_dff_A_9FNc9TVV7_0;
	wire w_dff_A_UuQOzaaV8_0;
	wire w_dff_A_p8mRBsUd9_0;
	wire w_dff_A_yBeS5tNQ7_2;
	wire w_dff_A_a9rIOCa60_0;
	wire w_dff_A_aDqauZ9T3_0;
	wire w_dff_A_u0dyAunK0_0;
	wire w_dff_A_KTsi93jF9_0;
	wire w_dff_A_iswhRiWp5_0;
	wire w_dff_A_z3jNHQMA0_0;
	wire w_dff_A_azFe6ujw4_1;
	wire w_dff_A_2cvsLWe78_0;
	jnot g000(.din(w_G102gat_0[1]),.dout(n43),.clk(gclk));
	jand g001(.dina(w_G108gat_0[2]),.dinb(w_n43_0[1]),.dout(n44),.clk(gclk));
	jnot g002(.din(w_G43gat_0[1]),.dout(n45),.clk(gclk));
	jor g003(.dina(w_n45_0[1]),.dinb(w_dff_B_Ml2pD0BU8_1),.dout(n46),.clk(gclk));
	jnot g004(.din(w_n46_0[2]),.dout(n47),.clk(gclk));
	jor g005(.dina(w_n47_0[1]),.dinb(w_n44_0[1]),.dout(n48),.clk(gclk));
	jnot g006(.din(w_G63gat_0[2]),.dout(n49),.clk(gclk));
	jand g007(.dina(w_G69gat_0[2]),.dinb(w_n49_0[1]),.dout(n50),.clk(gclk));
	jnot g008(.din(w_G11gat_0[2]),.dout(n51),.clk(gclk));
	jand g009(.dina(w_G17gat_0[2]),.dinb(w_n51_0[1]),.dout(n52),.clk(gclk));
	jor g010(.dina(n52),.dinb(n50),.dout(n53),.clk(gclk));
	jnot g011(.din(w_G24gat_0[2]),.dout(n54),.clk(gclk));
	jand g012(.dina(w_G30gat_0[2]),.dinb(w_n54_0[1]),.dout(n55),.clk(gclk));
	jnot g013(.din(w_G50gat_0[1]),.dout(n56),.clk(gclk));
	jand g014(.dina(w_G56gat_1[1]),.dinb(n56),.dout(n57),.clk(gclk));
	jor g015(.dina(w_n57_0[1]),.dinb(n55),.dout(n58),.clk(gclk));
	jor g016(.dina(n58),.dinb(n53),.dout(n59),.clk(gclk));
	jnot g017(.din(w_G1gat_0[2]),.dout(n60),.clk(gclk));
	jand g018(.dina(w_G4gat_0[2]),.dinb(w_n60_0[1]),.dout(n61),.clk(gclk));
	jnot g019(.din(w_G89gat_0[2]),.dout(n62),.clk(gclk));
	jand g020(.dina(w_G95gat_0[2]),.dinb(w_n62_0[1]),.dout(n63),.clk(gclk));
	jnot g021(.din(w_G76gat_0[2]),.dout(n64),.clk(gclk));
	jand g022(.dina(w_G82gat_0[2]),.dinb(w_n64_0[1]),.dout(n65),.clk(gclk));
	jor g023(.dina(n65),.dinb(n63),.dout(n66),.clk(gclk));
	jor g024(.dina(n66),.dinb(w_dff_B_13jNcIH78_1),.dout(n67),.clk(gclk));
	jor g025(.dina(n67),.dinb(n59),.dout(n68),.clk(gclk));
	jor g026(.dina(n68),.dinb(w_dff_B_YwTz4Rdk3_1),.dout(G223gat_fa_),.clk(gclk));
	jnot g027(.din(w_G21gat_0[2]),.dout(n70),.clk(gclk));
	jnot g028(.din(w_n44_0[0]),.dout(n71),.clk(gclk));
	jand g029(.dina(w_n46_0[1]),.dinb(n71),.dout(n72),.clk(gclk));
	jnot g030(.din(w_G69gat_0[1]),.dout(n73),.clk(gclk));
	jor g031(.dina(w_n73_0[1]),.dinb(w_G63gat_0[1]),.dout(n74),.clk(gclk));
	jnot g032(.din(w_G17gat_0[1]),.dout(n75),.clk(gclk));
	jor g033(.dina(w_n75_0[1]),.dinb(w_G11gat_0[1]),.dout(n76),.clk(gclk));
	jand g034(.dina(n76),.dinb(n74),.dout(n77),.clk(gclk));
	jnot g035(.din(w_G30gat_0[1]),.dout(n78),.clk(gclk));
	jor g036(.dina(w_n78_0[1]),.dinb(w_G24gat_0[1]),.dout(n79),.clk(gclk));
	jnot g037(.din(w_G56gat_1[0]),.dout(n80),.clk(gclk));
	jor g038(.dina(w_n80_0[1]),.dinb(w_G50gat_0[0]),.dout(n81),.clk(gclk));
	jand g039(.dina(w_n81_0[1]),.dinb(n79),.dout(n82),.clk(gclk));
	jand g040(.dina(n82),.dinb(n77),.dout(n83),.clk(gclk));
	jnot g041(.din(w_G4gat_0[1]),.dout(n84),.clk(gclk));
	jor g042(.dina(w_n84_0[1]),.dinb(w_G1gat_0[1]),.dout(n85),.clk(gclk));
	jnot g043(.din(w_G95gat_0[1]),.dout(n86),.clk(gclk));
	jor g044(.dina(w_n86_0[1]),.dinb(w_G89gat_0[1]),.dout(n87),.clk(gclk));
	jnot g045(.din(w_G82gat_0[1]),.dout(n88),.clk(gclk));
	jor g046(.dina(w_n88_0[1]),.dinb(w_G76gat_0[1]),.dout(n89),.clk(gclk));
	jand g047(.dina(n89),.dinb(n87),.dout(n90),.clk(gclk));
	jand g048(.dina(n90),.dinb(w_dff_B_7OeTX8tP1_1),.dout(n91),.clk(gclk));
	jand g049(.dina(n91),.dinb(n83),.dout(n92),.clk(gclk));
	jand g050(.dina(n92),.dinb(w_dff_B_iVWKt9F30_1),.dout(n93),.clk(gclk));
	jor g051(.dina(w_n93_3[2]),.dinb(w_n51_0[0]),.dout(n94),.clk(gclk));
	jand g052(.dina(n94),.dinb(w_G17gat_0[0]),.dout(n95),.clk(gclk));
	jand g053(.dina(w_n95_0[1]),.dinb(w_n70_0[1]),.dout(n96),.clk(gclk));
	jnot g054(.din(w_G99gat_0[2]),.dout(n97),.clk(gclk));
	jor g055(.dina(w_n93_3[1]),.dinb(w_n62_0[0]),.dout(n98),.clk(gclk));
	jand g056(.dina(n98),.dinb(w_G95gat_0[0]),.dout(n99),.clk(gclk));
	jand g057(.dina(n99),.dinb(w_dff_B_awY5TtCk8_1),.dout(n100),.clk(gclk));
	jor g058(.dina(n100),.dinb(n96),.dout(n101),.clk(gclk));
	jnot g059(.din(w_G73gat_0[2]),.dout(n102),.clk(gclk));
	jor g060(.dina(w_n93_3[0]),.dinb(w_n49_0[0]),.dout(n103),.clk(gclk));
	jand g061(.dina(n103),.dinb(w_G69gat_0[0]),.dout(n104),.clk(gclk));
	jand g062(.dina(w_n104_0[1]),.dinb(w_n102_0[1]),.dout(n105),.clk(gclk));
	jnot g063(.din(w_G34gat_0[2]),.dout(n106),.clk(gclk));
	jor g064(.dina(w_n93_2[2]),.dinb(w_n54_0[0]),.dout(n107),.clk(gclk));
	jand g065(.dina(n107),.dinb(w_G30gat_0[0]),.dout(n108),.clk(gclk));
	jand g066(.dina(w_n108_0[1]),.dinb(w_n106_0[1]),.dout(n109),.clk(gclk));
	jor g067(.dina(n109),.dinb(n105),.dout(n110),.clk(gclk));
	jnot g068(.din(w_G112gat_0[2]),.dout(n111),.clk(gclk));
	jor g069(.dina(w_n93_2[1]),.dinb(w_n43_0[0]),.dout(n112),.clk(gclk));
	jand g070(.dina(n112),.dinb(w_G108gat_0[1]),.dout(n113),.clk(gclk));
	jand g071(.dina(w_n113_0[1]),.dinb(w_n111_0[1]),.dout(n114),.clk(gclk));
	jor g072(.dina(w_dff_B_kNpHvdbT1_0),.dinb(n110),.dout(n115),.clk(gclk));
	jor g073(.dina(n115),.dinb(w_dff_B_tFxJeg604_1),.dout(n116),.clk(gclk));
	jnot g074(.din(w_G60gat_0[1]),.dout(n117),.clk(gclk));
	jxor g075(.dina(w_n93_2[0]),.dinb(w_n57_0[0]),.dout(n118),.clk(gclk));
	jand g076(.dina(n118),.dinb(w_G56gat_0[2]),.dout(n119),.clk(gclk));
	jand g077(.dina(w_n119_0[2]),.dinb(w_n117_0[1]),.dout(n120),.clk(gclk));
	jnot g078(.din(w_G86gat_0[2]),.dout(n121),.clk(gclk));
	jor g079(.dina(w_n93_1[2]),.dinb(w_n64_0[0]),.dout(n122),.clk(gclk));
	jand g080(.dina(n122),.dinb(w_G82gat_0[0]),.dout(n123),.clk(gclk));
	jand g081(.dina(w_n123_0[1]),.dinb(w_n121_0[1]),.dout(n124),.clk(gclk));
	jnot g082(.din(w_G8gat_0[2]),.dout(n125),.clk(gclk));
	jor g083(.dina(w_n93_1[1]),.dinb(w_n60_0[0]),.dout(n126),.clk(gclk));
	jand g084(.dina(n126),.dinb(w_G4gat_0[0]),.dout(n127),.clk(gclk));
	jand g085(.dina(w_n127_0[1]),.dinb(w_n125_0[1]),.dout(n128),.clk(gclk));
	jnot g086(.din(w_G47gat_0[2]),.dout(n129),.clk(gclk));
	jor g087(.dina(w_n93_1[0]),.dinb(w_n47_0[0]),.dout(n130),.clk(gclk));
	jand g088(.dina(n130),.dinb(w_G43gat_0[0]),.dout(n131),.clk(gclk));
	jand g089(.dina(w_n131_0[2]),.dinb(w_dff_B_vJDXMRpC0_1),.dout(n132),.clk(gclk));
	jor g090(.dina(n132),.dinb(n128),.dout(n133),.clk(gclk));
	jor g091(.dina(n133),.dinb(w_dff_B_NqK5r0uJ8_1),.dout(n134),.clk(gclk));
	jor g092(.dina(n134),.dinb(w_n120_0[1]),.dout(n135),.clk(gclk));
	jor g093(.dina(n135),.dinb(n116),.dout(G329gat_fa_),.clk(gclk));
	jand g094(.dina(w_G223gat_4),.dinb(w_G89gat_0[0]),.dout(n137),.clk(gclk));
	jor g095(.dina(n137),.dinb(w_n86_0[0]),.dout(n138),.clk(gclk));
	jand g096(.dina(w_G329gat_4),.dinb(w_G99gat_0[1]),.dout(n139),.clk(gclk));
	jor g097(.dina(n139),.dinb(w_n138_0[1]),.dout(n140),.clk(gclk));
	jor g098(.dina(w_n140_0[1]),.dinb(w_G105gat_0[1]),.dout(n141),.clk(gclk));
	jnot g099(.din(w_n141_0[1]),.dout(n142),.clk(gclk));
	jand g100(.dina(w_G329gat_3[2]),.dinb(w_G47gat_0[1]),.dout(n143),.clk(gclk));
	jnot g101(.din(n143),.dout(n144),.clk(gclk));
	jnot g102(.din(w_G53gat_0[1]),.dout(n145),.clk(gclk));
	jand g103(.dina(w_n131_0[1]),.dinb(w_n145_0[1]),.dout(n146),.clk(gclk));
	jand g104(.dina(w_dff_B_VFPT1eVQ5_0),.dinb(w_n144_0[1]),.dout(n147),.clk(gclk));
	jor g105(.dina(w_n147_0[1]),.dinb(n142),.dout(n148),.clk(gclk));
	jnot g106(.din(w_G40gat_0[1]),.dout(n149),.clk(gclk));
	jand g107(.dina(w_G223gat_3[2]),.dinb(w_G11gat_0[0]),.dout(n150),.clk(gclk));
	jor g108(.dina(n150),.dinb(w_n75_0[0]),.dout(n151),.clk(gclk));
	jor g109(.dina(w_n151_0[1]),.dinb(w_G21gat_0[1]),.dout(n152),.clk(gclk));
	jor g110(.dina(w_n138_0[0]),.dinb(w_G99gat_0[0]),.dout(n153),.clk(gclk));
	jand g111(.dina(n153),.dinb(n152),.dout(n154),.clk(gclk));
	jand g112(.dina(w_G223gat_3[1]),.dinb(w_G63gat_0[0]),.dout(n155),.clk(gclk));
	jor g113(.dina(n155),.dinb(w_n73_0[0]),.dout(n156),.clk(gclk));
	jor g114(.dina(w_n156_0[1]),.dinb(w_G73gat_0[1]),.dout(n157),.clk(gclk));
	jand g115(.dina(w_G223gat_3[0]),.dinb(w_G24gat_0[0]),.dout(n158),.clk(gclk));
	jor g116(.dina(n158),.dinb(w_n78_0[0]),.dout(n159),.clk(gclk));
	jor g117(.dina(w_n159_0[1]),.dinb(w_G34gat_0[1]),.dout(n160),.clk(gclk));
	jand g118(.dina(n160),.dinb(n157),.dout(n161),.clk(gclk));
	jnot g119(.din(w_G108gat_0[0]),.dout(n162),.clk(gclk));
	jand g120(.dina(w_G223gat_2[2]),.dinb(w_G102gat_0[0]),.dout(n163),.clk(gclk));
	jor g121(.dina(n163),.dinb(w_dff_B_KXeC1Orn6_1),.dout(n164),.clk(gclk));
	jor g122(.dina(w_n164_0[1]),.dinb(w_G112gat_0[1]),.dout(n165),.clk(gclk));
	jand g123(.dina(w_dff_B_rpyFMvjf6_0),.dinb(n161),.dout(n166),.clk(gclk));
	jand g124(.dina(n166),.dinb(w_dff_B_NkP5lfii7_1),.dout(n167),.clk(gclk));
	jnot g125(.din(w_n120_0[0]),.dout(n168),.clk(gclk));
	jand g126(.dina(w_G223gat_2[1]),.dinb(w_G76gat_0[0]),.dout(n169),.clk(gclk));
	jor g127(.dina(n169),.dinb(w_n88_0[0]),.dout(n170),.clk(gclk));
	jor g128(.dina(w_n170_0[1]),.dinb(w_G86gat_0[1]),.dout(n171),.clk(gclk));
	jand g129(.dina(w_G223gat_2[0]),.dinb(w_G1gat_0[0]),.dout(n172),.clk(gclk));
	jor g130(.dina(n172),.dinb(w_n84_0[0]),.dout(n173),.clk(gclk));
	jor g131(.dina(w_n173_0[1]),.dinb(w_G8gat_0[1]),.dout(n174),.clk(gclk));
	jand g132(.dina(w_G223gat_1[2]),.dinb(w_n46_0[0]),.dout(n175),.clk(gclk));
	jor g133(.dina(n175),.dinb(w_n45_0[0]),.dout(n176),.clk(gclk));
	jor g134(.dina(n176),.dinb(w_G47gat_0[0]),.dout(n177),.clk(gclk));
	jand g135(.dina(n177),.dinb(n174),.dout(n178),.clk(gclk));
	jand g136(.dina(n178),.dinb(w_dff_B_MGjLvvx48_1),.dout(n179),.clk(gclk));
	jand g137(.dina(n179),.dinb(w_dff_B_NQ6qWZcn7_1),.dout(n180),.clk(gclk));
	jand g138(.dina(n180),.dinb(n167),.dout(n181),.clk(gclk));
	jor g139(.dina(w_n181_2[2]),.dinb(w_n106_0[0]),.dout(n182),.clk(gclk));
	jand g140(.dina(n182),.dinb(w_n108_0[0]),.dout(n183),.clk(gclk));
	jand g141(.dina(w_n183_0[1]),.dinb(w_n149_0[1]),.dout(n184),.clk(gclk));
	jnot g142(.din(w_G66gat_0[2]),.dout(n185),.clk(gclk));
	jor g143(.dina(w_n181_2[1]),.dinb(w_n117_0[0]),.dout(n186),.clk(gclk));
	jand g144(.dina(n186),.dinb(w_n119_0[1]),.dout(n187),.clk(gclk));
	jand g145(.dina(n187),.dinb(w_n185_0[1]),.dout(n188),.clk(gclk));
	jor g146(.dina(n188),.dinb(n184),.dout(n189),.clk(gclk));
	jnot g147(.din(w_G14gat_0[2]),.dout(n190),.clk(gclk));
	jor g148(.dina(w_n181_2[0]),.dinb(w_n125_0[0]),.dout(n191),.clk(gclk));
	jand g149(.dina(n191),.dinb(w_n127_0[0]),.dout(n192),.clk(gclk));
	jand g150(.dina(n192),.dinb(w_dff_B_PlDjCZY22_1),.dout(n193),.clk(gclk));
	jnot g151(.din(w_G92gat_0[2]),.dout(n194),.clk(gclk));
	jor g152(.dina(w_n181_1[2]),.dinb(w_n121_0[0]),.dout(n195),.clk(gclk));
	jand g153(.dina(n195),.dinb(w_n123_0[0]),.dout(n196),.clk(gclk));
	jand g154(.dina(n196),.dinb(w_dff_B_XRoBwbH59_1),.dout(n197),.clk(gclk));
	jor g155(.dina(n197),.dinb(n193),.dout(n198),.clk(gclk));
	jor g156(.dina(n198),.dinb(n189),.dout(n199),.clk(gclk));
	jnot g157(.din(w_G79gat_0[1]),.dout(n200),.clk(gclk));
	jor g158(.dina(w_n181_1[1]),.dinb(w_n102_0[0]),.dout(n201),.clk(gclk));
	jand g159(.dina(n201),.dinb(w_n104_0[0]),.dout(n202),.clk(gclk));
	jand g160(.dina(w_n202_0[1]),.dinb(w_n200_0[1]),.dout(n203),.clk(gclk));
	jnot g161(.din(w_G115gat_0[1]),.dout(n204),.clk(gclk));
	jor g162(.dina(w_n181_1[0]),.dinb(w_n111_0[0]),.dout(n205),.clk(gclk));
	jand g163(.dina(n205),.dinb(w_n113_0[0]),.dout(n206),.clk(gclk));
	jand g164(.dina(w_n206_0[1]),.dinb(w_n204_0[1]),.dout(n207),.clk(gclk));
	jor g165(.dina(n207),.dinb(n203),.dout(n208),.clk(gclk));
	jnot g166(.din(w_G27gat_0[1]),.dout(n209),.clk(gclk));
	jor g167(.dina(w_n181_0[2]),.dinb(w_n70_0[0]),.dout(n210),.clk(gclk));
	jand g168(.dina(n210),.dinb(w_n95_0[0]),.dout(n211),.clk(gclk));
	jand g169(.dina(w_n211_0[1]),.dinb(w_n209_0[1]),.dout(n212),.clk(gclk));
	jor g170(.dina(w_dff_B_esJ086AR6_0),.dinb(n208),.dout(n213),.clk(gclk));
	jor g171(.dina(n213),.dinb(n199),.dout(n214),.clk(gclk));
	jor g172(.dina(n214),.dinb(w_dff_B_K8XvReoO8_1),.dout(G370gat_fa_),.clk(gclk));
	jnot g173(.din(w_n147_0[0]),.dout(n216),.clk(gclk));
	jand g174(.dina(n216),.dinb(w_n141_0[0]),.dout(n217),.clk(gclk));
	jand g175(.dina(w_G329gat_3[1]),.dinb(w_G34gat_0[0]),.dout(n218),.clk(gclk));
	jor g176(.dina(n218),.dinb(w_n159_0[0]),.dout(n219),.clk(gclk));
	jor g177(.dina(n219),.dinb(w_G40gat_0[0]),.dout(n220),.clk(gclk));
	jnot g178(.din(w_n119_0[0]),.dout(n221),.clk(gclk));
	jand g179(.dina(w_G329gat_3[0]),.dinb(w_G60gat_0[0]),.dout(n222),.clk(gclk));
	jor g180(.dina(w_n222_0[1]),.dinb(w_dff_B_NyDAsDHa5_1),.dout(n223),.clk(gclk));
	jor g181(.dina(n223),.dinb(w_G66gat_0[1]),.dout(n224),.clk(gclk));
	jand g182(.dina(n224),.dinb(n220),.dout(n225),.clk(gclk));
	jand g183(.dina(w_G329gat_2[2]),.dinb(w_G8gat_0[0]),.dout(n226),.clk(gclk));
	jor g184(.dina(n226),.dinb(w_n173_0[0]),.dout(n227),.clk(gclk));
	jor g185(.dina(w_n227_0[1]),.dinb(w_G14gat_0[1]),.dout(n228),.clk(gclk));
	jand g186(.dina(w_G329gat_2[1]),.dinb(w_G86gat_0[0]),.dout(n229),.clk(gclk));
	jor g187(.dina(n229),.dinb(w_n170_0[0]),.dout(n230),.clk(gclk));
	jor g188(.dina(w_n230_0[1]),.dinb(w_G92gat_0[1]),.dout(n231),.clk(gclk));
	jand g189(.dina(n231),.dinb(n228),.dout(n232),.clk(gclk));
	jand g190(.dina(n232),.dinb(n225),.dout(n233),.clk(gclk));
	jand g191(.dina(w_G329gat_2[0]),.dinb(w_G73gat_0[0]),.dout(n234),.clk(gclk));
	jor g192(.dina(n234),.dinb(w_n156_0[0]),.dout(n235),.clk(gclk));
	jor g193(.dina(n235),.dinb(w_G79gat_0[0]),.dout(n236),.clk(gclk));
	jand g194(.dina(w_G329gat_1[2]),.dinb(w_G112gat_0[0]),.dout(n237),.clk(gclk));
	jor g195(.dina(n237),.dinb(w_n164_0[0]),.dout(n238),.clk(gclk));
	jor g196(.dina(n238),.dinb(w_G115gat_0[0]),.dout(n239),.clk(gclk));
	jand g197(.dina(n239),.dinb(n236),.dout(n240),.clk(gclk));
	jand g198(.dina(w_G329gat_1[1]),.dinb(w_G21gat_0[0]),.dout(n241),.clk(gclk));
	jor g199(.dina(n241),.dinb(w_n151_0[0]),.dout(n242),.clk(gclk));
	jor g200(.dina(n242),.dinb(w_G27gat_0[0]),.dout(n243),.clk(gclk));
	jand g201(.dina(w_dff_B_zJt6HAym3_0),.dinb(n240),.dout(n244),.clk(gclk));
	jand g202(.dina(n244),.dinb(n233),.dout(n245),.clk(gclk));
	jand g203(.dina(n245),.dinb(w_dff_B_ZhxoKhHD8_1),.dout(n246),.clk(gclk));
	jor g204(.dina(w_n246_2[2]),.dinb(w_n209_0[0]),.dout(n247),.clk(gclk));
	jand g205(.dina(n247),.dinb(w_n211_0[0]),.dout(n248),.clk(gclk));
	jor g206(.dina(w_n246_2[1]),.dinb(w_n149_0[0]),.dout(n249),.clk(gclk));
	jand g207(.dina(n249),.dinb(w_n183_0[0]),.dout(n250),.clk(gclk));
	jor g208(.dina(w_n250_0[1]),.dinb(w_n248_0[1]),.dout(n251),.clk(gclk));
	jor g209(.dina(w_n246_2[0]),.dinb(w_n145_0[0]),.dout(n252),.clk(gclk));
	jand g210(.dina(w_n144_0[0]),.dinb(w_n131_0[0]),.dout(n253),.clk(gclk));
	jand g211(.dina(w_n253_0[1]),.dinb(n252),.dout(n254),.clk(gclk));
	jor g212(.dina(w_n246_1[2]),.dinb(w_n185_0[0]),.dout(n255),.clk(gclk));
	jand g213(.dina(w_G223gat_1[1]),.dinb(w_n81_0[0]),.dout(n256),.clk(gclk));
	jor g214(.dina(w_n222_0[0]),.dinb(w_dff_B_3iyEOD4r6_1),.dout(n257),.clk(gclk));
	jnot g215(.din(w_n257_0[1]),.dout(n258),.clk(gclk));
	jand g216(.dina(w_dff_B_8uzFWmwk8_0),.dinb(n255),.dout(n259),.clk(gclk));
	jand g217(.dina(n259),.dinb(w_G56gat_0[1]),.dout(n260),.clk(gclk));
	jor g218(.dina(n260),.dinb(w_n254_0[1]),.dout(n261),.clk(gclk));
	jor g219(.dina(n261),.dinb(w_n251_0[1]),.dout(G430gat_fa_),.clk(gclk));
	jand g220(.dina(w_G370gat_1[1]),.dinb(w_G92gat_0[0]),.dout(n263),.clk(gclk));
	jor g221(.dina(n263),.dinb(w_n230_0[0]),.dout(n264),.clk(gclk));
	jnot g222(.din(w_n264_0[1]),.dout(n265),.clk(gclk));
	jnot g223(.din(w_n140_0[0]),.dout(n266),.clk(gclk));
	jnot g224(.din(w_G105gat_0[0]),.dout(n267),.clk(gclk));
	jor g225(.dina(w_n246_1[1]),.dinb(w_dff_B_HKO3SEqS9_1),.dout(n268),.clk(gclk));
	jand g226(.dina(n268),.dinb(w_dff_B_FgqCtSzS2_1),.dout(n269),.clk(gclk));
	jor g227(.dina(w_n246_1[0]),.dinb(w_n200_0[0]),.dout(n270),.clk(gclk));
	jand g228(.dina(n270),.dinb(w_n202_0[0]),.dout(n271),.clk(gclk));
	jor g229(.dina(w_n246_0[2]),.dinb(w_n204_0[0]),.dout(n272),.clk(gclk));
	jand g230(.dina(n272),.dinb(w_n206_0[0]),.dout(n273),.clk(gclk));
	jor g231(.dina(n273),.dinb(w_n271_0[1]),.dout(n274),.clk(gclk));
	jor g232(.dina(n274),.dinb(w_n269_0[1]),.dout(n275),.clk(gclk));
	jor g233(.dina(n275),.dinb(w_n265_0[1]),.dout(n276),.clk(gclk));
	jor g234(.dina(n276),.dinb(w_G430gat_0),.dout(n277),.clk(gclk));
	jand g235(.dina(w_G370gat_1[0]),.dinb(w_G14gat_0[0]),.dout(n278),.clk(gclk));
	jor g236(.dina(n278),.dinb(w_n227_0[0]),.dout(n279),.clk(gclk));
	jand g237(.dina(w_dff_B_79cmHCEP3_0),.dinb(n277),.dout(G421gat),.clk(gclk));
	jnot g238(.din(w_n250_0[0]),.dout(n281),.clk(gclk));
	jand g239(.dina(w_G370gat_0[2]),.dinb(w_G53gat_0[0]),.dout(n282),.clk(gclk));
	jnot g240(.din(w_n253_0[0]),.dout(n283),.clk(gclk));
	jor g241(.dina(w_dff_B_iwDUkmAt4_0),.dinb(n282),.dout(n284),.clk(gclk));
	jand g242(.dina(w_G370gat_0[1]),.dinb(w_G66gat_0[0]),.dout(n285),.clk(gclk));
	jor g243(.dina(w_n257_0[0]),.dinb(n285),.dout(n286),.clk(gclk));
	jor g244(.dina(n286),.dinb(w_n80_0[0]),.dout(n287),.clk(gclk));
	jand g245(.dina(n287),.dinb(w_dff_B_eJEne66E0_1),.dout(n288),.clk(gclk));
	jand g246(.dina(w_n288_0[1]),.dinb(w_n281_0[1]),.dout(n289),.clk(gclk));
	jand g247(.dina(n289),.dinb(w_n271_0[0]),.dout(n290),.clk(gclk));
	jand g248(.dina(w_n265_0[0]),.dinb(w_n288_0[0]),.dout(n291),.clk(gclk));
	jor g249(.dina(n291),.dinb(w_n251_0[0]),.dout(n292),.clk(gclk));
	jor g250(.dina(n292),.dinb(w_n290_0[1]),.dout(G431gat),.clk(gclk));
	jand g251(.dina(w_n269_0[0]),.dinb(w_n264_0[0]),.dout(n294),.clk(gclk));
	jor g252(.dina(n294),.dinb(w_n254_0[0]),.dout(n295),.clk(gclk));
	jand g253(.dina(n295),.dinb(w_n281_0[0]),.dout(n296),.clk(gclk));
	jor g254(.dina(n296),.dinb(w_n248_0[0]),.dout(n297),.clk(gclk));
	jor g255(.dina(n297),.dinb(w_n290_0[0]),.dout(G432gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_9feHHqEP9_0),.doutb(w_dff_A_ZUmlp4ih2_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_dff_A_u2Wkcub51_0),.doutb(w_G4gat_0[1]),.doutc(w_dff_A_CPVaA3YE2_2),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_Le75QP4r4_0),.doutb(w_dff_A_tttNuUrm6_1),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G11gat_0(.douta(w_dff_A_X0lqFf1U5_0),.doutb(w_dff_A_asY2EJUK6_1),.doutc(w_G11gat_0[2]),.din(G11gat));
	jspl3 jspl3_w_G14gat_0(.douta(w_dff_A_X7CJlDZg1_0),.doutb(w_dff_A_zfRanZFb5_1),.doutc(w_G14gat_0[2]),.din(G14gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_dff_A_KATBrZG45_0),.doutb(w_G17gat_0[1]),.doutc(w_dff_A_2GQp74W96_2),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_dff_A_9ygUFtzK9_0),.doutb(w_dff_A_2UsyUsik1_1),.doutc(w_G21gat_0[2]),.din(G21gat));
	jspl3 jspl3_w_G24gat_0(.douta(w_dff_A_w7lt1dcp9_0),.doutb(w_dff_A_AuOKD7660_1),.doutc(w_G24gat_0[2]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_dff_A_mAgQsyME8_0),.doutb(w_G27gat_0[1]),.din(G27gat));
	jspl3 jspl3_w_G30gat_0(.douta(w_dff_A_TclB1t9Z4_0),.doutb(w_G30gat_0[1]),.doutc(w_dff_A_GkEWWy088_2),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_dff_A_qZdLlFXE3_0),.doutb(w_dff_A_z7fBMfWI3_1),.doutc(w_G34gat_0[2]),.din(G34gat));
	jspl jspl_w_G40gat_0(.douta(w_dff_A_KwV5G41l5_0),.doutb(w_G40gat_0[1]),.din(G40gat));
	jspl jspl_w_G43gat_0(.douta(w_dff_A_MieW2VVm4_0),.doutb(w_G43gat_0[1]),.din(G43gat));
	jspl3 jspl3_w_G47gat_0(.douta(w_dff_A_6LwEWqdP7_0),.doutb(w_dff_A_JLloTRJ83_1),.doutc(w_G47gat_0[2]),.din(G47gat));
	jspl jspl_w_G50gat_0(.douta(w_dff_A_sns6gJAF5_0),.doutb(w_G50gat_0[1]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_dff_A_rA6U099P1_0),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_G56gat_0[0]),.doutb(w_dff_A_t52nroUK4_1),.doutc(w_dff_A_HM7Xt9M00_2),.din(G56gat));
	jspl jspl_w_G56gat_1(.douta(w_G56gat_1[0]),.doutb(w_dff_A_dZOlZMLW4_1),.din(w_G56gat_0[0]));
	jspl jspl_w_G60gat_0(.douta(w_dff_A_Eb5WXesu6_0),.doutb(w_G60gat_0[1]),.din(G60gat));
	jspl3 jspl3_w_G63gat_0(.douta(w_dff_A_usOypx327_0),.doutb(w_dff_A_zdoTkP3m3_1),.doutc(w_G63gat_0[2]),.din(G63gat));
	jspl3 jspl3_w_G66gat_0(.douta(w_dff_A_pw1kHjUz2_0),.doutb(w_dff_A_EGfukxDR9_1),.doutc(w_G66gat_0[2]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_dff_A_7wRvwOcp8_0),.doutb(w_G69gat_0[1]),.doutc(w_dff_A_CDaLzzUH4_2),.din(G69gat));
	jspl3 jspl3_w_G73gat_0(.douta(w_dff_A_YZreO8RO2_0),.doutb(w_dff_A_EE1vAm416_1),.doutc(w_G73gat_0[2]),.din(G73gat));
	jspl3 jspl3_w_G76gat_0(.douta(w_dff_A_9dUrKNKd3_0),.doutb(w_dff_A_0ivgQ7UW7_1),.doutc(w_G76gat_0[2]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_dff_A_PkvW4NuJ6_0),.doutb(w_G79gat_0[1]),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_dff_A_NE6oXFhM3_0),.doutb(w_G82gat_0[1]),.doutc(w_dff_A_jCLSgv0p3_2),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_dff_A_8NTOvryK9_0),.doutb(w_dff_A_4RTxeQTv8_1),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G89gat_0(.douta(w_dff_A_lKn6yJlJ6_0),.doutb(w_dff_A_TRRJesDS2_1),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_FEf1B7nZ7_0),.doutb(w_dff_A_PWYb19Y21_1),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_dff_A_1s5F0kqf1_0),.doutb(w_G95gat_0[1]),.doutc(w_dff_A_m3tq5pOZ7_2),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_EV2WFCl09_0),.doutb(w_dff_A_xwKVzm7V8_1),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl jspl_w_G102gat_0(.douta(w_dff_A_70y3XZk07_0),.doutb(w_G102gat_0[1]),.din(G102gat));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_dff_A_UzWk0GRm9_1),.din(G105gat));
	jspl3 jspl3_w_G108gat_0(.douta(w_G108gat_0[0]),.doutb(w_dff_A_W3svUPV46_1),.doutc(w_dff_A_4i46PGmI0_2),.din(G108gat));
	jspl3 jspl3_w_G112gat_0(.douta(w_dff_A_IGg9SyEP8_0),.doutb(w_dff_A_Go6c1lDV5_1),.doutc(w_G112gat_0[2]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_dff_A_HRDrLIPA2_0),.doutb(w_G115gat_0[1]),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(w_G223gat_3[2]),.din(w_G223gat_0[2]));
	jspl jspl_w_G223gat_4(.douta(w_G223gat_4),.doutb(w_dff_A_SEMGl6Zg8_1),.din(w_G223gat_1[0]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl jspl_w_G329gat_4(.douta(w_G329gat_4),.doutb(w_dff_A_n8EDLT5F7_1),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_dff_A_yBeS5tNQ7_2),.din(w_G370gat_0[0]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(w_dff_A_azFe6ujw4_1),.din(G430gat_fa_));
	jspl jspl_w_n43_0(.douta(w_dff_A_YwwioSY85_0),.doutb(w_n43_0[1]),.din(n43));
	jspl jspl_w_n44_0(.douta(w_n44_0[0]),.doutb(w_dff_A_ebpXr9Hh7_1),.din(n44));
	jspl jspl_w_n45_0(.douta(w_dff_A_q6JCB2dB3_0),.doutb(w_n45_0[1]),.din(n45));
	jspl3 jspl3_w_n46_0(.douta(w_dff_A_B7Epgujb4_0),.doutb(w_dff_A_ywAkzHm66_1),.doutc(w_n46_0[2]),.din(n46));
	jspl jspl_w_n47_0(.douta(w_dff_A_nhp2kmJQ0_0),.doutb(w_n47_0[1]),.din(n47));
	jspl jspl_w_n49_0(.douta(w_dff_A_zUzEfCVk4_0),.doutb(w_n49_0[1]),.din(n49));
	jspl jspl_w_n51_0(.douta(w_dff_A_EODEH6fW7_0),.doutb(w_n51_0[1]),.din(n51));
	jspl jspl_w_n54_0(.douta(w_dff_A_2sB8qnBj9_0),.doutb(w_n54_0[1]),.din(n54));
	jspl jspl_w_n57_0(.douta(w_dff_A_rlN0UfkF4_0),.doutb(w_n57_0[1]),.din(n57));
	jspl jspl_w_n60_0(.douta(w_dff_A_9mFFV7fQ3_0),.doutb(w_n60_0[1]),.din(n60));
	jspl jspl_w_n62_0(.douta(w_dff_A_fk6MrzLy9_0),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n64_0(.douta(w_dff_A_kSn583jH5_0),.doutb(w_n64_0[1]),.din(n64));
	jspl jspl_w_n70_0(.douta(w_dff_A_dM4HeqPw5_0),.doutb(w_n70_0[1]),.din(w_dff_B_du5n4KHy9_2));
	jspl jspl_w_n73_0(.douta(w_dff_A_DfSg4lqe1_0),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n75_0(.douta(w_dff_A_jCXMQBrh3_0),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n78_0(.douta(w_dff_A_4tjV6s9y4_0),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n80_0(.douta(w_dff_A_KULj1DkY4_0),.doutb(w_n80_0[1]),.din(n80));
	jspl jspl_w_n81_0(.douta(w_dff_A_QWq5YH7x7_0),.doutb(w_n81_0[1]),.din(n81));
	jspl jspl_w_n84_0(.douta(w_dff_A_gGNBgYqU5_0),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_dff_A_VfX4Xf9w3_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_dff_A_kwJpDK9d3_0),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl3 jspl3_w_n93_1(.douta(w_n93_1[0]),.doutb(w_n93_1[1]),.doutc(w_n93_1[2]),.din(w_n93_0[0]));
	jspl3 jspl3_w_n93_2(.douta(w_n93_2[0]),.doutb(w_n93_2[1]),.doutc(w_n93_2[2]),.din(w_n93_0[1]));
	jspl3 jspl3_w_n93_3(.douta(w_n93_3[0]),.doutb(w_n93_3[1]),.doutc(w_n93_3[2]),.din(w_n93_0[2]));
	jspl jspl_w_n95_0(.douta(w_dff_A_cRMZYc3B1_0),.doutb(w_n95_0[1]),.din(n95));
	jspl jspl_w_n102_0(.douta(w_dff_A_xQEWaPFd4_0),.doutb(w_n102_0[1]),.din(w_dff_B_IF04gzgP6_2));
	jspl jspl_w_n104_0(.douta(w_dff_A_zUsGRMpU8_0),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n106_0(.douta(w_dff_A_V88cwFC23_0),.doutb(w_n106_0[1]),.din(w_dff_B_93DoIoKW3_2));
	jspl jspl_w_n108_0(.douta(w_dff_A_XMNTUH095_0),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n111_0(.douta(w_dff_A_mLXAvt4n0_0),.doutb(w_n111_0[1]),.din(w_dff_B_kRvHPEm09_2));
	jspl jspl_w_n113_0(.douta(w_dff_A_jvJV2ZFZ2_0),.doutb(w_n113_0[1]),.din(n113));
	jspl jspl_w_n117_0(.douta(w_dff_A_i5tkwe6P9_0),.doutb(w_n117_0[1]),.din(w_dff_B_A00qhiij1_2));
	jspl3 jspl3_w_n119_0(.douta(w_n119_0[0]),.doutb(w_dff_A_us47lpq66_1),.doutc(w_n119_0[2]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_dff_A_G9lrbznW0_1),.din(n120));
	jspl jspl_w_n121_0(.douta(w_dff_A_TNwq3u6B6_0),.doutb(w_n121_0[1]),.din(w_dff_B_aWMZslLJ7_2));
	jspl jspl_w_n123_0(.douta(w_dff_A_yXhG2H8g8_0),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n125_0(.douta(w_dff_A_sOSeQPg69_0),.doutb(w_n125_0[1]),.din(w_dff_B_jlkyKIwC3_2));
	jspl jspl_w_n127_0(.douta(w_dff_A_j1MTcUuX6_0),.doutb(w_n127_0[1]),.din(n127));
	jspl3 jspl3_w_n131_0(.douta(w_dff_A_fnI5mclx4_0),.doutb(w_n131_0[1]),.doutc(w_n131_0[2]),.din(n131));
	jspl jspl_w_n138_0(.douta(w_n138_0[0]),.doutb(w_dff_A_GzJpBzPy9_1),.din(n138));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n141_0(.douta(w_dff_A_iZIDpyIr3_0),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(n144));
	jspl jspl_w_n145_0(.douta(w_dff_A_MDnOkpYB1_0),.doutb(w_n145_0[1]),.din(w_dff_B_1M8i8mw79_2));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_dff_A_XQDfzSS13_1),.din(n147));
	jspl jspl_w_n149_0(.douta(w_dff_A_xnsN78VT8_0),.doutb(w_n149_0[1]),.din(w_dff_B_jl8Wcy995_2));
	jspl jspl_w_n151_0(.douta(w_dff_A_YjxOWqGe8_0),.doutb(w_n151_0[1]),.din(n151));
	jspl jspl_w_n156_0(.douta(w_dff_A_sKncualL7_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n159_0(.douta(w_dff_A_LLFs3lMj2_0),.doutb(w_n159_0[1]),.din(n159));
	jspl jspl_w_n164_0(.douta(w_dff_A_4GiB9DAe3_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n170_0(.douta(w_dff_A_HOZpH2xk1_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n173_0(.douta(w_dff_A_Z6xDi7py5_0),.doutb(w_n173_0[1]),.din(n173));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n181_2(.douta(w_n181_2[0]),.doutb(w_n181_2[1]),.doutc(w_n181_2[2]),.din(w_n181_0[1]));
	jspl jspl_w_n183_0(.douta(w_dff_A_8Dmcj8nY2_0),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n185_0(.douta(w_dff_A_zvdmaR5U2_0),.doutb(w_n185_0[1]),.din(w_dff_B_y54Z7sHy7_2));
	jspl jspl_w_n200_0(.douta(w_dff_A_UkbINEYs0_0),.doutb(w_n200_0[1]),.din(w_dff_B_jWf3GUkZ9_2));
	jspl jspl_w_n202_0(.douta(w_dff_A_4ovGi05V3_0),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n204_0(.douta(w_dff_A_seRwWBH32_0),.doutb(w_n204_0[1]),.din(w_dff_B_JHCPCgkZ6_2));
	jspl jspl_w_n206_0(.douta(w_dff_A_dbQqSDnz1_0),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n209_0(.douta(w_dff_A_qGfc80q32_0),.doutb(w_n209_0[1]),.din(w_dff_B_bgzYbinz7_2));
	jspl jspl_w_n211_0(.douta(w_dff_A_MtDsypUi6_0),.doutb(w_n211_0[1]),.din(n211));
	jspl jspl_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n227_0(.douta(w_dff_A_l6vhJiZM3_0),.doutb(w_n227_0[1]),.din(n227));
	jspl jspl_w_n230_0(.douta(w_dff_A_4hKeouNQ8_0),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl3 jspl3_w_n246_1(.douta(w_n246_1[0]),.doutb(w_n246_1[1]),.doutc(w_n246_1[2]),.din(w_n246_0[0]));
	jspl3 jspl3_w_n246_2(.douta(w_n246_2[0]),.doutb(w_n246_2[1]),.doutc(w_n246_2[2]),.din(w_n246_0[1]));
	jspl jspl_w_n248_0(.douta(w_dff_A_svtpdesh5_0),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_dff_A_ePfqqCRY9_0),.doutb(w_n251_0[1]),.din(w_dff_B_RfiQmJcF3_2));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_dff_A_e9JMKHNp3_1),.din(n253));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(w_dff_B_uui4NYYm0_2));
	jspl jspl_w_n257_0(.douta(w_dff_A_cQsYk8by8_0),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(w_dff_B_r4O0bDM98_2));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_dff_A_V53s9Bud7_1),.din(n269));
	jspl jspl_w_n271_0(.douta(w_dff_A_frZW8Ixb0_0),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.din(w_dff_B_oiWBOB7h9_2));
	jspl jspl_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.din(n288));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(n290));
	jdff dff_B_vwebLdyM5_0(.din(n279),.dout(w_dff_B_vwebLdyM5_0),.clk(gclk));
	jdff dff_B_oLBFTUv28_0(.din(w_dff_B_vwebLdyM5_0),.dout(w_dff_B_oLBFTUv28_0),.clk(gclk));
	jdff dff_B_SoG1fvF07_0(.din(w_dff_B_oLBFTUv28_0),.dout(w_dff_B_SoG1fvF07_0),.clk(gclk));
	jdff dff_B_79cmHCEP3_0(.din(w_dff_B_SoG1fvF07_0),.dout(w_dff_B_79cmHCEP3_0),.clk(gclk));
	jdff dff_B_wCIJXmYt4_0(.din(n258),.dout(w_dff_B_wCIJXmYt4_0),.clk(gclk));
	jdff dff_B_qxQuhH704_0(.din(w_dff_B_wCIJXmYt4_0),.dout(w_dff_B_qxQuhH704_0),.clk(gclk));
	jdff dff_B_gUf4KBF24_0(.din(w_dff_B_qxQuhH704_0),.dout(w_dff_B_gUf4KBF24_0),.clk(gclk));
	jdff dff_B_3oNaz6UP6_0(.din(w_dff_B_gUf4KBF24_0),.dout(w_dff_B_3oNaz6UP6_0),.clk(gclk));
	jdff dff_B_8uzFWmwk8_0(.din(w_dff_B_3oNaz6UP6_0),.dout(w_dff_B_8uzFWmwk8_0),.clk(gclk));
	jdff dff_B_r4O0bDM98_2(.din(n265),.dout(w_dff_B_r4O0bDM98_2),.clk(gclk));
	jdff dff_A_ePfqqCRY9_0(.dout(w_n251_0[0]),.din(w_dff_A_ePfqqCRY9_0),.clk(gclk));
	jdff dff_B_RfiQmJcF3_2(.din(n251),.dout(w_dff_B_RfiQmJcF3_2),.clk(gclk));
	jdff dff_A_V53s9Bud7_1(.dout(w_n269_0[1]),.din(w_dff_A_V53s9Bud7_1),.clk(gclk));
	jdff dff_B_43yBtcuU3_1(.din(n266),.dout(w_dff_B_43yBtcuU3_1),.clk(gclk));
	jdff dff_B_KVHQTPUU2_1(.din(w_dff_B_43yBtcuU3_1),.dout(w_dff_B_KVHQTPUU2_1),.clk(gclk));
	jdff dff_B_tOvj13OK4_1(.din(w_dff_B_KVHQTPUU2_1),.dout(w_dff_B_tOvj13OK4_1),.clk(gclk));
	jdff dff_B_qrDAUZOZ2_1(.din(w_dff_B_tOvj13OK4_1),.dout(w_dff_B_qrDAUZOZ2_1),.clk(gclk));
	jdff dff_B_FgqCtSzS2_1(.din(w_dff_B_qrDAUZOZ2_1),.dout(w_dff_B_FgqCtSzS2_1),.clk(gclk));
	jdff dff_B_KOSLGNRT6_1(.din(n267),.dout(w_dff_B_KOSLGNRT6_1),.clk(gclk));
	jdff dff_B_LmmiM9Xv9_1(.din(w_dff_B_KOSLGNRT6_1),.dout(w_dff_B_LmmiM9Xv9_1),.clk(gclk));
	jdff dff_B_LfGHjFt56_1(.din(w_dff_B_LmmiM9Xv9_1),.dout(w_dff_B_LfGHjFt56_1),.clk(gclk));
	jdff dff_B_CPy1CaQU2_1(.din(w_dff_B_LfGHjFt56_1),.dout(w_dff_B_CPy1CaQU2_1),.clk(gclk));
	jdff dff_B_25uQAo1M0_1(.din(w_dff_B_CPy1CaQU2_1),.dout(w_dff_B_25uQAo1M0_1),.clk(gclk));
	jdff dff_B_hSBrOcX19_1(.din(w_dff_B_25uQAo1M0_1),.dout(w_dff_B_hSBrOcX19_1),.clk(gclk));
	jdff dff_B_E0fz8Fo44_1(.din(w_dff_B_hSBrOcX19_1),.dout(w_dff_B_E0fz8Fo44_1),.clk(gclk));
	jdff dff_B_cMRFAcil9_1(.din(w_dff_B_E0fz8Fo44_1),.dout(w_dff_B_cMRFAcil9_1),.clk(gclk));
	jdff dff_B_WnVUmdgl8_1(.din(w_dff_B_cMRFAcil9_1),.dout(w_dff_B_WnVUmdgl8_1),.clk(gclk));
	jdff dff_B_wwQQdLiQ3_1(.din(w_dff_B_WnVUmdgl8_1),.dout(w_dff_B_wwQQdLiQ3_1),.clk(gclk));
	jdff dff_B_yN1SrVII7_1(.din(w_dff_B_wwQQdLiQ3_1),.dout(w_dff_B_yN1SrVII7_1),.clk(gclk));
	jdff dff_B_O01IHSQm2_1(.din(w_dff_B_yN1SrVII7_1),.dout(w_dff_B_O01IHSQm2_1),.clk(gclk));
	jdff dff_B_szApWXCv5_1(.din(w_dff_B_O01IHSQm2_1),.dout(w_dff_B_szApWXCv5_1),.clk(gclk));
	jdff dff_B_pOZNkinj4_1(.din(w_dff_B_szApWXCv5_1),.dout(w_dff_B_pOZNkinj4_1),.clk(gclk));
	jdff dff_B_zQrb1Bal0_1(.din(w_dff_B_pOZNkinj4_1),.dout(w_dff_B_zQrb1Bal0_1),.clk(gclk));
	jdff dff_B_ODz5wPXy6_1(.din(w_dff_B_zQrb1Bal0_1),.dout(w_dff_B_ODz5wPXy6_1),.clk(gclk));
	jdff dff_B_4KOH86ug3_1(.din(w_dff_B_ODz5wPXy6_1),.dout(w_dff_B_4KOH86ug3_1),.clk(gclk));
	jdff dff_B_CN6R47Uy5_1(.din(w_dff_B_4KOH86ug3_1),.dout(w_dff_B_CN6R47Uy5_1),.clk(gclk));
	jdff dff_B_HKO3SEqS9_1(.din(w_dff_B_CN6R47Uy5_1),.dout(w_dff_B_HKO3SEqS9_1),.clk(gclk));
	jdff dff_B_uui4NYYm0_2(.din(n254),.dout(w_dff_B_uui4NYYm0_2),.clk(gclk));
	jdff dff_A_XDeI3lnr5_0(.dout(w_n248_0[0]),.din(w_dff_A_XDeI3lnr5_0),.clk(gclk));
	jdff dff_A_e9DjkIqI4_0(.dout(w_dff_A_XDeI3lnr5_0),.din(w_dff_A_e9DjkIqI4_0),.clk(gclk));
	jdff dff_A_svtpdesh5_0(.dout(w_dff_A_e9DjkIqI4_0),.din(w_dff_A_svtpdesh5_0),.clk(gclk));
	jdff dff_B_eJEne66E0_1(.din(n284),.dout(w_dff_B_eJEne66E0_1),.clk(gclk));
	jdff dff_A_GZGs2fVn7_0(.dout(w_n257_0[0]),.din(w_dff_A_GZGs2fVn7_0),.clk(gclk));
	jdff dff_A_6UT3alEb7_0(.dout(w_dff_A_GZGs2fVn7_0),.din(w_dff_A_6UT3alEb7_0),.clk(gclk));
	jdff dff_A_ssRhug4y7_0(.dout(w_dff_A_6UT3alEb7_0),.din(w_dff_A_ssRhug4y7_0),.clk(gclk));
	jdff dff_A_2GaXWSBg2_0(.dout(w_dff_A_ssRhug4y7_0),.din(w_dff_A_2GaXWSBg2_0),.clk(gclk));
	jdff dff_A_cVOe3GPp0_0(.dout(w_dff_A_2GaXWSBg2_0),.din(w_dff_A_cVOe3GPp0_0),.clk(gclk));
	jdff dff_A_cQsYk8by8_0(.dout(w_dff_A_cVOe3GPp0_0),.din(w_dff_A_cQsYk8by8_0),.clk(gclk));
	jdff dff_B_d4byrfUW0_1(.din(n256),.dout(w_dff_B_d4byrfUW0_1),.clk(gclk));
	jdff dff_B_38Cgd16t7_1(.din(w_dff_B_d4byrfUW0_1),.dout(w_dff_B_38Cgd16t7_1),.clk(gclk));
	jdff dff_B_JDh6NcOG2_1(.din(w_dff_B_38Cgd16t7_1),.dout(w_dff_B_JDh6NcOG2_1),.clk(gclk));
	jdff dff_B_PCjPAHOB3_1(.din(w_dff_B_JDh6NcOG2_1),.dout(w_dff_B_PCjPAHOB3_1),.clk(gclk));
	jdff dff_B_PLk0RNOm6_1(.din(w_dff_B_PCjPAHOB3_1),.dout(w_dff_B_PLk0RNOm6_1),.clk(gclk));
	jdff dff_B_6Urc5rC95_1(.din(w_dff_B_PLk0RNOm6_1),.dout(w_dff_B_6Urc5rC95_1),.clk(gclk));
	jdff dff_B_3iyEOD4r6_1(.din(w_dff_B_6Urc5rC95_1),.dout(w_dff_B_3iyEOD4r6_1),.clk(gclk));
	jdff dff_B_E92dO7Rk5_0(.din(n283),.dout(w_dff_B_E92dO7Rk5_0),.clk(gclk));
	jdff dff_B_iO0msDPq8_0(.din(w_dff_B_E92dO7Rk5_0),.dout(w_dff_B_iO0msDPq8_0),.clk(gclk));
	jdff dff_B_vuu4jUCe9_0(.din(w_dff_B_iO0msDPq8_0),.dout(w_dff_B_vuu4jUCe9_0),.clk(gclk));
	jdff dff_B_iwDUkmAt4_0(.din(w_dff_B_vuu4jUCe9_0),.dout(w_dff_B_iwDUkmAt4_0),.clk(gclk));
	jdff dff_A_bwA1ag0Z4_1(.dout(w_n253_0[1]),.din(w_dff_A_bwA1ag0Z4_1),.clk(gclk));
	jdff dff_A_KlHbBqMD0_1(.dout(w_dff_A_bwA1ag0Z4_1),.din(w_dff_A_KlHbBqMD0_1),.clk(gclk));
	jdff dff_A_OITiqYk01_1(.dout(w_dff_A_KlHbBqMD0_1),.din(w_dff_A_OITiqYk01_1),.clk(gclk));
	jdff dff_A_75VzJehO6_1(.dout(w_dff_A_OITiqYk01_1),.din(w_dff_A_75VzJehO6_1),.clk(gclk));
	jdff dff_A_e9JMKHNp3_1(.dout(w_dff_A_75VzJehO6_1),.din(w_dff_A_e9JMKHNp3_1),.clk(gclk));
	jdff dff_B_K8XvReoO8_1(.din(n148),.dout(w_dff_B_K8XvReoO8_1),.clk(gclk));
	jdff dff_B_esJ086AR6_0(.din(n212),.dout(w_dff_B_esJ086AR6_0),.clk(gclk));
	jdff dff_A_IOZJOknJ8_0(.dout(w_n211_0[0]),.din(w_dff_A_IOZJOknJ8_0),.clk(gclk));
	jdff dff_A_8aKTlphy4_0(.dout(w_dff_A_IOZJOknJ8_0),.din(w_dff_A_8aKTlphy4_0),.clk(gclk));
	jdff dff_A_3fXteCz35_0(.dout(w_dff_A_8aKTlphy4_0),.din(w_dff_A_3fXteCz35_0),.clk(gclk));
	jdff dff_A_DR3j0Nzw8_0(.dout(w_dff_A_3fXteCz35_0),.din(w_dff_A_DR3j0Nzw8_0),.clk(gclk));
	jdff dff_A_ZNZawBni9_0(.dout(w_dff_A_DR3j0Nzw8_0),.din(w_dff_A_ZNZawBni9_0),.clk(gclk));
	jdff dff_A_MtDsypUi6_0(.dout(w_dff_A_ZNZawBni9_0),.din(w_dff_A_MtDsypUi6_0),.clk(gclk));
	jdff dff_A_ISmlcl4W5_0(.dout(w_n209_0[0]),.din(w_dff_A_ISmlcl4W5_0),.clk(gclk));
	jdff dff_A_QEWSt3uY8_0(.dout(w_dff_A_ISmlcl4W5_0),.din(w_dff_A_QEWSt3uY8_0),.clk(gclk));
	jdff dff_A_emJaql312_0(.dout(w_dff_A_QEWSt3uY8_0),.din(w_dff_A_emJaql312_0),.clk(gclk));
	jdff dff_A_tpC5tqD67_0(.dout(w_dff_A_emJaql312_0),.din(w_dff_A_tpC5tqD67_0),.clk(gclk));
	jdff dff_A_qGfc80q32_0(.dout(w_dff_A_tpC5tqD67_0),.din(w_dff_A_qGfc80q32_0),.clk(gclk));
	jdff dff_B_7WqDrcLp1_2(.din(n209),.dout(w_dff_B_7WqDrcLp1_2),.clk(gclk));
	jdff dff_B_9ID2y5OB1_2(.din(w_dff_B_7WqDrcLp1_2),.dout(w_dff_B_9ID2y5OB1_2),.clk(gclk));
	jdff dff_B_yfSETw2Y7_2(.din(w_dff_B_9ID2y5OB1_2),.dout(w_dff_B_yfSETw2Y7_2),.clk(gclk));
	jdff dff_B_z9yi05R28_2(.din(w_dff_B_yfSETw2Y7_2),.dout(w_dff_B_z9yi05R28_2),.clk(gclk));
	jdff dff_B_fFJEMfJy2_2(.din(w_dff_B_z9yi05R28_2),.dout(w_dff_B_fFJEMfJy2_2),.clk(gclk));
	jdff dff_B_Ri7WhaH01_2(.din(w_dff_B_fFJEMfJy2_2),.dout(w_dff_B_Ri7WhaH01_2),.clk(gclk));
	jdff dff_B_RGAJpQ5v8_2(.din(w_dff_B_Ri7WhaH01_2),.dout(w_dff_B_RGAJpQ5v8_2),.clk(gclk));
	jdff dff_B_PJRQGn585_2(.din(w_dff_B_RGAJpQ5v8_2),.dout(w_dff_B_PJRQGn585_2),.clk(gclk));
	jdff dff_B_88KCtT4B9_2(.din(w_dff_B_PJRQGn585_2),.dout(w_dff_B_88KCtT4B9_2),.clk(gclk));
	jdff dff_B_KXRq1A8e9_2(.din(w_dff_B_88KCtT4B9_2),.dout(w_dff_B_KXRq1A8e9_2),.clk(gclk));
	jdff dff_B_w7y06zHV5_2(.din(w_dff_B_KXRq1A8e9_2),.dout(w_dff_B_w7y06zHV5_2),.clk(gclk));
	jdff dff_B_BsuvV6W49_2(.din(w_dff_B_w7y06zHV5_2),.dout(w_dff_B_BsuvV6W49_2),.clk(gclk));
	jdff dff_B_ks6N9hNk0_2(.din(w_dff_B_BsuvV6W49_2),.dout(w_dff_B_ks6N9hNk0_2),.clk(gclk));
	jdff dff_B_bgzYbinz7_2(.din(w_dff_B_ks6N9hNk0_2),.dout(w_dff_B_bgzYbinz7_2),.clk(gclk));
	jdff dff_A_olLEk2cE6_0(.dout(w_n206_0[0]),.din(w_dff_A_olLEk2cE6_0),.clk(gclk));
	jdff dff_A_UbvmZKng4_0(.dout(w_dff_A_olLEk2cE6_0),.din(w_dff_A_UbvmZKng4_0),.clk(gclk));
	jdff dff_A_VRvNWvrO0_0(.dout(w_dff_A_UbvmZKng4_0),.din(w_dff_A_VRvNWvrO0_0),.clk(gclk));
	jdff dff_A_4fTmYll73_0(.dout(w_dff_A_VRvNWvrO0_0),.din(w_dff_A_4fTmYll73_0),.clk(gclk));
	jdff dff_A_OWTt24nJ5_0(.dout(w_dff_A_4fTmYll73_0),.din(w_dff_A_OWTt24nJ5_0),.clk(gclk));
	jdff dff_A_dbQqSDnz1_0(.dout(w_dff_A_OWTt24nJ5_0),.din(w_dff_A_dbQqSDnz1_0),.clk(gclk));
	jdff dff_A_RhOqGTS71_0(.dout(w_n204_0[0]),.din(w_dff_A_RhOqGTS71_0),.clk(gclk));
	jdff dff_A_Q5X4imaJ6_0(.dout(w_dff_A_RhOqGTS71_0),.din(w_dff_A_Q5X4imaJ6_0),.clk(gclk));
	jdff dff_A_kavg2DEy0_0(.dout(w_dff_A_Q5X4imaJ6_0),.din(w_dff_A_kavg2DEy0_0),.clk(gclk));
	jdff dff_A_0searHjC4_0(.dout(w_dff_A_kavg2DEy0_0),.din(w_dff_A_0searHjC4_0),.clk(gclk));
	jdff dff_A_seRwWBH32_0(.dout(w_dff_A_0searHjC4_0),.din(w_dff_A_seRwWBH32_0),.clk(gclk));
	jdff dff_B_ZgxHQ6Hk4_2(.din(n204),.dout(w_dff_B_ZgxHQ6Hk4_2),.clk(gclk));
	jdff dff_B_bzAcanZg5_2(.din(w_dff_B_ZgxHQ6Hk4_2),.dout(w_dff_B_bzAcanZg5_2),.clk(gclk));
	jdff dff_B_PA8Pnz9I4_2(.din(w_dff_B_bzAcanZg5_2),.dout(w_dff_B_PA8Pnz9I4_2),.clk(gclk));
	jdff dff_B_OGPoxPg14_2(.din(w_dff_B_PA8Pnz9I4_2),.dout(w_dff_B_OGPoxPg14_2),.clk(gclk));
	jdff dff_B_t73EmK7g8_2(.din(w_dff_B_OGPoxPg14_2),.dout(w_dff_B_t73EmK7g8_2),.clk(gclk));
	jdff dff_B_eg2rpMol3_2(.din(w_dff_B_t73EmK7g8_2),.dout(w_dff_B_eg2rpMol3_2),.clk(gclk));
	jdff dff_B_RYjBlcNS3_2(.din(w_dff_B_eg2rpMol3_2),.dout(w_dff_B_RYjBlcNS3_2),.clk(gclk));
	jdff dff_B_0GnCNoDc7_2(.din(w_dff_B_RYjBlcNS3_2),.dout(w_dff_B_0GnCNoDc7_2),.clk(gclk));
	jdff dff_B_xvkXV2VS7_2(.din(w_dff_B_0GnCNoDc7_2),.dout(w_dff_B_xvkXV2VS7_2),.clk(gclk));
	jdff dff_B_nFb1iLfC0_2(.din(w_dff_B_xvkXV2VS7_2),.dout(w_dff_B_nFb1iLfC0_2),.clk(gclk));
	jdff dff_B_JKd3r0gC1_2(.din(w_dff_B_nFb1iLfC0_2),.dout(w_dff_B_JKd3r0gC1_2),.clk(gclk));
	jdff dff_B_17S53n1d3_2(.din(w_dff_B_JKd3r0gC1_2),.dout(w_dff_B_17S53n1d3_2),.clk(gclk));
	jdff dff_B_IwNFJkjs7_2(.din(w_dff_B_17S53n1d3_2),.dout(w_dff_B_IwNFJkjs7_2),.clk(gclk));
	jdff dff_B_JHCPCgkZ6_2(.din(w_dff_B_IwNFJkjs7_2),.dout(w_dff_B_JHCPCgkZ6_2),.clk(gclk));
	jdff dff_B_GDaQqjpP7_1(.din(n194),.dout(w_dff_B_GDaQqjpP7_1),.clk(gclk));
	jdff dff_B_f2VOUnh55_1(.din(w_dff_B_GDaQqjpP7_1),.dout(w_dff_B_f2VOUnh55_1),.clk(gclk));
	jdff dff_B_LUQePqha0_1(.din(w_dff_B_f2VOUnh55_1),.dout(w_dff_B_LUQePqha0_1),.clk(gclk));
	jdff dff_B_SAF5a7wU9_1(.din(w_dff_B_LUQePqha0_1),.dout(w_dff_B_SAF5a7wU9_1),.clk(gclk));
	jdff dff_B_yKHAQ7bZ8_1(.din(w_dff_B_SAF5a7wU9_1),.dout(w_dff_B_yKHAQ7bZ8_1),.clk(gclk));
	jdff dff_B_X07PlIy63_1(.din(w_dff_B_yKHAQ7bZ8_1),.dout(w_dff_B_X07PlIy63_1),.clk(gclk));
	jdff dff_B_m65lksJo0_1(.din(w_dff_B_X07PlIy63_1),.dout(w_dff_B_m65lksJo0_1),.clk(gclk));
	jdff dff_B_0erNJKzh6_1(.din(w_dff_B_m65lksJo0_1),.dout(w_dff_B_0erNJKzh6_1),.clk(gclk));
	jdff dff_B_iZMOoaEc6_1(.din(w_dff_B_0erNJKzh6_1),.dout(w_dff_B_iZMOoaEc6_1),.clk(gclk));
	jdff dff_B_R9RicJHW6_1(.din(w_dff_B_iZMOoaEc6_1),.dout(w_dff_B_R9RicJHW6_1),.clk(gclk));
	jdff dff_B_aDb6Ttog1_1(.din(w_dff_B_R9RicJHW6_1),.dout(w_dff_B_aDb6Ttog1_1),.clk(gclk));
	jdff dff_B_m0F1ncWq9_1(.din(w_dff_B_aDb6Ttog1_1),.dout(w_dff_B_m0F1ncWq9_1),.clk(gclk));
	jdff dff_B_bw5EIPSK4_1(.din(w_dff_B_m0F1ncWq9_1),.dout(w_dff_B_bw5EIPSK4_1),.clk(gclk));
	jdff dff_B_XRoBwbH59_1(.din(w_dff_B_bw5EIPSK4_1),.dout(w_dff_B_XRoBwbH59_1),.clk(gclk));
	jdff dff_B_bwo9Ndcl8_1(.din(n190),.dout(w_dff_B_bwo9Ndcl8_1),.clk(gclk));
	jdff dff_B_O2ProZuN1_1(.din(w_dff_B_bwo9Ndcl8_1),.dout(w_dff_B_O2ProZuN1_1),.clk(gclk));
	jdff dff_B_tDQLSqeZ0_1(.din(w_dff_B_O2ProZuN1_1),.dout(w_dff_B_tDQLSqeZ0_1),.clk(gclk));
	jdff dff_B_rnxsM0XU5_1(.din(w_dff_B_tDQLSqeZ0_1),.dout(w_dff_B_rnxsM0XU5_1),.clk(gclk));
	jdff dff_B_hikrsU7Z5_1(.din(w_dff_B_rnxsM0XU5_1),.dout(w_dff_B_hikrsU7Z5_1),.clk(gclk));
	jdff dff_B_8IOPiCWU6_1(.din(w_dff_B_hikrsU7Z5_1),.dout(w_dff_B_8IOPiCWU6_1),.clk(gclk));
	jdff dff_B_4MbmWuke4_1(.din(w_dff_B_8IOPiCWU6_1),.dout(w_dff_B_4MbmWuke4_1),.clk(gclk));
	jdff dff_B_KTg1yAft1_1(.din(w_dff_B_4MbmWuke4_1),.dout(w_dff_B_KTg1yAft1_1),.clk(gclk));
	jdff dff_B_XEkyDelF6_1(.din(w_dff_B_KTg1yAft1_1),.dout(w_dff_B_XEkyDelF6_1),.clk(gclk));
	jdff dff_B_9z3QR0bs6_1(.din(w_dff_B_XEkyDelF6_1),.dout(w_dff_B_9z3QR0bs6_1),.clk(gclk));
	jdff dff_B_AftZ3Wo78_1(.din(w_dff_B_9z3QR0bs6_1),.dout(w_dff_B_AftZ3Wo78_1),.clk(gclk));
	jdff dff_B_7nSYDCnB8_1(.din(w_dff_B_AftZ3Wo78_1),.dout(w_dff_B_7nSYDCnB8_1),.clk(gclk));
	jdff dff_B_GotyeNsY1_1(.din(w_dff_B_7nSYDCnB8_1),.dout(w_dff_B_GotyeNsY1_1),.clk(gclk));
	jdff dff_B_PlDjCZY22_1(.din(w_dff_B_GotyeNsY1_1),.dout(w_dff_B_PlDjCZY22_1),.clk(gclk));
	jdff dff_A_PiFD3WSk3_0(.dout(w_n185_0[0]),.din(w_dff_A_PiFD3WSk3_0),.clk(gclk));
	jdff dff_A_OMLjdNpq0_0(.dout(w_dff_A_PiFD3WSk3_0),.din(w_dff_A_OMLjdNpq0_0),.clk(gclk));
	jdff dff_A_eBwg2Bxj9_0(.dout(w_dff_A_OMLjdNpq0_0),.din(w_dff_A_eBwg2Bxj9_0),.clk(gclk));
	jdff dff_A_TLy8opGb5_0(.dout(w_dff_A_eBwg2Bxj9_0),.din(w_dff_A_TLy8opGb5_0),.clk(gclk));
	jdff dff_A_zvdmaR5U2_0(.dout(w_dff_A_TLy8opGb5_0),.din(w_dff_A_zvdmaR5U2_0),.clk(gclk));
	jdff dff_B_QQbq5IlY3_2(.din(n185),.dout(w_dff_B_QQbq5IlY3_2),.clk(gclk));
	jdff dff_B_OZd97weI4_2(.din(w_dff_B_QQbq5IlY3_2),.dout(w_dff_B_OZd97weI4_2),.clk(gclk));
	jdff dff_B_P5IQ1JFW2_2(.din(w_dff_B_OZd97weI4_2),.dout(w_dff_B_P5IQ1JFW2_2),.clk(gclk));
	jdff dff_B_iunqsuTI3_2(.din(w_dff_B_P5IQ1JFW2_2),.dout(w_dff_B_iunqsuTI3_2),.clk(gclk));
	jdff dff_B_gtk4BpM27_2(.din(w_dff_B_iunqsuTI3_2),.dout(w_dff_B_gtk4BpM27_2),.clk(gclk));
	jdff dff_B_AOsJNhcZ1_2(.din(w_dff_B_gtk4BpM27_2),.dout(w_dff_B_AOsJNhcZ1_2),.clk(gclk));
	jdff dff_B_pzAcnuhG5_2(.din(w_dff_B_AOsJNhcZ1_2),.dout(w_dff_B_pzAcnuhG5_2),.clk(gclk));
	jdff dff_B_Dbx0aZZD7_2(.din(w_dff_B_pzAcnuhG5_2),.dout(w_dff_B_Dbx0aZZD7_2),.clk(gclk));
	jdff dff_B_MnC1J1qK4_2(.din(w_dff_B_Dbx0aZZD7_2),.dout(w_dff_B_MnC1J1qK4_2),.clk(gclk));
	jdff dff_B_dcRO4kWi7_2(.din(w_dff_B_MnC1J1qK4_2),.dout(w_dff_B_dcRO4kWi7_2),.clk(gclk));
	jdff dff_B_cjtuyWXx7_2(.din(w_dff_B_dcRO4kWi7_2),.dout(w_dff_B_cjtuyWXx7_2),.clk(gclk));
	jdff dff_B_iyYNJnsV9_2(.din(w_dff_B_cjtuyWXx7_2),.dout(w_dff_B_iyYNJnsV9_2),.clk(gclk));
	jdff dff_B_1JorpXEE6_2(.din(w_dff_B_iyYNJnsV9_2),.dout(w_dff_B_1JorpXEE6_2),.clk(gclk));
	jdff dff_B_y54Z7sHy7_2(.din(w_dff_B_1JorpXEE6_2),.dout(w_dff_B_y54Z7sHy7_2),.clk(gclk));
	jdff dff_B_oiWBOB7h9_2(.din(n281),.dout(w_dff_B_oiWBOB7h9_2),.clk(gclk));
	jdff dff_A_DgN3MSVq3_0(.dout(w_n149_0[0]),.din(w_dff_A_DgN3MSVq3_0),.clk(gclk));
	jdff dff_A_82TKdms76_0(.dout(w_dff_A_DgN3MSVq3_0),.din(w_dff_A_82TKdms76_0),.clk(gclk));
	jdff dff_A_3SzNbMJf1_0(.dout(w_dff_A_82TKdms76_0),.din(w_dff_A_3SzNbMJf1_0),.clk(gclk));
	jdff dff_A_jeePaV4h6_0(.dout(w_dff_A_3SzNbMJf1_0),.din(w_dff_A_jeePaV4h6_0),.clk(gclk));
	jdff dff_A_xnsN78VT8_0(.dout(w_dff_A_jeePaV4h6_0),.din(w_dff_A_xnsN78VT8_0),.clk(gclk));
	jdff dff_B_GIyhLYus5_2(.din(n149),.dout(w_dff_B_GIyhLYus5_2),.clk(gclk));
	jdff dff_B_PwQ2kG6V7_2(.din(w_dff_B_GIyhLYus5_2),.dout(w_dff_B_PwQ2kG6V7_2),.clk(gclk));
	jdff dff_B_ZbC8dhtR8_2(.din(w_dff_B_PwQ2kG6V7_2),.dout(w_dff_B_ZbC8dhtR8_2),.clk(gclk));
	jdff dff_B_2SXjRmGM2_2(.din(w_dff_B_ZbC8dhtR8_2),.dout(w_dff_B_2SXjRmGM2_2),.clk(gclk));
	jdff dff_B_LvX2UqvK5_2(.din(w_dff_B_2SXjRmGM2_2),.dout(w_dff_B_LvX2UqvK5_2),.clk(gclk));
	jdff dff_B_BKDMNEAh6_2(.din(w_dff_B_LvX2UqvK5_2),.dout(w_dff_B_BKDMNEAh6_2),.clk(gclk));
	jdff dff_B_O2oHx9JX0_2(.din(w_dff_B_BKDMNEAh6_2),.dout(w_dff_B_O2oHx9JX0_2),.clk(gclk));
	jdff dff_B_3IVECn2B0_2(.din(w_dff_B_O2oHx9JX0_2),.dout(w_dff_B_3IVECn2B0_2),.clk(gclk));
	jdff dff_B_B5gS4YMs9_2(.din(w_dff_B_3IVECn2B0_2),.dout(w_dff_B_B5gS4YMs9_2),.clk(gclk));
	jdff dff_B_Laq60N2c5_2(.din(w_dff_B_B5gS4YMs9_2),.dout(w_dff_B_Laq60N2c5_2),.clk(gclk));
	jdff dff_B_TO6m9H4P8_2(.din(w_dff_B_Laq60N2c5_2),.dout(w_dff_B_TO6m9H4P8_2),.clk(gclk));
	jdff dff_B_R8eM2w5n0_2(.din(w_dff_B_TO6m9H4P8_2),.dout(w_dff_B_R8eM2w5n0_2),.clk(gclk));
	jdff dff_B_cEebf5uW0_2(.din(w_dff_B_R8eM2w5n0_2),.dout(w_dff_B_cEebf5uW0_2),.clk(gclk));
	jdff dff_B_jl8Wcy995_2(.din(w_dff_B_cEebf5uW0_2),.dout(w_dff_B_jl8Wcy995_2),.clk(gclk));
	jdff dff_A_RM1anhUw6_0(.dout(w_n183_0[0]),.din(w_dff_A_RM1anhUw6_0),.clk(gclk));
	jdff dff_A_sKthbOZ28_0(.dout(w_dff_A_RM1anhUw6_0),.din(w_dff_A_sKthbOZ28_0),.clk(gclk));
	jdff dff_A_ZcZgjok87_0(.dout(w_dff_A_sKthbOZ28_0),.din(w_dff_A_ZcZgjok87_0),.clk(gclk));
	jdff dff_A_D2pY2psu8_0(.dout(w_dff_A_ZcZgjok87_0),.din(w_dff_A_D2pY2psu8_0),.clk(gclk));
	jdff dff_A_fMuf9xEt9_0(.dout(w_dff_A_D2pY2psu8_0),.din(w_dff_A_fMuf9xEt9_0),.clk(gclk));
	jdff dff_A_8Dmcj8nY2_0(.dout(w_dff_A_fMuf9xEt9_0),.din(w_dff_A_8Dmcj8nY2_0),.clk(gclk));
	jdff dff_A_UtKslg8F9_0(.dout(w_n271_0[0]),.din(w_dff_A_UtKslg8F9_0),.clk(gclk));
	jdff dff_A_1hTnlo0v1_0(.dout(w_dff_A_UtKslg8F9_0),.din(w_dff_A_1hTnlo0v1_0),.clk(gclk));
	jdff dff_A_frZW8Ixb0_0(.dout(w_dff_A_1hTnlo0v1_0),.din(w_dff_A_frZW8Ixb0_0),.clk(gclk));
	jdff dff_B_ZhxoKhHD8_1(.din(n217),.dout(w_dff_B_ZhxoKhHD8_1),.clk(gclk));
	jdff dff_B_zJt6HAym3_0(.din(n243),.dout(w_dff_B_zJt6HAym3_0),.clk(gclk));
	jdff dff_A_WPTe1u9q5_0(.dout(w_G27gat_0[0]),.din(w_dff_A_WPTe1u9q5_0),.clk(gclk));
	jdff dff_A_GSNYGnTk2_0(.dout(w_dff_A_WPTe1u9q5_0),.din(w_dff_A_GSNYGnTk2_0),.clk(gclk));
	jdff dff_A_kqEjlvSJ1_0(.dout(w_dff_A_GSNYGnTk2_0),.din(w_dff_A_kqEjlvSJ1_0),.clk(gclk));
	jdff dff_A_VCL4iba75_0(.dout(w_dff_A_kqEjlvSJ1_0),.din(w_dff_A_VCL4iba75_0),.clk(gclk));
	jdff dff_A_1w8blDM99_0(.dout(w_dff_A_VCL4iba75_0),.din(w_dff_A_1w8blDM99_0),.clk(gclk));
	jdff dff_A_qWk2rJrB6_0(.dout(w_dff_A_1w8blDM99_0),.din(w_dff_A_qWk2rJrB6_0),.clk(gclk));
	jdff dff_A_DzX34acp6_0(.dout(w_dff_A_qWk2rJrB6_0),.din(w_dff_A_DzX34acp6_0),.clk(gclk));
	jdff dff_A_aCCqTrBc7_0(.dout(w_dff_A_DzX34acp6_0),.din(w_dff_A_aCCqTrBc7_0),.clk(gclk));
	jdff dff_A_SWPagyCX3_0(.dout(w_dff_A_aCCqTrBc7_0),.din(w_dff_A_SWPagyCX3_0),.clk(gclk));
	jdff dff_A_QTPwGdp08_0(.dout(w_dff_A_SWPagyCX3_0),.din(w_dff_A_QTPwGdp08_0),.clk(gclk));
	jdff dff_A_Rq4e2tBh2_0(.dout(w_dff_A_QTPwGdp08_0),.din(w_dff_A_Rq4e2tBh2_0),.clk(gclk));
	jdff dff_A_NxpvU0VK7_0(.dout(w_dff_A_Rq4e2tBh2_0),.din(w_dff_A_NxpvU0VK7_0),.clk(gclk));
	jdff dff_A_wgEUhDkE2_0(.dout(w_dff_A_NxpvU0VK7_0),.din(w_dff_A_wgEUhDkE2_0),.clk(gclk));
	jdff dff_A_arkkcmbz7_0(.dout(w_dff_A_wgEUhDkE2_0),.din(w_dff_A_arkkcmbz7_0),.clk(gclk));
	jdff dff_A_mAgQsyME8_0(.dout(w_dff_A_arkkcmbz7_0),.din(w_dff_A_mAgQsyME8_0),.clk(gclk));
	jdff dff_A_kNAQRqxn5_0(.dout(w_G115gat_0[0]),.din(w_dff_A_kNAQRqxn5_0),.clk(gclk));
	jdff dff_A_vY8QnSd14_0(.dout(w_dff_A_kNAQRqxn5_0),.din(w_dff_A_vY8QnSd14_0),.clk(gclk));
	jdff dff_A_zzuNB8Ds1_0(.dout(w_dff_A_vY8QnSd14_0),.din(w_dff_A_zzuNB8Ds1_0),.clk(gclk));
	jdff dff_A_FAluccEs6_0(.dout(w_dff_A_zzuNB8Ds1_0),.din(w_dff_A_FAluccEs6_0),.clk(gclk));
	jdff dff_A_1gshwirA9_0(.dout(w_dff_A_FAluccEs6_0),.din(w_dff_A_1gshwirA9_0),.clk(gclk));
	jdff dff_A_dxkrPtun8_0(.dout(w_dff_A_1gshwirA9_0),.din(w_dff_A_dxkrPtun8_0),.clk(gclk));
	jdff dff_A_u6BXhCcu8_0(.dout(w_dff_A_dxkrPtun8_0),.din(w_dff_A_u6BXhCcu8_0),.clk(gclk));
	jdff dff_A_bsEdBsHB3_0(.dout(w_dff_A_u6BXhCcu8_0),.din(w_dff_A_bsEdBsHB3_0),.clk(gclk));
	jdff dff_A_UOSQooNn3_0(.dout(w_dff_A_bsEdBsHB3_0),.din(w_dff_A_UOSQooNn3_0),.clk(gclk));
	jdff dff_A_1B5QYVXI4_0(.dout(w_dff_A_UOSQooNn3_0),.din(w_dff_A_1B5QYVXI4_0),.clk(gclk));
	jdff dff_A_XJLVieiL0_0(.dout(w_dff_A_1B5QYVXI4_0),.din(w_dff_A_XJLVieiL0_0),.clk(gclk));
	jdff dff_A_jFB0XQEE4_0(.dout(w_dff_A_XJLVieiL0_0),.din(w_dff_A_jFB0XQEE4_0),.clk(gclk));
	jdff dff_A_UP0ZRpiA9_0(.dout(w_dff_A_jFB0XQEE4_0),.din(w_dff_A_UP0ZRpiA9_0),.clk(gclk));
	jdff dff_A_iuNc7Xhb9_0(.dout(w_dff_A_UP0ZRpiA9_0),.din(w_dff_A_iuNc7Xhb9_0),.clk(gclk));
	jdff dff_A_HRDrLIPA2_0(.dout(w_dff_A_iuNc7Xhb9_0),.din(w_dff_A_HRDrLIPA2_0),.clk(gclk));
	jdff dff_A_yzk0Ipx60_0(.dout(w_n230_0[0]),.din(w_dff_A_yzk0Ipx60_0),.clk(gclk));
	jdff dff_A_RAmVZyC48_0(.dout(w_dff_A_yzk0Ipx60_0),.din(w_dff_A_RAmVZyC48_0),.clk(gclk));
	jdff dff_A_n93NZ9wV0_0(.dout(w_dff_A_RAmVZyC48_0),.din(w_dff_A_n93NZ9wV0_0),.clk(gclk));
	jdff dff_A_ITq3EleO6_0(.dout(w_dff_A_n93NZ9wV0_0),.din(w_dff_A_ITq3EleO6_0),.clk(gclk));
	jdff dff_A_mCrN3Lj91_0(.dout(w_dff_A_ITq3EleO6_0),.din(w_dff_A_mCrN3Lj91_0),.clk(gclk));
	jdff dff_A_4hKeouNQ8_0(.dout(w_dff_A_mCrN3Lj91_0),.din(w_dff_A_4hKeouNQ8_0),.clk(gclk));
	jdff dff_A_CQcrHCBb6_0(.dout(w_G92gat_0[0]),.din(w_dff_A_CQcrHCBb6_0),.clk(gclk));
	jdff dff_A_C1l3zL6B5_0(.dout(w_dff_A_CQcrHCBb6_0),.din(w_dff_A_C1l3zL6B5_0),.clk(gclk));
	jdff dff_A_YD7hr8tY0_0(.dout(w_dff_A_C1l3zL6B5_0),.din(w_dff_A_YD7hr8tY0_0),.clk(gclk));
	jdff dff_A_i0KCF6q20_0(.dout(w_dff_A_YD7hr8tY0_0),.din(w_dff_A_i0KCF6q20_0),.clk(gclk));
	jdff dff_A_4dtMxGzU6_0(.dout(w_dff_A_i0KCF6q20_0),.din(w_dff_A_4dtMxGzU6_0),.clk(gclk));
	jdff dff_A_z1qq2N689_0(.dout(w_dff_A_4dtMxGzU6_0),.din(w_dff_A_z1qq2N689_0),.clk(gclk));
	jdff dff_A_cDTPGoMq9_0(.dout(w_dff_A_z1qq2N689_0),.din(w_dff_A_cDTPGoMq9_0),.clk(gclk));
	jdff dff_A_ieM7F0Qu8_0(.dout(w_dff_A_cDTPGoMq9_0),.din(w_dff_A_ieM7F0Qu8_0),.clk(gclk));
	jdff dff_A_z9Dm9cNI4_0(.dout(w_dff_A_ieM7F0Qu8_0),.din(w_dff_A_z9Dm9cNI4_0),.clk(gclk));
	jdff dff_A_bNf7nTdS6_0(.dout(w_dff_A_z9Dm9cNI4_0),.din(w_dff_A_bNf7nTdS6_0),.clk(gclk));
	jdff dff_A_67IY7bF71_0(.dout(w_dff_A_bNf7nTdS6_0),.din(w_dff_A_67IY7bF71_0),.clk(gclk));
	jdff dff_A_KCe3CFxT9_0(.dout(w_dff_A_67IY7bF71_0),.din(w_dff_A_KCe3CFxT9_0),.clk(gclk));
	jdff dff_A_V9xet9mD8_0(.dout(w_dff_A_KCe3CFxT9_0),.din(w_dff_A_V9xet9mD8_0),.clk(gclk));
	jdff dff_A_Ce1tMWSv9_0(.dout(w_dff_A_V9xet9mD8_0),.din(w_dff_A_Ce1tMWSv9_0),.clk(gclk));
	jdff dff_A_lorB278v7_0(.dout(w_dff_A_Ce1tMWSv9_0),.din(w_dff_A_lorB278v7_0),.clk(gclk));
	jdff dff_A_8sSn4NmT8_0(.dout(w_dff_A_lorB278v7_0),.din(w_dff_A_8sSn4NmT8_0),.clk(gclk));
	jdff dff_A_TPK5Ey768_0(.dout(w_dff_A_8sSn4NmT8_0),.din(w_dff_A_TPK5Ey768_0),.clk(gclk));
	jdff dff_A_1LZv9Un12_0(.dout(w_dff_A_TPK5Ey768_0),.din(w_dff_A_1LZv9Un12_0),.clk(gclk));
	jdff dff_A_loKggvBq6_0(.dout(w_dff_A_1LZv9Un12_0),.din(w_dff_A_loKggvBq6_0),.clk(gclk));
	jdff dff_A_FEf1B7nZ7_0(.dout(w_dff_A_loKggvBq6_0),.din(w_dff_A_FEf1B7nZ7_0),.clk(gclk));
	jdff dff_A_2uLs2c3S9_1(.dout(w_G92gat_0[1]),.din(w_dff_A_2uLs2c3S9_1),.clk(gclk));
	jdff dff_A_AhuKunsi1_1(.dout(w_dff_A_2uLs2c3S9_1),.din(w_dff_A_AhuKunsi1_1),.clk(gclk));
	jdff dff_A_pcFbUBcz9_1(.dout(w_dff_A_AhuKunsi1_1),.din(w_dff_A_pcFbUBcz9_1),.clk(gclk));
	jdff dff_A_s3eF31HN8_1(.dout(w_dff_A_pcFbUBcz9_1),.din(w_dff_A_s3eF31HN8_1),.clk(gclk));
	jdff dff_A_MsmPoJDb8_1(.dout(w_dff_A_s3eF31HN8_1),.din(w_dff_A_MsmPoJDb8_1),.clk(gclk));
	jdff dff_A_Xfxgwyf14_1(.dout(w_dff_A_MsmPoJDb8_1),.din(w_dff_A_Xfxgwyf14_1),.clk(gclk));
	jdff dff_A_FFB9MV8l1_1(.dout(w_dff_A_Xfxgwyf14_1),.din(w_dff_A_FFB9MV8l1_1),.clk(gclk));
	jdff dff_A_LVJrnfm42_1(.dout(w_dff_A_FFB9MV8l1_1),.din(w_dff_A_LVJrnfm42_1),.clk(gclk));
	jdff dff_A_14DWDvVg9_1(.dout(w_dff_A_LVJrnfm42_1),.din(w_dff_A_14DWDvVg9_1),.clk(gclk));
	jdff dff_A_3upgWeKT5_1(.dout(w_dff_A_14DWDvVg9_1),.din(w_dff_A_3upgWeKT5_1),.clk(gclk));
	jdff dff_A_kTp2LQFU5_1(.dout(w_dff_A_3upgWeKT5_1),.din(w_dff_A_kTp2LQFU5_1),.clk(gclk));
	jdff dff_A_b2buw0UU4_1(.dout(w_dff_A_kTp2LQFU5_1),.din(w_dff_A_b2buw0UU4_1),.clk(gclk));
	jdff dff_A_OGEALcHA6_1(.dout(w_dff_A_b2buw0UU4_1),.din(w_dff_A_OGEALcHA6_1),.clk(gclk));
	jdff dff_A_MxjzSkw00_1(.dout(w_dff_A_OGEALcHA6_1),.din(w_dff_A_MxjzSkw00_1),.clk(gclk));
	jdff dff_A_PWYb19Y21_1(.dout(w_dff_A_MxjzSkw00_1),.din(w_dff_A_PWYb19Y21_1),.clk(gclk));
	jdff dff_A_f59jYA8P5_0(.dout(w_n227_0[0]),.din(w_dff_A_f59jYA8P5_0),.clk(gclk));
	jdff dff_A_pRmMQpeE8_0(.dout(w_dff_A_f59jYA8P5_0),.din(w_dff_A_pRmMQpeE8_0),.clk(gclk));
	jdff dff_A_QIn5Lzi67_0(.dout(w_dff_A_pRmMQpeE8_0),.din(w_dff_A_QIn5Lzi67_0),.clk(gclk));
	jdff dff_A_AjrOsry46_0(.dout(w_dff_A_QIn5Lzi67_0),.din(w_dff_A_AjrOsry46_0),.clk(gclk));
	jdff dff_A_Qx88tkmG9_0(.dout(w_dff_A_AjrOsry46_0),.din(w_dff_A_Qx88tkmG9_0),.clk(gclk));
	jdff dff_A_l6vhJiZM3_0(.dout(w_dff_A_Qx88tkmG9_0),.din(w_dff_A_l6vhJiZM3_0),.clk(gclk));
	jdff dff_A_isqtWgis2_0(.dout(w_G14gat_0[0]),.din(w_dff_A_isqtWgis2_0),.clk(gclk));
	jdff dff_A_ITwmwsQp0_0(.dout(w_dff_A_isqtWgis2_0),.din(w_dff_A_ITwmwsQp0_0),.clk(gclk));
	jdff dff_A_wBFge4ko1_0(.dout(w_dff_A_ITwmwsQp0_0),.din(w_dff_A_wBFge4ko1_0),.clk(gclk));
	jdff dff_A_ZxDfTi8f3_0(.dout(w_dff_A_wBFge4ko1_0),.din(w_dff_A_ZxDfTi8f3_0),.clk(gclk));
	jdff dff_A_wwlGmWnf0_0(.dout(w_dff_A_ZxDfTi8f3_0),.din(w_dff_A_wwlGmWnf0_0),.clk(gclk));
	jdff dff_A_yTO17ioo5_0(.dout(w_dff_A_wwlGmWnf0_0),.din(w_dff_A_yTO17ioo5_0),.clk(gclk));
	jdff dff_A_Cw8fn0Qz3_0(.dout(w_dff_A_yTO17ioo5_0),.din(w_dff_A_Cw8fn0Qz3_0),.clk(gclk));
	jdff dff_A_Dgi3RNPu2_0(.dout(w_dff_A_Cw8fn0Qz3_0),.din(w_dff_A_Dgi3RNPu2_0),.clk(gclk));
	jdff dff_A_tOFYThyM9_0(.dout(w_dff_A_Dgi3RNPu2_0),.din(w_dff_A_tOFYThyM9_0),.clk(gclk));
	jdff dff_A_AUmjnKpy6_0(.dout(w_dff_A_tOFYThyM9_0),.din(w_dff_A_AUmjnKpy6_0),.clk(gclk));
	jdff dff_A_kz696BsN3_0(.dout(w_dff_A_AUmjnKpy6_0),.din(w_dff_A_kz696BsN3_0),.clk(gclk));
	jdff dff_A_PsC3Z56w8_0(.dout(w_dff_A_kz696BsN3_0),.din(w_dff_A_PsC3Z56w8_0),.clk(gclk));
	jdff dff_A_32rDj0y51_0(.dout(w_dff_A_PsC3Z56w8_0),.din(w_dff_A_32rDj0y51_0),.clk(gclk));
	jdff dff_A_awSD8oBC8_0(.dout(w_dff_A_32rDj0y51_0),.din(w_dff_A_awSD8oBC8_0),.clk(gclk));
	jdff dff_A_bMTPEd8B3_0(.dout(w_dff_A_awSD8oBC8_0),.din(w_dff_A_bMTPEd8B3_0),.clk(gclk));
	jdff dff_A_KgaLiSJk5_0(.dout(w_dff_A_bMTPEd8B3_0),.din(w_dff_A_KgaLiSJk5_0),.clk(gclk));
	jdff dff_A_SifZUAWh9_0(.dout(w_dff_A_KgaLiSJk5_0),.din(w_dff_A_SifZUAWh9_0),.clk(gclk));
	jdff dff_A_WB3qmmwu6_0(.dout(w_dff_A_SifZUAWh9_0),.din(w_dff_A_WB3qmmwu6_0),.clk(gclk));
	jdff dff_A_1mWI1GVB8_0(.dout(w_dff_A_WB3qmmwu6_0),.din(w_dff_A_1mWI1GVB8_0),.clk(gclk));
	jdff dff_A_X7CJlDZg1_0(.dout(w_dff_A_1mWI1GVB8_0),.din(w_dff_A_X7CJlDZg1_0),.clk(gclk));
	jdff dff_A_HjH7T54d8_1(.dout(w_G14gat_0[1]),.din(w_dff_A_HjH7T54d8_1),.clk(gclk));
	jdff dff_A_Jjd5WVeh4_1(.dout(w_dff_A_HjH7T54d8_1),.din(w_dff_A_Jjd5WVeh4_1),.clk(gclk));
	jdff dff_A_vzidcSnN8_1(.dout(w_dff_A_Jjd5WVeh4_1),.din(w_dff_A_vzidcSnN8_1),.clk(gclk));
	jdff dff_A_0BDYz8ZI6_1(.dout(w_dff_A_vzidcSnN8_1),.din(w_dff_A_0BDYz8ZI6_1),.clk(gclk));
	jdff dff_A_dSPJwEna1_1(.dout(w_dff_A_0BDYz8ZI6_1),.din(w_dff_A_dSPJwEna1_1),.clk(gclk));
	jdff dff_A_wA5Uq0Mn6_1(.dout(w_dff_A_dSPJwEna1_1),.din(w_dff_A_wA5Uq0Mn6_1),.clk(gclk));
	jdff dff_A_CmdJG8Ph9_1(.dout(w_dff_A_wA5Uq0Mn6_1),.din(w_dff_A_CmdJG8Ph9_1),.clk(gclk));
	jdff dff_A_CzKBE1lf3_1(.dout(w_dff_A_CmdJG8Ph9_1),.din(w_dff_A_CzKBE1lf3_1),.clk(gclk));
	jdff dff_A_J9fnEt7q1_1(.dout(w_dff_A_CzKBE1lf3_1),.din(w_dff_A_J9fnEt7q1_1),.clk(gclk));
	jdff dff_A_s4X9JNUG4_1(.dout(w_dff_A_J9fnEt7q1_1),.din(w_dff_A_s4X9JNUG4_1),.clk(gclk));
	jdff dff_A_6TGauh890_1(.dout(w_dff_A_s4X9JNUG4_1),.din(w_dff_A_6TGauh890_1),.clk(gclk));
	jdff dff_A_4bV3bnYD5_1(.dout(w_dff_A_6TGauh890_1),.din(w_dff_A_4bV3bnYD5_1),.clk(gclk));
	jdff dff_A_eSG4JE0Y4_1(.dout(w_dff_A_4bV3bnYD5_1),.din(w_dff_A_eSG4JE0Y4_1),.clk(gclk));
	jdff dff_A_cyGpAo5m7_1(.dout(w_dff_A_eSG4JE0Y4_1),.din(w_dff_A_cyGpAo5m7_1),.clk(gclk));
	jdff dff_A_zfRanZFb5_1(.dout(w_dff_A_cyGpAo5m7_1),.din(w_dff_A_zfRanZFb5_1),.clk(gclk));
	jdff dff_B_Vv1U1Xsw1_1(.din(n221),.dout(w_dff_B_Vv1U1Xsw1_1),.clk(gclk));
	jdff dff_B_8QAkKt3M0_1(.din(w_dff_B_Vv1U1Xsw1_1),.dout(w_dff_B_8QAkKt3M0_1),.clk(gclk));
	jdff dff_B_355MOtrO4_1(.din(w_dff_B_8QAkKt3M0_1),.dout(w_dff_B_355MOtrO4_1),.clk(gclk));
	jdff dff_B_it2znLd43_1(.din(w_dff_B_355MOtrO4_1),.dout(w_dff_B_it2znLd43_1),.clk(gclk));
	jdff dff_B_NyDAsDHa5_1(.din(w_dff_B_it2znLd43_1),.dout(w_dff_B_NyDAsDHa5_1),.clk(gclk));
	jdff dff_A_ly6rZopT4_0(.dout(w_G66gat_0[0]),.din(w_dff_A_ly6rZopT4_0),.clk(gclk));
	jdff dff_A_gyXE4MHt9_0(.dout(w_dff_A_ly6rZopT4_0),.din(w_dff_A_gyXE4MHt9_0),.clk(gclk));
	jdff dff_A_iWtpklWD3_0(.dout(w_dff_A_gyXE4MHt9_0),.din(w_dff_A_iWtpklWD3_0),.clk(gclk));
	jdff dff_A_ukOAbM1O3_0(.dout(w_dff_A_iWtpklWD3_0),.din(w_dff_A_ukOAbM1O3_0),.clk(gclk));
	jdff dff_A_KHlim5GW8_0(.dout(w_dff_A_ukOAbM1O3_0),.din(w_dff_A_KHlim5GW8_0),.clk(gclk));
	jdff dff_A_o4Gn8Rp16_0(.dout(w_dff_A_KHlim5GW8_0),.din(w_dff_A_o4Gn8Rp16_0),.clk(gclk));
	jdff dff_A_htKJlJg06_0(.dout(w_dff_A_o4Gn8Rp16_0),.din(w_dff_A_htKJlJg06_0),.clk(gclk));
	jdff dff_A_iyv5sVN33_0(.dout(w_dff_A_htKJlJg06_0),.din(w_dff_A_iyv5sVN33_0),.clk(gclk));
	jdff dff_A_jUuZdhSc6_0(.dout(w_dff_A_iyv5sVN33_0),.din(w_dff_A_jUuZdhSc6_0),.clk(gclk));
	jdff dff_A_qUxF57Qh6_0(.dout(w_dff_A_jUuZdhSc6_0),.din(w_dff_A_qUxF57Qh6_0),.clk(gclk));
	jdff dff_A_Q9c17TY98_0(.dout(w_dff_A_qUxF57Qh6_0),.din(w_dff_A_Q9c17TY98_0),.clk(gclk));
	jdff dff_A_xKPOWsTF8_0(.dout(w_dff_A_Q9c17TY98_0),.din(w_dff_A_xKPOWsTF8_0),.clk(gclk));
	jdff dff_A_C3dt0v0v1_0(.dout(w_dff_A_xKPOWsTF8_0),.din(w_dff_A_C3dt0v0v1_0),.clk(gclk));
	jdff dff_A_FZnNBvdh3_0(.dout(w_dff_A_C3dt0v0v1_0),.din(w_dff_A_FZnNBvdh3_0),.clk(gclk));
	jdff dff_A_xWYS2Qnl3_0(.dout(w_dff_A_FZnNBvdh3_0),.din(w_dff_A_xWYS2Qnl3_0),.clk(gclk));
	jdff dff_A_WUcUq3Y59_0(.dout(w_dff_A_xWYS2Qnl3_0),.din(w_dff_A_WUcUq3Y59_0),.clk(gclk));
	jdff dff_A_8TKz3JAl9_0(.dout(w_dff_A_WUcUq3Y59_0),.din(w_dff_A_8TKz3JAl9_0),.clk(gclk));
	jdff dff_A_hMc6BZEG9_0(.dout(w_dff_A_8TKz3JAl9_0),.din(w_dff_A_hMc6BZEG9_0),.clk(gclk));
	jdff dff_A_Qp1Rk47H9_0(.dout(w_dff_A_hMc6BZEG9_0),.din(w_dff_A_Qp1Rk47H9_0),.clk(gclk));
	jdff dff_A_pw1kHjUz2_0(.dout(w_dff_A_Qp1Rk47H9_0),.din(w_dff_A_pw1kHjUz2_0),.clk(gclk));
	jdff dff_A_6mPWo1Ja7_1(.dout(w_G66gat_0[1]),.din(w_dff_A_6mPWo1Ja7_1),.clk(gclk));
	jdff dff_A_b0eEEZzx3_1(.dout(w_dff_A_6mPWo1Ja7_1),.din(w_dff_A_b0eEEZzx3_1),.clk(gclk));
	jdff dff_A_RChVbdHd9_1(.dout(w_dff_A_b0eEEZzx3_1),.din(w_dff_A_RChVbdHd9_1),.clk(gclk));
	jdff dff_A_Ug4oAg0y9_1(.dout(w_dff_A_RChVbdHd9_1),.din(w_dff_A_Ug4oAg0y9_1),.clk(gclk));
	jdff dff_A_CpzthAVL9_1(.dout(w_dff_A_Ug4oAg0y9_1),.din(w_dff_A_CpzthAVL9_1),.clk(gclk));
	jdff dff_A_r3ILZe7g6_1(.dout(w_dff_A_CpzthAVL9_1),.din(w_dff_A_r3ILZe7g6_1),.clk(gclk));
	jdff dff_A_jco5sZSn2_1(.dout(w_dff_A_r3ILZe7g6_1),.din(w_dff_A_jco5sZSn2_1),.clk(gclk));
	jdff dff_A_tBcWuE1L0_1(.dout(w_dff_A_jco5sZSn2_1),.din(w_dff_A_tBcWuE1L0_1),.clk(gclk));
	jdff dff_A_f9fvTdNm4_1(.dout(w_dff_A_tBcWuE1L0_1),.din(w_dff_A_f9fvTdNm4_1),.clk(gclk));
	jdff dff_A_RzDsK4NF5_1(.dout(w_dff_A_f9fvTdNm4_1),.din(w_dff_A_RzDsK4NF5_1),.clk(gclk));
	jdff dff_A_ymJMnyH77_1(.dout(w_dff_A_RzDsK4NF5_1),.din(w_dff_A_ymJMnyH77_1),.clk(gclk));
	jdff dff_A_8JAKO9mK3_1(.dout(w_dff_A_ymJMnyH77_1),.din(w_dff_A_8JAKO9mK3_1),.clk(gclk));
	jdff dff_A_JpuSwqI38_1(.dout(w_dff_A_8JAKO9mK3_1),.din(w_dff_A_JpuSwqI38_1),.clk(gclk));
	jdff dff_A_TlcIV72U0_1(.dout(w_dff_A_JpuSwqI38_1),.din(w_dff_A_TlcIV72U0_1),.clk(gclk));
	jdff dff_A_EGfukxDR9_1(.dout(w_dff_A_TlcIV72U0_1),.din(w_dff_A_EGfukxDR9_1),.clk(gclk));
	jdff dff_A_IYKTXbQ26_0(.dout(w_G40gat_0[0]),.din(w_dff_A_IYKTXbQ26_0),.clk(gclk));
	jdff dff_A_3MUahvAy4_0(.dout(w_dff_A_IYKTXbQ26_0),.din(w_dff_A_3MUahvAy4_0),.clk(gclk));
	jdff dff_A_YYeBLsx88_0(.dout(w_dff_A_3MUahvAy4_0),.din(w_dff_A_YYeBLsx88_0),.clk(gclk));
	jdff dff_A_VYWMwE812_0(.dout(w_dff_A_YYeBLsx88_0),.din(w_dff_A_VYWMwE812_0),.clk(gclk));
	jdff dff_A_CmjLWyko3_0(.dout(w_dff_A_VYWMwE812_0),.din(w_dff_A_CmjLWyko3_0),.clk(gclk));
	jdff dff_A_9zRzmdzM7_0(.dout(w_dff_A_CmjLWyko3_0),.din(w_dff_A_9zRzmdzM7_0),.clk(gclk));
	jdff dff_A_SyYmKoxZ3_0(.dout(w_dff_A_9zRzmdzM7_0),.din(w_dff_A_SyYmKoxZ3_0),.clk(gclk));
	jdff dff_A_cU0uybh90_0(.dout(w_dff_A_SyYmKoxZ3_0),.din(w_dff_A_cU0uybh90_0),.clk(gclk));
	jdff dff_A_FClwhfiw9_0(.dout(w_dff_A_cU0uybh90_0),.din(w_dff_A_FClwhfiw9_0),.clk(gclk));
	jdff dff_A_gUxxbEq39_0(.dout(w_dff_A_FClwhfiw9_0),.din(w_dff_A_gUxxbEq39_0),.clk(gclk));
	jdff dff_A_Ee5Gfiu55_0(.dout(w_dff_A_gUxxbEq39_0),.din(w_dff_A_Ee5Gfiu55_0),.clk(gclk));
	jdff dff_A_MFKm1KjX7_0(.dout(w_dff_A_Ee5Gfiu55_0),.din(w_dff_A_MFKm1KjX7_0),.clk(gclk));
	jdff dff_A_1MGRnFlX9_0(.dout(w_dff_A_MFKm1KjX7_0),.din(w_dff_A_1MGRnFlX9_0),.clk(gclk));
	jdff dff_A_rBTwsf5d4_0(.dout(w_dff_A_1MGRnFlX9_0),.din(w_dff_A_rBTwsf5d4_0),.clk(gclk));
	jdff dff_A_KwV5G41l5_0(.dout(w_dff_A_rBTwsf5d4_0),.din(w_dff_A_KwV5G41l5_0),.clk(gclk));
	jdff dff_A_XQDfzSS13_1(.dout(w_n147_0[1]),.din(w_dff_A_XQDfzSS13_1),.clk(gclk));
	jdff dff_B_fpzEPT5I7_0(.din(n146),.dout(w_dff_B_fpzEPT5I7_0),.clk(gclk));
	jdff dff_B_m25x534I1_0(.din(w_dff_B_fpzEPT5I7_0),.dout(w_dff_B_m25x534I1_0),.clk(gclk));
	jdff dff_B_7DzAXQHl2_0(.din(w_dff_B_m25x534I1_0),.dout(w_dff_B_7DzAXQHl2_0),.clk(gclk));
	jdff dff_B_LUBtFMM42_0(.din(w_dff_B_7DzAXQHl2_0),.dout(w_dff_B_LUBtFMM42_0),.clk(gclk));
	jdff dff_B_JCNH5Y7g8_0(.din(w_dff_B_LUBtFMM42_0),.dout(w_dff_B_JCNH5Y7g8_0),.clk(gclk));
	jdff dff_B_VFPT1eVQ5_0(.din(w_dff_B_JCNH5Y7g8_0),.dout(w_dff_B_VFPT1eVQ5_0),.clk(gclk));
	jdff dff_A_cAgb6sJp5_0(.dout(w_n145_0[0]),.din(w_dff_A_cAgb6sJp5_0),.clk(gclk));
	jdff dff_A_UwRY90fB9_0(.dout(w_dff_A_cAgb6sJp5_0),.din(w_dff_A_UwRY90fB9_0),.clk(gclk));
	jdff dff_A_oy9L780f9_0(.dout(w_dff_A_UwRY90fB9_0),.din(w_dff_A_oy9L780f9_0),.clk(gclk));
	jdff dff_A_YZGk8nx20_0(.dout(w_dff_A_oy9L780f9_0),.din(w_dff_A_YZGk8nx20_0),.clk(gclk));
	jdff dff_A_XGUntYs56_0(.dout(w_dff_A_YZGk8nx20_0),.din(w_dff_A_XGUntYs56_0),.clk(gclk));
	jdff dff_A_83uB0iM15_0(.dout(w_dff_A_XGUntYs56_0),.din(w_dff_A_83uB0iM15_0),.clk(gclk));
	jdff dff_A_HlQglHUY2_0(.dout(w_dff_A_83uB0iM15_0),.din(w_dff_A_HlQglHUY2_0),.clk(gclk));
	jdff dff_A_bF9J1icF2_0(.dout(w_dff_A_HlQglHUY2_0),.din(w_dff_A_bF9J1icF2_0),.clk(gclk));
	jdff dff_A_vDrPrNMf5_0(.dout(w_dff_A_bF9J1icF2_0),.din(w_dff_A_vDrPrNMf5_0),.clk(gclk));
	jdff dff_A_zbeykTCV7_0(.dout(w_dff_A_vDrPrNMf5_0),.din(w_dff_A_zbeykTCV7_0),.clk(gclk));
	jdff dff_A_AsDAUV2P7_0(.dout(w_dff_A_zbeykTCV7_0),.din(w_dff_A_AsDAUV2P7_0),.clk(gclk));
	jdff dff_A_MDnOkpYB1_0(.dout(w_dff_A_AsDAUV2P7_0),.din(w_dff_A_MDnOkpYB1_0),.clk(gclk));
	jdff dff_B_A5e2h8VR1_2(.din(n145),.dout(w_dff_B_A5e2h8VR1_2),.clk(gclk));
	jdff dff_B_YI0AwNSz6_2(.din(w_dff_B_A5e2h8VR1_2),.dout(w_dff_B_YI0AwNSz6_2),.clk(gclk));
	jdff dff_B_2X8y0zbI3_2(.din(w_dff_B_YI0AwNSz6_2),.dout(w_dff_B_2X8y0zbI3_2),.clk(gclk));
	jdff dff_B_3tLIWoyx4_2(.din(w_dff_B_2X8y0zbI3_2),.dout(w_dff_B_3tLIWoyx4_2),.clk(gclk));
	jdff dff_B_ygig0ASU9_2(.din(w_dff_B_3tLIWoyx4_2),.dout(w_dff_B_ygig0ASU9_2),.clk(gclk));
	jdff dff_B_VUJKNZ2w6_2(.din(w_dff_B_ygig0ASU9_2),.dout(w_dff_B_VUJKNZ2w6_2),.clk(gclk));
	jdff dff_B_1M8i8mw79_2(.din(w_dff_B_VUJKNZ2w6_2),.dout(w_dff_B_1M8i8mw79_2),.clk(gclk));
	jdff dff_A_TehYMzBl8_0(.dout(w_G53gat_0[0]),.din(w_dff_A_TehYMzBl8_0),.clk(gclk));
	jdff dff_A_Fn7Iv4Cx7_0(.dout(w_dff_A_TehYMzBl8_0),.din(w_dff_A_Fn7Iv4Cx7_0),.clk(gclk));
	jdff dff_A_HE2idggS8_0(.dout(w_dff_A_Fn7Iv4Cx7_0),.din(w_dff_A_HE2idggS8_0),.clk(gclk));
	jdff dff_A_yrQ2Xsar7_0(.dout(w_dff_A_HE2idggS8_0),.din(w_dff_A_yrQ2Xsar7_0),.clk(gclk));
	jdff dff_A_2vSLHRkS3_0(.dout(w_dff_A_yrQ2Xsar7_0),.din(w_dff_A_2vSLHRkS3_0),.clk(gclk));
	jdff dff_A_2iqLDpq24_0(.dout(w_dff_A_2vSLHRkS3_0),.din(w_dff_A_2iqLDpq24_0),.clk(gclk));
	jdff dff_A_OsNwv2H67_0(.dout(w_dff_A_2iqLDpq24_0),.din(w_dff_A_OsNwv2H67_0),.clk(gclk));
	jdff dff_A_KBGWrlXH4_0(.dout(w_dff_A_OsNwv2H67_0),.din(w_dff_A_KBGWrlXH4_0),.clk(gclk));
	jdff dff_A_2c9lvAsF9_0(.dout(w_dff_A_KBGWrlXH4_0),.din(w_dff_A_2c9lvAsF9_0),.clk(gclk));
	jdff dff_A_4C9omT440_0(.dout(w_dff_A_2c9lvAsF9_0),.din(w_dff_A_4C9omT440_0),.clk(gclk));
	jdff dff_A_9n1BOoKH9_0(.dout(w_dff_A_4C9omT440_0),.din(w_dff_A_9n1BOoKH9_0),.clk(gclk));
	jdff dff_A_HDcVbxuz4_0(.dout(w_dff_A_9n1BOoKH9_0),.din(w_dff_A_HDcVbxuz4_0),.clk(gclk));
	jdff dff_A_3z2JhcZs3_0(.dout(w_dff_A_HDcVbxuz4_0),.din(w_dff_A_3z2JhcZs3_0),.clk(gclk));
	jdff dff_A_FMq6roSG4_0(.dout(w_dff_A_3z2JhcZs3_0),.din(w_dff_A_FMq6roSG4_0),.clk(gclk));
	jdff dff_A_7U1ypy1a6_0(.dout(w_dff_A_FMq6roSG4_0),.din(w_dff_A_7U1ypy1a6_0),.clk(gclk));
	jdff dff_A_WpQyq9FU3_0(.dout(w_dff_A_7U1ypy1a6_0),.din(w_dff_A_WpQyq9FU3_0),.clk(gclk));
	jdff dff_A_0X4VuQBb3_0(.dout(w_dff_A_WpQyq9FU3_0),.din(w_dff_A_0X4VuQBb3_0),.clk(gclk));
	jdff dff_A_4KdI0J6J9_0(.dout(w_dff_A_0X4VuQBb3_0),.din(w_dff_A_4KdI0J6J9_0),.clk(gclk));
	jdff dff_A_NXAvvox10_0(.dout(w_dff_A_4KdI0J6J9_0),.din(w_dff_A_NXAvvox10_0),.clk(gclk));
	jdff dff_A_rA6U099P1_0(.dout(w_dff_A_NXAvvox10_0),.din(w_dff_A_rA6U099P1_0),.clk(gclk));
	jdff dff_A_iZIDpyIr3_0(.dout(w_n141_0[0]),.din(w_dff_A_iZIDpyIr3_0),.clk(gclk));
	jdff dff_B_NqK5r0uJ8_1(.din(n124),.dout(w_dff_B_NqK5r0uJ8_1),.clk(gclk));
	jdff dff_B_KqJio3Rg4_1(.din(n129),.dout(w_dff_B_KqJio3Rg4_1),.clk(gclk));
	jdff dff_B_pYwWI0Mm8_1(.din(w_dff_B_KqJio3Rg4_1),.dout(w_dff_B_pYwWI0Mm8_1),.clk(gclk));
	jdff dff_B_ka8Zgljp4_1(.din(w_dff_B_pYwWI0Mm8_1),.dout(w_dff_B_ka8Zgljp4_1),.clk(gclk));
	jdff dff_B_Fyq44NgT7_1(.din(w_dff_B_ka8Zgljp4_1),.dout(w_dff_B_Fyq44NgT7_1),.clk(gclk));
	jdff dff_B_ZdKfvdf30_1(.din(w_dff_B_Fyq44NgT7_1),.dout(w_dff_B_ZdKfvdf30_1),.clk(gclk));
	jdff dff_B_447HS49Y5_1(.din(w_dff_B_ZdKfvdf30_1),.dout(w_dff_B_447HS49Y5_1),.clk(gclk));
	jdff dff_B_vJDXMRpC0_1(.din(w_dff_B_447HS49Y5_1),.dout(w_dff_B_vJDXMRpC0_1),.clk(gclk));
	jdff dff_A_ukWOq8tP3_0(.dout(w_n131_0[0]),.din(w_dff_A_ukWOq8tP3_0),.clk(gclk));
	jdff dff_A_YYqfWhRq9_0(.dout(w_dff_A_ukWOq8tP3_0),.din(w_dff_A_YYqfWhRq9_0),.clk(gclk));
	jdff dff_A_CXIqUqbt1_0(.dout(w_dff_A_YYqfWhRq9_0),.din(w_dff_A_CXIqUqbt1_0),.clk(gclk));
	jdff dff_A_Rmm5znAV3_0(.dout(w_dff_A_CXIqUqbt1_0),.din(w_dff_A_Rmm5znAV3_0),.clk(gclk));
	jdff dff_A_iLzFQlOm1_0(.dout(w_dff_A_Rmm5znAV3_0),.din(w_dff_A_iLzFQlOm1_0),.clk(gclk));
	jdff dff_A_o9WJ33q89_0(.dout(w_dff_A_iLzFQlOm1_0),.din(w_dff_A_o9WJ33q89_0),.clk(gclk));
	jdff dff_A_fnI5mclx4_0(.dout(w_dff_A_o9WJ33q89_0),.din(w_dff_A_fnI5mclx4_0),.clk(gclk));
	jdff dff_A_DcKErPU78_0(.dout(w_n127_0[0]),.din(w_dff_A_DcKErPU78_0),.clk(gclk));
	jdff dff_A_oBfutAC63_0(.dout(w_dff_A_DcKErPU78_0),.din(w_dff_A_oBfutAC63_0),.clk(gclk));
	jdff dff_A_BVrgXk641_0(.dout(w_dff_A_oBfutAC63_0),.din(w_dff_A_BVrgXk641_0),.clk(gclk));
	jdff dff_A_GtwakSja0_0(.dout(w_dff_A_BVrgXk641_0),.din(w_dff_A_GtwakSja0_0),.clk(gclk));
	jdff dff_A_8y8N3Guq4_0(.dout(w_dff_A_GtwakSja0_0),.din(w_dff_A_8y8N3Guq4_0),.clk(gclk));
	jdff dff_A_j1MTcUuX6_0(.dout(w_dff_A_8y8N3Guq4_0),.din(w_dff_A_j1MTcUuX6_0),.clk(gclk));
	jdff dff_A_BTCMwIhv4_0(.dout(w_n125_0[0]),.din(w_dff_A_BTCMwIhv4_0),.clk(gclk));
	jdff dff_A_0vTTxGiD2_0(.dout(w_dff_A_BTCMwIhv4_0),.din(w_dff_A_0vTTxGiD2_0),.clk(gclk));
	jdff dff_A_YR1Vi4Ty3_0(.dout(w_dff_A_0vTTxGiD2_0),.din(w_dff_A_YR1Vi4Ty3_0),.clk(gclk));
	jdff dff_A_uIcAZ2sq8_0(.dout(w_dff_A_YR1Vi4Ty3_0),.din(w_dff_A_uIcAZ2sq8_0),.clk(gclk));
	jdff dff_A_sOSeQPg69_0(.dout(w_dff_A_uIcAZ2sq8_0),.din(w_dff_A_sOSeQPg69_0),.clk(gclk));
	jdff dff_B_ppkxjZnz4_2(.din(n125),.dout(w_dff_B_ppkxjZnz4_2),.clk(gclk));
	jdff dff_B_MvqA1pyZ4_2(.din(w_dff_B_ppkxjZnz4_2),.dout(w_dff_B_MvqA1pyZ4_2),.clk(gclk));
	jdff dff_B_nYPoKPki5_2(.din(w_dff_B_MvqA1pyZ4_2),.dout(w_dff_B_nYPoKPki5_2),.clk(gclk));
	jdff dff_B_Z878v3sO5_2(.din(w_dff_B_nYPoKPki5_2),.dout(w_dff_B_Z878v3sO5_2),.clk(gclk));
	jdff dff_B_bzuIyA295_2(.din(w_dff_B_Z878v3sO5_2),.dout(w_dff_B_bzuIyA295_2),.clk(gclk));
	jdff dff_B_NgIky2cZ8_2(.din(w_dff_B_bzuIyA295_2),.dout(w_dff_B_NgIky2cZ8_2),.clk(gclk));
	jdff dff_B_jlkyKIwC3_2(.din(w_dff_B_NgIky2cZ8_2),.dout(w_dff_B_jlkyKIwC3_2),.clk(gclk));
	jdff dff_A_t0fwS1Fi4_0(.dout(w_n123_0[0]),.din(w_dff_A_t0fwS1Fi4_0),.clk(gclk));
	jdff dff_A_eBAMU7Fu8_0(.dout(w_dff_A_t0fwS1Fi4_0),.din(w_dff_A_eBAMU7Fu8_0),.clk(gclk));
	jdff dff_A_qiARuj7l3_0(.dout(w_dff_A_eBAMU7Fu8_0),.din(w_dff_A_qiARuj7l3_0),.clk(gclk));
	jdff dff_A_Fx7tNW6C3_0(.dout(w_dff_A_qiARuj7l3_0),.din(w_dff_A_Fx7tNW6C3_0),.clk(gclk));
	jdff dff_A_KQeLt5oc7_0(.dout(w_dff_A_Fx7tNW6C3_0),.din(w_dff_A_KQeLt5oc7_0),.clk(gclk));
	jdff dff_A_yXhG2H8g8_0(.dout(w_dff_A_KQeLt5oc7_0),.din(w_dff_A_yXhG2H8g8_0),.clk(gclk));
	jdff dff_A_PNEJJfWC8_0(.dout(w_n121_0[0]),.din(w_dff_A_PNEJJfWC8_0),.clk(gclk));
	jdff dff_A_iXm02h9u9_0(.dout(w_dff_A_PNEJJfWC8_0),.din(w_dff_A_iXm02h9u9_0),.clk(gclk));
	jdff dff_A_ZJXP5Yfj7_0(.dout(w_dff_A_iXm02h9u9_0),.din(w_dff_A_ZJXP5Yfj7_0),.clk(gclk));
	jdff dff_A_UGzvVhbG3_0(.dout(w_dff_A_ZJXP5Yfj7_0),.din(w_dff_A_UGzvVhbG3_0),.clk(gclk));
	jdff dff_A_TNwq3u6B6_0(.dout(w_dff_A_UGzvVhbG3_0),.din(w_dff_A_TNwq3u6B6_0),.clk(gclk));
	jdff dff_B_IOWr197e6_2(.din(n121),.dout(w_dff_B_IOWr197e6_2),.clk(gclk));
	jdff dff_B_OkO0mU4i5_2(.din(w_dff_B_IOWr197e6_2),.dout(w_dff_B_OkO0mU4i5_2),.clk(gclk));
	jdff dff_B_JbGIOMH40_2(.din(w_dff_B_OkO0mU4i5_2),.dout(w_dff_B_JbGIOMH40_2),.clk(gclk));
	jdff dff_B_L9v1PK3V0_2(.din(w_dff_B_JbGIOMH40_2),.dout(w_dff_B_L9v1PK3V0_2),.clk(gclk));
	jdff dff_B_uW5GfRcs4_2(.din(w_dff_B_L9v1PK3V0_2),.dout(w_dff_B_uW5GfRcs4_2),.clk(gclk));
	jdff dff_B_s9Nl5gDw7_2(.din(w_dff_B_uW5GfRcs4_2),.dout(w_dff_B_s9Nl5gDw7_2),.clk(gclk));
	jdff dff_B_aWMZslLJ7_2(.din(w_dff_B_s9Nl5gDw7_2),.dout(w_dff_B_aWMZslLJ7_2),.clk(gclk));
	jdff dff_B_tFxJeg604_1(.din(n101),.dout(w_dff_B_tFxJeg604_1),.clk(gclk));
	jdff dff_B_kNpHvdbT1_0(.din(n114),.dout(w_dff_B_kNpHvdbT1_0),.clk(gclk));
	jdff dff_A_wK59n6K32_0(.dout(w_n113_0[0]),.din(w_dff_A_wK59n6K32_0),.clk(gclk));
	jdff dff_A_Fot6INnu1_0(.dout(w_dff_A_wK59n6K32_0),.din(w_dff_A_Fot6INnu1_0),.clk(gclk));
	jdff dff_A_m4w3asQE4_0(.dout(w_dff_A_Fot6INnu1_0),.din(w_dff_A_m4w3asQE4_0),.clk(gclk));
	jdff dff_A_ep4zO53T7_0(.dout(w_dff_A_m4w3asQE4_0),.din(w_dff_A_ep4zO53T7_0),.clk(gclk));
	jdff dff_A_jNCJ47D70_0(.dout(w_dff_A_ep4zO53T7_0),.din(w_dff_A_jNCJ47D70_0),.clk(gclk));
	jdff dff_A_jvJV2ZFZ2_0(.dout(w_dff_A_jNCJ47D70_0),.din(w_dff_A_jvJV2ZFZ2_0),.clk(gclk));
	jdff dff_A_q0VOqsmD5_0(.dout(w_n111_0[0]),.din(w_dff_A_q0VOqsmD5_0),.clk(gclk));
	jdff dff_A_oYvf3OG94_0(.dout(w_dff_A_q0VOqsmD5_0),.din(w_dff_A_oYvf3OG94_0),.clk(gclk));
	jdff dff_A_qPPMUy726_0(.dout(w_dff_A_oYvf3OG94_0),.din(w_dff_A_qPPMUy726_0),.clk(gclk));
	jdff dff_A_7Lu1vTHu9_0(.dout(w_dff_A_qPPMUy726_0),.din(w_dff_A_7Lu1vTHu9_0),.clk(gclk));
	jdff dff_A_mLXAvt4n0_0(.dout(w_dff_A_7Lu1vTHu9_0),.din(w_dff_A_mLXAvt4n0_0),.clk(gclk));
	jdff dff_B_b4dbHZai5_2(.din(n111),.dout(w_dff_B_b4dbHZai5_2),.clk(gclk));
	jdff dff_B_eurmNImh1_2(.din(w_dff_B_b4dbHZai5_2),.dout(w_dff_B_eurmNImh1_2),.clk(gclk));
	jdff dff_B_Yp7sK7kU0_2(.din(w_dff_B_eurmNImh1_2),.dout(w_dff_B_Yp7sK7kU0_2),.clk(gclk));
	jdff dff_B_FEn4Q8Yo7_2(.din(w_dff_B_Yp7sK7kU0_2),.dout(w_dff_B_FEn4Q8Yo7_2),.clk(gclk));
	jdff dff_B_TVEWEfFY6_2(.din(w_dff_B_FEn4Q8Yo7_2),.dout(w_dff_B_TVEWEfFY6_2),.clk(gclk));
	jdff dff_B_MJmaSI9H1_2(.din(w_dff_B_TVEWEfFY6_2),.dout(w_dff_B_MJmaSI9H1_2),.clk(gclk));
	jdff dff_B_kRvHPEm09_2(.din(w_dff_B_MJmaSI9H1_2),.dout(w_dff_B_kRvHPEm09_2),.clk(gclk));
	jdff dff_A_iJzAqBOW0_0(.dout(w_n108_0[0]),.din(w_dff_A_iJzAqBOW0_0),.clk(gclk));
	jdff dff_A_UBAr06oW3_0(.dout(w_dff_A_iJzAqBOW0_0),.din(w_dff_A_UBAr06oW3_0),.clk(gclk));
	jdff dff_A_zLWEIj8B8_0(.dout(w_dff_A_UBAr06oW3_0),.din(w_dff_A_zLWEIj8B8_0),.clk(gclk));
	jdff dff_A_19qyuNKG3_0(.dout(w_dff_A_zLWEIj8B8_0),.din(w_dff_A_19qyuNKG3_0),.clk(gclk));
	jdff dff_A_eMNfuXmO1_0(.dout(w_dff_A_19qyuNKG3_0),.din(w_dff_A_eMNfuXmO1_0),.clk(gclk));
	jdff dff_A_XMNTUH095_0(.dout(w_dff_A_eMNfuXmO1_0),.din(w_dff_A_XMNTUH095_0),.clk(gclk));
	jdff dff_A_hB2DIHX84_0(.dout(w_n106_0[0]),.din(w_dff_A_hB2DIHX84_0),.clk(gclk));
	jdff dff_A_tUk0OBpo4_0(.dout(w_dff_A_hB2DIHX84_0),.din(w_dff_A_tUk0OBpo4_0),.clk(gclk));
	jdff dff_A_QdaKPHcP5_0(.dout(w_dff_A_tUk0OBpo4_0),.din(w_dff_A_QdaKPHcP5_0),.clk(gclk));
	jdff dff_A_Wkzy1KtS0_0(.dout(w_dff_A_QdaKPHcP5_0),.din(w_dff_A_Wkzy1KtS0_0),.clk(gclk));
	jdff dff_A_V88cwFC23_0(.dout(w_dff_A_Wkzy1KtS0_0),.din(w_dff_A_V88cwFC23_0),.clk(gclk));
	jdff dff_B_dA3SBpJ68_2(.din(n106),.dout(w_dff_B_dA3SBpJ68_2),.clk(gclk));
	jdff dff_B_G1ZeSt958_2(.din(w_dff_B_dA3SBpJ68_2),.dout(w_dff_B_G1ZeSt958_2),.clk(gclk));
	jdff dff_B_3aBa0O241_2(.din(w_dff_B_G1ZeSt958_2),.dout(w_dff_B_3aBa0O241_2),.clk(gclk));
	jdff dff_B_Wus2GaKB4_2(.din(w_dff_B_3aBa0O241_2),.dout(w_dff_B_Wus2GaKB4_2),.clk(gclk));
	jdff dff_B_5oAjXXeq8_2(.din(w_dff_B_Wus2GaKB4_2),.dout(w_dff_B_5oAjXXeq8_2),.clk(gclk));
	jdff dff_B_U9Vb01T34_2(.din(w_dff_B_5oAjXXeq8_2),.dout(w_dff_B_U9Vb01T34_2),.clk(gclk));
	jdff dff_B_93DoIoKW3_2(.din(w_dff_B_U9Vb01T34_2),.dout(w_dff_B_93DoIoKW3_2),.clk(gclk));
	jdff dff_B_4Hy0jiv52_1(.din(n97),.dout(w_dff_B_4Hy0jiv52_1),.clk(gclk));
	jdff dff_B_ecmWlFWi7_1(.din(w_dff_B_4Hy0jiv52_1),.dout(w_dff_B_ecmWlFWi7_1),.clk(gclk));
	jdff dff_B_hhc665Rx5_1(.din(w_dff_B_ecmWlFWi7_1),.dout(w_dff_B_hhc665Rx5_1),.clk(gclk));
	jdff dff_B_AnQhNxo99_1(.din(w_dff_B_hhc665Rx5_1),.dout(w_dff_B_AnQhNxo99_1),.clk(gclk));
	jdff dff_B_DQXU00sF7_1(.din(w_dff_B_AnQhNxo99_1),.dout(w_dff_B_DQXU00sF7_1),.clk(gclk));
	jdff dff_B_djL2IWfi4_1(.din(w_dff_B_DQXU00sF7_1),.dout(w_dff_B_djL2IWfi4_1),.clk(gclk));
	jdff dff_B_awY5TtCk8_1(.din(w_dff_B_djL2IWfi4_1),.dout(w_dff_B_awY5TtCk8_1),.clk(gclk));
	jdff dff_A_0gGFO1si5_0(.dout(w_n95_0[0]),.din(w_dff_A_0gGFO1si5_0),.clk(gclk));
	jdff dff_A_w5VXco6n2_0(.dout(w_dff_A_0gGFO1si5_0),.din(w_dff_A_w5VXco6n2_0),.clk(gclk));
	jdff dff_A_O5BubKlF6_0(.dout(w_dff_A_w5VXco6n2_0),.din(w_dff_A_O5BubKlF6_0),.clk(gclk));
	jdff dff_A_uvZBCxhN2_0(.dout(w_dff_A_O5BubKlF6_0),.din(w_dff_A_uvZBCxhN2_0),.clk(gclk));
	jdff dff_A_IbJJYA8K7_0(.dout(w_dff_A_uvZBCxhN2_0),.din(w_dff_A_IbJJYA8K7_0),.clk(gclk));
	jdff dff_A_cRMZYc3B1_0(.dout(w_dff_A_IbJJYA8K7_0),.din(w_dff_A_cRMZYc3B1_0),.clk(gclk));
	jdff dff_A_dAdDwizU1_0(.dout(w_n70_0[0]),.din(w_dff_A_dAdDwizU1_0),.clk(gclk));
	jdff dff_A_cIgXDEL30_0(.dout(w_dff_A_dAdDwizU1_0),.din(w_dff_A_cIgXDEL30_0),.clk(gclk));
	jdff dff_A_1e8abMSn7_0(.dout(w_dff_A_cIgXDEL30_0),.din(w_dff_A_1e8abMSn7_0),.clk(gclk));
	jdff dff_A_yCXfxgGn8_0(.dout(w_dff_A_1e8abMSn7_0),.din(w_dff_A_yCXfxgGn8_0),.clk(gclk));
	jdff dff_A_dM4HeqPw5_0(.dout(w_dff_A_yCXfxgGn8_0),.din(w_dff_A_dM4HeqPw5_0),.clk(gclk));
	jdff dff_B_7S11WjdZ4_2(.din(n70),.dout(w_dff_B_7S11WjdZ4_2),.clk(gclk));
	jdff dff_B_CXrh2OYW4_2(.din(w_dff_B_7S11WjdZ4_2),.dout(w_dff_B_CXrh2OYW4_2),.clk(gclk));
	jdff dff_B_6Cbbxs066_2(.din(w_dff_B_CXrh2OYW4_2),.dout(w_dff_B_6Cbbxs066_2),.clk(gclk));
	jdff dff_B_nZFvdqNt7_2(.din(w_dff_B_6Cbbxs066_2),.dout(w_dff_B_nZFvdqNt7_2),.clk(gclk));
	jdff dff_B_ubgIpsNP6_2(.din(w_dff_B_nZFvdqNt7_2),.dout(w_dff_B_ubgIpsNP6_2),.clk(gclk));
	jdff dff_B_WMzIhlvR0_2(.din(w_dff_B_ubgIpsNP6_2),.dout(w_dff_B_WMzIhlvR0_2),.clk(gclk));
	jdff dff_B_du5n4KHy9_2(.din(w_dff_B_WMzIhlvR0_2),.dout(w_dff_B_du5n4KHy9_2),.clk(gclk));
	jdff dff_A_HsvVj9Sr9_1(.dout(w_G105gat_0[1]),.din(w_dff_A_HsvVj9Sr9_1),.clk(gclk));
	jdff dff_A_GfVaUSdR8_1(.dout(w_dff_A_HsvVj9Sr9_1),.din(w_dff_A_GfVaUSdR8_1),.clk(gclk));
	jdff dff_A_TazNC8XV7_1(.dout(w_dff_A_GfVaUSdR8_1),.din(w_dff_A_TazNC8XV7_1),.clk(gclk));
	jdff dff_A_QCoJQIcB1_1(.dout(w_dff_A_TazNC8XV7_1),.din(w_dff_A_QCoJQIcB1_1),.clk(gclk));
	jdff dff_A_efO9Ivv29_1(.dout(w_dff_A_QCoJQIcB1_1),.din(w_dff_A_efO9Ivv29_1),.clk(gclk));
	jdff dff_A_TLOHSE780_1(.dout(w_dff_A_efO9Ivv29_1),.din(w_dff_A_TLOHSE780_1),.clk(gclk));
	jdff dff_A_gevF5jCx6_1(.dout(w_dff_A_TLOHSE780_1),.din(w_dff_A_gevF5jCx6_1),.clk(gclk));
	jdff dff_A_W2xbkyoo0_1(.dout(w_dff_A_gevF5jCx6_1),.din(w_dff_A_W2xbkyoo0_1),.clk(gclk));
	jdff dff_A_kPjP12Jp9_1(.dout(w_dff_A_W2xbkyoo0_1),.din(w_dff_A_kPjP12Jp9_1),.clk(gclk));
	jdff dff_A_DrfipQrw9_1(.dout(w_dff_A_kPjP12Jp9_1),.din(w_dff_A_DrfipQrw9_1),.clk(gclk));
	jdff dff_A_KAZwzF9R4_1(.dout(w_dff_A_DrfipQrw9_1),.din(w_dff_A_KAZwzF9R4_1),.clk(gclk));
	jdff dff_A_qrbowgNY3_1(.dout(w_dff_A_KAZwzF9R4_1),.din(w_dff_A_qrbowgNY3_1),.clk(gclk));
	jdff dff_A_RC5qWVzk6_1(.dout(w_dff_A_qrbowgNY3_1),.din(w_dff_A_RC5qWVzk6_1),.clk(gclk));
	jdff dff_A_SbUyfcqN9_1(.dout(w_dff_A_RC5qWVzk6_1),.din(w_dff_A_SbUyfcqN9_1),.clk(gclk));
	jdff dff_A_UzWk0GRm9_1(.dout(w_dff_A_SbUyfcqN9_1),.din(w_dff_A_UzWk0GRm9_1),.clk(gclk));
	jdff dff_A_rN8koomI5_0(.dout(w_n200_0[0]),.din(w_dff_A_rN8koomI5_0),.clk(gclk));
	jdff dff_A_PzEU658U9_0(.dout(w_dff_A_rN8koomI5_0),.din(w_dff_A_PzEU658U9_0),.clk(gclk));
	jdff dff_A_mOfbwand3_0(.dout(w_dff_A_PzEU658U9_0),.din(w_dff_A_mOfbwand3_0),.clk(gclk));
	jdff dff_A_AkUplPZz5_0(.dout(w_dff_A_mOfbwand3_0),.din(w_dff_A_AkUplPZz5_0),.clk(gclk));
	jdff dff_A_UkbINEYs0_0(.dout(w_dff_A_AkUplPZz5_0),.din(w_dff_A_UkbINEYs0_0),.clk(gclk));
	jdff dff_B_i0JwDmKu3_2(.din(n200),.dout(w_dff_B_i0JwDmKu3_2),.clk(gclk));
	jdff dff_B_nkkH4yCR3_2(.din(w_dff_B_i0JwDmKu3_2),.dout(w_dff_B_nkkH4yCR3_2),.clk(gclk));
	jdff dff_B_4zpay2Qy5_2(.din(w_dff_B_nkkH4yCR3_2),.dout(w_dff_B_4zpay2Qy5_2),.clk(gclk));
	jdff dff_B_1gHkALnk9_2(.din(w_dff_B_4zpay2Qy5_2),.dout(w_dff_B_1gHkALnk9_2),.clk(gclk));
	jdff dff_B_cqrnNfOR2_2(.din(w_dff_B_1gHkALnk9_2),.dout(w_dff_B_cqrnNfOR2_2),.clk(gclk));
	jdff dff_B_P2897u1Q3_2(.din(w_dff_B_cqrnNfOR2_2),.dout(w_dff_B_P2897u1Q3_2),.clk(gclk));
	jdff dff_B_IaRzRIba6_2(.din(w_dff_B_P2897u1Q3_2),.dout(w_dff_B_IaRzRIba6_2),.clk(gclk));
	jdff dff_B_Q13EOOKL1_2(.din(w_dff_B_IaRzRIba6_2),.dout(w_dff_B_Q13EOOKL1_2),.clk(gclk));
	jdff dff_B_1GMVD8i19_2(.din(w_dff_B_Q13EOOKL1_2),.dout(w_dff_B_1GMVD8i19_2),.clk(gclk));
	jdff dff_B_J8W4Nmss9_2(.din(w_dff_B_1GMVD8i19_2),.dout(w_dff_B_J8W4Nmss9_2),.clk(gclk));
	jdff dff_B_hbK7XanY0_2(.din(w_dff_B_J8W4Nmss9_2),.dout(w_dff_B_hbK7XanY0_2),.clk(gclk));
	jdff dff_B_180tNT1g1_2(.din(w_dff_B_hbK7XanY0_2),.dout(w_dff_B_180tNT1g1_2),.clk(gclk));
	jdff dff_B_KfyEUUMm8_2(.din(w_dff_B_180tNT1g1_2),.dout(w_dff_B_KfyEUUMm8_2),.clk(gclk));
	jdff dff_B_jWf3GUkZ9_2(.din(w_dff_B_KfyEUUMm8_2),.dout(w_dff_B_jWf3GUkZ9_2),.clk(gclk));
	jdff dff_A_QD8Sn8xn6_0(.dout(w_G79gat_0[0]),.din(w_dff_A_QD8Sn8xn6_0),.clk(gclk));
	jdff dff_A_hnXEFaRo3_0(.dout(w_dff_A_QD8Sn8xn6_0),.din(w_dff_A_hnXEFaRo3_0),.clk(gclk));
	jdff dff_A_ubLSppHX7_0(.dout(w_dff_A_hnXEFaRo3_0),.din(w_dff_A_ubLSppHX7_0),.clk(gclk));
	jdff dff_A_fChuHLr85_0(.dout(w_dff_A_ubLSppHX7_0),.din(w_dff_A_fChuHLr85_0),.clk(gclk));
	jdff dff_A_p5a7Vwgh8_0(.dout(w_dff_A_fChuHLr85_0),.din(w_dff_A_p5a7Vwgh8_0),.clk(gclk));
	jdff dff_A_gj7DxBKd2_0(.dout(w_dff_A_p5a7Vwgh8_0),.din(w_dff_A_gj7DxBKd2_0),.clk(gclk));
	jdff dff_A_xuEWtplg7_0(.dout(w_dff_A_gj7DxBKd2_0),.din(w_dff_A_xuEWtplg7_0),.clk(gclk));
	jdff dff_A_gHCh00wX9_0(.dout(w_dff_A_xuEWtplg7_0),.din(w_dff_A_gHCh00wX9_0),.clk(gclk));
	jdff dff_A_56IQBdFD6_0(.dout(w_dff_A_gHCh00wX9_0),.din(w_dff_A_56IQBdFD6_0),.clk(gclk));
	jdff dff_A_Ntc4VIEX7_0(.dout(w_dff_A_56IQBdFD6_0),.din(w_dff_A_Ntc4VIEX7_0),.clk(gclk));
	jdff dff_A_UCyxuw599_0(.dout(w_dff_A_Ntc4VIEX7_0),.din(w_dff_A_UCyxuw599_0),.clk(gclk));
	jdff dff_A_sPIJUNzg2_0(.dout(w_dff_A_UCyxuw599_0),.din(w_dff_A_sPIJUNzg2_0),.clk(gclk));
	jdff dff_A_fwbZKcqG5_0(.dout(w_dff_A_sPIJUNzg2_0),.din(w_dff_A_fwbZKcqG5_0),.clk(gclk));
	jdff dff_A_5Rzh4lej4_0(.dout(w_dff_A_fwbZKcqG5_0),.din(w_dff_A_5Rzh4lej4_0),.clk(gclk));
	jdff dff_A_PkvW4NuJ6_0(.dout(w_dff_A_5Rzh4lej4_0),.din(w_dff_A_PkvW4NuJ6_0),.clk(gclk));
	jdff dff_A_IQsc8pdn6_0(.dout(w_n202_0[0]),.din(w_dff_A_IQsc8pdn6_0),.clk(gclk));
	jdff dff_A_qx6bSRxL0_0(.dout(w_dff_A_IQsc8pdn6_0),.din(w_dff_A_qx6bSRxL0_0),.clk(gclk));
	jdff dff_A_1ZnpfZau8_0(.dout(w_dff_A_qx6bSRxL0_0),.din(w_dff_A_1ZnpfZau8_0),.clk(gclk));
	jdff dff_A_eYlnGbmT1_0(.dout(w_dff_A_1ZnpfZau8_0),.din(w_dff_A_eYlnGbmT1_0),.clk(gclk));
	jdff dff_A_YZFvLYFV8_0(.dout(w_dff_A_eYlnGbmT1_0),.din(w_dff_A_YZFvLYFV8_0),.clk(gclk));
	jdff dff_A_4ovGi05V3_0(.dout(w_dff_A_YZFvLYFV8_0),.din(w_dff_A_4ovGi05V3_0),.clk(gclk));
	jdff dff_B_NQ6qWZcn7_1(.din(n168),.dout(w_dff_B_NQ6qWZcn7_1),.clk(gclk));
	jdff dff_B_MGjLvvx48_1(.din(n171),.dout(w_dff_B_MGjLvvx48_1),.clk(gclk));
	jdff dff_A_azkryNac6_0(.dout(w_G47gat_0[0]),.din(w_dff_A_azkryNac6_0),.clk(gclk));
	jdff dff_A_NU4en6Er5_0(.dout(w_dff_A_azkryNac6_0),.din(w_dff_A_NU4en6Er5_0),.clk(gclk));
	jdff dff_A_4Obfc4wf3_0(.dout(w_dff_A_NU4en6Er5_0),.din(w_dff_A_4Obfc4wf3_0),.clk(gclk));
	jdff dff_A_TwTZHlF69_0(.dout(w_dff_A_4Obfc4wf3_0),.din(w_dff_A_TwTZHlF69_0),.clk(gclk));
	jdff dff_A_jyiK3bZm1_0(.dout(w_dff_A_TwTZHlF69_0),.din(w_dff_A_jyiK3bZm1_0),.clk(gclk));
	jdff dff_A_hGZTRHHC4_0(.dout(w_dff_A_jyiK3bZm1_0),.din(w_dff_A_hGZTRHHC4_0),.clk(gclk));
	jdff dff_A_CphBLeP64_0(.dout(w_dff_A_hGZTRHHC4_0),.din(w_dff_A_CphBLeP64_0),.clk(gclk));
	jdff dff_A_6LwEWqdP7_0(.dout(w_dff_A_CphBLeP64_0),.din(w_dff_A_6LwEWqdP7_0),.clk(gclk));
	jdff dff_A_d3psj1Pa9_1(.dout(w_G47gat_0[1]),.din(w_dff_A_d3psj1Pa9_1),.clk(gclk));
	jdff dff_A_jn0pbfpr1_1(.dout(w_dff_A_d3psj1Pa9_1),.din(w_dff_A_jn0pbfpr1_1),.clk(gclk));
	jdff dff_A_G66HetqF0_1(.dout(w_dff_A_jn0pbfpr1_1),.din(w_dff_A_G66HetqF0_1),.clk(gclk));
	jdff dff_A_2DcnsPvc6_1(.dout(w_dff_A_G66HetqF0_1),.din(w_dff_A_2DcnsPvc6_1),.clk(gclk));
	jdff dff_A_LL1Dh6kU8_1(.dout(w_dff_A_2DcnsPvc6_1),.din(w_dff_A_LL1Dh6kU8_1),.clk(gclk));
	jdff dff_A_my1kK3pL0_1(.dout(w_dff_A_LL1Dh6kU8_1),.din(w_dff_A_my1kK3pL0_1),.clk(gclk));
	jdff dff_A_ofCS9CID6_1(.dout(w_dff_A_my1kK3pL0_1),.din(w_dff_A_ofCS9CID6_1),.clk(gclk));
	jdff dff_A_T6pXnsGV7_1(.dout(w_dff_A_ofCS9CID6_1),.din(w_dff_A_T6pXnsGV7_1),.clk(gclk));
	jdff dff_A_AH4PL5i43_1(.dout(w_dff_A_T6pXnsGV7_1),.din(w_dff_A_AH4PL5i43_1),.clk(gclk));
	jdff dff_A_i4JLvFh20_1(.dout(w_dff_A_AH4PL5i43_1),.din(w_dff_A_i4JLvFh20_1),.clk(gclk));
	jdff dff_A_m22eKOdL3_1(.dout(w_dff_A_i4JLvFh20_1),.din(w_dff_A_m22eKOdL3_1),.clk(gclk));
	jdff dff_A_ETi4jrU66_1(.dout(w_dff_A_m22eKOdL3_1),.din(w_dff_A_ETi4jrU66_1),.clk(gclk));
	jdff dff_A_JLloTRJ83_1(.dout(w_dff_A_ETi4jrU66_1),.din(w_dff_A_JLloTRJ83_1),.clk(gclk));
	jdff dff_A_gnRA4fNu1_0(.dout(w_n173_0[0]),.din(w_dff_A_gnRA4fNu1_0),.clk(gclk));
	jdff dff_A_7cwWfYfj1_0(.dout(w_dff_A_gnRA4fNu1_0),.din(w_dff_A_7cwWfYfj1_0),.clk(gclk));
	jdff dff_A_tF4grip08_0(.dout(w_dff_A_7cwWfYfj1_0),.din(w_dff_A_tF4grip08_0),.clk(gclk));
	jdff dff_A_yEMOP4rc7_0(.dout(w_dff_A_tF4grip08_0),.din(w_dff_A_yEMOP4rc7_0),.clk(gclk));
	jdff dff_A_7o0mONMx5_0(.dout(w_dff_A_yEMOP4rc7_0),.din(w_dff_A_7o0mONMx5_0),.clk(gclk));
	jdff dff_A_Z6xDi7py5_0(.dout(w_dff_A_7o0mONMx5_0),.din(w_dff_A_Z6xDi7py5_0),.clk(gclk));
	jdff dff_A_keSjFFSW4_0(.dout(w_G8gat_0[0]),.din(w_dff_A_keSjFFSW4_0),.clk(gclk));
	jdff dff_A_FmMZyJLw4_0(.dout(w_dff_A_keSjFFSW4_0),.din(w_dff_A_FmMZyJLw4_0),.clk(gclk));
	jdff dff_A_GQSUqkXk1_0(.dout(w_dff_A_FmMZyJLw4_0),.din(w_dff_A_GQSUqkXk1_0),.clk(gclk));
	jdff dff_A_0GQ949Hm5_0(.dout(w_dff_A_GQSUqkXk1_0),.din(w_dff_A_0GQ949Hm5_0),.clk(gclk));
	jdff dff_A_5LXmG0EF7_0(.dout(w_dff_A_0GQ949Hm5_0),.din(w_dff_A_5LXmG0EF7_0),.clk(gclk));
	jdff dff_A_OkcAVjAQ3_0(.dout(w_dff_A_5LXmG0EF7_0),.din(w_dff_A_OkcAVjAQ3_0),.clk(gclk));
	jdff dff_A_7ZIDyrBl4_0(.dout(w_dff_A_OkcAVjAQ3_0),.din(w_dff_A_7ZIDyrBl4_0),.clk(gclk));
	jdff dff_A_tJnszgV80_0(.dout(w_dff_A_7ZIDyrBl4_0),.din(w_dff_A_tJnszgV80_0),.clk(gclk));
	jdff dff_A_5K6pCmpL2_0(.dout(w_dff_A_tJnszgV80_0),.din(w_dff_A_5K6pCmpL2_0),.clk(gclk));
	jdff dff_A_e9MGPYqX1_0(.dout(w_dff_A_5K6pCmpL2_0),.din(w_dff_A_e9MGPYqX1_0),.clk(gclk));
	jdff dff_A_MP349w4b3_0(.dout(w_dff_A_e9MGPYqX1_0),.din(w_dff_A_MP349w4b3_0),.clk(gclk));
	jdff dff_A_F67Yb6UX5_0(.dout(w_dff_A_MP349w4b3_0),.din(w_dff_A_F67Yb6UX5_0),.clk(gclk));
	jdff dff_A_Le75QP4r4_0(.dout(w_dff_A_F67Yb6UX5_0),.din(w_dff_A_Le75QP4r4_0),.clk(gclk));
	jdff dff_A_d0c6zVx68_1(.dout(w_G8gat_0[1]),.din(w_dff_A_d0c6zVx68_1),.clk(gclk));
	jdff dff_A_7n9lGIWn3_1(.dout(w_dff_A_d0c6zVx68_1),.din(w_dff_A_7n9lGIWn3_1),.clk(gclk));
	jdff dff_A_fBde5rFb6_1(.dout(w_dff_A_7n9lGIWn3_1),.din(w_dff_A_fBde5rFb6_1),.clk(gclk));
	jdff dff_A_I8xSQwyx5_1(.dout(w_dff_A_fBde5rFb6_1),.din(w_dff_A_I8xSQwyx5_1),.clk(gclk));
	jdff dff_A_sDy1bD010_1(.dout(w_dff_A_I8xSQwyx5_1),.din(w_dff_A_sDy1bD010_1),.clk(gclk));
	jdff dff_A_8JQYqsyZ2_1(.dout(w_dff_A_sDy1bD010_1),.din(w_dff_A_8JQYqsyZ2_1),.clk(gclk));
	jdff dff_A_zm39boY64_1(.dout(w_dff_A_8JQYqsyZ2_1),.din(w_dff_A_zm39boY64_1),.clk(gclk));
	jdff dff_A_tttNuUrm6_1(.dout(w_dff_A_zm39boY64_1),.din(w_dff_A_tttNuUrm6_1),.clk(gclk));
	jdff dff_A_Bn1RDwuN2_0(.dout(w_n170_0[0]),.din(w_dff_A_Bn1RDwuN2_0),.clk(gclk));
	jdff dff_A_0hA8ov3Z6_0(.dout(w_dff_A_Bn1RDwuN2_0),.din(w_dff_A_0hA8ov3Z6_0),.clk(gclk));
	jdff dff_A_4UeZc7LN8_0(.dout(w_dff_A_0hA8ov3Z6_0),.din(w_dff_A_4UeZc7LN8_0),.clk(gclk));
	jdff dff_A_1XKNu4IG7_0(.dout(w_dff_A_4UeZc7LN8_0),.din(w_dff_A_1XKNu4IG7_0),.clk(gclk));
	jdff dff_A_KphDdd8P5_0(.dout(w_dff_A_1XKNu4IG7_0),.din(w_dff_A_KphDdd8P5_0),.clk(gclk));
	jdff dff_A_HOZpH2xk1_0(.dout(w_dff_A_KphDdd8P5_0),.din(w_dff_A_HOZpH2xk1_0),.clk(gclk));
	jdff dff_A_wj4A0kFJ0_0(.dout(w_G86gat_0[0]),.din(w_dff_A_wj4A0kFJ0_0),.clk(gclk));
	jdff dff_A_lTb9FXNb9_0(.dout(w_dff_A_wj4A0kFJ0_0),.din(w_dff_A_lTb9FXNb9_0),.clk(gclk));
	jdff dff_A_yzggL9pr8_0(.dout(w_dff_A_lTb9FXNb9_0),.din(w_dff_A_yzggL9pr8_0),.clk(gclk));
	jdff dff_A_zhixABwN9_0(.dout(w_dff_A_yzggL9pr8_0),.din(w_dff_A_zhixABwN9_0),.clk(gclk));
	jdff dff_A_8r4FoLHq8_0(.dout(w_dff_A_zhixABwN9_0),.din(w_dff_A_8r4FoLHq8_0),.clk(gclk));
	jdff dff_A_HTtol3Ui3_0(.dout(w_dff_A_8r4FoLHq8_0),.din(w_dff_A_HTtol3Ui3_0),.clk(gclk));
	jdff dff_A_Fw3USXt87_0(.dout(w_dff_A_HTtol3Ui3_0),.din(w_dff_A_Fw3USXt87_0),.clk(gclk));
	jdff dff_A_oYqhOt2F2_0(.dout(w_dff_A_Fw3USXt87_0),.din(w_dff_A_oYqhOt2F2_0),.clk(gclk));
	jdff dff_A_H7KaN3Pn9_0(.dout(w_dff_A_oYqhOt2F2_0),.din(w_dff_A_H7KaN3Pn9_0),.clk(gclk));
	jdff dff_A_G3oHU4zl8_0(.dout(w_dff_A_H7KaN3Pn9_0),.din(w_dff_A_G3oHU4zl8_0),.clk(gclk));
	jdff dff_A_xGqxvpuB2_0(.dout(w_dff_A_G3oHU4zl8_0),.din(w_dff_A_xGqxvpuB2_0),.clk(gclk));
	jdff dff_A_YPeFjJbQ3_0(.dout(w_dff_A_xGqxvpuB2_0),.din(w_dff_A_YPeFjJbQ3_0),.clk(gclk));
	jdff dff_A_8NTOvryK9_0(.dout(w_dff_A_YPeFjJbQ3_0),.din(w_dff_A_8NTOvryK9_0),.clk(gclk));
	jdff dff_A_Wj9TiAki9_1(.dout(w_G86gat_0[1]),.din(w_dff_A_Wj9TiAki9_1),.clk(gclk));
	jdff dff_A_IxTDQcvy2_1(.dout(w_dff_A_Wj9TiAki9_1),.din(w_dff_A_IxTDQcvy2_1),.clk(gclk));
	jdff dff_A_0R3kRCOl1_1(.dout(w_dff_A_IxTDQcvy2_1),.din(w_dff_A_0R3kRCOl1_1),.clk(gclk));
	jdff dff_A_h5QL0kCJ5_1(.dout(w_dff_A_0R3kRCOl1_1),.din(w_dff_A_h5QL0kCJ5_1),.clk(gclk));
	jdff dff_A_LYIfWeTe0_1(.dout(w_dff_A_h5QL0kCJ5_1),.din(w_dff_A_LYIfWeTe0_1),.clk(gclk));
	jdff dff_A_ox9oGVPL0_1(.dout(w_dff_A_LYIfWeTe0_1),.din(w_dff_A_ox9oGVPL0_1),.clk(gclk));
	jdff dff_A_n0dbXPoS4_1(.dout(w_dff_A_ox9oGVPL0_1),.din(w_dff_A_n0dbXPoS4_1),.clk(gclk));
	jdff dff_A_4RTxeQTv8_1(.dout(w_dff_A_n0dbXPoS4_1),.din(w_dff_A_4RTxeQTv8_1),.clk(gclk));
	jdff dff_A_CMuI8L6j7_1(.dout(w_n120_0[1]),.din(w_dff_A_CMuI8L6j7_1),.clk(gclk));
	jdff dff_A_G9lrbznW0_1(.dout(w_dff_A_CMuI8L6j7_1),.din(w_dff_A_G9lrbznW0_1),.clk(gclk));
	jdff dff_A_KeFNm4pW6_1(.dout(w_n119_0[1]),.din(w_dff_A_KeFNm4pW6_1),.clk(gclk));
	jdff dff_A_kC62ZcDW3_1(.dout(w_dff_A_KeFNm4pW6_1),.din(w_dff_A_kC62ZcDW3_1),.clk(gclk));
	jdff dff_A_jcY5vvGb8_1(.dout(w_dff_A_kC62ZcDW3_1),.din(w_dff_A_jcY5vvGb8_1),.clk(gclk));
	jdff dff_A_wRopOt5L7_1(.dout(w_dff_A_jcY5vvGb8_1),.din(w_dff_A_wRopOt5L7_1),.clk(gclk));
	jdff dff_A_22tN93cK1_1(.dout(w_dff_A_wRopOt5L7_1),.din(w_dff_A_22tN93cK1_1),.clk(gclk));
	jdff dff_A_us47lpq66_1(.dout(w_dff_A_22tN93cK1_1),.din(w_dff_A_us47lpq66_1),.clk(gclk));
	jdff dff_A_AC2CS2hU4_0(.dout(w_n117_0[0]),.din(w_dff_A_AC2CS2hU4_0),.clk(gclk));
	jdff dff_A_shvZ5KCl4_0(.dout(w_dff_A_AC2CS2hU4_0),.din(w_dff_A_shvZ5KCl4_0),.clk(gclk));
	jdff dff_A_yPTK2SJA6_0(.dout(w_dff_A_shvZ5KCl4_0),.din(w_dff_A_yPTK2SJA6_0),.clk(gclk));
	jdff dff_A_BUk5ewy63_0(.dout(w_dff_A_yPTK2SJA6_0),.din(w_dff_A_BUk5ewy63_0),.clk(gclk));
	jdff dff_A_i5tkwe6P9_0(.dout(w_dff_A_BUk5ewy63_0),.din(w_dff_A_i5tkwe6P9_0),.clk(gclk));
	jdff dff_B_iEHWkATf7_2(.din(n117),.dout(w_dff_B_iEHWkATf7_2),.clk(gclk));
	jdff dff_B_eWavxSBs5_2(.din(w_dff_B_iEHWkATf7_2),.dout(w_dff_B_eWavxSBs5_2),.clk(gclk));
	jdff dff_B_GVnRsVxf0_2(.din(w_dff_B_eWavxSBs5_2),.dout(w_dff_B_GVnRsVxf0_2),.clk(gclk));
	jdff dff_B_flLocZ0f0_2(.din(w_dff_B_GVnRsVxf0_2),.dout(w_dff_B_flLocZ0f0_2),.clk(gclk));
	jdff dff_B_8H0gQXti6_2(.din(w_dff_B_flLocZ0f0_2),.dout(w_dff_B_8H0gQXti6_2),.clk(gclk));
	jdff dff_B_4MgC1ltu4_2(.din(w_dff_B_8H0gQXti6_2),.dout(w_dff_B_4MgC1ltu4_2),.clk(gclk));
	jdff dff_B_A00qhiij1_2(.din(w_dff_B_4MgC1ltu4_2),.dout(w_dff_B_A00qhiij1_2),.clk(gclk));
	jdff dff_A_lolXuHU57_0(.dout(w_G60gat_0[0]),.din(w_dff_A_lolXuHU57_0),.clk(gclk));
	jdff dff_A_druw62o49_0(.dout(w_dff_A_lolXuHU57_0),.din(w_dff_A_druw62o49_0),.clk(gclk));
	jdff dff_A_EWhHvAiG8_0(.dout(w_dff_A_druw62o49_0),.din(w_dff_A_EWhHvAiG8_0),.clk(gclk));
	jdff dff_A_Vjp4mi7i3_0(.dout(w_dff_A_EWhHvAiG8_0),.din(w_dff_A_Vjp4mi7i3_0),.clk(gclk));
	jdff dff_A_uHBZwbJl4_0(.dout(w_dff_A_Vjp4mi7i3_0),.din(w_dff_A_uHBZwbJl4_0),.clk(gclk));
	jdff dff_A_7h7Fu2Q37_0(.dout(w_dff_A_uHBZwbJl4_0),.din(w_dff_A_7h7Fu2Q37_0),.clk(gclk));
	jdff dff_A_aBwOw3bx5_0(.dout(w_dff_A_7h7Fu2Q37_0),.din(w_dff_A_aBwOw3bx5_0),.clk(gclk));
	jdff dff_A_L8UYUXoS7_0(.dout(w_dff_A_aBwOw3bx5_0),.din(w_dff_A_L8UYUXoS7_0),.clk(gclk));
	jdff dff_A_wOe423ER8_0(.dout(w_dff_A_L8UYUXoS7_0),.din(w_dff_A_wOe423ER8_0),.clk(gclk));
	jdff dff_A_VvECfKTc5_0(.dout(w_dff_A_wOe423ER8_0),.din(w_dff_A_VvECfKTc5_0),.clk(gclk));
	jdff dff_A_Ca2DWTUk9_0(.dout(w_dff_A_VvECfKTc5_0),.din(w_dff_A_Ca2DWTUk9_0),.clk(gclk));
	jdff dff_A_WYBF2niX3_0(.dout(w_dff_A_Ca2DWTUk9_0),.din(w_dff_A_WYBF2niX3_0),.clk(gclk));
	jdff dff_A_Eb5WXesu6_0(.dout(w_dff_A_WYBF2niX3_0),.din(w_dff_A_Eb5WXesu6_0),.clk(gclk));
	jdff dff_B_NkP5lfii7_1(.din(n154),.dout(w_dff_B_NkP5lfii7_1),.clk(gclk));
	jdff dff_B_rpyFMvjf6_0(.din(n165),.dout(w_dff_B_rpyFMvjf6_0),.clk(gclk));
	jdff dff_A_AV111u4x0_0(.dout(w_n164_0[0]),.din(w_dff_A_AV111u4x0_0),.clk(gclk));
	jdff dff_A_wo8KVVH63_0(.dout(w_dff_A_AV111u4x0_0),.din(w_dff_A_wo8KVVH63_0),.clk(gclk));
	jdff dff_A_ccHW2PQS0_0(.dout(w_dff_A_wo8KVVH63_0),.din(w_dff_A_ccHW2PQS0_0),.clk(gclk));
	jdff dff_A_Xhx1JmBs3_0(.dout(w_dff_A_ccHW2PQS0_0),.din(w_dff_A_Xhx1JmBs3_0),.clk(gclk));
	jdff dff_A_XsWQRDXO9_0(.dout(w_dff_A_Xhx1JmBs3_0),.din(w_dff_A_XsWQRDXO9_0),.clk(gclk));
	jdff dff_A_4GiB9DAe3_0(.dout(w_dff_A_XsWQRDXO9_0),.din(w_dff_A_4GiB9DAe3_0),.clk(gclk));
	jdff dff_B_ceKxluQL1_1(.din(n162),.dout(w_dff_B_ceKxluQL1_1),.clk(gclk));
	jdff dff_B_ixQvM5mF6_1(.din(w_dff_B_ceKxluQL1_1),.dout(w_dff_B_ixQvM5mF6_1),.clk(gclk));
	jdff dff_B_rwvNWt2F9_1(.din(w_dff_B_ixQvM5mF6_1),.dout(w_dff_B_rwvNWt2F9_1),.clk(gclk));
	jdff dff_B_DThuhYie8_1(.din(w_dff_B_rwvNWt2F9_1),.dout(w_dff_B_DThuhYie8_1),.clk(gclk));
	jdff dff_B_rOFVomLb6_1(.din(w_dff_B_DThuhYie8_1),.dout(w_dff_B_rOFVomLb6_1),.clk(gclk));
	jdff dff_B_KXeC1Orn6_1(.din(w_dff_B_rOFVomLb6_1),.dout(w_dff_B_KXeC1Orn6_1),.clk(gclk));
	jdff dff_A_k3fKdYD15_0(.dout(w_G112gat_0[0]),.din(w_dff_A_k3fKdYD15_0),.clk(gclk));
	jdff dff_A_whBlaFGt4_0(.dout(w_dff_A_k3fKdYD15_0),.din(w_dff_A_whBlaFGt4_0),.clk(gclk));
	jdff dff_A_CuHV83vG7_0(.dout(w_dff_A_whBlaFGt4_0),.din(w_dff_A_CuHV83vG7_0),.clk(gclk));
	jdff dff_A_HSg7n5MY5_0(.dout(w_dff_A_CuHV83vG7_0),.din(w_dff_A_HSg7n5MY5_0),.clk(gclk));
	jdff dff_A_cIuwW6t58_0(.dout(w_dff_A_HSg7n5MY5_0),.din(w_dff_A_cIuwW6t58_0),.clk(gclk));
	jdff dff_A_D1ma7eyi6_0(.dout(w_dff_A_cIuwW6t58_0),.din(w_dff_A_D1ma7eyi6_0),.clk(gclk));
	jdff dff_A_EdJiK31x6_0(.dout(w_dff_A_D1ma7eyi6_0),.din(w_dff_A_EdJiK31x6_0),.clk(gclk));
	jdff dff_A_r3BlC9AS4_0(.dout(w_dff_A_EdJiK31x6_0),.din(w_dff_A_r3BlC9AS4_0),.clk(gclk));
	jdff dff_A_Dsjj1ZWE9_0(.dout(w_dff_A_r3BlC9AS4_0),.din(w_dff_A_Dsjj1ZWE9_0),.clk(gclk));
	jdff dff_A_yUVK0bzL0_0(.dout(w_dff_A_Dsjj1ZWE9_0),.din(w_dff_A_yUVK0bzL0_0),.clk(gclk));
	jdff dff_A_bUhEWbP29_0(.dout(w_dff_A_yUVK0bzL0_0),.din(w_dff_A_bUhEWbP29_0),.clk(gclk));
	jdff dff_A_07xr8NJQ7_0(.dout(w_dff_A_bUhEWbP29_0),.din(w_dff_A_07xr8NJQ7_0),.clk(gclk));
	jdff dff_A_IGg9SyEP8_0(.dout(w_dff_A_07xr8NJQ7_0),.din(w_dff_A_IGg9SyEP8_0),.clk(gclk));
	jdff dff_A_A4cTJAJG0_1(.dout(w_G112gat_0[1]),.din(w_dff_A_A4cTJAJG0_1),.clk(gclk));
	jdff dff_A_VelxpJ7w3_1(.dout(w_dff_A_A4cTJAJG0_1),.din(w_dff_A_VelxpJ7w3_1),.clk(gclk));
	jdff dff_A_pbbzKgfQ3_1(.dout(w_dff_A_VelxpJ7w3_1),.din(w_dff_A_pbbzKgfQ3_1),.clk(gclk));
	jdff dff_A_CrRJtig80_1(.dout(w_dff_A_pbbzKgfQ3_1),.din(w_dff_A_CrRJtig80_1),.clk(gclk));
	jdff dff_A_16ISkeaI6_1(.dout(w_dff_A_CrRJtig80_1),.din(w_dff_A_16ISkeaI6_1),.clk(gclk));
	jdff dff_A_9HJ1m68B0_1(.dout(w_dff_A_16ISkeaI6_1),.din(w_dff_A_9HJ1m68B0_1),.clk(gclk));
	jdff dff_A_MRcXXCTX4_1(.dout(w_dff_A_9HJ1m68B0_1),.din(w_dff_A_MRcXXCTX4_1),.clk(gclk));
	jdff dff_A_Go6c1lDV5_1(.dout(w_dff_A_MRcXXCTX4_1),.din(w_dff_A_Go6c1lDV5_1),.clk(gclk));
	jdff dff_A_8zIyKzcm6_0(.dout(w_n159_0[0]),.din(w_dff_A_8zIyKzcm6_0),.clk(gclk));
	jdff dff_A_BXapyMDz5_0(.dout(w_dff_A_8zIyKzcm6_0),.din(w_dff_A_BXapyMDz5_0),.clk(gclk));
	jdff dff_A_FBcAiRaI0_0(.dout(w_dff_A_BXapyMDz5_0),.din(w_dff_A_FBcAiRaI0_0),.clk(gclk));
	jdff dff_A_jyNHHBvE5_0(.dout(w_dff_A_FBcAiRaI0_0),.din(w_dff_A_jyNHHBvE5_0),.clk(gclk));
	jdff dff_A_t01SNbxc5_0(.dout(w_dff_A_jyNHHBvE5_0),.din(w_dff_A_t01SNbxc5_0),.clk(gclk));
	jdff dff_A_LLFs3lMj2_0(.dout(w_dff_A_t01SNbxc5_0),.din(w_dff_A_LLFs3lMj2_0),.clk(gclk));
	jdff dff_A_O0hk1lCZ9_0(.dout(w_G34gat_0[0]),.din(w_dff_A_O0hk1lCZ9_0),.clk(gclk));
	jdff dff_A_iy7XwnFi0_0(.dout(w_dff_A_O0hk1lCZ9_0),.din(w_dff_A_iy7XwnFi0_0),.clk(gclk));
	jdff dff_A_9ClCkjFc1_0(.dout(w_dff_A_iy7XwnFi0_0),.din(w_dff_A_9ClCkjFc1_0),.clk(gclk));
	jdff dff_A_nDCd2ZVJ3_0(.dout(w_dff_A_9ClCkjFc1_0),.din(w_dff_A_nDCd2ZVJ3_0),.clk(gclk));
	jdff dff_A_PV5SEcjm8_0(.dout(w_dff_A_nDCd2ZVJ3_0),.din(w_dff_A_PV5SEcjm8_0),.clk(gclk));
	jdff dff_A_TfER06w00_0(.dout(w_dff_A_PV5SEcjm8_0),.din(w_dff_A_TfER06w00_0),.clk(gclk));
	jdff dff_A_azgze0TS8_0(.dout(w_dff_A_TfER06w00_0),.din(w_dff_A_azgze0TS8_0),.clk(gclk));
	jdff dff_A_4T1XvxtM9_0(.dout(w_dff_A_azgze0TS8_0),.din(w_dff_A_4T1XvxtM9_0),.clk(gclk));
	jdff dff_A_syqbI9W44_0(.dout(w_dff_A_4T1XvxtM9_0),.din(w_dff_A_syqbI9W44_0),.clk(gclk));
	jdff dff_A_NlPQNhwO8_0(.dout(w_dff_A_syqbI9W44_0),.din(w_dff_A_NlPQNhwO8_0),.clk(gclk));
	jdff dff_A_Cd7ZuZQ00_0(.dout(w_dff_A_NlPQNhwO8_0),.din(w_dff_A_Cd7ZuZQ00_0),.clk(gclk));
	jdff dff_A_ZMqb7ndf1_0(.dout(w_dff_A_Cd7ZuZQ00_0),.din(w_dff_A_ZMqb7ndf1_0),.clk(gclk));
	jdff dff_A_qZdLlFXE3_0(.dout(w_dff_A_ZMqb7ndf1_0),.din(w_dff_A_qZdLlFXE3_0),.clk(gclk));
	jdff dff_A_6QRAG9CT9_1(.dout(w_G34gat_0[1]),.din(w_dff_A_6QRAG9CT9_1),.clk(gclk));
	jdff dff_A_AcLiwcxi2_1(.dout(w_dff_A_6QRAG9CT9_1),.din(w_dff_A_AcLiwcxi2_1),.clk(gclk));
	jdff dff_A_qcwqUm645_1(.dout(w_dff_A_AcLiwcxi2_1),.din(w_dff_A_qcwqUm645_1),.clk(gclk));
	jdff dff_A_dYv6qkAD3_1(.dout(w_dff_A_qcwqUm645_1),.din(w_dff_A_dYv6qkAD3_1),.clk(gclk));
	jdff dff_A_dVLWKPsM2_1(.dout(w_dff_A_dYv6qkAD3_1),.din(w_dff_A_dVLWKPsM2_1),.clk(gclk));
	jdff dff_A_aGjZh8xo6_1(.dout(w_dff_A_dVLWKPsM2_1),.din(w_dff_A_aGjZh8xo6_1),.clk(gclk));
	jdff dff_A_uxhi2cct6_1(.dout(w_dff_A_aGjZh8xo6_1),.din(w_dff_A_uxhi2cct6_1),.clk(gclk));
	jdff dff_A_z7fBMfWI3_1(.dout(w_dff_A_uxhi2cct6_1),.din(w_dff_A_z7fBMfWI3_1),.clk(gclk));
	jdff dff_A_2oNqJcOO7_0(.dout(w_n156_0[0]),.din(w_dff_A_2oNqJcOO7_0),.clk(gclk));
	jdff dff_A_HRjeNp6v5_0(.dout(w_dff_A_2oNqJcOO7_0),.din(w_dff_A_HRjeNp6v5_0),.clk(gclk));
	jdff dff_A_aQ800rtG2_0(.dout(w_dff_A_HRjeNp6v5_0),.din(w_dff_A_aQ800rtG2_0),.clk(gclk));
	jdff dff_A_2zq3WU0W6_0(.dout(w_dff_A_aQ800rtG2_0),.din(w_dff_A_2zq3WU0W6_0),.clk(gclk));
	jdff dff_A_uV1tepnh5_0(.dout(w_dff_A_2zq3WU0W6_0),.din(w_dff_A_uV1tepnh5_0),.clk(gclk));
	jdff dff_A_sKncualL7_0(.dout(w_dff_A_uV1tepnh5_0),.din(w_dff_A_sKncualL7_0),.clk(gclk));
	jdff dff_A_5RRJF1ak2_1(.dout(w_n138_0[1]),.din(w_dff_A_5RRJF1ak2_1),.clk(gclk));
	jdff dff_A_L1yUcqb50_1(.dout(w_dff_A_5RRJF1ak2_1),.din(w_dff_A_L1yUcqb50_1),.clk(gclk));
	jdff dff_A_dkLUS4L14_1(.dout(w_dff_A_L1yUcqb50_1),.din(w_dff_A_dkLUS4L14_1),.clk(gclk));
	jdff dff_A_2m4pnNzZ3_1(.dout(w_dff_A_dkLUS4L14_1),.din(w_dff_A_2m4pnNzZ3_1),.clk(gclk));
	jdff dff_A_euCG29MY4_1(.dout(w_dff_A_2m4pnNzZ3_1),.din(w_dff_A_euCG29MY4_1),.clk(gclk));
	jdff dff_A_GzJpBzPy9_1(.dout(w_dff_A_euCG29MY4_1),.din(w_dff_A_GzJpBzPy9_1),.clk(gclk));
	jdff dff_A_TQUWBhtX2_0(.dout(w_G99gat_0[0]),.din(w_dff_A_TQUWBhtX2_0),.clk(gclk));
	jdff dff_A_vJIq0LWk4_0(.dout(w_dff_A_TQUWBhtX2_0),.din(w_dff_A_vJIq0LWk4_0),.clk(gclk));
	jdff dff_A_NYzJIYwp2_0(.dout(w_dff_A_vJIq0LWk4_0),.din(w_dff_A_NYzJIYwp2_0),.clk(gclk));
	jdff dff_A_duF1Fab66_0(.dout(w_dff_A_NYzJIYwp2_0),.din(w_dff_A_duF1Fab66_0),.clk(gclk));
	jdff dff_A_HqieGEOn9_0(.dout(w_dff_A_duF1Fab66_0),.din(w_dff_A_HqieGEOn9_0),.clk(gclk));
	jdff dff_A_STDLK6Qv8_0(.dout(w_dff_A_HqieGEOn9_0),.din(w_dff_A_STDLK6Qv8_0),.clk(gclk));
	jdff dff_A_nZgFW8Dk0_0(.dout(w_dff_A_STDLK6Qv8_0),.din(w_dff_A_nZgFW8Dk0_0),.clk(gclk));
	jdff dff_A_EV2WFCl09_0(.dout(w_dff_A_nZgFW8Dk0_0),.din(w_dff_A_EV2WFCl09_0),.clk(gclk));
	jdff dff_A_MvLqRxip3_1(.dout(w_G99gat_0[1]),.din(w_dff_A_MvLqRxip3_1),.clk(gclk));
	jdff dff_A_wLWdPZcw9_1(.dout(w_dff_A_MvLqRxip3_1),.din(w_dff_A_wLWdPZcw9_1),.clk(gclk));
	jdff dff_A_bLQHGVVf3_1(.dout(w_dff_A_wLWdPZcw9_1),.din(w_dff_A_bLQHGVVf3_1),.clk(gclk));
	jdff dff_A_VFNv39zM4_1(.dout(w_dff_A_bLQHGVVf3_1),.din(w_dff_A_VFNv39zM4_1),.clk(gclk));
	jdff dff_A_bvzu4eKc1_1(.dout(w_dff_A_VFNv39zM4_1),.din(w_dff_A_bvzu4eKc1_1),.clk(gclk));
	jdff dff_A_O7QdYVcU6_1(.dout(w_dff_A_bvzu4eKc1_1),.din(w_dff_A_O7QdYVcU6_1),.clk(gclk));
	jdff dff_A_NazXc7KQ6_1(.dout(w_dff_A_O7QdYVcU6_1),.din(w_dff_A_NazXc7KQ6_1),.clk(gclk));
	jdff dff_A_7yy3x1e71_1(.dout(w_dff_A_NazXc7KQ6_1),.din(w_dff_A_7yy3x1e71_1),.clk(gclk));
	jdff dff_A_xPBJ9FAM0_1(.dout(w_dff_A_7yy3x1e71_1),.din(w_dff_A_xPBJ9FAM0_1),.clk(gclk));
	jdff dff_A_fQLewJoZ8_1(.dout(w_dff_A_xPBJ9FAM0_1),.din(w_dff_A_fQLewJoZ8_1),.clk(gclk));
	jdff dff_A_9vng2tpv8_1(.dout(w_dff_A_fQLewJoZ8_1),.din(w_dff_A_9vng2tpv8_1),.clk(gclk));
	jdff dff_A_chPBt41z6_1(.dout(w_dff_A_9vng2tpv8_1),.din(w_dff_A_chPBt41z6_1),.clk(gclk));
	jdff dff_A_xwKVzm7V8_1(.dout(w_dff_A_chPBt41z6_1),.din(w_dff_A_xwKVzm7V8_1),.clk(gclk));
	jdff dff_A_BRBQYKct3_0(.dout(w_n151_0[0]),.din(w_dff_A_BRBQYKct3_0),.clk(gclk));
	jdff dff_A_7nwawlw80_0(.dout(w_dff_A_BRBQYKct3_0),.din(w_dff_A_7nwawlw80_0),.clk(gclk));
	jdff dff_A_IOns0ZG35_0(.dout(w_dff_A_7nwawlw80_0),.din(w_dff_A_IOns0ZG35_0),.clk(gclk));
	jdff dff_A_0UIFhdOv2_0(.dout(w_dff_A_IOns0ZG35_0),.din(w_dff_A_0UIFhdOv2_0),.clk(gclk));
	jdff dff_A_DZmf4tuv4_0(.dout(w_dff_A_0UIFhdOv2_0),.din(w_dff_A_DZmf4tuv4_0),.clk(gclk));
	jdff dff_A_YjxOWqGe8_0(.dout(w_dff_A_DZmf4tuv4_0),.din(w_dff_A_YjxOWqGe8_0),.clk(gclk));
	jdff dff_B_YwTz4Rdk3_1(.din(n48),.dout(w_dff_B_YwTz4Rdk3_1),.clk(gclk));
	jdff dff_B_13jNcIH78_1(.din(n61),.dout(w_dff_B_13jNcIH78_1),.clk(gclk));
	jdff dff_A_JInPuuqa8_0(.dout(w_n64_0[0]),.din(w_dff_A_JInPuuqa8_0),.clk(gclk));
	jdff dff_A_G1Aw1gSS7_0(.dout(w_dff_A_JInPuuqa8_0),.din(w_dff_A_G1Aw1gSS7_0),.clk(gclk));
	jdff dff_A_aNspGlsp1_0(.dout(w_dff_A_G1Aw1gSS7_0),.din(w_dff_A_aNspGlsp1_0),.clk(gclk));
	jdff dff_A_GDQYNaQN9_0(.dout(w_dff_A_aNspGlsp1_0),.din(w_dff_A_GDQYNaQN9_0),.clk(gclk));
	jdff dff_A_kSn583jH5_0(.dout(w_dff_A_GDQYNaQN9_0),.din(w_dff_A_kSn583jH5_0),.clk(gclk));
	jdff dff_A_TBubJOYM9_0(.dout(w_n62_0[0]),.din(w_dff_A_TBubJOYM9_0),.clk(gclk));
	jdff dff_A_8WMfvOJY9_0(.dout(w_dff_A_TBubJOYM9_0),.din(w_dff_A_8WMfvOJY9_0),.clk(gclk));
	jdff dff_A_B6ddvVpF3_0(.dout(w_dff_A_8WMfvOJY9_0),.din(w_dff_A_B6ddvVpF3_0),.clk(gclk));
	jdff dff_A_IaUakkkr1_0(.dout(w_dff_A_B6ddvVpF3_0),.din(w_dff_A_IaUakkkr1_0),.clk(gclk));
	jdff dff_A_fk6MrzLy9_0(.dout(w_dff_A_IaUakkkr1_0),.din(w_dff_A_fk6MrzLy9_0),.clk(gclk));
	jdff dff_A_UMoQmOdK2_0(.dout(w_n60_0[0]),.din(w_dff_A_UMoQmOdK2_0),.clk(gclk));
	jdff dff_A_qqnjVmhM7_0(.dout(w_dff_A_UMoQmOdK2_0),.din(w_dff_A_qqnjVmhM7_0),.clk(gclk));
	jdff dff_A_hrgFTxrx9_0(.dout(w_dff_A_qqnjVmhM7_0),.din(w_dff_A_hrgFTxrx9_0),.clk(gclk));
	jdff dff_A_7AlZQU0f4_0(.dout(w_dff_A_hrgFTxrx9_0),.din(w_dff_A_7AlZQU0f4_0),.clk(gclk));
	jdff dff_A_9mFFV7fQ3_0(.dout(w_dff_A_7AlZQU0f4_0),.din(w_dff_A_9mFFV7fQ3_0),.clk(gclk));
	jdff dff_A_XFRjWb0e7_0(.dout(w_n57_0[0]),.din(w_dff_A_XFRjWb0e7_0),.clk(gclk));
	jdff dff_A_AB5AJAx93_0(.dout(w_dff_A_XFRjWb0e7_0),.din(w_dff_A_AB5AJAx93_0),.clk(gclk));
	jdff dff_A_7sx2afBE9_0(.dout(w_dff_A_AB5AJAx93_0),.din(w_dff_A_7sx2afBE9_0),.clk(gclk));
	jdff dff_A_rlN0UfkF4_0(.dout(w_dff_A_7sx2afBE9_0),.din(w_dff_A_rlN0UfkF4_0),.clk(gclk));
	jdff dff_A_ZeyIuTAQ0_0(.dout(w_n54_0[0]),.din(w_dff_A_ZeyIuTAQ0_0),.clk(gclk));
	jdff dff_A_XfAAkZ0G4_0(.dout(w_dff_A_ZeyIuTAQ0_0),.din(w_dff_A_XfAAkZ0G4_0),.clk(gclk));
	jdff dff_A_s1kCKJxT9_0(.dout(w_dff_A_XfAAkZ0G4_0),.din(w_dff_A_s1kCKJxT9_0),.clk(gclk));
	jdff dff_A_JwZoJf724_0(.dout(w_dff_A_s1kCKJxT9_0),.din(w_dff_A_JwZoJf724_0),.clk(gclk));
	jdff dff_A_2sB8qnBj9_0(.dout(w_dff_A_JwZoJf724_0),.din(w_dff_A_2sB8qnBj9_0),.clk(gclk));
	jdff dff_A_dmo9lwF68_0(.dout(w_n51_0[0]),.din(w_dff_A_dmo9lwF68_0),.clk(gclk));
	jdff dff_A_cN0njtaj5_0(.dout(w_dff_A_dmo9lwF68_0),.din(w_dff_A_cN0njtaj5_0),.clk(gclk));
	jdff dff_A_uwlUsmnk9_0(.dout(w_dff_A_cN0njtaj5_0),.din(w_dff_A_uwlUsmnk9_0),.clk(gclk));
	jdff dff_A_CNqPklHs0_0(.dout(w_dff_A_uwlUsmnk9_0),.din(w_dff_A_CNqPklHs0_0),.clk(gclk));
	jdff dff_A_EODEH6fW7_0(.dout(w_dff_A_CNqPklHs0_0),.din(w_dff_A_EODEH6fW7_0),.clk(gclk));
	jdff dff_A_GjiScDiW3_0(.dout(w_n47_0[0]),.din(w_dff_A_GjiScDiW3_0),.clk(gclk));
	jdff dff_A_R73CpPBc0_0(.dout(w_dff_A_GjiScDiW3_0),.din(w_dff_A_R73CpPBc0_0),.clk(gclk));
	jdff dff_A_nhp2kmJQ0_0(.dout(w_dff_A_R73CpPBc0_0),.din(w_dff_A_nhp2kmJQ0_0),.clk(gclk));
	jdff dff_A_X3q7bKiM4_0(.dout(w_G21gat_0[0]),.din(w_dff_A_X3q7bKiM4_0),.clk(gclk));
	jdff dff_A_RNTOFx799_0(.dout(w_dff_A_X3q7bKiM4_0),.din(w_dff_A_RNTOFx799_0),.clk(gclk));
	jdff dff_A_SN7SJ5w29_0(.dout(w_dff_A_RNTOFx799_0),.din(w_dff_A_SN7SJ5w29_0),.clk(gclk));
	jdff dff_A_Y8ekKrsm4_0(.dout(w_dff_A_SN7SJ5w29_0),.din(w_dff_A_Y8ekKrsm4_0),.clk(gclk));
	jdff dff_A_IqGY3AHw1_0(.dout(w_dff_A_Y8ekKrsm4_0),.din(w_dff_A_IqGY3AHw1_0),.clk(gclk));
	jdff dff_A_bSHxnqms8_0(.dout(w_dff_A_IqGY3AHw1_0),.din(w_dff_A_bSHxnqms8_0),.clk(gclk));
	jdff dff_A_anc3jKno6_0(.dout(w_dff_A_bSHxnqms8_0),.din(w_dff_A_anc3jKno6_0),.clk(gclk));
	jdff dff_A_AOrQJtKy9_0(.dout(w_dff_A_anc3jKno6_0),.din(w_dff_A_AOrQJtKy9_0),.clk(gclk));
	jdff dff_A_YHIgEvW72_0(.dout(w_dff_A_AOrQJtKy9_0),.din(w_dff_A_YHIgEvW72_0),.clk(gclk));
	jdff dff_A_M8ITuz5Y3_0(.dout(w_dff_A_YHIgEvW72_0),.din(w_dff_A_M8ITuz5Y3_0),.clk(gclk));
	jdff dff_A_hXIi3Tfy1_0(.dout(w_dff_A_M8ITuz5Y3_0),.din(w_dff_A_hXIi3Tfy1_0),.clk(gclk));
	jdff dff_A_ReeXbjtY2_0(.dout(w_dff_A_hXIi3Tfy1_0),.din(w_dff_A_ReeXbjtY2_0),.clk(gclk));
	jdff dff_A_9ygUFtzK9_0(.dout(w_dff_A_ReeXbjtY2_0),.din(w_dff_A_9ygUFtzK9_0),.clk(gclk));
	jdff dff_A_cGZvoynY1_1(.dout(w_G21gat_0[1]),.din(w_dff_A_cGZvoynY1_1),.clk(gclk));
	jdff dff_A_TPD2k8Xz9_1(.dout(w_dff_A_cGZvoynY1_1),.din(w_dff_A_TPD2k8Xz9_1),.clk(gclk));
	jdff dff_A_TqNdzYTj2_1(.dout(w_dff_A_TPD2k8Xz9_1),.din(w_dff_A_TqNdzYTj2_1),.clk(gclk));
	jdff dff_A_ETYGaLcs1_1(.dout(w_dff_A_TqNdzYTj2_1),.din(w_dff_A_ETYGaLcs1_1),.clk(gclk));
	jdff dff_A_kkX8SL0T2_1(.dout(w_dff_A_ETYGaLcs1_1),.din(w_dff_A_kkX8SL0T2_1),.clk(gclk));
	jdff dff_A_1J93v6sV9_1(.dout(w_dff_A_kkX8SL0T2_1),.din(w_dff_A_1J93v6sV9_1),.clk(gclk));
	jdff dff_A_uMKEEnY32_1(.dout(w_dff_A_1J93v6sV9_1),.din(w_dff_A_uMKEEnY32_1),.clk(gclk));
	jdff dff_A_2UsyUsik1_1(.dout(w_dff_A_uMKEEnY32_1),.din(w_dff_A_2UsyUsik1_1),.clk(gclk));
	jdff dff_A_XHwaf2sQ1_0(.dout(w_n102_0[0]),.din(w_dff_A_XHwaf2sQ1_0),.clk(gclk));
	jdff dff_A_9NlhitPg0_0(.dout(w_dff_A_XHwaf2sQ1_0),.din(w_dff_A_9NlhitPg0_0),.clk(gclk));
	jdff dff_A_omjH5Oei0_0(.dout(w_dff_A_9NlhitPg0_0),.din(w_dff_A_omjH5Oei0_0),.clk(gclk));
	jdff dff_A_nhH959ff2_0(.dout(w_dff_A_omjH5Oei0_0),.din(w_dff_A_nhH959ff2_0),.clk(gclk));
	jdff dff_A_xQEWaPFd4_0(.dout(w_dff_A_nhH959ff2_0),.din(w_dff_A_xQEWaPFd4_0),.clk(gclk));
	jdff dff_B_ixIUlemi6_2(.din(n102),.dout(w_dff_B_ixIUlemi6_2),.clk(gclk));
	jdff dff_B_oN58kuea0_2(.din(w_dff_B_ixIUlemi6_2),.dout(w_dff_B_oN58kuea0_2),.clk(gclk));
	jdff dff_B_Q9b2boXO0_2(.din(w_dff_B_oN58kuea0_2),.dout(w_dff_B_Q9b2boXO0_2),.clk(gclk));
	jdff dff_B_vHmKgquF2_2(.din(w_dff_B_Q9b2boXO0_2),.dout(w_dff_B_vHmKgquF2_2),.clk(gclk));
	jdff dff_B_t6OXCiwM1_2(.din(w_dff_B_vHmKgquF2_2),.dout(w_dff_B_t6OXCiwM1_2),.clk(gclk));
	jdff dff_B_yn1gTL1Z5_2(.din(w_dff_B_t6OXCiwM1_2),.dout(w_dff_B_yn1gTL1Z5_2),.clk(gclk));
	jdff dff_B_IF04gzgP6_2(.din(w_dff_B_yn1gTL1Z5_2),.dout(w_dff_B_IF04gzgP6_2),.clk(gclk));
	jdff dff_A_bU10WHIn3_0(.dout(w_G73gat_0[0]),.din(w_dff_A_bU10WHIn3_0),.clk(gclk));
	jdff dff_A_hvrbYllE2_0(.dout(w_dff_A_bU10WHIn3_0),.din(w_dff_A_hvrbYllE2_0),.clk(gclk));
	jdff dff_A_TxrgJKPe2_0(.dout(w_dff_A_hvrbYllE2_0),.din(w_dff_A_TxrgJKPe2_0),.clk(gclk));
	jdff dff_A_3UCTd4K72_0(.dout(w_dff_A_TxrgJKPe2_0),.din(w_dff_A_3UCTd4K72_0),.clk(gclk));
	jdff dff_A_QMSVHAYt5_0(.dout(w_dff_A_3UCTd4K72_0),.din(w_dff_A_QMSVHAYt5_0),.clk(gclk));
	jdff dff_A_hyeI8XLQ6_0(.dout(w_dff_A_QMSVHAYt5_0),.din(w_dff_A_hyeI8XLQ6_0),.clk(gclk));
	jdff dff_A_Cz0JYlKT3_0(.dout(w_dff_A_hyeI8XLQ6_0),.din(w_dff_A_Cz0JYlKT3_0),.clk(gclk));
	jdff dff_A_h8TvgjHo5_0(.dout(w_dff_A_Cz0JYlKT3_0),.din(w_dff_A_h8TvgjHo5_0),.clk(gclk));
	jdff dff_A_GwkEOQSb7_0(.dout(w_dff_A_h8TvgjHo5_0),.din(w_dff_A_GwkEOQSb7_0),.clk(gclk));
	jdff dff_A_HivPc0ry6_0(.dout(w_dff_A_GwkEOQSb7_0),.din(w_dff_A_HivPc0ry6_0),.clk(gclk));
	jdff dff_A_NSJpxvh96_0(.dout(w_dff_A_HivPc0ry6_0),.din(w_dff_A_NSJpxvh96_0),.clk(gclk));
	jdff dff_A_PjSU1GIe5_0(.dout(w_dff_A_NSJpxvh96_0),.din(w_dff_A_PjSU1GIe5_0),.clk(gclk));
	jdff dff_A_YZreO8RO2_0(.dout(w_dff_A_PjSU1GIe5_0),.din(w_dff_A_YZreO8RO2_0),.clk(gclk));
	jdff dff_A_HUmFkQhw3_1(.dout(w_G73gat_0[1]),.din(w_dff_A_HUmFkQhw3_1),.clk(gclk));
	jdff dff_A_EKVT5ugf1_1(.dout(w_dff_A_HUmFkQhw3_1),.din(w_dff_A_EKVT5ugf1_1),.clk(gclk));
	jdff dff_A_AZ5gkIHl5_1(.dout(w_dff_A_EKVT5ugf1_1),.din(w_dff_A_AZ5gkIHl5_1),.clk(gclk));
	jdff dff_A_mj4enfqA6_1(.dout(w_dff_A_AZ5gkIHl5_1),.din(w_dff_A_mj4enfqA6_1),.clk(gclk));
	jdff dff_A_b3uE29Xi6_1(.dout(w_dff_A_mj4enfqA6_1),.din(w_dff_A_b3uE29Xi6_1),.clk(gclk));
	jdff dff_A_SfkfkjLP5_1(.dout(w_dff_A_b3uE29Xi6_1),.din(w_dff_A_SfkfkjLP5_1),.clk(gclk));
	jdff dff_A_ilKvU5Xf7_1(.dout(w_dff_A_SfkfkjLP5_1),.din(w_dff_A_ilKvU5Xf7_1),.clk(gclk));
	jdff dff_A_EE1vAm416_1(.dout(w_dff_A_ilKvU5Xf7_1),.din(w_dff_A_EE1vAm416_1),.clk(gclk));
	jdff dff_A_U9Sinh8X8_0(.dout(w_n104_0[0]),.din(w_dff_A_U9Sinh8X8_0),.clk(gclk));
	jdff dff_A_1CKWLqAN1_0(.dout(w_dff_A_U9Sinh8X8_0),.din(w_dff_A_1CKWLqAN1_0),.clk(gclk));
	jdff dff_A_1jdCjZXD7_0(.dout(w_dff_A_1CKWLqAN1_0),.din(w_dff_A_1jdCjZXD7_0),.clk(gclk));
	jdff dff_A_ScTkoQ8O2_0(.dout(w_dff_A_1jdCjZXD7_0),.din(w_dff_A_ScTkoQ8O2_0),.clk(gclk));
	jdff dff_A_4sJ3XD5G4_0(.dout(w_dff_A_ScTkoQ8O2_0),.din(w_dff_A_4sJ3XD5G4_0),.clk(gclk));
	jdff dff_A_zUsGRMpU8_0(.dout(w_dff_A_4sJ3XD5G4_0),.din(w_dff_A_zUsGRMpU8_0),.clk(gclk));
	jdff dff_B_iVWKt9F30_1(.din(n72),.dout(w_dff_B_iVWKt9F30_1),.clk(gclk));
	jdff dff_B_7OeTX8tP1_1(.din(n85),.dout(w_dff_B_7OeTX8tP1_1),.clk(gclk));
	jdff dff_A_cLYJzDLR9_0(.dout(w_n88_0[0]),.din(w_dff_A_cLYJzDLR9_0),.clk(gclk));
	jdff dff_A_9d8Zy8bX8_0(.dout(w_dff_A_cLYJzDLR9_0),.din(w_dff_A_9d8Zy8bX8_0),.clk(gclk));
	jdff dff_A_I8zY70O09_0(.dout(w_dff_A_9d8Zy8bX8_0),.din(w_dff_A_I8zY70O09_0),.clk(gclk));
	jdff dff_A_nKaof8P33_0(.dout(w_dff_A_I8zY70O09_0),.din(w_dff_A_nKaof8P33_0),.clk(gclk));
	jdff dff_A_AsYHRkx51_0(.dout(w_dff_A_nKaof8P33_0),.din(w_dff_A_AsYHRkx51_0),.clk(gclk));
	jdff dff_A_kwJpDK9d3_0(.dout(w_dff_A_AsYHRkx51_0),.din(w_dff_A_kwJpDK9d3_0),.clk(gclk));
	jdff dff_A_pJCoHLR02_0(.dout(w_G82gat_0[0]),.din(w_dff_A_pJCoHLR02_0),.clk(gclk));
	jdff dff_A_SeAMmSL87_0(.dout(w_dff_A_pJCoHLR02_0),.din(w_dff_A_SeAMmSL87_0),.clk(gclk));
	jdff dff_A_qakHzVMB1_0(.dout(w_dff_A_SeAMmSL87_0),.din(w_dff_A_qakHzVMB1_0),.clk(gclk));
	jdff dff_A_NZCBwXPu8_0(.dout(w_dff_A_qakHzVMB1_0),.din(w_dff_A_NZCBwXPu8_0),.clk(gclk));
	jdff dff_A_8Ff8nEbI3_0(.dout(w_dff_A_NZCBwXPu8_0),.din(w_dff_A_8Ff8nEbI3_0),.clk(gclk));
	jdff dff_A_6gIMxOOk2_0(.dout(w_dff_A_8Ff8nEbI3_0),.din(w_dff_A_6gIMxOOk2_0),.clk(gclk));
	jdff dff_A_NE6oXFhM3_0(.dout(w_dff_A_6gIMxOOk2_0),.din(w_dff_A_NE6oXFhM3_0),.clk(gclk));
	jdff dff_A_jCLSgv0p3_2(.dout(w_G82gat_0[2]),.din(w_dff_A_jCLSgv0p3_2),.clk(gclk));
	jdff dff_A_pRmSFdzO9_0(.dout(w_G76gat_0[0]),.din(w_dff_A_pRmSFdzO9_0),.clk(gclk));
	jdff dff_A_tW2aJNWD6_0(.dout(w_dff_A_pRmSFdzO9_0),.din(w_dff_A_tW2aJNWD6_0),.clk(gclk));
	jdff dff_A_eTIT3P1E9_0(.dout(w_dff_A_tW2aJNWD6_0),.din(w_dff_A_eTIT3P1E9_0),.clk(gclk));
	jdff dff_A_lbMIEfNe9_0(.dout(w_dff_A_eTIT3P1E9_0),.din(w_dff_A_lbMIEfNe9_0),.clk(gclk));
	jdff dff_A_iOnzaU6I2_0(.dout(w_dff_A_lbMIEfNe9_0),.din(w_dff_A_iOnzaU6I2_0),.clk(gclk));
	jdff dff_A_9dUrKNKd3_0(.dout(w_dff_A_iOnzaU6I2_0),.din(w_dff_A_9dUrKNKd3_0),.clk(gclk));
	jdff dff_A_0ivgQ7UW7_1(.dout(w_G76gat_0[1]),.din(w_dff_A_0ivgQ7UW7_1),.clk(gclk));
	jdff dff_A_sQG3aNIQ2_0(.dout(w_n86_0[0]),.din(w_dff_A_sQG3aNIQ2_0),.clk(gclk));
	jdff dff_A_NSLkkRcy3_0(.dout(w_dff_A_sQG3aNIQ2_0),.din(w_dff_A_NSLkkRcy3_0),.clk(gclk));
	jdff dff_A_NZvhiyj07_0(.dout(w_dff_A_NSLkkRcy3_0),.din(w_dff_A_NZvhiyj07_0),.clk(gclk));
	jdff dff_A_TtnypJFA6_0(.dout(w_dff_A_NZvhiyj07_0),.din(w_dff_A_TtnypJFA6_0),.clk(gclk));
	jdff dff_A_JuVeqah71_0(.dout(w_dff_A_TtnypJFA6_0),.din(w_dff_A_JuVeqah71_0),.clk(gclk));
	jdff dff_A_VfX4Xf9w3_0(.dout(w_dff_A_JuVeqah71_0),.din(w_dff_A_VfX4Xf9w3_0),.clk(gclk));
	jdff dff_A_9RG3yveU9_0(.dout(w_G95gat_0[0]),.din(w_dff_A_9RG3yveU9_0),.clk(gclk));
	jdff dff_A_27ER9Jzv1_0(.dout(w_dff_A_9RG3yveU9_0),.din(w_dff_A_27ER9Jzv1_0),.clk(gclk));
	jdff dff_A_tSk2aKxK9_0(.dout(w_dff_A_27ER9Jzv1_0),.din(w_dff_A_tSk2aKxK9_0),.clk(gclk));
	jdff dff_A_R0n8zemA2_0(.dout(w_dff_A_tSk2aKxK9_0),.din(w_dff_A_R0n8zemA2_0),.clk(gclk));
	jdff dff_A_wyeJougk1_0(.dout(w_dff_A_R0n8zemA2_0),.din(w_dff_A_wyeJougk1_0),.clk(gclk));
	jdff dff_A_rq5gl4iL9_0(.dout(w_dff_A_wyeJougk1_0),.din(w_dff_A_rq5gl4iL9_0),.clk(gclk));
	jdff dff_A_1s5F0kqf1_0(.dout(w_dff_A_rq5gl4iL9_0),.din(w_dff_A_1s5F0kqf1_0),.clk(gclk));
	jdff dff_A_m3tq5pOZ7_2(.dout(w_G95gat_0[2]),.din(w_dff_A_m3tq5pOZ7_2),.clk(gclk));
	jdff dff_A_bc99Wd5Z3_0(.dout(w_G89gat_0[0]),.din(w_dff_A_bc99Wd5Z3_0),.clk(gclk));
	jdff dff_A_vtgvAEaQ7_0(.dout(w_dff_A_bc99Wd5Z3_0),.din(w_dff_A_vtgvAEaQ7_0),.clk(gclk));
	jdff dff_A_jei1LsGN8_0(.dout(w_dff_A_vtgvAEaQ7_0),.din(w_dff_A_jei1LsGN8_0),.clk(gclk));
	jdff dff_A_sOO6HaqA6_0(.dout(w_dff_A_jei1LsGN8_0),.din(w_dff_A_sOO6HaqA6_0),.clk(gclk));
	jdff dff_A_d2JnQgsp2_0(.dout(w_dff_A_sOO6HaqA6_0),.din(w_dff_A_d2JnQgsp2_0),.clk(gclk));
	jdff dff_A_lKn6yJlJ6_0(.dout(w_dff_A_d2JnQgsp2_0),.din(w_dff_A_lKn6yJlJ6_0),.clk(gclk));
	jdff dff_A_TRRJesDS2_1(.dout(w_G89gat_0[1]),.din(w_dff_A_TRRJesDS2_1),.clk(gclk));
	jdff dff_A_xVmFd9Dm5_0(.dout(w_n84_0[0]),.din(w_dff_A_xVmFd9Dm5_0),.clk(gclk));
	jdff dff_A_uMGYBVYl1_0(.dout(w_dff_A_xVmFd9Dm5_0),.din(w_dff_A_uMGYBVYl1_0),.clk(gclk));
	jdff dff_A_EiSnpKIJ6_0(.dout(w_dff_A_uMGYBVYl1_0),.din(w_dff_A_EiSnpKIJ6_0),.clk(gclk));
	jdff dff_A_T7qDgt7E6_0(.dout(w_dff_A_EiSnpKIJ6_0),.din(w_dff_A_T7qDgt7E6_0),.clk(gclk));
	jdff dff_A_dOTcBzwc9_0(.dout(w_dff_A_T7qDgt7E6_0),.din(w_dff_A_dOTcBzwc9_0),.clk(gclk));
	jdff dff_A_gGNBgYqU5_0(.dout(w_dff_A_dOTcBzwc9_0),.din(w_dff_A_gGNBgYqU5_0),.clk(gclk));
	jdff dff_A_pcgnEsJ98_0(.dout(w_G4gat_0[0]),.din(w_dff_A_pcgnEsJ98_0),.clk(gclk));
	jdff dff_A_GmnGWvfI8_0(.dout(w_dff_A_pcgnEsJ98_0),.din(w_dff_A_GmnGWvfI8_0),.clk(gclk));
	jdff dff_A_VHqVsIXk3_0(.dout(w_dff_A_GmnGWvfI8_0),.din(w_dff_A_VHqVsIXk3_0),.clk(gclk));
	jdff dff_A_2D6P5aMx2_0(.dout(w_dff_A_VHqVsIXk3_0),.din(w_dff_A_2D6P5aMx2_0),.clk(gclk));
	jdff dff_A_WiWzKvF72_0(.dout(w_dff_A_2D6P5aMx2_0),.din(w_dff_A_WiWzKvF72_0),.clk(gclk));
	jdff dff_A_S1nC82Tx3_0(.dout(w_dff_A_WiWzKvF72_0),.din(w_dff_A_S1nC82Tx3_0),.clk(gclk));
	jdff dff_A_u2Wkcub51_0(.dout(w_dff_A_S1nC82Tx3_0),.din(w_dff_A_u2Wkcub51_0),.clk(gclk));
	jdff dff_A_CPVaA3YE2_2(.dout(w_G4gat_0[2]),.din(w_dff_A_CPVaA3YE2_2),.clk(gclk));
	jdff dff_A_hl3QBdk34_0(.dout(w_G1gat_0[0]),.din(w_dff_A_hl3QBdk34_0),.clk(gclk));
	jdff dff_A_M4NHu0WP6_0(.dout(w_dff_A_hl3QBdk34_0),.din(w_dff_A_M4NHu0WP6_0),.clk(gclk));
	jdff dff_A_2GBha37m9_0(.dout(w_dff_A_M4NHu0WP6_0),.din(w_dff_A_2GBha37m9_0),.clk(gclk));
	jdff dff_A_dTgi6XPn2_0(.dout(w_dff_A_2GBha37m9_0),.din(w_dff_A_dTgi6XPn2_0),.clk(gclk));
	jdff dff_A_7fGXVDn78_0(.dout(w_dff_A_dTgi6XPn2_0),.din(w_dff_A_7fGXVDn78_0),.clk(gclk));
	jdff dff_A_9feHHqEP9_0(.dout(w_dff_A_7fGXVDn78_0),.din(w_dff_A_9feHHqEP9_0),.clk(gclk));
	jdff dff_A_ZUmlp4ih2_1(.dout(w_G1gat_0[1]),.din(w_dff_A_ZUmlp4ih2_1),.clk(gclk));
	jdff dff_A_893RPwEf4_0(.dout(w_n81_0[0]),.din(w_dff_A_893RPwEf4_0),.clk(gclk));
	jdff dff_A_luoqwI3p0_0(.dout(w_dff_A_893RPwEf4_0),.din(w_dff_A_luoqwI3p0_0),.clk(gclk));
	jdff dff_A_dZEkaBhF4_0(.dout(w_dff_A_luoqwI3p0_0),.din(w_dff_A_dZEkaBhF4_0),.clk(gclk));
	jdff dff_A_QWq5YH7x7_0(.dout(w_dff_A_dZEkaBhF4_0),.din(w_dff_A_QWq5YH7x7_0),.clk(gclk));
	jdff dff_A_s3FmS4px5_0(.dout(w_n80_0[0]),.din(w_dff_A_s3FmS4px5_0),.clk(gclk));
	jdff dff_A_2z1I5Puz3_0(.dout(w_dff_A_s3FmS4px5_0),.din(w_dff_A_2z1I5Puz3_0),.clk(gclk));
	jdff dff_A_ULD4DwGY1_0(.dout(w_dff_A_2z1I5Puz3_0),.din(w_dff_A_ULD4DwGY1_0),.clk(gclk));
	jdff dff_A_VeGUxuiq8_0(.dout(w_dff_A_ULD4DwGY1_0),.din(w_dff_A_VeGUxuiq8_0),.clk(gclk));
	jdff dff_A_ZKU1lP1t1_0(.dout(w_dff_A_VeGUxuiq8_0),.din(w_dff_A_ZKU1lP1t1_0),.clk(gclk));
	jdff dff_A_NMfp3Yml3_0(.dout(w_dff_A_ZKU1lP1t1_0),.din(w_dff_A_NMfp3Yml3_0),.clk(gclk));
	jdff dff_A_5iMHirOA5_0(.dout(w_dff_A_NMfp3Yml3_0),.din(w_dff_A_5iMHirOA5_0),.clk(gclk));
	jdff dff_A_2jtw5R4j9_0(.dout(w_dff_A_5iMHirOA5_0),.din(w_dff_A_2jtw5R4j9_0),.clk(gclk));
	jdff dff_A_EcgTezgs3_0(.dout(w_dff_A_2jtw5R4j9_0),.din(w_dff_A_EcgTezgs3_0),.clk(gclk));
	jdff dff_A_wfQ7uCxp3_0(.dout(w_dff_A_EcgTezgs3_0),.din(w_dff_A_wfQ7uCxp3_0),.clk(gclk));
	jdff dff_A_GiJdxXtb8_0(.dout(w_dff_A_wfQ7uCxp3_0),.din(w_dff_A_GiJdxXtb8_0),.clk(gclk));
	jdff dff_A_bgcdtyLP4_0(.dout(w_dff_A_GiJdxXtb8_0),.din(w_dff_A_bgcdtyLP4_0),.clk(gclk));
	jdff dff_A_0bQ4fxyL7_0(.dout(w_dff_A_bgcdtyLP4_0),.din(w_dff_A_0bQ4fxyL7_0),.clk(gclk));
	jdff dff_A_eSJpdP357_0(.dout(w_dff_A_0bQ4fxyL7_0),.din(w_dff_A_eSJpdP357_0),.clk(gclk));
	jdff dff_A_C69Ak8SM2_0(.dout(w_dff_A_eSJpdP357_0),.din(w_dff_A_C69Ak8SM2_0),.clk(gclk));
	jdff dff_A_m4p2c9nk5_0(.dout(w_dff_A_C69Ak8SM2_0),.din(w_dff_A_m4p2c9nk5_0),.clk(gclk));
	jdff dff_A_A1f7VNc53_0(.dout(w_dff_A_m4p2c9nk5_0),.din(w_dff_A_A1f7VNc53_0),.clk(gclk));
	jdff dff_A_xY1SuJ7Y7_0(.dout(w_dff_A_A1f7VNc53_0),.din(w_dff_A_xY1SuJ7Y7_0),.clk(gclk));
	jdff dff_A_INVL3gxL2_0(.dout(w_dff_A_xY1SuJ7Y7_0),.din(w_dff_A_INVL3gxL2_0),.clk(gclk));
	jdff dff_A_mziMIdWz5_0(.dout(w_dff_A_INVL3gxL2_0),.din(w_dff_A_mziMIdWz5_0),.clk(gclk));
	jdff dff_A_KULj1DkY4_0(.dout(w_dff_A_mziMIdWz5_0),.din(w_dff_A_KULj1DkY4_0),.clk(gclk));
	jdff dff_A_dZOlZMLW4_1(.dout(w_G56gat_1[1]),.din(w_dff_A_dZOlZMLW4_1),.clk(gclk));
	jdff dff_A_LVGuxcLB1_1(.dout(w_G56gat_0[1]),.din(w_dff_A_LVGuxcLB1_1),.clk(gclk));
	jdff dff_A_wmTR8ict7_1(.dout(w_dff_A_LVGuxcLB1_1),.din(w_dff_A_wmTR8ict7_1),.clk(gclk));
	jdff dff_A_yFShnhJM9_1(.dout(w_dff_A_wmTR8ict7_1),.din(w_dff_A_yFShnhJM9_1),.clk(gclk));
	jdff dff_A_ZMA7FEMY9_1(.dout(w_dff_A_yFShnhJM9_1),.din(w_dff_A_ZMA7FEMY9_1),.clk(gclk));
	jdff dff_A_qhPKt9yi6_1(.dout(w_dff_A_ZMA7FEMY9_1),.din(w_dff_A_qhPKt9yi6_1),.clk(gclk));
	jdff dff_A_ySmVm7jB4_1(.dout(w_dff_A_qhPKt9yi6_1),.din(w_dff_A_ySmVm7jB4_1),.clk(gclk));
	jdff dff_A_oiBtZd8U0_1(.dout(w_dff_A_ySmVm7jB4_1),.din(w_dff_A_oiBtZd8U0_1),.clk(gclk));
	jdff dff_A_FBpKnxet5_1(.dout(w_dff_A_oiBtZd8U0_1),.din(w_dff_A_FBpKnxet5_1),.clk(gclk));
	jdff dff_A_fYIfsCf14_1(.dout(w_dff_A_FBpKnxet5_1),.din(w_dff_A_fYIfsCf14_1),.clk(gclk));
	jdff dff_A_xozF5Ach0_1(.dout(w_dff_A_fYIfsCf14_1),.din(w_dff_A_xozF5Ach0_1),.clk(gclk));
	jdff dff_A_pdTn0NBz5_1(.dout(w_dff_A_xozF5Ach0_1),.din(w_dff_A_pdTn0NBz5_1),.clk(gclk));
	jdff dff_A_UrBp0ROh1_1(.dout(w_dff_A_pdTn0NBz5_1),.din(w_dff_A_UrBp0ROh1_1),.clk(gclk));
	jdff dff_A_SbqqBJrZ8_1(.dout(w_dff_A_UrBp0ROh1_1),.din(w_dff_A_SbqqBJrZ8_1),.clk(gclk));
	jdff dff_A_PcM4HkA08_1(.dout(w_dff_A_SbqqBJrZ8_1),.din(w_dff_A_PcM4HkA08_1),.clk(gclk));
	jdff dff_A_Ht3awnJL8_1(.dout(w_dff_A_PcM4HkA08_1),.din(w_dff_A_Ht3awnJL8_1),.clk(gclk));
	jdff dff_A_2ixDfRJv6_1(.dout(w_dff_A_Ht3awnJL8_1),.din(w_dff_A_2ixDfRJv6_1),.clk(gclk));
	jdff dff_A_j3CELniN6_1(.dout(w_dff_A_2ixDfRJv6_1),.din(w_dff_A_j3CELniN6_1),.clk(gclk));
	jdff dff_A_p3oH2QIB6_1(.dout(w_dff_A_j3CELniN6_1),.din(w_dff_A_p3oH2QIB6_1),.clk(gclk));
	jdff dff_A_c91kfoCy9_1(.dout(w_dff_A_p3oH2QIB6_1),.din(w_dff_A_c91kfoCy9_1),.clk(gclk));
	jdff dff_A_x2trJ02B9_1(.dout(w_dff_A_c91kfoCy9_1),.din(w_dff_A_x2trJ02B9_1),.clk(gclk));
	jdff dff_A_KLpJZTcl2_1(.dout(w_dff_A_x2trJ02B9_1),.din(w_dff_A_KLpJZTcl2_1),.clk(gclk));
	jdff dff_A_t52nroUK4_1(.dout(w_dff_A_KLpJZTcl2_1),.din(w_dff_A_t52nroUK4_1),.clk(gclk));
	jdff dff_A_68hQuQow0_2(.dout(w_G56gat_0[2]),.din(w_dff_A_68hQuQow0_2),.clk(gclk));
	jdff dff_A_UAyRo1Zw5_2(.dout(w_dff_A_68hQuQow0_2),.din(w_dff_A_UAyRo1Zw5_2),.clk(gclk));
	jdff dff_A_cZX06fTd3_2(.dout(w_dff_A_UAyRo1Zw5_2),.din(w_dff_A_cZX06fTd3_2),.clk(gclk));
	jdff dff_A_rhNdrFvP2_2(.dout(w_dff_A_cZX06fTd3_2),.din(w_dff_A_rhNdrFvP2_2),.clk(gclk));
	jdff dff_A_84alNLuP1_2(.dout(w_dff_A_rhNdrFvP2_2),.din(w_dff_A_84alNLuP1_2),.clk(gclk));
	jdff dff_A_3RBbZaOv7_2(.dout(w_dff_A_84alNLuP1_2),.din(w_dff_A_3RBbZaOv7_2),.clk(gclk));
	jdff dff_A_HM7Xt9M00_2(.dout(w_dff_A_3RBbZaOv7_2),.din(w_dff_A_HM7Xt9M00_2),.clk(gclk));
	jdff dff_A_sns6gJAF5_0(.dout(w_G50gat_0[0]),.din(w_dff_A_sns6gJAF5_0),.clk(gclk));
	jdff dff_A_ygNnZWiE9_0(.dout(w_n78_0[0]),.din(w_dff_A_ygNnZWiE9_0),.clk(gclk));
	jdff dff_A_UYxhPOTK9_0(.dout(w_dff_A_ygNnZWiE9_0),.din(w_dff_A_UYxhPOTK9_0),.clk(gclk));
	jdff dff_A_OstBHuum1_0(.dout(w_dff_A_UYxhPOTK9_0),.din(w_dff_A_OstBHuum1_0),.clk(gclk));
	jdff dff_A_LXonWnii7_0(.dout(w_dff_A_OstBHuum1_0),.din(w_dff_A_LXonWnii7_0),.clk(gclk));
	jdff dff_A_ReADckMX0_0(.dout(w_dff_A_LXonWnii7_0),.din(w_dff_A_ReADckMX0_0),.clk(gclk));
	jdff dff_A_4tjV6s9y4_0(.dout(w_dff_A_ReADckMX0_0),.din(w_dff_A_4tjV6s9y4_0),.clk(gclk));
	jdff dff_A_44Q1Hx1w5_0(.dout(w_G30gat_0[0]),.din(w_dff_A_44Q1Hx1w5_0),.clk(gclk));
	jdff dff_A_ErKFxt4K2_0(.dout(w_dff_A_44Q1Hx1w5_0),.din(w_dff_A_ErKFxt4K2_0),.clk(gclk));
	jdff dff_A_l0mWy9y61_0(.dout(w_dff_A_ErKFxt4K2_0),.din(w_dff_A_l0mWy9y61_0),.clk(gclk));
	jdff dff_A_QmPZJawy2_0(.dout(w_dff_A_l0mWy9y61_0),.din(w_dff_A_QmPZJawy2_0),.clk(gclk));
	jdff dff_A_mVgvovWA6_0(.dout(w_dff_A_QmPZJawy2_0),.din(w_dff_A_mVgvovWA6_0),.clk(gclk));
	jdff dff_A_s7Pv9KOO4_0(.dout(w_dff_A_mVgvovWA6_0),.din(w_dff_A_s7Pv9KOO4_0),.clk(gclk));
	jdff dff_A_TclB1t9Z4_0(.dout(w_dff_A_s7Pv9KOO4_0),.din(w_dff_A_TclB1t9Z4_0),.clk(gclk));
	jdff dff_A_GkEWWy088_2(.dout(w_G30gat_0[2]),.din(w_dff_A_GkEWWy088_2),.clk(gclk));
	jdff dff_A_VhMnQ70e8_0(.dout(w_G24gat_0[0]),.din(w_dff_A_VhMnQ70e8_0),.clk(gclk));
	jdff dff_A_RbLgk9ah9_0(.dout(w_dff_A_VhMnQ70e8_0),.din(w_dff_A_RbLgk9ah9_0),.clk(gclk));
	jdff dff_A_NcyuVqO52_0(.dout(w_dff_A_RbLgk9ah9_0),.din(w_dff_A_NcyuVqO52_0),.clk(gclk));
	jdff dff_A_FKAcYUAm7_0(.dout(w_dff_A_NcyuVqO52_0),.din(w_dff_A_FKAcYUAm7_0),.clk(gclk));
	jdff dff_A_cLWxCmsI0_0(.dout(w_dff_A_FKAcYUAm7_0),.din(w_dff_A_cLWxCmsI0_0),.clk(gclk));
	jdff dff_A_w7lt1dcp9_0(.dout(w_dff_A_cLWxCmsI0_0),.din(w_dff_A_w7lt1dcp9_0),.clk(gclk));
	jdff dff_A_AuOKD7660_1(.dout(w_G24gat_0[1]),.din(w_dff_A_AuOKD7660_1),.clk(gclk));
	jdff dff_A_LaLU8o9Q5_0(.dout(w_n75_0[0]),.din(w_dff_A_LaLU8o9Q5_0),.clk(gclk));
	jdff dff_A_CCVTszga5_0(.dout(w_dff_A_LaLU8o9Q5_0),.din(w_dff_A_CCVTszga5_0),.clk(gclk));
	jdff dff_A_52ov8LUL3_0(.dout(w_dff_A_CCVTszga5_0),.din(w_dff_A_52ov8LUL3_0),.clk(gclk));
	jdff dff_A_tN7AdNdI6_0(.dout(w_dff_A_52ov8LUL3_0),.din(w_dff_A_tN7AdNdI6_0),.clk(gclk));
	jdff dff_A_HE4889sh5_0(.dout(w_dff_A_tN7AdNdI6_0),.din(w_dff_A_HE4889sh5_0),.clk(gclk));
	jdff dff_A_jCXMQBrh3_0(.dout(w_dff_A_HE4889sh5_0),.din(w_dff_A_jCXMQBrh3_0),.clk(gclk));
	jdff dff_A_1r8vJFC17_0(.dout(w_G17gat_0[0]),.din(w_dff_A_1r8vJFC17_0),.clk(gclk));
	jdff dff_A_5hpQmw7i6_0(.dout(w_dff_A_1r8vJFC17_0),.din(w_dff_A_5hpQmw7i6_0),.clk(gclk));
	jdff dff_A_Y53OLZNa4_0(.dout(w_dff_A_5hpQmw7i6_0),.din(w_dff_A_Y53OLZNa4_0),.clk(gclk));
	jdff dff_A_VqdGLU0k9_0(.dout(w_dff_A_Y53OLZNa4_0),.din(w_dff_A_VqdGLU0k9_0),.clk(gclk));
	jdff dff_A_VUb1qwie9_0(.dout(w_dff_A_VqdGLU0k9_0),.din(w_dff_A_VUb1qwie9_0),.clk(gclk));
	jdff dff_A_i1HZzGEE2_0(.dout(w_dff_A_VUb1qwie9_0),.din(w_dff_A_i1HZzGEE2_0),.clk(gclk));
	jdff dff_A_KATBrZG45_0(.dout(w_dff_A_i1HZzGEE2_0),.din(w_dff_A_KATBrZG45_0),.clk(gclk));
	jdff dff_A_2GQp74W96_2(.dout(w_G17gat_0[2]),.din(w_dff_A_2GQp74W96_2),.clk(gclk));
	jdff dff_A_oZF4Mh1o2_0(.dout(w_G11gat_0[0]),.din(w_dff_A_oZF4Mh1o2_0),.clk(gclk));
	jdff dff_A_DC01FJdH6_0(.dout(w_dff_A_oZF4Mh1o2_0),.din(w_dff_A_DC01FJdH6_0),.clk(gclk));
	jdff dff_A_2N3DnU7i7_0(.dout(w_dff_A_DC01FJdH6_0),.din(w_dff_A_2N3DnU7i7_0),.clk(gclk));
	jdff dff_A_gyI1bUZ51_0(.dout(w_dff_A_2N3DnU7i7_0),.din(w_dff_A_gyI1bUZ51_0),.clk(gclk));
	jdff dff_A_e7Fk9voQ8_0(.dout(w_dff_A_gyI1bUZ51_0),.din(w_dff_A_e7Fk9voQ8_0),.clk(gclk));
	jdff dff_A_X0lqFf1U5_0(.dout(w_dff_A_e7Fk9voQ8_0),.din(w_dff_A_X0lqFf1U5_0),.clk(gclk));
	jdff dff_A_asY2EJUK6_1(.dout(w_G11gat_0[1]),.din(w_dff_A_asY2EJUK6_1),.clk(gclk));
	jdff dff_A_iICP0BMf4_0(.dout(w_n73_0[0]),.din(w_dff_A_iICP0BMf4_0),.clk(gclk));
	jdff dff_A_5Q2BFT2c6_0(.dout(w_dff_A_iICP0BMf4_0),.din(w_dff_A_5Q2BFT2c6_0),.clk(gclk));
	jdff dff_A_cSSoVR0x0_0(.dout(w_dff_A_5Q2BFT2c6_0),.din(w_dff_A_cSSoVR0x0_0),.clk(gclk));
	jdff dff_A_tH7PkBp22_0(.dout(w_dff_A_cSSoVR0x0_0),.din(w_dff_A_tH7PkBp22_0),.clk(gclk));
	jdff dff_A_BvclH8Jb5_0(.dout(w_dff_A_tH7PkBp22_0),.din(w_dff_A_BvclH8Jb5_0),.clk(gclk));
	jdff dff_A_DfSg4lqe1_0(.dout(w_dff_A_BvclH8Jb5_0),.din(w_dff_A_DfSg4lqe1_0),.clk(gclk));
	jdff dff_A_pOArUeeG7_0(.dout(w_G69gat_0[0]),.din(w_dff_A_pOArUeeG7_0),.clk(gclk));
	jdff dff_A_kAOLIRaY0_0(.dout(w_dff_A_pOArUeeG7_0),.din(w_dff_A_kAOLIRaY0_0),.clk(gclk));
	jdff dff_A_A8Ooo5bE8_0(.dout(w_dff_A_kAOLIRaY0_0),.din(w_dff_A_A8Ooo5bE8_0),.clk(gclk));
	jdff dff_A_hKHameyp3_0(.dout(w_dff_A_A8Ooo5bE8_0),.din(w_dff_A_hKHameyp3_0),.clk(gclk));
	jdff dff_A_Jtk8u1bt3_0(.dout(w_dff_A_hKHameyp3_0),.din(w_dff_A_Jtk8u1bt3_0),.clk(gclk));
	jdff dff_A_UnP2Bxod0_0(.dout(w_dff_A_Jtk8u1bt3_0),.din(w_dff_A_UnP2Bxod0_0),.clk(gclk));
	jdff dff_A_7wRvwOcp8_0(.dout(w_dff_A_UnP2Bxod0_0),.din(w_dff_A_7wRvwOcp8_0),.clk(gclk));
	jdff dff_A_CDaLzzUH4_2(.dout(w_G69gat_0[2]),.din(w_dff_A_CDaLzzUH4_2),.clk(gclk));
	jdff dff_A_EMEt9F877_0(.dout(w_n46_0[0]),.din(w_dff_A_EMEt9F877_0),.clk(gclk));
	jdff dff_A_vP4Y4k477_0(.dout(w_dff_A_EMEt9F877_0),.din(w_dff_A_vP4Y4k477_0),.clk(gclk));
	jdff dff_A_ZQ72B3iZ6_0(.dout(w_dff_A_vP4Y4k477_0),.din(w_dff_A_ZQ72B3iZ6_0),.clk(gclk));
	jdff dff_A_B7Epgujb4_0(.dout(w_dff_A_ZQ72B3iZ6_0),.din(w_dff_A_B7Epgujb4_0),.clk(gclk));
	jdff dff_A_ywAkzHm66_1(.dout(w_n46_0[1]),.din(w_dff_A_ywAkzHm66_1),.clk(gclk));
	jdff dff_B_Ml2pD0BU8_1(.din(G37gat),.dout(w_dff_B_Ml2pD0BU8_1),.clk(gclk));
	jdff dff_A_Gv5iyWLq3_0(.dout(w_n45_0[0]),.din(w_dff_A_Gv5iyWLq3_0),.clk(gclk));
	jdff dff_A_OQjvPBdC0_0(.dout(w_dff_A_Gv5iyWLq3_0),.din(w_dff_A_OQjvPBdC0_0),.clk(gclk));
	jdff dff_A_FDkYign09_0(.dout(w_dff_A_OQjvPBdC0_0),.din(w_dff_A_FDkYign09_0),.clk(gclk));
	jdff dff_A_Q0N3R1ey1_0(.dout(w_dff_A_FDkYign09_0),.din(w_dff_A_Q0N3R1ey1_0),.clk(gclk));
	jdff dff_A_sOhfZZak9_0(.dout(w_dff_A_Q0N3R1ey1_0),.din(w_dff_A_sOhfZZak9_0),.clk(gclk));
	jdff dff_A_q6JCB2dB3_0(.dout(w_dff_A_sOhfZZak9_0),.din(w_dff_A_q6JCB2dB3_0),.clk(gclk));
	jdff dff_A_XNVAdMtj9_0(.dout(w_G43gat_0[0]),.din(w_dff_A_XNVAdMtj9_0),.clk(gclk));
	jdff dff_A_GRRshK6s2_0(.dout(w_dff_A_XNVAdMtj9_0),.din(w_dff_A_GRRshK6s2_0),.clk(gclk));
	jdff dff_A_gyc3Z5Gb4_0(.dout(w_dff_A_GRRshK6s2_0),.din(w_dff_A_gyc3Z5Gb4_0),.clk(gclk));
	jdff dff_A_PXIAEZS05_0(.dout(w_dff_A_gyc3Z5Gb4_0),.din(w_dff_A_PXIAEZS05_0),.clk(gclk));
	jdff dff_A_qgQcvee10_0(.dout(w_dff_A_PXIAEZS05_0),.din(w_dff_A_qgQcvee10_0),.clk(gclk));
	jdff dff_A_wbdwtidA6_0(.dout(w_dff_A_qgQcvee10_0),.din(w_dff_A_wbdwtidA6_0),.clk(gclk));
	jdff dff_A_MieW2VVm4_0(.dout(w_dff_A_wbdwtidA6_0),.din(w_dff_A_MieW2VVm4_0),.clk(gclk));
	jdff dff_A_ebpXr9Hh7_1(.dout(w_n44_0[1]),.din(w_dff_A_ebpXr9Hh7_1),.clk(gclk));
	jdff dff_A_NucbvHI39_1(.dout(w_G108gat_0[1]),.din(w_dff_A_NucbvHI39_1),.clk(gclk));
	jdff dff_A_iWOI8SEZ1_1(.dout(w_dff_A_NucbvHI39_1),.din(w_dff_A_iWOI8SEZ1_1),.clk(gclk));
	jdff dff_A_MbjdOFz08_1(.dout(w_dff_A_iWOI8SEZ1_1),.din(w_dff_A_MbjdOFz08_1),.clk(gclk));
	jdff dff_A_gvY4XCXn2_1(.dout(w_dff_A_MbjdOFz08_1),.din(w_dff_A_gvY4XCXn2_1),.clk(gclk));
	jdff dff_A_SH013tnM8_1(.dout(w_dff_A_gvY4XCXn2_1),.din(w_dff_A_SH013tnM8_1),.clk(gclk));
	jdff dff_A_IAtl95gj8_1(.dout(w_dff_A_SH013tnM8_1),.din(w_dff_A_IAtl95gj8_1),.clk(gclk));
	jdff dff_A_W3svUPV46_1(.dout(w_dff_A_IAtl95gj8_1),.din(w_dff_A_W3svUPV46_1),.clk(gclk));
	jdff dff_A_4i46PGmI0_2(.dout(w_G108gat_0[2]),.din(w_dff_A_4i46PGmI0_2),.clk(gclk));
	jdff dff_A_xAe2rTE61_0(.dout(w_n43_0[0]),.din(w_dff_A_xAe2rTE61_0),.clk(gclk));
	jdff dff_A_2znjptDJ4_0(.dout(w_dff_A_xAe2rTE61_0),.din(w_dff_A_2znjptDJ4_0),.clk(gclk));
	jdff dff_A_UfIjYvQB1_0(.dout(w_dff_A_2znjptDJ4_0),.din(w_dff_A_UfIjYvQB1_0),.clk(gclk));
	jdff dff_A_TNcbctzq1_0(.dout(w_dff_A_UfIjYvQB1_0),.din(w_dff_A_TNcbctzq1_0),.clk(gclk));
	jdff dff_A_YwwioSY85_0(.dout(w_dff_A_TNcbctzq1_0),.din(w_dff_A_YwwioSY85_0),.clk(gclk));
	jdff dff_A_N65usaMv8_0(.dout(w_G102gat_0[0]),.din(w_dff_A_N65usaMv8_0),.clk(gclk));
	jdff dff_A_45DDNgtQ3_0(.dout(w_dff_A_N65usaMv8_0),.din(w_dff_A_45DDNgtQ3_0),.clk(gclk));
	jdff dff_A_o6ixDT2s2_0(.dout(w_dff_A_45DDNgtQ3_0),.din(w_dff_A_o6ixDT2s2_0),.clk(gclk));
	jdff dff_A_pz45IahK8_0(.dout(w_dff_A_o6ixDT2s2_0),.din(w_dff_A_pz45IahK8_0),.clk(gclk));
	jdff dff_A_JaxLAtvC3_0(.dout(w_dff_A_pz45IahK8_0),.din(w_dff_A_JaxLAtvC3_0),.clk(gclk));
	jdff dff_A_70y3XZk07_0(.dout(w_dff_A_JaxLAtvC3_0),.din(w_dff_A_70y3XZk07_0),.clk(gclk));
	jdff dff_A_WfdLipTW7_0(.dout(w_n49_0[0]),.din(w_dff_A_WfdLipTW7_0),.clk(gclk));
	jdff dff_A_cnpsrrmk0_0(.dout(w_dff_A_WfdLipTW7_0),.din(w_dff_A_cnpsrrmk0_0),.clk(gclk));
	jdff dff_A_mWIZI3vw2_0(.dout(w_dff_A_cnpsrrmk0_0),.din(w_dff_A_mWIZI3vw2_0),.clk(gclk));
	jdff dff_A_9vXIbKq39_0(.dout(w_dff_A_mWIZI3vw2_0),.din(w_dff_A_9vXIbKq39_0),.clk(gclk));
	jdff dff_A_zUzEfCVk4_0(.dout(w_dff_A_9vXIbKq39_0),.din(w_dff_A_zUzEfCVk4_0),.clk(gclk));
	jdff dff_A_81gjaSbA7_0(.dout(w_G63gat_0[0]),.din(w_dff_A_81gjaSbA7_0),.clk(gclk));
	jdff dff_A_ojfR0qZ85_0(.dout(w_dff_A_81gjaSbA7_0),.din(w_dff_A_ojfR0qZ85_0),.clk(gclk));
	jdff dff_A_bgSF60ae4_0(.dout(w_dff_A_ojfR0qZ85_0),.din(w_dff_A_bgSF60ae4_0),.clk(gclk));
	jdff dff_A_7z1ywyqd3_0(.dout(w_dff_A_bgSF60ae4_0),.din(w_dff_A_7z1ywyqd3_0),.clk(gclk));
	jdff dff_A_ObiHwby38_0(.dout(w_dff_A_7z1ywyqd3_0),.din(w_dff_A_ObiHwby38_0),.clk(gclk));
	jdff dff_A_usOypx327_0(.dout(w_dff_A_ObiHwby38_0),.din(w_dff_A_usOypx327_0),.clk(gclk));
	jdff dff_A_zdoTkP3m3_1(.dout(w_G63gat_0[1]),.din(w_dff_A_zdoTkP3m3_1),.clk(gclk));
	jdff dff_A_SEMGl6Zg8_1(.dout(w_dff_A_FgI7NOuD4_0),.din(w_dff_A_SEMGl6Zg8_1),.clk(gclk));
	jdff dff_A_FgI7NOuD4_0(.dout(w_dff_A_W85J9Emz9_0),.din(w_dff_A_FgI7NOuD4_0),.clk(gclk));
	jdff dff_A_W85J9Emz9_0(.dout(w_dff_A_6RXb5wTr2_0),.din(w_dff_A_W85J9Emz9_0),.clk(gclk));
	jdff dff_A_6RXb5wTr2_0(.dout(w_dff_A_yAs7j40J5_0),.din(w_dff_A_6RXb5wTr2_0),.clk(gclk));
	jdff dff_A_yAs7j40J5_0(.dout(w_dff_A_nxGMixCD4_0),.din(w_dff_A_yAs7j40J5_0),.clk(gclk));
	jdff dff_A_nxGMixCD4_0(.dout(w_dff_A_iBZzaS8T9_0),.din(w_dff_A_nxGMixCD4_0),.clk(gclk));
	jdff dff_A_iBZzaS8T9_0(.dout(w_dff_A_fo5d3vHc4_0),.din(w_dff_A_iBZzaS8T9_0),.clk(gclk));
	jdff dff_A_fo5d3vHc4_0(.dout(w_dff_A_cxMmrtHl2_0),.din(w_dff_A_fo5d3vHc4_0),.clk(gclk));
	jdff dff_A_cxMmrtHl2_0(.dout(w_dff_A_jEd241Z64_0),.din(w_dff_A_cxMmrtHl2_0),.clk(gclk));
	jdff dff_A_jEd241Z64_0(.dout(w_dff_A_uHCETZMJ0_0),.din(w_dff_A_jEd241Z64_0),.clk(gclk));
	jdff dff_A_uHCETZMJ0_0(.dout(w_dff_A_mIpwl0R25_0),.din(w_dff_A_uHCETZMJ0_0),.clk(gclk));
	jdff dff_A_mIpwl0R25_0(.dout(w_dff_A_KSXBSmRr2_0),.din(w_dff_A_mIpwl0R25_0),.clk(gclk));
	jdff dff_A_KSXBSmRr2_0(.dout(w_dff_A_HrY8qfug8_0),.din(w_dff_A_KSXBSmRr2_0),.clk(gclk));
	jdff dff_A_HrY8qfug8_0(.dout(w_dff_A_F6lggsDY0_0),.din(w_dff_A_HrY8qfug8_0),.clk(gclk));
	jdff dff_A_F6lggsDY0_0(.dout(w_dff_A_5ANkbwFV0_0),.din(w_dff_A_F6lggsDY0_0),.clk(gclk));
	jdff dff_A_5ANkbwFV0_0(.dout(w_dff_A_bl0NvcbN2_0),.din(w_dff_A_5ANkbwFV0_0),.clk(gclk));
	jdff dff_A_bl0NvcbN2_0(.dout(w_dff_A_fU2MW94j0_0),.din(w_dff_A_bl0NvcbN2_0),.clk(gclk));
	jdff dff_A_fU2MW94j0_0(.dout(w_dff_A_N81KYzpx5_0),.din(w_dff_A_fU2MW94j0_0),.clk(gclk));
	jdff dff_A_N81KYzpx5_0(.dout(w_dff_A_8gq10dYw0_0),.din(w_dff_A_N81KYzpx5_0),.clk(gclk));
	jdff dff_A_8gq10dYw0_0(.dout(w_dff_A_7QgaQTST6_0),.din(w_dff_A_8gq10dYw0_0),.clk(gclk));
	jdff dff_A_7QgaQTST6_0(.dout(G223gat),.din(w_dff_A_7QgaQTST6_0),.clk(gclk));
	jdff dff_A_n8EDLT5F7_1(.dout(w_dff_A_g5CDUu0d0_0),.din(w_dff_A_n8EDLT5F7_1),.clk(gclk));
	jdff dff_A_g5CDUu0d0_0(.dout(w_dff_A_QGRhmXyi2_0),.din(w_dff_A_g5CDUu0d0_0),.clk(gclk));
	jdff dff_A_QGRhmXyi2_0(.dout(w_dff_A_046ZAo3f0_0),.din(w_dff_A_QGRhmXyi2_0),.clk(gclk));
	jdff dff_A_046ZAo3f0_0(.dout(w_dff_A_p08ej82O1_0),.din(w_dff_A_046ZAo3f0_0),.clk(gclk));
	jdff dff_A_p08ej82O1_0(.dout(w_dff_A_CSDyzqPJ5_0),.din(w_dff_A_p08ej82O1_0),.clk(gclk));
	jdff dff_A_CSDyzqPJ5_0(.dout(w_dff_A_NrCqfr6e4_0),.din(w_dff_A_CSDyzqPJ5_0),.clk(gclk));
	jdff dff_A_NrCqfr6e4_0(.dout(w_dff_A_yhzrV6pF0_0),.din(w_dff_A_NrCqfr6e4_0),.clk(gclk));
	jdff dff_A_yhzrV6pF0_0(.dout(w_dff_A_lrl24h1E3_0),.din(w_dff_A_yhzrV6pF0_0),.clk(gclk));
	jdff dff_A_lrl24h1E3_0(.dout(w_dff_A_43gH8nQM2_0),.din(w_dff_A_lrl24h1E3_0),.clk(gclk));
	jdff dff_A_43gH8nQM2_0(.dout(w_dff_A_qXojXBgN6_0),.din(w_dff_A_43gH8nQM2_0),.clk(gclk));
	jdff dff_A_qXojXBgN6_0(.dout(w_dff_A_9FNc9TVV7_0),.din(w_dff_A_qXojXBgN6_0),.clk(gclk));
	jdff dff_A_9FNc9TVV7_0(.dout(w_dff_A_UuQOzaaV8_0),.din(w_dff_A_9FNc9TVV7_0),.clk(gclk));
	jdff dff_A_UuQOzaaV8_0(.dout(w_dff_A_p8mRBsUd9_0),.din(w_dff_A_UuQOzaaV8_0),.clk(gclk));
	jdff dff_A_p8mRBsUd9_0(.dout(G329gat),.din(w_dff_A_p8mRBsUd9_0),.clk(gclk));
	jdff dff_A_yBeS5tNQ7_2(.dout(w_dff_A_a9rIOCa60_0),.din(w_dff_A_yBeS5tNQ7_2),.clk(gclk));
	jdff dff_A_a9rIOCa60_0(.dout(w_dff_A_aDqauZ9T3_0),.din(w_dff_A_a9rIOCa60_0),.clk(gclk));
	jdff dff_A_aDqauZ9T3_0(.dout(w_dff_A_u0dyAunK0_0),.din(w_dff_A_aDqauZ9T3_0),.clk(gclk));
	jdff dff_A_u0dyAunK0_0(.dout(w_dff_A_KTsi93jF9_0),.din(w_dff_A_u0dyAunK0_0),.clk(gclk));
	jdff dff_A_KTsi93jF9_0(.dout(w_dff_A_iswhRiWp5_0),.din(w_dff_A_KTsi93jF9_0),.clk(gclk));
	jdff dff_A_iswhRiWp5_0(.dout(w_dff_A_z3jNHQMA0_0),.din(w_dff_A_iswhRiWp5_0),.clk(gclk));
	jdff dff_A_z3jNHQMA0_0(.dout(G370gat),.din(w_dff_A_z3jNHQMA0_0),.clk(gclk));
	jdff dff_A_azFe6ujw4_1(.dout(w_dff_A_2cvsLWe78_0),.din(w_dff_A_azFe6ujw4_1),.clk(gclk));
	jdff dff_A_2cvsLWe78_0(.dout(G430gat),.din(w_dff_A_2cvsLWe78_0),.clk(gclk));
endmodule

