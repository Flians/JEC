/*

c1355:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jcb: 6
	jdff: 449
	jand: 65

Summary:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jcb: 6
	jdff: 449
	jand: 65
*/

module c1355(gclk, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat, G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat, G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat, G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat, G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat, G1352gat, G1353gat, G1354gat, G1355gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G15gat;
	input G22gat;
	input G29gat;
	input G36gat;
	input G43gat;
	input G50gat;
	input G57gat;
	input G64gat;
	input G71gat;
	input G78gat;
	input G85gat;
	input G92gat;
	input G99gat;
	input G106gat;
	input G113gat;
	input G120gat;
	input G127gat;
	input G134gat;
	input G141gat;
	input G148gat;
	input G155gat;
	input G162gat;
	input G169gat;
	input G176gat;
	input G183gat;
	input G190gat;
	input G197gat;
	input G204gat;
	input G211gat;
	input G218gat;
	input G225gat;
	input G226gat;
	input G227gat;
	input G228gat;
	input G229gat;
	input G230gat;
	input G231gat;
	input G232gat;
	input G233gat;
	output G1324gat;
	output G1325gat;
	output G1326gat;
	output G1327gat;
	output G1328gat;
	output G1329gat;
	output G1330gat;
	output G1331gat;
	output G1332gat;
	output G1333gat;
	output G1334gat;
	output G1335gat;
	output G1336gat;
	output G1337gat;
	output G1338gat;
	output G1339gat;
	output G1340gat;
	output G1341gat;
	output G1342gat;
	output G1343gat;
	output G1344gat;
	output G1345gat;
	output G1346gat;
	output G1347gat;
	output G1348gat;
	output G1349gat;
	output G1350gat;
	output G1351gat;
	output G1352gat;
	output G1353gat;
	output G1354gat;
	output G1355gat;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n179;
	wire n180;
	wire n182;
	wire n183;
	wire n185;
	wire n186;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n194;
	wire n196;
	wire n198;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n206;
	wire n208;
	wire n210;
	wire n212;
	wire n213;
	wire n215;
	wire n217;
	wire n219;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n234;
	wire n236;
	wire n238;
	wire n240;
	wire n241;
	wire n242;
	wire n244;
	wire n246;
	wire n248;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n255;
	wire n257;
	wire n259;
	wire n261;
	wire n262;
	wire n264;
	wire n266;
	wire n268;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G8gat_0;
	wire [2:0] w_G15gat_0;
	wire [2:0] w_G22gat_0;
	wire [2:0] w_G29gat_0;
	wire [2:0] w_G36gat_0;
	wire [2:0] w_G43gat_0;
	wire [2:0] w_G50gat_0;
	wire [2:0] w_G57gat_0;
	wire [2:0] w_G64gat_0;
	wire [2:0] w_G71gat_0;
	wire [2:0] w_G78gat_0;
	wire [2:0] w_G85gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G99gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G113gat_0;
	wire [2:0] w_G120gat_0;
	wire [2:0] w_G127gat_0;
	wire [2:0] w_G134gat_0;
	wire [2:0] w_G141gat_0;
	wire [2:0] w_G148gat_0;
	wire [2:0] w_G155gat_0;
	wire [2:0] w_G162gat_0;
	wire [2:0] w_G169gat_0;
	wire [2:0] w_G176gat_0;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G190gat_0;
	wire [2:0] w_G197gat_0;
	wire [2:0] w_G204gat_0;
	wire [2:0] w_G211gat_0;
	wire [2:0] w_G218gat_0;
	wire [2:0] w_G233gat_0;
	wire [2:0] w_G233gat_1;
	wire [1:0] w_n79_0;
	wire [1:0] w_n85_0;
	wire [2:0] w_n87_0;
	wire [1:0] w_n87_1;
	wire [2:0] w_n88_0;
	wire [2:0] w_n88_1;
	wire [1:0] w_n94_0;
	wire [2:0] w_n97_0;
	wire [1:0] w_n97_1;
	wire [1:0] w_n101_0;
	wire [2:0] w_n103_0;
	wire [1:0] w_n103_1;
	wire [1:0] w_n109_0;
	wire [1:0] w_n115_0;
	wire [2:0] w_n117_0;
	wire [1:0] w_n117_1;
	wire [2:0] w_n118_0;
	wire [2:0] w_n118_1;
	wire [1:0] w_n119_0;
	wire [1:0] w_n125_0;
	wire [1:0] w_n131_0;
	wire [2:0] w_n133_0;
	wire [1:0] w_n133_1;
	wire [2:0] w_n142_0;
	wire [1:0] w_n142_1;
	wire [2:0] w_n150_0;
	wire [1:0] w_n150_1;
	wire [2:0] w_n156_0;
	wire [2:0] w_n164_0;
	wire [1:0] w_n164_1;
	wire [2:0] w_n165_0;
	wire [2:0] w_n165_1;
	wire [2:0] w_n173_0;
	wire [1:0] w_n173_1;
	wire [1:0] w_n174_0;
	wire [2:0] w_n176_0;
	wire [1:0] w_n176_1;
	wire [2:0] w_n179_0;
	wire [2:0] w_n179_1;
	wire [2:0] w_n182_0;
	wire [2:0] w_n182_1;
	wire [2:0] w_n185_0;
	wire [2:0] w_n185_1;
	wire [2:0] w_n188_0;
	wire [2:0] w_n188_1;
	wire [1:0] w_n190_0;
	wire [2:0] w_n191_0;
	wire [1:0] w_n191_1;
	wire [2:0] w_n200_0;
	wire [2:0] w_n200_1;
	wire [1:0] w_n201_0;
	wire [2:0] w_n203_0;
	wire [1:0] w_n203_1;
	wire [2:0] w_n212_0;
	wire [1:0] w_n212_1;
	wire [1:0] w_n221_0;
	wire [1:0] w_n229_0;
	wire [1:0] w_n230_0;
	wire [2:0] w_n231_0;
	wire [1:0] w_n231_1;
	wire [1:0] w_n240_0;
	wire [2:0] w_n241_0;
	wire [1:0] w_n241_1;
	wire [1:0] w_n251_0;
	wire [2:0] w_n252_0;
	wire [1:0] w_n252_1;
	wire [2:0] w_n261_0;
	wire [1:0] w_n261_1;
	wire w_dff_A_vdPcnTFX3_0;
	wire w_dff_B_r8FJVIJ24_2;
	wire w_dff_A_hRCJFKgL4_1;
	wire w_dff_B_UWBylWK54_2;
	wire w_dff_B_7Cck4rhx1_2;
	wire w_dff_B_BNLlAz3j6_2;
	wire w_dff_B_qUrfu9jW1_0;
	wire w_dff_B_owl8iB525_1;
	wire w_dff_A_lGAB4W7I8_0;
	wire w_dff_A_UTvZTO7I7_0;
	wire w_dff_A_dpigLNVm3_0;
	wire w_dff_A_qSiySCfX4_0;
	wire w_dff_A_gU9C9yEW4_0;
	wire w_dff_A_uw7ucNNN1_0;
	wire w_dff_A_7Be8AeBF8_1;
	wire w_dff_A_Ui5HdkiS3_1;
	wire w_dff_A_QrBhabZh9_1;
	wire w_dff_A_bKsqmj1W5_1;
	wire w_dff_A_d6agRoYl7_0;
	wire w_dff_A_NZ7vswYn4_0;
	wire w_dff_A_DTeIsMUa0_0;
	wire w_dff_A_Yw9zhwJZ6_0;
	wire w_dff_A_Yh9lxLTl9_1;
	wire w_dff_A_GaqwIUbM1_1;
	wire w_dff_A_iEzGq03t6_1;
	wire w_dff_A_FezvLLFD3_1;
	wire w_dff_A_HVymXHBn8_0;
	wire w_dff_A_3jIiPkuY9_0;
	wire w_dff_A_sJw7kvzQ3_0;
	wire w_dff_A_p1148UTE1_0;
	wire w_dff_A_OOM77HGc5_1;
	wire w_dff_A_hfqDjlSn7_1;
	wire w_dff_A_XpX6X2mh5_1;
	wire w_dff_A_jylKDbSY7_1;
	wire w_dff_B_BgaXxk1H8_1;
	wire w_dff_A_TmkUtfMt5_0;
	wire w_dff_A_2vQDDBMR5_0;
	wire w_dff_A_K9FeKXkR0_0;
	wire w_dff_A_cOd908YV2_0;
	wire w_dff_A_YygD2thL4_2;
	wire w_dff_A_w1kJl7rA1_2;
	wire w_dff_A_auMrjeNo8_2;
	wire w_dff_A_DcTjdZYh3_2;
	wire w_dff_A_Inlo5oks1_0;
	wire w_dff_A_qPeFRIWT1_0;
	wire w_dff_A_3Mvle7Tq3_0;
	wire w_dff_A_JkHF1v2x3_0;
	wire w_dff_A_2VwTkvX12_1;
	wire w_dff_A_0zWqIJsV5_1;
	wire w_dff_A_1jIi0ivv1_1;
	wire w_dff_A_Sge4AOLm8_1;
	wire w_dff_B_IehodlcR5_2;
	wire w_dff_B_A8fCb3Nv3_2;
	wire w_dff_A_0ZLYMpt93_0;
	wire w_dff_A_qu6ztY5D1_0;
	wire w_dff_A_flIgCFXO2_0;
	wire w_dff_A_oAScp9vP1_0;
	wire w_dff_A_cci19hNq5_2;
	wire w_dff_A_3HIlSwSn5_2;
	wire w_dff_A_4Ju04hih4_2;
	wire w_dff_A_yFAt378D6_2;
	wire w_dff_A_c8UqvpQi4_1;
	wire w_dff_A_Y9q25Hs56_1;
	wire w_dff_A_5NEjFakf1_1;
	wire w_dff_A_j2oGcDX49_1;
	wire w_dff_A_54LPtYOM0_2;
	wire w_dff_A_TBZ1rb6v5_2;
	wire w_dff_A_0sagchlM8_2;
	wire w_dff_A_43cGsIwN6_2;
	wire w_dff_A_QRus6GbE7_0;
	wire w_dff_A_HR8rokqC6_1;
	wire w_dff_A_QpLUy2g79_1;
	wire w_dff_A_H1abPuNI0_1;
	wire w_dff_A_0ViuaRIr7_1;
	wire w_dff_A_PEgZkBLG6_2;
	wire w_dff_A_EEsZ9AwR2_2;
	wire w_dff_A_LzL16HWy4_2;
	wire w_dff_A_pQGFEaYd0_2;
	wire w_dff_A_GHrb1CeX8_1;
	wire w_dff_A_HzaJ06GZ9_1;
	wire w_dff_A_1AgXO7ki6_1;
	wire w_dff_A_aulwWU2G9_1;
	wire w_dff_A_qBWieEza7_1;
	wire w_dff_A_rjjrpJgt2_2;
	wire w_dff_A_zc9hvvMt9_2;
	wire w_dff_A_NEYxA4Vr7_2;
	wire w_dff_A_9gXtwih81_2;
	wire w_dff_A_yru3O2PL1_0;
	wire w_dff_B_FOpXhkhO3_1;
	wire w_dff_B_w00ffTJc9_0;
	wire w_dff_B_1n0vBH7l2_1;
	wire w_dff_A_ET4d4aUP5_2;
	wire w_dff_A_RNt34pof7_2;
	wire w_dff_A_RE71uI073_2;
	wire w_dff_A_z5ik1pbm6_0;
	wire w_dff_A_JtFH7GZw0_0;
	wire w_dff_A_hlD9GBci7_0;
	wire w_dff_A_DxHEB6cJ1_0;
	wire w_dff_A_imgJg5xS1_2;
	wire w_dff_A_v3McqeVC7_2;
	wire w_dff_A_KycxdNdu5_2;
	wire w_dff_A_CjlEWrLC3_2;
	wire w_dff_A_NOx3pkQq9_1;
	wire w_dff_A_YhQXZeI68_0;
	wire w_dff_A_1iUUqMce3_0;
	wire w_dff_A_sulxPjQc9_0;
	wire w_dff_A_ZRU7skZH6_0;
	wire w_dff_A_86JC351g8_0;
	wire w_dff_A_jQ4qLKjT1_0;
	wire w_dff_A_qi7AQSsh8_0;
	wire w_dff_A_I6dWuaU49_0;
	wire w_dff_A_MtHr3Kaq5_0;
	wire w_dff_A_RnARyNcU7_0;
	wire w_dff_A_ZySGaYA15_0;
	wire w_dff_A_d9WF0F7t5_0;
	wire w_dff_A_0CGjDb7w0_0;
	wire w_dff_A_0IJJrDDU9_0;
	wire w_dff_A_efdEqy2z8_0;
	wire w_dff_A_zBCtljCk0_0;
	wire w_dff_A_q2raEr044_0;
	wire w_dff_A_VMvjioiq2_0;
	wire w_dff_A_n7wLgPXX5_0;
	wire w_dff_A_6ofuZSxw0_0;
	wire w_dff_A_5SFFyfvI3_1;
	wire w_dff_A_BfXk90y80_2;
	wire w_dff_A_bedMVhhi9_0;
	wire w_dff_A_N0P3wn1K3_0;
	wire w_dff_A_OFLk40Xe9_0;
	wire w_dff_A_GSWiFwCq8_0;
	wire w_dff_A_SDCfabFB9_0;
	wire w_dff_A_KXgaq1yM2_0;
	wire w_dff_A_LK6DEAa72_0;
	wire w_dff_A_C9oQZRvw3_0;
	wire w_dff_A_WEFQwI8F3_0;
	wire w_dff_A_eodqpG4e5_0;
	wire w_dff_A_ktA7mwbm7_0;
	wire w_dff_A_5DkprJcj8_0;
	wire w_dff_A_9lv3Amie2_0;
	wire w_dff_A_tuJ8xmcg2_0;
	wire w_dff_A_BLnz5Epy3_0;
	wire w_dff_A_IssG3zlj8_0;
	wire w_dff_A_Jnsshwon5_0;
	wire w_dff_A_2m3yCjbj1_0;
	wire w_dff_A_ApktT6vx1_0;
	wire w_dff_A_q7DjgNRJ8_0;
	wire w_dff_B_9LmMrDv48_2;
	wire w_dff_B_E1H7gFcr9_2;
	wire w_dff_A_B6URFRbq9_0;
	wire w_dff_A_NddPX5cX2_0;
	wire w_dff_A_ABv4K3DA1_0;
	wire w_dff_A_TuXQfG4X9_0;
	wire w_dff_A_8dVzED9r0_2;
	wire w_dff_A_KlEUMlVr0_2;
	wire w_dff_A_dum3mdWz3_2;
	wire w_dff_A_OTPAWWJ69_2;
	wire w_dff_A_CKvDnEw04_1;
	wire w_dff_B_q9oyvLJJ6_0;
	wire w_dff_A_lOLlEOb58_0;
	wire w_dff_A_mM24LcMB6_0;
	wire w_dff_A_6vkJHhZs1_0;
	wire w_dff_A_cwU9WSZM9_0;
	wire w_dff_A_uK3IhWNC8_0;
	wire w_dff_A_nOG9BSCP4_0;
	wire w_dff_A_Y5lBGqJ05_0;
	wire w_dff_A_VIJiJCyq6_0;
	wire w_dff_A_xrVHGazt6_0;
	wire w_dff_A_IH5t9iYx6_0;
	wire w_dff_A_UGnvSxT39_0;
	wire w_dff_A_xpi9CXyb3_0;
	wire w_dff_A_frFC1J7Q2_0;
	wire w_dff_A_fJuxviOY2_0;
	wire w_dff_A_47to3FvV1_0;
	wire w_dff_A_OircruCZ0_0;
	wire w_dff_A_6WLlouUT9_0;
	wire w_dff_A_RpfDDlFo6_0;
	wire w_dff_A_VHaVAnIW9_0;
	wire w_dff_A_gHSCOu0H3_0;
	wire w_dff_A_xE6xDtaC4_0;
	wire w_dff_A_J5WdBcqk6_0;
	wire w_dff_A_lnajIqec4_0;
	wire w_dff_A_sf4y9oYY9_0;
	wire w_dff_A_VhGPRo4X9_0;
	wire w_dff_A_tF6ERLtR4_0;
	wire w_dff_A_YYzIuxGT1_0;
	wire w_dff_A_bq72miS85_0;
	wire w_dff_A_WWjmO0TC2_0;
	wire w_dff_A_A1pMQ3Hm9_0;
	wire w_dff_A_p7USBnxT4_0;
	wire w_dff_A_UapwwjJo4_0;
	wire w_dff_A_B0ewAVea1_0;
	wire w_dff_A_JaToxVeE5_0;
	wire w_dff_A_9DIBqpjA1_0;
	wire w_dff_A_R3jQqNUW5_0;
	wire w_dff_A_oLRS4jul9_0;
	wire w_dff_A_Zd8H5dRg1_0;
	wire w_dff_A_j66GuRiM8_0;
	wire w_dff_A_W3c8usBA7_0;
	wire w_dff_A_9nyimzTq6_0;
	wire w_dff_A_vtR8LFjb2_0;
	wire w_dff_A_NHUrFMKO0_0;
	wire w_dff_A_S7GBDa9p6_0;
	wire w_dff_A_GcX1QMaQ6_0;
	wire w_dff_A_ct0PvfPt1_0;
	wire w_dff_A_PFr7EWCL5_0;
	wire w_dff_A_80VcY0VA5_0;
	wire w_dff_A_AbDVtYd55_0;
	wire w_dff_A_aihb3rzW4_0;
	wire w_dff_A_JHNkrrkt6_0;
	wire w_dff_A_EffmJLfU4_0;
	wire w_dff_A_L6XCZfzh4_0;
	wire w_dff_A_0XEFr1mJ0_0;
	wire w_dff_A_ZDWXEuLp0_0;
	wire w_dff_A_wJBJlFIN9_0;
	wire w_dff_A_fyAQG2qW5_0;
	wire w_dff_A_U61K6byg2_0;
	wire w_dff_A_bby7G3um4_0;
	wire w_dff_A_lp3Apxky4_0;
	wire w_dff_A_gP1fpRqZ8_0;
	wire w_dff_A_LlpRzyEu7_0;
	wire w_dff_A_Ju18mdtB7_0;
	wire w_dff_A_jKuVhO7H9_0;
	wire w_dff_A_RFGsi2yE6_0;
	wire w_dff_A_yVntB7KN0_0;
	wire w_dff_A_AJQpFf6c2_0;
	wire w_dff_A_7Ebkt2Cy9_0;
	wire w_dff_A_g0UO8wW58_0;
	wire w_dff_A_QGzJNjho4_0;
	wire w_dff_A_FoARUN5b2_0;
	wire w_dff_A_Ij0lj3FY2_0;
	wire w_dff_A_uXUcPjyI4_0;
	wire w_dff_A_NOZUmB3r9_0;
	wire w_dff_A_unqp0OXJ2_0;
	wire w_dff_A_LyHyXneI0_0;
	wire w_dff_A_vVsZFM9R9_0;
	wire w_dff_A_mdjorY9t5_0;
	wire w_dff_A_Nm8hYCEe7_0;
	wire w_dff_A_16R7wHZT0_0;
	wire w_dff_A_9qXqSa537_1;
	wire w_dff_B_NbjDkQI86_0;
	wire w_dff_A_KiFH5kca6_0;
	wire w_dff_A_WXZVXrH93_0;
	wire w_dff_A_WcAG9DI67_0;
	wire w_dff_A_mg8rkEyR8_0;
	wire w_dff_A_TNOiG2DB9_0;
	wire w_dff_A_U71FEFkk9_0;
	wire w_dff_A_kYSyubT59_0;
	wire w_dff_A_wIbPCJM10_0;
	wire w_dff_A_4bjXMHAC1_0;
	wire w_dff_A_888GxPFd1_0;
	wire w_dff_A_EAvaAVwd9_0;
	wire w_dff_A_Y83I1f5Q7_0;
	wire w_dff_A_tDnMmOMw2_0;
	wire w_dff_A_f43pz4dJ4_0;
	wire w_dff_A_ZBiGlx7o4_0;
	wire w_dff_A_z6Pxcvfe2_0;
	wire w_dff_A_Un8zDzAg9_0;
	wire w_dff_A_XbydEyyt1_0;
	wire w_dff_A_wKgpVQdz7_0;
	wire w_dff_A_UeBD4cLQ8_0;
	wire w_dff_A_lNzLxEo71_0;
	wire w_dff_A_21Nq3TIT9_0;
	wire w_dff_A_bKM8lDHK4_0;
	wire w_dff_A_nZ63Rjea4_0;
	wire w_dff_A_ocj7L1Z45_0;
	wire w_dff_A_YO9xdqZR3_0;
	wire w_dff_A_nkADfmy61_0;
	wire w_dff_A_2CLsx5uI0_0;
	wire w_dff_A_QXrEgSM40_0;
	wire w_dff_A_QOW4o5NL8_0;
	wire w_dff_A_9UWkVhLH5_0;
	wire w_dff_A_ayISePTn6_0;
	wire w_dff_A_OZi5rbvL0_0;
	wire w_dff_A_QQojFK2U1_0;
	wire w_dff_A_M1uRzLfT9_0;
	wire w_dff_A_Q3zomeuh1_0;
	wire w_dff_A_emCous512_0;
	wire w_dff_A_T9HaHUw18_0;
	wire w_dff_A_zfRI8mNA3_0;
	wire w_dff_A_62ez2TRR5_0;
	wire w_dff_A_4OA0Gfg71_0;
	wire w_dff_A_hVfAd7SZ0_0;
	wire w_dff_A_fj8u79Wu6_0;
	wire w_dff_A_iq55yZHa1_0;
	wire w_dff_A_tbexwx929_0;
	wire w_dff_A_I1gdxe1m7_0;
	wire w_dff_A_1LiiKV618_0;
	wire w_dff_A_dihKoGgo0_0;
	wire w_dff_A_ILkwBy1f5_0;
	wire w_dff_A_TMb2lijH8_0;
	wire w_dff_A_CTXvQAYN3_0;
	wire w_dff_A_7OBGOj2w8_0;
	wire w_dff_A_hni43xyM4_0;
	wire w_dff_A_VwyN0akb0_0;
	wire w_dff_A_AVSdgegI6_0;
	wire w_dff_A_52PZheCw3_0;
	wire w_dff_A_8J6VeEuK7_0;
	wire w_dff_A_V6g4VQdq1_0;
	wire w_dff_A_E0BAUg2T6_0;
	wire w_dff_A_8JaEixeq4_0;
	wire w_dff_A_WCYXH9172_0;
	wire w_dff_A_tuEIIjdG2_0;
	wire w_dff_A_DiQ4yvs05_0;
	wire w_dff_A_6394ptkw4_0;
	wire w_dff_A_hs4t52pc0_0;
	wire w_dff_A_GZX8HBgJ8_0;
	wire w_dff_A_Pai67DP20_0;
	wire w_dff_A_UIW96QiQ1_0;
	wire w_dff_A_xcG2OLcu9_0;
	wire w_dff_A_wQEy2KyV0_0;
	wire w_dff_A_5nYDEzEt4_0;
	wire w_dff_A_ksfwVJTC7_0;
	wire w_dff_A_odu2dyA62_0;
	wire w_dff_A_Xz7dIdf21_0;
	wire w_dff_A_6Wv0SJQa4_0;
	wire w_dff_A_5a8LTbLo0_0;
	wire w_dff_A_4QBemBD09_0;
	wire w_dff_A_pupSgkaY3_0;
	wire w_dff_A_k2FiQ56T2_0;
	wire w_dff_A_Hq3tDri10_0;
	wire w_dff_A_0D4s2Gdo9_1;
	wire w_dff_A_6uaFYpQ50_1;
	wire w_dff_A_08ryss2d4_1;
	wire w_dff_A_yaIGEDZr2_1;
	wire w_dff_A_WGMDp3wy0_2;
	wire w_dff_A_nNydAWo07_2;
	wire w_dff_A_QC21nsqe6_2;
	wire w_dff_A_2jSnBeHT6_2;
	wire w_dff_A_GA9OqbVz5_1;
	wire w_dff_B_Xo319tDN4_1;
	wire w_dff_A_hSz9sN5M7_0;
	wire w_dff_A_yIlyZ2qw9_0;
	wire w_dff_A_6A89NvFf1_0;
	wire w_dff_A_XHVa2PdQ6_0;
	wire w_dff_A_GSgHsgiB4_0;
	wire w_dff_A_ZUy2e09b2_0;
	wire w_dff_A_5GamDoKq7_0;
	wire w_dff_A_RVpORlXa0_0;
	wire w_dff_A_0zdwHsLo0_0;
	wire w_dff_A_N9GJF8Yq0_0;
	wire w_dff_A_7ogGRhSk8_0;
	wire w_dff_A_epMiw4AP8_0;
	wire w_dff_A_kJhRpB537_0;
	wire w_dff_A_n6irMDDe0_0;
	wire w_dff_A_fFBhEhC89_0;
	wire w_dff_A_7FKm4skU2_0;
	wire w_dff_A_CZbXNoCq5_0;
	wire w_dff_A_s69AW2Fs6_0;
	wire w_dff_A_0LwUw7DL4_0;
	wire w_dff_A_NTUOQ2Dc1_0;
	wire w_dff_A_nH2CFQxK8_0;
	wire w_dff_A_P0pATZpu5_0;
	wire w_dff_A_CmV82uFf5_0;
	wire w_dff_A_ArnMqjTV9_0;
	wire w_dff_A_7vLI3jZR5_0;
	wire w_dff_A_cU3b97YW4_0;
	wire w_dff_A_vg3w83hV5_0;
	wire w_dff_A_ffnDFGgU1_0;
	wire w_dff_A_RpaAdJF60_0;
	wire w_dff_A_Xitz6zWQ0_0;
	wire w_dff_A_LxsrAVop3_0;
	wire w_dff_A_dWQcn0NB0_0;
	wire w_dff_A_cv1xoxRd8_0;
	wire w_dff_A_Lqqu33rW4_0;
	wire w_dff_A_ZOxxSYZV7_0;
	wire w_dff_A_vpAUhqgM5_0;
	wire w_dff_A_jPksLCYx7_0;
	wire w_dff_A_J9EUjqCr9_0;
	wire w_dff_A_seiQmn7Y2_0;
	wire w_dff_A_hQ93Wxpt5_0;
	wire w_dff_A_QdfBtJXe6_0;
	wire w_dff_A_k9ev0bn76_0;
	wire w_dff_A_6qXIiSgi8_0;
	wire w_dff_A_G9wTVSPf9_0;
	wire w_dff_A_CTfT16IF5_0;
	wire w_dff_A_ElqjSLiE6_0;
	wire w_dff_A_TzOVK7Js5_0;
	wire w_dff_A_d84snmT29_0;
	wire w_dff_A_6VTyIUdl5_0;
	wire w_dff_A_8EXb0oLX9_0;
	wire w_dff_A_DwujNDRM0_0;
	wire w_dff_A_nOS9wDOF4_0;
	wire w_dff_A_Td4g39v61_0;
	wire w_dff_A_qA4dQDjZ3_0;
	wire w_dff_A_Vy1OX6oJ6_0;
	wire w_dff_A_ViCNu6qF5_0;
	wire w_dff_A_pQiwXVJ70_0;
	wire w_dff_A_lhkC14OG6_0;
	wire w_dff_A_JT5YBbSq8_0;
	wire w_dff_A_mWGmOgUG6_0;
	wire w_dff_A_4Lr9U9Wf4_0;
	wire w_dff_A_5bLXqItI0_0;
	wire w_dff_A_qLA6ovTt7_0;
	wire w_dff_A_mXyI7v1d2_0;
	wire w_dff_A_eLZtMan07_0;
	wire w_dff_A_rP3JqqWt2_0;
	wire w_dff_A_JjetcthL6_0;
	wire w_dff_A_a0MzTrRl1_0;
	wire w_dff_A_q2xmU7879_0;
	wire w_dff_A_8iNtpnhp8_0;
	wire w_dff_A_DrKOrulf4_0;
	wire w_dff_A_dqEL3aSt9_0;
	wire w_dff_A_5fshzP8e3_0;
	wire w_dff_A_iw9woJxl2_0;
	wire w_dff_A_3mtbQBH67_0;
	wire w_dff_A_omcknDYr7_0;
	wire w_dff_A_PiXkER0f4_0;
	wire w_dff_A_pbI64Yim0_0;
	wire w_dff_A_9qY27C2D5_0;
	wire w_dff_A_M4t8SJ0K9_0;
	wire w_dff_A_aEnsqv513_0;
	wire w_dff_A_Dbdk0u5X4_0;
	wire w_dff_A_zoXouxbX3_0;
	wire w_dff_A_nI7xrFNy1_0;
	wire w_dff_A_fXfTq2In2_0;
	wire w_dff_A_LKggevtQ5_0;
	wire w_dff_A_o9NgQYoj2_0;
	wire w_dff_A_aydRc4zT7_0;
	wire w_dff_A_VO7Uf5QN5_0;
	wire w_dff_A_ePkpiFcd3_0;
	wire w_dff_A_Hy9M0DwN2_0;
	wire w_dff_A_7PMAeOua3_0;
	wire w_dff_A_9fg9i70z2_0;
	wire w_dff_A_aoAzma2Y8_0;
	wire w_dff_A_um6aLhpZ4_0;
	wire w_dff_A_gPhuAdES2_0;
	wire w_dff_A_4kILrvpf1_0;
	wire w_dff_A_XtZcJDB85_0;
	wire w_dff_A_3utV0gN68_0;
	wire w_dff_A_EBGdVPH94_0;
	wire w_dff_A_N1sW4CcE8_0;
	wire w_dff_A_oOJ2sYzY8_0;
	wire w_dff_A_nMV08u7c0_0;
	wire w_dff_A_Ga2VoN8N9_0;
	wire w_dff_A_JvPUZ4wM5_0;
	wire w_dff_A_Pe3402fb4_0;
	wire w_dff_A_5qBKOiqD8_0;
	wire w_dff_A_0uWmPsc89_0;
	wire w_dff_A_lZx38iLY4_0;
	wire w_dff_A_Mih6RlS80_0;
	wire w_dff_A_0lyfOHWN2_0;
	wire w_dff_A_wlwr0xjB8_0;
	wire w_dff_A_qfBUllui9_0;
	wire w_dff_A_L11IOaEB3_0;
	wire w_dff_A_1EMa7xGF8_0;
	wire w_dff_A_vvwYoSry0_0;
	wire w_dff_A_svDUcBLl9_0;
	wire w_dff_A_ItiD22yw2_0;
	wire w_dff_A_a15osvgB0_0;
	wire w_dff_A_rrUk5ZKY3_0;
	jxor g000(.dina(w_G85gat_0[2]),.dinb(w_G57gat_0[2]),.dout(n74),.clk(gclk));
	jxor g001(.dina(w_G29gat_0[2]),.dinb(w_G1gat_0[2]),.dout(n75),.clk(gclk));
	jxor g002(.dina(n75),.dinb(n74),.dout(n76),.clk(gclk));
	jxor g003(.dina(w_G162gat_0[2]),.dinb(w_G155gat_0[2]),.dout(n77),.clk(gclk));
	jxor g004(.dina(w_G148gat_0[2]),.dinb(w_G141gat_0[2]),.dout(n78),.clk(gclk));
	jxor g005(.dina(n78),.dinb(n77),.dout(n79),.clk(gclk));
	jxor g006(.dina(w_n79_0[1]),.dinb(n76),.dout(n80),.clk(gclk));
	jand g007(.dina(w_G233gat_1[2]),.dinb(G225gat),.dout(n81),.clk(gclk));
	jnot g008(.din(n81),.dout(n82),.clk(gclk));
	jxor g009(.dina(w_G134gat_0[2]),.dinb(w_G127gat_0[2]),.dout(n83),.clk(gclk));
	jxor g010(.dina(w_G120gat_0[2]),.dinb(w_G113gat_0[2]),.dout(n84),.clk(gclk));
	jxor g011(.dina(n84),.dinb(n83),.dout(n85),.clk(gclk));
	jxor g012(.dina(w_n85_0[1]),.dinb(n82),.dout(n86),.clk(gclk));
	jxor g013(.dina(n86),.dinb(n80),.dout(n87),.clk(gclk));
	jnot g014(.din(w_n87_1[1]),.dout(n88),.clk(gclk));
	jxor g015(.dina(w_G218gat_0[2]),.dinb(w_G190gat_0[2]),.dout(n89),.clk(gclk));
	jxor g016(.dina(w_G162gat_0[1]),.dinb(w_G134gat_0[1]),.dout(n90),.clk(gclk));
	jxor g017(.dina(n90),.dinb(n89),.dout(n91),.clk(gclk));
	jxor g018(.dina(w_G106gat_0[2]),.dinb(w_G99gat_0[2]),.dout(n92),.clk(gclk));
	jxor g019(.dina(w_G92gat_0[2]),.dinb(w_G85gat_0[1]),.dout(n93),.clk(gclk));
	jxor g020(.dina(n93),.dinb(n92),.dout(n94),.clk(gclk));
	jxor g021(.dina(w_n94_0[1]),.dinb(n91),.dout(n95),.clk(gclk));
	jnot g022(.din(G232gat),.dout(n96),.clk(gclk));
	jnot g023(.din(w_G233gat_1[1]),.dout(n97),.clk(gclk));
	jcb g024(.dina(w_n97_1[1]),.dinb(n96),.dout(n98));
	jxor g025(.dina(w_G50gat_0[2]),.dinb(w_G43gat_0[2]),.dout(n99),.clk(gclk));
	jxor g026(.dina(w_G36gat_0[2]),.dinb(w_G29gat_0[1]),.dout(n100),.clk(gclk));
	jxor g027(.dina(n100),.dinb(n99),.dout(n101),.clk(gclk));
	jxor g028(.dina(w_n101_0[1]),.dinb(w_dff_B_Xo319tDN4_1),.dout(n102),.clk(gclk));
	jxor g029(.dina(n102),.dinb(n95),.dout(n103),.clk(gclk));
	jxor g030(.dina(w_G211gat_0[2]),.dinb(w_G183gat_0[2]),.dout(n104),.clk(gclk));
	jxor g031(.dina(w_G155gat_0[1]),.dinb(w_G127gat_0[1]),.dout(n105),.clk(gclk));
	jxor g032(.dina(n105),.dinb(n104),.dout(n106),.clk(gclk));
	jxor g033(.dina(w_G78gat_0[2]),.dinb(w_G71gat_0[2]),.dout(n107),.clk(gclk));
	jxor g034(.dina(w_G64gat_0[2]),.dinb(w_G57gat_0[1]),.dout(n108),.clk(gclk));
	jxor g035(.dina(n108),.dinb(n107),.dout(n109),.clk(gclk));
	jxor g036(.dina(w_n109_0[1]),.dinb(n106),.dout(n110),.clk(gclk));
	jnot g037(.din(G231gat),.dout(n111),.clk(gclk));
	jcb g038(.dina(w_n97_1[0]),.dinb(n111),.dout(n112));
	jxor g039(.dina(w_G22gat_0[2]),.dinb(w_G15gat_0[2]),.dout(n113),.clk(gclk));
	jxor g040(.dina(w_G8gat_0[2]),.dinb(w_G1gat_0[1]),.dout(n114),.clk(gclk));
	jxor g041(.dina(n114),.dinb(n113),.dout(n115),.clk(gclk));
	jxor g042(.dina(w_n115_0[1]),.dinb(w_dff_B_1n0vBH7l2_1),.dout(n116),.clk(gclk));
	jxor g043(.dina(n116),.dinb(n110),.dout(n117),.clk(gclk));
	jnot g044(.din(w_n117_1[1]),.dout(n118),.clk(gclk));
	jand g045(.dina(w_n118_1[2]),.dinb(w_n103_1[1]),.dout(n119),.clk(gclk));
	jxor g046(.dina(w_G92gat_0[1]),.dinb(w_G64gat_0[1]),.dout(n120),.clk(gclk));
	jxor g047(.dina(w_G36gat_0[1]),.dinb(w_G8gat_0[1]),.dout(n121),.clk(gclk));
	jxor g048(.dina(n121),.dinb(n120),.dout(n122),.clk(gclk));
	jxor g049(.dina(w_G190gat_0[1]),.dinb(w_G183gat_0[1]),.dout(n123),.clk(gclk));
	jxor g050(.dina(w_G176gat_0[2]),.dinb(w_G169gat_0[2]),.dout(n124),.clk(gclk));
	jxor g051(.dina(n124),.dinb(n123),.dout(n125),.clk(gclk));
	jxor g052(.dina(w_n125_0[1]),.dinb(n122),.dout(n126),.clk(gclk));
	jand g053(.dina(w_G233gat_1[0]),.dinb(G226gat),.dout(n127),.clk(gclk));
	jnot g054(.din(n127),.dout(n128),.clk(gclk));
	jxor g055(.dina(w_G218gat_0[1]),.dinb(w_G211gat_0[1]),.dout(n129),.clk(gclk));
	jxor g056(.dina(w_G204gat_0[2]),.dinb(w_G197gat_0[2]),.dout(n130),.clk(gclk));
	jxor g057(.dina(n130),.dinb(n129),.dout(n131),.clk(gclk));
	jxor g058(.dina(w_n131_0[1]),.dinb(n128),.dout(n132),.clk(gclk));
	jxor g059(.dina(n132),.dinb(n126),.dout(n133),.clk(gclk));
	jxor g060(.dina(w_n133_1[1]),.dinb(w_n87_1[0]),.dout(n134),.clk(gclk));
	jxor g061(.dina(w_G99gat_0[1]),.dinb(w_G71gat_0[1]),.dout(n135),.clk(gclk));
	jxor g062(.dina(w_G43gat_0[1]),.dinb(w_G15gat_0[1]),.dout(n136),.clk(gclk));
	jxor g063(.dina(n136),.dinb(n135),.dout(n137),.clk(gclk));
	jxor g064(.dina(n137),.dinb(w_n125_0[0]),.dout(n138),.clk(gclk));
	jnot g065(.din(G227gat),.dout(n139),.clk(gclk));
	jcb g066(.dina(w_n97_0[2]),.dinb(n139),.dout(n140));
	jxor g067(.dina(w_dff_B_NbjDkQI86_0),.dinb(w_n85_0[0]),.dout(n141),.clk(gclk));
	jxor g068(.dina(n141),.dinb(n138),.dout(n142),.clk(gclk));
	jxor g069(.dina(w_G106gat_0[1]),.dinb(w_G78gat_0[1]),.dout(n143),.clk(gclk));
	jxor g070(.dina(w_G50gat_0[1]),.dinb(w_G22gat_0[1]),.dout(n144),.clk(gclk));
	jxor g071(.dina(n144),.dinb(n143),.dout(n145),.clk(gclk));
	jxor g072(.dina(n145),.dinb(w_n131_0[0]),.dout(n146),.clk(gclk));
	jnot g073(.din(G228gat),.dout(n147),.clk(gclk));
	jcb g074(.dina(w_n97_0[1]),.dinb(n147),.dout(n148));
	jxor g075(.dina(w_dff_B_q9oyvLJJ6_0),.dinb(w_n79_0[0]),.dout(n149),.clk(gclk));
	jxor g076(.dina(n149),.dinb(n146),.dout(n150),.clk(gclk));
	jand g077(.dina(w_n150_1[1]),.dinb(w_n142_1[1]),.dout(n151),.clk(gclk));
	jand g078(.dina(n151),.dinb(n134),.dout(n152),.clk(gclk));
	jxor g079(.dina(w_n150_1[0]),.dinb(w_n142_1[0]),.dout(n153),.clk(gclk));
	jand g080(.dina(n153),.dinb(w_n87_0[2]),.dout(n154),.clk(gclk));
	jand g081(.dina(n154),.dinb(w_n133_1[0]),.dout(n155),.clk(gclk));
	jcb g082(.dina(n155),.dinb(w_dff_B_owl8iB525_1),.dout(n156));
	jxor g083(.dina(w_G197gat_0[1]),.dinb(w_G169gat_0[1]),.dout(n157),.clk(gclk));
	jxor g084(.dina(w_G141gat_0[1]),.dinb(w_G113gat_0[1]),.dout(n158),.clk(gclk));
	jxor g085(.dina(n158),.dinb(n157),.dout(n159),.clk(gclk));
	jxor g086(.dina(n159),.dinb(w_n115_0[0]),.dout(n160),.clk(gclk));
	jand g087(.dina(w_G233gat_0[2]),.dinb(G229gat),.dout(n161),.clk(gclk));
	jnot g088(.din(n161),.dout(n162),.clk(gclk));
	jxor g089(.dina(n162),.dinb(w_n101_0[0]),.dout(n163),.clk(gclk));
	jxor g090(.dina(n163),.dinb(n160),.dout(n164),.clk(gclk));
	jnot g091(.din(w_n164_1[1]),.dout(n165),.clk(gclk));
	jxor g092(.dina(w_G204gat_0[1]),.dinb(w_G176gat_0[1]),.dout(n166),.clk(gclk));
	jxor g093(.dina(w_G148gat_0[1]),.dinb(w_G120gat_0[1]),.dout(n167),.clk(gclk));
	jxor g094(.dina(n167),.dinb(n166),.dout(n168),.clk(gclk));
	jxor g095(.dina(n168),.dinb(w_n109_0[0]),.dout(n169),.clk(gclk));
	jand g096(.dina(w_G233gat_0[1]),.dinb(G230gat),.dout(n170),.clk(gclk));
	jnot g097(.din(n170),.dout(n171),.clk(gclk));
	jxor g098(.dina(n171),.dinb(w_n94_0[0]),.dout(n172),.clk(gclk));
	jxor g099(.dina(n172),.dinb(n169),.dout(n173),.clk(gclk));
	jand g100(.dina(w_n173_1[1]),.dinb(w_n165_1[2]),.dout(n174),.clk(gclk));
	jand g101(.dina(w_n174_0[1]),.dinb(w_n156_0[2]),.dout(n175),.clk(gclk));
	jand g102(.dina(n175),.dinb(w_n119_0[1]),.dout(n176),.clk(gclk));
	jand g103(.dina(w_n176_1[1]),.dinb(w_n88_1[2]),.dout(n177),.clk(gclk));
	jxor g104(.dina(n177),.dinb(w_G1gat_0[0]),.dout(G1324gat),.clk(gclk));
	jnot g105(.din(w_n133_0[2]),.dout(n179),.clk(gclk));
	jand g106(.dina(w_n176_1[0]),.dinb(w_n179_1[2]),.dout(n180),.clk(gclk));
	jxor g107(.dina(n180),.dinb(w_G8gat_0[0]),.dout(G1325gat),.clk(gclk));
	jnot g108(.din(w_n142_0[2]),.dout(n182),.clk(gclk));
	jand g109(.dina(w_n176_0[2]),.dinb(w_n182_1[2]),.dout(n183),.clk(gclk));
	jxor g110(.dina(n183),.dinb(w_G15gat_0[0]),.dout(G1326gat),.clk(gclk));
	jnot g111(.din(w_n150_0[2]),.dout(n185),.clk(gclk));
	jand g112(.dina(w_n176_0[1]),.dinb(w_n185_1[2]),.dout(n186),.clk(gclk));
	jxor g113(.dina(n186),.dinb(w_G22gat_0[0]),.dout(G1327gat),.clk(gclk));
	jnot g114(.din(w_n103_1[0]),.dout(n188),.clk(gclk));
	jand g115(.dina(w_n117_1[0]),.dinb(w_n188_1[2]),.dout(n189),.clk(gclk));
	jand g116(.dina(w_dff_B_qUrfu9jW1_0),.dinb(w_n156_0[1]),.dout(n190),.clk(gclk));
	jand g117(.dina(w_n190_0[1]),.dinb(w_n174_0[0]),.dout(n191),.clk(gclk));
	jand g118(.dina(w_n191_1[1]),.dinb(w_n88_1[1]),.dout(n192),.clk(gclk));
	jxor g119(.dina(n192),.dinb(w_G29gat_0[0]),.dout(G1328gat),.clk(gclk));
	jand g120(.dina(w_n191_1[0]),.dinb(w_n179_1[1]),.dout(n194),.clk(gclk));
	jxor g121(.dina(n194),.dinb(w_G36gat_0[0]),.dout(G1329gat),.clk(gclk));
	jand g122(.dina(w_n191_0[2]),.dinb(w_n182_1[1]),.dout(n196),.clk(gclk));
	jxor g123(.dina(n196),.dinb(w_G43gat_0[0]),.dout(G1330gat),.clk(gclk));
	jand g124(.dina(w_n191_0[1]),.dinb(w_n185_1[1]),.dout(n198),.clk(gclk));
	jxor g125(.dina(n198),.dinb(w_G50gat_0[0]),.dout(G1331gat),.clk(gclk));
	jnot g126(.din(w_n173_1[0]),.dout(n200),.clk(gclk));
	jand g127(.dina(w_n200_1[2]),.dinb(w_n164_1[0]),.dout(n201),.clk(gclk));
	jand g128(.dina(w_n156_0[0]),.dinb(w_n119_0[0]),.dout(n202),.clk(gclk));
	jand g129(.dina(n202),.dinb(w_n201_0[1]),.dout(n203),.clk(gclk));
	jand g130(.dina(w_n203_1[1]),.dinb(w_n88_1[0]),.dout(n204),.clk(gclk));
	jxor g131(.dina(n204),.dinb(w_G57gat_0[0]),.dout(G1332gat),.clk(gclk));
	jand g132(.dina(w_n203_1[0]),.dinb(w_n179_1[0]),.dout(n206),.clk(gclk));
	jxor g133(.dina(n206),.dinb(w_G64gat_0[0]),.dout(G1333gat),.clk(gclk));
	jand g134(.dina(w_n203_0[2]),.dinb(w_n182_1[0]),.dout(n208),.clk(gclk));
	jxor g135(.dina(n208),.dinb(w_G71gat_0[0]),.dout(G1334gat),.clk(gclk));
	jand g136(.dina(w_n203_0[1]),.dinb(w_n185_1[0]),.dout(n210),.clk(gclk));
	jxor g137(.dina(n210),.dinb(w_G78gat_0[0]),.dout(G1335gat),.clk(gclk));
	jand g138(.dina(w_n201_0[0]),.dinb(w_n190_0[0]),.dout(n212),.clk(gclk));
	jand g139(.dina(w_n212_1[1]),.dinb(w_n88_0[2]),.dout(n213),.clk(gclk));
	jxor g140(.dina(n213),.dinb(w_G85gat_0[0]),.dout(G1336gat),.clk(gclk));
	jand g141(.dina(w_n212_1[0]),.dinb(w_n179_0[2]),.dout(n215),.clk(gclk));
	jxor g142(.dina(n215),.dinb(w_G92gat_0[0]),.dout(G1337gat),.clk(gclk));
	jand g143(.dina(w_n212_0[2]),.dinb(w_n182_0[2]),.dout(n217),.clk(gclk));
	jxor g144(.dina(n217),.dinb(w_G99gat_0[0]),.dout(G1338gat),.clk(gclk));
	jand g145(.dina(w_n212_0[1]),.dinb(w_n185_0[2]),.dout(n219),.clk(gclk));
	jxor g146(.dina(n219),.dinb(w_G106gat_0[0]),.dout(G1339gat),.clk(gclk));
	jand g147(.dina(w_n150_0[1]),.dinb(w_n182_0[1]),.dout(n221),.clk(gclk));
	jand g148(.dina(w_n133_0[1]),.dinb(w_n88_0[1]),.dout(n222),.clk(gclk));
	jxor g149(.dina(w_n117_0[2]),.dinb(w_n103_0[2]),.dout(n223),.clk(gclk));
	jand g150(.dina(n223),.dinb(w_n164_0[2]),.dout(n224),.clk(gclk));
	jand g151(.dina(n224),.dinb(w_n173_0[2]),.dout(n225),.clk(gclk));
	jxor g152(.dina(w_n173_0[1]),.dinb(w_n164_0[1]),.dout(n226),.clk(gclk));
	jand g153(.dina(w_n117_0[1]),.dinb(w_n103_0[1]),.dout(n227),.clk(gclk));
	jand g154(.dina(n227),.dinb(n226),.dout(n228),.clk(gclk));
	jcb g155(.dina(w_dff_B_w00ffTJc9_0),.dinb(n225),.dout(n229));
	jand g156(.dina(w_n229_0[1]),.dinb(w_dff_B_BgaXxk1H8_1),.dout(n230),.clk(gclk));
	jand g157(.dina(w_n230_0[1]),.dinb(w_n221_0[1]),.dout(n231),.clk(gclk));
	jand g158(.dina(w_n231_1[1]),.dinb(w_n165_1[1]),.dout(n232),.clk(gclk));
	jxor g159(.dina(n232),.dinb(w_G113gat_0[0]),.dout(G1340gat),.clk(gclk));
	jand g160(.dina(w_n231_1[0]),.dinb(w_n200_1[1]),.dout(n234),.clk(gclk));
	jxor g161(.dina(n234),.dinb(w_G120gat_0[0]),.dout(G1341gat),.clk(gclk));
	jand g162(.dina(w_n231_0[2]),.dinb(w_n118_1[1]),.dout(n236),.clk(gclk));
	jxor g163(.dina(n236),.dinb(w_G127gat_0[0]),.dout(G1342gat),.clk(gclk));
	jand g164(.dina(w_n231_0[1]),.dinb(w_n188_1[1]),.dout(n238),.clk(gclk));
	jxor g165(.dina(n238),.dinb(w_G134gat_0[0]),.dout(G1343gat),.clk(gclk));
	jand g166(.dina(w_n185_0[1]),.dinb(w_n142_0[1]),.dout(n240),.clk(gclk));
	jand g167(.dina(w_n230_0[0]),.dinb(w_n240_0[1]),.dout(n241),.clk(gclk));
	jand g168(.dina(w_n241_1[1]),.dinb(w_n165_1[0]),.dout(n242),.clk(gclk));
	jxor g169(.dina(n242),.dinb(w_G141gat_0[0]),.dout(G1344gat),.clk(gclk));
	jand g170(.dina(w_n241_1[0]),.dinb(w_n200_1[0]),.dout(n244),.clk(gclk));
	jxor g171(.dina(n244),.dinb(w_G148gat_0[0]),.dout(G1345gat),.clk(gclk));
	jand g172(.dina(w_n241_0[2]),.dinb(w_n118_1[0]),.dout(n246),.clk(gclk));
	jxor g173(.dina(n246),.dinb(w_G155gat_0[0]),.dout(G1346gat),.clk(gclk));
	jand g174(.dina(w_n241_0[1]),.dinb(w_n188_1[0]),.dout(n248),.clk(gclk));
	jxor g175(.dina(n248),.dinb(w_G162gat_0[0]),.dout(G1347gat),.clk(gclk));
	jand g176(.dina(w_n179_0[1]),.dinb(w_n87_0[1]),.dout(n250),.clk(gclk));
	jand g177(.dina(w_n229_0[0]),.dinb(w_dff_B_FOpXhkhO3_1),.dout(n251),.clk(gclk));
	jand g178(.dina(w_n251_0[1]),.dinb(w_n221_0[0]),.dout(n252),.clk(gclk));
	jand g179(.dina(w_n252_1[1]),.dinb(w_n165_0[2]),.dout(n253),.clk(gclk));
	jxor g180(.dina(n253),.dinb(w_G169gat_0[0]),.dout(G1348gat),.clk(gclk));
	jand g181(.dina(w_n252_1[0]),.dinb(w_n200_0[2]),.dout(n255),.clk(gclk));
	jxor g182(.dina(n255),.dinb(w_G176gat_0[0]),.dout(G1349gat),.clk(gclk));
	jand g183(.dina(w_n252_0[2]),.dinb(w_n118_0[2]),.dout(n257),.clk(gclk));
	jxor g184(.dina(n257),.dinb(w_G183gat_0[0]),.dout(G1350gat),.clk(gclk));
	jand g185(.dina(w_n252_0[1]),.dinb(w_n188_0[2]),.dout(n259),.clk(gclk));
	jxor g186(.dina(n259),.dinb(w_G190gat_0[0]),.dout(G1351gat),.clk(gclk));
	jand g187(.dina(w_n251_0[0]),.dinb(w_n240_0[0]),.dout(n261),.clk(gclk));
	jand g188(.dina(w_n261_1[1]),.dinb(w_n165_0[1]),.dout(n262),.clk(gclk));
	jxor g189(.dina(n262),.dinb(w_G197gat_0[0]),.dout(G1352gat),.clk(gclk));
	jand g190(.dina(w_n261_1[0]),.dinb(w_n200_0[1]),.dout(n264),.clk(gclk));
	jxor g191(.dina(n264),.dinb(w_G204gat_0[0]),.dout(G1353gat),.clk(gclk));
	jand g192(.dina(w_n261_0[2]),.dinb(w_n118_0[1]),.dout(n266),.clk(gclk));
	jxor g193(.dina(n266),.dinb(w_G211gat_0[0]),.dout(G1354gat),.clk(gclk));
	jand g194(.dina(w_n261_0[1]),.dinb(w_n188_0[1]),.dout(n268),.clk(gclk));
	jxor g195(.dina(n268),.dinb(w_G218gat_0[0]),.dout(G1355gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_eodqpG4e5_0),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_RnARyNcU7_0),.doutb(w_G8gat_0[1]),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G15gat_0(.douta(w_dff_A_62ez2TRR5_0),.doutb(w_G15gat_0[1]),.doutc(w_G15gat_0[2]),.din(G15gat));
	jspl3 jspl3_w_G22gat_0(.douta(w_dff_A_W3c8usBA7_0),.doutb(w_G22gat_0[1]),.doutc(w_G22gat_0[2]),.din(G22gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_dff_A_NTUOQ2Dc1_0),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl3 jspl3_w_G36gat_0(.douta(w_dff_A_N9GJF8Yq0_0),.doutb(w_G36gat_0[1]),.doutc(w_G36gat_0[2]),.din(G36gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_dff_A_hQ93Wxpt5_0),.doutb(w_G43gat_0[1]),.doutc(w_G43gat_0[2]),.din(G43gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_dff_A_Xitz6zWQ0_0),.doutb(w_G50gat_0[1]),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl3 jspl3_w_G57gat_0(.douta(w_dff_A_q7DjgNRJ8_0),.doutb(w_G57gat_0[1]),.doutc(w_G57gat_0[2]),.din(G57gat));
	jspl3 jspl3_w_G64gat_0(.douta(w_dff_A_6ofuZSxw0_0),.doutb(w_G64gat_0[1]),.doutc(w_G64gat_0[2]),.din(G64gat));
	jspl3 jspl3_w_G71gat_0(.douta(w_dff_A_TMb2lijH8_0),.doutb(w_G71gat_0[1]),.doutc(w_G71gat_0[2]),.din(G71gat));
	jspl3 jspl3_w_G78gat_0(.douta(w_dff_A_aihb3rzW4_0),.doutb(w_G78gat_0[1]),.doutc(w_G78gat_0[2]),.din(G78gat));
	jspl3 jspl3_w_G85gat_0(.douta(w_dff_A_mWGmOgUG6_0),.doutb(w_G85gat_0[1]),.doutc(w_G85gat_0[2]),.din(G85gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_8EXb0oLX9_0),.doutb(w_G92gat_0[1]),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_M4t8SJ0K9_0),.doutb(w_G99gat_0[1]),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_8iNtpnhp8_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G113gat_0(.douta(w_dff_A_UeBD4cLQ8_0),.doutb(w_G113gat_0[1]),.doutc(w_G113gat_0[2]),.din(G113gat));
	jspl3 jspl3_w_G120gat_0(.douta(w_dff_A_888GxPFd1_0),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G127gat_0(.douta(w_dff_A_QOW4o5NL8_0),.doutb(w_G127gat_0[1]),.doutc(w_G127gat_0[2]),.din(G127gat));
	jspl3 jspl3_w_G134gat_0(.douta(w_dff_A_EBGdVPH94_0),.doutb(w_G134gat_0[1]),.doutc(w_G134gat_0[2]),.din(G134gat));
	jspl3 jspl3_w_G141gat_0(.douta(w_dff_A_gHSCOu0H3_0),.doutb(w_G141gat_0[1]),.doutc(w_G141gat_0[2]),.din(G141gat));
	jspl3 jspl3_w_G148gat_0(.douta(w_dff_A_IH5t9iYx6_0),.doutb(w_G148gat_0[1]),.doutc(w_G148gat_0[2]),.din(G148gat));
	jspl3 jspl3_w_G155gat_0(.douta(w_dff_A_A1pMQ3Hm9_0),.doutb(w_G155gat_0[1]),.doutc(w_G155gat_0[2]),.din(G155gat));
	jspl3 jspl3_w_G162gat_0(.douta(w_dff_A_ePkpiFcd3_0),.doutb(w_G162gat_0[1]),.doutc(w_G162gat_0[2]),.din(G162gat));
	jspl3 jspl3_w_G169gat_0(.douta(w_dff_A_wQEy2KyV0_0),.doutb(w_G169gat_0[1]),.doutc(w_G169gat_0[2]),.din(G169gat));
	jspl3 jspl3_w_G176gat_0(.douta(w_dff_A_8JaEixeq4_0),.doutb(w_G176gat_0[1]),.doutc(w_G176gat_0[2]),.din(G176gat));
	jspl3 jspl3_w_G183gat_0(.douta(w_dff_A_Hq3tDri10_0),.doutb(w_G183gat_0[1]),.doutc(w_G183gat_0[2]),.din(G183gat));
	jspl3 jspl3_w_G190gat_0(.douta(w_dff_A_rrUk5ZKY3_0),.doutb(w_G190gat_0[1]),.doutc(w_G190gat_0[2]),.din(G190gat));
	jspl3 jspl3_w_G197gat_0(.douta(w_dff_A_QGzJNjho4_0),.doutb(w_G197gat_0[1]),.doutc(w_G197gat_0[2]),.din(G197gat));
	jspl3 jspl3_w_G204gat_0(.douta(w_dff_A_lp3Apxky4_0),.doutb(w_G204gat_0[1]),.doutc(w_G204gat_0[2]),.din(G204gat));
	jspl3 jspl3_w_G211gat_0(.douta(w_dff_A_16R7wHZT0_0),.doutb(w_G211gat_0[1]),.doutc(w_G211gat_0[2]),.din(G211gat));
	jspl3 jspl3_w_G218gat_0(.douta(w_dff_A_Mih6RlS80_0),.doutb(w_G218gat_0[1]),.doutc(w_G218gat_0[2]),.din(G218gat));
	jspl3 jspl3_w_G233gat_0(.douta(w_G233gat_0[0]),.doutb(w_G233gat_0[1]),.doutc(w_G233gat_0[2]),.din(G233gat));
	jspl3 jspl3_w_G233gat_1(.douta(w_G233gat_1[0]),.doutb(w_G233gat_1[1]),.doutc(w_G233gat_1[2]),.din(w_G233gat_0[0]));
	jspl jspl_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.din(n79));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl3 jspl3_w_n87_0(.douta(w_n87_0[0]),.doutb(w_dff_A_5SFFyfvI3_1),.doutc(w_dff_A_BfXk90y80_2),.din(n87));
	jspl jspl_w_n87_1(.douta(w_n87_1[0]),.doutb(w_n87_1[1]),.din(w_n87_0[0]));
	jspl3 jspl3_w_n88_0(.douta(w_dff_A_cOd908YV2_0),.doutb(w_n88_0[1]),.doutc(w_dff_A_DcTjdZYh3_2),.din(n88));
	jspl3 jspl3_w_n88_1(.douta(w_n88_1[0]),.doutb(w_n88_1[1]),.doutc(w_n88_1[2]),.din(w_n88_0[0]));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.doutc(w_n97_0[2]),.din(n97));
	jspl jspl_w_n97_1(.douta(w_n97_1[0]),.doutb(w_n97_1[1]),.din(w_n97_0[0]));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.doutc(w_n103_0[2]),.din(n103));
	jspl jspl_w_n103_1(.douta(w_n103_1[0]),.doutb(w_dff_A_GA9OqbVz5_1),.din(w_n103_0[0]));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl jspl_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.din(n115));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n117_1(.douta(w_dff_A_yru3O2PL1_0),.doutb(w_n117_1[1]),.din(w_n117_0[0]));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_dff_A_qBWieEza7_1),.doutc(w_dff_A_9gXtwih81_2),.din(n118));
	jspl3 jspl3_w_n118_1(.douta(w_dff_A_p1148UTE1_0),.doutb(w_dff_A_jylKDbSY7_1),.doutc(w_n118_1[2]),.din(w_n118_0[0]));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_dff_A_hRCJFKgL4_1),.din(w_dff_B_UWBylWK54_2));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n133_0(.douta(w_n133_0[0]),.doutb(w_dff_A_NOx3pkQq9_1),.doutc(w_n133_0[2]),.din(n133));
	jspl jspl_w_n133_1(.douta(w_dff_A_UTvZTO7I7_0),.doutb(w_n133_1[1]),.din(w_n133_0[0]));
	jspl3 jspl3_w_n142_0(.douta(w_n142_0[0]),.doutb(w_dff_A_9qXqSa537_1),.doutc(w_n142_0[2]),.din(n142));
	jspl jspl_w_n142_1(.douta(w_n142_1[0]),.doutb(w_n142_1[1]),.din(w_n142_0[0]));
	jspl3 jspl3_w_n150_0(.douta(w_n150_0[0]),.doutb(w_dff_A_CKvDnEw04_1),.doutc(w_n150_0[2]),.din(n150));
	jspl jspl_w_n150_1(.douta(w_n150_1[0]),.doutb(w_n150_1[1]),.din(w_n150_0[0]));
	jspl3 jspl3_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.doutc(w_n156_0[2]),.din(n156));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_dff_A_ET4d4aUP5_2),.din(n164));
	jspl jspl_w_n164_1(.douta(w_dff_A_QRus6GbE7_0),.doutb(w_n164_1[1]),.din(w_n164_0[0]));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_j2oGcDX49_1),.doutc(w_dff_A_43cGsIwN6_2),.din(n165));
	jspl3 jspl3_w_n165_1(.douta(w_dff_A_uw7ucNNN1_0),.doutb(w_dff_A_bKsqmj1W5_1),.doutc(w_n165_1[2]),.din(w_n165_0[0]));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_dff_A_RE71uI073_2),.din(n173));
	jspl jspl_w_n173_1(.douta(w_n173_1[0]),.doutb(w_dff_A_GHrb1CeX8_1),.din(w_n173_0[0]));
	jspl jspl_w_n174_0(.douta(w_dff_A_vdPcnTFX3_0),.doutb(w_n174_0[1]),.din(w_dff_B_r8FJVIJ24_2));
	jspl3 jspl3_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.doutc(w_n176_0[2]),.din(n176));
	jspl jspl_w_n176_1(.douta(w_n176_1[0]),.doutb(w_n176_1[1]),.din(w_n176_0[0]));
	jspl3 jspl3_w_n179_0(.douta(w_dff_A_DxHEB6cJ1_0),.doutb(w_n179_0[1]),.doutc(w_dff_A_CjlEWrLC3_2),.din(n179));
	jspl3 jspl3_w_n179_1(.douta(w_n179_1[0]),.doutb(w_n179_1[1]),.doutc(w_n179_1[2]),.din(w_n179_0[0]));
	jspl3 jspl3_w_n182_0(.douta(w_dff_A_oAScp9vP1_0),.doutb(w_n182_0[1]),.doutc(w_dff_A_yFAt378D6_2),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n185_0(.douta(w_dff_A_TuXQfG4X9_0),.doutb(w_n185_0[1]),.doutc(w_dff_A_OTPAWWJ69_2),.din(n185));
	jspl3 jspl3_w_n185_1(.douta(w_n185_1[0]),.doutb(w_n185_1[1]),.doutc(w_n185_1[2]),.din(w_n185_0[0]));
	jspl3 jspl3_w_n188_0(.douta(w_n188_0[0]),.doutb(w_dff_A_yaIGEDZr2_1),.doutc(w_dff_A_2jSnBeHT6_2),.din(n188));
	jspl3 jspl3_w_n188_1(.douta(w_dff_A_JkHF1v2x3_0),.doutb(w_dff_A_Sge4AOLm8_1),.doutc(w_n188_1[2]),.din(w_n188_0[0]));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n191_1(.douta(w_n191_1[0]),.doutb(w_n191_1[1]),.din(w_n191_0[0]));
	jspl3 jspl3_w_n200_0(.douta(w_n200_0[0]),.doutb(w_dff_A_0ViuaRIr7_1),.doutc(w_dff_A_pQGFEaYd0_2),.din(n200));
	jspl3 jspl3_w_n200_1(.douta(w_dff_A_Yw9zhwJZ6_0),.doutb(w_dff_A_FezvLLFD3_1),.doutc(w_n200_1[2]),.din(w_n200_0[0]));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(w_dff_B_BNLlAz3j6_2));
	jspl3 jspl3_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.doutc(w_n203_0[2]),.din(n203));
	jspl jspl_w_n203_1(.douta(w_n203_1[0]),.doutb(w_n203_1[1]),.din(w_n203_0[0]));
	jspl3 jspl3_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.doutc(w_n212_0[2]),.din(n212));
	jspl jspl_w_n212_1(.douta(w_n212_1[0]),.doutb(w_n212_1[1]),.din(w_n212_0[0]));
	jspl jspl_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.din(w_dff_B_A8fCb3Nv3_2));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.din(n229));
	jspl jspl_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.doutc(w_n231_0[2]),.din(n231));
	jspl jspl_w_n231_1(.douta(w_n231_1[0]),.doutb(w_n231_1[1]),.din(w_n231_0[0]));
	jspl jspl_w_n240_0(.douta(w_n240_0[0]),.doutb(w_n240_0[1]),.din(w_dff_B_E1H7gFcr9_2));
	jspl3 jspl3_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.doutc(w_n241_0[2]),.din(n241));
	jspl jspl_w_n241_1(.douta(w_n241_1[0]),.doutb(w_n241_1[1]),.din(w_n241_0[0]));
	jspl jspl_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.din(n251));
	jspl3 jspl3_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.doutc(w_n252_0[2]),.din(n252));
	jspl jspl_w_n252_1(.douta(w_n252_1[0]),.doutb(w_n252_1[1]),.din(w_n252_0[0]));
	jspl3 jspl3_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.doutc(w_n261_0[2]),.din(n261));
	jspl jspl_w_n261_1(.douta(w_n261_1[0]),.doutb(w_n261_1[1]),.din(w_n261_0[0]));
	jdff dff_A_vdPcnTFX3_0(.dout(w_n174_0[0]),.din(w_dff_A_vdPcnTFX3_0),.clk(gclk));
	jdff dff_B_r8FJVIJ24_2(.din(n174),.dout(w_dff_B_r8FJVIJ24_2),.clk(gclk));
	jdff dff_A_hRCJFKgL4_1(.dout(w_n119_0[1]),.din(w_dff_A_hRCJFKgL4_1),.clk(gclk));
	jdff dff_B_UWBylWK54_2(.din(n119),.dout(w_dff_B_UWBylWK54_2),.clk(gclk));
	jdff dff_B_7Cck4rhx1_2(.din(n201),.dout(w_dff_B_7Cck4rhx1_2),.clk(gclk));
	jdff dff_B_BNLlAz3j6_2(.din(w_dff_B_7Cck4rhx1_2),.dout(w_dff_B_BNLlAz3j6_2),.clk(gclk));
	jdff dff_B_qUrfu9jW1_0(.din(n189),.dout(w_dff_B_qUrfu9jW1_0),.clk(gclk));
	jdff dff_B_owl8iB525_1(.din(n152),.dout(w_dff_B_owl8iB525_1),.clk(gclk));
	jdff dff_A_lGAB4W7I8_0(.dout(w_n133_1[0]),.din(w_dff_A_lGAB4W7I8_0),.clk(gclk));
	jdff dff_A_UTvZTO7I7_0(.dout(w_dff_A_lGAB4W7I8_0),.din(w_dff_A_UTvZTO7I7_0),.clk(gclk));
	jdff dff_A_dpigLNVm3_0(.dout(w_n165_1[0]),.din(w_dff_A_dpigLNVm3_0),.clk(gclk));
	jdff dff_A_qSiySCfX4_0(.dout(w_dff_A_dpigLNVm3_0),.din(w_dff_A_qSiySCfX4_0),.clk(gclk));
	jdff dff_A_gU9C9yEW4_0(.dout(w_dff_A_qSiySCfX4_0),.din(w_dff_A_gU9C9yEW4_0),.clk(gclk));
	jdff dff_A_uw7ucNNN1_0(.dout(w_dff_A_gU9C9yEW4_0),.din(w_dff_A_uw7ucNNN1_0),.clk(gclk));
	jdff dff_A_7Be8AeBF8_1(.dout(w_n165_1[1]),.din(w_dff_A_7Be8AeBF8_1),.clk(gclk));
	jdff dff_A_Ui5HdkiS3_1(.dout(w_dff_A_7Be8AeBF8_1),.din(w_dff_A_Ui5HdkiS3_1),.clk(gclk));
	jdff dff_A_QrBhabZh9_1(.dout(w_dff_A_Ui5HdkiS3_1),.din(w_dff_A_QrBhabZh9_1),.clk(gclk));
	jdff dff_A_bKsqmj1W5_1(.dout(w_dff_A_QrBhabZh9_1),.din(w_dff_A_bKsqmj1W5_1),.clk(gclk));
	jdff dff_A_d6agRoYl7_0(.dout(w_n200_1[0]),.din(w_dff_A_d6agRoYl7_0),.clk(gclk));
	jdff dff_A_NZ7vswYn4_0(.dout(w_dff_A_d6agRoYl7_0),.din(w_dff_A_NZ7vswYn4_0),.clk(gclk));
	jdff dff_A_DTeIsMUa0_0(.dout(w_dff_A_NZ7vswYn4_0),.din(w_dff_A_DTeIsMUa0_0),.clk(gclk));
	jdff dff_A_Yw9zhwJZ6_0(.dout(w_dff_A_DTeIsMUa0_0),.din(w_dff_A_Yw9zhwJZ6_0),.clk(gclk));
	jdff dff_A_Yh9lxLTl9_1(.dout(w_n200_1[1]),.din(w_dff_A_Yh9lxLTl9_1),.clk(gclk));
	jdff dff_A_GaqwIUbM1_1(.dout(w_dff_A_Yh9lxLTl9_1),.din(w_dff_A_GaqwIUbM1_1),.clk(gclk));
	jdff dff_A_iEzGq03t6_1(.dout(w_dff_A_GaqwIUbM1_1),.din(w_dff_A_iEzGq03t6_1),.clk(gclk));
	jdff dff_A_FezvLLFD3_1(.dout(w_dff_A_iEzGq03t6_1),.din(w_dff_A_FezvLLFD3_1),.clk(gclk));
	jdff dff_A_HVymXHBn8_0(.dout(w_n118_1[0]),.din(w_dff_A_HVymXHBn8_0),.clk(gclk));
	jdff dff_A_3jIiPkuY9_0(.dout(w_dff_A_HVymXHBn8_0),.din(w_dff_A_3jIiPkuY9_0),.clk(gclk));
	jdff dff_A_sJw7kvzQ3_0(.dout(w_dff_A_3jIiPkuY9_0),.din(w_dff_A_sJw7kvzQ3_0),.clk(gclk));
	jdff dff_A_p1148UTE1_0(.dout(w_dff_A_sJw7kvzQ3_0),.din(w_dff_A_p1148UTE1_0),.clk(gclk));
	jdff dff_A_OOM77HGc5_1(.dout(w_n118_1[1]),.din(w_dff_A_OOM77HGc5_1),.clk(gclk));
	jdff dff_A_hfqDjlSn7_1(.dout(w_dff_A_OOM77HGc5_1),.din(w_dff_A_hfqDjlSn7_1),.clk(gclk));
	jdff dff_A_XpX6X2mh5_1(.dout(w_dff_A_hfqDjlSn7_1),.din(w_dff_A_XpX6X2mh5_1),.clk(gclk));
	jdff dff_A_jylKDbSY7_1(.dout(w_dff_A_XpX6X2mh5_1),.din(w_dff_A_jylKDbSY7_1),.clk(gclk));
	jdff dff_B_BgaXxk1H8_1(.din(n222),.dout(w_dff_B_BgaXxk1H8_1),.clk(gclk));
	jdff dff_A_TmkUtfMt5_0(.dout(w_n88_0[0]),.din(w_dff_A_TmkUtfMt5_0),.clk(gclk));
	jdff dff_A_2vQDDBMR5_0(.dout(w_dff_A_TmkUtfMt5_0),.din(w_dff_A_2vQDDBMR5_0),.clk(gclk));
	jdff dff_A_K9FeKXkR0_0(.dout(w_dff_A_2vQDDBMR5_0),.din(w_dff_A_K9FeKXkR0_0),.clk(gclk));
	jdff dff_A_cOd908YV2_0(.dout(w_dff_A_K9FeKXkR0_0),.din(w_dff_A_cOd908YV2_0),.clk(gclk));
	jdff dff_A_YygD2thL4_2(.dout(w_n88_0[2]),.din(w_dff_A_YygD2thL4_2),.clk(gclk));
	jdff dff_A_w1kJl7rA1_2(.dout(w_dff_A_YygD2thL4_2),.din(w_dff_A_w1kJl7rA1_2),.clk(gclk));
	jdff dff_A_auMrjeNo8_2(.dout(w_dff_A_w1kJl7rA1_2),.din(w_dff_A_auMrjeNo8_2),.clk(gclk));
	jdff dff_A_DcTjdZYh3_2(.dout(w_dff_A_auMrjeNo8_2),.din(w_dff_A_DcTjdZYh3_2),.clk(gclk));
	jdff dff_A_Inlo5oks1_0(.dout(w_n188_1[0]),.din(w_dff_A_Inlo5oks1_0),.clk(gclk));
	jdff dff_A_qPeFRIWT1_0(.dout(w_dff_A_Inlo5oks1_0),.din(w_dff_A_qPeFRIWT1_0),.clk(gclk));
	jdff dff_A_3Mvle7Tq3_0(.dout(w_dff_A_qPeFRIWT1_0),.din(w_dff_A_3Mvle7Tq3_0),.clk(gclk));
	jdff dff_A_JkHF1v2x3_0(.dout(w_dff_A_3Mvle7Tq3_0),.din(w_dff_A_JkHF1v2x3_0),.clk(gclk));
	jdff dff_A_2VwTkvX12_1(.dout(w_n188_1[1]),.din(w_dff_A_2VwTkvX12_1),.clk(gclk));
	jdff dff_A_0zWqIJsV5_1(.dout(w_dff_A_2VwTkvX12_1),.din(w_dff_A_0zWqIJsV5_1),.clk(gclk));
	jdff dff_A_1jIi0ivv1_1(.dout(w_dff_A_0zWqIJsV5_1),.din(w_dff_A_1jIi0ivv1_1),.clk(gclk));
	jdff dff_A_Sge4AOLm8_1(.dout(w_dff_A_1jIi0ivv1_1),.din(w_dff_A_Sge4AOLm8_1),.clk(gclk));
	jdff dff_B_IehodlcR5_2(.din(n221),.dout(w_dff_B_IehodlcR5_2),.clk(gclk));
	jdff dff_B_A8fCb3Nv3_2(.din(w_dff_B_IehodlcR5_2),.dout(w_dff_B_A8fCb3Nv3_2),.clk(gclk));
	jdff dff_A_0ZLYMpt93_0(.dout(w_n182_0[0]),.din(w_dff_A_0ZLYMpt93_0),.clk(gclk));
	jdff dff_A_qu6ztY5D1_0(.dout(w_dff_A_0ZLYMpt93_0),.din(w_dff_A_qu6ztY5D1_0),.clk(gclk));
	jdff dff_A_flIgCFXO2_0(.dout(w_dff_A_qu6ztY5D1_0),.din(w_dff_A_flIgCFXO2_0),.clk(gclk));
	jdff dff_A_oAScp9vP1_0(.dout(w_dff_A_flIgCFXO2_0),.din(w_dff_A_oAScp9vP1_0),.clk(gclk));
	jdff dff_A_cci19hNq5_2(.dout(w_n182_0[2]),.din(w_dff_A_cci19hNq5_2),.clk(gclk));
	jdff dff_A_3HIlSwSn5_2(.dout(w_dff_A_cci19hNq5_2),.din(w_dff_A_3HIlSwSn5_2),.clk(gclk));
	jdff dff_A_4Ju04hih4_2(.dout(w_dff_A_3HIlSwSn5_2),.din(w_dff_A_4Ju04hih4_2),.clk(gclk));
	jdff dff_A_yFAt378D6_2(.dout(w_dff_A_4Ju04hih4_2),.din(w_dff_A_yFAt378D6_2),.clk(gclk));
	jdff dff_A_c8UqvpQi4_1(.dout(w_n165_0[1]),.din(w_dff_A_c8UqvpQi4_1),.clk(gclk));
	jdff dff_A_Y9q25Hs56_1(.dout(w_dff_A_c8UqvpQi4_1),.din(w_dff_A_Y9q25Hs56_1),.clk(gclk));
	jdff dff_A_5NEjFakf1_1(.dout(w_dff_A_Y9q25Hs56_1),.din(w_dff_A_5NEjFakf1_1),.clk(gclk));
	jdff dff_A_j2oGcDX49_1(.dout(w_dff_A_5NEjFakf1_1),.din(w_dff_A_j2oGcDX49_1),.clk(gclk));
	jdff dff_A_54LPtYOM0_2(.dout(w_n165_0[2]),.din(w_dff_A_54LPtYOM0_2),.clk(gclk));
	jdff dff_A_TBZ1rb6v5_2(.dout(w_dff_A_54LPtYOM0_2),.din(w_dff_A_TBZ1rb6v5_2),.clk(gclk));
	jdff dff_A_0sagchlM8_2(.dout(w_dff_A_TBZ1rb6v5_2),.din(w_dff_A_0sagchlM8_2),.clk(gclk));
	jdff dff_A_43cGsIwN6_2(.dout(w_dff_A_0sagchlM8_2),.din(w_dff_A_43cGsIwN6_2),.clk(gclk));
	jdff dff_A_QRus6GbE7_0(.dout(w_n164_1[0]),.din(w_dff_A_QRus6GbE7_0),.clk(gclk));
	jdff dff_A_HR8rokqC6_1(.dout(w_n200_0[1]),.din(w_dff_A_HR8rokqC6_1),.clk(gclk));
	jdff dff_A_QpLUy2g79_1(.dout(w_dff_A_HR8rokqC6_1),.din(w_dff_A_QpLUy2g79_1),.clk(gclk));
	jdff dff_A_H1abPuNI0_1(.dout(w_dff_A_QpLUy2g79_1),.din(w_dff_A_H1abPuNI0_1),.clk(gclk));
	jdff dff_A_0ViuaRIr7_1(.dout(w_dff_A_H1abPuNI0_1),.din(w_dff_A_0ViuaRIr7_1),.clk(gclk));
	jdff dff_A_PEgZkBLG6_2(.dout(w_n200_0[2]),.din(w_dff_A_PEgZkBLG6_2),.clk(gclk));
	jdff dff_A_EEsZ9AwR2_2(.dout(w_dff_A_PEgZkBLG6_2),.din(w_dff_A_EEsZ9AwR2_2),.clk(gclk));
	jdff dff_A_LzL16HWy4_2(.dout(w_dff_A_EEsZ9AwR2_2),.din(w_dff_A_LzL16HWy4_2),.clk(gclk));
	jdff dff_A_pQGFEaYd0_2(.dout(w_dff_A_LzL16HWy4_2),.din(w_dff_A_pQGFEaYd0_2),.clk(gclk));
	jdff dff_A_GHrb1CeX8_1(.dout(w_n173_1[1]),.din(w_dff_A_GHrb1CeX8_1),.clk(gclk));
	jdff dff_A_HzaJ06GZ9_1(.dout(w_n118_0[1]),.din(w_dff_A_HzaJ06GZ9_1),.clk(gclk));
	jdff dff_A_1AgXO7ki6_1(.dout(w_dff_A_HzaJ06GZ9_1),.din(w_dff_A_1AgXO7ki6_1),.clk(gclk));
	jdff dff_A_aulwWU2G9_1(.dout(w_dff_A_1AgXO7ki6_1),.din(w_dff_A_aulwWU2G9_1),.clk(gclk));
	jdff dff_A_qBWieEza7_1(.dout(w_dff_A_aulwWU2G9_1),.din(w_dff_A_qBWieEza7_1),.clk(gclk));
	jdff dff_A_rjjrpJgt2_2(.dout(w_n118_0[2]),.din(w_dff_A_rjjrpJgt2_2),.clk(gclk));
	jdff dff_A_zc9hvvMt9_2(.dout(w_dff_A_rjjrpJgt2_2),.din(w_dff_A_zc9hvvMt9_2),.clk(gclk));
	jdff dff_A_NEYxA4Vr7_2(.dout(w_dff_A_zc9hvvMt9_2),.din(w_dff_A_NEYxA4Vr7_2),.clk(gclk));
	jdff dff_A_9gXtwih81_2(.dout(w_dff_A_NEYxA4Vr7_2),.din(w_dff_A_9gXtwih81_2),.clk(gclk));
	jdff dff_A_yru3O2PL1_0(.dout(w_n117_1[0]),.din(w_dff_A_yru3O2PL1_0),.clk(gclk));
	jdff dff_B_FOpXhkhO3_1(.din(n250),.dout(w_dff_B_FOpXhkhO3_1),.clk(gclk));
	jdff dff_B_w00ffTJc9_0(.din(n228),.dout(w_dff_B_w00ffTJc9_0),.clk(gclk));
	jdff dff_B_1n0vBH7l2_1(.din(n112),.dout(w_dff_B_1n0vBH7l2_1),.clk(gclk));
	jdff dff_A_ET4d4aUP5_2(.dout(w_n164_0[2]),.din(w_dff_A_ET4d4aUP5_2),.clk(gclk));
	jdff dff_A_RNt34pof7_2(.dout(w_n173_0[2]),.din(w_dff_A_RNt34pof7_2),.clk(gclk));
	jdff dff_A_RE71uI073_2(.dout(w_dff_A_RNt34pof7_2),.din(w_dff_A_RE71uI073_2),.clk(gclk));
	jdff dff_A_z5ik1pbm6_0(.dout(w_n179_0[0]),.din(w_dff_A_z5ik1pbm6_0),.clk(gclk));
	jdff dff_A_JtFH7GZw0_0(.dout(w_dff_A_z5ik1pbm6_0),.din(w_dff_A_JtFH7GZw0_0),.clk(gclk));
	jdff dff_A_hlD9GBci7_0(.dout(w_dff_A_JtFH7GZw0_0),.din(w_dff_A_hlD9GBci7_0),.clk(gclk));
	jdff dff_A_DxHEB6cJ1_0(.dout(w_dff_A_hlD9GBci7_0),.din(w_dff_A_DxHEB6cJ1_0),.clk(gclk));
	jdff dff_A_imgJg5xS1_2(.dout(w_n179_0[2]),.din(w_dff_A_imgJg5xS1_2),.clk(gclk));
	jdff dff_A_v3McqeVC7_2(.dout(w_dff_A_imgJg5xS1_2),.din(w_dff_A_v3McqeVC7_2),.clk(gclk));
	jdff dff_A_KycxdNdu5_2(.dout(w_dff_A_v3McqeVC7_2),.din(w_dff_A_KycxdNdu5_2),.clk(gclk));
	jdff dff_A_CjlEWrLC3_2(.dout(w_dff_A_KycxdNdu5_2),.din(w_dff_A_CjlEWrLC3_2),.clk(gclk));
	jdff dff_A_NOx3pkQq9_1(.dout(w_n133_0[1]),.din(w_dff_A_NOx3pkQq9_1),.clk(gclk));
	jdff dff_A_YhQXZeI68_0(.dout(w_G8gat_0[0]),.din(w_dff_A_YhQXZeI68_0),.clk(gclk));
	jdff dff_A_1iUUqMce3_0(.dout(w_dff_A_YhQXZeI68_0),.din(w_dff_A_1iUUqMce3_0),.clk(gclk));
	jdff dff_A_sulxPjQc9_0(.dout(w_dff_A_1iUUqMce3_0),.din(w_dff_A_sulxPjQc9_0),.clk(gclk));
	jdff dff_A_ZRU7skZH6_0(.dout(w_dff_A_sulxPjQc9_0),.din(w_dff_A_ZRU7skZH6_0),.clk(gclk));
	jdff dff_A_86JC351g8_0(.dout(w_dff_A_ZRU7skZH6_0),.din(w_dff_A_86JC351g8_0),.clk(gclk));
	jdff dff_A_jQ4qLKjT1_0(.dout(w_dff_A_86JC351g8_0),.din(w_dff_A_jQ4qLKjT1_0),.clk(gclk));
	jdff dff_A_qi7AQSsh8_0(.dout(w_dff_A_jQ4qLKjT1_0),.din(w_dff_A_qi7AQSsh8_0),.clk(gclk));
	jdff dff_A_I6dWuaU49_0(.dout(w_dff_A_qi7AQSsh8_0),.din(w_dff_A_I6dWuaU49_0),.clk(gclk));
	jdff dff_A_MtHr3Kaq5_0(.dout(w_dff_A_I6dWuaU49_0),.din(w_dff_A_MtHr3Kaq5_0),.clk(gclk));
	jdff dff_A_RnARyNcU7_0(.dout(w_dff_A_MtHr3Kaq5_0),.din(w_dff_A_RnARyNcU7_0),.clk(gclk));
	jdff dff_A_ZySGaYA15_0(.dout(w_G64gat_0[0]),.din(w_dff_A_ZySGaYA15_0),.clk(gclk));
	jdff dff_A_d9WF0F7t5_0(.dout(w_dff_A_ZySGaYA15_0),.din(w_dff_A_d9WF0F7t5_0),.clk(gclk));
	jdff dff_A_0CGjDb7w0_0(.dout(w_dff_A_d9WF0F7t5_0),.din(w_dff_A_0CGjDb7w0_0),.clk(gclk));
	jdff dff_A_0IJJrDDU9_0(.dout(w_dff_A_0CGjDb7w0_0),.din(w_dff_A_0IJJrDDU9_0),.clk(gclk));
	jdff dff_A_efdEqy2z8_0(.dout(w_dff_A_0IJJrDDU9_0),.din(w_dff_A_efdEqy2z8_0),.clk(gclk));
	jdff dff_A_zBCtljCk0_0(.dout(w_dff_A_efdEqy2z8_0),.din(w_dff_A_zBCtljCk0_0),.clk(gclk));
	jdff dff_A_q2raEr044_0(.dout(w_dff_A_zBCtljCk0_0),.din(w_dff_A_q2raEr044_0),.clk(gclk));
	jdff dff_A_VMvjioiq2_0(.dout(w_dff_A_q2raEr044_0),.din(w_dff_A_VMvjioiq2_0),.clk(gclk));
	jdff dff_A_n7wLgPXX5_0(.dout(w_dff_A_VMvjioiq2_0),.din(w_dff_A_n7wLgPXX5_0),.clk(gclk));
	jdff dff_A_6ofuZSxw0_0(.dout(w_dff_A_n7wLgPXX5_0),.din(w_dff_A_6ofuZSxw0_0),.clk(gclk));
	jdff dff_A_5SFFyfvI3_1(.dout(w_n87_0[1]),.din(w_dff_A_5SFFyfvI3_1),.clk(gclk));
	jdff dff_A_BfXk90y80_2(.dout(w_n87_0[2]),.din(w_dff_A_BfXk90y80_2),.clk(gclk));
	jdff dff_A_bedMVhhi9_0(.dout(w_G1gat_0[0]),.din(w_dff_A_bedMVhhi9_0),.clk(gclk));
	jdff dff_A_N0P3wn1K3_0(.dout(w_dff_A_bedMVhhi9_0),.din(w_dff_A_N0P3wn1K3_0),.clk(gclk));
	jdff dff_A_OFLk40Xe9_0(.dout(w_dff_A_N0P3wn1K3_0),.din(w_dff_A_OFLk40Xe9_0),.clk(gclk));
	jdff dff_A_GSWiFwCq8_0(.dout(w_dff_A_OFLk40Xe9_0),.din(w_dff_A_GSWiFwCq8_0),.clk(gclk));
	jdff dff_A_SDCfabFB9_0(.dout(w_dff_A_GSWiFwCq8_0),.din(w_dff_A_SDCfabFB9_0),.clk(gclk));
	jdff dff_A_KXgaq1yM2_0(.dout(w_dff_A_SDCfabFB9_0),.din(w_dff_A_KXgaq1yM2_0),.clk(gclk));
	jdff dff_A_LK6DEAa72_0(.dout(w_dff_A_KXgaq1yM2_0),.din(w_dff_A_LK6DEAa72_0),.clk(gclk));
	jdff dff_A_C9oQZRvw3_0(.dout(w_dff_A_LK6DEAa72_0),.din(w_dff_A_C9oQZRvw3_0),.clk(gclk));
	jdff dff_A_WEFQwI8F3_0(.dout(w_dff_A_C9oQZRvw3_0),.din(w_dff_A_WEFQwI8F3_0),.clk(gclk));
	jdff dff_A_eodqpG4e5_0(.dout(w_dff_A_WEFQwI8F3_0),.din(w_dff_A_eodqpG4e5_0),.clk(gclk));
	jdff dff_A_ktA7mwbm7_0(.dout(w_G57gat_0[0]),.din(w_dff_A_ktA7mwbm7_0),.clk(gclk));
	jdff dff_A_5DkprJcj8_0(.dout(w_dff_A_ktA7mwbm7_0),.din(w_dff_A_5DkprJcj8_0),.clk(gclk));
	jdff dff_A_9lv3Amie2_0(.dout(w_dff_A_5DkprJcj8_0),.din(w_dff_A_9lv3Amie2_0),.clk(gclk));
	jdff dff_A_tuJ8xmcg2_0(.dout(w_dff_A_9lv3Amie2_0),.din(w_dff_A_tuJ8xmcg2_0),.clk(gclk));
	jdff dff_A_BLnz5Epy3_0(.dout(w_dff_A_tuJ8xmcg2_0),.din(w_dff_A_BLnz5Epy3_0),.clk(gclk));
	jdff dff_A_IssG3zlj8_0(.dout(w_dff_A_BLnz5Epy3_0),.din(w_dff_A_IssG3zlj8_0),.clk(gclk));
	jdff dff_A_Jnsshwon5_0(.dout(w_dff_A_IssG3zlj8_0),.din(w_dff_A_Jnsshwon5_0),.clk(gclk));
	jdff dff_A_2m3yCjbj1_0(.dout(w_dff_A_Jnsshwon5_0),.din(w_dff_A_2m3yCjbj1_0),.clk(gclk));
	jdff dff_A_ApktT6vx1_0(.dout(w_dff_A_2m3yCjbj1_0),.din(w_dff_A_ApktT6vx1_0),.clk(gclk));
	jdff dff_A_q7DjgNRJ8_0(.dout(w_dff_A_ApktT6vx1_0),.din(w_dff_A_q7DjgNRJ8_0),.clk(gclk));
	jdff dff_B_9LmMrDv48_2(.din(n240),.dout(w_dff_B_9LmMrDv48_2),.clk(gclk));
	jdff dff_B_E1H7gFcr9_2(.din(w_dff_B_9LmMrDv48_2),.dout(w_dff_B_E1H7gFcr9_2),.clk(gclk));
	jdff dff_A_B6URFRbq9_0(.dout(w_n185_0[0]),.din(w_dff_A_B6URFRbq9_0),.clk(gclk));
	jdff dff_A_NddPX5cX2_0(.dout(w_dff_A_B6URFRbq9_0),.din(w_dff_A_NddPX5cX2_0),.clk(gclk));
	jdff dff_A_ABv4K3DA1_0(.dout(w_dff_A_NddPX5cX2_0),.din(w_dff_A_ABv4K3DA1_0),.clk(gclk));
	jdff dff_A_TuXQfG4X9_0(.dout(w_dff_A_ABv4K3DA1_0),.din(w_dff_A_TuXQfG4X9_0),.clk(gclk));
	jdff dff_A_8dVzED9r0_2(.dout(w_n185_0[2]),.din(w_dff_A_8dVzED9r0_2),.clk(gclk));
	jdff dff_A_KlEUMlVr0_2(.dout(w_dff_A_8dVzED9r0_2),.din(w_dff_A_KlEUMlVr0_2),.clk(gclk));
	jdff dff_A_dum3mdWz3_2(.dout(w_dff_A_KlEUMlVr0_2),.din(w_dff_A_dum3mdWz3_2),.clk(gclk));
	jdff dff_A_OTPAWWJ69_2(.dout(w_dff_A_dum3mdWz3_2),.din(w_dff_A_OTPAWWJ69_2),.clk(gclk));
	jdff dff_A_CKvDnEw04_1(.dout(w_n150_0[1]),.din(w_dff_A_CKvDnEw04_1),.clk(gclk));
	jdff dff_B_q9oyvLJJ6_0(.din(n148),.dout(w_dff_B_q9oyvLJJ6_0),.clk(gclk));
	jdff dff_A_lOLlEOb58_0(.dout(w_G148gat_0[0]),.din(w_dff_A_lOLlEOb58_0),.clk(gclk));
	jdff dff_A_mM24LcMB6_0(.dout(w_dff_A_lOLlEOb58_0),.din(w_dff_A_mM24LcMB6_0),.clk(gclk));
	jdff dff_A_6vkJHhZs1_0(.dout(w_dff_A_mM24LcMB6_0),.din(w_dff_A_6vkJHhZs1_0),.clk(gclk));
	jdff dff_A_cwU9WSZM9_0(.dout(w_dff_A_6vkJHhZs1_0),.din(w_dff_A_cwU9WSZM9_0),.clk(gclk));
	jdff dff_A_uK3IhWNC8_0(.dout(w_dff_A_cwU9WSZM9_0),.din(w_dff_A_uK3IhWNC8_0),.clk(gclk));
	jdff dff_A_nOG9BSCP4_0(.dout(w_dff_A_uK3IhWNC8_0),.din(w_dff_A_nOG9BSCP4_0),.clk(gclk));
	jdff dff_A_Y5lBGqJ05_0(.dout(w_dff_A_nOG9BSCP4_0),.din(w_dff_A_Y5lBGqJ05_0),.clk(gclk));
	jdff dff_A_VIJiJCyq6_0(.dout(w_dff_A_Y5lBGqJ05_0),.din(w_dff_A_VIJiJCyq6_0),.clk(gclk));
	jdff dff_A_xrVHGazt6_0(.dout(w_dff_A_VIJiJCyq6_0),.din(w_dff_A_xrVHGazt6_0),.clk(gclk));
	jdff dff_A_IH5t9iYx6_0(.dout(w_dff_A_xrVHGazt6_0),.din(w_dff_A_IH5t9iYx6_0),.clk(gclk));
	jdff dff_A_UGnvSxT39_0(.dout(w_G141gat_0[0]),.din(w_dff_A_UGnvSxT39_0),.clk(gclk));
	jdff dff_A_xpi9CXyb3_0(.dout(w_dff_A_UGnvSxT39_0),.din(w_dff_A_xpi9CXyb3_0),.clk(gclk));
	jdff dff_A_frFC1J7Q2_0(.dout(w_dff_A_xpi9CXyb3_0),.din(w_dff_A_frFC1J7Q2_0),.clk(gclk));
	jdff dff_A_fJuxviOY2_0(.dout(w_dff_A_frFC1J7Q2_0),.din(w_dff_A_fJuxviOY2_0),.clk(gclk));
	jdff dff_A_47to3FvV1_0(.dout(w_dff_A_fJuxviOY2_0),.din(w_dff_A_47to3FvV1_0),.clk(gclk));
	jdff dff_A_OircruCZ0_0(.dout(w_dff_A_47to3FvV1_0),.din(w_dff_A_OircruCZ0_0),.clk(gclk));
	jdff dff_A_6WLlouUT9_0(.dout(w_dff_A_OircruCZ0_0),.din(w_dff_A_6WLlouUT9_0),.clk(gclk));
	jdff dff_A_RpfDDlFo6_0(.dout(w_dff_A_6WLlouUT9_0),.din(w_dff_A_RpfDDlFo6_0),.clk(gclk));
	jdff dff_A_VHaVAnIW9_0(.dout(w_dff_A_RpfDDlFo6_0),.din(w_dff_A_VHaVAnIW9_0),.clk(gclk));
	jdff dff_A_gHSCOu0H3_0(.dout(w_dff_A_VHaVAnIW9_0),.din(w_dff_A_gHSCOu0H3_0),.clk(gclk));
	jdff dff_A_xE6xDtaC4_0(.dout(w_G155gat_0[0]),.din(w_dff_A_xE6xDtaC4_0),.clk(gclk));
	jdff dff_A_J5WdBcqk6_0(.dout(w_dff_A_xE6xDtaC4_0),.din(w_dff_A_J5WdBcqk6_0),.clk(gclk));
	jdff dff_A_lnajIqec4_0(.dout(w_dff_A_J5WdBcqk6_0),.din(w_dff_A_lnajIqec4_0),.clk(gclk));
	jdff dff_A_sf4y9oYY9_0(.dout(w_dff_A_lnajIqec4_0),.din(w_dff_A_sf4y9oYY9_0),.clk(gclk));
	jdff dff_A_VhGPRo4X9_0(.dout(w_dff_A_sf4y9oYY9_0),.din(w_dff_A_VhGPRo4X9_0),.clk(gclk));
	jdff dff_A_tF6ERLtR4_0(.dout(w_dff_A_VhGPRo4X9_0),.din(w_dff_A_tF6ERLtR4_0),.clk(gclk));
	jdff dff_A_YYzIuxGT1_0(.dout(w_dff_A_tF6ERLtR4_0),.din(w_dff_A_YYzIuxGT1_0),.clk(gclk));
	jdff dff_A_bq72miS85_0(.dout(w_dff_A_YYzIuxGT1_0),.din(w_dff_A_bq72miS85_0),.clk(gclk));
	jdff dff_A_WWjmO0TC2_0(.dout(w_dff_A_bq72miS85_0),.din(w_dff_A_WWjmO0TC2_0),.clk(gclk));
	jdff dff_A_A1pMQ3Hm9_0(.dout(w_dff_A_WWjmO0TC2_0),.din(w_dff_A_A1pMQ3Hm9_0),.clk(gclk));
	jdff dff_A_p7USBnxT4_0(.dout(w_G22gat_0[0]),.din(w_dff_A_p7USBnxT4_0),.clk(gclk));
	jdff dff_A_UapwwjJo4_0(.dout(w_dff_A_p7USBnxT4_0),.din(w_dff_A_UapwwjJo4_0),.clk(gclk));
	jdff dff_A_B0ewAVea1_0(.dout(w_dff_A_UapwwjJo4_0),.din(w_dff_A_B0ewAVea1_0),.clk(gclk));
	jdff dff_A_JaToxVeE5_0(.dout(w_dff_A_B0ewAVea1_0),.din(w_dff_A_JaToxVeE5_0),.clk(gclk));
	jdff dff_A_9DIBqpjA1_0(.dout(w_dff_A_JaToxVeE5_0),.din(w_dff_A_9DIBqpjA1_0),.clk(gclk));
	jdff dff_A_R3jQqNUW5_0(.dout(w_dff_A_9DIBqpjA1_0),.din(w_dff_A_R3jQqNUW5_0),.clk(gclk));
	jdff dff_A_oLRS4jul9_0(.dout(w_dff_A_R3jQqNUW5_0),.din(w_dff_A_oLRS4jul9_0),.clk(gclk));
	jdff dff_A_Zd8H5dRg1_0(.dout(w_dff_A_oLRS4jul9_0),.din(w_dff_A_Zd8H5dRg1_0),.clk(gclk));
	jdff dff_A_j66GuRiM8_0(.dout(w_dff_A_Zd8H5dRg1_0),.din(w_dff_A_j66GuRiM8_0),.clk(gclk));
	jdff dff_A_W3c8usBA7_0(.dout(w_dff_A_j66GuRiM8_0),.din(w_dff_A_W3c8usBA7_0),.clk(gclk));
	jdff dff_A_9nyimzTq6_0(.dout(w_G78gat_0[0]),.din(w_dff_A_9nyimzTq6_0),.clk(gclk));
	jdff dff_A_vtR8LFjb2_0(.dout(w_dff_A_9nyimzTq6_0),.din(w_dff_A_vtR8LFjb2_0),.clk(gclk));
	jdff dff_A_NHUrFMKO0_0(.dout(w_dff_A_vtR8LFjb2_0),.din(w_dff_A_NHUrFMKO0_0),.clk(gclk));
	jdff dff_A_S7GBDa9p6_0(.dout(w_dff_A_NHUrFMKO0_0),.din(w_dff_A_S7GBDa9p6_0),.clk(gclk));
	jdff dff_A_GcX1QMaQ6_0(.dout(w_dff_A_S7GBDa9p6_0),.din(w_dff_A_GcX1QMaQ6_0),.clk(gclk));
	jdff dff_A_ct0PvfPt1_0(.dout(w_dff_A_GcX1QMaQ6_0),.din(w_dff_A_ct0PvfPt1_0),.clk(gclk));
	jdff dff_A_PFr7EWCL5_0(.dout(w_dff_A_ct0PvfPt1_0),.din(w_dff_A_PFr7EWCL5_0),.clk(gclk));
	jdff dff_A_80VcY0VA5_0(.dout(w_dff_A_PFr7EWCL5_0),.din(w_dff_A_80VcY0VA5_0),.clk(gclk));
	jdff dff_A_AbDVtYd55_0(.dout(w_dff_A_80VcY0VA5_0),.din(w_dff_A_AbDVtYd55_0),.clk(gclk));
	jdff dff_A_aihb3rzW4_0(.dout(w_dff_A_AbDVtYd55_0),.din(w_dff_A_aihb3rzW4_0),.clk(gclk));
	jdff dff_A_JHNkrrkt6_0(.dout(w_G204gat_0[0]),.din(w_dff_A_JHNkrrkt6_0),.clk(gclk));
	jdff dff_A_EffmJLfU4_0(.dout(w_dff_A_JHNkrrkt6_0),.din(w_dff_A_EffmJLfU4_0),.clk(gclk));
	jdff dff_A_L6XCZfzh4_0(.dout(w_dff_A_EffmJLfU4_0),.din(w_dff_A_L6XCZfzh4_0),.clk(gclk));
	jdff dff_A_0XEFr1mJ0_0(.dout(w_dff_A_L6XCZfzh4_0),.din(w_dff_A_0XEFr1mJ0_0),.clk(gclk));
	jdff dff_A_ZDWXEuLp0_0(.dout(w_dff_A_0XEFr1mJ0_0),.din(w_dff_A_ZDWXEuLp0_0),.clk(gclk));
	jdff dff_A_wJBJlFIN9_0(.dout(w_dff_A_ZDWXEuLp0_0),.din(w_dff_A_wJBJlFIN9_0),.clk(gclk));
	jdff dff_A_fyAQG2qW5_0(.dout(w_dff_A_wJBJlFIN9_0),.din(w_dff_A_fyAQG2qW5_0),.clk(gclk));
	jdff dff_A_U61K6byg2_0(.dout(w_dff_A_fyAQG2qW5_0),.din(w_dff_A_U61K6byg2_0),.clk(gclk));
	jdff dff_A_bby7G3um4_0(.dout(w_dff_A_U61K6byg2_0),.din(w_dff_A_bby7G3um4_0),.clk(gclk));
	jdff dff_A_lp3Apxky4_0(.dout(w_dff_A_bby7G3um4_0),.din(w_dff_A_lp3Apxky4_0),.clk(gclk));
	jdff dff_A_gP1fpRqZ8_0(.dout(w_G197gat_0[0]),.din(w_dff_A_gP1fpRqZ8_0),.clk(gclk));
	jdff dff_A_LlpRzyEu7_0(.dout(w_dff_A_gP1fpRqZ8_0),.din(w_dff_A_LlpRzyEu7_0),.clk(gclk));
	jdff dff_A_Ju18mdtB7_0(.dout(w_dff_A_LlpRzyEu7_0),.din(w_dff_A_Ju18mdtB7_0),.clk(gclk));
	jdff dff_A_jKuVhO7H9_0(.dout(w_dff_A_Ju18mdtB7_0),.din(w_dff_A_jKuVhO7H9_0),.clk(gclk));
	jdff dff_A_RFGsi2yE6_0(.dout(w_dff_A_jKuVhO7H9_0),.din(w_dff_A_RFGsi2yE6_0),.clk(gclk));
	jdff dff_A_yVntB7KN0_0(.dout(w_dff_A_RFGsi2yE6_0),.din(w_dff_A_yVntB7KN0_0),.clk(gclk));
	jdff dff_A_AJQpFf6c2_0(.dout(w_dff_A_yVntB7KN0_0),.din(w_dff_A_AJQpFf6c2_0),.clk(gclk));
	jdff dff_A_7Ebkt2Cy9_0(.dout(w_dff_A_AJQpFf6c2_0),.din(w_dff_A_7Ebkt2Cy9_0),.clk(gclk));
	jdff dff_A_g0UO8wW58_0(.dout(w_dff_A_7Ebkt2Cy9_0),.din(w_dff_A_g0UO8wW58_0),.clk(gclk));
	jdff dff_A_QGzJNjho4_0(.dout(w_dff_A_g0UO8wW58_0),.din(w_dff_A_QGzJNjho4_0),.clk(gclk));
	jdff dff_A_FoARUN5b2_0(.dout(w_G211gat_0[0]),.din(w_dff_A_FoARUN5b2_0),.clk(gclk));
	jdff dff_A_Ij0lj3FY2_0(.dout(w_dff_A_FoARUN5b2_0),.din(w_dff_A_Ij0lj3FY2_0),.clk(gclk));
	jdff dff_A_uXUcPjyI4_0(.dout(w_dff_A_Ij0lj3FY2_0),.din(w_dff_A_uXUcPjyI4_0),.clk(gclk));
	jdff dff_A_NOZUmB3r9_0(.dout(w_dff_A_uXUcPjyI4_0),.din(w_dff_A_NOZUmB3r9_0),.clk(gclk));
	jdff dff_A_unqp0OXJ2_0(.dout(w_dff_A_NOZUmB3r9_0),.din(w_dff_A_unqp0OXJ2_0),.clk(gclk));
	jdff dff_A_LyHyXneI0_0(.dout(w_dff_A_unqp0OXJ2_0),.din(w_dff_A_LyHyXneI0_0),.clk(gclk));
	jdff dff_A_vVsZFM9R9_0(.dout(w_dff_A_LyHyXneI0_0),.din(w_dff_A_vVsZFM9R9_0),.clk(gclk));
	jdff dff_A_mdjorY9t5_0(.dout(w_dff_A_vVsZFM9R9_0),.din(w_dff_A_mdjorY9t5_0),.clk(gclk));
	jdff dff_A_Nm8hYCEe7_0(.dout(w_dff_A_mdjorY9t5_0),.din(w_dff_A_Nm8hYCEe7_0),.clk(gclk));
	jdff dff_A_16R7wHZT0_0(.dout(w_dff_A_Nm8hYCEe7_0),.din(w_dff_A_16R7wHZT0_0),.clk(gclk));
	jdff dff_A_9qXqSa537_1(.dout(w_n142_0[1]),.din(w_dff_A_9qXqSa537_1),.clk(gclk));
	jdff dff_B_NbjDkQI86_0(.din(n140),.dout(w_dff_B_NbjDkQI86_0),.clk(gclk));
	jdff dff_A_KiFH5kca6_0(.dout(w_G120gat_0[0]),.din(w_dff_A_KiFH5kca6_0),.clk(gclk));
	jdff dff_A_WXZVXrH93_0(.dout(w_dff_A_KiFH5kca6_0),.din(w_dff_A_WXZVXrH93_0),.clk(gclk));
	jdff dff_A_WcAG9DI67_0(.dout(w_dff_A_WXZVXrH93_0),.din(w_dff_A_WcAG9DI67_0),.clk(gclk));
	jdff dff_A_mg8rkEyR8_0(.dout(w_dff_A_WcAG9DI67_0),.din(w_dff_A_mg8rkEyR8_0),.clk(gclk));
	jdff dff_A_TNOiG2DB9_0(.dout(w_dff_A_mg8rkEyR8_0),.din(w_dff_A_TNOiG2DB9_0),.clk(gclk));
	jdff dff_A_U71FEFkk9_0(.dout(w_dff_A_TNOiG2DB9_0),.din(w_dff_A_U71FEFkk9_0),.clk(gclk));
	jdff dff_A_kYSyubT59_0(.dout(w_dff_A_U71FEFkk9_0),.din(w_dff_A_kYSyubT59_0),.clk(gclk));
	jdff dff_A_wIbPCJM10_0(.dout(w_dff_A_kYSyubT59_0),.din(w_dff_A_wIbPCJM10_0),.clk(gclk));
	jdff dff_A_4bjXMHAC1_0(.dout(w_dff_A_wIbPCJM10_0),.din(w_dff_A_4bjXMHAC1_0),.clk(gclk));
	jdff dff_A_888GxPFd1_0(.dout(w_dff_A_4bjXMHAC1_0),.din(w_dff_A_888GxPFd1_0),.clk(gclk));
	jdff dff_A_EAvaAVwd9_0(.dout(w_G113gat_0[0]),.din(w_dff_A_EAvaAVwd9_0),.clk(gclk));
	jdff dff_A_Y83I1f5Q7_0(.dout(w_dff_A_EAvaAVwd9_0),.din(w_dff_A_Y83I1f5Q7_0),.clk(gclk));
	jdff dff_A_tDnMmOMw2_0(.dout(w_dff_A_Y83I1f5Q7_0),.din(w_dff_A_tDnMmOMw2_0),.clk(gclk));
	jdff dff_A_f43pz4dJ4_0(.dout(w_dff_A_tDnMmOMw2_0),.din(w_dff_A_f43pz4dJ4_0),.clk(gclk));
	jdff dff_A_ZBiGlx7o4_0(.dout(w_dff_A_f43pz4dJ4_0),.din(w_dff_A_ZBiGlx7o4_0),.clk(gclk));
	jdff dff_A_z6Pxcvfe2_0(.dout(w_dff_A_ZBiGlx7o4_0),.din(w_dff_A_z6Pxcvfe2_0),.clk(gclk));
	jdff dff_A_Un8zDzAg9_0(.dout(w_dff_A_z6Pxcvfe2_0),.din(w_dff_A_Un8zDzAg9_0),.clk(gclk));
	jdff dff_A_XbydEyyt1_0(.dout(w_dff_A_Un8zDzAg9_0),.din(w_dff_A_XbydEyyt1_0),.clk(gclk));
	jdff dff_A_wKgpVQdz7_0(.dout(w_dff_A_XbydEyyt1_0),.din(w_dff_A_wKgpVQdz7_0),.clk(gclk));
	jdff dff_A_UeBD4cLQ8_0(.dout(w_dff_A_wKgpVQdz7_0),.din(w_dff_A_UeBD4cLQ8_0),.clk(gclk));
	jdff dff_A_lNzLxEo71_0(.dout(w_G127gat_0[0]),.din(w_dff_A_lNzLxEo71_0),.clk(gclk));
	jdff dff_A_21Nq3TIT9_0(.dout(w_dff_A_lNzLxEo71_0),.din(w_dff_A_21Nq3TIT9_0),.clk(gclk));
	jdff dff_A_bKM8lDHK4_0(.dout(w_dff_A_21Nq3TIT9_0),.din(w_dff_A_bKM8lDHK4_0),.clk(gclk));
	jdff dff_A_nZ63Rjea4_0(.dout(w_dff_A_bKM8lDHK4_0),.din(w_dff_A_nZ63Rjea4_0),.clk(gclk));
	jdff dff_A_ocj7L1Z45_0(.dout(w_dff_A_nZ63Rjea4_0),.din(w_dff_A_ocj7L1Z45_0),.clk(gclk));
	jdff dff_A_YO9xdqZR3_0(.dout(w_dff_A_ocj7L1Z45_0),.din(w_dff_A_YO9xdqZR3_0),.clk(gclk));
	jdff dff_A_nkADfmy61_0(.dout(w_dff_A_YO9xdqZR3_0),.din(w_dff_A_nkADfmy61_0),.clk(gclk));
	jdff dff_A_2CLsx5uI0_0(.dout(w_dff_A_nkADfmy61_0),.din(w_dff_A_2CLsx5uI0_0),.clk(gclk));
	jdff dff_A_QXrEgSM40_0(.dout(w_dff_A_2CLsx5uI0_0),.din(w_dff_A_QXrEgSM40_0),.clk(gclk));
	jdff dff_A_QOW4o5NL8_0(.dout(w_dff_A_QXrEgSM40_0),.din(w_dff_A_QOW4o5NL8_0),.clk(gclk));
	jdff dff_A_9UWkVhLH5_0(.dout(w_G15gat_0[0]),.din(w_dff_A_9UWkVhLH5_0),.clk(gclk));
	jdff dff_A_ayISePTn6_0(.dout(w_dff_A_9UWkVhLH5_0),.din(w_dff_A_ayISePTn6_0),.clk(gclk));
	jdff dff_A_OZi5rbvL0_0(.dout(w_dff_A_ayISePTn6_0),.din(w_dff_A_OZi5rbvL0_0),.clk(gclk));
	jdff dff_A_QQojFK2U1_0(.dout(w_dff_A_OZi5rbvL0_0),.din(w_dff_A_QQojFK2U1_0),.clk(gclk));
	jdff dff_A_M1uRzLfT9_0(.dout(w_dff_A_QQojFK2U1_0),.din(w_dff_A_M1uRzLfT9_0),.clk(gclk));
	jdff dff_A_Q3zomeuh1_0(.dout(w_dff_A_M1uRzLfT9_0),.din(w_dff_A_Q3zomeuh1_0),.clk(gclk));
	jdff dff_A_emCous512_0(.dout(w_dff_A_Q3zomeuh1_0),.din(w_dff_A_emCous512_0),.clk(gclk));
	jdff dff_A_T9HaHUw18_0(.dout(w_dff_A_emCous512_0),.din(w_dff_A_T9HaHUw18_0),.clk(gclk));
	jdff dff_A_zfRI8mNA3_0(.dout(w_dff_A_T9HaHUw18_0),.din(w_dff_A_zfRI8mNA3_0),.clk(gclk));
	jdff dff_A_62ez2TRR5_0(.dout(w_dff_A_zfRI8mNA3_0),.din(w_dff_A_62ez2TRR5_0),.clk(gclk));
	jdff dff_A_4OA0Gfg71_0(.dout(w_G71gat_0[0]),.din(w_dff_A_4OA0Gfg71_0),.clk(gclk));
	jdff dff_A_hVfAd7SZ0_0(.dout(w_dff_A_4OA0Gfg71_0),.din(w_dff_A_hVfAd7SZ0_0),.clk(gclk));
	jdff dff_A_fj8u79Wu6_0(.dout(w_dff_A_hVfAd7SZ0_0),.din(w_dff_A_fj8u79Wu6_0),.clk(gclk));
	jdff dff_A_iq55yZHa1_0(.dout(w_dff_A_fj8u79Wu6_0),.din(w_dff_A_iq55yZHa1_0),.clk(gclk));
	jdff dff_A_tbexwx929_0(.dout(w_dff_A_iq55yZHa1_0),.din(w_dff_A_tbexwx929_0),.clk(gclk));
	jdff dff_A_I1gdxe1m7_0(.dout(w_dff_A_tbexwx929_0),.din(w_dff_A_I1gdxe1m7_0),.clk(gclk));
	jdff dff_A_1LiiKV618_0(.dout(w_dff_A_I1gdxe1m7_0),.din(w_dff_A_1LiiKV618_0),.clk(gclk));
	jdff dff_A_dihKoGgo0_0(.dout(w_dff_A_1LiiKV618_0),.din(w_dff_A_dihKoGgo0_0),.clk(gclk));
	jdff dff_A_ILkwBy1f5_0(.dout(w_dff_A_dihKoGgo0_0),.din(w_dff_A_ILkwBy1f5_0),.clk(gclk));
	jdff dff_A_TMb2lijH8_0(.dout(w_dff_A_ILkwBy1f5_0),.din(w_dff_A_TMb2lijH8_0),.clk(gclk));
	jdff dff_A_CTXvQAYN3_0(.dout(w_G176gat_0[0]),.din(w_dff_A_CTXvQAYN3_0),.clk(gclk));
	jdff dff_A_7OBGOj2w8_0(.dout(w_dff_A_CTXvQAYN3_0),.din(w_dff_A_7OBGOj2w8_0),.clk(gclk));
	jdff dff_A_hni43xyM4_0(.dout(w_dff_A_7OBGOj2w8_0),.din(w_dff_A_hni43xyM4_0),.clk(gclk));
	jdff dff_A_VwyN0akb0_0(.dout(w_dff_A_hni43xyM4_0),.din(w_dff_A_VwyN0akb0_0),.clk(gclk));
	jdff dff_A_AVSdgegI6_0(.dout(w_dff_A_VwyN0akb0_0),.din(w_dff_A_AVSdgegI6_0),.clk(gclk));
	jdff dff_A_52PZheCw3_0(.dout(w_dff_A_AVSdgegI6_0),.din(w_dff_A_52PZheCw3_0),.clk(gclk));
	jdff dff_A_8J6VeEuK7_0(.dout(w_dff_A_52PZheCw3_0),.din(w_dff_A_8J6VeEuK7_0),.clk(gclk));
	jdff dff_A_V6g4VQdq1_0(.dout(w_dff_A_8J6VeEuK7_0),.din(w_dff_A_V6g4VQdq1_0),.clk(gclk));
	jdff dff_A_E0BAUg2T6_0(.dout(w_dff_A_V6g4VQdq1_0),.din(w_dff_A_E0BAUg2T6_0),.clk(gclk));
	jdff dff_A_8JaEixeq4_0(.dout(w_dff_A_E0BAUg2T6_0),.din(w_dff_A_8JaEixeq4_0),.clk(gclk));
	jdff dff_A_WCYXH9172_0(.dout(w_G169gat_0[0]),.din(w_dff_A_WCYXH9172_0),.clk(gclk));
	jdff dff_A_tuEIIjdG2_0(.dout(w_dff_A_WCYXH9172_0),.din(w_dff_A_tuEIIjdG2_0),.clk(gclk));
	jdff dff_A_DiQ4yvs05_0(.dout(w_dff_A_tuEIIjdG2_0),.din(w_dff_A_DiQ4yvs05_0),.clk(gclk));
	jdff dff_A_6394ptkw4_0(.dout(w_dff_A_DiQ4yvs05_0),.din(w_dff_A_6394ptkw4_0),.clk(gclk));
	jdff dff_A_hs4t52pc0_0(.dout(w_dff_A_6394ptkw4_0),.din(w_dff_A_hs4t52pc0_0),.clk(gclk));
	jdff dff_A_GZX8HBgJ8_0(.dout(w_dff_A_hs4t52pc0_0),.din(w_dff_A_GZX8HBgJ8_0),.clk(gclk));
	jdff dff_A_Pai67DP20_0(.dout(w_dff_A_GZX8HBgJ8_0),.din(w_dff_A_Pai67DP20_0),.clk(gclk));
	jdff dff_A_UIW96QiQ1_0(.dout(w_dff_A_Pai67DP20_0),.din(w_dff_A_UIW96QiQ1_0),.clk(gclk));
	jdff dff_A_xcG2OLcu9_0(.dout(w_dff_A_UIW96QiQ1_0),.din(w_dff_A_xcG2OLcu9_0),.clk(gclk));
	jdff dff_A_wQEy2KyV0_0(.dout(w_dff_A_xcG2OLcu9_0),.din(w_dff_A_wQEy2KyV0_0),.clk(gclk));
	jdff dff_A_5nYDEzEt4_0(.dout(w_G183gat_0[0]),.din(w_dff_A_5nYDEzEt4_0),.clk(gclk));
	jdff dff_A_ksfwVJTC7_0(.dout(w_dff_A_5nYDEzEt4_0),.din(w_dff_A_ksfwVJTC7_0),.clk(gclk));
	jdff dff_A_odu2dyA62_0(.dout(w_dff_A_ksfwVJTC7_0),.din(w_dff_A_odu2dyA62_0),.clk(gclk));
	jdff dff_A_Xz7dIdf21_0(.dout(w_dff_A_odu2dyA62_0),.din(w_dff_A_Xz7dIdf21_0),.clk(gclk));
	jdff dff_A_6Wv0SJQa4_0(.dout(w_dff_A_Xz7dIdf21_0),.din(w_dff_A_6Wv0SJQa4_0),.clk(gclk));
	jdff dff_A_5a8LTbLo0_0(.dout(w_dff_A_6Wv0SJQa4_0),.din(w_dff_A_5a8LTbLo0_0),.clk(gclk));
	jdff dff_A_4QBemBD09_0(.dout(w_dff_A_5a8LTbLo0_0),.din(w_dff_A_4QBemBD09_0),.clk(gclk));
	jdff dff_A_pupSgkaY3_0(.dout(w_dff_A_4QBemBD09_0),.din(w_dff_A_pupSgkaY3_0),.clk(gclk));
	jdff dff_A_k2FiQ56T2_0(.dout(w_dff_A_pupSgkaY3_0),.din(w_dff_A_k2FiQ56T2_0),.clk(gclk));
	jdff dff_A_Hq3tDri10_0(.dout(w_dff_A_k2FiQ56T2_0),.din(w_dff_A_Hq3tDri10_0),.clk(gclk));
	jdff dff_A_0D4s2Gdo9_1(.dout(w_n188_0[1]),.din(w_dff_A_0D4s2Gdo9_1),.clk(gclk));
	jdff dff_A_6uaFYpQ50_1(.dout(w_dff_A_0D4s2Gdo9_1),.din(w_dff_A_6uaFYpQ50_1),.clk(gclk));
	jdff dff_A_08ryss2d4_1(.dout(w_dff_A_6uaFYpQ50_1),.din(w_dff_A_08ryss2d4_1),.clk(gclk));
	jdff dff_A_yaIGEDZr2_1(.dout(w_dff_A_08ryss2d4_1),.din(w_dff_A_yaIGEDZr2_1),.clk(gclk));
	jdff dff_A_WGMDp3wy0_2(.dout(w_n188_0[2]),.din(w_dff_A_WGMDp3wy0_2),.clk(gclk));
	jdff dff_A_nNydAWo07_2(.dout(w_dff_A_WGMDp3wy0_2),.din(w_dff_A_nNydAWo07_2),.clk(gclk));
	jdff dff_A_QC21nsqe6_2(.dout(w_dff_A_nNydAWo07_2),.din(w_dff_A_QC21nsqe6_2),.clk(gclk));
	jdff dff_A_2jSnBeHT6_2(.dout(w_dff_A_QC21nsqe6_2),.din(w_dff_A_2jSnBeHT6_2),.clk(gclk));
	jdff dff_A_GA9OqbVz5_1(.dout(w_n103_1[1]),.din(w_dff_A_GA9OqbVz5_1),.clk(gclk));
	jdff dff_B_Xo319tDN4_1(.din(n98),.dout(w_dff_B_Xo319tDN4_1),.clk(gclk));
	jdff dff_A_hSz9sN5M7_0(.dout(w_G36gat_0[0]),.din(w_dff_A_hSz9sN5M7_0),.clk(gclk));
	jdff dff_A_yIlyZ2qw9_0(.dout(w_dff_A_hSz9sN5M7_0),.din(w_dff_A_yIlyZ2qw9_0),.clk(gclk));
	jdff dff_A_6A89NvFf1_0(.dout(w_dff_A_yIlyZ2qw9_0),.din(w_dff_A_6A89NvFf1_0),.clk(gclk));
	jdff dff_A_XHVa2PdQ6_0(.dout(w_dff_A_6A89NvFf1_0),.din(w_dff_A_XHVa2PdQ6_0),.clk(gclk));
	jdff dff_A_GSgHsgiB4_0(.dout(w_dff_A_XHVa2PdQ6_0),.din(w_dff_A_GSgHsgiB4_0),.clk(gclk));
	jdff dff_A_ZUy2e09b2_0(.dout(w_dff_A_GSgHsgiB4_0),.din(w_dff_A_ZUy2e09b2_0),.clk(gclk));
	jdff dff_A_5GamDoKq7_0(.dout(w_dff_A_ZUy2e09b2_0),.din(w_dff_A_5GamDoKq7_0),.clk(gclk));
	jdff dff_A_RVpORlXa0_0(.dout(w_dff_A_5GamDoKq7_0),.din(w_dff_A_RVpORlXa0_0),.clk(gclk));
	jdff dff_A_0zdwHsLo0_0(.dout(w_dff_A_RVpORlXa0_0),.din(w_dff_A_0zdwHsLo0_0),.clk(gclk));
	jdff dff_A_N9GJF8Yq0_0(.dout(w_dff_A_0zdwHsLo0_0),.din(w_dff_A_N9GJF8Yq0_0),.clk(gclk));
	jdff dff_A_7ogGRhSk8_0(.dout(w_G29gat_0[0]),.din(w_dff_A_7ogGRhSk8_0),.clk(gclk));
	jdff dff_A_epMiw4AP8_0(.dout(w_dff_A_7ogGRhSk8_0),.din(w_dff_A_epMiw4AP8_0),.clk(gclk));
	jdff dff_A_kJhRpB537_0(.dout(w_dff_A_epMiw4AP8_0),.din(w_dff_A_kJhRpB537_0),.clk(gclk));
	jdff dff_A_n6irMDDe0_0(.dout(w_dff_A_kJhRpB537_0),.din(w_dff_A_n6irMDDe0_0),.clk(gclk));
	jdff dff_A_fFBhEhC89_0(.dout(w_dff_A_n6irMDDe0_0),.din(w_dff_A_fFBhEhC89_0),.clk(gclk));
	jdff dff_A_7FKm4skU2_0(.dout(w_dff_A_fFBhEhC89_0),.din(w_dff_A_7FKm4skU2_0),.clk(gclk));
	jdff dff_A_CZbXNoCq5_0(.dout(w_dff_A_7FKm4skU2_0),.din(w_dff_A_CZbXNoCq5_0),.clk(gclk));
	jdff dff_A_s69AW2Fs6_0(.dout(w_dff_A_CZbXNoCq5_0),.din(w_dff_A_s69AW2Fs6_0),.clk(gclk));
	jdff dff_A_0LwUw7DL4_0(.dout(w_dff_A_s69AW2Fs6_0),.din(w_dff_A_0LwUw7DL4_0),.clk(gclk));
	jdff dff_A_NTUOQ2Dc1_0(.dout(w_dff_A_0LwUw7DL4_0),.din(w_dff_A_NTUOQ2Dc1_0),.clk(gclk));
	jdff dff_A_nH2CFQxK8_0(.dout(w_G50gat_0[0]),.din(w_dff_A_nH2CFQxK8_0),.clk(gclk));
	jdff dff_A_P0pATZpu5_0(.dout(w_dff_A_nH2CFQxK8_0),.din(w_dff_A_P0pATZpu5_0),.clk(gclk));
	jdff dff_A_CmV82uFf5_0(.dout(w_dff_A_P0pATZpu5_0),.din(w_dff_A_CmV82uFf5_0),.clk(gclk));
	jdff dff_A_ArnMqjTV9_0(.dout(w_dff_A_CmV82uFf5_0),.din(w_dff_A_ArnMqjTV9_0),.clk(gclk));
	jdff dff_A_7vLI3jZR5_0(.dout(w_dff_A_ArnMqjTV9_0),.din(w_dff_A_7vLI3jZR5_0),.clk(gclk));
	jdff dff_A_cU3b97YW4_0(.dout(w_dff_A_7vLI3jZR5_0),.din(w_dff_A_cU3b97YW4_0),.clk(gclk));
	jdff dff_A_vg3w83hV5_0(.dout(w_dff_A_cU3b97YW4_0),.din(w_dff_A_vg3w83hV5_0),.clk(gclk));
	jdff dff_A_ffnDFGgU1_0(.dout(w_dff_A_vg3w83hV5_0),.din(w_dff_A_ffnDFGgU1_0),.clk(gclk));
	jdff dff_A_RpaAdJF60_0(.dout(w_dff_A_ffnDFGgU1_0),.din(w_dff_A_RpaAdJF60_0),.clk(gclk));
	jdff dff_A_Xitz6zWQ0_0(.dout(w_dff_A_RpaAdJF60_0),.din(w_dff_A_Xitz6zWQ0_0),.clk(gclk));
	jdff dff_A_LxsrAVop3_0(.dout(w_G43gat_0[0]),.din(w_dff_A_LxsrAVop3_0),.clk(gclk));
	jdff dff_A_dWQcn0NB0_0(.dout(w_dff_A_LxsrAVop3_0),.din(w_dff_A_dWQcn0NB0_0),.clk(gclk));
	jdff dff_A_cv1xoxRd8_0(.dout(w_dff_A_dWQcn0NB0_0),.din(w_dff_A_cv1xoxRd8_0),.clk(gclk));
	jdff dff_A_Lqqu33rW4_0(.dout(w_dff_A_cv1xoxRd8_0),.din(w_dff_A_Lqqu33rW4_0),.clk(gclk));
	jdff dff_A_ZOxxSYZV7_0(.dout(w_dff_A_Lqqu33rW4_0),.din(w_dff_A_ZOxxSYZV7_0),.clk(gclk));
	jdff dff_A_vpAUhqgM5_0(.dout(w_dff_A_ZOxxSYZV7_0),.din(w_dff_A_vpAUhqgM5_0),.clk(gclk));
	jdff dff_A_jPksLCYx7_0(.dout(w_dff_A_vpAUhqgM5_0),.din(w_dff_A_jPksLCYx7_0),.clk(gclk));
	jdff dff_A_J9EUjqCr9_0(.dout(w_dff_A_jPksLCYx7_0),.din(w_dff_A_J9EUjqCr9_0),.clk(gclk));
	jdff dff_A_seiQmn7Y2_0(.dout(w_dff_A_J9EUjqCr9_0),.din(w_dff_A_seiQmn7Y2_0),.clk(gclk));
	jdff dff_A_hQ93Wxpt5_0(.dout(w_dff_A_seiQmn7Y2_0),.din(w_dff_A_hQ93Wxpt5_0),.clk(gclk));
	jdff dff_A_QdfBtJXe6_0(.dout(w_G92gat_0[0]),.din(w_dff_A_QdfBtJXe6_0),.clk(gclk));
	jdff dff_A_k9ev0bn76_0(.dout(w_dff_A_QdfBtJXe6_0),.din(w_dff_A_k9ev0bn76_0),.clk(gclk));
	jdff dff_A_6qXIiSgi8_0(.dout(w_dff_A_k9ev0bn76_0),.din(w_dff_A_6qXIiSgi8_0),.clk(gclk));
	jdff dff_A_G9wTVSPf9_0(.dout(w_dff_A_6qXIiSgi8_0),.din(w_dff_A_G9wTVSPf9_0),.clk(gclk));
	jdff dff_A_CTfT16IF5_0(.dout(w_dff_A_G9wTVSPf9_0),.din(w_dff_A_CTfT16IF5_0),.clk(gclk));
	jdff dff_A_ElqjSLiE6_0(.dout(w_dff_A_CTfT16IF5_0),.din(w_dff_A_ElqjSLiE6_0),.clk(gclk));
	jdff dff_A_TzOVK7Js5_0(.dout(w_dff_A_ElqjSLiE6_0),.din(w_dff_A_TzOVK7Js5_0),.clk(gclk));
	jdff dff_A_d84snmT29_0(.dout(w_dff_A_TzOVK7Js5_0),.din(w_dff_A_d84snmT29_0),.clk(gclk));
	jdff dff_A_6VTyIUdl5_0(.dout(w_dff_A_d84snmT29_0),.din(w_dff_A_6VTyIUdl5_0),.clk(gclk));
	jdff dff_A_8EXb0oLX9_0(.dout(w_dff_A_6VTyIUdl5_0),.din(w_dff_A_8EXb0oLX9_0),.clk(gclk));
	jdff dff_A_DwujNDRM0_0(.dout(w_G85gat_0[0]),.din(w_dff_A_DwujNDRM0_0),.clk(gclk));
	jdff dff_A_nOS9wDOF4_0(.dout(w_dff_A_DwujNDRM0_0),.din(w_dff_A_nOS9wDOF4_0),.clk(gclk));
	jdff dff_A_Td4g39v61_0(.dout(w_dff_A_nOS9wDOF4_0),.din(w_dff_A_Td4g39v61_0),.clk(gclk));
	jdff dff_A_qA4dQDjZ3_0(.dout(w_dff_A_Td4g39v61_0),.din(w_dff_A_qA4dQDjZ3_0),.clk(gclk));
	jdff dff_A_Vy1OX6oJ6_0(.dout(w_dff_A_qA4dQDjZ3_0),.din(w_dff_A_Vy1OX6oJ6_0),.clk(gclk));
	jdff dff_A_ViCNu6qF5_0(.dout(w_dff_A_Vy1OX6oJ6_0),.din(w_dff_A_ViCNu6qF5_0),.clk(gclk));
	jdff dff_A_pQiwXVJ70_0(.dout(w_dff_A_ViCNu6qF5_0),.din(w_dff_A_pQiwXVJ70_0),.clk(gclk));
	jdff dff_A_lhkC14OG6_0(.dout(w_dff_A_pQiwXVJ70_0),.din(w_dff_A_lhkC14OG6_0),.clk(gclk));
	jdff dff_A_JT5YBbSq8_0(.dout(w_dff_A_lhkC14OG6_0),.din(w_dff_A_JT5YBbSq8_0),.clk(gclk));
	jdff dff_A_mWGmOgUG6_0(.dout(w_dff_A_JT5YBbSq8_0),.din(w_dff_A_mWGmOgUG6_0),.clk(gclk));
	jdff dff_A_4Lr9U9Wf4_0(.dout(w_G106gat_0[0]),.din(w_dff_A_4Lr9U9Wf4_0),.clk(gclk));
	jdff dff_A_5bLXqItI0_0(.dout(w_dff_A_4Lr9U9Wf4_0),.din(w_dff_A_5bLXqItI0_0),.clk(gclk));
	jdff dff_A_qLA6ovTt7_0(.dout(w_dff_A_5bLXqItI0_0),.din(w_dff_A_qLA6ovTt7_0),.clk(gclk));
	jdff dff_A_mXyI7v1d2_0(.dout(w_dff_A_qLA6ovTt7_0),.din(w_dff_A_mXyI7v1d2_0),.clk(gclk));
	jdff dff_A_eLZtMan07_0(.dout(w_dff_A_mXyI7v1d2_0),.din(w_dff_A_eLZtMan07_0),.clk(gclk));
	jdff dff_A_rP3JqqWt2_0(.dout(w_dff_A_eLZtMan07_0),.din(w_dff_A_rP3JqqWt2_0),.clk(gclk));
	jdff dff_A_JjetcthL6_0(.dout(w_dff_A_rP3JqqWt2_0),.din(w_dff_A_JjetcthL6_0),.clk(gclk));
	jdff dff_A_a0MzTrRl1_0(.dout(w_dff_A_JjetcthL6_0),.din(w_dff_A_a0MzTrRl1_0),.clk(gclk));
	jdff dff_A_q2xmU7879_0(.dout(w_dff_A_a0MzTrRl1_0),.din(w_dff_A_q2xmU7879_0),.clk(gclk));
	jdff dff_A_8iNtpnhp8_0(.dout(w_dff_A_q2xmU7879_0),.din(w_dff_A_8iNtpnhp8_0),.clk(gclk));
	jdff dff_A_DrKOrulf4_0(.dout(w_G99gat_0[0]),.din(w_dff_A_DrKOrulf4_0),.clk(gclk));
	jdff dff_A_dqEL3aSt9_0(.dout(w_dff_A_DrKOrulf4_0),.din(w_dff_A_dqEL3aSt9_0),.clk(gclk));
	jdff dff_A_5fshzP8e3_0(.dout(w_dff_A_dqEL3aSt9_0),.din(w_dff_A_5fshzP8e3_0),.clk(gclk));
	jdff dff_A_iw9woJxl2_0(.dout(w_dff_A_5fshzP8e3_0),.din(w_dff_A_iw9woJxl2_0),.clk(gclk));
	jdff dff_A_3mtbQBH67_0(.dout(w_dff_A_iw9woJxl2_0),.din(w_dff_A_3mtbQBH67_0),.clk(gclk));
	jdff dff_A_omcknDYr7_0(.dout(w_dff_A_3mtbQBH67_0),.din(w_dff_A_omcknDYr7_0),.clk(gclk));
	jdff dff_A_PiXkER0f4_0(.dout(w_dff_A_omcknDYr7_0),.din(w_dff_A_PiXkER0f4_0),.clk(gclk));
	jdff dff_A_pbI64Yim0_0(.dout(w_dff_A_PiXkER0f4_0),.din(w_dff_A_pbI64Yim0_0),.clk(gclk));
	jdff dff_A_9qY27C2D5_0(.dout(w_dff_A_pbI64Yim0_0),.din(w_dff_A_9qY27C2D5_0),.clk(gclk));
	jdff dff_A_M4t8SJ0K9_0(.dout(w_dff_A_9qY27C2D5_0),.din(w_dff_A_M4t8SJ0K9_0),.clk(gclk));
	jdff dff_A_aEnsqv513_0(.dout(w_G162gat_0[0]),.din(w_dff_A_aEnsqv513_0),.clk(gclk));
	jdff dff_A_Dbdk0u5X4_0(.dout(w_dff_A_aEnsqv513_0),.din(w_dff_A_Dbdk0u5X4_0),.clk(gclk));
	jdff dff_A_zoXouxbX3_0(.dout(w_dff_A_Dbdk0u5X4_0),.din(w_dff_A_zoXouxbX3_0),.clk(gclk));
	jdff dff_A_nI7xrFNy1_0(.dout(w_dff_A_zoXouxbX3_0),.din(w_dff_A_nI7xrFNy1_0),.clk(gclk));
	jdff dff_A_fXfTq2In2_0(.dout(w_dff_A_nI7xrFNy1_0),.din(w_dff_A_fXfTq2In2_0),.clk(gclk));
	jdff dff_A_LKggevtQ5_0(.dout(w_dff_A_fXfTq2In2_0),.din(w_dff_A_LKggevtQ5_0),.clk(gclk));
	jdff dff_A_o9NgQYoj2_0(.dout(w_dff_A_LKggevtQ5_0),.din(w_dff_A_o9NgQYoj2_0),.clk(gclk));
	jdff dff_A_aydRc4zT7_0(.dout(w_dff_A_o9NgQYoj2_0),.din(w_dff_A_aydRc4zT7_0),.clk(gclk));
	jdff dff_A_VO7Uf5QN5_0(.dout(w_dff_A_aydRc4zT7_0),.din(w_dff_A_VO7Uf5QN5_0),.clk(gclk));
	jdff dff_A_ePkpiFcd3_0(.dout(w_dff_A_VO7Uf5QN5_0),.din(w_dff_A_ePkpiFcd3_0),.clk(gclk));
	jdff dff_A_Hy9M0DwN2_0(.dout(w_G134gat_0[0]),.din(w_dff_A_Hy9M0DwN2_0),.clk(gclk));
	jdff dff_A_7PMAeOua3_0(.dout(w_dff_A_Hy9M0DwN2_0),.din(w_dff_A_7PMAeOua3_0),.clk(gclk));
	jdff dff_A_9fg9i70z2_0(.dout(w_dff_A_7PMAeOua3_0),.din(w_dff_A_9fg9i70z2_0),.clk(gclk));
	jdff dff_A_aoAzma2Y8_0(.dout(w_dff_A_9fg9i70z2_0),.din(w_dff_A_aoAzma2Y8_0),.clk(gclk));
	jdff dff_A_um6aLhpZ4_0(.dout(w_dff_A_aoAzma2Y8_0),.din(w_dff_A_um6aLhpZ4_0),.clk(gclk));
	jdff dff_A_gPhuAdES2_0(.dout(w_dff_A_um6aLhpZ4_0),.din(w_dff_A_gPhuAdES2_0),.clk(gclk));
	jdff dff_A_4kILrvpf1_0(.dout(w_dff_A_gPhuAdES2_0),.din(w_dff_A_4kILrvpf1_0),.clk(gclk));
	jdff dff_A_XtZcJDB85_0(.dout(w_dff_A_4kILrvpf1_0),.din(w_dff_A_XtZcJDB85_0),.clk(gclk));
	jdff dff_A_3utV0gN68_0(.dout(w_dff_A_XtZcJDB85_0),.din(w_dff_A_3utV0gN68_0),.clk(gclk));
	jdff dff_A_EBGdVPH94_0(.dout(w_dff_A_3utV0gN68_0),.din(w_dff_A_EBGdVPH94_0),.clk(gclk));
	jdff dff_A_N1sW4CcE8_0(.dout(w_G218gat_0[0]),.din(w_dff_A_N1sW4CcE8_0),.clk(gclk));
	jdff dff_A_oOJ2sYzY8_0(.dout(w_dff_A_N1sW4CcE8_0),.din(w_dff_A_oOJ2sYzY8_0),.clk(gclk));
	jdff dff_A_nMV08u7c0_0(.dout(w_dff_A_oOJ2sYzY8_0),.din(w_dff_A_nMV08u7c0_0),.clk(gclk));
	jdff dff_A_Ga2VoN8N9_0(.dout(w_dff_A_nMV08u7c0_0),.din(w_dff_A_Ga2VoN8N9_0),.clk(gclk));
	jdff dff_A_JvPUZ4wM5_0(.dout(w_dff_A_Ga2VoN8N9_0),.din(w_dff_A_JvPUZ4wM5_0),.clk(gclk));
	jdff dff_A_Pe3402fb4_0(.dout(w_dff_A_JvPUZ4wM5_0),.din(w_dff_A_Pe3402fb4_0),.clk(gclk));
	jdff dff_A_5qBKOiqD8_0(.dout(w_dff_A_Pe3402fb4_0),.din(w_dff_A_5qBKOiqD8_0),.clk(gclk));
	jdff dff_A_0uWmPsc89_0(.dout(w_dff_A_5qBKOiqD8_0),.din(w_dff_A_0uWmPsc89_0),.clk(gclk));
	jdff dff_A_lZx38iLY4_0(.dout(w_dff_A_0uWmPsc89_0),.din(w_dff_A_lZx38iLY4_0),.clk(gclk));
	jdff dff_A_Mih6RlS80_0(.dout(w_dff_A_lZx38iLY4_0),.din(w_dff_A_Mih6RlS80_0),.clk(gclk));
	jdff dff_A_0lyfOHWN2_0(.dout(w_G190gat_0[0]),.din(w_dff_A_0lyfOHWN2_0),.clk(gclk));
	jdff dff_A_wlwr0xjB8_0(.dout(w_dff_A_0lyfOHWN2_0),.din(w_dff_A_wlwr0xjB8_0),.clk(gclk));
	jdff dff_A_qfBUllui9_0(.dout(w_dff_A_wlwr0xjB8_0),.din(w_dff_A_qfBUllui9_0),.clk(gclk));
	jdff dff_A_L11IOaEB3_0(.dout(w_dff_A_qfBUllui9_0),.din(w_dff_A_L11IOaEB3_0),.clk(gclk));
	jdff dff_A_1EMa7xGF8_0(.dout(w_dff_A_L11IOaEB3_0),.din(w_dff_A_1EMa7xGF8_0),.clk(gclk));
	jdff dff_A_vvwYoSry0_0(.dout(w_dff_A_1EMa7xGF8_0),.din(w_dff_A_vvwYoSry0_0),.clk(gclk));
	jdff dff_A_svDUcBLl9_0(.dout(w_dff_A_vvwYoSry0_0),.din(w_dff_A_svDUcBLl9_0),.clk(gclk));
	jdff dff_A_ItiD22yw2_0(.dout(w_dff_A_svDUcBLl9_0),.din(w_dff_A_ItiD22yw2_0),.clk(gclk));
	jdff dff_A_a15osvgB0_0(.dout(w_dff_A_ItiD22yw2_0),.din(w_dff_A_a15osvgB0_0),.clk(gclk));
	jdff dff_A_rrUk5ZKY3_0(.dout(w_dff_A_a15osvgB0_0),.din(w_dff_A_rrUk5ZKY3_0),.clk(gclk));
endmodule

