/*

c3540:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jdff: 1943
	jand: 535
	jor: 374

Summary:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jdff: 1943
	jand: 535
	jor: 374
*/

module c3540(gclk, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402);
	input gclk;
	input G1;
	input G13;
	input G20;
	input G33;
	input G41;
	input G45;
	input G50;
	input G58;
	input G68;
	input G77;
	input G87;
	input G97;
	input G107;
	input G116;
	input G124;
	input G125;
	input G128;
	input G132;
	input G137;
	input G143;
	input G150;
	input G159;
	input G169;
	input G179;
	input G190;
	input G200;
	input G213;
	input G222;
	input G223;
	input G226;
	input G232;
	input G238;
	input G244;
	input G250;
	input G257;
	input G264;
	input G270;
	input G274;
	input G283;
	input G294;
	input G303;
	input G311;
	input G317;
	input G322;
	input G326;
	input G329;
	input G330;
	input G343;
	input G1698;
	input G2897;
	output G353;
	output G355;
	output G361;
	output G358;
	output G351;
	output G372;
	output G369;
	output G399;
	output G364;
	output G396;
	output G384;
	output G367;
	output G387;
	output G393;
	output G390;
	output G378;
	output G375;
	output G381;
	output G407;
	output G409;
	output G405;
	output G402;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [2:0] w_G1_2;
	wire [1:0] w_G1_3;
	wire [2:0] w_G13_0;
	wire [1:0] w_G13_1;
	wire [2:0] w_G20_0;
	wire [2:0] w_G20_1;
	wire [2:0] w_G20_2;
	wire [2:0] w_G20_3;
	wire [2:0] w_G20_4;
	wire [2:0] w_G20_5;
	wire [2:0] w_G20_6;
	wire [1:0] w_G20_7;
	wire [2:0] w_G33_0;
	wire [2:0] w_G33_1;
	wire [2:0] w_G33_2;
	wire [2:0] w_G33_3;
	wire [2:0] w_G33_4;
	wire [2:0] w_G33_5;
	wire [2:0] w_G33_6;
	wire [2:0] w_G33_7;
	wire [2:0] w_G33_8;
	wire [2:0] w_G33_9;
	wire [2:0] w_G33_10;
	wire [2:0] w_G33_11;
	wire [2:0] w_G41_0;
	wire [1:0] w_G41_1;
	wire [2:0] w_G45_0;
	wire [2:0] w_G45_1;
	wire [2:0] w_G50_0;
	wire [2:0] w_G50_1;
	wire [2:0] w_G50_2;
	wire [2:0] w_G50_3;
	wire [2:0] w_G50_4;
	wire [2:0] w_G50_5;
	wire [2:0] w_G58_0;
	wire [2:0] w_G58_1;
	wire [2:0] w_G58_2;
	wire [2:0] w_G58_3;
	wire [2:0] w_G58_4;
	wire [1:0] w_G58_5;
	wire [2:0] w_G68_0;
	wire [2:0] w_G68_1;
	wire [2:0] w_G68_2;
	wire [2:0] w_G68_3;
	wire [2:0] w_G68_4;
	wire [1:0] w_G68_5;
	wire [2:0] w_G77_0;
	wire [2:0] w_G77_1;
	wire [2:0] w_G77_2;
	wire [2:0] w_G77_3;
	wire [2:0] w_G77_4;
	wire [1:0] w_G77_5;
	wire [2:0] w_G87_0;
	wire [2:0] w_G87_1;
	wire [2:0] w_G87_2;
	wire [2:0] w_G87_3;
	wire [2:0] w_G97_0;
	wire [2:0] w_G97_1;
	wire [2:0] w_G97_2;
	wire [2:0] w_G97_3;
	wire [2:0] w_G97_4;
	wire [1:0] w_G97_5;
	wire [2:0] w_G107_0;
	wire [2:0] w_G107_1;
	wire [2:0] w_G107_2;
	wire [2:0] w_G107_3;
	wire [2:0] w_G107_4;
	wire [1:0] w_G107_5;
	wire [2:0] w_G116_0;
	wire [2:0] w_G116_1;
	wire [2:0] w_G116_2;
	wire [2:0] w_G116_3;
	wire [2:0] w_G116_4;
	wire [1:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [2:0] w_G132_0;
	wire [1:0] w_G132_1;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G143_0;
	wire [2:0] w_G143_1;
	wire [1:0] w_G143_2;
	wire [2:0] w_G150_0;
	wire [2:0] w_G150_1;
	wire [2:0] w_G150_2;
	wire [1:0] w_G150_3;
	wire [2:0] w_G159_0;
	wire [2:0] w_G159_1;
	wire [2:0] w_G159_2;
	wire [2:0] w_G159_3;
	wire [2:0] w_G169_0;
	wire [1:0] w_G169_1;
	wire [2:0] w_G179_0;
	wire [2:0] w_G179_1;
	wire [2:0] w_G179_2;
	wire [2:0] w_G190_0;
	wire [2:0] w_G190_1;
	wire [2:0] w_G190_2;
	wire [2:0] w_G190_3;
	wire [1:0] w_G190_4;
	wire [2:0] w_G200_0;
	wire [2:0] w_G200_1;
	wire [2:0] w_G200_2;
	wire [2:0] w_G200_3;
	wire [2:0] w_G200_4;
	wire [2:0] w_G213_0;
	wire [1:0] w_G223_0;
	wire [2:0] w_G226_0;
	wire [1:0] w_G226_1;
	wire [2:0] w_G232_0;
	wire [2:0] w_G232_1;
	wire [2:0] w_G238_0;
	wire [2:0] w_G238_1;
	wire [2:0] w_G244_0;
	wire [2:0] w_G244_1;
	wire [2:0] w_G250_0;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [2:0] w_G264_0;
	wire [1:0] w_G264_1;
	wire [2:0] w_G270_0;
	wire [2:0] w_G274_0;
	wire [2:0] w_G283_0;
	wire [2:0] w_G283_1;
	wire [2:0] w_G283_2;
	wire [2:0] w_G283_3;
	wire [2:0] w_G294_0;
	wire [2:0] w_G294_1;
	wire [2:0] w_G294_2;
	wire [1:0] w_G294_3;
	wire [2:0] w_G303_0;
	wire [2:0] w_G303_1;
	wire [2:0] w_G303_2;
	wire [2:0] w_G311_0;
	wire [2:0] w_G311_1;
	wire [2:0] w_G317_0;
	wire [1:0] w_G317_1;
	wire [2:0] w_G322_0;
	wire [1:0] w_G326_0;
	wire [1:0] w_G330_0;
	wire [1:0] w_G343_0;
	wire [2:0] w_G1698_0;
	wire w_G355_0;
	wire G355_fa_;
	wire [1:0] w_G396_0;
	wire G396_fa_;
	wire w_G384_0;
	wire G384_fa_;
	wire [1:0] w_G387_0;
	wire G387_fa_;
	wire [2:0] w_n72_0;
	wire [1:0] w_n72_1;
	wire [2:0] w_n73_0;
	wire [2:0] w_n73_1;
	wire [2:0] w_n73_2;
	wire [2:0] w_n74_0;
	wire [1:0] w_n74_1;
	wire [2:0] w_n75_0;
	wire [1:0] w_n75_1;
	wire [1:0] w_n76_0;
	wire [1:0] w_n77_0;
	wire [2:0] w_n79_0;
	wire [2:0] w_n80_0;
	wire [1:0] w_n80_1;
	wire [2:0] w_n81_0;
	wire [2:0] w_n85_0;
	wire [1:0] w_n86_0;
	wire [2:0] w_n88_0;
	wire [1:0] w_n88_1;
	wire [2:0] w_n91_0;
	wire [2:0] w_n91_1;
	wire [1:0] w_n93_0;
	wire [2:0] w_n97_0;
	wire [2:0] w_n97_1;
	wire [1:0] w_n97_2;
	wire [2:0] w_n98_0;
	wire [2:0] w_n98_1;
	wire [1:0] w_n98_2;
	wire [2:0] w_n103_0;
	wire [2:0] w_n105_0;
	wire [2:0] w_n105_1;
	wire [1:0] w_n105_2;
	wire [1:0] w_n106_0;
	wire [2:0] w_n112_0;
	wire [2:0] w_n112_1;
	wire [2:0] w_n112_2;
	wire [2:0] w_n112_3;
	wire [2:0] w_n112_4;
	wire [2:0] w_n112_5;
	wire [2:0] w_n113_0;
	wire [2:0] w_n113_1;
	wire [2:0] w_n113_2;
	wire [1:0] w_n113_3;
	wire [2:0] w_n114_0;
	wire [2:0] w_n114_1;
	wire [2:0] w_n115_0;
	wire [1:0] w_n115_1;
	wire [1:0] w_n116_0;
	wire [2:0] w_n118_0;
	wire [2:0] w_n121_0;
	wire [2:0] w_n122_0;
	wire [1:0] w_n122_1;
	wire [2:0] w_n123_0;
	wire [2:0] w_n123_1;
	wire [1:0] w_n131_0;
	wire [1:0] w_n135_0;
	wire [2:0] w_n137_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n144_0;
	wire [2:0] w_n146_0;
	wire [2:0] w_n146_1;
	wire [2:0] w_n146_2;
	wire [2:0] w_n146_3;
	wire [2:0] w_n147_0;
	wire [2:0] w_n148_0;
	wire [2:0] w_n148_1;
	wire [2:0] w_n148_2;
	wire [2:0] w_n148_3;
	wire [2:0] w_n148_4;
	wire [2:0] w_n148_5;
	wire [2:0] w_n148_6;
	wire [2:0] w_n148_7;
	wire [2:0] w_n148_8;
	wire [2:0] w_n148_9;
	wire [2:0] w_n149_0;
	wire [2:0] w_n149_1;
	wire [1:0] w_n149_2;
	wire [2:0] w_n151_0;
	wire [2:0] w_n151_1;
	wire [2:0] w_n151_2;
	wire [2:0] w_n151_3;
	wire [2:0] w_n151_4;
	wire [2:0] w_n152_0;
	wire [2:0] w_n152_1;
	wire [2:0] w_n152_2;
	wire [1:0] w_n152_3;
	wire [1:0] w_n154_0;
	wire [2:0] w_n155_0;
	wire [2:0] w_n155_1;
	wire [2:0] w_n155_2;
	wire [1:0] w_n155_3;
	wire [2:0] w_n157_0;
	wire [2:0] w_n161_0;
	wire [1:0] w_n161_1;
	wire [2:0] w_n162_0;
	wire [1:0] w_n163_0;
	wire [2:0] w_n166_0;
	wire [2:0] w_n166_1;
	wire [2:0] w_n166_2;
	wire [1:0] w_n166_3;
	wire [2:0] w_n170_0;
	wire [1:0] w_n172_0;
	wire [2:0] w_n179_0;
	wire [2:0] w_n179_1;
	wire [1:0] w_n180_0;
	wire [2:0] w_n185_0;
	wire [2:0] w_n185_1;
	wire [2:0] w_n185_2;
	wire [2:0] w_n185_3;
	wire [2:0] w_n189_0;
	wire [2:0] w_n189_1;
	wire [1:0] w_n189_2;
	wire [2:0] w_n190_0;
	wire [2:0] w_n190_1;
	wire [2:0] w_n191_0;
	wire [1:0] w_n195_0;
	wire [2:0] w_n196_0;
	wire [2:0] w_n196_1;
	wire [2:0] w_n196_2;
	wire [2:0] w_n197_0;
	wire [1:0] w_n197_1;
	wire [2:0] w_n199_0;
	wire [1:0] w_n199_1;
	wire [1:0] w_n201_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n206_0;
	wire [2:0] w_n210_0;
	wire [1:0] w_n213_0;
	wire [1:0] w_n214_0;
	wire [1:0] w_n218_0;
	wire [1:0] w_n219_0;
	wire [2:0] w_n221_0;
	wire [1:0] w_n228_0;
	wire [2:0] w_n229_0;
	wire [1:0] w_n230_0;
	wire [2:0] w_n231_0;
	wire [2:0] w_n234_0;
	wire [1:0] w_n241_0;
	wire [2:0] w_n242_0;
	wire [2:0] w_n243_0;
	wire [2:0] w_n246_0;
	wire [1:0] w_n246_1;
	wire [1:0] w_n249_0;
	wire [1:0] w_n255_0;
	wire [1:0] w_n257_0;
	wire [1:0] w_n259_0;
	wire [1:0] w_n261_0;
	wire [1:0] w_n262_0;
	wire [2:0] w_n269_0;
	wire [2:0] w_n269_1;
	wire [1:0] w_n270_0;
	wire [2:0] w_n271_0;
	wire [2:0] w_n271_1;
	wire [2:0] w_n274_0;
	wire [1:0] w_n278_0;
	wire [1:0] w_n279_0;
	wire [1:0] w_n281_0;
	wire [2:0] w_n288_0;
	wire [1:0] w_n288_1;
	wire [1:0] w_n296_0;
	wire [1:0] w_n298_0;
	wire [1:0] w_n300_0;
	wire [1:0] w_n303_0;
	wire [2:0] w_n312_0;
	wire [1:0] w_n312_1;
	wire [1:0] w_n315_0;
	wire [1:0] w_n320_0;
	wire [1:0] w_n324_0;
	wire [1:0] w_n328_0;
	wire [1:0] w_n334_0;
	wire [1:0] w_n339_0;
	wire [2:0] w_n346_0;
	wire [1:0] w_n346_1;
	wire [2:0] w_n355_0;
	wire [1:0] w_n355_1;
	wire [1:0] w_n362_0;
	wire [2:0] w_n367_0;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n374_0;
	wire [1:0] w_n381_0;
	wire [2:0] w_n382_0;
	wire [1:0] w_n382_1;
	wire [2:0] w_n385_0;
	wire [1:0] w_n385_1;
	wire [2:0] w_n387_0;
	wire [1:0] w_n387_1;
	wire [1:0] w_n390_0;
	wire [2:0] w_n401_0;
	wire [2:0] w_n404_0;
	wire [1:0] w_n405_0;
	wire [2:0] w_n407_0;
	wire [2:0] w_n407_1;
	wire [1:0] w_n407_2;
	wire [1:0] w_n412_0;
	wire [2:0] w_n420_0;
	wire [1:0] w_n420_1;
	wire [2:0] w_n425_0;
	wire [2:0] w_n425_1;
	wire [1:0] w_n426_0;
	wire [1:0] w_n430_0;
	wire [2:0] w_n436_0;
	wire [2:0] w_n439_0;
	wire [1:0] w_n439_1;
	wire [1:0] w_n445_0;
	wire [1:0] w_n446_0;
	wire [2:0] w_n455_0;
	wire [2:0] w_n462_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n474_0;
	wire [1:0] w_n475_0;
	wire [1:0] w_n478_0;
	wire [1:0] w_n479_0;
	wire [1:0] w_n483_0;
	wire [1:0] w_n484_0;
	wire [2:0] w_n492_0;
	wire [1:0] w_n507_0;
	wire [1:0] w_n508_0;
	wire [1:0] w_n511_0;
	wire [1:0] w_n512_0;
	wire [1:0] w_n516_0;
	wire [1:0] w_n517_0;
	wire [2:0] w_n519_0;
	wire [2:0] w_n519_1;
	wire [1:0] w_n523_0;
	wire [1:0] w_n524_0;
	wire [1:0] w_n528_0;
	wire [1:0] w_n532_0;
	wire [1:0] w_n534_0;
	wire [2:0] w_n536_0;
	wire [1:0] w_n539_0;
	wire [1:0] w_n541_0;
	wire [2:0] w_n542_0;
	wire [1:0] w_n543_0;
	wire [2:0] w_n548_0;
	wire [1:0] w_n550_0;
	wire [2:0] w_n552_0;
	wire [1:0] w_n552_1;
	wire [2:0] w_n553_0;
	wire [2:0] w_n553_1;
	wire [2:0] w_n553_2;
	wire [2:0] w_n554_0;
	wire [2:0] w_n554_1;
	wire [2:0] w_n554_2;
	wire [2:0] w_n554_3;
	wire [1:0] w_n556_0;
	wire [1:0] w_n557_0;
	wire [2:0] w_n561_0;
	wire [2:0] w_n563_0;
	wire [1:0] w_n564_0;
	wire [1:0] w_n565_0;
	wire [1:0] w_n567_0;
	wire [2:0] w_n571_0;
	wire [2:0] w_n572_0;
	wire [2:0] w_n573_0;
	wire [2:0] w_n576_0;
	wire [1:0] w_n576_1;
	wire [2:0] w_n588_0;
	wire [1:0] w_n588_1;
	wire [2:0] w_n589_0;
	wire [2:0] w_n589_1;
	wire [2:0] w_n591_0;
	wire [1:0] w_n591_1;
	wire [2:0] w_n592_0;
	wire [2:0] w_n592_1;
	wire [1:0] w_n592_2;
	wire [2:0] w_n593_0;
	wire [1:0] w_n602_0;
	wire [2:0] w_n603_0;
	wire [2:0] w_n603_1;
	wire [1:0] w_n603_2;
	wire [2:0] w_n604_0;
	wire [2:0] w_n604_1;
	wire [1:0] w_n604_2;
	wire [2:0] w_n605_0;
	wire [2:0] w_n605_1;
	wire [2:0] w_n608_0;
	wire [2:0] w_n608_1;
	wire [2:0] w_n612_0;
	wire [2:0] w_n612_1;
	wire [2:0] w_n612_2;
	wire [2:0] w_n612_3;
	wire [1:0] w_n612_4;
	wire [2:0] w_n613_0;
	wire [1:0] w_n613_1;
	wire [1:0] w_n615_0;
	wire [1:0] w_n616_0;
	wire [2:0] w_n617_0;
	wire [2:0] w_n617_1;
	wire [2:0] w_n617_2;
	wire [2:0] w_n617_3;
	wire [2:0] w_n617_4;
	wire [2:0] w_n617_5;
	wire [1:0] w_n617_6;
	wire [1:0] w_n619_0;
	wire [1:0] w_n622_0;
	wire [2:0] w_n623_0;
	wire [2:0] w_n623_1;
	wire [2:0] w_n623_2;
	wire [2:0] w_n623_3;
	wire [2:0] w_n623_4;
	wire [1:0] w_n623_5;
	wire [1:0] w_n626_0;
	wire [2:0] w_n627_0;
	wire [2:0] w_n627_1;
	wire [2:0] w_n627_2;
	wire [2:0] w_n627_3;
	wire [2:0] w_n627_4;
	wire [2:0] w_n627_5;
	wire [2:0] w_n627_6;
	wire [1:0] w_n627_7;
	wire [2:0] w_n631_0;
	wire [2:0] w_n631_1;
	wire [2:0] w_n631_2;
	wire [2:0] w_n631_3;
	wire [2:0] w_n631_4;
	wire [2:0] w_n631_5;
	wire [2:0] w_n631_6;
	wire [1:0] w_n631_7;
	wire [2:0] w_n634_0;
	wire [2:0] w_n634_1;
	wire [2:0] w_n634_2;
	wire [2:0] w_n634_3;
	wire [1:0] w_n634_4;
	wire [2:0] w_n636_0;
	wire [2:0] w_n636_1;
	wire [2:0] w_n636_2;
	wire [2:0] w_n636_3;
	wire [2:0] w_n636_4;
	wire [2:0] w_n636_5;
	wire [2:0] w_n636_6;
	wire [1:0] w_n636_7;
	wire [1:0] w_n639_0;
	wire [2:0] w_n640_0;
	wire [2:0] w_n640_1;
	wire [2:0] w_n640_2;
	wire [2:0] w_n640_3;
	wire [2:0] w_n640_4;
	wire [2:0] w_n640_5;
	wire [2:0] w_n640_6;
	wire [1:0] w_n640_7;
	wire [2:0] w_n642_0;
	wire [2:0] w_n642_1;
	wire [2:0] w_n642_2;
	wire [2:0] w_n642_3;
	wire [2:0] w_n642_4;
	wire [2:0] w_n642_5;
	wire [2:0] w_n642_6;
	wire [1:0] w_n642_7;
	wire [1:0] w_n654_0;
	wire [1:0] w_n657_0;
	wire [1:0] w_n661_0;
	wire [2:0] w_n672_0;
	wire [1:0] w_n672_1;
	wire [2:0] w_n675_0;
	wire [1:0] w_n676_0;
	wire [1:0] w_n680_0;
	wire [1:0] w_n692_0;
	wire [2:0] w_n696_0;
	wire [2:0] w_n696_1;
	wire [1:0] w_n717_0;
	wire [1:0] w_n728_0;
	wire [2:0] w_n743_0;
	wire [1:0] w_n743_1;
	wire [1:0] w_n750_0;
	wire [1:0] w_n754_0;
	wire [2:0] w_n758_0;
	wire [1:0] w_n758_1;
	wire [1:0] w_n759_0;
	wire [1:0] w_n760_0;
	wire [2:0] w_n764_0;
	wire [2:0] w_n764_1;
	wire [1:0] w_n769_0;
	wire [2:0] w_n771_0;
	wire [1:0] w_n779_0;
	wire [1:0] w_n797_0;
	wire [1:0] w_n801_0;
	wire [1:0] w_n816_0;
	wire [1:0] w_n823_0;
	wire [1:0] w_n825_0;
	wire [2:0] w_n853_0;
	wire [2:0] w_n855_0;
	wire [2:0] w_n861_0;
	wire [1:0] w_n861_1;
	wire [1:0] w_n863_0;
	wire [1:0] w_n864_0;
	wire [1:0] w_n899_0;
	wire [1:0] w_n909_0;
	wire [2:0] w_n937_0;
	wire [1:0] w_n940_0;
	wire [1:0] w_n962_0;
	wire [2:0] w_n988_0;
	wire [1:0] w_n990_0;
	wire [2:0] w_n991_0;
	wire [1:0] w_n992_0;
	wire [2:0] w_n994_0;
	wire [2:0] w_n996_0;
	wire [1:0] w_n999_0;
	wire [2:0] w_n1001_0;
	wire [2:0] w_n1002_0;
	wire [1:0] w_n1003_0;
	wire [2:0] w_n1049_0;
	wire [1:0] w_n1052_0;
	wire [1:0] w_n1057_0;
	wire [1:0] w_n1059_0;
	wire [1:0] w_n1088_0;
	wire [2:0] w_n1114_0;
	wire [2:0] w_n1162_0;
	wire [1:0] w_n1164_0;
	wire [1:0] w_n1172_0;
	wire [1:0] w_n1175_0;
	wire [1:0] w_n1183_0;
	wire [1:0] w_n1184_0;
	wire [1:0] w_n1187_0;
	wire w_dff_B_27IG3dus8_1;
	wire w_dff_B_brpxkulE2_0;
	wire w_dff_B_OdmNiY9Q7_0;
	wire w_dff_A_oKzhe3GQ7_1;
	wire w_dff_A_KZg6e6nu4_1;
	wire w_dff_A_b2IsJz1y0_0;
	wire w_dff_B_P1MteBTm6_1;
	wire w_dff_B_VcQ3QnV95_0;
	wire w_dff_B_0KF7IW7h5_0;
	wire w_dff_B_khbgpzw24_0;
	wire w_dff_B_UkrzfmdC8_0;
	wire w_dff_B_kaCxY0zh4_0;
	wire w_dff_B_1nhceMPk4_0;
	wire w_dff_B_SHGn3OUc7_0;
	wire w_dff_B_tCOiiRT90_0;
	wire w_dff_B_T8MWrgiF9_0;
	wire w_dff_B_CQkULghC5_0;
	wire w_dff_B_EWujXDTd0_0;
	wire w_dff_B_LX6rMsV55_0;
	wire w_dff_B_0gYPtSiV2_0;
	wire w_dff_B_m3YYBuz63_0;
	wire w_dff_B_xvy5vnMy1_0;
	wire w_dff_B_5L7Inghj0_0;
	wire w_dff_B_rHWr3kVT1_0;
	wire w_dff_B_y3xYfgSg7_0;
	wire w_dff_B_HMSjkaM36_0;
	wire w_dff_B_XrsLfFOK7_0;
	wire w_dff_B_tNTamC3K6_0;
	wire w_dff_B_9rLj559m2_0;
	wire w_dff_B_Fy6euJsy2_0;
	wire w_dff_B_05mxwore0_0;
	wire w_dff_B_FkBCJ4Gk0_0;
	wire w_dff_B_17rdGTZ48_0;
	wire w_dff_B_mgTPp4yG5_0;
	wire w_dff_B_qqINFvwM6_0;
	wire w_dff_B_07cq4XHF0_1;
	wire w_dff_B_oehH8Av27_0;
	wire w_dff_B_LsPz2THP9_0;
	wire w_dff_B_eQEFrEFx6_0;
	wire w_dff_B_gbjR7sTU1_0;
	wire w_dff_B_8e36eyeG0_0;
	wire w_dff_B_iDQYgquA2_0;
	wire w_dff_B_S6qopbMi1_0;
	wire w_dff_B_y1uw5VNx6_0;
	wire w_dff_B_jNbPZpET7_0;
	wire w_dff_B_90YbSXgM0_0;
	wire w_dff_B_HLxDSfFW2_0;
	wire w_dff_B_tZULgeE83_0;
	wire w_dff_B_N0U1Ql070_0;
	wire w_dff_B_5JVTNJGQ0_0;
	wire w_dff_B_ZqvK0iFu6_0;
	wire w_dff_B_QDRAx9Hn9_0;
	wire w_dff_B_C6syMAPg1_0;
	wire w_dff_B_9O43Ezeg7_0;
	wire w_dff_B_bvj5x9wr1_0;
	wire w_dff_A_Wp42wl8u7_1;
	wire w_dff_A_L1JiYjgh4_1;
	wire w_dff_B_6KOFtQeg5_0;
	wire w_dff_A_3432eBZr8_0;
	wire w_dff_B_meZ7zUbD1_1;
	wire w_dff_A_cxfiEA5b1_0;
	wire w_dff_B_bxV1Hvf69_1;
	wire w_dff_B_dCbiIkUu2_1;
	wire w_dff_B_ltsCm6fP4_1;
	wire w_dff_B_snMa3UHB8_1;
	wire w_dff_B_86oEXe4D6_1;
	wire w_dff_B_EH4oItPu9_1;
	wire w_dff_B_hLXk1Tdo1_1;
	wire w_dff_B_vbuZhOVL4_1;
	wire w_dff_B_KvLiyaVF0_1;
	wire w_dff_B_tmHNNuv62_1;
	wire w_dff_B_5dTyv3FO1_1;
	wire w_dff_B_7R0XxOkQ1_1;
	wire w_dff_B_Js4S65zn1_1;
	wire w_dff_B_BjpQtCIc2_1;
	wire w_dff_B_27XFPe0M5_1;
	wire w_dff_B_WgMwadz85_1;
	wire w_dff_B_RKoL6UN74_1;
	wire w_dff_B_At1DnCxB3_1;
	wire w_dff_B_x7bO9Ypj8_1;
	wire w_dff_B_I4BoaXlS4_1;
	wire w_dff_B_qSe9mCK36_1;
	wire w_dff_B_8Y0PSoG76_1;
	wire w_dff_B_7CIeihSw2_1;
	wire w_dff_B_RHlzz7bS4_1;
	wire w_dff_B_0GIqr2mo9_1;
	wire w_dff_B_zk7gRSOB7_1;
	wire w_dff_A_lED9eLgz9_0;
	wire w_dff_B_a5t1mwIU9_1;
	wire w_dff_B_pqHyahDE9_1;
	wire w_dff_B_8PLgku0F9_1;
	wire w_dff_B_YQwWnxHW1_1;
	wire w_dff_B_eOVT77cD4_1;
	wire w_dff_B_EsSZhU0t7_1;
	wire w_dff_B_7W6IxzaU9_1;
	wire w_dff_B_5pwmVud73_1;
	wire w_dff_B_iyKO1Vem0_1;
	wire w_dff_B_sY70pu2D3_1;
	wire w_dff_B_FRzAIkLh2_1;
	wire w_dff_B_Rxfz5tES0_1;
	wire w_dff_B_O3zsCVqI7_1;
	wire w_dff_B_BBvpIZVz0_1;
	wire w_dff_B_iYYAhPtH2_1;
	wire w_dff_B_hJxebwXO2_1;
	wire w_dff_B_1rOe19vF7_1;
	wire w_dff_B_Flku22kH6_1;
	wire w_dff_B_d8xbczx92_1;
	wire w_dff_B_wtKDcpXr5_1;
	wire w_dff_B_jiHOXbbj5_1;
	wire w_dff_B_V6P9iNHF9_1;
	wire w_dff_B_MZbxAC849_1;
	wire w_dff_B_xNCmMBk97_1;
	wire w_dff_B_bvOcEYhx9_1;
	wire w_dff_B_Sba8qWKe1_1;
	wire w_dff_B_4zqwHMcn3_1;
	wire w_dff_B_89NlKiQx0_1;
	wire w_dff_A_Kz26MWjc3_0;
	wire w_dff_A_1pFUqW7z5_0;
	wire w_dff_A_ynV1tQbq2_0;
	wire w_dff_A_2p23fOaE8_0;
	wire w_dff_A_Ddh77EIo3_0;
	wire w_dff_A_uwHyYCaN4_0;
	wire w_dff_A_1TDUvT3S2_0;
	wire w_dff_A_qccnRTgA4_0;
	wire w_dff_A_jFumDGFP9_0;
	wire w_dff_A_DQgbQ5ou2_0;
	wire w_dff_A_HGepiMnx9_0;
	wire w_dff_A_Va2RIp0d2_0;
	wire w_dff_A_ZSVgJwjz6_0;
	wire w_dff_A_mSp6CN364_0;
	wire w_dff_A_4n7xRdXz6_0;
	wire w_dff_A_Hy90Dgah0_0;
	wire w_dff_A_2rnEDkGI8_0;
	wire w_dff_A_QzfuWymG6_0;
	wire w_dff_A_0QdGZfhF6_0;
	wire w_dff_A_8u3wyKNW2_0;
	wire w_dff_A_TTIOfwLJ6_0;
	wire w_dff_A_42VEkzUd0_0;
	wire w_dff_A_wmnia9FE7_0;
	wire w_dff_A_CT01YOIy2_0;
	wire w_dff_A_pm5yIr7C7_1;
	wire w_dff_A_wZnauLqZ3_1;
	wire w_dff_A_b2x55jkc4_1;
	wire w_dff_A_8FfXxIw29_1;
	wire w_dff_A_FDRDn6rK2_1;
	wire w_dff_A_oR8cAYML1_1;
	wire w_dff_A_hG1efiug5_1;
	wire w_dff_A_gQjEEydM9_1;
	wire w_dff_A_HHybKUxy7_1;
	wire w_dff_A_QXJHZhwo8_1;
	wire w_dff_A_pFKJmAwX6_1;
	wire w_dff_A_9a8RfQD82_1;
	wire w_dff_A_d3DqCKDa1_1;
	wire w_dff_A_8snGbMCi7_1;
	wire w_dff_A_1P8R3ZrU3_1;
	wire w_dff_A_0pCg8Ewb9_1;
	wire w_dff_A_45atGmSj6_1;
	wire w_dff_A_u41i3XLP8_1;
	wire w_dff_A_2upM7GSy5_1;
	wire w_dff_A_At8SYZXR9_1;
	wire w_dff_A_3acnhz7g5_1;
	wire w_dff_A_tHSp7MYp2_1;
	wire w_dff_A_53yDP0x22_1;
	wire w_dff_A_8p9Ep5ph6_1;
	wire w_dff_A_9rvIgHbL5_1;
	wire w_dff_A_kY51oWpU0_0;
	wire w_dff_B_HqIxwYqi2_1;
	wire w_dff_B_3QW2tG859_0;
	wire w_dff_B_O3ot9kj41_0;
	wire w_dff_B_03xtniDy3_0;
	wire w_dff_B_y9O1gk6A7_0;
	wire w_dff_B_yPoaqPFV1_0;
	wire w_dff_B_KqbWPMAA7_0;
	wire w_dff_B_1c3CAWR25_0;
	wire w_dff_B_w0GE4BjP7_0;
	wire w_dff_B_0r2lgX6Z4_0;
	wire w_dff_B_DuAUmMZp2_0;
	wire w_dff_B_HxY5XDOG6_0;
	wire w_dff_B_XqlUH8W71_0;
	wire w_dff_B_zWQ86AaD6_0;
	wire w_dff_B_CxBiZ04u6_0;
	wire w_dff_B_fapM1V6I5_0;
	wire w_dff_B_0HFPlUPS2_1;
	wire w_dff_B_qyrcYnYh3_1;
	wire w_dff_B_tA2cNRR86_1;
	wire w_dff_B_jfKWCVpc4_1;
	wire w_dff_B_OAVFaoik4_1;
	wire w_dff_B_3SVCqB2k5_1;
	wire w_dff_B_zSzYDKI31_1;
	wire w_dff_B_cvIotsGl6_1;
	wire w_dff_B_jkOunhVU9_1;
	wire w_dff_B_rbq2gHyU0_0;
	wire w_dff_B_cPSoNOer7_0;
	wire w_dff_B_G3VsxjGG6_0;
	wire w_dff_B_KrTOm0AB8_0;
	wire w_dff_B_3o3G4KE37_0;
	wire w_dff_B_gwqg9ZZ57_0;
	wire w_dff_B_LUT0e8DE8_0;
	wire w_dff_B_9yTnoITB3_0;
	wire w_dff_B_tpz87DSL5_1;
	wire w_dff_B_cLwlpkND2_1;
	wire w_dff_B_4u4Xii5w3_1;
	wire w_dff_B_eukirPuF1_0;
	wire w_dff_B_N2TiApL38_0;
	wire w_dff_B_5vmXC67r0_0;
	wire w_dff_B_GlwAPsGr3_0;
	wire w_dff_B_UpLf7Cvj0_1;
	wire w_dff_B_N3LKBBhK5_1;
	wire w_dff_B_SqTZABBO3_0;
	wire w_dff_B_geNj874Y9_1;
	wire w_dff_B_yVxRmE8s9_1;
	wire w_dff_B_lDAau8753_1;
	wire w_dff_B_SGJTEFsZ7_1;
	wire w_dff_B_c4nG2qid7_1;
	wire w_dff_B_nawDsiCY0_1;
	wire w_dff_B_wxIQ6v6t5_1;
	wire w_dff_B_sBac9MlJ7_1;
	wire w_dff_B_wflMoR4i4_0;
	wire w_dff_B_tJBu7D9I1_0;
	wire w_dff_B_qtNdDxOv6_0;
	wire w_dff_B_MtutydP07_0;
	wire w_dff_B_ZfoTuBf89_1;
	wire w_dff_B_MNVBHVb13_1;
	wire w_dff_B_QdTlWOPy6_1;
	wire w_dff_B_fq5VyQy93_1;
	wire w_dff_B_UR8JTR1B3_1;
	wire w_dff_A_ouZz7z5y9_1;
	wire w_dff_A_LEONILnR6_1;
	wire w_dff_A_iGsM9aDg2_1;
	wire w_dff_A_Jc0GopvY0_1;
	wire w_dff_A_N46omXvs3_1;
	wire w_dff_A_Ci7AUCfM4_0;
	wire w_dff_B_M7G7dGwZ6_1;
	wire w_dff_B_Z2wHRDtU8_1;
	wire w_dff_B_Mkgb4XIy6_1;
	wire w_dff_B_ggWbuOSW4_1;
	wire w_dff_B_PJlIltPn0_1;
	wire w_dff_B_2wUF6utT3_1;
	wire w_dff_A_kOmwN3a39_1;
	wire w_dff_A_HvaXIMe72_1;
	wire w_dff_A_Xh1K58Al4_1;
	wire w_dff_B_BkXH2J6l7_0;
	wire w_dff_B_yH6i9vbF7_0;
	wire w_dff_B_RLfVDbH87_0;
	wire w_dff_B_fmOTz5GE4_0;
	wire w_dff_B_Z5qrbyLp9_0;
	wire w_dff_B_QhpdVcFt4_0;
	wire w_dff_B_rPYqRfFP4_0;
	wire w_dff_B_HpupBuZ24_0;
	wire w_dff_A_VoEFyJdg8_0;
	wire w_dff_A_be0PVgZO0_0;
	wire w_dff_A_X0rfnNi28_1;
	wire w_dff_A_RStRHZ5r4_1;
	wire w_dff_B_WRO4cqmB1_0;
	wire w_dff_B_NZiGFut64_0;
	wire w_dff_B_CD8o9nVP1_0;
	wire w_dff_B_r1dpAwhO4_0;
	wire w_dff_B_dlwqYE0v5_0;
	wire w_dff_B_4gFb7LAe8_0;
	wire w_dff_B_rqk3hDLC2_0;
	wire w_dff_B_AJAqmFDh4_0;
	wire w_dff_B_QS0ZtmA05_0;
	wire w_dff_B_s0mZ4UlJ2_0;
	wire w_dff_B_1ETCG16F7_0;
	wire w_dff_B_CflVqS060_1;
	wire w_dff_B_0Sh2KuhN6_1;
	wire w_dff_B_IdX0IT347_1;
	wire w_dff_B_qWSCPjmn4_1;
	wire w_dff_B_iqyfaPSa7_1;
	wire w_dff_B_1Bg5NWFk1_0;
	wire w_dff_B_DMifZ2951_1;
	wire w_dff_B_R4fIqzS48_1;
	wire w_dff_B_t4O3bn2m0_1;
	wire w_dff_B_pMOYEzSd0_1;
	wire w_dff_B_H4wbGmLC0_1;
	wire w_dff_B_ECYdSkgf0_0;
	wire w_dff_A_xryQdEie7_1;
	wire w_dff_B_GRyt55l36_2;
	wire w_dff_B_uFvxpkhR8_2;
	wire w_dff_B_GGlOXZyL8_2;
	wire w_dff_A_gsJdNsID4_1;
	wire w_dff_A_hlvTrcX62_1;
	wire w_dff_A_reohEdbc8_0;
	wire w_dff_A_HgkOWHrE4_1;
	wire w_dff_A_XItf8W6e8_1;
	wire w_dff_A_0wblCObB8_1;
	wire w_dff_A_v1fpQzmh4_0;
	wire w_dff_B_6QtczEZz2_0;
	wire w_dff_B_MA6gwNRH6_0;
	wire w_dff_B_PjZIbyet8_0;
	wire w_dff_B_CPQM883m4_0;
	wire w_dff_A_MuEtCERx8_2;
	wire w_dff_A_vEisUAsu2_2;
	wire w_dff_A_CtVzTCe36_1;
	wire w_dff_B_nO6CwKfE5_1;
	wire w_dff_B_jlWztoAt0_1;
	wire w_dff_B_Ltzkq9aT6_1;
	wire w_dff_B_BzDzznrh5_1;
	wire w_dff_B_iBNBekbK7_1;
	wire w_dff_A_BCacFK5p1_0;
	wire w_dff_A_aXqDb7Dy9_0;
	wire w_dff_A_kO1rFbt35_1;
	wire w_dff_B_HbqcTied8_0;
	wire w_dff_B_Hlt852rt5_0;
	wire w_dff_B_v9TyYiHT8_0;
	wire w_dff_B_QigrX8J72_0;
	wire w_dff_B_sFDQ1TAz3_0;
	wire w_dff_B_5FHqcI0s9_0;
	wire w_dff_B_5DfRk7g22_0;
	wire w_dff_B_bd4qKzwn7_0;
	wire w_dff_B_6cZt0YIi7_1;
	wire w_dff_B_C05oqTQr5_1;
	wire w_dff_B_tybHPE6C0_0;
	wire w_dff_A_7QBH7DgZ4_2;
	wire w_dff_B_TASpClio3_2;
	wire w_dff_B_bujkl3Rf1_1;
	wire w_dff_B_woEMQmxf1_1;
	wire w_dff_B_7ZSJceom5_1;
	wire w_dff_B_nXJrMS4Q5_1;
	wire w_dff_B_3vBlmhip4_0;
	wire w_dff_A_PugzPvyA2_0;
	wire w_dff_A_sFVymup87_2;
	wire w_dff_A_goNGes1R7_1;
	wire w_dff_A_nTIZuExK6_1;
	wire w_dff_A_hMSCEz6U5_1;
	wire w_dff_A_F7LThMu61_1;
	wire w_dff_A_xJ1nBBsq8_2;
	wire w_dff_A_lbkfI0PV4_2;
	wire w_dff_A_ViR2xfxe9_2;
	wire w_dff_A_U84xEFrr8_2;
	wire w_dff_B_bTXCXE3W2_0;
	wire w_dff_A_0J4OVUoY9_1;
	wire w_dff_B_ivslArfX2_1;
	wire w_dff_B_2acrcGUW7_1;
	wire w_dff_B_1JNOJRPv9_1;
	wire w_dff_B_4bYsWbFL6_0;
	wire w_dff_B_60i9nVvj7_1;
	wire w_dff_B_M0D7D2sP4_0;
	wire w_dff_A_b3zYzCpI2_0;
	wire w_dff_A_1B2TbiEd3_0;
	wire w_dff_A_aEkXezqP0_0;
	wire w_dff_B_GkG2VC3M5_1;
	wire w_dff_B_z0hCELaH0_1;
	wire w_dff_B_FH0il0nK3_1;
	wire w_dff_B_oHTSJ5C89_1;
	wire w_dff_B_pK2sato87_1;
	wire w_dff_B_Bt9QAkTd5_1;
	wire w_dff_B_jDrwD3dI6_0;
	wire w_dff_B_JUvPulu93_0;
	wire w_dff_B_EVI7LtAT4_1;
	wire w_dff_B_1KlVEaGy7_1;
	wire w_dff_B_WMVZfwea1_1;
	wire w_dff_B_csNboiwg8_1;
	wire w_dff_B_uN3yNqMX3_1;
	wire w_dff_B_RgDzYCTb1_1;
	wire w_dff_A_5MRBFqNf2_1;
	wire w_dff_A_miPFumjC5_1;
	wire w_dff_A_vySj1KXD5_2;
	wire w_dff_A_h8BRsSgY3_2;
	wire w_dff_B_91mPsrla4_0;
	wire w_dff_B_HZLESQmS3_0;
	wire w_dff_B_iiAPVMOV7_0;
	wire w_dff_B_izibPMR73_0;
	wire w_dff_A_n3ud26WU8_1;
	wire w_dff_A_jYdxiSC18_1;
	wire w_dff_A_ejReBi1n1_2;
	wire w_dff_A_OgC83iMD6_2;
	wire w_dff_B_XA4MjNtg9_1;
	wire w_dff_B_MFdEChYk2_1;
	wire w_dff_B_BOKcaclG7_1;
	wire w_dff_B_5xXmWcjF8_0;
	wire w_dff_B_lMaU6M2E7_0;
	wire w_dff_B_ZDlQ6QMx7_0;
	wire w_dff_B_KGN0Cfxo1_0;
	wire w_dff_B_Nsxm4RzF0_0;
	wire w_dff_B_4csAsGzu2_0;
	wire w_dff_B_QDoeX3ui6_1;
	wire w_dff_B_6RDoPbTe0_1;
	wire w_dff_B_SfLpZ49O7_0;
	wire w_dff_A_yZq3Id2l3_0;
	wire w_dff_B_3TlZntCp2_1;
	wire w_dff_B_iHQo5wAi7_1;
	wire w_dff_B_MPZkSopX3_1;
	wire w_dff_B_jB04fN5o7_1;
	wire w_dff_B_pKX3Z6ci2_1;
	wire w_dff_B_41U9DHKJ6_1;
	wire w_dff_B_9KRSL5N54_1;
	wire w_dff_B_VokvmHoW1_1;
	wire w_dff_B_XDbCX56u3_1;
	wire w_dff_B_o7ogLalW2_1;
	wire w_dff_B_60dAyajg5_1;
	wire w_dff_B_aLyvrF5y2_1;
	wire w_dff_B_E3kh8RIO8_1;
	wire w_dff_B_icDZmfxm3_1;
	wire w_dff_B_JiIMEmpI1_0;
	wire w_dff_A_CPktjDSG5_2;
	wire w_dff_A_qp1sAGMq6_0;
	wire w_dff_A_4qe0AaBu3_0;
	wire w_dff_A_G158mUnH8_0;
	wire w_dff_A_LdP0sqej6_0;
	wire w_dff_B_IhUb9nu18_0;
	wire w_dff_B_jj7AxzEY2_0;
	wire w_dff_A_R9T0BBH90_0;
	wire w_dff_B_CaZgp0CW2_0;
	wire w_dff_B_xcyXUC0e7_0;
	wire w_dff_B_pBuz2pDf9_0;
	wire w_dff_B_SVihhk5e3_0;
	wire w_dff_B_anfcVjYq8_0;
	wire w_dff_B_7vlzAMVs7_1;
	wire w_dff_B_Wtje1SaE7_1;
	wire w_dff_B_8U9rPPQx0_1;
	wire w_dff_B_7KrCzawj1_1;
	wire w_dff_B_BFovSasJ9_1;
	wire w_dff_A_3K811a2e5_1;
	wire w_dff_A_oOUnMqgv3_1;
	wire w_dff_B_vF6pt99o2_1;
	wire w_dff_B_WnKyF0ti2_1;
	wire w_dff_B_AyWMX6dN8_1;
	wire w_dff_B_FFFNZjvU1_1;
	wire w_dff_B_gz7dj8DM7_1;
	wire w_dff_A_dueqaJgq7_0;
	wire w_dff_A_OzKVJmt60_1;
	wire w_dff_A_0n0CCISK2_1;
	wire w_dff_A_gRyxMBcX9_1;
	wire w_dff_A_wrgjO4ru4_2;
	wire w_dff_A_BL9huDU75_2;
	wire w_dff_A_iqe8B1jB8_2;
	wire w_dff_A_64ftG2JB1_2;
	wire w_dff_A_z0DziQVH6_1;
	wire w_dff_B_jijveFSS1_0;
	wire w_dff_A_lGm10NeH2_0;
	wire w_dff_A_Cfx5oZ4z1_0;
	wire w_dff_A_KnaJJwVi3_2;
	wire w_dff_A_ul9kiYTC7_2;
	wire w_dff_B_RxDJlPs49_1;
	wire w_dff_B_SfGEYDQO1_1;
	wire w_dff_B_imB7NkY34_0;
	wire w_dff_B_TYKlVe3n2_0;
	wire w_dff_A_P2HetoOa5_1;
	wire w_dff_A_oerN6jKl5_2;
	wire w_dff_B_r4P1rwqF3_1;
	wire w_dff_B_umOvivqc3_0;
	wire w_dff_A_ySobaZ7d0_0;
	wire w_dff_A_4xonIQ2c6_1;
	wire w_dff_A_VOB1MuIG0_1;
	wire w_dff_B_3YAnUPyw5_1;
	wire w_dff_B_CwgtMlEH9_1;
	wire w_dff_A_auWLdSP48_0;
	wire w_dff_A_MMhFJs1l8_0;
	wire w_dff_A_Ci1lgWHE0_0;
	wire w_dff_A_NyrFAQ7A8_0;
	wire w_dff_A_7zXK7Z0j7_0;
	wire w_dff_A_b1O6bxue3_1;
	wire w_dff_B_QKGI8h3V0_0;
	wire w_dff_B_pKNYMOUG6_0;
	wire w_dff_B_llGLiG5a1_2;
	wire w_dff_B_e8e0s9Tw7_2;
	wire w_dff_A_gNDVYk1S1_0;
	wire w_dff_A_OexgeZbJ0_0;
	wire w_dff_A_wHFAAAM29_0;
	wire w_dff_B_r7I87ypp4_0;
	wire w_dff_B_XBhVLbD39_0;
	wire w_dff_B_scrVZ7927_0;
	wire w_dff_B_AqESJkoR8_0;
	wire w_dff_B_T07KtoY26_1;
	wire w_dff_B_t9fHK07t4_1;
	wire w_dff_B_A4QDMoH20_2;
	wire w_dff_B_vwMSbg3t9_1;
	wire w_dff_B_z7x30knv6_1;
	wire w_dff_B_9Ye4cWSA9_0;
	wire w_dff_A_twfCMpHp6_1;
	wire w_dff_A_FoTsNkAw5_1;
	wire w_dff_A_jxubB8fU3_1;
	wire w_dff_A_lRwSU2RU9_2;
	wire w_dff_A_bd3qanCL6_2;
	wire w_dff_A_cwbGpK2Z3_2;
	wire w_dff_B_82kYTqqJ9_1;
	wire w_dff_B_h10GtyIo3_1;
	wire w_dff_B_EJ1B3EeP0_1;
	wire w_dff_B_hSFoL9Vx7_1;
	wire w_dff_B_JttXkiGp9_1;
	wire w_dff_B_XCGnxZHc1_1;
	wire w_dff_B_hLJtlJJF9_0;
	wire w_dff_B_gkg3k09p5_1;
	wire w_dff_B_Gc1DhZXX9_1;
	wire w_dff_B_ItcZGkKB8_0;
	wire w_dff_A_XwDnaQlt8_0;
	wire w_dff_B_LMCkRrVG6_3;
	wire w_dff_B_H1HY01fP6_3;
	wire w_dff_B_ZmiO3i2x6_3;
	wire w_dff_A_v49lq3ym8_0;
	wire w_dff_B_Spb4oRM94_2;
	wire w_dff_B_iymQpDhf8_2;
	wire w_dff_B_iGSNmT5R3_2;
	wire w_dff_B_nxT6o9XU7_0;
	wire w_dff_B_NKXEqKka3_1;
	wire w_dff_B_8uaxFcVp8_1;
	wire w_dff_B_n5lwAc6J4_1;
	wire w_dff_B_fa6AkwhY3_1;
	wire w_dff_A_UIxmzBzU1_1;
	wire w_dff_A_REiphj4s6_1;
	wire w_dff_A_Dg7xY4Fv9_1;
	wire w_dff_A_PuunYYEp3_2;
	wire w_dff_A_qFR6XBNy6_2;
	wire w_dff_B_csnaLUaJ0_1;
	wire w_dff_B_SEmiHP4u7_0;
	wire w_dff_A_81pCt3ZJ1_0;
	wire w_dff_B_wNpOitCb0_3;
	wire w_dff_B_GH2siCI67_3;
	wire w_dff_B_rX8Nivot9_3;
	wire w_dff_A_eVb0pw6a8_1;
	wire w_dff_A_izTLcR693_1;
	wire w_dff_A_1HXeJx3I1_1;
	wire w_dff_A_ItvJ0AUZ0_1;
	wire w_dff_A_4pTrGx9u1_1;
	wire w_dff_A_Xcd62Tim0_1;
	wire w_dff_A_kV4MqbCa6_1;
	wire w_dff_A_pftuPXJG7_1;
	wire w_dff_A_ujHVhFXE2_0;
	wire w_dff_A_Ag613vyg4_0;
	wire w_dff_A_dg8jophn1_0;
	wire w_dff_A_uHQJX5Vw1_0;
	wire w_dff_A_vPuHMoXa2_0;
	wire w_dff_A_eoNa2PPz0_0;
	wire w_dff_A_PmPtq17c4_0;
	wire w_dff_A_6nzvRsWK0_0;
	wire w_dff_A_Qi2CfUyN8_0;
	wire w_dff_A_Kdl1A3t00_0;
	wire w_dff_A_A0bUwg7l5_0;
	wire w_dff_A_ylJrylbW4_2;
	wire w_dff_A_LaKsi5FD4_2;
	wire w_dff_A_KivU3g2Y0_2;
	wire w_dff_A_J1tWehzc5_2;
	wire w_dff_A_T1KNWnat5_2;
	wire w_dff_A_iJjgRdQp3_2;
	wire w_dff_A_ji8CAmEm2_2;
	wire w_dff_A_LszETj6i5_2;
	wire w_dff_A_CfZyoAll3_2;
	wire w_dff_A_9vAQujb96_2;
	wire w_dff_A_W5fxPdRt2_2;
	wire w_dff_A_Ben8Znh69_1;
	wire w_dff_A_g596W5QG4_1;
	wire w_dff_A_EkXCf4t16_1;
	wire w_dff_A_OBzN97CG2_1;
	wire w_dff_A_Ziy1fTaz3_1;
	wire w_dff_A_Rh16nUJt7_1;
	wire w_dff_A_ogfxIjFq3_1;
	wire w_dff_A_V9S1PCU52_1;
	wire w_dff_A_utYsbCW66_1;
	wire w_dff_A_VPWo4PEw8_1;
	wire w_dff_A_yUSiJE2a0_1;
	wire w_dff_A_S8IxAVDR1_2;
	wire w_dff_A_LXrKOMXU9_2;
	wire w_dff_A_sa20jRqe0_2;
	wire w_dff_A_y1zRS86h4_2;
	wire w_dff_A_S2S9Tqky1_2;
	wire w_dff_A_vvbmvctz9_2;
	wire w_dff_A_pOHd292y6_2;
	wire w_dff_A_FpweQpZM3_2;
	wire w_dff_A_zH2JcY4f7_2;
	wire w_dff_A_MFZomLcF0_2;
	wire w_dff_A_YCIlTHLf2_2;
	wire w_dff_B_h5FG6BeU4_0;
	wire w_dff_B_ISAkrs8o5_0;
	wire w_dff_B_CUucMEAh7_0;
	wire w_dff_B_hy5ZWvia2_0;
	wire w_dff_B_CqHJVKye5_0;
	wire w_dff_A_iUfvIEz78_0;
	wire w_dff_A_7vTYN9o84_0;
	wire w_dff_A_afHYqFxH2_1;
	wire w_dff_A_zsQunHwU7_1;
	wire w_dff_A_Dp2CALI72_1;
	wire w_dff_A_AWNgwUnV3_2;
	wire w_dff_A_CCeIWJGa4_2;
	wire w_dff_A_AQIsk6hs2_2;
	wire w_dff_B_nMMtbWXq2_2;
	wire w_dff_B_US2VQ0nN2_2;
	wire w_dff_B_j0ovojQ30_2;
	wire w_dff_B_6rRYUcVr6_2;
	wire w_dff_B_jQEs3KYQ8_2;
	wire w_dff_B_UkCu8P9U7_2;
	wire w_dff_B_X6l0t1JA9_2;
	wire w_dff_B_kEvGkueG5_2;
	wire w_dff_B_5RQQ68ig4_2;
	wire w_dff_B_NutjzFEL9_2;
	wire w_dff_B_rCqzEXuV5_2;
	wire w_dff_B_thoodCAy6_2;
	wire w_dff_B_S2SNhrZX6_2;
	wire w_dff_A_hTgHDsrK5_1;
	wire w_dff_B_LDRONa5J9_0;
	wire w_dff_B_8uFYQU0E4_0;
	wire w_dff_B_k2RQ2kjo3_0;
	wire w_dff_B_beaLWjaP9_0;
	wire w_dff_B_bg2628tI6_0;
	wire w_dff_B_1sI4oKiB0_0;
	wire w_dff_B_XgRgISjX1_0;
	wire w_dff_B_VuOjOOvv5_0;
	wire w_dff_B_Lq59G3kr3_0;
	wire w_dff_B_mnHUxTSm7_0;
	wire w_dff_B_jzkxmxX52_0;
	wire w_dff_B_kddCkst46_1;
	wire w_dff_B_ORN9O6023_1;
	wire w_dff_B_5yDNasKG3_1;
	wire w_dff_B_GuNW2e8p9_1;
	wire w_dff_A_4YM7diBN0_1;
	wire w_dff_A_byatC4aG6_1;
	wire w_dff_A_hHFRDDwG8_2;
	wire w_dff_A_JY0B51aq6_1;
	wire w_dff_A_LJCRtSSc7_1;
	wire w_dff_A_2wjzWZAY2_1;
	wire w_dff_A_E9E5rxLQ7_1;
	wire w_dff_A_WqWUz2897_2;
	wire w_dff_A_WoNmbVIo1_2;
	wire w_dff_A_hCTVNgxW4_2;
	wire w_dff_A_UPue7mKt7_2;
	wire w_dff_A_VPKwfkVC7_1;
	wire w_dff_A_JH9MCF8f4_0;
	wire w_dff_A_BxsKgBGG5_0;
	wire w_dff_A_BhkLDNvD8_0;
	wire w_dff_A_xk3kCVKM2_0;
	wire w_dff_A_ynk5dqSb2_2;
	wire w_dff_A_Ku9B3Y2T2_2;
	wire w_dff_A_ZBccMnZ21_2;
	wire w_dff_A_iBOwVAhb4_1;
	wire w_dff_B_nx93J3LY3_1;
	wire w_dff_B_YnLdvlym2_1;
	wire w_dff_B_ui9JvqB01_1;
	wire w_dff_B_07FqMLME8_0;
	wire w_dff_A_dNdWUtir8_1;
	wire w_dff_A_HGXab7lh5_2;
	wire w_dff_A_3k1m8a2A3_0;
	wire w_dff_B_9LjZadz51_3;
	wire w_dff_B_V6JONzVg6_3;
	wire w_dff_B_Nv8zABFN6_3;
	wire w_dff_B_GdT3MNyE9_1;
	wire w_dff_B_LpNfrY359_0;
	wire w_dff_A_iO2LrXBq8_0;
	wire w_dff_A_SLH6Xzgr1_1;
	wire w_dff_A_60JJg4zp8_1;
	wire w_dff_A_jRhn2qcD5_1;
	wire w_dff_A_ti8Wxqyt9_1;
	wire w_dff_A_6ZpunHw50_1;
	wire w_dff_A_tDWTM7ME4_1;
	wire w_dff_A_iA6ky1Cq2_1;
	wire w_dff_A_D22jo48r6_1;
	wire w_dff_A_rkOouUbH5_2;
	wire w_dff_A_CfidJJKC8_2;
	wire w_dff_B_TULLagoq1_0;
	wire w_dff_B_cPx4GLvs2_0;
	wire w_dff_B_f1Dh1Z274_0;
	wire w_dff_B_sc5ECryo4_0;
	wire w_dff_A_IUdNnhry2_0;
	wire w_dff_B_KM6fBycT4_0;
	wire w_dff_B_QrDDYXQC2_0;
	wire w_dff_B_Knx9thml1_0;
	wire w_dff_B_uZqli6Na3_0;
	wire w_dff_B_wPggN8AG0_0;
	wire w_dff_A_6HEAOcvv8_2;
	wire w_dff_A_wkG5dVVG0_1;
	wire w_dff_A_I4QRRSBC3_1;
	wire w_dff_A_gAq1C1p84_2;
	wire w_dff_A_RqxBxNm63_2;
	wire w_dff_A_Tgsmx2AP1_0;
	wire w_dff_A_2gKLDoFq8_1;
	wire w_dff_A_Jq6HlDRh1_1;
	wire w_dff_A_xygUTBYQ0_1;
	wire w_dff_A_KWWvRnfy9_1;
	wire w_dff_B_kRL33Kwb6_1;
	wire w_dff_B_X5McmxHP1_1;
	wire w_dff_A_Ql0JBR2b8_1;
	wire w_dff_B_tzQ4OxgE2_1;
	wire w_dff_B_IkMZBkBp9_0;
	wire w_dff_B_6AA9bqyU6_0;
	wire w_dff_B_kQIUHOkP2_0;
	wire w_dff_B_DmEc0be85_1;
	wire w_dff_A_yZBgr7T34_0;
	wire w_dff_A_i2cl3Bp49_0;
	wire w_dff_B_rUgMDvnS7_1;
	wire w_dff_B_wq0pYMBx5_1;
	wire w_dff_A_pmyIkI1G1_0;
	wire w_dff_A_E2BCCOSl0_0;
	wire w_dff_B_eHtuai9V9_0;
	wire w_dff_B_DaWjeVjL0_1;
	wire w_dff_B_bgCGocnM4_1;
	wire w_dff_B_nwC5A8HM1_1;
	wire w_dff_B_g2sFFUCp9_1;
	wire w_dff_B_ZlgEJhOi6_0;
	wire w_dff_B_4GyJWtJN6_0;
	wire w_dff_B_pwH9jyPc2_1;
	wire w_dff_B_GXNaKhtp0_1;
	wire w_dff_B_KQl9HTF33_1;
	wire w_dff_A_Rva1AEKD2_1;
	wire w_dff_A_fcI5NC2f2_1;
	wire w_dff_B_OqO96hog7_1;
	wire w_dff_B_sob5fowR5_1;
	wire w_dff_A_DfSwjIls9_0;
	wire w_dff_A_GcD66brr2_0;
	wire w_dff_A_Hl1mrqai0_0;
	wire w_dff_A_sYv13dku0_0;
	wire w_dff_B_QXqYkzoH9_0;
	wire w_dff_A_Y1zkbMin2_1;
	wire w_dff_A_VGVZ5Om46_1;
	wire w_dff_A_bdTsspxu3_2;
	wire w_dff_A_0wvv5lHZ5_2;
	wire w_dff_A_7l3Pgq8W7_2;
	wire w_dff_A_Aw8GGBk42_2;
	wire w_dff_B_O8CWMqll9_1;
	wire w_dff_B_p1GlhHg72_1;
	wire w_dff_B_6p6SfMK66_1;
	wire w_dff_A_NVMS29z04_0;
	wire w_dff_B_aFDTMb6B2_2;
	wire w_dff_A_iZRRhRrA3_1;
	wire w_dff_A_mjNH1ppj0_1;
	wire w_dff_A_f4ZUCAnr5_1;
	wire w_dff_B_iyPl7ZmR6_2;
	wire w_dff_B_KYm3OC3V3_2;
	wire w_dff_B_MDlhKS9x1_1;
	wire w_dff_B_okKJV17k9_1;
	wire w_dff_B_fXFLWVgQ2_1;
	wire w_dff_B_sKt8HdsP3_0;
	wire w_dff_B_BmUIe2270_0;
	wire w_dff_A_se3X5d4g7_2;
	wire w_dff_B_Sggb8bRB2_1;
	wire w_dff_B_j1vmASJy6_1;
	wire w_dff_B_1IiMTn0s3_1;
	wire w_dff_A_UtVkimCc4_1;
	wire w_dff_A_R3DlfM8k2_1;
	wire w_dff_A_Zz5ApCGF9_1;
	wire w_dff_A_wbXxIzL69_2;
	wire w_dff_A_UhyvKCbr2_2;
	wire w_dff_A_ZMc46jzT5_2;
	wire w_dff_A_efmkBkH97_2;
	wire w_dff_A_k7Tm4JLD1_1;
	wire w_dff_A_NQWsafb08_1;
	wire w_dff_A_Q7OJ38FA2_1;
	wire w_dff_A_6lOqnehS9_2;
	wire w_dff_A_j7xJR0ii1_2;
	wire w_dff_A_T3yNR4nP6_0;
	wire w_dff_A_cOaJiuwx8_0;
	wire w_dff_A_tYBCD6H65_2;
	wire w_dff_A_jZYY5mXL9_2;
	wire w_dff_A_qGQbUysa8_2;
	wire w_dff_A_Bkc40ouF1_2;
	wire w_dff_A_MDo3JADq1_1;
	wire w_dff_A_kd626oGo4_1;
	wire w_dff_A_wySSWbT54_1;
	wire w_dff_A_pOseXtjT4_0;
	wire w_dff_A_ErXiBYYZ2_0;
	wire w_dff_A_cR9FzrOM6_1;
	wire w_dff_A_B5q9nHKd8_0;
	wire w_dff_A_9fkugbRV3_2;
	wire w_dff_A_ALYf8q0U3_2;
	wire w_dff_A_FhmdJnKA2_2;
	wire w_dff_A_T6Lcc6IH2_2;
	wire w_dff_A_X1hUSW124_0;
	wire w_dff_A_ogpRhe583_0;
	wire w_dff_A_3yl5nL2Z1_0;
	wire w_dff_A_lSMlxxfa2_0;
	wire w_dff_B_JFbHVnB53_0;
	wire w_dff_B_vGkxd8xS3_0;
	wire w_dff_B_r4LG1yPQ1_0;
	wire w_dff_B_xLr7nSLd4_0;
	wire w_dff_B_QhMunovb1_0;
	wire w_dff_B_5HwZXw286_0;
	wire w_dff_B_8PHEd5ke3_0;
	wire w_dff_B_HgA4b9FY1_0;
	wire w_dff_B_Ppn9qytr3_0;
	wire w_dff_A_pBq5s4Ky8_2;
	wire w_dff_A_LWd1eegR5_2;
	wire w_dff_A_qpMqPPcq4_2;
	wire w_dff_A_TgSkigYm6_2;
	wire w_dff_A_U1yV6sTq2_2;
	wire w_dff_A_cxDIl5xZ8_2;
	wire w_dff_A_ae2eSZrV7_2;
	wire w_dff_A_tv0YYWOD6_2;
	wire w_dff_A_QIOLY1di5_0;
	wire w_dff_A_Js16njrf8_0;
	wire w_dff_A_WyZX4gsb9_0;
	wire w_dff_A_7dGQOBZh0_0;
	wire w_dff_B_nCPTWesU8_1;
	wire w_dff_B_FVLNdNhN9_1;
	wire w_dff_B_DDUVIJFg5_1;
	wire w_dff_B_oi0MVyjt8_1;
	wire w_dff_B_BzC8fKGl8_1;
	wire w_dff_B_ipLwlcnj3_0;
	wire w_dff_A_hARDuVkP8_0;
	wire w_dff_A_QcckcgpA9_0;
	wire w_dff_A_zRY7bSLT2_0;
	wire w_dff_A_a7FNnu3y0_0;
	wire w_dff_A_FTZodH591_2;
	wire w_dff_A_xytoGJ765_2;
	wire w_dff_A_K9gIku7k7_0;
	wire w_dff_A_zKMlK3M14_2;
	wire w_dff_A_TeDTVq7P5_2;
	wire w_dff_B_1L2my1Ce8_1;
	wire w_dff_B_bHxLWWnm0_0;
	wire w_dff_A_PdTwVXbF9_1;
	wire w_dff_B_lMcfsCfC6_3;
	wire w_dff_B_a15zM2mw9_3;
	wire w_dff_B_VxTUBMna6_3;
	wire w_dff_B_XrhrrlvU0_1;
	wire w_dff_B_TVNJnW056_1;
	wire w_dff_B_r2gcMh6c5_1;
	wire w_dff_B_jVLjZUPy4_1;
	wire w_dff_A_7umLYpXk7_1;
	wire w_dff_A_jxYs8qcu1_1;
	wire w_dff_A_A7uLTU6D5_1;
	wire w_dff_A_RZGU9K3y6_2;
	wire w_dff_A_QAexC1sc5_2;
	wire w_dff_A_fg08Ldde0_1;
	wire w_dff_B_3B131pBc4_3;
	wire w_dff_B_QIrx4NMT7_3;
	wire w_dff_B_ob9irtai4_3;
	wire w_dff_B_1aarbTzk5_3;
	wire w_dff_B_bPHmTA1B5_3;
	wire w_dff_B_OJom1FYt1_3;
	wire w_dff_A_1jvSdNCV3_0;
	wire w_dff_A_qnf9fads5_1;
	wire w_dff_A_a7wtfoCu3_1;
	wire w_dff_A_Tu0gHDuX6_0;
	wire w_dff_A_NYxeNxQl8_0;
	wire w_dff_A_cIHiKiZJ6_1;
	wire w_dff_B_10MjFtWH4_3;
	wire w_dff_B_FaIakyj15_3;
	wire w_dff_A_S6zJZXWQ4_1;
	wire w_dff_A_5WXIHceh4_1;
	wire w_dff_A_voKTqiQL6_1;
	wire w_dff_A_xVhRKMLI4_1;
	wire w_dff_A_bXRGpFUT9_1;
	wire w_dff_A_ZQoEcb4V4_2;
	wire w_dff_A_1O6QwAK35_2;
	wire w_dff_A_voqPKDHg0_2;
	wire w_dff_A_qJaP0EbY2_2;
	wire w_dff_A_ZwW0hqYD3_2;
	wire w_dff_A_Y6d7z2k86_0;
	wire w_dff_A_VSlrG3Dt9_0;
	wire w_dff_A_q4g8PyAu0_0;
	wire w_dff_A_Lcjr7Jkd0_2;
	wire w_dff_A_PQWol2Sk5_2;
	wire w_dff_A_E87Knj2C7_2;
	wire w_dff_A_0z4pOVe93_2;
	wire w_dff_A_E8BBP3RC2_1;
	wire w_dff_A_YDRcNMc83_1;
	wire w_dff_A_YtGq8GRF4_1;
	wire w_dff_A_t519heTb5_0;
	wire w_dff_A_pQn8Bwgt4_0;
	wire w_dff_A_sftDko8u2_0;
	wire w_dff_A_c0tZk3tN5_0;
	wire w_dff_A_UIfhTpSR6_1;
	wire w_dff_A_Os20HUNC9_1;
	wire w_dff_A_nE77gkUE2_1;
	wire w_dff_A_kTjxzvWT2_1;
	wire w_dff_A_BgoFfZ3G5_1;
	wire w_dff_B_YOTbRa345_1;
	wire w_dff_B_VXotR1C14_0;
	wire w_dff_A_sZBHAwzC5_0;
	wire w_dff_A_OjuoUKn81_0;
	wire w_dff_A_6kKoFWxY3_0;
	wire w_dff_A_6QzVYnv16_0;
	wire w_dff_A_WpFUIipS7_0;
	wire w_dff_A_XapG0G1E1_0;
	wire w_dff_A_k8AR201x1_1;
	wire w_dff_A_hjzNrcIA2_1;
	wire w_dff_A_3IWXGl4Q0_1;
	wire w_dff_A_B9U87A7P4_0;
	wire w_dff_A_8HWxLwAr6_1;
	wire w_dff_A_jajZH1VY4_1;
	wire w_dff_A_cgO3RsdM6_1;
	wire w_dff_A_jgi2bvqi1_1;
	wire w_dff_A_NrGcdwvs9_1;
	wire w_dff_A_rbiAdqSD1_1;
	wire w_dff_A_Bv9YZrCL5_1;
	wire w_dff_A_SVEJQEdk3_1;
	wire w_dff_A_ockTjTGj2_1;
	wire w_dff_A_j1AoV3UV3_2;
	wire w_dff_A_PsH6dYKB1_2;
	wire w_dff_A_NNb2mDc57_2;
	wire w_dff_A_LEOZPeAq6_2;
	wire w_dff_A_RLuNULWX6_2;
	wire w_dff_A_hnkDfjQ26_2;
	wire w_dff_A_cCghVtay5_2;
	wire w_dff_A_4V9nTFmm2_0;
	wire w_dff_A_BmjXFYCM9_0;
	wire w_dff_A_zyh5SjHl5_1;
	wire w_dff_A_SoJMaa6U8_1;
	wire w_dff_A_UqmQbHpi3_1;
	wire w_dff_B_hcZHqHtM7_3;
	wire w_dff_B_pBdD8D9U3_3;
	wire w_dff_B_ZMOIlzt87_3;
	wire w_dff_A_rz8ZnS6y4_0;
	wire w_dff_A_3WnZy8Of3_0;
	wire w_dff_A_EqDyQK220_0;
	wire w_dff_A_XyPl7Lk52_0;
	wire w_dff_A_qpkrdL6F0_0;
	wire w_dff_A_aJLsqmqe2_0;
	wire w_dff_A_2IN7JSSE6_0;
	wire w_dff_A_milrLsVw7_0;
	wire w_dff_A_eDV0uxhS1_0;
	wire w_dff_A_94mwUmcO2_2;
	wire w_dff_A_0IwzuOTi7_2;
	wire w_dff_A_Isvsff5S9_2;
	wire w_dff_A_cxIVGy278_2;
	wire w_dff_A_PltvLy5v7_2;
	wire w_dff_A_bLHjKvDv5_2;
	wire w_dff_A_YfFfKuRT3_2;
	wire w_dff_A_ZCgrvjX68_2;
	wire w_dff_A_DNgoaVjB0_2;
	wire w_dff_A_AleqX0qi5_1;
	wire w_dff_A_0ODAtrUi0_1;
	wire w_dff_A_ILahda5L6_1;
	wire w_dff_A_x1atrqor5_1;
	wire w_dff_A_PoO6PUAm4_1;
	wire w_dff_A_MXYQ7IB02_1;
	wire w_dff_A_KIRTliAh7_1;
	wire w_dff_A_YM0Ge1Vw3_1;
	wire w_dff_A_QQY4p0rR0_1;
	wire w_dff_A_euVF13K51_1;
	wire w_dff_A_krnNoCNg3_1;
	wire w_dff_A_lUaj8Hsi0_1;
	wire w_dff_A_pmUtW7ki4_1;
	wire w_dff_A_ZyVloKti1_2;
	wire w_dff_A_6HQUVwQJ4_2;
	wire w_dff_A_fnaKOyxR0_2;
	wire w_dff_A_EAZ32BHi9_2;
	wire w_dff_A_bK1TnP9p4_2;
	wire w_dff_A_7hze8iR17_2;
	wire w_dff_A_qCgzmTEy5_0;
	wire w_dff_A_hmWkYl082_0;
	wire w_dff_A_ke3cuQ8i2_0;
	wire w_dff_A_oQQHS6Mo0_0;
	wire w_dff_A_3o3Aga818_0;
	wire w_dff_A_4PtGJqYM5_0;
	wire w_dff_A_S6x8R5Mw2_0;
	wire w_dff_A_Gn1AnE2P9_0;
	wire w_dff_A_pbjlvNlT9_0;
	wire w_dff_A_J6QaOLpY5_0;
	wire w_dff_A_it7GQ7Dp9_0;
	wire w_dff_A_Y9PeBElv4_0;
	wire w_dff_A_8ee8hWvj7_0;
	wire w_dff_A_eDriXEU77_1;
	wire w_dff_A_vbppFX2z4_1;
	wire w_dff_A_r9m11Sp88_1;
	wire w_dff_A_S2lH40NS3_1;
	wire w_dff_A_hwFI4iZB9_1;
	wire w_dff_A_lNkq2tnW6_1;
	wire w_dff_A_17g9O5Q45_1;
	wire w_dff_A_BHDPSEJu9_1;
	wire w_dff_A_es2IyWpY0_1;
	wire w_dff_A_e1hrWvYU6_1;
	wire w_dff_A_VZd0gpUa7_1;
	wire w_dff_A_epIckd794_1;
	wire w_dff_A_rmQ2P6ob1_1;
	wire w_dff_A_4rI3Hm1b7_1;
	wire w_dff_A_JcjRvWF04_1;
	wire w_dff_A_Sk17eZjh8_1;
	wire w_dff_A_Z5GJ55JZ7_1;
	wire w_dff_A_Jlmq51Zr9_1;
	wire w_dff_A_y4ktkX414_1;
	wire w_dff_A_zP91gkby3_1;
	wire w_dff_A_gn9FCwl94_1;
	wire w_dff_A_EU8P0IAU4_1;
	wire w_dff_A_Z7lBfSnI7_1;
	wire w_dff_A_vyM2sOR99_1;
	wire w_dff_A_Br01DCnm4_1;
	wire w_dff_A_fSXR1oKu2_1;
	wire w_dff_A_fqyNz2KY1_2;
	wire w_dff_A_eD5IR1Xa5_2;
	wire w_dff_A_nTNjntaC7_2;
	wire w_dff_A_1QqJ9wCN0_2;
	wire w_dff_A_cwOhX6n43_2;
	wire w_dff_A_BRkAedmK3_2;
	wire w_dff_A_oSt0Z7Fn2_2;
	wire w_dff_A_GaKWSEUJ3_2;
	wire w_dff_A_6jzFGnfY0_2;
	wire w_dff_A_lxyL6k5x6_2;
	wire w_dff_A_5WFaK1hc7_2;
	wire w_dff_A_0qz3eAIP3_2;
	wire w_dff_A_qItjlHxo7_2;
	wire w_dff_A_2Lxs9L7N3_0;
	wire w_dff_A_teYQVboa8_0;
	wire w_dff_A_h56ZK11V3_0;
	wire w_dff_A_6yVyZMe51_0;
	wire w_dff_A_FrwTlVFw6_1;
	wire w_dff_A_GjQKIh0o2_1;
	wire w_dff_B_sOUDt0Jw2_0;
	wire w_dff_A_sEsirQ287_0;
	wire w_dff_A_tjhWdLt39_0;
	wire w_dff_A_wb8Hnplw2_2;
	wire w_dff_A_jEUckHfx1_2;
	wire w_dff_A_bOcYBU0u4_2;
	wire w_dff_A_ho90xERe3_2;
	wire w_dff_A_XAQQnvFH0_2;
	wire w_dff_A_5l6bkAPs5_2;
	wire w_dff_A_LBbokkSq4_2;
	wire w_dff_A_4flnU5zK4_2;
	wire w_dff_A_zv0BLC0m7_0;
	wire w_dff_A_foqsK1iu2_0;
	wire w_dff_A_b2z0fmQw0_2;
	wire w_dff_A_K3AGBwzM7_2;
	wire w_dff_A_Qm3iBtMs3_0;
	wire w_dff_A_Bqe3jeLH4_0;
	wire w_dff_A_oKToOtMw2_0;
	wire w_dff_A_rE5M3qzY2_0;
	wire w_dff_A_BtVjkjIy1_0;
	wire w_dff_A_VkJ1vD6E1_0;
	wire w_dff_A_qcHqbGIZ2_0;
	wire w_dff_A_XgjECKGW1_0;
	wire w_dff_A_NfkWhLiY8_0;
	wire w_dff_A_J59My1ut6_0;
	wire w_dff_A_Cc4Z5JpJ0_0;
	wire w_dff_A_OHnnts5a2_0;
	wire w_dff_A_cnEcAlP81_0;
	wire w_dff_A_5VOD5gPl1_0;
	wire w_dff_A_uUFNsoGC3_0;
	wire w_dff_A_q04vrTA72_0;
	wire w_dff_A_6sHJM5Xy7_0;
	wire w_dff_A_0Vx3tG7G7_0;
	wire w_dff_A_Dpu2HDyE5_0;
	wire w_dff_A_RVW5JvzM4_0;
	wire w_dff_A_nRPaJcOi2_0;
	wire w_dff_A_38n0BuBO0_0;
	wire w_dff_A_5EtYuR3P8_0;
	wire w_dff_A_2Z8Vb7209_0;
	wire w_dff_A_WuP3LnJy6_0;
	wire w_dff_A_gLushfnS0_2;
	wire w_dff_A_EkWjSkVG5_2;
	wire w_dff_A_0FM0OZMY3_2;
	wire w_dff_A_2ztTpdvS4_2;
	wire w_dff_A_ABqeBcBg4_2;
	wire w_dff_A_o4yGNFE28_2;
	wire w_dff_A_3vwKYx7W8_2;
	wire w_dff_A_e5zBkha42_2;
	wire w_dff_A_PXx4x6xd0_2;
	wire w_dff_A_hJFt0JUq5_2;
	wire w_dff_A_NOqUuvhp9_2;
	wire w_dff_A_oK4zSfYn4_2;
	wire w_dff_A_v2epItUz6_2;
	wire w_dff_A_efDEuNxq6_0;
	wire w_dff_A_SbLLWM3N7_0;
	wire w_dff_A_tBKkmNvp4_0;
	wire w_dff_A_y3PO73Gt2_0;
	wire w_dff_A_otLYebaF9_0;
	wire w_dff_A_jUt24f707_0;
	wire w_dff_A_7wzqqj0K4_0;
	wire w_dff_A_g7s5hUKJ2_0;
	wire w_dff_A_HF26pmmT6_0;
	wire w_dff_A_KIjRKvEF8_0;
	wire w_dff_A_BR7yUBq60_0;
	wire w_dff_A_Msh28AIK4_0;
	wire w_dff_A_4H3XaxPj6_0;
	wire w_dff_A_VeR9ydHJ0_0;
	wire w_dff_A_DYaQg0vp6_0;
	wire w_dff_A_Tlt9Iy7U2_0;
	wire w_dff_A_4dWGbo2M2_0;
	wire w_dff_A_uVqKDdK71_0;
	wire w_dff_A_NIIAfPAZ6_0;
	wire w_dff_A_FtjmGpGm0_0;
	wire w_dff_A_u6fPMMaP3_0;
	wire w_dff_A_FVLSn8r61_0;
	wire w_dff_A_QFC8lswS0_0;
	wire w_dff_A_dbpOmaep7_0;
	wire w_dff_A_7yC2WvL09_0;
	wire w_dff_A_NKSqx6L97_0;
	wire w_dff_A_h4aSon9b3_0;
	wire w_dff_A_26u5r4nr6_0;
	wire w_dff_A_KUQs97An9_0;
	wire w_dff_A_sgipNb9P9_0;
	wire w_dff_A_wb61tip46_2;
	wire w_dff_A_eAITEikv4_2;
	wire w_dff_A_JILv7yJU2_2;
	wire w_dff_A_lyF7RBDh0_2;
	wire w_dff_A_FIvS8d8q9_2;
	wire w_dff_A_M10eiDHh9_2;
	wire w_dff_A_lNKpBkY69_2;
	wire w_dff_A_wNh1CPYe6_2;
	wire w_dff_A_eWsVhYOj0_2;
	wire w_dff_A_Ex1egs7k1_2;
	wire w_dff_A_e4fD6PVS9_2;
	wire w_dff_A_wbSx4lJH0_2;
	wire w_dff_A_Kfs7AARq6_2;
	wire w_dff_A_RDXHd6ax8_2;
	wire w_dff_A_PLUdXRwP9_2;
	wire w_dff_A_u2zHD1e91_2;
	wire w_dff_A_n6nBEFBo6_1;
	wire w_dff_A_E5pJEshh8_1;
	wire w_dff_A_MLM49nvu0_1;
	wire w_dff_A_KAKvmEud6_1;
	wire w_dff_A_UmJBnRF14_1;
	wire w_dff_A_q1cvYpYO2_1;
	wire w_dff_A_9hmZZOMP7_1;
	wire w_dff_A_T3VMcTWS5_1;
	wire w_dff_A_0DJNY8V99_1;
	wire w_dff_A_0di6ejzZ1_1;
	wire w_dff_A_Q6Dq8Ah13_1;
	wire w_dff_A_RXvEj56w3_1;
	wire w_dff_A_tHQQdhbh2_1;
	wire w_dff_A_cMUk0oNq2_1;
	wire w_dff_A_6R3kS48e5_1;
	wire w_dff_A_c5SsrmG99_2;
	wire w_dff_A_EAFlgYlb7_2;
	wire w_dff_A_ZwSopGnD6_2;
	wire w_dff_A_8r5WNWsq5_2;
	wire w_dff_A_SRQIDQ7D6_2;
	wire w_dff_A_XIXWfR327_2;
	wire w_dff_A_lItuLGzC4_2;
	wire w_dff_A_ZzE4B1hQ3_2;
	wire w_dff_A_RzWSvsP64_2;
	wire w_dff_A_8t7XT2I58_2;
	wire w_dff_A_Wyu1IZHA3_2;
	wire w_dff_A_zCFOVLXZ8_2;
	wire w_dff_A_kgQl7vYj7_2;
	wire w_dff_A_oIS23WKq9_2;
	wire w_dff_A_tOxrVneJ3_2;
	wire w_dff_A_Et3t0F1f3_2;
	wire w_dff_A_byAoXEJY4_0;
	wire w_dff_B_jnmeR2JH2_1;
	wire w_dff_A_y0drUesM0_0;
	wire w_dff_A_oKWf7lUA3_2;
	wire w_dff_A_GMUR2CPS4_1;
	wire w_dff_A_z8LJpB2h8_1;
	wire w_dff_B_z3m5Avw11_2;
	wire w_dff_B_5I69Vif71_1;
	wire w_dff_B_2IrSLCfN1_1;
	wire w_dff_A_3lsDjhPM0_1;
	wire w_dff_A_zACDLaCd8_1;
	wire w_dff_A_H7rNPwfV6_1;
	wire w_dff_A_KERD0IRv4_1;
	wire w_dff_A_YzTLrI8s4_1;
	wire w_dff_A_UHbBUwz78_1;
	wire w_dff_A_a4r3djru3_2;
	wire w_dff_A_qexzSkda6_1;
	wire w_dff_B_BY0d8Vvj8_1;
	wire w_dff_B_RrKfitDe2_1;
	wire w_dff_B_blmEti2I9_1;
	wire w_dff_B_5UrRsifg7_1;
	wire w_dff_B_SftRxwdb3_0;
	wire w_dff_B_7bGxVacK4_0;
	wire w_dff_A_f247w4bX7_1;
	wire w_dff_A_ZekLadoH4_1;
	wire w_dff_A_Tuc3xxEz9_1;
	wire w_dff_A_452Wf0t57_2;
	wire w_dff_A_b1BQvMIP9_2;
	wire w_dff_B_FlaDmVrW3_0;
	wire w_dff_A_Evo67m0p9_0;
	wire w_dff_A_BXlryQIW5_0;
	wire w_dff_A_fZIAVK5L5_1;
	wire w_dff_A_iUA9Ib5T0_1;
	wire w_dff_A_2N6qgzwC1_0;
	wire w_dff_A_12RyQrOQ0_1;
	wire w_dff_A_iBXOt02u3_0;
	wire w_dff_A_m5tUA2gX7_2;
	wire w_dff_A_4h93hrzN3_2;
	wire w_dff_A_1oddAwu36_2;
	wire w_dff_A_m1kh582q3_2;
	wire w_dff_A_O5xTzMGe8_1;
	wire w_dff_A_u587GSUF0_2;
	wire w_dff_A_y5BjkwQk8_2;
	wire w_dff_A_5GiiMNAY6_2;
	wire w_dff_A_oNKs1aL00_1;
	wire w_dff_A_MSnj6Roc5_2;
	wire w_dff_A_oDxiCE6K5_2;
	wire w_dff_B_ncTjER867_2;
	wire w_dff_B_UiuHreiG2_2;
	wire w_dff_A_Q0cECAjb6_0;
	wire w_dff_A_heQ81J368_0;
	wire w_dff_A_AlW9APjx6_0;
	wire w_dff_A_AzYgYmxN5_0;
	wire w_dff_A_4R66MgMk3_1;
	wire w_dff_A_YzT3lXEH0_1;
	wire w_dff_A_dRsxdNdo2_1;
	wire w_dff_A_3XLrzspX8_1;
	wire w_dff_A_OYmyEwU07_1;
	wire w_dff_A_Xyt08d892_1;
	wire w_dff_B_5oDl5aKy0_1;
	wire w_dff_A_0p8q4oEL4_0;
	wire w_dff_A_rPI04wTs3_0;
	wire w_dff_A_4JHMJTxp3_1;
	wire w_dff_A_EOEzw3Vb1_1;
	wire w_dff_A_AYPTE2zr5_1;
	wire w_dff_A_z1MRiI3L0_1;
	wire w_dff_A_zfeHizBJ6_1;
	wire w_dff_A_hwWaFAFZ0_2;
	wire w_dff_A_CC0y3FIr4_2;
	wire w_dff_B_8wZLjwLq1_0;
	wire w_dff_A_freTjB7M9_1;
	wire w_dff_B_tmtaSXRO8_1;
	wire w_dff_A_sJNSF0Ru5_1;
	wire w_dff_A_ZsxRKSK08_0;
	wire w_dff_A_m4ejHiAa8_2;
	wire w_dff_A_NeBlkTsm6_2;
	wire w_dff_B_ShiCuMxf1_0;
	wire w_dff_B_LVfRVNFb1_1;
	wire w_dff_B_1acgoLbH7_1;
	wire w_dff_A_xefzw0Xr8_1;
	wire w_dff_A_WS3oRN2k1_2;
	wire w_dff_A_7SSjdnDc8_2;
	wire w_dff_A_xiYrl7Po4_2;
	wire w_dff_A_4vEzungA6_2;
	wire w_dff_A_jQrP0qoc7_2;
	wire w_dff_A_OPmw6A1f2_0;
	wire w_dff_A_FsF9GHw87_0;
	wire w_dff_A_LEHBkyB51_0;
	wire w_dff_A_VFWpqNBh3_1;
	wire w_dff_A_hKnFbtoY1_1;
	wire w_dff_B_yf8mo9is2_3;
	wire w_dff_B_msZ2tOuf0_3;
	wire w_dff_A_enXX1quV3_0;
	wire w_dff_A_jqIH72iD9_0;
	wire w_dff_A_GOOIVse66_0;
	wire w_dff_A_NLwXJCfA3_0;
	wire w_dff_A_f6ABZmXF8_0;
	wire w_dff_A_jEYlmuyq8_0;
	wire w_dff_A_4pgYoo2E4_0;
	wire w_dff_A_VI4Ow6M03_0;
	wire w_dff_A_aiaFnVaD1_0;
	wire w_dff_A_HI4z6a6C1_0;
	wire w_dff_A_9HLKkSpm3_0;
	wire w_dff_A_91jmAvar1_0;
	wire w_dff_A_gGprMvpd8_0;
	wire w_dff_A_VRV9qAWt3_0;
	wire w_dff_A_UZPuOWI86_0;
	wire w_dff_A_4aWkU8mK7_0;
	wire w_dff_A_lu5uwDg92_0;
	wire w_dff_A_KoQiKot56_0;
	wire w_dff_A_UWsNxs513_0;
	wire w_dff_A_kz12i0ey7_0;
	wire w_dff_A_9D9xGHVi8_0;
	wire w_dff_A_KgJyM3XM4_0;
	wire w_dff_A_iIEJL7x26_1;
	wire w_dff_A_cdQ8lvh06_1;
	wire w_dff_A_OwvypD2H7_1;
	wire w_dff_A_14bn1H3V2_1;
	wire w_dff_A_H6Iufzoy3_1;
	wire w_dff_A_NxuSkR1F8_0;
	wire w_dff_A_qXdsbkWq8_0;
	wire w_dff_A_lkOogajD3_0;
	wire w_dff_A_6ibv6KxW6_0;
	wire w_dff_A_0ooMxjBe8_2;
	wire w_dff_A_WfffUTBY0_2;
	wire w_dff_A_QXkNSAJn4_2;
	wire w_dff_A_5qQQlvTO6_2;
	wire w_dff_A_5IqAVncz2_2;
	wire w_dff_A_MFGIaPWm2_2;
	wire w_dff_A_bK8Nu5iM8_1;
	wire w_dff_A_7LcNbOki3_1;
	wire w_dff_A_fpDwdSui3_1;
	wire w_dff_A_H37i0v2h2_1;
	wire w_dff_A_yC9TF1hH3_1;
	wire w_dff_A_PIWTNxa47_1;
	wire w_dff_A_l6eqF4jg5_1;
	wire w_dff_A_Nt9qYN4z2_2;
	wire w_dff_A_RWubiC2U0_2;
	wire w_dff_A_7yhEceqI7_2;
	wire w_dff_A_w3NQBbIP8_2;
	wire w_dff_A_m20jSWco6_2;
	wire w_dff_A_pcLx0mV21_2;
	wire w_dff_A_Q5eaKtoA0_2;
	wire w_dff_A_7xrzCvZ98_0;
	wire w_dff_A_WHdKEeti2_2;
	wire w_dff_A_xfuiYykq1_0;
	wire w_dff_A_jXlgNbp25_0;
	wire w_dff_A_k8cXiJ2y9_1;
	wire w_dff_A_xBHXsD235_1;
	wire w_dff_A_7HMNrkS60_1;
	wire w_dff_A_9ajb0Fgk1_1;
	wire w_dff_A_hfgBgHRV7_1;
	wire w_dff_A_L3eaQgWY6_1;
	wire w_dff_A_4BPmvvzp9_1;
	wire w_dff_A_dyn12HjZ2_1;
	wire w_dff_A_HyiWPJhq6_1;
	wire w_dff_A_m10HyTs41_1;
	wire w_dff_A_XXE2nEhX0_1;
	wire w_dff_A_ptdNnmc79_1;
	wire w_dff_A_Q8B1EI8U6_1;
	wire w_dff_A_28R9RAxr3_1;
	wire w_dff_A_ppYdNBXJ7_1;
	wire w_dff_A_8yOL4Dgw9_1;
	wire w_dff_A_oRsplpzq6_1;
	wire w_dff_A_mvZgpjTa2_1;
	wire w_dff_A_vPeGR7Cb2_1;
	wire w_dff_B_M01Athst6_0;
	wire w_dff_B_hX57umbd8_1;
	wire w_dff_B_AzoIUIvS6_1;
	wire w_dff_A_PBSqfgil2_0;
	wire w_dff_A_cYysVxzc5_0;
	wire w_dff_A_RiNEh80W2_0;
	wire w_dff_A_jOo9fuYz8_0;
	wire w_dff_A_Imtw7rXu0_0;
	wire w_dff_A_h4Q5cbvG7_0;
	wire w_dff_A_cZDb5ZWs9_0;
	wire w_dff_A_eCBS0RGn4_0;
	wire w_dff_A_pBjB8zcm8_0;
	wire w_dff_A_CcQV7sao7_1;
	wire w_dff_A_907yCrwn3_1;
	wire w_dff_A_5gty9tSV0_1;
	wire w_dff_A_jKKD54u20_0;
	wire w_dff_A_g5QmKHKA5_1;
	wire w_dff_B_0hyWijOB1_0;
	wire w_dff_A_8lUREGvv9_0;
	wire w_dff_A_X9o9EagP8_0;
	wire w_dff_B_YJgMbXiN0_0;
	wire w_dff_A_rDKXslHr0_0;
	wire w_dff_A_gTv3yu3c8_1;
	wire w_dff_B_8oMyJe3n5_0;
	wire w_dff_B_dx20306R1_1;
	wire w_dff_A_IdEcDTYM4_1;
	wire w_dff_A_25vdNoTz2_1;
	wire w_dff_A_xs3jEeia8_1;
	wire w_dff_A_K1vDXWvX4_1;
	wire w_dff_A_VN3q0wQ22_1;
	wire w_dff_A_Eg5R2SEy7_1;
	wire w_dff_A_qZwwkgyD6_1;
	wire w_dff_A_xEzVN75u1_2;
	wire w_dff_A_xg4r9KJb0_2;
	wire w_dff_A_IZgxIELf9_2;
	wire w_dff_A_VD87RK157_2;
	wire w_dff_A_V41USIAe6_2;
	wire w_dff_A_Hrh71dSF0_2;
	wire w_dff_A_LDnZStKM2_2;
	wire w_dff_B_eIoYXnst0_0;
	wire w_dff_B_HPMsywrA8_1;
	wire w_dff_A_gxRNkctz1_1;
	wire w_dff_B_f909SO4t3_1;
	wire w_dff_A_V7oCZJGo4_0;
	wire w_dff_A_i4efet1B6_0;
	wire w_dff_A_5OOqrkCz7_0;
	wire w_dff_A_xED5Ylry2_1;
	wire w_dff_A_FmN24kVt6_1;
	wire w_dff_A_szOXg0XM3_1;
	wire w_dff_A_k4uqZuK57_2;
	wire w_dff_A_mEmlEm6s2_1;
	wire w_dff_A_pg5ld5f74_2;
	wire w_dff_A_3GIROOwX0_1;
	wire w_dff_A_Vd13r1yy1_1;
	wire w_dff_A_kigN5drF4_0;
	wire w_dff_A_Mcvi3e8f7_0;
	wire w_dff_A_NoZTrR2V0_1;
	wire w_dff_A_p17GX4UV7_1;
	wire w_dff_A_n0VUd9i96_0;
	wire w_dff_A_sWlRsFGD9_2;
	wire w_dff_A_K9aNkitx6_0;
	wire w_dff_A_diXvnU778_0;
	wire w_dff_A_Y2GmgOsp7_0;
	wire w_dff_A_ytftHHj82_2;
	wire w_dff_A_Y4JxR3WW4_2;
	wire w_dff_A_m5Q5lf740_2;
	wire w_dff_A_aA3KFQK93_0;
	wire w_dff_A_sEnV04eU0_1;
	wire w_dff_A_OnhiM6jf3_1;
	wire w_dff_A_QxyDXSi28_1;
	wire w_dff_A_fSTzQJGM8_1;
	wire w_dff_A_vs3ZJwGa9_1;
	wire w_dff_A_F4dMoCGY8_0;
	wire w_dff_A_JAB0NABu1_0;
	wire w_dff_A_YTISlkpo1_0;
	wire w_dff_A_j389pyct4_1;
	wire w_dff_A_yhiv0qnJ2_1;
	wire w_dff_A_RpaMBR3p5_1;
	wire w_dff_A_8jcRzIF35_0;
	wire w_dff_A_0kfJlfHL3_0;
	wire w_dff_A_myBV1axo5_0;
	wire w_dff_A_gzwjnW8H8_0;
	wire w_dff_B_Mur7JrsD8_1;
	wire w_dff_A_4cmS3fqh7_1;
	wire w_dff_A_BA5H7OT31_1;
	wire w_dff_A_xrb7684A8_0;
	wire w_dff_A_vkj7UK126_0;
	wire w_dff_A_FRSK5cPf6_0;
	wire w_dff_A_buMYHT8l8_1;
	wire w_dff_A_qesgmJmZ7_1;
	wire w_dff_A_CIgBAP6t9_1;
	wire w_dff_A_HEpS09PU5_1;
	wire w_dff_A_OO5hki6w7_0;
	wire w_dff_A_IgAXfZzA0_0;
	wire w_dff_A_Q36Cbjon5_0;
	wire w_dff_A_ud7KC6Dr5_2;
	wire w_dff_A_KoVECPo00_2;
	wire w_dff_A_DVvo8ZCm3_2;
	wire w_dff_A_phx9anFf7_2;
	wire w_dff_A_kYlrdnQQ1_1;
	wire w_dff_A_tYn1OjxC8_1;
	wire w_dff_A_WHrdW1Ds3_1;
	wire w_dff_A_4UQrobXj6_1;
	wire w_dff_A_22UFqUHs9_2;
	wire w_dff_A_wQqteubQ1_2;
	wire w_dff_B_QdJvX37F8_1;
	wire w_dff_A_OOS4yCBy7_1;
	wire w_dff_A_ep0BYdZp7_0;
	wire w_dff_B_b3AJGpTB4_2;
	wire w_dff_A_oB7QLt3h5_0;
	wire w_dff_A_7vqWpU2b0_0;
	wire w_dff_A_8lZq8ZH51_0;
	wire w_dff_A_iYKKcq6s5_0;
	wire w_dff_A_epM4ApjK4_1;
	wire w_dff_A_d6qjtnqe1_0;
	wire w_dff_A_sE9iFuPG8_0;
	wire w_dff_A_jhqvHvKy5_0;
	wire w_dff_A_RA3arEWY5_1;
	wire w_dff_B_wMQgszaN9_0;
	wire w_dff_B_rjK55iLY6_1;
	wire w_dff_A_XQVY9OJj8_0;
	wire w_dff_A_WKwum4yB3_0;
	wire w_dff_A_Fhdl4g5f6_0;
	wire w_dff_A_kStMTVvA0_0;
	wire w_dff_A_0eUypARF3_1;
	wire w_dff_A_zKYKHmZ62_0;
	wire w_dff_A_dL83xHsC3_0;
	wire w_dff_A_dReq60Ge5_2;
	wire w_dff_A_LoneYxIj4_2;
	wire w_dff_A_EIUmMT0j9_2;
	wire w_dff_A_hxoan87X8_2;
	wire w_dff_B_ZpafX9QN3_2;
	wire w_dff_B_Vq8gzTDt7_2;
	wire w_dff_A_k9xFSACD7_0;
	wire w_dff_A_EPeBne8a8_0;
	wire w_dff_A_pLaXYgni3_0;
	wire w_dff_A_PVD5866S1_0;
	wire w_dff_A_rkCxOl9m8_0;
	wire w_dff_A_diV3Ue6L8_0;
	wire w_dff_A_SYSv08G87_0;
	wire w_dff_B_Pfjezq0K0_1;
	wire w_dff_B_Lh5p2nfy2_1;
	wire w_dff_A_l2Iq00g77_0;
	wire w_dff_A_Veso47nX9_0;
	wire w_dff_A_q6XlzzcL2_0;
	wire w_dff_A_WKO8z8L31_1;
	wire w_dff_A_puhMWKVZ2_1;
	wire w_dff_A_Pd07LdMc2_0;
	wire w_dff_A_E9VK3GGi0_0;
	wire w_dff_A_dERL1esi8_0;
	wire w_dff_A_4xdXvQ5i9_1;
	wire w_dff_A_Nj1xB4c89_0;
	wire w_dff_A_Zk9P2qZg2_0;
	wire w_dff_A_b8kFfbc09_0;
	wire w_dff_A_gflqMBrW2_0;
	wire w_dff_A_gmoFzwOH9_1;
	wire w_dff_A_S3Ofe1LR7_1;
	wire w_dff_A_ancPBdLJ4_1;
	wire w_dff_A_edXna7eJ5_2;
	wire w_dff_A_7iP5EJLw6_2;
	wire w_dff_A_LxrKDjch3_1;
	wire w_dff_A_ohRw46K36_0;
	wire w_dff_A_3JjXdUhZ0_0;
	wire w_dff_A_NhpZJ60q4_1;
	wire w_dff_A_DwDP3ax58_1;
	wire w_dff_A_a661qqWF4_0;
	wire w_dff_A_gin0FYtn7_0;
	wire w_dff_A_vm3CoLng7_0;
	wire w_dff_A_nop1cqlb2_1;
	wire w_dff_A_qi5N4hBn9_1;
	wire w_dff_A_JHrJ7IEG6_1;
	wire w_dff_A_e8sfntoC4_1;
	wire w_dff_A_NdYvpb6L3_0;
	wire w_dff_A_Ky48hNU60_0;
	wire w_dff_A_OrDQkYHF2_0;
	wire w_dff_A_Rq2WqyD75_1;
	wire w_dff_A_WgHVasRv6_1;
	wire w_dff_A_BEM9gBeJ0_1;
	wire w_dff_A_vdMaJsxe1_2;
	wire w_dff_B_JFQs6Cz90_1;
	wire w_dff_A_myor13xe4_0;
	wire w_dff_A_0xjxALv33_0;
	wire w_dff_A_Cqq1PXCx8_0;
	wire w_dff_A_fMhCZthv7_0;
	wire w_dff_A_tHjXO9qn9_0;
	wire w_dff_A_w7jeGZ1o2_0;
	wire w_dff_A_04AmFTHf6_0;
	wire w_dff_A_dvjVEWxA4_1;
	wire w_dff_A_Vj3zXUSD7_2;
	wire w_dff_A_zEvWIwJo2_2;
	wire w_dff_A_S5qBGsov9_2;
	wire w_dff_A_DvuEtOEI0_2;
	wire w_dff_A_AC7C3EdM4_2;
	wire w_dff_A_zNAJmdNo3_2;
	wire w_dff_A_tSw5gpj66_2;
	wire w_dff_A_h3hOAETZ3_0;
	wire w_dff_A_eTefsioD9_0;
	wire w_dff_A_NYW3Xivn3_0;
	wire w_dff_A_vTaEXAVh6_0;
	wire w_dff_A_lU4zRC4C0_0;
	wire w_dff_A_KmYiWHCA8_0;
	wire w_dff_A_gp0OvPEx3_0;
	wire w_dff_A_KuEorIls1_1;
	wire w_dff_A_1pNUcVq28_1;
	wire w_dff_A_8WEsy4756_1;
	wire w_dff_A_aeTsSMyu8_1;
	wire w_dff_A_t2h3zT050_1;
	wire w_dff_A_D5ioe1ut3_0;
	wire w_dff_A_UiqxvAbc6_0;
	wire w_dff_B_XO0IhvhS0_2;
	wire w_dff_A_OaCuvt4G3_0;
	wire w_dff_A_zh0VzruW5_2;
	wire w_dff_A_iEPVGXbc1_1;
	wire w_dff_A_AFPinfUT7_0;
	wire w_dff_A_6560CfKM2_1;
	wire w_dff_A_r7UpT6j45_0;
	wire w_dff_A_jYX9ILcw5_2;
	wire w_dff_B_2j51IpD02_3;
	wire w_dff_B_6ZjQg0y14_3;
	wire w_dff_B_0K4ozC484_3;
	wire w_dff_B_Kx6Og7Dy1_3;
	wire w_dff_B_3i5XDcRf5_3;
	wire w_dff_A_SdzZ5niv9_0;
	wire w_dff_A_Op3Y7Qyk3_0;
	wire w_dff_A_6Bh61tbJ4_0;
	wire w_dff_A_zBWmPbHG3_0;
	wire w_dff_A_Y1JWnzVp6_0;
	wire w_dff_A_qFpA9wC00_0;
	wire w_dff_A_0Cd7dMhP4_0;
	wire w_dff_A_tEBnN8hb4_1;
	wire w_dff_A_Q9Jvy1F31_1;
	wire w_dff_A_BvBckVrT2_1;
	wire w_dff_A_ZPJlTqa26_1;
	wire w_dff_A_svGUg6Zs8_1;
	wire w_dff_A_PDTYNlM86_1;
	wire w_dff_A_hueIkzjX5_1;
	wire w_dff_A_7goX015T1_0;
	wire w_dff_A_ztx9r2Kk8_0;
	wire w_dff_A_8lMDIxq95_0;
	wire w_dff_A_VZusJvtW5_0;
	wire w_dff_A_LLg45RjN1_0;
	wire w_dff_A_dPZsFRWr1_0;
	wire w_dff_A_9SVGVaCc9_0;
	wire w_dff_B_ZzgSafiw8_0;
	wire w_dff_A_JQXtkOfm4_1;
	wire w_dff_A_jlBU6s221_0;
	wire w_dff_A_3zB2eNgH8_0;
	wire w_dff_A_lQeOl7ID9_2;
	wire w_dff_A_bCeVzPG46_0;
	wire w_dff_A_ySZaPlsh8_0;
	wire w_dff_A_vaFRwjF51_2;
	wire w_dff_A_LwmgBJME5_2;
	wire w_dff_A_9SLDHbAe5_2;
	wire w_dff_A_migydITg8_2;
	wire w_dff_A_W57appsB7_0;
	wire w_dff_A_rvJlGxMM5_1;
	wire w_dff_A_J1r9uf2M9_1;
	wire w_dff_A_hmRUict03_1;
	wire w_dff_A_aqb3i7Wl7_1;
	wire w_dff_A_HHjywFP82_2;
	wire w_dff_A_Zb3xwYVa1_2;
	wire w_dff_A_fba0B7RA2_2;
	wire w_dff_A_0WhyBnTx4_2;
	wire w_dff_A_zOTSQUUw9_2;
	wire w_dff_A_xy0sGcsL6_2;
	wire w_dff_A_vPPBpKop8_2;
	wire w_dff_A_mELiXizb9_2;
	wire w_dff_A_I8vtH30z0_1;
	wire w_dff_A_UNJo7RyV4_1;
	wire w_dff_A_zpj0968i2_1;
	wire w_dff_A_8g564uFz5_2;
	wire w_dff_A_yvp6lg1U7_2;
	wire w_dff_A_41vnu8CB0_2;
	wire w_dff_A_FyrA18Hj7_0;
	wire w_dff_A_RA2zgpyC4_0;
	wire w_dff_A_KAbfLiU74_0;
	wire w_dff_A_LCf4WESU9_1;
	wire w_dff_A_627OoBlb1_0;
	wire w_dff_A_kurh59Sd5_0;
	wire w_dff_A_eX8x4eDb8_2;
	wire w_dff_A_0bJBcDI72_2;
	wire w_dff_A_8CcwNKW05_2;
	wire w_dff_A_qyr4YAAL0_0;
	wire w_dff_A_4NSeATNu0_0;
	wire w_dff_A_wlDyDHq85_0;
	wire w_dff_A_Rx4qNfI10_1;
	wire w_dff_A_B5O5RWX09_1;
	wire w_dff_A_0ZObVAKv4_2;
	wire w_dff_A_STJGStVK6_2;
	wire w_dff_A_fdHaWDMG5_2;
	wire w_dff_A_3ugz4ekH2_1;
	wire w_dff_A_GckQdKlQ9_0;
	wire w_dff_A_bpt5RxmD3_1;
	wire w_dff_A_gPbxcvWN4_0;
	wire w_dff_A_cdRuprlC3_2;
	wire w_dff_A_Aan9hUfF7_2;
	wire w_dff_A_9F1ay21P3_2;
	wire w_dff_A_RNnn8wkf2_2;
	wire w_dff_A_iHywy3nW6_2;
	wire w_dff_A_xLbWa16Q8_1;
	wire w_dff_A_H1BMiCLW6_0;
	wire w_dff_A_a8iaffyV9_2;
	wire w_dff_A_PrKjblqV4_0;
	wire w_dff_B_5J6oeO852_2;
	wire w_dff_B_EMpldElG0_2;
	wire w_dff_A_iE1iT1Y11_0;
	wire w_dff_A_ZAgSLwp21_0;
	wire w_dff_A_VSsmvDUq1_0;
	wire w_dff_A_3PEqnBcy6_2;
	wire w_dff_A_NM1O3RPj3_2;
	wire w_dff_A_CVpa9cST4_2;
	wire w_dff_A_UPHWAMW62_2;
	wire w_dff_A_TknSeaS27_1;
	wire w_dff_A_VQWbXmd77_1;
	wire w_dff_A_LbIR4ecf3_1;
	wire w_dff_A_UERcl1tV7_2;
	wire w_dff_A_g5BCQ1hB0_0;
	wire w_dff_A_UJGM8GXu6_1;
	wire w_dff_A_5F5KU4zg0_0;
	wire w_dff_B_WNMm4euq5_0;
	wire w_dff_A_glHElJOj6_0;
	wire w_dff_A_1pW9fGce3_0;
	wire w_dff_A_h6y2HzJO2_0;
	wire w_dff_A_BVbQtBU74_2;
	wire w_dff_A_IZ76Ei1m6_2;
	wire w_dff_A_4s0TyoYc9_0;
	wire w_dff_B_HqtnbwdP0_0;
	wire w_dff_A_E0S8gfdK9_2;
	wire w_dff_A_wjUr3Scq4_0;
	wire w_dff_A_ZwyCD0fH4_1;
	wire w_dff_A_1pje1mkK3_0;
	wire w_dff_A_vUIlcnRK2_2;
	wire w_dff_A_T6R9xgvp5_2;
	wire w_dff_A_JyxtuiHL2_2;
	wire w_dff_A_a8nK50Vz3_0;
	wire w_dff_A_6srOqm5Z0_0;
	wire w_dff_A_js40K4Sf9_1;
	wire w_dff_A_jMjaoHUR0_1;
	wire w_dff_A_dXhCYzvS6_1;
	wire w_dff_A_LKBQMA7Q4_1;
	wire w_dff_A_VuZYIoto5_2;
	wire w_dff_A_QYvsE2TM0_2;
	wire w_dff_A_zXJtZd5W5_2;
	wire w_dff_A_BhSiJ9au1_0;
	wire w_dff_A_Kgb8rgQL7_1;
	wire w_dff_A_QsEFNNHz1_0;
	wire w_dff_A_g1sQxtI67_0;
	wire w_dff_A_HHFWPCEd1_1;
	wire w_dff_A_Pf8WR8ke6_1;
	wire w_dff_B_rwCQmGns8_1;
	wire w_dff_A_XmqvYvIZ1_0;
	wire w_dff_A_0vFtVP2w7_0;
	wire w_dff_A_tiDUSUyz2_2;
	wire w_dff_A_wPVodFzS2_2;
	wire w_dff_A_m9AQBAfc0_1;
	wire w_dff_A_yrtdOxd48_1;
	wire w_dff_A_NaGJkzdY8_1;
	wire w_dff_A_VMQDtKWt8_2;
	wire w_dff_A_wIbuJ4LX4_2;
	wire w_dff_A_kEIBVVPy7_2;
	wire w_dff_A_WYs0vfay0_1;
	wire w_dff_A_nPtrMTIV5_1;
	wire w_dff_A_xBne4DBd4_1;
	wire w_dff_A_ck8EZlDh9_2;
	wire w_dff_A_kOAxi8ve7_0;
	wire w_dff_A_lN1JJFlD5_0;
	wire w_dff_A_k6eV8qlH9_1;
	wire w_dff_A_nxMrEFUv2_1;
	wire w_dff_A_cHbsuxtE2_1;
	wire w_dff_A_ygpYplsT6_1;
	wire w_dff_A_QvNaOfpl1_2;
	wire w_dff_A_71vYR1RX5_2;
	wire w_dff_A_Cc3xYaea6_2;
	wire w_dff_A_DghhoA0d2_0;
	wire w_dff_A_z9ZgqKo90_0;
	wire w_dff_A_pyR7l0nS8_1;
	wire w_dff_A_UaOFlXuZ9_1;
	wire w_dff_A_vFYBr6sJ7_1;
	wire w_dff_A_xklEYXbG0_1;
	wire w_dff_A_AXuFwqn41_2;
	wire w_dff_A_ppap3l3i7_2;
	wire w_dff_A_RXzNqvLP6_2;
	wire w_dff_A_YpwrCHtT1_2;
	wire w_dff_A_0uRYzCfa2_1;
	wire w_dff_A_3G10Qk7Z1_1;
	wire w_dff_A_iWfDf8LR3_2;
	wire w_dff_A_MFQzdhd58_2;
	wire w_dff_A_Dp18gep98_1;
	wire w_dff_A_HThULbC84_1;
	wire w_dff_A_F456LDT18_0;
	wire w_dff_A_Wo6mhXIz9_1;
	wire w_dff_A_RKU5LgTY8_2;
	wire w_dff_A_EE6LrMLh2_2;
	wire w_dff_A_3Vq1cj8a2_2;
	wire w_dff_A_aYuOSGG61_2;
	wire w_dff_A_1sYSLJKw4_2;
	wire w_dff_A_euNSTRCr8_2;
	wire w_dff_A_GKmywLFy8_2;
	wire w_dff_A_6zatj6M01_0;
	wire w_dff_A_7tAftBDu2_1;
	wire w_dff_A_9AnwOYgO0_2;
	wire w_dff_A_pi8XySmV6_1;
	wire w_dff_A_EsjesbNK5_2;
	wire w_dff_A_DlJf6hDJ7_2;
	wire w_dff_A_X0OT3Diz9_0;
	wire w_dff_A_X0OpRtEZ5_2;
	wire w_dff_A_pjgwWpzJ1_0;
	wire w_dff_A_3ji1y7E47_1;
	wire w_dff_A_SvNwvbPR2_1;
	wire w_dff_A_9d0Oyzz15_1;
	wire w_dff_A_jB4hXWJ21_1;
	wire w_dff_A_TYEQOXSd2_1;
	wire w_dff_A_nLw5oAua9_1;
	wire w_dff_A_N37N5do51_2;
	wire w_dff_A_YnphOlLj9_2;
	wire w_dff_A_iOPizZua7_2;
	wire w_dff_A_XnwGzwWC9_2;
	wire w_dff_A_DJD2xBfu6_2;
	wire w_dff_A_7t4Mkimw9_2;
	wire w_dff_A_ecrH86MZ3_0;
	wire w_dff_A_CIUS7Gav5_0;
	wire w_dff_A_N15nrHCM4_0;
	wire w_dff_A_hN2WiKWB3_0;
	wire w_dff_A_E2uRmedZ7_0;
	wire w_dff_A_RNPboyHt6_0;
	wire w_dff_A_5SRtP6CE7_0;
	wire w_dff_A_oYAU9c182_1;
	wire w_dff_A_9gtS7jRs7_1;
	wire w_dff_A_kOz5WkqB0_1;
	wire w_dff_A_KNOXphIj4_1;
	wire w_dff_A_9Yn9EafO9_1;
	wire w_dff_A_ms5jV2pR2_1;
	wire w_dff_A_5ltwZ2ye2_1;
	wire w_dff_A_Lt7Qfty51_2;
	wire w_dff_A_e0zbmbUP5_2;
	wire w_dff_A_Q7INts5y4_2;
	wire w_dff_A_VyNIVmih6_2;
	wire w_dff_A_K4nfzJYu7_2;
	wire w_dff_A_mo6qCbGr2_2;
	wire w_dff_A_vkYHzYam5_2;
	wire w_dff_A_BaeaEVsM2_2;
	wire w_dff_A_XgtW6qji8_0;
	wire w_dff_A_JpAMYWHg4_0;
	wire w_dff_A_qEcFQfSS3_0;
	wire w_dff_A_ic3agfWW8_0;
	wire w_dff_A_5YXSH2j93_0;
	wire w_dff_A_mWGi77gq4_0;
	wire w_dff_A_YapfiCWH5_0;
	wire w_dff_A_RuDMLY429_0;
	wire w_dff_A_rvHqpQg65_0;
	wire w_dff_A_tVYmYUbc7_0;
	wire w_dff_A_6tRvnHb68_0;
	wire w_dff_A_zr3ABjfk5_0;
	wire w_dff_A_VX4ll8OB7_0;
	wire w_dff_A_SjsoBwiK5_0;
	wire w_dff_A_n03ppBW46_0;
	wire w_dff_A_MlGXvFTp3_0;
	wire w_dff_A_YFvttSyB0_0;
	wire w_dff_A_nhOyjTGc7_0;
	wire w_dff_A_fKUsN38t3_0;
	wire w_dff_A_BEZMkJS57_0;
	wire w_dff_A_G3Xvkq2P1_0;
	wire w_dff_A_mwAJJ9ZA1_0;
	wire w_dff_A_DfmZ2fx43_0;
	wire w_dff_A_zeiEugJd5_0;
	wire w_dff_A_D1cH4P2b3_1;
	wire w_dff_A_lymXg1rU4_0;
	wire w_dff_A_qVXL5q4A7_0;
	wire w_dff_A_zTTihcWl2_0;
	wire w_dff_A_7ofWyn2G2_0;
	wire w_dff_A_uprW2tFx8_0;
	wire w_dff_A_IjpJGnU97_0;
	wire w_dff_A_q5DJKGA85_0;
	wire w_dff_A_Q8i2HS3Z9_0;
	wire w_dff_A_IkOcXU3g5_0;
	wire w_dff_A_ktK1BNft1_0;
	wire w_dff_A_FfhpUuu83_0;
	wire w_dff_A_tRfRM30g0_0;
	wire w_dff_A_vjNtIkT79_0;
	wire w_dff_A_q70ixND62_0;
	wire w_dff_A_XcsLJeh18_0;
	wire w_dff_A_YEJIxoIy0_0;
	wire w_dff_A_z38LIswg3_0;
	wire w_dff_A_LNiISBmP2_0;
	wire w_dff_A_Etbi6mcC9_0;
	wire w_dff_A_H922DeuZ8_0;
	wire w_dff_A_ZeJnYqn39_0;
	wire w_dff_A_oA6LAxVK4_0;
	wire w_dff_A_VcUXKZc98_0;
	wire w_dff_A_ZYKz2ojx0_2;
	wire w_dff_A_MAt5EeXn0_0;
	wire w_dff_A_Seo4hX7x7_0;
	wire w_dff_A_k6NaR4C44_0;
	wire w_dff_A_V4yQwgQX0_0;
	wire w_dff_A_d0MVzWK97_0;
	wire w_dff_A_0RpYHYl57_0;
	wire w_dff_A_JKHJmjux9_0;
	wire w_dff_A_IMs5XXbX2_0;
	wire w_dff_A_Oep19O2I7_0;
	wire w_dff_A_N6eXX0fK0_0;
	wire w_dff_A_8RXTpRqG7_0;
	wire w_dff_A_65zzfM8Q4_0;
	wire w_dff_A_8bIyJC0G2_0;
	wire w_dff_A_rIsbS6QB5_0;
	wire w_dff_A_0A1jKdQI8_0;
	wire w_dff_A_zRU7muaP3_0;
	wire w_dff_A_ewYtief36_0;
	wire w_dff_A_unEFxqqU1_0;
	wire w_dff_A_oOPWcNbr2_0;
	wire w_dff_A_w0LqHfb65_0;
	wire w_dff_A_c5kn6LU27_2;
	wire w_dff_A_xSALYtp61_0;
	wire w_dff_A_56wXPuXI2_0;
	wire w_dff_A_ihb6mLs17_0;
	wire w_dff_A_QVzgLuCv6_0;
	wire w_dff_A_MDTFNVlg6_0;
	wire w_dff_A_tAWKkV5u1_0;
	wire w_dff_A_VA54F3DT2_0;
	wire w_dff_A_4tCAIW6u7_0;
	wire w_dff_A_D68iNJyj2_0;
	wire w_dff_A_upEdZ1dj3_0;
	wire w_dff_A_07hJC3vz0_0;
	wire w_dff_A_0oCyMF9c1_0;
	wire w_dff_A_u3tYelhM2_0;
	wire w_dff_A_XhLoKl765_0;
	wire w_dff_A_8oeRjjOv6_0;
	wire w_dff_A_Kw1uMcA16_0;
	wire w_dff_A_cm0DJlYr7_0;
	wire w_dff_A_lWjHae9i7_0;
	wire w_dff_A_U4l3J0JQ7_0;
	wire w_dff_A_87c0mXR40_0;
	wire w_dff_A_py3qjAlO6_0;
	wire w_dff_A_8lkpG9yj5_0;
	wire w_dff_A_CvdrDH3z9_0;
	wire w_dff_A_mPRw3Kex9_2;
	wire w_dff_A_y1Q6LEgZ9_0;
	wire w_dff_A_p1bPyM9u7_0;
	wire w_dff_A_rbSnQTIY6_0;
	wire w_dff_A_i3upuMjk4_0;
	wire w_dff_A_UR7UTR4p5_0;
	wire w_dff_A_0u8mcTUR9_0;
	wire w_dff_A_p4ScEj226_0;
	wire w_dff_A_jdihPNqz1_0;
	wire w_dff_A_h2Cz38b28_0;
	wire w_dff_A_GKAkkJ7B6_0;
	wire w_dff_A_jJa7iNCX4_0;
	wire w_dff_A_618NVufX0_0;
	wire w_dff_A_SLEXvMko7_0;
	wire w_dff_A_I20KqZEp7_0;
	wire w_dff_A_kh6Uzcp47_0;
	wire w_dff_A_B59Nuf1J2_0;
	wire w_dff_A_oAY020Le8_0;
	wire w_dff_A_2ALw7X1a9_0;
	wire w_dff_A_pStHHbCW0_0;
	wire w_dff_A_8x7lEdjR2_0;
	wire w_dff_A_8f0RZSV56_0;
	wire w_dff_A_SvdPApWS4_0;
	wire w_dff_A_6ONkQnMn0_0;
	wire w_dff_A_FbzfaOjn5_2;
	wire w_dff_A_KzvB2uNu4_0;
	wire w_dff_A_xWbtP3id0_0;
	wire w_dff_A_pTl5v5kN3_0;
	wire w_dff_A_3TPtL5WN2_0;
	wire w_dff_A_I48EkiSa1_0;
	wire w_dff_A_yTLimDf87_0;
	wire w_dff_A_PNAbjEge8_0;
	wire w_dff_A_dpNyKKEl7_0;
	wire w_dff_A_cp4P7mBH1_0;
	wire w_dff_A_mygSIe9a7_0;
	wire w_dff_A_o7rzffrE2_0;
	wire w_dff_A_nPRB9dci2_0;
	wire w_dff_A_kgTTyovo2_0;
	wire w_dff_A_Ep6aoRix8_2;
	wire w_dff_A_eP3wTA3N7_0;
	wire w_dff_A_OtAf2P787_0;
	wire w_dff_A_WTY8soBG5_0;
	wire w_dff_A_LdX8lXc20_0;
	wire w_dff_A_D608efx06_0;
	wire w_dff_A_LIJAooz69_0;
	wire w_dff_A_VX24oOND5_0;
	wire w_dff_A_SOGSA02F6_0;
	wire w_dff_A_pfdz49sz5_0;
	wire w_dff_A_YnUcfUw68_0;
	wire w_dff_A_iA9WOhAQ2_0;
	wire w_dff_A_vQ0SPl6k0_2;
	wire w_dff_A_JrM6IIrg5_0;
	wire w_dff_A_pklSCn3U3_0;
	wire w_dff_A_TdQOTeQf5_0;
	wire w_dff_A_Pa2E6NBo5_0;
	wire w_dff_A_VI4Dtggs0_0;
	wire w_dff_A_Opq9hlDY1_0;
	wire w_dff_A_0lqtm2la8_0;
	wire w_dff_A_i57QZi4A1_0;
	wire w_dff_A_R1LmDXZA0_0;
	wire w_dff_A_JI7qBb718_0;
	wire w_dff_A_3k4lhRIx4_2;
	wire w_dff_A_nXDml4y44_0;
	wire w_dff_A_Nu36lPLI6_0;
	wire w_dff_A_GFS75Zp92_0;
	wire w_dff_A_xzkZ9uSh1_0;
	wire w_dff_A_TDvoZI8F5_0;
	wire w_dff_A_pEEQiuzB3_0;
	wire w_dff_A_TYhu1Dlb1_0;
	wire w_dff_A_aD5WL3mf0_0;
	wire w_dff_A_C4xbmaE17_0;
	wire w_dff_A_TdpNpc2m6_0;
	wire w_dff_A_OFRPwL4t5_2;
	wire w_dff_A_a9A7N3kO2_0;
	wire w_dff_A_yAxqF3cL1_0;
	wire w_dff_A_QgCylUag0_0;
	wire w_dff_A_Xhk2UlNL3_0;
	wire w_dff_A_WcPydgds6_0;
	wire w_dff_A_emA5oVt34_0;
	wire w_dff_A_euiRlEsq7_0;
	wire w_dff_A_yydSEIER9_0;
	wire w_dff_A_dEJtFI0h0_0;
	wire w_dff_A_LumBvitA5_0;
	wire w_dff_A_ErMg6Nz96_1;
	wire w_dff_A_qUxcG1CY5_0;
	wire w_dff_A_je4DMXyj0_0;
	wire w_dff_A_qMh23JUk2_0;
	wire w_dff_A_36H58dk06_0;
	wire w_dff_A_geHM8Gn20_0;
	wire w_dff_A_2EzwbEhp6_0;
	wire w_dff_A_TWQT8v469_0;
	wire w_dff_A_FbrOxECu5_2;
	wire w_dff_A_sRBNHj852_0;
	wire w_dff_A_n7NXOdYh2_0;
	wire w_dff_A_8lrdO1GS6_0;
	wire w_dff_A_lCop0IM32_0;
	wire w_dff_A_0lqkBuEO4_2;
	wire w_dff_A_sd6gKFIT9_0;
	wire w_dff_A_fvywW1pb5_0;
	wire w_dff_A_uM599SED7_0;
	wire w_dff_A_FzYIJVPg9_0;
	wire w_dff_A_VD26nmsp6_1;
	wire w_dff_A_6bseNoBV9_0;
	wire w_dff_A_V3JHIXrH3_0;
	wire w_dff_A_6Q8Zs9tx2_0;
	wire w_dff_A_tLq9uSYe7_0;
	wire w_dff_A_RN59Cewo1_0;
	wire w_dff_A_znlqw13Q4_0;
	wire w_dff_A_ij4JhiJs2_1;
	wire w_dff_A_6l9hh6411_0;
	wire w_dff_A_mUwWp1dw2_0;
	wire w_dff_A_Q8xVQi4b3_0;
	wire w_dff_A_UIyIURTM6_0;
	wire w_dff_A_C43idKl58_0;
	wire w_dff_A_9yDN0YMg2_1;
	wire w_dff_A_dVn5qsyl7_0;
	wire w_dff_A_zscp8Mq69_0;
	wire w_dff_A_kfqeLiiM7_0;
	wire w_dff_A_lmLOe4yt4_0;
	wire w_dff_A_wSPhLArv2_1;
	wire w_dff_A_3420XUV54_0;
	wire w_dff_A_3MaFdEDz7_0;
	wire w_dff_A_2VxUnDSH8_1;
	wire w_dff_A_OAhS0AMB1_0;
	wire w_dff_A_XEXW3dEe3_0;
	wire w_dff_A_bKJIWztW0_0;
	wire w_dff_A_CC4x2ebW6_0;
	wire w_dff_A_9QSoc5cq7_1;
	wire w_dff_A_5Bcl7rAn0_2;
	jnot g0000(.din(w_G77_5[1]),.dout(n72),.clk(gclk));
	jnot g0001(.din(w_G50_5[2]),.dout(n73),.clk(gclk));
	jnot g0002(.din(w_G58_5[1]),.dout(n74),.clk(gclk));
	jnot g0003(.din(w_G68_5[1]),.dout(n75),.clk(gclk));
	jand g0004(.dina(w_n75_1[1]),.dinb(w_n74_1[1]),.dout(n76),.clk(gclk));
	jand g0005(.dina(w_n76_0[1]),.dinb(w_n73_2[2]),.dout(n77),.clk(gclk));
	jand g0006(.dina(w_n77_0[1]),.dinb(w_n72_1[1]),.dout(w_dff_A_BaeaEVsM2_2),.clk(gclk));
	jnot g0007(.din(w_G97_5[1]),.dout(n79),.clk(gclk));
	jnot g0008(.din(w_G107_5[1]),.dout(n80),.clk(gclk));
	jand g0009(.dina(w_n80_1[1]),.dinb(w_n79_0[2]),.dout(n81),.clk(gclk));
	jnot g0010(.din(w_n81_0[2]),.dout(n82),.clk(gclk));
	jand g0011(.dina(n82),.dinb(w_G87_3[2]),.dout(n83),.clk(gclk));
	jnot g0012(.din(n83),.dout(G355_fa_),.clk(gclk));
	jand g0013(.dina(w_G20_7[1]),.dinb(w_G1_3[1]),.dout(n85),.clk(gclk));
	jnot g0014(.din(w_G226_1[1]),.dout(n86),.clk(gclk));
	jor g0015(.dina(w_n86_0[1]),.dinb(w_n73_2[1]),.dout(n87),.clk(gclk));
	jnot g0016(.din(w_G264_1[1]),.dout(n88),.clk(gclk));
	jor g0017(.dina(w_n88_1[1]),.dinb(w_n80_1[0]),.dout(n89),.clk(gclk));
	jand g0018(.dina(n89),.dinb(n87),.dout(n90),.clk(gclk));
	jnot g0019(.din(w_G257_1[2]),.dout(n91),.clk(gclk));
	jor g0020(.dina(w_n91_1[2]),.dinb(w_n79_0[1]),.dout(n92),.clk(gclk));
	jnot g0021(.din(w_G238_1[2]),.dout(n93),.clk(gclk));
	jor g0022(.dina(w_n93_0[1]),.dinb(w_n75_1[0]),.dout(n94),.clk(gclk));
	jand g0023(.dina(n94),.dinb(n92),.dout(n95),.clk(gclk));
	jand g0024(.dina(n95),.dinb(n90),.dout(n96),.clk(gclk));
	jnot g0025(.din(w_G87_3[1]),.dout(n97),.clk(gclk));
	jnot g0026(.din(w_G250_0[2]),.dout(n98),.clk(gclk));
	jor g0027(.dina(w_n98_2[1]),.dinb(w_n97_2[1]),.dout(n99),.clk(gclk));
	jnot g0028(.din(w_G232_1[2]),.dout(n100),.clk(gclk));
	jor g0029(.dina(n100),.dinb(w_n74_1[0]),.dout(n101),.clk(gclk));
	jand g0030(.dina(n101),.dinb(n99),.dout(n102),.clk(gclk));
	jnot g0031(.din(w_G244_1[2]),.dout(n103),.clk(gclk));
	jor g0032(.dina(w_n103_0[2]),.dinb(w_n72_1[0]),.dout(n104),.clk(gclk));
	jnot g0033(.din(w_G116_4[2]),.dout(n105),.clk(gclk));
	jnot g0034(.din(w_G270_0[2]),.dout(n106),.clk(gclk));
	jor g0035(.dina(w_n106_0[1]),.dinb(w_n105_2[1]),.dout(n107),.clk(gclk));
	jand g0036(.dina(n107),.dinb(n104),.dout(n108),.clk(gclk));
	jand g0037(.dina(n108),.dinb(n102),.dout(n109),.clk(gclk));
	jand g0038(.dina(n109),.dinb(n96),.dout(n110),.clk(gclk));
	jor g0039(.dina(n110),.dinb(w_n85_0[2]),.dout(n111),.clk(gclk));
	jnot g0040(.din(w_G20_7[0]),.dout(n112),.clk(gclk));
	jnot g0041(.din(w_G1_3[0]),.dout(n113),.clk(gclk));
	jnot g0042(.din(w_G13_1[1]),.dout(n114),.clk(gclk));
	jor g0043(.dina(w_n114_1[2]),.dinb(w_n113_3[1]),.dout(n115),.clk(gclk));
	jor g0044(.dina(w_n115_1[1]),.dinb(w_n112_5[2]),.dout(n116),.clk(gclk));
	jnot g0045(.din(w_n76_0[0]),.dout(n117),.clk(gclk));
	jand g0046(.dina(n117),.dinb(w_G50_5[1]),.dout(n118),.clk(gclk));
	jnot g0047(.din(w_n118_0[2]),.dout(n119),.clk(gclk));
	jor g0048(.dina(n119),.dinb(w_n116_0[1]),.dout(n120),.clk(gclk));
	jand g0049(.dina(w_n114_1[1]),.dinb(w_G1_2[2]),.dout(n121),.clk(gclk));
	jand g0050(.dina(w_n121_0[2]),.dinb(w_G20_6[2]),.dout(n122),.clk(gclk));
	jnot g0051(.din(w_n122_1[1]),.dout(n123),.clk(gclk));
	jand g0052(.dina(w_n88_1[0]),.dinb(w_n91_1[1]),.dout(n124),.clk(gclk));
	jor g0053(.dina(n124),.dinb(w_n98_2[0]),.dout(n125),.clk(gclk));
	jor g0054(.dina(w_dff_B_OdmNiY9Q7_0),.dinb(w_n123_1[2]),.dout(n126),.clk(gclk));
	jand g0055(.dina(w_dff_B_brpxkulE2_0),.dinb(n120),.dout(n127),.clk(gclk));
	jand g0056(.dina(n127),.dinb(w_dff_B_27IG3dus8_1),.dout(w_dff_A_ZYKz2ojx0_2),.clk(gclk));
	jxor g0057(.dina(w_G270_0[1]),.dinb(w_G264_1[0]),.dout(n129),.clk(gclk));
	jxor g0058(.dina(w_G257_1[1]),.dinb(w_n98_1[2]),.dout(n130),.clk(gclk));
	jxor g0059(.dina(n130),.dinb(w_dff_B_3TlZntCp2_1),.dout(n131),.clk(gclk));
	jnot g0060(.din(w_n131_0[1]),.dout(n132),.clk(gclk));
	jxor g0061(.dina(w_G244_1[1]),.dinb(w_G238_1[1]),.dout(n133),.clk(gclk));
	jxor g0062(.dina(w_G232_1[1]),.dinb(w_n86_0[0]),.dout(n134),.clk(gclk));
	jxor g0063(.dina(n134),.dinb(w_dff_B_vF6pt99o2_1),.dout(n135),.clk(gclk));
	jxor g0064(.dina(w_n135_0[1]),.dinb(n132),.dout(w_dff_A_c5kn6LU27_2),.clk(gclk));
	jxor g0065(.dina(w_G68_5[0]),.dinb(w_G58_5[0]),.dout(n137),.clk(gclk));
	jnot g0066(.din(w_n137_0[2]),.dout(n138),.clk(gclk));
	jxor g0067(.dina(w_G77_5[0]),.dinb(w_G50_5[0]),.dout(n139),.clk(gclk));
	jxor g0068(.dina(w_dff_B_9Ye4cWSA9_0),.dinb(n138),.dout(n140),.clk(gclk));
	jnot g0069(.din(w_n140_0[1]),.dout(n141),.clk(gclk));
	jxor g0070(.dina(w_G116_4[1]),.dinb(w_G107_5[0]),.dout(n142),.clk(gclk));
	jxor g0071(.dina(w_G97_5[0]),.dinb(w_n97_2[0]),.dout(n143),.clk(gclk));
	jxor g0072(.dina(n143),.dinb(w_dff_B_bujkl3Rf1_1),.dout(n144),.clk(gclk));
	jxor g0073(.dina(w_n144_0[1]),.dinb(n141),.dout(w_dff_A_mPRw3Kex9_2),.clk(gclk));
	jnot g0074(.din(w_G169_1[1]),.dout(n146),.clk(gclk));
	jand g0075(.dina(w_G13_1[0]),.dinb(w_G1_2[1]),.dout(n147),.clk(gclk));
	jnot g0076(.din(w_G33_11[2]),.dout(n148),.clk(gclk));
	jnot g0077(.din(w_G41_1[1]),.dout(n149),.clk(gclk));
	jor g0078(.dina(w_n149_2[1]),.dinb(w_n148_9[2]),.dout(n150),.clk(gclk));
	jand g0079(.dina(n150),.dinb(w_n147_0[2]),.dout(n151),.clk(gclk));
	jand g0080(.dina(w_G1698_0[2]),.dinb(w_n148_9[1]),.dout(n152),.clk(gclk));
	jand g0081(.dina(w_n152_3[1]),.dinb(w_G244_1[0]),.dout(n153),.clk(gclk));
	jnot g0082(.din(w_G1698_0[1]),.dout(n154),.clk(gclk));
	jand g0083(.dina(w_n154_0[1]),.dinb(w_n148_9[0]),.dout(n155),.clk(gclk));
	jand g0084(.dina(w_n155_3[1]),.dinb(w_G238_1[0]),.dout(n156),.clk(gclk));
	jand g0085(.dina(w_G116_4[0]),.dinb(w_G33_11[1]),.dout(n157),.clk(gclk));
	jor g0086(.dina(w_n157_0[2]),.dinb(n156),.dout(n158),.clk(gclk));
	jor g0087(.dina(n158),.dinb(w_dff_B_rwCQmGns8_1),.dout(n159),.clk(gclk));
	jand g0088(.dina(n159),.dinb(w_n151_4[2]),.dout(n160),.clk(gclk));
	jnot g0089(.din(w_G45_1[2]),.dout(n161),.clk(gclk));
	jor g0090(.dina(w_n161_1[1]),.dinb(w_G1_2[0]),.dout(n162),.clk(gclk));
	jand g0091(.dina(w_n162_0[2]),.dinb(w_n98_1[1]),.dout(n163),.clk(gclk));
	jnot g0092(.din(w_n163_0[1]),.dout(n164),.clk(gclk));
	jand g0093(.dina(w_G41_1[0]),.dinb(w_G33_11[0]),.dout(n165),.clk(gclk));
	jor g0094(.dina(w_dff_B_HqtnbwdP0_0),.dinb(w_n115_1[0]),.dout(n166),.clk(gclk));
	jor g0095(.dina(w_n162_0[1]),.dinb(w_G274_0[2]),.dout(n167),.clk(gclk));
	jand g0096(.dina(n167),.dinb(w_n166_3[1]),.dout(n168),.clk(gclk));
	jand g0097(.dina(n168),.dinb(n164),.dout(n169),.clk(gclk));
	jor g0098(.dina(w_dff_B_WNMm4euq5_0),.dinb(n160),.dout(n170),.clk(gclk));
	jand g0099(.dina(w_n170_0[2]),.dinb(w_n146_3[2]),.dout(n171),.clk(gclk));
	jand g0100(.dina(w_G97_4[2]),.dinb(w_G33_10[2]),.dout(n172),.clk(gclk));
	jand g0101(.dina(w_G68_4[2]),.dinb(w_n148_8[2]),.dout(n173),.clk(gclk));
	jor g0102(.dina(n173),.dinb(w_G20_6[1]),.dout(n174),.clk(gclk));
	jor g0103(.dina(n174),.dinb(w_n172_0[1]),.dout(n175),.clk(gclk));
	jnot g0104(.din(n175),.dout(n176),.clk(gclk));
	jor g0105(.dina(w_n112_5[1]),.dinb(w_n113_3[0]),.dout(n177),.clk(gclk));
	jor g0106(.dina(n177),.dinb(w_n148_8[1]),.dout(n178),.clk(gclk));
	jand g0107(.dina(n178),.dinb(w_n115_0[2]),.dout(n179),.clk(gclk));
	jand g0108(.dina(w_n81_0[1]),.dinb(w_n97_1[2]),.dout(n180),.clk(gclk));
	jand g0109(.dina(w_n180_0[1]),.dinb(w_G20_6[0]),.dout(n181),.clk(gclk));
	jor g0110(.dina(n181),.dinb(w_n179_1[2]),.dout(n182),.clk(gclk));
	jor g0111(.dina(n182),.dinb(n176),.dout(n183),.clk(gclk));
	jand g0112(.dina(w_G20_5[2]),.dinb(w_n113_2[2]),.dout(n184),.clk(gclk));
	jand g0113(.dina(n184),.dinb(w_G13_0[2]),.dout(n185),.clk(gclk));
	jand g0114(.dina(w_n185_3[2]),.dinb(w_n97_1[1]),.dout(n186),.clk(gclk));
	jnot g0115(.din(n186),.dout(n187),.clk(gclk));
	jand g0116(.dina(w_n85_0[1]),.dinb(w_G33_10[1]),.dout(n188),.clk(gclk));
	jor g0117(.dina(n188),.dinb(w_n147_0[1]),.dout(n189),.clk(gclk));
	jor g0118(.dina(w_n185_3[1]),.dinb(w_n189_2[1]),.dout(n190),.clk(gclk));
	jand g0119(.dina(w_G33_10[0]),.dinb(w_n113_2[1]),.dout(n191),.clk(gclk));
	jor g0120(.dina(w_n191_0[2]),.dinb(w_n97_1[0]),.dout(n192),.clk(gclk));
	jor g0121(.dina(w_dff_B_ZzgSafiw8_0),.dinb(w_n190_1[2]),.dout(n193),.clk(gclk));
	jand g0122(.dina(n193),.dinb(n187),.dout(n194),.clk(gclk));
	jand g0123(.dina(n194),.dinb(n183),.dout(n195),.clk(gclk));
	jnot g0124(.din(w_G179_2[2]),.dout(n196),.clk(gclk));
	jor g0125(.dina(w_n154_0[0]),.dinb(w_G33_9[2]),.dout(n197),.clk(gclk));
	jor g0126(.dina(w_n197_1[1]),.dinb(w_n103_0[1]),.dout(n198),.clk(gclk));
	jor g0127(.dina(w_G1698_0[0]),.dinb(w_G33_9[1]),.dout(n199),.clk(gclk));
	jor g0128(.dina(w_n199_1[1]),.dinb(w_n93_0[0]),.dout(n200),.clk(gclk));
	jnot g0129(.din(w_n157_0[1]),.dout(n201),.clk(gclk));
	jand g0130(.dina(w_n201_0[1]),.dinb(n200),.dout(n202),.clk(gclk));
	jand g0131(.dina(n202),.dinb(n198),.dout(n203),.clk(gclk));
	jor g0132(.dina(n203),.dinb(w_n166_3[0]),.dout(n204),.clk(gclk));
	jnot g0133(.din(w_G274_0[1]),.dout(n205),.clk(gclk));
	jand g0134(.dina(w_G45_1[1]),.dinb(w_n113_2[0]),.dout(n206),.clk(gclk));
	jand g0135(.dina(w_n206_0[1]),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jor g0136(.dina(n207),.dinb(w_n151_4[1]),.dout(n208),.clk(gclk));
	jor g0137(.dina(n208),.dinb(w_n163_0[0]),.dout(n209),.clk(gclk));
	jand g0138(.dina(n209),.dinb(n204),.dout(n210),.clk(gclk));
	jand g0139(.dina(w_n210_0[2]),.dinb(w_n196_2[2]),.dout(n211),.clk(gclk));
	jor g0140(.dina(n211),.dinb(w_n195_0[1]),.dout(n212),.clk(gclk));
	jor g0141(.dina(n212),.dinb(n171),.dout(n213),.clk(gclk));
	jnot g0142(.din(w_n195_0[0]),.dout(n214),.clk(gclk));
	jand g0143(.dina(w_n210_0[1]),.dinb(w_G190_4[1]),.dout(n215),.clk(gclk));
	jand g0144(.dina(w_n170_0[1]),.dinb(w_G200_4[2]),.dout(n216),.clk(gclk));
	jor g0145(.dina(n216),.dinb(w_dff_B_JFQs6Cz90_1),.dout(n217),.clk(gclk));
	jor g0146(.dina(n217),.dinb(w_n214_0[1]),.dout(n218),.clk(gclk));
	jand g0147(.dina(w_n218_0[1]),.dinb(w_n213_0[1]),.dout(n219),.clk(gclk));
	jor g0148(.dina(w_n197_1[0]),.dinb(w_n98_1[0]),.dout(n220),.clk(gclk));
	jand g0149(.dina(w_G283_3[2]),.dinb(w_G33_9[0]),.dout(n221),.clk(gclk));
	jnot g0150(.din(w_n221_0[2]),.dout(n222),.clk(gclk));
	jor g0151(.dina(w_n199_1[0]),.dinb(w_n103_0[0]),.dout(n223),.clk(gclk));
	jand g0152(.dina(n223),.dinb(n222),.dout(n224),.clk(gclk));
	jand g0153(.dina(n224),.dinb(n220),.dout(n225),.clk(gclk));
	jor g0154(.dina(n225),.dinb(w_n166_2[2]),.dout(n226),.clk(gclk));
	jor g0155(.dina(w_n151_4[0]),.dinb(w_n205_0[0]),.dout(n227),.clk(gclk));
	jor g0156(.dina(w_n162_0[0]),.dinb(w_G41_0[2]),.dout(n228),.clk(gclk));
	jor g0157(.dina(w_n228_0[1]),.dinb(n227),.dout(n229),.clk(gclk));
	jand g0158(.dina(w_n206_0[0]),.dinb(w_n149_2[0]),.dout(n230),.clk(gclk));
	jor g0159(.dina(w_n230_0[1]),.dinb(w_n151_3[2]),.dout(n231),.clk(gclk));
	jor g0160(.dina(w_n231_0[2]),.dinb(w_n91_1[0]),.dout(n232),.clk(gclk));
	jand g0161(.dina(n232),.dinb(w_n229_0[2]),.dout(n233),.clk(gclk));
	jand g0162(.dina(n233),.dinb(w_dff_B_Lh5p2nfy2_1),.dout(n234),.clk(gclk));
	jor g0163(.dina(w_n234_0[2]),.dinb(w_n146_3[1]),.dout(n235),.clk(gclk));
	jand g0164(.dina(w_n152_3[0]),.dinb(w_G250_0[1]),.dout(n236),.clk(gclk));
	jand g0165(.dina(w_n155_3[0]),.dinb(w_G244_0[2]),.dout(n237),.clk(gclk));
	jor g0166(.dina(n237),.dinb(w_n221_0[1]),.dout(n238),.clk(gclk));
	jor g0167(.dina(n238),.dinb(w_dff_B_Pfjezq0K0_1),.dout(n239),.clk(gclk));
	jand g0168(.dina(n239),.dinb(w_n151_3[1]),.dout(n240),.clk(gclk));
	jand g0169(.dina(w_n166_2[1]),.dinb(w_G274_0[0]),.dout(n241),.clk(gclk));
	jand g0170(.dina(w_n230_0[0]),.dinb(w_n241_0[1]),.dout(n242),.clk(gclk));
	jand g0171(.dina(w_n228_0[0]),.dinb(w_n166_2[0]),.dout(n243),.clk(gclk));
	jand g0172(.dina(w_n243_0[2]),.dinb(w_G257_1[0]),.dout(n244),.clk(gclk));
	jor g0173(.dina(n244),.dinb(w_n242_0[2]),.dout(n245),.clk(gclk));
	jor g0174(.dina(n245),.dinb(n240),.dout(n246),.clk(gclk));
	jor g0175(.dina(w_n246_1[1]),.dinb(w_n196_2[1]),.dout(n247),.clk(gclk));
	jand g0176(.dina(n247),.dinb(n235),.dout(n248),.clk(gclk));
	jand g0177(.dina(w_G107_4[2]),.dinb(w_G33_8[2]),.dout(n249),.clk(gclk));
	jand g0178(.dina(w_G77_4[2]),.dinb(w_n148_8[0]),.dout(n250),.clk(gclk));
	jor g0179(.dina(n250),.dinb(w_G20_5[1]),.dout(n251),.clk(gclk));
	jor g0180(.dina(n251),.dinb(w_n249_0[1]),.dout(n252),.clk(gclk));
	jand g0181(.dina(w_G107_4[1]),.dinb(w_G97_4[1]),.dout(n253),.clk(gclk));
	jor g0182(.dina(n253),.dinb(w_n112_5[0]),.dout(n254),.clk(gclk));
	jor g0183(.dina(n254),.dinb(w_n81_0[0]),.dout(n255),.clk(gclk));
	jand g0184(.dina(w_n255_0[1]),.dinb(n252),.dout(n256),.clk(gclk));
	jand g0185(.dina(n256),.dinb(w_n189_2[0]),.dout(n257),.clk(gclk));
	jnot g0186(.din(w_n257_0[1]),.dout(n258),.clk(gclk));
	jand g0187(.dina(w_n185_3[0]),.dinb(w_n79_0[0]),.dout(n259),.clk(gclk));
	jnot g0188(.din(w_n259_0[1]),.dout(n260),.clk(gclk));
	jnot g0189(.din(w_n191_0[1]),.dout(n261),.clk(gclk));
	jand g0190(.dina(w_n261_0[1]),.dinb(w_G97_4[0]),.dout(n262),.clk(gclk));
	jnot g0191(.din(w_n262_0[1]),.dout(n263),.clk(gclk));
	jor g0192(.dina(n263),.dinb(w_n190_1[1]),.dout(n264),.clk(gclk));
	jand g0193(.dina(n264),.dinb(w_dff_B_rjK55iLY6_1),.dout(n265),.clk(gclk));
	jand g0194(.dina(n265),.dinb(n258),.dout(n266),.clk(gclk));
	jor g0195(.dina(w_dff_B_wMQgszaN9_0),.dinb(n248),.dout(n267),.clk(gclk));
	jand g0196(.dina(w_n246_1[0]),.dinb(w_G200_4[1]),.dout(n268),.clk(gclk));
	jor g0197(.dina(w_n112_4[2]),.dinb(w_G1_1[2]),.dout(n269),.clk(gclk));
	jor g0198(.dina(w_n269_1[2]),.dinb(w_n114_1[0]),.dout(n270),.clk(gclk));
	jand g0199(.dina(w_n270_0[1]),.dinb(w_n179_1[1]),.dout(n271),.clk(gclk));
	jand g0200(.dina(w_n262_0[0]),.dinb(w_n271_1[2]),.dout(n272),.clk(gclk));
	jor g0201(.dina(n272),.dinb(w_n259_0[0]),.dout(n273),.clk(gclk));
	jor g0202(.dina(n273),.dinb(w_n257_0[0]),.dout(n274),.clk(gclk));
	jand g0203(.dina(w_n234_0[1]),.dinb(w_G190_4[0]),.dout(n275),.clk(gclk));
	jor g0204(.dina(n275),.dinb(w_n274_0[2]),.dout(n276),.clk(gclk));
	jor g0205(.dina(n276),.dinb(w_dff_B_QdJvX37F8_1),.dout(n277),.clk(gclk));
	jand g0206(.dina(n277),.dinb(n267),.dout(n278),.clk(gclk));
	jand g0207(.dina(w_n278_0[1]),.dinb(w_n219_0[1]),.dout(n279),.clk(gclk));
	jand g0208(.dina(w_n152_2[2]),.dinb(w_G264_0[2]),.dout(n280),.clk(gclk));
	jand g0209(.dina(w_G303_2[2]),.dinb(w_G33_8[1]),.dout(n281),.clk(gclk));
	jand g0210(.dina(w_n155_2[2]),.dinb(w_G257_0[2]),.dout(n282),.clk(gclk));
	jor g0211(.dina(n282),.dinb(w_n281_0[1]),.dout(n283),.clk(gclk));
	jor g0212(.dina(n283),.dinb(w_dff_B_Mur7JrsD8_1),.dout(n284),.clk(gclk));
	jand g0213(.dina(n284),.dinb(w_n151_3[0]),.dout(n285),.clk(gclk));
	jand g0214(.dina(w_n243_0[1]),.dinb(w_G270_0[0]),.dout(n286),.clk(gclk));
	jor g0215(.dina(n286),.dinb(w_n242_0[1]),.dout(n287),.clk(gclk));
	jor g0216(.dina(n287),.dinb(n285),.dout(n288),.clk(gclk));
	jand g0217(.dina(w_n288_1[1]),.dinb(w_n146_3[0]),.dout(n289),.clk(gclk));
	jand g0218(.dina(w_G97_3[2]),.dinb(w_n148_7[2]),.dout(n290),.clk(gclk));
	jor g0219(.dina(n290),.dinb(w_G20_5[0]),.dout(n291),.clk(gclk));
	jor g0220(.dina(n291),.dinb(w_n221_0[0]),.dout(n292),.clk(gclk));
	jand g0221(.dina(w_n105_2[0]),.dinb(w_G20_4[2]),.dout(n293),.clk(gclk));
	jnot g0222(.din(n293),.dout(n294),.clk(gclk));
	jand g0223(.dina(n294),.dinb(w_n189_1[2]),.dout(n295),.clk(gclk));
	jand g0224(.dina(n295),.dinb(n292),.dout(n296),.clk(gclk));
	jnot g0225(.din(w_n296_0[1]),.dout(n297),.clk(gclk));
	jand g0226(.dina(w_n185_2[2]),.dinb(w_n105_1[2]),.dout(n298),.clk(gclk));
	jnot g0227(.din(w_n298_0[1]),.dout(n299),.clk(gclk));
	jor g0228(.dina(w_n191_0[0]),.dinb(w_n105_1[1]),.dout(n300),.clk(gclk));
	jor g0229(.dina(w_n300_0[1]),.dinb(w_n190_1[0]),.dout(n301),.clk(gclk));
	jand g0230(.dina(n301),.dinb(n299),.dout(n302),.clk(gclk));
	jand g0231(.dina(n302),.dinb(n297),.dout(n303),.clk(gclk));
	jor g0232(.dina(w_n197_0[2]),.dinb(w_n88_0[2]),.dout(n304),.clk(gclk));
	jnot g0233(.din(w_n281_0[0]),.dout(n305),.clk(gclk));
	jor g0234(.dina(w_n199_0[2]),.dinb(w_n91_0[2]),.dout(n306),.clk(gclk));
	jand g0235(.dina(n306),.dinb(n305),.dout(n307),.clk(gclk));
	jand g0236(.dina(n307),.dinb(n304),.dout(n308),.clk(gclk));
	jor g0237(.dina(n308),.dinb(w_n166_1[2]),.dout(n309),.clk(gclk));
	jor g0238(.dina(w_n231_0[1]),.dinb(w_n106_0[0]),.dout(n310),.clk(gclk));
	jand g0239(.dina(n310),.dinb(w_n229_0[1]),.dout(n311),.clk(gclk));
	jand g0240(.dina(n311),.dinb(w_dff_B_f909SO4t3_1),.dout(n312),.clk(gclk));
	jand g0241(.dina(w_n312_1[1]),.dinb(w_n196_2[0]),.dout(n313),.clk(gclk));
	jor g0242(.dina(n313),.dinb(w_n303_0[1]),.dout(n314),.clk(gclk));
	jor g0243(.dina(n314),.dinb(w_dff_B_HPMsywrA8_1),.dout(n315),.clk(gclk));
	jand g0244(.dina(w_n288_1[0]),.dinb(w_G200_4[0]),.dout(n316),.clk(gclk));
	jnot g0245(.din(w_n300_0[0]),.dout(n317),.clk(gclk));
	jand g0246(.dina(w_dff_B_eIoYXnst0_0),.dinb(w_n271_1[1]),.dout(n318),.clk(gclk));
	jor g0247(.dina(n318),.dinb(w_n298_0[0]),.dout(n319),.clk(gclk));
	jor g0248(.dina(n319),.dinb(w_n296_0[0]),.dout(n320),.clk(gclk));
	jand g0249(.dina(w_n312_1[0]),.dinb(w_G190_3[2]),.dout(n321),.clk(gclk));
	jor g0250(.dina(n321),.dinb(w_n320_0[1]),.dout(n322),.clk(gclk));
	jor g0251(.dina(n322),.dinb(w_dff_B_dx20306R1_1),.dout(n323),.clk(gclk));
	jand g0252(.dina(n323),.dinb(w_n315_0[1]),.dout(n324),.clk(gclk));
	jor g0253(.dina(w_n97_0[2]),.dinb(w_G33_8[0]),.dout(n325),.clk(gclk));
	jand g0254(.dina(n325),.dinb(w_n112_4[1]),.dout(n326),.clk(gclk));
	jand g0255(.dina(n326),.dinb(w_n201_0[0]),.dout(n327),.clk(gclk));
	jor g0256(.dina(n327),.dinb(w_n179_1[0]),.dout(n328),.clk(gclk));
	jor g0257(.dina(w_n328_0[1]),.dinb(w_G20_4[1]),.dout(n329),.clk(gclk));
	jand g0258(.dina(n329),.dinb(w_G107_4[0]),.dout(n330),.clk(gclk));
	jand g0259(.dina(w_n328_0[0]),.dinb(w_n270_0[0]),.dout(n331),.clk(gclk));
	jor g0260(.dina(w_dff_B_8oMyJe3n5_0),.dinb(n330),.dout(n332),.clk(gclk));
	jand g0261(.dina(w_n261_0[0]),.dinb(w_G107_3[2]),.dout(n333),.clk(gclk));
	jand g0262(.dina(w_dff_B_YJgMbXiN0_0),.dinb(w_n271_1[0]),.dout(n334),.clk(gclk));
	jnot g0263(.din(w_n334_0[1]),.dout(n335),.clk(gclk));
	jand g0264(.dina(w_dff_B_0hyWijOB1_0),.dinb(n332),.dout(n336),.clk(gclk));
	jor g0265(.dina(w_n197_0[1]),.dinb(w_n91_0[1]),.dout(n337),.clk(gclk));
	jor g0266(.dina(w_n199_0[1]),.dinb(w_n98_0[2]),.dout(n338),.clk(gclk));
	jand g0267(.dina(w_G294_3[1]),.dinb(w_G33_7[2]),.dout(n339),.clk(gclk));
	jnot g0268(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jand g0269(.dina(n340),.dinb(n338),.dout(n341),.clk(gclk));
	jand g0270(.dina(n341),.dinb(n337),.dout(n342),.clk(gclk));
	jor g0271(.dina(n342),.dinb(w_n166_1[1]),.dout(n343),.clk(gclk));
	jor g0272(.dina(w_n231_0[0]),.dinb(w_n88_0[1]),.dout(n344),.clk(gclk));
	jand g0273(.dina(n344),.dinb(w_n229_0[0]),.dout(n345),.clk(gclk));
	jand g0274(.dina(n345),.dinb(w_dff_B_AzoIUIvS6_1),.dout(n346),.clk(gclk));
	jand g0275(.dina(w_n346_1[1]),.dinb(w_n196_1[2]),.dout(n347),.clk(gclk));
	jand g0276(.dina(w_n152_2[1]),.dinb(w_G257_0[1]),.dout(n348),.clk(gclk));
	jand g0277(.dina(w_n155_2[1]),.dinb(w_G250_0[0]),.dout(n349),.clk(gclk));
	jor g0278(.dina(w_n339_0[0]),.dinb(n349),.dout(n350),.clk(gclk));
	jor g0279(.dina(n350),.dinb(w_dff_B_hX57umbd8_1),.dout(n351),.clk(gclk));
	jand g0280(.dina(n351),.dinb(w_n151_2[2]),.dout(n352),.clk(gclk));
	jand g0281(.dina(w_n243_0[0]),.dinb(w_G264_0[1]),.dout(n353),.clk(gclk));
	jor g0282(.dina(n353),.dinb(w_n242_0[0]),.dout(n354),.clk(gclk));
	jor g0283(.dina(n354),.dinb(n352),.dout(n355),.clk(gclk));
	jand g0284(.dina(w_n355_1[1]),.dinb(w_n146_2[2]),.dout(n356),.clk(gclk));
	jor g0285(.dina(n356),.dinb(n347),.dout(n357),.clk(gclk));
	jor g0286(.dina(n357),.dinb(n336),.dout(n358),.clk(gclk));
	jand g0287(.dina(w_G87_3[0]),.dinb(w_n148_7[1]),.dout(n359),.clk(gclk));
	jor g0288(.dina(n359),.dinb(w_G20_4[0]),.dout(n360),.clk(gclk));
	jor g0289(.dina(n360),.dinb(w_n157_0[0]),.dout(n361),.clk(gclk));
	jand g0290(.dina(n361),.dinb(w_n189_1[1]),.dout(n362),.clk(gclk));
	jand g0291(.dina(w_n362_0[1]),.dinb(w_n112_4[0]),.dout(n363),.clk(gclk));
	jor g0292(.dina(n363),.dinb(w_n80_0[2]),.dout(n364),.clk(gclk));
	jor g0293(.dina(w_n362_0[0]),.dinb(w_n185_2[1]),.dout(n365),.clk(gclk));
	jand g0294(.dina(w_dff_B_M01Athst6_0),.dinb(n364),.dout(n366),.clk(gclk));
	jor g0295(.dina(w_n334_0[0]),.dinb(n366),.dout(n367),.clk(gclk));
	jor g0296(.dina(w_n355_1[0]),.dinb(w_G190_3[1]),.dout(n368),.clk(gclk));
	jor g0297(.dina(w_n346_1[0]),.dinb(w_G200_3[2]),.dout(n369),.clk(gclk));
	jand g0298(.dina(n369),.dinb(n368),.dout(n370),.clk(gclk));
	jor g0299(.dina(n370),.dinb(w_n367_0[2]),.dout(n371),.clk(gclk));
	jand g0300(.dina(w_n371_0[1]),.dinb(n358),.dout(n372),.clk(gclk));
	jand g0301(.dina(w_n372_0[1]),.dinb(w_n324_0[1]),.dout(n373),.clk(gclk));
	jand g0302(.dina(n373),.dinb(w_n279_0[1]),.dout(n374),.clk(gclk));
	jand g0303(.dina(w_n155_2[0]),.dinb(w_G232_1[0]),.dout(n375),.clk(gclk));
	jand g0304(.dina(w_n152_2[0]),.dinb(w_G238_0[2]),.dout(n376),.clk(gclk));
	jor g0305(.dina(n376),.dinb(w_n249_0[0]),.dout(n377),.clk(gclk));
	jor g0306(.dina(n377),.dinb(w_dff_B_5oDl5aKy0_1),.dout(n378),.clk(gclk));
	jand g0307(.dina(n378),.dinb(w_n151_2[1]),.dout(n379),.clk(gclk));
	jand g0308(.dina(w_n161_1[0]),.dinb(w_n149_1[2]),.dout(n380),.clk(gclk));
	jor g0309(.dina(n380),.dinb(w_G1_1[1]),.dout(n381),.clk(gclk));
	jand g0310(.dina(w_n381_0[1]),.dinb(w_n166_1[0]),.dout(n382),.clk(gclk));
	jand g0311(.dina(w_n382_1[1]),.dinb(w_G244_0[1]),.dout(n383),.clk(gclk));
	jnot g0312(.din(w_n381_0[0]),.dout(n384),.clk(gclk));
	jand g0313(.dina(n384),.dinb(w_n241_0[0]),.dout(n385),.clk(gclk));
	jor g0314(.dina(w_n385_1[1]),.dinb(n383),.dout(n386),.clk(gclk));
	jor g0315(.dina(n386),.dinb(n379),.dout(n387),.clk(gclk));
	jand g0316(.dina(w_n387_1[1]),.dinb(w_n146_2[1]),.dout(n388),.clk(gclk));
	jnot g0317(.din(n388),.dout(n389),.clk(gclk));
	jand g0318(.dina(w_G87_2[2]),.dinb(w_G33_7[1]),.dout(n390),.clk(gclk));
	jand g0319(.dina(w_G58_4[2]),.dinb(w_n148_7[0]),.dout(n391),.clk(gclk));
	jor g0320(.dina(n391),.dinb(w_G20_3[2]),.dout(n392),.clk(gclk));
	jor g0321(.dina(n392),.dinb(w_n390_0[1]),.dout(n393),.clk(gclk));
	jor g0322(.dina(w_G77_4[1]),.dinb(w_n112_3[2]),.dout(n394),.clk(gclk));
	jand g0323(.dina(w_dff_B_FlaDmVrW3_0),.dinb(w_n189_1[0]),.dout(n395),.clk(gclk));
	jand g0324(.dina(n395),.dinb(n393),.dout(n396),.clk(gclk));
	jand g0325(.dina(w_n185_2[0]),.dinb(w_n72_0[2]),.dout(n397),.clk(gclk));
	jand g0326(.dina(w_n269_1[1]),.dinb(w_G77_4[0]),.dout(n398),.clk(gclk));
	jand g0327(.dina(w_dff_B_7bGxVacK4_0),.dinb(w_n271_0[2]),.dout(n399),.clk(gclk));
	jor g0328(.dina(n399),.dinb(w_dff_B_5UrRsifg7_1),.dout(n400),.clk(gclk));
	jor g0329(.dina(n400),.dinb(w_dff_B_RrKfitDe2_1),.dout(n401),.clk(gclk));
	jor g0330(.dina(w_n387_1[0]),.dinb(w_G179_2[1]),.dout(n402),.clk(gclk));
	jand g0331(.dina(n402),.dinb(w_n401_0[2]),.dout(n403),.clk(gclk));
	jand g0332(.dina(n403),.dinb(n389),.dout(n404),.clk(gclk));
	jnot g0333(.din(w_n404_0[2]),.dout(n405),.clk(gclk));
	jand g0334(.dina(w_n387_0[2]),.dinb(w_G200_3[1]),.dout(n406),.clk(gclk));
	jnot g0335(.din(w_G190_3[0]),.dout(n407),.clk(gclk));
	jor g0336(.dina(w_n387_0[1]),.dinb(w_n407_2[1]),.dout(n408),.clk(gclk));
	jnot g0337(.din(n408),.dout(n409),.clk(gclk));
	jor g0338(.dina(n409),.dinb(w_n401_0[1]),.dout(n410),.clk(gclk));
	jor g0339(.dina(n410),.dinb(w_dff_B_2IrSLCfN1_1),.dout(n411),.clk(gclk));
	jand g0340(.dina(n411),.dinb(w_n405_0[1]),.dout(n412),.clk(gclk));
	jand g0341(.dina(w_n155_1[2]),.dinb(w_G226_1[0]),.dout(n413),.clk(gclk));
	jand g0342(.dina(w_n152_1[2]),.dinb(w_G232_0[2]),.dout(n414),.clk(gclk));
	jor g0343(.dina(n414),.dinb(w_n172_0[0]),.dout(n415),.clk(gclk));
	jor g0344(.dina(n415),.dinb(w_dff_B_DmEc0be85_1),.dout(n416),.clk(gclk));
	jand g0345(.dina(n416),.dinb(w_n151_2[0]),.dout(n417),.clk(gclk));
	jand g0346(.dina(w_n382_1[0]),.dinb(w_G238_0[1]),.dout(n418),.clk(gclk));
	jor g0347(.dina(n418),.dinb(w_n385_1[0]),.dout(n419),.clk(gclk));
	jor g0348(.dina(n419),.dinb(n417),.dout(n420),.clk(gclk));
	jand g0349(.dina(w_n420_1[1]),.dinb(w_n146_2[0]),.dout(n421),.clk(gclk));
	jnot g0350(.din(n421),.dout(n422),.clk(gclk));
	jand g0351(.dina(w_n269_1[0]),.dinb(w_G68_4[1]),.dout(n423),.clk(gclk));
	jand g0352(.dina(w_dff_B_kQIUHOkP2_0),.dinb(w_n271_0[1]),.dout(n424),.clk(gclk));
	jand g0353(.dina(w_n148_6[2]),.dinb(w_n114_0[2]),.dout(n425),.clk(gclk));
	jnot g0354(.din(w_n425_1[2]),.dout(n426),.clk(gclk));
	jand g0355(.dina(w_n426_0[1]),.dinb(w_n85_0[0]),.dout(n427),.clk(gclk));
	jor g0356(.dina(n427),.dinb(w_n185_1[2]),.dout(n428),.clk(gclk));
	jand g0357(.dina(n428),.dinb(w_n75_0[2]),.dout(n429),.clk(gclk));
	jand g0358(.dina(w_G77_3[2]),.dinb(w_G33_7[0]),.dout(n430),.clk(gclk));
	jand g0359(.dina(w_G50_4[2]),.dinb(w_n148_6[1]),.dout(n431),.clk(gclk));
	jor g0360(.dina(n431),.dinb(w_n430_0[1]),.dout(n432),.clk(gclk));
	jand g0361(.dina(n432),.dinb(w_n112_3[1]),.dout(n433),.clk(gclk));
	jand g0362(.dina(n433),.dinb(w_n189_0[2]),.dout(n434),.clk(gclk));
	jor g0363(.dina(w_dff_B_IkMZBkBp9_0),.dinb(n429),.dout(n435),.clk(gclk));
	jor g0364(.dina(n435),.dinb(w_dff_B_tzQ4OxgE2_1),.dout(n436),.clk(gclk));
	jor g0365(.dina(w_n420_1[0]),.dinb(w_G179_2[0]),.dout(n437),.clk(gclk));
	jand g0366(.dina(n437),.dinb(w_n436_0[2]),.dout(n438),.clk(gclk));
	jand g0367(.dina(n438),.dinb(n422),.dout(n439),.clk(gclk));
	jnot g0368(.din(w_n439_1[1]),.dout(n440),.clk(gclk));
	jand g0369(.dina(w_n420_0[2]),.dinb(w_G200_3[0]),.dout(n441),.clk(gclk));
	jor g0370(.dina(w_n420_0[1]),.dinb(w_n407_2[0]),.dout(n442),.clk(gclk));
	jnot g0371(.din(n442),.dout(n443),.clk(gclk));
	jor g0372(.dina(n443),.dinb(w_n436_0[1]),.dout(n444),.clk(gclk));
	jor g0373(.dina(n444),.dinb(w_dff_B_X5McmxHP1_1),.dout(n445),.clk(gclk));
	jand g0374(.dina(w_n445_0[1]),.dinb(n440),.dout(n446),.clk(gclk));
	jand g0375(.dina(w_n446_0[1]),.dinb(w_n412_0[1]),.dout(n447),.clk(gclk));
	jand g0376(.dina(w_n152_1[1]),.dinb(w_G223_0[1]),.dout(n448),.clk(gclk));
	jand g0377(.dina(w_n155_1[1]),.dinb(w_dff_B_6p6SfMK66_1),.dout(n449),.clk(gclk));
	jor g0378(.dina(n449),.dinb(w_n430_0[0]),.dout(n450),.clk(gclk));
	jor g0379(.dina(n450),.dinb(w_dff_B_O8CWMqll9_1),.dout(n451),.clk(gclk));
	jand g0380(.dina(n451),.dinb(w_n151_1[2]),.dout(n452),.clk(gclk));
	jand g0381(.dina(w_n382_0[2]),.dinb(w_G226_0[2]),.dout(n453),.clk(gclk));
	jor g0382(.dina(n453),.dinb(w_n385_0[2]),.dout(n454),.clk(gclk));
	jor g0383(.dina(n454),.dinb(n452),.dout(n455),.clk(gclk));
	jand g0384(.dina(w_n455_0[2]),.dinb(w_n146_1[2]),.dout(n456),.clk(gclk));
	jand g0385(.dina(w_n269_0[2]),.dinb(w_G50_4[1]),.dout(n457),.clk(gclk));
	jnot g0386(.din(n457),.dout(n458),.clk(gclk));
	jor g0387(.dina(n458),.dinb(w_n190_0[2]),.dout(n459),.clk(gclk));
	jor g0388(.dina(w_n77_0[0]),.dinb(w_n112_3[0]),.dout(n460),.clk(gclk));
	jnot g0389(.din(w_G150_3[1]),.dout(n461),.clk(gclk));
	jand g0390(.dina(w_n148_6[0]),.dinb(w_n112_2[2]),.dout(n462),.clk(gclk));
	jnot g0391(.din(w_n462_0[2]),.dout(n463),.clk(gclk));
	jor g0392(.dina(n463),.dinb(w_dff_B_1IiMTn0s3_1),.dout(n464),.clk(gclk));
	jand g0393(.dina(w_G33_6[2]),.dinb(w_n112_2[1]),.dout(n465),.clk(gclk));
	jand g0394(.dina(w_n465_0[1]),.dinb(w_G58_4[1]),.dout(n466),.clk(gclk));
	jnot g0395(.din(n466),.dout(n467),.clk(gclk));
	jand g0396(.dina(n467),.dinb(n464),.dout(n468),.clk(gclk));
	jand g0397(.dina(n468),.dinb(w_dff_B_Sggb8bRB2_1),.dout(n469),.clk(gclk));
	jor g0398(.dina(n469),.dinb(w_n179_0[2]),.dout(n470),.clk(gclk));
	jand g0399(.dina(w_n185_1[1]),.dinb(w_n73_2[0]),.dout(n471),.clk(gclk));
	jnot g0400(.din(n471),.dout(n472),.clk(gclk));
	jand g0401(.dina(w_dff_B_BmUIe2270_0),.dinb(n470),.dout(n473),.clk(gclk));
	jand g0402(.dina(n473),.dinb(w_dff_B_fXFLWVgQ2_1),.dout(n474),.clk(gclk));
	jnot g0403(.din(w_n455_0[1]),.dout(n475),.clk(gclk));
	jand g0404(.dina(w_n475_0[1]),.dinb(w_n196_1[1]),.dout(n476),.clk(gclk));
	jor g0405(.dina(n476),.dinb(w_n474_0[1]),.dout(n477),.clk(gclk));
	jor g0406(.dina(n477),.dinb(w_dff_B_sob5fowR5_1),.dout(n478),.clk(gclk));
	jnot g0407(.din(w_n474_0[0]),.dout(n479),.clk(gclk));
	jand g0408(.dina(w_n475_0[0]),.dinb(w_G190_2[2]),.dout(n480),.clk(gclk));
	jand g0409(.dina(w_n455_0[0]),.dinb(w_G200_2[2]),.dout(n481),.clk(gclk));
	jor g0410(.dina(w_dff_B_QXqYkzoH9_0),.dinb(n480),.dout(n482),.clk(gclk));
	jor g0411(.dina(n482),.dinb(w_n479_0[1]),.dout(n483),.clk(gclk));
	jand g0412(.dina(w_n483_0[1]),.dinb(w_n478_0[1]),.dout(n484),.clk(gclk));
	jand g0413(.dina(w_n152_1[0]),.dinb(w_G226_0[1]),.dout(n485),.clk(gclk));
	jand g0414(.dina(w_n155_1[0]),.dinb(w_G223_0[0]),.dout(n486),.clk(gclk));
	jor g0415(.dina(n486),.dinb(w_n390_0[0]),.dout(n487),.clk(gclk));
	jor g0416(.dina(n487),.dinb(w_dff_B_DaWjeVjL0_1),.dout(n488),.clk(gclk));
	jand g0417(.dina(n488),.dinb(w_n151_1[1]),.dout(n489),.clk(gclk));
	jand g0418(.dina(w_n382_0[1]),.dinb(w_G232_0[1]),.dout(n490),.clk(gclk));
	jor g0419(.dina(n490),.dinb(w_n385_0[1]),.dout(n491),.clk(gclk));
	jor g0420(.dina(n491),.dinb(n489),.dout(n492),.clk(gclk));
	jand g0421(.dina(w_n492_0[2]),.dinb(w_n146_1[1]),.dout(n493),.clk(gclk));
	jand g0422(.dina(w_n269_0[1]),.dinb(w_G58_4[0]),.dout(n494),.clk(gclk));
	jnot g0423(.din(n494),.dout(n495),.clk(gclk));
	jor g0424(.dina(n495),.dinb(w_n190_0[1]),.dout(n496),.clk(gclk));
	jor g0425(.dina(w_n137_0[1]),.dinb(w_n112_2[0]),.dout(n497),.clk(gclk));
	jand g0426(.dina(w_n462_0[1]),.dinb(w_G159_3[2]),.dout(n498),.clk(gclk));
	jand g0427(.dina(w_n465_0[0]),.dinb(w_G68_4[0]),.dout(n499),.clk(gclk));
	jor g0428(.dina(n499),.dinb(n498),.dout(n500),.clk(gclk));
	jnot g0429(.din(n500),.dout(n501),.clk(gclk));
	jand g0430(.dina(n501),.dinb(w_dff_B_KQl9HTF33_1),.dout(n502),.clk(gclk));
	jor g0431(.dina(n502),.dinb(w_n179_0[1]),.dout(n503),.clk(gclk));
	jand g0432(.dina(w_n185_1[0]),.dinb(w_n74_0[2]),.dout(n504),.clk(gclk));
	jnot g0433(.din(n504),.dout(n505),.clk(gclk));
	jand g0434(.dina(w_dff_B_4GyJWtJN6_0),.dinb(n503),.dout(n506),.clk(gclk));
	jand g0435(.dina(n506),.dinb(w_dff_B_g2sFFUCp9_1),.dout(n507),.clk(gclk));
	jnot g0436(.din(w_n492_0[1]),.dout(n508),.clk(gclk));
	jand g0437(.dina(w_n508_0[1]),.dinb(w_n196_1[0]),.dout(n509),.clk(gclk));
	jor g0438(.dina(n509),.dinb(w_n507_0[1]),.dout(n510),.clk(gclk));
	jor g0439(.dina(n510),.dinb(w_dff_B_wq0pYMBx5_1),.dout(n511),.clk(gclk));
	jnot g0440(.din(w_n507_0[0]),.dout(n512),.clk(gclk));
	jand g0441(.dina(w_n508_0[0]),.dinb(w_G190_2[1]),.dout(n513),.clk(gclk));
	jand g0442(.dina(w_n492_0[0]),.dinb(w_G200_2[1]),.dout(n514),.clk(gclk));
	jor g0443(.dina(w_dff_B_eHtuai9V9_0),.dinb(n513),.dout(n515),.clk(gclk));
	jor g0444(.dina(n515),.dinb(w_n512_0[1]),.dout(n516),.clk(gclk));
	jand g0445(.dina(w_n516_0[1]),.dinb(w_n511_0[1]),.dout(n517),.clk(gclk));
	jand g0446(.dina(w_n517_0[1]),.dinb(w_n484_0[1]),.dout(n518),.clk(gclk));
	jand g0447(.dina(n518),.dinb(n447),.dout(n519),.clk(gclk));
	jand g0448(.dina(w_n519_1[2]),.dinb(w_n374_0[1]),.dout(w_dff_A_FbzfaOjn5_2),.clk(gclk));
	jor g0449(.dina(w_n355_0[2]),.dinb(w_G179_1[2]),.dout(n521),.clk(gclk));
	jor g0450(.dina(w_n346_0[2]),.dinb(w_G169_1[0]),.dout(n522),.clk(gclk));
	jand g0451(.dina(n522),.dinb(n521),.dout(n523),.clk(gclk));
	jand g0452(.dina(w_n523_0[1]),.dinb(w_n367_0[1]),.dout(n524),.clk(gclk));
	jor g0453(.dina(w_n312_0[2]),.dinb(w_G169_0[2]),.dout(n525),.clk(gclk));
	jor g0454(.dina(w_n288_0[2]),.dinb(w_G179_1[1]),.dout(n526),.clk(gclk));
	jand g0455(.dina(n526),.dinb(w_n320_0[0]),.dout(n527),.clk(gclk));
	jand g0456(.dina(n527),.dinb(w_dff_B_tmtaSXRO8_1),.dout(n528),.clk(gclk));
	jand g0457(.dina(w_n371_0[0]),.dinb(w_n528_0[1]),.dout(n529),.clk(gclk));
	jor g0458(.dina(n529),.dinb(w_n524_0[1]),.dout(n530),.clk(gclk));
	jand g0459(.dina(n530),.dinb(w_n279_0[0]),.dout(n531),.clk(gclk));
	jnot g0460(.din(w_n213_0[0]),.dout(n532),.clk(gclk));
	jand g0461(.dina(w_n246_0[2]),.dinb(w_G169_0[1]),.dout(n533),.clk(gclk));
	jand g0462(.dina(w_n234_0[0]),.dinb(w_G179_1[0]),.dout(n534),.clk(gclk));
	jor g0463(.dina(w_n534_0[1]),.dinb(n533),.dout(n535),.clk(gclk));
	jand g0464(.dina(w_n274_0[1]),.dinb(n535),.dout(n536),.clk(gclk));
	jand g0465(.dina(w_n536_0[2]),.dinb(w_n218_0[0]),.dout(n537),.clk(gclk));
	jor g0466(.dina(n537),.dinb(w_n532_0[1]),.dout(n538),.clk(gclk));
	jor g0467(.dina(w_dff_B_8wZLjwLq1_0),.dinb(n531),.dout(n539),.clk(gclk));
	jand g0468(.dina(w_n539_0[1]),.dinb(w_n519_1[1]),.dout(n540),.clk(gclk));
	jnot g0469(.din(w_n478_0[0]),.dout(n541),.clk(gclk));
	jnot g0470(.din(w_n511_0[0]),.dout(n542),.clk(gclk));
	jor g0471(.dina(w_n439_1[0]),.dinb(w_n404_0[1]),.dout(n543),.clk(gclk));
	jand g0472(.dina(w_n543_0[1]),.dinb(w_n445_0[0]),.dout(n544),.clk(gclk));
	jor g0473(.dina(n544),.dinb(w_n542_0[2]),.dout(n545),.clk(gclk));
	jand g0474(.dina(n545),.dinb(w_n516_0[0]),.dout(n546),.clk(gclk));
	jor g0475(.dina(n546),.dinb(w_n541_0[1]),.dout(n547),.clk(gclk));
	jand g0476(.dina(n547),.dinb(w_n483_0[0]),.dout(n548),.clk(gclk));
	jor g0477(.dina(w_n548_0[2]),.dinb(w_dff_B_P1MteBTm6_1),.dout(w_dff_A_Ep6aoRix8_2),.clk(gclk));
	jand g0478(.dina(w_n112_1[2]),.dinb(w_G13_0[1]),.dout(n550),.clk(gclk));
	jand g0479(.dina(w_G213_0[2]),.dinb(w_n113_1[2]),.dout(n551),.clk(gclk));
	jand g0480(.dina(n551),.dinb(w_n550_0[1]),.dout(n552),.clk(gclk));
	jand g0481(.dina(w_n552_1[1]),.dinb(w_G343_0[1]),.dout(n553),.clk(gclk));
	jnot g0482(.din(w_n553_2[2]),.dout(n554),.clk(gclk));
	jand g0483(.dina(w_n554_3[2]),.dinb(w_n524_0[0]),.dout(n555),.clk(gclk));
	jand g0484(.dina(w_n554_3[1]),.dinb(w_n528_0[0]),.dout(n556),.clk(gclk));
	jand g0485(.dina(w_n553_2[1]),.dinb(w_n367_0[0]),.dout(n557),.clk(gclk));
	jnot g0486(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jand g0487(.dina(n558),.dinb(w_n372_0[0]),.dout(n559),.clk(gclk));
	jand g0488(.dina(w_n557_0[0]),.dinb(w_n523_0[0]),.dout(n560),.clk(gclk));
	jor g0489(.dina(w_dff_B_pKNYMOUG6_0),.dinb(n559),.dout(n561),.clk(gclk));
	jand g0490(.dina(w_n561_0[2]),.dinb(w_n556_0[1]),.dout(n562),.clk(gclk));
	jor g0491(.dina(n562),.dinb(w_dff_B_BOKcaclG7_1),.dout(n563),.clk(gclk));
	jnot g0492(.din(w_n561_0[1]),.dout(n564),.clk(gclk));
	jnot g0493(.din(w_G330_0[1]),.dout(n565),.clk(gclk));
	jnot g0494(.din(w_n324_0[0]),.dout(n566),.clk(gclk));
	jor g0495(.dina(w_n554_3[0]),.dinb(w_n303_0[0]),.dout(n567),.clk(gclk));
	jnot g0496(.din(w_n567_0[1]),.dout(n568),.clk(gclk));
	jor g0497(.dina(w_dff_B_CqHJVKye5_0),.dinb(n566),.dout(n569),.clk(gclk));
	jor g0498(.dina(w_n567_0[0]),.dinb(w_n315_0[0]),.dout(n570),.clk(gclk));
	jand g0499(.dina(w_dff_B_ISAkrs8o5_0),.dinb(n569),.dout(n571),.clk(gclk));
	jor g0500(.dina(w_n571_0[2]),.dinb(w_n565_0[1]),.dout(n572),.clk(gclk));
	jor g0501(.dina(w_n572_0[2]),.dinb(w_n564_0[1]),.dout(n573),.clk(gclk));
	jnot g0502(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jor g0503(.dina(n574),.dinb(w_n563_0[2]),.dout(w_dff_A_vQ0SPl6k0_2),.clk(gclk));
	jand g0504(.dina(w_n554_2[2]),.dinb(w_n539_0[0]),.dout(n576),.clk(gclk));
	jor g0505(.dina(w_n553_2[0]),.dinb(w_n374_0[0]),.dout(n577),.clk(gclk));
	jand g0506(.dina(w_n346_0[1]),.dinb(w_n210_0[0]),.dout(n578),.clk(gclk));
	jand g0507(.dina(n578),.dinb(w_n312_0[1]),.dout(n579),.clk(gclk));
	jand g0508(.dina(n579),.dinb(w_n534_0[0]),.dout(n580),.clk(gclk));
	jand g0509(.dina(w_n288_0[1]),.dinb(w_n196_0[2]),.dout(n581),.clk(gclk));
	jand g0510(.dina(w_n355_0[1]),.dinb(w_n246_0[1]),.dout(n582),.clk(gclk));
	jand g0511(.dina(n582),.dinb(w_n170_0[0]),.dout(n583),.clk(gclk));
	jand g0512(.dina(n583),.dinb(w_dff_B_1acgoLbH7_1),.dout(n584),.clk(gclk));
	jor g0513(.dina(n584),.dinb(w_n554_2[1]),.dout(n585),.clk(gclk));
	jor g0514(.dina(n585),.dinb(w_dff_B_LVfRVNFb1_1),.dout(n586),.clk(gclk));
	jand g0515(.dina(n586),.dinb(w_G330_0[0]),.dout(n587),.clk(gclk));
	jand g0516(.dina(w_dff_B_ShiCuMxf1_0),.dinb(n577),.dout(n588),.clk(gclk));
	jor g0517(.dina(w_n588_1[1]),.dinb(w_n576_1[1]),.dout(n589),.clk(gclk));
	jand g0518(.dina(w_n589_1[2]),.dinb(w_n113_1[1]),.dout(n590),.clk(gclk));
	jand g0519(.dina(w_n122_1[0]),.dinb(w_n149_1[1]),.dout(n591),.clk(gclk));
	jnot g0520(.din(w_n591_1[1]),.dout(n592),.clk(gclk));
	jand g0521(.dina(w_n180_0[0]),.dinb(w_n105_1[0]),.dout(n593),.clk(gclk));
	jand g0522(.dina(w_n593_0[2]),.dinb(w_G1_1[0]),.dout(n594),.clk(gclk));
	jand g0523(.dina(n594),.dinb(w_n592_2[1]),.dout(n595),.clk(gclk));
	jand g0524(.dina(w_n591_1[0]),.dinb(w_n118_0[1]),.dout(n596),.clk(gclk));
	jor g0525(.dina(w_dff_B_EWujXDTd0_0),.dinb(n595),.dout(n597),.clk(gclk));
	jor g0526(.dina(w_dff_B_CQkULghC5_0),.dinb(n590),.dout(w_dff_A_3k4lhRIx4_2),.clk(gclk));
	jand g0527(.dina(w_n571_0[1]),.dinb(w_n565_0[0]),.dout(n599),.clk(gclk));
	jnot g0528(.din(n599),.dout(n600),.clk(gclk));
	jand g0529(.dina(w_n550_0[0]),.dinb(w_G45_1[0]),.dout(n601),.clk(gclk));
	jor g0530(.dina(n601),.dinb(w_n113_1[0]),.dout(n602),.clk(gclk));
	jnot g0531(.din(w_n602_0[1]),.dout(n603),.clk(gclk));
	jand g0532(.dina(w_n603_2[1]),.dinb(w_n592_2[0]),.dout(n604),.clk(gclk));
	jnot g0533(.din(w_n604_2[1]),.dout(n605),.clk(gclk));
	jand g0534(.dina(w_n605_1[2]),.dinb(w_n572_0[1]),.dout(n606),.clk(gclk));
	jand g0535(.dina(n606),.dinb(n600),.dout(n607),.clk(gclk));
	jand g0536(.dina(w_n462_0[0]),.dinb(w_n114_0[1]),.dout(n608),.clk(gclk));
	jand g0537(.dina(w_n608_1[2]),.dinb(w_n571_0[0]),.dout(n609),.clk(gclk));
	jnot g0538(.din(n609),.dout(n610),.clk(gclk));
	jand g0539(.dina(w_n146_1[0]),.dinb(w_G20_3[1]),.dout(n611),.clk(gclk));
	jor g0540(.dina(n611),.dinb(w_n115_0[1]),.dout(n612),.clk(gclk));
	jand g0541(.dina(w_G179_0[2]),.dinb(w_G20_3[0]),.dout(n613),.clk(gclk));
	jnot g0542(.din(w_n613_1[1]),.dout(n614),.clk(gclk));
	jand g0543(.dina(w_G200_2[0]),.dinb(w_G20_2[2]),.dout(n615),.clk(gclk));
	jand g0544(.dina(w_n615_0[1]),.dinb(n614),.dout(n616),.clk(gclk));
	jand g0545(.dina(w_n616_0[1]),.dinb(w_G190_2[0]),.dout(n617),.clk(gclk));
	jand g0546(.dina(w_n617_6[1]),.dinb(w_G303_2[1]),.dout(n618),.clk(gclk));
	jand g0547(.dina(w_n407_1[2]),.dinb(w_G20_2[1]),.dout(n619),.clk(gclk));
	jnot g0548(.din(w_n619_0[1]),.dout(n620),.clk(gclk));
	jor g0549(.dina(w_n615_0[0]),.dinb(w_n613_1[0]),.dout(n621),.clk(gclk));
	jnot g0550(.din(n621),.dout(n622),.clk(gclk));
	jand g0551(.dina(w_n622_0[1]),.dinb(n620),.dout(n623),.clk(gclk));
	jand g0552(.dina(w_n623_5[1]),.dinb(w_G294_3[0]),.dout(n624),.clk(gclk));
	jnot g0553(.din(w_G200_1[2]),.dout(n625),.clk(gclk));
	jand g0554(.dina(w_n613_0[2]),.dinb(n625),.dout(n626),.clk(gclk));
	jand g0555(.dina(w_n626_0[1]),.dinb(w_G190_1[2]),.dout(n627),.clk(gclk));
	jand g0556(.dina(w_n627_7[1]),.dinb(w_G322_0[2]),.dout(n628),.clk(gclk));
	jor g0557(.dina(w_dff_B_SEmiHP4u7_0),.dinb(n624),.dout(n629),.clk(gclk));
	jor g0558(.dina(n629),.dinb(w_dff_B_csnaLUaJ0_1),.dout(n630),.clk(gclk));
	jand g0559(.dina(w_n622_0[0]),.dinb(w_n619_0[0]),.dout(n631),.clk(gclk));
	jand g0560(.dina(w_n631_7[1]),.dinb(w_dff_B_fa6AkwhY3_1),.dout(n632),.clk(gclk));
	jor g0561(.dina(n632),.dinb(w_n148_5[2]),.dout(n633),.clk(gclk));
	jand g0562(.dina(w_n616_0[0]),.dinb(w_n407_1[1]),.dout(n634),.clk(gclk));
	jand g0563(.dina(w_n634_4[1]),.dinb(w_G283_3[1]),.dout(n635),.clk(gclk));
	jand g0564(.dina(w_n626_0[0]),.dinb(w_n407_1[0]),.dout(n636),.clk(gclk));
	jand g0565(.dina(w_n636_7[1]),.dinb(w_G311_1[2]),.dout(n637),.clk(gclk));
	jor g0566(.dina(w_dff_B_nxT6o9XU7_0),.dinb(n635),.dout(n638),.clk(gclk));
	jand g0567(.dina(w_n613_0[1]),.dinb(w_G200_1[1]),.dout(n639),.clk(gclk));
	jand g0568(.dina(w_n639_0[1]),.dinb(w_G190_1[1]),.dout(n640),.clk(gclk));
	jand g0569(.dina(w_n640_7[1]),.dinb(w_G326_0[1]),.dout(n641),.clk(gclk));
	jand g0570(.dina(w_n639_0[0]),.dinb(w_n407_0[2]),.dout(n642),.clk(gclk));
	jand g0571(.dina(w_n642_7[1]),.dinb(w_G317_1[1]),.dout(n643),.clk(gclk));
	jor g0572(.dina(n643),.dinb(n641),.dout(n644),.clk(gclk));
	jor g0573(.dina(w_dff_B_ItcZGkKB8_0),.dinb(n638),.dout(n645),.clk(gclk));
	jor g0574(.dina(n645),.dinb(w_dff_B_Gc1DhZXX9_1),.dout(n646),.clk(gclk));
	jor g0575(.dina(n646),.dinb(w_dff_B_gkg3k09p5_1),.dout(n647),.clk(gclk));
	jand g0576(.dina(w_n631_7[0]),.dinb(w_G159_3[1]),.dout(n648),.clk(gclk));
	jand g0577(.dina(w_n640_7[0]),.dinb(w_G50_4[0]),.dout(n649),.clk(gclk));
	jand g0578(.dina(w_n642_7[0]),.dinb(w_G68_3[2]),.dout(n650),.clk(gclk));
	jor g0579(.dina(n650),.dinb(n649),.dout(n651),.clk(gclk));
	jor g0580(.dina(n651),.dinb(n648),.dout(n652),.clk(gclk));
	jnot g0581(.din(n652),.dout(n653),.clk(gclk));
	jand g0582(.dina(w_n617_6[0]),.dinb(w_G87_2[1]),.dout(n654),.clk(gclk));
	jnot g0583(.din(w_n654_0[1]),.dout(n655),.clk(gclk));
	jand g0584(.dina(n655),.dinb(w_n148_5[1]),.dout(n656),.clk(gclk));
	jand g0585(.dina(w_n634_4[0]),.dinb(w_G107_3[1]),.dout(n657),.clk(gclk));
	jand g0586(.dina(w_n636_7[0]),.dinb(w_G77_3[1]),.dout(n658),.clk(gclk));
	jor g0587(.dina(w_dff_B_hLJtlJJF9_0),.dinb(w_n657_0[1]),.dout(n659),.clk(gclk));
	jand g0588(.dina(w_n627_7[0]),.dinb(w_G58_3[2]),.dout(n660),.clk(gclk));
	jand g0589(.dina(w_n623_5[0]),.dinb(w_G97_3[1]),.dout(n661),.clk(gclk));
	jor g0590(.dina(w_n661_0[1]),.dinb(w_dff_B_XCGnxZHc1_1),.dout(n662),.clk(gclk));
	jor g0591(.dina(n662),.dinb(n659),.dout(n663),.clk(gclk));
	jnot g0592(.din(n663),.dout(n664),.clk(gclk));
	jand g0593(.dina(n664),.dinb(w_dff_B_JttXkiGp9_1),.dout(n665),.clk(gclk));
	jand g0594(.dina(n665),.dinb(w_dff_B_hSFoL9Vx7_1),.dout(n666),.clk(gclk));
	jnot g0595(.din(n666),.dout(n667),.clk(gclk));
	jand g0596(.dina(n667),.dinb(w_dff_B_h10GtyIo3_1),.dout(n668),.clk(gclk));
	jor g0597(.dina(n668),.dinb(w_n612_4[1]),.dout(n669),.clk(gclk));
	jnot g0598(.din(w_n608_1[1]),.dout(n670),.clk(gclk));
	jand g0599(.dina(w_n612_4[0]),.dinb(n670),.dout(n671),.clk(gclk));
	jnot g0600(.din(n671),.dout(n672),.clk(gclk));
	jand g0601(.dina(w_n140_0[0]),.dinb(w_G45_0[2]),.dout(n673),.clk(gclk));
	jand g0602(.dina(w_n118_0[0]),.dinb(w_n161_0[2]),.dout(n674),.clk(gclk));
	jand g0603(.dina(w_n122_0[2]),.dinb(w_G33_6[1]),.dout(n675),.clk(gclk));
	jnot g0604(.din(w_n675_0[2]),.dout(n676),.clk(gclk));
	jor g0605(.dina(w_n676_0[1]),.dinb(n674),.dout(n677),.clk(gclk));
	jor g0606(.dina(n677),.dinb(w_dff_B_z7x30knv6_1),.dout(n678),.clk(gclk));
	jand g0607(.dina(w_n123_1[1]),.dinb(w_n105_0[2]),.dout(n679),.clk(gclk));
	jand g0608(.dina(w_n122_0[1]),.dinb(w_n148_5[0]),.dout(n680),.clk(gclk));
	jand g0609(.dina(w_n680_0[1]),.dinb(w_G355_0),.dout(n681),.clk(gclk));
	jor g0610(.dina(n681),.dinb(w_dff_B_t9fHK07t4_1),.dout(n682),.clk(gclk));
	jnot g0611(.din(n682),.dout(n683),.clk(gclk));
	jand g0612(.dina(n683),.dinb(w_dff_B_T07KtoY26_1),.dout(n684),.clk(gclk));
	jor g0613(.dina(n684),.dinb(w_n672_1[1]),.dout(n685),.clk(gclk));
	jand g0614(.dina(n685),.dinb(w_n604_2[0]),.dout(n686),.clk(gclk));
	jand g0615(.dina(w_dff_B_AqESJkoR8_0),.dinb(n669),.dout(n687),.clk(gclk));
	jand g0616(.dina(w_dff_B_XBhVLbD39_0),.dinb(n610),.dout(n688),.clk(gclk));
	jor g0617(.dina(n688),.dinb(n607),.dout(G396_fa_),.clk(gclk));
	jnot g0618(.din(w_n588_1[0]),.dout(n690),.clk(gclk));
	jnot g0619(.din(w_n401_0[0]),.dout(n691),.clk(gclk));
	jor g0620(.dina(w_n554_2[0]),.dinb(n691),.dout(n692),.clk(gclk));
	jand g0621(.dina(w_n692_0[1]),.dinb(w_n412_0[0]),.dout(n693),.clk(gclk));
	jor g0622(.dina(w_n692_0[0]),.dinb(w_n405_0[0]),.dout(n694),.clk(gclk));
	jnot g0623(.din(n694),.dout(n695),.clk(gclk));
	jor g0624(.dina(n695),.dinb(n693),.dout(n696),.clk(gclk));
	jxor g0625(.dina(w_n696_1[2]),.dinb(w_n576_1[0]),.dout(n697),.clk(gclk));
	jnot g0626(.din(n697),.dout(n698),.clk(gclk));
	jand g0627(.dina(n698),.dinb(w_dff_B_jnmeR2JH2_1),.dout(n699),.clk(gclk));
	jor g0628(.dina(w_n991_0[2]),.dinb(w_n604_1[2]),.dout(n701),.clk(gclk));
	jor g0629(.dina(w_dff_B_sOUDt0Jw2_0),.dinb(n699),.dout(n702),.clk(gclk));
	jnot g0630(.din(w_n696_1[1]),.dout(n703),.clk(gclk));
	jand g0631(.dina(n703),.dinb(w_n425_1[1]),.dout(n704),.clk(gclk));
	jnot g0632(.din(n704),.dout(n705),.clk(gclk));
	jand g0633(.dina(w_n631_6[2]),.dinb(w_G132_1[1]),.dout(n706),.clk(gclk));
	jand g0634(.dina(w_n623_4[2]),.dinb(w_G58_3[1]),.dout(n707),.clk(gclk));
	jand g0635(.dina(w_n642_6[2]),.dinb(w_G150_3[0]),.dout(n708),.clk(gclk));
	jor g0636(.dina(w_dff_B_VXotR1C14_0),.dinb(n707),.dout(n709),.clk(gclk));
	jor g0637(.dina(n709),.dinb(w_dff_B_YOTbRa345_1),.dout(n710),.clk(gclk));
	jand g0638(.dina(w_n617_5[2]),.dinb(w_G50_3[2]),.dout(n711),.clk(gclk));
	jor g0639(.dina(n711),.dinb(w_G33_6[0]),.dout(n712),.clk(gclk));
	jand g0640(.dina(w_n636_6[2]),.dinb(w_G159_3[0]),.dout(n713),.clk(gclk));
	jand g0641(.dina(w_n627_6[2]),.dinb(w_G143_2[1]),.dout(n714),.clk(gclk));
	jor g0642(.dina(n714),.dinb(n713),.dout(n715),.clk(gclk));
	jand g0643(.dina(w_n640_6[2]),.dinb(w_G137_1[2]),.dout(n716),.clk(gclk));
	jand g0644(.dina(w_n634_3[2]),.dinb(w_G68_3[1]),.dout(n717),.clk(gclk));
	jor g0645(.dina(w_n717_0[1]),.dinb(w_dff_B_jVLjZUPy4_1),.dout(n718),.clk(gclk));
	jor g0646(.dina(n718),.dinb(w_dff_B_r2gcMh6c5_1),.dout(n719),.clk(gclk));
	jor g0647(.dina(n719),.dinb(w_dff_B_TVNJnW056_1),.dout(n720),.clk(gclk));
	jor g0648(.dina(n720),.dinb(w_dff_B_XrhrrlvU0_1),.dout(n721),.clk(gclk));
	jand g0649(.dina(w_n631_6[1]),.dinb(w_G311_1[1]),.dout(n722),.clk(gclk));
	jand g0650(.dina(w_n617_5[1]),.dinb(w_G107_3[0]),.dout(n723),.clk(gclk));
	jand g0651(.dina(w_n642_6[1]),.dinb(w_G283_3[0]),.dout(n724),.clk(gclk));
	jor g0652(.dina(w_dff_B_bHxLWWnm0_0),.dinb(n723),.dout(n725),.clk(gclk));
	jor g0653(.dina(n725),.dinb(w_dff_B_1L2my1Ce8_1),.dout(n726),.clk(gclk));
	jnot g0654(.din(n726),.dout(n727),.clk(gclk));
	jand g0655(.dina(w_n634_3[1]),.dinb(w_G87_2[0]),.dout(n728),.clk(gclk));
	jnot g0656(.din(w_n728_0[1]),.dout(n729),.clk(gclk));
	jand g0657(.dina(n729),.dinb(w_G33_5[2]),.dout(n730),.clk(gclk));
	jand g0658(.dina(w_n636_6[1]),.dinb(w_G116_3[2]),.dout(n731),.clk(gclk));
	jand g0659(.dina(w_n627_6[1]),.dinb(w_G294_2[2]),.dout(n732),.clk(gclk));
	jor g0660(.dina(n732),.dinb(n731),.dout(n733),.clk(gclk));
	jand g0661(.dina(w_n640_6[1]),.dinb(w_G303_2[0]),.dout(n734),.clk(gclk));
	jor g0662(.dina(w_dff_B_ipLwlcnj3_0),.dinb(w_n661_0[0]),.dout(n735),.clk(gclk));
	jor g0663(.dina(n735),.dinb(w_dff_B_BzC8fKGl8_1),.dout(n736),.clk(gclk));
	jnot g0664(.din(n736),.dout(n737),.clk(gclk));
	jand g0665(.dina(n737),.dinb(w_dff_B_oi0MVyjt8_1),.dout(n738),.clk(gclk));
	jand g0666(.dina(n738),.dinb(w_dff_B_DDUVIJFg5_1),.dout(n739),.clk(gclk));
	jnot g0667(.din(n739),.dout(n740),.clk(gclk));
	jand g0668(.dina(n740),.dinb(w_dff_B_FVLNdNhN9_1),.dout(n741),.clk(gclk));
	jor g0669(.dina(n741),.dinb(w_n612_3[2]),.dout(n742),.clk(gclk));
	jand g0670(.dina(w_n612_3[1]),.dinb(w_n426_0[0]),.dout(n743),.clk(gclk));
	jand g0671(.dina(w_n743_1[1]),.dinb(w_n72_0[1]),.dout(n744),.clk(gclk));
	jor g0672(.dina(w_dff_B_Ppn9qytr3_0),.dinb(w_n605_1[1]),.dout(n745),.clk(gclk));
	jnot g0673(.din(n745),.dout(n746),.clk(gclk));
	jand g0674(.dina(w_dff_B_8PHEd5ke3_0),.dinb(n742),.dout(n747),.clk(gclk));
	jand g0675(.dina(w_dff_B_r4LG1yPQ1_0),.dinb(n705),.dout(n748),.clk(gclk));
	jnot g0676(.din(n748),.dout(n749),.clk(gclk));
	jand g0677(.dina(n749),.dinb(n702),.dout(n750),.clk(gclk));
	jnot g0678(.din(w_n750_0[1]),.dout(G384_fa_),.clk(gclk));
	jnot g0679(.din(w_n552_1[0]),.dout(n752),.clk(gclk));
	jand g0680(.dina(w_dff_B_HpupBuZ24_0),.dinb(w_n542_0[1]),.dout(n753),.clk(gclk));
	jand g0681(.dina(w_n552_0[2]),.dinb(w_n512_0[0]),.dout(n754),.clk(gclk));
	jnot g0682(.din(w_n754_0[1]),.dout(n755),.clk(gclk));
	jand g0683(.dina(n755),.dinb(w_n517_0[0]),.dout(n756),.clk(gclk));
	jand g0684(.dina(w_n754_0[0]),.dinb(w_n542_0[0]),.dout(n757),.clk(gclk));
	jor g0685(.dina(n757),.dinb(n756),.dout(n758),.clk(gclk));
	jand g0686(.dina(w_n696_1[0]),.dinb(w_n576_0[2]),.dout(n759),.clk(gclk));
	jand g0687(.dina(w_n553_1[2]),.dinb(w_n436_0[0]),.dout(n760),.clk(gclk));
	jnot g0688(.din(w_n760_0[1]),.dout(n761),.clk(gclk));
	jand g0689(.dina(w_dff_B_sc5ECryo4_0),.dinb(w_n446_0[0]),.dout(n762),.clk(gclk));
	jand g0690(.dina(w_n760_0[0]),.dinb(w_n439_0[2]),.dout(n763),.clk(gclk));
	jor g0691(.dina(w_dff_B_cPx4GLvs2_0),.dinb(n762),.dout(n764),.clk(gclk));
	jand g0692(.dina(w_n764_1[2]),.dinb(w_n759_0[1]),.dout(n765),.clk(gclk));
	jor g0693(.dina(w_n764_1[1]),.dinb(w_n439_0[1]),.dout(n766),.clk(gclk));
	jand g0694(.dina(w_n554_1[2]),.dinb(w_n543_0[0]),.dout(n767),.clk(gclk));
	jand g0695(.dina(w_dff_B_CPQM883m4_0),.dinb(n766),.dout(n768),.clk(gclk));
	jor g0696(.dina(w_dff_B_6QtczEZz2_0),.dinb(n765),.dout(n769),.clk(gclk));
	jand g0697(.dina(w_n769_0[1]),.dinb(w_n758_1[1]),.dout(n770),.clk(gclk));
	jor g0698(.dina(n770),.dinb(w_dff_B_2wUF6utT3_1),.dout(n771),.clk(gclk));
	jnot g0699(.din(w_n771_0[2]),.dout(n772),.clk(gclk));
	jand g0700(.dina(w_n576_0[1]),.dinb(w_n519_1[0]),.dout(n773),.clk(gclk));
	jor g0701(.dina(n773),.dinb(w_n548_0[1]),.dout(n774),.clk(gclk));
	jand g0702(.dina(w_n764_1[0]),.dinb(w_n696_0[2]),.dout(n775),.clk(gclk));
	jand g0703(.dina(n775),.dinb(w_n758_1[0]),.dout(n776),.clk(gclk));
	jxor g0704(.dina(n776),.dinb(w_n519_0[2]),.dout(n777),.clk(gclk));
	jand g0705(.dina(n777),.dinb(w_n588_0[2]),.dout(n778),.clk(gclk));
	jxor g0706(.dina(n778),.dinb(w_dff_B_meZ7zUbD1_1),.dout(n779),.clk(gclk));
	jnot g0707(.din(w_n779_0[1]),.dout(n780),.clk(gclk));
	jor g0708(.dina(w_dff_B_6KOFtQeg5_0),.dinb(n772),.dout(n781),.clk(gclk));
	jor g0709(.dina(w_n779_0[0]),.dinb(w_n771_0[1]),.dout(n782),.clk(gclk));
	jnot g0710(.din(w_n121_0[1]),.dout(n783),.clk(gclk));
	jand g0711(.dina(n783),.dinb(w_n116_0[0]),.dout(n784),.clk(gclk));
	jand g0712(.dina(w_dff_B_bvj5x9wr1_0),.dinb(n782),.dout(n785),.clk(gclk));
	jand g0713(.dina(n785),.dinb(n781),.dout(n786),.clk(gclk));
	jand g0714(.dina(w_G77_3[0]),.dinb(w_G50_3[1]),.dout(n787),.clk(gclk));
	jand g0715(.dina(n787),.dinb(w_n137_0[0]),.dout(n788),.clk(gclk));
	jand g0716(.dina(w_G68_3[0]),.dinb(w_n73_1[2]),.dout(n789),.clk(gclk));
	jor g0717(.dina(n789),.dinb(n788),.dout(n790),.clk(gclk));
	jand g0718(.dina(n790),.dinb(w_n121_0[0]),.dout(n791),.clk(gclk));
	jnot g0719(.din(w_n255_0[0]),.dout(n792),.clk(gclk));
	jand g0720(.dina(w_n147_0[0]),.dinb(w_G116_3[1]),.dout(n793),.clk(gclk));
	jand g0721(.dina(w_dff_B_LsPz2THP9_0),.dinb(n792),.dout(n794),.clk(gclk));
	jor g0722(.dina(n794),.dinb(w_dff_B_07cq4XHF0_1),.dout(n795),.clk(gclk));
	jor g0723(.dina(w_dff_B_qqINFvwM6_0),.dinb(n786),.dout(w_dff_A_FbrOxECu5_2),.clk(gclk));
	jand g0724(.dina(w_n553_1[1]),.dinb(w_n214_0[0]),.dout(n797),.clk(gclk));
	jnot g0725(.din(w_n797_0[1]),.dout(n798),.clk(gclk));
	jand g0726(.dina(w_dff_B_jj7AxzEY2_0),.dinb(w_n219_0[0]),.dout(n799),.clk(gclk));
	jand g0727(.dina(w_n797_0[0]),.dinb(w_n532_0[0]),.dout(n800),.clk(gclk));
	jor g0728(.dina(w_dff_B_IhUb9nu18_0),.dinb(n799),.dout(n801),.clk(gclk));
	jnot g0729(.din(w_n801_0[1]),.dout(n802),.clk(gclk));
	jand g0730(.dina(n802),.dinb(w_n608_1[0]),.dout(n803),.clk(gclk));
	jnot g0731(.din(n803),.dout(n804),.clk(gclk));
	jand g0732(.dina(w_n631_6[0]),.dinb(w_G317_1[0]),.dout(n805),.clk(gclk));
	jand g0733(.dina(w_n623_4[1]),.dinb(w_G107_2[2]),.dout(n806),.clk(gclk));
	jand g0734(.dina(w_n642_6[0]),.dinb(w_G294_2[1]),.dout(n807),.clk(gclk));
	jor g0735(.dina(w_dff_B_JiIMEmpI1_0),.dinb(n806),.dout(n808),.clk(gclk));
	jor g0736(.dina(n808),.dinb(w_dff_B_icDZmfxm3_1),.dout(n809),.clk(gclk));
	jand g0737(.dina(w_n617_5[0]),.dinb(w_G116_3[0]),.dout(n810),.clk(gclk));
	jor g0738(.dina(n810),.dinb(w_n148_4[2]),.dout(n811),.clk(gclk));
	jand g0739(.dina(w_n636_6[0]),.dinb(w_G283_2[2]),.dout(n812),.clk(gclk));
	jand g0740(.dina(w_n627_6[0]),.dinb(w_G303_1[2]),.dout(n813),.clk(gclk));
	jor g0741(.dina(n813),.dinb(n812),.dout(n814),.clk(gclk));
	jand g0742(.dina(w_n640_6[0]),.dinb(w_G311_1[0]),.dout(n815),.clk(gclk));
	jand g0743(.dina(w_n634_3[0]),.dinb(w_G97_3[0]),.dout(n816),.clk(gclk));
	jor g0744(.dina(w_n816_0[1]),.dinb(w_dff_B_E3kh8RIO8_1),.dout(n817),.clk(gclk));
	jor g0745(.dina(n817),.dinb(w_dff_B_aLyvrF5y2_1),.dout(n818),.clk(gclk));
	jor g0746(.dina(n818),.dinb(w_dff_B_60dAyajg5_1),.dout(n819),.clk(gclk));
	jor g0747(.dina(n819),.dinb(w_dff_B_o7ogLalW2_1),.dout(n820),.clk(gclk));
	jand g0748(.dina(w_n631_5[2]),.dinb(w_G137_1[1]),.dout(n821),.clk(gclk));
	jnot g0749(.din(n821),.dout(n822),.clk(gclk));
	jand g0750(.dina(w_n623_4[0]),.dinb(w_G68_2[2]),.dout(n823),.clk(gclk));
	jnot g0751(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jand g0752(.dina(w_n634_2[2]),.dinb(w_G77_2[2]),.dout(n825),.clk(gclk));
	jnot g0753(.din(w_n825_0[1]),.dout(n826),.clk(gclk));
	jand g0754(.dina(n826),.dinb(n824),.dout(n827),.clk(gclk));
	jand g0755(.dina(n827),.dinb(w_dff_B_XDbCX56u3_1),.dout(n828),.clk(gclk));
	jand g0756(.dina(w_n642_5[2]),.dinb(w_G159_2[2]),.dout(n829),.clk(gclk));
	jor g0757(.dina(n829),.dinb(w_G33_5[1]),.dout(n830),.clk(gclk));
	jand g0758(.dina(w_n640_5[2]),.dinb(w_G143_2[0]),.dout(n831),.clk(gclk));
	jand g0759(.dina(w_n627_5[2]),.dinb(w_G150_2[2]),.dout(n832),.clk(gclk));
	jor g0760(.dina(n832),.dinb(n831),.dout(n833),.clk(gclk));
	jand g0761(.dina(w_n636_5[2]),.dinb(w_G50_3[0]),.dout(n834),.clk(gclk));
	jand g0762(.dina(w_n617_4[2]),.dinb(w_G58_3[0]),.dout(n835),.clk(gclk));
	jor g0763(.dina(n835),.dinb(w_dff_B_VokvmHoW1_1),.dout(n836),.clk(gclk));
	jor g0764(.dina(n836),.dinb(w_dff_B_9KRSL5N54_1),.dout(n837),.clk(gclk));
	jor g0765(.dina(n837),.dinb(w_dff_B_41U9DHKJ6_1),.dout(n838),.clk(gclk));
	jnot g0766(.din(n838),.dout(n839),.clk(gclk));
	jand g0767(.dina(n839),.dinb(w_dff_B_jB04fN5o7_1),.dout(n840),.clk(gclk));
	jnot g0768(.din(n840),.dout(n841),.clk(gclk));
	jand g0769(.dina(n841),.dinb(w_dff_B_MPZkSopX3_1),.dout(n842),.clk(gclk));
	jor g0770(.dina(n842),.dinb(w_n612_3[0]),.dout(n843),.clk(gclk));
	jand g0771(.dina(w_n675_0[1]),.dinb(w_n131_0[0]),.dout(n844),.clk(gclk));
	jand g0772(.dina(w_n123_1[0]),.dinb(w_G87_1[2]),.dout(n845),.clk(gclk));
	jor g0773(.dina(w_dff_B_SfLpZ49O7_0),.dinb(w_n672_1[0]),.dout(n846),.clk(gclk));
	jor g0774(.dina(n846),.dinb(w_dff_B_6RDoPbTe0_1),.dout(n847),.clk(gclk));
	jand g0775(.dina(n847),.dinb(w_n604_1[1]),.dout(n848),.clk(gclk));
	jand g0776(.dina(w_dff_B_4csAsGzu2_0),.dinb(n843),.dout(n849),.clk(gclk));
	jand g0777(.dina(w_dff_B_lMaU6M2E7_0),.dinb(n804),.dout(n850),.clk(gclk));
	jnot g0778(.din(w_n589_1[1]),.dout(n851),.clk(gclk));
	jxor g0779(.dina(w_n561_0[0]),.dinb(w_n556_0[0]),.dout(n852),.clk(gclk));
	jxor g0780(.dina(w_dff_B_QKGI8h3V0_0),.dinb(w_n572_0[0]),.dout(n853),.clk(gclk));
	jnot g0781(.din(w_n853_0[2]),.dout(n854),.clk(gclk));
	jand g0782(.dina(n854),.dinb(n851),.dout(n855),.clk(gclk));
	jnot g0783(.din(w_n278_0[0]),.dout(n856),.clk(gclk));
	jand g0784(.dina(w_n553_1[0]),.dinb(w_n274_0[0]),.dout(n857),.clk(gclk));
	jor g0785(.dina(w_dff_B_izibPMR73_0),.dinb(n856),.dout(n858),.clk(gclk));
	jand g0786(.dina(w_n553_0[2]),.dinb(w_n536_0[1]),.dout(n859),.clk(gclk));
	jnot g0787(.din(n859),.dout(n860),.clk(gclk));
	jand g0788(.dina(w_dff_B_91mPsrla4_0),.dinb(n858),.dout(n861),.clk(gclk));
	jxor g0789(.dina(w_n861_1[1]),.dinb(w_n573_0[1]),.dout(n862),.clk(gclk));
	jxor g0790(.dina(n862),.dinb(w_n563_0[1]),.dout(n863),.clk(gclk));
	jand g0791(.dina(w_n863_0[1]),.dinb(w_n855_0[2]),.dout(n864),.clk(gclk));
	jor g0792(.dina(w_n864_0[1]),.dinb(w_n589_1[0]),.dout(n865),.clk(gclk));
	jand g0793(.dina(n865),.dinb(w_n591_0[2]),.dout(n866),.clk(gclk));
	jor g0794(.dina(n866),.dinb(w_n602_0[0]),.dout(n867),.clk(gclk));
	jand g0795(.dina(w_n554_1[1]),.dinb(w_n536_0[0]),.dout(n868),.clk(gclk));
	jnot g0796(.din(w_n861_1[0]),.dout(n869),.clk(gclk));
	jand g0797(.dina(n869),.dinb(w_n563_0[0]),.dout(n870),.clk(gclk));
	jor g0798(.dina(n870),.dinb(w_dff_B_RgDzYCTb1_1),.dout(n871),.clk(gclk));
	jor g0799(.dina(w_n861_0[2]),.dinb(w_n573_0[0]),.dout(n872),.clk(gclk));
	jxor g0800(.dina(n872),.dinb(w_n801_0[0]),.dout(n873),.clk(gclk));
	jxor g0801(.dina(n873),.dinb(w_dff_B_EVI7LtAT4_1),.dout(n874),.clk(gclk));
	jnot g0802(.din(n874),.dout(n875),.clk(gclk));
	jand g0803(.dina(w_dff_B_JUvPulu93_0),.dinb(n867),.dout(n876),.clk(gclk));
	jor g0804(.dina(n876),.dinb(w_dff_B_Bt9QAkTd5_1),.dout(G387_fa_),.clk(gclk));
	jand g0805(.dina(w_n853_0[1]),.dinb(w_n589_0[2]),.dout(n878),.clk(gclk));
	jor g0806(.dina(w_n855_0[1]),.dinb(w_n592_1[2]),.dout(n879),.clk(gclk));
	jor g0807(.dina(n879),.dinb(w_dff_B_CwgtMlEH9_1),.dout(n880),.clk(gclk));
	jor g0808(.dina(w_n853_0[0]),.dinb(w_n603_2[0]),.dout(n881),.clk(gclk));
	jand g0809(.dina(w_n608_0[2]),.dinb(w_n564_0[0]),.dout(n882),.clk(gclk));
	jand g0810(.dina(w_n631_5[1]),.dinb(w_G326_0[0]),.dout(n883),.clk(gclk));
	jand g0811(.dina(w_n623_3[2]),.dinb(w_G283_2[1]),.dout(n884),.clk(gclk));
	jand g0812(.dina(w_n627_5[1]),.dinb(w_G317_0[2]),.dout(n885),.clk(gclk));
	jor g0813(.dina(w_dff_B_umOvivqc3_0),.dinb(n884),.dout(n886),.clk(gclk));
	jor g0814(.dina(n886),.dinb(w_dff_B_r4P1rwqF3_1),.dout(n887),.clk(gclk));
	jand g0815(.dina(w_n617_4[1]),.dinb(w_G294_2[0]),.dout(n888),.clk(gclk));
	jor g0816(.dina(n888),.dinb(w_n148_4[1]),.dout(n889),.clk(gclk));
	jand g0817(.dina(w_n634_2[1]),.dinb(w_G116_2[2]),.dout(n890),.clk(gclk));
	jand g0818(.dina(w_n636_5[1]),.dinb(w_G303_1[1]),.dout(n891),.clk(gclk));
	jor g0819(.dina(w_dff_B_TYKlVe3n2_0),.dinb(n890),.dout(n892),.clk(gclk));
	jand g0820(.dina(w_n640_5[1]),.dinb(w_G322_0[1]),.dout(n893),.clk(gclk));
	jand g0821(.dina(w_n642_5[1]),.dinb(w_G311_0[2]),.dout(n894),.clk(gclk));
	jor g0822(.dina(n894),.dinb(n893),.dout(n895),.clk(gclk));
	jor g0823(.dina(w_dff_B_imB7NkY34_0),.dinb(n892),.dout(n896),.clk(gclk));
	jor g0824(.dina(n896),.dinb(w_dff_B_SfGEYDQO1_1),.dout(n897),.clk(gclk));
	jor g0825(.dina(n897),.dinb(w_dff_B_RxDJlPs49_1),.dout(n898),.clk(gclk));
	jand g0826(.dina(w_n623_3[1]),.dinb(w_G87_1[1]),.dout(n899),.clk(gclk));
	jand g0827(.dina(w_n642_5[0]),.dinb(w_G58_2[2]),.dout(n900),.clk(gclk));
	jor g0828(.dina(w_dff_B_jijveFSS1_0),.dinb(w_n816_0[0]),.dout(n901),.clk(gclk));
	jor g0829(.dina(n901),.dinb(w_n899_0[1]),.dout(n902),.clk(gclk));
	jand g0830(.dina(w_n631_5[0]),.dinb(w_G150_2[1]),.dout(n903),.clk(gclk));
	jor g0831(.dina(n903),.dinb(w_G33_5[0]),.dout(n904),.clk(gclk));
	jand g0832(.dina(w_n640_5[0]),.dinb(w_G159_2[1]),.dout(n905),.clk(gclk));
	jand g0833(.dina(w_n636_5[0]),.dinb(w_G68_2[1]),.dout(n906),.clk(gclk));
	jor g0834(.dina(n906),.dinb(n905),.dout(n907),.clk(gclk));
	jand g0835(.dina(w_n627_5[0]),.dinb(w_G50_2[2]),.dout(n908),.clk(gclk));
	jand g0836(.dina(w_n617_4[0]),.dinb(w_G77_2[1]),.dout(n909),.clk(gclk));
	jor g0837(.dina(w_n909_0[1]),.dinb(w_dff_B_gz7dj8DM7_1),.dout(n910),.clk(gclk));
	jor g0838(.dina(n910),.dinb(w_dff_B_FFFNZjvU1_1),.dout(n911),.clk(gclk));
	jor g0839(.dina(n911),.dinb(w_dff_B_AyWMX6dN8_1),.dout(n912),.clk(gclk));
	jor g0840(.dina(n912),.dinb(w_dff_B_WnKyF0ti2_1),.dout(n913),.clk(gclk));
	jand g0841(.dina(n913),.dinb(n898),.dout(n914),.clk(gclk));
	jor g0842(.dina(n914),.dinb(w_n612_2[2]),.dout(n915),.clk(gclk));
	jand g0843(.dina(w_n135_0[0]),.dinb(w_G45_0[1]),.dout(n916),.clk(gclk));
	jand g0844(.dina(w_G77_2[0]),.dinb(w_G68_2[0]),.dout(n917),.clk(gclk));
	jnot g0845(.din(n917),.dout(n918),.clk(gclk));
	jand g0846(.dina(w_G58_2[1]),.dinb(w_n161_0[1]),.dout(n919),.clk(gclk));
	jand g0847(.dina(n919),.dinb(w_n73_1[1]),.dout(n920),.clk(gclk));
	jand g0848(.dina(n920),.dinb(w_dff_B_BFovSasJ9_1),.dout(n921),.clk(gclk));
	jand g0849(.dina(n921),.dinb(w_n593_0[1]),.dout(n922),.clk(gclk));
	jor g0850(.dina(n922),.dinb(w_n676_0[0]),.dout(n923),.clk(gclk));
	jor g0851(.dina(n923),.dinb(w_dff_B_7KrCzawj1_1),.dout(n924),.clk(gclk));
	jand g0852(.dina(w_n123_0[2]),.dinb(w_n80_0[1]),.dout(n925),.clk(gclk));
	jnot g0853(.din(w_n593_0[0]),.dout(n926),.clk(gclk));
	jand g0854(.dina(w_n680_0[0]),.dinb(n926),.dout(n927),.clk(gclk));
	jor g0855(.dina(n927),.dinb(w_dff_B_Wtje1SaE7_1),.dout(n928),.clk(gclk));
	jnot g0856(.din(n928),.dout(n929),.clk(gclk));
	jand g0857(.dina(n929),.dinb(w_dff_B_7vlzAMVs7_1),.dout(n930),.clk(gclk));
	jor g0858(.dina(n930),.dinb(w_n672_0[2]),.dout(n931),.clk(gclk));
	jand g0859(.dina(n931),.dinb(w_n604_1[0]),.dout(n932),.clk(gclk));
	jand g0860(.dina(n932),.dinb(n915),.dout(n933),.clk(gclk));
	jnot g0861(.din(n933),.dout(n934),.clk(gclk));
	jor g0862(.dina(w_dff_B_anfcVjYq8_0),.dinb(n882),.dout(n935),.clk(gclk));
	jand g0863(.dina(w_dff_B_pBuz2pDf9_0),.dinb(n881),.dout(n936),.clk(gclk));
	jand g0864(.dina(w_dff_B_xcyXUC0e7_0),.dinb(n880),.dout(n937),.clk(gclk));
	jnot g0865(.din(w_n937_0[2]),.dout(w_dff_A_VD26nmsp6_1),.clk(gclk));
	jnot g0866(.din(w_n855_0[0]),.dout(n939),.clk(gclk));
	jnot g0867(.din(w_n863_0[0]),.dout(n940),.clk(gclk));
	jand g0868(.dina(w_n940_0[1]),.dinb(n939),.dout(n941),.clk(gclk));
	jor g0869(.dina(w_n864_0[0]),.dinb(w_n592_1[1]),.dout(n942),.clk(gclk));
	jor g0870(.dina(n942),.dinb(n941),.dout(n943),.clk(gclk));
	jor g0871(.dina(w_n940_0[0]),.dinb(w_n603_1[2]),.dout(n944),.clk(gclk));
	jand g0872(.dina(w_n861_0[1]),.dinb(w_n608_0[1]),.dout(n945),.clk(gclk));
	jnot g0873(.din(n945),.dout(n946),.clk(gclk));
	jand g0874(.dina(w_n623_3[0]),.dinb(w_G116_2[1]),.dout(n947),.clk(gclk));
	jand g0875(.dina(w_n617_3[2]),.dinb(w_G283_2[0]),.dout(n948),.clk(gclk));
	jand g0876(.dina(w_n642_4[2]),.dinb(w_G303_1[0]),.dout(n949),.clk(gclk));
	jor g0877(.dina(w_dff_B_M0D7D2sP4_0),.dinb(n948),.dout(n950),.clk(gclk));
	jor g0878(.dina(n950),.dinb(w_dff_B_60i9nVvj7_1),.dout(n951),.clk(gclk));
	jand g0879(.dina(w_n631_4[2]),.dinb(w_G322_0[0]),.dout(n952),.clk(gclk));
	jor g0880(.dina(n952),.dinb(w_n148_4[0]),.dout(n953),.clk(gclk));
	jand g0881(.dina(w_n636_4[2]),.dinb(w_G294_1[2]),.dout(n954),.clk(gclk));
	jand g0882(.dina(w_n627_4[2]),.dinb(w_G311_0[1]),.dout(n955),.clk(gclk));
	jor g0883(.dina(n955),.dinb(n954),.dout(n956),.clk(gclk));
	jand g0884(.dina(w_n640_4[2]),.dinb(w_G317_0[1]),.dout(n957),.clk(gclk));
	jor g0885(.dina(w_dff_B_4bYsWbFL6_0),.dinb(w_n657_0[0]),.dout(n958),.clk(gclk));
	jor g0886(.dina(n958),.dinb(w_dff_B_1JNOJRPv9_1),.dout(n959),.clk(gclk));
	jor g0887(.dina(n959),.dinb(w_dff_B_2acrcGUW7_1),.dout(n960),.clk(gclk));
	jor g0888(.dina(n960),.dinb(w_dff_B_ivslArfX2_1),.dout(n961),.clk(gclk));
	jand g0889(.dina(w_n623_2[2]),.dinb(w_G77_1[2]),.dout(n962),.clk(gclk));
	jand g0890(.dina(w_n617_3[1]),.dinb(w_G68_1[2]),.dout(n963),.clk(gclk));
	jand g0891(.dina(w_n642_4[1]),.dinb(w_G50_2[1]),.dout(n964),.clk(gclk));
	jor g0892(.dina(w_dff_B_bTXCXE3W2_0),.dinb(n963),.dout(n965),.clk(gclk));
	jor g0893(.dina(n965),.dinb(w_n962_0[1]),.dout(n966),.clk(gclk));
	jand g0894(.dina(w_n631_4[1]),.dinb(w_G143_1[2]),.dout(n967),.clk(gclk));
	jor g0895(.dina(n967),.dinb(w_G33_4[2]),.dout(n968),.clk(gclk));
	jand g0896(.dina(w_n636_4[1]),.dinb(w_G58_2[0]),.dout(n969),.clk(gclk));
	jand g0897(.dina(w_n627_4[1]),.dinb(w_G159_2[0]),.dout(n970),.clk(gclk));
	jor g0898(.dina(n970),.dinb(n969),.dout(n971),.clk(gclk));
	jand g0899(.dina(w_n640_4[1]),.dinb(w_G150_2[0]),.dout(n972),.clk(gclk));
	jor g0900(.dina(w_dff_B_3vBlmhip4_0),.dinb(w_n728_0[0]),.dout(n973),.clk(gclk));
	jor g0901(.dina(n973),.dinb(w_dff_B_nXJrMS4Q5_1),.dout(n974),.clk(gclk));
	jor g0902(.dina(n974),.dinb(w_dff_B_7ZSJceom5_1),.dout(n975),.clk(gclk));
	jor g0903(.dina(n975),.dinb(w_dff_B_woEMQmxf1_1),.dout(n976),.clk(gclk));
	jand g0904(.dina(n976),.dinb(n961),.dout(n977),.clk(gclk));
	jor g0905(.dina(n977),.dinb(w_n612_2[1]),.dout(n978),.clk(gclk));
	jand g0906(.dina(w_n675_0[0]),.dinb(w_n144_0[0]),.dout(n979),.clk(gclk));
	jand g0907(.dina(w_n123_0[1]),.dinb(w_G97_2[2]),.dout(n980),.clk(gclk));
	jor g0908(.dina(w_dff_B_tybHPE6C0_0),.dinb(w_n672_0[1]),.dout(n981),.clk(gclk));
	jor g0909(.dina(n981),.dinb(w_dff_B_C05oqTQr5_1),.dout(n982),.clk(gclk));
	jand g0910(.dina(n982),.dinb(w_n604_0[2]),.dout(n983),.clk(gclk));
	jand g0911(.dina(w_dff_B_bd4qKzwn7_0),.dinb(n978),.dout(n984),.clk(gclk));
	jand g0912(.dina(w_dff_B_5FHqcI0s9_0),.dinb(n946),.dout(n985),.clk(gclk));
	jnot g0913(.din(n985),.dout(n986),.clk(gclk));
	jand g0914(.dina(w_dff_B_Hlt852rt5_0),.dinb(n944),.dout(n987),.clk(gclk));
	jand g0915(.dina(n987),.dinb(n943),.dout(n988),.clk(gclk));
	jnot g0916(.din(w_n988_0[2]),.dout(w_dff_A_ij4JhiJs2_1),.clk(gclk));
	jnot g0917(.din(w_n758_0[2]),.dout(n990),.clk(gclk));
	jand g0918(.dina(w_n696_0[1]),.dinb(w_n588_0[1]),.dout(n991),.clk(gclk));
	jand g0919(.dina(w_n991_0[1]),.dinb(w_n764_0[2]),.dout(n992),.clk(gclk));
	jxor g0920(.dina(w_n992_0[1]),.dinb(w_n990_0[1]),.dout(n993),.clk(gclk));
	jxor g0921(.dina(n993),.dinb(w_n769_0[0]),.dout(n994),.clk(gclk));
	jand g0922(.dina(w_n589_0[1]),.dinb(w_n519_0[1]),.dout(n995),.clk(gclk));
	jor g0923(.dina(n995),.dinb(w_n548_0[0]),.dout(n996),.clk(gclk));
	jand g0924(.dina(w_n554_1[0]),.dinb(w_n404_0[0]),.dout(n997),.clk(gclk));
	jor g0925(.dina(w_dff_B_wPggN8AG0_0),.dinb(w_n759_0[0]),.dout(n998),.clk(gclk));
	jnot g0926(.din(w_n764_0[1]),.dout(n999),.clk(gclk));
	jxor g0927(.dina(w_n991_0[0]),.dinb(w_n999_0[1]),.dout(n1000),.clk(gclk));
	jxor g0928(.dina(n1000),.dinb(n998),.dout(n1001),.clk(gclk));
	jor g0929(.dina(w_n1001_0[2]),.dinb(w_n996_0[2]),.dout(n1002),.clk(gclk));
	jor g0930(.dina(w_n1002_0[2]),.dinb(w_n994_0[2]),.dout(n1003),.clk(gclk));
	jnot g0931(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jand g0932(.dina(w_n1002_0[1]),.dinb(w_n994_0[1]),.dout(n1005),.clk(gclk));
	jor g0933(.dina(n1005),.dinb(w_n592_1[0]),.dout(n1006),.clk(gclk));
	jor g0934(.dina(n1006),.dinb(n1004),.dout(n1007),.clk(gclk));
	jor g0935(.dina(w_n994_0[0]),.dinb(w_n603_1[1]),.dout(n1008),.clk(gclk));
	jand g0936(.dina(w_n990_0[0]),.dinb(w_n425_1[0]),.dout(n1009),.clk(gclk));
	jnot g0937(.din(n1009),.dout(n1010),.clk(gclk));
	jand g0938(.dina(w_n631_4[0]),.dinb(w_G125_0[1]),.dout(n1011),.clk(gclk));
	jand g0939(.dina(w_n623_2[1]),.dinb(w_G159_1[2]),.dout(n1012),.clk(gclk));
	jand g0940(.dina(w_n642_4[0]),.dinb(w_G137_1[0]),.dout(n1013),.clk(gclk));
	jor g0941(.dina(w_dff_B_ECYdSkgf0_0),.dinb(n1012),.dout(n1014),.clk(gclk));
	jor g0942(.dina(n1014),.dinb(w_dff_B_H4wbGmLC0_1),.dout(n1015),.clk(gclk));
	jand g0943(.dina(w_n617_3[0]),.dinb(w_G150_1[2]),.dout(n1016),.clk(gclk));
	jor g0944(.dina(n1016),.dinb(w_G33_4[1]),.dout(n1017),.clk(gclk));
	jand g0945(.dina(w_n636_4[0]),.dinb(w_G143_1[1]),.dout(n1018),.clk(gclk));
	jand g0946(.dina(w_n627_4[0]),.dinb(w_G132_1[0]),.dout(n1019),.clk(gclk));
	jor g0947(.dina(n1019),.dinb(n1018),.dout(n1020),.clk(gclk));
	jand g0948(.dina(w_n640_4[0]),.dinb(w_G128_0[2]),.dout(n1021),.clk(gclk));
	jand g0949(.dina(w_n634_2[0]),.dinb(w_G50_2[0]),.dout(n1022),.clk(gclk));
	jor g0950(.dina(n1022),.dinb(w_dff_B_pMOYEzSd0_1),.dout(n1023),.clk(gclk));
	jor g0951(.dina(n1023),.dinb(w_dff_B_t4O3bn2m0_1),.dout(n1024),.clk(gclk));
	jor g0952(.dina(n1024),.dinb(w_dff_B_R4fIqzS48_1),.dout(n1025),.clk(gclk));
	jor g0953(.dina(n1025),.dinb(w_dff_B_DMifZ2951_1),.dout(n1026),.clk(gclk));
	jand g0954(.dina(w_n631_3[2]),.dinb(w_G294_1[1]),.dout(n1027),.clk(gclk));
	jand g0955(.dina(w_n642_3[2]),.dinb(w_G107_2[1]),.dout(n1028),.clk(gclk));
	jor g0956(.dina(w_dff_B_1Bg5NWFk1_0),.dinb(w_n962_0[0]),.dout(n1029),.clk(gclk));
	jor g0957(.dina(n1029),.dinb(w_dff_B_iqyfaPSa7_1),.dout(n1030),.clk(gclk));
	jand g0958(.dina(w_n640_3[2]),.dinb(w_G283_1[2]),.dout(n1031),.clk(gclk));
	jor g0959(.dina(n1031),.dinb(w_n148_3[2]),.dout(n1032),.clk(gclk));
	jand g0960(.dina(w_n636_3[2]),.dinb(w_G97_2[1]),.dout(n1033),.clk(gclk));
	jand g0961(.dina(w_n627_3[2]),.dinb(w_G116_2[0]),.dout(n1034),.clk(gclk));
	jor g0962(.dina(n1034),.dinb(n1033),.dout(n1035),.clk(gclk));
	jor g0963(.dina(w_n717_0[0]),.dinb(w_n654_0[0]),.dout(n1036),.clk(gclk));
	jor g0964(.dina(n1036),.dinb(w_dff_B_qWSCPjmn4_1),.dout(n1037),.clk(gclk));
	jor g0965(.dina(n1037),.dinb(w_dff_B_IdX0IT347_1),.dout(n1038),.clk(gclk));
	jor g0966(.dina(n1038),.dinb(w_dff_B_CflVqS060_1),.dout(n1039),.clk(gclk));
	jand g0967(.dina(n1039),.dinb(n1026),.dout(n1040),.clk(gclk));
	jor g0968(.dina(n1040),.dinb(w_n612_2[0]),.dout(n1041),.clk(gclk));
	jand g0969(.dina(w_n743_1[0]),.dinb(w_n74_0[1]),.dout(n1042),.clk(gclk));
	jor g0970(.dina(w_dff_B_1ETCG16F7_0),.dinb(w_n605_1[0]),.dout(n1043),.clk(gclk));
	jnot g0971(.din(n1043),.dout(n1044),.clk(gclk));
	jand g0972(.dina(w_dff_B_QS0ZtmA05_0),.dinb(n1041),.dout(n1045),.clk(gclk));
	jand g0973(.dina(w_dff_B_rqk3hDLC2_0),.dinb(n1010),.dout(n1046),.clk(gclk));
	jnot g0974(.din(n1046),.dout(n1047),.clk(gclk));
	jand g0975(.dina(w_dff_B_NZiGFut64_0),.dinb(n1008),.dout(n1048),.clk(gclk));
	jand g0976(.dina(w_dff_B_WRO4cqmB1_0),.dinb(n1007),.dout(n1049),.clk(gclk));
	jnot g0977(.din(w_n1049_0[2]),.dout(w_dff_A_9yDN0YMg2_1),.clk(gclk));
	jand g0978(.dina(w_n992_0[0]),.dinb(w_n758_0[1]),.dout(n1051),.clk(gclk));
	jand g0979(.dina(w_n552_0[1]),.dinb(w_n479_0[0]),.dout(n1052),.clk(gclk));
	jnot g0980(.din(w_n1052_0[1]),.dout(n1053),.clk(gclk));
	jand g0981(.dina(n1053),.dinb(w_n484_0[0]),.dout(n1054),.clk(gclk));
	jand g0982(.dina(w_n1052_0[0]),.dinb(w_n541_0[0]),.dout(n1055),.clk(gclk));
	jor g0983(.dina(n1055),.dinb(n1054),.dout(n1056),.clk(gclk));
	jnot g0984(.din(n1056),.dout(n1057),.clk(gclk));
	jxor g0985(.dina(w_n1057_0[1]),.dinb(w_n771_0[0]),.dout(n1058),.clk(gclk));
	jxor g0986(.dina(n1058),.dinb(w_dff_B_UR8JTR1B3_1),.dout(n1059),.clk(gclk));
	jor g0987(.dina(w_n1059_0[1]),.dinb(w_n603_1[0]),.dout(n1060),.clk(gclk));
	jnot g0988(.din(w_n996_0[1]),.dout(n1061),.clk(gclk));
	jand g0989(.dina(w_n1003_0[0]),.dinb(w_dff_B_MNVBHVb13_1),.dout(n1062),.clk(gclk));
	jor g0990(.dina(n1062),.dinb(w_n592_0[2]),.dout(n1063),.clk(gclk));
	jor g0991(.dina(n1063),.dinb(w_n1059_0[0]),.dout(n1064),.clk(gclk));
	jand g0992(.dina(w_n1057_0[0]),.dinb(w_n425_0[2]),.dout(n1065),.clk(gclk));
	jnot g0993(.din(w_n612_1[2]),.dout(n1066),.clk(gclk));
	jand g0994(.dina(w_n642_3[1]),.dinb(w_G132_0[2]),.dout(n1067),.clk(gclk));
	jand g0995(.dina(w_n627_3[1]),.dinb(w_G128_0[1]),.dout(n1068),.clk(gclk));
	jand g0996(.dina(w_n636_3[1]),.dinb(w_G137_0[2]),.dout(n1069),.clk(gclk));
	jor g0997(.dina(n1069),.dinb(n1068),.dout(n1070),.clk(gclk));
	jor g0998(.dina(n1070),.dinb(w_dff_B_ZfoTuBf89_1),.dout(n1071),.clk(gclk));
	jnot g0999(.din(n1071),.dout(n1072),.clk(gclk));
	jand g1000(.dina(w_n623_2[0]),.dinb(w_G150_1[1]),.dout(n1073),.clk(gclk));
	jnot g1001(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1002(.dina(w_n149_1[0]),.dinb(w_n148_3[1]),.dout(n1075),.clk(gclk));
	jand g1003(.dina(w_dff_B_MtutydP07_0),.dinb(n1074),.dout(n1076),.clk(gclk));
	jand g1004(.dina(w_n640_3[1]),.dinb(w_G125_0[0]),.dout(n1077),.clk(gclk));
	jand g1005(.dina(w_n617_2[2]),.dinb(w_G143_1[0]),.dout(n1078),.clk(gclk));
	jor g1006(.dina(n1078),.dinb(w_dff_B_sBac9MlJ7_1),.dout(n1079),.clk(gclk));
	jand g1007(.dina(w_n631_3[1]),.dinb(w_dff_B_wxIQ6v6t5_1),.dout(n1080),.clk(gclk));
	jand g1008(.dina(w_n634_1[2]),.dinb(w_G159_1[1]),.dout(n1081),.clk(gclk));
	jor g1009(.dina(n1081),.dinb(n1080),.dout(n1082),.clk(gclk));
	jor g1010(.dina(n1082),.dinb(n1079),.dout(n1083),.clk(gclk));
	jnot g1011(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1012(.dina(n1084),.dinb(w_dff_B_lDAau8753_1),.dout(n1085),.clk(gclk));
	jand g1013(.dina(n1085),.dinb(w_dff_B_yVxRmE8s9_1),.dout(n1086),.clk(gclk));
	jand g1014(.dina(w_n627_3[0]),.dinb(w_G107_2[0]),.dout(n1087),.clk(gclk));
	jand g1015(.dina(w_n634_1[1]),.dinb(w_G58_1[2]),.dout(n1088),.clk(gclk));
	jand g1016(.dina(w_n636_3[0]),.dinb(w_G87_1[0]),.dout(n1089),.clk(gclk));
	jor g1017(.dina(w_dff_B_SqTZABBO3_0),.dinb(w_n1088_0[1]),.dout(n1090),.clk(gclk));
	jor g1018(.dina(n1090),.dinb(w_dff_B_N3LKBBhK5_1),.dout(n1091),.clk(gclk));
	jnot g1019(.din(n1091),.dout(n1092),.clk(gclk));
	jand g1020(.dina(w_n642_3[0]),.dinb(w_G97_2[0]),.dout(n1093),.clk(gclk));
	jnot g1021(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1022(.dina(w_n149_0[2]),.dinb(w_G33_4[0]),.dout(n1095),.clk(gclk));
	jand g1023(.dina(w_dff_B_GlwAPsGr3_0),.dinb(n1094),.dout(n1096),.clk(gclk));
	jand g1024(.dina(w_n631_3[0]),.dinb(w_G283_1[1]),.dout(n1097),.clk(gclk));
	jor g1025(.dina(n1097),.dinb(w_n823_0[0]),.dout(n1098),.clk(gclk));
	jand g1026(.dina(w_n640_3[0]),.dinb(w_G116_1[2]),.dout(n1099),.clk(gclk));
	jor g1027(.dina(w_dff_B_eukirPuF1_0),.dinb(w_n909_0[0]),.dout(n1100),.clk(gclk));
	jor g1028(.dina(n1100),.dinb(n1098),.dout(n1101),.clk(gclk));
	jnot g1029(.din(n1101),.dout(n1102),.clk(gclk));
	jand g1030(.dina(n1102),.dinb(w_dff_B_4u4Xii5w3_1),.dout(n1103),.clk(gclk));
	jand g1031(.dina(n1103),.dinb(w_dff_B_tpz87DSL5_1),.dout(n1104),.clk(gclk));
	jand g1032(.dina(w_n73_1[0]),.dinb(w_G41_0[1]),.dout(n1105),.clk(gclk));
	jor g1033(.dina(w_dff_B_9yTnoITB3_0),.dinb(n1104),.dout(n1106),.clk(gclk));
	jor g1034(.dina(n1106),.dinb(w_dff_B_jkOunhVU9_1),.dout(n1107),.clk(gclk));
	jand g1035(.dina(n1107),.dinb(w_dff_B_cvIotsGl6_1),.dout(n1108),.clk(gclk));
	jand g1036(.dina(w_n743_0[2]),.dinb(w_n73_0[2]),.dout(n1109),.clk(gclk));
	jor g1037(.dina(w_dff_B_fapM1V6I5_0),.dinb(w_n605_0[2]),.dout(n1110),.clk(gclk));
	jor g1038(.dina(w_dff_B_zWQ86AaD6_0),.dinb(n1108),.dout(n1111),.clk(gclk));
	jor g1039(.dina(w_dff_B_w0GE4BjP7_0),.dinb(n1065),.dout(n1112),.clk(gclk));
	jand g1040(.dina(w_dff_B_KqbWPMAA7_0),.dinb(n1064),.dout(n1113),.clk(gclk));
	jand g1041(.dina(n1113),.dinb(w_dff_B_HqIxwYqi2_1),.dout(n1114),.clk(gclk));
	jnot g1042(.din(w_n1114_0[2]),.dout(w_dff_A_wSPhLArv2_1),.clk(gclk));
	jand g1043(.dina(w_n1001_0[1]),.dinb(w_n996_0[0]),.dout(n1116),.clk(gclk));
	jnot g1044(.din(n1116),.dout(n1117),.clk(gclk));
	jand g1045(.dina(w_n1002_0[0]),.dinb(w_n591_0[1]),.dout(n1118),.clk(gclk));
	jand g1046(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jnot g1047(.din(n1119),.dout(n1120),.clk(gclk));
	jor g1048(.dina(w_n1001_0[0]),.dinb(w_n603_0[2]),.dout(n1121),.clk(gclk));
	jand g1049(.dina(w_n999_0[0]),.dinb(w_n425_0[1]),.dout(n1122),.clk(gclk));
	jnot g1050(.din(n1122),.dout(n1123),.clk(gclk));
	jand g1051(.dina(w_n623_1[2]),.dinb(w_G50_1[2]),.dout(n1124),.clk(gclk));
	jand g1052(.dina(w_n617_2[1]),.dinb(w_G159_1[0]),.dout(n1125),.clk(gclk));
	jand g1053(.dina(w_n642_2[2]),.dinb(w_G143_0[2]),.dout(n1126),.clk(gclk));
	jor g1054(.dina(w_dff_B_LpNfrY359_0),.dinb(n1125),.dout(n1127),.clk(gclk));
	jor g1055(.dina(n1127),.dinb(w_dff_B_GdT3MNyE9_1),.dout(n1128),.clk(gclk));
	jand g1056(.dina(w_n631_2[2]),.dinb(w_G128_0[0]),.dout(n1129),.clk(gclk));
	jor g1057(.dina(n1129),.dinb(w_G33_3[2]),.dout(n1130),.clk(gclk));
	jand g1058(.dina(w_n636_2[2]),.dinb(w_G150_1[0]),.dout(n1131),.clk(gclk));
	jand g1059(.dina(w_n627_2[2]),.dinb(w_G137_0[1]),.dout(n1132),.clk(gclk));
	jor g1060(.dina(n1132),.dinb(n1131),.dout(n1133),.clk(gclk));
	jand g1061(.dina(w_n640_2[2]),.dinb(w_G132_0[1]),.dout(n1134),.clk(gclk));
	jor g1062(.dina(w_dff_B_07FqMLME8_0),.dinb(w_n1088_0[0]),.dout(n1135),.clk(gclk));
	jor g1063(.dina(n1135),.dinb(w_dff_B_ui9JvqB01_1),.dout(n1136),.clk(gclk));
	jor g1064(.dina(n1136),.dinb(w_dff_B_YnLdvlym2_1),.dout(n1137),.clk(gclk));
	jor g1065(.dina(n1137),.dinb(w_dff_B_nx93J3LY3_1),.dout(n1138),.clk(gclk));
	jand g1066(.dina(w_n617_2[0]),.dinb(w_G97_1[2]),.dout(n1139),.clk(gclk));
	jand g1067(.dina(w_n640_2[1]),.dinb(w_G294_1[0]),.dout(n1140),.clk(gclk));
	jand g1068(.dina(w_n642_2[1]),.dinb(w_G116_1[1]),.dout(n1141),.clk(gclk));
	jor g1069(.dina(n1141),.dinb(n1140),.dout(n1142),.clk(gclk));
	jor g1070(.dina(n1142),.dinb(n1139),.dout(n1143),.clk(gclk));
	jand g1071(.dina(w_n631_2[1]),.dinb(w_G303_0[2]),.dout(n1144),.clk(gclk));
	jor g1072(.dina(n1144),.dinb(w_n148_3[0]),.dout(n1145),.clk(gclk));
	jand g1073(.dina(w_n636_2[1]),.dinb(w_G107_1[2]),.dout(n1146),.clk(gclk));
	jand g1074(.dina(w_n627_2[1]),.dinb(w_G283_1[0]),.dout(n1147),.clk(gclk));
	jor g1075(.dina(n1147),.dinb(n1146),.dout(n1148),.clk(gclk));
	jor g1076(.dina(w_n899_0[0]),.dinb(w_n825_0[0]),.dout(n1149),.clk(gclk));
	jor g1077(.dina(n1149),.dinb(w_dff_B_GuNW2e8p9_1),.dout(n1150),.clk(gclk));
	jor g1078(.dina(n1150),.dinb(w_dff_B_5yDNasKG3_1),.dout(n1151),.clk(gclk));
	jor g1079(.dina(n1151),.dinb(w_dff_B_ORN9O6023_1),.dout(n1152),.clk(gclk));
	jand g1080(.dina(n1152),.dinb(n1138),.dout(n1153),.clk(gclk));
	jor g1081(.dina(n1153),.dinb(w_n612_1[1]),.dout(n1154),.clk(gclk));
	jand g1082(.dina(w_n743_0[1]),.dinb(w_n75_0[1]),.dout(n1155),.clk(gclk));
	jor g1083(.dina(w_dff_B_jzkxmxX52_0),.dinb(w_n605_0[1]),.dout(n1156),.clk(gclk));
	jnot g1084(.din(n1156),.dout(n1157),.clk(gclk));
	jand g1085(.dina(w_dff_B_Lq59G3kr3_0),.dinb(n1154),.dout(n1158),.clk(gclk));
	jand g1086(.dina(w_dff_B_XgRgISjX1_0),.dinb(n1123),.dout(n1159),.clk(gclk));
	jnot g1087(.din(n1159),.dout(n1160),.clk(gclk));
	jand g1088(.dina(n1160),.dinb(n1121),.dout(n1161),.clk(gclk));
	jand g1089(.dina(w_dff_B_8uFYQU0E4_0),.dinb(n1120),.dout(n1162),.clk(gclk));
	jnot g1090(.din(w_n1162_0[2]),.dout(w_dff_A_2VxUnDSH8_1),.clk(gclk));
	jand g1091(.dina(w_n1114_0[1]),.dinb(w_n1049_0[1]),.dout(n1164),.clk(gclk));
	jnot g1092(.din(w_G387_0[1]),.dout(n1165),.clk(gclk));
	jnot g1093(.din(w_G396_0[1]),.dout(n1166),.clk(gclk));
	jand g1094(.dina(w_n937_0[1]),.dinb(w_dff_B_pqHyahDE9_1),.dout(n1167),.clk(gclk));
	jand g1095(.dina(n1167),.dinb(w_n750_0[0]),.dout(n1168),.clk(gclk));
	jand g1096(.dina(n1168),.dinb(w_n988_0[1]),.dout(n1169),.clk(gclk));
	jand g1097(.dina(n1169),.dinb(w_n1162_0[1]),.dout(n1170),.clk(gclk));
	jand g1098(.dina(n1170),.dinb(n1165),.dout(n1171),.clk(gclk));
	jand g1099(.dina(n1171),.dinb(w_n1164_0[1]),.dout(n1172),.clk(gclk));
	jnot g1100(.din(w_n1172_0[1]),.dout(w_dff_A_9QSoc5cq7_1),.clk(gclk));
	jnot g1101(.din(w_G213_0[1]),.dout(n1174),.clk(gclk));
	jnot g1102(.din(w_G343_0[0]),.dout(n1175),.clk(gclk));
	jand g1103(.dina(w_n1164_0[0]),.dinb(w_n1175_0[1]),.dout(n1176),.clk(gclk));
	jor g1104(.dina(n1176),.dinb(w_dff_B_zk7gRSOB7_1),.dout(n1177),.clk(gclk));
	jor g1105(.dina(n1177),.dinb(w_n1172_0[0]),.dout(G409),.clk(gclk));
	jxor g1106(.dina(w_n1162_0[0]),.dinb(w_G384_0),.dout(n1179),.clk(gclk));
	jxor g1107(.dina(w_n937_0[0]),.dinb(w_G396_0[0]),.dout(n1180),.clk(gclk));
	jxor g1108(.dina(w_n988_0[0]),.dinb(w_G387_0[0]),.dout(n1181),.clk(gclk));
	jxor g1109(.dina(n1181),.dinb(w_dff_B_iBNBekbK7_1),.dout(n1182),.clk(gclk));
	jxor g1110(.dina(n1182),.dinb(w_dff_B_jlWztoAt0_1),.dout(n1183),.clk(gclk));
	jand g1111(.dina(w_n1175_0[0]),.dinb(w_G213_0[0]),.dout(n1184),.clk(gclk));
	jnot g1112(.din(w_n1184_0[1]),.dout(n1185),.clk(gclk));
	jor g1113(.dina(n1185),.dinb(w_dff_B_89NlKiQx0_1),.dout(n1186),.clk(gclk));
	jxor g1114(.dina(w_n1114_0[0]),.dinb(w_n1049_0[0]),.dout(n1187),.clk(gclk));
	jor g1115(.dina(w_n1187_0[1]),.dinb(w_n1184_0[0]),.dout(n1188),.clk(gclk));
	jand g1116(.dina(n1188),.dinb(w_dff_B_bvOcEYhx9_1),.dout(n1189),.clk(gclk));
	jxor g1117(.dina(n1189),.dinb(w_n1183_0[1]),.dout(G405),.clk(gclk));
	jxor g1118(.dina(w_n1187_0[0]),.dinb(w_n1183_0[0]),.dout(w_dff_A_5Bcl7rAn0_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_dff_A_pjgwWpzJ1_0),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_dff_A_jhqvHvKy5_0),.doutb(w_dff_A_RA3arEWY5_1),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G1_2(.douta(w_dff_A_X0OT3Diz9_0),.doutb(w_G1_2[1]),.doutc(w_dff_A_X0OpRtEZ5_2),.din(w_G1_0[1]));
	jspl jspl_w_G1_3(.douta(w_G1_3[0]),.doutb(w_G1_3[1]),.din(w_G1_0[2]));
	jspl3 jspl3_w_G13_0(.douta(w_G13_0[0]),.doutb(w_dff_A_pi8XySmV6_1),.doutc(w_dff_A_DlJf6hDJ7_2),.din(G13));
	jspl jspl_w_G13_1(.douta(w_G13_1[0]),.doutb(w_G13_1[1]),.din(w_G13_0[0]));
	jspl3 jspl3_w_G20_0(.douta(w_dff_A_PrKjblqV4_0),.doutb(w_G20_0[1]),.doutc(w_G20_0[2]),.din(G20));
	jspl3 jspl3_w_G20_1(.douta(w_G20_1[0]),.doutb(w_G20_1[1]),.doutc(w_dff_A_a8iaffyV9_2),.din(w_G20_0[0]));
	jspl3 jspl3_w_G20_2(.douta(w_G20_2[0]),.doutb(w_dff_A_3ugz4ekH2_1),.doutc(w_G20_2[2]),.din(w_G20_0[1]));
	jspl3 jspl3_w_G20_3(.douta(w_G20_3[0]),.doutb(w_dff_A_oNKs1aL00_1),.doutc(w_dff_A_oDxiCE6K5_2),.din(w_G20_0[2]));
	jspl3 jspl3_w_G20_4(.douta(w_dff_A_aA3KFQK93_0),.doutb(w_dff_A_fSTzQJGM8_1),.doutc(w_G20_4[2]),.din(w_G20_1[0]));
	jspl3 jspl3_w_G20_5(.douta(w_dff_A_W57appsB7_0),.doutb(w_dff_A_rvJlGxMM5_1),.doutc(w_G20_5[2]),.din(w_G20_1[1]));
	jspl3 jspl3_w_G20_6(.douta(w_dff_A_H1BMiCLW6_0),.doutb(w_G20_6[1]),.doutc(w_G20_6[2]),.din(w_G20_1[2]));
	jspl jspl_w_G20_7(.douta(w_G20_7[0]),.doutb(w_G20_7[1]),.din(w_G20_2[0]));
	jspl3 jspl3_w_G33_0(.douta(w_dff_A_6zatj6M01_0),.doutb(w_G33_0[1]),.doutc(w_G33_0[2]),.din(G33));
	jspl3 jspl3_w_G33_1(.douta(w_G33_1[0]),.doutb(w_dff_A_BgoFfZ3G5_1),.doutc(w_G33_1[2]),.din(w_G33_0[0]));
	jspl3 jspl3_w_G33_2(.douta(w_G33_2[0]),.doutb(w_G33_2[1]),.doutc(w_G33_2[2]),.din(w_G33_0[1]));
	jspl3 jspl3_w_G33_3(.douta(w_G33_3[0]),.doutb(w_G33_3[1]),.doutc(w_dff_A_GKmywLFy8_2),.din(w_G33_0[2]));
	jspl3 jspl3_w_G33_4(.douta(w_G33_4[0]),.doutb(w_dff_A_F7LThMu61_1),.doutc(w_dff_A_U84xEFrr8_2),.din(w_G33_1[0]));
	jspl3 jspl3_w_G33_5(.douta(w_dff_A_K9gIku7k7_0),.doutb(w_G33_5[1]),.doutc(w_dff_A_TeDTVq7P5_2),.din(w_G33_1[1]));
	jspl3 jspl3_w_G33_6(.douta(w_dff_A_c0tZk3tN5_0),.doutb(w_dff_A_Os20HUNC9_1),.doutc(w_G33_6[2]),.din(w_G33_1[2]));
	jspl3 jspl3_w_G33_7(.douta(w_G33_7[0]),.doutb(w_G33_7[1]),.doutc(w_G33_7[2]),.din(w_G33_2[0]));
	jspl3 jspl3_w_G33_8(.douta(w_dff_A_SYSv08G87_0),.doutb(w_G33_8[1]),.doutc(w_G33_8[2]),.din(w_G33_2[1]));
	jspl3 jspl3_w_G33_9(.douta(w_G33_9[0]),.doutb(w_G33_9[1]),.doutc(w_dff_A_zh0VzruW5_2),.din(w_G33_2[2]));
	jspl3 jspl3_w_G33_10(.douta(w_dff_A_g5BCQ1hB0_0),.doutb(w_dff_A_UJGM8GXu6_1),.doutc(w_G33_10[2]),.din(w_G33_3[0]));
	jspl3 jspl3_w_G33_11(.douta(w_G33_11[0]),.doutb(w_G33_11[1]),.doutc(w_G33_11[2]),.din(w_G33_3[1]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_dff_A_Wo6mhXIz9_1),.doutc(w_dff_A_EE6LrMLh2_2),.din(G41));
	jspl jspl_w_G41_1(.douta(w_G41_1[0]),.doutb(w_G41_1[1]),.din(w_G41_0[0]));
	jspl3 jspl3_w_G45_0(.douta(w_G45_0[0]),.doutb(w_dff_A_LKBQMA7Q4_1),.doutc(w_dff_A_zXJtZd5W5_2),.din(G45));
	jspl3 jspl3_w_G45_1(.douta(w_dff_A_6srOqm5Z0_0),.doutb(w_dff_A_js40K4Sf9_1),.doutc(w_G45_1[2]),.din(w_G45_0[0]));
	jspl3 jspl3_w_G50_0(.douta(w_G50_0[0]),.doutb(w_dff_A_YtGq8GRF4_1),.doutc(w_G50_0[2]),.din(G50));
	jspl3 jspl3_w_G50_1(.douta(w_dff_A_B5q9nHKd8_0),.doutb(w_G50_1[1]),.doutc(w_dff_A_T6Lcc6IH2_2),.din(w_G50_0[0]));
	jspl3 jspl3_w_G50_2(.douta(w_dff_A_dueqaJgq7_0),.doutb(w_G50_2[1]),.doutc(w_G50_2[2]),.din(w_G50_0[1]));
	jspl3 jspl3_w_G50_3(.douta(w_dff_A_q4g8PyAu0_0),.doutb(w_G50_3[1]),.doutc(w_dff_A_0z4pOVe93_2),.din(w_G50_0[2]));
	jspl3 jspl3_w_G50_4(.douta(w_dff_A_ErXiBYYZ2_0),.doutb(w_dff_A_cR9FzrOM6_1),.doutc(w_G50_4[2]),.din(w_G50_1[0]));
	jspl3 jspl3_w_G50_5(.douta(w_G50_5[0]),.doutb(w_dff_A_wySSWbT54_1),.doutc(w_G50_5[2]),.din(w_G50_1[1]));
	jspl3 jspl3_w_G58_0(.douta(w_G58_0[0]),.doutb(w_dff_A_O5xTzMGe8_1),.doutc(w_dff_A_5GiiMNAY6_2),.din(G58));
	jspl3 jspl3_w_G58_1(.douta(w_dff_A_iBXOt02u3_0),.doutb(w_G58_1[1]),.doutc(w_dff_A_m1kh582q3_2),.din(w_G58_0[0]));
	jspl3 jspl3_w_G58_2(.douta(w_dff_A_Cfx5oZ4z1_0),.doutb(w_G58_2[1]),.doutc(w_dff_A_ul9kiYTC7_2),.din(w_G58_0[1]));
	jspl3 jspl3_w_G58_3(.douta(w_dff_A_B9U87A7P4_0),.doutb(w_dff_A_8HWxLwAr6_1),.doutc(w_G58_3[2]),.din(w_G58_0[2]));
	jspl3 jspl3_w_G58_4(.douta(w_dff_A_2N6qgzwC1_0),.doutb(w_dff_A_12RyQrOQ0_1),.doutc(w_G58_4[2]),.din(w_G58_1[0]));
	jspl jspl_w_G58_5(.douta(w_G58_5[0]),.doutb(w_G58_5[1]),.din(w_G58_1[1]));
	jspl3 jspl3_w_G68_0(.douta(w_G68_0[0]),.doutb(w_G68_0[1]),.doutc(w_dff_A_iHywy3nW6_2),.din(G68));
	jspl3 jspl3_w_G68_1(.douta(w_dff_A_gPbxcvWN4_0),.doutb(w_G68_1[1]),.doutc(w_dff_A_RNnn8wkf2_2),.din(w_G68_0[0]));
	jspl3 jspl3_w_G68_2(.douta(w_G68_2[0]),.doutb(w_dff_A_gRyxMBcX9_1),.doutc(w_dff_A_64ftG2JB1_2),.din(w_G68_0[1]));
	jspl3 jspl3_w_G68_3(.douta(w_G68_3[0]),.doutb(w_dff_A_A7uLTU6D5_1),.doutc(w_dff_A_QAexC1sc5_2),.din(w_G68_0[2]));
	jspl3 jspl3_w_G68_4(.douta(w_dff_A_GckQdKlQ9_0),.doutb(w_dff_A_bpt5RxmD3_1),.doutc(w_G68_4[2]),.din(w_G68_1[0]));
	jspl jspl_w_G68_5(.douta(w_G68_5[0]),.doutb(w_G68_5[1]),.din(w_G68_1[1]));
	jspl3 jspl3_w_G77_0(.douta(w_G77_0[0]),.doutb(w_G77_0[1]),.doutc(w_G77_0[2]),.din(G77));
	jspl3 jspl3_w_G77_1(.douta(w_dff_A_dL83xHsC3_0),.doutb(w_G77_1[1]),.doutc(w_dff_A_hxoan87X8_2),.din(w_G77_0[0]));
	jspl3 jspl3_w_G77_2(.douta(w_G77_2[0]),.doutb(w_dff_A_E9E5rxLQ7_1),.doutc(w_dff_A_UPue7mKt7_2),.din(w_G77_0[1]));
	jspl3 jspl3_w_G77_3(.douta(w_G77_3[0]),.doutb(w_dff_A_f4ZUCAnr5_1),.doutc(w_G77_3[2]),.din(w_G77_0[2]));
	jspl3 jspl3_w_G77_4(.douta(w_dff_A_zKYKHmZ62_0),.doutb(w_G77_4[1]),.doutc(w_G77_4[2]),.din(w_G77_1[0]));
	jspl jspl_w_G77_5(.douta(w_G77_5[0]),.doutb(w_G77_5[1]),.din(w_G77_1[1]));
	jspl3 jspl3_w_G87_0(.douta(w_dff_A_wlDyDHq85_0),.doutb(w_G87_0[1]),.doutc(w_G87_0[2]),.din(G87));
	jspl3 jspl3_w_G87_1(.douta(w_G87_1[0]),.doutb(w_dff_A_byatC4aG6_1),.doutc(w_dff_A_hHFRDDwG8_2),.din(w_G87_0[0]));
	jspl3 jspl3_w_G87_2(.douta(w_dff_A_AzYgYmxN5_0),.doutb(w_dff_A_3XLrzspX8_1),.doutc(w_G87_2[2]),.din(w_G87_0[1]));
	jspl3 jspl3_w_G87_3(.douta(w_dff_A_kurh59Sd5_0),.doutb(w_G87_3[1]),.doutc(w_dff_A_8CcwNKW05_2),.din(w_G87_0[2]));
	jspl3 jspl3_w_G97_0(.douta(w_G97_0[0]),.doutb(w_dff_A_LbIR4ecf3_1),.doutc(w_dff_A_UERcl1tV7_2),.din(G97));
	jspl3 jspl3_w_G97_1(.douta(w_G97_1[0]),.doutb(w_G97_1[1]),.doutc(w_dff_A_UPHWAMW62_2),.din(w_G97_0[0]));
	jspl3 jspl3_w_G97_2(.douta(w_G97_2[0]),.doutb(w_G97_2[1]),.doutc(w_dff_A_7QBH7DgZ4_2),.din(w_G97_0[1]));
	jspl3 jspl3_w_G97_3(.douta(w_dff_A_YTISlkpo1_0),.doutb(w_dff_A_RpaMBR3p5_1),.doutc(w_G97_3[2]),.din(w_G97_0[2]));
	jspl3 jspl3_w_G97_4(.douta(w_dff_A_VSsmvDUq1_0),.doutb(w_G97_4[1]),.doutc(w_G97_4[2]),.din(w_G97_1[0]));
	jspl jspl_w_G97_5(.douta(w_dff_A_KAbfLiU74_0),.doutb(w_G97_5[1]),.din(w_G97_1[1]));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_dff_A_zpj0968i2_1),.doutc(w_dff_A_41vnu8CB0_2),.din(G107));
	jspl3 jspl3_w_G107_1(.douta(w_G107_1[0]),.doutb(w_G107_1[1]),.doutc(w_dff_A_mELiXizb9_2),.din(w_G107_0[0]));
	jspl3 jspl3_w_G107_2(.douta(w_G107_2[0]),.doutb(w_G107_2[1]),.doutc(w_dff_A_CPktjDSG5_2),.din(w_G107_0[1]));
	jspl3 jspl3_w_G107_3(.douta(w_dff_A_rDKXslHr0_0),.doutb(w_dff_A_gTv3yu3c8_1),.doutc(w_G107_3[2]),.din(w_G107_0[2]));
	jspl3 jspl3_w_G107_4(.douta(w_dff_A_diV3Ue6L8_0),.doutb(w_G107_4[1]),.doutc(w_G107_4[2]),.din(w_G107_1[0]));
	jspl jspl_w_G107_5(.douta(w_G107_5[0]),.doutb(w_G107_5[1]),.din(w_G107_1[1]));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_dff_A_xBne4DBd4_1),.doutc(w_dff_A_ck8EZlDh9_2),.din(G116));
	jspl3 jspl3_w_G116_1(.douta(w_G116_1[0]),.doutb(w_dff_A_NaGJkzdY8_1),.doutc(w_dff_A_kEIBVVPy7_2),.din(w_G116_0[0]));
	jspl3 jspl3_w_G116_2(.douta(w_G116_2[0]),.doutb(w_dff_A_P2HetoOa5_1),.doutc(w_dff_A_oerN6jKl5_2),.din(w_G116_0[1]));
	jspl3 jspl3_w_G116_3(.douta(w_dff_A_a7FNnu3y0_0),.doutb(w_G116_3[1]),.doutc(w_dff_A_xytoGJ765_2),.din(w_G116_0[2]));
	jspl3 jspl3_w_G116_4(.douta(w_G116_4[0]),.doutb(w_G116_4[1]),.doutc(w_G116_4[2]),.din(w_G116_1[0]));
	jspl jspl_w_G125_0(.douta(w_G125_0[0]),.doutb(w_dff_A_xryQdEie7_1),.din(w_dff_B_GGlOXZyL8_2));
	jspl3 jspl3_w_G128_0(.douta(w_dff_A_3k1m8a2A3_0),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(w_dff_B_Nv8zABFN6_3));
	jspl3 jspl3_w_G132_0(.douta(w_G132_0[0]),.doutb(w_G132_0[1]),.doutc(w_G132_0[2]),.din(w_dff_B_ZMOIlzt87_3));
	jspl jspl_w_G132_1(.douta(w_G132_1[0]),.doutb(w_dff_A_UqmQbHpi3_1),.din(w_G132_0[0]));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(w_dff_B_ob9irtai4_3));
	jspl3 jspl3_w_G137_1(.douta(w_G137_1[0]),.doutb(w_dff_A_fg08Ldde0_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(w_dff_B_OJom1FYt1_3));
	jspl3 jspl3_w_G143_1(.douta(w_dff_A_PugzPvyA2_0),.doutb(w_G143_1[1]),.doutc(w_dff_A_sFVymup87_2),.din(w_G143_0[0]));
	jspl jspl_w_G143_2(.douta(w_G143_2[0]),.doutb(w_G143_2[1]),.din(w_G143_0[1]));
	jspl3 jspl3_w_G150_0(.douta(w_dff_A_XapG0G1E1_0),.doutb(w_dff_A_3IWXGl4Q0_1),.doutc(w_G150_0[2]),.din(G150));
	jspl3 jspl3_w_G150_1(.douta(w_G150_1[0]),.doutb(w_dff_A_dNdWUtir8_1),.doutc(w_dff_A_HGXab7lh5_2),.din(w_G150_0[0]));
	jspl3 jspl3_w_G150_2(.douta(w_G150_2[0]),.doutb(w_dff_A_z0DziQVH6_1),.doutc(w_G150_2[2]),.din(w_G150_0[1]));
	jspl jspl_w_G150_3(.douta(w_dff_A_6kKoFWxY3_0),.doutb(w_G150_3[1]),.din(w_G150_0[2]));
	jspl3 jspl3_w_G159_0(.douta(w_dff_A_NYxeNxQl8_0),.doutb(w_dff_A_cIHiKiZJ6_1),.doutc(w_G159_0[2]),.din(w_dff_B_FaIakyj15_3));
	jspl3 jspl3_w_G159_1(.douta(w_G159_1[0]),.doutb(w_G159_1[1]),.doutc(w_G159_1[2]),.din(w_G159_0[0]));
	jspl3 jspl3_w_G159_2(.douta(w_G159_2[0]),.doutb(w_G159_2[1]),.doutc(w_G159_2[2]),.din(w_G159_0[1]));
	jspl3 jspl3_w_G159_3(.douta(w_dff_A_1jvSdNCV3_0),.doutb(w_dff_A_a7wtfoCu3_1),.doutc(w_G159_3[2]),.din(w_G159_0[2]));
	jspl3 jspl3_w_G169_0(.douta(w_G169_0[0]),.doutb(w_dff_A_5ltwZ2ye2_1),.doutc(w_dff_A_vkYHzYam5_2),.din(G169));
	jspl jspl_w_G169_1(.douta(w_dff_A_5SRtP6CE7_0),.doutb(w_G169_1[1]),.din(w_G169_0[0]));
	jspl3 jspl3_w_G179_0(.douta(w_dff_A_9SVGVaCc9_0),.doutb(w_G179_0[1]),.doutc(w_G179_0[2]),.din(G179));
	jspl3 jspl3_w_G179_1(.douta(w_G179_1[0]),.doutb(w_G179_1[1]),.doutc(w_G179_1[2]),.din(w_G179_0[0]));
	jspl3 jspl3_w_G179_2(.douta(w_dff_A_0Cd7dMhP4_0),.doutb(w_dff_A_hueIkzjX5_1),.doutc(w_G179_2[2]),.din(w_G179_0[1]));
	jspl3 jspl3_w_G190_0(.douta(w_dff_A_gp0OvPEx3_0),.doutb(w_dff_A_8WEsy4756_1),.doutc(w_G190_0[2]),.din(G190));
	jspl3 jspl3_w_G190_1(.douta(w_dff_A_lU4zRC4C0_0),.doutb(w_G190_1[1]),.doutc(w_G190_1[2]),.din(w_G190_0[0]));
	jspl3 jspl3_w_G190_2(.douta(w_G190_2[0]),.doutb(w_dff_A_bXRGpFUT9_1),.doutc(w_dff_A_ZwW0hqYD3_2),.din(w_G190_0[1]));
	jspl3 jspl3_w_G190_3(.douta(w_G190_3[0]),.doutb(w_dff_A_qZwwkgyD6_1),.doutc(w_dff_A_LDnZStKM2_2),.din(w_G190_0[2]));
	jspl jspl_w_G190_4(.douta(w_dff_A_h3hOAETZ3_0),.doutb(w_G190_4[1]),.din(w_G190_1[0]));
	jspl3 jspl3_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.doutc(w_dff_A_tSw5gpj66_2),.din(G200));
	jspl3 jspl3_w_G200_1(.douta(w_dff_A_04AmFTHf6_0),.doutb(w_dff_A_dvjVEWxA4_1),.doutc(w_G200_1[2]),.din(w_G200_0[0]));
	jspl3 jspl3_w_G200_2(.douta(w_G200_2[0]),.doutb(w_dff_A_ockTjTGj2_1),.doutc(w_dff_A_cCghVtay5_2),.din(w_G200_0[1]));
	jspl3 jspl3_w_G200_3(.douta(w_G200_3[0]),.doutb(w_G200_3[1]),.doutc(w_G200_3[2]),.din(w_G200_0[2]));
	jspl3 jspl3_w_G200_4(.douta(w_G200_4[0]),.doutb(w_G200_4[1]),.doutc(w_G200_4[2]),.din(w_G200_1[0]));
	jspl3 jspl3_w_G213_0(.douta(w_dff_A_7xrzCvZ98_0),.doutb(w_G213_0[1]),.doutc(w_dff_A_WHdKEeti2_2),.din(G213));
	jspl jspl_w_G223_0(.douta(w_G223_0[0]),.doutb(w_G223_0[1]),.din(w_dff_B_KYm3OC3V3_2));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_dff_A_VGVZ5Om46_1),.doutc(w_dff_A_Aw8GGBk42_2),.din(G226));
	jspl jspl_w_G226_1(.douta(w_dff_A_i2cl3Bp49_0),.doutb(w_G226_1[1]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G232_0(.douta(w_G232_0[0]),.doutb(w_dff_A_zfeHizBJ6_1),.doutc(w_dff_A_CC0y3FIr4_2),.din(G232));
	jspl3 jspl3_w_G232_1(.douta(w_dff_A_rPI04wTs3_0),.doutb(w_dff_A_4JHMJTxp3_1),.doutc(w_G232_1[2]),.din(w_G232_0[0]));
	jspl3 jspl3_w_G238_0(.douta(w_G238_0[0]),.doutb(w_dff_A_ygpYplsT6_1),.doutc(w_dff_A_71vYR1RX5_2),.din(G238));
	jspl3 jspl3_w_G238_1(.douta(w_dff_A_lN1JJFlD5_0),.doutb(w_G238_1[1]),.doutc(w_G238_1[2]),.din(w_G238_0[0]));
	jspl3 jspl3_w_G244_0(.douta(w_G244_0[0]),.doutb(w_dff_A_xklEYXbG0_1),.doutc(w_dff_A_ppap3l3i7_2),.din(G244));
	jspl3 jspl3_w_G244_1(.douta(w_dff_A_z9ZgqKo90_0),.doutb(w_G244_1[1]),.doutc(w_G244_1[2]),.din(w_G244_0[0]));
	jspl3 jspl3_w_G250_0(.douta(w_dff_A_g1sQxtI67_0),.doutb(w_dff_A_Pf8WR8ke6_1),.doutc(w_G250_0[2]),.din(G250));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_dff_A_ancPBdLJ4_1),.doutc(w_dff_A_7iP5EJLw6_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_gflqMBrW2_0),.doutb(w_dff_A_gmoFzwOH9_1),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G264_0(.douta(w_G264_0[0]),.doutb(w_dff_A_4UQrobXj6_1),.doutc(w_dff_A_wQqteubQ1_2),.din(G264));
	jspl jspl_w_G264_1(.douta(w_G264_1[0]),.doutb(w_G264_1[1]),.din(w_G264_0[0]));
	jspl3 jspl3_w_G270_0(.douta(w_dff_A_gzwjnW8H8_0),.doutb(w_G270_0[1]),.doutc(w_G270_0[2]),.din(G270));
	jspl3 jspl3_w_G274_0(.douta(w_dff_A_h6y2HzJO2_0),.doutb(w_G274_0[1]),.doutc(w_dff_A_IZ76Ei1m6_2),.din(G274));
	jspl3 jspl3_w_G283_0(.douta(w_dff_A_OrDQkYHF2_0),.doutb(w_dff_A_BEM9gBeJ0_1),.doutc(w_G283_0[2]),.din(G283));
	jspl3 jspl3_w_G283_1(.douta(w_G283_1[0]),.doutb(w_dff_A_VPKwfkVC7_1),.doutc(w_G283_1[2]),.din(w_G283_0[0]));
	jspl3 jspl3_w_G283_2(.douta(w_dff_A_ySobaZ7d0_0),.doutb(w_dff_A_4xonIQ2c6_1),.doutc(w_G283_2[2]),.din(w_G283_0[1]));
	jspl3 jspl3_w_G283_3(.douta(w_dff_A_vm3CoLng7_0),.doutb(w_dff_A_e8sfntoC4_1),.doutc(w_G283_3[2]),.din(w_G283_0[2]));
	jspl3 jspl3_w_G294_0(.douta(w_dff_A_pBjB8zcm8_0),.doutb(w_dff_A_5gty9tSV0_1),.doutc(w_G294_0[2]),.din(G294));
	jspl3 jspl3_w_G294_1(.douta(w_G294_1[0]),.doutb(w_dff_A_iBOwVAhb4_1),.doutc(w_G294_1[2]),.din(w_G294_0[0]));
	jspl3 jspl3_w_G294_2(.douta(w_dff_A_hARDuVkP8_0),.doutb(w_G294_2[1]),.doutc(w_G294_2[2]),.din(w_G294_0[1]));
	jspl jspl_w_G294_3(.douta(w_dff_A_h4Q5cbvG7_0),.doutb(w_G294_3[1]),.din(w_G294_0[2]));
	jspl3 jspl3_w_G303_0(.douta(w_dff_A_Q36Cbjon5_0),.doutb(w_G303_0[1]),.doutc(w_dff_A_phx9anFf7_2),.din(G303));
	jspl3 jspl3_w_G303_1(.douta(w_G303_1[0]),.doutb(w_G303_1[1]),.doutc(w_G303_1[2]),.din(w_G303_0[0]));
	jspl3 jspl3_w_G303_2(.douta(w_dff_A_FRSK5cPf6_0),.doutb(w_dff_A_HEpS09PU5_1),.doutc(w_G303_2[2]),.din(w_G303_0[1]));
	jspl3 jspl3_w_G311_0(.douta(w_G311_0[0]),.doutb(w_G311_0[1]),.doutc(w_G311_0[2]),.din(w_dff_B_VxTUBMna6_3));
	jspl3 jspl3_w_G311_1(.douta(w_G311_1[0]),.doutb(w_dff_A_PdTwVXbF9_1),.doutc(w_G311_1[2]),.din(w_G311_0[0]));
	jspl3 jspl3_w_G317_0(.douta(w_G317_0[0]),.doutb(w_G317_0[1]),.doutc(w_G317_0[2]),.din(w_dff_B_ZmiO3i2x6_3));
	jspl jspl_w_G317_1(.douta(w_dff_A_XwDnaQlt8_0),.doutb(w_G317_1[1]),.din(w_G317_0[0]));
	jspl3 jspl3_w_G322_0(.douta(w_dff_A_81pCt3ZJ1_0),.doutb(w_G322_0[1]),.doutc(w_G322_0[2]),.din(w_dff_B_rX8Nivot9_3));
	jspl jspl_w_G326_0(.douta(w_dff_A_v49lq3ym8_0),.doutb(w_G326_0[1]),.din(w_dff_B_iGSNmT5R3_2));
	jspl jspl_w_G330_0(.douta(w_dff_A_gGprMvpd8_0),.doutb(w_G330_0[1]),.din(G330));
	jspl jspl_w_G343_0(.douta(w_G343_0[0]),.doutb(w_dff_A_mvZgpjTa2_1),.din(G343));
	jspl3 jspl3_w_G1698_0(.douta(w_G1698_0[0]),.doutb(w_G1698_0[1]),.doutc(w_dff_A_Cc3xYaea6_2),.din(G1698));
	jspl jspl_w_G355_0(.douta(w_G355_0),.doutb(w_dff_A_D1cH4P2b3_1),.din(G355_fa_));
	jspl3 jspl3_w_G396_0(.douta(w_dff_A_wHFAAAM29_0),.doutb(w_G396_0[1]),.doutc(w_dff_A_OFRPwL4t5_2),.din(G396_fa_));
	jspl jspl_w_G384_0(.douta(w_dff_A_ogpRhe583_0),.doutb(w_dff_A_ErMg6Nz96_1),.din(G384_fa_));
	jspl3 jspl3_w_G387_0(.douta(w_G387_0[0]),.doutb(w_G387_0[1]),.doutc(w_dff_A_0lqkBuEO4_2),.din(G387_fa_));
	jspl3 jspl3_w_n72_0(.douta(w_n72_0[0]),.doutb(w_dff_A_Tuc3xxEz9_1),.doutc(w_dff_A_b1BQvMIP9_2),.din(n72));
	jspl jspl_w_n72_1(.douta(w_n72_1[0]),.doutb(w_dff_A_KZg6e6nu4_1),.din(w_n72_0[0]));
	jspl3 jspl3_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.doutc(w_dff_A_Bkc40ouF1_2),.din(n73));
	jspl3 jspl3_w_n73_1(.douta(w_n73_1[0]),.doutb(w_dff_A_3K811a2e5_1),.doutc(w_n73_1[2]),.din(w_n73_0[0]));
	jspl3 jspl3_w_n73_2(.douta(w_dff_A_cOaJiuwx8_0),.doutb(w_n73_2[1]),.doutc(w_dff_A_tYBCD6H65_2),.din(w_n73_0[1]));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_dff_A_Q7OJ38FA2_1),.doutc(w_dff_A_j7xJR0ii1_2),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_dff_A_Zz5ApCGF9_1),.doutc(w_dff_A_efmkBkH97_2),.din(n75));
	jspl jspl_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.din(w_n75_0[0]));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.din(n76));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl3 jspl3_w_n79_0(.douta(w_dff_A_RA2zgpyC4_0),.doutb(w_n79_0[1]),.doutc(w_n79_0[2]),.din(n79));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_dff_A_aqb3i7Wl7_1),.doutc(w_dff_A_zOTSQUUw9_2),.din(n80));
	jspl jspl_w_n80_1(.douta(w_n80_1[0]),.doutb(w_n80_1[1]),.din(w_n80_0[0]));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_ySZaPlsh8_0),.doutb(w_n85_0[1]),.doutc(w_dff_A_migydITg8_2),.din(n85));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n88_0(.douta(w_n88_0[0]),.doutb(w_dff_A_szOXg0XM3_1),.doutc(w_dff_A_k4uqZuK57_2),.din(n88));
	jspl jspl_w_n88_1(.douta(w_n88_1[0]),.doutb(w_n88_1[1]),.din(w_n88_0[0]));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_dff_A_4xdXvQ5i9_1),.doutc(w_n91_0[2]),.din(n91));
	jspl3 jspl3_w_n91_1(.douta(w_dff_A_dERL1esi8_0),.doutb(w_n91_1[1]),.doutc(w_n91_1[2]),.din(w_n91_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n97_0(.douta(w_dff_A_627OoBlb1_0),.doutb(w_n97_0[1]),.doutc(w_n97_0[2]),.din(n97));
	jspl3 jspl3_w_n97_1(.douta(w_n97_1[0]),.doutb(w_dff_A_LCf4WESU9_1),.doutc(w_n97_1[2]),.din(w_n97_0[0]));
	jspl jspl_w_n97_2(.douta(w_n97_2[0]),.doutb(w_n97_2[1]),.din(w_n97_0[1]));
	jspl3 jspl3_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.doutc(w_n98_0[2]),.din(n98));
	jspl3 jspl3_w_n98_1(.douta(w_dff_A_BhSiJ9au1_0),.doutb(w_dff_A_Kgb8rgQL7_1),.doutc(w_n98_1[2]),.din(w_n98_0[0]));
	jspl jspl_w_n98_2(.douta(w_dff_A_b2IsJz1y0_0),.doutb(w_n98_2[1]),.din(w_n98_0[1]));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_iEPVGXbc1_1),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n105_0(.douta(w_dff_A_Y2GmgOsp7_0),.doutb(w_n105_0[1]),.doutc(w_dff_A_m5Q5lf740_2),.din(n105));
	jspl3 jspl3_w_n105_1(.douta(w_dff_A_n0VUd9i96_0),.doutb(w_n105_1[1]),.doutc(w_dff_A_sWlRsFGD9_2),.din(w_n105_0[0]));
	jspl jspl_w_n105_2(.douta(w_n105_2[0]),.doutb(w_n105_2[1]),.din(w_n105_0[1]));
	jspl jspl_w_n106_0(.douta(w_dff_A_5OOqrkCz7_0),.doutb(w_n106_0[1]),.din(n106));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl3 jspl3_w_n112_3(.douta(w_dff_A_BXlryQIW5_0),.doutb(w_dff_A_iUA9Ib5T0_1),.doutc(w_n112_3[2]),.din(w_n112_0[2]));
	jspl3 jspl3_w_n112_4(.douta(w_dff_A_iYKKcq6s5_0),.doutb(w_dff_A_epM4ApjK4_1),.doutc(w_n112_4[2]),.din(w_n112_1[0]));
	jspl3 jspl3_w_n112_5(.douta(w_n112_5[0]),.doutb(w_n112_5[1]),.doutc(w_dff_A_fdHaWDMG5_2),.din(w_n112_1[1]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.doutc(w_n113_0[2]),.din(n113));
	jspl3 jspl3_w_n113_1(.douta(w_dff_A_jXlgNbp25_0),.doutb(w_dff_A_ppYdNBXJ7_1),.doutc(w_n113_1[2]),.din(w_n113_0[0]));
	jspl3 jspl3_w_n113_2(.douta(w_n113_2[0]),.doutb(w_n113_2[1]),.doutc(w_n113_2[2]),.din(w_n113_0[1]));
	jspl jspl_w_n113_3(.douta(w_n113_3[0]),.doutb(w_n113_3[1]),.din(w_n113_0[2]));
	jspl3 jspl3_w_n114_0(.douta(w_n114_0[0]),.doutb(w_dff_A_ZwyCD0fH4_1),.doutc(w_n114_0[2]),.din(n114));
	jspl3 jspl3_w_n114_1(.douta(w_dff_A_wjUr3Scq4_0),.doutb(w_n114_1[1]),.doutc(w_n114_1[2]),.din(w_n114_0[0]));
	jspl3 jspl3_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.doutc(w_dff_A_E0S8gfdK9_2),.din(n115));
	jspl jspl_w_n115_1(.douta(w_n115_1[0]),.doutb(w_n115_1[1]),.din(w_n115_0[0]));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_dff_A_L1JiYjgh4_1),.din(n116));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl3 jspl3_w_n121_0(.douta(w_dff_A_byAoXEJY4_0),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.doutc(w_n122_0[2]),.din(n122));
	jspl jspl_w_n122_1(.douta(w_n122_1[0]),.doutb(w_n122_1[1]),.din(w_n122_0[0]));
	jspl3 jspl3_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.doutc(w_n123_0[2]),.din(n123));
	jspl3 jspl3_w_n123_1(.douta(w_n123_1[0]),.doutb(w_n123_1[1]),.doutc(w_n123_1[2]),.din(w_n123_0[0]));
	jspl jspl_w_n131_0(.douta(w_dff_A_yZq3Id2l3_0),.doutb(w_n131_0[1]),.din(n131));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_dff_A_oOUnMqgv3_1),.din(n135));
	jspl3 jspl3_w_n137_0(.douta(w_n137_0[0]),.doutb(w_n137_0[1]),.doutc(w_n137_0[2]),.din(n137));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(w_dff_B_TASpClio3_2));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_nLw5oAua9_1),.doutc(w_dff_A_7t4Mkimw9_2),.din(n146));
	jspl3 jspl3_w_n146_1(.douta(w_n146_1[0]),.doutb(w_dff_A_pmUtW7ki4_1),.doutc(w_dff_A_7hze8iR17_2),.din(w_n146_0[0]));
	jspl3 jspl3_w_n146_2(.douta(w_n146_2[0]),.doutb(w_n146_2[1]),.doutc(w_n146_2[2]),.din(w_n146_0[1]));
	jspl3 jspl3_w_n146_3(.douta(w_n146_3[0]),.doutb(w_n146_3[1]),.doutc(w_n146_3[2]),.din(w_n146_0[2]));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_dff_A_7tAftBDu2_1),.doutc(w_dff_A_9AnwOYgO0_2),.din(n147));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_dff_A_6yVyZMe51_0),.doutb(w_dff_A_GjQKIh0o2_1),.doutc(w_n148_1[2]),.din(w_n148_0[0]));
	jspl3 jspl3_w_n148_2(.douta(w_n148_2[0]),.doutb(w_n148_2[1]),.doutc(w_n148_2[2]),.din(w_n148_0[1]));
	jspl3 jspl3_w_n148_3(.douta(w_dff_A_xk3kCVKM2_0),.doutb(w_n148_3[1]),.doutc(w_dff_A_ZBccMnZ21_2),.din(w_n148_0[2]));
	jspl3 jspl3_w_n148_4(.douta(w_n148_4[0]),.doutb(w_n148_4[1]),.doutc(w_n148_4[2]),.din(w_n148_1[0]));
	jspl3 jspl3_w_n148_5(.douta(w_n148_5[0]),.doutb(w_dff_A_Dg7xY4Fv9_1),.doutc(w_dff_A_qFR6XBNy6_2),.din(w_n148_1[1]));
	jspl3 jspl3_w_n148_6(.douta(w_n148_6[0]),.doutb(w_n148_6[1]),.doutc(w_n148_6[2]),.din(w_n148_1[2]));
	jspl3 jspl3_w_n148_7(.douta(w_n148_7[0]),.doutb(w_n148_7[1]),.doutc(w_n148_7[2]),.din(w_n148_2[0]));
	jspl3 jspl3_w_n148_8(.douta(w_n148_8[0]),.doutb(w_dff_A_xLbWa16Q8_1),.doutc(w_n148_8[2]),.din(w_n148_2[1]));
	jspl3 jspl3_w_n148_9(.douta(w_n148_9[0]),.doutb(w_n148_9[1]),.doutc(w_n148_9[2]),.din(w_n148_2[2]));
	jspl3 jspl3_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.doutc(w_n149_0[2]),.din(n149));
	jspl3 jspl3_w_n149_1(.douta(w_n149_1[0]),.doutb(w_dff_A_Xyt08d892_1),.doutc(w_n149_1[2]),.din(w_n149_0[0]));
	jspl jspl_w_n149_2(.douta(w_dff_A_F456LDT18_0),.doutb(w_n149_2[1]),.din(w_n149_0[1]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_HThULbC84_1),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_dff_A_3G10Qk7Z1_1),.doutc(w_dff_A_MFQzdhd58_2),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_n151_2[0]),.doutb(w_n151_2[1]),.doutc(w_n151_2[2]),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_dff_A_q6XlzzcL2_0),.doutb(w_dff_A_puhMWKVZ2_1),.doutc(w_n151_3[2]),.din(w_n151_0[2]));
	jspl3 jspl3_w_n151_4(.douta(w_n151_4[0]),.doutb(w_n151_4[1]),.doutc(w_dff_A_YpwrCHtT1_2),.din(w_n151_1[0]));
	jspl3 jspl3_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.doutc(w_n152_0[2]),.din(n152));
	jspl3 jspl3_w_n152_1(.douta(w_n152_1[0]),.doutb(w_n152_1[1]),.doutc(w_n152_1[2]),.din(w_n152_0[0]));
	jspl3 jspl3_w_n152_2(.douta(w_n152_2[0]),.doutb(w_n152_2[1]),.doutc(w_n152_2[2]),.din(w_n152_0[1]));
	jspl jspl_w_n152_3(.douta(w_n152_3[0]),.doutb(w_n152_3[1]),.din(w_n152_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(n154));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl3 jspl3_w_n155_1(.douta(w_n155_1[0]),.doutb(w_n155_1[1]),.doutc(w_n155_1[2]),.din(w_n155_0[0]));
	jspl3 jspl3_w_n155_2(.douta(w_n155_2[0]),.doutb(w_n155_2[1]),.doutc(w_n155_2[2]),.din(w_n155_0[1]));
	jspl jspl_w_n155_3(.douta(w_n155_3[0]),.doutb(w_n155_3[1]),.din(w_n155_0[2]));
	jspl3 jspl3_w_n157_0(.douta(w_dff_A_0vFtVP2w7_0),.doutb(w_n157_0[1]),.doutc(w_dff_A_wPVodFzS2_2),.din(n157));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_dff_A_JyxtuiHL2_2),.din(n161));
	jspl jspl_w_n161_1(.douta(w_n161_1[0]),.doutb(w_n161_1[1]),.din(w_n161_0[0]));
	jspl3 jspl3_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.doutc(w_n162_0[2]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_dff_A_1pje1mkK3_0),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_dff_A_mEmlEm6s2_1),.doutc(w_dff_A_pg5ld5f74_2),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_dff_A_vdMaJsxe1_2),.din(w_n166_0[1]));
	jspl jspl_w_n166_3(.douta(w_dff_A_4s0TyoYc9_0),.doutb(w_n166_3[1]),.din(w_n166_0[2]));
	jspl3 jspl3_w_n170_0(.douta(w_dff_A_5F5KU4zg0_0),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(w_dff_B_EMpldElG0_2));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_dff_A_B5O5RWX09_1),.doutc(w_dff_A_STJGStVK6_2),.din(n179));
	jspl3 jspl3_w_n179_1(.douta(w_n179_1[0]),.doutb(w_n179_1[1]),.doutc(w_n179_1[2]),.din(w_n179_0[0]));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.doutc(w_n185_0[2]),.din(n185));
	jspl3 jspl3_w_n185_1(.douta(w_n185_1[0]),.doutb(w_n185_1[1]),.doutc(w_dff_A_se3X5d4g7_2),.din(w_n185_0[0]));
	jspl3 jspl3_w_n185_2(.douta(w_n185_2[0]),.doutb(w_dff_A_p17GX4UV7_1),.doutc(w_n185_2[2]),.din(w_n185_0[1]));
	jspl3 jspl3_w_n185_3(.douta(w_n185_3[0]),.doutb(w_n185_3[1]),.doutc(w_n185_3[2]),.din(w_n185_0[2]));
	jspl3 jspl3_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.doutc(w_dff_A_lQeOl7ID9_2),.din(n189));
	jspl3 jspl3_w_n189_1(.douta(w_n189_1[0]),.doutb(w_dff_A_vs3ZJwGa9_1),.doutc(w_n189_1[2]),.din(w_n189_0[0]));
	jspl jspl_w_n189_2(.douta(w_dff_A_3zB2eNgH8_0),.doutb(w_n189_2[1]),.din(w_n189_0[1]));
	jspl3 jspl3_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.doutc(w_n190_0[2]),.din(n190));
	jspl3 jspl3_w_n190_1(.douta(w_n190_1[0]),.doutb(w_dff_A_JQXtkOfm4_1),.doutc(w_n190_1[2]),.din(w_n190_0[0]));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_dff_A_r7UpT6j45_0),.doutb(w_n196_0[1]),.doutc(w_dff_A_jYX9ILcw5_2),.din(w_dff_B_3i5XDcRf5_3));
	jspl3 jspl3_w_n196_1(.douta(w_dff_A_jKKD54u20_0),.doutb(w_dff_A_g5QmKHKA5_1),.doutc(w_n196_1[2]),.din(w_n196_0[0]));
	jspl3 jspl3_w_n196_2(.douta(w_dff_A_AFPinfUT7_0),.doutb(w_dff_A_6560CfKM2_1),.doutc(w_n196_2[2]),.din(w_n196_0[1]));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_n197_1[0]),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n199_1(.douta(w_n199_1[0]),.doutb(w_n199_1[1]),.din(w_n199_0[0]));
	jspl jspl_w_n201_0(.douta(w_dff_A_OaCuvt4G3_0),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n205_0(.douta(w_dff_A_UiqxvAbc6_0),.doutb(w_n205_0[1]),.din(w_dff_B_XO0IhvhS0_2));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl3 jspl3_w_n210_0(.douta(w_dff_A_D5ioe1ut3_0),.doutb(w_n210_0[1]),.doutc(w_n210_0[2]),.din(n210));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_dff_A_t2h3zT050_1),.din(n213));
	jspl jspl_w_n214_0(.douta(w_n214_0[0]),.doutb(w_dff_A_aeTsSMyu8_1),.din(n214));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl3 jspl3_w_n221_0(.douta(w_dff_A_3JjXdUhZ0_0),.doutb(w_dff_A_DwDP3ax58_1),.doutc(w_n221_0[2]),.din(n221));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_dff_A_LxrKDjch3_1),.din(n228));
	jspl3 jspl3_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.doutc(w_n229_0[2]),.din(n229));
	jspl jspl_w_n230_0(.douta(w_dff_A_l2Iq00g77_0),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.doutc(w_n231_0[2]),.din(n231));
	jspl3 jspl3_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.doutc(w_n234_0[2]),.din(n234));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(n241));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl jspl_w_n246_1(.douta(w_n246_1[0]),.doutb(w_n246_1[1]),.din(w_n246_0[0]));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_Vq8gzTDt7_2));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_dff_A_0eUypARF3_1),.din(n255));
	jspl jspl_w_n257_0(.douta(w_dff_A_kStMTVvA0_0),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n259_0(.douta(w_dff_A_Fhdl4g5f6_0),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n262_0(.douta(w_dff_A_XQVY9OJj8_0),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.doutc(w_n269_1[2]),.din(w_n269_0[0]));
	jspl jspl_w_n270_0(.douta(w_dff_A_ep0BYdZp7_0),.doutb(w_n270_0[1]),.din(w_dff_B_b3AJGpTB4_2));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_n271_1[0]),.doutb(w_n271_1[1]),.doutc(w_n271_1[2]),.din(w_n271_0[0]));
	jspl3 jspl3_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_OOS4yCBy7_1),.doutc(w_n274_0[2]),.din(n274));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(n278));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(n279));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_dff_A_BA5H7OT31_1),.din(n281));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n288_1(.douta(w_n288_1[0]),.doutb(w_n288_1[1]),.din(w_n288_0[0]));
	jspl jspl_w_n296_0(.douta(w_dff_A_diXvnU778_0),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n298_0(.douta(w_dff_A_Mcvi3e8f7_0),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_dff_A_Vd13r1yy1_1),.din(n300));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_3GIROOwX0_1),.din(n303));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_dff_A_gxRNkctz1_1),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n334_0(.douta(w_dff_A_X9o9EagP8_0),.doutb(w_n334_0[1]),.din(n334));
	jspl jspl_w_n339_0(.douta(w_dff_A_cYysVxzc5_0),.doutb(w_n339_0[1]),.din(n339));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl jspl_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.din(w_n355_0[0]));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_dff_A_vPeGR7Cb2_1),.din(n374));
	jspl jspl_w_n381_0(.douta(w_n381_0[0]),.doutb(w_n381_0[1]),.din(n381));
	jspl3 jspl3_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.doutc(w_n382_0[2]),.din(n382));
	jspl jspl_w_n382_1(.douta(w_n382_1[0]),.doutb(w_n382_1[1]),.din(w_n382_0[0]));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl jspl_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(w_dff_B_UiuHreiG2_2));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_dff_A_qexzSkda6_1),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n407_0(.douta(w_n407_0[0]),.doutb(w_dff_A_UHbBUwz78_1),.doutc(w_dff_A_a4r3djru3_2),.din(n407));
	jspl3 jspl3_w_n407_1(.douta(w_dff_A_BmjXFYCM9_0),.doutb(w_dff_A_SoJMaa6U8_1),.doutc(w_n407_1[2]),.din(w_n407_0[0]));
	jspl jspl_w_n407_2(.douta(w_n407_2[0]),.doutb(w_n407_2[1]),.din(w_n407_0[1]));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(n412));
	jspl3 jspl3_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jspl jspl_w_n420_1(.douta(w_n420_1[0]),.doutb(w_n420_1[1]),.din(w_n420_0[0]));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_dff_A_fSXR1oKu2_1),.doutc(w_dff_A_qItjlHxo7_2),.din(n425));
	jspl3 jspl3_w_n425_1(.douta(w_dff_A_8ee8hWvj7_0),.doutb(w_dff_A_rmQ2P6ob1_1),.doutc(w_n425_1[2]),.din(w_n425_0[0]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl jspl_w_n430_0(.douta(w_dff_A_NVMS29z04_0),.doutb(w_n430_0[1]),.din(w_dff_B_aFDTMb6B2_2));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_dff_A_Ql0JBR2b8_1),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_dff_A_KWWvRnfy9_1),.doutc(w_n439_0[2]),.din(n439));
	jspl jspl_w_n439_1(.douta(w_n439_1[0]),.doutb(w_n439_1[1]),.din(w_n439_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl3 jspl3_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.doutc(w_n455_0[2]),.din(n455));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(n474));
	jspl jspl_w_n475_0(.douta(w_n475_0[0]),.doutb(w_n475_0[1]),.din(n475));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(n479));
	jspl jspl_w_n483_0(.douta(w_dff_A_sYv13dku0_0),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl3 jspl3_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.doutc(w_n492_0[2]),.din(n492));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n516_0(.douta(w_dff_A_E2BCCOSl0_0),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n519_0(.douta(w_n519_0[0]),.doutb(w_dff_A_I4QRRSBC3_1),.doutc(w_dff_A_RqxBxNm63_2),.din(n519));
	jspl3 jspl3_w_n519_1(.douta(w_dff_A_cxfiEA5b1_0),.doutb(w_n519_1[1]),.doutc(w_n519_1[2]),.din(w_n519_0[0]));
	jspl jspl_w_n523_0(.douta(w_dff_A_ZsxRKSK08_0),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_dff_A_sJNSF0Ru5_1),.din(n524));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_dff_A_freTjB7M9_1),.din(n532));
	jspl jspl_w_n534_0(.douta(w_dff_A_enXX1quV3_0),.doutb(w_n534_0[1]),.din(n534));
	jspl3 jspl3_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.doutc(w_n536_0[2]),.din(n536));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_dff_A_fcI5NC2f2_1),.din(n541));
	jspl3 jspl3_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.doutc(w_n542_0[2]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n548_0(.douta(w_dff_A_Tgsmx2AP1_0),.doutb(w_n548_0[1]),.doutc(w_n548_0[2]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl3 jspl3_w_n552_0(.douta(w_n552_0[0]),.doutb(w_dff_A_l6eqF4jg5_1),.doutc(w_dff_A_Q5eaKtoA0_2),.din(n552));
	jspl jspl_w_n552_1(.douta(w_n552_1[0]),.doutb(w_n552_1[1]),.din(w_n552_0[0]));
	jspl3 jspl3_w_n553_0(.douta(w_dff_A_6ibv6KxW6_0),.doutb(w_n553_0[1]),.doutc(w_dff_A_MFGIaPWm2_2),.din(n553));
	jspl3 jspl3_w_n553_1(.douta(w_n553_1[0]),.doutb(w_n553_1[1]),.doutc(w_n553_1[2]),.din(w_n553_0[0]));
	jspl3 jspl3_w_n553_2(.douta(w_dff_A_KgJyM3XM4_0),.doutb(w_dff_A_H6Iufzoy3_1),.doutc(w_n553_2[2]),.din(w_n553_0[1]));
	jspl3 jspl3_w_n554_0(.douta(w_dff_A_LEHBkyB51_0),.doutb(w_dff_A_hKnFbtoY1_1),.doutc(w_n554_0[2]),.din(w_dff_B_msZ2tOuf0_3));
	jspl3 jspl3_w_n554_1(.douta(w_n554_1[0]),.doutb(w_n554_1[1]),.doutc(w_dff_A_6HEAOcvv8_2),.din(w_n554_0[0]));
	jspl3 jspl3_w_n554_2(.douta(w_n554_2[0]),.doutb(w_dff_A_xefzw0Xr8_1),.doutc(w_dff_A_jQrP0qoc7_2),.din(w_n554_0[1]));
	jspl3 jspl3_w_n554_3(.douta(w_n554_3[0]),.doutb(w_dff_A_Dp2CALI72_1),.doutc(w_dff_A_AQIsk6hs2_2),.din(w_n554_0[2]));
	jspl jspl_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.din(w_dff_B_e8e0s9Tw7_2));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl3 jspl3_w_n563_0(.douta(w_n563_0[0]),.doutb(w_dff_A_jYdxiSC18_1),.doutc(w_dff_A_OgC83iMD6_2),.din(n563));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_VOB1MuIG0_1),.din(n564));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(w_dff_B_S2SNhrZX6_2));
	jspl jspl_w_n567_0(.douta(w_dff_A_7vTYN9o84_0),.doutb(w_n567_0[1]),.din(n567));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_n571_0[2]),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n576_1(.douta(w_n576_1[0]),.doutb(w_n576_1[1]),.din(w_n576_0[0]));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_dff_A_NeBlkTsm6_2),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n589_0(.douta(w_n589_0[0]),.doutb(w_n589_0[1]),.doutc(w_n589_0[2]),.din(n589));
	jspl3 jspl3_w_n589_1(.douta(w_dff_A_Ci1lgWHE0_0),.doutb(w_n589_1[1]),.doutc(w_n589_1[2]),.din(w_n589_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_dff_A_6R3kS48e5_1),.doutc(w_dff_A_Et3t0F1f3_2),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_dff_A_sgipNb9P9_0),.doutb(w_n592_0[1]),.doutc(w_dff_A_u2zHD1e91_2),.din(n592));
	jspl3 jspl3_w_n592_1(.douta(w_dff_A_7zXK7Z0j7_0),.doutb(w_dff_A_b1O6bxue3_1),.doutc(w_n592_1[2]),.din(w_n592_0[0]));
	jspl jspl_w_n592_2(.douta(w_n592_2[0]),.doutb(w_n592_2[1]),.din(w_n592_0[1]));
	jspl3 jspl3_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.doutc(w_n593_0[2]),.din(n593));
	jspl jspl_w_n602_0(.douta(w_dff_A_4dWGbo2M2_0),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n603_0(.douta(w_dff_A_WuP3LnJy6_0),.doutb(w_n603_0[1]),.doutc(w_dff_A_v2epItUz6_2),.din(n603));
	jspl3 jspl3_w_n603_1(.douta(w_dff_A_aEkXezqP0_0),.doutb(w_n603_1[1]),.doutc(w_n603_1[2]),.din(w_n603_0[0]));
	jspl jspl_w_n603_2(.douta(w_dff_A_Cc4Z5JpJ0_0),.doutb(w_n603_2[1]),.din(w_n603_0[1]));
	jspl3 jspl3_w_n604_0(.douta(w_dff_A_foqsK1iu2_0),.doutb(w_n604_0[1]),.doutc(w_dff_A_K3AGBwzM7_2),.din(n604));
	jspl3 jspl3_w_n604_1(.douta(w_dff_A_tjhWdLt39_0),.doutb(w_n604_1[1]),.doutc(w_dff_A_4flnU5zK4_2),.din(w_n604_0[0]));
	jspl jspl_w_n604_2(.douta(w_dff_A_7dGQOBZh0_0),.doutb(w_n604_2[1]),.din(w_n604_0[1]));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_dff_A_tv0YYWOD6_2),.din(w_n605_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_dff_A_yUSiJE2a0_1),.doutc(w_dff_A_YCIlTHLf2_2),.din(n608));
	jspl3 jspl3_w_n608_1(.douta(w_dff_A_A0bUwg7l5_0),.doutb(w_n608_1[1]),.doutc(w_dff_A_W5fxPdRt2_2),.din(w_n608_0[0]));
	jspl3 jspl3_w_n612_0(.douta(w_n612_0[0]),.doutb(w_dff_A_KIRTliAh7_1),.doutc(w_n612_0[2]),.din(n612));
	jspl3 jspl3_w_n612_1(.douta(w_dff_A_iO2LrXBq8_0),.doutb(w_dff_A_iA6ky1Cq2_1),.doutc(w_n612_1[2]),.din(w_n612_0[0]));
	jspl3 jspl3_w_n612_2(.douta(w_n612_2[0]),.doutb(w_n612_2[1]),.doutc(w_n612_2[2]),.din(w_n612_0[1]));
	jspl3 jspl3_w_n612_3(.douta(w_dff_A_eDV0uxhS1_0),.doutb(w_n612_3[1]),.doutc(w_dff_A_DNgoaVjB0_2),.din(w_n612_0[2]));
	jspl jspl_w_n612_4(.douta(w_n612_4[0]),.doutb(w_dff_A_pftuPXJG7_1),.din(w_n612_1[0]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl jspl_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.din(w_n613_0[0]));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_dff_A_jajZH1VY4_1),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl3 jspl3_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.doutc(w_n617_1[2]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n617_2(.douta(w_n617_2[0]),.doutb(w_n617_2[1]),.doutc(w_n617_2[2]),.din(w_n617_0[1]));
	jspl3 jspl3_w_n617_3(.douta(w_n617_3[0]),.doutb(w_n617_3[1]),.doutc(w_n617_3[2]),.din(w_n617_0[2]));
	jspl3 jspl3_w_n617_4(.douta(w_n617_4[0]),.doutb(w_n617_4[1]),.doutc(w_n617_4[2]),.din(w_n617_1[0]));
	jspl3 jspl3_w_n617_5(.douta(w_n617_5[0]),.doutb(w_n617_5[1]),.doutc(w_n617_5[2]),.din(w_n617_1[1]));
	jspl jspl_w_n617_6(.douta(w_n617_6[0]),.doutb(w_n617_6[1]),.din(w_n617_1[2]));
	jspl jspl_w_n619_0(.douta(w_dff_A_4V9nTFmm2_0),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl3 jspl3_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.doutc(w_n623_0[2]),.din(n623));
	jspl3 jspl3_w_n623_1(.douta(w_n623_1[0]),.doutb(w_n623_1[1]),.doutc(w_n623_1[2]),.din(w_n623_0[0]));
	jspl3 jspl3_w_n623_2(.douta(w_n623_2[0]),.doutb(w_n623_2[1]),.doutc(w_n623_2[2]),.din(w_n623_0[1]));
	jspl3 jspl3_w_n623_3(.douta(w_n623_3[0]),.doutb(w_n623_3[1]),.doutc(w_n623_3[2]),.din(w_n623_0[2]));
	jspl3 jspl3_w_n623_4(.douta(w_n623_4[0]),.doutb(w_n623_4[1]),.doutc(w_n623_4[2]),.din(w_n623_1[0]));
	jspl jspl_w_n623_5(.douta(w_n623_5[0]),.doutb(w_n623_5[1]),.din(w_n623_1[1]));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(n626));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl3 jspl3_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.doutc(w_n627_1[2]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n627_2(.douta(w_n627_2[0]),.doutb(w_n627_2[1]),.doutc(w_n627_2[2]),.din(w_n627_0[1]));
	jspl3 jspl3_w_n627_3(.douta(w_n627_3[0]),.doutb(w_n627_3[1]),.doutc(w_n627_3[2]),.din(w_n627_0[2]));
	jspl3 jspl3_w_n627_4(.douta(w_n627_4[0]),.doutb(w_n627_4[1]),.doutc(w_n627_4[2]),.din(w_n627_1[0]));
	jspl3 jspl3_w_n627_5(.douta(w_n627_5[0]),.doutb(w_n627_5[1]),.doutc(w_n627_5[2]),.din(w_n627_1[1]));
	jspl3 jspl3_w_n627_6(.douta(w_n627_6[0]),.doutb(w_n627_6[1]),.doutc(w_n627_6[2]),.din(w_n627_1[2]));
	jspl jspl_w_n627_7(.douta(w_n627_7[0]),.doutb(w_n627_7[1]),.din(w_n627_2[0]));
	jspl3 jspl3_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.doutc(w_n631_0[2]),.din(n631));
	jspl3 jspl3_w_n631_1(.douta(w_n631_1[0]),.doutb(w_n631_1[1]),.doutc(w_n631_1[2]),.din(w_n631_0[0]));
	jspl3 jspl3_w_n631_2(.douta(w_n631_2[0]),.doutb(w_n631_2[1]),.doutc(w_n631_2[2]),.din(w_n631_0[1]));
	jspl3 jspl3_w_n631_3(.douta(w_n631_3[0]),.doutb(w_n631_3[1]),.doutc(w_n631_3[2]),.din(w_n631_0[2]));
	jspl3 jspl3_w_n631_4(.douta(w_n631_4[0]),.doutb(w_n631_4[1]),.doutc(w_n631_4[2]),.din(w_n631_1[0]));
	jspl3 jspl3_w_n631_5(.douta(w_n631_5[0]),.doutb(w_n631_5[1]),.doutc(w_n631_5[2]),.din(w_n631_1[1]));
	jspl3 jspl3_w_n631_6(.douta(w_n631_6[0]),.doutb(w_n631_6[1]),.doutc(w_n631_6[2]),.din(w_n631_1[2]));
	jspl jspl_w_n631_7(.douta(w_n631_7[0]),.doutb(w_n631_7[1]),.din(w_n631_2[0]));
	jspl3 jspl3_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.doutc(w_n634_0[2]),.din(n634));
	jspl3 jspl3_w_n634_1(.douta(w_n634_1[0]),.doutb(w_n634_1[1]),.doutc(w_n634_1[2]),.din(w_n634_0[0]));
	jspl3 jspl3_w_n634_2(.douta(w_n634_2[0]),.doutb(w_n634_2[1]),.doutc(w_n634_2[2]),.din(w_n634_0[1]));
	jspl3 jspl3_w_n634_3(.douta(w_n634_3[0]),.doutb(w_n634_3[1]),.doutc(w_n634_3[2]),.din(w_n634_0[2]));
	jspl jspl_w_n634_4(.douta(w_n634_4[0]),.doutb(w_n634_4[1]),.din(w_n634_1[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n636_1(.douta(w_n636_1[0]),.doutb(w_n636_1[1]),.doutc(w_n636_1[2]),.din(w_n636_0[0]));
	jspl3 jspl3_w_n636_2(.douta(w_n636_2[0]),.doutb(w_n636_2[1]),.doutc(w_n636_2[2]),.din(w_n636_0[1]));
	jspl3 jspl3_w_n636_3(.douta(w_n636_3[0]),.doutb(w_n636_3[1]),.doutc(w_n636_3[2]),.din(w_n636_0[2]));
	jspl3 jspl3_w_n636_4(.douta(w_n636_4[0]),.doutb(w_n636_4[1]),.doutc(w_n636_4[2]),.din(w_n636_1[0]));
	jspl3 jspl3_w_n636_5(.douta(w_n636_5[0]),.doutb(w_n636_5[1]),.doutc(w_n636_5[2]),.din(w_n636_1[1]));
	jspl3 jspl3_w_n636_6(.douta(w_n636_6[0]),.doutb(w_n636_6[1]),.doutc(w_n636_6[2]),.din(w_n636_1[2]));
	jspl jspl_w_n636_7(.douta(w_n636_7[0]),.doutb(w_n636_7[1]),.din(w_n636_2[0]));
	jspl jspl_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.din(n639));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl3 jspl3_w_n640_2(.douta(w_n640_2[0]),.doutb(w_n640_2[1]),.doutc(w_n640_2[2]),.din(w_n640_0[1]));
	jspl3 jspl3_w_n640_3(.douta(w_n640_3[0]),.doutb(w_n640_3[1]),.doutc(w_n640_3[2]),.din(w_n640_0[2]));
	jspl3 jspl3_w_n640_4(.douta(w_n640_4[0]),.doutb(w_n640_4[1]),.doutc(w_n640_4[2]),.din(w_n640_1[0]));
	jspl3 jspl3_w_n640_5(.douta(w_n640_5[0]),.doutb(w_n640_5[1]),.doutc(w_n640_5[2]),.din(w_n640_1[1]));
	jspl3 jspl3_w_n640_6(.douta(w_n640_6[0]),.doutb(w_n640_6[1]),.doutc(w_n640_6[2]),.din(w_n640_1[2]));
	jspl jspl_w_n640_7(.douta(w_n640_7[0]),.doutb(w_n640_7[1]),.din(w_n640_2[0]));
	jspl3 jspl3_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.doutc(w_n642_0[2]),.din(n642));
	jspl3 jspl3_w_n642_1(.douta(w_n642_1[0]),.doutb(w_n642_1[1]),.doutc(w_n642_1[2]),.din(w_n642_0[0]));
	jspl3 jspl3_w_n642_2(.douta(w_n642_2[0]),.doutb(w_n642_2[1]),.doutc(w_n642_2[2]),.din(w_n642_0[1]));
	jspl3 jspl3_w_n642_3(.douta(w_n642_3[0]),.doutb(w_n642_3[1]),.doutc(w_n642_3[2]),.din(w_n642_0[2]));
	jspl3 jspl3_w_n642_4(.douta(w_n642_4[0]),.doutb(w_n642_4[1]),.doutc(w_n642_4[2]),.din(w_n642_1[0]));
	jspl3 jspl3_w_n642_5(.douta(w_n642_5[0]),.doutb(w_n642_5[1]),.doutc(w_n642_5[2]),.din(w_n642_1[1]));
	jspl3 jspl3_w_n642_6(.douta(w_n642_6[0]),.doutb(w_n642_6[1]),.doutc(w_n642_6[2]),.din(w_n642_1[2]));
	jspl jspl_w_n642_7(.douta(w_n642_7[0]),.doutb(w_n642_7[1]),.din(w_n642_2[0]));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(n654));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl3 jspl3_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.doutc(w_dff_A_cwbGpK2Z3_2),.din(n672));
	jspl jspl_w_n672_1(.douta(w_n672_1[0]),.doutb(w_dff_A_jxubB8fU3_1),.din(w_n672_0[0]));
	jspl3 jspl3_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.doutc(w_n675_0[2]),.din(n675));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(w_dff_B_A4QDMoH20_2));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_dff_A_z8LJpB2h8_1),.din(w_dff_B_z3m5Avw11_2));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_dff_A_GMUR2CPS4_1),.doutc(w_n696_0[2]),.din(n696));
	jspl3 jspl3_w_n696_1(.douta(w_dff_A_y0drUesM0_0),.doutb(w_n696_1[1]),.doutc(w_dff_A_oKWf7lUA3_2),.din(w_n696_0[0]));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.doutc(w_n743_0[2]),.din(n743));
	jspl jspl_w_n743_1(.douta(w_n743_1[0]),.doutb(w_n743_1[1]),.din(w_n743_0[0]));
	jspl jspl_w_n750_0(.douta(w_dff_A_lSMlxxfa2_0),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n754_0(.douta(w_dff_A_v1fpQzmh4_0),.doutb(w_n754_0[1]),.din(n754));
	jspl3 jspl3_w_n758_0(.douta(w_dff_A_reohEdbc8_0),.doutb(w_dff_A_0wblCObB8_1),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n758_1(.douta(w_n758_1[0]),.doutb(w_dff_A_Xh1K58Al4_1),.din(w_n758_0[0]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_dff_A_IUdNnhry2_0),.doutb(w_n760_0[1]),.din(n760));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_dff_A_CfidJJKC8_2),.din(n764));
	jspl3 jspl3_w_n764_1(.douta(w_n764_1[0]),.doutb(w_n764_1[1]),.doutc(w_dff_A_vEisUAsu2_2),.din(w_n764_0[0]));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_n771_0[2]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_dff_A_3432eBZr8_0),.doutb(w_n779_0[1]),.din(n779));
	jspl jspl_w_n797_0(.douta(w_dff_A_R9T0BBH90_0),.doutb(w_n797_0[1]),.din(n797));
	jspl jspl_w_n801_0(.douta(w_dff_A_LdP0sqej6_0),.doutb(w_n801_0[1]),.din(n801));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl3 jspl3_w_n853_0(.douta(w_n853_0[0]),.doutb(w_n853_0[1]),.doutc(w_n853_0[2]),.din(n853));
	jspl3 jspl3_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.doutc(w_n855_0[2]),.din(n855));
	jspl3 jspl3_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.doutc(w_dff_A_h8BRsSgY3_2),.din(n861));
	jspl jspl_w_n861_1(.douta(w_n861_1[0]),.doutb(w_dff_A_miPFumjC5_1),.din(w_n861_0[0]));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.din(n863));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_dff_A_4YM7diBN0_1),.din(n899));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl3 jspl3_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.doutc(w_n937_0[2]),.din(n937));
	jspl jspl_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.din(n940));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_dff_A_0J4OVUoY9_1),.din(n962));
	jspl3 jspl3_w_n988_0(.douta(w_dff_A_aXqDb7Dy9_0),.doutb(w_dff_A_kO1rFbt35_1),.doutc(w_n988_0[2]),.din(n988));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_dff_A_hlvTrcX62_1),.din(n990));
	jspl3 jspl3_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.doutc(w_n991_0[2]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_dff_A_D22jo48r6_1),.din(n999));
	jspl3 jspl3_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.doutc(w_n1001_0[2]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.doutc(w_n1002_0[2]),.din(n1002));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl3 jspl3_w_n1049_0(.douta(w_dff_A_be0PVgZO0_0),.doutb(w_dff_A_RStRHZ5r4_1),.doutc(w_n1049_0[2]),.din(n1049));
	jspl jspl_w_n1052_0(.douta(w_dff_A_Ci7AUCfM4_0),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_dff_A_N46omXvs3_1),.din(n1057));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(n1059));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl3 jspl3_w_n1162_0(.douta(w_n1162_0[0]),.doutb(w_dff_A_hTgHDsrK5_1),.doutc(w_n1162_0[2]),.din(n1162));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(n1164));
	jspl jspl_w_n1172_0(.douta(w_dff_A_lED9eLgz9_0),.doutb(w_n1172_0[1]),.din(n1172));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_dff_A_9rvIgHbL5_1),.din(n1175));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_dff_A_CtVzTCe36_1),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_dff_A_CT01YOIy2_0),.doutb(w_n1184_0[1]),.din(n1184));
	jspl jspl_w_n1187_0(.douta(w_dff_A_kY51oWpU0_0),.doutb(w_n1187_0[1]),.din(n1187));
	jdff dff_B_27IG3dus8_1(.din(n111),.dout(w_dff_B_27IG3dus8_1),.clk(gclk));
	jdff dff_B_brpxkulE2_0(.din(n126),.dout(w_dff_B_brpxkulE2_0),.clk(gclk));
	jdff dff_B_OdmNiY9Q7_0(.din(n125),.dout(w_dff_B_OdmNiY9Q7_0),.clk(gclk));
	jdff dff_A_oKzhe3GQ7_1(.dout(w_n72_1[1]),.din(w_dff_A_oKzhe3GQ7_1),.clk(gclk));
	jdff dff_A_KZg6e6nu4_1(.dout(w_dff_A_oKzhe3GQ7_1),.din(w_dff_A_KZg6e6nu4_1),.clk(gclk));
	jdff dff_A_b2IsJz1y0_0(.dout(w_n98_2[0]),.din(w_dff_A_b2IsJz1y0_0),.clk(gclk));
	jdff dff_B_P1MteBTm6_1(.din(n540),.dout(w_dff_B_P1MteBTm6_1),.clk(gclk));
	jdff dff_B_VcQ3QnV95_0(.din(n597),.dout(w_dff_B_VcQ3QnV95_0),.clk(gclk));
	jdff dff_B_0KF7IW7h5_0(.din(w_dff_B_VcQ3QnV95_0),.dout(w_dff_B_0KF7IW7h5_0),.clk(gclk));
	jdff dff_B_khbgpzw24_0(.din(w_dff_B_0KF7IW7h5_0),.dout(w_dff_B_khbgpzw24_0),.clk(gclk));
	jdff dff_B_UkrzfmdC8_0(.din(w_dff_B_khbgpzw24_0),.dout(w_dff_B_UkrzfmdC8_0),.clk(gclk));
	jdff dff_B_kaCxY0zh4_0(.din(w_dff_B_UkrzfmdC8_0),.dout(w_dff_B_kaCxY0zh4_0),.clk(gclk));
	jdff dff_B_1nhceMPk4_0(.din(w_dff_B_kaCxY0zh4_0),.dout(w_dff_B_1nhceMPk4_0),.clk(gclk));
	jdff dff_B_SHGn3OUc7_0(.din(w_dff_B_1nhceMPk4_0),.dout(w_dff_B_SHGn3OUc7_0),.clk(gclk));
	jdff dff_B_tCOiiRT90_0(.din(w_dff_B_SHGn3OUc7_0),.dout(w_dff_B_tCOiiRT90_0),.clk(gclk));
	jdff dff_B_T8MWrgiF9_0(.din(w_dff_B_tCOiiRT90_0),.dout(w_dff_B_T8MWrgiF9_0),.clk(gclk));
	jdff dff_B_CQkULghC5_0(.din(w_dff_B_T8MWrgiF9_0),.dout(w_dff_B_CQkULghC5_0),.clk(gclk));
	jdff dff_B_EWujXDTd0_0(.din(n596),.dout(w_dff_B_EWujXDTd0_0),.clk(gclk));
	jdff dff_B_LX6rMsV55_0(.din(n795),.dout(w_dff_B_LX6rMsV55_0),.clk(gclk));
	jdff dff_B_0gYPtSiV2_0(.din(w_dff_B_LX6rMsV55_0),.dout(w_dff_B_0gYPtSiV2_0),.clk(gclk));
	jdff dff_B_m3YYBuz63_0(.din(w_dff_B_0gYPtSiV2_0),.dout(w_dff_B_m3YYBuz63_0),.clk(gclk));
	jdff dff_B_xvy5vnMy1_0(.din(w_dff_B_m3YYBuz63_0),.dout(w_dff_B_xvy5vnMy1_0),.clk(gclk));
	jdff dff_B_5L7Inghj0_0(.din(w_dff_B_xvy5vnMy1_0),.dout(w_dff_B_5L7Inghj0_0),.clk(gclk));
	jdff dff_B_rHWr3kVT1_0(.din(w_dff_B_5L7Inghj0_0),.dout(w_dff_B_rHWr3kVT1_0),.clk(gclk));
	jdff dff_B_y3xYfgSg7_0(.din(w_dff_B_rHWr3kVT1_0),.dout(w_dff_B_y3xYfgSg7_0),.clk(gclk));
	jdff dff_B_HMSjkaM36_0(.din(w_dff_B_y3xYfgSg7_0),.dout(w_dff_B_HMSjkaM36_0),.clk(gclk));
	jdff dff_B_XrsLfFOK7_0(.din(w_dff_B_HMSjkaM36_0),.dout(w_dff_B_XrsLfFOK7_0),.clk(gclk));
	jdff dff_B_tNTamC3K6_0(.din(w_dff_B_XrsLfFOK7_0),.dout(w_dff_B_tNTamC3K6_0),.clk(gclk));
	jdff dff_B_9rLj559m2_0(.din(w_dff_B_tNTamC3K6_0),.dout(w_dff_B_9rLj559m2_0),.clk(gclk));
	jdff dff_B_Fy6euJsy2_0(.din(w_dff_B_9rLj559m2_0),.dout(w_dff_B_Fy6euJsy2_0),.clk(gclk));
	jdff dff_B_05mxwore0_0(.din(w_dff_B_Fy6euJsy2_0),.dout(w_dff_B_05mxwore0_0),.clk(gclk));
	jdff dff_B_FkBCJ4Gk0_0(.din(w_dff_B_05mxwore0_0),.dout(w_dff_B_FkBCJ4Gk0_0),.clk(gclk));
	jdff dff_B_17rdGTZ48_0(.din(w_dff_B_FkBCJ4Gk0_0),.dout(w_dff_B_17rdGTZ48_0),.clk(gclk));
	jdff dff_B_mgTPp4yG5_0(.din(w_dff_B_17rdGTZ48_0),.dout(w_dff_B_mgTPp4yG5_0),.clk(gclk));
	jdff dff_B_qqINFvwM6_0(.din(w_dff_B_mgTPp4yG5_0),.dout(w_dff_B_qqINFvwM6_0),.clk(gclk));
	jdff dff_B_07cq4XHF0_1(.din(n791),.dout(w_dff_B_07cq4XHF0_1),.clk(gclk));
	jdff dff_B_oehH8Av27_0(.din(n793),.dout(w_dff_B_oehH8Av27_0),.clk(gclk));
	jdff dff_B_LsPz2THP9_0(.din(w_dff_B_oehH8Av27_0),.dout(w_dff_B_LsPz2THP9_0),.clk(gclk));
	jdff dff_B_eQEFrEFx6_0(.din(n784),.dout(w_dff_B_eQEFrEFx6_0),.clk(gclk));
	jdff dff_B_gbjR7sTU1_0(.din(w_dff_B_eQEFrEFx6_0),.dout(w_dff_B_gbjR7sTU1_0),.clk(gclk));
	jdff dff_B_8e36eyeG0_0(.din(w_dff_B_gbjR7sTU1_0),.dout(w_dff_B_8e36eyeG0_0),.clk(gclk));
	jdff dff_B_iDQYgquA2_0(.din(w_dff_B_8e36eyeG0_0),.dout(w_dff_B_iDQYgquA2_0),.clk(gclk));
	jdff dff_B_S6qopbMi1_0(.din(w_dff_B_iDQYgquA2_0),.dout(w_dff_B_S6qopbMi1_0),.clk(gclk));
	jdff dff_B_y1uw5VNx6_0(.din(w_dff_B_S6qopbMi1_0),.dout(w_dff_B_y1uw5VNx6_0),.clk(gclk));
	jdff dff_B_jNbPZpET7_0(.din(w_dff_B_y1uw5VNx6_0),.dout(w_dff_B_jNbPZpET7_0),.clk(gclk));
	jdff dff_B_90YbSXgM0_0(.din(w_dff_B_jNbPZpET7_0),.dout(w_dff_B_90YbSXgM0_0),.clk(gclk));
	jdff dff_B_HLxDSfFW2_0(.din(w_dff_B_90YbSXgM0_0),.dout(w_dff_B_HLxDSfFW2_0),.clk(gclk));
	jdff dff_B_tZULgeE83_0(.din(w_dff_B_HLxDSfFW2_0),.dout(w_dff_B_tZULgeE83_0),.clk(gclk));
	jdff dff_B_N0U1Ql070_0(.din(w_dff_B_tZULgeE83_0),.dout(w_dff_B_N0U1Ql070_0),.clk(gclk));
	jdff dff_B_5JVTNJGQ0_0(.din(w_dff_B_N0U1Ql070_0),.dout(w_dff_B_5JVTNJGQ0_0),.clk(gclk));
	jdff dff_B_ZqvK0iFu6_0(.din(w_dff_B_5JVTNJGQ0_0),.dout(w_dff_B_ZqvK0iFu6_0),.clk(gclk));
	jdff dff_B_QDRAx9Hn9_0(.din(w_dff_B_ZqvK0iFu6_0),.dout(w_dff_B_QDRAx9Hn9_0),.clk(gclk));
	jdff dff_B_C6syMAPg1_0(.din(w_dff_B_QDRAx9Hn9_0),.dout(w_dff_B_C6syMAPg1_0),.clk(gclk));
	jdff dff_B_9O43Ezeg7_0(.din(w_dff_B_C6syMAPg1_0),.dout(w_dff_B_9O43Ezeg7_0),.clk(gclk));
	jdff dff_B_bvj5x9wr1_0(.din(w_dff_B_9O43Ezeg7_0),.dout(w_dff_B_bvj5x9wr1_0),.clk(gclk));
	jdff dff_A_Wp42wl8u7_1(.dout(w_n116_0[1]),.din(w_dff_A_Wp42wl8u7_1),.clk(gclk));
	jdff dff_A_L1JiYjgh4_1(.dout(w_dff_A_Wp42wl8u7_1),.din(w_dff_A_L1JiYjgh4_1),.clk(gclk));
	jdff dff_B_6KOFtQeg5_0(.din(n780),.dout(w_dff_B_6KOFtQeg5_0),.clk(gclk));
	jdff dff_A_3432eBZr8_0(.dout(w_n779_0[0]),.din(w_dff_A_3432eBZr8_0),.clk(gclk));
	jdff dff_B_meZ7zUbD1_1(.din(n774),.dout(w_dff_B_meZ7zUbD1_1),.clk(gclk));
	jdff dff_A_cxfiEA5b1_0(.dout(w_n519_1[0]),.din(w_dff_A_cxfiEA5b1_0),.clk(gclk));
	jdff dff_B_bxV1Hvf69_1(.din(n1174),.dout(w_dff_B_bxV1Hvf69_1),.clk(gclk));
	jdff dff_B_dCbiIkUu2_1(.din(w_dff_B_bxV1Hvf69_1),.dout(w_dff_B_dCbiIkUu2_1),.clk(gclk));
	jdff dff_B_ltsCm6fP4_1(.din(w_dff_B_dCbiIkUu2_1),.dout(w_dff_B_ltsCm6fP4_1),.clk(gclk));
	jdff dff_B_snMa3UHB8_1(.din(w_dff_B_ltsCm6fP4_1),.dout(w_dff_B_snMa3UHB8_1),.clk(gclk));
	jdff dff_B_86oEXe4D6_1(.din(w_dff_B_snMa3UHB8_1),.dout(w_dff_B_86oEXe4D6_1),.clk(gclk));
	jdff dff_B_EH4oItPu9_1(.din(w_dff_B_86oEXe4D6_1),.dout(w_dff_B_EH4oItPu9_1),.clk(gclk));
	jdff dff_B_hLXk1Tdo1_1(.din(w_dff_B_EH4oItPu9_1),.dout(w_dff_B_hLXk1Tdo1_1),.clk(gclk));
	jdff dff_B_vbuZhOVL4_1(.din(w_dff_B_hLXk1Tdo1_1),.dout(w_dff_B_vbuZhOVL4_1),.clk(gclk));
	jdff dff_B_KvLiyaVF0_1(.din(w_dff_B_vbuZhOVL4_1),.dout(w_dff_B_KvLiyaVF0_1),.clk(gclk));
	jdff dff_B_tmHNNuv62_1(.din(w_dff_B_KvLiyaVF0_1),.dout(w_dff_B_tmHNNuv62_1),.clk(gclk));
	jdff dff_B_5dTyv3FO1_1(.din(w_dff_B_tmHNNuv62_1),.dout(w_dff_B_5dTyv3FO1_1),.clk(gclk));
	jdff dff_B_7R0XxOkQ1_1(.din(w_dff_B_5dTyv3FO1_1),.dout(w_dff_B_7R0XxOkQ1_1),.clk(gclk));
	jdff dff_B_Js4S65zn1_1(.din(w_dff_B_7R0XxOkQ1_1),.dout(w_dff_B_Js4S65zn1_1),.clk(gclk));
	jdff dff_B_BjpQtCIc2_1(.din(w_dff_B_Js4S65zn1_1),.dout(w_dff_B_BjpQtCIc2_1),.clk(gclk));
	jdff dff_B_27XFPe0M5_1(.din(w_dff_B_BjpQtCIc2_1),.dout(w_dff_B_27XFPe0M5_1),.clk(gclk));
	jdff dff_B_WgMwadz85_1(.din(w_dff_B_27XFPe0M5_1),.dout(w_dff_B_WgMwadz85_1),.clk(gclk));
	jdff dff_B_RKoL6UN74_1(.din(w_dff_B_WgMwadz85_1),.dout(w_dff_B_RKoL6UN74_1),.clk(gclk));
	jdff dff_B_At1DnCxB3_1(.din(w_dff_B_RKoL6UN74_1),.dout(w_dff_B_At1DnCxB3_1),.clk(gclk));
	jdff dff_B_x7bO9Ypj8_1(.din(w_dff_B_At1DnCxB3_1),.dout(w_dff_B_x7bO9Ypj8_1),.clk(gclk));
	jdff dff_B_I4BoaXlS4_1(.din(w_dff_B_x7bO9Ypj8_1),.dout(w_dff_B_I4BoaXlS4_1),.clk(gclk));
	jdff dff_B_qSe9mCK36_1(.din(w_dff_B_I4BoaXlS4_1),.dout(w_dff_B_qSe9mCK36_1),.clk(gclk));
	jdff dff_B_8Y0PSoG76_1(.din(w_dff_B_qSe9mCK36_1),.dout(w_dff_B_8Y0PSoG76_1),.clk(gclk));
	jdff dff_B_7CIeihSw2_1(.din(w_dff_B_8Y0PSoG76_1),.dout(w_dff_B_7CIeihSw2_1),.clk(gclk));
	jdff dff_B_RHlzz7bS4_1(.din(w_dff_B_7CIeihSw2_1),.dout(w_dff_B_RHlzz7bS4_1),.clk(gclk));
	jdff dff_B_0GIqr2mo9_1(.din(w_dff_B_RHlzz7bS4_1),.dout(w_dff_B_0GIqr2mo9_1),.clk(gclk));
	jdff dff_B_zk7gRSOB7_1(.din(w_dff_B_0GIqr2mo9_1),.dout(w_dff_B_zk7gRSOB7_1),.clk(gclk));
	jdff dff_A_lED9eLgz9_0(.dout(w_n1172_0[0]),.din(w_dff_A_lED9eLgz9_0),.clk(gclk));
	jdff dff_B_a5t1mwIU9_1(.din(n1166),.dout(w_dff_B_a5t1mwIU9_1),.clk(gclk));
	jdff dff_B_pqHyahDE9_1(.din(w_dff_B_a5t1mwIU9_1),.dout(w_dff_B_pqHyahDE9_1),.clk(gclk));
	jdff dff_B_8PLgku0F9_1(.din(n1186),.dout(w_dff_B_8PLgku0F9_1),.clk(gclk));
	jdff dff_B_YQwWnxHW1_1(.din(w_dff_B_8PLgku0F9_1),.dout(w_dff_B_YQwWnxHW1_1),.clk(gclk));
	jdff dff_B_eOVT77cD4_1(.din(w_dff_B_YQwWnxHW1_1),.dout(w_dff_B_eOVT77cD4_1),.clk(gclk));
	jdff dff_B_EsSZhU0t7_1(.din(w_dff_B_eOVT77cD4_1),.dout(w_dff_B_EsSZhU0t7_1),.clk(gclk));
	jdff dff_B_7W6IxzaU9_1(.din(w_dff_B_EsSZhU0t7_1),.dout(w_dff_B_7W6IxzaU9_1),.clk(gclk));
	jdff dff_B_5pwmVud73_1(.din(w_dff_B_7W6IxzaU9_1),.dout(w_dff_B_5pwmVud73_1),.clk(gclk));
	jdff dff_B_iyKO1Vem0_1(.din(w_dff_B_5pwmVud73_1),.dout(w_dff_B_iyKO1Vem0_1),.clk(gclk));
	jdff dff_B_sY70pu2D3_1(.din(w_dff_B_iyKO1Vem0_1),.dout(w_dff_B_sY70pu2D3_1),.clk(gclk));
	jdff dff_B_FRzAIkLh2_1(.din(w_dff_B_sY70pu2D3_1),.dout(w_dff_B_FRzAIkLh2_1),.clk(gclk));
	jdff dff_B_Rxfz5tES0_1(.din(w_dff_B_FRzAIkLh2_1),.dout(w_dff_B_Rxfz5tES0_1),.clk(gclk));
	jdff dff_B_O3zsCVqI7_1(.din(w_dff_B_Rxfz5tES0_1),.dout(w_dff_B_O3zsCVqI7_1),.clk(gclk));
	jdff dff_B_BBvpIZVz0_1(.din(w_dff_B_O3zsCVqI7_1),.dout(w_dff_B_BBvpIZVz0_1),.clk(gclk));
	jdff dff_B_iYYAhPtH2_1(.din(w_dff_B_BBvpIZVz0_1),.dout(w_dff_B_iYYAhPtH2_1),.clk(gclk));
	jdff dff_B_hJxebwXO2_1(.din(w_dff_B_iYYAhPtH2_1),.dout(w_dff_B_hJxebwXO2_1),.clk(gclk));
	jdff dff_B_1rOe19vF7_1(.din(w_dff_B_hJxebwXO2_1),.dout(w_dff_B_1rOe19vF7_1),.clk(gclk));
	jdff dff_B_Flku22kH6_1(.din(w_dff_B_1rOe19vF7_1),.dout(w_dff_B_Flku22kH6_1),.clk(gclk));
	jdff dff_B_d8xbczx92_1(.din(w_dff_B_Flku22kH6_1),.dout(w_dff_B_d8xbczx92_1),.clk(gclk));
	jdff dff_B_wtKDcpXr5_1(.din(w_dff_B_d8xbczx92_1),.dout(w_dff_B_wtKDcpXr5_1),.clk(gclk));
	jdff dff_B_jiHOXbbj5_1(.din(w_dff_B_wtKDcpXr5_1),.dout(w_dff_B_jiHOXbbj5_1),.clk(gclk));
	jdff dff_B_V6P9iNHF9_1(.din(w_dff_B_jiHOXbbj5_1),.dout(w_dff_B_V6P9iNHF9_1),.clk(gclk));
	jdff dff_B_MZbxAC849_1(.din(w_dff_B_V6P9iNHF9_1),.dout(w_dff_B_MZbxAC849_1),.clk(gclk));
	jdff dff_B_xNCmMBk97_1(.din(w_dff_B_MZbxAC849_1),.dout(w_dff_B_xNCmMBk97_1),.clk(gclk));
	jdff dff_B_bvOcEYhx9_1(.din(w_dff_B_xNCmMBk97_1),.dout(w_dff_B_bvOcEYhx9_1),.clk(gclk));
	jdff dff_B_Sba8qWKe1_1(.din(G2897),.dout(w_dff_B_Sba8qWKe1_1),.clk(gclk));
	jdff dff_B_4zqwHMcn3_1(.din(w_dff_B_Sba8qWKe1_1),.dout(w_dff_B_4zqwHMcn3_1),.clk(gclk));
	jdff dff_B_89NlKiQx0_1(.din(w_dff_B_4zqwHMcn3_1),.dout(w_dff_B_89NlKiQx0_1),.clk(gclk));
	jdff dff_A_Kz26MWjc3_0(.dout(w_n1184_0[0]),.din(w_dff_A_Kz26MWjc3_0),.clk(gclk));
	jdff dff_A_1pFUqW7z5_0(.dout(w_dff_A_Kz26MWjc3_0),.din(w_dff_A_1pFUqW7z5_0),.clk(gclk));
	jdff dff_A_ynV1tQbq2_0(.dout(w_dff_A_1pFUqW7z5_0),.din(w_dff_A_ynV1tQbq2_0),.clk(gclk));
	jdff dff_A_2p23fOaE8_0(.dout(w_dff_A_ynV1tQbq2_0),.din(w_dff_A_2p23fOaE8_0),.clk(gclk));
	jdff dff_A_Ddh77EIo3_0(.dout(w_dff_A_2p23fOaE8_0),.din(w_dff_A_Ddh77EIo3_0),.clk(gclk));
	jdff dff_A_uwHyYCaN4_0(.dout(w_dff_A_Ddh77EIo3_0),.din(w_dff_A_uwHyYCaN4_0),.clk(gclk));
	jdff dff_A_1TDUvT3S2_0(.dout(w_dff_A_uwHyYCaN4_0),.din(w_dff_A_1TDUvT3S2_0),.clk(gclk));
	jdff dff_A_qccnRTgA4_0(.dout(w_dff_A_1TDUvT3S2_0),.din(w_dff_A_qccnRTgA4_0),.clk(gclk));
	jdff dff_A_jFumDGFP9_0(.dout(w_dff_A_qccnRTgA4_0),.din(w_dff_A_jFumDGFP9_0),.clk(gclk));
	jdff dff_A_DQgbQ5ou2_0(.dout(w_dff_A_jFumDGFP9_0),.din(w_dff_A_DQgbQ5ou2_0),.clk(gclk));
	jdff dff_A_HGepiMnx9_0(.dout(w_dff_A_DQgbQ5ou2_0),.din(w_dff_A_HGepiMnx9_0),.clk(gclk));
	jdff dff_A_Va2RIp0d2_0(.dout(w_dff_A_HGepiMnx9_0),.din(w_dff_A_Va2RIp0d2_0),.clk(gclk));
	jdff dff_A_ZSVgJwjz6_0(.dout(w_dff_A_Va2RIp0d2_0),.din(w_dff_A_ZSVgJwjz6_0),.clk(gclk));
	jdff dff_A_mSp6CN364_0(.dout(w_dff_A_ZSVgJwjz6_0),.din(w_dff_A_mSp6CN364_0),.clk(gclk));
	jdff dff_A_4n7xRdXz6_0(.dout(w_dff_A_mSp6CN364_0),.din(w_dff_A_4n7xRdXz6_0),.clk(gclk));
	jdff dff_A_Hy90Dgah0_0(.dout(w_dff_A_4n7xRdXz6_0),.din(w_dff_A_Hy90Dgah0_0),.clk(gclk));
	jdff dff_A_2rnEDkGI8_0(.dout(w_dff_A_Hy90Dgah0_0),.din(w_dff_A_2rnEDkGI8_0),.clk(gclk));
	jdff dff_A_QzfuWymG6_0(.dout(w_dff_A_2rnEDkGI8_0),.din(w_dff_A_QzfuWymG6_0),.clk(gclk));
	jdff dff_A_0QdGZfhF6_0(.dout(w_dff_A_QzfuWymG6_0),.din(w_dff_A_0QdGZfhF6_0),.clk(gclk));
	jdff dff_A_8u3wyKNW2_0(.dout(w_dff_A_0QdGZfhF6_0),.din(w_dff_A_8u3wyKNW2_0),.clk(gclk));
	jdff dff_A_TTIOfwLJ6_0(.dout(w_dff_A_8u3wyKNW2_0),.din(w_dff_A_TTIOfwLJ6_0),.clk(gclk));
	jdff dff_A_42VEkzUd0_0(.dout(w_dff_A_TTIOfwLJ6_0),.din(w_dff_A_42VEkzUd0_0),.clk(gclk));
	jdff dff_A_wmnia9FE7_0(.dout(w_dff_A_42VEkzUd0_0),.din(w_dff_A_wmnia9FE7_0),.clk(gclk));
	jdff dff_A_CT01YOIy2_0(.dout(w_dff_A_wmnia9FE7_0),.din(w_dff_A_CT01YOIy2_0),.clk(gclk));
	jdff dff_A_pm5yIr7C7_1(.dout(w_n1175_0[1]),.din(w_dff_A_pm5yIr7C7_1),.clk(gclk));
	jdff dff_A_wZnauLqZ3_1(.dout(w_dff_A_pm5yIr7C7_1),.din(w_dff_A_wZnauLqZ3_1),.clk(gclk));
	jdff dff_A_b2x55jkc4_1(.dout(w_dff_A_wZnauLqZ3_1),.din(w_dff_A_b2x55jkc4_1),.clk(gclk));
	jdff dff_A_8FfXxIw29_1(.dout(w_dff_A_b2x55jkc4_1),.din(w_dff_A_8FfXxIw29_1),.clk(gclk));
	jdff dff_A_FDRDn6rK2_1(.dout(w_dff_A_8FfXxIw29_1),.din(w_dff_A_FDRDn6rK2_1),.clk(gclk));
	jdff dff_A_oR8cAYML1_1(.dout(w_dff_A_FDRDn6rK2_1),.din(w_dff_A_oR8cAYML1_1),.clk(gclk));
	jdff dff_A_hG1efiug5_1(.dout(w_dff_A_oR8cAYML1_1),.din(w_dff_A_hG1efiug5_1),.clk(gclk));
	jdff dff_A_gQjEEydM9_1(.dout(w_dff_A_hG1efiug5_1),.din(w_dff_A_gQjEEydM9_1),.clk(gclk));
	jdff dff_A_HHybKUxy7_1(.dout(w_dff_A_gQjEEydM9_1),.din(w_dff_A_HHybKUxy7_1),.clk(gclk));
	jdff dff_A_QXJHZhwo8_1(.dout(w_dff_A_HHybKUxy7_1),.din(w_dff_A_QXJHZhwo8_1),.clk(gclk));
	jdff dff_A_pFKJmAwX6_1(.dout(w_dff_A_QXJHZhwo8_1),.din(w_dff_A_pFKJmAwX6_1),.clk(gclk));
	jdff dff_A_9a8RfQD82_1(.dout(w_dff_A_pFKJmAwX6_1),.din(w_dff_A_9a8RfQD82_1),.clk(gclk));
	jdff dff_A_d3DqCKDa1_1(.dout(w_dff_A_9a8RfQD82_1),.din(w_dff_A_d3DqCKDa1_1),.clk(gclk));
	jdff dff_A_8snGbMCi7_1(.dout(w_dff_A_d3DqCKDa1_1),.din(w_dff_A_8snGbMCi7_1),.clk(gclk));
	jdff dff_A_1P8R3ZrU3_1(.dout(w_dff_A_8snGbMCi7_1),.din(w_dff_A_1P8R3ZrU3_1),.clk(gclk));
	jdff dff_A_0pCg8Ewb9_1(.dout(w_dff_A_1P8R3ZrU3_1),.din(w_dff_A_0pCg8Ewb9_1),.clk(gclk));
	jdff dff_A_45atGmSj6_1(.dout(w_dff_A_0pCg8Ewb9_1),.din(w_dff_A_45atGmSj6_1),.clk(gclk));
	jdff dff_A_u41i3XLP8_1(.dout(w_dff_A_45atGmSj6_1),.din(w_dff_A_u41i3XLP8_1),.clk(gclk));
	jdff dff_A_2upM7GSy5_1(.dout(w_dff_A_u41i3XLP8_1),.din(w_dff_A_2upM7GSy5_1),.clk(gclk));
	jdff dff_A_At8SYZXR9_1(.dout(w_dff_A_2upM7GSy5_1),.din(w_dff_A_At8SYZXR9_1),.clk(gclk));
	jdff dff_A_3acnhz7g5_1(.dout(w_dff_A_At8SYZXR9_1),.din(w_dff_A_3acnhz7g5_1),.clk(gclk));
	jdff dff_A_tHSp7MYp2_1(.dout(w_dff_A_3acnhz7g5_1),.din(w_dff_A_tHSp7MYp2_1),.clk(gclk));
	jdff dff_A_53yDP0x22_1(.dout(w_dff_A_tHSp7MYp2_1),.din(w_dff_A_53yDP0x22_1),.clk(gclk));
	jdff dff_A_8p9Ep5ph6_1(.dout(w_dff_A_53yDP0x22_1),.din(w_dff_A_8p9Ep5ph6_1),.clk(gclk));
	jdff dff_A_9rvIgHbL5_1(.dout(w_dff_A_8p9Ep5ph6_1),.din(w_dff_A_9rvIgHbL5_1),.clk(gclk));
	jdff dff_A_kY51oWpU0_0(.dout(w_n1187_0[0]),.din(w_dff_A_kY51oWpU0_0),.clk(gclk));
	jdff dff_B_HqIxwYqi2_1(.din(n1060),.dout(w_dff_B_HqIxwYqi2_1),.clk(gclk));
	jdff dff_B_3QW2tG859_0(.din(n1112),.dout(w_dff_B_3QW2tG859_0),.clk(gclk));
	jdff dff_B_O3ot9kj41_0(.din(w_dff_B_3QW2tG859_0),.dout(w_dff_B_O3ot9kj41_0),.clk(gclk));
	jdff dff_B_03xtniDy3_0(.din(w_dff_B_O3ot9kj41_0),.dout(w_dff_B_03xtniDy3_0),.clk(gclk));
	jdff dff_B_y9O1gk6A7_0(.din(w_dff_B_03xtniDy3_0),.dout(w_dff_B_y9O1gk6A7_0),.clk(gclk));
	jdff dff_B_yPoaqPFV1_0(.din(w_dff_B_y9O1gk6A7_0),.dout(w_dff_B_yPoaqPFV1_0),.clk(gclk));
	jdff dff_B_KqbWPMAA7_0(.din(w_dff_B_yPoaqPFV1_0),.dout(w_dff_B_KqbWPMAA7_0),.clk(gclk));
	jdff dff_B_1c3CAWR25_0(.din(n1111),.dout(w_dff_B_1c3CAWR25_0),.clk(gclk));
	jdff dff_B_w0GE4BjP7_0(.din(w_dff_B_1c3CAWR25_0),.dout(w_dff_B_w0GE4BjP7_0),.clk(gclk));
	jdff dff_B_0r2lgX6Z4_0(.din(n1110),.dout(w_dff_B_0r2lgX6Z4_0),.clk(gclk));
	jdff dff_B_DuAUmMZp2_0(.din(w_dff_B_0r2lgX6Z4_0),.dout(w_dff_B_DuAUmMZp2_0),.clk(gclk));
	jdff dff_B_HxY5XDOG6_0(.din(w_dff_B_DuAUmMZp2_0),.dout(w_dff_B_HxY5XDOG6_0),.clk(gclk));
	jdff dff_B_XqlUH8W71_0(.din(w_dff_B_HxY5XDOG6_0),.dout(w_dff_B_XqlUH8W71_0),.clk(gclk));
	jdff dff_B_zWQ86AaD6_0(.din(w_dff_B_XqlUH8W71_0),.dout(w_dff_B_zWQ86AaD6_0),.clk(gclk));
	jdff dff_B_CxBiZ04u6_0(.din(n1109),.dout(w_dff_B_CxBiZ04u6_0),.clk(gclk));
	jdff dff_B_fapM1V6I5_0(.din(w_dff_B_CxBiZ04u6_0),.dout(w_dff_B_fapM1V6I5_0),.clk(gclk));
	jdff dff_B_0HFPlUPS2_1(.din(n1066),.dout(w_dff_B_0HFPlUPS2_1),.clk(gclk));
	jdff dff_B_qyrcYnYh3_1(.din(w_dff_B_0HFPlUPS2_1),.dout(w_dff_B_qyrcYnYh3_1),.clk(gclk));
	jdff dff_B_tA2cNRR86_1(.din(w_dff_B_qyrcYnYh3_1),.dout(w_dff_B_tA2cNRR86_1),.clk(gclk));
	jdff dff_B_jfKWCVpc4_1(.din(w_dff_B_tA2cNRR86_1),.dout(w_dff_B_jfKWCVpc4_1),.clk(gclk));
	jdff dff_B_OAVFaoik4_1(.din(w_dff_B_jfKWCVpc4_1),.dout(w_dff_B_OAVFaoik4_1),.clk(gclk));
	jdff dff_B_3SVCqB2k5_1(.din(w_dff_B_OAVFaoik4_1),.dout(w_dff_B_3SVCqB2k5_1),.clk(gclk));
	jdff dff_B_zSzYDKI31_1(.din(w_dff_B_3SVCqB2k5_1),.dout(w_dff_B_zSzYDKI31_1),.clk(gclk));
	jdff dff_B_cvIotsGl6_1(.din(w_dff_B_zSzYDKI31_1),.dout(w_dff_B_cvIotsGl6_1),.clk(gclk));
	jdff dff_B_jkOunhVU9_1(.din(n1086),.dout(w_dff_B_jkOunhVU9_1),.clk(gclk));
	jdff dff_B_rbq2gHyU0_0(.din(n1105),.dout(w_dff_B_rbq2gHyU0_0),.clk(gclk));
	jdff dff_B_cPSoNOer7_0(.din(w_dff_B_rbq2gHyU0_0),.dout(w_dff_B_cPSoNOer7_0),.clk(gclk));
	jdff dff_B_G3VsxjGG6_0(.din(w_dff_B_cPSoNOer7_0),.dout(w_dff_B_G3VsxjGG6_0),.clk(gclk));
	jdff dff_B_KrTOm0AB8_0(.din(w_dff_B_G3VsxjGG6_0),.dout(w_dff_B_KrTOm0AB8_0),.clk(gclk));
	jdff dff_B_3o3G4KE37_0(.din(w_dff_B_KrTOm0AB8_0),.dout(w_dff_B_3o3G4KE37_0),.clk(gclk));
	jdff dff_B_gwqg9ZZ57_0(.din(w_dff_B_3o3G4KE37_0),.dout(w_dff_B_gwqg9ZZ57_0),.clk(gclk));
	jdff dff_B_LUT0e8DE8_0(.din(w_dff_B_gwqg9ZZ57_0),.dout(w_dff_B_LUT0e8DE8_0),.clk(gclk));
	jdff dff_B_9yTnoITB3_0(.din(w_dff_B_LUT0e8DE8_0),.dout(w_dff_B_9yTnoITB3_0),.clk(gclk));
	jdff dff_B_tpz87DSL5_1(.din(n1092),.dout(w_dff_B_tpz87DSL5_1),.clk(gclk));
	jdff dff_B_cLwlpkND2_1(.din(n1096),.dout(w_dff_B_cLwlpkND2_1),.clk(gclk));
	jdff dff_B_4u4Xii5w3_1(.din(w_dff_B_cLwlpkND2_1),.dout(w_dff_B_4u4Xii5w3_1),.clk(gclk));
	jdff dff_B_eukirPuF1_0(.din(n1099),.dout(w_dff_B_eukirPuF1_0),.clk(gclk));
	jdff dff_B_N2TiApL38_0(.din(n1095),.dout(w_dff_B_N2TiApL38_0),.clk(gclk));
	jdff dff_B_5vmXC67r0_0(.din(w_dff_B_N2TiApL38_0),.dout(w_dff_B_5vmXC67r0_0),.clk(gclk));
	jdff dff_B_GlwAPsGr3_0(.din(w_dff_B_5vmXC67r0_0),.dout(w_dff_B_GlwAPsGr3_0),.clk(gclk));
	jdff dff_B_UpLf7Cvj0_1(.din(n1087),.dout(w_dff_B_UpLf7Cvj0_1),.clk(gclk));
	jdff dff_B_N3LKBBhK5_1(.din(w_dff_B_UpLf7Cvj0_1),.dout(w_dff_B_N3LKBBhK5_1),.clk(gclk));
	jdff dff_B_SqTZABBO3_0(.din(n1089),.dout(w_dff_B_SqTZABBO3_0),.clk(gclk));
	jdff dff_B_geNj874Y9_1(.din(n1072),.dout(w_dff_B_geNj874Y9_1),.clk(gclk));
	jdff dff_B_yVxRmE8s9_1(.din(w_dff_B_geNj874Y9_1),.dout(w_dff_B_yVxRmE8s9_1),.clk(gclk));
	jdff dff_B_lDAau8753_1(.din(n1076),.dout(w_dff_B_lDAau8753_1),.clk(gclk));
	jdff dff_B_SGJTEFsZ7_1(.din(G124),.dout(w_dff_B_SGJTEFsZ7_1),.clk(gclk));
	jdff dff_B_c4nG2qid7_1(.din(w_dff_B_SGJTEFsZ7_1),.dout(w_dff_B_c4nG2qid7_1),.clk(gclk));
	jdff dff_B_nawDsiCY0_1(.din(w_dff_B_c4nG2qid7_1),.dout(w_dff_B_nawDsiCY0_1),.clk(gclk));
	jdff dff_B_wxIQ6v6t5_1(.din(w_dff_B_nawDsiCY0_1),.dout(w_dff_B_wxIQ6v6t5_1),.clk(gclk));
	jdff dff_B_sBac9MlJ7_1(.din(n1077),.dout(w_dff_B_sBac9MlJ7_1),.clk(gclk));
	jdff dff_B_wflMoR4i4_0(.din(n1075),.dout(w_dff_B_wflMoR4i4_0),.clk(gclk));
	jdff dff_B_tJBu7D9I1_0(.din(w_dff_B_wflMoR4i4_0),.dout(w_dff_B_tJBu7D9I1_0),.clk(gclk));
	jdff dff_B_qtNdDxOv6_0(.din(w_dff_B_tJBu7D9I1_0),.dout(w_dff_B_qtNdDxOv6_0),.clk(gclk));
	jdff dff_B_MtutydP07_0(.din(w_dff_B_qtNdDxOv6_0),.dout(w_dff_B_MtutydP07_0),.clk(gclk));
	jdff dff_B_ZfoTuBf89_1(.din(n1067),.dout(w_dff_B_ZfoTuBf89_1),.clk(gclk));
	jdff dff_B_MNVBHVb13_1(.din(n1061),.dout(w_dff_B_MNVBHVb13_1),.clk(gclk));
	jdff dff_B_QdTlWOPy6_1(.din(n1051),.dout(w_dff_B_QdTlWOPy6_1),.clk(gclk));
	jdff dff_B_fq5VyQy93_1(.din(w_dff_B_QdTlWOPy6_1),.dout(w_dff_B_fq5VyQy93_1),.clk(gclk));
	jdff dff_B_UR8JTR1B3_1(.din(w_dff_B_fq5VyQy93_1),.dout(w_dff_B_UR8JTR1B3_1),.clk(gclk));
	jdff dff_A_ouZz7z5y9_1(.dout(w_n1057_0[1]),.din(w_dff_A_ouZz7z5y9_1),.clk(gclk));
	jdff dff_A_LEONILnR6_1(.dout(w_dff_A_ouZz7z5y9_1),.din(w_dff_A_LEONILnR6_1),.clk(gclk));
	jdff dff_A_iGsM9aDg2_1(.dout(w_dff_A_LEONILnR6_1),.din(w_dff_A_iGsM9aDg2_1),.clk(gclk));
	jdff dff_A_Jc0GopvY0_1(.dout(w_dff_A_iGsM9aDg2_1),.din(w_dff_A_Jc0GopvY0_1),.clk(gclk));
	jdff dff_A_N46omXvs3_1(.dout(w_dff_A_Jc0GopvY0_1),.din(w_dff_A_N46omXvs3_1),.clk(gclk));
	jdff dff_A_Ci7AUCfM4_0(.dout(w_n1052_0[0]),.din(w_dff_A_Ci7AUCfM4_0),.clk(gclk));
	jdff dff_B_M7G7dGwZ6_1(.din(n753),.dout(w_dff_B_M7G7dGwZ6_1),.clk(gclk));
	jdff dff_B_Z2wHRDtU8_1(.din(w_dff_B_M7G7dGwZ6_1),.dout(w_dff_B_Z2wHRDtU8_1),.clk(gclk));
	jdff dff_B_Mkgb4XIy6_1(.din(w_dff_B_Z2wHRDtU8_1),.dout(w_dff_B_Mkgb4XIy6_1),.clk(gclk));
	jdff dff_B_ggWbuOSW4_1(.din(w_dff_B_Mkgb4XIy6_1),.dout(w_dff_B_ggWbuOSW4_1),.clk(gclk));
	jdff dff_B_PJlIltPn0_1(.din(w_dff_B_ggWbuOSW4_1),.dout(w_dff_B_PJlIltPn0_1),.clk(gclk));
	jdff dff_B_2wUF6utT3_1(.din(w_dff_B_PJlIltPn0_1),.dout(w_dff_B_2wUF6utT3_1),.clk(gclk));
	jdff dff_A_kOmwN3a39_1(.dout(w_n758_1[1]),.din(w_dff_A_kOmwN3a39_1),.clk(gclk));
	jdff dff_A_HvaXIMe72_1(.dout(w_dff_A_kOmwN3a39_1),.din(w_dff_A_HvaXIMe72_1),.clk(gclk));
	jdff dff_A_Xh1K58Al4_1(.dout(w_dff_A_HvaXIMe72_1),.din(w_dff_A_Xh1K58Al4_1),.clk(gclk));
	jdff dff_B_BkXH2J6l7_0(.din(n752),.dout(w_dff_B_BkXH2J6l7_0),.clk(gclk));
	jdff dff_B_yH6i9vbF7_0(.din(w_dff_B_BkXH2J6l7_0),.dout(w_dff_B_yH6i9vbF7_0),.clk(gclk));
	jdff dff_B_RLfVDbH87_0(.din(w_dff_B_yH6i9vbF7_0),.dout(w_dff_B_RLfVDbH87_0),.clk(gclk));
	jdff dff_B_fmOTz5GE4_0(.din(w_dff_B_RLfVDbH87_0),.dout(w_dff_B_fmOTz5GE4_0),.clk(gclk));
	jdff dff_B_Z5qrbyLp9_0(.din(w_dff_B_fmOTz5GE4_0),.dout(w_dff_B_Z5qrbyLp9_0),.clk(gclk));
	jdff dff_B_QhpdVcFt4_0(.din(w_dff_B_Z5qrbyLp9_0),.dout(w_dff_B_QhpdVcFt4_0),.clk(gclk));
	jdff dff_B_rPYqRfFP4_0(.din(w_dff_B_QhpdVcFt4_0),.dout(w_dff_B_rPYqRfFP4_0),.clk(gclk));
	jdff dff_B_HpupBuZ24_0(.din(w_dff_B_rPYqRfFP4_0),.dout(w_dff_B_HpupBuZ24_0),.clk(gclk));
	jdff dff_A_VoEFyJdg8_0(.dout(w_n1049_0[0]),.din(w_dff_A_VoEFyJdg8_0),.clk(gclk));
	jdff dff_A_be0PVgZO0_0(.dout(w_dff_A_VoEFyJdg8_0),.din(w_dff_A_be0PVgZO0_0),.clk(gclk));
	jdff dff_A_X0rfnNi28_1(.dout(w_n1049_0[1]),.din(w_dff_A_X0rfnNi28_1),.clk(gclk));
	jdff dff_A_RStRHZ5r4_1(.dout(w_dff_A_X0rfnNi28_1),.din(w_dff_A_RStRHZ5r4_1),.clk(gclk));
	jdff dff_B_WRO4cqmB1_0(.din(n1048),.dout(w_dff_B_WRO4cqmB1_0),.clk(gclk));
	jdff dff_B_NZiGFut64_0(.din(n1047),.dout(w_dff_B_NZiGFut64_0),.clk(gclk));
	jdff dff_B_CD8o9nVP1_0(.din(n1045),.dout(w_dff_B_CD8o9nVP1_0),.clk(gclk));
	jdff dff_B_r1dpAwhO4_0(.din(w_dff_B_CD8o9nVP1_0),.dout(w_dff_B_r1dpAwhO4_0),.clk(gclk));
	jdff dff_B_dlwqYE0v5_0(.din(w_dff_B_r1dpAwhO4_0),.dout(w_dff_B_dlwqYE0v5_0),.clk(gclk));
	jdff dff_B_4gFb7LAe8_0(.din(w_dff_B_dlwqYE0v5_0),.dout(w_dff_B_4gFb7LAe8_0),.clk(gclk));
	jdff dff_B_rqk3hDLC2_0(.din(w_dff_B_4gFb7LAe8_0),.dout(w_dff_B_rqk3hDLC2_0),.clk(gclk));
	jdff dff_B_AJAqmFDh4_0(.din(n1044),.dout(w_dff_B_AJAqmFDh4_0),.clk(gclk));
	jdff dff_B_QS0ZtmA05_0(.din(w_dff_B_AJAqmFDh4_0),.dout(w_dff_B_QS0ZtmA05_0),.clk(gclk));
	jdff dff_B_s0mZ4UlJ2_0(.din(n1042),.dout(w_dff_B_s0mZ4UlJ2_0),.clk(gclk));
	jdff dff_B_1ETCG16F7_0(.din(w_dff_B_s0mZ4UlJ2_0),.dout(w_dff_B_1ETCG16F7_0),.clk(gclk));
	jdff dff_B_CflVqS060_1(.din(n1030),.dout(w_dff_B_CflVqS060_1),.clk(gclk));
	jdff dff_B_0Sh2KuhN6_1(.din(n1032),.dout(w_dff_B_0Sh2KuhN6_1),.clk(gclk));
	jdff dff_B_IdX0IT347_1(.din(w_dff_B_0Sh2KuhN6_1),.dout(w_dff_B_IdX0IT347_1),.clk(gclk));
	jdff dff_B_qWSCPjmn4_1(.din(n1035),.dout(w_dff_B_qWSCPjmn4_1),.clk(gclk));
	jdff dff_B_iqyfaPSa7_1(.din(n1027),.dout(w_dff_B_iqyfaPSa7_1),.clk(gclk));
	jdff dff_B_1Bg5NWFk1_0(.din(n1028),.dout(w_dff_B_1Bg5NWFk1_0),.clk(gclk));
	jdff dff_B_DMifZ2951_1(.din(n1015),.dout(w_dff_B_DMifZ2951_1),.clk(gclk));
	jdff dff_B_R4fIqzS48_1(.din(n1017),.dout(w_dff_B_R4fIqzS48_1),.clk(gclk));
	jdff dff_B_t4O3bn2m0_1(.din(n1020),.dout(w_dff_B_t4O3bn2m0_1),.clk(gclk));
	jdff dff_B_pMOYEzSd0_1(.din(n1021),.dout(w_dff_B_pMOYEzSd0_1),.clk(gclk));
	jdff dff_B_H4wbGmLC0_1(.din(n1011),.dout(w_dff_B_H4wbGmLC0_1),.clk(gclk));
	jdff dff_B_ECYdSkgf0_0(.din(n1013),.dout(w_dff_B_ECYdSkgf0_0),.clk(gclk));
	jdff dff_A_xryQdEie7_1(.dout(w_G125_0[1]),.din(w_dff_A_xryQdEie7_1),.clk(gclk));
	jdff dff_B_GRyt55l36_2(.din(G125),.dout(w_dff_B_GRyt55l36_2),.clk(gclk));
	jdff dff_B_uFvxpkhR8_2(.din(w_dff_B_GRyt55l36_2),.dout(w_dff_B_uFvxpkhR8_2),.clk(gclk));
	jdff dff_B_GGlOXZyL8_2(.din(w_dff_B_uFvxpkhR8_2),.dout(w_dff_B_GGlOXZyL8_2),.clk(gclk));
	jdff dff_A_gsJdNsID4_1(.dout(w_n990_0[1]),.din(w_dff_A_gsJdNsID4_1),.clk(gclk));
	jdff dff_A_hlvTrcX62_1(.dout(w_dff_A_gsJdNsID4_1),.din(w_dff_A_hlvTrcX62_1),.clk(gclk));
	jdff dff_A_reohEdbc8_0(.dout(w_n758_0[0]),.din(w_dff_A_reohEdbc8_0),.clk(gclk));
	jdff dff_A_HgkOWHrE4_1(.dout(w_n758_0[1]),.din(w_dff_A_HgkOWHrE4_1),.clk(gclk));
	jdff dff_A_XItf8W6e8_1(.dout(w_dff_A_HgkOWHrE4_1),.din(w_dff_A_XItf8W6e8_1),.clk(gclk));
	jdff dff_A_0wblCObB8_1(.dout(w_dff_A_XItf8W6e8_1),.din(w_dff_A_0wblCObB8_1),.clk(gclk));
	jdff dff_A_v1fpQzmh4_0(.dout(w_n754_0[0]),.din(w_dff_A_v1fpQzmh4_0),.clk(gclk));
	jdff dff_B_6QtczEZz2_0(.din(n768),.dout(w_dff_B_6QtczEZz2_0),.clk(gclk));
	jdff dff_B_MA6gwNRH6_0(.din(n767),.dout(w_dff_B_MA6gwNRH6_0),.clk(gclk));
	jdff dff_B_PjZIbyet8_0(.din(w_dff_B_MA6gwNRH6_0),.dout(w_dff_B_PjZIbyet8_0),.clk(gclk));
	jdff dff_B_CPQM883m4_0(.din(w_dff_B_PjZIbyet8_0),.dout(w_dff_B_CPQM883m4_0),.clk(gclk));
	jdff dff_A_MuEtCERx8_2(.dout(w_n764_1[2]),.din(w_dff_A_MuEtCERx8_2),.clk(gclk));
	jdff dff_A_vEisUAsu2_2(.dout(w_dff_A_MuEtCERx8_2),.din(w_dff_A_vEisUAsu2_2),.clk(gclk));
	jdff dff_A_CtVzTCe36_1(.dout(w_n1183_0[1]),.din(w_dff_A_CtVzTCe36_1),.clk(gclk));
	jdff dff_B_nO6CwKfE5_1(.din(n1179),.dout(w_dff_B_nO6CwKfE5_1),.clk(gclk));
	jdff dff_B_jlWztoAt0_1(.din(w_dff_B_nO6CwKfE5_1),.dout(w_dff_B_jlWztoAt0_1),.clk(gclk));
	jdff dff_B_Ltzkq9aT6_1(.din(n1180),.dout(w_dff_B_Ltzkq9aT6_1),.clk(gclk));
	jdff dff_B_BzDzznrh5_1(.din(w_dff_B_Ltzkq9aT6_1),.dout(w_dff_B_BzDzznrh5_1),.clk(gclk));
	jdff dff_B_iBNBekbK7_1(.din(w_dff_B_BzDzznrh5_1),.dout(w_dff_B_iBNBekbK7_1),.clk(gclk));
	jdff dff_A_BCacFK5p1_0(.dout(w_n988_0[0]),.din(w_dff_A_BCacFK5p1_0),.clk(gclk));
	jdff dff_A_aXqDb7Dy9_0(.dout(w_dff_A_BCacFK5p1_0),.din(w_dff_A_aXqDb7Dy9_0),.clk(gclk));
	jdff dff_A_kO1rFbt35_1(.dout(w_n988_0[1]),.din(w_dff_A_kO1rFbt35_1),.clk(gclk));
	jdff dff_B_HbqcTied8_0(.din(n986),.dout(w_dff_B_HbqcTied8_0),.clk(gclk));
	jdff dff_B_Hlt852rt5_0(.din(w_dff_B_HbqcTied8_0),.dout(w_dff_B_Hlt852rt5_0),.clk(gclk));
	jdff dff_B_v9TyYiHT8_0(.din(n984),.dout(w_dff_B_v9TyYiHT8_0),.clk(gclk));
	jdff dff_B_QigrX8J72_0(.din(w_dff_B_v9TyYiHT8_0),.dout(w_dff_B_QigrX8J72_0),.clk(gclk));
	jdff dff_B_sFDQ1TAz3_0(.din(w_dff_B_QigrX8J72_0),.dout(w_dff_B_sFDQ1TAz3_0),.clk(gclk));
	jdff dff_B_5FHqcI0s9_0(.din(w_dff_B_sFDQ1TAz3_0),.dout(w_dff_B_5FHqcI0s9_0),.clk(gclk));
	jdff dff_B_5DfRk7g22_0(.din(n983),.dout(w_dff_B_5DfRk7g22_0),.clk(gclk));
	jdff dff_B_bd4qKzwn7_0(.din(w_dff_B_5DfRk7g22_0),.dout(w_dff_B_bd4qKzwn7_0),.clk(gclk));
	jdff dff_B_6cZt0YIi7_1(.din(n979),.dout(w_dff_B_6cZt0YIi7_1),.clk(gclk));
	jdff dff_B_C05oqTQr5_1(.din(w_dff_B_6cZt0YIi7_1),.dout(w_dff_B_C05oqTQr5_1),.clk(gclk));
	jdff dff_B_tybHPE6C0_0(.din(n980),.dout(w_dff_B_tybHPE6C0_0),.clk(gclk));
	jdff dff_A_7QBH7DgZ4_2(.dout(w_G97_2[2]),.din(w_dff_A_7QBH7DgZ4_2),.clk(gclk));
	jdff dff_B_TASpClio3_2(.din(n144),.dout(w_dff_B_TASpClio3_2),.clk(gclk));
	jdff dff_B_bujkl3Rf1_1(.din(n142),.dout(w_dff_B_bujkl3Rf1_1),.clk(gclk));
	jdff dff_B_woEMQmxf1_1(.din(n966),.dout(w_dff_B_woEMQmxf1_1),.clk(gclk));
	jdff dff_B_7ZSJceom5_1(.din(n968),.dout(w_dff_B_7ZSJceom5_1),.clk(gclk));
	jdff dff_B_nXJrMS4Q5_1(.din(n971),.dout(w_dff_B_nXJrMS4Q5_1),.clk(gclk));
	jdff dff_B_3vBlmhip4_0(.din(n972),.dout(w_dff_B_3vBlmhip4_0),.clk(gclk));
	jdff dff_A_PugzPvyA2_0(.dout(w_G143_1[0]),.din(w_dff_A_PugzPvyA2_0),.clk(gclk));
	jdff dff_A_sFVymup87_2(.dout(w_G143_1[2]),.din(w_dff_A_sFVymup87_2),.clk(gclk));
	jdff dff_A_goNGes1R7_1(.dout(w_G33_4[1]),.din(w_dff_A_goNGes1R7_1),.clk(gclk));
	jdff dff_A_nTIZuExK6_1(.dout(w_dff_A_goNGes1R7_1),.din(w_dff_A_nTIZuExK6_1),.clk(gclk));
	jdff dff_A_hMSCEz6U5_1(.dout(w_dff_A_nTIZuExK6_1),.din(w_dff_A_hMSCEz6U5_1),.clk(gclk));
	jdff dff_A_F7LThMu61_1(.dout(w_dff_A_hMSCEz6U5_1),.din(w_dff_A_F7LThMu61_1),.clk(gclk));
	jdff dff_A_xJ1nBBsq8_2(.dout(w_G33_4[2]),.din(w_dff_A_xJ1nBBsq8_2),.clk(gclk));
	jdff dff_A_lbkfI0PV4_2(.dout(w_dff_A_xJ1nBBsq8_2),.din(w_dff_A_lbkfI0PV4_2),.clk(gclk));
	jdff dff_A_ViR2xfxe9_2(.dout(w_dff_A_lbkfI0PV4_2),.din(w_dff_A_ViR2xfxe9_2),.clk(gclk));
	jdff dff_A_U84xEFrr8_2(.dout(w_dff_A_ViR2xfxe9_2),.din(w_dff_A_U84xEFrr8_2),.clk(gclk));
	jdff dff_B_bTXCXE3W2_0(.din(n964),.dout(w_dff_B_bTXCXE3W2_0),.clk(gclk));
	jdff dff_A_0J4OVUoY9_1(.dout(w_n962_0[1]),.din(w_dff_A_0J4OVUoY9_1),.clk(gclk));
	jdff dff_B_ivslArfX2_1(.din(n951),.dout(w_dff_B_ivslArfX2_1),.clk(gclk));
	jdff dff_B_2acrcGUW7_1(.din(n953),.dout(w_dff_B_2acrcGUW7_1),.clk(gclk));
	jdff dff_B_1JNOJRPv9_1(.din(n956),.dout(w_dff_B_1JNOJRPv9_1),.clk(gclk));
	jdff dff_B_4bYsWbFL6_0(.din(n957),.dout(w_dff_B_4bYsWbFL6_0),.clk(gclk));
	jdff dff_B_60i9nVvj7_1(.din(n947),.dout(w_dff_B_60i9nVvj7_1),.clk(gclk));
	jdff dff_B_M0D7D2sP4_0(.din(n949),.dout(w_dff_B_M0D7D2sP4_0),.clk(gclk));
	jdff dff_A_b3zYzCpI2_0(.dout(w_n603_1[0]),.din(w_dff_A_b3zYzCpI2_0),.clk(gclk));
	jdff dff_A_1B2TbiEd3_0(.dout(w_dff_A_b3zYzCpI2_0),.din(w_dff_A_1B2TbiEd3_0),.clk(gclk));
	jdff dff_A_aEkXezqP0_0(.dout(w_dff_A_1B2TbiEd3_0),.din(w_dff_A_aEkXezqP0_0),.clk(gclk));
	jdff dff_B_GkG2VC3M5_1(.din(n850),.dout(w_dff_B_GkG2VC3M5_1),.clk(gclk));
	jdff dff_B_z0hCELaH0_1(.din(w_dff_B_GkG2VC3M5_1),.dout(w_dff_B_z0hCELaH0_1),.clk(gclk));
	jdff dff_B_FH0il0nK3_1(.din(w_dff_B_z0hCELaH0_1),.dout(w_dff_B_FH0il0nK3_1),.clk(gclk));
	jdff dff_B_oHTSJ5C89_1(.din(w_dff_B_FH0il0nK3_1),.dout(w_dff_B_oHTSJ5C89_1),.clk(gclk));
	jdff dff_B_pK2sato87_1(.din(w_dff_B_oHTSJ5C89_1),.dout(w_dff_B_pK2sato87_1),.clk(gclk));
	jdff dff_B_Bt9QAkTd5_1(.din(w_dff_B_pK2sato87_1),.dout(w_dff_B_Bt9QAkTd5_1),.clk(gclk));
	jdff dff_B_jDrwD3dI6_0(.din(n875),.dout(w_dff_B_jDrwD3dI6_0),.clk(gclk));
	jdff dff_B_JUvPulu93_0(.din(w_dff_B_jDrwD3dI6_0),.dout(w_dff_B_JUvPulu93_0),.clk(gclk));
	jdff dff_B_EVI7LtAT4_1(.din(n871),.dout(w_dff_B_EVI7LtAT4_1),.clk(gclk));
	jdff dff_B_1KlVEaGy7_1(.din(n868),.dout(w_dff_B_1KlVEaGy7_1),.clk(gclk));
	jdff dff_B_WMVZfwea1_1(.din(w_dff_B_1KlVEaGy7_1),.dout(w_dff_B_WMVZfwea1_1),.clk(gclk));
	jdff dff_B_csNboiwg8_1(.din(w_dff_B_WMVZfwea1_1),.dout(w_dff_B_csNboiwg8_1),.clk(gclk));
	jdff dff_B_uN3yNqMX3_1(.din(w_dff_B_csNboiwg8_1),.dout(w_dff_B_uN3yNqMX3_1),.clk(gclk));
	jdff dff_B_RgDzYCTb1_1(.din(w_dff_B_uN3yNqMX3_1),.dout(w_dff_B_RgDzYCTb1_1),.clk(gclk));
	jdff dff_A_5MRBFqNf2_1(.dout(w_n861_1[1]),.din(w_dff_A_5MRBFqNf2_1),.clk(gclk));
	jdff dff_A_miPFumjC5_1(.dout(w_dff_A_5MRBFqNf2_1),.din(w_dff_A_miPFumjC5_1),.clk(gclk));
	jdff dff_A_vySj1KXD5_2(.dout(w_n861_0[2]),.din(w_dff_A_vySj1KXD5_2),.clk(gclk));
	jdff dff_A_h8BRsSgY3_2(.dout(w_dff_A_vySj1KXD5_2),.din(w_dff_A_h8BRsSgY3_2),.clk(gclk));
	jdff dff_B_91mPsrla4_0(.din(n860),.dout(w_dff_B_91mPsrla4_0),.clk(gclk));
	jdff dff_B_HZLESQmS3_0(.din(n857),.dout(w_dff_B_HZLESQmS3_0),.clk(gclk));
	jdff dff_B_iiAPVMOV7_0(.din(w_dff_B_HZLESQmS3_0),.dout(w_dff_B_iiAPVMOV7_0),.clk(gclk));
	jdff dff_B_izibPMR73_0(.din(w_dff_B_iiAPVMOV7_0),.dout(w_dff_B_izibPMR73_0),.clk(gclk));
	jdff dff_A_n3ud26WU8_1(.dout(w_n563_0[1]),.din(w_dff_A_n3ud26WU8_1),.clk(gclk));
	jdff dff_A_jYdxiSC18_1(.dout(w_dff_A_n3ud26WU8_1),.din(w_dff_A_jYdxiSC18_1),.clk(gclk));
	jdff dff_A_ejReBi1n1_2(.dout(w_n563_0[2]),.din(w_dff_A_ejReBi1n1_2),.clk(gclk));
	jdff dff_A_OgC83iMD6_2(.dout(w_dff_A_ejReBi1n1_2),.din(w_dff_A_OgC83iMD6_2),.clk(gclk));
	jdff dff_B_XA4MjNtg9_1(.din(n555),.dout(w_dff_B_XA4MjNtg9_1),.clk(gclk));
	jdff dff_B_MFdEChYk2_1(.din(w_dff_B_XA4MjNtg9_1),.dout(w_dff_B_MFdEChYk2_1),.clk(gclk));
	jdff dff_B_BOKcaclG7_1(.din(w_dff_B_MFdEChYk2_1),.dout(w_dff_B_BOKcaclG7_1),.clk(gclk));
	jdff dff_B_5xXmWcjF8_0(.din(n849),.dout(w_dff_B_5xXmWcjF8_0),.clk(gclk));
	jdff dff_B_lMaU6M2E7_0(.din(w_dff_B_5xXmWcjF8_0),.dout(w_dff_B_lMaU6M2E7_0),.clk(gclk));
	jdff dff_B_ZDlQ6QMx7_0(.din(n848),.dout(w_dff_B_ZDlQ6QMx7_0),.clk(gclk));
	jdff dff_B_KGN0Cfxo1_0(.din(w_dff_B_ZDlQ6QMx7_0),.dout(w_dff_B_KGN0Cfxo1_0),.clk(gclk));
	jdff dff_B_Nsxm4RzF0_0(.din(w_dff_B_KGN0Cfxo1_0),.dout(w_dff_B_Nsxm4RzF0_0),.clk(gclk));
	jdff dff_B_4csAsGzu2_0(.din(w_dff_B_Nsxm4RzF0_0),.dout(w_dff_B_4csAsGzu2_0),.clk(gclk));
	jdff dff_B_QDoeX3ui6_1(.din(n844),.dout(w_dff_B_QDoeX3ui6_1),.clk(gclk));
	jdff dff_B_6RDoPbTe0_1(.din(w_dff_B_QDoeX3ui6_1),.dout(w_dff_B_6RDoPbTe0_1),.clk(gclk));
	jdff dff_B_SfLpZ49O7_0(.din(n845),.dout(w_dff_B_SfLpZ49O7_0),.clk(gclk));
	jdff dff_A_yZq3Id2l3_0(.dout(w_n131_0[0]),.din(w_dff_A_yZq3Id2l3_0),.clk(gclk));
	jdff dff_B_3TlZntCp2_1(.din(n129),.dout(w_dff_B_3TlZntCp2_1),.clk(gclk));
	jdff dff_B_iHQo5wAi7_1(.din(n820),.dout(w_dff_B_iHQo5wAi7_1),.clk(gclk));
	jdff dff_B_MPZkSopX3_1(.din(w_dff_B_iHQo5wAi7_1),.dout(w_dff_B_MPZkSopX3_1),.clk(gclk));
	jdff dff_B_jB04fN5o7_1(.din(n828),.dout(w_dff_B_jB04fN5o7_1),.clk(gclk));
	jdff dff_B_pKX3Z6ci2_1(.din(n830),.dout(w_dff_B_pKX3Z6ci2_1),.clk(gclk));
	jdff dff_B_41U9DHKJ6_1(.din(w_dff_B_pKX3Z6ci2_1),.dout(w_dff_B_41U9DHKJ6_1),.clk(gclk));
	jdff dff_B_9KRSL5N54_1(.din(n833),.dout(w_dff_B_9KRSL5N54_1),.clk(gclk));
	jdff dff_B_VokvmHoW1_1(.din(n834),.dout(w_dff_B_VokvmHoW1_1),.clk(gclk));
	jdff dff_B_XDbCX56u3_1(.din(n822),.dout(w_dff_B_XDbCX56u3_1),.clk(gclk));
	jdff dff_B_o7ogLalW2_1(.din(n809),.dout(w_dff_B_o7ogLalW2_1),.clk(gclk));
	jdff dff_B_60dAyajg5_1(.din(n811),.dout(w_dff_B_60dAyajg5_1),.clk(gclk));
	jdff dff_B_aLyvrF5y2_1(.din(n814),.dout(w_dff_B_aLyvrF5y2_1),.clk(gclk));
	jdff dff_B_E3kh8RIO8_1(.din(n815),.dout(w_dff_B_E3kh8RIO8_1),.clk(gclk));
	jdff dff_B_icDZmfxm3_1(.din(n805),.dout(w_dff_B_icDZmfxm3_1),.clk(gclk));
	jdff dff_B_JiIMEmpI1_0(.din(n807),.dout(w_dff_B_JiIMEmpI1_0),.clk(gclk));
	jdff dff_A_CPktjDSG5_2(.dout(w_G107_2[2]),.din(w_dff_A_CPktjDSG5_2),.clk(gclk));
	jdff dff_A_qp1sAGMq6_0(.dout(w_n801_0[0]),.din(w_dff_A_qp1sAGMq6_0),.clk(gclk));
	jdff dff_A_4qe0AaBu3_0(.dout(w_dff_A_qp1sAGMq6_0),.din(w_dff_A_4qe0AaBu3_0),.clk(gclk));
	jdff dff_A_G158mUnH8_0(.dout(w_dff_A_4qe0AaBu3_0),.din(w_dff_A_G158mUnH8_0),.clk(gclk));
	jdff dff_A_LdP0sqej6_0(.dout(w_dff_A_G158mUnH8_0),.din(w_dff_A_LdP0sqej6_0),.clk(gclk));
	jdff dff_B_IhUb9nu18_0(.din(n800),.dout(w_dff_B_IhUb9nu18_0),.clk(gclk));
	jdff dff_B_jj7AxzEY2_0(.din(n798),.dout(w_dff_B_jj7AxzEY2_0),.clk(gclk));
	jdff dff_A_R9T0BBH90_0(.dout(w_n797_0[0]),.din(w_dff_A_R9T0BBH90_0),.clk(gclk));
	jdff dff_B_CaZgp0CW2_0(.din(n936),.dout(w_dff_B_CaZgp0CW2_0),.clk(gclk));
	jdff dff_B_xcyXUC0e7_0(.din(w_dff_B_CaZgp0CW2_0),.dout(w_dff_B_xcyXUC0e7_0),.clk(gclk));
	jdff dff_B_pBuz2pDf9_0(.din(n935),.dout(w_dff_B_pBuz2pDf9_0),.clk(gclk));
	jdff dff_B_SVihhk5e3_0(.din(n934),.dout(w_dff_B_SVihhk5e3_0),.clk(gclk));
	jdff dff_B_anfcVjYq8_0(.din(w_dff_B_SVihhk5e3_0),.dout(w_dff_B_anfcVjYq8_0),.clk(gclk));
	jdff dff_B_7vlzAMVs7_1(.din(n924),.dout(w_dff_B_7vlzAMVs7_1),.clk(gclk));
	jdff dff_B_Wtje1SaE7_1(.din(n925),.dout(w_dff_B_Wtje1SaE7_1),.clk(gclk));
	jdff dff_B_8U9rPPQx0_1(.din(n916),.dout(w_dff_B_8U9rPPQx0_1),.clk(gclk));
	jdff dff_B_7KrCzawj1_1(.din(w_dff_B_8U9rPPQx0_1),.dout(w_dff_B_7KrCzawj1_1),.clk(gclk));
	jdff dff_B_BFovSasJ9_1(.din(n918),.dout(w_dff_B_BFovSasJ9_1),.clk(gclk));
	jdff dff_A_3K811a2e5_1(.dout(w_n73_1[1]),.din(w_dff_A_3K811a2e5_1),.clk(gclk));
	jdff dff_A_oOUnMqgv3_1(.dout(w_n135_0[1]),.din(w_dff_A_oOUnMqgv3_1),.clk(gclk));
	jdff dff_B_vF6pt99o2_1(.din(n133),.dout(w_dff_B_vF6pt99o2_1),.clk(gclk));
	jdff dff_B_WnKyF0ti2_1(.din(n902),.dout(w_dff_B_WnKyF0ti2_1),.clk(gclk));
	jdff dff_B_AyWMX6dN8_1(.din(n904),.dout(w_dff_B_AyWMX6dN8_1),.clk(gclk));
	jdff dff_B_FFFNZjvU1_1(.din(n907),.dout(w_dff_B_FFFNZjvU1_1),.clk(gclk));
	jdff dff_B_gz7dj8DM7_1(.din(n908),.dout(w_dff_B_gz7dj8DM7_1),.clk(gclk));
	jdff dff_A_dueqaJgq7_0(.dout(w_G50_2[0]),.din(w_dff_A_dueqaJgq7_0),.clk(gclk));
	jdff dff_A_OzKVJmt60_1(.dout(w_G68_2[1]),.din(w_dff_A_OzKVJmt60_1),.clk(gclk));
	jdff dff_A_0n0CCISK2_1(.dout(w_dff_A_OzKVJmt60_1),.din(w_dff_A_0n0CCISK2_1),.clk(gclk));
	jdff dff_A_gRyxMBcX9_1(.dout(w_dff_A_0n0CCISK2_1),.din(w_dff_A_gRyxMBcX9_1),.clk(gclk));
	jdff dff_A_wrgjO4ru4_2(.dout(w_G68_2[2]),.din(w_dff_A_wrgjO4ru4_2),.clk(gclk));
	jdff dff_A_BL9huDU75_2(.dout(w_dff_A_wrgjO4ru4_2),.din(w_dff_A_BL9huDU75_2),.clk(gclk));
	jdff dff_A_iqe8B1jB8_2(.dout(w_dff_A_BL9huDU75_2),.din(w_dff_A_iqe8B1jB8_2),.clk(gclk));
	jdff dff_A_64ftG2JB1_2(.dout(w_dff_A_iqe8B1jB8_2),.din(w_dff_A_64ftG2JB1_2),.clk(gclk));
	jdff dff_A_z0DziQVH6_1(.dout(w_G150_2[1]),.din(w_dff_A_z0DziQVH6_1),.clk(gclk));
	jdff dff_B_jijveFSS1_0(.din(n900),.dout(w_dff_B_jijveFSS1_0),.clk(gclk));
	jdff dff_A_lGm10NeH2_0(.dout(w_G58_2[0]),.din(w_dff_A_lGm10NeH2_0),.clk(gclk));
	jdff dff_A_Cfx5oZ4z1_0(.dout(w_dff_A_lGm10NeH2_0),.din(w_dff_A_Cfx5oZ4z1_0),.clk(gclk));
	jdff dff_A_KnaJJwVi3_2(.dout(w_G58_2[2]),.din(w_dff_A_KnaJJwVi3_2),.clk(gclk));
	jdff dff_A_ul9kiYTC7_2(.dout(w_dff_A_KnaJJwVi3_2),.din(w_dff_A_ul9kiYTC7_2),.clk(gclk));
	jdff dff_B_RxDJlPs49_1(.din(n887),.dout(w_dff_B_RxDJlPs49_1),.clk(gclk));
	jdff dff_B_SfGEYDQO1_1(.din(n889),.dout(w_dff_B_SfGEYDQO1_1),.clk(gclk));
	jdff dff_B_imB7NkY34_0(.din(n895),.dout(w_dff_B_imB7NkY34_0),.clk(gclk));
	jdff dff_B_TYKlVe3n2_0(.din(n891),.dout(w_dff_B_TYKlVe3n2_0),.clk(gclk));
	jdff dff_A_P2HetoOa5_1(.dout(w_G116_2[1]),.din(w_dff_A_P2HetoOa5_1),.clk(gclk));
	jdff dff_A_oerN6jKl5_2(.dout(w_G116_2[2]),.din(w_dff_A_oerN6jKl5_2),.clk(gclk));
	jdff dff_B_r4P1rwqF3_1(.din(n883),.dout(w_dff_B_r4P1rwqF3_1),.clk(gclk));
	jdff dff_B_umOvivqc3_0(.din(n885),.dout(w_dff_B_umOvivqc3_0),.clk(gclk));
	jdff dff_A_ySobaZ7d0_0(.dout(w_G283_2[0]),.din(w_dff_A_ySobaZ7d0_0),.clk(gclk));
	jdff dff_A_4xonIQ2c6_1(.dout(w_G283_2[1]),.din(w_dff_A_4xonIQ2c6_1),.clk(gclk));
	jdff dff_A_VOB1MuIG0_1(.dout(w_n564_0[1]),.din(w_dff_A_VOB1MuIG0_1),.clk(gclk));
	jdff dff_B_3YAnUPyw5_1(.din(n878),.dout(w_dff_B_3YAnUPyw5_1),.clk(gclk));
	jdff dff_B_CwgtMlEH9_1(.din(w_dff_B_3YAnUPyw5_1),.dout(w_dff_B_CwgtMlEH9_1),.clk(gclk));
	jdff dff_A_auWLdSP48_0(.dout(w_n589_1[0]),.din(w_dff_A_auWLdSP48_0),.clk(gclk));
	jdff dff_A_MMhFJs1l8_0(.dout(w_dff_A_auWLdSP48_0),.din(w_dff_A_MMhFJs1l8_0),.clk(gclk));
	jdff dff_A_Ci1lgWHE0_0(.dout(w_dff_A_MMhFJs1l8_0),.din(w_dff_A_Ci1lgWHE0_0),.clk(gclk));
	jdff dff_A_NyrFAQ7A8_0(.dout(w_n592_1[0]),.din(w_dff_A_NyrFAQ7A8_0),.clk(gclk));
	jdff dff_A_7zXK7Z0j7_0(.dout(w_dff_A_NyrFAQ7A8_0),.din(w_dff_A_7zXK7Z0j7_0),.clk(gclk));
	jdff dff_A_b1O6bxue3_1(.dout(w_n592_1[1]),.din(w_dff_A_b1O6bxue3_1),.clk(gclk));
	jdff dff_B_QKGI8h3V0_0(.din(n852),.dout(w_dff_B_QKGI8h3V0_0),.clk(gclk));
	jdff dff_B_pKNYMOUG6_0(.din(n560),.dout(w_dff_B_pKNYMOUG6_0),.clk(gclk));
	jdff dff_B_llGLiG5a1_2(.din(n556),.dout(w_dff_B_llGLiG5a1_2),.clk(gclk));
	jdff dff_B_e8e0s9Tw7_2(.din(w_dff_B_llGLiG5a1_2),.dout(w_dff_B_e8e0s9Tw7_2),.clk(gclk));
	jdff dff_A_gNDVYk1S1_0(.dout(w_G396_0[0]),.din(w_dff_A_gNDVYk1S1_0),.clk(gclk));
	jdff dff_A_OexgeZbJ0_0(.dout(w_dff_A_gNDVYk1S1_0),.din(w_dff_A_OexgeZbJ0_0),.clk(gclk));
	jdff dff_A_wHFAAAM29_0(.dout(w_dff_A_OexgeZbJ0_0),.din(w_dff_A_wHFAAAM29_0),.clk(gclk));
	jdff dff_B_r7I87ypp4_0(.din(n687),.dout(w_dff_B_r7I87ypp4_0),.clk(gclk));
	jdff dff_B_XBhVLbD39_0(.din(w_dff_B_r7I87ypp4_0),.dout(w_dff_B_XBhVLbD39_0),.clk(gclk));
	jdff dff_B_scrVZ7927_0(.din(n686),.dout(w_dff_B_scrVZ7927_0),.clk(gclk));
	jdff dff_B_AqESJkoR8_0(.din(w_dff_B_scrVZ7927_0),.dout(w_dff_B_AqESJkoR8_0),.clk(gclk));
	jdff dff_B_T07KtoY26_1(.din(n678),.dout(w_dff_B_T07KtoY26_1),.clk(gclk));
	jdff dff_B_t9fHK07t4_1(.din(n679),.dout(w_dff_B_t9fHK07t4_1),.clk(gclk));
	jdff dff_B_A4QDMoH20_2(.din(n680),.dout(w_dff_B_A4QDMoH20_2),.clk(gclk));
	jdff dff_B_vwMSbg3t9_1(.din(n673),.dout(w_dff_B_vwMSbg3t9_1),.clk(gclk));
	jdff dff_B_z7x30knv6_1(.din(w_dff_B_vwMSbg3t9_1),.dout(w_dff_B_z7x30knv6_1),.clk(gclk));
	jdff dff_B_9Ye4cWSA9_0(.din(n139),.dout(w_dff_B_9Ye4cWSA9_0),.clk(gclk));
	jdff dff_A_twfCMpHp6_1(.dout(w_n672_1[1]),.din(w_dff_A_twfCMpHp6_1),.clk(gclk));
	jdff dff_A_FoTsNkAw5_1(.dout(w_dff_A_twfCMpHp6_1),.din(w_dff_A_FoTsNkAw5_1),.clk(gclk));
	jdff dff_A_jxubB8fU3_1(.dout(w_dff_A_FoTsNkAw5_1),.din(w_dff_A_jxubB8fU3_1),.clk(gclk));
	jdff dff_A_lRwSU2RU9_2(.dout(w_n672_0[2]),.din(w_dff_A_lRwSU2RU9_2),.clk(gclk));
	jdff dff_A_bd3qanCL6_2(.dout(w_dff_A_lRwSU2RU9_2),.din(w_dff_A_bd3qanCL6_2),.clk(gclk));
	jdff dff_A_cwbGpK2Z3_2(.dout(w_dff_A_bd3qanCL6_2),.din(w_dff_A_cwbGpK2Z3_2),.clk(gclk));
	jdff dff_B_82kYTqqJ9_1(.din(n647),.dout(w_dff_B_82kYTqqJ9_1),.clk(gclk));
	jdff dff_B_h10GtyIo3_1(.din(w_dff_B_82kYTqqJ9_1),.dout(w_dff_B_h10GtyIo3_1),.clk(gclk));
	jdff dff_B_EJ1B3EeP0_1(.din(n653),.dout(w_dff_B_EJ1B3EeP0_1),.clk(gclk));
	jdff dff_B_hSFoL9Vx7_1(.din(w_dff_B_EJ1B3EeP0_1),.dout(w_dff_B_hSFoL9Vx7_1),.clk(gclk));
	jdff dff_B_JttXkiGp9_1(.din(n656),.dout(w_dff_B_JttXkiGp9_1),.clk(gclk));
	jdff dff_B_XCGnxZHc1_1(.din(n660),.dout(w_dff_B_XCGnxZHc1_1),.clk(gclk));
	jdff dff_B_hLJtlJJF9_0(.din(n658),.dout(w_dff_B_hLJtlJJF9_0),.clk(gclk));
	jdff dff_B_gkg3k09p5_1(.din(n630),.dout(w_dff_B_gkg3k09p5_1),.clk(gclk));
	jdff dff_B_Gc1DhZXX9_1(.din(n633),.dout(w_dff_B_Gc1DhZXX9_1),.clk(gclk));
	jdff dff_B_ItcZGkKB8_0(.din(n644),.dout(w_dff_B_ItcZGkKB8_0),.clk(gclk));
	jdff dff_A_XwDnaQlt8_0(.dout(w_G317_1[0]),.din(w_dff_A_XwDnaQlt8_0),.clk(gclk));
	jdff dff_B_LMCkRrVG6_3(.din(G317),.dout(w_dff_B_LMCkRrVG6_3),.clk(gclk));
	jdff dff_B_H1HY01fP6_3(.din(w_dff_B_LMCkRrVG6_3),.dout(w_dff_B_H1HY01fP6_3),.clk(gclk));
	jdff dff_B_ZmiO3i2x6_3(.din(w_dff_B_H1HY01fP6_3),.dout(w_dff_B_ZmiO3i2x6_3),.clk(gclk));
	jdff dff_A_v49lq3ym8_0(.dout(w_G326_0[0]),.din(w_dff_A_v49lq3ym8_0),.clk(gclk));
	jdff dff_B_Spb4oRM94_2(.din(G326),.dout(w_dff_B_Spb4oRM94_2),.clk(gclk));
	jdff dff_B_iymQpDhf8_2(.din(w_dff_B_Spb4oRM94_2),.dout(w_dff_B_iymQpDhf8_2),.clk(gclk));
	jdff dff_B_iGSNmT5R3_2(.din(w_dff_B_iymQpDhf8_2),.dout(w_dff_B_iGSNmT5R3_2),.clk(gclk));
	jdff dff_B_nxT6o9XU7_0(.din(n637),.dout(w_dff_B_nxT6o9XU7_0),.clk(gclk));
	jdff dff_B_NKXEqKka3_1(.din(G329),.dout(w_dff_B_NKXEqKka3_1),.clk(gclk));
	jdff dff_B_8uaxFcVp8_1(.din(w_dff_B_NKXEqKka3_1),.dout(w_dff_B_8uaxFcVp8_1),.clk(gclk));
	jdff dff_B_n5lwAc6J4_1(.din(w_dff_B_8uaxFcVp8_1),.dout(w_dff_B_n5lwAc6J4_1),.clk(gclk));
	jdff dff_B_fa6AkwhY3_1(.din(w_dff_B_n5lwAc6J4_1),.dout(w_dff_B_fa6AkwhY3_1),.clk(gclk));
	jdff dff_A_UIxmzBzU1_1(.dout(w_n148_5[1]),.din(w_dff_A_UIxmzBzU1_1),.clk(gclk));
	jdff dff_A_REiphj4s6_1(.dout(w_dff_A_UIxmzBzU1_1),.din(w_dff_A_REiphj4s6_1),.clk(gclk));
	jdff dff_A_Dg7xY4Fv9_1(.dout(w_dff_A_REiphj4s6_1),.din(w_dff_A_Dg7xY4Fv9_1),.clk(gclk));
	jdff dff_A_PuunYYEp3_2(.dout(w_n148_5[2]),.din(w_dff_A_PuunYYEp3_2),.clk(gclk));
	jdff dff_A_qFR6XBNy6_2(.dout(w_dff_A_PuunYYEp3_2),.din(w_dff_A_qFR6XBNy6_2),.clk(gclk));
	jdff dff_B_csnaLUaJ0_1(.din(n618),.dout(w_dff_B_csnaLUaJ0_1),.clk(gclk));
	jdff dff_B_SEmiHP4u7_0(.din(n628),.dout(w_dff_B_SEmiHP4u7_0),.clk(gclk));
	jdff dff_A_81pCt3ZJ1_0(.dout(w_G322_0[0]),.din(w_dff_A_81pCt3ZJ1_0),.clk(gclk));
	jdff dff_B_wNpOitCb0_3(.din(G322),.dout(w_dff_B_wNpOitCb0_3),.clk(gclk));
	jdff dff_B_GH2siCI67_3(.din(w_dff_B_wNpOitCb0_3),.dout(w_dff_B_GH2siCI67_3),.clk(gclk));
	jdff dff_B_rX8Nivot9_3(.din(w_dff_B_GH2siCI67_3),.dout(w_dff_B_rX8Nivot9_3),.clk(gclk));
	jdff dff_A_eVb0pw6a8_1(.dout(w_n612_4[1]),.din(w_dff_A_eVb0pw6a8_1),.clk(gclk));
	jdff dff_A_izTLcR693_1(.dout(w_dff_A_eVb0pw6a8_1),.din(w_dff_A_izTLcR693_1),.clk(gclk));
	jdff dff_A_1HXeJx3I1_1(.dout(w_dff_A_izTLcR693_1),.din(w_dff_A_1HXeJx3I1_1),.clk(gclk));
	jdff dff_A_ItvJ0AUZ0_1(.dout(w_dff_A_1HXeJx3I1_1),.din(w_dff_A_ItvJ0AUZ0_1),.clk(gclk));
	jdff dff_A_4pTrGx9u1_1(.dout(w_dff_A_ItvJ0AUZ0_1),.din(w_dff_A_4pTrGx9u1_1),.clk(gclk));
	jdff dff_A_Xcd62Tim0_1(.dout(w_dff_A_4pTrGx9u1_1),.din(w_dff_A_Xcd62Tim0_1),.clk(gclk));
	jdff dff_A_kV4MqbCa6_1(.dout(w_dff_A_Xcd62Tim0_1),.din(w_dff_A_kV4MqbCa6_1),.clk(gclk));
	jdff dff_A_pftuPXJG7_1(.dout(w_dff_A_kV4MqbCa6_1),.din(w_dff_A_pftuPXJG7_1),.clk(gclk));
	jdff dff_A_ujHVhFXE2_0(.dout(w_n608_1[0]),.din(w_dff_A_ujHVhFXE2_0),.clk(gclk));
	jdff dff_A_Ag613vyg4_0(.dout(w_dff_A_ujHVhFXE2_0),.din(w_dff_A_Ag613vyg4_0),.clk(gclk));
	jdff dff_A_dg8jophn1_0(.dout(w_dff_A_Ag613vyg4_0),.din(w_dff_A_dg8jophn1_0),.clk(gclk));
	jdff dff_A_uHQJX5Vw1_0(.dout(w_dff_A_dg8jophn1_0),.din(w_dff_A_uHQJX5Vw1_0),.clk(gclk));
	jdff dff_A_vPuHMoXa2_0(.dout(w_dff_A_uHQJX5Vw1_0),.din(w_dff_A_vPuHMoXa2_0),.clk(gclk));
	jdff dff_A_eoNa2PPz0_0(.dout(w_dff_A_vPuHMoXa2_0),.din(w_dff_A_eoNa2PPz0_0),.clk(gclk));
	jdff dff_A_PmPtq17c4_0(.dout(w_dff_A_eoNa2PPz0_0),.din(w_dff_A_PmPtq17c4_0),.clk(gclk));
	jdff dff_A_6nzvRsWK0_0(.dout(w_dff_A_PmPtq17c4_0),.din(w_dff_A_6nzvRsWK0_0),.clk(gclk));
	jdff dff_A_Qi2CfUyN8_0(.dout(w_dff_A_6nzvRsWK0_0),.din(w_dff_A_Qi2CfUyN8_0),.clk(gclk));
	jdff dff_A_Kdl1A3t00_0(.dout(w_dff_A_Qi2CfUyN8_0),.din(w_dff_A_Kdl1A3t00_0),.clk(gclk));
	jdff dff_A_A0bUwg7l5_0(.dout(w_dff_A_Kdl1A3t00_0),.din(w_dff_A_A0bUwg7l5_0),.clk(gclk));
	jdff dff_A_ylJrylbW4_2(.dout(w_n608_1[2]),.din(w_dff_A_ylJrylbW4_2),.clk(gclk));
	jdff dff_A_LaKsi5FD4_2(.dout(w_dff_A_ylJrylbW4_2),.din(w_dff_A_LaKsi5FD4_2),.clk(gclk));
	jdff dff_A_KivU3g2Y0_2(.dout(w_dff_A_LaKsi5FD4_2),.din(w_dff_A_KivU3g2Y0_2),.clk(gclk));
	jdff dff_A_J1tWehzc5_2(.dout(w_dff_A_KivU3g2Y0_2),.din(w_dff_A_J1tWehzc5_2),.clk(gclk));
	jdff dff_A_T1KNWnat5_2(.dout(w_dff_A_J1tWehzc5_2),.din(w_dff_A_T1KNWnat5_2),.clk(gclk));
	jdff dff_A_iJjgRdQp3_2(.dout(w_dff_A_T1KNWnat5_2),.din(w_dff_A_iJjgRdQp3_2),.clk(gclk));
	jdff dff_A_ji8CAmEm2_2(.dout(w_dff_A_iJjgRdQp3_2),.din(w_dff_A_ji8CAmEm2_2),.clk(gclk));
	jdff dff_A_LszETj6i5_2(.dout(w_dff_A_ji8CAmEm2_2),.din(w_dff_A_LszETj6i5_2),.clk(gclk));
	jdff dff_A_CfZyoAll3_2(.dout(w_dff_A_LszETj6i5_2),.din(w_dff_A_CfZyoAll3_2),.clk(gclk));
	jdff dff_A_9vAQujb96_2(.dout(w_dff_A_CfZyoAll3_2),.din(w_dff_A_9vAQujb96_2),.clk(gclk));
	jdff dff_A_W5fxPdRt2_2(.dout(w_dff_A_9vAQujb96_2),.din(w_dff_A_W5fxPdRt2_2),.clk(gclk));
	jdff dff_A_Ben8Znh69_1(.dout(w_n608_0[1]),.din(w_dff_A_Ben8Znh69_1),.clk(gclk));
	jdff dff_A_g596W5QG4_1(.dout(w_dff_A_Ben8Znh69_1),.din(w_dff_A_g596W5QG4_1),.clk(gclk));
	jdff dff_A_EkXCf4t16_1(.dout(w_dff_A_g596W5QG4_1),.din(w_dff_A_EkXCf4t16_1),.clk(gclk));
	jdff dff_A_OBzN97CG2_1(.dout(w_dff_A_EkXCf4t16_1),.din(w_dff_A_OBzN97CG2_1),.clk(gclk));
	jdff dff_A_Ziy1fTaz3_1(.dout(w_dff_A_OBzN97CG2_1),.din(w_dff_A_Ziy1fTaz3_1),.clk(gclk));
	jdff dff_A_Rh16nUJt7_1(.dout(w_dff_A_Ziy1fTaz3_1),.din(w_dff_A_Rh16nUJt7_1),.clk(gclk));
	jdff dff_A_ogfxIjFq3_1(.dout(w_dff_A_Rh16nUJt7_1),.din(w_dff_A_ogfxIjFq3_1),.clk(gclk));
	jdff dff_A_V9S1PCU52_1(.dout(w_dff_A_ogfxIjFq3_1),.din(w_dff_A_V9S1PCU52_1),.clk(gclk));
	jdff dff_A_utYsbCW66_1(.dout(w_dff_A_V9S1PCU52_1),.din(w_dff_A_utYsbCW66_1),.clk(gclk));
	jdff dff_A_VPWo4PEw8_1(.dout(w_dff_A_utYsbCW66_1),.din(w_dff_A_VPWo4PEw8_1),.clk(gclk));
	jdff dff_A_yUSiJE2a0_1(.dout(w_dff_A_VPWo4PEw8_1),.din(w_dff_A_yUSiJE2a0_1),.clk(gclk));
	jdff dff_A_S8IxAVDR1_2(.dout(w_n608_0[2]),.din(w_dff_A_S8IxAVDR1_2),.clk(gclk));
	jdff dff_A_LXrKOMXU9_2(.dout(w_dff_A_S8IxAVDR1_2),.din(w_dff_A_LXrKOMXU9_2),.clk(gclk));
	jdff dff_A_sa20jRqe0_2(.dout(w_dff_A_LXrKOMXU9_2),.din(w_dff_A_sa20jRqe0_2),.clk(gclk));
	jdff dff_A_y1zRS86h4_2(.dout(w_dff_A_sa20jRqe0_2),.din(w_dff_A_y1zRS86h4_2),.clk(gclk));
	jdff dff_A_S2S9Tqky1_2(.dout(w_dff_A_y1zRS86h4_2),.din(w_dff_A_S2S9Tqky1_2),.clk(gclk));
	jdff dff_A_vvbmvctz9_2(.dout(w_dff_A_S2S9Tqky1_2),.din(w_dff_A_vvbmvctz9_2),.clk(gclk));
	jdff dff_A_pOHd292y6_2(.dout(w_dff_A_vvbmvctz9_2),.din(w_dff_A_pOHd292y6_2),.clk(gclk));
	jdff dff_A_FpweQpZM3_2(.dout(w_dff_A_pOHd292y6_2),.din(w_dff_A_FpweQpZM3_2),.clk(gclk));
	jdff dff_A_zH2JcY4f7_2(.dout(w_dff_A_FpweQpZM3_2),.din(w_dff_A_zH2JcY4f7_2),.clk(gclk));
	jdff dff_A_MFZomLcF0_2(.dout(w_dff_A_zH2JcY4f7_2),.din(w_dff_A_MFZomLcF0_2),.clk(gclk));
	jdff dff_A_YCIlTHLf2_2(.dout(w_dff_A_MFZomLcF0_2),.din(w_dff_A_YCIlTHLf2_2),.clk(gclk));
	jdff dff_B_h5FG6BeU4_0(.din(n570),.dout(w_dff_B_h5FG6BeU4_0),.clk(gclk));
	jdff dff_B_ISAkrs8o5_0(.din(w_dff_B_h5FG6BeU4_0),.dout(w_dff_B_ISAkrs8o5_0),.clk(gclk));
	jdff dff_B_CUucMEAh7_0(.din(n568),.dout(w_dff_B_CUucMEAh7_0),.clk(gclk));
	jdff dff_B_hy5ZWvia2_0(.din(w_dff_B_CUucMEAh7_0),.dout(w_dff_B_hy5ZWvia2_0),.clk(gclk));
	jdff dff_B_CqHJVKye5_0(.din(w_dff_B_hy5ZWvia2_0),.dout(w_dff_B_CqHJVKye5_0),.clk(gclk));
	jdff dff_A_iUfvIEz78_0(.dout(w_n567_0[0]),.din(w_dff_A_iUfvIEz78_0),.clk(gclk));
	jdff dff_A_7vTYN9o84_0(.dout(w_dff_A_iUfvIEz78_0),.din(w_dff_A_7vTYN9o84_0),.clk(gclk));
	jdff dff_A_afHYqFxH2_1(.dout(w_n554_3[1]),.din(w_dff_A_afHYqFxH2_1),.clk(gclk));
	jdff dff_A_zsQunHwU7_1(.dout(w_dff_A_afHYqFxH2_1),.din(w_dff_A_zsQunHwU7_1),.clk(gclk));
	jdff dff_A_Dp2CALI72_1(.dout(w_dff_A_zsQunHwU7_1),.din(w_dff_A_Dp2CALI72_1),.clk(gclk));
	jdff dff_A_AWNgwUnV3_2(.dout(w_n554_3[2]),.din(w_dff_A_AWNgwUnV3_2),.clk(gclk));
	jdff dff_A_CCeIWJGa4_2(.dout(w_dff_A_AWNgwUnV3_2),.din(w_dff_A_CCeIWJGa4_2),.clk(gclk));
	jdff dff_A_AQIsk6hs2_2(.dout(w_dff_A_CCeIWJGa4_2),.din(w_dff_A_AQIsk6hs2_2),.clk(gclk));
	jdff dff_B_nMMtbWXq2_2(.din(n565),.dout(w_dff_B_nMMtbWXq2_2),.clk(gclk));
	jdff dff_B_US2VQ0nN2_2(.din(w_dff_B_nMMtbWXq2_2),.dout(w_dff_B_US2VQ0nN2_2),.clk(gclk));
	jdff dff_B_j0ovojQ30_2(.din(w_dff_B_US2VQ0nN2_2),.dout(w_dff_B_j0ovojQ30_2),.clk(gclk));
	jdff dff_B_6rRYUcVr6_2(.din(w_dff_B_j0ovojQ30_2),.dout(w_dff_B_6rRYUcVr6_2),.clk(gclk));
	jdff dff_B_jQEs3KYQ8_2(.din(w_dff_B_6rRYUcVr6_2),.dout(w_dff_B_jQEs3KYQ8_2),.clk(gclk));
	jdff dff_B_UkCu8P9U7_2(.din(w_dff_B_jQEs3KYQ8_2),.dout(w_dff_B_UkCu8P9U7_2),.clk(gclk));
	jdff dff_B_X6l0t1JA9_2(.din(w_dff_B_UkCu8P9U7_2),.dout(w_dff_B_X6l0t1JA9_2),.clk(gclk));
	jdff dff_B_kEvGkueG5_2(.din(w_dff_B_X6l0t1JA9_2),.dout(w_dff_B_kEvGkueG5_2),.clk(gclk));
	jdff dff_B_5RQQ68ig4_2(.din(w_dff_B_kEvGkueG5_2),.dout(w_dff_B_5RQQ68ig4_2),.clk(gclk));
	jdff dff_B_NutjzFEL9_2(.din(w_dff_B_5RQQ68ig4_2),.dout(w_dff_B_NutjzFEL9_2),.clk(gclk));
	jdff dff_B_rCqzEXuV5_2(.din(w_dff_B_NutjzFEL9_2),.dout(w_dff_B_rCqzEXuV5_2),.clk(gclk));
	jdff dff_B_thoodCAy6_2(.din(w_dff_B_rCqzEXuV5_2),.dout(w_dff_B_thoodCAy6_2),.clk(gclk));
	jdff dff_B_S2SNhrZX6_2(.din(w_dff_B_thoodCAy6_2),.dout(w_dff_B_S2SNhrZX6_2),.clk(gclk));
	jdff dff_A_hTgHDsrK5_1(.dout(w_n1162_0[1]),.din(w_dff_A_hTgHDsrK5_1),.clk(gclk));
	jdff dff_B_LDRONa5J9_0(.din(n1161),.dout(w_dff_B_LDRONa5J9_0),.clk(gclk));
	jdff dff_B_8uFYQU0E4_0(.din(w_dff_B_LDRONa5J9_0),.dout(w_dff_B_8uFYQU0E4_0),.clk(gclk));
	jdff dff_B_k2RQ2kjo3_0(.din(n1158),.dout(w_dff_B_k2RQ2kjo3_0),.clk(gclk));
	jdff dff_B_beaLWjaP9_0(.din(w_dff_B_k2RQ2kjo3_0),.dout(w_dff_B_beaLWjaP9_0),.clk(gclk));
	jdff dff_B_bg2628tI6_0(.din(w_dff_B_beaLWjaP9_0),.dout(w_dff_B_bg2628tI6_0),.clk(gclk));
	jdff dff_B_1sI4oKiB0_0(.din(w_dff_B_bg2628tI6_0),.dout(w_dff_B_1sI4oKiB0_0),.clk(gclk));
	jdff dff_B_XgRgISjX1_0(.din(w_dff_B_1sI4oKiB0_0),.dout(w_dff_B_XgRgISjX1_0),.clk(gclk));
	jdff dff_B_VuOjOOvv5_0(.din(n1157),.dout(w_dff_B_VuOjOOvv5_0),.clk(gclk));
	jdff dff_B_Lq59G3kr3_0(.din(w_dff_B_VuOjOOvv5_0),.dout(w_dff_B_Lq59G3kr3_0),.clk(gclk));
	jdff dff_B_mnHUxTSm7_0(.din(n1155),.dout(w_dff_B_mnHUxTSm7_0),.clk(gclk));
	jdff dff_B_jzkxmxX52_0(.din(w_dff_B_mnHUxTSm7_0),.dout(w_dff_B_jzkxmxX52_0),.clk(gclk));
	jdff dff_B_kddCkst46_1(.din(n1143),.dout(w_dff_B_kddCkst46_1),.clk(gclk));
	jdff dff_B_ORN9O6023_1(.din(w_dff_B_kddCkst46_1),.dout(w_dff_B_ORN9O6023_1),.clk(gclk));
	jdff dff_B_5yDNasKG3_1(.din(n1145),.dout(w_dff_B_5yDNasKG3_1),.clk(gclk));
	jdff dff_B_GuNW2e8p9_1(.din(n1148),.dout(w_dff_B_GuNW2e8p9_1),.clk(gclk));
	jdff dff_A_4YM7diBN0_1(.dout(w_n899_0[1]),.din(w_dff_A_4YM7diBN0_1),.clk(gclk));
	jdff dff_A_byatC4aG6_1(.dout(w_G87_1[1]),.din(w_dff_A_byatC4aG6_1),.clk(gclk));
	jdff dff_A_hHFRDDwG8_2(.dout(w_G87_1[2]),.din(w_dff_A_hHFRDDwG8_2),.clk(gclk));
	jdff dff_A_JY0B51aq6_1(.dout(w_G77_2[1]),.din(w_dff_A_JY0B51aq6_1),.clk(gclk));
	jdff dff_A_LJCRtSSc7_1(.dout(w_dff_A_JY0B51aq6_1),.din(w_dff_A_LJCRtSSc7_1),.clk(gclk));
	jdff dff_A_2wjzWZAY2_1(.dout(w_dff_A_LJCRtSSc7_1),.din(w_dff_A_2wjzWZAY2_1),.clk(gclk));
	jdff dff_A_E9E5rxLQ7_1(.dout(w_dff_A_2wjzWZAY2_1),.din(w_dff_A_E9E5rxLQ7_1),.clk(gclk));
	jdff dff_A_WqWUz2897_2(.dout(w_G77_2[2]),.din(w_dff_A_WqWUz2897_2),.clk(gclk));
	jdff dff_A_WoNmbVIo1_2(.dout(w_dff_A_WqWUz2897_2),.din(w_dff_A_WoNmbVIo1_2),.clk(gclk));
	jdff dff_A_hCTVNgxW4_2(.dout(w_dff_A_WoNmbVIo1_2),.din(w_dff_A_hCTVNgxW4_2),.clk(gclk));
	jdff dff_A_UPue7mKt7_2(.dout(w_dff_A_hCTVNgxW4_2),.din(w_dff_A_UPue7mKt7_2),.clk(gclk));
	jdff dff_A_VPKwfkVC7_1(.dout(w_G283_1[1]),.din(w_dff_A_VPKwfkVC7_1),.clk(gclk));
	jdff dff_A_JH9MCF8f4_0(.dout(w_n148_3[0]),.din(w_dff_A_JH9MCF8f4_0),.clk(gclk));
	jdff dff_A_BxsKgBGG5_0(.dout(w_dff_A_JH9MCF8f4_0),.din(w_dff_A_BxsKgBGG5_0),.clk(gclk));
	jdff dff_A_BhkLDNvD8_0(.dout(w_dff_A_BxsKgBGG5_0),.din(w_dff_A_BhkLDNvD8_0),.clk(gclk));
	jdff dff_A_xk3kCVKM2_0(.dout(w_dff_A_BhkLDNvD8_0),.din(w_dff_A_xk3kCVKM2_0),.clk(gclk));
	jdff dff_A_ynk5dqSb2_2(.dout(w_n148_3[2]),.din(w_dff_A_ynk5dqSb2_2),.clk(gclk));
	jdff dff_A_Ku9B3Y2T2_2(.dout(w_dff_A_ynk5dqSb2_2),.din(w_dff_A_Ku9B3Y2T2_2),.clk(gclk));
	jdff dff_A_ZBccMnZ21_2(.dout(w_dff_A_Ku9B3Y2T2_2),.din(w_dff_A_ZBccMnZ21_2),.clk(gclk));
	jdff dff_A_iBOwVAhb4_1(.dout(w_G294_1[1]),.din(w_dff_A_iBOwVAhb4_1),.clk(gclk));
	jdff dff_B_nx93J3LY3_1(.din(n1128),.dout(w_dff_B_nx93J3LY3_1),.clk(gclk));
	jdff dff_B_YnLdvlym2_1(.din(n1130),.dout(w_dff_B_YnLdvlym2_1),.clk(gclk));
	jdff dff_B_ui9JvqB01_1(.din(n1133),.dout(w_dff_B_ui9JvqB01_1),.clk(gclk));
	jdff dff_B_07FqMLME8_0(.din(n1134),.dout(w_dff_B_07FqMLME8_0),.clk(gclk));
	jdff dff_A_dNdWUtir8_1(.dout(w_G150_1[1]),.din(w_dff_A_dNdWUtir8_1),.clk(gclk));
	jdff dff_A_HGXab7lh5_2(.dout(w_G150_1[2]),.din(w_dff_A_HGXab7lh5_2),.clk(gclk));
	jdff dff_A_3k1m8a2A3_0(.dout(w_G128_0[0]),.din(w_dff_A_3k1m8a2A3_0),.clk(gclk));
	jdff dff_B_9LjZadz51_3(.din(G128),.dout(w_dff_B_9LjZadz51_3),.clk(gclk));
	jdff dff_B_V6JONzVg6_3(.din(w_dff_B_9LjZadz51_3),.dout(w_dff_B_V6JONzVg6_3),.clk(gclk));
	jdff dff_B_Nv8zABFN6_3(.din(w_dff_B_V6JONzVg6_3),.dout(w_dff_B_Nv8zABFN6_3),.clk(gclk));
	jdff dff_B_GdT3MNyE9_1(.din(n1124),.dout(w_dff_B_GdT3MNyE9_1),.clk(gclk));
	jdff dff_B_LpNfrY359_0(.din(n1126),.dout(w_dff_B_LpNfrY359_0),.clk(gclk));
	jdff dff_A_iO2LrXBq8_0(.dout(w_n612_1[0]),.din(w_dff_A_iO2LrXBq8_0),.clk(gclk));
	jdff dff_A_SLH6Xzgr1_1(.dout(w_n612_1[1]),.din(w_dff_A_SLH6Xzgr1_1),.clk(gclk));
	jdff dff_A_60JJg4zp8_1(.dout(w_dff_A_SLH6Xzgr1_1),.din(w_dff_A_60JJg4zp8_1),.clk(gclk));
	jdff dff_A_jRhn2qcD5_1(.dout(w_dff_A_60JJg4zp8_1),.din(w_dff_A_jRhn2qcD5_1),.clk(gclk));
	jdff dff_A_ti8Wxqyt9_1(.dout(w_dff_A_jRhn2qcD5_1),.din(w_dff_A_ti8Wxqyt9_1),.clk(gclk));
	jdff dff_A_6ZpunHw50_1(.dout(w_dff_A_ti8Wxqyt9_1),.din(w_dff_A_6ZpunHw50_1),.clk(gclk));
	jdff dff_A_tDWTM7ME4_1(.dout(w_dff_A_6ZpunHw50_1),.din(w_dff_A_tDWTM7ME4_1),.clk(gclk));
	jdff dff_A_iA6ky1Cq2_1(.dout(w_dff_A_tDWTM7ME4_1),.din(w_dff_A_iA6ky1Cq2_1),.clk(gclk));
	jdff dff_A_D22jo48r6_1(.dout(w_n999_0[1]),.din(w_dff_A_D22jo48r6_1),.clk(gclk));
	jdff dff_A_rkOouUbH5_2(.dout(w_n764_0[2]),.din(w_dff_A_rkOouUbH5_2),.clk(gclk));
	jdff dff_A_CfidJJKC8_2(.dout(w_dff_A_rkOouUbH5_2),.din(w_dff_A_CfidJJKC8_2),.clk(gclk));
	jdff dff_B_TULLagoq1_0(.din(n763),.dout(w_dff_B_TULLagoq1_0),.clk(gclk));
	jdff dff_B_cPx4GLvs2_0(.din(w_dff_B_TULLagoq1_0),.dout(w_dff_B_cPx4GLvs2_0),.clk(gclk));
	jdff dff_B_f1Dh1Z274_0(.din(n761),.dout(w_dff_B_f1Dh1Z274_0),.clk(gclk));
	jdff dff_B_sc5ECryo4_0(.din(w_dff_B_f1Dh1Z274_0),.dout(w_dff_B_sc5ECryo4_0),.clk(gclk));
	jdff dff_A_IUdNnhry2_0(.dout(w_n760_0[0]),.din(w_dff_A_IUdNnhry2_0),.clk(gclk));
	jdff dff_B_KM6fBycT4_0(.din(n997),.dout(w_dff_B_KM6fBycT4_0),.clk(gclk));
	jdff dff_B_QrDDYXQC2_0(.din(w_dff_B_KM6fBycT4_0),.dout(w_dff_B_QrDDYXQC2_0),.clk(gclk));
	jdff dff_B_Knx9thml1_0(.din(w_dff_B_QrDDYXQC2_0),.dout(w_dff_B_Knx9thml1_0),.clk(gclk));
	jdff dff_B_uZqli6Na3_0(.din(w_dff_B_Knx9thml1_0),.dout(w_dff_B_uZqli6Na3_0),.clk(gclk));
	jdff dff_B_wPggN8AG0_0(.din(w_dff_B_uZqli6Na3_0),.dout(w_dff_B_wPggN8AG0_0),.clk(gclk));
	jdff dff_A_6HEAOcvv8_2(.dout(w_n554_1[2]),.din(w_dff_A_6HEAOcvv8_2),.clk(gclk));
	jdff dff_A_wkG5dVVG0_1(.dout(w_n519_0[1]),.din(w_dff_A_wkG5dVVG0_1),.clk(gclk));
	jdff dff_A_I4QRRSBC3_1(.dout(w_dff_A_wkG5dVVG0_1),.din(w_dff_A_I4QRRSBC3_1),.clk(gclk));
	jdff dff_A_gAq1C1p84_2(.dout(w_n519_0[2]),.din(w_dff_A_gAq1C1p84_2),.clk(gclk));
	jdff dff_A_RqxBxNm63_2(.dout(w_dff_A_gAq1C1p84_2),.din(w_dff_A_RqxBxNm63_2),.clk(gclk));
	jdff dff_A_Tgsmx2AP1_0(.dout(w_n548_0[0]),.din(w_dff_A_Tgsmx2AP1_0),.clk(gclk));
	jdff dff_A_2gKLDoFq8_1(.dout(w_n439_0[1]),.din(w_dff_A_2gKLDoFq8_1),.clk(gclk));
	jdff dff_A_Jq6HlDRh1_1(.dout(w_dff_A_2gKLDoFq8_1),.din(w_dff_A_Jq6HlDRh1_1),.clk(gclk));
	jdff dff_A_xygUTBYQ0_1(.dout(w_dff_A_Jq6HlDRh1_1),.din(w_dff_A_xygUTBYQ0_1),.clk(gclk));
	jdff dff_A_KWWvRnfy9_1(.dout(w_dff_A_xygUTBYQ0_1),.din(w_dff_A_KWWvRnfy9_1),.clk(gclk));
	jdff dff_B_kRL33Kwb6_1(.din(n441),.dout(w_dff_B_kRL33Kwb6_1),.clk(gclk));
	jdff dff_B_X5McmxHP1_1(.din(w_dff_B_kRL33Kwb6_1),.dout(w_dff_B_X5McmxHP1_1),.clk(gclk));
	jdff dff_A_Ql0JBR2b8_1(.dout(w_n436_0[1]),.din(w_dff_A_Ql0JBR2b8_1),.clk(gclk));
	jdff dff_B_tzQ4OxgE2_1(.din(n424),.dout(w_dff_B_tzQ4OxgE2_1),.clk(gclk));
	jdff dff_B_IkMZBkBp9_0(.din(n434),.dout(w_dff_B_IkMZBkBp9_0),.clk(gclk));
	jdff dff_B_6AA9bqyU6_0(.din(n423),.dout(w_dff_B_6AA9bqyU6_0),.clk(gclk));
	jdff dff_B_kQIUHOkP2_0(.din(w_dff_B_6AA9bqyU6_0),.dout(w_dff_B_kQIUHOkP2_0),.clk(gclk));
	jdff dff_B_DmEc0be85_1(.din(n413),.dout(w_dff_B_DmEc0be85_1),.clk(gclk));
	jdff dff_A_yZBgr7T34_0(.dout(w_G226_1[0]),.din(w_dff_A_yZBgr7T34_0),.clk(gclk));
	jdff dff_A_i2cl3Bp49_0(.dout(w_dff_A_yZBgr7T34_0),.din(w_dff_A_i2cl3Bp49_0),.clk(gclk));
	jdff dff_B_rUgMDvnS7_1(.din(n493),.dout(w_dff_B_rUgMDvnS7_1),.clk(gclk));
	jdff dff_B_wq0pYMBx5_1(.din(w_dff_B_rUgMDvnS7_1),.dout(w_dff_B_wq0pYMBx5_1),.clk(gclk));
	jdff dff_A_pmyIkI1G1_0(.dout(w_n516_0[0]),.din(w_dff_A_pmyIkI1G1_0),.clk(gclk));
	jdff dff_A_E2BCCOSl0_0(.dout(w_dff_A_pmyIkI1G1_0),.din(w_dff_A_E2BCCOSl0_0),.clk(gclk));
	jdff dff_B_eHtuai9V9_0(.din(n514),.dout(w_dff_B_eHtuai9V9_0),.clk(gclk));
	jdff dff_B_DaWjeVjL0_1(.din(n485),.dout(w_dff_B_DaWjeVjL0_1),.clk(gclk));
	jdff dff_B_bgCGocnM4_1(.din(n496),.dout(w_dff_B_bgCGocnM4_1),.clk(gclk));
	jdff dff_B_nwC5A8HM1_1(.din(w_dff_B_bgCGocnM4_1),.dout(w_dff_B_nwC5A8HM1_1),.clk(gclk));
	jdff dff_B_g2sFFUCp9_1(.din(w_dff_B_nwC5A8HM1_1),.dout(w_dff_B_g2sFFUCp9_1),.clk(gclk));
	jdff dff_B_ZlgEJhOi6_0(.din(n505),.dout(w_dff_B_ZlgEJhOi6_0),.clk(gclk));
	jdff dff_B_4GyJWtJN6_0(.din(w_dff_B_ZlgEJhOi6_0),.dout(w_dff_B_4GyJWtJN6_0),.clk(gclk));
	jdff dff_B_pwH9jyPc2_1(.din(n497),.dout(w_dff_B_pwH9jyPc2_1),.clk(gclk));
	jdff dff_B_GXNaKhtp0_1(.din(w_dff_B_pwH9jyPc2_1),.dout(w_dff_B_GXNaKhtp0_1),.clk(gclk));
	jdff dff_B_KQl9HTF33_1(.din(w_dff_B_GXNaKhtp0_1),.dout(w_dff_B_KQl9HTF33_1),.clk(gclk));
	jdff dff_A_Rva1AEKD2_1(.dout(w_n541_0[1]),.din(w_dff_A_Rva1AEKD2_1),.clk(gclk));
	jdff dff_A_fcI5NC2f2_1(.dout(w_dff_A_Rva1AEKD2_1),.din(w_dff_A_fcI5NC2f2_1),.clk(gclk));
	jdff dff_B_OqO96hog7_1(.din(n456),.dout(w_dff_B_OqO96hog7_1),.clk(gclk));
	jdff dff_B_sob5fowR5_1(.din(w_dff_B_OqO96hog7_1),.dout(w_dff_B_sob5fowR5_1),.clk(gclk));
	jdff dff_A_DfSwjIls9_0(.dout(w_n483_0[0]),.din(w_dff_A_DfSwjIls9_0),.clk(gclk));
	jdff dff_A_GcD66brr2_0(.dout(w_dff_A_DfSwjIls9_0),.din(w_dff_A_GcD66brr2_0),.clk(gclk));
	jdff dff_A_Hl1mrqai0_0(.dout(w_dff_A_GcD66brr2_0),.din(w_dff_A_Hl1mrqai0_0),.clk(gclk));
	jdff dff_A_sYv13dku0_0(.dout(w_dff_A_Hl1mrqai0_0),.din(w_dff_A_sYv13dku0_0),.clk(gclk));
	jdff dff_B_QXqYkzoH9_0(.din(n481),.dout(w_dff_B_QXqYkzoH9_0),.clk(gclk));
	jdff dff_A_Y1zkbMin2_1(.dout(w_G226_0[1]),.din(w_dff_A_Y1zkbMin2_1),.clk(gclk));
	jdff dff_A_VGVZ5Om46_1(.dout(w_dff_A_Y1zkbMin2_1),.din(w_dff_A_VGVZ5Om46_1),.clk(gclk));
	jdff dff_A_bdTsspxu3_2(.dout(w_G226_0[2]),.din(w_dff_A_bdTsspxu3_2),.clk(gclk));
	jdff dff_A_0wvv5lHZ5_2(.dout(w_dff_A_bdTsspxu3_2),.din(w_dff_A_0wvv5lHZ5_2),.clk(gclk));
	jdff dff_A_7l3Pgq8W7_2(.dout(w_dff_A_0wvv5lHZ5_2),.din(w_dff_A_7l3Pgq8W7_2),.clk(gclk));
	jdff dff_A_Aw8GGBk42_2(.dout(w_dff_A_7l3Pgq8W7_2),.din(w_dff_A_Aw8GGBk42_2),.clk(gclk));
	jdff dff_B_O8CWMqll9_1(.din(n448),.dout(w_dff_B_O8CWMqll9_1),.clk(gclk));
	jdff dff_B_p1GlhHg72_1(.din(G222),.dout(w_dff_B_p1GlhHg72_1),.clk(gclk));
	jdff dff_B_6p6SfMK66_1(.din(w_dff_B_p1GlhHg72_1),.dout(w_dff_B_6p6SfMK66_1),.clk(gclk));
	jdff dff_A_NVMS29z04_0(.dout(w_n430_0[0]),.din(w_dff_A_NVMS29z04_0),.clk(gclk));
	jdff dff_B_aFDTMb6B2_2(.din(n430),.dout(w_dff_B_aFDTMb6B2_2),.clk(gclk));
	jdff dff_A_iZRRhRrA3_1(.dout(w_G77_3[1]),.din(w_dff_A_iZRRhRrA3_1),.clk(gclk));
	jdff dff_A_mjNH1ppj0_1(.dout(w_dff_A_iZRRhRrA3_1),.din(w_dff_A_mjNH1ppj0_1),.clk(gclk));
	jdff dff_A_f4ZUCAnr5_1(.dout(w_dff_A_mjNH1ppj0_1),.din(w_dff_A_f4ZUCAnr5_1),.clk(gclk));
	jdff dff_B_iyPl7ZmR6_2(.din(G223),.dout(w_dff_B_iyPl7ZmR6_2),.clk(gclk));
	jdff dff_B_KYm3OC3V3_2(.din(w_dff_B_iyPl7ZmR6_2),.dout(w_dff_B_KYm3OC3V3_2),.clk(gclk));
	jdff dff_B_MDlhKS9x1_1(.din(n459),.dout(w_dff_B_MDlhKS9x1_1),.clk(gclk));
	jdff dff_B_okKJV17k9_1(.din(w_dff_B_MDlhKS9x1_1),.dout(w_dff_B_okKJV17k9_1),.clk(gclk));
	jdff dff_B_fXFLWVgQ2_1(.din(w_dff_B_okKJV17k9_1),.dout(w_dff_B_fXFLWVgQ2_1),.clk(gclk));
	jdff dff_B_sKt8HdsP3_0(.din(n472),.dout(w_dff_B_sKt8HdsP3_0),.clk(gclk));
	jdff dff_B_BmUIe2270_0(.din(w_dff_B_sKt8HdsP3_0),.dout(w_dff_B_BmUIe2270_0),.clk(gclk));
	jdff dff_A_se3X5d4g7_2(.dout(w_n185_1[2]),.din(w_dff_A_se3X5d4g7_2),.clk(gclk));
	jdff dff_B_Sggb8bRB2_1(.din(n460),.dout(w_dff_B_Sggb8bRB2_1),.clk(gclk));
	jdff dff_B_j1vmASJy6_1(.din(n461),.dout(w_dff_B_j1vmASJy6_1),.clk(gclk));
	jdff dff_B_1IiMTn0s3_1(.din(w_dff_B_j1vmASJy6_1),.dout(w_dff_B_1IiMTn0s3_1),.clk(gclk));
	jdff dff_A_UtVkimCc4_1(.dout(w_n75_0[1]),.din(w_dff_A_UtVkimCc4_1),.clk(gclk));
	jdff dff_A_R3DlfM8k2_1(.dout(w_dff_A_UtVkimCc4_1),.din(w_dff_A_R3DlfM8k2_1),.clk(gclk));
	jdff dff_A_Zz5ApCGF9_1(.dout(w_dff_A_R3DlfM8k2_1),.din(w_dff_A_Zz5ApCGF9_1),.clk(gclk));
	jdff dff_A_wbXxIzL69_2(.dout(w_n75_0[2]),.din(w_dff_A_wbXxIzL69_2),.clk(gclk));
	jdff dff_A_UhyvKCbr2_2(.dout(w_dff_A_wbXxIzL69_2),.din(w_dff_A_UhyvKCbr2_2),.clk(gclk));
	jdff dff_A_ZMc46jzT5_2(.dout(w_dff_A_UhyvKCbr2_2),.din(w_dff_A_ZMc46jzT5_2),.clk(gclk));
	jdff dff_A_efmkBkH97_2(.dout(w_dff_A_ZMc46jzT5_2),.din(w_dff_A_efmkBkH97_2),.clk(gclk));
	jdff dff_A_k7Tm4JLD1_1(.dout(w_n74_0[1]),.din(w_dff_A_k7Tm4JLD1_1),.clk(gclk));
	jdff dff_A_NQWsafb08_1(.dout(w_dff_A_k7Tm4JLD1_1),.din(w_dff_A_NQWsafb08_1),.clk(gclk));
	jdff dff_A_Q7OJ38FA2_1(.dout(w_dff_A_NQWsafb08_1),.din(w_dff_A_Q7OJ38FA2_1),.clk(gclk));
	jdff dff_A_6lOqnehS9_2(.dout(w_n74_0[2]),.din(w_dff_A_6lOqnehS9_2),.clk(gclk));
	jdff dff_A_j7xJR0ii1_2(.dout(w_dff_A_6lOqnehS9_2),.din(w_dff_A_j7xJR0ii1_2),.clk(gclk));
	jdff dff_A_T3yNR4nP6_0(.dout(w_n73_2[0]),.din(w_dff_A_T3yNR4nP6_0),.clk(gclk));
	jdff dff_A_cOaJiuwx8_0(.dout(w_dff_A_T3yNR4nP6_0),.din(w_dff_A_cOaJiuwx8_0),.clk(gclk));
	jdff dff_A_tYBCD6H65_2(.dout(w_n73_2[2]),.din(w_dff_A_tYBCD6H65_2),.clk(gclk));
	jdff dff_A_jZYY5mXL9_2(.dout(w_n73_0[2]),.din(w_dff_A_jZYY5mXL9_2),.clk(gclk));
	jdff dff_A_qGQbUysa8_2(.dout(w_dff_A_jZYY5mXL9_2),.din(w_dff_A_qGQbUysa8_2),.clk(gclk));
	jdff dff_A_Bkc40ouF1_2(.dout(w_dff_A_qGQbUysa8_2),.din(w_dff_A_Bkc40ouF1_2),.clk(gclk));
	jdff dff_A_MDo3JADq1_1(.dout(w_G50_5[1]),.din(w_dff_A_MDo3JADq1_1),.clk(gclk));
	jdff dff_A_kd626oGo4_1(.dout(w_dff_A_MDo3JADq1_1),.din(w_dff_A_kd626oGo4_1),.clk(gclk));
	jdff dff_A_wySSWbT54_1(.dout(w_dff_A_kd626oGo4_1),.din(w_dff_A_wySSWbT54_1),.clk(gclk));
	jdff dff_A_pOseXtjT4_0(.dout(w_G50_4[0]),.din(w_dff_A_pOseXtjT4_0),.clk(gclk));
	jdff dff_A_ErXiBYYZ2_0(.dout(w_dff_A_pOseXtjT4_0),.din(w_dff_A_ErXiBYYZ2_0),.clk(gclk));
	jdff dff_A_cR9FzrOM6_1(.dout(w_G50_4[1]),.din(w_dff_A_cR9FzrOM6_1),.clk(gclk));
	jdff dff_A_B5q9nHKd8_0(.dout(w_G50_1[0]),.din(w_dff_A_B5q9nHKd8_0),.clk(gclk));
	jdff dff_A_9fkugbRV3_2(.dout(w_G50_1[2]),.din(w_dff_A_9fkugbRV3_2),.clk(gclk));
	jdff dff_A_ALYf8q0U3_2(.dout(w_dff_A_9fkugbRV3_2),.din(w_dff_A_ALYf8q0U3_2),.clk(gclk));
	jdff dff_A_FhmdJnKA2_2(.dout(w_dff_A_ALYf8q0U3_2),.din(w_dff_A_FhmdJnKA2_2),.clk(gclk));
	jdff dff_A_T6Lcc6IH2_2(.dout(w_dff_A_FhmdJnKA2_2),.din(w_dff_A_T6Lcc6IH2_2),.clk(gclk));
	jdff dff_A_X1hUSW124_0(.dout(w_G384_0),.din(w_dff_A_X1hUSW124_0),.clk(gclk));
	jdff dff_A_ogpRhe583_0(.dout(w_dff_A_X1hUSW124_0),.din(w_dff_A_ogpRhe583_0),.clk(gclk));
	jdff dff_A_3yl5nL2Z1_0(.dout(w_n750_0[0]),.din(w_dff_A_3yl5nL2Z1_0),.clk(gclk));
	jdff dff_A_lSMlxxfa2_0(.dout(w_dff_A_3yl5nL2Z1_0),.din(w_dff_A_lSMlxxfa2_0),.clk(gclk));
	jdff dff_B_JFbHVnB53_0(.din(n747),.dout(w_dff_B_JFbHVnB53_0),.clk(gclk));
	jdff dff_B_vGkxd8xS3_0(.din(w_dff_B_JFbHVnB53_0),.dout(w_dff_B_vGkxd8xS3_0),.clk(gclk));
	jdff dff_B_r4LG1yPQ1_0(.din(w_dff_B_vGkxd8xS3_0),.dout(w_dff_B_r4LG1yPQ1_0),.clk(gclk));
	jdff dff_B_xLr7nSLd4_0(.din(n746),.dout(w_dff_B_xLr7nSLd4_0),.clk(gclk));
	jdff dff_B_QhMunovb1_0(.din(w_dff_B_xLr7nSLd4_0),.dout(w_dff_B_QhMunovb1_0),.clk(gclk));
	jdff dff_B_5HwZXw286_0(.din(w_dff_B_QhMunovb1_0),.dout(w_dff_B_5HwZXw286_0),.clk(gclk));
	jdff dff_B_8PHEd5ke3_0(.din(w_dff_B_5HwZXw286_0),.dout(w_dff_B_8PHEd5ke3_0),.clk(gclk));
	jdff dff_B_HgA4b9FY1_0(.din(n744),.dout(w_dff_B_HgA4b9FY1_0),.clk(gclk));
	jdff dff_B_Ppn9qytr3_0(.din(w_dff_B_HgA4b9FY1_0),.dout(w_dff_B_Ppn9qytr3_0),.clk(gclk));
	jdff dff_A_pBq5s4Ky8_2(.dout(w_n605_1[2]),.din(w_dff_A_pBq5s4Ky8_2),.clk(gclk));
	jdff dff_A_LWd1eegR5_2(.dout(w_dff_A_pBq5s4Ky8_2),.din(w_dff_A_LWd1eegR5_2),.clk(gclk));
	jdff dff_A_qpMqPPcq4_2(.dout(w_dff_A_LWd1eegR5_2),.din(w_dff_A_qpMqPPcq4_2),.clk(gclk));
	jdff dff_A_TgSkigYm6_2(.dout(w_dff_A_qpMqPPcq4_2),.din(w_dff_A_TgSkigYm6_2),.clk(gclk));
	jdff dff_A_U1yV6sTq2_2(.dout(w_dff_A_TgSkigYm6_2),.din(w_dff_A_U1yV6sTq2_2),.clk(gclk));
	jdff dff_A_cxDIl5xZ8_2(.dout(w_dff_A_U1yV6sTq2_2),.din(w_dff_A_cxDIl5xZ8_2),.clk(gclk));
	jdff dff_A_ae2eSZrV7_2(.dout(w_dff_A_cxDIl5xZ8_2),.din(w_dff_A_ae2eSZrV7_2),.clk(gclk));
	jdff dff_A_tv0YYWOD6_2(.dout(w_dff_A_ae2eSZrV7_2),.din(w_dff_A_tv0YYWOD6_2),.clk(gclk));
	jdff dff_A_QIOLY1di5_0(.dout(w_n604_2[0]),.din(w_dff_A_QIOLY1di5_0),.clk(gclk));
	jdff dff_A_Js16njrf8_0(.dout(w_dff_A_QIOLY1di5_0),.din(w_dff_A_Js16njrf8_0),.clk(gclk));
	jdff dff_A_WyZX4gsb9_0(.dout(w_dff_A_Js16njrf8_0),.din(w_dff_A_WyZX4gsb9_0),.clk(gclk));
	jdff dff_A_7dGQOBZh0_0(.dout(w_dff_A_WyZX4gsb9_0),.din(w_dff_A_7dGQOBZh0_0),.clk(gclk));
	jdff dff_B_nCPTWesU8_1(.din(n721),.dout(w_dff_B_nCPTWesU8_1),.clk(gclk));
	jdff dff_B_FVLNdNhN9_1(.din(w_dff_B_nCPTWesU8_1),.dout(w_dff_B_FVLNdNhN9_1),.clk(gclk));
	jdff dff_B_DDUVIJFg5_1(.din(n727),.dout(w_dff_B_DDUVIJFg5_1),.clk(gclk));
	jdff dff_B_oi0MVyjt8_1(.din(n730),.dout(w_dff_B_oi0MVyjt8_1),.clk(gclk));
	jdff dff_B_BzC8fKGl8_1(.din(n733),.dout(w_dff_B_BzC8fKGl8_1),.clk(gclk));
	jdff dff_B_ipLwlcnj3_0(.din(n734),.dout(w_dff_B_ipLwlcnj3_0),.clk(gclk));
	jdff dff_A_hARDuVkP8_0(.dout(w_G294_2[0]),.din(w_dff_A_hARDuVkP8_0),.clk(gclk));
	jdff dff_A_QcckcgpA9_0(.dout(w_G116_3[0]),.din(w_dff_A_QcckcgpA9_0),.clk(gclk));
	jdff dff_A_zRY7bSLT2_0(.dout(w_dff_A_QcckcgpA9_0),.din(w_dff_A_zRY7bSLT2_0),.clk(gclk));
	jdff dff_A_a7FNnu3y0_0(.dout(w_dff_A_zRY7bSLT2_0),.din(w_dff_A_a7FNnu3y0_0),.clk(gclk));
	jdff dff_A_FTZodH591_2(.dout(w_G116_3[2]),.din(w_dff_A_FTZodH591_2),.clk(gclk));
	jdff dff_A_xytoGJ765_2(.dout(w_dff_A_FTZodH591_2),.din(w_dff_A_xytoGJ765_2),.clk(gclk));
	jdff dff_A_K9gIku7k7_0(.dout(w_G33_5[0]),.din(w_dff_A_K9gIku7k7_0),.clk(gclk));
	jdff dff_A_zKMlK3M14_2(.dout(w_G33_5[2]),.din(w_dff_A_zKMlK3M14_2),.clk(gclk));
	jdff dff_A_TeDTVq7P5_2(.dout(w_dff_A_zKMlK3M14_2),.din(w_dff_A_TeDTVq7P5_2),.clk(gclk));
	jdff dff_B_1L2my1Ce8_1(.din(n722),.dout(w_dff_B_1L2my1Ce8_1),.clk(gclk));
	jdff dff_B_bHxLWWnm0_0(.din(n724),.dout(w_dff_B_bHxLWWnm0_0),.clk(gclk));
	jdff dff_A_PdTwVXbF9_1(.dout(w_G311_1[1]),.din(w_dff_A_PdTwVXbF9_1),.clk(gclk));
	jdff dff_B_lMcfsCfC6_3(.din(G311),.dout(w_dff_B_lMcfsCfC6_3),.clk(gclk));
	jdff dff_B_a15zM2mw9_3(.din(w_dff_B_lMcfsCfC6_3),.dout(w_dff_B_a15zM2mw9_3),.clk(gclk));
	jdff dff_B_VxTUBMna6_3(.din(w_dff_B_a15zM2mw9_3),.dout(w_dff_B_VxTUBMna6_3),.clk(gclk));
	jdff dff_B_XrhrrlvU0_1(.din(n710),.dout(w_dff_B_XrhrrlvU0_1),.clk(gclk));
	jdff dff_B_TVNJnW056_1(.din(n712),.dout(w_dff_B_TVNJnW056_1),.clk(gclk));
	jdff dff_B_r2gcMh6c5_1(.din(n715),.dout(w_dff_B_r2gcMh6c5_1),.clk(gclk));
	jdff dff_B_jVLjZUPy4_1(.din(n716),.dout(w_dff_B_jVLjZUPy4_1),.clk(gclk));
	jdff dff_A_7umLYpXk7_1(.dout(w_G68_3[1]),.din(w_dff_A_7umLYpXk7_1),.clk(gclk));
	jdff dff_A_jxYs8qcu1_1(.dout(w_dff_A_7umLYpXk7_1),.din(w_dff_A_jxYs8qcu1_1),.clk(gclk));
	jdff dff_A_A7uLTU6D5_1(.dout(w_dff_A_jxYs8qcu1_1),.din(w_dff_A_A7uLTU6D5_1),.clk(gclk));
	jdff dff_A_RZGU9K3y6_2(.dout(w_G68_3[2]),.din(w_dff_A_RZGU9K3y6_2),.clk(gclk));
	jdff dff_A_QAexC1sc5_2(.dout(w_dff_A_RZGU9K3y6_2),.din(w_dff_A_QAexC1sc5_2),.clk(gclk));
	jdff dff_A_fg08Ldde0_1(.dout(w_G137_1[1]),.din(w_dff_A_fg08Ldde0_1),.clk(gclk));
	jdff dff_B_3B131pBc4_3(.din(G137),.dout(w_dff_B_3B131pBc4_3),.clk(gclk));
	jdff dff_B_QIrx4NMT7_3(.din(w_dff_B_3B131pBc4_3),.dout(w_dff_B_QIrx4NMT7_3),.clk(gclk));
	jdff dff_B_ob9irtai4_3(.din(w_dff_B_QIrx4NMT7_3),.dout(w_dff_B_ob9irtai4_3),.clk(gclk));
	jdff dff_B_1aarbTzk5_3(.din(G143),.dout(w_dff_B_1aarbTzk5_3),.clk(gclk));
	jdff dff_B_bPHmTA1B5_3(.din(w_dff_B_1aarbTzk5_3),.dout(w_dff_B_bPHmTA1B5_3),.clk(gclk));
	jdff dff_B_OJom1FYt1_3(.din(w_dff_B_bPHmTA1B5_3),.dout(w_dff_B_OJom1FYt1_3),.clk(gclk));
	jdff dff_A_1jvSdNCV3_0(.dout(w_G159_3[0]),.din(w_dff_A_1jvSdNCV3_0),.clk(gclk));
	jdff dff_A_qnf9fads5_1(.dout(w_G159_3[1]),.din(w_dff_A_qnf9fads5_1),.clk(gclk));
	jdff dff_A_a7wtfoCu3_1(.dout(w_dff_A_qnf9fads5_1),.din(w_dff_A_a7wtfoCu3_1),.clk(gclk));
	jdff dff_A_Tu0gHDuX6_0(.dout(w_G159_0[0]),.din(w_dff_A_Tu0gHDuX6_0),.clk(gclk));
	jdff dff_A_NYxeNxQl8_0(.dout(w_dff_A_Tu0gHDuX6_0),.din(w_dff_A_NYxeNxQl8_0),.clk(gclk));
	jdff dff_A_cIHiKiZJ6_1(.dout(w_G159_0[1]),.din(w_dff_A_cIHiKiZJ6_1),.clk(gclk));
	jdff dff_B_10MjFtWH4_3(.din(G159),.dout(w_dff_B_10MjFtWH4_3),.clk(gclk));
	jdff dff_B_FaIakyj15_3(.din(w_dff_B_10MjFtWH4_3),.dout(w_dff_B_FaIakyj15_3),.clk(gclk));
	jdff dff_A_S6zJZXWQ4_1(.dout(w_G190_2[1]),.din(w_dff_A_S6zJZXWQ4_1),.clk(gclk));
	jdff dff_A_5WXIHceh4_1(.dout(w_dff_A_S6zJZXWQ4_1),.din(w_dff_A_5WXIHceh4_1),.clk(gclk));
	jdff dff_A_voKTqiQL6_1(.dout(w_dff_A_5WXIHceh4_1),.din(w_dff_A_voKTqiQL6_1),.clk(gclk));
	jdff dff_A_xVhRKMLI4_1(.dout(w_dff_A_voKTqiQL6_1),.din(w_dff_A_xVhRKMLI4_1),.clk(gclk));
	jdff dff_A_bXRGpFUT9_1(.dout(w_dff_A_xVhRKMLI4_1),.din(w_dff_A_bXRGpFUT9_1),.clk(gclk));
	jdff dff_A_ZQoEcb4V4_2(.dout(w_G190_2[2]),.din(w_dff_A_ZQoEcb4V4_2),.clk(gclk));
	jdff dff_A_1O6QwAK35_2(.dout(w_dff_A_ZQoEcb4V4_2),.din(w_dff_A_1O6QwAK35_2),.clk(gclk));
	jdff dff_A_voqPKDHg0_2(.dout(w_dff_A_1O6QwAK35_2),.din(w_dff_A_voqPKDHg0_2),.clk(gclk));
	jdff dff_A_qJaP0EbY2_2(.dout(w_dff_A_voqPKDHg0_2),.din(w_dff_A_qJaP0EbY2_2),.clk(gclk));
	jdff dff_A_ZwW0hqYD3_2(.dout(w_dff_A_qJaP0EbY2_2),.din(w_dff_A_ZwW0hqYD3_2),.clk(gclk));
	jdff dff_A_Y6d7z2k86_0(.dout(w_G50_3[0]),.din(w_dff_A_Y6d7z2k86_0),.clk(gclk));
	jdff dff_A_VSlrG3Dt9_0(.dout(w_dff_A_Y6d7z2k86_0),.din(w_dff_A_VSlrG3Dt9_0),.clk(gclk));
	jdff dff_A_q4g8PyAu0_0(.dout(w_dff_A_VSlrG3Dt9_0),.din(w_dff_A_q4g8PyAu0_0),.clk(gclk));
	jdff dff_A_Lcjr7Jkd0_2(.dout(w_G50_3[2]),.din(w_dff_A_Lcjr7Jkd0_2),.clk(gclk));
	jdff dff_A_PQWol2Sk5_2(.dout(w_dff_A_Lcjr7Jkd0_2),.din(w_dff_A_PQWol2Sk5_2),.clk(gclk));
	jdff dff_A_E87Knj2C7_2(.dout(w_dff_A_PQWol2Sk5_2),.din(w_dff_A_E87Knj2C7_2),.clk(gclk));
	jdff dff_A_0z4pOVe93_2(.dout(w_dff_A_E87Knj2C7_2),.din(w_dff_A_0z4pOVe93_2),.clk(gclk));
	jdff dff_A_E8BBP3RC2_1(.dout(w_G50_0[1]),.din(w_dff_A_E8BBP3RC2_1),.clk(gclk));
	jdff dff_A_YDRcNMc83_1(.dout(w_dff_A_E8BBP3RC2_1),.din(w_dff_A_YDRcNMc83_1),.clk(gclk));
	jdff dff_A_YtGq8GRF4_1(.dout(w_dff_A_YDRcNMc83_1),.din(w_dff_A_YtGq8GRF4_1),.clk(gclk));
	jdff dff_A_t519heTb5_0(.dout(w_G33_6[0]),.din(w_dff_A_t519heTb5_0),.clk(gclk));
	jdff dff_A_pQn8Bwgt4_0(.dout(w_dff_A_t519heTb5_0),.din(w_dff_A_pQn8Bwgt4_0),.clk(gclk));
	jdff dff_A_sftDko8u2_0(.dout(w_dff_A_pQn8Bwgt4_0),.din(w_dff_A_sftDko8u2_0),.clk(gclk));
	jdff dff_A_c0tZk3tN5_0(.dout(w_dff_A_sftDko8u2_0),.din(w_dff_A_c0tZk3tN5_0),.clk(gclk));
	jdff dff_A_UIfhTpSR6_1(.dout(w_G33_6[1]),.din(w_dff_A_UIfhTpSR6_1),.clk(gclk));
	jdff dff_A_Os20HUNC9_1(.dout(w_dff_A_UIfhTpSR6_1),.din(w_dff_A_Os20HUNC9_1),.clk(gclk));
	jdff dff_A_nE77gkUE2_1(.dout(w_G33_1[1]),.din(w_dff_A_nE77gkUE2_1),.clk(gclk));
	jdff dff_A_kTjxzvWT2_1(.dout(w_dff_A_nE77gkUE2_1),.din(w_dff_A_kTjxzvWT2_1),.clk(gclk));
	jdff dff_A_BgoFfZ3G5_1(.dout(w_dff_A_kTjxzvWT2_1),.din(w_dff_A_BgoFfZ3G5_1),.clk(gclk));
	jdff dff_B_YOTbRa345_1(.din(n706),.dout(w_dff_B_YOTbRa345_1),.clk(gclk));
	jdff dff_B_VXotR1C14_0(.din(n708),.dout(w_dff_B_VXotR1C14_0),.clk(gclk));
	jdff dff_A_sZBHAwzC5_0(.dout(w_G150_3[0]),.din(w_dff_A_sZBHAwzC5_0),.clk(gclk));
	jdff dff_A_OjuoUKn81_0(.dout(w_dff_A_sZBHAwzC5_0),.din(w_dff_A_OjuoUKn81_0),.clk(gclk));
	jdff dff_A_6kKoFWxY3_0(.dout(w_dff_A_OjuoUKn81_0),.din(w_dff_A_6kKoFWxY3_0),.clk(gclk));
	jdff dff_A_6QzVYnv16_0(.dout(w_G150_0[0]),.din(w_dff_A_6QzVYnv16_0),.clk(gclk));
	jdff dff_A_WpFUIipS7_0(.dout(w_dff_A_6QzVYnv16_0),.din(w_dff_A_WpFUIipS7_0),.clk(gclk));
	jdff dff_A_XapG0G1E1_0(.dout(w_dff_A_WpFUIipS7_0),.din(w_dff_A_XapG0G1E1_0),.clk(gclk));
	jdff dff_A_k8AR201x1_1(.dout(w_G150_0[1]),.din(w_dff_A_k8AR201x1_1),.clk(gclk));
	jdff dff_A_hjzNrcIA2_1(.dout(w_dff_A_k8AR201x1_1),.din(w_dff_A_hjzNrcIA2_1),.clk(gclk));
	jdff dff_A_3IWXGl4Q0_1(.dout(w_dff_A_hjzNrcIA2_1),.din(w_dff_A_3IWXGl4Q0_1),.clk(gclk));
	jdff dff_A_B9U87A7P4_0(.dout(w_G58_3[0]),.din(w_dff_A_B9U87A7P4_0),.clk(gclk));
	jdff dff_A_8HWxLwAr6_1(.dout(w_G58_3[1]),.din(w_dff_A_8HWxLwAr6_1),.clk(gclk));
	jdff dff_A_jajZH1VY4_1(.dout(w_n615_0[1]),.din(w_dff_A_jajZH1VY4_1),.clk(gclk));
	jdff dff_A_cgO3RsdM6_1(.dout(w_G200_2[1]),.din(w_dff_A_cgO3RsdM6_1),.clk(gclk));
	jdff dff_A_jgi2bvqi1_1(.dout(w_dff_A_cgO3RsdM6_1),.din(w_dff_A_jgi2bvqi1_1),.clk(gclk));
	jdff dff_A_NrGcdwvs9_1(.dout(w_dff_A_jgi2bvqi1_1),.din(w_dff_A_NrGcdwvs9_1),.clk(gclk));
	jdff dff_A_rbiAdqSD1_1(.dout(w_dff_A_NrGcdwvs9_1),.din(w_dff_A_rbiAdqSD1_1),.clk(gclk));
	jdff dff_A_Bv9YZrCL5_1(.dout(w_dff_A_rbiAdqSD1_1),.din(w_dff_A_Bv9YZrCL5_1),.clk(gclk));
	jdff dff_A_SVEJQEdk3_1(.dout(w_dff_A_Bv9YZrCL5_1),.din(w_dff_A_SVEJQEdk3_1),.clk(gclk));
	jdff dff_A_ockTjTGj2_1(.dout(w_dff_A_SVEJQEdk3_1),.din(w_dff_A_ockTjTGj2_1),.clk(gclk));
	jdff dff_A_j1AoV3UV3_2(.dout(w_G200_2[2]),.din(w_dff_A_j1AoV3UV3_2),.clk(gclk));
	jdff dff_A_PsH6dYKB1_2(.dout(w_dff_A_j1AoV3UV3_2),.din(w_dff_A_PsH6dYKB1_2),.clk(gclk));
	jdff dff_A_NNb2mDc57_2(.dout(w_dff_A_PsH6dYKB1_2),.din(w_dff_A_NNb2mDc57_2),.clk(gclk));
	jdff dff_A_LEOZPeAq6_2(.dout(w_dff_A_NNb2mDc57_2),.din(w_dff_A_LEOZPeAq6_2),.clk(gclk));
	jdff dff_A_RLuNULWX6_2(.dout(w_dff_A_LEOZPeAq6_2),.din(w_dff_A_RLuNULWX6_2),.clk(gclk));
	jdff dff_A_hnkDfjQ26_2(.dout(w_dff_A_RLuNULWX6_2),.din(w_dff_A_hnkDfjQ26_2),.clk(gclk));
	jdff dff_A_cCghVtay5_2(.dout(w_dff_A_hnkDfjQ26_2),.din(w_dff_A_cCghVtay5_2),.clk(gclk));
	jdff dff_A_4V9nTFmm2_0(.dout(w_n619_0[0]),.din(w_dff_A_4V9nTFmm2_0),.clk(gclk));
	jdff dff_A_BmjXFYCM9_0(.dout(w_n407_1[0]),.din(w_dff_A_BmjXFYCM9_0),.clk(gclk));
	jdff dff_A_zyh5SjHl5_1(.dout(w_n407_1[1]),.din(w_dff_A_zyh5SjHl5_1),.clk(gclk));
	jdff dff_A_SoJMaa6U8_1(.dout(w_dff_A_zyh5SjHl5_1),.din(w_dff_A_SoJMaa6U8_1),.clk(gclk));
	jdff dff_A_UqmQbHpi3_1(.dout(w_G132_1[1]),.din(w_dff_A_UqmQbHpi3_1),.clk(gclk));
	jdff dff_B_hcZHqHtM7_3(.din(G132),.dout(w_dff_B_hcZHqHtM7_3),.clk(gclk));
	jdff dff_B_pBdD8D9U3_3(.din(w_dff_B_hcZHqHtM7_3),.dout(w_dff_B_pBdD8D9U3_3),.clk(gclk));
	jdff dff_B_ZMOIlzt87_3(.din(w_dff_B_pBdD8D9U3_3),.dout(w_dff_B_ZMOIlzt87_3),.clk(gclk));
	jdff dff_A_rz8ZnS6y4_0(.dout(w_n612_3[0]),.din(w_dff_A_rz8ZnS6y4_0),.clk(gclk));
	jdff dff_A_3WnZy8Of3_0(.dout(w_dff_A_rz8ZnS6y4_0),.din(w_dff_A_3WnZy8Of3_0),.clk(gclk));
	jdff dff_A_EqDyQK220_0(.dout(w_dff_A_3WnZy8Of3_0),.din(w_dff_A_EqDyQK220_0),.clk(gclk));
	jdff dff_A_XyPl7Lk52_0(.dout(w_dff_A_EqDyQK220_0),.din(w_dff_A_XyPl7Lk52_0),.clk(gclk));
	jdff dff_A_qpkrdL6F0_0(.dout(w_dff_A_XyPl7Lk52_0),.din(w_dff_A_qpkrdL6F0_0),.clk(gclk));
	jdff dff_A_aJLsqmqe2_0(.dout(w_dff_A_qpkrdL6F0_0),.din(w_dff_A_aJLsqmqe2_0),.clk(gclk));
	jdff dff_A_2IN7JSSE6_0(.dout(w_dff_A_aJLsqmqe2_0),.din(w_dff_A_2IN7JSSE6_0),.clk(gclk));
	jdff dff_A_milrLsVw7_0(.dout(w_dff_A_2IN7JSSE6_0),.din(w_dff_A_milrLsVw7_0),.clk(gclk));
	jdff dff_A_eDV0uxhS1_0(.dout(w_dff_A_milrLsVw7_0),.din(w_dff_A_eDV0uxhS1_0),.clk(gclk));
	jdff dff_A_94mwUmcO2_2(.dout(w_n612_3[2]),.din(w_dff_A_94mwUmcO2_2),.clk(gclk));
	jdff dff_A_0IwzuOTi7_2(.dout(w_dff_A_94mwUmcO2_2),.din(w_dff_A_0IwzuOTi7_2),.clk(gclk));
	jdff dff_A_Isvsff5S9_2(.dout(w_dff_A_0IwzuOTi7_2),.din(w_dff_A_Isvsff5S9_2),.clk(gclk));
	jdff dff_A_cxIVGy278_2(.dout(w_dff_A_Isvsff5S9_2),.din(w_dff_A_cxIVGy278_2),.clk(gclk));
	jdff dff_A_PltvLy5v7_2(.dout(w_dff_A_cxIVGy278_2),.din(w_dff_A_PltvLy5v7_2),.clk(gclk));
	jdff dff_A_bLHjKvDv5_2(.dout(w_dff_A_PltvLy5v7_2),.din(w_dff_A_bLHjKvDv5_2),.clk(gclk));
	jdff dff_A_YfFfKuRT3_2(.dout(w_dff_A_bLHjKvDv5_2),.din(w_dff_A_YfFfKuRT3_2),.clk(gclk));
	jdff dff_A_ZCgrvjX68_2(.dout(w_dff_A_YfFfKuRT3_2),.din(w_dff_A_ZCgrvjX68_2),.clk(gclk));
	jdff dff_A_DNgoaVjB0_2(.dout(w_dff_A_ZCgrvjX68_2),.din(w_dff_A_DNgoaVjB0_2),.clk(gclk));
	jdff dff_A_AleqX0qi5_1(.dout(w_n612_0[1]),.din(w_dff_A_AleqX0qi5_1),.clk(gclk));
	jdff dff_A_0ODAtrUi0_1(.dout(w_dff_A_AleqX0qi5_1),.din(w_dff_A_0ODAtrUi0_1),.clk(gclk));
	jdff dff_A_ILahda5L6_1(.dout(w_dff_A_0ODAtrUi0_1),.din(w_dff_A_ILahda5L6_1),.clk(gclk));
	jdff dff_A_x1atrqor5_1(.dout(w_dff_A_ILahda5L6_1),.din(w_dff_A_x1atrqor5_1),.clk(gclk));
	jdff dff_A_PoO6PUAm4_1(.dout(w_dff_A_x1atrqor5_1),.din(w_dff_A_PoO6PUAm4_1),.clk(gclk));
	jdff dff_A_MXYQ7IB02_1(.dout(w_dff_A_PoO6PUAm4_1),.din(w_dff_A_MXYQ7IB02_1),.clk(gclk));
	jdff dff_A_KIRTliAh7_1(.dout(w_dff_A_MXYQ7IB02_1),.din(w_dff_A_KIRTliAh7_1),.clk(gclk));
	jdff dff_A_YM0Ge1Vw3_1(.dout(w_n146_1[1]),.din(w_dff_A_YM0Ge1Vw3_1),.clk(gclk));
	jdff dff_A_QQY4p0rR0_1(.dout(w_dff_A_YM0Ge1Vw3_1),.din(w_dff_A_QQY4p0rR0_1),.clk(gclk));
	jdff dff_A_euVF13K51_1(.dout(w_dff_A_QQY4p0rR0_1),.din(w_dff_A_euVF13K51_1),.clk(gclk));
	jdff dff_A_krnNoCNg3_1(.dout(w_dff_A_euVF13K51_1),.din(w_dff_A_krnNoCNg3_1),.clk(gclk));
	jdff dff_A_lUaj8Hsi0_1(.dout(w_dff_A_krnNoCNg3_1),.din(w_dff_A_lUaj8Hsi0_1),.clk(gclk));
	jdff dff_A_pmUtW7ki4_1(.dout(w_dff_A_lUaj8Hsi0_1),.din(w_dff_A_pmUtW7ki4_1),.clk(gclk));
	jdff dff_A_ZyVloKti1_2(.dout(w_n146_1[2]),.din(w_dff_A_ZyVloKti1_2),.clk(gclk));
	jdff dff_A_6HQUVwQJ4_2(.dout(w_dff_A_ZyVloKti1_2),.din(w_dff_A_6HQUVwQJ4_2),.clk(gclk));
	jdff dff_A_fnaKOyxR0_2(.dout(w_dff_A_6HQUVwQJ4_2),.din(w_dff_A_fnaKOyxR0_2),.clk(gclk));
	jdff dff_A_EAZ32BHi9_2(.dout(w_dff_A_fnaKOyxR0_2),.din(w_dff_A_EAZ32BHi9_2),.clk(gclk));
	jdff dff_A_bK1TnP9p4_2(.dout(w_dff_A_EAZ32BHi9_2),.din(w_dff_A_bK1TnP9p4_2),.clk(gclk));
	jdff dff_A_7hze8iR17_2(.dout(w_dff_A_bK1TnP9p4_2),.din(w_dff_A_7hze8iR17_2),.clk(gclk));
	jdff dff_A_qCgzmTEy5_0(.dout(w_n425_1[0]),.din(w_dff_A_qCgzmTEy5_0),.clk(gclk));
	jdff dff_A_hmWkYl082_0(.dout(w_dff_A_qCgzmTEy5_0),.din(w_dff_A_hmWkYl082_0),.clk(gclk));
	jdff dff_A_ke3cuQ8i2_0(.dout(w_dff_A_hmWkYl082_0),.din(w_dff_A_ke3cuQ8i2_0),.clk(gclk));
	jdff dff_A_oQQHS6Mo0_0(.dout(w_dff_A_ke3cuQ8i2_0),.din(w_dff_A_oQQHS6Mo0_0),.clk(gclk));
	jdff dff_A_3o3Aga818_0(.dout(w_dff_A_oQQHS6Mo0_0),.din(w_dff_A_3o3Aga818_0),.clk(gclk));
	jdff dff_A_4PtGJqYM5_0(.dout(w_dff_A_3o3Aga818_0),.din(w_dff_A_4PtGJqYM5_0),.clk(gclk));
	jdff dff_A_S6x8R5Mw2_0(.dout(w_dff_A_4PtGJqYM5_0),.din(w_dff_A_S6x8R5Mw2_0),.clk(gclk));
	jdff dff_A_Gn1AnE2P9_0(.dout(w_dff_A_S6x8R5Mw2_0),.din(w_dff_A_Gn1AnE2P9_0),.clk(gclk));
	jdff dff_A_pbjlvNlT9_0(.dout(w_dff_A_Gn1AnE2P9_0),.din(w_dff_A_pbjlvNlT9_0),.clk(gclk));
	jdff dff_A_J6QaOLpY5_0(.dout(w_dff_A_pbjlvNlT9_0),.din(w_dff_A_J6QaOLpY5_0),.clk(gclk));
	jdff dff_A_it7GQ7Dp9_0(.dout(w_dff_A_J6QaOLpY5_0),.din(w_dff_A_it7GQ7Dp9_0),.clk(gclk));
	jdff dff_A_Y9PeBElv4_0(.dout(w_dff_A_it7GQ7Dp9_0),.din(w_dff_A_Y9PeBElv4_0),.clk(gclk));
	jdff dff_A_8ee8hWvj7_0(.dout(w_dff_A_Y9PeBElv4_0),.din(w_dff_A_8ee8hWvj7_0),.clk(gclk));
	jdff dff_A_eDriXEU77_1(.dout(w_n425_1[1]),.din(w_dff_A_eDriXEU77_1),.clk(gclk));
	jdff dff_A_vbppFX2z4_1(.dout(w_dff_A_eDriXEU77_1),.din(w_dff_A_vbppFX2z4_1),.clk(gclk));
	jdff dff_A_r9m11Sp88_1(.dout(w_dff_A_vbppFX2z4_1),.din(w_dff_A_r9m11Sp88_1),.clk(gclk));
	jdff dff_A_S2lH40NS3_1(.dout(w_dff_A_r9m11Sp88_1),.din(w_dff_A_S2lH40NS3_1),.clk(gclk));
	jdff dff_A_hwFI4iZB9_1(.dout(w_dff_A_S2lH40NS3_1),.din(w_dff_A_hwFI4iZB9_1),.clk(gclk));
	jdff dff_A_lNkq2tnW6_1(.dout(w_dff_A_hwFI4iZB9_1),.din(w_dff_A_lNkq2tnW6_1),.clk(gclk));
	jdff dff_A_17g9O5Q45_1(.dout(w_dff_A_lNkq2tnW6_1),.din(w_dff_A_17g9O5Q45_1),.clk(gclk));
	jdff dff_A_BHDPSEJu9_1(.dout(w_dff_A_17g9O5Q45_1),.din(w_dff_A_BHDPSEJu9_1),.clk(gclk));
	jdff dff_A_es2IyWpY0_1(.dout(w_dff_A_BHDPSEJu9_1),.din(w_dff_A_es2IyWpY0_1),.clk(gclk));
	jdff dff_A_e1hrWvYU6_1(.dout(w_dff_A_es2IyWpY0_1),.din(w_dff_A_e1hrWvYU6_1),.clk(gclk));
	jdff dff_A_VZd0gpUa7_1(.dout(w_dff_A_e1hrWvYU6_1),.din(w_dff_A_VZd0gpUa7_1),.clk(gclk));
	jdff dff_A_epIckd794_1(.dout(w_dff_A_VZd0gpUa7_1),.din(w_dff_A_epIckd794_1),.clk(gclk));
	jdff dff_A_rmQ2P6ob1_1(.dout(w_dff_A_epIckd794_1),.din(w_dff_A_rmQ2P6ob1_1),.clk(gclk));
	jdff dff_A_4rI3Hm1b7_1(.dout(w_n425_0[1]),.din(w_dff_A_4rI3Hm1b7_1),.clk(gclk));
	jdff dff_A_JcjRvWF04_1(.dout(w_dff_A_4rI3Hm1b7_1),.din(w_dff_A_JcjRvWF04_1),.clk(gclk));
	jdff dff_A_Sk17eZjh8_1(.dout(w_dff_A_JcjRvWF04_1),.din(w_dff_A_Sk17eZjh8_1),.clk(gclk));
	jdff dff_A_Z5GJ55JZ7_1(.dout(w_dff_A_Sk17eZjh8_1),.din(w_dff_A_Z5GJ55JZ7_1),.clk(gclk));
	jdff dff_A_Jlmq51Zr9_1(.dout(w_dff_A_Z5GJ55JZ7_1),.din(w_dff_A_Jlmq51Zr9_1),.clk(gclk));
	jdff dff_A_y4ktkX414_1(.dout(w_dff_A_Jlmq51Zr9_1),.din(w_dff_A_y4ktkX414_1),.clk(gclk));
	jdff dff_A_zP91gkby3_1(.dout(w_dff_A_y4ktkX414_1),.din(w_dff_A_zP91gkby3_1),.clk(gclk));
	jdff dff_A_gn9FCwl94_1(.dout(w_dff_A_zP91gkby3_1),.din(w_dff_A_gn9FCwl94_1),.clk(gclk));
	jdff dff_A_EU8P0IAU4_1(.dout(w_dff_A_gn9FCwl94_1),.din(w_dff_A_EU8P0IAU4_1),.clk(gclk));
	jdff dff_A_Z7lBfSnI7_1(.dout(w_dff_A_EU8P0IAU4_1),.din(w_dff_A_Z7lBfSnI7_1),.clk(gclk));
	jdff dff_A_vyM2sOR99_1(.dout(w_dff_A_Z7lBfSnI7_1),.din(w_dff_A_vyM2sOR99_1),.clk(gclk));
	jdff dff_A_Br01DCnm4_1(.dout(w_dff_A_vyM2sOR99_1),.din(w_dff_A_Br01DCnm4_1),.clk(gclk));
	jdff dff_A_fSXR1oKu2_1(.dout(w_dff_A_Br01DCnm4_1),.din(w_dff_A_fSXR1oKu2_1),.clk(gclk));
	jdff dff_A_fqyNz2KY1_2(.dout(w_n425_0[2]),.din(w_dff_A_fqyNz2KY1_2),.clk(gclk));
	jdff dff_A_eD5IR1Xa5_2(.dout(w_dff_A_fqyNz2KY1_2),.din(w_dff_A_eD5IR1Xa5_2),.clk(gclk));
	jdff dff_A_nTNjntaC7_2(.dout(w_dff_A_eD5IR1Xa5_2),.din(w_dff_A_nTNjntaC7_2),.clk(gclk));
	jdff dff_A_1QqJ9wCN0_2(.dout(w_dff_A_nTNjntaC7_2),.din(w_dff_A_1QqJ9wCN0_2),.clk(gclk));
	jdff dff_A_cwOhX6n43_2(.dout(w_dff_A_1QqJ9wCN0_2),.din(w_dff_A_cwOhX6n43_2),.clk(gclk));
	jdff dff_A_BRkAedmK3_2(.dout(w_dff_A_cwOhX6n43_2),.din(w_dff_A_BRkAedmK3_2),.clk(gclk));
	jdff dff_A_oSt0Z7Fn2_2(.dout(w_dff_A_BRkAedmK3_2),.din(w_dff_A_oSt0Z7Fn2_2),.clk(gclk));
	jdff dff_A_GaKWSEUJ3_2(.dout(w_dff_A_oSt0Z7Fn2_2),.din(w_dff_A_GaKWSEUJ3_2),.clk(gclk));
	jdff dff_A_6jzFGnfY0_2(.dout(w_dff_A_GaKWSEUJ3_2),.din(w_dff_A_6jzFGnfY0_2),.clk(gclk));
	jdff dff_A_lxyL6k5x6_2(.dout(w_dff_A_6jzFGnfY0_2),.din(w_dff_A_lxyL6k5x6_2),.clk(gclk));
	jdff dff_A_5WFaK1hc7_2(.dout(w_dff_A_lxyL6k5x6_2),.din(w_dff_A_5WFaK1hc7_2),.clk(gclk));
	jdff dff_A_0qz3eAIP3_2(.dout(w_dff_A_5WFaK1hc7_2),.din(w_dff_A_0qz3eAIP3_2),.clk(gclk));
	jdff dff_A_qItjlHxo7_2(.dout(w_dff_A_0qz3eAIP3_2),.din(w_dff_A_qItjlHxo7_2),.clk(gclk));
	jdff dff_A_2Lxs9L7N3_0(.dout(w_n148_1[0]),.din(w_dff_A_2Lxs9L7N3_0),.clk(gclk));
	jdff dff_A_teYQVboa8_0(.dout(w_dff_A_2Lxs9L7N3_0),.din(w_dff_A_teYQVboa8_0),.clk(gclk));
	jdff dff_A_h56ZK11V3_0(.dout(w_dff_A_teYQVboa8_0),.din(w_dff_A_h56ZK11V3_0),.clk(gclk));
	jdff dff_A_6yVyZMe51_0(.dout(w_dff_A_h56ZK11V3_0),.din(w_dff_A_6yVyZMe51_0),.clk(gclk));
	jdff dff_A_FrwTlVFw6_1(.dout(w_n148_1[1]),.din(w_dff_A_FrwTlVFw6_1),.clk(gclk));
	jdff dff_A_GjQKIh0o2_1(.dout(w_dff_A_FrwTlVFw6_1),.din(w_dff_A_GjQKIh0o2_1),.clk(gclk));
	jdff dff_B_sOUDt0Jw2_0(.din(n701),.dout(w_dff_B_sOUDt0Jw2_0),.clk(gclk));
	jdff dff_A_sEsirQ287_0(.dout(w_n604_1[0]),.din(w_dff_A_sEsirQ287_0),.clk(gclk));
	jdff dff_A_tjhWdLt39_0(.dout(w_dff_A_sEsirQ287_0),.din(w_dff_A_tjhWdLt39_0),.clk(gclk));
	jdff dff_A_wb8Hnplw2_2(.dout(w_n604_1[2]),.din(w_dff_A_wb8Hnplw2_2),.clk(gclk));
	jdff dff_A_jEUckHfx1_2(.dout(w_dff_A_wb8Hnplw2_2),.din(w_dff_A_jEUckHfx1_2),.clk(gclk));
	jdff dff_A_bOcYBU0u4_2(.dout(w_dff_A_jEUckHfx1_2),.din(w_dff_A_bOcYBU0u4_2),.clk(gclk));
	jdff dff_A_ho90xERe3_2(.dout(w_dff_A_bOcYBU0u4_2),.din(w_dff_A_ho90xERe3_2),.clk(gclk));
	jdff dff_A_XAQQnvFH0_2(.dout(w_dff_A_ho90xERe3_2),.din(w_dff_A_XAQQnvFH0_2),.clk(gclk));
	jdff dff_A_5l6bkAPs5_2(.dout(w_dff_A_XAQQnvFH0_2),.din(w_dff_A_5l6bkAPs5_2),.clk(gclk));
	jdff dff_A_LBbokkSq4_2(.dout(w_dff_A_5l6bkAPs5_2),.din(w_dff_A_LBbokkSq4_2),.clk(gclk));
	jdff dff_A_4flnU5zK4_2(.dout(w_dff_A_LBbokkSq4_2),.din(w_dff_A_4flnU5zK4_2),.clk(gclk));
	jdff dff_A_zv0BLC0m7_0(.dout(w_n604_0[0]),.din(w_dff_A_zv0BLC0m7_0),.clk(gclk));
	jdff dff_A_foqsK1iu2_0(.dout(w_dff_A_zv0BLC0m7_0),.din(w_dff_A_foqsK1iu2_0),.clk(gclk));
	jdff dff_A_b2z0fmQw0_2(.dout(w_n604_0[2]),.din(w_dff_A_b2z0fmQw0_2),.clk(gclk));
	jdff dff_A_K3AGBwzM7_2(.dout(w_dff_A_b2z0fmQw0_2),.din(w_dff_A_K3AGBwzM7_2),.clk(gclk));
	jdff dff_A_Qm3iBtMs3_0(.dout(w_n603_2[0]),.din(w_dff_A_Qm3iBtMs3_0),.clk(gclk));
	jdff dff_A_Bqe3jeLH4_0(.dout(w_dff_A_Qm3iBtMs3_0),.din(w_dff_A_Bqe3jeLH4_0),.clk(gclk));
	jdff dff_A_oKToOtMw2_0(.dout(w_dff_A_Bqe3jeLH4_0),.din(w_dff_A_oKToOtMw2_0),.clk(gclk));
	jdff dff_A_rE5M3qzY2_0(.dout(w_dff_A_oKToOtMw2_0),.din(w_dff_A_rE5M3qzY2_0),.clk(gclk));
	jdff dff_A_BtVjkjIy1_0(.dout(w_dff_A_rE5M3qzY2_0),.din(w_dff_A_BtVjkjIy1_0),.clk(gclk));
	jdff dff_A_VkJ1vD6E1_0(.dout(w_dff_A_BtVjkjIy1_0),.din(w_dff_A_VkJ1vD6E1_0),.clk(gclk));
	jdff dff_A_qcHqbGIZ2_0(.dout(w_dff_A_VkJ1vD6E1_0),.din(w_dff_A_qcHqbGIZ2_0),.clk(gclk));
	jdff dff_A_XgjECKGW1_0(.dout(w_dff_A_qcHqbGIZ2_0),.din(w_dff_A_XgjECKGW1_0),.clk(gclk));
	jdff dff_A_NfkWhLiY8_0(.dout(w_dff_A_XgjECKGW1_0),.din(w_dff_A_NfkWhLiY8_0),.clk(gclk));
	jdff dff_A_J59My1ut6_0(.dout(w_dff_A_NfkWhLiY8_0),.din(w_dff_A_J59My1ut6_0),.clk(gclk));
	jdff dff_A_Cc4Z5JpJ0_0(.dout(w_dff_A_J59My1ut6_0),.din(w_dff_A_Cc4Z5JpJ0_0),.clk(gclk));
	jdff dff_A_OHnnts5a2_0(.dout(w_n603_0[0]),.din(w_dff_A_OHnnts5a2_0),.clk(gclk));
	jdff dff_A_cnEcAlP81_0(.dout(w_dff_A_OHnnts5a2_0),.din(w_dff_A_cnEcAlP81_0),.clk(gclk));
	jdff dff_A_5VOD5gPl1_0(.dout(w_dff_A_cnEcAlP81_0),.din(w_dff_A_5VOD5gPl1_0),.clk(gclk));
	jdff dff_A_uUFNsoGC3_0(.dout(w_dff_A_5VOD5gPl1_0),.din(w_dff_A_uUFNsoGC3_0),.clk(gclk));
	jdff dff_A_q04vrTA72_0(.dout(w_dff_A_uUFNsoGC3_0),.din(w_dff_A_q04vrTA72_0),.clk(gclk));
	jdff dff_A_6sHJM5Xy7_0(.dout(w_dff_A_q04vrTA72_0),.din(w_dff_A_6sHJM5Xy7_0),.clk(gclk));
	jdff dff_A_0Vx3tG7G7_0(.dout(w_dff_A_6sHJM5Xy7_0),.din(w_dff_A_0Vx3tG7G7_0),.clk(gclk));
	jdff dff_A_Dpu2HDyE5_0(.dout(w_dff_A_0Vx3tG7G7_0),.din(w_dff_A_Dpu2HDyE5_0),.clk(gclk));
	jdff dff_A_RVW5JvzM4_0(.dout(w_dff_A_Dpu2HDyE5_0),.din(w_dff_A_RVW5JvzM4_0),.clk(gclk));
	jdff dff_A_nRPaJcOi2_0(.dout(w_dff_A_RVW5JvzM4_0),.din(w_dff_A_nRPaJcOi2_0),.clk(gclk));
	jdff dff_A_38n0BuBO0_0(.dout(w_dff_A_nRPaJcOi2_0),.din(w_dff_A_38n0BuBO0_0),.clk(gclk));
	jdff dff_A_5EtYuR3P8_0(.dout(w_dff_A_38n0BuBO0_0),.din(w_dff_A_5EtYuR3P8_0),.clk(gclk));
	jdff dff_A_2Z8Vb7209_0(.dout(w_dff_A_5EtYuR3P8_0),.din(w_dff_A_2Z8Vb7209_0),.clk(gclk));
	jdff dff_A_WuP3LnJy6_0(.dout(w_dff_A_2Z8Vb7209_0),.din(w_dff_A_WuP3LnJy6_0),.clk(gclk));
	jdff dff_A_gLushfnS0_2(.dout(w_n603_0[2]),.din(w_dff_A_gLushfnS0_2),.clk(gclk));
	jdff dff_A_EkWjSkVG5_2(.dout(w_dff_A_gLushfnS0_2),.din(w_dff_A_EkWjSkVG5_2),.clk(gclk));
	jdff dff_A_0FM0OZMY3_2(.dout(w_dff_A_EkWjSkVG5_2),.din(w_dff_A_0FM0OZMY3_2),.clk(gclk));
	jdff dff_A_2ztTpdvS4_2(.dout(w_dff_A_0FM0OZMY3_2),.din(w_dff_A_2ztTpdvS4_2),.clk(gclk));
	jdff dff_A_ABqeBcBg4_2(.dout(w_dff_A_2ztTpdvS4_2),.din(w_dff_A_ABqeBcBg4_2),.clk(gclk));
	jdff dff_A_o4yGNFE28_2(.dout(w_dff_A_ABqeBcBg4_2),.din(w_dff_A_o4yGNFE28_2),.clk(gclk));
	jdff dff_A_3vwKYx7W8_2(.dout(w_dff_A_o4yGNFE28_2),.din(w_dff_A_3vwKYx7W8_2),.clk(gclk));
	jdff dff_A_e5zBkha42_2(.dout(w_dff_A_3vwKYx7W8_2),.din(w_dff_A_e5zBkha42_2),.clk(gclk));
	jdff dff_A_PXx4x6xd0_2(.dout(w_dff_A_e5zBkha42_2),.din(w_dff_A_PXx4x6xd0_2),.clk(gclk));
	jdff dff_A_hJFt0JUq5_2(.dout(w_dff_A_PXx4x6xd0_2),.din(w_dff_A_hJFt0JUq5_2),.clk(gclk));
	jdff dff_A_NOqUuvhp9_2(.dout(w_dff_A_hJFt0JUq5_2),.din(w_dff_A_NOqUuvhp9_2),.clk(gclk));
	jdff dff_A_oK4zSfYn4_2(.dout(w_dff_A_NOqUuvhp9_2),.din(w_dff_A_oK4zSfYn4_2),.clk(gclk));
	jdff dff_A_v2epItUz6_2(.dout(w_dff_A_oK4zSfYn4_2),.din(w_dff_A_v2epItUz6_2),.clk(gclk));
	jdff dff_A_efDEuNxq6_0(.dout(w_n602_0[0]),.din(w_dff_A_efDEuNxq6_0),.clk(gclk));
	jdff dff_A_SbLLWM3N7_0(.dout(w_dff_A_efDEuNxq6_0),.din(w_dff_A_SbLLWM3N7_0),.clk(gclk));
	jdff dff_A_tBKkmNvp4_0(.dout(w_dff_A_SbLLWM3N7_0),.din(w_dff_A_tBKkmNvp4_0),.clk(gclk));
	jdff dff_A_y3PO73Gt2_0(.dout(w_dff_A_tBKkmNvp4_0),.din(w_dff_A_y3PO73Gt2_0),.clk(gclk));
	jdff dff_A_otLYebaF9_0(.dout(w_dff_A_y3PO73Gt2_0),.din(w_dff_A_otLYebaF9_0),.clk(gclk));
	jdff dff_A_jUt24f707_0(.dout(w_dff_A_otLYebaF9_0),.din(w_dff_A_jUt24f707_0),.clk(gclk));
	jdff dff_A_7wzqqj0K4_0(.dout(w_dff_A_jUt24f707_0),.din(w_dff_A_7wzqqj0K4_0),.clk(gclk));
	jdff dff_A_g7s5hUKJ2_0(.dout(w_dff_A_7wzqqj0K4_0),.din(w_dff_A_g7s5hUKJ2_0),.clk(gclk));
	jdff dff_A_HF26pmmT6_0(.dout(w_dff_A_g7s5hUKJ2_0),.din(w_dff_A_HF26pmmT6_0),.clk(gclk));
	jdff dff_A_KIjRKvEF8_0(.dout(w_dff_A_HF26pmmT6_0),.din(w_dff_A_KIjRKvEF8_0),.clk(gclk));
	jdff dff_A_BR7yUBq60_0(.dout(w_dff_A_KIjRKvEF8_0),.din(w_dff_A_BR7yUBq60_0),.clk(gclk));
	jdff dff_A_Msh28AIK4_0(.dout(w_dff_A_BR7yUBq60_0),.din(w_dff_A_Msh28AIK4_0),.clk(gclk));
	jdff dff_A_4H3XaxPj6_0(.dout(w_dff_A_Msh28AIK4_0),.din(w_dff_A_4H3XaxPj6_0),.clk(gclk));
	jdff dff_A_VeR9ydHJ0_0(.dout(w_dff_A_4H3XaxPj6_0),.din(w_dff_A_VeR9ydHJ0_0),.clk(gclk));
	jdff dff_A_DYaQg0vp6_0(.dout(w_dff_A_VeR9ydHJ0_0),.din(w_dff_A_DYaQg0vp6_0),.clk(gclk));
	jdff dff_A_Tlt9Iy7U2_0(.dout(w_dff_A_DYaQg0vp6_0),.din(w_dff_A_Tlt9Iy7U2_0),.clk(gclk));
	jdff dff_A_4dWGbo2M2_0(.dout(w_dff_A_Tlt9Iy7U2_0),.din(w_dff_A_4dWGbo2M2_0),.clk(gclk));
	jdff dff_A_uVqKDdK71_0(.dout(w_n592_0[0]),.din(w_dff_A_uVqKDdK71_0),.clk(gclk));
	jdff dff_A_NIIAfPAZ6_0(.dout(w_dff_A_uVqKDdK71_0),.din(w_dff_A_NIIAfPAZ6_0),.clk(gclk));
	jdff dff_A_FtjmGpGm0_0(.dout(w_dff_A_NIIAfPAZ6_0),.din(w_dff_A_FtjmGpGm0_0),.clk(gclk));
	jdff dff_A_u6fPMMaP3_0(.dout(w_dff_A_FtjmGpGm0_0),.din(w_dff_A_u6fPMMaP3_0),.clk(gclk));
	jdff dff_A_FVLSn8r61_0(.dout(w_dff_A_u6fPMMaP3_0),.din(w_dff_A_FVLSn8r61_0),.clk(gclk));
	jdff dff_A_QFC8lswS0_0(.dout(w_dff_A_FVLSn8r61_0),.din(w_dff_A_QFC8lswS0_0),.clk(gclk));
	jdff dff_A_dbpOmaep7_0(.dout(w_dff_A_QFC8lswS0_0),.din(w_dff_A_dbpOmaep7_0),.clk(gclk));
	jdff dff_A_7yC2WvL09_0(.dout(w_dff_A_dbpOmaep7_0),.din(w_dff_A_7yC2WvL09_0),.clk(gclk));
	jdff dff_A_NKSqx6L97_0(.dout(w_dff_A_7yC2WvL09_0),.din(w_dff_A_NKSqx6L97_0),.clk(gclk));
	jdff dff_A_h4aSon9b3_0(.dout(w_dff_A_NKSqx6L97_0),.din(w_dff_A_h4aSon9b3_0),.clk(gclk));
	jdff dff_A_26u5r4nr6_0(.dout(w_dff_A_h4aSon9b3_0),.din(w_dff_A_26u5r4nr6_0),.clk(gclk));
	jdff dff_A_KUQs97An9_0(.dout(w_dff_A_26u5r4nr6_0),.din(w_dff_A_KUQs97An9_0),.clk(gclk));
	jdff dff_A_sgipNb9P9_0(.dout(w_dff_A_KUQs97An9_0),.din(w_dff_A_sgipNb9P9_0),.clk(gclk));
	jdff dff_A_wb61tip46_2(.dout(w_n592_0[2]),.din(w_dff_A_wb61tip46_2),.clk(gclk));
	jdff dff_A_eAITEikv4_2(.dout(w_dff_A_wb61tip46_2),.din(w_dff_A_eAITEikv4_2),.clk(gclk));
	jdff dff_A_JILv7yJU2_2(.dout(w_dff_A_eAITEikv4_2),.din(w_dff_A_JILv7yJU2_2),.clk(gclk));
	jdff dff_A_lyF7RBDh0_2(.dout(w_dff_A_JILv7yJU2_2),.din(w_dff_A_lyF7RBDh0_2),.clk(gclk));
	jdff dff_A_FIvS8d8q9_2(.dout(w_dff_A_lyF7RBDh0_2),.din(w_dff_A_FIvS8d8q9_2),.clk(gclk));
	jdff dff_A_M10eiDHh9_2(.dout(w_dff_A_FIvS8d8q9_2),.din(w_dff_A_M10eiDHh9_2),.clk(gclk));
	jdff dff_A_lNKpBkY69_2(.dout(w_dff_A_M10eiDHh9_2),.din(w_dff_A_lNKpBkY69_2),.clk(gclk));
	jdff dff_A_wNh1CPYe6_2(.dout(w_dff_A_lNKpBkY69_2),.din(w_dff_A_wNh1CPYe6_2),.clk(gclk));
	jdff dff_A_eWsVhYOj0_2(.dout(w_dff_A_wNh1CPYe6_2),.din(w_dff_A_eWsVhYOj0_2),.clk(gclk));
	jdff dff_A_Ex1egs7k1_2(.dout(w_dff_A_eWsVhYOj0_2),.din(w_dff_A_Ex1egs7k1_2),.clk(gclk));
	jdff dff_A_e4fD6PVS9_2(.dout(w_dff_A_Ex1egs7k1_2),.din(w_dff_A_e4fD6PVS9_2),.clk(gclk));
	jdff dff_A_wbSx4lJH0_2(.dout(w_dff_A_e4fD6PVS9_2),.din(w_dff_A_wbSx4lJH0_2),.clk(gclk));
	jdff dff_A_Kfs7AARq6_2(.dout(w_dff_A_wbSx4lJH0_2),.din(w_dff_A_Kfs7AARq6_2),.clk(gclk));
	jdff dff_A_RDXHd6ax8_2(.dout(w_dff_A_Kfs7AARq6_2),.din(w_dff_A_RDXHd6ax8_2),.clk(gclk));
	jdff dff_A_PLUdXRwP9_2(.dout(w_dff_A_RDXHd6ax8_2),.din(w_dff_A_PLUdXRwP9_2),.clk(gclk));
	jdff dff_A_u2zHD1e91_2(.dout(w_dff_A_PLUdXRwP9_2),.din(w_dff_A_u2zHD1e91_2),.clk(gclk));
	jdff dff_A_n6nBEFBo6_1(.dout(w_n591_0[1]),.din(w_dff_A_n6nBEFBo6_1),.clk(gclk));
	jdff dff_A_E5pJEshh8_1(.dout(w_dff_A_n6nBEFBo6_1),.din(w_dff_A_E5pJEshh8_1),.clk(gclk));
	jdff dff_A_MLM49nvu0_1(.dout(w_dff_A_E5pJEshh8_1),.din(w_dff_A_MLM49nvu0_1),.clk(gclk));
	jdff dff_A_KAKvmEud6_1(.dout(w_dff_A_MLM49nvu0_1),.din(w_dff_A_KAKvmEud6_1),.clk(gclk));
	jdff dff_A_UmJBnRF14_1(.dout(w_dff_A_KAKvmEud6_1),.din(w_dff_A_UmJBnRF14_1),.clk(gclk));
	jdff dff_A_q1cvYpYO2_1(.dout(w_dff_A_UmJBnRF14_1),.din(w_dff_A_q1cvYpYO2_1),.clk(gclk));
	jdff dff_A_9hmZZOMP7_1(.dout(w_dff_A_q1cvYpYO2_1),.din(w_dff_A_9hmZZOMP7_1),.clk(gclk));
	jdff dff_A_T3VMcTWS5_1(.dout(w_dff_A_9hmZZOMP7_1),.din(w_dff_A_T3VMcTWS5_1),.clk(gclk));
	jdff dff_A_0DJNY8V99_1(.dout(w_dff_A_T3VMcTWS5_1),.din(w_dff_A_0DJNY8V99_1),.clk(gclk));
	jdff dff_A_0di6ejzZ1_1(.dout(w_dff_A_0DJNY8V99_1),.din(w_dff_A_0di6ejzZ1_1),.clk(gclk));
	jdff dff_A_Q6Dq8Ah13_1(.dout(w_dff_A_0di6ejzZ1_1),.din(w_dff_A_Q6Dq8Ah13_1),.clk(gclk));
	jdff dff_A_RXvEj56w3_1(.dout(w_dff_A_Q6Dq8Ah13_1),.din(w_dff_A_RXvEj56w3_1),.clk(gclk));
	jdff dff_A_tHQQdhbh2_1(.dout(w_dff_A_RXvEj56w3_1),.din(w_dff_A_tHQQdhbh2_1),.clk(gclk));
	jdff dff_A_cMUk0oNq2_1(.dout(w_dff_A_tHQQdhbh2_1),.din(w_dff_A_cMUk0oNq2_1),.clk(gclk));
	jdff dff_A_6R3kS48e5_1(.dout(w_dff_A_cMUk0oNq2_1),.din(w_dff_A_6R3kS48e5_1),.clk(gclk));
	jdff dff_A_c5SsrmG99_2(.dout(w_n591_0[2]),.din(w_dff_A_c5SsrmG99_2),.clk(gclk));
	jdff dff_A_EAFlgYlb7_2(.dout(w_dff_A_c5SsrmG99_2),.din(w_dff_A_EAFlgYlb7_2),.clk(gclk));
	jdff dff_A_ZwSopGnD6_2(.dout(w_dff_A_EAFlgYlb7_2),.din(w_dff_A_ZwSopGnD6_2),.clk(gclk));
	jdff dff_A_8r5WNWsq5_2(.dout(w_dff_A_ZwSopGnD6_2),.din(w_dff_A_8r5WNWsq5_2),.clk(gclk));
	jdff dff_A_SRQIDQ7D6_2(.dout(w_dff_A_8r5WNWsq5_2),.din(w_dff_A_SRQIDQ7D6_2),.clk(gclk));
	jdff dff_A_XIXWfR327_2(.dout(w_dff_A_SRQIDQ7D6_2),.din(w_dff_A_XIXWfR327_2),.clk(gclk));
	jdff dff_A_lItuLGzC4_2(.dout(w_dff_A_XIXWfR327_2),.din(w_dff_A_lItuLGzC4_2),.clk(gclk));
	jdff dff_A_ZzE4B1hQ3_2(.dout(w_dff_A_lItuLGzC4_2),.din(w_dff_A_ZzE4B1hQ3_2),.clk(gclk));
	jdff dff_A_RzWSvsP64_2(.dout(w_dff_A_ZzE4B1hQ3_2),.din(w_dff_A_RzWSvsP64_2),.clk(gclk));
	jdff dff_A_8t7XT2I58_2(.dout(w_dff_A_RzWSvsP64_2),.din(w_dff_A_8t7XT2I58_2),.clk(gclk));
	jdff dff_A_Wyu1IZHA3_2(.dout(w_dff_A_8t7XT2I58_2),.din(w_dff_A_Wyu1IZHA3_2),.clk(gclk));
	jdff dff_A_zCFOVLXZ8_2(.dout(w_dff_A_Wyu1IZHA3_2),.din(w_dff_A_zCFOVLXZ8_2),.clk(gclk));
	jdff dff_A_kgQl7vYj7_2(.dout(w_dff_A_zCFOVLXZ8_2),.din(w_dff_A_kgQl7vYj7_2),.clk(gclk));
	jdff dff_A_oIS23WKq9_2(.dout(w_dff_A_kgQl7vYj7_2),.din(w_dff_A_oIS23WKq9_2),.clk(gclk));
	jdff dff_A_tOxrVneJ3_2(.dout(w_dff_A_oIS23WKq9_2),.din(w_dff_A_tOxrVneJ3_2),.clk(gclk));
	jdff dff_A_Et3t0F1f3_2(.dout(w_dff_A_tOxrVneJ3_2),.din(w_dff_A_Et3t0F1f3_2),.clk(gclk));
	jdff dff_A_byAoXEJY4_0(.dout(w_n121_0[0]),.din(w_dff_A_byAoXEJY4_0),.clk(gclk));
	jdff dff_B_jnmeR2JH2_1(.din(n690),.dout(w_dff_B_jnmeR2JH2_1),.clk(gclk));
	jdff dff_A_y0drUesM0_0(.dout(w_n696_1[0]),.din(w_dff_A_y0drUesM0_0),.clk(gclk));
	jdff dff_A_oKWf7lUA3_2(.dout(w_n696_1[2]),.din(w_dff_A_oKWf7lUA3_2),.clk(gclk));
	jdff dff_A_GMUR2CPS4_1(.dout(w_n696_0[1]),.din(w_dff_A_GMUR2CPS4_1),.clk(gclk));
	jdff dff_A_z8LJpB2h8_1(.dout(w_n692_0[1]),.din(w_dff_A_z8LJpB2h8_1),.clk(gclk));
	jdff dff_B_z3m5Avw11_2(.din(n692),.dout(w_dff_B_z3m5Avw11_2),.clk(gclk));
	jdff dff_B_5I69Vif71_1(.din(n406),.dout(w_dff_B_5I69Vif71_1),.clk(gclk));
	jdff dff_B_2IrSLCfN1_1(.din(w_dff_B_5I69Vif71_1),.dout(w_dff_B_2IrSLCfN1_1),.clk(gclk));
	jdff dff_A_3lsDjhPM0_1(.dout(w_n407_0[1]),.din(w_dff_A_3lsDjhPM0_1),.clk(gclk));
	jdff dff_A_zACDLaCd8_1(.dout(w_dff_A_3lsDjhPM0_1),.din(w_dff_A_zACDLaCd8_1),.clk(gclk));
	jdff dff_A_H7rNPwfV6_1(.dout(w_dff_A_zACDLaCd8_1),.din(w_dff_A_H7rNPwfV6_1),.clk(gclk));
	jdff dff_A_KERD0IRv4_1(.dout(w_dff_A_H7rNPwfV6_1),.din(w_dff_A_KERD0IRv4_1),.clk(gclk));
	jdff dff_A_YzTLrI8s4_1(.dout(w_dff_A_KERD0IRv4_1),.din(w_dff_A_YzTLrI8s4_1),.clk(gclk));
	jdff dff_A_UHbBUwz78_1(.dout(w_dff_A_YzTLrI8s4_1),.din(w_dff_A_UHbBUwz78_1),.clk(gclk));
	jdff dff_A_a4r3djru3_2(.dout(w_n407_0[2]),.din(w_dff_A_a4r3djru3_2),.clk(gclk));
	jdff dff_A_qexzSkda6_1(.dout(w_n401_0[1]),.din(w_dff_A_qexzSkda6_1),.clk(gclk));
	jdff dff_B_BY0d8Vvj8_1(.din(n396),.dout(w_dff_B_BY0d8Vvj8_1),.clk(gclk));
	jdff dff_B_RrKfitDe2_1(.din(w_dff_B_BY0d8Vvj8_1),.dout(w_dff_B_RrKfitDe2_1),.clk(gclk));
	jdff dff_B_blmEti2I9_1(.din(n397),.dout(w_dff_B_blmEti2I9_1),.clk(gclk));
	jdff dff_B_5UrRsifg7_1(.din(w_dff_B_blmEti2I9_1),.dout(w_dff_B_5UrRsifg7_1),.clk(gclk));
	jdff dff_B_SftRxwdb3_0(.din(n398),.dout(w_dff_B_SftRxwdb3_0),.clk(gclk));
	jdff dff_B_7bGxVacK4_0(.din(w_dff_B_SftRxwdb3_0),.dout(w_dff_B_7bGxVacK4_0),.clk(gclk));
	jdff dff_A_f247w4bX7_1(.dout(w_n72_0[1]),.din(w_dff_A_f247w4bX7_1),.clk(gclk));
	jdff dff_A_ZekLadoH4_1(.dout(w_dff_A_f247w4bX7_1),.din(w_dff_A_ZekLadoH4_1),.clk(gclk));
	jdff dff_A_Tuc3xxEz9_1(.dout(w_dff_A_ZekLadoH4_1),.din(w_dff_A_Tuc3xxEz9_1),.clk(gclk));
	jdff dff_A_452Wf0t57_2(.dout(w_n72_0[2]),.din(w_dff_A_452Wf0t57_2),.clk(gclk));
	jdff dff_A_b1BQvMIP9_2(.dout(w_dff_A_452Wf0t57_2),.din(w_dff_A_b1BQvMIP9_2),.clk(gclk));
	jdff dff_B_FlaDmVrW3_0(.din(n394),.dout(w_dff_B_FlaDmVrW3_0),.clk(gclk));
	jdff dff_A_Evo67m0p9_0(.dout(w_n112_3[0]),.din(w_dff_A_Evo67m0p9_0),.clk(gclk));
	jdff dff_A_BXlryQIW5_0(.dout(w_dff_A_Evo67m0p9_0),.din(w_dff_A_BXlryQIW5_0),.clk(gclk));
	jdff dff_A_fZIAVK5L5_1(.dout(w_n112_3[1]),.din(w_dff_A_fZIAVK5L5_1),.clk(gclk));
	jdff dff_A_iUA9Ib5T0_1(.dout(w_dff_A_fZIAVK5L5_1),.din(w_dff_A_iUA9Ib5T0_1),.clk(gclk));
	jdff dff_A_2N6qgzwC1_0(.dout(w_G58_4[0]),.din(w_dff_A_2N6qgzwC1_0),.clk(gclk));
	jdff dff_A_12RyQrOQ0_1(.dout(w_G58_4[1]),.din(w_dff_A_12RyQrOQ0_1),.clk(gclk));
	jdff dff_A_iBXOt02u3_0(.dout(w_G58_1[0]),.din(w_dff_A_iBXOt02u3_0),.clk(gclk));
	jdff dff_A_m5tUA2gX7_2(.dout(w_G58_1[2]),.din(w_dff_A_m5tUA2gX7_2),.clk(gclk));
	jdff dff_A_4h93hrzN3_2(.dout(w_dff_A_m5tUA2gX7_2),.din(w_dff_A_4h93hrzN3_2),.clk(gclk));
	jdff dff_A_1oddAwu36_2(.dout(w_dff_A_4h93hrzN3_2),.din(w_dff_A_1oddAwu36_2),.clk(gclk));
	jdff dff_A_m1kh582q3_2(.dout(w_dff_A_1oddAwu36_2),.din(w_dff_A_m1kh582q3_2),.clk(gclk));
	jdff dff_A_O5xTzMGe8_1(.dout(w_G58_0[1]),.din(w_dff_A_O5xTzMGe8_1),.clk(gclk));
	jdff dff_A_u587GSUF0_2(.dout(w_G58_0[2]),.din(w_dff_A_u587GSUF0_2),.clk(gclk));
	jdff dff_A_y5BjkwQk8_2(.dout(w_dff_A_u587GSUF0_2),.din(w_dff_A_y5BjkwQk8_2),.clk(gclk));
	jdff dff_A_5GiiMNAY6_2(.dout(w_dff_A_y5BjkwQk8_2),.din(w_dff_A_5GiiMNAY6_2),.clk(gclk));
	jdff dff_A_oNKs1aL00_1(.dout(w_G20_3[1]),.din(w_dff_A_oNKs1aL00_1),.clk(gclk));
	jdff dff_A_MSnj6Roc5_2(.dout(w_G20_3[2]),.din(w_dff_A_MSnj6Roc5_2),.clk(gclk));
	jdff dff_A_oDxiCE6K5_2(.dout(w_dff_A_MSnj6Roc5_2),.din(w_dff_A_oDxiCE6K5_2),.clk(gclk));
	jdff dff_B_ncTjER867_2(.din(n390),.dout(w_dff_B_ncTjER867_2),.clk(gclk));
	jdff dff_B_UiuHreiG2_2(.din(w_dff_B_ncTjER867_2),.dout(w_dff_B_UiuHreiG2_2),.clk(gclk));
	jdff dff_A_Q0cECAjb6_0(.dout(w_G87_2[0]),.din(w_dff_A_Q0cECAjb6_0),.clk(gclk));
	jdff dff_A_heQ81J368_0(.dout(w_dff_A_Q0cECAjb6_0),.din(w_dff_A_heQ81J368_0),.clk(gclk));
	jdff dff_A_AlW9APjx6_0(.dout(w_dff_A_heQ81J368_0),.din(w_dff_A_AlW9APjx6_0),.clk(gclk));
	jdff dff_A_AzYgYmxN5_0(.dout(w_dff_A_AlW9APjx6_0),.din(w_dff_A_AzYgYmxN5_0),.clk(gclk));
	jdff dff_A_4R66MgMk3_1(.dout(w_G87_2[1]),.din(w_dff_A_4R66MgMk3_1),.clk(gclk));
	jdff dff_A_YzT3lXEH0_1(.dout(w_dff_A_4R66MgMk3_1),.din(w_dff_A_YzT3lXEH0_1),.clk(gclk));
	jdff dff_A_dRsxdNdo2_1(.dout(w_dff_A_YzT3lXEH0_1),.din(w_dff_A_dRsxdNdo2_1),.clk(gclk));
	jdff dff_A_3XLrzspX8_1(.dout(w_dff_A_dRsxdNdo2_1),.din(w_dff_A_3XLrzspX8_1),.clk(gclk));
	jdff dff_A_OYmyEwU07_1(.dout(w_n149_1[1]),.din(w_dff_A_OYmyEwU07_1),.clk(gclk));
	jdff dff_A_Xyt08d892_1(.dout(w_dff_A_OYmyEwU07_1),.din(w_dff_A_Xyt08d892_1),.clk(gclk));
	jdff dff_B_5oDl5aKy0_1(.din(n375),.dout(w_dff_B_5oDl5aKy0_1),.clk(gclk));
	jdff dff_A_0p8q4oEL4_0(.dout(w_G232_1[0]),.din(w_dff_A_0p8q4oEL4_0),.clk(gclk));
	jdff dff_A_rPI04wTs3_0(.dout(w_dff_A_0p8q4oEL4_0),.din(w_dff_A_rPI04wTs3_0),.clk(gclk));
	jdff dff_A_4JHMJTxp3_1(.dout(w_G232_1[1]),.din(w_dff_A_4JHMJTxp3_1),.clk(gclk));
	jdff dff_A_EOEzw3Vb1_1(.dout(w_G232_0[1]),.din(w_dff_A_EOEzw3Vb1_1),.clk(gclk));
	jdff dff_A_AYPTE2zr5_1(.dout(w_dff_A_EOEzw3Vb1_1),.din(w_dff_A_AYPTE2zr5_1),.clk(gclk));
	jdff dff_A_z1MRiI3L0_1(.dout(w_dff_A_AYPTE2zr5_1),.din(w_dff_A_z1MRiI3L0_1),.clk(gclk));
	jdff dff_A_zfeHizBJ6_1(.dout(w_dff_A_z1MRiI3L0_1),.din(w_dff_A_zfeHizBJ6_1),.clk(gclk));
	jdff dff_A_hwWaFAFZ0_2(.dout(w_G232_0[2]),.din(w_dff_A_hwWaFAFZ0_2),.clk(gclk));
	jdff dff_A_CC0y3FIr4_2(.dout(w_dff_A_hwWaFAFZ0_2),.din(w_dff_A_CC0y3FIr4_2),.clk(gclk));
	jdff dff_B_8wZLjwLq1_0(.din(n538),.dout(w_dff_B_8wZLjwLq1_0),.clk(gclk));
	jdff dff_A_freTjB7M9_1(.dout(w_n532_0[1]),.din(w_dff_A_freTjB7M9_1),.clk(gclk));
	jdff dff_B_tmtaSXRO8_1(.din(n525),.dout(w_dff_B_tmtaSXRO8_1),.clk(gclk));
	jdff dff_A_sJNSF0Ru5_1(.dout(w_n524_0[1]),.din(w_dff_A_sJNSF0Ru5_1),.clk(gclk));
	jdff dff_A_ZsxRKSK08_0(.dout(w_n523_0[0]),.din(w_dff_A_ZsxRKSK08_0),.clk(gclk));
	jdff dff_A_m4ejHiAa8_2(.dout(w_n588_0[2]),.din(w_dff_A_m4ejHiAa8_2),.clk(gclk));
	jdff dff_A_NeBlkTsm6_2(.dout(w_dff_A_m4ejHiAa8_2),.din(w_dff_A_NeBlkTsm6_2),.clk(gclk));
	jdff dff_B_ShiCuMxf1_0(.din(n587),.dout(w_dff_B_ShiCuMxf1_0),.clk(gclk));
	jdff dff_B_LVfRVNFb1_1(.din(n580),.dout(w_dff_B_LVfRVNFb1_1),.clk(gclk));
	jdff dff_B_1acgoLbH7_1(.din(n581),.dout(w_dff_B_1acgoLbH7_1),.clk(gclk));
	jdff dff_A_xefzw0Xr8_1(.dout(w_n554_2[1]),.din(w_dff_A_xefzw0Xr8_1),.clk(gclk));
	jdff dff_A_WS3oRN2k1_2(.dout(w_n554_2[2]),.din(w_dff_A_WS3oRN2k1_2),.clk(gclk));
	jdff dff_A_7SSjdnDc8_2(.dout(w_dff_A_WS3oRN2k1_2),.din(w_dff_A_7SSjdnDc8_2),.clk(gclk));
	jdff dff_A_xiYrl7Po4_2(.dout(w_dff_A_7SSjdnDc8_2),.din(w_dff_A_xiYrl7Po4_2),.clk(gclk));
	jdff dff_A_4vEzungA6_2(.dout(w_dff_A_xiYrl7Po4_2),.din(w_dff_A_4vEzungA6_2),.clk(gclk));
	jdff dff_A_jQrP0qoc7_2(.dout(w_dff_A_4vEzungA6_2),.din(w_dff_A_jQrP0qoc7_2),.clk(gclk));
	jdff dff_A_OPmw6A1f2_0(.dout(w_n554_0[0]),.din(w_dff_A_OPmw6A1f2_0),.clk(gclk));
	jdff dff_A_FsF9GHw87_0(.dout(w_dff_A_OPmw6A1f2_0),.din(w_dff_A_FsF9GHw87_0),.clk(gclk));
	jdff dff_A_LEHBkyB51_0(.dout(w_dff_A_FsF9GHw87_0),.din(w_dff_A_LEHBkyB51_0),.clk(gclk));
	jdff dff_A_VFWpqNBh3_1(.dout(w_n554_0[1]),.din(w_dff_A_VFWpqNBh3_1),.clk(gclk));
	jdff dff_A_hKnFbtoY1_1(.dout(w_dff_A_VFWpqNBh3_1),.din(w_dff_A_hKnFbtoY1_1),.clk(gclk));
	jdff dff_B_yf8mo9is2_3(.din(n554),.dout(w_dff_B_yf8mo9is2_3),.clk(gclk));
	jdff dff_B_msZ2tOuf0_3(.din(w_dff_B_yf8mo9is2_3),.dout(w_dff_B_msZ2tOuf0_3),.clk(gclk));
	jdff dff_A_enXX1quV3_0(.dout(w_n534_0[0]),.din(w_dff_A_enXX1quV3_0),.clk(gclk));
	jdff dff_A_jqIH72iD9_0(.dout(w_G330_0[0]),.din(w_dff_A_jqIH72iD9_0),.clk(gclk));
	jdff dff_A_GOOIVse66_0(.dout(w_dff_A_jqIH72iD9_0),.din(w_dff_A_GOOIVse66_0),.clk(gclk));
	jdff dff_A_NLwXJCfA3_0(.dout(w_dff_A_GOOIVse66_0),.din(w_dff_A_NLwXJCfA3_0),.clk(gclk));
	jdff dff_A_f6ABZmXF8_0(.dout(w_dff_A_NLwXJCfA3_0),.din(w_dff_A_f6ABZmXF8_0),.clk(gclk));
	jdff dff_A_jEYlmuyq8_0(.dout(w_dff_A_f6ABZmXF8_0),.din(w_dff_A_jEYlmuyq8_0),.clk(gclk));
	jdff dff_A_4pgYoo2E4_0(.dout(w_dff_A_jEYlmuyq8_0),.din(w_dff_A_4pgYoo2E4_0),.clk(gclk));
	jdff dff_A_VI4Ow6M03_0(.dout(w_dff_A_4pgYoo2E4_0),.din(w_dff_A_VI4Ow6M03_0),.clk(gclk));
	jdff dff_A_aiaFnVaD1_0(.dout(w_dff_A_VI4Ow6M03_0),.din(w_dff_A_aiaFnVaD1_0),.clk(gclk));
	jdff dff_A_HI4z6a6C1_0(.dout(w_dff_A_aiaFnVaD1_0),.din(w_dff_A_HI4z6a6C1_0),.clk(gclk));
	jdff dff_A_9HLKkSpm3_0(.dout(w_dff_A_HI4z6a6C1_0),.din(w_dff_A_9HLKkSpm3_0),.clk(gclk));
	jdff dff_A_91jmAvar1_0(.dout(w_dff_A_9HLKkSpm3_0),.din(w_dff_A_91jmAvar1_0),.clk(gclk));
	jdff dff_A_gGprMvpd8_0(.dout(w_dff_A_91jmAvar1_0),.din(w_dff_A_gGprMvpd8_0),.clk(gclk));
	jdff dff_A_VRV9qAWt3_0(.dout(w_n553_2[0]),.din(w_dff_A_VRV9qAWt3_0),.clk(gclk));
	jdff dff_A_UZPuOWI86_0(.dout(w_dff_A_VRV9qAWt3_0),.din(w_dff_A_UZPuOWI86_0),.clk(gclk));
	jdff dff_A_4aWkU8mK7_0(.dout(w_dff_A_UZPuOWI86_0),.din(w_dff_A_4aWkU8mK7_0),.clk(gclk));
	jdff dff_A_lu5uwDg92_0(.dout(w_dff_A_4aWkU8mK7_0),.din(w_dff_A_lu5uwDg92_0),.clk(gclk));
	jdff dff_A_KoQiKot56_0(.dout(w_dff_A_lu5uwDg92_0),.din(w_dff_A_KoQiKot56_0),.clk(gclk));
	jdff dff_A_UWsNxs513_0(.dout(w_dff_A_KoQiKot56_0),.din(w_dff_A_UWsNxs513_0),.clk(gclk));
	jdff dff_A_kz12i0ey7_0(.dout(w_dff_A_UWsNxs513_0),.din(w_dff_A_kz12i0ey7_0),.clk(gclk));
	jdff dff_A_9D9xGHVi8_0(.dout(w_dff_A_kz12i0ey7_0),.din(w_dff_A_9D9xGHVi8_0),.clk(gclk));
	jdff dff_A_KgJyM3XM4_0(.dout(w_dff_A_9D9xGHVi8_0),.din(w_dff_A_KgJyM3XM4_0),.clk(gclk));
	jdff dff_A_iIEJL7x26_1(.dout(w_n553_2[1]),.din(w_dff_A_iIEJL7x26_1),.clk(gclk));
	jdff dff_A_cdQ8lvh06_1(.dout(w_dff_A_iIEJL7x26_1),.din(w_dff_A_cdQ8lvh06_1),.clk(gclk));
	jdff dff_A_OwvypD2H7_1(.dout(w_dff_A_cdQ8lvh06_1),.din(w_dff_A_OwvypD2H7_1),.clk(gclk));
	jdff dff_A_14bn1H3V2_1(.dout(w_dff_A_OwvypD2H7_1),.din(w_dff_A_14bn1H3V2_1),.clk(gclk));
	jdff dff_A_H6Iufzoy3_1(.dout(w_dff_A_14bn1H3V2_1),.din(w_dff_A_H6Iufzoy3_1),.clk(gclk));
	jdff dff_A_NxuSkR1F8_0(.dout(w_n553_0[0]),.din(w_dff_A_NxuSkR1F8_0),.clk(gclk));
	jdff dff_A_qXdsbkWq8_0(.dout(w_dff_A_NxuSkR1F8_0),.din(w_dff_A_qXdsbkWq8_0),.clk(gclk));
	jdff dff_A_lkOogajD3_0(.dout(w_dff_A_qXdsbkWq8_0),.din(w_dff_A_lkOogajD3_0),.clk(gclk));
	jdff dff_A_6ibv6KxW6_0(.dout(w_dff_A_lkOogajD3_0),.din(w_dff_A_6ibv6KxW6_0),.clk(gclk));
	jdff dff_A_0ooMxjBe8_2(.dout(w_n553_0[2]),.din(w_dff_A_0ooMxjBe8_2),.clk(gclk));
	jdff dff_A_WfffUTBY0_2(.dout(w_dff_A_0ooMxjBe8_2),.din(w_dff_A_WfffUTBY0_2),.clk(gclk));
	jdff dff_A_QXkNSAJn4_2(.dout(w_dff_A_WfffUTBY0_2),.din(w_dff_A_QXkNSAJn4_2),.clk(gclk));
	jdff dff_A_5qQQlvTO6_2(.dout(w_dff_A_QXkNSAJn4_2),.din(w_dff_A_5qQQlvTO6_2),.clk(gclk));
	jdff dff_A_5IqAVncz2_2(.dout(w_dff_A_5qQQlvTO6_2),.din(w_dff_A_5IqAVncz2_2),.clk(gclk));
	jdff dff_A_MFGIaPWm2_2(.dout(w_dff_A_5IqAVncz2_2),.din(w_dff_A_MFGIaPWm2_2),.clk(gclk));
	jdff dff_A_bK8Nu5iM8_1(.dout(w_n552_0[1]),.din(w_dff_A_bK8Nu5iM8_1),.clk(gclk));
	jdff dff_A_7LcNbOki3_1(.dout(w_dff_A_bK8Nu5iM8_1),.din(w_dff_A_7LcNbOki3_1),.clk(gclk));
	jdff dff_A_fpDwdSui3_1(.dout(w_dff_A_7LcNbOki3_1),.din(w_dff_A_fpDwdSui3_1),.clk(gclk));
	jdff dff_A_H37i0v2h2_1(.dout(w_dff_A_fpDwdSui3_1),.din(w_dff_A_H37i0v2h2_1),.clk(gclk));
	jdff dff_A_yC9TF1hH3_1(.dout(w_dff_A_H37i0v2h2_1),.din(w_dff_A_yC9TF1hH3_1),.clk(gclk));
	jdff dff_A_PIWTNxa47_1(.dout(w_dff_A_yC9TF1hH3_1),.din(w_dff_A_PIWTNxa47_1),.clk(gclk));
	jdff dff_A_l6eqF4jg5_1(.dout(w_dff_A_PIWTNxa47_1),.din(w_dff_A_l6eqF4jg5_1),.clk(gclk));
	jdff dff_A_Nt9qYN4z2_2(.dout(w_n552_0[2]),.din(w_dff_A_Nt9qYN4z2_2),.clk(gclk));
	jdff dff_A_RWubiC2U0_2(.dout(w_dff_A_Nt9qYN4z2_2),.din(w_dff_A_RWubiC2U0_2),.clk(gclk));
	jdff dff_A_7yhEceqI7_2(.dout(w_dff_A_RWubiC2U0_2),.din(w_dff_A_7yhEceqI7_2),.clk(gclk));
	jdff dff_A_w3NQBbIP8_2(.dout(w_dff_A_7yhEceqI7_2),.din(w_dff_A_w3NQBbIP8_2),.clk(gclk));
	jdff dff_A_m20jSWco6_2(.dout(w_dff_A_w3NQBbIP8_2),.din(w_dff_A_m20jSWco6_2),.clk(gclk));
	jdff dff_A_pcLx0mV21_2(.dout(w_dff_A_m20jSWco6_2),.din(w_dff_A_pcLx0mV21_2),.clk(gclk));
	jdff dff_A_Q5eaKtoA0_2(.dout(w_dff_A_pcLx0mV21_2),.din(w_dff_A_Q5eaKtoA0_2),.clk(gclk));
	jdff dff_A_7xrzCvZ98_0(.dout(w_G213_0[0]),.din(w_dff_A_7xrzCvZ98_0),.clk(gclk));
	jdff dff_A_WHdKEeti2_2(.dout(w_G213_0[2]),.din(w_dff_A_WHdKEeti2_2),.clk(gclk));
	jdff dff_A_xfuiYykq1_0(.dout(w_n113_1[0]),.din(w_dff_A_xfuiYykq1_0),.clk(gclk));
	jdff dff_A_jXlgNbp25_0(.dout(w_dff_A_xfuiYykq1_0),.din(w_dff_A_jXlgNbp25_0),.clk(gclk));
	jdff dff_A_k8cXiJ2y9_1(.dout(w_n113_1[1]),.din(w_dff_A_k8cXiJ2y9_1),.clk(gclk));
	jdff dff_A_xBHXsD235_1(.dout(w_dff_A_k8cXiJ2y9_1),.din(w_dff_A_xBHXsD235_1),.clk(gclk));
	jdff dff_A_7HMNrkS60_1(.dout(w_dff_A_xBHXsD235_1),.din(w_dff_A_7HMNrkS60_1),.clk(gclk));
	jdff dff_A_9ajb0Fgk1_1(.dout(w_dff_A_7HMNrkS60_1),.din(w_dff_A_9ajb0Fgk1_1),.clk(gclk));
	jdff dff_A_hfgBgHRV7_1(.dout(w_dff_A_9ajb0Fgk1_1),.din(w_dff_A_hfgBgHRV7_1),.clk(gclk));
	jdff dff_A_L3eaQgWY6_1(.dout(w_dff_A_hfgBgHRV7_1),.din(w_dff_A_L3eaQgWY6_1),.clk(gclk));
	jdff dff_A_4BPmvvzp9_1(.dout(w_dff_A_L3eaQgWY6_1),.din(w_dff_A_4BPmvvzp9_1),.clk(gclk));
	jdff dff_A_dyn12HjZ2_1(.dout(w_dff_A_4BPmvvzp9_1),.din(w_dff_A_dyn12HjZ2_1),.clk(gclk));
	jdff dff_A_HyiWPJhq6_1(.dout(w_dff_A_dyn12HjZ2_1),.din(w_dff_A_HyiWPJhq6_1),.clk(gclk));
	jdff dff_A_m10HyTs41_1(.dout(w_dff_A_HyiWPJhq6_1),.din(w_dff_A_m10HyTs41_1),.clk(gclk));
	jdff dff_A_XXE2nEhX0_1(.dout(w_dff_A_m10HyTs41_1),.din(w_dff_A_XXE2nEhX0_1),.clk(gclk));
	jdff dff_A_ptdNnmc79_1(.dout(w_dff_A_XXE2nEhX0_1),.din(w_dff_A_ptdNnmc79_1),.clk(gclk));
	jdff dff_A_Q8B1EI8U6_1(.dout(w_dff_A_ptdNnmc79_1),.din(w_dff_A_Q8B1EI8U6_1),.clk(gclk));
	jdff dff_A_28R9RAxr3_1(.dout(w_dff_A_Q8B1EI8U6_1),.din(w_dff_A_28R9RAxr3_1),.clk(gclk));
	jdff dff_A_ppYdNBXJ7_1(.dout(w_dff_A_28R9RAxr3_1),.din(w_dff_A_ppYdNBXJ7_1),.clk(gclk));
	jdff dff_A_8yOL4Dgw9_1(.dout(w_G343_0[1]),.din(w_dff_A_8yOL4Dgw9_1),.clk(gclk));
	jdff dff_A_oRsplpzq6_1(.dout(w_dff_A_8yOL4Dgw9_1),.din(w_dff_A_oRsplpzq6_1),.clk(gclk));
	jdff dff_A_mvZgpjTa2_1(.dout(w_dff_A_oRsplpzq6_1),.din(w_dff_A_mvZgpjTa2_1),.clk(gclk));
	jdff dff_A_vPeGR7Cb2_1(.dout(w_n374_0[1]),.din(w_dff_A_vPeGR7Cb2_1),.clk(gclk));
	jdff dff_B_M01Athst6_0(.din(n365),.dout(w_dff_B_M01Athst6_0),.clk(gclk));
	jdff dff_B_hX57umbd8_1(.din(n348),.dout(w_dff_B_hX57umbd8_1),.clk(gclk));
	jdff dff_B_AzoIUIvS6_1(.din(n343),.dout(w_dff_B_AzoIUIvS6_1),.clk(gclk));
	jdff dff_A_PBSqfgil2_0(.dout(w_n339_0[0]),.din(w_dff_A_PBSqfgil2_0),.clk(gclk));
	jdff dff_A_cYysVxzc5_0(.dout(w_dff_A_PBSqfgil2_0),.din(w_dff_A_cYysVxzc5_0),.clk(gclk));
	jdff dff_A_RiNEh80W2_0(.dout(w_G294_3[0]),.din(w_dff_A_RiNEh80W2_0),.clk(gclk));
	jdff dff_A_jOo9fuYz8_0(.dout(w_dff_A_RiNEh80W2_0),.din(w_dff_A_jOo9fuYz8_0),.clk(gclk));
	jdff dff_A_Imtw7rXu0_0(.dout(w_dff_A_jOo9fuYz8_0),.din(w_dff_A_Imtw7rXu0_0),.clk(gclk));
	jdff dff_A_h4Q5cbvG7_0(.dout(w_dff_A_Imtw7rXu0_0),.din(w_dff_A_h4Q5cbvG7_0),.clk(gclk));
	jdff dff_A_cZDb5ZWs9_0(.dout(w_G294_0[0]),.din(w_dff_A_cZDb5ZWs9_0),.clk(gclk));
	jdff dff_A_eCBS0RGn4_0(.dout(w_dff_A_cZDb5ZWs9_0),.din(w_dff_A_eCBS0RGn4_0),.clk(gclk));
	jdff dff_A_pBjB8zcm8_0(.dout(w_dff_A_eCBS0RGn4_0),.din(w_dff_A_pBjB8zcm8_0),.clk(gclk));
	jdff dff_A_CcQV7sao7_1(.dout(w_G294_0[1]),.din(w_dff_A_CcQV7sao7_1),.clk(gclk));
	jdff dff_A_907yCrwn3_1(.dout(w_dff_A_CcQV7sao7_1),.din(w_dff_A_907yCrwn3_1),.clk(gclk));
	jdff dff_A_5gty9tSV0_1(.dout(w_dff_A_907yCrwn3_1),.din(w_dff_A_5gty9tSV0_1),.clk(gclk));
	jdff dff_A_jKKD54u20_0(.dout(w_n196_1[0]),.din(w_dff_A_jKKD54u20_0),.clk(gclk));
	jdff dff_A_g5QmKHKA5_1(.dout(w_n196_1[1]),.din(w_dff_A_g5QmKHKA5_1),.clk(gclk));
	jdff dff_B_0hyWijOB1_0(.din(n335),.dout(w_dff_B_0hyWijOB1_0),.clk(gclk));
	jdff dff_A_8lUREGvv9_0(.dout(w_n334_0[0]),.din(w_dff_A_8lUREGvv9_0),.clk(gclk));
	jdff dff_A_X9o9EagP8_0(.dout(w_dff_A_8lUREGvv9_0),.din(w_dff_A_X9o9EagP8_0),.clk(gclk));
	jdff dff_B_YJgMbXiN0_0(.din(n333),.dout(w_dff_B_YJgMbXiN0_0),.clk(gclk));
	jdff dff_A_rDKXslHr0_0(.dout(w_G107_3[0]),.din(w_dff_A_rDKXslHr0_0),.clk(gclk));
	jdff dff_A_gTv3yu3c8_1(.dout(w_G107_3[1]),.din(w_dff_A_gTv3yu3c8_1),.clk(gclk));
	jdff dff_B_8oMyJe3n5_0(.din(n331),.dout(w_dff_B_8oMyJe3n5_0),.clk(gclk));
	jdff dff_B_dx20306R1_1(.din(n316),.dout(w_dff_B_dx20306R1_1),.clk(gclk));
	jdff dff_A_IdEcDTYM4_1(.dout(w_G190_3[1]),.din(w_dff_A_IdEcDTYM4_1),.clk(gclk));
	jdff dff_A_25vdNoTz2_1(.dout(w_dff_A_IdEcDTYM4_1),.din(w_dff_A_25vdNoTz2_1),.clk(gclk));
	jdff dff_A_xs3jEeia8_1(.dout(w_dff_A_25vdNoTz2_1),.din(w_dff_A_xs3jEeia8_1),.clk(gclk));
	jdff dff_A_K1vDXWvX4_1(.dout(w_dff_A_xs3jEeia8_1),.din(w_dff_A_K1vDXWvX4_1),.clk(gclk));
	jdff dff_A_VN3q0wQ22_1(.dout(w_dff_A_K1vDXWvX4_1),.din(w_dff_A_VN3q0wQ22_1),.clk(gclk));
	jdff dff_A_Eg5R2SEy7_1(.dout(w_dff_A_VN3q0wQ22_1),.din(w_dff_A_Eg5R2SEy7_1),.clk(gclk));
	jdff dff_A_qZwwkgyD6_1(.dout(w_dff_A_Eg5R2SEy7_1),.din(w_dff_A_qZwwkgyD6_1),.clk(gclk));
	jdff dff_A_xEzVN75u1_2(.dout(w_G190_3[2]),.din(w_dff_A_xEzVN75u1_2),.clk(gclk));
	jdff dff_A_xg4r9KJb0_2(.dout(w_dff_A_xEzVN75u1_2),.din(w_dff_A_xg4r9KJb0_2),.clk(gclk));
	jdff dff_A_IZgxIELf9_2(.dout(w_dff_A_xg4r9KJb0_2),.din(w_dff_A_IZgxIELf9_2),.clk(gclk));
	jdff dff_A_VD87RK157_2(.dout(w_dff_A_IZgxIELf9_2),.din(w_dff_A_VD87RK157_2),.clk(gclk));
	jdff dff_A_V41USIAe6_2(.dout(w_dff_A_VD87RK157_2),.din(w_dff_A_V41USIAe6_2),.clk(gclk));
	jdff dff_A_Hrh71dSF0_2(.dout(w_dff_A_V41USIAe6_2),.din(w_dff_A_Hrh71dSF0_2),.clk(gclk));
	jdff dff_A_LDnZStKM2_2(.dout(w_dff_A_Hrh71dSF0_2),.din(w_dff_A_LDnZStKM2_2),.clk(gclk));
	jdff dff_B_eIoYXnst0_0(.din(n317),.dout(w_dff_B_eIoYXnst0_0),.clk(gclk));
	jdff dff_B_HPMsywrA8_1(.din(n289),.dout(w_dff_B_HPMsywrA8_1),.clk(gclk));
	jdff dff_A_gxRNkctz1_1(.dout(w_n312_0[1]),.din(w_dff_A_gxRNkctz1_1),.clk(gclk));
	jdff dff_B_f909SO4t3_1(.din(n309),.dout(w_dff_B_f909SO4t3_1),.clk(gclk));
	jdff dff_A_V7oCZJGo4_0(.dout(w_n106_0[0]),.din(w_dff_A_V7oCZJGo4_0),.clk(gclk));
	jdff dff_A_i4efet1B6_0(.dout(w_dff_A_V7oCZJGo4_0),.din(w_dff_A_i4efet1B6_0),.clk(gclk));
	jdff dff_A_5OOqrkCz7_0(.dout(w_dff_A_i4efet1B6_0),.din(w_dff_A_5OOqrkCz7_0),.clk(gclk));
	jdff dff_A_xED5Ylry2_1(.dout(w_n88_0[1]),.din(w_dff_A_xED5Ylry2_1),.clk(gclk));
	jdff dff_A_FmN24kVt6_1(.dout(w_dff_A_xED5Ylry2_1),.din(w_dff_A_FmN24kVt6_1),.clk(gclk));
	jdff dff_A_szOXg0XM3_1(.dout(w_dff_A_FmN24kVt6_1),.din(w_dff_A_szOXg0XM3_1),.clk(gclk));
	jdff dff_A_k4uqZuK57_2(.dout(w_n88_0[2]),.din(w_dff_A_k4uqZuK57_2),.clk(gclk));
	jdff dff_A_mEmlEm6s2_1(.dout(w_n166_1[1]),.din(w_dff_A_mEmlEm6s2_1),.clk(gclk));
	jdff dff_A_pg5ld5f74_2(.dout(w_n166_1[2]),.din(w_dff_A_pg5ld5f74_2),.clk(gclk));
	jdff dff_A_3GIROOwX0_1(.dout(w_n303_0[1]),.din(w_dff_A_3GIROOwX0_1),.clk(gclk));
	jdff dff_A_Vd13r1yy1_1(.dout(w_n300_0[1]),.din(w_dff_A_Vd13r1yy1_1),.clk(gclk));
	jdff dff_A_kigN5drF4_0(.dout(w_n298_0[0]),.din(w_dff_A_kigN5drF4_0),.clk(gclk));
	jdff dff_A_Mcvi3e8f7_0(.dout(w_dff_A_kigN5drF4_0),.din(w_dff_A_Mcvi3e8f7_0),.clk(gclk));
	jdff dff_A_NoZTrR2V0_1(.dout(w_n185_2[1]),.din(w_dff_A_NoZTrR2V0_1),.clk(gclk));
	jdff dff_A_p17GX4UV7_1(.dout(w_dff_A_NoZTrR2V0_1),.din(w_dff_A_p17GX4UV7_1),.clk(gclk));
	jdff dff_A_n0VUd9i96_0(.dout(w_n105_1[0]),.din(w_dff_A_n0VUd9i96_0),.clk(gclk));
	jdff dff_A_sWlRsFGD9_2(.dout(w_n105_1[2]),.din(w_dff_A_sWlRsFGD9_2),.clk(gclk));
	jdff dff_A_K9aNkitx6_0(.dout(w_n296_0[0]),.din(w_dff_A_K9aNkitx6_0),.clk(gclk));
	jdff dff_A_diXvnU778_0(.dout(w_dff_A_K9aNkitx6_0),.din(w_dff_A_diXvnU778_0),.clk(gclk));
	jdff dff_A_Y2GmgOsp7_0(.dout(w_n105_0[0]),.din(w_dff_A_Y2GmgOsp7_0),.clk(gclk));
	jdff dff_A_ytftHHj82_2(.dout(w_n105_0[2]),.din(w_dff_A_ytftHHj82_2),.clk(gclk));
	jdff dff_A_Y4JxR3WW4_2(.dout(w_dff_A_ytftHHj82_2),.din(w_dff_A_Y4JxR3WW4_2),.clk(gclk));
	jdff dff_A_m5Q5lf740_2(.dout(w_dff_A_Y4JxR3WW4_2),.din(w_dff_A_m5Q5lf740_2),.clk(gclk));
	jdff dff_A_aA3KFQK93_0(.dout(w_G20_4[0]),.din(w_dff_A_aA3KFQK93_0),.clk(gclk));
	jdff dff_A_sEnV04eU0_1(.dout(w_G20_4[1]),.din(w_dff_A_sEnV04eU0_1),.clk(gclk));
	jdff dff_A_OnhiM6jf3_1(.dout(w_dff_A_sEnV04eU0_1),.din(w_dff_A_OnhiM6jf3_1),.clk(gclk));
	jdff dff_A_QxyDXSi28_1(.dout(w_dff_A_OnhiM6jf3_1),.din(w_dff_A_QxyDXSi28_1),.clk(gclk));
	jdff dff_A_fSTzQJGM8_1(.dout(w_dff_A_QxyDXSi28_1),.din(w_dff_A_fSTzQJGM8_1),.clk(gclk));
	jdff dff_A_vs3ZJwGa9_1(.dout(w_n189_1[1]),.din(w_dff_A_vs3ZJwGa9_1),.clk(gclk));
	jdff dff_A_F4dMoCGY8_0(.dout(w_G97_3[0]),.din(w_dff_A_F4dMoCGY8_0),.clk(gclk));
	jdff dff_A_JAB0NABu1_0(.dout(w_dff_A_F4dMoCGY8_0),.din(w_dff_A_JAB0NABu1_0),.clk(gclk));
	jdff dff_A_YTISlkpo1_0(.dout(w_dff_A_JAB0NABu1_0),.din(w_dff_A_YTISlkpo1_0),.clk(gclk));
	jdff dff_A_j389pyct4_1(.dout(w_G97_3[1]),.din(w_dff_A_j389pyct4_1),.clk(gclk));
	jdff dff_A_yhiv0qnJ2_1(.dout(w_dff_A_j389pyct4_1),.din(w_dff_A_yhiv0qnJ2_1),.clk(gclk));
	jdff dff_A_RpaMBR3p5_1(.dout(w_dff_A_yhiv0qnJ2_1),.din(w_dff_A_RpaMBR3p5_1),.clk(gclk));
	jdff dff_A_8jcRzIF35_0(.dout(w_G270_0[0]),.din(w_dff_A_8jcRzIF35_0),.clk(gclk));
	jdff dff_A_0kfJlfHL3_0(.dout(w_dff_A_8jcRzIF35_0),.din(w_dff_A_0kfJlfHL3_0),.clk(gclk));
	jdff dff_A_myBV1axo5_0(.dout(w_dff_A_0kfJlfHL3_0),.din(w_dff_A_myBV1axo5_0),.clk(gclk));
	jdff dff_A_gzwjnW8H8_0(.dout(w_dff_A_myBV1axo5_0),.din(w_dff_A_gzwjnW8H8_0),.clk(gclk));
	jdff dff_B_Mur7JrsD8_1(.din(n280),.dout(w_dff_B_Mur7JrsD8_1),.clk(gclk));
	jdff dff_A_4cmS3fqh7_1(.dout(w_n281_0[1]),.din(w_dff_A_4cmS3fqh7_1),.clk(gclk));
	jdff dff_A_BA5H7OT31_1(.dout(w_dff_A_4cmS3fqh7_1),.din(w_dff_A_BA5H7OT31_1),.clk(gclk));
	jdff dff_A_xrb7684A8_0(.dout(w_G303_2[0]),.din(w_dff_A_xrb7684A8_0),.clk(gclk));
	jdff dff_A_vkj7UK126_0(.dout(w_dff_A_xrb7684A8_0),.din(w_dff_A_vkj7UK126_0),.clk(gclk));
	jdff dff_A_FRSK5cPf6_0(.dout(w_dff_A_vkj7UK126_0),.din(w_dff_A_FRSK5cPf6_0),.clk(gclk));
	jdff dff_A_buMYHT8l8_1(.dout(w_G303_2[1]),.din(w_dff_A_buMYHT8l8_1),.clk(gclk));
	jdff dff_A_qesgmJmZ7_1(.dout(w_dff_A_buMYHT8l8_1),.din(w_dff_A_qesgmJmZ7_1),.clk(gclk));
	jdff dff_A_CIgBAP6t9_1(.dout(w_dff_A_qesgmJmZ7_1),.din(w_dff_A_CIgBAP6t9_1),.clk(gclk));
	jdff dff_A_HEpS09PU5_1(.dout(w_dff_A_CIgBAP6t9_1),.din(w_dff_A_HEpS09PU5_1),.clk(gclk));
	jdff dff_A_OO5hki6w7_0(.dout(w_G303_0[0]),.din(w_dff_A_OO5hki6w7_0),.clk(gclk));
	jdff dff_A_IgAXfZzA0_0(.dout(w_dff_A_OO5hki6w7_0),.din(w_dff_A_IgAXfZzA0_0),.clk(gclk));
	jdff dff_A_Q36Cbjon5_0(.dout(w_dff_A_IgAXfZzA0_0),.din(w_dff_A_Q36Cbjon5_0),.clk(gclk));
	jdff dff_A_ud7KC6Dr5_2(.dout(w_G303_0[2]),.din(w_dff_A_ud7KC6Dr5_2),.clk(gclk));
	jdff dff_A_KoVECPo00_2(.dout(w_dff_A_ud7KC6Dr5_2),.din(w_dff_A_KoVECPo00_2),.clk(gclk));
	jdff dff_A_DVvo8ZCm3_2(.dout(w_dff_A_KoVECPo00_2),.din(w_dff_A_DVvo8ZCm3_2),.clk(gclk));
	jdff dff_A_phx9anFf7_2(.dout(w_dff_A_DVvo8ZCm3_2),.din(w_dff_A_phx9anFf7_2),.clk(gclk));
	jdff dff_A_kYlrdnQQ1_1(.dout(w_G264_0[1]),.din(w_dff_A_kYlrdnQQ1_1),.clk(gclk));
	jdff dff_A_tYn1OjxC8_1(.dout(w_dff_A_kYlrdnQQ1_1),.din(w_dff_A_tYn1OjxC8_1),.clk(gclk));
	jdff dff_A_WHrdW1Ds3_1(.dout(w_dff_A_tYn1OjxC8_1),.din(w_dff_A_WHrdW1Ds3_1),.clk(gclk));
	jdff dff_A_4UQrobXj6_1(.dout(w_dff_A_WHrdW1Ds3_1),.din(w_dff_A_4UQrobXj6_1),.clk(gclk));
	jdff dff_A_22UFqUHs9_2(.dout(w_G264_0[2]),.din(w_dff_A_22UFqUHs9_2),.clk(gclk));
	jdff dff_A_wQqteubQ1_2(.dout(w_dff_A_22UFqUHs9_2),.din(w_dff_A_wQqteubQ1_2),.clk(gclk));
	jdff dff_B_QdJvX37F8_1(.din(n268),.dout(w_dff_B_QdJvX37F8_1),.clk(gclk));
	jdff dff_A_OOS4yCBy7_1(.dout(w_n274_0[1]),.din(w_dff_A_OOS4yCBy7_1),.clk(gclk));
	jdff dff_A_ep0BYdZp7_0(.dout(w_n270_0[0]),.din(w_dff_A_ep0BYdZp7_0),.clk(gclk));
	jdff dff_B_b3AJGpTB4_2(.din(n270),.dout(w_dff_B_b3AJGpTB4_2),.clk(gclk));
	jdff dff_A_oB7QLt3h5_0(.dout(w_n112_4[0]),.din(w_dff_A_oB7QLt3h5_0),.clk(gclk));
	jdff dff_A_7vqWpU2b0_0(.dout(w_dff_A_oB7QLt3h5_0),.din(w_dff_A_7vqWpU2b0_0),.clk(gclk));
	jdff dff_A_8lZq8ZH51_0(.dout(w_dff_A_7vqWpU2b0_0),.din(w_dff_A_8lZq8ZH51_0),.clk(gclk));
	jdff dff_A_iYKKcq6s5_0(.dout(w_dff_A_8lZq8ZH51_0),.din(w_dff_A_iYKKcq6s5_0),.clk(gclk));
	jdff dff_A_epM4ApjK4_1(.dout(w_n112_4[1]),.din(w_dff_A_epM4ApjK4_1),.clk(gclk));
	jdff dff_A_d6qjtnqe1_0(.dout(w_G1_1[0]),.din(w_dff_A_d6qjtnqe1_0),.clk(gclk));
	jdff dff_A_sE9iFuPG8_0(.dout(w_dff_A_d6qjtnqe1_0),.din(w_dff_A_sE9iFuPG8_0),.clk(gclk));
	jdff dff_A_jhqvHvKy5_0(.dout(w_dff_A_sE9iFuPG8_0),.din(w_dff_A_jhqvHvKy5_0),.clk(gclk));
	jdff dff_A_RA3arEWY5_1(.dout(w_G1_1[1]),.din(w_dff_A_RA3arEWY5_1),.clk(gclk));
	jdff dff_B_wMQgszaN9_0(.din(n266),.dout(w_dff_B_wMQgszaN9_0),.clk(gclk));
	jdff dff_B_rjK55iLY6_1(.din(n260),.dout(w_dff_B_rjK55iLY6_1),.clk(gclk));
	jdff dff_A_XQVY9OJj8_0(.dout(w_n262_0[0]),.din(w_dff_A_XQVY9OJj8_0),.clk(gclk));
	jdff dff_A_WKwum4yB3_0(.dout(w_n259_0[0]),.din(w_dff_A_WKwum4yB3_0),.clk(gclk));
	jdff dff_A_Fhdl4g5f6_0(.dout(w_dff_A_WKwum4yB3_0),.din(w_dff_A_Fhdl4g5f6_0),.clk(gclk));
	jdff dff_A_kStMTVvA0_0(.dout(w_n257_0[0]),.din(w_dff_A_kStMTVvA0_0),.clk(gclk));
	jdff dff_A_0eUypARF3_1(.dout(w_n255_0[1]),.din(w_dff_A_0eUypARF3_1),.clk(gclk));
	jdff dff_A_zKYKHmZ62_0(.dout(w_G77_4[0]),.din(w_dff_A_zKYKHmZ62_0),.clk(gclk));
	jdff dff_A_dL83xHsC3_0(.dout(w_G77_1[0]),.din(w_dff_A_dL83xHsC3_0),.clk(gclk));
	jdff dff_A_dReq60Ge5_2(.dout(w_G77_1[2]),.din(w_dff_A_dReq60Ge5_2),.clk(gclk));
	jdff dff_A_LoneYxIj4_2(.dout(w_dff_A_dReq60Ge5_2),.din(w_dff_A_LoneYxIj4_2),.clk(gclk));
	jdff dff_A_EIUmMT0j9_2(.dout(w_dff_A_LoneYxIj4_2),.din(w_dff_A_EIUmMT0j9_2),.clk(gclk));
	jdff dff_A_hxoan87X8_2(.dout(w_dff_A_EIUmMT0j9_2),.din(w_dff_A_hxoan87X8_2),.clk(gclk));
	jdff dff_B_ZpafX9QN3_2(.din(n249),.dout(w_dff_B_ZpafX9QN3_2),.clk(gclk));
	jdff dff_B_Vq8gzTDt7_2(.din(w_dff_B_ZpafX9QN3_2),.dout(w_dff_B_Vq8gzTDt7_2),.clk(gclk));
	jdff dff_A_k9xFSACD7_0(.dout(w_G107_4[0]),.din(w_dff_A_k9xFSACD7_0),.clk(gclk));
	jdff dff_A_EPeBne8a8_0(.dout(w_dff_A_k9xFSACD7_0),.din(w_dff_A_EPeBne8a8_0),.clk(gclk));
	jdff dff_A_pLaXYgni3_0(.dout(w_dff_A_EPeBne8a8_0),.din(w_dff_A_pLaXYgni3_0),.clk(gclk));
	jdff dff_A_PVD5866S1_0(.dout(w_dff_A_pLaXYgni3_0),.din(w_dff_A_PVD5866S1_0),.clk(gclk));
	jdff dff_A_rkCxOl9m8_0(.dout(w_dff_A_PVD5866S1_0),.din(w_dff_A_rkCxOl9m8_0),.clk(gclk));
	jdff dff_A_diV3Ue6L8_0(.dout(w_dff_A_rkCxOl9m8_0),.din(w_dff_A_diV3Ue6L8_0),.clk(gclk));
	jdff dff_A_SYSv08G87_0(.dout(w_G33_8[0]),.din(w_dff_A_SYSv08G87_0),.clk(gclk));
	jdff dff_B_Pfjezq0K0_1(.din(n236),.dout(w_dff_B_Pfjezq0K0_1),.clk(gclk));
	jdff dff_B_Lh5p2nfy2_1(.din(n226),.dout(w_dff_B_Lh5p2nfy2_1),.clk(gclk));
	jdff dff_A_l2Iq00g77_0(.dout(w_n230_0[0]),.din(w_dff_A_l2Iq00g77_0),.clk(gclk));
	jdff dff_A_Veso47nX9_0(.dout(w_n151_3[0]),.din(w_dff_A_Veso47nX9_0),.clk(gclk));
	jdff dff_A_q6XlzzcL2_0(.dout(w_dff_A_Veso47nX9_0),.din(w_dff_A_q6XlzzcL2_0),.clk(gclk));
	jdff dff_A_WKO8z8L31_1(.dout(w_n151_3[1]),.din(w_dff_A_WKO8z8L31_1),.clk(gclk));
	jdff dff_A_puhMWKVZ2_1(.dout(w_dff_A_WKO8z8L31_1),.din(w_dff_A_puhMWKVZ2_1),.clk(gclk));
	jdff dff_A_Pd07LdMc2_0(.dout(w_n91_1[0]),.din(w_dff_A_Pd07LdMc2_0),.clk(gclk));
	jdff dff_A_E9VK3GGi0_0(.dout(w_dff_A_Pd07LdMc2_0),.din(w_dff_A_E9VK3GGi0_0),.clk(gclk));
	jdff dff_A_dERL1esi8_0(.dout(w_dff_A_E9VK3GGi0_0),.din(w_dff_A_dERL1esi8_0),.clk(gclk));
	jdff dff_A_4xdXvQ5i9_1(.dout(w_n91_0[1]),.din(w_dff_A_4xdXvQ5i9_1),.clk(gclk));
	jdff dff_A_Nj1xB4c89_0(.dout(w_G257_1[0]),.din(w_dff_A_Nj1xB4c89_0),.clk(gclk));
	jdff dff_A_Zk9P2qZg2_0(.dout(w_dff_A_Nj1xB4c89_0),.din(w_dff_A_Zk9P2qZg2_0),.clk(gclk));
	jdff dff_A_b8kFfbc09_0(.dout(w_dff_A_Zk9P2qZg2_0),.din(w_dff_A_b8kFfbc09_0),.clk(gclk));
	jdff dff_A_gflqMBrW2_0(.dout(w_dff_A_b8kFfbc09_0),.din(w_dff_A_gflqMBrW2_0),.clk(gclk));
	jdff dff_A_gmoFzwOH9_1(.dout(w_G257_1[1]),.din(w_dff_A_gmoFzwOH9_1),.clk(gclk));
	jdff dff_A_S3Ofe1LR7_1(.dout(w_G257_0[1]),.din(w_dff_A_S3Ofe1LR7_1),.clk(gclk));
	jdff dff_A_ancPBdLJ4_1(.dout(w_dff_A_S3Ofe1LR7_1),.din(w_dff_A_ancPBdLJ4_1),.clk(gclk));
	jdff dff_A_edXna7eJ5_2(.dout(w_G257_0[2]),.din(w_dff_A_edXna7eJ5_2),.clk(gclk));
	jdff dff_A_7iP5EJLw6_2(.dout(w_dff_A_edXna7eJ5_2),.din(w_dff_A_7iP5EJLw6_2),.clk(gclk));
	jdff dff_A_LxrKDjch3_1(.dout(w_n228_0[1]),.din(w_dff_A_LxrKDjch3_1),.clk(gclk));
	jdff dff_A_ohRw46K36_0(.dout(w_n221_0[0]),.din(w_dff_A_ohRw46K36_0),.clk(gclk));
	jdff dff_A_3JjXdUhZ0_0(.dout(w_dff_A_ohRw46K36_0),.din(w_dff_A_3JjXdUhZ0_0),.clk(gclk));
	jdff dff_A_NhpZJ60q4_1(.dout(w_n221_0[1]),.din(w_dff_A_NhpZJ60q4_1),.clk(gclk));
	jdff dff_A_DwDP3ax58_1(.dout(w_dff_A_NhpZJ60q4_1),.din(w_dff_A_DwDP3ax58_1),.clk(gclk));
	jdff dff_A_a661qqWF4_0(.dout(w_G283_3[0]),.din(w_dff_A_a661qqWF4_0),.clk(gclk));
	jdff dff_A_gin0FYtn7_0(.dout(w_dff_A_a661qqWF4_0),.din(w_dff_A_gin0FYtn7_0),.clk(gclk));
	jdff dff_A_vm3CoLng7_0(.dout(w_dff_A_gin0FYtn7_0),.din(w_dff_A_vm3CoLng7_0),.clk(gclk));
	jdff dff_A_nop1cqlb2_1(.dout(w_G283_3[1]),.din(w_dff_A_nop1cqlb2_1),.clk(gclk));
	jdff dff_A_qi5N4hBn9_1(.dout(w_dff_A_nop1cqlb2_1),.din(w_dff_A_qi5N4hBn9_1),.clk(gclk));
	jdff dff_A_JHrJ7IEG6_1(.dout(w_dff_A_qi5N4hBn9_1),.din(w_dff_A_JHrJ7IEG6_1),.clk(gclk));
	jdff dff_A_e8sfntoC4_1(.dout(w_dff_A_JHrJ7IEG6_1),.din(w_dff_A_e8sfntoC4_1),.clk(gclk));
	jdff dff_A_NdYvpb6L3_0(.dout(w_G283_0[0]),.din(w_dff_A_NdYvpb6L3_0),.clk(gclk));
	jdff dff_A_Ky48hNU60_0(.dout(w_dff_A_NdYvpb6L3_0),.din(w_dff_A_Ky48hNU60_0),.clk(gclk));
	jdff dff_A_OrDQkYHF2_0(.dout(w_dff_A_Ky48hNU60_0),.din(w_dff_A_OrDQkYHF2_0),.clk(gclk));
	jdff dff_A_Rq2WqyD75_1(.dout(w_G283_0[1]),.din(w_dff_A_Rq2WqyD75_1),.clk(gclk));
	jdff dff_A_WgHVasRv6_1(.dout(w_dff_A_Rq2WqyD75_1),.din(w_dff_A_WgHVasRv6_1),.clk(gclk));
	jdff dff_A_BEM9gBeJ0_1(.dout(w_dff_A_WgHVasRv6_1),.din(w_dff_A_BEM9gBeJ0_1),.clk(gclk));
	jdff dff_A_vdMaJsxe1_2(.dout(w_n166_2[2]),.din(w_dff_A_vdMaJsxe1_2),.clk(gclk));
	jdff dff_B_JFQs6Cz90_1(.din(n215),.dout(w_dff_B_JFQs6Cz90_1),.clk(gclk));
	jdff dff_A_myor13xe4_0(.dout(w_G200_1[0]),.din(w_dff_A_myor13xe4_0),.clk(gclk));
	jdff dff_A_0xjxALv33_0(.dout(w_dff_A_myor13xe4_0),.din(w_dff_A_0xjxALv33_0),.clk(gclk));
	jdff dff_A_Cqq1PXCx8_0(.dout(w_dff_A_0xjxALv33_0),.din(w_dff_A_Cqq1PXCx8_0),.clk(gclk));
	jdff dff_A_fMhCZthv7_0(.dout(w_dff_A_Cqq1PXCx8_0),.din(w_dff_A_fMhCZthv7_0),.clk(gclk));
	jdff dff_A_tHjXO9qn9_0(.dout(w_dff_A_fMhCZthv7_0),.din(w_dff_A_tHjXO9qn9_0),.clk(gclk));
	jdff dff_A_w7jeGZ1o2_0(.dout(w_dff_A_tHjXO9qn9_0),.din(w_dff_A_w7jeGZ1o2_0),.clk(gclk));
	jdff dff_A_04AmFTHf6_0(.dout(w_dff_A_w7jeGZ1o2_0),.din(w_dff_A_04AmFTHf6_0),.clk(gclk));
	jdff dff_A_dvjVEWxA4_1(.dout(w_G200_1[1]),.din(w_dff_A_dvjVEWxA4_1),.clk(gclk));
	jdff dff_A_Vj3zXUSD7_2(.dout(w_G200_0[2]),.din(w_dff_A_Vj3zXUSD7_2),.clk(gclk));
	jdff dff_A_zEvWIwJo2_2(.dout(w_dff_A_Vj3zXUSD7_2),.din(w_dff_A_zEvWIwJo2_2),.clk(gclk));
	jdff dff_A_S5qBGsov9_2(.dout(w_dff_A_zEvWIwJo2_2),.din(w_dff_A_S5qBGsov9_2),.clk(gclk));
	jdff dff_A_DvuEtOEI0_2(.dout(w_dff_A_S5qBGsov9_2),.din(w_dff_A_DvuEtOEI0_2),.clk(gclk));
	jdff dff_A_AC7C3EdM4_2(.dout(w_dff_A_DvuEtOEI0_2),.din(w_dff_A_AC7C3EdM4_2),.clk(gclk));
	jdff dff_A_zNAJmdNo3_2(.dout(w_dff_A_AC7C3EdM4_2),.din(w_dff_A_zNAJmdNo3_2),.clk(gclk));
	jdff dff_A_tSw5gpj66_2(.dout(w_dff_A_zNAJmdNo3_2),.din(w_dff_A_tSw5gpj66_2),.clk(gclk));
	jdff dff_A_h3hOAETZ3_0(.dout(w_G190_4[0]),.din(w_dff_A_h3hOAETZ3_0),.clk(gclk));
	jdff dff_A_eTefsioD9_0(.dout(w_G190_1[0]),.din(w_dff_A_eTefsioD9_0),.clk(gclk));
	jdff dff_A_NYW3Xivn3_0(.dout(w_dff_A_eTefsioD9_0),.din(w_dff_A_NYW3Xivn3_0),.clk(gclk));
	jdff dff_A_vTaEXAVh6_0(.dout(w_dff_A_NYW3Xivn3_0),.din(w_dff_A_vTaEXAVh6_0),.clk(gclk));
	jdff dff_A_lU4zRC4C0_0(.dout(w_dff_A_vTaEXAVh6_0),.din(w_dff_A_lU4zRC4C0_0),.clk(gclk));
	jdff dff_A_KmYiWHCA8_0(.dout(w_G190_0[0]),.din(w_dff_A_KmYiWHCA8_0),.clk(gclk));
	jdff dff_A_gp0OvPEx3_0(.dout(w_dff_A_KmYiWHCA8_0),.din(w_dff_A_gp0OvPEx3_0),.clk(gclk));
	jdff dff_A_KuEorIls1_1(.dout(w_G190_0[1]),.din(w_dff_A_KuEorIls1_1),.clk(gclk));
	jdff dff_A_1pNUcVq28_1(.dout(w_dff_A_KuEorIls1_1),.din(w_dff_A_1pNUcVq28_1),.clk(gclk));
	jdff dff_A_8WEsy4756_1(.dout(w_dff_A_1pNUcVq28_1),.din(w_dff_A_8WEsy4756_1),.clk(gclk));
	jdff dff_A_aeTsSMyu8_1(.dout(w_n214_0[1]),.din(w_dff_A_aeTsSMyu8_1),.clk(gclk));
	jdff dff_A_t2h3zT050_1(.dout(w_n213_0[1]),.din(w_dff_A_t2h3zT050_1),.clk(gclk));
	jdff dff_A_D5ioe1ut3_0(.dout(w_n210_0[0]),.din(w_dff_A_D5ioe1ut3_0),.clk(gclk));
	jdff dff_A_UiqxvAbc6_0(.dout(w_n205_0[0]),.din(w_dff_A_UiqxvAbc6_0),.clk(gclk));
	jdff dff_B_XO0IhvhS0_2(.din(n205),.dout(w_dff_B_XO0IhvhS0_2),.clk(gclk));
	jdff dff_A_OaCuvt4G3_0(.dout(w_n201_0[0]),.din(w_dff_A_OaCuvt4G3_0),.clk(gclk));
	jdff dff_A_zh0VzruW5_2(.dout(w_G33_9[2]),.din(w_dff_A_zh0VzruW5_2),.clk(gclk));
	jdff dff_A_iEPVGXbc1_1(.dout(w_n103_0[1]),.din(w_dff_A_iEPVGXbc1_1),.clk(gclk));
	jdff dff_A_AFPinfUT7_0(.dout(w_n196_2[0]),.din(w_dff_A_AFPinfUT7_0),.clk(gclk));
	jdff dff_A_6560CfKM2_1(.dout(w_n196_2[1]),.din(w_dff_A_6560CfKM2_1),.clk(gclk));
	jdff dff_A_r7UpT6j45_0(.dout(w_n196_0[0]),.din(w_dff_A_r7UpT6j45_0),.clk(gclk));
	jdff dff_A_jYX9ILcw5_2(.dout(w_n196_0[2]),.din(w_dff_A_jYX9ILcw5_2),.clk(gclk));
	jdff dff_B_2j51IpD02_3(.din(n196),.dout(w_dff_B_2j51IpD02_3),.clk(gclk));
	jdff dff_B_6ZjQg0y14_3(.din(w_dff_B_2j51IpD02_3),.dout(w_dff_B_6ZjQg0y14_3),.clk(gclk));
	jdff dff_B_0K4ozC484_3(.din(w_dff_B_6ZjQg0y14_3),.dout(w_dff_B_0K4ozC484_3),.clk(gclk));
	jdff dff_B_Kx6Og7Dy1_3(.din(w_dff_B_0K4ozC484_3),.dout(w_dff_B_Kx6Og7Dy1_3),.clk(gclk));
	jdff dff_B_3i5XDcRf5_3(.din(w_dff_B_Kx6Og7Dy1_3),.dout(w_dff_B_3i5XDcRf5_3),.clk(gclk));
	jdff dff_A_SdzZ5niv9_0(.dout(w_G179_2[0]),.din(w_dff_A_SdzZ5niv9_0),.clk(gclk));
	jdff dff_A_Op3Y7Qyk3_0(.dout(w_dff_A_SdzZ5niv9_0),.din(w_dff_A_Op3Y7Qyk3_0),.clk(gclk));
	jdff dff_A_6Bh61tbJ4_0(.dout(w_dff_A_Op3Y7Qyk3_0),.din(w_dff_A_6Bh61tbJ4_0),.clk(gclk));
	jdff dff_A_zBWmPbHG3_0(.dout(w_dff_A_6Bh61tbJ4_0),.din(w_dff_A_zBWmPbHG3_0),.clk(gclk));
	jdff dff_A_Y1JWnzVp6_0(.dout(w_dff_A_zBWmPbHG3_0),.din(w_dff_A_Y1JWnzVp6_0),.clk(gclk));
	jdff dff_A_qFpA9wC00_0(.dout(w_dff_A_Y1JWnzVp6_0),.din(w_dff_A_qFpA9wC00_0),.clk(gclk));
	jdff dff_A_0Cd7dMhP4_0(.dout(w_dff_A_qFpA9wC00_0),.din(w_dff_A_0Cd7dMhP4_0),.clk(gclk));
	jdff dff_A_tEBnN8hb4_1(.dout(w_G179_2[1]),.din(w_dff_A_tEBnN8hb4_1),.clk(gclk));
	jdff dff_A_Q9Jvy1F31_1(.dout(w_dff_A_tEBnN8hb4_1),.din(w_dff_A_Q9Jvy1F31_1),.clk(gclk));
	jdff dff_A_BvBckVrT2_1(.dout(w_dff_A_Q9Jvy1F31_1),.din(w_dff_A_BvBckVrT2_1),.clk(gclk));
	jdff dff_A_ZPJlTqa26_1(.dout(w_dff_A_BvBckVrT2_1),.din(w_dff_A_ZPJlTqa26_1),.clk(gclk));
	jdff dff_A_svGUg6Zs8_1(.dout(w_dff_A_ZPJlTqa26_1),.din(w_dff_A_svGUg6Zs8_1),.clk(gclk));
	jdff dff_A_PDTYNlM86_1(.dout(w_dff_A_svGUg6Zs8_1),.din(w_dff_A_PDTYNlM86_1),.clk(gclk));
	jdff dff_A_hueIkzjX5_1(.dout(w_dff_A_PDTYNlM86_1),.din(w_dff_A_hueIkzjX5_1),.clk(gclk));
	jdff dff_A_7goX015T1_0(.dout(w_G179_0[0]),.din(w_dff_A_7goX015T1_0),.clk(gclk));
	jdff dff_A_ztx9r2Kk8_0(.dout(w_dff_A_7goX015T1_0),.din(w_dff_A_ztx9r2Kk8_0),.clk(gclk));
	jdff dff_A_8lMDIxq95_0(.dout(w_dff_A_ztx9r2Kk8_0),.din(w_dff_A_8lMDIxq95_0),.clk(gclk));
	jdff dff_A_VZusJvtW5_0(.dout(w_dff_A_8lMDIxq95_0),.din(w_dff_A_VZusJvtW5_0),.clk(gclk));
	jdff dff_A_LLg45RjN1_0(.dout(w_dff_A_VZusJvtW5_0),.din(w_dff_A_LLg45RjN1_0),.clk(gclk));
	jdff dff_A_dPZsFRWr1_0(.dout(w_dff_A_LLg45RjN1_0),.din(w_dff_A_dPZsFRWr1_0),.clk(gclk));
	jdff dff_A_9SVGVaCc9_0(.dout(w_dff_A_dPZsFRWr1_0),.din(w_dff_A_9SVGVaCc9_0),.clk(gclk));
	jdff dff_B_ZzgSafiw8_0(.din(n192),.dout(w_dff_B_ZzgSafiw8_0),.clk(gclk));
	jdff dff_A_JQXtkOfm4_1(.dout(w_n190_1[1]),.din(w_dff_A_JQXtkOfm4_1),.clk(gclk));
	jdff dff_A_jlBU6s221_0(.dout(w_n189_2[0]),.din(w_dff_A_jlBU6s221_0),.clk(gclk));
	jdff dff_A_3zB2eNgH8_0(.dout(w_dff_A_jlBU6s221_0),.din(w_dff_A_3zB2eNgH8_0),.clk(gclk));
	jdff dff_A_lQeOl7ID9_2(.dout(w_n189_0[2]),.din(w_dff_A_lQeOl7ID9_2),.clk(gclk));
	jdff dff_A_bCeVzPG46_0(.dout(w_n85_0[0]),.din(w_dff_A_bCeVzPG46_0),.clk(gclk));
	jdff dff_A_ySZaPlsh8_0(.dout(w_dff_A_bCeVzPG46_0),.din(w_dff_A_ySZaPlsh8_0),.clk(gclk));
	jdff dff_A_vaFRwjF51_2(.dout(w_n85_0[2]),.din(w_dff_A_vaFRwjF51_2),.clk(gclk));
	jdff dff_A_LwmgBJME5_2(.dout(w_dff_A_vaFRwjF51_2),.din(w_dff_A_LwmgBJME5_2),.clk(gclk));
	jdff dff_A_9SLDHbAe5_2(.dout(w_dff_A_LwmgBJME5_2),.din(w_dff_A_9SLDHbAe5_2),.clk(gclk));
	jdff dff_A_migydITg8_2(.dout(w_dff_A_9SLDHbAe5_2),.din(w_dff_A_migydITg8_2),.clk(gclk));
	jdff dff_A_W57appsB7_0(.dout(w_G20_5[0]),.din(w_dff_A_W57appsB7_0),.clk(gclk));
	jdff dff_A_rvJlGxMM5_1(.dout(w_G20_5[1]),.din(w_dff_A_rvJlGxMM5_1),.clk(gclk));
	jdff dff_A_J1r9uf2M9_1(.dout(w_n80_0[1]),.din(w_dff_A_J1r9uf2M9_1),.clk(gclk));
	jdff dff_A_hmRUict03_1(.dout(w_dff_A_J1r9uf2M9_1),.din(w_dff_A_hmRUict03_1),.clk(gclk));
	jdff dff_A_aqb3i7Wl7_1(.dout(w_dff_A_hmRUict03_1),.din(w_dff_A_aqb3i7Wl7_1),.clk(gclk));
	jdff dff_A_HHjywFP82_2(.dout(w_n80_0[2]),.din(w_dff_A_HHjywFP82_2),.clk(gclk));
	jdff dff_A_Zb3xwYVa1_2(.dout(w_dff_A_HHjywFP82_2),.din(w_dff_A_Zb3xwYVa1_2),.clk(gclk));
	jdff dff_A_fba0B7RA2_2(.dout(w_dff_A_Zb3xwYVa1_2),.din(w_dff_A_fba0B7RA2_2),.clk(gclk));
	jdff dff_A_0WhyBnTx4_2(.dout(w_dff_A_fba0B7RA2_2),.din(w_dff_A_0WhyBnTx4_2),.clk(gclk));
	jdff dff_A_zOTSQUUw9_2(.dout(w_dff_A_0WhyBnTx4_2),.din(w_dff_A_zOTSQUUw9_2),.clk(gclk));
	jdff dff_A_xy0sGcsL6_2(.dout(w_G107_1[2]),.din(w_dff_A_xy0sGcsL6_2),.clk(gclk));
	jdff dff_A_vPPBpKop8_2(.dout(w_dff_A_xy0sGcsL6_2),.din(w_dff_A_vPPBpKop8_2),.clk(gclk));
	jdff dff_A_mELiXizb9_2(.dout(w_dff_A_vPPBpKop8_2),.din(w_dff_A_mELiXizb9_2),.clk(gclk));
	jdff dff_A_I8vtH30z0_1(.dout(w_G107_0[1]),.din(w_dff_A_I8vtH30z0_1),.clk(gclk));
	jdff dff_A_UNJo7RyV4_1(.dout(w_dff_A_I8vtH30z0_1),.din(w_dff_A_UNJo7RyV4_1),.clk(gclk));
	jdff dff_A_zpj0968i2_1(.dout(w_dff_A_UNJo7RyV4_1),.din(w_dff_A_zpj0968i2_1),.clk(gclk));
	jdff dff_A_8g564uFz5_2(.dout(w_G107_0[2]),.din(w_dff_A_8g564uFz5_2),.clk(gclk));
	jdff dff_A_yvp6lg1U7_2(.dout(w_dff_A_8g564uFz5_2),.din(w_dff_A_yvp6lg1U7_2),.clk(gclk));
	jdff dff_A_41vnu8CB0_2(.dout(w_dff_A_yvp6lg1U7_2),.din(w_dff_A_41vnu8CB0_2),.clk(gclk));
	jdff dff_A_FyrA18Hj7_0(.dout(w_n79_0[0]),.din(w_dff_A_FyrA18Hj7_0),.clk(gclk));
	jdff dff_A_RA2zgpyC4_0(.dout(w_dff_A_FyrA18Hj7_0),.din(w_dff_A_RA2zgpyC4_0),.clk(gclk));
	jdff dff_A_KAbfLiU74_0(.dout(w_G97_5[0]),.din(w_dff_A_KAbfLiU74_0),.clk(gclk));
	jdff dff_A_LCf4WESU9_1(.dout(w_n97_1[1]),.din(w_dff_A_LCf4WESU9_1),.clk(gclk));
	jdff dff_A_627OoBlb1_0(.dout(w_n97_0[0]),.din(w_dff_A_627OoBlb1_0),.clk(gclk));
	jdff dff_A_kurh59Sd5_0(.dout(w_G87_3[0]),.din(w_dff_A_kurh59Sd5_0),.clk(gclk));
	jdff dff_A_eX8x4eDb8_2(.dout(w_G87_3[2]),.din(w_dff_A_eX8x4eDb8_2),.clk(gclk));
	jdff dff_A_0bJBcDI72_2(.dout(w_dff_A_eX8x4eDb8_2),.din(w_dff_A_0bJBcDI72_2),.clk(gclk));
	jdff dff_A_8CcwNKW05_2(.dout(w_dff_A_0bJBcDI72_2),.din(w_dff_A_8CcwNKW05_2),.clk(gclk));
	jdff dff_A_qyr4YAAL0_0(.dout(w_G87_0[0]),.din(w_dff_A_qyr4YAAL0_0),.clk(gclk));
	jdff dff_A_4NSeATNu0_0(.dout(w_dff_A_qyr4YAAL0_0),.din(w_dff_A_4NSeATNu0_0),.clk(gclk));
	jdff dff_A_wlDyDHq85_0(.dout(w_dff_A_4NSeATNu0_0),.din(w_dff_A_wlDyDHq85_0),.clk(gclk));
	jdff dff_A_Rx4qNfI10_1(.dout(w_n179_0[1]),.din(w_dff_A_Rx4qNfI10_1),.clk(gclk));
	jdff dff_A_B5O5RWX09_1(.dout(w_dff_A_Rx4qNfI10_1),.din(w_dff_A_B5O5RWX09_1),.clk(gclk));
	jdff dff_A_0ZObVAKv4_2(.dout(w_n179_0[2]),.din(w_dff_A_0ZObVAKv4_2),.clk(gclk));
	jdff dff_A_STJGStVK6_2(.dout(w_dff_A_0ZObVAKv4_2),.din(w_dff_A_STJGStVK6_2),.clk(gclk));
	jdff dff_A_fdHaWDMG5_2(.dout(w_n112_5[2]),.din(w_dff_A_fdHaWDMG5_2),.clk(gclk));
	jdff dff_A_3ugz4ekH2_1(.dout(w_G20_2[1]),.din(w_dff_A_3ugz4ekH2_1),.clk(gclk));
	jdff dff_A_GckQdKlQ9_0(.dout(w_G68_4[0]),.din(w_dff_A_GckQdKlQ9_0),.clk(gclk));
	jdff dff_A_bpt5RxmD3_1(.dout(w_G68_4[1]),.din(w_dff_A_bpt5RxmD3_1),.clk(gclk));
	jdff dff_A_gPbxcvWN4_0(.dout(w_G68_1[0]),.din(w_dff_A_gPbxcvWN4_0),.clk(gclk));
	jdff dff_A_cdRuprlC3_2(.dout(w_G68_1[2]),.din(w_dff_A_cdRuprlC3_2),.clk(gclk));
	jdff dff_A_Aan9hUfF7_2(.dout(w_dff_A_cdRuprlC3_2),.din(w_dff_A_Aan9hUfF7_2),.clk(gclk));
	jdff dff_A_9F1ay21P3_2(.dout(w_dff_A_Aan9hUfF7_2),.din(w_dff_A_9F1ay21P3_2),.clk(gclk));
	jdff dff_A_RNnn8wkf2_2(.dout(w_dff_A_9F1ay21P3_2),.din(w_dff_A_RNnn8wkf2_2),.clk(gclk));
	jdff dff_A_iHywy3nW6_2(.dout(w_G68_0[2]),.din(w_dff_A_iHywy3nW6_2),.clk(gclk));
	jdff dff_A_xLbWa16Q8_1(.dout(w_n148_8[1]),.din(w_dff_A_xLbWa16Q8_1),.clk(gclk));
	jdff dff_A_H1BMiCLW6_0(.dout(w_G20_6[0]),.din(w_dff_A_H1BMiCLW6_0),.clk(gclk));
	jdff dff_A_a8iaffyV9_2(.dout(w_G20_1[2]),.din(w_dff_A_a8iaffyV9_2),.clk(gclk));
	jdff dff_A_PrKjblqV4_0(.dout(w_G20_0[0]),.din(w_dff_A_PrKjblqV4_0),.clk(gclk));
	jdff dff_B_5J6oeO852_2(.din(n172),.dout(w_dff_B_5J6oeO852_2),.clk(gclk));
	jdff dff_B_EMpldElG0_2(.din(w_dff_B_5J6oeO852_2),.dout(w_dff_B_EMpldElG0_2),.clk(gclk));
	jdff dff_A_iE1iT1Y11_0(.dout(w_G97_4[0]),.din(w_dff_A_iE1iT1Y11_0),.clk(gclk));
	jdff dff_A_ZAgSLwp21_0(.dout(w_dff_A_iE1iT1Y11_0),.din(w_dff_A_ZAgSLwp21_0),.clk(gclk));
	jdff dff_A_VSsmvDUq1_0(.dout(w_dff_A_ZAgSLwp21_0),.din(w_dff_A_VSsmvDUq1_0),.clk(gclk));
	jdff dff_A_3PEqnBcy6_2(.dout(w_G97_1[2]),.din(w_dff_A_3PEqnBcy6_2),.clk(gclk));
	jdff dff_A_NM1O3RPj3_2(.dout(w_dff_A_3PEqnBcy6_2),.din(w_dff_A_NM1O3RPj3_2),.clk(gclk));
	jdff dff_A_CVpa9cST4_2(.dout(w_dff_A_NM1O3RPj3_2),.din(w_dff_A_CVpa9cST4_2),.clk(gclk));
	jdff dff_A_UPHWAMW62_2(.dout(w_dff_A_CVpa9cST4_2),.din(w_dff_A_UPHWAMW62_2),.clk(gclk));
	jdff dff_A_TknSeaS27_1(.dout(w_G97_0[1]),.din(w_dff_A_TknSeaS27_1),.clk(gclk));
	jdff dff_A_VQWbXmd77_1(.dout(w_dff_A_TknSeaS27_1),.din(w_dff_A_VQWbXmd77_1),.clk(gclk));
	jdff dff_A_LbIR4ecf3_1(.dout(w_dff_A_VQWbXmd77_1),.din(w_dff_A_LbIR4ecf3_1),.clk(gclk));
	jdff dff_A_UERcl1tV7_2(.dout(w_G97_0[2]),.din(w_dff_A_UERcl1tV7_2),.clk(gclk));
	jdff dff_A_g5BCQ1hB0_0(.dout(w_G33_10[0]),.din(w_dff_A_g5BCQ1hB0_0),.clk(gclk));
	jdff dff_A_UJGM8GXu6_1(.dout(w_G33_10[1]),.din(w_dff_A_UJGM8GXu6_1),.clk(gclk));
	jdff dff_A_5F5KU4zg0_0(.dout(w_n170_0[0]),.din(w_dff_A_5F5KU4zg0_0),.clk(gclk));
	jdff dff_B_WNMm4euq5_0(.din(n169),.dout(w_dff_B_WNMm4euq5_0),.clk(gclk));
	jdff dff_A_glHElJOj6_0(.dout(w_G274_0[0]),.din(w_dff_A_glHElJOj6_0),.clk(gclk));
	jdff dff_A_1pW9fGce3_0(.dout(w_dff_A_glHElJOj6_0),.din(w_dff_A_1pW9fGce3_0),.clk(gclk));
	jdff dff_A_h6y2HzJO2_0(.dout(w_dff_A_1pW9fGce3_0),.din(w_dff_A_h6y2HzJO2_0),.clk(gclk));
	jdff dff_A_BVbQtBU74_2(.dout(w_G274_0[2]),.din(w_dff_A_BVbQtBU74_2),.clk(gclk));
	jdff dff_A_IZ76Ei1m6_2(.dout(w_dff_A_BVbQtBU74_2),.din(w_dff_A_IZ76Ei1m6_2),.clk(gclk));
	jdff dff_A_4s0TyoYc9_0(.dout(w_n166_3[0]),.din(w_dff_A_4s0TyoYc9_0),.clk(gclk));
	jdff dff_B_HqtnbwdP0_0(.din(n165),.dout(w_dff_B_HqtnbwdP0_0),.clk(gclk));
	jdff dff_A_E0S8gfdK9_2(.dout(w_n115_0[2]),.din(w_dff_A_E0S8gfdK9_2),.clk(gclk));
	jdff dff_A_wjUr3Scq4_0(.dout(w_n114_1[0]),.din(w_dff_A_wjUr3Scq4_0),.clk(gclk));
	jdff dff_A_ZwyCD0fH4_1(.dout(w_n114_0[1]),.din(w_dff_A_ZwyCD0fH4_1),.clk(gclk));
	jdff dff_A_1pje1mkK3_0(.dout(w_n163_0[0]),.din(w_dff_A_1pje1mkK3_0),.clk(gclk));
	jdff dff_A_vUIlcnRK2_2(.dout(w_n161_0[2]),.din(w_dff_A_vUIlcnRK2_2),.clk(gclk));
	jdff dff_A_T6R9xgvp5_2(.dout(w_dff_A_vUIlcnRK2_2),.din(w_dff_A_T6R9xgvp5_2),.clk(gclk));
	jdff dff_A_JyxtuiHL2_2(.dout(w_dff_A_T6R9xgvp5_2),.din(w_dff_A_JyxtuiHL2_2),.clk(gclk));
	jdff dff_A_a8nK50Vz3_0(.dout(w_G45_1[0]),.din(w_dff_A_a8nK50Vz3_0),.clk(gclk));
	jdff dff_A_6srOqm5Z0_0(.dout(w_dff_A_a8nK50Vz3_0),.din(w_dff_A_6srOqm5Z0_0),.clk(gclk));
	jdff dff_A_js40K4Sf9_1(.dout(w_G45_1[1]),.din(w_dff_A_js40K4Sf9_1),.clk(gclk));
	jdff dff_A_jMjaoHUR0_1(.dout(w_G45_0[1]),.din(w_dff_A_jMjaoHUR0_1),.clk(gclk));
	jdff dff_A_dXhCYzvS6_1(.dout(w_dff_A_jMjaoHUR0_1),.din(w_dff_A_dXhCYzvS6_1),.clk(gclk));
	jdff dff_A_LKBQMA7Q4_1(.dout(w_dff_A_dXhCYzvS6_1),.din(w_dff_A_LKBQMA7Q4_1),.clk(gclk));
	jdff dff_A_VuZYIoto5_2(.dout(w_G45_0[2]),.din(w_dff_A_VuZYIoto5_2),.clk(gclk));
	jdff dff_A_QYvsE2TM0_2(.dout(w_dff_A_VuZYIoto5_2),.din(w_dff_A_QYvsE2TM0_2),.clk(gclk));
	jdff dff_A_zXJtZd5W5_2(.dout(w_dff_A_QYvsE2TM0_2),.din(w_dff_A_zXJtZd5W5_2),.clk(gclk));
	jdff dff_A_BhSiJ9au1_0(.dout(w_n98_1[0]),.din(w_dff_A_BhSiJ9au1_0),.clk(gclk));
	jdff dff_A_Kgb8rgQL7_1(.dout(w_n98_1[1]),.din(w_dff_A_Kgb8rgQL7_1),.clk(gclk));
	jdff dff_A_QsEFNNHz1_0(.dout(w_G250_0[0]),.din(w_dff_A_QsEFNNHz1_0),.clk(gclk));
	jdff dff_A_g1sQxtI67_0(.dout(w_dff_A_QsEFNNHz1_0),.din(w_dff_A_g1sQxtI67_0),.clk(gclk));
	jdff dff_A_HHFWPCEd1_1(.dout(w_G250_0[1]),.din(w_dff_A_HHFWPCEd1_1),.clk(gclk));
	jdff dff_A_Pf8WR8ke6_1(.dout(w_dff_A_HHFWPCEd1_1),.din(w_dff_A_Pf8WR8ke6_1),.clk(gclk));
	jdff dff_B_rwCQmGns8_1(.din(n153),.dout(w_dff_B_rwCQmGns8_1),.clk(gclk));
	jdff dff_A_XmqvYvIZ1_0(.dout(w_n157_0[0]),.din(w_dff_A_XmqvYvIZ1_0),.clk(gclk));
	jdff dff_A_0vFtVP2w7_0(.dout(w_dff_A_XmqvYvIZ1_0),.din(w_dff_A_0vFtVP2w7_0),.clk(gclk));
	jdff dff_A_tiDUSUyz2_2(.dout(w_n157_0[2]),.din(w_dff_A_tiDUSUyz2_2),.clk(gclk));
	jdff dff_A_wPVodFzS2_2(.dout(w_dff_A_tiDUSUyz2_2),.din(w_dff_A_wPVodFzS2_2),.clk(gclk));
	jdff dff_A_m9AQBAfc0_1(.dout(w_G116_1[1]),.din(w_dff_A_m9AQBAfc0_1),.clk(gclk));
	jdff dff_A_yrtdOxd48_1(.dout(w_dff_A_m9AQBAfc0_1),.din(w_dff_A_yrtdOxd48_1),.clk(gclk));
	jdff dff_A_NaGJkzdY8_1(.dout(w_dff_A_yrtdOxd48_1),.din(w_dff_A_NaGJkzdY8_1),.clk(gclk));
	jdff dff_A_VMQDtKWt8_2(.dout(w_G116_1[2]),.din(w_dff_A_VMQDtKWt8_2),.clk(gclk));
	jdff dff_A_wIbuJ4LX4_2(.dout(w_dff_A_VMQDtKWt8_2),.din(w_dff_A_wIbuJ4LX4_2),.clk(gclk));
	jdff dff_A_kEIBVVPy7_2(.dout(w_dff_A_wIbuJ4LX4_2),.din(w_dff_A_kEIBVVPy7_2),.clk(gclk));
	jdff dff_A_WYs0vfay0_1(.dout(w_G116_0[1]),.din(w_dff_A_WYs0vfay0_1),.clk(gclk));
	jdff dff_A_nPtrMTIV5_1(.dout(w_dff_A_WYs0vfay0_1),.din(w_dff_A_nPtrMTIV5_1),.clk(gclk));
	jdff dff_A_xBne4DBd4_1(.dout(w_dff_A_nPtrMTIV5_1),.din(w_dff_A_xBne4DBd4_1),.clk(gclk));
	jdff dff_A_ck8EZlDh9_2(.dout(w_G116_0[2]),.din(w_dff_A_ck8EZlDh9_2),.clk(gclk));
	jdff dff_A_kOAxi8ve7_0(.dout(w_G238_1[0]),.din(w_dff_A_kOAxi8ve7_0),.clk(gclk));
	jdff dff_A_lN1JJFlD5_0(.dout(w_dff_A_kOAxi8ve7_0),.din(w_dff_A_lN1JJFlD5_0),.clk(gclk));
	jdff dff_A_k6eV8qlH9_1(.dout(w_G238_0[1]),.din(w_dff_A_k6eV8qlH9_1),.clk(gclk));
	jdff dff_A_nxMrEFUv2_1(.dout(w_dff_A_k6eV8qlH9_1),.din(w_dff_A_nxMrEFUv2_1),.clk(gclk));
	jdff dff_A_cHbsuxtE2_1(.dout(w_dff_A_nxMrEFUv2_1),.din(w_dff_A_cHbsuxtE2_1),.clk(gclk));
	jdff dff_A_ygpYplsT6_1(.dout(w_dff_A_cHbsuxtE2_1),.din(w_dff_A_ygpYplsT6_1),.clk(gclk));
	jdff dff_A_QvNaOfpl1_2(.dout(w_G238_0[2]),.din(w_dff_A_QvNaOfpl1_2),.clk(gclk));
	jdff dff_A_71vYR1RX5_2(.dout(w_dff_A_QvNaOfpl1_2),.din(w_dff_A_71vYR1RX5_2),.clk(gclk));
	jdff dff_A_Cc3xYaea6_2(.dout(w_G1698_0[2]),.din(w_dff_A_Cc3xYaea6_2),.clk(gclk));
	jdff dff_A_DghhoA0d2_0(.dout(w_G244_1[0]),.din(w_dff_A_DghhoA0d2_0),.clk(gclk));
	jdff dff_A_z9ZgqKo90_0(.dout(w_dff_A_DghhoA0d2_0),.din(w_dff_A_z9ZgqKo90_0),.clk(gclk));
	jdff dff_A_pyR7l0nS8_1(.dout(w_G244_0[1]),.din(w_dff_A_pyR7l0nS8_1),.clk(gclk));
	jdff dff_A_UaOFlXuZ9_1(.dout(w_dff_A_pyR7l0nS8_1),.din(w_dff_A_UaOFlXuZ9_1),.clk(gclk));
	jdff dff_A_vFYBr6sJ7_1(.dout(w_dff_A_UaOFlXuZ9_1),.din(w_dff_A_vFYBr6sJ7_1),.clk(gclk));
	jdff dff_A_xklEYXbG0_1(.dout(w_dff_A_vFYBr6sJ7_1),.din(w_dff_A_xklEYXbG0_1),.clk(gclk));
	jdff dff_A_AXuFwqn41_2(.dout(w_G244_0[2]),.din(w_dff_A_AXuFwqn41_2),.clk(gclk));
	jdff dff_A_ppap3l3i7_2(.dout(w_dff_A_AXuFwqn41_2),.din(w_dff_A_ppap3l3i7_2),.clk(gclk));
	jdff dff_A_RXzNqvLP6_2(.dout(w_n151_4[2]),.din(w_dff_A_RXzNqvLP6_2),.clk(gclk));
	jdff dff_A_YpwrCHtT1_2(.dout(w_dff_A_RXzNqvLP6_2),.din(w_dff_A_YpwrCHtT1_2),.clk(gclk));
	jdff dff_A_0uRYzCfa2_1(.dout(w_n151_1[1]),.din(w_dff_A_0uRYzCfa2_1),.clk(gclk));
	jdff dff_A_3G10Qk7Z1_1(.dout(w_dff_A_0uRYzCfa2_1),.din(w_dff_A_3G10Qk7Z1_1),.clk(gclk));
	jdff dff_A_iWfDf8LR3_2(.dout(w_n151_1[2]),.din(w_dff_A_iWfDf8LR3_2),.clk(gclk));
	jdff dff_A_MFQzdhd58_2(.dout(w_dff_A_iWfDf8LR3_2),.din(w_dff_A_MFQzdhd58_2),.clk(gclk));
	jdff dff_A_Dp18gep98_1(.dout(w_n151_0[1]),.din(w_dff_A_Dp18gep98_1),.clk(gclk));
	jdff dff_A_HThULbC84_1(.dout(w_dff_A_Dp18gep98_1),.din(w_dff_A_HThULbC84_1),.clk(gclk));
	jdff dff_A_F456LDT18_0(.dout(w_n149_2[0]),.din(w_dff_A_F456LDT18_0),.clk(gclk));
	jdff dff_A_Wo6mhXIz9_1(.dout(w_G41_0[1]),.din(w_dff_A_Wo6mhXIz9_1),.clk(gclk));
	jdff dff_A_RKU5LgTY8_2(.dout(w_G41_0[2]),.din(w_dff_A_RKU5LgTY8_2),.clk(gclk));
	jdff dff_A_EE6LrMLh2_2(.dout(w_dff_A_RKU5LgTY8_2),.din(w_dff_A_EE6LrMLh2_2),.clk(gclk));
	jdff dff_A_3Vq1cj8a2_2(.dout(w_G33_3[2]),.din(w_dff_A_3Vq1cj8a2_2),.clk(gclk));
	jdff dff_A_aYuOSGG61_2(.dout(w_dff_A_3Vq1cj8a2_2),.din(w_dff_A_aYuOSGG61_2),.clk(gclk));
	jdff dff_A_1sYSLJKw4_2(.dout(w_dff_A_aYuOSGG61_2),.din(w_dff_A_1sYSLJKw4_2),.clk(gclk));
	jdff dff_A_euNSTRCr8_2(.dout(w_dff_A_1sYSLJKw4_2),.din(w_dff_A_euNSTRCr8_2),.clk(gclk));
	jdff dff_A_GKmywLFy8_2(.dout(w_dff_A_euNSTRCr8_2),.din(w_dff_A_GKmywLFy8_2),.clk(gclk));
	jdff dff_A_6zatj6M01_0(.dout(w_G33_0[0]),.din(w_dff_A_6zatj6M01_0),.clk(gclk));
	jdff dff_A_7tAftBDu2_1(.dout(w_n147_0[1]),.din(w_dff_A_7tAftBDu2_1),.clk(gclk));
	jdff dff_A_9AnwOYgO0_2(.dout(w_n147_0[2]),.din(w_dff_A_9AnwOYgO0_2),.clk(gclk));
	jdff dff_A_pi8XySmV6_1(.dout(w_G13_0[1]),.din(w_dff_A_pi8XySmV6_1),.clk(gclk));
	jdff dff_A_EsjesbNK5_2(.dout(w_G13_0[2]),.din(w_dff_A_EsjesbNK5_2),.clk(gclk));
	jdff dff_A_DlJf6hDJ7_2(.dout(w_dff_A_EsjesbNK5_2),.din(w_dff_A_DlJf6hDJ7_2),.clk(gclk));
	jdff dff_A_X0OT3Diz9_0(.dout(w_G1_2[0]),.din(w_dff_A_X0OT3Diz9_0),.clk(gclk));
	jdff dff_A_X0OpRtEZ5_2(.dout(w_G1_2[2]),.din(w_dff_A_X0OpRtEZ5_2),.clk(gclk));
	jdff dff_A_pjgwWpzJ1_0(.dout(w_G1_0[0]),.din(w_dff_A_pjgwWpzJ1_0),.clk(gclk));
	jdff dff_A_3ji1y7E47_1(.dout(w_n146_0[1]),.din(w_dff_A_3ji1y7E47_1),.clk(gclk));
	jdff dff_A_SvNwvbPR2_1(.dout(w_dff_A_3ji1y7E47_1),.din(w_dff_A_SvNwvbPR2_1),.clk(gclk));
	jdff dff_A_9d0Oyzz15_1(.dout(w_dff_A_SvNwvbPR2_1),.din(w_dff_A_9d0Oyzz15_1),.clk(gclk));
	jdff dff_A_jB4hXWJ21_1(.dout(w_dff_A_9d0Oyzz15_1),.din(w_dff_A_jB4hXWJ21_1),.clk(gclk));
	jdff dff_A_TYEQOXSd2_1(.dout(w_dff_A_jB4hXWJ21_1),.din(w_dff_A_TYEQOXSd2_1),.clk(gclk));
	jdff dff_A_nLw5oAua9_1(.dout(w_dff_A_TYEQOXSd2_1),.din(w_dff_A_nLw5oAua9_1),.clk(gclk));
	jdff dff_A_N37N5do51_2(.dout(w_n146_0[2]),.din(w_dff_A_N37N5do51_2),.clk(gclk));
	jdff dff_A_YnphOlLj9_2(.dout(w_dff_A_N37N5do51_2),.din(w_dff_A_YnphOlLj9_2),.clk(gclk));
	jdff dff_A_iOPizZua7_2(.dout(w_dff_A_YnphOlLj9_2),.din(w_dff_A_iOPizZua7_2),.clk(gclk));
	jdff dff_A_XnwGzwWC9_2(.dout(w_dff_A_iOPizZua7_2),.din(w_dff_A_XnwGzwWC9_2),.clk(gclk));
	jdff dff_A_DJD2xBfu6_2(.dout(w_dff_A_XnwGzwWC9_2),.din(w_dff_A_DJD2xBfu6_2),.clk(gclk));
	jdff dff_A_7t4Mkimw9_2(.dout(w_dff_A_DJD2xBfu6_2),.din(w_dff_A_7t4Mkimw9_2),.clk(gclk));
	jdff dff_A_ecrH86MZ3_0(.dout(w_G169_1[0]),.din(w_dff_A_ecrH86MZ3_0),.clk(gclk));
	jdff dff_A_CIUS7Gav5_0(.dout(w_dff_A_ecrH86MZ3_0),.din(w_dff_A_CIUS7Gav5_0),.clk(gclk));
	jdff dff_A_N15nrHCM4_0(.dout(w_dff_A_CIUS7Gav5_0),.din(w_dff_A_N15nrHCM4_0),.clk(gclk));
	jdff dff_A_hN2WiKWB3_0(.dout(w_dff_A_N15nrHCM4_0),.din(w_dff_A_hN2WiKWB3_0),.clk(gclk));
	jdff dff_A_E2uRmedZ7_0(.dout(w_dff_A_hN2WiKWB3_0),.din(w_dff_A_E2uRmedZ7_0),.clk(gclk));
	jdff dff_A_RNPboyHt6_0(.dout(w_dff_A_E2uRmedZ7_0),.din(w_dff_A_RNPboyHt6_0),.clk(gclk));
	jdff dff_A_5SRtP6CE7_0(.dout(w_dff_A_RNPboyHt6_0),.din(w_dff_A_5SRtP6CE7_0),.clk(gclk));
	jdff dff_A_oYAU9c182_1(.dout(w_G169_0[1]),.din(w_dff_A_oYAU9c182_1),.clk(gclk));
	jdff dff_A_9gtS7jRs7_1(.dout(w_dff_A_oYAU9c182_1),.din(w_dff_A_9gtS7jRs7_1),.clk(gclk));
	jdff dff_A_kOz5WkqB0_1(.dout(w_dff_A_9gtS7jRs7_1),.din(w_dff_A_kOz5WkqB0_1),.clk(gclk));
	jdff dff_A_KNOXphIj4_1(.dout(w_dff_A_kOz5WkqB0_1),.din(w_dff_A_KNOXphIj4_1),.clk(gclk));
	jdff dff_A_9Yn9EafO9_1(.dout(w_dff_A_KNOXphIj4_1),.din(w_dff_A_9Yn9EafO9_1),.clk(gclk));
	jdff dff_A_ms5jV2pR2_1(.dout(w_dff_A_9Yn9EafO9_1),.din(w_dff_A_ms5jV2pR2_1),.clk(gclk));
	jdff dff_A_5ltwZ2ye2_1(.dout(w_dff_A_ms5jV2pR2_1),.din(w_dff_A_5ltwZ2ye2_1),.clk(gclk));
	jdff dff_A_Lt7Qfty51_2(.dout(w_G169_0[2]),.din(w_dff_A_Lt7Qfty51_2),.clk(gclk));
	jdff dff_A_e0zbmbUP5_2(.dout(w_dff_A_Lt7Qfty51_2),.din(w_dff_A_e0zbmbUP5_2),.clk(gclk));
	jdff dff_A_Q7INts5y4_2(.dout(w_dff_A_e0zbmbUP5_2),.din(w_dff_A_Q7INts5y4_2),.clk(gclk));
	jdff dff_A_VyNIVmih6_2(.dout(w_dff_A_Q7INts5y4_2),.din(w_dff_A_VyNIVmih6_2),.clk(gclk));
	jdff dff_A_K4nfzJYu7_2(.dout(w_dff_A_VyNIVmih6_2),.din(w_dff_A_K4nfzJYu7_2),.clk(gclk));
	jdff dff_A_mo6qCbGr2_2(.dout(w_dff_A_K4nfzJYu7_2),.din(w_dff_A_mo6qCbGr2_2),.clk(gclk));
	jdff dff_A_vkYHzYam5_2(.dout(w_dff_A_mo6qCbGr2_2),.din(w_dff_A_vkYHzYam5_2),.clk(gclk));
	jdff dff_A_BaeaEVsM2_2(.dout(w_dff_A_XgtW6qji8_0),.din(w_dff_A_BaeaEVsM2_2),.clk(gclk));
	jdff dff_A_XgtW6qji8_0(.dout(w_dff_A_JpAMYWHg4_0),.din(w_dff_A_XgtW6qji8_0),.clk(gclk));
	jdff dff_A_JpAMYWHg4_0(.dout(w_dff_A_qEcFQfSS3_0),.din(w_dff_A_JpAMYWHg4_0),.clk(gclk));
	jdff dff_A_qEcFQfSS3_0(.dout(w_dff_A_ic3agfWW8_0),.din(w_dff_A_qEcFQfSS3_0),.clk(gclk));
	jdff dff_A_ic3agfWW8_0(.dout(w_dff_A_5YXSH2j93_0),.din(w_dff_A_ic3agfWW8_0),.clk(gclk));
	jdff dff_A_5YXSH2j93_0(.dout(w_dff_A_mWGi77gq4_0),.din(w_dff_A_5YXSH2j93_0),.clk(gclk));
	jdff dff_A_mWGi77gq4_0(.dout(w_dff_A_YapfiCWH5_0),.din(w_dff_A_mWGi77gq4_0),.clk(gclk));
	jdff dff_A_YapfiCWH5_0(.dout(w_dff_A_RuDMLY429_0),.din(w_dff_A_YapfiCWH5_0),.clk(gclk));
	jdff dff_A_RuDMLY429_0(.dout(w_dff_A_rvHqpQg65_0),.din(w_dff_A_RuDMLY429_0),.clk(gclk));
	jdff dff_A_rvHqpQg65_0(.dout(w_dff_A_tVYmYUbc7_0),.din(w_dff_A_rvHqpQg65_0),.clk(gclk));
	jdff dff_A_tVYmYUbc7_0(.dout(w_dff_A_6tRvnHb68_0),.din(w_dff_A_tVYmYUbc7_0),.clk(gclk));
	jdff dff_A_6tRvnHb68_0(.dout(w_dff_A_zr3ABjfk5_0),.din(w_dff_A_6tRvnHb68_0),.clk(gclk));
	jdff dff_A_zr3ABjfk5_0(.dout(w_dff_A_VX4ll8OB7_0),.din(w_dff_A_zr3ABjfk5_0),.clk(gclk));
	jdff dff_A_VX4ll8OB7_0(.dout(w_dff_A_SjsoBwiK5_0),.din(w_dff_A_VX4ll8OB7_0),.clk(gclk));
	jdff dff_A_SjsoBwiK5_0(.dout(w_dff_A_n03ppBW46_0),.din(w_dff_A_SjsoBwiK5_0),.clk(gclk));
	jdff dff_A_n03ppBW46_0(.dout(w_dff_A_MlGXvFTp3_0),.din(w_dff_A_n03ppBW46_0),.clk(gclk));
	jdff dff_A_MlGXvFTp3_0(.dout(w_dff_A_YFvttSyB0_0),.din(w_dff_A_MlGXvFTp3_0),.clk(gclk));
	jdff dff_A_YFvttSyB0_0(.dout(w_dff_A_nhOyjTGc7_0),.din(w_dff_A_YFvttSyB0_0),.clk(gclk));
	jdff dff_A_nhOyjTGc7_0(.dout(w_dff_A_fKUsN38t3_0),.din(w_dff_A_nhOyjTGc7_0),.clk(gclk));
	jdff dff_A_fKUsN38t3_0(.dout(w_dff_A_BEZMkJS57_0),.din(w_dff_A_fKUsN38t3_0),.clk(gclk));
	jdff dff_A_BEZMkJS57_0(.dout(w_dff_A_G3Xvkq2P1_0),.din(w_dff_A_BEZMkJS57_0),.clk(gclk));
	jdff dff_A_G3Xvkq2P1_0(.dout(w_dff_A_mwAJJ9ZA1_0),.din(w_dff_A_G3Xvkq2P1_0),.clk(gclk));
	jdff dff_A_mwAJJ9ZA1_0(.dout(w_dff_A_DfmZ2fx43_0),.din(w_dff_A_mwAJJ9ZA1_0),.clk(gclk));
	jdff dff_A_DfmZ2fx43_0(.dout(w_dff_A_zeiEugJd5_0),.din(w_dff_A_DfmZ2fx43_0),.clk(gclk));
	jdff dff_A_zeiEugJd5_0(.dout(G353),.din(w_dff_A_zeiEugJd5_0),.clk(gclk));
	jdff dff_A_D1cH4P2b3_1(.dout(w_dff_A_lymXg1rU4_0),.din(w_dff_A_D1cH4P2b3_1),.clk(gclk));
	jdff dff_A_lymXg1rU4_0(.dout(w_dff_A_qVXL5q4A7_0),.din(w_dff_A_lymXg1rU4_0),.clk(gclk));
	jdff dff_A_qVXL5q4A7_0(.dout(w_dff_A_zTTihcWl2_0),.din(w_dff_A_qVXL5q4A7_0),.clk(gclk));
	jdff dff_A_zTTihcWl2_0(.dout(w_dff_A_7ofWyn2G2_0),.din(w_dff_A_zTTihcWl2_0),.clk(gclk));
	jdff dff_A_7ofWyn2G2_0(.dout(w_dff_A_uprW2tFx8_0),.din(w_dff_A_7ofWyn2G2_0),.clk(gclk));
	jdff dff_A_uprW2tFx8_0(.dout(w_dff_A_IjpJGnU97_0),.din(w_dff_A_uprW2tFx8_0),.clk(gclk));
	jdff dff_A_IjpJGnU97_0(.dout(w_dff_A_q5DJKGA85_0),.din(w_dff_A_IjpJGnU97_0),.clk(gclk));
	jdff dff_A_q5DJKGA85_0(.dout(w_dff_A_Q8i2HS3Z9_0),.din(w_dff_A_q5DJKGA85_0),.clk(gclk));
	jdff dff_A_Q8i2HS3Z9_0(.dout(w_dff_A_IkOcXU3g5_0),.din(w_dff_A_Q8i2HS3Z9_0),.clk(gclk));
	jdff dff_A_IkOcXU3g5_0(.dout(w_dff_A_ktK1BNft1_0),.din(w_dff_A_IkOcXU3g5_0),.clk(gclk));
	jdff dff_A_ktK1BNft1_0(.dout(w_dff_A_FfhpUuu83_0),.din(w_dff_A_ktK1BNft1_0),.clk(gclk));
	jdff dff_A_FfhpUuu83_0(.dout(w_dff_A_tRfRM30g0_0),.din(w_dff_A_FfhpUuu83_0),.clk(gclk));
	jdff dff_A_tRfRM30g0_0(.dout(w_dff_A_vjNtIkT79_0),.din(w_dff_A_tRfRM30g0_0),.clk(gclk));
	jdff dff_A_vjNtIkT79_0(.dout(w_dff_A_q70ixND62_0),.din(w_dff_A_vjNtIkT79_0),.clk(gclk));
	jdff dff_A_q70ixND62_0(.dout(w_dff_A_XcsLJeh18_0),.din(w_dff_A_q70ixND62_0),.clk(gclk));
	jdff dff_A_XcsLJeh18_0(.dout(w_dff_A_YEJIxoIy0_0),.din(w_dff_A_XcsLJeh18_0),.clk(gclk));
	jdff dff_A_YEJIxoIy0_0(.dout(w_dff_A_z38LIswg3_0),.din(w_dff_A_YEJIxoIy0_0),.clk(gclk));
	jdff dff_A_z38LIswg3_0(.dout(w_dff_A_LNiISBmP2_0),.din(w_dff_A_z38LIswg3_0),.clk(gclk));
	jdff dff_A_LNiISBmP2_0(.dout(w_dff_A_Etbi6mcC9_0),.din(w_dff_A_LNiISBmP2_0),.clk(gclk));
	jdff dff_A_Etbi6mcC9_0(.dout(w_dff_A_H922DeuZ8_0),.din(w_dff_A_Etbi6mcC9_0),.clk(gclk));
	jdff dff_A_H922DeuZ8_0(.dout(w_dff_A_ZeJnYqn39_0),.din(w_dff_A_H922DeuZ8_0),.clk(gclk));
	jdff dff_A_ZeJnYqn39_0(.dout(w_dff_A_oA6LAxVK4_0),.din(w_dff_A_ZeJnYqn39_0),.clk(gclk));
	jdff dff_A_oA6LAxVK4_0(.dout(w_dff_A_VcUXKZc98_0),.din(w_dff_A_oA6LAxVK4_0),.clk(gclk));
	jdff dff_A_VcUXKZc98_0(.dout(G355),.din(w_dff_A_VcUXKZc98_0),.clk(gclk));
	jdff dff_A_ZYKz2ojx0_2(.dout(w_dff_A_MAt5EeXn0_0),.din(w_dff_A_ZYKz2ojx0_2),.clk(gclk));
	jdff dff_A_MAt5EeXn0_0(.dout(w_dff_A_Seo4hX7x7_0),.din(w_dff_A_MAt5EeXn0_0),.clk(gclk));
	jdff dff_A_Seo4hX7x7_0(.dout(w_dff_A_k6NaR4C44_0),.din(w_dff_A_Seo4hX7x7_0),.clk(gclk));
	jdff dff_A_k6NaR4C44_0(.dout(w_dff_A_V4yQwgQX0_0),.din(w_dff_A_k6NaR4C44_0),.clk(gclk));
	jdff dff_A_V4yQwgQX0_0(.dout(w_dff_A_d0MVzWK97_0),.din(w_dff_A_V4yQwgQX0_0),.clk(gclk));
	jdff dff_A_d0MVzWK97_0(.dout(w_dff_A_0RpYHYl57_0),.din(w_dff_A_d0MVzWK97_0),.clk(gclk));
	jdff dff_A_0RpYHYl57_0(.dout(w_dff_A_JKHJmjux9_0),.din(w_dff_A_0RpYHYl57_0),.clk(gclk));
	jdff dff_A_JKHJmjux9_0(.dout(w_dff_A_IMs5XXbX2_0),.din(w_dff_A_JKHJmjux9_0),.clk(gclk));
	jdff dff_A_IMs5XXbX2_0(.dout(w_dff_A_Oep19O2I7_0),.din(w_dff_A_IMs5XXbX2_0),.clk(gclk));
	jdff dff_A_Oep19O2I7_0(.dout(w_dff_A_N6eXX0fK0_0),.din(w_dff_A_Oep19O2I7_0),.clk(gclk));
	jdff dff_A_N6eXX0fK0_0(.dout(w_dff_A_8RXTpRqG7_0),.din(w_dff_A_N6eXX0fK0_0),.clk(gclk));
	jdff dff_A_8RXTpRqG7_0(.dout(w_dff_A_65zzfM8Q4_0),.din(w_dff_A_8RXTpRqG7_0),.clk(gclk));
	jdff dff_A_65zzfM8Q4_0(.dout(w_dff_A_8bIyJC0G2_0),.din(w_dff_A_65zzfM8Q4_0),.clk(gclk));
	jdff dff_A_8bIyJC0G2_0(.dout(w_dff_A_rIsbS6QB5_0),.din(w_dff_A_8bIyJC0G2_0),.clk(gclk));
	jdff dff_A_rIsbS6QB5_0(.dout(w_dff_A_0A1jKdQI8_0),.din(w_dff_A_rIsbS6QB5_0),.clk(gclk));
	jdff dff_A_0A1jKdQI8_0(.dout(w_dff_A_zRU7muaP3_0),.din(w_dff_A_0A1jKdQI8_0),.clk(gclk));
	jdff dff_A_zRU7muaP3_0(.dout(w_dff_A_ewYtief36_0),.din(w_dff_A_zRU7muaP3_0),.clk(gclk));
	jdff dff_A_ewYtief36_0(.dout(w_dff_A_unEFxqqU1_0),.din(w_dff_A_ewYtief36_0),.clk(gclk));
	jdff dff_A_unEFxqqU1_0(.dout(w_dff_A_oOPWcNbr2_0),.din(w_dff_A_unEFxqqU1_0),.clk(gclk));
	jdff dff_A_oOPWcNbr2_0(.dout(w_dff_A_w0LqHfb65_0),.din(w_dff_A_oOPWcNbr2_0),.clk(gclk));
	jdff dff_A_w0LqHfb65_0(.dout(G361),.din(w_dff_A_w0LqHfb65_0),.clk(gclk));
	jdff dff_A_c5kn6LU27_2(.dout(w_dff_A_xSALYtp61_0),.din(w_dff_A_c5kn6LU27_2),.clk(gclk));
	jdff dff_A_xSALYtp61_0(.dout(w_dff_A_56wXPuXI2_0),.din(w_dff_A_xSALYtp61_0),.clk(gclk));
	jdff dff_A_56wXPuXI2_0(.dout(w_dff_A_ihb6mLs17_0),.din(w_dff_A_56wXPuXI2_0),.clk(gclk));
	jdff dff_A_ihb6mLs17_0(.dout(w_dff_A_QVzgLuCv6_0),.din(w_dff_A_ihb6mLs17_0),.clk(gclk));
	jdff dff_A_QVzgLuCv6_0(.dout(w_dff_A_MDTFNVlg6_0),.din(w_dff_A_QVzgLuCv6_0),.clk(gclk));
	jdff dff_A_MDTFNVlg6_0(.dout(w_dff_A_tAWKkV5u1_0),.din(w_dff_A_MDTFNVlg6_0),.clk(gclk));
	jdff dff_A_tAWKkV5u1_0(.dout(w_dff_A_VA54F3DT2_0),.din(w_dff_A_tAWKkV5u1_0),.clk(gclk));
	jdff dff_A_VA54F3DT2_0(.dout(w_dff_A_4tCAIW6u7_0),.din(w_dff_A_VA54F3DT2_0),.clk(gclk));
	jdff dff_A_4tCAIW6u7_0(.dout(w_dff_A_D68iNJyj2_0),.din(w_dff_A_4tCAIW6u7_0),.clk(gclk));
	jdff dff_A_D68iNJyj2_0(.dout(w_dff_A_upEdZ1dj3_0),.din(w_dff_A_D68iNJyj2_0),.clk(gclk));
	jdff dff_A_upEdZ1dj3_0(.dout(w_dff_A_07hJC3vz0_0),.din(w_dff_A_upEdZ1dj3_0),.clk(gclk));
	jdff dff_A_07hJC3vz0_0(.dout(w_dff_A_0oCyMF9c1_0),.din(w_dff_A_07hJC3vz0_0),.clk(gclk));
	jdff dff_A_0oCyMF9c1_0(.dout(w_dff_A_u3tYelhM2_0),.din(w_dff_A_0oCyMF9c1_0),.clk(gclk));
	jdff dff_A_u3tYelhM2_0(.dout(w_dff_A_XhLoKl765_0),.din(w_dff_A_u3tYelhM2_0),.clk(gclk));
	jdff dff_A_XhLoKl765_0(.dout(w_dff_A_8oeRjjOv6_0),.din(w_dff_A_XhLoKl765_0),.clk(gclk));
	jdff dff_A_8oeRjjOv6_0(.dout(w_dff_A_Kw1uMcA16_0),.din(w_dff_A_8oeRjjOv6_0),.clk(gclk));
	jdff dff_A_Kw1uMcA16_0(.dout(w_dff_A_cm0DJlYr7_0),.din(w_dff_A_Kw1uMcA16_0),.clk(gclk));
	jdff dff_A_cm0DJlYr7_0(.dout(w_dff_A_lWjHae9i7_0),.din(w_dff_A_cm0DJlYr7_0),.clk(gclk));
	jdff dff_A_lWjHae9i7_0(.dout(w_dff_A_U4l3J0JQ7_0),.din(w_dff_A_lWjHae9i7_0),.clk(gclk));
	jdff dff_A_U4l3J0JQ7_0(.dout(w_dff_A_87c0mXR40_0),.din(w_dff_A_U4l3J0JQ7_0),.clk(gclk));
	jdff dff_A_87c0mXR40_0(.dout(w_dff_A_py3qjAlO6_0),.din(w_dff_A_87c0mXR40_0),.clk(gclk));
	jdff dff_A_py3qjAlO6_0(.dout(w_dff_A_8lkpG9yj5_0),.din(w_dff_A_py3qjAlO6_0),.clk(gclk));
	jdff dff_A_8lkpG9yj5_0(.dout(w_dff_A_CvdrDH3z9_0),.din(w_dff_A_8lkpG9yj5_0),.clk(gclk));
	jdff dff_A_CvdrDH3z9_0(.dout(G358),.din(w_dff_A_CvdrDH3z9_0),.clk(gclk));
	jdff dff_A_mPRw3Kex9_2(.dout(w_dff_A_y1Q6LEgZ9_0),.din(w_dff_A_mPRw3Kex9_2),.clk(gclk));
	jdff dff_A_y1Q6LEgZ9_0(.dout(w_dff_A_p1bPyM9u7_0),.din(w_dff_A_y1Q6LEgZ9_0),.clk(gclk));
	jdff dff_A_p1bPyM9u7_0(.dout(w_dff_A_rbSnQTIY6_0),.din(w_dff_A_p1bPyM9u7_0),.clk(gclk));
	jdff dff_A_rbSnQTIY6_0(.dout(w_dff_A_i3upuMjk4_0),.din(w_dff_A_rbSnQTIY6_0),.clk(gclk));
	jdff dff_A_i3upuMjk4_0(.dout(w_dff_A_UR7UTR4p5_0),.din(w_dff_A_i3upuMjk4_0),.clk(gclk));
	jdff dff_A_UR7UTR4p5_0(.dout(w_dff_A_0u8mcTUR9_0),.din(w_dff_A_UR7UTR4p5_0),.clk(gclk));
	jdff dff_A_0u8mcTUR9_0(.dout(w_dff_A_p4ScEj226_0),.din(w_dff_A_0u8mcTUR9_0),.clk(gclk));
	jdff dff_A_p4ScEj226_0(.dout(w_dff_A_jdihPNqz1_0),.din(w_dff_A_p4ScEj226_0),.clk(gclk));
	jdff dff_A_jdihPNqz1_0(.dout(w_dff_A_h2Cz38b28_0),.din(w_dff_A_jdihPNqz1_0),.clk(gclk));
	jdff dff_A_h2Cz38b28_0(.dout(w_dff_A_GKAkkJ7B6_0),.din(w_dff_A_h2Cz38b28_0),.clk(gclk));
	jdff dff_A_GKAkkJ7B6_0(.dout(w_dff_A_jJa7iNCX4_0),.din(w_dff_A_GKAkkJ7B6_0),.clk(gclk));
	jdff dff_A_jJa7iNCX4_0(.dout(w_dff_A_618NVufX0_0),.din(w_dff_A_jJa7iNCX4_0),.clk(gclk));
	jdff dff_A_618NVufX0_0(.dout(w_dff_A_SLEXvMko7_0),.din(w_dff_A_618NVufX0_0),.clk(gclk));
	jdff dff_A_SLEXvMko7_0(.dout(w_dff_A_I20KqZEp7_0),.din(w_dff_A_SLEXvMko7_0),.clk(gclk));
	jdff dff_A_I20KqZEp7_0(.dout(w_dff_A_kh6Uzcp47_0),.din(w_dff_A_I20KqZEp7_0),.clk(gclk));
	jdff dff_A_kh6Uzcp47_0(.dout(w_dff_A_B59Nuf1J2_0),.din(w_dff_A_kh6Uzcp47_0),.clk(gclk));
	jdff dff_A_B59Nuf1J2_0(.dout(w_dff_A_oAY020Le8_0),.din(w_dff_A_B59Nuf1J2_0),.clk(gclk));
	jdff dff_A_oAY020Le8_0(.dout(w_dff_A_2ALw7X1a9_0),.din(w_dff_A_oAY020Le8_0),.clk(gclk));
	jdff dff_A_2ALw7X1a9_0(.dout(w_dff_A_pStHHbCW0_0),.din(w_dff_A_2ALw7X1a9_0),.clk(gclk));
	jdff dff_A_pStHHbCW0_0(.dout(w_dff_A_8x7lEdjR2_0),.din(w_dff_A_pStHHbCW0_0),.clk(gclk));
	jdff dff_A_8x7lEdjR2_0(.dout(w_dff_A_8f0RZSV56_0),.din(w_dff_A_8x7lEdjR2_0),.clk(gclk));
	jdff dff_A_8f0RZSV56_0(.dout(w_dff_A_SvdPApWS4_0),.din(w_dff_A_8f0RZSV56_0),.clk(gclk));
	jdff dff_A_SvdPApWS4_0(.dout(w_dff_A_6ONkQnMn0_0),.din(w_dff_A_SvdPApWS4_0),.clk(gclk));
	jdff dff_A_6ONkQnMn0_0(.dout(G351),.din(w_dff_A_6ONkQnMn0_0),.clk(gclk));
	jdff dff_A_FbzfaOjn5_2(.dout(w_dff_A_KzvB2uNu4_0),.din(w_dff_A_FbzfaOjn5_2),.clk(gclk));
	jdff dff_A_KzvB2uNu4_0(.dout(w_dff_A_xWbtP3id0_0),.din(w_dff_A_KzvB2uNu4_0),.clk(gclk));
	jdff dff_A_xWbtP3id0_0(.dout(w_dff_A_pTl5v5kN3_0),.din(w_dff_A_xWbtP3id0_0),.clk(gclk));
	jdff dff_A_pTl5v5kN3_0(.dout(w_dff_A_3TPtL5WN2_0),.din(w_dff_A_pTl5v5kN3_0),.clk(gclk));
	jdff dff_A_3TPtL5WN2_0(.dout(w_dff_A_I48EkiSa1_0),.din(w_dff_A_3TPtL5WN2_0),.clk(gclk));
	jdff dff_A_I48EkiSa1_0(.dout(w_dff_A_yTLimDf87_0),.din(w_dff_A_I48EkiSa1_0),.clk(gclk));
	jdff dff_A_yTLimDf87_0(.dout(w_dff_A_PNAbjEge8_0),.din(w_dff_A_yTLimDf87_0),.clk(gclk));
	jdff dff_A_PNAbjEge8_0(.dout(w_dff_A_dpNyKKEl7_0),.din(w_dff_A_PNAbjEge8_0),.clk(gclk));
	jdff dff_A_dpNyKKEl7_0(.dout(w_dff_A_cp4P7mBH1_0),.din(w_dff_A_dpNyKKEl7_0),.clk(gclk));
	jdff dff_A_cp4P7mBH1_0(.dout(w_dff_A_mygSIe9a7_0),.din(w_dff_A_cp4P7mBH1_0),.clk(gclk));
	jdff dff_A_mygSIe9a7_0(.dout(w_dff_A_o7rzffrE2_0),.din(w_dff_A_mygSIe9a7_0),.clk(gclk));
	jdff dff_A_o7rzffrE2_0(.dout(w_dff_A_nPRB9dci2_0),.din(w_dff_A_o7rzffrE2_0),.clk(gclk));
	jdff dff_A_nPRB9dci2_0(.dout(w_dff_A_kgTTyovo2_0),.din(w_dff_A_nPRB9dci2_0),.clk(gclk));
	jdff dff_A_kgTTyovo2_0(.dout(G372),.din(w_dff_A_kgTTyovo2_0),.clk(gclk));
	jdff dff_A_Ep6aoRix8_2(.dout(w_dff_A_eP3wTA3N7_0),.din(w_dff_A_Ep6aoRix8_2),.clk(gclk));
	jdff dff_A_eP3wTA3N7_0(.dout(w_dff_A_OtAf2P787_0),.din(w_dff_A_eP3wTA3N7_0),.clk(gclk));
	jdff dff_A_OtAf2P787_0(.dout(w_dff_A_WTY8soBG5_0),.din(w_dff_A_OtAf2P787_0),.clk(gclk));
	jdff dff_A_WTY8soBG5_0(.dout(w_dff_A_LdX8lXc20_0),.din(w_dff_A_WTY8soBG5_0),.clk(gclk));
	jdff dff_A_LdX8lXc20_0(.dout(w_dff_A_D608efx06_0),.din(w_dff_A_LdX8lXc20_0),.clk(gclk));
	jdff dff_A_D608efx06_0(.dout(w_dff_A_LIJAooz69_0),.din(w_dff_A_D608efx06_0),.clk(gclk));
	jdff dff_A_LIJAooz69_0(.dout(w_dff_A_VX24oOND5_0),.din(w_dff_A_LIJAooz69_0),.clk(gclk));
	jdff dff_A_VX24oOND5_0(.dout(w_dff_A_SOGSA02F6_0),.din(w_dff_A_VX24oOND5_0),.clk(gclk));
	jdff dff_A_SOGSA02F6_0(.dout(w_dff_A_pfdz49sz5_0),.din(w_dff_A_SOGSA02F6_0),.clk(gclk));
	jdff dff_A_pfdz49sz5_0(.dout(w_dff_A_YnUcfUw68_0),.din(w_dff_A_pfdz49sz5_0),.clk(gclk));
	jdff dff_A_YnUcfUw68_0(.dout(w_dff_A_iA9WOhAQ2_0),.din(w_dff_A_YnUcfUw68_0),.clk(gclk));
	jdff dff_A_iA9WOhAQ2_0(.dout(G369),.din(w_dff_A_iA9WOhAQ2_0),.clk(gclk));
	jdff dff_A_vQ0SPl6k0_2(.dout(w_dff_A_JrM6IIrg5_0),.din(w_dff_A_vQ0SPl6k0_2),.clk(gclk));
	jdff dff_A_JrM6IIrg5_0(.dout(w_dff_A_pklSCn3U3_0),.din(w_dff_A_JrM6IIrg5_0),.clk(gclk));
	jdff dff_A_pklSCn3U3_0(.dout(w_dff_A_TdQOTeQf5_0),.din(w_dff_A_pklSCn3U3_0),.clk(gclk));
	jdff dff_A_TdQOTeQf5_0(.dout(w_dff_A_Pa2E6NBo5_0),.din(w_dff_A_TdQOTeQf5_0),.clk(gclk));
	jdff dff_A_Pa2E6NBo5_0(.dout(w_dff_A_VI4Dtggs0_0),.din(w_dff_A_Pa2E6NBo5_0),.clk(gclk));
	jdff dff_A_VI4Dtggs0_0(.dout(w_dff_A_Opq9hlDY1_0),.din(w_dff_A_VI4Dtggs0_0),.clk(gclk));
	jdff dff_A_Opq9hlDY1_0(.dout(w_dff_A_0lqtm2la8_0),.din(w_dff_A_Opq9hlDY1_0),.clk(gclk));
	jdff dff_A_0lqtm2la8_0(.dout(w_dff_A_i57QZi4A1_0),.din(w_dff_A_0lqtm2la8_0),.clk(gclk));
	jdff dff_A_i57QZi4A1_0(.dout(w_dff_A_R1LmDXZA0_0),.din(w_dff_A_i57QZi4A1_0),.clk(gclk));
	jdff dff_A_R1LmDXZA0_0(.dout(w_dff_A_JI7qBb718_0),.din(w_dff_A_R1LmDXZA0_0),.clk(gclk));
	jdff dff_A_JI7qBb718_0(.dout(G399),.din(w_dff_A_JI7qBb718_0),.clk(gclk));
	jdff dff_A_3k4lhRIx4_2(.dout(w_dff_A_nXDml4y44_0),.din(w_dff_A_3k4lhRIx4_2),.clk(gclk));
	jdff dff_A_nXDml4y44_0(.dout(w_dff_A_Nu36lPLI6_0),.din(w_dff_A_nXDml4y44_0),.clk(gclk));
	jdff dff_A_Nu36lPLI6_0(.dout(w_dff_A_GFS75Zp92_0),.din(w_dff_A_Nu36lPLI6_0),.clk(gclk));
	jdff dff_A_GFS75Zp92_0(.dout(w_dff_A_xzkZ9uSh1_0),.din(w_dff_A_GFS75Zp92_0),.clk(gclk));
	jdff dff_A_xzkZ9uSh1_0(.dout(w_dff_A_TDvoZI8F5_0),.din(w_dff_A_xzkZ9uSh1_0),.clk(gclk));
	jdff dff_A_TDvoZI8F5_0(.dout(w_dff_A_pEEQiuzB3_0),.din(w_dff_A_TDvoZI8F5_0),.clk(gclk));
	jdff dff_A_pEEQiuzB3_0(.dout(w_dff_A_TYhu1Dlb1_0),.din(w_dff_A_pEEQiuzB3_0),.clk(gclk));
	jdff dff_A_TYhu1Dlb1_0(.dout(w_dff_A_aD5WL3mf0_0),.din(w_dff_A_TYhu1Dlb1_0),.clk(gclk));
	jdff dff_A_aD5WL3mf0_0(.dout(w_dff_A_C4xbmaE17_0),.din(w_dff_A_aD5WL3mf0_0),.clk(gclk));
	jdff dff_A_C4xbmaE17_0(.dout(w_dff_A_TdpNpc2m6_0),.din(w_dff_A_C4xbmaE17_0),.clk(gclk));
	jdff dff_A_TdpNpc2m6_0(.dout(G364),.din(w_dff_A_TdpNpc2m6_0),.clk(gclk));
	jdff dff_A_OFRPwL4t5_2(.dout(w_dff_A_a9A7N3kO2_0),.din(w_dff_A_OFRPwL4t5_2),.clk(gclk));
	jdff dff_A_a9A7N3kO2_0(.dout(w_dff_A_yAxqF3cL1_0),.din(w_dff_A_a9A7N3kO2_0),.clk(gclk));
	jdff dff_A_yAxqF3cL1_0(.dout(w_dff_A_QgCylUag0_0),.din(w_dff_A_yAxqF3cL1_0),.clk(gclk));
	jdff dff_A_QgCylUag0_0(.dout(w_dff_A_Xhk2UlNL3_0),.din(w_dff_A_QgCylUag0_0),.clk(gclk));
	jdff dff_A_Xhk2UlNL3_0(.dout(w_dff_A_WcPydgds6_0),.din(w_dff_A_Xhk2UlNL3_0),.clk(gclk));
	jdff dff_A_WcPydgds6_0(.dout(w_dff_A_emA5oVt34_0),.din(w_dff_A_WcPydgds6_0),.clk(gclk));
	jdff dff_A_emA5oVt34_0(.dout(w_dff_A_euiRlEsq7_0),.din(w_dff_A_emA5oVt34_0),.clk(gclk));
	jdff dff_A_euiRlEsq7_0(.dout(w_dff_A_yydSEIER9_0),.din(w_dff_A_euiRlEsq7_0),.clk(gclk));
	jdff dff_A_yydSEIER9_0(.dout(w_dff_A_dEJtFI0h0_0),.din(w_dff_A_yydSEIER9_0),.clk(gclk));
	jdff dff_A_dEJtFI0h0_0(.dout(w_dff_A_LumBvitA5_0),.din(w_dff_A_dEJtFI0h0_0),.clk(gclk));
	jdff dff_A_LumBvitA5_0(.dout(G396),.din(w_dff_A_LumBvitA5_0),.clk(gclk));
	jdff dff_A_ErMg6Nz96_1(.dout(w_dff_A_qUxcG1CY5_0),.din(w_dff_A_ErMg6Nz96_1),.clk(gclk));
	jdff dff_A_qUxcG1CY5_0(.dout(w_dff_A_je4DMXyj0_0),.din(w_dff_A_qUxcG1CY5_0),.clk(gclk));
	jdff dff_A_je4DMXyj0_0(.dout(w_dff_A_qMh23JUk2_0),.din(w_dff_A_je4DMXyj0_0),.clk(gclk));
	jdff dff_A_qMh23JUk2_0(.dout(w_dff_A_36H58dk06_0),.din(w_dff_A_qMh23JUk2_0),.clk(gclk));
	jdff dff_A_36H58dk06_0(.dout(w_dff_A_geHM8Gn20_0),.din(w_dff_A_36H58dk06_0),.clk(gclk));
	jdff dff_A_geHM8Gn20_0(.dout(w_dff_A_2EzwbEhp6_0),.din(w_dff_A_geHM8Gn20_0),.clk(gclk));
	jdff dff_A_2EzwbEhp6_0(.dout(w_dff_A_TWQT8v469_0),.din(w_dff_A_2EzwbEhp6_0),.clk(gclk));
	jdff dff_A_TWQT8v469_0(.dout(G384),.din(w_dff_A_TWQT8v469_0),.clk(gclk));
	jdff dff_A_FbrOxECu5_2(.dout(w_dff_A_sRBNHj852_0),.din(w_dff_A_FbrOxECu5_2),.clk(gclk));
	jdff dff_A_sRBNHj852_0(.dout(w_dff_A_n7NXOdYh2_0),.din(w_dff_A_sRBNHj852_0),.clk(gclk));
	jdff dff_A_n7NXOdYh2_0(.dout(w_dff_A_8lrdO1GS6_0),.din(w_dff_A_n7NXOdYh2_0),.clk(gclk));
	jdff dff_A_8lrdO1GS6_0(.dout(w_dff_A_lCop0IM32_0),.din(w_dff_A_8lrdO1GS6_0),.clk(gclk));
	jdff dff_A_lCop0IM32_0(.dout(G367),.din(w_dff_A_lCop0IM32_0),.clk(gclk));
	jdff dff_A_0lqkBuEO4_2(.dout(w_dff_A_sd6gKFIT9_0),.din(w_dff_A_0lqkBuEO4_2),.clk(gclk));
	jdff dff_A_sd6gKFIT9_0(.dout(w_dff_A_fvywW1pb5_0),.din(w_dff_A_sd6gKFIT9_0),.clk(gclk));
	jdff dff_A_fvywW1pb5_0(.dout(w_dff_A_uM599SED7_0),.din(w_dff_A_fvywW1pb5_0),.clk(gclk));
	jdff dff_A_uM599SED7_0(.dout(w_dff_A_FzYIJVPg9_0),.din(w_dff_A_uM599SED7_0),.clk(gclk));
	jdff dff_A_FzYIJVPg9_0(.dout(G387),.din(w_dff_A_FzYIJVPg9_0),.clk(gclk));
	jdff dff_A_VD26nmsp6_1(.dout(w_dff_A_6bseNoBV9_0),.din(w_dff_A_VD26nmsp6_1),.clk(gclk));
	jdff dff_A_6bseNoBV9_0(.dout(w_dff_A_V3JHIXrH3_0),.din(w_dff_A_6bseNoBV9_0),.clk(gclk));
	jdff dff_A_V3JHIXrH3_0(.dout(w_dff_A_6Q8Zs9tx2_0),.din(w_dff_A_V3JHIXrH3_0),.clk(gclk));
	jdff dff_A_6Q8Zs9tx2_0(.dout(w_dff_A_tLq9uSYe7_0),.din(w_dff_A_6Q8Zs9tx2_0),.clk(gclk));
	jdff dff_A_tLq9uSYe7_0(.dout(w_dff_A_RN59Cewo1_0),.din(w_dff_A_tLq9uSYe7_0),.clk(gclk));
	jdff dff_A_RN59Cewo1_0(.dout(w_dff_A_znlqw13Q4_0),.din(w_dff_A_RN59Cewo1_0),.clk(gclk));
	jdff dff_A_znlqw13Q4_0(.dout(G393),.din(w_dff_A_znlqw13Q4_0),.clk(gclk));
	jdff dff_A_ij4JhiJs2_1(.dout(w_dff_A_6l9hh6411_0),.din(w_dff_A_ij4JhiJs2_1),.clk(gclk));
	jdff dff_A_6l9hh6411_0(.dout(w_dff_A_mUwWp1dw2_0),.din(w_dff_A_6l9hh6411_0),.clk(gclk));
	jdff dff_A_mUwWp1dw2_0(.dout(w_dff_A_Q8xVQi4b3_0),.din(w_dff_A_mUwWp1dw2_0),.clk(gclk));
	jdff dff_A_Q8xVQi4b3_0(.dout(w_dff_A_UIyIURTM6_0),.din(w_dff_A_Q8xVQi4b3_0),.clk(gclk));
	jdff dff_A_UIyIURTM6_0(.dout(w_dff_A_C43idKl58_0),.din(w_dff_A_UIyIURTM6_0),.clk(gclk));
	jdff dff_A_C43idKl58_0(.dout(G390),.din(w_dff_A_C43idKl58_0),.clk(gclk));
	jdff dff_A_9yDN0YMg2_1(.dout(w_dff_A_dVn5qsyl7_0),.din(w_dff_A_9yDN0YMg2_1),.clk(gclk));
	jdff dff_A_dVn5qsyl7_0(.dout(w_dff_A_zscp8Mq69_0),.din(w_dff_A_dVn5qsyl7_0),.clk(gclk));
	jdff dff_A_zscp8Mq69_0(.dout(w_dff_A_kfqeLiiM7_0),.din(w_dff_A_zscp8Mq69_0),.clk(gclk));
	jdff dff_A_kfqeLiiM7_0(.dout(w_dff_A_lmLOe4yt4_0),.din(w_dff_A_kfqeLiiM7_0),.clk(gclk));
	jdff dff_A_lmLOe4yt4_0(.dout(G378),.din(w_dff_A_lmLOe4yt4_0),.clk(gclk));
	jdff dff_A_wSPhLArv2_1(.dout(w_dff_A_3420XUV54_0),.din(w_dff_A_wSPhLArv2_1),.clk(gclk));
	jdff dff_A_3420XUV54_0(.dout(w_dff_A_3MaFdEDz7_0),.din(w_dff_A_3420XUV54_0),.clk(gclk));
	jdff dff_A_3MaFdEDz7_0(.dout(G375),.din(w_dff_A_3MaFdEDz7_0),.clk(gclk));
	jdff dff_A_2VxUnDSH8_1(.dout(w_dff_A_OAhS0AMB1_0),.din(w_dff_A_2VxUnDSH8_1),.clk(gclk));
	jdff dff_A_OAhS0AMB1_0(.dout(w_dff_A_XEXW3dEe3_0),.din(w_dff_A_OAhS0AMB1_0),.clk(gclk));
	jdff dff_A_XEXW3dEe3_0(.dout(w_dff_A_bKJIWztW0_0),.din(w_dff_A_XEXW3dEe3_0),.clk(gclk));
	jdff dff_A_bKJIWztW0_0(.dout(w_dff_A_CC4x2ebW6_0),.din(w_dff_A_bKJIWztW0_0),.clk(gclk));
	jdff dff_A_CC4x2ebW6_0(.dout(G381),.din(w_dff_A_CC4x2ebW6_0),.clk(gclk));
	jdff dff_A_9QSoc5cq7_1(.dout(G407),.din(w_dff_A_9QSoc5cq7_1),.clk(gclk));
	jdff dff_A_5Bcl7rAn0_2(.dout(G402),.din(w_dff_A_5Bcl7rAn0_2),.clk(gclk));
endmodule

