// Benchmark "top" written by ABC on Wed May 27 23:35:00 2020

module top ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , a16 ,
    a17 , a18 , a19 , a20 , a21 , a22 , a23 , a24 ,
    a25 , a26 , a27 , a28 , a29 , a30 , a31 , a32 ,
    a33 , a34 , a35 , a36 , a37 , a38 , a39 , a40 ,
    a41 , a42 , a43 , a44 , a45 , a46 , a47 , a48 ,
    a49 , a50 , a51 , a52 , a53 , a54 , a55 , a56 ,
    a57 , a58 , a59 , a60 , a61 , a62 , a63 , b0 ,
    b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 , b9 ,
    b10 , b11 , b12 , b13 , b14 , b15 , b16 , b17 ,
    b18 , b19 , b20 , b21 , b22 , b23 , b24 , b25 ,
    b26 , b27 , b28 , b29 , b30 , b31 , b32 , b33 ,
    b34 , b35 , b36 , b37 , b38 , b39 , b40 , b41 ,
    b42 , b43 , b44 , b45 , b46 , b47 , b48 , b49 ,
    b50 , b51 , b52 , b53 , b54 , b55 , b56 , b57 ,
    b58 , b59 , b60 , b61 , b62 , b63 ,
    quotient0 , quotient1 , quotient2 , quotient3 ,
    quotient4 , quotient5 , quotient6 , quotient7 ,
    quotient8 , quotient9 , quotient10 , quotient11 ,
    quotient12 , quotient13 , quotient14 , quotient15 ,
    quotient16 , quotient17 , quotient18 , quotient19 ,
    quotient20 , quotient21 , quotient22 , quotient23 ,
    quotient24 , quotient25 , quotient26 , quotient27 ,
    quotient28 , quotient29 , quotient30 , quotient31 ,
    quotient32 , quotient33 , quotient34 , quotient35 ,
    quotient36 , quotient37 , quotient38 , quotient39 ,
    quotient40 , quotient41 , quotient42 , quotient43 ,
    quotient44 , quotient45 , quotient46 , quotient47 ,
    quotient48 , quotient49 , quotient50 , quotient51 ,
    quotient52 , quotient53 , quotient54 , quotient55 ,
    quotient56 , quotient57 , quotient58 , quotient59 ,
    quotient60 , quotient61 , quotient62 , quotient63 ,
    remainder0 , remainder1 , remainder2 , remainder3 ,
    remainder4 , remainder5 , remainder6 , remainder7 ,
    remainder8 , remainder9 , remainder10 , remainder11 ,
    remainder12 , remainder13 , remainder14 , remainder15 ,
    remainder16 , remainder17 , remainder18 , remainder19 ,
    remainder20 , remainder21 , remainder22 , remainder23 ,
    remainder24 , remainder25 , remainder26 , remainder27 ,
    remainder28 , remainder29 , remainder30 , remainder31 ,
    remainder32 , remainder33 , remainder34 , remainder35 ,
    remainder36 , remainder37 , remainder38 , remainder39 ,
    remainder40 , remainder41 , remainder42 , remainder43 ,
    remainder44 , remainder45 , remainder46 , remainder47 ,
    remainder48 , remainder49 , remainder50 , remainder51 ,
    remainder52 , remainder53 , remainder54 , remainder55 ,
    remainder56 , remainder57 , remainder58 , remainder59 ,
    remainder60 , remainder61 , remainder62 , remainder63   );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    a16 , a17 , a18 , a19 , a20 , a21 , a22 , a23 ,
    a24 , a25 , a26 , a27 , a28 , a29 , a30 , a31 ,
    a32 , a33 , a34 , a35 , a36 , a37 , a38 , a39 ,
    a40 , a41 , a42 , a43 , a44 , a45 , a46 , a47 ,
    a48 , a49 , a50 , a51 , a52 , a53 , a54 , a55 ,
    a56 , a57 , a58 , a59 , a60 , a61 , a62 , a63 ,
    b0 , b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 ,
    b9 , b10 , b11 , b12 , b13 , b14 , b15 , b16 ,
    b17 , b18 , b19 , b20 , b21 , b22 , b23 , b24 ,
    b25 , b26 , b27 , b28 , b29 , b30 , b31 , b32 ,
    b33 , b34 , b35 , b36 , b37 , b38 , b39 , b40 ,
    b41 , b42 , b43 , b44 , b45 , b46 , b47 , b48 ,
    b49 , b50 , b51 , b52 , b53 , b54 , b55 , b56 ,
    b57 , b58 , b59 , b60 , b61 , b62 , b63 ;
  output quotient0 , quotient1 , quotient2 , quotient3 ,
    quotient4 , quotient5 , quotient6 , quotient7 ,
    quotient8 , quotient9 , quotient10 , quotient11 ,
    quotient12 , quotient13 , quotient14 , quotient15 ,
    quotient16 , quotient17 , quotient18 , quotient19 ,
    quotient20 , quotient21 , quotient22 , quotient23 ,
    quotient24 , quotient25 , quotient26 , quotient27 ,
    quotient28 , quotient29 , quotient30 , quotient31 ,
    quotient32 , quotient33 , quotient34 , quotient35 ,
    quotient36 , quotient37 , quotient38 , quotient39 ,
    quotient40 , quotient41 , quotient42 , quotient43 ,
    quotient44 , quotient45 , quotient46 , quotient47 ,
    quotient48 , quotient49 , quotient50 , quotient51 ,
    quotient52 , quotient53 , quotient54 , quotient55 ,
    quotient56 , quotient57 , quotient58 , quotient59 ,
    quotient60 , quotient61 , quotient62 , quotient63 ,
    remainder0 , remainder1 , remainder2 , remainder3 ,
    remainder4 , remainder5 , remainder6 , remainder7 ,
    remainder8 , remainder9 , remainder10 , remainder11 ,
    remainder12 , remainder13 , remainder14 , remainder15 ,
    remainder16 , remainder17 , remainder18 , remainder19 ,
    remainder20 , remainder21 , remainder22 , remainder23 ,
    remainder24 , remainder25 , remainder26 , remainder27 ,
    remainder28 , remainder29 , remainder30 , remainder31 ,
    remainder32 , remainder33 , remainder34 , remainder35 ,
    remainder36 , remainder37 , remainder38 , remainder39 ,
    remainder40 , remainder41 , remainder42 , remainder43 ,
    remainder44 , remainder45 , remainder46 , remainder47 ,
    remainder48 , remainder49 , remainder50 , remainder51 ,
    remainder52 , remainder53 , remainder54 , remainder55 ,
    remainder56 , remainder57 , remainder58 , remainder59 ,
    remainder60 , remainder61 , remainder62 , remainder63 ;
  wire n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n458, n459,
    n460, n461, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n546, n547, n548, n551, n554,
    n555, n556, n557, n558, n559, n563, n564, n565, n566, n567, n569, n571,
    n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638, n641, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938, n939, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1161, n1162, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1553, n1554, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1620, n1621, n1623, n1624, n1625, n1626, n1630,
    n1632, n1633, n1638, n1639, n1643, n1644, n1648, n1649, n1653, n1654,
    n1658, n1659, n1663, n1664, n1668, n1669, n1673, n1674, n1678, n1679,
    n1683, n1684, n1688, n1694, n1695, n1696, n1698, n1701, n1702, n1703,
    n1704, n1705, n1706, n1708, n1709, n1711, n1712, n1714, n1715, n1717,
    n1718, n1720, n1721, n1723, n1724, n1726, n1727, n1729, n1730, n1732,
    n1733, n1735, n1736, n1738, n1739, n1741, n1742, n1744, n1745, n1746,
    n1747, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1830, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
    n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
    n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
    n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
    n1973, n1974, n1975, n1976, n1977, n1979, n1980, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2040,
    n2045, n2054, n2060, n2065, n2070, n2075, n2080, n2085, n2090, n2095,
    n2100, n2105, n2110, n2115, n2120, n2125, n2133, n2138, n2139, n2140,
    n2196, n2197, n2280, n2282, n2283, n2284, n2285, n2288, n2289, n2292,
    n2293, n2298, n2299, n2300, n2442, n2445, n2446, n2457, n2458, n2459,
    n2460, n2461, n2468, n2470, n2471, n2472, n2547, n2649, n2650, n2651,
    n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2851, n2852, n2855,
    n2860, n2861, n2953, n3111, n3118, n3119, n3120, n3320, n3321, n3322,
    n3400, n3401, n3402, n3403, n3544, n3545, n3548, n3553, n3554, n3658,
    n3716, n3838, n3839, n3840, n3847, n3848, n3849, n4073, n4074, n4075,
    n4295, n4301, n4302, n4303, n4533, n4534, n4535, n4536, n4539, n4545,
    n4546, n4547, n4642, n4798, n4799, n4800, n5046, n5052, n5053, n5054,
    n5307, n5308, n5311, n5317, n5318, n5319, n5591, n5592, n5593, n5692,
    n5693, n5694, n5701, n5702, n5703, n5704, n5899, n5900, n5903, n5908,
    n5909, n6049, n6286, n6293, n6294, n6295, n6403, n6404, n6599, n6600,
    n6601, n6715, n6716, n6929, n6930, n6933, n6938, n6939, n7091, n7354,
    n7355, n7356, n7363, n7364, n7365, n7722, n7723, n7883, n7960, n8203,
    n8204, n8369, n8458, n8658, n8659, n8660, n8667, n8668, n8669, n9015,
    n9016, n9017, n9354, n9360, n9361, n9362, n9719, n9720, n9721, n9866,
    n9867, n9868, n9869, n10100, n10101, n10102, n10459, n10460, n10463,
    n10469, n10470, n10471, n10607, n10853, n10854, n10855, n11254, n11255,
    n11256, n11637, n11638, n11641, n11647, n11648, n11649, n11794, n12061,
    n12062, n12063, n12211, n12214, n12215, n12216, n12485, n12486, n12487,
    n12894, n12895, n12898, n12904, n12905, n12906, n13060, n13081, n13342,
    n13343, n13344, n13501, n13502, n13503, n13504, n13837, n13838, n14053,
    n14054, n14055, n14061, n14440, n14447, n14448, n14449, n14612, n14903,
    n14904, n14905, n15090, n15381, n15382, n15383, n15840, n15845, n15846,
    n15847, n16024, n16325, n16326, n16327, n16812, n16813, n16814, n17307,
    n17308, n17309, n17810, n17811, n17812, n18009, n18364, n18365, n18490,
    n18497, n18498, n18499, n18501, n18502, n18511, n18568, n18575, n18577,
    n18578, n18579, n18592, n18593, n18596, n18651, n18652, n18653, n18720,
    n18735, n18737, n18738, n18739, n18768, n18798, n18801, n18802, n18803,
    n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
    n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
    n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
    n18938, n18939, n18943, n19007, n19037, n19039, n19040, n19041, n19139,
    n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
    n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
    n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
    n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19219, n19220,
    n19221, n19223, n19255, n19307, n19310, n19311, n19313, n19314, n19315,
    n19316, n19317, n19327, n19400, n19445, n19447, n19448, n19449, n19574,
    n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
    n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
    n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
    n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
    n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
    n19620, n19678, n19679, n19680, n19682, n19713, n19718, n19723, n19729,
    n19735, n19741, n19747, n19753, n19759, n19765, n19771, n19779, n19787,
    n19788, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
    n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19813, n19814,
    n19815, n19817, n19818, n19819, n19821, n19822, n19823, n19825, n19826,
    n19827, n19829, n19830, n19831, n19833, n19834, n19835, n19837, n19838,
    n19839, n19841, n19842, n19843, n19845, n19846, n19847, n19849, n19850,
    n19851, n19853, n19854, n19855, n19856, n19858, n19859, n19860, n19891,
    n19892, n19893, n19894, n19896, n19897, n19899, n19900, n19901, n19904,
    n19905, n19906, n19909, n19910, n19911, n19914, n19915, n19916, n19919,
    n19920, n19921, n19924, n19925, n19926, n19929, n19930, n19931, n19934,
    n19935, n19936, n19939, n19940, n19941, n19944, n19945, n19946, n19949,
    n19950, n19951, n19954, n19955, n19956, n19959, n19960, n19961, n19963,
    n19964, n19965, n19966, n19967, n19968, n19970, n19971, n19978, n19981,
    n19984, n19987, n19990, n19993, n19996, n19999, n20002, n20005, n20008,
    n20011, n20014, n20019, n20094, n20097, n20098, n20099, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
    n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
    n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
    n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
    n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20166,
    n20167, n20227, n20233, n20239, n20245, n20251, n20257, n20263, n20269,
    n20275, n20281, n20287, n20293, n20299, n20305, n20313, n20321, n20322,
    n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
    n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
    n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
    n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
    n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
    n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
    n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
    n20386, n20387, n20388, n20390, n20391, n20396, n20397, n20398, n20400,
    n20401, n20402, n20404, n20405, n20406, n20408, n20409, n20410, n20412,
    n20413, n20414, n20416, n20417, n20418, n20420, n20421, n20422, n20424,
    n20425, n20426, n20428, n20429, n20430, n20432, n20433, n20434, n20436,
    n20437, n20438, n20440, n20441, n20442, n20444, n20445, n20446, n20448,
    n20449, n20450, n20452, n20453, n20454, n20456, n20457, n20458, n20460,
    n20461, n20462, n20496, n20497, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20508, n20509, n20511, n20512, n20513, n20514,
    n20516, n20517, n20518, n20519, n20521, n20522, n20523, n20524, n20526,
    n20527, n20528, n20529, n20531, n20532, n20533, n20534, n20536, n20537,
    n20538, n20539, n20541, n20542, n20543, n20544, n20546, n20547, n20548,
    n20549, n20551, n20552, n20553, n20554, n20556, n20557, n20558, n20559,
    n20561, n20562, n20563, n20564, n20566, n20567, n20568, n20569, n20571,
    n20572, n20573, n20574, n20576, n20577, n20578, n20579, n20581, n20582,
    n20583, n20584, n20586, n20587, n20588, n20589, n20590, n20591, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
    n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
    n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
    n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
    n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
    n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
    n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
    n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
    n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
    n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
    n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
    n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
    n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
    n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
    n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
    n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
    n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
    n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
    n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
    n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
    n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
    n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
    n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
    n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
    n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
    n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
    n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
    n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
    n20909, n20910, n20911, n20912, n20913, n20914, n20917, n20918, n20919,
    n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
    n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
    n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
    n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
    n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
    n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
    n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
    n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
    n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
    n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
    n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
    n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
    n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21066,
    n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
    n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
    n21085, n21086, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
    n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
    n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
    n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
    n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
    n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
    n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
    n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
    n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
    n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
    n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
    n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
    n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
    n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
    n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
    n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
    n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
    n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
    n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
    n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
    n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
    n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
    n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
    n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
    n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
    n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
    n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
    n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
    n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
    n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
    n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
    n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
    n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
    n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
    n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
    n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
    n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
    n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
    n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
    n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
    n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
    n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
    n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
    n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
    n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
    n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
    n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
    n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
    n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
    n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
    n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
    n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
    n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
    n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
    n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
    n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
    n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598,
    n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
    n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
    n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
    n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
    n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
    n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
    n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
    n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670,
    n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
    n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,
    n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
    n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
    n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
    n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
    n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
    n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
    n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
    n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
    n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
    n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
    n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
    n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
    n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805,
    n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814,
    n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
    n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
    n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
    n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
    n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
    n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
    n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877,
    n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
    n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
    n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
    n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
    n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
    n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
    n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
    n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949,
    n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958,
    n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
    n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
    n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
    n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
    n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
    n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
    n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021,
    n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030,
    n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
    n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,
    n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
    n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
    n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
    n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
    n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093,
    n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102,
    n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
    n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
    n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
    n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
    n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
    n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
    n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165,
    n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174,
    n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
    n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
    n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
    n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
    n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
    n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
    n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237,
    n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
    n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
    n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
    n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
    n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
    n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
    n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
    n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309,
    n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318,
    n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
    n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
    n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
    n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
    n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
    n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372,
    n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381,
    n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390,
    n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
    n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
    n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
    n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
    n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
    n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
    n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453,
    n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462,
    n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
    n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
    n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
    n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
    n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
    n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
    n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525,
    n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534,
    n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
    n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
    n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
    n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
    n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
    n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588,
    n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597,
    n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606,
    n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
    n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,
    n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
    n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
    n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
    n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669,
    n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678,
    n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
    n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
    n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
    n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
    n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
    n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
    n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741,
    n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750,
    n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
    n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
    n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
    n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
    n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
    n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804,
    n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813,
    n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822,
    n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
    n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
    n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
    n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
    n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
    n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876,
    n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885,
    n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894,
    n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
    n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
    n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
    n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930,
    n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
    n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948,
    n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957,
    n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966,
    n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
    n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,
    n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
    n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002,
    n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
    n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020,
    n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029,
    n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038,
    n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
    n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
    n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
    n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074,
    n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
    n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092,
    n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101,
    n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110,
    n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119,
    n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128,
    n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
    n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146,
    n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
    n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164,
    n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173,
    n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182,
    n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191,
    n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200,
    n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
    n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218,
    n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
    n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236,
    n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245,
    n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254,
    n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
    n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272,
    n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
    n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290,
    n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
    n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308,
    n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317,
    n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326,
    n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
    n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,
    n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
    n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362,
    n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
    n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380,
    n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389,
    n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398,
    n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
    n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416,
    n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
    n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434,
    n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
    n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452,
    n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461,
    n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470,
    n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479,
    n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488,
    n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
    n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506,
    n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
    n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524,
    n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533,
    n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542,
    n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551,
    n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560,
    n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
    n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578,
    n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
    n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596,
    n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605,
    n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614,
    n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
    n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632,
    n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
    n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650,
    n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
    n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668,
    n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677,
    n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686,
    n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
    n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704,
    n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
    n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
    n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
    n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740,
    n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
    n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758,
    n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
    n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776,
    n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
    n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
    n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
    n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812,
    n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821,
    n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830,
    n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
    n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,
    n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
    n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
    n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
    n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884,
    n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
    n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
    n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
    n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
    n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
    n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
    n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956,
    n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
    n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974,
    n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
    n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,
    n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
    n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010,
    n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
    n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028,
    n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
    n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046,
    n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
    n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
    n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
    n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082,
    n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
    n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100,
    n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
    n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118,
    n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
    n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
    n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
    n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
    n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
    n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172,
    n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181,
    n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190,
    n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
    n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
    n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
    n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226,
    n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
    n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244,
    n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253,
    n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262,
    n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271,
    n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280,
    n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
    n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298,
    n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
    n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316,
    n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325,
    n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334,
    n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343,
    n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352,
    n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
    n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370,
    n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
    n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388,
    n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397,
    n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406,
    n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
    n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
    n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
    n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
    n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
    n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460,
    n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469,
    n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478,
    n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
    n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,
    n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
    n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
    n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
    n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532,
    n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541,
    n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550,
    n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559,
    n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568,
    n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
    n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586,
    n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
    n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604,
    n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613,
    n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622,
    n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631,
    n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640,
    n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
    n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
    n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
    n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676,
    n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685,
    n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694,
    n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
    n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712,
    n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
    n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
    n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
    n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748,
    n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757,
    n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766,
    n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775,
    n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784,
    n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
    n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
    n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
    n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820,
    n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829,
    n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838,
    n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847,
    n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856,
    n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
    n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
    n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
    n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892,
    n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901,
    n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910,
    n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
    n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,
    n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
    n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
    n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
    n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
    n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973,
    n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982,
    n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991,
    n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,
    n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
    n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
    n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
    n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036,
    n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045,
    n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054,
    n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063,
    n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
    n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
    n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
    n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
    n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108,
    n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117,
    n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126,
    n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135,
    n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
    n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
    n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
    n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
    n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180,
    n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189,
    n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198,
    n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207,
    n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
    n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
    n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
    n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
    n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252,
    n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261,
    n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270,
    n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279,
    n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
    n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
    n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
    n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
    n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324,
    n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333,
    n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342,
    n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351,
    n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,
    n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
    n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
    n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
    n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396,
    n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405,
    n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414,
    n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423,
    n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
    n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
    n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
    n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
    n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468,
    n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477,
    n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486,
    n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495,
    n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,
    n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
    n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
    n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
    n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540,
    n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549,
    n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558,
    n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567,
    n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576,
    n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
    n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
    n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
    n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612,
    n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621,
    n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630,
    n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639,
    n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648,
    n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
    n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
    n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
    n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684,
    n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693,
    n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702,
    n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711,
    n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720,
    n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
    n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
    n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
    n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756,
    n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765,
    n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774,
    n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783,
    n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,
    n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
    n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810,
    n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
    n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828,
    n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837,
    n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846,
    n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855,
    n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864,
    n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
    n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882,
    n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
    n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900,
    n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909,
    n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918,
    n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927,
    n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936,
    n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
    n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954,
    n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
    n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972,
    n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981,
    n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990,
    n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999,
    n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008,
    n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
    n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
    n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044,
    n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062,
    n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
    n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
    n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
    n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116,
    n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125,
    n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134,
    n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143,
    n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
    n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
    n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
    n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
    n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188,
    n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197,
    n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206,
    n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215,
    n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
    n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
    n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
    n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
    n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260,
    n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269,
    n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278,
    n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287,
    n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296,
    n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
    n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314,
    n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
    n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332,
    n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341,
    n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350,
    n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359,
    n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,
    n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
    n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
    n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
    n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404,
    n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413,
    n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422,
    n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431,
    n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,
    n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
    n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
    n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
    n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476,
    n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485,
    n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494,
    n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503,
    n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512,
    n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
    n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
    n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
    n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548,
    n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557,
    n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566,
    n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575,
    n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584,
    n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
    n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
    n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
    n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620,
    n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629,
    n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638,
    n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647,
    n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656,
    n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
    n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
    n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
    n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692,
    n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
    n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710,
    n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719,
    n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728,
    n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
    n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
    n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
    n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
    n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773,
    n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782,
    n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791,
    n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800,
    n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
    n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
    n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
    n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836,
    n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845,
    n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854,
    n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863,
    n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872,
    n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
    n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
    n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899,
    n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908,
    n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917,
    n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926,
    n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935,
    n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944,
    n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
    n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
    n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971,
    n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980,
    n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989,
    n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998,
    n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007,
    n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016,
    n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
    n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
    n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043,
    n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052,
    n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061,
    n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070,
    n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079,
    n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088,
    n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
    n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
    n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
    n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124,
    n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133,
    n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142,
    n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151,
    n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,
    n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
    n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
    n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
    n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196,
    n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205,
    n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214,
    n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223,
    n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232,
    n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
    n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
    n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259,
    n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268,
    n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277,
    n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286,
    n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295,
    n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304,
    n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
    n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322,
    n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
    n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340,
    n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349,
    n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358,
    n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367,
    n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376,
    n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
    n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394,
    n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
    n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412,
    n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421,
    n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430,
    n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439,
    n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448,
    n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
    n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466,
    n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475,
    n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484,
    n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493,
    n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502,
    n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511,
    n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520,
    n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
    n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
    n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
    n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556,
    n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565,
    n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574,
    n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583,
    n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592,
    n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
    n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
    n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
    n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628,
    n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637,
    n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646,
    n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655,
    n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664,
    n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
    n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
    n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
    n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700,
    n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709,
    n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718,
    n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727,
    n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736,
    n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
    n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754,
    n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
    n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772,
    n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781,
    n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790,
    n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799,
    n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808,
    n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
    n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
    n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
    n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844,
    n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853,
    n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862,
    n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871,
    n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880,
    n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
    n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898,
    n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
    n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916,
    n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925,
    n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934,
    n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943,
    n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952,
    n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
    n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
    n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
    n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988,
    n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997,
    n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006,
    n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015,
    n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024,
    n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
    n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
    n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
    n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060,
    n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069,
    n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078,
    n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087,
    n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096,
    n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
    n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
    n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
    n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132,
    n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141,
    n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150,
    n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159,
    n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168,
    n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
    n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
    n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
    n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204,
    n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213,
    n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222,
    n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231,
    n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240,
    n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
    n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258,
    n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
    n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276,
    n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285,
    n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294,
    n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303,
    n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312,
    n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
    n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
    n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
    n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348,
    n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
    n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366,
    n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375,
    n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384,
    n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
    n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
    n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
    n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
    n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
    n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447,
    n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
    n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
    n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
    n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
    n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492,
    n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501,
    n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510,
    n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
    n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528,
    n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
    n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546,
    n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
    n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564,
    n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573,
    n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582,
    n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591,
    n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600,
    n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
    n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
    n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
    n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636,
    n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645,
    n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654,
    n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663,
    n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672,
    n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
    n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690,
    n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
    n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708,
    n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717,
    n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726,
    n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735,
    n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744,
    n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
    n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762,
    n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
    n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780,
    n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789,
    n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798,
    n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807,
    n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816,
    n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
    n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834,
    n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
    n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852,
    n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861,
    n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870,
    n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879,
    n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888,
    n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
    n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906,
    n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
    n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924,
    n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933,
    n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942,
    n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951,
    n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960,
    n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
    n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978,
    n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987,
    n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996,
    n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005,
    n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014,
    n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023,
    n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032,
    n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
    n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050,
    n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059,
    n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068,
    n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077,
    n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086,
    n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095,
    n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104,
    n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
    n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122,
    n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131,
    n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140,
    n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149,
    n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158,
    n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167,
    n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176,
    n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
    n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194,
    n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
    n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212,
    n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221,
    n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230,
    n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239,
    n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248,
    n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
    n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266,
    n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
    n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284,
    n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293,
    n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302,
    n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311,
    n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320,
    n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
    n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338,
    n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347,
    n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356,
    n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365,
    n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374,
    n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383,
    n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392,
    n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
    n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410,
    n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419,
    n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428,
    n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437,
    n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446,
    n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455,
    n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464,
    n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
    n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482,
    n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491,
    n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500,
    n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509,
    n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518,
    n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527,
    n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536,
    n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
    n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554,
    n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563,
    n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572,
    n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581,
    n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590,
    n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599,
    n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608,
    n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
    n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
    n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635,
    n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644,
    n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653,
    n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662,
    n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671,
    n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680,
    n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
    n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698,
    n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
    n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716,
    n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725,
    n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
    n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743,
    n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752,
    n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
    n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770,
    n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779,
    n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788,
    n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797,
    n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806,
    n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815,
    n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824,
    n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
    n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842,
    n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851,
    n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860,
    n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869,
    n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878,
    n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887,
    n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896,
    n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
    n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914,
    n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
    n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932,
    n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941,
    n29942, n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950,
    n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959,
    n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968,
    n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
    n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986,
    n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995,
    n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004,
    n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013,
    n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022,
    n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031,
    n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040,
    n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
    n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058,
    n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067,
    n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076,
    n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085,
    n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094,
    n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103,
    n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112,
    n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
    n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130,
    n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139,
    n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148,
    n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157,
    n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166,
    n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175,
    n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184,
    n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
    n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202,
    n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211,
    n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220,
    n30221, n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229,
    n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238,
    n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247,
    n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256,
    n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
    n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274,
    n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283,
    n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292,
    n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301,
    n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310,
    n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319,
    n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328,
    n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
    n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346,
    n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355,
    n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364,
    n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373,
    n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382,
    n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391,
    n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400,
    n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
    n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418,
    n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427,
    n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436,
    n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445,
    n30446, n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454,
    n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463,
    n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472,
    n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
    n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490,
    n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499,
    n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508,
    n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517,
    n30518, n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526,
    n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535,
    n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544,
    n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
    n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562,
    n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571,
    n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580,
    n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589,
    n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598,
    n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607,
    n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616,
    n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
    n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634,
    n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643,
    n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652,
    n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661,
    n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670,
    n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679,
    n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688,
    n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
    n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706,
    n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715,
    n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724,
    n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733,
    n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742,
    n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751,
    n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760,
    n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
    n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778,
    n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787,
    n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796,
    n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805,
    n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814,
    n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823,
    n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832,
    n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
    n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850,
    n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859,
    n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868,
    n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877,
    n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886,
    n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895,
    n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904,
    n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
    n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922,
    n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931,
    n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940,
    n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949,
    n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958,
    n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967,
    n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976,
    n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
    n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994,
    n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003,
    n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012,
    n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021,
    n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030,
    n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039,
    n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048,
    n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
    n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066,
    n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075,
    n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084,
    n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093,
    n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
    n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111,
    n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120,
    n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
    n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138,
    n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147,
    n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156,
    n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165,
    n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174,
    n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183,
    n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192,
    n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
    n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210,
    n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219,
    n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228,
    n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237,
    n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246,
    n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255,
    n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264,
    n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
    n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282,
    n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291,
    n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300,
    n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309,
    n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318,
    n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327,
    n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336,
    n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
    n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354,
    n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363,
    n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372,
    n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381,
    n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390,
    n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399,
    n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408,
    n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
    n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426,
    n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435,
    n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444,
    n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453,
    n31454, n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462,
    n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471,
    n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480,
    n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
    n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498,
    n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507,
    n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516,
    n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525,
    n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534,
    n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543,
    n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552,
    n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
    n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570,
    n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579,
    n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588,
    n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597,
    n31598, n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606,
    n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615,
    n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624,
    n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
    n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642,
    n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651,
    n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660,
    n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669,
    n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678,
    n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687,
    n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696,
    n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
    n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714,
    n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723,
    n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732,
    n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741,
    n31742, n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750,
    n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759,
    n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768,
    n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
    n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786,
    n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795,
    n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804,
    n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813,
    n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822,
    n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831,
    n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840,
    n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
    n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858,
    n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867,
    n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876,
    n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885,
    n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894,
    n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903,
    n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912,
    n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
    n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930,
    n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939,
    n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948,
    n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957,
    n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966,
    n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975,
    n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984,
    n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
    n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002,
    n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011,
    n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020,
    n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029,
    n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038,
    n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047,
    n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056,
    n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
    n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074,
    n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083,
    n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092,
    n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101,
    n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110,
    n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119,
    n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128,
    n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
    n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146,
    n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155,
    n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164,
    n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173,
    n32174, n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182,
    n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191,
    n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200,
    n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
    n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218,
    n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227,
    n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236,
    n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245,
    n32246, n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254,
    n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263,
    n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272,
    n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
    n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290,
    n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299,
    n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308,
    n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317,
    n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326,
    n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335,
    n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344,
    n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
    n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362,
    n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371,
    n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380,
    n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389,
    n32390, n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398,
    n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407,
    n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416,
    n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
    n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434,
    n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443,
    n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452,
    n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461,
    n32462, n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470,
    n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479,
    n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488,
    n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
    n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506,
    n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515,
    n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524,
    n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533,
    n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542,
    n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551,
    n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560,
    n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
    n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578,
    n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587,
    n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596,
    n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605,
    n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614,
    n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623,
    n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632,
    n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
    n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650,
    n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659,
    n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668,
    n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677,
    n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
    n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695,
    n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704,
    n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
    n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722,
    n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731,
    n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740,
    n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749,
    n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758,
    n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767,
    n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776,
    n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
    n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794,
    n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803,
    n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812,
    n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821,
    n32822, n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830,
    n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839,
    n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848,
    n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
    n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866,
    n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875,
    n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884,
    n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893,
    n32894, n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
    n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911,
    n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920,
    n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
    n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938,
    n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947,
    n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956,
    n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965,
    n32966, n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974,
    n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983,
    n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992,
    n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
    n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010,
    n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019,
    n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028,
    n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037,
    n33038, n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046,
    n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055,
    n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064,
    n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
    n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082,
    n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091,
    n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100,
    n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109,
    n33110, n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118,
    n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127,
    n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136,
    n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
    n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154,
    n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163,
    n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172,
    n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181,
    n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190,
    n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199,
    n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208,
    n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
    n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226,
    n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235,
    n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244,
    n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253,
    n33254, n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262,
    n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271,
    n33272, n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280,
    n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
    n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298,
    n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307,
    n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316,
    n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325,
    n33326, n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334,
    n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343,
    n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352,
    n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
    n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370,
    n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379,
    n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388,
    n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397,
    n33398, n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406,
    n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415,
    n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424,
    n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
    n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442,
    n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451,
    n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460,
    n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469,
    n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478,
    n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487,
    n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496,
    n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
    n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514,
    n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523,
    n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532,
    n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541,
    n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550,
    n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559,
    n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568,
    n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
    n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586,
    n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595,
    n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604,
    n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613,
    n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622,
    n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631,
    n33632, n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640,
    n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
    n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658,
    n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667,
    n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676,
    n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685,
    n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
    n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703,
    n33704, n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712,
    n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
    n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730,
    n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739,
    n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748,
    n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757,
    n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
    n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775,
    n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784,
    n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
    n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802,
    n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811,
    n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820,
    n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829,
    n33830, n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
    n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847,
    n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856,
    n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
    n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874,
    n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883,
    n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892,
    n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901,
    n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
    n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919,
    n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928,
    n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
    n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946,
    n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955,
    n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964,
    n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972, n33973,
    n33974, n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982,
    n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991,
    n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000,
    n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
    n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018,
    n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027,
    n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036,
    n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044, n34045,
    n34046, n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054,
    n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063,
    n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072,
    n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
    n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090,
    n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099,
    n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108,
    n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116, n34117,
    n34118, n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
    n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135,
    n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144,
    n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
    n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162,
    n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171,
    n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180,
    n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189,
    n34190, n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198,
    n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207,
    n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216,
    n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
    n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234,
    n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243,
    n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252,
    n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261,
    n34262, n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270,
    n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279,
    n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288,
    n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
    n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306,
    n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315,
    n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324,
    n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333,
    n34334, n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342,
    n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351,
    n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360,
    n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
    n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378,
    n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387,
    n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396,
    n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405,
    n34406, n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414,
    n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423,
    n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432,
    n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
    n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450,
    n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459,
    n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468,
    n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477,
    n34478, n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486,
    n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495,
    n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504,
    n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
    n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522,
    n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531,
    n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540,
    n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549,
    n34550, n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558,
    n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567,
    n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576,
    n34577, n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
    n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594,
    n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603,
    n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612,
    n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620, n34621,
    n34622, n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630,
    n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639,
    n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648,
    n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
    n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666,
    n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675,
    n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684,
    n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693,
    n34694, n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702,
    n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711,
    n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720,
    n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
    n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738,
    n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747,
    n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756,
    n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765,
    n34766, n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774,
    n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783,
    n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792,
    n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
    n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810,
    n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819,
    n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828,
    n34829, n34830, n34831, n34832, n34833, n34834, n34835, n34836, n34837,
    n34838, n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846,
    n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855,
    n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864,
    n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
    n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882,
    n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891,
    n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900,
    n34901, n34902, n34903, n34904, n34905, n34906, n34907, n34908, n34909,
    n34910, n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918,
    n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927,
    n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936,
    n34937, n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
    n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954,
    n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963,
    n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972,
    n34973, n34974, n34975, n34976, n34977, n34978, n34979, n34980, n34981,
    n34982, n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990,
    n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999,
    n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008,
    n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
    n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026,
    n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035,
    n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044,
    n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053,
    n35054, n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062,
    n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071,
    n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080,
    n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
    n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098,
    n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107,
    n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116,
    n35117, n35118, n35119, n35120, n35121, n35122, n35123, n35124, n35125,
    n35126, n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134,
    n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143,
    n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152,
    n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
    n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170,
    n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179,
    n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188,
    n35189, n35190, n35191, n35192, n35193, n35194, n35195, n35196, n35197,
    n35198, n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206,
    n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215,
    n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224,
    n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
    n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242,
    n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251,
    n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260,
    n35261, n35262, n35263, n35264, n35265, n35266, n35267, n35268, n35269,
    n35270, n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278,
    n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287,
    n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296,
    n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
    n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314,
    n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323,
    n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332,
    n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340, n35341,
    n35342, n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350,
    n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359,
    n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368,
    n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
    n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386,
    n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395,
    n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404,
    n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412, n35413,
    n35414, n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422,
    n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431,
    n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440,
    n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
    n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458,
    n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467,
    n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476,
    n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484, n35485,
    n35486, n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494,
    n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503,
    n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512,
    n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
    n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530,
    n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539,
    n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548,
    n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556, n35557,
    n35558, n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566,
    n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575,
    n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584,
    n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
    n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602,
    n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611,
    n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620,
    n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629,
    n35630, n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638,
    n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647,
    n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656,
    n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
    n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674,
    n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683,
    n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692,
    n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701,
    n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710,
    n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719,
    n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728,
    n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
    n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746,
    n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755,
    n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764,
    n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772, n35773,
    n35774, n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782,
    n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791,
    n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800,
    n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
    n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818,
    n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827,
    n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836,
    n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844, n35845,
    n35846, n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854,
    n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863,
    n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872,
    n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
    n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890,
    n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899,
    n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908,
    n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916, n35917,
    n35918, n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926,
    n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935,
    n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944,
    n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
    n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962,
    n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971,
    n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980,
    n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988, n35989,
    n35990, n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998,
    n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007,
    n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016,
    n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
    n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034,
    n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043,
    n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052,
    n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060, n36061,
    n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070,
    n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079,
    n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088,
    n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
    n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106,
    n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115,
    n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124,
    n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133,
    n36134, n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142,
    n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151,
    n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160,
    n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
    n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178,
    n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187,
    n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196,
    n36197, n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205,
    n36206, n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214,
    n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223,
    n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232,
    n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
    n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250,
    n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259,
    n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268,
    n36269, n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277,
    n36278, n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286,
    n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295,
    n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304,
    n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
    n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322,
    n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331,
    n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340,
    n36341, n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349,
    n36350, n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358,
    n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367,
    n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376,
    n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
    n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394,
    n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403,
    n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412,
    n36413, n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421,
    n36422, n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430,
    n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439,
    n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448,
    n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
    n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466,
    n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475,
    n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484,
    n36485, n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493,
    n36494, n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502,
    n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511,
    n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520,
    n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
    n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538,
    n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547,
    n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556,
    n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565,
    n36566, n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574,
    n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583,
    n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592,
    n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
    n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610,
    n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619,
    n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628,
    n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637,
    n36638, n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646,
    n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655,
    n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664,
    n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
    n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682,
    n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691,
    n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700,
    n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708, n36709,
    n36710, n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718,
    n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727,
    n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736,
    n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
    n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754,
    n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763,
    n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772,
    n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781,
    n36782, n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790,
    n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799,
    n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808,
    n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
    n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826,
    n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835,
    n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844,
    n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852, n36853,
    n36854, n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862,
    n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871,
    n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880,
    n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
    n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898,
    n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907,
    n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916,
    n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925,
    n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934,
    n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943,
    n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952,
    n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
    n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970,
    n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979,
    n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988,
    n36989, n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997,
    n36998, n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006,
    n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015,
    n37016, n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024,
    n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
    n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042,
    n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051,
    n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060,
    n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069,
    n37070, n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078,
    n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087,
    n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096,
    n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
    n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114,
    n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123,
    n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132,
    n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141,
    n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150,
    n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159,
    n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168,
    n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
    n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186,
    n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195,
    n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204,
    n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213,
    n37214, n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222,
    n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231,
    n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240,
    n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
    n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258,
    n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267,
    n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276,
    n37277, n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37285,
    n37286, n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294,
    n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303,
    n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312,
    n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
    n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330,
    n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339,
    n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348,
    n37349, n37350, n37351, n37352, n37353, n37354, n37355, n37356, n37357,
    n37358, n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366,
    n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375,
    n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384,
    n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
    n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402,
    n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411,
    n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420,
    n37421, n37422, n37423, n37424, n37425, n37426, n37427, n37428, n37429,
    n37430, n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438,
    n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447,
    n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456,
    n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
    n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474,
    n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483,
    n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492,
    n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500, n37501,
    n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510,
    n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519,
    n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528,
    n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
    n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546,
    n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555,
    n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564,
    n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573,
    n37574, n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582,
    n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591,
    n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600,
    n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
    n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618,
    n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627,
    n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636,
    n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645,
    n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654,
    n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663,
    n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672,
    n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
    n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690,
    n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699,
    n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708,
    n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717,
    n37718, n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726,
    n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735,
    n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744,
    n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
    n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762,
    n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771,
    n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780,
    n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789,
    n37790, n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798,
    n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807,
    n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816,
    n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
    n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834,
    n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843,
    n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852,
    n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861,
    n37862, n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870,
    n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879,
    n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888,
    n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
    n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906,
    n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915,
    n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924,
    n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933,
    n37934, n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942,
    n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951,
    n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960,
    n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
    n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978,
    n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987,
    n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996,
    n37997, n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005,
    n38006, n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014,
    n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023,
    n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032,
    n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
    n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050,
    n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059,
    n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068,
    n38069, n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077,
    n38078, n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086,
    n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095,
    n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104,
    n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
    n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122,
    n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131,
    n38132, n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140,
    n38141, n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149,
    n38150, n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158,
    n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167,
    n38168, n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176,
    n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
    n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194,
    n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203,
    n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212,
    n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221,
    n38222, n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230,
    n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239,
    n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248,
    n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
    n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266,
    n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275,
    n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284,
    n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293,
    n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302,
    n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311,
    n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320,
    n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
    n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338,
    n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347,
    n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356,
    n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365,
    n38366, n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374,
    n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383,
    n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392,
    n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
    n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410,
    n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419,
    n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428,
    n38429, n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437,
    n38438, n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446,
    n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455,
    n38456, n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464,
    n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
    n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482,
    n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491,
    n38492, n38493, n38494, n38495, n38496, n38497, n38498, n38499, n38500,
    n38501, n38502, n38503, n38504, n38505, n38506, n38507, n38508, n38509,
    n38510, n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518,
    n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527,
    n38528, n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536,
    n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
    n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554,
    n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563,
    n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571, n38572,
    n38573, n38574, n38575, n38576, n38577, n38578, n38579, n38580, n38581,
    n38582, n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590,
    n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599,
    n38600, n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608,
    n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
    n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626,
    n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635,
    n38636, n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644,
    n38645, n38646, n38647, n38648, n38649, n38650, n38651, n38652, n38653,
    n38654, n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662,
    n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671,
    n38672, n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680,
    n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
    n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698,
    n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707,
    n38708, n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716,
    n38717, n38718, n38719, n38720, n38721, n38722, n38723, n38724, n38725,
    n38726, n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734,
    n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743,
    n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752,
    n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
    n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770,
    n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779,
    n38780, n38781, n38782, n38783, n38784, n38785, n38786, n38787, n38788,
    n38789, n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797,
    n38798, n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806,
    n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815,
    n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824,
    n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
    n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842,
    n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851,
    n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860,
    n38861, n38862, n38863, n38864, n38865, n38866, n38867, n38868, n38869,
    n38870, n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878,
    n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887,
    n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896,
    n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
    n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914,
    n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923,
    n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932,
    n38933, n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941,
    n38942, n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950,
    n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959,
    n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968,
    n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
    n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986,
    n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995,
    n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004,
    n39005, n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013,
    n39014, n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022,
    n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031,
    n39032, n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040,
    n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
    n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058,
    n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067,
    n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076,
    n39077, n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085,
    n39086, n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094,
    n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103,
    n39104, n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112,
    n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
    n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130,
    n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139,
    n39140, n39141, n39142, n39143, n39144, n39145, n39146, n39147, n39148,
    n39149, n39150, n39151, n39152, n39153, n39154, n39155, n39156, n39157,
    n39158, n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166,
    n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175,
    n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184,
    n39185, n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
    n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202,
    n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211,
    n39212, n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220,
    n39221, n39222, n39223, n39224, n39225, n39226, n39227, n39228, n39229,
    n39230, n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238,
    n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247,
    n39248, n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256,
    n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
    n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274,
    n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283,
    n39284, n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292,
    n39293, n39294, n39295, n39296, n39297, n39298, n39299, n39300, n39301,
    n39302, n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310,
    n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319,
    n39320, n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328,
    n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337,
    n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346,
    n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355,
    n39356, n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364,
    n39365, n39366, n39367, n39368, n39369, n39370, n39371, n39372, n39373,
    n39374, n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382,
    n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391,
    n39392, n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400,
    n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409,
    n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418,
    n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427,
    n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436,
    n39437, n39438, n39439, n39440, n39441, n39442, n39443, n39444, n39445,
    n39446, n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454,
    n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463,
    n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472,
    n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481,
    n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490,
    n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499,
    n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508,
    n39509, n39510, n39511, n39512, n39513, n39514, n39515, n39516, n39517,
    n39518, n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526,
    n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535,
    n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
    n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
    n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562,
    n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571,
    n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580,
    n39581, n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589,
    n39590, n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598,
    n39599, n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607,
    n39608, n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616,
    n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
    n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634,
    n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643,
    n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652,
    n39653, n39654, n39655, n39656, n39657, n39658, n39659, n39660, n39661,
    n39662, n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670,
    n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679,
    n39680, n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688,
    n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697,
    n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706,
    n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715,
    n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724,
    n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732, n39733,
    n39734, n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742,
    n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751,
    n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760,
    n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769,
    n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778,
    n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787,
    n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796,
    n39797, n39798, n39799, n39800, n39801, n39802, n39803, n39804, n39805,
    n39806, n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814,
    n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823,
    n39824, n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832,
    n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
    n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850,
    n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859,
    n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868,
    n39869, n39870, n39871, n39872, n39873, n39874, n39875, n39876, n39877,
    n39878, n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886,
    n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895,
    n39896, n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904,
    n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
    n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922,
    n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931,
    n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940,
    n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948, n39949,
    n39950, n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958,
    n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967,
    n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976,
    n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
    n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994,
    n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003,
    n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012,
    n40013, n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021,
    n40022, n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030,
    n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039,
    n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048,
    n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
    n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066,
    n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075,
    n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084,
    n40085, n40086, n40087, n40088, n40089, n40090, n40091, n40092, n40093,
    n40094, n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102,
    n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111,
    n40112, n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120,
    n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
    n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138,
    n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147,
    n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156,
    n40157, n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165,
    n40166, n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174,
    n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183,
    n40184, n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192,
    n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
    n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210,
    n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219,
    n40220, n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228,
    n40229, n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237,
    n40238, n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246,
    n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255,
    n40256, n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264,
    n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273,
    n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282,
    n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291,
    n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300,
    n40301, n40302, n40303, n40304, n40305, n40306, n40307, n40308, n40309,
    n40310, n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318,
    n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327,
    n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336,
    n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345,
    n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354,
    n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363,
    n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372,
    n40373, n40374, n40375, n40376, n40377, n40378, n40379, n40380, n40381,
    n40382, n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390,
    n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399,
    n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408,
    n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417,
    n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426,
    n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435,
    n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444,
    n40445, n40446, n40447, n40448, n40449, n40450, n40451, n40452, n40453,
    n40454, n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462,
    n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471,
    n40472, n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480,
    n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489,
    n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498,
    n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507,
    n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516,
    n40517, n40518, n40519, n40520, n40521, n40522, n40523, n40524, n40525,
    n40526, n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534,
    n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543,
    n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552,
    n40553, n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561,
    n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570,
    n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579,
    n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588,
    n40589, n40590, n40591, n40592, n40593, n40594, n40595, n40596, n40597,
    n40598, n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606,
    n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615,
    n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624,
    n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
    n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642,
    n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651,
    n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660,
    n40661, n40662, n40663, n40664, n40665, n40666, n40667, n40668, n40669,
    n40670, n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678,
    n40679, n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687,
    n40688, n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696,
    n40697, n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705,
    n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714,
    n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723,
    n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732,
    n40733, n40734, n40735, n40736, n40737, n40738, n40739, n40740, n40741,
    n40742, n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750,
    n40751, n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759,
    n40760, n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768,
    n40769, n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777,
    n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786,
    n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795,
    n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804,
    n40805, n40806, n40807, n40808, n40809, n40810, n40811, n40812, n40813,
    n40814, n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822,
    n40823, n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831,
    n40832, n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840,
    n40841, n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849,
    n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858,
    n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867,
    n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876,
    n40877, n40878, n40879, n40880, n40881, n40882, n40883, n40884, n40885,
    n40886, n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894,
    n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903,
    n40904, n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912,
    n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921,
    n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930,
    n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939,
    n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948,
    n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957,
    n40958, n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966,
    n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975,
    n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984,
    n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
    n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002,
    n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011,
    n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020,
    n41021, n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029,
    n41030, n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038,
    n41039, n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047,
    n41048, n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056,
    n41057, n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065,
    n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074,
    n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083,
    n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092,
    n41093, n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101,
    n41102, n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110,
    n41111, n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119,
    n41120, n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128,
    n41129, n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137,
    n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146,
    n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155,
    n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164,
    n41165, n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173,
    n41174, n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182,
    n41183, n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191,
    n41192, n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200,
    n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209,
    n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218,
    n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227,
    n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236,
    n41237, n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245,
    n41246, n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254,
    n41255, n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263,
    n41264, n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272,
    n41273, n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281,
    n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290,
    n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299,
    n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308,
    n41309, n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317,
    n41318, n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326,
    n41327, n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335,
    n41336, n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344,
    n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353,
    n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362,
    n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371,
    n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380,
    n41381, n41382, n41383, n41384, n41385, n41386, n41387, n41388, n41389,
    n41390, n41391, n41392, n41393, n41394, n41395, n41396, n41397, n41398,
    n41399, n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407,
    n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416,
    n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425,
    n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434,
    n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443,
    n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452,
    n41453, n41454, n41455, n41456, n41457, n41458, n41459, n41460, n41461,
    n41462, n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470,
    n41471, n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479,
    n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488,
    n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497,
    n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506,
    n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515,
    n41516, n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524,
    n41525, n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533,
    n41534, n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542,
    n41543, n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551,
    n41552, n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560,
    n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569,
    n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578,
    n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587,
    n41588, n41589, n41590, n41591, n41592, n41593, n41594, n41595, n41596,
    n41597, n41598, n41599, n41600, n41601, n41602, n41603, n41604, n41605,
    n41606, n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614,
    n41615, n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623,
    n41624, n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632,
    n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641,
    n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650,
    n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659,
    n41660, n41661, n41662, n41663, n41664, n41665, n41666, n41667, n41668,
    n41669, n41670, n41671, n41672, n41673, n41674, n41675, n41676, n41677,
    n41678, n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686,
    n41687, n41688, n41689, n41690, n41691, n41692, n41693, n41694, n41695,
    n41696, n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704,
    n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713,
    n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722,
    n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731,
    n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739, n41740,
    n41741, n41742, n41743, n41744, n41745, n41746, n41747, n41748, n41749,
    n41750, n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758,
    n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767,
    n41768, n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776,
    n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785,
    n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794,
    n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803,
    n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812,
    n41813, n41814, n41815, n41816, n41817, n41818, n41819, n41820, n41821,
    n41822, n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830,
    n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838, n41839,
    n41840, n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848,
    n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857,
    n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866,
    n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875,
    n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884,
    n41885, n41886, n41887, n41888, n41889, n41890, n41891, n41892, n41893,
    n41894, n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902,
    n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911,
    n41912, n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920,
    n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929,
    n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938,
    n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947,
    n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956,
    n41957, n41958, n41959, n41960, n41961, n41962, n41963, n41964, n41965,
    n41966, n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974,
    n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983,
    n41984, n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992,
    n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001,
    n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010,
    n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019,
    n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028,
    n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036, n42037,
    n42038, n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046,
    n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054, n42055,
    n42056, n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064,
    n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073,
    n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082,
    n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091,
    n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100,
    n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42108, n42109,
    n42110, n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118,
    n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126, n42127,
    n42128, n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136,
    n42137, n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145,
    n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154,
    n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163,
    n42164, n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172,
    n42173, n42174, n42175, n42176, n42177, n42178, n42179, n42180, n42181,
    n42182, n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190,
    n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198, n42199,
    n42200, n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208,
    n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217,
    n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226,
    n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235,
    n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244,
    n42245, n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253,
    n42254, n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262,
    n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270, n42271,
    n42272, n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280,
    n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289,
    n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298,
    n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307,
    n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316,
    n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324, n42325,
    n42326, n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334,
    n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342, n42343,
    n42344, n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352,
    n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361,
    n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370,
    n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379,
    n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388,
    n42389, n42390, n42391, n42392, n42393, n42394, n42395, n42396, n42397,
    n42398, n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406,
    n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414, n42415,
    n42416, n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424,
    n42425, n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433,
    n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442,
    n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451,
    n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460,
    n42461, n42462, n42463, n42464, n42465, n42466, n42467, n42468, n42469,
    n42470, n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478,
    n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486, n42487,
    n42488, n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496,
    n42497, n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505,
    n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514,
    n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523,
    n42524, n42525, n42526, n42527, n42528, n42529, n42530, n42531, n42532,
    n42533, n42534, n42535, n42536, n42537, n42538, n42539, n42540, n42541,
    n42542, n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550,
    n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558, n42559,
    n42560, n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568,
    n42569, n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577,
    n42578, n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586,
    n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595,
    n42596, n42597, n42598, n42599, n42600, n42601, n42602, n42603, n42604,
    n42605, n42606, n42607, n42608, n42609, n42610, n42611, n42612, n42613,
    n42614, n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622,
    n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630, n42631,
    n42632, n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640,
    n42641, n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649,
    n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658,
    n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667,
    n42668, n42669, n42670, n42671, n42672, n42673, n42674, n42675, n42676,
    n42677, n42678, n42679, n42680, n42681, n42682, n42683, n42684, n42685,
    n42686, n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694,
    n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702, n42703,
    n42704, n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712,
    n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721,
    n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730,
    n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739,
    n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748,
    n42749, n42750, n42751, n42752, n42753, n42754, n42755, n42756, n42757,
    n42758, n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766,
    n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775,
    n42776, n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784,
    n42785, n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793,
    n42794, n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802,
    n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811,
    n42812, n42813, n42814, n42815, n42816, n42817, n42818, n42819, n42820,
    n42821, n42822, n42823, n42824, n42825, n42826, n42827, n42828, n42829,
    n42830, n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838,
    n42839, n42840, n42841, n42842, n42843, n42844, n42845, n42846, n42847,
    n42848, n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856,
    n42857, n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865,
    n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874,
    n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883,
    n42884, n42885, n42886, n42887, n42888, n42889, n42890, n42891, n42892,
    n42893, n42894, n42895, n42896, n42897, n42898, n42899, n42900, n42901,
    n42902, n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910,
    n42911, n42912, n42913, n42914, n42915, n42916, n42917, n42918, n42919,
    n42920, n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928,
    n42929, n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937,
    n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946,
    n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955,
    n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963, n42964,
    n42965, n42966, n42967, n42968, n42969, n42970, n42971, n42972, n42973,
    n42974, n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982,
    n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991,
    n42992, n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000,
    n43001, n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009,
    n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018,
    n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027,
    n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035, n43036,
    n43037, n43038, n43039, n43040, n43041, n43042, n43043, n43044, n43045,
    n43046, n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054,
    n43055, n43056, n43057, n43058, n43059, n43060, n43061, n43062, n43063,
    n43064, n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072,
    n43073, n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081,
    n43082, n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090,
    n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099,
    n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107, n43108,
    n43109, n43110, n43111, n43112, n43113, n43114, n43115, n43116, n43117,
    n43118, n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126,
    n43127, n43128, n43129, n43130, n43131, n43132, n43133, n43134, n43135,
    n43136, n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144,
    n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153,
    n43154, n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162,
    n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171,
    n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179, n43180,
    n43181, n43182, n43183, n43184, n43185, n43186, n43187, n43188, n43189,
    n43190, n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198,
    n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206, n43207,
    n43208, n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216,
    n43217, n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225,
    n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234,
    n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243,
    n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251, n43252,
    n43253, n43254, n43255, n43256, n43257, n43258, n43259, n43260, n43261,
    n43262, n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270,
    n43271, n43272, n43273, n43275, n43276, n43277, n43278, n43280, n43281,
    n43282, n43283, n43285, n43286, n43287, n43289, n43290, n43291, n43293,
    n43294, n43295, n43297, n43298, n43299, n43301, n43302, n43303, n43305,
    n43306, n43307, n43309, n43310, n43311, n43313, n43314, n43315, n43317,
    n43318, n43319, n43321, n43322, n43323, n43325, n43326, n43327, n43329,
    n43330, n43331, n43333, n43334, n43335, n43337, n43338, n43339, n43341,
    n43342, n43343, n43345, n43346, n43347, n43349, n43350, n43351, n43353,
    n43354, n43355, n43357, n43358, n43359, n43361, n43362, n43363, n43365,
    n43366, n43367, n43369, n43370, n43371, n43373, n43374, n43375, n43377,
    n43378, n43379, n43381, n43382, n43383, n43385, n43386, n43387, n43389,
    n43390, n43391, n43393, n43394, n43395, n43397, n43398, n43399, n43401,
    n43402, n43403, n43405, n43406, n43407, n43409, n43410, n43411, n43413,
    n43414, n43415, n43417, n43418, n43419, n43421, n43422, n43423, n43425,
    n43426, n43427, n43429, n43430, n43431, n43433, n43434, n43435, n43437,
    n43438, n43439, n43441, n43442, n43443, n43445, n43446, n43447, n43449,
    n43450, n43451, n43453, n43454, n43455, n43457, n43458, n43459, n43461,
    n43462, n43463, n43465, n43466, n43467, n43469, n43470, n43471, n43473,
    n43474, n43475, n43477, n43478, n43479, n43481, n43482, n43483, n43485,
    n43486, n43487, n43489, n43490, n43491, n43493, n43494, n43495, n43497,
    n43498, n43499, n43501, n43502, n43503, n43505, n43506, n43507, n43509,
    n43510, n43511, n43513, n43514, n43515, n43517, n43518, n43519, n43521,
    n43522, n43523, n43525, n43526;
  jnot g00000(.din(b61 ), .dout(n256));
  jnot g00001(.din(a62 ), .dout(n257));
  jnot g00002(.din(b1 ), .dout(n258));
  jand g00003(.dina(b0 ), .dinb(n257), .dout(n259));
  jnot g00004(.din(n259), .dout(n260));
  jand g00005(.dina(n260), .dinb(n258), .dout(n261));
  jor  g00006(.dina(b63 ), .dinb(b62 ), .dout(n262));
  jor  g00007(.dina(n262), .dinb(b61 ), .dout(n263));
  jor  g00008(.dina(n263), .dinb(b60 ), .dout(n264));
  jor  g00009(.dina(b56 ), .dinb(b53 ), .dout(n265));
  jor  g00010(.dina(b59 ), .dinb(b52 ), .dout(n266));
  jor  g00011(.dina(n266), .dinb(n265), .dout(n267));
  jor  g00012(.dina(b58 ), .dinb(b57 ), .dout(n268));
  jor  g00013(.dina(b55 ), .dinb(b54 ), .dout(n269));
  jor  g00014(.dina(n269), .dinb(n268), .dout(n270));
  jor  g00015(.dina(n270), .dinb(n267), .dout(n271));
  jor  g00016(.dina(n271), .dinb(n264), .dout(n272));
  jor  g00017(.dina(b47 ), .dinb(b46 ), .dout(n273));
  jor  g00018(.dina(n273), .dinb(b45 ), .dout(n274));
  jor  g00019(.dina(b51 ), .dinb(b50 ), .dout(n275));
  jor  g00020(.dina(b49 ), .dinb(b48 ), .dout(n276));
  jor  g00021(.dina(n276), .dinb(b44 ), .dout(n277));
  jor  g00022(.dina(n277), .dinb(n275), .dout(n278));
  jor  g00023(.dina(n278), .dinb(n274), .dout(n279));
  jor  g00024(.dina(n279), .dinb(n272), .dout(n280));
  jnot g00025(.din(b42 ), .dout(n281));
  jnot g00026(.din(b43 ), .dout(n282));
  jand g00027(.dina(n282), .dinb(n281), .dout(n283));
  jnot g00028(.din(b40 ), .dout(n284));
  jnot g00029(.din(b41 ), .dout(n285));
  jand g00030(.dina(n285), .dinb(n284), .dout(n286));
  jand g00031(.dina(n286), .dinb(n283), .dout(n287));
  jnot g00032(.din(n287), .dout(n288));
  jor  g00033(.dina(n288), .dinb(n280), .dout(n289));
  jnot g00034(.din(b38 ), .dout(n290));
  jnot g00035(.din(b39 ), .dout(n291));
  jand g00036(.dina(n291), .dinb(n290), .dout(n292));
  jnot g00037(.din(b36 ), .dout(n293));
  jnot g00038(.din(b37 ), .dout(n294));
  jand g00039(.dina(n294), .dinb(n293), .dout(n295));
  jand g00040(.dina(n295), .dinb(n292), .dout(n296));
  jnot g00041(.din(b33 ), .dout(n297));
  jnot g00042(.din(b34 ), .dout(n298));
  jand g00043(.dina(n298), .dinb(n297), .dout(n299));
  jnot g00044(.din(b32 ), .dout(n300));
  jnot g00045(.din(b35 ), .dout(n301));
  jand g00046(.dina(n301), .dinb(n300), .dout(n302));
  jand g00047(.dina(n302), .dinb(n299), .dout(n303));
  jand g00048(.dina(n303), .dinb(n296), .dout(n304));
  jnot g00049(.din(n304), .dout(n305));
  jor  g00050(.dina(n305), .dinb(n289), .dout(n306));
  jor  g00051(.dina(b27 ), .dinb(b26 ), .dout(n307));
  jor  g00052(.dina(b25 ), .dinb(b24 ), .dout(n308));
  jor  g00053(.dina(n308), .dinb(n307), .dout(n309));
  jor  g00054(.dina(b31 ), .dinb(b30 ), .dout(n310));
  jor  g00055(.dina(b29 ), .dinb(b28 ), .dout(n311));
  jor  g00056(.dina(n311), .dinb(n310), .dout(n312));
  jor  g00057(.dina(n312), .dinb(n309), .dout(n313));
  jor  g00058(.dina(b22 ), .dinb(b21 ), .dout(n314));
  jor  g00059(.dina(n314), .dinb(b20 ), .dout(n315));
  jor  g00060(.dina(n315), .dinb(b23 ), .dout(n316));
  jor  g00061(.dina(n316), .dinb(n313), .dout(n317));
  jor  g00062(.dina(n317), .dinb(n306), .dout(n318));
  jor  g00063(.dina(b19 ), .dinb(b18 ), .dout(n319));
  jor  g00064(.dina(b17 ), .dinb(b16 ), .dout(n320));
  jor  g00065(.dina(n320), .dinb(n319), .dout(n321));
  jor  g00066(.dina(n321), .dinb(n318), .dout(n322));
  jnot g00067(.din(b8 ), .dout(n323));
  jnot g00068(.din(b9 ), .dout(n324));
  jnot g00069(.din(b10 ), .dout(n325));
  jand g00070(.dina(n325), .dinb(n324), .dout(n326));
  jand g00071(.dina(n326), .dinb(n323), .dout(n327));
  jnot g00072(.din(n327), .dout(n328));
  jor  g00073(.dina(b15 ), .dinb(b14 ), .dout(n329));
  jor  g00074(.dina(b13 ), .dinb(b12 ), .dout(n330));
  jor  g00075(.dina(n330), .dinb(n329), .dout(n331));
  jor  g00076(.dina(n331), .dinb(b11 ), .dout(n332));
  jor  g00077(.dina(n332), .dinb(n328), .dout(n333));
  jnot g00078(.din(b6 ), .dout(n334));
  jnot g00079(.din(b7 ), .dout(n335));
  jand g00080(.dina(n335), .dinb(n334), .dout(n336));
  jnot g00081(.din(b4 ), .dout(n337));
  jnot g00082(.din(b5 ), .dout(n338));
  jand g00083(.dina(n338), .dinb(n337), .dout(n339));
  jand g00084(.dina(n339), .dinb(n336), .dout(n340));
  jnot g00085(.din(n340), .dout(n341));
  jor  g00086(.dina(n341), .dinb(n333), .dout(n342));
  jor  g00087(.dina(n342), .dinb(n322), .dout(n343));
  jnot g00088(.din(b3 ), .dout(n344));
  jand g00089(.dina(n344), .dinb(b0 ), .dout(n345));
  jnot g00090(.din(a63 ), .dout(n346));
  jand g00091(.dina(b0 ), .dinb(n346), .dout(n347));
  jnot g00092(.din(b2 ), .dout(n348));
  jand g00093(.dina(n348), .dinb(n258), .dout(n349));
  jnot g00094(.din(n349), .dout(n350));
  jor  g00095(.dina(n350), .dinb(n347), .dout(n351));
  jnot g00096(.din(n351), .dout(n352));
  jand g00097(.dina(n352), .dinb(n345), .dout(n353));
  jnot g00098(.din(n353), .dout(n354));
  jor  g00099(.dina(n354), .dinb(n343), .dout(n355));
  jand g00100(.dina(n259), .dinb(b1 ), .dout(n356));
  jor  g00101(.dina(n356), .dinb(n346), .dout(n357));
  jnot g00102(.din(n357), .dout(n358));
  jand g00103(.dina(n358), .dinb(n355), .dout(n359));
  jor  g00104(.dina(n359), .dinb(n261), .dout(n360));
  jand g00105(.dina(n344), .dinb(n348), .dout(n361));
  jnot g00106(.din(b57 ), .dout(n362));
  jnot g00107(.din(b58 ), .dout(n363));
  jand g00108(.dina(n363), .dinb(n362), .dout(n364));
  jnot g00109(.din(b59 ), .dout(n365));
  jnot g00110(.din(b60 ), .dout(n366));
  jnot g00111(.din(b62 ), .dout(n367));
  jnot g00112(.din(b63 ), .dout(n368));
  jand g00113(.dina(n368), .dinb(n367), .dout(n369));
  jand g00114(.dina(n369), .dinb(n256), .dout(n370));
  jand g00115(.dina(n370), .dinb(n366), .dout(n371));
  jand g00116(.dina(n371), .dinb(n365), .dout(n372));
  jand g00117(.dina(n372), .dinb(n364), .dout(n373));
  jnot g00118(.din(b53 ), .dout(n374));
  jnot g00119(.din(b56 ), .dout(n375));
  jnot g00120(.din(b54 ), .dout(n376));
  jnot g00121(.din(b55 ), .dout(n377));
  jand g00122(.dina(n377), .dinb(n376), .dout(n378));
  jand g00123(.dina(n378), .dinb(n375), .dout(n379));
  jand g00124(.dina(n379), .dinb(n374), .dout(n380));
  jand g00125(.dina(n380), .dinb(n373), .dout(n381));
  jnot g00126(.din(n275), .dout(n382));
  jnot g00127(.din(b49 ), .dout(n383));
  jnot g00128(.din(b52 ), .dout(n384));
  jand g00129(.dina(n384), .dinb(n383), .dout(n385));
  jand g00130(.dina(n385), .dinb(n382), .dout(n386));
  jand g00131(.dina(n386), .dinb(n381), .dout(n387));
  jand g00132(.dina(n293), .dinb(n301), .dout(n388));
  jand g00133(.dina(n290), .dinb(n294), .dout(n389));
  jand g00134(.dina(n389), .dinb(n388), .dout(n390));
  jand g00135(.dina(n284), .dinb(n291), .dout(n391));
  jand g00136(.dina(n391), .dinb(n299), .dout(n392));
  jand g00137(.dina(n392), .dinb(n390), .dout(n393));
  jnot g00138(.din(n274), .dout(n394));
  jand g00139(.dina(n281), .dinb(n285), .dout(n395));
  jnot g00140(.din(b48 ), .dout(n396));
  jnot g00141(.din(b44 ), .dout(n397));
  jand g00142(.dina(n397), .dinb(n282), .dout(n398));
  jand g00143(.dina(n398), .dinb(n396), .dout(n399));
  jand g00144(.dina(n399), .dinb(n395), .dout(n400));
  jand g00145(.dina(n400), .dinb(n394), .dout(n401));
  jand g00146(.dina(n401), .dinb(n393), .dout(n402));
  jand g00147(.dina(n402), .dinb(n387), .dout(n403));
  jnot g00148(.din(n314), .dout(n404));
  jnot g00149(.din(b23 ), .dout(n405));
  jnot g00150(.din(b24 ), .dout(n406));
  jand g00151(.dina(n406), .dinb(n405), .dout(n407));
  jand g00152(.dina(n407), .dinb(n404), .dout(n408));
  jnot g00153(.din(b27 ), .dout(n409));
  jnot g00154(.din(b28 ), .dout(n410));
  jand g00155(.dina(n410), .dinb(n409), .dout(n411));
  jnot g00156(.din(b25 ), .dout(n412));
  jnot g00157(.din(b26 ), .dout(n413));
  jand g00158(.dina(n413), .dinb(n412), .dout(n414));
  jand g00159(.dina(n414), .dinb(n411), .dout(n415));
  jnot g00160(.din(b19 ), .dout(n416));
  jnot g00161(.din(b20 ), .dout(n417));
  jand g00162(.dina(n417), .dinb(n416), .dout(n418));
  jand g00163(.dina(n418), .dinb(n415), .dout(n419));
  jand g00164(.dina(n419), .dinb(n408), .dout(n420));
  jnot g00165(.din(b17 ), .dout(n421));
  jnot g00166(.din(b18 ), .dout(n422));
  jand g00167(.dina(n422), .dinb(n421), .dout(n423));
  jnot g00168(.din(b31 ), .dout(n424));
  jand g00169(.dina(n300), .dinb(n424), .dout(n425));
  jnot g00170(.din(b29 ), .dout(n426));
  jnot g00171(.din(b30 ), .dout(n427));
  jand g00172(.dina(n427), .dinb(n426), .dout(n428));
  jand g00173(.dina(n428), .dinb(n425), .dout(n429));
  jand g00174(.dina(n429), .dinb(n423), .dout(n430));
  jand g00175(.dina(n430), .dinb(n420), .dout(n431));
  jnot g00176(.din(b15 ), .dout(n432));
  jnot g00177(.din(b16 ), .dout(n433));
  jand g00178(.dina(n433), .dinb(n432), .dout(n434));
  jnot g00179(.din(b13 ), .dout(n435));
  jnot g00180(.din(b14 ), .dout(n436));
  jand g00181(.dina(n436), .dinb(n435), .dout(n437));
  jand g00182(.dina(n437), .dinb(n434), .dout(n438));
  jnot g00183(.din(b11 ), .dout(n439));
  jnot g00184(.din(b12 ), .dout(n440));
  jand g00185(.dina(n440), .dinb(n439), .dout(n441));
  jand g00186(.dina(n441), .dinb(n326), .dout(n442));
  jand g00187(.dina(n442), .dinb(n438), .dout(n443));
  jand g00188(.dina(n443), .dinb(n431), .dout(n444));
  jand g00189(.dina(n444), .dinb(n403), .dout(n445));
  jand g00190(.dina(n334), .dinb(n338), .dout(n446));
  jand g00191(.dina(n323), .dinb(n335), .dout(n447));
  jand g00192(.dina(n447), .dinb(n446), .dout(n448));
  jand g00193(.dina(n337), .dinb(b0 ), .dout(n449));
  jand g00194(.dina(n449), .dinb(n448), .dout(n450));
  jand g00195(.dina(n450), .dinb(n445), .dout(n451));
  jand g00196(.dina(n451), .dinb(n361), .dout(n452));
  jand g00197(.dina(n452), .dinb(n360), .dout(n453));
  jor  g00198(.dina(n453), .dinb(n257), .dout(n454));
  jor  g00199(.dina(n313), .dinb(n306), .dout(n455));
  jor  g00200(.dina(n321), .dinb(n316), .dout(n456));
  jnot g00201(.din(n342), .dout(n458));
  jand g00202(.dina(n361), .dinb(n458), .dout(n459));
  jnot g00203(.din(n459), .dout(n460));
  jor  g00204(.dina(n460), .dinb(n322), .dout(n461));
  jnot g00205(.din(a61 ), .dout(n467));
  jand g00206(.dina(b0 ), .dinb(n467), .dout(n468));
  jand g00207(.dina(n468), .dinb(b1 ), .dout(n469));
  jor  g00208(.dina(n469), .dinb(n454), .dout(n470));
  jnot g00209(.din(n468), .dout(n471));
  jand g00210(.dina(n471), .dinb(n258), .dout(n472));
  jnot g00211(.din(n472), .dout(n473));
  jand g00212(.dina(n473), .dinb(n470), .dout(n474));
  jor  g00213(.dina(n474), .dinb(b2 ), .dout(n475));
  jnot g00214(.din(n461), .dout(n476));
  jnot g00215(.din(n261), .dout(n477));
  jand g00216(.dina(n358), .dinb(n477), .dout(n478));
  jand g00217(.dina(n478), .dinb(n476), .dout(n479));
  jor  g00218(.dina(n479), .dinb(n346), .dout(n480));
  jnot g00219(.din(n480), .dout(n481));
  jand g00220(.dina(n481), .dinb(n355), .dout(n482));
  jnot g00221(.din(n482), .dout(n483));
  jand g00222(.dina(n474), .dinb(b2 ), .dout(n484));
  jor  g00223(.dina(n484), .dinb(n483), .dout(n485));
  jand g00224(.dina(n485), .dinb(n475), .dout(n486));
  jor  g00225(.dina(n322), .dinb(n333), .dout(n487));
  jand g00226(.dina(n345), .dinb(n340), .dout(n488));
  jnot g00227(.din(n488), .dout(n489));
  jor  g00228(.dina(n489), .dinb(n487), .dout(n490));
  jor  g00229(.dina(n490), .dinb(n486), .dout(n491));
  jand g00230(.dina(n491), .dinb(a61 ), .dout(n492));
  jnot g00231(.din(n486), .dout(n493));
  jand g00232(.dina(n337), .dinb(n344), .dout(n494));
  jand g00233(.dina(n494), .dinb(n448), .dout(n495));
  jand g00234(.dina(n495), .dinb(n445), .dout(n496));
  jand g00235(.dina(n496), .dinb(n468), .dout(n497));
  jand g00236(.dina(n497), .dinb(n493), .dout(n498));
  jor  g00237(.dina(n498), .dinb(n492), .dout(n499));
  jnot g00238(.din(n343), .dout(n500));
  jnot g00239(.din(n484), .dout(n501));
  jand g00240(.dina(n496), .dinb(n475), .dout(n502));
  jand g00241(.dina(n502), .dinb(n501), .dout(n503));
  jor  g00242(.dina(n503), .dinb(n483), .dout(n504));
  jand g00243(.dina(n504), .dinb(b3 ), .dout(n505));
  jnot g00244(.din(n505), .dout(n506));
  jnot g00245(.din(n504), .dout(n507));
  jand g00246(.dina(n507), .dinb(n344), .dout(n508));
  jnot g00247(.din(n454), .dout(n509));
  jnot g00248(.din(b47 ), .dout(n510));
  jand g00249(.dina(n396), .dinb(n510), .dout(n511));
  jand g00250(.dina(n511), .dinb(n387), .dout(n512));
  jnot g00251(.din(b45 ), .dout(n513));
  jnot g00252(.din(b46 ), .dout(n514));
  jand g00253(.dina(n514), .dinb(n513), .dout(n515));
  jand g00254(.dina(n515), .dinb(n512), .dout(n516));
  jand g00255(.dina(n516), .dinb(n398), .dout(n517));
  jand g00256(.dina(n517), .dinb(n395), .dout(n518));
  jxor g00257(.dina(n468), .dinb(b1 ), .dout(n520));
  jand g00258(.dina(n520), .dinb(n495), .dout(n521));
  jand g00259(.dina(n521), .dinb(n444), .dout(n522));
  jand g00260(.dina(n522), .dinb(n403), .dout(n523));
  jnot g00261(.din(n523), .dout(n524));
  jor  g00262(.dina(n524), .dinb(n486), .dout(n525));
  jand g00263(.dina(n525), .dinb(n509), .dout(n526));
  jand g00264(.dina(n520), .dinb(n496), .dout(n527));
  jand g00265(.dina(n527), .dinb(n454), .dout(n528));
  jand g00266(.dina(n528), .dinb(n493), .dout(n529));
  jor  g00267(.dina(n529), .dinb(n526), .dout(n530));
  jand g00268(.dina(n530), .dinb(n348), .dout(n531));
  jor  g00269(.dina(n530), .dinb(n348), .dout(n532));
  jnot g00270(.din(a60 ), .dout(n533));
  jand g00271(.dina(b0 ), .dinb(n533), .dout(n534));
  jand g00272(.dina(n534), .dinb(b1 ), .dout(n535));
  jnot g00273(.din(n535), .dout(n536));
  jand g00274(.dina(n536), .dinb(n499), .dout(n537));
  jnot g00275(.din(n534), .dout(n538));
  jand g00276(.dina(n538), .dinb(n258), .dout(n539));
  jor  g00277(.dina(n539), .dinb(n537), .dout(n540));
  jand g00278(.dina(n540), .dinb(n532), .dout(n541));
  jor  g00279(.dina(n541), .dinb(n531), .dout(n542));
  jor  g00280(.dina(n542), .dinb(n508), .dout(n543));
  jand g00281(.dina(n543), .dinb(n506), .dout(n544));
  jand g00282(.dina(n544), .dinb(n500), .dout(quotient60 ));
  jxor g00283(.dina(n534), .dinb(b1 ), .dout(n546));
  jand g00284(.dina(n546), .dinb(quotient60 ), .dout(n547));
  jxor g00285(.dina(n547), .dinb(n499), .dout(n548));
  jand g00286(.dina(n2457), .dinb(n408), .dout(n551));
  jand g00287(.dina(n447), .dinb(n443), .dout(n554));
  jand g00288(.dina(n554), .dinb(n988), .dout(n555));
  jand g00289(.dina(n555), .dinb(n446), .dout(n556));
  jnot g00290(.din(n556), .dout(n557));
  jnot g00291(.din(quotient60 ), .dout(n558));
  jand g00292(.dina(n540), .dinb(n348), .dout(n559));
  jnot g00293(.din(n532), .dout(n563));
  jnot g00294(.din(n540), .dout(n564));
  jand g00295(.dina(n564), .dinb(n563), .dout(n565));
  jor  g00296(.dina(n565), .dinb(n542), .dout(n566));
  jor  g00297(.dina(n566), .dinb(n558), .dout(n567));
  jor  g00298(.dina(n18592), .dinb(b3 ), .dout(n569));
  jand g00299(.dina(n548), .dinb(n348), .dout(n571));
  jnot g00300(.din(n571), .dout(n572));
  jor  g00301(.dina(n548), .dinb(n348), .dout(n573));
  jnot g00302(.din(n573), .dout(n574));
  jand g00303(.dina(n544), .dinb(n451), .dout(n575));
  jor  g00304(.dina(n575), .dinb(n533), .dout(n576));
  jnot g00305(.din(n333), .dout(n577));
  jand g00306(.dina(n375), .dinb(n374), .dout(n578));
  jand g00307(.dina(n365), .dinb(n384), .dout(n579));
  jand g00308(.dina(n579), .dinb(n578), .dout(n580));
  jand g00309(.dina(n378), .dinb(n364), .dout(n581));
  jand g00310(.dina(n581), .dinb(n580), .dout(n582));
  jand g00311(.dina(n582), .dinb(n371), .dout(n583));
  jand g00312(.dina(n383), .dinb(n396), .dout(n584));
  jand g00313(.dina(n584), .dinb(n397), .dout(n585));
  jand g00314(.dina(n585), .dinb(n382), .dout(n586));
  jand g00315(.dina(n586), .dinb(n394), .dout(n587));
  jand g00316(.dina(n587), .dinb(n583), .dout(n588));
  jand g00317(.dina(n287), .dinb(n588), .dout(n589));
  jand g00318(.dina(n304), .dinb(n589), .dout(n590));
  jnot g00319(.din(n313), .dout(n591));
  jand g00320(.dina(n591), .dinb(n590), .dout(n592));
  jnot g00321(.din(n456), .dout(n593));
  jand g00322(.dina(n593), .dinb(n592), .dout(n594));
  jand g00323(.dina(n594), .dinb(n577), .dout(n595));
  jand g00324(.dina(n534), .dinb(n340), .dout(n596));
  jand g00325(.dina(n596), .dinb(n595), .dout(n597));
  jand g00326(.dina(n597), .dinb(n544), .dout(n598));
  jnot g00327(.din(n598), .dout(n599));
  jand g00328(.dina(n599), .dinb(n576), .dout(n600));
  jnot g00329(.din(a59 ), .dout(n601));
  jand g00330(.dina(b0 ), .dinb(n601), .dout(n602));
  jand g00331(.dina(n602), .dinb(b1 ), .dout(n603));
  jor  g00332(.dina(n603), .dinb(n600), .dout(n604));
  jnot g00333(.din(n602), .dout(n605));
  jand g00334(.dina(n605), .dinb(n258), .dout(n606));
  jnot g00335(.din(n606), .dout(n607));
  jand g00336(.dina(n607), .dinb(n604), .dout(n608));
  jor  g00337(.dina(n608), .dinb(n574), .dout(n609));
  jand g00338(.dina(n609), .dinb(n572), .dout(n610));
  jor  g00339(.dina(n610), .dinb(n18596), .dout(n611));
  jand g00340(.dina(n611), .dinb(n569), .dout(n612));
  jor  g00341(.dina(n612), .dinb(b4 ), .dout(n613));
  jand g00342(.dina(n558), .dinb(n507), .dout(n614));
  jand g00343(.dina(n508), .dinb(n500), .dout(n615));
  jand g00344(.dina(n615), .dinb(n542), .dout(n616));
  jor  g00345(.dina(n616), .dinb(n614), .dout(n617));
  jnot g00346(.din(n617), .dout(n618));
  jand g00347(.dina(n612), .dinb(b4 ), .dout(n619));
  jor  g00348(.dina(n619), .dinb(n618), .dout(n620));
  jand g00349(.dina(n620), .dinb(n613), .dout(n621));
  jor  g00350(.dina(n621), .dinb(n557), .dout(n622));
  jnot g00351(.din(n608), .dout(n623));
  jand g00352(.dina(n623), .dinb(n348), .dout(n624));
  jor  g00353(.dina(n624), .dinb(n622), .dout(n625));
  jand g00354(.dina(n625), .dinb(n548), .dout(n626));
  jnot g00355(.din(n610), .dout(n627));
  jand g00356(.dina(n608), .dinb(n574), .dout(n628));
  jor  g00357(.dina(n628), .dinb(n627), .dout(n629));
  jor  g00358(.dina(n629), .dinb(n622), .dout(n630));
  jnot g00359(.din(n630), .dout(n631));
  jor  g00360(.dina(n631), .dinb(n626), .dout(n632));
  jnot g00361(.din(n619), .dout(n633));
  jand g00362(.dina(n633), .dinb(n556), .dout(n634));
  jand g00363(.dina(n634), .dinb(n613), .dout(n635));
  jor  g00364(.dina(n635), .dinb(n618), .dout(n636));
  jnot g00365(.din(n636), .dout(n637));
  jand g00366(.dina(n637), .dinb(n556), .dout(n638));
  jand g00367(.dina(n595), .dinb(n336), .dout(n641));
  jand g00368(.dina(n627), .dinb(n344), .dout(n643));
  jor  g00369(.dina(n643), .dinb(n622), .dout(n644));
  jand g00370(.dina(n644), .dinb(n18593), .dout(n645));
  jnot g00371(.din(n645), .dout(n646));
  jnot g00372(.din(n612), .dout(n647));
  jand g00373(.dina(n610), .dinb(n18596), .dout(n648));
  jor  g00374(.dina(n648), .dinb(n647), .dout(n649));
  jor  g00375(.dina(n649), .dinb(n622), .dout(n650));
  jand g00376(.dina(n650), .dinb(n646), .dout(n651));
  jand g00377(.dina(n632), .dinb(n344), .dout(n654));
  jxor g00378(.dina(n602), .dinb(n258), .dout(n655));
  jor  g00379(.dina(n655), .dinb(n622), .dout(n656));
  jxor g00380(.dina(n656), .dinb(n600), .dout(n657));
  jand g00381(.dina(n657), .dinb(n348), .dout(n658));
  jand g00382(.dina(n595), .dinb(b0 ), .dout(n659));
  jand g00383(.dina(n659), .dinb(n335), .dout(n660));
  jand g00384(.dina(n660), .dinb(n446), .dout(n661));
  jnot g00385(.din(n661), .dout(n662));
  jor  g00386(.dina(n662), .dinb(n621), .dout(n663));
  jand g00387(.dina(n663), .dinb(a59 ), .dout(n664));
  jand g00388(.dina(n602), .dinb(n448), .dout(n665));
  jand g00389(.dina(n665), .dinb(n445), .dout(n666));
  jnot g00390(.din(n666), .dout(n667));
  jor  g00391(.dina(n667), .dinb(n621), .dout(n668));
  jnot g00392(.din(n668), .dout(n669));
  jor  g00393(.dina(n669), .dinb(n664), .dout(n670));
  jand g00394(.dina(n670), .dinb(n258), .dout(n671));
  jnot g00395(.din(a58 ), .dout(n672));
  jand g00396(.dina(b0 ), .dinb(n672), .dout(n673));
  jnot g00397(.din(n673), .dout(n674));
  jxor g00398(.dina(n670), .dinb(n258), .dout(n675));
  jand g00399(.dina(n675), .dinb(n674), .dout(n676));
  jor  g00400(.dina(n676), .dinb(n671), .dout(n677));
  jxor g00401(.dina(n657), .dinb(n348), .dout(n678));
  jand g00402(.dina(n678), .dinb(n677), .dout(n679));
  jor  g00403(.dina(n679), .dinb(n658), .dout(n680));
  jxor g00404(.dina(n632), .dinb(n344), .dout(n681));
  jand g00405(.dina(n681), .dinb(n680), .dout(n682));
  jor  g00406(.dina(n682), .dinb(n654), .dout(n683));
  jxor g00407(.dina(n651), .dinb(b4 ), .dout(n684));
  jand g00408(.dina(n684), .dinb(n683), .dout(n685));
  jor  g00409(.dina(n685), .dinb(n18653), .dout(n686));
  jxor g00410(.dina(n636), .dinb(b5 ), .dout(n687));
  jand g00411(.dina(n687), .dinb(n686), .dout(n688));
  jand g00412(.dina(n688), .dinb(n641), .dout(n689));
  jor  g00413(.dina(n689), .dinb(n638), .dout(quotient58 ));
  jnot g00414(.din(quotient58 ), .dout(n691));
  jand g00415(.dina(n691), .dinb(n632), .dout(n692));
  jxor g00416(.dina(n681), .dinb(n680), .dout(n693));
  jand g00417(.dina(n693), .dinb(quotient58 ), .dout(n694));
  jor  g00418(.dina(n694), .dinb(n692), .dout(n695));
  jxor g00419(.dina(n687), .dinb(n686), .dout(n696));
  jor  g00420(.dina(n696), .dinb(n691), .dout(n697));
  jnot g00421(.din(n689), .dout(n698));
  jand g00422(.dina(n698), .dinb(n636), .dout(n699));
  jnot g00423(.din(n699), .dout(n700));
  jand g00424(.dina(n700), .dinb(n697), .dout(n701));
  jand g00425(.dina(n701), .dinb(n334), .dout(n702));
  jnot g00426(.din(n701), .dout(n703));
  jand g00427(.dina(n703), .dinb(b6 ), .dout(n704));
  jnot g00428(.din(n704), .dout(n705));
  jand g00429(.dina(n691), .dinb(n18652), .dout(n706));
  jxor g00430(.dina(n684), .dinb(n683), .dout(n707));
  jand g00431(.dina(n707), .dinb(quotient58 ), .dout(n708));
  jor  g00432(.dina(n708), .dinb(n706), .dout(n709));
  jand g00433(.dina(n709), .dinb(n338), .dout(n710));
  jand g00434(.dina(n695), .dinb(n337), .dout(n711));
  jand g00435(.dina(n691), .dinb(n657), .dout(n712));
  jxor g00436(.dina(n678), .dinb(n677), .dout(n713));
  jand g00437(.dina(n713), .dinb(quotient58 ), .dout(n714));
  jor  g00438(.dina(n714), .dinb(n712), .dout(n715));
  jand g00439(.dina(n715), .dinb(n344), .dout(n716));
  jnot g00440(.din(n670), .dout(n717));
  jor  g00441(.dina(quotient58 ), .dinb(n717), .dout(n718));
  jxor g00442(.dina(n675), .dinb(n674), .dout(n719));
  jnot g00443(.din(n719), .dout(n720));
  jor  g00444(.dina(n720), .dinb(n691), .dout(n721));
  jand g00445(.dina(n721), .dinb(n718), .dout(n722));
  jand g00446(.dina(quotient58 ), .dinb(b0 ), .dout(n725));
  jor  g00447(.dina(n725), .dinb(n672), .dout(n726));
  jand g00448(.dina(quotient58 ), .dinb(n673), .dout(n727));
  jnot g00449(.din(n727), .dout(n728));
  jand g00450(.dina(n728), .dinb(n726), .dout(n729));
  jnot g00451(.din(n729), .dout(n730));
  jand g00452(.dina(n730), .dinb(n258), .dout(n731));
  jnot g00453(.din(a57 ), .dout(n732));
  jand g00454(.dina(b0 ), .dinb(n732), .dout(n733));
  jnot g00455(.din(n733), .dout(n734));
  jxor g00456(.dina(n729), .dinb(b1 ), .dout(n735));
  jand g00457(.dina(n735), .dinb(n734), .dout(n736));
  jor  g00458(.dina(n736), .dinb(n731), .dout(n737));
  jxor g00459(.dina(n722), .dinb(b2 ), .dout(n738));
  jand g00460(.dina(n738), .dinb(n737), .dout(n739));
  jor  g00461(.dina(n739), .dinb(n18739), .dout(n740));
  jxor g00462(.dina(n715), .dinb(n344), .dout(n741));
  jand g00463(.dina(n741), .dinb(n740), .dout(n742));
  jor  g00464(.dina(n742), .dinb(n716), .dout(n743));
  jxor g00465(.dina(n695), .dinb(n337), .dout(n744));
  jand g00466(.dina(n744), .dinb(n743), .dout(n745));
  jor  g00467(.dina(n745), .dinb(n711), .dout(n746));
  jxor g00468(.dina(n709), .dinb(n338), .dout(n747));
  jand g00469(.dina(n747), .dinb(n746), .dout(n748));
  jor  g00470(.dina(n748), .dinb(n710), .dout(n749));
  jand g00471(.dina(n749), .dinb(n705), .dout(n750));
  jor  g00472(.dina(n750), .dinb(n702), .dout(n751));
  jand g00473(.dina(n751), .dinb(n555), .dout(quotient57 ));
  jnot g00474(.din(quotient57 ), .dout(n753));
  jand g00475(.dina(n753), .dinb(n695), .dout(n754));
  jxor g00476(.dina(n744), .dinb(n743), .dout(n755));
  jand g00477(.dina(n755), .dinb(quotient57 ), .dout(n756));
  jor  g00478(.dina(n756), .dinb(n754), .dout(n757));
  jand g00479(.dina(n753), .dinb(n701), .dout(n758));
  jand g00480(.dina(n702), .dinb(n555), .dout(n759));
  jand g00481(.dina(n759), .dinb(n749), .dout(n760));
  jor  g00482(.dina(n760), .dinb(n758), .dout(n761));
  jand g00483(.dina(n761), .dinb(n335), .dout(n762));
  jand g00484(.dina(n753), .dinb(n709), .dout(n763));
  jxor g00485(.dina(n747), .dinb(n746), .dout(n764));
  jand g00486(.dina(n764), .dinb(quotient57 ), .dout(n765));
  jor  g00487(.dina(n765), .dinb(n763), .dout(n766));
  jand g00488(.dina(n766), .dinb(n334), .dout(n767));
  jand g00489(.dina(n757), .dinb(n338), .dout(n768));
  jand g00490(.dina(n753), .dinb(n715), .dout(n769));
  jxor g00491(.dina(n741), .dinb(n740), .dout(n770));
  jand g00492(.dina(n770), .dinb(quotient57 ), .dout(n771));
  jor  g00493(.dina(n771), .dinb(n769), .dout(n772));
  jand g00494(.dina(n772), .dinb(n337), .dout(n773));
  jand g00495(.dina(n753), .dinb(n18738), .dout(n774));
  jxor g00496(.dina(n738), .dinb(n737), .dout(n775));
  jand g00497(.dina(n775), .dinb(quotient57 ), .dout(n776));
  jor  g00498(.dina(n776), .dinb(n774), .dout(n777));
  jand g00499(.dina(n777), .dinb(n344), .dout(n778));
  jand g00500(.dina(n753), .dinb(n730), .dout(n779));
  jxor g00501(.dina(n735), .dinb(n734), .dout(n780));
  jand g00502(.dina(n780), .dinb(quotient57 ), .dout(n781));
  jor  g00503(.dina(n781), .dinb(n779), .dout(n782));
  jand g00504(.dina(n782), .dinb(n348), .dout(n783));
  jand g00505(.dina(n751), .dinb(n660), .dout(n784));
  jor  g00506(.dina(n784), .dinb(n732), .dout(n785));
  jand g00507(.dina(n733), .dinb(n555), .dout(n786));
  jand g00508(.dina(n786), .dinb(n751), .dout(n787));
  jnot g00509(.din(n787), .dout(n788));
  jand g00510(.dina(n788), .dinb(n785), .dout(n789));
  jnot g00511(.din(n789), .dout(n790));
  jand g00512(.dina(n790), .dinb(n258), .dout(n791));
  jnot g00513(.din(a56 ), .dout(n792));
  jand g00514(.dina(b0 ), .dinb(n792), .dout(n793));
  jnot g00515(.din(n793), .dout(n794));
  jxor g00516(.dina(n789), .dinb(b1 ), .dout(n795));
  jand g00517(.dina(n795), .dinb(n794), .dout(n796));
  jor  g00518(.dina(n796), .dinb(n791), .dout(n797));
  jxor g00519(.dina(n782), .dinb(n348), .dout(n798));
  jand g00520(.dina(n798), .dinb(n797), .dout(n799));
  jor  g00521(.dina(n799), .dinb(n783), .dout(n800));
  jxor g00522(.dina(n777), .dinb(n344), .dout(n801));
  jand g00523(.dina(n801), .dinb(n800), .dout(n802));
  jor  g00524(.dina(n802), .dinb(n778), .dout(n803));
  jxor g00525(.dina(n772), .dinb(n337), .dout(n804));
  jand g00526(.dina(n804), .dinb(n803), .dout(n805));
  jor  g00527(.dina(n805), .dinb(n773), .dout(n806));
  jxor g00528(.dina(n757), .dinb(n338), .dout(n807));
  jand g00529(.dina(n807), .dinb(n806), .dout(n808));
  jor  g00530(.dina(n808), .dinb(n768), .dout(n809));
  jxor g00531(.dina(n766), .dinb(n334), .dout(n810));
  jand g00532(.dina(n810), .dinb(n809), .dout(n811));
  jor  g00533(.dina(n811), .dinb(n767), .dout(n812));
  jnot g00534(.din(n761), .dout(n813));
  jand g00535(.dina(n813), .dinb(b7 ), .dout(n814));
  jnot g00536(.din(n814), .dout(n815));
  jand g00537(.dina(n815), .dinb(n812), .dout(n816));
  jor  g00538(.dina(n816), .dinb(n762), .dout(n817));
  jand g00539(.dina(n817), .dinb(n595), .dout(quotient56 ));
  jnot g00540(.din(quotient56 ), .dout(n819));
  jand g00541(.dina(n819), .dinb(n757), .dout(n820));
  jxor g00542(.dina(n807), .dinb(n806), .dout(n821));
  jand g00543(.dina(n821), .dinb(quotient56 ), .dout(n822));
  jor  g00544(.dina(n822), .dinb(n820), .dout(n823));
  jand g00545(.dina(n819), .dinb(n761), .dout(n824));
  jand g00546(.dina(n762), .dinb(n595), .dout(n825));
  jand g00547(.dina(n825), .dinb(n812), .dout(n826));
  jor  g00548(.dina(n826), .dinb(n824), .dout(n827));
  jand g00549(.dina(n827), .dinb(n595), .dout(n828));
  jand g00550(.dina(n819), .dinb(n766), .dout(n829));
  jxor g00551(.dina(n810), .dinb(n809), .dout(n830));
  jand g00552(.dina(n830), .dinb(quotient56 ), .dout(n831));
  jor  g00553(.dina(n831), .dinb(n829), .dout(n832));
  jand g00554(.dina(n832), .dinb(n335), .dout(n833));
  jand g00555(.dina(n823), .dinb(n334), .dout(n834));
  jand g00556(.dina(n819), .dinb(n772), .dout(n835));
  jxor g00557(.dina(n804), .dinb(n803), .dout(n836));
  jand g00558(.dina(n836), .dinb(quotient56 ), .dout(n837));
  jor  g00559(.dina(n837), .dinb(n835), .dout(n838));
  jand g00560(.dina(n838), .dinb(n338), .dout(n839));
  jand g00561(.dina(n819), .dinb(n777), .dout(n840));
  jxor g00562(.dina(n801), .dinb(n800), .dout(n841));
  jand g00563(.dina(n841), .dinb(quotient56 ), .dout(n842));
  jor  g00564(.dina(n842), .dinb(n840), .dout(n843));
  jand g00565(.dina(n843), .dinb(n337), .dout(n844));
  jand g00566(.dina(n819), .dinb(n782), .dout(n845));
  jxor g00567(.dina(n798), .dinb(n797), .dout(n846));
  jand g00568(.dina(n846), .dinb(quotient56 ), .dout(n847));
  jor  g00569(.dina(n847), .dinb(n845), .dout(n848));
  jand g00570(.dina(n848), .dinb(n344), .dout(n849));
  jand g00571(.dina(n819), .dinb(n790), .dout(n850));
  jxor g00572(.dina(n795), .dinb(n794), .dout(n851));
  jand g00573(.dina(n851), .dinb(quotient56 ), .dout(n852));
  jor  g00574(.dina(n852), .dinb(n850), .dout(n853));
  jand g00575(.dina(n853), .dinb(n348), .dout(n854));
  jand g00576(.dina(n441), .dinb(b0 ), .dout(n856));
  jand g00577(.dina(n856), .dinb(n327), .dout(n857));
  jand g00578(.dina(n857), .dinb(n989), .dout(n858));
  jand g00579(.dina(n858), .dinb(n817), .dout(n859));
  jor  g00580(.dina(n859), .dinb(n792), .dout(n860));
  jand g00581(.dina(n659), .dinb(n792), .dout(n861));
  jand g00582(.dina(n861), .dinb(n817), .dout(n862));
  jnot g00583(.din(n862), .dout(n863));
  jand g00584(.dina(n863), .dinb(n860), .dout(n864));
  jor  g00585(.dina(n864), .dinb(b1 ), .dout(n865));
  jnot g00586(.din(n865), .dout(n866));
  jnot g00587(.din(a55 ), .dout(n867));
  jand g00588(.dina(b0 ), .dinb(n867), .dout(n868));
  jnot g00589(.din(n868), .dout(n869));
  jxor g00590(.dina(n864), .dinb(b1 ), .dout(n870));
  jand g00591(.dina(n870), .dinb(n869), .dout(n871));
  jor  g00592(.dina(n871), .dinb(n866), .dout(n872));
  jxor g00593(.dina(n853), .dinb(n348), .dout(n873));
  jand g00594(.dina(n873), .dinb(n872), .dout(n874));
  jor  g00595(.dina(n874), .dinb(n854), .dout(n875));
  jxor g00596(.dina(n848), .dinb(n344), .dout(n876));
  jand g00597(.dina(n876), .dinb(n875), .dout(n877));
  jor  g00598(.dina(n877), .dinb(n849), .dout(n878));
  jxor g00599(.dina(n843), .dinb(n337), .dout(n879));
  jand g00600(.dina(n879), .dinb(n878), .dout(n880));
  jor  g00601(.dina(n880), .dinb(n844), .dout(n881));
  jxor g00602(.dina(n838), .dinb(n338), .dout(n882));
  jand g00603(.dina(n882), .dinb(n881), .dout(n883));
  jor  g00604(.dina(n883), .dinb(n839), .dout(n884));
  jxor g00605(.dina(n823), .dinb(n334), .dout(n885));
  jand g00606(.dina(n885), .dinb(n884), .dout(n886));
  jor  g00607(.dina(n886), .dinb(n834), .dout(n887));
  jxor g00608(.dina(n832), .dinb(n335), .dout(n888));
  jand g00609(.dina(n888), .dinb(n887), .dout(n889));
  jor  g00610(.dina(n889), .dinb(n833), .dout(n890));
  jxor g00611(.dina(n827), .dinb(b8 ), .dout(n891));
  jnot g00612(.din(n891), .dout(n892));
  jand g00613(.dina(n892), .dinb(n890), .dout(n893));
  jand g00614(.dina(n893), .dinb(n445), .dout(n894));
  jor  g00615(.dina(n894), .dinb(n828), .dout(quotient55 ));
  jnot g00616(.din(quotient55 ), .dout(n896));
  jand g00617(.dina(n896), .dinb(n823), .dout(n897));
  jxor g00618(.dina(n885), .dinb(n884), .dout(n898));
  jand g00619(.dina(n898), .dinb(quotient55 ), .dout(n899));
  jor  g00620(.dina(n899), .dinb(n897), .dout(n900));
  jxor g00621(.dina(n892), .dinb(n890), .dout(n901));
  jor  g00622(.dina(n901), .dinb(n896), .dout(n902));
  jor  g00623(.dina(n894), .dinb(n827), .dout(n903));
  jand g00624(.dina(n903), .dinb(n902), .dout(n904));
  jnot g00625(.din(n904), .dout(n905));
  jand g00626(.dina(n905), .dinb(b9 ), .dout(n906));
  jnot g00627(.din(n906), .dout(n907));
  jand g00628(.dina(n904), .dinb(n324), .dout(n908));
  jand g00629(.dina(n896), .dinb(n832), .dout(n909));
  jxor g00630(.dina(n888), .dinb(n887), .dout(n910));
  jand g00631(.dina(n910), .dinb(quotient55 ), .dout(n911));
  jor  g00632(.dina(n911), .dinb(n909), .dout(n912));
  jand g00633(.dina(n912), .dinb(n323), .dout(n913));
  jand g00634(.dina(n900), .dinb(n335), .dout(n914));
  jand g00635(.dina(n896), .dinb(n838), .dout(n915));
  jxor g00636(.dina(n882), .dinb(n881), .dout(n916));
  jand g00637(.dina(n916), .dinb(quotient55 ), .dout(n917));
  jor  g00638(.dina(n917), .dinb(n915), .dout(n918));
  jand g00639(.dina(n918), .dinb(n334), .dout(n919));
  jand g00640(.dina(n896), .dinb(n843), .dout(n920));
  jxor g00641(.dina(n879), .dinb(n878), .dout(n921));
  jand g00642(.dina(n921), .dinb(quotient55 ), .dout(n922));
  jor  g00643(.dina(n922), .dinb(n920), .dout(n923));
  jand g00644(.dina(n923), .dinb(n338), .dout(n924));
  jand g00645(.dina(n896), .dinb(n848), .dout(n925));
  jxor g00646(.dina(n876), .dinb(n875), .dout(n926));
  jand g00647(.dina(n926), .dinb(quotient55 ), .dout(n927));
  jor  g00648(.dina(n927), .dinb(n925), .dout(n928));
  jand g00649(.dina(n928), .dinb(n337), .dout(n929));
  jand g00650(.dina(n896), .dinb(n853), .dout(n930));
  jxor g00651(.dina(n873), .dinb(n872), .dout(n931));
  jand g00652(.dina(n931), .dinb(quotient55 ), .dout(n932));
  jor  g00653(.dina(n932), .dinb(n930), .dout(n933));
  jand g00654(.dina(n933), .dinb(n344), .dout(n934));
  jor  g00655(.dina(quotient55 ), .dinb(n864), .dout(n935));
  jxor g00656(.dina(n870), .dinb(n869), .dout(n936));
  jnot g00657(.din(n936), .dout(n937));
  jor  g00658(.dina(n937), .dinb(n896), .dout(n938));
  jand g00659(.dina(n938), .dinb(n935), .dout(n939));
  jand g00660(.dina(quotient55 ), .dinb(b0 ), .dout(n942));
  jor  g00661(.dina(n942), .dinb(n867), .dout(n943));
  jand g00662(.dina(quotient55 ), .dinb(n868), .dout(n944));
  jnot g00663(.din(n944), .dout(n945));
  jand g00664(.dina(n945), .dinb(n943), .dout(n946));
  jnot g00665(.din(n946), .dout(n947));
  jand g00666(.dina(n947), .dinb(n258), .dout(n948));
  jnot g00667(.din(a54 ), .dout(n949));
  jand g00668(.dina(b0 ), .dinb(n949), .dout(n950));
  jnot g00669(.din(n950), .dout(n951));
  jxor g00670(.dina(n946), .dinb(b1 ), .dout(n952));
  jand g00671(.dina(n952), .dinb(n951), .dout(n953));
  jor  g00672(.dina(n953), .dinb(n948), .dout(n954));
  jxor g00673(.dina(n939), .dinb(b2 ), .dout(n955));
  jand g00674(.dina(n955), .dinb(n954), .dout(n956));
  jor  g00675(.dina(n956), .dinb(n19041), .dout(n957));
  jxor g00676(.dina(n933), .dinb(n344), .dout(n958));
  jand g00677(.dina(n958), .dinb(n957), .dout(n959));
  jor  g00678(.dina(n959), .dinb(n934), .dout(n960));
  jxor g00679(.dina(n928), .dinb(n337), .dout(n961));
  jand g00680(.dina(n961), .dinb(n960), .dout(n962));
  jor  g00681(.dina(n962), .dinb(n929), .dout(n963));
  jxor g00682(.dina(n923), .dinb(n338), .dout(n964));
  jand g00683(.dina(n964), .dinb(n963), .dout(n965));
  jor  g00684(.dina(n965), .dinb(n924), .dout(n966));
  jxor g00685(.dina(n918), .dinb(n334), .dout(n967));
  jand g00686(.dina(n967), .dinb(n966), .dout(n968));
  jor  g00687(.dina(n968), .dinb(n919), .dout(n969));
  jxor g00688(.dina(n900), .dinb(n335), .dout(n970));
  jand g00689(.dina(n970), .dinb(n969), .dout(n971));
  jor  g00690(.dina(n971), .dinb(n914), .dout(n972));
  jxor g00691(.dina(n912), .dinb(n323), .dout(n973));
  jand g00692(.dina(n973), .dinb(n972), .dout(n974));
  jor  g00693(.dina(n974), .dinb(n913), .dout(n975));
  jor  g00694(.dina(n975), .dinb(n908), .dout(n976));
  jand g00695(.dina(n976), .dinb(n907), .dout(n977));
  jand g00696(.dina(n594), .dinb(n439), .dout(n978));
  jnot g00697(.din(n331), .dout(n979));
  jand g00698(.dina(n979), .dinb(n325), .dout(n980));
  jand g00699(.dina(n980), .dinb(n978), .dout(n981));
  jand g00700(.dina(n981), .dinb(n977), .dout(quotient54 ));
  jnot g00701(.din(quotient54 ), .dout(n983));
  jand g00702(.dina(n983), .dinb(n900), .dout(n984));
  jxor g00703(.dina(n970), .dinb(n969), .dout(n985));
  jand g00704(.dina(n985), .dinb(quotient54 ), .dout(n986));
  jor  g00705(.dina(n986), .dinb(n984), .dout(n987));
  jand g00706(.dina(n431), .dinb(n403), .dout(n988));
  jand g00707(.dina(n988), .dinb(n438), .dout(n989));
  jand g00708(.dina(n989), .dinb(n441), .dout(n990));
  jnot g00709(.din(n990), .dout(n991));
  jand g00710(.dina(n983), .dinb(n904), .dout(n992));
  jand g00711(.dina(n981), .dinb(n908), .dout(n993));
  jand g00712(.dina(n993), .dinb(n975), .dout(n994));
  jor  g00713(.dina(n994), .dinb(n992), .dout(n995));
  jand g00714(.dina(n995), .dinb(n325), .dout(n996));
  jnot g00715(.din(n996), .dout(n997));
  jand g00716(.dina(n983), .dinb(n912), .dout(n998));
  jxor g00717(.dina(n973), .dinb(n972), .dout(n999));
  jand g00718(.dina(n999), .dinb(quotient54 ), .dout(n1000));
  jor  g00719(.dina(n1000), .dinb(n998), .dout(n1001));
  jand g00720(.dina(n1001), .dinb(n324), .dout(n1002));
  jnot g00721(.din(n1002), .dout(n1003));
  jand g00722(.dina(n987), .dinb(n323), .dout(n1004));
  jnot g00723(.din(n1004), .dout(n1005));
  jand g00724(.dina(n983), .dinb(n918), .dout(n1006));
  jxor g00725(.dina(n967), .dinb(n966), .dout(n1007));
  jand g00726(.dina(n1007), .dinb(quotient54 ), .dout(n1008));
  jor  g00727(.dina(n1008), .dinb(n1006), .dout(n1009));
  jand g00728(.dina(n1009), .dinb(n335), .dout(n1010));
  jnot g00729(.din(n1010), .dout(n1011));
  jand g00730(.dina(n983), .dinb(n923), .dout(n1012));
  jxor g00731(.dina(n964), .dinb(n963), .dout(n1013));
  jand g00732(.dina(n1013), .dinb(quotient54 ), .dout(n1014));
  jor  g00733(.dina(n1014), .dinb(n1012), .dout(n1015));
  jand g00734(.dina(n1015), .dinb(n334), .dout(n1016));
  jnot g00735(.din(n1016), .dout(n1017));
  jand g00736(.dina(n983), .dinb(n928), .dout(n1018));
  jxor g00737(.dina(n961), .dinb(n960), .dout(n1019));
  jand g00738(.dina(n1019), .dinb(quotient54 ), .dout(n1020));
  jor  g00739(.dina(n1020), .dinb(n1018), .dout(n1021));
  jand g00740(.dina(n1021), .dinb(n338), .dout(n1022));
  jnot g00741(.din(n1022), .dout(n1023));
  jand g00742(.dina(n983), .dinb(n933), .dout(n1024));
  jxor g00743(.dina(n958), .dinb(n957), .dout(n1025));
  jand g00744(.dina(n1025), .dinb(quotient54 ), .dout(n1026));
  jor  g00745(.dina(n1026), .dinb(n1024), .dout(n1027));
  jand g00746(.dina(n1027), .dinb(n337), .dout(n1028));
  jnot g00747(.din(n1028), .dout(n1029));
  jand g00748(.dina(n983), .dinb(n19040), .dout(n1030));
  jxor g00749(.dina(n955), .dinb(n954), .dout(n1031));
  jand g00750(.dina(n1031), .dinb(quotient54 ), .dout(n1032));
  jor  g00751(.dina(n1032), .dinb(n1030), .dout(n1033));
  jand g00752(.dina(n1033), .dinb(n344), .dout(n1034));
  jnot g00753(.din(n1034), .dout(n1035));
  jand g00754(.dina(n983), .dinb(n947), .dout(n1036));
  jxor g00755(.dina(n952), .dinb(n951), .dout(n1037));
  jand g00756(.dina(n1037), .dinb(quotient54 ), .dout(n1038));
  jor  g00757(.dina(n1038), .dinb(n1036), .dout(n1039));
  jand g00758(.dina(n1039), .dinb(n348), .dout(n1040));
  jnot g00759(.din(n1040), .dout(n1041));
  jand g00760(.dina(n325), .dinb(b0 ), .dout(n1042));
  jand g00761(.dina(n1042), .dinb(n990), .dout(n1043));
  jand g00762(.dina(n1043), .dinb(n977), .dout(n1044));
  jor  g00763(.dina(n1044), .dinb(n949), .dout(n1045));
  jand g00764(.dina(n981), .dinb(n950), .dout(n1046));
  jand g00765(.dina(n1046), .dinb(n977), .dout(n1047));
  jnot g00766(.din(n1047), .dout(n1048));
  jand g00767(.dina(n1048), .dinb(n1045), .dout(n1049));
  jor  g00768(.dina(n1049), .dinb(b1 ), .dout(n1050));
  jnot g00769(.din(a53 ), .dout(n1051));
  jand g00770(.dina(b0 ), .dinb(n1051), .dout(n1052));
  jxor g00771(.dina(n1049), .dinb(n258), .dout(n1053));
  jor  g00772(.dina(n1053), .dinb(n1052), .dout(n1054));
  jand g00773(.dina(n1054), .dinb(n1050), .dout(n1055));
  jxor g00774(.dina(n1039), .dinb(n348), .dout(n1056));
  jnot g00775(.din(n1056), .dout(n1057));
  jor  g00776(.dina(n1057), .dinb(n1055), .dout(n1058));
  jand g00777(.dina(n1058), .dinb(n1041), .dout(n1059));
  jxor g00778(.dina(n1033), .dinb(n344), .dout(n1060));
  jnot g00779(.din(n1060), .dout(n1061));
  jor  g00780(.dina(n1061), .dinb(n1059), .dout(n1062));
  jand g00781(.dina(n1062), .dinb(n1035), .dout(n1063));
  jxor g00782(.dina(n1027), .dinb(n337), .dout(n1064));
  jnot g00783(.din(n1064), .dout(n1065));
  jor  g00784(.dina(n1065), .dinb(n1063), .dout(n1066));
  jand g00785(.dina(n1066), .dinb(n1029), .dout(n1067));
  jxor g00786(.dina(n1021), .dinb(n338), .dout(n1068));
  jnot g00787(.din(n1068), .dout(n1069));
  jor  g00788(.dina(n1069), .dinb(n1067), .dout(n1070));
  jand g00789(.dina(n1070), .dinb(n1023), .dout(n1071));
  jxor g00790(.dina(n1015), .dinb(n334), .dout(n1072));
  jnot g00791(.din(n1072), .dout(n1073));
  jor  g00792(.dina(n1073), .dinb(n1071), .dout(n1074));
  jand g00793(.dina(n1074), .dinb(n1017), .dout(n1075));
  jxor g00794(.dina(n1009), .dinb(n335), .dout(n1076));
  jnot g00795(.din(n1076), .dout(n1077));
  jor  g00796(.dina(n1077), .dinb(n1075), .dout(n1078));
  jand g00797(.dina(n1078), .dinb(n1011), .dout(n1079));
  jxor g00798(.dina(n987), .dinb(n323), .dout(n1080));
  jnot g00799(.din(n1080), .dout(n1081));
  jor  g00800(.dina(n1081), .dinb(n1079), .dout(n1082));
  jand g00801(.dina(n1082), .dinb(n1005), .dout(n1083));
  jxor g00802(.dina(n1001), .dinb(n324), .dout(n1084));
  jnot g00803(.din(n1084), .dout(n1085));
  jor  g00804(.dina(n1085), .dinb(n1083), .dout(n1086));
  jand g00805(.dina(n1086), .dinb(n1003), .dout(n1087));
  jnot g00806(.din(n995), .dout(n1088));
  jand g00807(.dina(n1088), .dinb(b10 ), .dout(n1089));
  jor  g00808(.dina(n1089), .dinb(n1087), .dout(n1090));
  jand g00809(.dina(n1090), .dinb(n997), .dout(n1091));
  jor  g00810(.dina(n1091), .dinb(n991), .dout(n1092));
  jand g00811(.dina(n1092), .dinb(n987), .dout(n1093));
  jnot g00812(.din(n1092), .dout(quotient53 ));
  jnot g00813(.din(n1050), .dout(n1095));
  jnot g00814(.din(n1052), .dout(n1096));
  jxor g00815(.dina(n1049), .dinb(b1 ), .dout(n1097));
  jand g00816(.dina(n1097), .dinb(n1096), .dout(n1098));
  jor  g00817(.dina(n1098), .dinb(n1095), .dout(n1099));
  jand g00818(.dina(n1056), .dinb(n1099), .dout(n1100));
  jor  g00819(.dina(n1100), .dinb(n1040), .dout(n1101));
  jand g00820(.dina(n1060), .dinb(n1101), .dout(n1102));
  jor  g00821(.dina(n1102), .dinb(n1034), .dout(n1103));
  jand g00822(.dina(n1064), .dinb(n1103), .dout(n1104));
  jor  g00823(.dina(n1104), .dinb(n1028), .dout(n1105));
  jand g00824(.dina(n1068), .dinb(n1105), .dout(n1106));
  jor  g00825(.dina(n1106), .dinb(n1022), .dout(n1107));
  jand g00826(.dina(n1072), .dinb(n1107), .dout(n1108));
  jor  g00827(.dina(n1108), .dinb(n1016), .dout(n1109));
  jand g00828(.dina(n1076), .dinb(n1109), .dout(n1110));
  jor  g00829(.dina(n1110), .dinb(n1010), .dout(n1111));
  jxor g00830(.dina(n1080), .dinb(n1111), .dout(n1112));
  jand g00831(.dina(n1112), .dinb(quotient53 ), .dout(n1113));
  jor  g00832(.dina(n1113), .dinb(n1093), .dout(n1114));
  jand g00833(.dina(n1092), .dinb(n995), .dout(n1115));
  jand g00834(.dina(n1080), .dinb(n1111), .dout(n1116));
  jor  g00835(.dina(n1116), .dinb(n1004), .dout(n1117));
  jand g00836(.dina(n1084), .dinb(n1117), .dout(n1118));
  jor  g00837(.dina(n1118), .dinb(n1002), .dout(n1119));
  jand g00838(.dina(n996), .dinb(n990), .dout(n1120));
  jand g00839(.dina(n1120), .dinb(n1119), .dout(n1121));
  jor  g00840(.dina(n1121), .dinb(n1115), .dout(n1122));
  jand g00841(.dina(n1122), .dinb(n990), .dout(n1123));
  jand g00842(.dina(n1092), .dinb(n1001), .dout(n1124));
  jxor g00843(.dina(n1084), .dinb(n1117), .dout(n1125));
  jand g00844(.dina(n1125), .dinb(quotient53 ), .dout(n1126));
  jor  g00845(.dina(n1126), .dinb(n1124), .dout(n1127));
  jand g00846(.dina(n1127), .dinb(n325), .dout(n1128));
  jand g00847(.dina(n1114), .dinb(n324), .dout(n1129));
  jand g00848(.dina(n1092), .dinb(n1009), .dout(n1130));
  jxor g00849(.dina(n1076), .dinb(n1109), .dout(n1131));
  jand g00850(.dina(n1131), .dinb(quotient53 ), .dout(n1132));
  jor  g00851(.dina(n1132), .dinb(n1130), .dout(n1133));
  jand g00852(.dina(n1133), .dinb(n323), .dout(n1134));
  jand g00853(.dina(n1092), .dinb(n1015), .dout(n1135));
  jxor g00854(.dina(n1072), .dinb(n1107), .dout(n1136));
  jand g00855(.dina(n1136), .dinb(quotient53 ), .dout(n1137));
  jor  g00856(.dina(n1137), .dinb(n1135), .dout(n1138));
  jand g00857(.dina(n1138), .dinb(n335), .dout(n1139));
  jand g00858(.dina(n1092), .dinb(n1021), .dout(n1140));
  jxor g00859(.dina(n1068), .dinb(n1105), .dout(n1141));
  jand g00860(.dina(n1141), .dinb(quotient53 ), .dout(n1142));
  jor  g00861(.dina(n1142), .dinb(n1140), .dout(n1143));
  jand g00862(.dina(n1143), .dinb(n334), .dout(n1144));
  jand g00863(.dina(n1092), .dinb(n1027), .dout(n1145));
  jxor g00864(.dina(n1064), .dinb(n1103), .dout(n1146));
  jand g00865(.dina(n1146), .dinb(quotient53 ), .dout(n1147));
  jor  g00866(.dina(n1147), .dinb(n1145), .dout(n1148));
  jand g00867(.dina(n1148), .dinb(n338), .dout(n1149));
  jand g00868(.dina(n1092), .dinb(n1033), .dout(n1150));
  jxor g00869(.dina(n1060), .dinb(n1101), .dout(n1151));
  jand g00870(.dina(n1151), .dinb(quotient53 ), .dout(n1152));
  jor  g00871(.dina(n1152), .dinb(n1150), .dout(n1153));
  jand g00872(.dina(n1153), .dinb(n337), .dout(n1154));
  jand g00873(.dina(n1092), .dinb(n1039), .dout(n1155));
  jxor g00874(.dina(n1056), .dinb(n1099), .dout(n1156));
  jand g00875(.dina(n1156), .dinb(quotient53 ), .dout(n1157));
  jor  g00876(.dina(n1157), .dinb(n1155), .dout(n1158));
  jand g00877(.dina(n1158), .dinb(n344), .dout(n1159));
  jxor g00878(.dina(n1097), .dinb(n1096), .dout(n1161));
  jand g00879(.dina(n1161), .dinb(quotient53 ), .dout(n1162));
  jnot g00880(.din(n1089), .dout(n1167));
  jand g00881(.dina(n1167), .dinb(n1119), .dout(n1168));
  jor  g00882(.dina(n1168), .dinb(n996), .dout(n1169));
  jand g00883(.dina(n979), .dinb(b0 ), .dout(n1170));
  jand g00884(.dina(n1170), .dinb(n978), .dout(n1171));
  jand g00885(.dina(n1171), .dinb(n1169), .dout(n1172));
  jor  g00886(.dina(n1172), .dinb(n1051), .dout(n1173));
  jor  g00887(.dina(n1092), .dinb(n1096), .dout(n1174));
  jand g00888(.dina(n1174), .dinb(n1173), .dout(n1175));
  jor  g00889(.dina(n1175), .dinb(b1 ), .dout(n1176));
  jnot g00890(.din(n1176), .dout(n1177));
  jnot g00891(.din(a52 ), .dout(n1178));
  jand g00892(.dina(b0 ), .dinb(n1178), .dout(n1179));
  jnot g00893(.din(n1179), .dout(n1180));
  jxor g00894(.dina(n1175), .dinb(b1 ), .dout(n1181));
  jand g00895(.dina(n1181), .dinb(n1180), .dout(n1182));
  jor  g00896(.dina(n1182), .dinb(n1177), .dout(n1183));
  jand g00897(.dina(n19327), .dinb(n1183), .dout(n1185));
  jor  g00898(.dina(n1185), .dinb(n19311), .dout(n1186));
  jxor g00899(.dina(n1158), .dinb(n344), .dout(n1187));
  jand g00900(.dina(n1187), .dinb(n1186), .dout(n1188));
  jor  g00901(.dina(n1188), .dinb(n1159), .dout(n1189));
  jxor g00902(.dina(n1153), .dinb(n337), .dout(n1190));
  jand g00903(.dina(n1190), .dinb(n1189), .dout(n1191));
  jor  g00904(.dina(n1191), .dinb(n1154), .dout(n1192));
  jxor g00905(.dina(n1148), .dinb(n338), .dout(n1193));
  jand g00906(.dina(n1193), .dinb(n1192), .dout(n1194));
  jor  g00907(.dina(n1194), .dinb(n1149), .dout(n1195));
  jxor g00908(.dina(n1143), .dinb(n334), .dout(n1196));
  jand g00909(.dina(n1196), .dinb(n1195), .dout(n1197));
  jor  g00910(.dina(n1197), .dinb(n1144), .dout(n1198));
  jxor g00911(.dina(n1138), .dinb(n335), .dout(n1199));
  jand g00912(.dina(n1199), .dinb(n1198), .dout(n1200));
  jor  g00913(.dina(n1200), .dinb(n1139), .dout(n1201));
  jxor g00914(.dina(n1133), .dinb(n323), .dout(n1202));
  jand g00915(.dina(n1202), .dinb(n1201), .dout(n1203));
  jor  g00916(.dina(n1203), .dinb(n1134), .dout(n1204));
  jxor g00917(.dina(n1114), .dinb(n324), .dout(n1205));
  jand g00918(.dina(n1205), .dinb(n1204), .dout(n1206));
  jor  g00919(.dina(n1206), .dinb(n1129), .dout(n1207));
  jxor g00920(.dina(n1127), .dinb(n325), .dout(n1208));
  jand g00921(.dina(n1208), .dinb(n1207), .dout(n1209));
  jor  g00922(.dina(n1209), .dinb(n1128), .dout(n1210));
  jxor g00923(.dina(n1122), .dinb(b11 ), .dout(n1211));
  jnot g00924(.din(n1211), .dout(n1212));
  jand g00925(.dina(n1212), .dinb(n1210), .dout(n1213));
  jand g00926(.dina(n979), .dinb(n594), .dout(n1214));
  jand g00927(.dina(n1214), .dinb(n1213), .dout(n1215));
  jor  g00928(.dina(n1215), .dinb(n1123), .dout(quotient52 ));
  jnot g00929(.din(quotient52 ), .dout(n1217));
  jand g00930(.dina(n1217), .dinb(n1114), .dout(n1218));
  jxor g00931(.dina(n1205), .dinb(n1204), .dout(n1219));
  jand g00932(.dina(n1219), .dinb(quotient52 ), .dout(n1220));
  jor  g00933(.dina(n1220), .dinb(n1218), .dout(n1221));
  jxor g00934(.dina(n1212), .dinb(n1210), .dout(n1222));
  jor  g00935(.dina(n1222), .dinb(n1217), .dout(n1223));
  jor  g00936(.dina(n1215), .dinb(n1122), .dout(n1224));
  jand g00937(.dina(n1224), .dinb(n1223), .dout(n1225));
  jnot g00938(.din(n1225), .dout(n1226));
  jand g00939(.dina(n1226), .dinb(b12 ), .dout(n1227));
  jnot g00940(.din(n1227), .dout(n1228));
  jand g00941(.dina(n1225), .dinb(n440), .dout(n1229));
  jand g00942(.dina(n1217), .dinb(n1127), .dout(n1230));
  jxor g00943(.dina(n1208), .dinb(n1207), .dout(n1231));
  jand g00944(.dina(n1231), .dinb(quotient52 ), .dout(n1232));
  jor  g00945(.dina(n1232), .dinb(n1230), .dout(n1233));
  jand g00946(.dina(n1233), .dinb(n439), .dout(n1234));
  jand g00947(.dina(n1221), .dinb(n325), .dout(n1235));
  jand g00948(.dina(n1217), .dinb(n1133), .dout(n1236));
  jxor g00949(.dina(n1202), .dinb(n1201), .dout(n1237));
  jand g00950(.dina(n1237), .dinb(quotient52 ), .dout(n1238));
  jor  g00951(.dina(n1238), .dinb(n1236), .dout(n1239));
  jand g00952(.dina(n1239), .dinb(n324), .dout(n1240));
  jand g00953(.dina(n1217), .dinb(n1138), .dout(n1241));
  jxor g00954(.dina(n1199), .dinb(n1198), .dout(n1242));
  jand g00955(.dina(n1242), .dinb(quotient52 ), .dout(n1243));
  jor  g00956(.dina(n1243), .dinb(n1241), .dout(n1244));
  jand g00957(.dina(n1244), .dinb(n323), .dout(n1245));
  jand g00958(.dina(n1217), .dinb(n1143), .dout(n1246));
  jxor g00959(.dina(n1196), .dinb(n1195), .dout(n1247));
  jand g00960(.dina(n1247), .dinb(quotient52 ), .dout(n1248));
  jor  g00961(.dina(n1248), .dinb(n1246), .dout(n1249));
  jand g00962(.dina(n1249), .dinb(n335), .dout(n1250));
  jand g00963(.dina(n1217), .dinb(n1148), .dout(n1251));
  jxor g00964(.dina(n1193), .dinb(n1192), .dout(n1252));
  jand g00965(.dina(n1252), .dinb(quotient52 ), .dout(n1253));
  jor  g00966(.dina(n1253), .dinb(n1251), .dout(n1254));
  jand g00967(.dina(n1254), .dinb(n334), .dout(n1255));
  jand g00968(.dina(n1217), .dinb(n1153), .dout(n1256));
  jxor g00969(.dina(n1190), .dinb(n1189), .dout(n1257));
  jand g00970(.dina(n1257), .dinb(quotient52 ), .dout(n1258));
  jor  g00971(.dina(n1258), .dinb(n1256), .dout(n1259));
  jand g00972(.dina(n1259), .dinb(n338), .dout(n1260));
  jand g00973(.dina(n1217), .dinb(n1158), .dout(n1261));
  jxor g00974(.dina(n1187), .dinb(n1186), .dout(n1262));
  jand g00975(.dina(n1262), .dinb(quotient52 ), .dout(n1263));
  jor  g00976(.dina(n1263), .dinb(n1261), .dout(n1264));
  jand g00977(.dina(n1264), .dinb(n337), .dout(n1265));
  jand g00978(.dina(n1217), .dinb(n19310), .dout(n1266));
  jxor g00979(.dina(n19327), .dinb(n1183), .dout(n1267));
  jand g00980(.dina(n1267), .dinb(quotient52 ), .dout(n1268));
  jor  g00981(.dina(n1268), .dinb(n1266), .dout(n1269));
  jand g00982(.dina(n1269), .dinb(n344), .dout(n1270));
  jor  g00983(.dina(quotient52 ), .dinb(n1175), .dout(n1271));
  jxor g00984(.dina(n1181), .dinb(n1180), .dout(n1272));
  jnot g00985(.din(n1272), .dout(n1273));
  jor  g00986(.dina(n1273), .dinb(n1217), .dout(n1274));
  jand g00987(.dina(n1274), .dinb(n1271), .dout(n1275));
  jand g00988(.dina(quotient52 ), .dinb(b0 ), .dout(n1278));
  jor  g00989(.dina(n1278), .dinb(n1178), .dout(n1279));
  jand g00990(.dina(quotient52 ), .dinb(n1179), .dout(n1280));
  jnot g00991(.din(n1280), .dout(n1281));
  jand g00992(.dina(n1281), .dinb(n1279), .dout(n1282));
  jnot g00993(.din(n1282), .dout(n1283));
  jand g00994(.dina(n1283), .dinb(n258), .dout(n1284));
  jnot g00995(.din(a51 ), .dout(n1285));
  jand g00996(.dina(b0 ), .dinb(n1285), .dout(n1286));
  jnot g00997(.din(n1286), .dout(n1287));
  jxor g00998(.dina(n1282), .dinb(b1 ), .dout(n1288));
  jand g00999(.dina(n1288), .dinb(n1287), .dout(n1289));
  jor  g01000(.dina(n1289), .dinb(n1284), .dout(n1290));
  jxor g01001(.dina(n1275), .dinb(b2 ), .dout(n1291));
  jand g01002(.dina(n1291), .dinb(n1290), .dout(n1292));
  jor  g01003(.dina(n1292), .dinb(n19449), .dout(n1293));
  jxor g01004(.dina(n1269), .dinb(n344), .dout(n1294));
  jand g01005(.dina(n1294), .dinb(n1293), .dout(n1295));
  jor  g01006(.dina(n1295), .dinb(n1270), .dout(n1296));
  jxor g01007(.dina(n1264), .dinb(n337), .dout(n1297));
  jand g01008(.dina(n1297), .dinb(n1296), .dout(n1298));
  jor  g01009(.dina(n1298), .dinb(n1265), .dout(n1299));
  jxor g01010(.dina(n1259), .dinb(n338), .dout(n1300));
  jand g01011(.dina(n1300), .dinb(n1299), .dout(n1301));
  jor  g01012(.dina(n1301), .dinb(n1260), .dout(n1302));
  jxor g01013(.dina(n1254), .dinb(n334), .dout(n1303));
  jand g01014(.dina(n1303), .dinb(n1302), .dout(n1304));
  jor  g01015(.dina(n1304), .dinb(n1255), .dout(n1305));
  jxor g01016(.dina(n1249), .dinb(n335), .dout(n1306));
  jand g01017(.dina(n1306), .dinb(n1305), .dout(n1307));
  jor  g01018(.dina(n1307), .dinb(n1250), .dout(n1308));
  jxor g01019(.dina(n1244), .dinb(n323), .dout(n1309));
  jand g01020(.dina(n1309), .dinb(n1308), .dout(n1310));
  jor  g01021(.dina(n1310), .dinb(n1245), .dout(n1311));
  jxor g01022(.dina(n1239), .dinb(n324), .dout(n1312));
  jand g01023(.dina(n1312), .dinb(n1311), .dout(n1313));
  jor  g01024(.dina(n1313), .dinb(n1240), .dout(n1314));
  jxor g01025(.dina(n1221), .dinb(n325), .dout(n1315));
  jand g01026(.dina(n1315), .dinb(n1314), .dout(n1316));
  jor  g01027(.dina(n1316), .dinb(n1235), .dout(n1317));
  jxor g01028(.dina(n1233), .dinb(n439), .dout(n1318));
  jand g01029(.dina(n1318), .dinb(n1317), .dout(n1319));
  jor  g01030(.dina(n1319), .dinb(n1234), .dout(n1320));
  jor  g01031(.dina(n1320), .dinb(n1229), .dout(n1321));
  jand g01032(.dina(n1321), .dinb(n1228), .dout(n1322));
  jand g01033(.dina(n1322), .dinb(n989), .dout(quotient51 ));
  jnot g01034(.din(quotient51 ), .dout(n1324));
  jand g01035(.dina(n1324), .dinb(n1221), .dout(n1325));
  jxor g01036(.dina(n1315), .dinb(n1314), .dout(n1326));
  jand g01037(.dina(n1326), .dinb(quotient51 ), .dout(n1327));
  jor  g01038(.dina(n1327), .dinb(n1325), .dout(n1328));
  jnot g01039(.din(n329), .dout(n1329));
  jand g01040(.dina(n1329), .dinb(n594), .dout(n1330));
  jnot g01041(.din(n1330), .dout(n1331));
  jand g01042(.dina(n1324), .dinb(n1225), .dout(n1332));
  jand g01043(.dina(n1229), .dinb(n989), .dout(n1333));
  jand g01044(.dina(n1333), .dinb(n1320), .dout(n1334));
  jor  g01045(.dina(n1334), .dinb(n1332), .dout(n1335));
  jand g01046(.dina(n1335), .dinb(n435), .dout(n1336));
  jnot g01047(.din(n1336), .dout(n1337));
  jand g01048(.dina(n1324), .dinb(n1233), .dout(n1338));
  jxor g01049(.dina(n1318), .dinb(n1317), .dout(n1339));
  jand g01050(.dina(n1339), .dinb(quotient51 ), .dout(n1340));
  jor  g01051(.dina(n1340), .dinb(n1338), .dout(n1341));
  jand g01052(.dina(n1341), .dinb(n440), .dout(n1342));
  jnot g01053(.din(n1342), .dout(n1343));
  jand g01054(.dina(n1328), .dinb(n439), .dout(n1344));
  jnot g01055(.din(n1344), .dout(n1345));
  jand g01056(.dina(n1324), .dinb(n1239), .dout(n1346));
  jxor g01057(.dina(n1312), .dinb(n1311), .dout(n1347));
  jand g01058(.dina(n1347), .dinb(quotient51 ), .dout(n1348));
  jor  g01059(.dina(n1348), .dinb(n1346), .dout(n1349));
  jand g01060(.dina(n1349), .dinb(n325), .dout(n1350));
  jnot g01061(.din(n1350), .dout(n1351));
  jand g01062(.dina(n1324), .dinb(n1244), .dout(n1352));
  jxor g01063(.dina(n1309), .dinb(n1308), .dout(n1353));
  jand g01064(.dina(n1353), .dinb(quotient51 ), .dout(n1354));
  jor  g01065(.dina(n1354), .dinb(n1352), .dout(n1355));
  jand g01066(.dina(n1355), .dinb(n324), .dout(n1356));
  jnot g01067(.din(n1356), .dout(n1357));
  jand g01068(.dina(n1324), .dinb(n1249), .dout(n1358));
  jxor g01069(.dina(n1306), .dinb(n1305), .dout(n1359));
  jand g01070(.dina(n1359), .dinb(quotient51 ), .dout(n1360));
  jor  g01071(.dina(n1360), .dinb(n1358), .dout(n1361));
  jand g01072(.dina(n1361), .dinb(n323), .dout(n1362));
  jnot g01073(.din(n1362), .dout(n1363));
  jand g01074(.dina(n1324), .dinb(n1254), .dout(n1364));
  jxor g01075(.dina(n1303), .dinb(n1302), .dout(n1365));
  jand g01076(.dina(n1365), .dinb(quotient51 ), .dout(n1366));
  jor  g01077(.dina(n1366), .dinb(n1364), .dout(n1367));
  jand g01078(.dina(n1367), .dinb(n335), .dout(n1368));
  jnot g01079(.din(n1368), .dout(n1369));
  jand g01080(.dina(n1324), .dinb(n1259), .dout(n1370));
  jxor g01081(.dina(n1300), .dinb(n1299), .dout(n1371));
  jand g01082(.dina(n1371), .dinb(quotient51 ), .dout(n1372));
  jor  g01083(.dina(n1372), .dinb(n1370), .dout(n1373));
  jand g01084(.dina(n1373), .dinb(n334), .dout(n1374));
  jnot g01085(.din(n1374), .dout(n1375));
  jand g01086(.dina(n1324), .dinb(n1264), .dout(n1376));
  jxor g01087(.dina(n1297), .dinb(n1296), .dout(n1377));
  jand g01088(.dina(n1377), .dinb(quotient51 ), .dout(n1378));
  jor  g01089(.dina(n1378), .dinb(n1376), .dout(n1379));
  jand g01090(.dina(n1379), .dinb(n338), .dout(n1380));
  jnot g01091(.din(n1380), .dout(n1381));
  jand g01092(.dina(n1324), .dinb(n1269), .dout(n1382));
  jxor g01093(.dina(n1294), .dinb(n1293), .dout(n1383));
  jand g01094(.dina(n1383), .dinb(quotient51 ), .dout(n1384));
  jor  g01095(.dina(n1384), .dinb(n1382), .dout(n1385));
  jand g01096(.dina(n1385), .dinb(n337), .dout(n1386));
  jnot g01097(.din(n1386), .dout(n1387));
  jand g01098(.dina(n1324), .dinb(n19448), .dout(n1388));
  jxor g01099(.dina(n1291), .dinb(n1290), .dout(n1389));
  jand g01100(.dina(n1389), .dinb(quotient51 ), .dout(n1390));
  jor  g01101(.dina(n1390), .dinb(n1388), .dout(n1391));
  jand g01102(.dina(n1391), .dinb(n344), .dout(n1392));
  jnot g01103(.din(n1392), .dout(n1393));
  jand g01104(.dina(n1324), .dinb(n1283), .dout(n1394));
  jxor g01105(.dina(n1288), .dinb(n1287), .dout(n1395));
  jand g01106(.dina(n1395), .dinb(quotient51 ), .dout(n1396));
  jor  g01107(.dina(n1396), .dinb(n1394), .dout(n1397));
  jand g01108(.dina(n1397), .dinb(n348), .dout(n1398));
  jnot g01109(.din(n1398), .dout(n1399));
  jand g01110(.dina(n435), .dinb(b0 ), .dout(n1400));
  jand g01111(.dina(n1400), .dinb(n1330), .dout(n1401));
  jand g01112(.dina(n1401), .dinb(n1322), .dout(n1402));
  jor  g01113(.dina(n1402), .dinb(n1285), .dout(n1403));
  jand g01114(.dina(n1286), .dinb(n989), .dout(n1404));
  jand g01115(.dina(n1404), .dinb(n1322), .dout(n1405));
  jnot g01116(.din(n1405), .dout(n1406));
  jand g01117(.dina(n1406), .dinb(n1403), .dout(n1407));
  jor  g01118(.dina(n1407), .dinb(b1 ), .dout(n1408));
  jnot g01119(.din(a50 ), .dout(n1409));
  jand g01120(.dina(b0 ), .dinb(n1409), .dout(n1410));
  jxor g01121(.dina(n1407), .dinb(n258), .dout(n1411));
  jor  g01122(.dina(n1411), .dinb(n1410), .dout(n1412));
  jand g01123(.dina(n1412), .dinb(n1408), .dout(n1413));
  jxor g01124(.dina(n1397), .dinb(n348), .dout(n1414));
  jnot g01125(.din(n1414), .dout(n1415));
  jor  g01126(.dina(n1415), .dinb(n1413), .dout(n1416));
  jand g01127(.dina(n1416), .dinb(n1399), .dout(n1417));
  jxor g01128(.dina(n1391), .dinb(n344), .dout(n1418));
  jnot g01129(.din(n1418), .dout(n1419));
  jor  g01130(.dina(n1419), .dinb(n1417), .dout(n1420));
  jand g01131(.dina(n1420), .dinb(n1393), .dout(n1421));
  jxor g01132(.dina(n1385), .dinb(n337), .dout(n1422));
  jnot g01133(.din(n1422), .dout(n1423));
  jor  g01134(.dina(n1423), .dinb(n1421), .dout(n1424));
  jand g01135(.dina(n1424), .dinb(n1387), .dout(n1425));
  jxor g01136(.dina(n1379), .dinb(n338), .dout(n1426));
  jnot g01137(.din(n1426), .dout(n1427));
  jor  g01138(.dina(n1427), .dinb(n1425), .dout(n1428));
  jand g01139(.dina(n1428), .dinb(n1381), .dout(n1429));
  jxor g01140(.dina(n1373), .dinb(n334), .dout(n1430));
  jnot g01141(.din(n1430), .dout(n1431));
  jor  g01142(.dina(n1431), .dinb(n1429), .dout(n1432));
  jand g01143(.dina(n1432), .dinb(n1375), .dout(n1433));
  jxor g01144(.dina(n1367), .dinb(n335), .dout(n1434));
  jnot g01145(.din(n1434), .dout(n1435));
  jor  g01146(.dina(n1435), .dinb(n1433), .dout(n1436));
  jand g01147(.dina(n1436), .dinb(n1369), .dout(n1437));
  jxor g01148(.dina(n1361), .dinb(n323), .dout(n1438));
  jnot g01149(.din(n1438), .dout(n1439));
  jor  g01150(.dina(n1439), .dinb(n1437), .dout(n1440));
  jand g01151(.dina(n1440), .dinb(n1363), .dout(n1441));
  jxor g01152(.dina(n1355), .dinb(n324), .dout(n1442));
  jnot g01153(.din(n1442), .dout(n1443));
  jor  g01154(.dina(n1443), .dinb(n1441), .dout(n1444));
  jand g01155(.dina(n1444), .dinb(n1357), .dout(n1445));
  jxor g01156(.dina(n1349), .dinb(n325), .dout(n1446));
  jnot g01157(.din(n1446), .dout(n1447));
  jor  g01158(.dina(n1447), .dinb(n1445), .dout(n1448));
  jand g01159(.dina(n1448), .dinb(n1351), .dout(n1449));
  jxor g01160(.dina(n1328), .dinb(n439), .dout(n1450));
  jnot g01161(.din(n1450), .dout(n1451));
  jor  g01162(.dina(n1451), .dinb(n1449), .dout(n1452));
  jand g01163(.dina(n1452), .dinb(n1345), .dout(n1453));
  jxor g01164(.dina(n1341), .dinb(n440), .dout(n1454));
  jnot g01165(.din(n1454), .dout(n1455));
  jor  g01166(.dina(n1455), .dinb(n1453), .dout(n1456));
  jand g01167(.dina(n1456), .dinb(n1343), .dout(n1457));
  jnot g01168(.din(n1335), .dout(n1458));
  jand g01169(.dina(n1458), .dinb(b13 ), .dout(n1459));
  jor  g01170(.dina(n1459), .dinb(n1457), .dout(n1460));
  jand g01171(.dina(n1460), .dinb(n1337), .dout(n1461));
  jor  g01172(.dina(n1461), .dinb(n1331), .dout(n1462));
  jand g01173(.dina(n1462), .dinb(n1328), .dout(n1463));
  jnot g01174(.din(n1462), .dout(quotient50 ));
  jnot g01175(.din(n1408), .dout(n1465));
  jnot g01176(.din(n1410), .dout(n1466));
  jxor g01177(.dina(n1407), .dinb(b1 ), .dout(n1467));
  jand g01178(.dina(n1467), .dinb(n1466), .dout(n1468));
  jor  g01179(.dina(n1468), .dinb(n1465), .dout(n1469));
  jand g01180(.dina(n1414), .dinb(n1469), .dout(n1470));
  jor  g01181(.dina(n1470), .dinb(n1398), .dout(n1471));
  jand g01182(.dina(n1418), .dinb(n1471), .dout(n1472));
  jor  g01183(.dina(n1472), .dinb(n1392), .dout(n1473));
  jand g01184(.dina(n1422), .dinb(n1473), .dout(n1474));
  jor  g01185(.dina(n1474), .dinb(n1386), .dout(n1475));
  jand g01186(.dina(n1426), .dinb(n1475), .dout(n1476));
  jor  g01187(.dina(n1476), .dinb(n1380), .dout(n1477));
  jand g01188(.dina(n1430), .dinb(n1477), .dout(n1478));
  jor  g01189(.dina(n1478), .dinb(n1374), .dout(n1479));
  jand g01190(.dina(n1434), .dinb(n1479), .dout(n1480));
  jor  g01191(.dina(n1480), .dinb(n1368), .dout(n1481));
  jand g01192(.dina(n1438), .dinb(n1481), .dout(n1482));
  jor  g01193(.dina(n1482), .dinb(n1362), .dout(n1483));
  jand g01194(.dina(n1442), .dinb(n1483), .dout(n1484));
  jor  g01195(.dina(n1484), .dinb(n1356), .dout(n1485));
  jand g01196(.dina(n1446), .dinb(n1485), .dout(n1486));
  jor  g01197(.dina(n1486), .dinb(n1350), .dout(n1487));
  jxor g01198(.dina(n1450), .dinb(n1487), .dout(n1488));
  jand g01199(.dina(n1488), .dinb(quotient50 ), .dout(n1489));
  jor  g01200(.dina(n1489), .dinb(n1463), .dout(n1490));
  jand g01201(.dina(n1462), .dinb(n1335), .dout(n1491));
  jand g01202(.dina(n1450), .dinb(n1487), .dout(n1492));
  jor  g01203(.dina(n1492), .dinb(n1344), .dout(n1493));
  jand g01204(.dina(n1454), .dinb(n1493), .dout(n1494));
  jor  g01205(.dina(n1494), .dinb(n1342), .dout(n1495));
  jand g01206(.dina(n1336), .dinb(n1330), .dout(n1496));
  jand g01207(.dina(n1496), .dinb(n1495), .dout(n1497));
  jor  g01208(.dina(n1497), .dinb(n1491), .dout(n1498));
  jand g01209(.dina(n1498), .dinb(n1330), .dout(n1499));
  jand g01210(.dina(n988), .dinb(n434), .dout(n1500));
  jand g01211(.dina(n1462), .dinb(n1341), .dout(n1501));
  jxor g01212(.dina(n1454), .dinb(n1493), .dout(n1502));
  jand g01213(.dina(n1502), .dinb(quotient50 ), .dout(n1503));
  jor  g01214(.dina(n1503), .dinb(n1501), .dout(n1504));
  jand g01215(.dina(n1504), .dinb(n435), .dout(n1505));
  jand g01216(.dina(n1490), .dinb(n440), .dout(n1506));
  jand g01217(.dina(n1462), .dinb(n1349), .dout(n1507));
  jxor g01218(.dina(n1446), .dinb(n1485), .dout(n1508));
  jand g01219(.dina(n1508), .dinb(quotient50 ), .dout(n1509));
  jor  g01220(.dina(n1509), .dinb(n1507), .dout(n1510));
  jand g01221(.dina(n1510), .dinb(n439), .dout(n1511));
  jand g01222(.dina(n1462), .dinb(n1355), .dout(n1512));
  jxor g01223(.dina(n1442), .dinb(n1483), .dout(n1513));
  jand g01224(.dina(n1513), .dinb(quotient50 ), .dout(n1514));
  jor  g01225(.dina(n1514), .dinb(n1512), .dout(n1515));
  jand g01226(.dina(n1515), .dinb(n325), .dout(n1516));
  jand g01227(.dina(n1462), .dinb(n1361), .dout(n1517));
  jxor g01228(.dina(n1438), .dinb(n1481), .dout(n1518));
  jand g01229(.dina(n1518), .dinb(quotient50 ), .dout(n1519));
  jor  g01230(.dina(n1519), .dinb(n1517), .dout(n1520));
  jand g01231(.dina(n1520), .dinb(n324), .dout(n1521));
  jand g01232(.dina(n1462), .dinb(n1367), .dout(n1522));
  jxor g01233(.dina(n1434), .dinb(n1479), .dout(n1523));
  jand g01234(.dina(n1523), .dinb(quotient50 ), .dout(n1524));
  jor  g01235(.dina(n1524), .dinb(n1522), .dout(n1525));
  jand g01236(.dina(n1525), .dinb(n323), .dout(n1526));
  jand g01237(.dina(n1462), .dinb(n1373), .dout(n1527));
  jxor g01238(.dina(n1430), .dinb(n1477), .dout(n1528));
  jand g01239(.dina(n1528), .dinb(quotient50 ), .dout(n1529));
  jor  g01240(.dina(n1529), .dinb(n1527), .dout(n1530));
  jand g01241(.dina(n1530), .dinb(n335), .dout(n1531));
  jand g01242(.dina(n1462), .dinb(n1379), .dout(n1532));
  jxor g01243(.dina(n1426), .dinb(n1475), .dout(n1533));
  jand g01244(.dina(n1533), .dinb(quotient50 ), .dout(n1534));
  jor  g01245(.dina(n1534), .dinb(n1532), .dout(n1535));
  jand g01246(.dina(n1535), .dinb(n334), .dout(n1536));
  jand g01247(.dina(n1462), .dinb(n1385), .dout(n1537));
  jxor g01248(.dina(n1422), .dinb(n1473), .dout(n1538));
  jand g01249(.dina(n1538), .dinb(quotient50 ), .dout(n1539));
  jor  g01250(.dina(n1539), .dinb(n1537), .dout(n1540));
  jand g01251(.dina(n1540), .dinb(n338), .dout(n1541));
  jand g01252(.dina(n1462), .dinb(n1391), .dout(n1542));
  jxor g01253(.dina(n1418), .dinb(n1471), .dout(n1543));
  jand g01254(.dina(n1543), .dinb(quotient50 ), .dout(n1544));
  jor  g01255(.dina(n1544), .dinb(n1542), .dout(n1545));
  jand g01256(.dina(n1545), .dinb(n337), .dout(n1546));
  jand g01257(.dina(n1462), .dinb(n1397), .dout(n1547));
  jxor g01258(.dina(n1414), .dinb(n1469), .dout(n1548));
  jand g01259(.dina(n1548), .dinb(quotient50 ), .dout(n1549));
  jor  g01260(.dina(n1549), .dinb(n1547), .dout(n1550));
  jand g01261(.dina(n1550), .dinb(n344), .dout(n1551));
  jxor g01262(.dina(n1467), .dinb(n1466), .dout(n1553));
  jand g01263(.dina(n1553), .dinb(quotient50 ), .dout(n1554));
  jnot g01264(.din(n1459), .dout(n1559));
  jand g01265(.dina(n1559), .dinb(n1495), .dout(n1560));
  jor  g01266(.dina(n1560), .dinb(n1336), .dout(n1561));
  jand g01267(.dina(n988), .dinb(b0 ), .dout(n1562));
  jand g01268(.dina(n1562), .dinb(n433), .dout(n1563));
  jand g01269(.dina(n1563), .dinb(n1329), .dout(n1564));
  jand g01270(.dina(n1564), .dinb(n1561), .dout(n1565));
  jor  g01271(.dina(n1565), .dinb(n1409), .dout(n1566));
  jor  g01272(.dina(n1462), .dinb(n1466), .dout(n1567));
  jand g01273(.dina(n1567), .dinb(n1566), .dout(n1568));
  jor  g01274(.dina(n1568), .dinb(b1 ), .dout(n1569));
  jnot g01275(.din(n1569), .dout(n1570));
  jnot g01276(.din(a49 ), .dout(n1571));
  jand g01277(.dina(b0 ), .dinb(n1571), .dout(n1572));
  jnot g01278(.din(n1572), .dout(n1573));
  jxor g01279(.dina(n1568), .dinb(b1 ), .dout(n1574));
  jand g01280(.dina(n1574), .dinb(n1573), .dout(n1575));
  jor  g01281(.dina(n1575), .dinb(n1570), .dout(n1576));
  jand g01282(.dina(n19808), .dinb(n1576), .dout(n1578));
  jor  g01283(.dina(n1578), .dinb(n19792), .dout(n1579));
  jxor g01284(.dina(n1550), .dinb(n344), .dout(n1580));
  jand g01285(.dina(n1580), .dinb(n1579), .dout(n1581));
  jor  g01286(.dina(n1581), .dinb(n1551), .dout(n1582));
  jxor g01287(.dina(n1545), .dinb(n337), .dout(n1583));
  jand g01288(.dina(n1583), .dinb(n1582), .dout(n1584));
  jor  g01289(.dina(n1584), .dinb(n1546), .dout(n1585));
  jxor g01290(.dina(n1540), .dinb(n338), .dout(n1586));
  jand g01291(.dina(n1586), .dinb(n1585), .dout(n1587));
  jor  g01292(.dina(n1587), .dinb(n1541), .dout(n1588));
  jxor g01293(.dina(n1535), .dinb(n334), .dout(n1589));
  jand g01294(.dina(n1589), .dinb(n1588), .dout(n1590));
  jor  g01295(.dina(n1590), .dinb(n1536), .dout(n1591));
  jxor g01296(.dina(n1530), .dinb(n335), .dout(n1592));
  jand g01297(.dina(n1592), .dinb(n1591), .dout(n1593));
  jor  g01298(.dina(n1593), .dinb(n1531), .dout(n1594));
  jxor g01299(.dina(n1525), .dinb(n323), .dout(n1595));
  jand g01300(.dina(n1595), .dinb(n1594), .dout(n1596));
  jor  g01301(.dina(n1596), .dinb(n1526), .dout(n1597));
  jxor g01302(.dina(n1520), .dinb(n324), .dout(n1598));
  jand g01303(.dina(n1598), .dinb(n1597), .dout(n1599));
  jor  g01304(.dina(n1599), .dinb(n1521), .dout(n1600));
  jxor g01305(.dina(n1515), .dinb(n325), .dout(n1601));
  jand g01306(.dina(n1601), .dinb(n1600), .dout(n1602));
  jor  g01307(.dina(n1602), .dinb(n1516), .dout(n1603));
  jxor g01308(.dina(n1510), .dinb(n439), .dout(n1604));
  jand g01309(.dina(n1604), .dinb(n1603), .dout(n1605));
  jor  g01310(.dina(n1605), .dinb(n1511), .dout(n1606));
  jxor g01311(.dina(n1490), .dinb(n440), .dout(n1607));
  jand g01312(.dina(n1607), .dinb(n1606), .dout(n1608));
  jor  g01313(.dina(n1608), .dinb(n1506), .dout(n1609));
  jxor g01314(.dina(n1504), .dinb(n435), .dout(n1610));
  jand g01315(.dina(n1610), .dinb(n1609), .dout(n1611));
  jor  g01316(.dina(n1611), .dinb(n1505), .dout(n1612));
  jxor g01317(.dina(n1498), .dinb(b14 ), .dout(n1613));
  jnot g01318(.din(n1613), .dout(n1614));
  jand g01319(.dina(n1614), .dinb(n1612), .dout(n1615));
  jand g01320(.dina(n1615), .dinb(n1500), .dout(n1616));
  jor  g01321(.dina(n1616), .dinb(n1499), .dout(quotient49 ));
  jxor g01322(.dina(n1607), .dinb(n1606), .dout(n1620));
  jand g01323(.dina(n1620), .dinb(quotient49 ), .dout(n1621));
  jxor g01324(.dina(n1614), .dinb(n1612), .dout(n1623));
  jor  g01325(.dina(n1623), .dinb(n19900), .dout(n1624));
  jor  g01326(.dina(n1616), .dinb(n1498), .dout(n1625));
  jand g01327(.dina(n1625), .dinb(n1624), .dout(n1626));
  jand g01328(.dina(n1626), .dinb(n432), .dout(n1630));
  jxor g01329(.dina(n1610), .dinb(n1609), .dout(n1632));
  jand g01330(.dina(n1632), .dinb(quotient49 ), .dout(n1633));
  jxor g01331(.dina(n1604), .dinb(n1603), .dout(n1638));
  jand g01332(.dina(n1638), .dinb(quotient49 ), .dout(n1639));
  jxor g01333(.dina(n1601), .dinb(n1600), .dout(n1643));
  jand g01334(.dina(n1643), .dinb(quotient49 ), .dout(n1644));
  jxor g01335(.dina(n1598), .dinb(n1597), .dout(n1648));
  jand g01336(.dina(n1648), .dinb(quotient49 ), .dout(n1649));
  jxor g01337(.dina(n1595), .dinb(n1594), .dout(n1653));
  jand g01338(.dina(n1653), .dinb(quotient49 ), .dout(n1654));
  jxor g01339(.dina(n1592), .dinb(n1591), .dout(n1658));
  jand g01340(.dina(n1658), .dinb(quotient49 ), .dout(n1659));
  jxor g01341(.dina(n1589), .dinb(n1588), .dout(n1663));
  jand g01342(.dina(n1663), .dinb(quotient49 ), .dout(n1664));
  jxor g01343(.dina(n1586), .dinb(n1585), .dout(n1668));
  jand g01344(.dina(n1668), .dinb(quotient49 ), .dout(n1669));
  jxor g01345(.dina(n1583), .dinb(n1582), .dout(n1673));
  jand g01346(.dina(n1673), .dinb(quotient49 ), .dout(n1674));
  jxor g01347(.dina(n1580), .dinb(n1579), .dout(n1678));
  jand g01348(.dina(n1678), .dinb(quotient49 ), .dout(n1679));
  jxor g01349(.dina(n19808), .dinb(n1576), .dout(n1683));
  jand g01350(.dina(n1683), .dinb(quotient49 ), .dout(n1684));
  jxor g01351(.dina(n1574), .dinb(n1573), .dout(n1688));
  jand g01352(.dina(quotient49 ), .dinb(b0 ), .dout(n1694));
  jor  g01353(.dina(n1694), .dinb(n1571), .dout(n1695));
  jand g01354(.dina(quotient49 ), .dinb(n1572), .dout(n1696));
  jand g01355(.dina(n19968), .dinb(n1695), .dout(n1698));
  jnot g01356(.din(a48 ), .dout(n1701));
  jand g01357(.dina(b0 ), .dinb(n1701), .dout(n1702));
  jnot g01358(.din(n1702), .dout(n1703));
  jxor g01359(.dina(n1698), .dinb(b1 ), .dout(n1704));
  jand g01360(.dina(n1704), .dinb(n1703), .dout(n1705));
  jor  g01361(.dina(n1705), .dinb(n19971), .dout(n1706));
  jand g01362(.dina(n19978), .dinb(n1706), .dout(n1708));
  jor  g01363(.dina(n1708), .dinb(n19965), .dout(n1709));
  jand g01364(.dina(n19981), .dinb(n1709), .dout(n1711));
  jor  g01365(.dina(n1711), .dinb(n19960), .dout(n1712));
  jand g01366(.dina(n19984), .dinb(n1712), .dout(n1714));
  jor  g01367(.dina(n1714), .dinb(n19955), .dout(n1715));
  jand g01368(.dina(n19987), .dinb(n1715), .dout(n1717));
  jor  g01369(.dina(n1717), .dinb(n19950), .dout(n1718));
  jand g01370(.dina(n19990), .dinb(n1718), .dout(n1720));
  jor  g01371(.dina(n1720), .dinb(n19945), .dout(n1721));
  jand g01372(.dina(n19993), .dinb(n1721), .dout(n1723));
  jor  g01373(.dina(n1723), .dinb(n19940), .dout(n1724));
  jand g01374(.dina(n19996), .dinb(n1724), .dout(n1726));
  jor  g01375(.dina(n1726), .dinb(n19935), .dout(n1727));
  jand g01376(.dina(n19999), .dinb(n1727), .dout(n1729));
  jor  g01377(.dina(n1729), .dinb(n19930), .dout(n1730));
  jand g01378(.dina(n20002), .dinb(n1730), .dout(n1732));
  jor  g01379(.dina(n1732), .dinb(n19925), .dout(n1733));
  jand g01380(.dina(n20005), .dinb(n1733), .dout(n1735));
  jor  g01381(.dina(n1735), .dinb(n19920), .dout(n1736));
  jand g01382(.dina(n20008), .dinb(n1736), .dout(n1738));
  jor  g01383(.dina(n1738), .dinb(n19915), .dout(n1739));
  jand g01384(.dina(n20011), .dinb(n1739), .dout(n1741));
  jor  g01385(.dina(n1741), .dinb(n19910), .dout(n1742));
  jand g01386(.dina(n20014), .dinb(n1742), .dout(n1744));
  jor  g01387(.dina(n1744), .dinb(n19905), .dout(n1745));
  jor  g01388(.dina(n1745), .dinb(n1630), .dout(n1746));
  jand g01389(.dina(n1746), .dinb(n19897), .dout(n1747));
  jand g01390(.dina(n1747), .dinb(n594), .dout(quotient48 ));
  jnot g01391(.din(quotient48 ), .dout(n1749));
  jand g01392(.dina(n1749), .dinb(n19909), .dout(n1750));
  jxor g01393(.dina(n20011), .dinb(n1739), .dout(n1751));
  jand g01394(.dina(n1751), .dinb(quotient48 ), .dout(n1752));
  jor  g01395(.dina(n1752), .dinb(n1750), .dout(n1753));
  jand g01396(.dina(n1749), .dinb(n1626), .dout(n1754));
  jand g01397(.dina(n1630), .dinb(n594), .dout(n1755));
  jand g01398(.dina(n1755), .dinb(n1745), .dout(n1756));
  jor  g01399(.dina(n1756), .dinb(n1754), .dout(n1757));
  jand g01400(.dina(n1757), .dinb(n433), .dout(n1758));
  jand g01401(.dina(n1749), .dinb(n19904), .dout(n1759));
  jxor g01402(.dina(n20014), .dinb(n1742), .dout(n1760));
  jand g01403(.dina(n1760), .dinb(quotient48 ), .dout(n1761));
  jor  g01404(.dina(n1761), .dinb(n1759), .dout(n1762));
  jand g01405(.dina(n1762), .dinb(n432), .dout(n1763));
  jand g01406(.dina(n1753), .dinb(n436), .dout(n1764));
  jand g01407(.dina(n1749), .dinb(n19914), .dout(n1765));
  jxor g01408(.dina(n20008), .dinb(n1736), .dout(n1766));
  jand g01409(.dina(n1766), .dinb(quotient48 ), .dout(n1767));
  jor  g01410(.dina(n1767), .dinb(n1765), .dout(n1768));
  jand g01411(.dina(n1768), .dinb(n435), .dout(n1769));
  jand g01412(.dina(n1749), .dinb(n19919), .dout(n1770));
  jxor g01413(.dina(n20005), .dinb(n1733), .dout(n1771));
  jand g01414(.dina(n1771), .dinb(quotient48 ), .dout(n1772));
  jor  g01415(.dina(n1772), .dinb(n1770), .dout(n1773));
  jand g01416(.dina(n1773), .dinb(n440), .dout(n1774));
  jand g01417(.dina(n1749), .dinb(n19924), .dout(n1775));
  jxor g01418(.dina(n20002), .dinb(n1730), .dout(n1776));
  jand g01419(.dina(n1776), .dinb(quotient48 ), .dout(n1777));
  jor  g01420(.dina(n1777), .dinb(n1775), .dout(n1778));
  jand g01421(.dina(n1778), .dinb(n439), .dout(n1779));
  jand g01422(.dina(n1749), .dinb(n19929), .dout(n1780));
  jxor g01423(.dina(n19999), .dinb(n1727), .dout(n1781));
  jand g01424(.dina(n1781), .dinb(quotient48 ), .dout(n1782));
  jor  g01425(.dina(n1782), .dinb(n1780), .dout(n1783));
  jand g01426(.dina(n1783), .dinb(n325), .dout(n1784));
  jand g01427(.dina(n1749), .dinb(n19934), .dout(n1785));
  jxor g01428(.dina(n19996), .dinb(n1724), .dout(n1786));
  jand g01429(.dina(n1786), .dinb(quotient48 ), .dout(n1787));
  jor  g01430(.dina(n1787), .dinb(n1785), .dout(n1788));
  jand g01431(.dina(n1788), .dinb(n324), .dout(n1789));
  jand g01432(.dina(n1749), .dinb(n19939), .dout(n1790));
  jxor g01433(.dina(n19993), .dinb(n1721), .dout(n1791));
  jand g01434(.dina(n1791), .dinb(quotient48 ), .dout(n1792));
  jor  g01435(.dina(n1792), .dinb(n1790), .dout(n1793));
  jand g01436(.dina(n1793), .dinb(n323), .dout(n1794));
  jand g01437(.dina(n1749), .dinb(n19944), .dout(n1795));
  jxor g01438(.dina(n19990), .dinb(n1718), .dout(n1796));
  jand g01439(.dina(n1796), .dinb(quotient48 ), .dout(n1797));
  jor  g01440(.dina(n1797), .dinb(n1795), .dout(n1798));
  jand g01441(.dina(n1798), .dinb(n335), .dout(n1799));
  jand g01442(.dina(n1749), .dinb(n19949), .dout(n1800));
  jxor g01443(.dina(n19987), .dinb(n1715), .dout(n1801));
  jand g01444(.dina(n1801), .dinb(quotient48 ), .dout(n1802));
  jor  g01445(.dina(n1802), .dinb(n1800), .dout(n1803));
  jand g01446(.dina(n1803), .dinb(n334), .dout(n1804));
  jand g01447(.dina(n1749), .dinb(n19954), .dout(n1805));
  jxor g01448(.dina(n19984), .dinb(n1712), .dout(n1806));
  jand g01449(.dina(n1806), .dinb(quotient48 ), .dout(n1807));
  jor  g01450(.dina(n1807), .dinb(n1805), .dout(n1808));
  jand g01451(.dina(n1808), .dinb(n338), .dout(n1809));
  jand g01452(.dina(n1749), .dinb(n19959), .dout(n1810));
  jxor g01453(.dina(n19981), .dinb(n1709), .dout(n1811));
  jand g01454(.dina(n1811), .dinb(quotient48 ), .dout(n1812));
  jor  g01455(.dina(n1812), .dinb(n1810), .dout(n1813));
  jand g01456(.dina(n1813), .dinb(n337), .dout(n1814));
  jand g01457(.dina(n1749), .dinb(n19964), .dout(n1815));
  jxor g01458(.dina(n19978), .dinb(n1706), .dout(n1816));
  jand g01459(.dina(n1816), .dinb(quotient48 ), .dout(n1817));
  jor  g01460(.dina(n1817), .dinb(n1815), .dout(n1818));
  jand g01461(.dina(n1818), .dinb(n344), .dout(n1819));
  jand g01462(.dina(n1749), .dinb(n19970), .dout(n1820));
  jxor g01463(.dina(n1704), .dinb(n1703), .dout(n1821));
  jand g01464(.dina(n1821), .dinb(quotient48 ), .dout(n1822));
  jor  g01465(.dina(n1822), .dinb(n1820), .dout(n1823));
  jand g01466(.dina(n1823), .dinb(n348), .dout(n1824));
  jand g01467(.dina(n1747), .dinb(n1563), .dout(n1825));
  jor  g01468(.dina(n1825), .dinb(n1701), .dout(n1826));
  jand g01469(.dina(n1702), .dinb(n594), .dout(n1827));
  jand g01470(.dina(n1827), .dinb(n1747), .dout(n1828));
  jand g01471(.dina(n20164), .dinb(n1826), .dout(n1830));
  jnot g01472(.din(a47 ), .dout(n1833));
  jand g01473(.dina(b0 ), .dinb(n1833), .dout(n1834));
  jnot g01474(.din(n1834), .dout(n1835));
  jxor g01475(.dina(n1830), .dinb(b1 ), .dout(n1836));
  jand g01476(.dina(n1836), .dinb(n1835), .dout(n1837));
  jor  g01477(.dina(n1837), .dinb(n20167), .dout(n1838));
  jxor g01478(.dina(n1823), .dinb(n348), .dout(n1839));
  jand g01479(.dina(n1839), .dinb(n1838), .dout(n1840));
  jor  g01480(.dina(n1840), .dinb(n1824), .dout(n1841));
  jxor g01481(.dina(n1818), .dinb(n344), .dout(n1842));
  jand g01482(.dina(n1842), .dinb(n1841), .dout(n1843));
  jor  g01483(.dina(n1843), .dinb(n1819), .dout(n1844));
  jxor g01484(.dina(n1813), .dinb(n337), .dout(n1845));
  jand g01485(.dina(n1845), .dinb(n1844), .dout(n1846));
  jor  g01486(.dina(n1846), .dinb(n1814), .dout(n1847));
  jxor g01487(.dina(n1808), .dinb(n338), .dout(n1848));
  jand g01488(.dina(n1848), .dinb(n1847), .dout(n1849));
  jor  g01489(.dina(n1849), .dinb(n1809), .dout(n1850));
  jxor g01490(.dina(n1803), .dinb(n334), .dout(n1851));
  jand g01491(.dina(n1851), .dinb(n1850), .dout(n1852));
  jor  g01492(.dina(n1852), .dinb(n1804), .dout(n1853));
  jxor g01493(.dina(n1798), .dinb(n335), .dout(n1854));
  jand g01494(.dina(n1854), .dinb(n1853), .dout(n1855));
  jor  g01495(.dina(n1855), .dinb(n1799), .dout(n1856));
  jxor g01496(.dina(n1793), .dinb(n323), .dout(n1857));
  jand g01497(.dina(n1857), .dinb(n1856), .dout(n1858));
  jor  g01498(.dina(n1858), .dinb(n1794), .dout(n1859));
  jxor g01499(.dina(n1788), .dinb(n324), .dout(n1860));
  jand g01500(.dina(n1860), .dinb(n1859), .dout(n1861));
  jor  g01501(.dina(n1861), .dinb(n1789), .dout(n1862));
  jxor g01502(.dina(n1783), .dinb(n325), .dout(n1863));
  jand g01503(.dina(n1863), .dinb(n1862), .dout(n1864));
  jor  g01504(.dina(n1864), .dinb(n1784), .dout(n1865));
  jxor g01505(.dina(n1778), .dinb(n439), .dout(n1866));
  jand g01506(.dina(n1866), .dinb(n1865), .dout(n1867));
  jor  g01507(.dina(n1867), .dinb(n1779), .dout(n1868));
  jxor g01508(.dina(n1773), .dinb(n440), .dout(n1869));
  jand g01509(.dina(n1869), .dinb(n1868), .dout(n1870));
  jor  g01510(.dina(n1870), .dinb(n1774), .dout(n1871));
  jxor g01511(.dina(n1768), .dinb(n435), .dout(n1872));
  jand g01512(.dina(n1872), .dinb(n1871), .dout(n1873));
  jor  g01513(.dina(n1873), .dinb(n1769), .dout(n1874));
  jxor g01514(.dina(n1753), .dinb(n436), .dout(n1875));
  jand g01515(.dina(n1875), .dinb(n1874), .dout(n1876));
  jor  g01516(.dina(n1876), .dinb(n1764), .dout(n1877));
  jxor g01517(.dina(n1762), .dinb(n432), .dout(n1878));
  jand g01518(.dina(n1878), .dinb(n1877), .dout(n1879));
  jor  g01519(.dina(n1879), .dinb(n1763), .dout(n1880));
  jnot g01520(.din(n1757), .dout(n1881));
  jand g01521(.dina(n1881), .dinb(b16 ), .dout(n1882));
  jnot g01522(.din(n1882), .dout(n1883));
  jand g01523(.dina(n1883), .dinb(n1880), .dout(n1884));
  jor  g01524(.dina(n1884), .dinb(n1758), .dout(n1885));
  jand g01525(.dina(n1885), .dinb(n988), .dout(quotient47 ));
  jnot g01526(.din(quotient47 ), .dout(n1887));
  jand g01527(.dina(n1887), .dinb(n1753), .dout(n1888));
  jxor g01528(.dina(n1875), .dinb(n1874), .dout(n1889));
  jand g01529(.dina(n1889), .dinb(quotient47 ), .dout(n1890));
  jor  g01530(.dina(n1890), .dinb(n1888), .dout(n1891));
  jand g01531(.dina(n1887), .dinb(n1757), .dout(n1892));
  jand g01532(.dina(n1758), .dinb(n988), .dout(n1893));
  jand g01533(.dina(n1893), .dinb(n1880), .dout(n1894));
  jor  g01534(.dina(n1894), .dinb(n1892), .dout(n1895));
  jand g01535(.dina(n1895), .dinb(n988), .dout(n1896));
  jor  g01536(.dina(n319), .dinb(n318), .dout(n1897));
  jand g01537(.dina(n1887), .dinb(n1762), .dout(n1899));
  jxor g01538(.dina(n1878), .dinb(n1877), .dout(n1900));
  jand g01539(.dina(n1900), .dinb(quotient47 ), .dout(n1901));
  jor  g01540(.dina(n1901), .dinb(n1899), .dout(n1902));
  jand g01541(.dina(n1902), .dinb(n433), .dout(n1903));
  jand g01542(.dina(n1891), .dinb(n432), .dout(n1904));
  jand g01543(.dina(n1887), .dinb(n1768), .dout(n1905));
  jxor g01544(.dina(n1872), .dinb(n1871), .dout(n1906));
  jand g01545(.dina(n1906), .dinb(quotient47 ), .dout(n1907));
  jor  g01546(.dina(n1907), .dinb(n1905), .dout(n1908));
  jand g01547(.dina(n1908), .dinb(n436), .dout(n1909));
  jand g01548(.dina(n1887), .dinb(n1773), .dout(n1910));
  jxor g01549(.dina(n1869), .dinb(n1868), .dout(n1911));
  jand g01550(.dina(n1911), .dinb(quotient47 ), .dout(n1912));
  jor  g01551(.dina(n1912), .dinb(n1910), .dout(n1913));
  jand g01552(.dina(n1913), .dinb(n435), .dout(n1914));
  jand g01553(.dina(n1887), .dinb(n1778), .dout(n1915));
  jxor g01554(.dina(n1866), .dinb(n1865), .dout(n1916));
  jand g01555(.dina(n1916), .dinb(quotient47 ), .dout(n1917));
  jor  g01556(.dina(n1917), .dinb(n1915), .dout(n1918));
  jand g01557(.dina(n1918), .dinb(n440), .dout(n1919));
  jand g01558(.dina(n1887), .dinb(n1783), .dout(n1920));
  jxor g01559(.dina(n1863), .dinb(n1862), .dout(n1921));
  jand g01560(.dina(n1921), .dinb(quotient47 ), .dout(n1922));
  jor  g01561(.dina(n1922), .dinb(n1920), .dout(n1923));
  jand g01562(.dina(n1923), .dinb(n439), .dout(n1924));
  jand g01563(.dina(n1887), .dinb(n1788), .dout(n1925));
  jxor g01564(.dina(n1860), .dinb(n1859), .dout(n1926));
  jand g01565(.dina(n1926), .dinb(quotient47 ), .dout(n1927));
  jor  g01566(.dina(n1927), .dinb(n1925), .dout(n1928));
  jand g01567(.dina(n1928), .dinb(n325), .dout(n1929));
  jand g01568(.dina(n1887), .dinb(n1793), .dout(n1930));
  jxor g01569(.dina(n1857), .dinb(n1856), .dout(n1931));
  jand g01570(.dina(n1931), .dinb(quotient47 ), .dout(n1932));
  jor  g01571(.dina(n1932), .dinb(n1930), .dout(n1933));
  jand g01572(.dina(n1933), .dinb(n324), .dout(n1934));
  jand g01573(.dina(n1887), .dinb(n1798), .dout(n1935));
  jxor g01574(.dina(n1854), .dinb(n1853), .dout(n1936));
  jand g01575(.dina(n1936), .dinb(quotient47 ), .dout(n1937));
  jor  g01576(.dina(n1937), .dinb(n1935), .dout(n1938));
  jand g01577(.dina(n1938), .dinb(n323), .dout(n1939));
  jand g01578(.dina(n1887), .dinb(n1803), .dout(n1940));
  jxor g01579(.dina(n1851), .dinb(n1850), .dout(n1941));
  jand g01580(.dina(n1941), .dinb(quotient47 ), .dout(n1942));
  jor  g01581(.dina(n1942), .dinb(n1940), .dout(n1943));
  jand g01582(.dina(n1943), .dinb(n335), .dout(n1944));
  jand g01583(.dina(n1887), .dinb(n1808), .dout(n1945));
  jxor g01584(.dina(n1848), .dinb(n1847), .dout(n1946));
  jand g01585(.dina(n1946), .dinb(quotient47 ), .dout(n1947));
  jor  g01586(.dina(n1947), .dinb(n1945), .dout(n1948));
  jand g01587(.dina(n1948), .dinb(n334), .dout(n1949));
  jand g01588(.dina(n1887), .dinb(n1813), .dout(n1950));
  jxor g01589(.dina(n1845), .dinb(n1844), .dout(n1951));
  jand g01590(.dina(n1951), .dinb(quotient47 ), .dout(n1952));
  jor  g01591(.dina(n1952), .dinb(n1950), .dout(n1953));
  jand g01592(.dina(n1953), .dinb(n338), .dout(n1954));
  jand g01593(.dina(n1887), .dinb(n1818), .dout(n1955));
  jxor g01594(.dina(n1842), .dinb(n1841), .dout(n1956));
  jand g01595(.dina(n1956), .dinb(quotient47 ), .dout(n1957));
  jor  g01596(.dina(n1957), .dinb(n1955), .dout(n1958));
  jand g01597(.dina(n1958), .dinb(n337), .dout(n1959));
  jand g01598(.dina(n1887), .dinb(n1823), .dout(n1960));
  jxor g01599(.dina(n1839), .dinb(n1838), .dout(n1961));
  jand g01600(.dina(n1961), .dinb(quotient47 ), .dout(n1962));
  jor  g01601(.dina(n1962), .dinb(n1960), .dout(n1963));
  jand g01602(.dina(n1963), .dinb(n344), .dout(n1964));
  jand g01603(.dina(n1887), .dinb(n20166), .dout(n1965));
  jxor g01604(.dina(n1836), .dinb(n1835), .dout(n1966));
  jand g01605(.dina(n1966), .dinb(quotient47 ), .dout(n1967));
  jor  g01606(.dina(n1967), .dinb(n1965), .dout(n1968));
  jand g01607(.dina(n1968), .dinb(n348), .dout(n1969));
  jnot g01608(.din(n318), .dout(n1970));
  jand g01609(.dina(n1970), .dinb(b0 ), .dout(n1971));
  jand g01610(.dina(n1971), .dinb(n416), .dout(n1972));
  jand g01611(.dina(n1972), .dinb(n423), .dout(n1973));
  jand g01612(.dina(n1973), .dinb(n1885), .dout(n1974));
  jor  g01613(.dina(n1974), .dinb(n1833), .dout(n1975));
  jand g01614(.dina(n1562), .dinb(n1833), .dout(n1976));
  jand g01615(.dina(n1976), .dinb(n1885), .dout(n1977));
  jand g01616(.dina(n20388), .dinb(n1975), .dout(n1979));
  jor  g01617(.dina(n1979), .dinb(b1 ), .dout(n1980));
  jnot g01618(.din(a46 ), .dout(n1982));
  jand g01619(.dina(b0 ), .dinb(n1982), .dout(n1983));
  jnot g01620(.din(n1983), .dout(n1984));
  jxor g01621(.dina(n1979), .dinb(b1 ), .dout(n1985));
  jand g01622(.dina(n1985), .dinb(n1984), .dout(n1986));
  jor  g01623(.dina(n1986), .dinb(n20391), .dout(n1987));
  jxor g01624(.dina(n1968), .dinb(n348), .dout(n1988));
  jand g01625(.dina(n1988), .dinb(n1987), .dout(n1989));
  jor  g01626(.dina(n1989), .dinb(n1969), .dout(n1990));
  jxor g01627(.dina(n1963), .dinb(n344), .dout(n1991));
  jand g01628(.dina(n1991), .dinb(n1990), .dout(n1992));
  jor  g01629(.dina(n1992), .dinb(n1964), .dout(n1993));
  jxor g01630(.dina(n1958), .dinb(n337), .dout(n1994));
  jand g01631(.dina(n1994), .dinb(n1993), .dout(n1995));
  jor  g01632(.dina(n1995), .dinb(n1959), .dout(n1996));
  jxor g01633(.dina(n1953), .dinb(n338), .dout(n1997));
  jand g01634(.dina(n1997), .dinb(n1996), .dout(n1998));
  jor  g01635(.dina(n1998), .dinb(n1954), .dout(n1999));
  jxor g01636(.dina(n1948), .dinb(n334), .dout(n2000));
  jand g01637(.dina(n2000), .dinb(n1999), .dout(n2001));
  jor  g01638(.dina(n2001), .dinb(n1949), .dout(n2002));
  jxor g01639(.dina(n1943), .dinb(n335), .dout(n2003));
  jand g01640(.dina(n2003), .dinb(n2002), .dout(n2004));
  jor  g01641(.dina(n2004), .dinb(n1944), .dout(n2005));
  jxor g01642(.dina(n1938), .dinb(n323), .dout(n2006));
  jand g01643(.dina(n2006), .dinb(n2005), .dout(n2007));
  jor  g01644(.dina(n2007), .dinb(n1939), .dout(n2008));
  jxor g01645(.dina(n1933), .dinb(n324), .dout(n2009));
  jand g01646(.dina(n2009), .dinb(n2008), .dout(n2010));
  jor  g01647(.dina(n2010), .dinb(n1934), .dout(n2011));
  jxor g01648(.dina(n1928), .dinb(n325), .dout(n2012));
  jand g01649(.dina(n2012), .dinb(n2011), .dout(n2013));
  jor  g01650(.dina(n2013), .dinb(n1929), .dout(n2014));
  jxor g01651(.dina(n1923), .dinb(n439), .dout(n2015));
  jand g01652(.dina(n2015), .dinb(n2014), .dout(n2016));
  jor  g01653(.dina(n2016), .dinb(n1924), .dout(n2017));
  jxor g01654(.dina(n1918), .dinb(n440), .dout(n2018));
  jand g01655(.dina(n2018), .dinb(n2017), .dout(n2019));
  jor  g01656(.dina(n2019), .dinb(n1919), .dout(n2020));
  jxor g01657(.dina(n1913), .dinb(n435), .dout(n2021));
  jand g01658(.dina(n2021), .dinb(n2020), .dout(n2022));
  jor  g01659(.dina(n2022), .dinb(n1914), .dout(n2023));
  jxor g01660(.dina(n1908), .dinb(n436), .dout(n2024));
  jand g01661(.dina(n2024), .dinb(n2023), .dout(n2025));
  jor  g01662(.dina(n2025), .dinb(n1909), .dout(n2026));
  jxor g01663(.dina(n1891), .dinb(n432), .dout(n2027));
  jand g01664(.dina(n2027), .dinb(n2026), .dout(n2028));
  jor  g01665(.dina(n2028), .dinb(n1904), .dout(n2029));
  jxor g01666(.dina(n1902), .dinb(n433), .dout(n2030));
  jand g01667(.dina(n2030), .dinb(n2029), .dout(n2031));
  jor  g01668(.dina(n2031), .dinb(n1903), .dout(n2032));
  jxor g01669(.dina(n1895), .dinb(b17 ), .dout(n2033));
  jor  g01670(.dina(n20497), .dinb(n1896), .dout(quotient46 ));
  jxor g01671(.dina(n2027), .dinb(n2026), .dout(n2040));
  jnot g01672(.din(n1896), .dout(n2045));
  jxor g01673(.dina(n2030), .dinb(n2029), .dout(n2054));
  jxor g01674(.dina(n2024), .dinb(n2023), .dout(n2060));
  jxor g01675(.dina(n2021), .dinb(n2020), .dout(n2065));
  jxor g01676(.dina(n2018), .dinb(n2017), .dout(n2070));
  jxor g01677(.dina(n2015), .dinb(n2014), .dout(n2075));
  jxor g01678(.dina(n2012), .dinb(n2011), .dout(n2080));
  jxor g01679(.dina(n2009), .dinb(n2008), .dout(n2085));
  jxor g01680(.dina(n2006), .dinb(n2005), .dout(n2090));
  jxor g01681(.dina(n2003), .dinb(n2002), .dout(n2095));
  jxor g01682(.dina(n2000), .dinb(n1999), .dout(n2100));
  jxor g01683(.dina(n1997), .dinb(n1996), .dout(n2105));
  jxor g01684(.dina(n1994), .dinb(n1993), .dout(n2110));
  jxor g01685(.dina(n1991), .dinb(n1990), .dout(n2115));
  jxor g01686(.dina(n1988), .dinb(n1987), .dout(n2120));
  jxor g01687(.dina(n1985), .dinb(n1984), .dout(n2125));
  jand g01688(.dina(quotient46 ), .dinb(n1983), .dout(n2133));
  jnot g01689(.din(a45 ), .dout(n2138));
  jand g01690(.dina(b0 ), .dinb(n2138), .dout(n2139));
  jnot g01691(.din(n2139), .dout(n2140));
  jand g01692(.dina(n429), .dinb(n403), .dout(n2196));
  jand g01693(.dina(n2196), .dinb(n420), .dout(n2197));
  jand g01694(.dina(n2197), .dinb(n20650), .dout(quotient45 ));
  jand g01695(.dina(n20652), .dinb(n20587), .dout(n2280));
  jand g01696(.dina(n20751), .dinb(quotient45 ), .dout(n2282));
  jor  g01697(.dina(n2282), .dinb(n2280), .dout(n2283));
  jand g01698(.dina(n2283), .dinb(n344), .dout(n2284));
  jand g01699(.dina(n20652), .dinb(n20593), .dout(n2285));
  jor  g01700(.dina(n20758), .dinb(n2285), .dout(n2288));
  jand g01701(.dina(n2288), .dinb(n348), .dout(n2289));
  jand g01702(.dina(n2197), .dinb(n2139), .dout(n2292));
  jand g01703(.dina(n2292), .dinb(n20650), .dout(n2293));
  jnot g01704(.din(a44 ), .dout(n2298));
  jand g01705(.dina(b0 ), .dinb(n2298), .dout(n2299));
  jnot g01706(.din(n2299), .dout(n2300));
  jand g01707(.dina(n20968), .dinb(n1970), .dout(quotient44 ));
  jand g01708(.dina(n20913), .dinb(n2283), .dout(n2442));
  jor  g01709(.dina(n21061), .dinb(n2442), .dout(n2445));
  jand g01710(.dina(n2445), .dinb(n337), .dout(n2446));
  jand g01711(.dina(n2196), .dinb(n415), .dout(n2457));
  jnot g01712(.din(n315), .dout(n2458));
  jand g01713(.dina(n407), .dinb(b0 ), .dout(n2459));
  jand g01714(.dina(n2459), .dinb(n2458), .dout(n2460));
  jand g01715(.dina(n2460), .dinb(n2457), .dout(n2461));
  jor  g01716(.dina(n21091), .dinb(b1 ), .dout(n2468));
  jnot g01717(.din(a43 ), .dout(n2470));
  jand g01718(.dina(b0 ), .dinb(n2470), .dout(n2471));
  jnot g01719(.din(n2471), .dout(n2472));
  jor  g01720(.dina(n21212), .dinb(n21213), .dout(quotient43 ));
  jnot g01721(.din(b21 ), .dout(n2547));
  jnot g01722(.din(a42 ), .dout(n2649));
  jand g01723(.dina(b0 ), .dinb(n2649), .dout(n2650));
  jnot g01724(.din(n2650), .dout(n2651));
  jnot g01725(.din(b22 ), .dout(n2714));
  jor  g01726(.dina(n310), .dinb(n306), .dout(n2715));
  jor  g01727(.dina(n2715), .dinb(n311), .dout(n2716));
  jor  g01728(.dina(n309), .dinb(b23 ), .dout(n2717));
  jor  g01729(.dina(n2717), .dinb(n2716), .dout(n2718));
  jnot g01730(.din(n2718), .dout(n2719));
  jand g01731(.dina(n2719), .dinb(n2714), .dout(n2720));
  jand g01732(.dina(n2720), .dinb(n21389), .dout(quotient42 ));
  jand g01733(.dina(n2714), .dinb(b0 ), .dout(n2851));
  jand g01734(.dina(n2851), .dinb(n2719), .dout(n2852));
  jand g01735(.dina(n2720), .dinb(n2650), .dout(n2855));
  jnot g01736(.din(a41 ), .dout(n2860));
  jand g01737(.dina(b0 ), .dinb(n2860), .dout(n2861));
  jnot g01738(.din(n21694), .dout(quotient41 ));
  jnot g01739(.din(n2861), .dout(n2953));
  jand g01740(.dina(n2719), .dinb(b0 ), .dout(n3111));
  jnot g01741(.din(a40 ), .dout(n3118));
  jand g01742(.dina(b0 ), .dinb(n3118), .dout(n3119));
  jnot g01743(.din(n3119), .dout(n3120));
  jor  g01744(.dina(n22045), .dinb(n21751), .dout(quotient40 ));
  jnot g01745(.din(a39 ), .dout(n3320));
  jand g01746(.dina(b0 ), .dinb(n3320), .dout(n3321));
  jnot g01747(.din(n3321), .dout(n3322));
  jand g01748(.dina(n22237), .dinb(n2457), .dout(quotient39 ));
  jnot g01749(.din(n307), .dout(n3400));
  jnot g01750(.din(n2716), .dout(n3401));
  jand g01751(.dina(n3401), .dinb(n3400), .dout(n3402));
  jnot g01752(.din(n3402), .dout(n3403));
  jand g01753(.dina(n412), .dinb(b0 ), .dout(n3544));
  jand g01754(.dina(n3544), .dinb(n3402), .dout(n3545));
  jand g01755(.dina(n3321), .dinb(n2457), .dout(n3548));
  jnot g01756(.din(a38 ), .dout(n3553));
  jand g01757(.dina(b0 ), .dinb(n3553), .dout(n3554));
  jnot g01758(.din(n22584), .dout(quotient38 ));
  jnot g01759(.din(n3554), .dout(n3658));
  jand g01760(.dina(n2196), .dinb(n411), .dout(n3716));
  jand g01761(.dina(n2196), .dinb(b0 ), .dout(n3838));
  jand g01762(.dina(n3838), .dinb(n410), .dout(n3839));
  jand g01763(.dina(n3839), .dinb(n3400), .dout(n3840));
  jnot g01764(.din(a37 ), .dout(n3847));
  jand g01765(.dina(b0 ), .dinb(n3847), .dout(n3848));
  jnot g01766(.din(n3848), .dout(n3849));
  jor  g01767(.dina(n22967), .dinb(n22968), .dout(quotient37 ));
  jnot g01768(.din(a36 ), .dout(n4073));
  jand g01769(.dina(b0 ), .dinb(n4073), .dout(n4074));
  jnot g01770(.din(n4074), .dout(n4075));
  jand g01771(.dina(n23192), .dinb(n3401), .dout(quotient36 ));
  jand g01772(.dina(n4074), .dinb(n3401), .dout(n4295));
  jnot g01773(.din(a35 ), .dout(n4301));
  jand g01774(.dina(b0 ), .dinb(n4301), .dout(n4302));
  jnot g01775(.din(n4302), .dout(n4303));
  jand g01776(.dina(n23538), .dinb(n2196), .dout(quotient35 ));
  jand g01777(.dina(n589), .dinb(b0 ), .dout(n4533));
  jand g01778(.dina(n304), .dinb(n424), .dout(n4534));
  jand g01779(.dina(n4534), .dinb(n4533), .dout(n4535));
  jand g01780(.dina(n4535), .dinb(n428), .dout(n4536));
  jand g01781(.dina(n3838), .dinb(n4301), .dout(n4539));
  jnot g01782(.din(a34 ), .dout(n4545));
  jand g01783(.dina(b0 ), .dinb(n4545), .dout(n4546));
  jnot g01784(.din(n4546), .dout(n4547));
  jor  g01785(.dina(n24007), .dinb(n24008), .dout(quotient34 ));
  jand g01786(.dina(n403), .dinb(n425), .dout(n4642));
  jnot g01787(.din(a33 ), .dout(n4798));
  jand g01788(.dina(b0 ), .dinb(n4798), .dout(n4799));
  jnot g01789(.din(n4799), .dout(n4800));
  jand g01790(.dina(n24256), .dinb(n4642), .dout(quotient33 ));
  jand g01791(.dina(n4799), .dinb(n4642), .dout(n5046));
  jnot g01792(.din(a32 ), .dout(n5052));
  jand g01793(.dina(b0 ), .dinb(n5052), .dout(n5053));
  jnot g01794(.din(n5053), .dout(n5054));
  jand g01795(.dina(n24638), .dinb(n590), .dout(quotient32 ));
  jand g01796(.dina(n300), .dinb(b0 ), .dout(n5307));
  jand g01797(.dina(n5307), .dinb(n403), .dout(n5308));
  jand g01798(.dina(n5053), .dinb(n590), .dout(n5311));
  jnot g01799(.din(a31 ), .dout(n5317));
  jand g01800(.dina(b0 ), .dinb(n5317), .dout(n5318));
  jnot g01801(.din(n5318), .dout(n5319));
  jor  g01802(.dina(n25167), .dinb(n24645), .dout(quotient31 ));
  jnot g01803(.din(a30 ), .dout(n5591));
  jand g01804(.dina(b0 ), .dinb(n5591), .dout(n5592));
  jnot g01805(.din(n5592), .dout(n5593));
  jand g01806(.dina(n296), .dinb(n301), .dout(n5692));
  jand g01807(.dina(n5692), .dinb(n298), .dout(n5693));
  jand g01808(.dina(n5693), .dinb(n589), .dout(n5694));
  jand g01809(.dina(n5694), .dinb(n25431), .dout(quotient30 ));
  jand g01810(.dina(n518), .dinb(n391), .dout(n5701));
  jand g01811(.dina(n5701), .dinb(n389), .dout(n5702));
  jand g01812(.dina(n5702), .dinb(n388), .dout(n5703));
  jnot g01813(.din(n5703), .dout(n5704));
  jand g01814(.dina(n298), .dinb(b0 ), .dout(n5899));
  jand g01815(.dina(n5899), .dinb(n5703), .dout(n5900));
  jand g01816(.dina(n5694), .dinb(n5592), .dout(n5903));
  jnot g01817(.din(a29 ), .dout(n5908));
  jand g01818(.dina(b0 ), .dinb(n5908), .dout(n5909));
  jnot g01819(.din(n25904), .dout(quotient29 ));
  jnot g01820(.din(n5909), .dout(n6049));
  jand g01821(.dina(n5692), .dinb(n4533), .dout(n6286));
  jnot g01822(.din(a28 ), .dout(n6293));
  jand g01823(.dina(b0 ), .dinb(n6293), .dout(n6294));
  jnot g01824(.din(n6294), .dout(n6295));
  jand g01825(.dina(n296), .dinb(n589), .dout(n6403));
  jnot g01826(.din(n6403), .dout(n6404));
  jor  g01827(.dina(n26413), .dinb(n26412), .dout(quotient28 ));
  jnot g01828(.din(a27 ), .dout(n6599));
  jand g01829(.dina(b0 ), .dinb(n6599), .dout(n6600));
  jnot g01830(.din(n6600), .dout(n6601));
  jand g01831(.dina(n26709), .dinb(n5702), .dout(quotient27 ));
  jand g01832(.dina(n292), .dinb(n589), .dout(n6715));
  jnot g01833(.din(n6715), .dout(n6716));
  jand g01834(.dina(n292), .dinb(n294), .dout(n6929));
  jand g01835(.dina(n6929), .dinb(n4533), .dout(n6930));
  jand g01836(.dina(n6600), .dinb(n5702), .dout(n6933));
  jnot g01837(.din(a26 ), .dout(n6938));
  jand g01838(.dina(b0 ), .dinb(n6938), .dout(n6939));
  jnot g01839(.din(n27224), .dout(quotient26 ));
  jnot g01840(.din(n6939), .dout(n7091));
  jand g01841(.dina(n284), .dinb(b0 ), .dout(n7354));
  jand g01842(.dina(n7354), .dinb(n518), .dout(n7355));
  jand g01843(.dina(n7355), .dinb(n292), .dout(n7356));
  jnot g01844(.din(a25 ), .dout(n7363));
  jand g01845(.dina(b0 ), .dinb(n7363), .dout(n7364));
  jnot g01846(.din(n7364), .dout(n7365));
  jor  g01847(.dina(n27775), .dinb(n27776), .dout(quotient25 ));
  jnot g01848(.din(a24 ), .dout(n7722));
  jand g01849(.dina(b0 ), .dinb(n7722), .dout(n7723));
  jnot g01850(.din(n28167), .dout(quotient24 ));
  jnot g01851(.din(n7723), .dout(n7883));
  jnot g01852(.din(n518), .dout(n7960));
  jnot g01853(.din(a23 ), .dout(n8203));
  jand g01854(.dina(b0 ), .dinb(n8203), .dout(n8204));
  jnot g01855(.din(n28653), .dout(quotient23 ));
  jnot g01856(.din(n8204), .dout(n8369));
  jand g01857(.dina(n283), .dinb(n588), .dout(n8458));
  jand g01858(.dina(n282), .dinb(b0 ), .dout(n8658));
  jand g01859(.dina(n8658), .dinb(n588), .dout(n8659));
  jand g01860(.dina(n8659), .dinb(n395), .dout(n8660));
  jnot g01861(.din(a22 ), .dout(n8667));
  jand g01862(.dina(b0 ), .dinb(n8667), .dout(n8668));
  jnot g01863(.din(n8668), .dout(n8669));
  jor  g01864(.dina(n29245), .dinb(n29246), .dout(quotient22 ));
  jnot g01865(.din(a21 ), .dout(n9015));
  jand g01866(.dina(b0 ), .dinb(n9015), .dout(n9016));
  jnot g01867(.din(n9016), .dout(n9017));
  jand g01868(.dina(n29590), .dinb(n517), .dout(quotient21 ));
  jand g01869(.dina(n9016), .dinb(n517), .dout(n9354));
  jnot g01870(.din(a20 ), .dout(n9360));
  jand g01871(.dina(b0 ), .dinb(n9360), .dout(n9361));
  jnot g01872(.din(n9361), .dout(n9362));
  jor  g01873(.dina(n29597), .dinb(n30294), .dout(quotient20 ));
  jnot g01874(.din(a19 ), .dout(n9719));
  jand g01875(.dina(b0 ), .dinb(n9719), .dout(n9720));
  jnot g01876(.din(n9720), .dout(n9721));
  jor  g01877(.dina(n30823), .dinb(n30821), .dout(quotient19 ));
  jnot g01878(.din(n273), .dout(n9866));
  jand g01879(.dina(n382), .dinb(n583), .dout(n9867));
  jand g01880(.dina(n9867), .dinb(n584), .dout(n9868));
  jand g01881(.dina(n9868), .dinb(n9866), .dout(n9869));
  jnot g01882(.din(a18 ), .dout(n10100));
  jand g01883(.dina(b0 ), .dinb(n10100), .dout(n10101));
  jnot g01884(.din(n10101), .dout(n10102));
  jand g01885(.dina(n31190), .dinb(n9869), .dout(quotient18 ));
  jand g01886(.dina(n514), .dinb(b0 ), .dout(n10459));
  jand g01887(.dina(n10459), .dinb(n512), .dout(n10460));
  jand g01888(.dina(n10101), .dinb(n9869), .dout(n10463));
  jnot g01889(.din(a17 ), .dout(n10469));
  jand g01890(.dina(b0 ), .dinb(n10469), .dout(n10470));
  jnot g01891(.din(n10470), .dout(n10471));
  jnot g01892(.din(n512), .dout(n10607));
  jor  g01893(.dina(n31197), .dinb(n31946), .dout(quotient17 ));
  jnot g01894(.din(a16 ), .dout(n10853));
  jand g01895(.dina(b0 ), .dinb(n10853), .dout(n10854));
  jnot g01896(.din(n10854), .dout(n10855));
  jor  g01897(.dina(n31942), .dinb(n32518), .dout(quotient16 ));
  jnot g01898(.din(a15 ), .dout(n11254));
  jand g01899(.dina(b0 ), .dinb(n11254), .dout(n11255));
  jnot g01900(.din(n11255), .dout(n11256));
  jand g01901(.dina(n32902), .dinb(n387), .dout(quotient15 ));
  jand g01902(.dina(n383), .dinb(b0 ), .dout(n11637));
  jand g01903(.dina(n11637), .dinb(n9867), .dout(n11638));
  jand g01904(.dina(n11255), .dinb(n387), .dout(n11641));
  jnot g01905(.din(a14 ), .dout(n11647));
  jand g01906(.dina(b0 ), .dinb(n11647), .dout(n11648));
  jnot g01907(.din(n11648), .dout(n11649));
  jnot g01908(.din(n9867), .dout(n11794));
  jor  g01909(.dina(n33694), .dinb(n33693), .dout(quotient14 ));
  jnot g01910(.din(a13 ), .dout(n12061));
  jand g01911(.dina(b0 ), .dinb(n12061), .dout(n12062));
  jnot g01912(.din(n12062), .dout(n12063));
  jnot g01913(.din(b50 ), .dout(n12211));
  jnot g01914(.din(b51 ), .dout(n12214));
  jand g01915(.dina(n384), .dinb(n12214), .dout(n12215));
  jand g01916(.dina(n12215), .dinb(n381), .dout(n12216));
  jor  g01917(.dina(n34298), .dinb(n34300), .dout(quotient13 ));
  jnot g01918(.din(a12 ), .dout(n12485));
  jand g01919(.dina(b0 ), .dinb(n12485), .dout(n12486));
  jnot g01920(.din(n12486), .dout(n12487));
  jand g01921(.dina(n34715), .dinb(n583), .dout(quotient12 ));
  jand g01922(.dina(n384), .dinb(b0 ), .dout(n12894));
  jand g01923(.dina(n12894), .dinb(n381), .dout(n12895));
  jand g01924(.dina(n12486), .dinb(n583), .dout(n12898));
  jnot g01925(.din(a11 ), .dout(n12904));
  jand g01926(.dina(b0 ), .dinb(n12904), .dout(n12905));
  jnot g01927(.din(n12905), .dout(n12906));
  jnot g01928(.din(n381), .dout(n13060));
  jor  g01929(.dina(n35555), .dinb(n35554), .dout(quotient11 ));
  jand g01930(.dina(n35560), .dinb(n381), .dout(n13081));
  jnot g01931(.din(a10 ), .dout(n13342));
  jand g01932(.dina(b0 ), .dinb(n13342), .dout(n13343));
  jnot g01933(.din(n13343), .dout(n13344));
  jxor g01934(.dina(n35560), .dinb(n374), .dout(n13501));
  jand g01935(.dina(n13501), .dinb(n35982), .dout(n13502));
  jand g01936(.dina(n379), .dinb(n373), .dout(n13503));
  jand g01937(.dina(n13503), .dinb(n13502), .dout(n13504));
  jor  g01938(.dina(n13504), .dinb(n13081), .dout(quotient10 ));
  jnot g01939(.din(a9 ), .dout(n13837));
  jand g01940(.dina(b0 ), .dinb(n13837), .dout(n13838));
  jand g01941(.dina(n373), .dinb(n375), .dout(n14053));
  jand g01942(.dina(n14053), .dinb(n377), .dout(n14054));
  jnot g01943(.din(n14054), .dout(n14055));
  jnot g01944(.din(n36745), .dout(quotient9 ));
  jnot g01945(.din(n13838), .dout(n14061));
  jand g01946(.dina(n14054), .dinb(b0 ), .dout(n14440));
  jnot g01947(.din(a8 ), .dout(n14447));
  jand g01948(.dina(b0 ), .dinb(n14447), .dout(n14448));
  jnot g01949(.din(n14448), .dout(n14449));
  jnot g01950(.din(n14053), .dout(n14612));
  jor  g01951(.dina(n37519), .dinb(n37524), .dout(quotient8 ));
  jnot g01952(.din(a7 ), .dout(n14903));
  jand g01953(.dina(b0 ), .dinb(n14903), .dout(n14904));
  jnot g01954(.din(n14904), .dout(n14905));
  jor  g01955(.dina(n38197), .dinb(n38196), .dout(quotient7 ));
  jand g01956(.dina(n372), .dinb(n363), .dout(n15090));
  jnot g01957(.din(a6 ), .dout(n15381));
  jand g01958(.dina(b0 ), .dinb(n15381), .dout(n15382));
  jnot g01959(.din(n15382), .dout(n15383));
  jand g01960(.dina(n38894), .dinb(n15090), .dout(quotient6 ));
  jand g01961(.dina(n15090), .dinb(b0 ), .dout(n15840));
  jnot g01962(.din(a5 ), .dout(n15845));
  jand g01963(.dina(b0 ), .dinb(n15845), .dout(n15846));
  jnot g01964(.din(n15846), .dout(n15847));
  jnot g01965(.din(n372), .dout(n16024));
  jand g01966(.dina(n39592), .dinb(n39591), .dout(quotient5 ));
  jnot g01967(.din(a4 ), .dout(n16325));
  jand g01968(.dina(b0 ), .dinb(n16325), .dout(n16326));
  jnot g01969(.din(n16326), .dout(n16327));
  jand g01970(.dina(n40305), .dinb(n40304), .dout(quotient4 ));
  jnot g01971(.din(a3 ), .dout(n16812));
  jand g01972(.dina(b0 ), .dinb(n16812), .dout(n16813));
  jnot g01973(.din(n16813), .dout(n16814));
  jand g01974(.dina(n41030), .dinb(n41029), .dout(quotient3 ));
  jnot g01975(.din(a2 ), .dout(n17307));
  jand g01976(.dina(b0 ), .dinb(n17307), .dout(n17308));
  jnot g01977(.din(n17308), .dout(n17309));
  jand g01978(.dina(n41769), .dinb(n41768), .dout(quotient2 ));
  jnot g01979(.din(a1 ), .dout(n17810));
  jand g01980(.dina(b0 ), .dinb(n17810), .dout(n17811));
  jnot g01981(.din(n17811), .dout(n17812));
  jand g01982(.dina(n42519), .dinb(n42518), .dout(quotient1 ));
  jor  g01983(.dina(n42529), .dinb(n256), .dout(n18009));
  jnot g01984(.din(b0 ), .dout(n18364));
  jor  g01985(.dina(n18364), .dinb(a0 ), .dout(n18365));
  jand g01986(.dina(n43266), .dinb(n18009), .dout(n18490));
  jor  g01987(.dina(n42524), .dinb(n42530), .dout(n18497));
  jor  g01988(.dina(n18497), .dinb(n18490), .dout(n18498));
  jor  g01989(.dina(n42523), .dinb(n367), .dout(n18499));
  jand g01990(.dina(n43143), .dinb(n18499), .dout(n18501));
  jand g01991(.dina(n18501), .dinb(n18498), .dout(n18502));
  jor  g01992(.dina(n42515), .dinb(n18502), .dout(quotient0 ));
  jnot g01993(.din(n622), .dout(quotient59 ));
  jand g01994(.dina(n496), .dinb(n493), .dout(quotient61 ));
  jand g01995(.dina(n476), .dinb(n360), .dout(quotient62 ));
  jand g01996(.dina(n494), .dinb(n352), .dout(n18511));
  jand g01997(.dina(n18511), .dinb(n556), .dout(quotient63 ));
  jand g01998(.dina(n544), .dinb(n500), .dout(n18568));
  jnot g01999(.din(n530), .dout(n18575));
  jnot g02000(.din(n559), .dout(n18577));
  jand g02001(.dina(n18577), .dinb(n18568), .dout(n18578));
  jor  g02002(.dina(n18578), .dinb(n18575), .dout(n18579));
  jand g02003(.dina(n567), .dinb(n18579), .dout(n18592));
  jnot g02004(.din(n18592), .dout(n18593));
  jand g02005(.dina(n18592), .dinb(b3 ), .dout(n18596));
  jnot g02006(.din(n650), .dout(n18651));
  jor  g02007(.dina(n18651), .dinb(n645), .dout(n18652));
  jand g02008(.dina(n18652), .dinb(n337), .dout(n18653));
  jor  g02009(.dina(n689), .dinb(n638), .dout(n18720));
  jand g02010(.dina(n691), .dinb(n670), .dout(n18735));
  jand g02011(.dina(n719), .dinb(n18720), .dout(n18737));
  jor  g02012(.dina(n18737), .dinb(n18735), .dout(n18738));
  jand g02013(.dina(n18738), .dinb(n348), .dout(n18739));
  jand g02014(.dina(n751), .dinb(n555), .dout(n18768));
  jor  g02015(.dina(n18768), .dinb(n729), .dout(n18798));
  jnot g02016(.din(n781), .dout(n18801));
  jand g02017(.dina(n18801), .dinb(n18798), .dout(n18802));
  jor  g02018(.dina(n18802), .dinb(b2 ), .dout(n18803));
  jnot g02019(.din(n858), .dout(n18911));
  jnot g02020(.din(n762), .dout(n18912));
  jnot g02021(.din(n767), .dout(n18913));
  jnot g02022(.din(n768), .dout(n18914));
  jnot g02023(.din(n773), .dout(n18915));
  jnot g02024(.din(n778), .dout(n18916));
  jnot g02025(.din(n791), .dout(n18917));
  jxor g02026(.dina(n789), .dinb(n258), .dout(n18918));
  jor  g02027(.dina(n18918), .dinb(n793), .dout(n18919));
  jand g02028(.dina(n18919), .dinb(n18917), .dout(n18920));
  jnot g02029(.din(n798), .dout(n18921));
  jor  g02030(.dina(n18921), .dinb(n18920), .dout(n18922));
  jand g02031(.dina(n18922), .dinb(n18803), .dout(n18923));
  jnot g02032(.din(n801), .dout(n18924));
  jor  g02033(.dina(n18924), .dinb(n18923), .dout(n18925));
  jand g02034(.dina(n18925), .dinb(n18916), .dout(n18926));
  jnot g02035(.din(n804), .dout(n18927));
  jor  g02036(.dina(n18927), .dinb(n18926), .dout(n18928));
  jand g02037(.dina(n18928), .dinb(n18915), .dout(n18929));
  jnot g02038(.din(n807), .dout(n18930));
  jor  g02039(.dina(n18930), .dinb(n18929), .dout(n18931));
  jand g02040(.dina(n18931), .dinb(n18914), .dout(n18932));
  jnot g02041(.din(n810), .dout(n18933));
  jor  g02042(.dina(n18933), .dinb(n18932), .dout(n18934));
  jand g02043(.dina(n18934), .dinb(n18913), .dout(n18935));
  jor  g02044(.dina(n814), .dinb(n18935), .dout(n18936));
  jand g02045(.dina(n18936), .dinb(n18912), .dout(n18937));
  jor  g02046(.dina(n18937), .dinb(n18911), .dout(n18938));
  jand g02047(.dina(n18938), .dinb(a56 ), .dout(n18939));
  jor  g02048(.dina(n862), .dinb(n18939), .dout(n18943));
  jor  g02049(.dina(n894), .dinb(n828), .dout(n19007));
  jand g02050(.dina(n896), .dinb(n18943), .dout(n19037));
  jand g02051(.dina(n936), .dinb(n19007), .dout(n19039));
  jor  g02052(.dina(n19039), .dinb(n19037), .dout(n19040));
  jand g02053(.dina(n19040), .dinb(n348), .dout(n19041));
  jnot g02054(.din(n908), .dout(n19139));
  jnot g02055(.din(n913), .dout(n19140));
  jnot g02056(.din(n914), .dout(n19141));
  jnot g02057(.din(n919), .dout(n19142));
  jnot g02058(.din(n924), .dout(n19143));
  jnot g02059(.din(n929), .dout(n19144));
  jnot g02060(.din(n934), .dout(n19145));
  jnot g02061(.din(n19041), .dout(n19146));
  jnot g02062(.din(n948), .dout(n19147));
  jxor g02063(.dina(n946), .dinb(n258), .dout(n19148));
  jor  g02064(.dina(n19148), .dinb(n950), .dout(n19149));
  jand g02065(.dina(n19149), .dinb(n19147), .dout(n19150));
  jnot g02066(.din(n955), .dout(n19151));
  jor  g02067(.dina(n19151), .dinb(n19150), .dout(n19152));
  jand g02068(.dina(n19152), .dinb(n19146), .dout(n19153));
  jnot g02069(.din(n958), .dout(n19154));
  jor  g02070(.dina(n19154), .dinb(n19153), .dout(n19155));
  jand g02071(.dina(n19155), .dinb(n19145), .dout(n19156));
  jnot g02072(.din(n961), .dout(n19157));
  jor  g02073(.dina(n19157), .dinb(n19156), .dout(n19158));
  jand g02074(.dina(n19158), .dinb(n19144), .dout(n19159));
  jnot g02075(.din(n964), .dout(n19160));
  jor  g02076(.dina(n19160), .dinb(n19159), .dout(n19161));
  jand g02077(.dina(n19161), .dinb(n19143), .dout(n19162));
  jnot g02078(.din(n967), .dout(n19163));
  jor  g02079(.dina(n19163), .dinb(n19162), .dout(n19164));
  jand g02080(.dina(n19164), .dinb(n19142), .dout(n19165));
  jnot g02081(.din(n970), .dout(n19166));
  jor  g02082(.dina(n19166), .dinb(n19165), .dout(n19167));
  jand g02083(.dina(n19167), .dinb(n19141), .dout(n19168));
  jnot g02084(.din(n973), .dout(n19169));
  jor  g02085(.dina(n19169), .dinb(n19168), .dout(n19170));
  jand g02086(.dina(n19170), .dinb(n19140), .dout(n19171));
  jor  g02087(.dina(n906), .dinb(n19171), .dout(n19172));
  jand g02088(.dina(n19172), .dinb(n19139), .dout(n19173));
  jnot g02089(.din(n1043), .dout(n19219));
  jor  g02090(.dina(n19173), .dinb(n19219), .dout(n19220));
  jand g02091(.dina(n19220), .dinb(a54 ), .dout(n19221));
  jor  g02092(.dina(n1047), .dinb(n19221), .dout(n19223));
  jand g02093(.dina(n1169), .dinb(n990), .dout(n19255));
  jand g02094(.dina(n1092), .dinb(n19223), .dout(n19307));
  jor  g02095(.dina(n1162), .dinb(n19307), .dout(n19310));
  jand g02096(.dina(n19310), .dinb(n348), .dout(n19311));
  jnot g02097(.din(n1171), .dout(n19313));
  jor  g02098(.dina(n1091), .dinb(n19313), .dout(n19314));
  jand g02099(.dina(n19314), .dinb(a53 ), .dout(n19315));
  jand g02100(.dina(n19255), .dinb(n1052), .dout(n19316));
  jor  g02101(.dina(n19316), .dinb(n19315), .dout(n19317));
  jxor g02102(.dina(n19310), .dinb(n348), .dout(n19327));
  jor  g02103(.dina(n1215), .dinb(n1123), .dout(n19400));
  jand g02104(.dina(n1217), .dinb(n19317), .dout(n19445));
  jand g02105(.dina(n1272), .dinb(n19400), .dout(n19447));
  jor  g02106(.dina(n19447), .dinb(n19445), .dout(n19448));
  jand g02107(.dina(n19448), .dinb(n348), .dout(n19449));
  jnot g02108(.din(n1229), .dout(n19574));
  jnot g02109(.din(n1234), .dout(n19575));
  jnot g02110(.din(n1235), .dout(n19576));
  jnot g02111(.din(n1240), .dout(n19577));
  jnot g02112(.din(n1245), .dout(n19578));
  jnot g02113(.din(n1250), .dout(n19579));
  jnot g02114(.din(n1255), .dout(n19580));
  jnot g02115(.din(n1260), .dout(n19581));
  jnot g02116(.din(n1265), .dout(n19582));
  jnot g02117(.din(n1270), .dout(n19583));
  jnot g02118(.din(n19449), .dout(n19584));
  jnot g02119(.din(n1284), .dout(n19585));
  jxor g02120(.dina(n1282), .dinb(n258), .dout(n19586));
  jor  g02121(.dina(n19586), .dinb(n1286), .dout(n19587));
  jand g02122(.dina(n19587), .dinb(n19585), .dout(n19588));
  jnot g02123(.din(n1291), .dout(n19589));
  jor  g02124(.dina(n19589), .dinb(n19588), .dout(n19590));
  jand g02125(.dina(n19590), .dinb(n19584), .dout(n19591));
  jnot g02126(.din(n1294), .dout(n19592));
  jor  g02127(.dina(n19592), .dinb(n19591), .dout(n19593));
  jand g02128(.dina(n19593), .dinb(n19583), .dout(n19594));
  jnot g02129(.din(n1297), .dout(n19595));
  jor  g02130(.dina(n19595), .dinb(n19594), .dout(n19596));
  jand g02131(.dina(n19596), .dinb(n19582), .dout(n19597));
  jnot g02132(.din(n1300), .dout(n19598));
  jor  g02133(.dina(n19598), .dinb(n19597), .dout(n19599));
  jand g02134(.dina(n19599), .dinb(n19581), .dout(n19600));
  jnot g02135(.din(n1303), .dout(n19601));
  jor  g02136(.dina(n19601), .dinb(n19600), .dout(n19602));
  jand g02137(.dina(n19602), .dinb(n19580), .dout(n19603));
  jnot g02138(.din(n1306), .dout(n19604));
  jor  g02139(.dina(n19604), .dinb(n19603), .dout(n19605));
  jand g02140(.dina(n19605), .dinb(n19579), .dout(n19606));
  jnot g02141(.din(n1309), .dout(n19607));
  jor  g02142(.dina(n19607), .dinb(n19606), .dout(n19608));
  jand g02143(.dina(n19608), .dinb(n19578), .dout(n19609));
  jnot g02144(.din(n1312), .dout(n19610));
  jor  g02145(.dina(n19610), .dinb(n19609), .dout(n19611));
  jand g02146(.dina(n19611), .dinb(n19577), .dout(n19612));
  jnot g02147(.din(n1315), .dout(n19613));
  jor  g02148(.dina(n19613), .dinb(n19612), .dout(n19614));
  jand g02149(.dina(n19614), .dinb(n19576), .dout(n19615));
  jnot g02150(.din(n1318), .dout(n19616));
  jor  g02151(.dina(n19616), .dinb(n19615), .dout(n19617));
  jand g02152(.dina(n19617), .dinb(n19575), .dout(n19618));
  jor  g02153(.dina(n1227), .dinb(n19618), .dout(n19619));
  jand g02154(.dina(n19619), .dinb(n19574), .dout(n19620));
  jnot g02155(.din(n1401), .dout(n19678));
  jor  g02156(.dina(n19620), .dinb(n19678), .dout(n19679));
  jand g02157(.dina(n19679), .dinb(a51 ), .dout(n19680));
  jor  g02158(.dina(n1405), .dinb(n19680), .dout(n19682));
  jnot g02159(.din(n1498), .dout(n19713));
  jand g02160(.dina(n1561), .dinb(n1330), .dout(n19718));
  jnot g02161(.din(n1505), .dout(n19723));
  jnot g02162(.din(n1506), .dout(n19729));
  jnot g02163(.din(n1511), .dout(n19735));
  jnot g02164(.din(n1516), .dout(n19741));
  jnot g02165(.din(n1521), .dout(n19747));
  jnot g02166(.din(n1526), .dout(n19753));
  jnot g02167(.din(n1531), .dout(n19759));
  jnot g02168(.din(n1536), .dout(n19765));
  jnot g02169(.din(n1541), .dout(n19771));
  jnot g02170(.din(n1546), .dout(n19779));
  jnot g02171(.din(n1551), .dout(n19787));
  jand g02172(.dina(n1462), .dinb(n19682), .dout(n19788));
  jor  g02173(.dina(n1554), .dinb(n19788), .dout(n19791));
  jand g02174(.dina(n19791), .dinb(n348), .dout(n19792));
  jnot g02175(.din(n19792), .dout(n19793));
  jnot g02176(.din(n1564), .dout(n19794));
  jor  g02177(.dina(n1461), .dinb(n19794), .dout(n19795));
  jand g02178(.dina(n19795), .dinb(a50 ), .dout(n19796));
  jand g02179(.dina(n19718), .dinb(n1410), .dout(n19797));
  jor  g02180(.dina(n19797), .dinb(n19796), .dout(n19798));
  jxor g02181(.dina(n1568), .dinb(n258), .dout(n19805));
  jor  g02182(.dina(n19805), .dinb(n1572), .dout(n19806));
  jand g02183(.dina(n19806), .dinb(n1569), .dout(n19807));
  jxor g02184(.dina(n19791), .dinb(n348), .dout(n19808));
  jnot g02185(.din(n19808), .dout(n19809));
  jor  g02186(.dina(n19809), .dinb(n19807), .dout(n19810));
  jand g02187(.dina(n19810), .dinb(n19793), .dout(n19811));
  jnot g02188(.din(n1580), .dout(n19813));
  jor  g02189(.dina(n19813), .dinb(n19811), .dout(n19814));
  jand g02190(.dina(n19814), .dinb(n19787), .dout(n19815));
  jnot g02191(.din(n1583), .dout(n19817));
  jor  g02192(.dina(n19817), .dinb(n19815), .dout(n19818));
  jand g02193(.dina(n19818), .dinb(n19779), .dout(n19819));
  jnot g02194(.din(n1586), .dout(n19821));
  jor  g02195(.dina(n19821), .dinb(n19819), .dout(n19822));
  jand g02196(.dina(n19822), .dinb(n19771), .dout(n19823));
  jnot g02197(.din(n1589), .dout(n19825));
  jor  g02198(.dina(n19825), .dinb(n19823), .dout(n19826));
  jand g02199(.dina(n19826), .dinb(n19765), .dout(n19827));
  jnot g02200(.din(n1592), .dout(n19829));
  jor  g02201(.dina(n19829), .dinb(n19827), .dout(n19830));
  jand g02202(.dina(n19830), .dinb(n19759), .dout(n19831));
  jnot g02203(.din(n1595), .dout(n19833));
  jor  g02204(.dina(n19833), .dinb(n19831), .dout(n19834));
  jand g02205(.dina(n19834), .dinb(n19753), .dout(n19835));
  jnot g02206(.din(n1598), .dout(n19837));
  jor  g02207(.dina(n19837), .dinb(n19835), .dout(n19838));
  jand g02208(.dina(n19838), .dinb(n19747), .dout(n19839));
  jnot g02209(.din(n1601), .dout(n19841));
  jor  g02210(.dina(n19841), .dinb(n19839), .dout(n19842));
  jand g02211(.dina(n19842), .dinb(n19741), .dout(n19843));
  jnot g02212(.din(n1604), .dout(n19845));
  jor  g02213(.dina(n19845), .dinb(n19843), .dout(n19846));
  jand g02214(.dina(n19846), .dinb(n19735), .dout(n19847));
  jnot g02215(.din(n1607), .dout(n19849));
  jor  g02216(.dina(n19849), .dinb(n19847), .dout(n19850));
  jand g02217(.dina(n19850), .dinb(n19729), .dout(n19851));
  jnot g02218(.din(n1610), .dout(n19853));
  jor  g02219(.dina(n19853), .dinb(n19851), .dout(n19854));
  jand g02220(.dina(n19854), .dinb(n19723), .dout(n19855));
  jnot g02221(.din(n1500), .dout(n19856));
  jor  g02222(.dina(n1613), .dinb(n19856), .dout(n19858));
  jor  g02223(.dina(n19858), .dinb(n19855), .dout(n19859));
  jand g02224(.dina(n19859), .dinb(n19713), .dout(n19860));
  jor  g02225(.dina(n1499), .dinb(n1616), .dout(n19891));
  jxor g02226(.dina(n1613), .dinb(n1612), .dout(n19892));
  jand g02227(.dina(n19892), .dinb(n19891), .dout(n19893));
  jor  g02228(.dina(n19893), .dinb(n19860), .dout(n19894));
  jand g02229(.dina(n19894), .dinb(b15 ), .dout(n19896));
  jnot g02230(.din(n19896), .dout(n19897));
  jnot g02231(.din(n1499), .dout(n19899));
  jand g02232(.dina(n19899), .dinb(n19859), .dout(n19900));
  jand g02233(.dina(n19900), .dinb(n1504), .dout(n19901));
  jor  g02234(.dina(n1633), .dinb(n19901), .dout(n19904));
  jand g02235(.dina(n19904), .dinb(n436), .dout(n19905));
  jand g02236(.dina(n19900), .dinb(n1490), .dout(n19906));
  jor  g02237(.dina(n1621), .dinb(n19906), .dout(n19909));
  jand g02238(.dina(n19909), .dinb(n435), .dout(n19910));
  jand g02239(.dina(n19900), .dinb(n1510), .dout(n19911));
  jor  g02240(.dina(n1639), .dinb(n19911), .dout(n19914));
  jand g02241(.dina(n19914), .dinb(n440), .dout(n19915));
  jand g02242(.dina(n19900), .dinb(n1515), .dout(n19916));
  jor  g02243(.dina(n1644), .dinb(n19916), .dout(n19919));
  jand g02244(.dina(n19919), .dinb(n439), .dout(n19920));
  jand g02245(.dina(n19900), .dinb(n1520), .dout(n19921));
  jor  g02246(.dina(n1649), .dinb(n19921), .dout(n19924));
  jand g02247(.dina(n19924), .dinb(n325), .dout(n19925));
  jand g02248(.dina(n19900), .dinb(n1525), .dout(n19926));
  jor  g02249(.dina(n1654), .dinb(n19926), .dout(n19929));
  jand g02250(.dina(n19929), .dinb(n324), .dout(n19930));
  jand g02251(.dina(n19900), .dinb(n1530), .dout(n19931));
  jor  g02252(.dina(n1659), .dinb(n19931), .dout(n19934));
  jand g02253(.dina(n19934), .dinb(n323), .dout(n19935));
  jand g02254(.dina(n19900), .dinb(n1535), .dout(n19936));
  jor  g02255(.dina(n1664), .dinb(n19936), .dout(n19939));
  jand g02256(.dina(n19939), .dinb(n335), .dout(n19940));
  jand g02257(.dina(n19900), .dinb(n1540), .dout(n19941));
  jor  g02258(.dina(n1669), .dinb(n19941), .dout(n19944));
  jand g02259(.dina(n19944), .dinb(n334), .dout(n19945));
  jand g02260(.dina(n19900), .dinb(n1545), .dout(n19946));
  jor  g02261(.dina(n1674), .dinb(n19946), .dout(n19949));
  jand g02262(.dina(n19949), .dinb(n338), .dout(n19950));
  jand g02263(.dina(n19900), .dinb(n1550), .dout(n19951));
  jor  g02264(.dina(n1679), .dinb(n19951), .dout(n19954));
  jand g02265(.dina(n19954), .dinb(n337), .dout(n19955));
  jand g02266(.dina(n19900), .dinb(n19791), .dout(n19956));
  jor  g02267(.dina(n1684), .dinb(n19956), .dout(n19959));
  jand g02268(.dina(n19959), .dinb(n344), .dout(n19960));
  jand g02269(.dina(n19900), .dinb(n19798), .dout(n19961));
  jand g02270(.dina(n1688), .dinb(n19891), .dout(n19963));
  jor  g02271(.dina(n19963), .dinb(n19961), .dout(n19964));
  jand g02272(.dina(n19964), .dinb(n348), .dout(n19965));
  jor  g02273(.dina(n19900), .dinb(n18364), .dout(n19966));
  jand g02274(.dina(n19966), .dinb(a49 ), .dout(n19967));
  jor  g02275(.dina(n19900), .dinb(n1573), .dout(n19968));
  jor  g02276(.dina(n1696), .dinb(n19967), .dout(n19970));
  jand g02277(.dina(n19970), .dinb(n258), .dout(n19971));
  jxor g02278(.dina(n19964), .dinb(n348), .dout(n19978));
  jxor g02279(.dina(n19959), .dinb(n344), .dout(n19981));
  jxor g02280(.dina(n19954), .dinb(n337), .dout(n19984));
  jxor g02281(.dina(n19949), .dinb(n338), .dout(n19987));
  jxor g02282(.dina(n19944), .dinb(n334), .dout(n19990));
  jxor g02283(.dina(n19939), .dinb(n335), .dout(n19993));
  jxor g02284(.dina(n19934), .dinb(n323), .dout(n19996));
  jxor g02285(.dina(n19929), .dinb(n324), .dout(n19999));
  jxor g02286(.dina(n19924), .dinb(n325), .dout(n20002));
  jxor g02287(.dina(n19919), .dinb(n439), .dout(n20005));
  jxor g02288(.dina(n19914), .dinb(n440), .dout(n20008));
  jxor g02289(.dina(n19909), .dinb(n435), .dout(n20011));
  jxor g02290(.dina(n19904), .dinb(n436), .dout(n20014));
  jand g02291(.dina(n1747), .dinb(n594), .dout(n20019));
  jor  g02292(.dina(n20019), .dinb(n1698), .dout(n20094));
  jnot g02293(.din(n1822), .dout(n20097));
  jand g02294(.dina(n20097), .dinb(n20094), .dout(n20098));
  jor  g02295(.dina(n20098), .dinb(b2 ), .dout(n20099));
  jnot g02296(.din(n1563), .dout(n20101));
  jnot g02297(.din(n1630), .dout(n20102));
  jnot g02298(.din(n19905), .dout(n20103));
  jnot g02299(.din(n19910), .dout(n20104));
  jnot g02300(.din(n19915), .dout(n20105));
  jnot g02301(.din(n19920), .dout(n20106));
  jnot g02302(.din(n19925), .dout(n20107));
  jnot g02303(.din(n19930), .dout(n20108));
  jnot g02304(.din(n19935), .dout(n20109));
  jnot g02305(.din(n19940), .dout(n20110));
  jnot g02306(.din(n19945), .dout(n20111));
  jnot g02307(.din(n19950), .dout(n20112));
  jnot g02308(.din(n19955), .dout(n20113));
  jnot g02309(.din(n19960), .dout(n20114));
  jnot g02310(.din(n19965), .dout(n20115));
  jnot g02311(.din(n19971), .dout(n20116));
  jxor g02312(.dina(n1698), .dinb(n258), .dout(n20117));
  jor  g02313(.dina(n20117), .dinb(n1702), .dout(n20118));
  jand g02314(.dina(n20118), .dinb(n20116), .dout(n20119));
  jnot g02315(.din(n19978), .dout(n20120));
  jor  g02316(.dina(n20120), .dinb(n20119), .dout(n20121));
  jand g02317(.dina(n20121), .dinb(n20115), .dout(n20122));
  jnot g02318(.din(n19981), .dout(n20123));
  jor  g02319(.dina(n20123), .dinb(n20122), .dout(n20124));
  jand g02320(.dina(n20124), .dinb(n20114), .dout(n20125));
  jnot g02321(.din(n19984), .dout(n20126));
  jor  g02322(.dina(n20126), .dinb(n20125), .dout(n20127));
  jand g02323(.dina(n20127), .dinb(n20113), .dout(n20128));
  jnot g02324(.din(n19987), .dout(n20129));
  jor  g02325(.dina(n20129), .dinb(n20128), .dout(n20130));
  jand g02326(.dina(n20130), .dinb(n20112), .dout(n20131));
  jnot g02327(.din(n19990), .dout(n20132));
  jor  g02328(.dina(n20132), .dinb(n20131), .dout(n20133));
  jand g02329(.dina(n20133), .dinb(n20111), .dout(n20134));
  jnot g02330(.din(n19993), .dout(n20135));
  jor  g02331(.dina(n20135), .dinb(n20134), .dout(n20136));
  jand g02332(.dina(n20136), .dinb(n20110), .dout(n20137));
  jnot g02333(.din(n19996), .dout(n20138));
  jor  g02334(.dina(n20138), .dinb(n20137), .dout(n20139));
  jand g02335(.dina(n20139), .dinb(n20109), .dout(n20140));
  jnot g02336(.din(n19999), .dout(n20141));
  jor  g02337(.dina(n20141), .dinb(n20140), .dout(n20142));
  jand g02338(.dina(n20142), .dinb(n20108), .dout(n20143));
  jnot g02339(.din(n20002), .dout(n20144));
  jor  g02340(.dina(n20144), .dinb(n20143), .dout(n20145));
  jand g02341(.dina(n20145), .dinb(n20107), .dout(n20146));
  jnot g02342(.din(n20005), .dout(n20147));
  jor  g02343(.dina(n20147), .dinb(n20146), .dout(n20148));
  jand g02344(.dina(n20148), .dinb(n20106), .dout(n20149));
  jnot g02345(.din(n20008), .dout(n20150));
  jor  g02346(.dina(n20150), .dinb(n20149), .dout(n20151));
  jand g02347(.dina(n20151), .dinb(n20105), .dout(n20152));
  jnot g02348(.din(n20011), .dout(n20153));
  jor  g02349(.dina(n20153), .dinb(n20152), .dout(n20154));
  jand g02350(.dina(n20154), .dinb(n20104), .dout(n20155));
  jnot g02351(.din(n20014), .dout(n20156));
  jor  g02352(.dina(n20156), .dinb(n20155), .dout(n20157));
  jand g02353(.dina(n20157), .dinb(n20103), .dout(n20158));
  jand g02354(.dina(n20158), .dinb(n20102), .dout(n20159));
  jor  g02355(.dina(n20159), .dinb(n19896), .dout(n20160));
  jor  g02356(.dina(n20160), .dinb(n20101), .dout(n20161));
  jand g02357(.dina(n20161), .dinb(a48 ), .dout(n20162));
  jnot g02358(.din(n1827), .dout(n20163));
  jor  g02359(.dina(n20160), .dinb(n20163), .dout(n20164));
  jor  g02360(.dina(n1828), .dinb(n20162), .dout(n20166));
  jand g02361(.dina(n20166), .dinb(n258), .dout(n20167));
  jnot g02362(.din(n1895), .dout(n20227));
  jnot g02363(.din(n1903), .dout(n20233));
  jnot g02364(.din(n1904), .dout(n20239));
  jnot g02365(.din(n1909), .dout(n20245));
  jnot g02366(.din(n1914), .dout(n20251));
  jnot g02367(.din(n1919), .dout(n20257));
  jnot g02368(.din(n1924), .dout(n20263));
  jnot g02369(.din(n1929), .dout(n20269));
  jnot g02370(.din(n1934), .dout(n20275));
  jnot g02371(.din(n1939), .dout(n20281));
  jnot g02372(.din(n1944), .dout(n20287));
  jnot g02373(.din(n1949), .dout(n20293));
  jnot g02374(.din(n1954), .dout(n20299));
  jnot g02375(.din(n1959), .dout(n20305));
  jnot g02376(.din(n1964), .dout(n20313));
  jnot g02377(.din(n1969), .dout(n20321));
  jnot g02378(.din(n1973), .dout(n20322));
  jnot g02379(.din(n1758), .dout(n20323));
  jnot g02380(.din(n1763), .dout(n20324));
  jnot g02381(.din(n1764), .dout(n20325));
  jnot g02382(.din(n1769), .dout(n20326));
  jnot g02383(.din(n1774), .dout(n20327));
  jnot g02384(.din(n1779), .dout(n20328));
  jnot g02385(.din(n1784), .dout(n20329));
  jnot g02386(.din(n1789), .dout(n20330));
  jnot g02387(.din(n1794), .dout(n20331));
  jnot g02388(.din(n1799), .dout(n20332));
  jnot g02389(.din(n1804), .dout(n20333));
  jnot g02390(.din(n1809), .dout(n20334));
  jnot g02391(.din(n1814), .dout(n20335));
  jnot g02392(.din(n1819), .dout(n20336));
  jnot g02393(.din(n20167), .dout(n20337));
  jxor g02394(.dina(n1830), .dinb(n258), .dout(n20338));
  jor  g02395(.dina(n20338), .dinb(n1834), .dout(n20339));
  jand g02396(.dina(n20339), .dinb(n20337), .dout(n20340));
  jnot g02397(.din(n1839), .dout(n20341));
  jor  g02398(.dina(n20341), .dinb(n20340), .dout(n20342));
  jand g02399(.dina(n20342), .dinb(n20099), .dout(n20343));
  jnot g02400(.din(n1842), .dout(n20344));
  jor  g02401(.dina(n20344), .dinb(n20343), .dout(n20345));
  jand g02402(.dina(n20345), .dinb(n20336), .dout(n20346));
  jnot g02403(.din(n1845), .dout(n20347));
  jor  g02404(.dina(n20347), .dinb(n20346), .dout(n20348));
  jand g02405(.dina(n20348), .dinb(n20335), .dout(n20349));
  jnot g02406(.din(n1848), .dout(n20350));
  jor  g02407(.dina(n20350), .dinb(n20349), .dout(n20351));
  jand g02408(.dina(n20351), .dinb(n20334), .dout(n20352));
  jnot g02409(.din(n1851), .dout(n20353));
  jor  g02410(.dina(n20353), .dinb(n20352), .dout(n20354));
  jand g02411(.dina(n20354), .dinb(n20333), .dout(n20355));
  jnot g02412(.din(n1854), .dout(n20356));
  jor  g02413(.dina(n20356), .dinb(n20355), .dout(n20357));
  jand g02414(.dina(n20357), .dinb(n20332), .dout(n20358));
  jnot g02415(.din(n1857), .dout(n20359));
  jor  g02416(.dina(n20359), .dinb(n20358), .dout(n20360));
  jand g02417(.dina(n20360), .dinb(n20331), .dout(n20361));
  jnot g02418(.din(n1860), .dout(n20362));
  jor  g02419(.dina(n20362), .dinb(n20361), .dout(n20363));
  jand g02420(.dina(n20363), .dinb(n20330), .dout(n20364));
  jnot g02421(.din(n1863), .dout(n20365));
  jor  g02422(.dina(n20365), .dinb(n20364), .dout(n20366));
  jand g02423(.dina(n20366), .dinb(n20329), .dout(n20367));
  jnot g02424(.din(n1866), .dout(n20368));
  jor  g02425(.dina(n20368), .dinb(n20367), .dout(n20369));
  jand g02426(.dina(n20369), .dinb(n20328), .dout(n20370));
  jnot g02427(.din(n1869), .dout(n20371));
  jor  g02428(.dina(n20371), .dinb(n20370), .dout(n20372));
  jand g02429(.dina(n20372), .dinb(n20327), .dout(n20373));
  jnot g02430(.din(n1872), .dout(n20374));
  jor  g02431(.dina(n20374), .dinb(n20373), .dout(n20375));
  jand g02432(.dina(n20375), .dinb(n20326), .dout(n20376));
  jnot g02433(.din(n1875), .dout(n20377));
  jor  g02434(.dina(n20377), .dinb(n20376), .dout(n20378));
  jand g02435(.dina(n20378), .dinb(n20325), .dout(n20379));
  jnot g02436(.din(n1878), .dout(n20380));
  jor  g02437(.dina(n20380), .dinb(n20379), .dout(n20381));
  jand g02438(.dina(n20381), .dinb(n20324), .dout(n20382));
  jor  g02439(.dina(n1882), .dinb(n20382), .dout(n20383));
  jand g02440(.dina(n20383), .dinb(n20323), .dout(n20384));
  jor  g02441(.dina(n20384), .dinb(n20322), .dout(n20385));
  jand g02442(.dina(n20385), .dinb(a47 ), .dout(n20386));
  jnot g02443(.din(n1976), .dout(n20387));
  jor  g02444(.dina(n20384), .dinb(n20387), .dout(n20388));
  jor  g02445(.dina(n1977), .dinb(n20386), .dout(n20390));
  jand g02446(.dina(n20390), .dinb(n258), .dout(n20391));
  jxor g02447(.dina(n1979), .dinb(n258), .dout(n20396));
  jor  g02448(.dina(n20396), .dinb(n1983), .dout(n20397));
  jand g02449(.dina(n20397), .dinb(n1980), .dout(n20398));
  jnot g02450(.din(n1988), .dout(n20400));
  jor  g02451(.dina(n20400), .dinb(n20398), .dout(n20401));
  jand g02452(.dina(n20401), .dinb(n20321), .dout(n20402));
  jnot g02453(.din(n1991), .dout(n20404));
  jor  g02454(.dina(n20404), .dinb(n20402), .dout(n20405));
  jand g02455(.dina(n20405), .dinb(n20313), .dout(n20406));
  jnot g02456(.din(n1994), .dout(n20408));
  jor  g02457(.dina(n20408), .dinb(n20406), .dout(n20409));
  jand g02458(.dina(n20409), .dinb(n20305), .dout(n20410));
  jnot g02459(.din(n1997), .dout(n20412));
  jor  g02460(.dina(n20412), .dinb(n20410), .dout(n20413));
  jand g02461(.dina(n20413), .dinb(n20299), .dout(n20414));
  jnot g02462(.din(n2000), .dout(n20416));
  jor  g02463(.dina(n20416), .dinb(n20414), .dout(n20417));
  jand g02464(.dina(n20417), .dinb(n20293), .dout(n20418));
  jnot g02465(.din(n2003), .dout(n20420));
  jor  g02466(.dina(n20420), .dinb(n20418), .dout(n20421));
  jand g02467(.dina(n20421), .dinb(n20287), .dout(n20422));
  jnot g02468(.din(n2006), .dout(n20424));
  jor  g02469(.dina(n20424), .dinb(n20422), .dout(n20425));
  jand g02470(.dina(n20425), .dinb(n20281), .dout(n20426));
  jnot g02471(.din(n2009), .dout(n20428));
  jor  g02472(.dina(n20428), .dinb(n20426), .dout(n20429));
  jand g02473(.dina(n20429), .dinb(n20275), .dout(n20430));
  jnot g02474(.din(n2012), .dout(n20432));
  jor  g02475(.dina(n20432), .dinb(n20430), .dout(n20433));
  jand g02476(.dina(n20433), .dinb(n20269), .dout(n20434));
  jnot g02477(.din(n2015), .dout(n20436));
  jor  g02478(.dina(n20436), .dinb(n20434), .dout(n20437));
  jand g02479(.dina(n20437), .dinb(n20263), .dout(n20438));
  jnot g02480(.din(n2018), .dout(n20440));
  jor  g02481(.dina(n20440), .dinb(n20438), .dout(n20441));
  jand g02482(.dina(n20441), .dinb(n20257), .dout(n20442));
  jnot g02483(.din(n2021), .dout(n20444));
  jor  g02484(.dina(n20444), .dinb(n20442), .dout(n20445));
  jand g02485(.dina(n20445), .dinb(n20251), .dout(n20446));
  jnot g02486(.din(n2024), .dout(n20448));
  jor  g02487(.dina(n20448), .dinb(n20446), .dout(n20449));
  jand g02488(.dina(n20449), .dinb(n20245), .dout(n20450));
  jnot g02489(.din(n2027), .dout(n20452));
  jor  g02490(.dina(n20452), .dinb(n20450), .dout(n20453));
  jand g02491(.dina(n20453), .dinb(n20239), .dout(n20454));
  jnot g02492(.din(n2030), .dout(n20456));
  jor  g02493(.dina(n20456), .dinb(n20454), .dout(n20457));
  jand g02494(.dina(n20457), .dinb(n20233), .dout(n20458));
  jor  g02495(.dina(n2033), .dinb(n1897), .dout(n20460));
  jor  g02496(.dina(n20460), .dinb(n20458), .dout(n20461));
  jand g02497(.dina(n20461), .dinb(n20227), .dout(n20462));
  jnot g02498(.din(n20460), .dout(n20496));
  jand g02499(.dina(n20496), .dinb(n2032), .dout(n20497));
  jor  g02500(.dina(n1896), .dinb(n20497), .dout(n20499));
  jxor g02501(.dina(n2033), .dinb(n2032), .dout(n20500));
  jand g02502(.dina(n20500), .dinb(n20499), .dout(n20501));
  jor  g02503(.dina(n20501), .dinb(n20462), .dout(n20502));
  jnot g02504(.din(n20502), .dout(n20503));
  jand g02505(.dina(n20502), .dinb(b18 ), .dout(n20504));
  jnot g02506(.din(n20504), .dout(n20505));
  jand g02507(.dina(n20503), .dinb(n422), .dout(n20506));
  jand g02508(.dina(n2045), .dinb(n20461), .dout(n20508));
  jand g02509(.dina(n20508), .dinb(n1902), .dout(n20509));
  jand g02510(.dina(n2054), .dinb(n20499), .dout(n20511));
  jor  g02511(.dina(n20511), .dinb(n20509), .dout(n20512));
  jand g02512(.dina(n20512), .dinb(n421), .dout(n20513));
  jand g02513(.dina(n20508), .dinb(n1891), .dout(n20514));
  jand g02514(.dina(n2040), .dinb(n20499), .dout(n20516));
  jor  g02515(.dina(n20516), .dinb(n20514), .dout(n20517));
  jand g02516(.dina(n20517), .dinb(n433), .dout(n20518));
  jand g02517(.dina(n20508), .dinb(n1908), .dout(n20519));
  jand g02518(.dina(n2060), .dinb(n20499), .dout(n20521));
  jor  g02519(.dina(n20521), .dinb(n20519), .dout(n20522));
  jand g02520(.dina(n20522), .dinb(n432), .dout(n20523));
  jand g02521(.dina(n20508), .dinb(n1913), .dout(n20524));
  jand g02522(.dina(n2065), .dinb(n20499), .dout(n20526));
  jor  g02523(.dina(n20526), .dinb(n20524), .dout(n20527));
  jand g02524(.dina(n20527), .dinb(n436), .dout(n20528));
  jand g02525(.dina(n20508), .dinb(n1918), .dout(n20529));
  jand g02526(.dina(n2070), .dinb(n20499), .dout(n20531));
  jor  g02527(.dina(n20531), .dinb(n20529), .dout(n20532));
  jand g02528(.dina(n20532), .dinb(n435), .dout(n20533));
  jand g02529(.dina(n20508), .dinb(n1923), .dout(n20534));
  jand g02530(.dina(n2075), .dinb(n20499), .dout(n20536));
  jor  g02531(.dina(n20536), .dinb(n20534), .dout(n20537));
  jand g02532(.dina(n20537), .dinb(n440), .dout(n20538));
  jand g02533(.dina(n20508), .dinb(n1928), .dout(n20539));
  jand g02534(.dina(n2080), .dinb(n20499), .dout(n20541));
  jor  g02535(.dina(n20541), .dinb(n20539), .dout(n20542));
  jand g02536(.dina(n20542), .dinb(n439), .dout(n20543));
  jand g02537(.dina(n20508), .dinb(n1933), .dout(n20544));
  jand g02538(.dina(n2085), .dinb(n20499), .dout(n20546));
  jor  g02539(.dina(n20546), .dinb(n20544), .dout(n20547));
  jand g02540(.dina(n20547), .dinb(n325), .dout(n20548));
  jand g02541(.dina(n20508), .dinb(n1938), .dout(n20549));
  jand g02542(.dina(n2090), .dinb(n20499), .dout(n20551));
  jor  g02543(.dina(n20551), .dinb(n20549), .dout(n20552));
  jand g02544(.dina(n20552), .dinb(n324), .dout(n20553));
  jand g02545(.dina(n20508), .dinb(n1943), .dout(n20554));
  jand g02546(.dina(n2095), .dinb(n20499), .dout(n20556));
  jor  g02547(.dina(n20556), .dinb(n20554), .dout(n20557));
  jand g02548(.dina(n20557), .dinb(n323), .dout(n20558));
  jand g02549(.dina(n20508), .dinb(n1948), .dout(n20559));
  jand g02550(.dina(n2100), .dinb(n20499), .dout(n20561));
  jor  g02551(.dina(n20561), .dinb(n20559), .dout(n20562));
  jand g02552(.dina(n20562), .dinb(n335), .dout(n20563));
  jand g02553(.dina(n20508), .dinb(n1953), .dout(n20564));
  jand g02554(.dina(n2105), .dinb(n20499), .dout(n20566));
  jor  g02555(.dina(n20566), .dinb(n20564), .dout(n20567));
  jand g02556(.dina(n20567), .dinb(n334), .dout(n20568));
  jand g02557(.dina(n20508), .dinb(n1958), .dout(n20569));
  jand g02558(.dina(n2110), .dinb(n20499), .dout(n20571));
  jor  g02559(.dina(n20571), .dinb(n20569), .dout(n20572));
  jand g02560(.dina(n20572), .dinb(n338), .dout(n20573));
  jand g02561(.dina(n20508), .dinb(n1963), .dout(n20574));
  jand g02562(.dina(n2115), .dinb(n20499), .dout(n20576));
  jor  g02563(.dina(n20576), .dinb(n20574), .dout(n20577));
  jand g02564(.dina(n20577), .dinb(n337), .dout(n20578));
  jand g02565(.dina(n20508), .dinb(n1968), .dout(n20579));
  jand g02566(.dina(n2120), .dinb(n20499), .dout(n20581));
  jor  g02567(.dina(n20581), .dinb(n20579), .dout(n20582));
  jand g02568(.dina(n20582), .dinb(n344), .dout(n20583));
  jand g02569(.dina(n20508), .dinb(n20390), .dout(n20584));
  jand g02570(.dina(n2125), .dinb(n20499), .dout(n20586));
  jor  g02571(.dina(n20586), .dinb(n20584), .dout(n20587));
  jand g02572(.dina(n20587), .dinb(n348), .dout(n20588));
  jor  g02573(.dina(n20508), .dinb(n18364), .dout(n20589));
  jand g02574(.dina(n20589), .dinb(a46 ), .dout(n20590));
  jor  g02575(.dina(n20508), .dinb(n1984), .dout(n20591));
  jor  g02576(.dina(n2133), .dinb(n20590), .dout(n20593));
  jand g02577(.dina(n20593), .dinb(n258), .dout(n20594));
  jand g02578(.dina(n20499), .dinb(b0 ), .dout(n20595));
  jor  g02579(.dina(n20595), .dinb(n1982), .dout(n20596));
  jand g02580(.dina(n20591), .dinb(n20596), .dout(n20597));
  jxor g02581(.dina(n20597), .dinb(b1 ), .dout(n20598));
  jand g02582(.dina(n20598), .dinb(n2140), .dout(n20599));
  jor  g02583(.dina(n20599), .dinb(n20594), .dout(n20600));
  jxor g02584(.dina(n20587), .dinb(n348), .dout(n20601));
  jand g02585(.dina(n20601), .dinb(n20600), .dout(n20602));
  jor  g02586(.dina(n20602), .dinb(n20588), .dout(n20603));
  jxor g02587(.dina(n20582), .dinb(n344), .dout(n20604));
  jand g02588(.dina(n20604), .dinb(n20603), .dout(n20605));
  jor  g02589(.dina(n20605), .dinb(n20583), .dout(n20606));
  jxor g02590(.dina(n20577), .dinb(n337), .dout(n20607));
  jand g02591(.dina(n20607), .dinb(n20606), .dout(n20608));
  jor  g02592(.dina(n20608), .dinb(n20578), .dout(n20609));
  jxor g02593(.dina(n20572), .dinb(n338), .dout(n20610));
  jand g02594(.dina(n20610), .dinb(n20609), .dout(n20611));
  jor  g02595(.dina(n20611), .dinb(n20573), .dout(n20612));
  jxor g02596(.dina(n20567), .dinb(n334), .dout(n20613));
  jand g02597(.dina(n20613), .dinb(n20612), .dout(n20614));
  jor  g02598(.dina(n20614), .dinb(n20568), .dout(n20615));
  jxor g02599(.dina(n20562), .dinb(n335), .dout(n20616));
  jand g02600(.dina(n20616), .dinb(n20615), .dout(n20617));
  jor  g02601(.dina(n20617), .dinb(n20563), .dout(n20618));
  jxor g02602(.dina(n20557), .dinb(n323), .dout(n20619));
  jand g02603(.dina(n20619), .dinb(n20618), .dout(n20620));
  jor  g02604(.dina(n20620), .dinb(n20558), .dout(n20621));
  jxor g02605(.dina(n20552), .dinb(n324), .dout(n20622));
  jand g02606(.dina(n20622), .dinb(n20621), .dout(n20623));
  jor  g02607(.dina(n20623), .dinb(n20553), .dout(n20624));
  jxor g02608(.dina(n20547), .dinb(n325), .dout(n20625));
  jand g02609(.dina(n20625), .dinb(n20624), .dout(n20626));
  jor  g02610(.dina(n20626), .dinb(n20548), .dout(n20627));
  jxor g02611(.dina(n20542), .dinb(n439), .dout(n20628));
  jand g02612(.dina(n20628), .dinb(n20627), .dout(n20629));
  jor  g02613(.dina(n20629), .dinb(n20543), .dout(n20630));
  jxor g02614(.dina(n20537), .dinb(n440), .dout(n20631));
  jand g02615(.dina(n20631), .dinb(n20630), .dout(n20632));
  jor  g02616(.dina(n20632), .dinb(n20538), .dout(n20633));
  jxor g02617(.dina(n20532), .dinb(n435), .dout(n20634));
  jand g02618(.dina(n20634), .dinb(n20633), .dout(n20635));
  jor  g02619(.dina(n20635), .dinb(n20533), .dout(n20636));
  jxor g02620(.dina(n20527), .dinb(n436), .dout(n20637));
  jand g02621(.dina(n20637), .dinb(n20636), .dout(n20638));
  jor  g02622(.dina(n20638), .dinb(n20528), .dout(n20639));
  jxor g02623(.dina(n20522), .dinb(n432), .dout(n20640));
  jand g02624(.dina(n20640), .dinb(n20639), .dout(n20641));
  jor  g02625(.dina(n20641), .dinb(n20523), .dout(n20642));
  jxor g02626(.dina(n20517), .dinb(n433), .dout(n20643));
  jand g02627(.dina(n20643), .dinb(n20642), .dout(n20644));
  jor  g02628(.dina(n20644), .dinb(n20518), .dout(n20645));
  jxor g02629(.dina(n20512), .dinb(n421), .dout(n20646));
  jand g02630(.dina(n20646), .dinb(n20645), .dout(n20647));
  jor  g02631(.dina(n20647), .dinb(n20513), .dout(n20648));
  jor  g02632(.dina(n20648), .dinb(n20506), .dout(n20649));
  jand g02633(.dina(n20649), .dinb(n20505), .dout(n20650));
  jand g02634(.dina(n20650), .dinb(n2197), .dout(n20651));
  jnot g02635(.din(n20651), .dout(n20652));
  jand g02636(.dina(n20652), .dinb(n20503), .dout(n20653));
  jand g02637(.dina(n20506), .dinb(n2197), .dout(n20654));
  jand g02638(.dina(n20654), .dinb(n20648), .dout(n20655));
  jor  g02639(.dina(n20655), .dinb(n20653), .dout(n20656));
  jand g02640(.dina(n20656), .dinb(n416), .dout(n20657));
  jnot g02641(.din(n20657), .dout(n20658));
  jand g02642(.dina(n20652), .dinb(n20512), .dout(n20659));
  jxor g02643(.dina(n20646), .dinb(n20645), .dout(n20660));
  jand g02644(.dina(n20660), .dinb(n20651), .dout(n20661));
  jor  g02645(.dina(n20661), .dinb(n20659), .dout(n20662));
  jand g02646(.dina(n20662), .dinb(n422), .dout(n20663));
  jnot g02647(.din(n20663), .dout(n20664));
  jand g02648(.dina(n20652), .dinb(n20517), .dout(n20665));
  jxor g02649(.dina(n20643), .dinb(n20642), .dout(n20666));
  jand g02650(.dina(n20666), .dinb(n20651), .dout(n20667));
  jor  g02651(.dina(n20667), .dinb(n20665), .dout(n20668));
  jand g02652(.dina(n20668), .dinb(n421), .dout(n20669));
  jnot g02653(.din(n20669), .dout(n20670));
  jand g02654(.dina(n20652), .dinb(n20522), .dout(n20671));
  jxor g02655(.dina(n20640), .dinb(n20639), .dout(n20672));
  jand g02656(.dina(n20672), .dinb(n20651), .dout(n20673));
  jor  g02657(.dina(n20673), .dinb(n20671), .dout(n20674));
  jand g02658(.dina(n20674), .dinb(n433), .dout(n20675));
  jnot g02659(.din(n20675), .dout(n20676));
  jand g02660(.dina(n20652), .dinb(n20527), .dout(n20677));
  jxor g02661(.dina(n20637), .dinb(n20636), .dout(n20678));
  jand g02662(.dina(n20678), .dinb(n20651), .dout(n20679));
  jor  g02663(.dina(n20679), .dinb(n20677), .dout(n20680));
  jand g02664(.dina(n20680), .dinb(n432), .dout(n20681));
  jnot g02665(.din(n20681), .dout(n20682));
  jand g02666(.dina(n20652), .dinb(n20532), .dout(n20683));
  jxor g02667(.dina(n20634), .dinb(n20633), .dout(n20684));
  jand g02668(.dina(n20684), .dinb(n20651), .dout(n20685));
  jor  g02669(.dina(n20685), .dinb(n20683), .dout(n20686));
  jand g02670(.dina(n20686), .dinb(n436), .dout(n20687));
  jnot g02671(.din(n20687), .dout(n20688));
  jand g02672(.dina(n20652), .dinb(n20537), .dout(n20689));
  jxor g02673(.dina(n20631), .dinb(n20630), .dout(n20690));
  jand g02674(.dina(n20690), .dinb(n20651), .dout(n20691));
  jor  g02675(.dina(n20691), .dinb(n20689), .dout(n20692));
  jand g02676(.dina(n20692), .dinb(n435), .dout(n20693));
  jnot g02677(.din(n20693), .dout(n20694));
  jand g02678(.dina(n20652), .dinb(n20542), .dout(n20695));
  jxor g02679(.dina(n20628), .dinb(n20627), .dout(n20696));
  jand g02680(.dina(n20696), .dinb(n20651), .dout(n20697));
  jor  g02681(.dina(n20697), .dinb(n20695), .dout(n20698));
  jand g02682(.dina(n20698), .dinb(n440), .dout(n20699));
  jnot g02683(.din(n20699), .dout(n20700));
  jand g02684(.dina(n20652), .dinb(n20547), .dout(n20701));
  jxor g02685(.dina(n20625), .dinb(n20624), .dout(n20702));
  jand g02686(.dina(n20702), .dinb(n20651), .dout(n20703));
  jor  g02687(.dina(n20703), .dinb(n20701), .dout(n20704));
  jand g02688(.dina(n20704), .dinb(n439), .dout(n20705));
  jnot g02689(.din(n20705), .dout(n20706));
  jand g02690(.dina(n20652), .dinb(n20552), .dout(n20707));
  jxor g02691(.dina(n20622), .dinb(n20621), .dout(n20708));
  jand g02692(.dina(n20708), .dinb(n20651), .dout(n20709));
  jor  g02693(.dina(n20709), .dinb(n20707), .dout(n20710));
  jand g02694(.dina(n20710), .dinb(n325), .dout(n20711));
  jnot g02695(.din(n20711), .dout(n20712));
  jand g02696(.dina(n20652), .dinb(n20557), .dout(n20713));
  jxor g02697(.dina(n20619), .dinb(n20618), .dout(n20714));
  jand g02698(.dina(n20714), .dinb(n20651), .dout(n20715));
  jor  g02699(.dina(n20715), .dinb(n20713), .dout(n20716));
  jand g02700(.dina(n20716), .dinb(n324), .dout(n20717));
  jnot g02701(.din(n20717), .dout(n20718));
  jand g02702(.dina(n20652), .dinb(n20562), .dout(n20719));
  jxor g02703(.dina(n20616), .dinb(n20615), .dout(n20720));
  jand g02704(.dina(n20720), .dinb(n20651), .dout(n20721));
  jor  g02705(.dina(n20721), .dinb(n20719), .dout(n20722));
  jand g02706(.dina(n20722), .dinb(n323), .dout(n20723));
  jnot g02707(.din(n20723), .dout(n20724));
  jand g02708(.dina(n20652), .dinb(n20567), .dout(n20725));
  jxor g02709(.dina(n20613), .dinb(n20612), .dout(n20726));
  jand g02710(.dina(n20726), .dinb(n20651), .dout(n20727));
  jor  g02711(.dina(n20727), .dinb(n20725), .dout(n20728));
  jand g02712(.dina(n20728), .dinb(n335), .dout(n20729));
  jnot g02713(.din(n20729), .dout(n20730));
  jand g02714(.dina(n20652), .dinb(n20572), .dout(n20731));
  jxor g02715(.dina(n20610), .dinb(n20609), .dout(n20732));
  jand g02716(.dina(n20732), .dinb(n20651), .dout(n20733));
  jor  g02717(.dina(n20733), .dinb(n20731), .dout(n20734));
  jand g02718(.dina(n20734), .dinb(n334), .dout(n20735));
  jnot g02719(.din(n20735), .dout(n20736));
  jand g02720(.dina(n20652), .dinb(n20577), .dout(n20737));
  jxor g02721(.dina(n20607), .dinb(n20606), .dout(n20738));
  jand g02722(.dina(n20738), .dinb(n20651), .dout(n20739));
  jor  g02723(.dina(n20739), .dinb(n20737), .dout(n20740));
  jand g02724(.dina(n20740), .dinb(n338), .dout(n20741));
  jnot g02725(.din(n20741), .dout(n20742));
  jand g02726(.dina(n20652), .dinb(n20582), .dout(n20743));
  jxor g02727(.dina(n20604), .dinb(n20603), .dout(n20744));
  jand g02728(.dina(n20744), .dinb(n20651), .dout(n20745));
  jor  g02729(.dina(n20745), .dinb(n20743), .dout(n20746));
  jand g02730(.dina(n20746), .dinb(n337), .dout(n20747));
  jnot g02731(.din(n20747), .dout(n20748));
  jnot g02732(.din(n20587), .dout(n20749));
  jor  g02733(.dina(n20651), .dinb(n20749), .dout(n20750));
  jxor g02734(.dina(n20601), .dinb(n20600), .dout(n20751));
  jnot g02735(.din(n20751), .dout(n20752));
  jor  g02736(.dina(n20752), .dinb(n20652), .dout(n20753));
  jand g02737(.dina(n20753), .dinb(n20750), .dout(n20754));
  jor  g02738(.dina(n20754), .dinb(b3 ), .dout(n20755));
  jor  g02739(.dina(n20651), .dinb(n20597), .dout(n20756));
  jxor g02740(.dina(n20598), .dinb(n2140), .dout(n20757));
  jand g02741(.dina(n20757), .dinb(n20651), .dout(n20758));
  jnot g02742(.din(n20758), .dout(n20759));
  jand g02743(.dina(n20759), .dinb(n20756), .dout(n20760));
  jor  g02744(.dina(n20760), .dinb(b2 ), .dout(n20761));
  jand g02745(.dina(n20650), .dinb(n1972), .dout(n20762));
  jor  g02746(.dina(n20762), .dinb(n2138), .dout(n20763));
  jnot g02747(.din(n2292), .dout(n20764));
  jnot g02748(.din(n20506), .dout(n20765));
  jnot g02749(.din(n20513), .dout(n20766));
  jnot g02750(.din(n20518), .dout(n20767));
  jnot g02751(.din(n20523), .dout(n20768));
  jnot g02752(.din(n20528), .dout(n20769));
  jnot g02753(.din(n20533), .dout(n20770));
  jnot g02754(.din(n20538), .dout(n20771));
  jnot g02755(.din(n20543), .dout(n20772));
  jnot g02756(.din(n20548), .dout(n20773));
  jnot g02757(.din(n20553), .dout(n20774));
  jnot g02758(.din(n20558), .dout(n20775));
  jnot g02759(.din(n20563), .dout(n20776));
  jnot g02760(.din(n20568), .dout(n20777));
  jnot g02761(.din(n20573), .dout(n20778));
  jnot g02762(.din(n20578), .dout(n20779));
  jnot g02763(.din(n20583), .dout(n20780));
  jnot g02764(.din(n20588), .dout(n20781));
  jnot g02765(.din(n20594), .dout(n20782));
  jxor g02766(.dina(n20597), .dinb(n258), .dout(n20783));
  jor  g02767(.dina(n20783), .dinb(n2139), .dout(n20784));
  jand g02768(.dina(n20784), .dinb(n20782), .dout(n20785));
  jnot g02769(.din(n20601), .dout(n20786));
  jor  g02770(.dina(n20786), .dinb(n20785), .dout(n20787));
  jand g02771(.dina(n20787), .dinb(n20781), .dout(n20788));
  jnot g02772(.din(n20604), .dout(n20789));
  jor  g02773(.dina(n20789), .dinb(n20788), .dout(n20790));
  jand g02774(.dina(n20790), .dinb(n20780), .dout(n20791));
  jnot g02775(.din(n20607), .dout(n20792));
  jor  g02776(.dina(n20792), .dinb(n20791), .dout(n20793));
  jand g02777(.dina(n20793), .dinb(n20779), .dout(n20794));
  jnot g02778(.din(n20610), .dout(n20795));
  jor  g02779(.dina(n20795), .dinb(n20794), .dout(n20796));
  jand g02780(.dina(n20796), .dinb(n20778), .dout(n20797));
  jnot g02781(.din(n20613), .dout(n20798));
  jor  g02782(.dina(n20798), .dinb(n20797), .dout(n20799));
  jand g02783(.dina(n20799), .dinb(n20777), .dout(n20800));
  jnot g02784(.din(n20616), .dout(n20801));
  jor  g02785(.dina(n20801), .dinb(n20800), .dout(n20802));
  jand g02786(.dina(n20802), .dinb(n20776), .dout(n20803));
  jnot g02787(.din(n20619), .dout(n20804));
  jor  g02788(.dina(n20804), .dinb(n20803), .dout(n20805));
  jand g02789(.dina(n20805), .dinb(n20775), .dout(n20806));
  jnot g02790(.din(n20622), .dout(n20807));
  jor  g02791(.dina(n20807), .dinb(n20806), .dout(n20808));
  jand g02792(.dina(n20808), .dinb(n20774), .dout(n20809));
  jnot g02793(.din(n20625), .dout(n20810));
  jor  g02794(.dina(n20810), .dinb(n20809), .dout(n20811));
  jand g02795(.dina(n20811), .dinb(n20773), .dout(n20812));
  jnot g02796(.din(n20628), .dout(n20813));
  jor  g02797(.dina(n20813), .dinb(n20812), .dout(n20814));
  jand g02798(.dina(n20814), .dinb(n20772), .dout(n20815));
  jnot g02799(.din(n20631), .dout(n20816));
  jor  g02800(.dina(n20816), .dinb(n20815), .dout(n20817));
  jand g02801(.dina(n20817), .dinb(n20771), .dout(n20818));
  jnot g02802(.din(n20634), .dout(n20819));
  jor  g02803(.dina(n20819), .dinb(n20818), .dout(n20820));
  jand g02804(.dina(n20820), .dinb(n20770), .dout(n20821));
  jnot g02805(.din(n20637), .dout(n20822));
  jor  g02806(.dina(n20822), .dinb(n20821), .dout(n20823));
  jand g02807(.dina(n20823), .dinb(n20769), .dout(n20824));
  jnot g02808(.din(n20640), .dout(n20825));
  jor  g02809(.dina(n20825), .dinb(n20824), .dout(n20826));
  jand g02810(.dina(n20826), .dinb(n20768), .dout(n20827));
  jnot g02811(.din(n20643), .dout(n20828));
  jor  g02812(.dina(n20828), .dinb(n20827), .dout(n20829));
  jand g02813(.dina(n20829), .dinb(n20767), .dout(n20830));
  jnot g02814(.din(n20646), .dout(n20831));
  jor  g02815(.dina(n20831), .dinb(n20830), .dout(n20832));
  jand g02816(.dina(n20832), .dinb(n20766), .dout(n20833));
  jand g02817(.dina(n20833), .dinb(n20765), .dout(n20834));
  jor  g02818(.dina(n20834), .dinb(n20504), .dout(n20835));
  jor  g02819(.dina(n20835), .dinb(n20764), .dout(n20836));
  jand g02820(.dina(n20836), .dinb(n20763), .dout(n20837));
  jor  g02821(.dina(n20837), .dinb(b1 ), .dout(n20838));
  jxor g02822(.dina(n20837), .dinb(n258), .dout(n20839));
  jor  g02823(.dina(n20839), .dinb(n2299), .dout(n20840));
  jand g02824(.dina(n20840), .dinb(n20838), .dout(n20841));
  jxor g02825(.dina(n20760), .dinb(n348), .dout(n20842));
  jor  g02826(.dina(n20842), .dinb(n20841), .dout(n20843));
  jand g02827(.dina(n20843), .dinb(n20761), .dout(n20844));
  jxor g02828(.dina(n20754), .dinb(b3 ), .dout(n20845));
  jnot g02829(.din(n20845), .dout(n20846));
  jor  g02830(.dina(n20846), .dinb(n20844), .dout(n20847));
  jand g02831(.dina(n20847), .dinb(n20755), .dout(n20848));
  jxor g02832(.dina(n20746), .dinb(n337), .dout(n20849));
  jnot g02833(.din(n20849), .dout(n20850));
  jor  g02834(.dina(n20850), .dinb(n20848), .dout(n20851));
  jand g02835(.dina(n20851), .dinb(n20748), .dout(n20852));
  jxor g02836(.dina(n20740), .dinb(n338), .dout(n20853));
  jnot g02837(.din(n20853), .dout(n20854));
  jor  g02838(.dina(n20854), .dinb(n20852), .dout(n20855));
  jand g02839(.dina(n20855), .dinb(n20742), .dout(n20856));
  jxor g02840(.dina(n20734), .dinb(n334), .dout(n20857));
  jnot g02841(.din(n20857), .dout(n20858));
  jor  g02842(.dina(n20858), .dinb(n20856), .dout(n20859));
  jand g02843(.dina(n20859), .dinb(n20736), .dout(n20860));
  jxor g02844(.dina(n20728), .dinb(n335), .dout(n20861));
  jnot g02845(.din(n20861), .dout(n20862));
  jor  g02846(.dina(n20862), .dinb(n20860), .dout(n20863));
  jand g02847(.dina(n20863), .dinb(n20730), .dout(n20864));
  jxor g02848(.dina(n20722), .dinb(n323), .dout(n20865));
  jnot g02849(.din(n20865), .dout(n20866));
  jor  g02850(.dina(n20866), .dinb(n20864), .dout(n20867));
  jand g02851(.dina(n20867), .dinb(n20724), .dout(n20868));
  jxor g02852(.dina(n20716), .dinb(n324), .dout(n20869));
  jnot g02853(.din(n20869), .dout(n20870));
  jor  g02854(.dina(n20870), .dinb(n20868), .dout(n20871));
  jand g02855(.dina(n20871), .dinb(n20718), .dout(n20872));
  jxor g02856(.dina(n20710), .dinb(n325), .dout(n20873));
  jnot g02857(.din(n20873), .dout(n20874));
  jor  g02858(.dina(n20874), .dinb(n20872), .dout(n20875));
  jand g02859(.dina(n20875), .dinb(n20712), .dout(n20876));
  jxor g02860(.dina(n20704), .dinb(n439), .dout(n20877));
  jnot g02861(.din(n20877), .dout(n20878));
  jor  g02862(.dina(n20878), .dinb(n20876), .dout(n20879));
  jand g02863(.dina(n20879), .dinb(n20706), .dout(n20880));
  jxor g02864(.dina(n20698), .dinb(n440), .dout(n20881));
  jnot g02865(.din(n20881), .dout(n20882));
  jor  g02866(.dina(n20882), .dinb(n20880), .dout(n20883));
  jand g02867(.dina(n20883), .dinb(n20700), .dout(n20884));
  jxor g02868(.dina(n20692), .dinb(n435), .dout(n20885));
  jnot g02869(.din(n20885), .dout(n20886));
  jor  g02870(.dina(n20886), .dinb(n20884), .dout(n20887));
  jand g02871(.dina(n20887), .dinb(n20694), .dout(n20888));
  jxor g02872(.dina(n20686), .dinb(n436), .dout(n20889));
  jnot g02873(.din(n20889), .dout(n20890));
  jor  g02874(.dina(n20890), .dinb(n20888), .dout(n20891));
  jand g02875(.dina(n20891), .dinb(n20688), .dout(n20892));
  jxor g02876(.dina(n20680), .dinb(n432), .dout(n20893));
  jnot g02877(.din(n20893), .dout(n20894));
  jor  g02878(.dina(n20894), .dinb(n20892), .dout(n20895));
  jand g02879(.dina(n20895), .dinb(n20682), .dout(n20896));
  jxor g02880(.dina(n20674), .dinb(n433), .dout(n20897));
  jnot g02881(.din(n20897), .dout(n20898));
  jor  g02882(.dina(n20898), .dinb(n20896), .dout(n20899));
  jand g02883(.dina(n20899), .dinb(n20676), .dout(n20900));
  jxor g02884(.dina(n20668), .dinb(n421), .dout(n20901));
  jnot g02885(.din(n20901), .dout(n20902));
  jor  g02886(.dina(n20902), .dinb(n20900), .dout(n20903));
  jand g02887(.dina(n20903), .dinb(n20670), .dout(n20904));
  jxor g02888(.dina(n20662), .dinb(n422), .dout(n20905));
  jnot g02889(.din(n20905), .dout(n20906));
  jor  g02890(.dina(n20906), .dinb(n20904), .dout(n20907));
  jand g02891(.dina(n20907), .dinb(n20664), .dout(n20908));
  jnot g02892(.din(n20656), .dout(n20909));
  jand g02893(.dina(n20909), .dinb(b19 ), .dout(n20910));
  jor  g02894(.dina(n20910), .dinb(n20908), .dout(n20911));
  jand g02895(.dina(n20911), .dinb(n20658), .dout(n20912));
  jor  g02896(.dina(n20912), .dinb(n318), .dout(n20913));
  jand g02897(.dina(n20913), .dinb(n20656), .dout(n20914));
  jnot g02898(.din(n1972), .dout(n20917));
  jor  g02899(.dina(n20835), .dinb(n20917), .dout(n20918));
  jand g02900(.dina(n20918), .dinb(a45 ), .dout(n20919));
  jor  g02901(.dina(n2293), .dinb(n20919), .dout(n20921));
  jand g02902(.dina(n20921), .dinb(n258), .dout(n20922));
  jxor g02903(.dina(n20837), .dinb(b1 ), .dout(n20923));
  jand g02904(.dina(n20923), .dinb(n2300), .dout(n20924));
  jor  g02905(.dina(n20924), .dinb(n20922), .dout(n20925));
  jxor g02906(.dina(n20760), .dinb(b2 ), .dout(n20926));
  jand g02907(.dina(n20926), .dinb(n20925), .dout(n20927));
  jor  g02908(.dina(n20927), .dinb(n2289), .dout(n20928));
  jand g02909(.dina(n20845), .dinb(n20928), .dout(n20929));
  jor  g02910(.dina(n20929), .dinb(n2284), .dout(n20930));
  jand g02911(.dina(n20849), .dinb(n20930), .dout(n20931));
  jor  g02912(.dina(n20931), .dinb(n20747), .dout(n20932));
  jand g02913(.dina(n20853), .dinb(n20932), .dout(n20933));
  jor  g02914(.dina(n20933), .dinb(n20741), .dout(n20934));
  jand g02915(.dina(n20857), .dinb(n20934), .dout(n20935));
  jor  g02916(.dina(n20935), .dinb(n20735), .dout(n20936));
  jand g02917(.dina(n20861), .dinb(n20936), .dout(n20937));
  jor  g02918(.dina(n20937), .dinb(n20729), .dout(n20938));
  jand g02919(.dina(n20865), .dinb(n20938), .dout(n20939));
  jor  g02920(.dina(n20939), .dinb(n20723), .dout(n20940));
  jand g02921(.dina(n20869), .dinb(n20940), .dout(n20941));
  jor  g02922(.dina(n20941), .dinb(n20717), .dout(n20942));
  jand g02923(.dina(n20873), .dinb(n20942), .dout(n20943));
  jor  g02924(.dina(n20943), .dinb(n20711), .dout(n20944));
  jand g02925(.dina(n20877), .dinb(n20944), .dout(n20945));
  jor  g02926(.dina(n20945), .dinb(n20705), .dout(n20946));
  jand g02927(.dina(n20881), .dinb(n20946), .dout(n20947));
  jor  g02928(.dina(n20947), .dinb(n20699), .dout(n20948));
  jand g02929(.dina(n20885), .dinb(n20948), .dout(n20949));
  jor  g02930(.dina(n20949), .dinb(n20693), .dout(n20950));
  jand g02931(.dina(n20889), .dinb(n20950), .dout(n20951));
  jor  g02932(.dina(n20951), .dinb(n20687), .dout(n20952));
  jand g02933(.dina(n20893), .dinb(n20952), .dout(n20953));
  jor  g02934(.dina(n20953), .dinb(n20681), .dout(n20954));
  jand g02935(.dina(n20897), .dinb(n20954), .dout(n20955));
  jor  g02936(.dina(n20955), .dinb(n20675), .dout(n20956));
  jand g02937(.dina(n20901), .dinb(n20956), .dout(n20957));
  jor  g02938(.dina(n20957), .dinb(n20669), .dout(n20958));
  jand g02939(.dina(n20905), .dinb(n20958), .dout(n20959));
  jor  g02940(.dina(n20959), .dinb(n20663), .dout(n20960));
  jand g02941(.dina(n20657), .dinb(n1970), .dout(n20961));
  jand g02942(.dina(n20961), .dinb(n20960), .dout(n20962));
  jor  g02943(.dina(n20962), .dinb(n20914), .dout(n20963));
  jnot g02944(.din(n20963), .dout(n20964));
  jand g02945(.dina(n20913), .dinb(n20662), .dout(n20965));
  jnot g02946(.din(n20910), .dout(n20966));
  jand g02947(.dina(n20966), .dinb(n20960), .dout(n20967));
  jor  g02948(.dina(n20967), .dinb(n20657), .dout(n20968));
  jand g02949(.dina(n20968), .dinb(n1970), .dout(n20969));
  jxor g02950(.dina(n20905), .dinb(n20958), .dout(n20970));
  jand g02951(.dina(n20970), .dinb(n20969), .dout(n20971));
  jor  g02952(.dina(n20971), .dinb(n20965), .dout(n20972));
  jand g02953(.dina(n20972), .dinb(n416), .dout(n20973));
  jnot g02954(.din(n20973), .dout(n20974));
  jand g02955(.dina(n20913), .dinb(n20668), .dout(n20975));
  jxor g02956(.dina(n20901), .dinb(n20956), .dout(n20976));
  jand g02957(.dina(n20976), .dinb(n20969), .dout(n20977));
  jor  g02958(.dina(n20977), .dinb(n20975), .dout(n20978));
  jand g02959(.dina(n20978), .dinb(n422), .dout(n20979));
  jnot g02960(.din(n20979), .dout(n20980));
  jand g02961(.dina(n20913), .dinb(n20674), .dout(n20981));
  jxor g02962(.dina(n20897), .dinb(n20954), .dout(n20982));
  jand g02963(.dina(n20982), .dinb(n20969), .dout(n20983));
  jor  g02964(.dina(n20983), .dinb(n20981), .dout(n20984));
  jand g02965(.dina(n20984), .dinb(n421), .dout(n20985));
  jnot g02966(.din(n20985), .dout(n20986));
  jand g02967(.dina(n20913), .dinb(n20680), .dout(n20987));
  jxor g02968(.dina(n20893), .dinb(n20952), .dout(n20988));
  jand g02969(.dina(n20988), .dinb(n20969), .dout(n20989));
  jor  g02970(.dina(n20989), .dinb(n20987), .dout(n20990));
  jand g02971(.dina(n20990), .dinb(n433), .dout(n20991));
  jnot g02972(.din(n20991), .dout(n20992));
  jand g02973(.dina(n20913), .dinb(n20686), .dout(n20993));
  jxor g02974(.dina(n20889), .dinb(n20950), .dout(n20994));
  jand g02975(.dina(n20994), .dinb(n20969), .dout(n20995));
  jor  g02976(.dina(n20995), .dinb(n20993), .dout(n20996));
  jand g02977(.dina(n20996), .dinb(n432), .dout(n20997));
  jnot g02978(.din(n20997), .dout(n20998));
  jand g02979(.dina(n20913), .dinb(n20692), .dout(n20999));
  jxor g02980(.dina(n20885), .dinb(n20948), .dout(n21000));
  jand g02981(.dina(n21000), .dinb(n20969), .dout(n21001));
  jor  g02982(.dina(n21001), .dinb(n20999), .dout(n21002));
  jand g02983(.dina(n21002), .dinb(n436), .dout(n21003));
  jnot g02984(.din(n21003), .dout(n21004));
  jand g02985(.dina(n20913), .dinb(n20698), .dout(n21005));
  jxor g02986(.dina(n20881), .dinb(n20946), .dout(n21006));
  jand g02987(.dina(n21006), .dinb(n20969), .dout(n21007));
  jor  g02988(.dina(n21007), .dinb(n21005), .dout(n21008));
  jand g02989(.dina(n21008), .dinb(n435), .dout(n21009));
  jnot g02990(.din(n21009), .dout(n21010));
  jand g02991(.dina(n20913), .dinb(n20704), .dout(n21011));
  jxor g02992(.dina(n20877), .dinb(n20944), .dout(n21012));
  jand g02993(.dina(n21012), .dinb(n20969), .dout(n21013));
  jor  g02994(.dina(n21013), .dinb(n21011), .dout(n21014));
  jand g02995(.dina(n21014), .dinb(n440), .dout(n21015));
  jnot g02996(.din(n21015), .dout(n21016));
  jand g02997(.dina(n20913), .dinb(n20710), .dout(n21017));
  jxor g02998(.dina(n20873), .dinb(n20942), .dout(n21018));
  jand g02999(.dina(n21018), .dinb(n20969), .dout(n21019));
  jor  g03000(.dina(n21019), .dinb(n21017), .dout(n21020));
  jand g03001(.dina(n21020), .dinb(n439), .dout(n21021));
  jnot g03002(.din(n21021), .dout(n21022));
  jand g03003(.dina(n20913), .dinb(n20716), .dout(n21023));
  jxor g03004(.dina(n20869), .dinb(n20940), .dout(n21024));
  jand g03005(.dina(n21024), .dinb(n20969), .dout(n21025));
  jor  g03006(.dina(n21025), .dinb(n21023), .dout(n21026));
  jand g03007(.dina(n21026), .dinb(n325), .dout(n21027));
  jnot g03008(.din(n21027), .dout(n21028));
  jand g03009(.dina(n20913), .dinb(n20722), .dout(n21029));
  jxor g03010(.dina(n20865), .dinb(n20938), .dout(n21030));
  jand g03011(.dina(n21030), .dinb(n20969), .dout(n21031));
  jor  g03012(.dina(n21031), .dinb(n21029), .dout(n21032));
  jand g03013(.dina(n21032), .dinb(n324), .dout(n21033));
  jnot g03014(.din(n21033), .dout(n21034));
  jand g03015(.dina(n20913), .dinb(n20728), .dout(n21035));
  jxor g03016(.dina(n20861), .dinb(n20936), .dout(n21036));
  jand g03017(.dina(n21036), .dinb(n20969), .dout(n21037));
  jor  g03018(.dina(n21037), .dinb(n21035), .dout(n21038));
  jand g03019(.dina(n21038), .dinb(n323), .dout(n21039));
  jnot g03020(.din(n21039), .dout(n21040));
  jand g03021(.dina(n20913), .dinb(n20734), .dout(n21041));
  jxor g03022(.dina(n20857), .dinb(n20934), .dout(n21042));
  jand g03023(.dina(n21042), .dinb(n20969), .dout(n21043));
  jor  g03024(.dina(n21043), .dinb(n21041), .dout(n21044));
  jand g03025(.dina(n21044), .dinb(n335), .dout(n21045));
  jnot g03026(.din(n21045), .dout(n21046));
  jand g03027(.dina(n20913), .dinb(n20740), .dout(n21047));
  jxor g03028(.dina(n20853), .dinb(n20932), .dout(n21048));
  jand g03029(.dina(n21048), .dinb(n20969), .dout(n21049));
  jor  g03030(.dina(n21049), .dinb(n21047), .dout(n21050));
  jand g03031(.dina(n21050), .dinb(n334), .dout(n21051));
  jnot g03032(.din(n21051), .dout(n21052));
  jand g03033(.dina(n20913), .dinb(n20746), .dout(n21053));
  jxor g03034(.dina(n20849), .dinb(n20930), .dout(n21054));
  jand g03035(.dina(n21054), .dinb(n20969), .dout(n21055));
  jor  g03036(.dina(n21055), .dinb(n21053), .dout(n21056));
  jand g03037(.dina(n21056), .dinb(n338), .dout(n21057));
  jnot g03038(.din(n21057), .dout(n21058));
  jor  g03039(.dina(n20969), .dinb(n20754), .dout(n21059));
  jxor g03040(.dina(n20845), .dinb(n20928), .dout(n21060));
  jand g03041(.dina(n21060), .dinb(n20969), .dout(n21061));
  jnot g03042(.din(n21061), .dout(n21062));
  jand g03043(.dina(n21062), .dinb(n21059), .dout(n21063));
  jnot g03044(.din(n2446), .dout(n21066));
  jor  g03045(.dina(n20969), .dinb(n20760), .dout(n21067));
  jxor g03046(.dina(n20926), .dinb(n20925), .dout(n21068));
  jnot g03047(.din(n21068), .dout(n21069));
  jor  g03048(.dina(n21069), .dinb(n20913), .dout(n21070));
  jand g03049(.dina(n21070), .dinb(n21067), .dout(n21071));
  jnot g03050(.din(n21071), .dout(n21072));
  jand g03051(.dina(n21072), .dinb(n344), .dout(n21073));
  jnot g03052(.din(n21073), .dout(n21074));
  jand g03053(.dina(n20913), .dinb(n20921), .dout(n21075));
  jxor g03054(.dina(n20923), .dinb(n2300), .dout(n21076));
  jand g03055(.dina(n21076), .dinb(n20969), .dout(n21077));
  jor  g03056(.dina(n21077), .dinb(n21075), .dout(n21078));
  jand g03057(.dina(n21078), .dinb(n348), .dout(n21079));
  jnot g03058(.din(n21079), .dout(n21080));
  jnot g03059(.din(n2461), .dout(n21081));
  jor  g03060(.dina(n20912), .dinb(n21081), .dout(n21082));
  jand g03061(.dina(n21082), .dinb(a44 ), .dout(n21083));
  jand g03062(.dina(n20969), .dinb(n2299), .dout(n21084));
  jor  g03063(.dina(n21084), .dinb(n21083), .dout(n21085));
  jand g03064(.dina(n21085), .dinb(n258), .dout(n21086));
  jand g03065(.dina(n20968), .dinb(n2461), .dout(n21088));
  jor  g03066(.dina(n21088), .dinb(n2298), .dout(n21089));
  jor  g03067(.dina(n20913), .dinb(n2300), .dout(n21090));
  jand g03068(.dina(n21090), .dinb(n21089), .dout(n21091));
  jxor g03069(.dina(n21091), .dinb(n258), .dout(n21092));
  jor  g03070(.dina(n21092), .dinb(n2471), .dout(n21093));
  jand g03071(.dina(n21093), .dinb(n2468), .dout(n21094));
  jxor g03072(.dina(n21078), .dinb(n348), .dout(n21095));
  jnot g03073(.din(n21095), .dout(n21096));
  jor  g03074(.dina(n21096), .dinb(n21094), .dout(n21097));
  jand g03075(.dina(n21097), .dinb(n21080), .dout(n21098));
  jxor g03076(.dina(n21071), .dinb(b3 ), .dout(n21099));
  jnot g03077(.din(n21099), .dout(n21100));
  jor  g03078(.dina(n21100), .dinb(n21098), .dout(n21101));
  jand g03079(.dina(n21101), .dinb(n21074), .dout(n21102));
  jxor g03080(.dina(n21063), .dinb(b4 ), .dout(n21103));
  jnot g03081(.din(n21103), .dout(n21104));
  jor  g03082(.dina(n21104), .dinb(n21102), .dout(n21105));
  jand g03083(.dina(n21105), .dinb(n21066), .dout(n21106));
  jxor g03084(.dina(n21056), .dinb(n338), .dout(n21107));
  jnot g03085(.din(n21107), .dout(n21108));
  jor  g03086(.dina(n21108), .dinb(n21106), .dout(n21109));
  jand g03087(.dina(n21109), .dinb(n21058), .dout(n21110));
  jxor g03088(.dina(n21050), .dinb(n334), .dout(n21111));
  jnot g03089(.din(n21111), .dout(n21112));
  jor  g03090(.dina(n21112), .dinb(n21110), .dout(n21113));
  jand g03091(.dina(n21113), .dinb(n21052), .dout(n21114));
  jxor g03092(.dina(n21044), .dinb(n335), .dout(n21115));
  jnot g03093(.din(n21115), .dout(n21116));
  jor  g03094(.dina(n21116), .dinb(n21114), .dout(n21117));
  jand g03095(.dina(n21117), .dinb(n21046), .dout(n21118));
  jxor g03096(.dina(n21038), .dinb(n323), .dout(n21119));
  jnot g03097(.din(n21119), .dout(n21120));
  jor  g03098(.dina(n21120), .dinb(n21118), .dout(n21121));
  jand g03099(.dina(n21121), .dinb(n21040), .dout(n21122));
  jxor g03100(.dina(n21032), .dinb(n324), .dout(n21123));
  jnot g03101(.din(n21123), .dout(n21124));
  jor  g03102(.dina(n21124), .dinb(n21122), .dout(n21125));
  jand g03103(.dina(n21125), .dinb(n21034), .dout(n21126));
  jxor g03104(.dina(n21026), .dinb(n325), .dout(n21127));
  jnot g03105(.din(n21127), .dout(n21128));
  jor  g03106(.dina(n21128), .dinb(n21126), .dout(n21129));
  jand g03107(.dina(n21129), .dinb(n21028), .dout(n21130));
  jxor g03108(.dina(n21020), .dinb(n439), .dout(n21131));
  jnot g03109(.din(n21131), .dout(n21132));
  jor  g03110(.dina(n21132), .dinb(n21130), .dout(n21133));
  jand g03111(.dina(n21133), .dinb(n21022), .dout(n21134));
  jxor g03112(.dina(n21014), .dinb(n440), .dout(n21135));
  jnot g03113(.din(n21135), .dout(n21136));
  jor  g03114(.dina(n21136), .dinb(n21134), .dout(n21137));
  jand g03115(.dina(n21137), .dinb(n21016), .dout(n21138));
  jxor g03116(.dina(n21008), .dinb(n435), .dout(n21139));
  jnot g03117(.din(n21139), .dout(n21140));
  jor  g03118(.dina(n21140), .dinb(n21138), .dout(n21141));
  jand g03119(.dina(n21141), .dinb(n21010), .dout(n21142));
  jxor g03120(.dina(n21002), .dinb(n436), .dout(n21143));
  jnot g03121(.din(n21143), .dout(n21144));
  jor  g03122(.dina(n21144), .dinb(n21142), .dout(n21145));
  jand g03123(.dina(n21145), .dinb(n21004), .dout(n21146));
  jxor g03124(.dina(n20996), .dinb(n432), .dout(n21147));
  jnot g03125(.din(n21147), .dout(n21148));
  jor  g03126(.dina(n21148), .dinb(n21146), .dout(n21149));
  jand g03127(.dina(n21149), .dinb(n20998), .dout(n21150));
  jxor g03128(.dina(n20990), .dinb(n433), .dout(n21151));
  jnot g03129(.din(n21151), .dout(n21152));
  jor  g03130(.dina(n21152), .dinb(n21150), .dout(n21153));
  jand g03131(.dina(n21153), .dinb(n20992), .dout(n21154));
  jxor g03132(.dina(n20984), .dinb(n421), .dout(n21155));
  jnot g03133(.din(n21155), .dout(n21156));
  jor  g03134(.dina(n21156), .dinb(n21154), .dout(n21157));
  jand g03135(.dina(n21157), .dinb(n20986), .dout(n21158));
  jxor g03136(.dina(n20978), .dinb(n422), .dout(n21159));
  jnot g03137(.din(n21159), .dout(n21160));
  jor  g03138(.dina(n21160), .dinb(n21158), .dout(n21161));
  jand g03139(.dina(n21161), .dinb(n20980), .dout(n21162));
  jxor g03140(.dina(n20972), .dinb(n416), .dout(n21163));
  jnot g03141(.din(n21163), .dout(n21164));
  jor  g03142(.dina(n21164), .dinb(n21162), .dout(n21165));
  jand g03143(.dina(n21165), .dinb(n20974), .dout(n21166));
  jnot g03144(.din(n551), .dout(n21167));
  jxor g03145(.dina(n20963), .dinb(b20 ), .dout(n21168));
  jor  g03146(.dina(n21168), .dinb(n21167), .dout(n21169));
  jor  g03147(.dina(n21169), .dinb(n21166), .dout(n21170));
  jand g03148(.dina(n21170), .dinb(n20964), .dout(n21171));
  jxor g03149(.dina(n21091), .dinb(b1 ), .dout(n21172));
  jand g03150(.dina(n21172), .dinb(n2472), .dout(n21173));
  jor  g03151(.dina(n21173), .dinb(n21086), .dout(n21174));
  jand g03152(.dina(n21095), .dinb(n21174), .dout(n21175));
  jor  g03153(.dina(n21175), .dinb(n21079), .dout(n21176));
  jand g03154(.dina(n21099), .dinb(n21176), .dout(n21177));
  jor  g03155(.dina(n21177), .dinb(n21073), .dout(n21178));
  jand g03156(.dina(n21103), .dinb(n21178), .dout(n21179));
  jor  g03157(.dina(n21179), .dinb(n2446), .dout(n21180));
  jand g03158(.dina(n21107), .dinb(n21180), .dout(n21181));
  jor  g03159(.dina(n21181), .dinb(n21057), .dout(n21182));
  jand g03160(.dina(n21111), .dinb(n21182), .dout(n21183));
  jor  g03161(.dina(n21183), .dinb(n21051), .dout(n21184));
  jand g03162(.dina(n21115), .dinb(n21184), .dout(n21185));
  jor  g03163(.dina(n21185), .dinb(n21045), .dout(n21186));
  jand g03164(.dina(n21119), .dinb(n21186), .dout(n21187));
  jor  g03165(.dina(n21187), .dinb(n21039), .dout(n21188));
  jand g03166(.dina(n21123), .dinb(n21188), .dout(n21189));
  jor  g03167(.dina(n21189), .dinb(n21033), .dout(n21190));
  jand g03168(.dina(n21127), .dinb(n21190), .dout(n21191));
  jor  g03169(.dina(n21191), .dinb(n21027), .dout(n21192));
  jand g03170(.dina(n21131), .dinb(n21192), .dout(n21193));
  jor  g03171(.dina(n21193), .dinb(n21021), .dout(n21194));
  jand g03172(.dina(n21135), .dinb(n21194), .dout(n21195));
  jor  g03173(.dina(n21195), .dinb(n21015), .dout(n21196));
  jand g03174(.dina(n21139), .dinb(n21196), .dout(n21197));
  jor  g03175(.dina(n21197), .dinb(n21009), .dout(n21198));
  jand g03176(.dina(n21143), .dinb(n21198), .dout(n21199));
  jor  g03177(.dina(n21199), .dinb(n21003), .dout(n21200));
  jand g03178(.dina(n21147), .dinb(n21200), .dout(n21201));
  jor  g03179(.dina(n21201), .dinb(n20997), .dout(n21202));
  jand g03180(.dina(n21151), .dinb(n21202), .dout(n21203));
  jor  g03181(.dina(n21203), .dinb(n20991), .dout(n21204));
  jand g03182(.dina(n21155), .dinb(n21204), .dout(n21205));
  jor  g03183(.dina(n21205), .dinb(n20985), .dout(n21206));
  jand g03184(.dina(n21159), .dinb(n21206), .dout(n21207));
  jor  g03185(.dina(n21207), .dinb(n20979), .dout(n21208));
  jand g03186(.dina(n21163), .dinb(n21208), .dout(n21209));
  jor  g03187(.dina(n21209), .dinb(n20973), .dout(n21210));
  jnot g03188(.din(n21169), .dout(n21211));
  jand g03189(.dina(n21211), .dinb(n21210), .dout(n21212));
  jand g03190(.dina(n20963), .dinb(n1970), .dout(n21213));
  jor  g03191(.dina(n21213), .dinb(n21212), .dout(n21214));
  jxor g03192(.dina(n21168), .dinb(n21210), .dout(n21215));
  jand g03193(.dina(n21215), .dinb(n21214), .dout(n21216));
  jor  g03194(.dina(n21216), .dinb(n21171), .dout(n21217));
  jnot g03195(.din(n21217), .dout(n21218));
  jand g03196(.dina(n21217), .dinb(b21 ), .dout(n21219));
  jnot g03197(.din(n21219), .dout(n21220));
  jand g03198(.dina(n21218), .dinb(n2547), .dout(n21221));
  jnot g03199(.din(n21213), .dout(n21222));
  jand g03200(.dina(n21222), .dinb(n21170), .dout(n21223));
  jand g03201(.dina(n21223), .dinb(n20972), .dout(n21224));
  jxor g03202(.dina(n21163), .dinb(n21208), .dout(n21225));
  jand g03203(.dina(n21225), .dinb(n21214), .dout(n21226));
  jor  g03204(.dina(n21226), .dinb(n21224), .dout(n21227));
  jand g03205(.dina(n21227), .dinb(n417), .dout(n21228));
  jand g03206(.dina(n21223), .dinb(n20978), .dout(n21229));
  jxor g03207(.dina(n21159), .dinb(n21206), .dout(n21230));
  jand g03208(.dina(n21230), .dinb(n21214), .dout(n21231));
  jor  g03209(.dina(n21231), .dinb(n21229), .dout(n21232));
  jand g03210(.dina(n21232), .dinb(n416), .dout(n21233));
  jand g03211(.dina(n21223), .dinb(n20984), .dout(n21234));
  jxor g03212(.dina(n21155), .dinb(n21204), .dout(n21235));
  jand g03213(.dina(n21235), .dinb(n21214), .dout(n21236));
  jor  g03214(.dina(n21236), .dinb(n21234), .dout(n21237));
  jand g03215(.dina(n21237), .dinb(n422), .dout(n21238));
  jand g03216(.dina(n21223), .dinb(n20990), .dout(n21239));
  jxor g03217(.dina(n21151), .dinb(n21202), .dout(n21240));
  jand g03218(.dina(n21240), .dinb(n21214), .dout(n21241));
  jor  g03219(.dina(n21241), .dinb(n21239), .dout(n21242));
  jand g03220(.dina(n21242), .dinb(n421), .dout(n21243));
  jand g03221(.dina(n21223), .dinb(n20996), .dout(n21244));
  jxor g03222(.dina(n21147), .dinb(n21200), .dout(n21245));
  jand g03223(.dina(n21245), .dinb(n21214), .dout(n21246));
  jor  g03224(.dina(n21246), .dinb(n21244), .dout(n21247));
  jand g03225(.dina(n21247), .dinb(n433), .dout(n21248));
  jand g03226(.dina(n21223), .dinb(n21002), .dout(n21249));
  jxor g03227(.dina(n21143), .dinb(n21198), .dout(n21250));
  jand g03228(.dina(n21250), .dinb(n21214), .dout(n21251));
  jor  g03229(.dina(n21251), .dinb(n21249), .dout(n21252));
  jand g03230(.dina(n21252), .dinb(n432), .dout(n21253));
  jand g03231(.dina(n21223), .dinb(n21008), .dout(n21254));
  jxor g03232(.dina(n21139), .dinb(n21196), .dout(n21255));
  jand g03233(.dina(n21255), .dinb(n21214), .dout(n21256));
  jor  g03234(.dina(n21256), .dinb(n21254), .dout(n21257));
  jand g03235(.dina(n21257), .dinb(n436), .dout(n21258));
  jand g03236(.dina(n21223), .dinb(n21014), .dout(n21259));
  jxor g03237(.dina(n21135), .dinb(n21194), .dout(n21260));
  jand g03238(.dina(n21260), .dinb(n21214), .dout(n21261));
  jor  g03239(.dina(n21261), .dinb(n21259), .dout(n21262));
  jand g03240(.dina(n21262), .dinb(n435), .dout(n21263));
  jand g03241(.dina(n21223), .dinb(n21020), .dout(n21264));
  jxor g03242(.dina(n21131), .dinb(n21192), .dout(n21265));
  jand g03243(.dina(n21265), .dinb(n21214), .dout(n21266));
  jor  g03244(.dina(n21266), .dinb(n21264), .dout(n21267));
  jand g03245(.dina(n21267), .dinb(n440), .dout(n21268));
  jand g03246(.dina(n21223), .dinb(n21026), .dout(n21269));
  jxor g03247(.dina(n21127), .dinb(n21190), .dout(n21270));
  jand g03248(.dina(n21270), .dinb(n21214), .dout(n21271));
  jor  g03249(.dina(n21271), .dinb(n21269), .dout(n21272));
  jand g03250(.dina(n21272), .dinb(n439), .dout(n21273));
  jand g03251(.dina(n21223), .dinb(n21032), .dout(n21274));
  jxor g03252(.dina(n21123), .dinb(n21188), .dout(n21275));
  jand g03253(.dina(n21275), .dinb(n21214), .dout(n21276));
  jor  g03254(.dina(n21276), .dinb(n21274), .dout(n21277));
  jand g03255(.dina(n21277), .dinb(n325), .dout(n21278));
  jand g03256(.dina(n21223), .dinb(n21038), .dout(n21279));
  jxor g03257(.dina(n21119), .dinb(n21186), .dout(n21280));
  jand g03258(.dina(n21280), .dinb(n21214), .dout(n21281));
  jor  g03259(.dina(n21281), .dinb(n21279), .dout(n21282));
  jand g03260(.dina(n21282), .dinb(n324), .dout(n21283));
  jand g03261(.dina(n21223), .dinb(n21044), .dout(n21284));
  jxor g03262(.dina(n21115), .dinb(n21184), .dout(n21285));
  jand g03263(.dina(n21285), .dinb(n21214), .dout(n21286));
  jor  g03264(.dina(n21286), .dinb(n21284), .dout(n21287));
  jand g03265(.dina(n21287), .dinb(n323), .dout(n21288));
  jand g03266(.dina(n21223), .dinb(n21050), .dout(n21289));
  jxor g03267(.dina(n21111), .dinb(n21182), .dout(n21290));
  jand g03268(.dina(n21290), .dinb(n21214), .dout(n21291));
  jor  g03269(.dina(n21291), .dinb(n21289), .dout(n21292));
  jand g03270(.dina(n21292), .dinb(n335), .dout(n21293));
  jand g03271(.dina(n21223), .dinb(n21056), .dout(n21294));
  jxor g03272(.dina(n21107), .dinb(n21180), .dout(n21295));
  jand g03273(.dina(n21295), .dinb(n21214), .dout(n21296));
  jor  g03274(.dina(n21296), .dinb(n21294), .dout(n21297));
  jand g03275(.dina(n21297), .dinb(n334), .dout(n21298));
  jand g03276(.dina(n21223), .dinb(n2445), .dout(n21299));
  jxor g03277(.dina(n21103), .dinb(n21178), .dout(n21300));
  jand g03278(.dina(n21300), .dinb(n21214), .dout(n21301));
  jor  g03279(.dina(n21301), .dinb(n21299), .dout(n21302));
  jand g03280(.dina(n21302), .dinb(n338), .dout(n21303));
  jand g03281(.dina(n21223), .dinb(n21072), .dout(n21304));
  jxor g03282(.dina(n21099), .dinb(n21176), .dout(n21305));
  jand g03283(.dina(n21305), .dinb(n21214), .dout(n21306));
  jor  g03284(.dina(n21306), .dinb(n21304), .dout(n21307));
  jand g03285(.dina(n21307), .dinb(n337), .dout(n21308));
  jand g03286(.dina(n21223), .dinb(n21078), .dout(n21309));
  jxor g03287(.dina(n21095), .dinb(n21174), .dout(n21310));
  jand g03288(.dina(n21310), .dinb(n21214), .dout(n21311));
  jor  g03289(.dina(n21311), .dinb(n21309), .dout(n21312));
  jand g03290(.dina(n21312), .dinb(n344), .dout(n21313));
  jand g03291(.dina(n21223), .dinb(n21085), .dout(n21314));
  jxor g03292(.dina(n21172), .dinb(n2472), .dout(n21315));
  jand g03293(.dina(n21315), .dinb(n21214), .dout(n21316));
  jor  g03294(.dina(n21316), .dinb(n21314), .dout(n21317));
  jand g03295(.dina(n21317), .dinb(n348), .dout(n21318));
  jor  g03296(.dina(n21223), .dinb(n18364), .dout(n21319));
  jand g03297(.dina(n21319), .dinb(a43 ), .dout(n21320));
  jor  g03298(.dina(n21223), .dinb(n2472), .dout(n21321));
  jnot g03299(.din(n21321), .dout(n21322));
  jor  g03300(.dina(n21322), .dinb(n21320), .dout(n21323));
  jand g03301(.dina(n21323), .dinb(n258), .dout(n21324));
  jand g03302(.dina(n21214), .dinb(b0 ), .dout(n21325));
  jor  g03303(.dina(n21325), .dinb(n2470), .dout(n21326));
  jand g03304(.dina(n21321), .dinb(n21326), .dout(n21327));
  jxor g03305(.dina(n21327), .dinb(b1 ), .dout(n21328));
  jand g03306(.dina(n21328), .dinb(n2651), .dout(n21329));
  jor  g03307(.dina(n21329), .dinb(n21324), .dout(n21330));
  jxor g03308(.dina(n21317), .dinb(n348), .dout(n21331));
  jand g03309(.dina(n21331), .dinb(n21330), .dout(n21332));
  jor  g03310(.dina(n21332), .dinb(n21318), .dout(n21333));
  jxor g03311(.dina(n21312), .dinb(n344), .dout(n21334));
  jand g03312(.dina(n21334), .dinb(n21333), .dout(n21335));
  jor  g03313(.dina(n21335), .dinb(n21313), .dout(n21336));
  jxor g03314(.dina(n21307), .dinb(n337), .dout(n21337));
  jand g03315(.dina(n21337), .dinb(n21336), .dout(n21338));
  jor  g03316(.dina(n21338), .dinb(n21308), .dout(n21339));
  jxor g03317(.dina(n21302), .dinb(n338), .dout(n21340));
  jand g03318(.dina(n21340), .dinb(n21339), .dout(n21341));
  jor  g03319(.dina(n21341), .dinb(n21303), .dout(n21342));
  jxor g03320(.dina(n21297), .dinb(n334), .dout(n21343));
  jand g03321(.dina(n21343), .dinb(n21342), .dout(n21344));
  jor  g03322(.dina(n21344), .dinb(n21298), .dout(n21345));
  jxor g03323(.dina(n21292), .dinb(n335), .dout(n21346));
  jand g03324(.dina(n21346), .dinb(n21345), .dout(n21347));
  jor  g03325(.dina(n21347), .dinb(n21293), .dout(n21348));
  jxor g03326(.dina(n21287), .dinb(n323), .dout(n21349));
  jand g03327(.dina(n21349), .dinb(n21348), .dout(n21350));
  jor  g03328(.dina(n21350), .dinb(n21288), .dout(n21351));
  jxor g03329(.dina(n21282), .dinb(n324), .dout(n21352));
  jand g03330(.dina(n21352), .dinb(n21351), .dout(n21353));
  jor  g03331(.dina(n21353), .dinb(n21283), .dout(n21354));
  jxor g03332(.dina(n21277), .dinb(n325), .dout(n21355));
  jand g03333(.dina(n21355), .dinb(n21354), .dout(n21356));
  jor  g03334(.dina(n21356), .dinb(n21278), .dout(n21357));
  jxor g03335(.dina(n21272), .dinb(n439), .dout(n21358));
  jand g03336(.dina(n21358), .dinb(n21357), .dout(n21359));
  jor  g03337(.dina(n21359), .dinb(n21273), .dout(n21360));
  jxor g03338(.dina(n21267), .dinb(n440), .dout(n21361));
  jand g03339(.dina(n21361), .dinb(n21360), .dout(n21362));
  jor  g03340(.dina(n21362), .dinb(n21268), .dout(n21363));
  jxor g03341(.dina(n21262), .dinb(n435), .dout(n21364));
  jand g03342(.dina(n21364), .dinb(n21363), .dout(n21365));
  jor  g03343(.dina(n21365), .dinb(n21263), .dout(n21366));
  jxor g03344(.dina(n21257), .dinb(n436), .dout(n21367));
  jand g03345(.dina(n21367), .dinb(n21366), .dout(n21368));
  jor  g03346(.dina(n21368), .dinb(n21258), .dout(n21369));
  jxor g03347(.dina(n21252), .dinb(n432), .dout(n21370));
  jand g03348(.dina(n21370), .dinb(n21369), .dout(n21371));
  jor  g03349(.dina(n21371), .dinb(n21253), .dout(n21372));
  jxor g03350(.dina(n21247), .dinb(n433), .dout(n21373));
  jand g03351(.dina(n21373), .dinb(n21372), .dout(n21374));
  jor  g03352(.dina(n21374), .dinb(n21248), .dout(n21375));
  jxor g03353(.dina(n21242), .dinb(n421), .dout(n21376));
  jand g03354(.dina(n21376), .dinb(n21375), .dout(n21377));
  jor  g03355(.dina(n21377), .dinb(n21243), .dout(n21378));
  jxor g03356(.dina(n21237), .dinb(n422), .dout(n21379));
  jand g03357(.dina(n21379), .dinb(n21378), .dout(n21380));
  jor  g03358(.dina(n21380), .dinb(n21238), .dout(n21381));
  jxor g03359(.dina(n21232), .dinb(n416), .dout(n21382));
  jand g03360(.dina(n21382), .dinb(n21381), .dout(n21383));
  jor  g03361(.dina(n21383), .dinb(n21233), .dout(n21384));
  jxor g03362(.dina(n21227), .dinb(n417), .dout(n21385));
  jand g03363(.dina(n21385), .dinb(n21384), .dout(n21386));
  jor  g03364(.dina(n21386), .dinb(n21228), .dout(n21387));
  jor  g03365(.dina(n21387), .dinb(n21221), .dout(n21388));
  jand g03366(.dina(n21388), .dinb(n21220), .dout(n21389));
  jand g03367(.dina(n21389), .dinb(n2720), .dout(n21390));
  jnot g03368(.din(n21390), .dout(n21391));
  jand g03369(.dina(n21391), .dinb(n21218), .dout(n21392));
  jand g03370(.dina(n21221), .dinb(n2720), .dout(n21393));
  jand g03371(.dina(n21393), .dinb(n21387), .dout(n21394));
  jor  g03372(.dina(n21394), .dinb(n21392), .dout(n21395));
  jand g03373(.dina(n21395), .dinb(n2714), .dout(n21396));
  jnot g03374(.din(n21396), .dout(n21397));
  jand g03375(.dina(n21391), .dinb(n21227), .dout(n21398));
  jxor g03376(.dina(n21385), .dinb(n21384), .dout(n21399));
  jand g03377(.dina(n21399), .dinb(n21390), .dout(n21400));
  jor  g03378(.dina(n21400), .dinb(n21398), .dout(n21401));
  jand g03379(.dina(n21401), .dinb(n2547), .dout(n21402));
  jnot g03380(.din(n21402), .dout(n21403));
  jand g03381(.dina(n21391), .dinb(n21232), .dout(n21404));
  jxor g03382(.dina(n21382), .dinb(n21381), .dout(n21405));
  jand g03383(.dina(n21405), .dinb(n21390), .dout(n21406));
  jor  g03384(.dina(n21406), .dinb(n21404), .dout(n21407));
  jand g03385(.dina(n21407), .dinb(n417), .dout(n21408));
  jnot g03386(.din(n21408), .dout(n21409));
  jand g03387(.dina(n21391), .dinb(n21237), .dout(n21410));
  jxor g03388(.dina(n21379), .dinb(n21378), .dout(n21411));
  jand g03389(.dina(n21411), .dinb(n21390), .dout(n21412));
  jor  g03390(.dina(n21412), .dinb(n21410), .dout(n21413));
  jand g03391(.dina(n21413), .dinb(n416), .dout(n21414));
  jnot g03392(.din(n21414), .dout(n21415));
  jand g03393(.dina(n21391), .dinb(n21242), .dout(n21416));
  jxor g03394(.dina(n21376), .dinb(n21375), .dout(n21417));
  jand g03395(.dina(n21417), .dinb(n21390), .dout(n21418));
  jor  g03396(.dina(n21418), .dinb(n21416), .dout(n21419));
  jand g03397(.dina(n21419), .dinb(n422), .dout(n21420));
  jnot g03398(.din(n21420), .dout(n21421));
  jand g03399(.dina(n21391), .dinb(n21247), .dout(n21422));
  jxor g03400(.dina(n21373), .dinb(n21372), .dout(n21423));
  jand g03401(.dina(n21423), .dinb(n21390), .dout(n21424));
  jor  g03402(.dina(n21424), .dinb(n21422), .dout(n21425));
  jand g03403(.dina(n21425), .dinb(n421), .dout(n21426));
  jnot g03404(.din(n21426), .dout(n21427));
  jand g03405(.dina(n21391), .dinb(n21252), .dout(n21428));
  jxor g03406(.dina(n21370), .dinb(n21369), .dout(n21429));
  jand g03407(.dina(n21429), .dinb(n21390), .dout(n21430));
  jor  g03408(.dina(n21430), .dinb(n21428), .dout(n21431));
  jand g03409(.dina(n21431), .dinb(n433), .dout(n21432));
  jnot g03410(.din(n21432), .dout(n21433));
  jand g03411(.dina(n21391), .dinb(n21257), .dout(n21434));
  jxor g03412(.dina(n21367), .dinb(n21366), .dout(n21435));
  jand g03413(.dina(n21435), .dinb(n21390), .dout(n21436));
  jor  g03414(.dina(n21436), .dinb(n21434), .dout(n21437));
  jand g03415(.dina(n21437), .dinb(n432), .dout(n21438));
  jnot g03416(.din(n21438), .dout(n21439));
  jand g03417(.dina(n21391), .dinb(n21262), .dout(n21440));
  jxor g03418(.dina(n21364), .dinb(n21363), .dout(n21441));
  jand g03419(.dina(n21441), .dinb(n21390), .dout(n21442));
  jor  g03420(.dina(n21442), .dinb(n21440), .dout(n21443));
  jand g03421(.dina(n21443), .dinb(n436), .dout(n21444));
  jnot g03422(.din(n21444), .dout(n21445));
  jand g03423(.dina(n21391), .dinb(n21267), .dout(n21446));
  jxor g03424(.dina(n21361), .dinb(n21360), .dout(n21447));
  jand g03425(.dina(n21447), .dinb(n21390), .dout(n21448));
  jor  g03426(.dina(n21448), .dinb(n21446), .dout(n21449));
  jand g03427(.dina(n21449), .dinb(n435), .dout(n21450));
  jnot g03428(.din(n21450), .dout(n21451));
  jand g03429(.dina(n21391), .dinb(n21272), .dout(n21452));
  jxor g03430(.dina(n21358), .dinb(n21357), .dout(n21453));
  jand g03431(.dina(n21453), .dinb(n21390), .dout(n21454));
  jor  g03432(.dina(n21454), .dinb(n21452), .dout(n21455));
  jand g03433(.dina(n21455), .dinb(n440), .dout(n21456));
  jnot g03434(.din(n21456), .dout(n21457));
  jand g03435(.dina(n21391), .dinb(n21277), .dout(n21458));
  jxor g03436(.dina(n21355), .dinb(n21354), .dout(n21459));
  jand g03437(.dina(n21459), .dinb(n21390), .dout(n21460));
  jor  g03438(.dina(n21460), .dinb(n21458), .dout(n21461));
  jand g03439(.dina(n21461), .dinb(n439), .dout(n21462));
  jnot g03440(.din(n21462), .dout(n21463));
  jand g03441(.dina(n21391), .dinb(n21282), .dout(n21464));
  jxor g03442(.dina(n21352), .dinb(n21351), .dout(n21465));
  jand g03443(.dina(n21465), .dinb(n21390), .dout(n21466));
  jor  g03444(.dina(n21466), .dinb(n21464), .dout(n21467));
  jand g03445(.dina(n21467), .dinb(n325), .dout(n21468));
  jnot g03446(.din(n21468), .dout(n21469));
  jand g03447(.dina(n21391), .dinb(n21287), .dout(n21470));
  jxor g03448(.dina(n21349), .dinb(n21348), .dout(n21471));
  jand g03449(.dina(n21471), .dinb(n21390), .dout(n21472));
  jor  g03450(.dina(n21472), .dinb(n21470), .dout(n21473));
  jand g03451(.dina(n21473), .dinb(n324), .dout(n21474));
  jnot g03452(.din(n21474), .dout(n21475));
  jand g03453(.dina(n21391), .dinb(n21292), .dout(n21476));
  jxor g03454(.dina(n21346), .dinb(n21345), .dout(n21477));
  jand g03455(.dina(n21477), .dinb(n21390), .dout(n21478));
  jor  g03456(.dina(n21478), .dinb(n21476), .dout(n21479));
  jand g03457(.dina(n21479), .dinb(n323), .dout(n21480));
  jnot g03458(.din(n21480), .dout(n21481));
  jand g03459(.dina(n21391), .dinb(n21297), .dout(n21482));
  jxor g03460(.dina(n21343), .dinb(n21342), .dout(n21483));
  jand g03461(.dina(n21483), .dinb(n21390), .dout(n21484));
  jor  g03462(.dina(n21484), .dinb(n21482), .dout(n21485));
  jand g03463(.dina(n21485), .dinb(n335), .dout(n21486));
  jnot g03464(.din(n21486), .dout(n21487));
  jand g03465(.dina(n21391), .dinb(n21302), .dout(n21488));
  jxor g03466(.dina(n21340), .dinb(n21339), .dout(n21489));
  jand g03467(.dina(n21489), .dinb(n21390), .dout(n21490));
  jor  g03468(.dina(n21490), .dinb(n21488), .dout(n21491));
  jand g03469(.dina(n21491), .dinb(n334), .dout(n21492));
  jnot g03470(.din(n21492), .dout(n21493));
  jand g03471(.dina(n21391), .dinb(n21307), .dout(n21494));
  jxor g03472(.dina(n21337), .dinb(n21336), .dout(n21495));
  jand g03473(.dina(n21495), .dinb(n21390), .dout(n21496));
  jor  g03474(.dina(n21496), .dinb(n21494), .dout(n21497));
  jand g03475(.dina(n21497), .dinb(n338), .dout(n21498));
  jnot g03476(.din(n21498), .dout(n21499));
  jand g03477(.dina(n21391), .dinb(n21312), .dout(n21500));
  jxor g03478(.dina(n21334), .dinb(n21333), .dout(n21501));
  jand g03479(.dina(n21501), .dinb(n21390), .dout(n21502));
  jor  g03480(.dina(n21502), .dinb(n21500), .dout(n21503));
  jand g03481(.dina(n21503), .dinb(n337), .dout(n21504));
  jnot g03482(.din(n21504), .dout(n21505));
  jnot g03483(.din(n21317), .dout(n21506));
  jor  g03484(.dina(n21390), .dinb(n21506), .dout(n21507));
  jxor g03485(.dina(n21331), .dinb(n21330), .dout(n21508));
  jnot g03486(.din(n21508), .dout(n21509));
  jor  g03487(.dina(n21509), .dinb(n21391), .dout(n21510));
  jand g03488(.dina(n21510), .dinb(n21507), .dout(n21511));
  jor  g03489(.dina(n21511), .dinb(b3 ), .dout(n21512));
  jor  g03490(.dina(n21390), .dinb(n21327), .dout(n21513));
  jxor g03491(.dina(n21328), .dinb(n2651), .dout(n21514));
  jand g03492(.dina(n21514), .dinb(n21390), .dout(n21515));
  jnot g03493(.din(n21515), .dout(n21516));
  jand g03494(.dina(n21516), .dinb(n21513), .dout(n21517));
  jor  g03495(.dina(n21517), .dinb(b2 ), .dout(n21518));
  jand g03496(.dina(n21389), .dinb(n2852), .dout(n21519));
  jor  g03497(.dina(n21519), .dinb(n2649), .dout(n21520));
  jnot g03498(.din(n2855), .dout(n21521));
  jnot g03499(.din(n21221), .dout(n21522));
  jnot g03500(.din(n21228), .dout(n21523));
  jnot g03501(.din(n21233), .dout(n21524));
  jnot g03502(.din(n21238), .dout(n21525));
  jnot g03503(.din(n21243), .dout(n21526));
  jnot g03504(.din(n21248), .dout(n21527));
  jnot g03505(.din(n21253), .dout(n21528));
  jnot g03506(.din(n21258), .dout(n21529));
  jnot g03507(.din(n21263), .dout(n21530));
  jnot g03508(.din(n21268), .dout(n21531));
  jnot g03509(.din(n21273), .dout(n21532));
  jnot g03510(.din(n21278), .dout(n21533));
  jnot g03511(.din(n21283), .dout(n21534));
  jnot g03512(.din(n21288), .dout(n21535));
  jnot g03513(.din(n21293), .dout(n21536));
  jnot g03514(.din(n21298), .dout(n21537));
  jnot g03515(.din(n21303), .dout(n21538));
  jnot g03516(.din(n21308), .dout(n21539));
  jnot g03517(.din(n21313), .dout(n21540));
  jnot g03518(.din(n21318), .dout(n21541));
  jnot g03519(.din(n21324), .dout(n21542));
  jxor g03520(.dina(n21327), .dinb(n258), .dout(n21543));
  jor  g03521(.dina(n21543), .dinb(n2650), .dout(n21544));
  jand g03522(.dina(n21544), .dinb(n21542), .dout(n21545));
  jnot g03523(.din(n21331), .dout(n21546));
  jor  g03524(.dina(n21546), .dinb(n21545), .dout(n21547));
  jand g03525(.dina(n21547), .dinb(n21541), .dout(n21548));
  jnot g03526(.din(n21334), .dout(n21549));
  jor  g03527(.dina(n21549), .dinb(n21548), .dout(n21550));
  jand g03528(.dina(n21550), .dinb(n21540), .dout(n21551));
  jnot g03529(.din(n21337), .dout(n21552));
  jor  g03530(.dina(n21552), .dinb(n21551), .dout(n21553));
  jand g03531(.dina(n21553), .dinb(n21539), .dout(n21554));
  jnot g03532(.din(n21340), .dout(n21555));
  jor  g03533(.dina(n21555), .dinb(n21554), .dout(n21556));
  jand g03534(.dina(n21556), .dinb(n21538), .dout(n21557));
  jnot g03535(.din(n21343), .dout(n21558));
  jor  g03536(.dina(n21558), .dinb(n21557), .dout(n21559));
  jand g03537(.dina(n21559), .dinb(n21537), .dout(n21560));
  jnot g03538(.din(n21346), .dout(n21561));
  jor  g03539(.dina(n21561), .dinb(n21560), .dout(n21562));
  jand g03540(.dina(n21562), .dinb(n21536), .dout(n21563));
  jnot g03541(.din(n21349), .dout(n21564));
  jor  g03542(.dina(n21564), .dinb(n21563), .dout(n21565));
  jand g03543(.dina(n21565), .dinb(n21535), .dout(n21566));
  jnot g03544(.din(n21352), .dout(n21567));
  jor  g03545(.dina(n21567), .dinb(n21566), .dout(n21568));
  jand g03546(.dina(n21568), .dinb(n21534), .dout(n21569));
  jnot g03547(.din(n21355), .dout(n21570));
  jor  g03548(.dina(n21570), .dinb(n21569), .dout(n21571));
  jand g03549(.dina(n21571), .dinb(n21533), .dout(n21572));
  jnot g03550(.din(n21358), .dout(n21573));
  jor  g03551(.dina(n21573), .dinb(n21572), .dout(n21574));
  jand g03552(.dina(n21574), .dinb(n21532), .dout(n21575));
  jnot g03553(.din(n21361), .dout(n21576));
  jor  g03554(.dina(n21576), .dinb(n21575), .dout(n21577));
  jand g03555(.dina(n21577), .dinb(n21531), .dout(n21578));
  jnot g03556(.din(n21364), .dout(n21579));
  jor  g03557(.dina(n21579), .dinb(n21578), .dout(n21580));
  jand g03558(.dina(n21580), .dinb(n21530), .dout(n21581));
  jnot g03559(.din(n21367), .dout(n21582));
  jor  g03560(.dina(n21582), .dinb(n21581), .dout(n21583));
  jand g03561(.dina(n21583), .dinb(n21529), .dout(n21584));
  jnot g03562(.din(n21370), .dout(n21585));
  jor  g03563(.dina(n21585), .dinb(n21584), .dout(n21586));
  jand g03564(.dina(n21586), .dinb(n21528), .dout(n21587));
  jnot g03565(.din(n21373), .dout(n21588));
  jor  g03566(.dina(n21588), .dinb(n21587), .dout(n21589));
  jand g03567(.dina(n21589), .dinb(n21527), .dout(n21590));
  jnot g03568(.din(n21376), .dout(n21591));
  jor  g03569(.dina(n21591), .dinb(n21590), .dout(n21592));
  jand g03570(.dina(n21592), .dinb(n21526), .dout(n21593));
  jnot g03571(.din(n21379), .dout(n21594));
  jor  g03572(.dina(n21594), .dinb(n21593), .dout(n21595));
  jand g03573(.dina(n21595), .dinb(n21525), .dout(n21596));
  jnot g03574(.din(n21382), .dout(n21597));
  jor  g03575(.dina(n21597), .dinb(n21596), .dout(n21598));
  jand g03576(.dina(n21598), .dinb(n21524), .dout(n21599));
  jnot g03577(.din(n21385), .dout(n21600));
  jor  g03578(.dina(n21600), .dinb(n21599), .dout(n21601));
  jand g03579(.dina(n21601), .dinb(n21523), .dout(n21602));
  jand g03580(.dina(n21602), .dinb(n21522), .dout(n21603));
  jor  g03581(.dina(n21603), .dinb(n21219), .dout(n21604));
  jor  g03582(.dina(n21604), .dinb(n21521), .dout(n21605));
  jand g03583(.dina(n21605), .dinb(n21520), .dout(n21606));
  jor  g03584(.dina(n21606), .dinb(b1 ), .dout(n21607));
  jxor g03585(.dina(n21606), .dinb(n258), .dout(n21608));
  jor  g03586(.dina(n21608), .dinb(n2861), .dout(n21609));
  jand g03587(.dina(n21609), .dinb(n21607), .dout(n21610));
  jxor g03588(.dina(n21517), .dinb(n348), .dout(n21611));
  jor  g03589(.dina(n21611), .dinb(n21610), .dout(n21612));
  jand g03590(.dina(n21612), .dinb(n21518), .dout(n21613));
  jxor g03591(.dina(n21511), .dinb(b3 ), .dout(n21614));
  jnot g03592(.din(n21614), .dout(n21615));
  jor  g03593(.dina(n21615), .dinb(n21613), .dout(n21616));
  jand g03594(.dina(n21616), .dinb(n21512), .dout(n21617));
  jxor g03595(.dina(n21503), .dinb(n337), .dout(n21618));
  jnot g03596(.din(n21618), .dout(n21619));
  jor  g03597(.dina(n21619), .dinb(n21617), .dout(n21620));
  jand g03598(.dina(n21620), .dinb(n21505), .dout(n21621));
  jxor g03599(.dina(n21497), .dinb(n338), .dout(n21622));
  jnot g03600(.din(n21622), .dout(n21623));
  jor  g03601(.dina(n21623), .dinb(n21621), .dout(n21624));
  jand g03602(.dina(n21624), .dinb(n21499), .dout(n21625));
  jxor g03603(.dina(n21491), .dinb(n334), .dout(n21626));
  jnot g03604(.din(n21626), .dout(n21627));
  jor  g03605(.dina(n21627), .dinb(n21625), .dout(n21628));
  jand g03606(.dina(n21628), .dinb(n21493), .dout(n21629));
  jxor g03607(.dina(n21485), .dinb(n335), .dout(n21630));
  jnot g03608(.din(n21630), .dout(n21631));
  jor  g03609(.dina(n21631), .dinb(n21629), .dout(n21632));
  jand g03610(.dina(n21632), .dinb(n21487), .dout(n21633));
  jxor g03611(.dina(n21479), .dinb(n323), .dout(n21634));
  jnot g03612(.din(n21634), .dout(n21635));
  jor  g03613(.dina(n21635), .dinb(n21633), .dout(n21636));
  jand g03614(.dina(n21636), .dinb(n21481), .dout(n21637));
  jxor g03615(.dina(n21473), .dinb(n324), .dout(n21638));
  jnot g03616(.din(n21638), .dout(n21639));
  jor  g03617(.dina(n21639), .dinb(n21637), .dout(n21640));
  jand g03618(.dina(n21640), .dinb(n21475), .dout(n21641));
  jxor g03619(.dina(n21467), .dinb(n325), .dout(n21642));
  jnot g03620(.din(n21642), .dout(n21643));
  jor  g03621(.dina(n21643), .dinb(n21641), .dout(n21644));
  jand g03622(.dina(n21644), .dinb(n21469), .dout(n21645));
  jxor g03623(.dina(n21461), .dinb(n439), .dout(n21646));
  jnot g03624(.din(n21646), .dout(n21647));
  jor  g03625(.dina(n21647), .dinb(n21645), .dout(n21648));
  jand g03626(.dina(n21648), .dinb(n21463), .dout(n21649));
  jxor g03627(.dina(n21455), .dinb(n440), .dout(n21650));
  jnot g03628(.din(n21650), .dout(n21651));
  jor  g03629(.dina(n21651), .dinb(n21649), .dout(n21652));
  jand g03630(.dina(n21652), .dinb(n21457), .dout(n21653));
  jxor g03631(.dina(n21449), .dinb(n435), .dout(n21654));
  jnot g03632(.din(n21654), .dout(n21655));
  jor  g03633(.dina(n21655), .dinb(n21653), .dout(n21656));
  jand g03634(.dina(n21656), .dinb(n21451), .dout(n21657));
  jxor g03635(.dina(n21443), .dinb(n436), .dout(n21658));
  jnot g03636(.din(n21658), .dout(n21659));
  jor  g03637(.dina(n21659), .dinb(n21657), .dout(n21660));
  jand g03638(.dina(n21660), .dinb(n21445), .dout(n21661));
  jxor g03639(.dina(n21437), .dinb(n432), .dout(n21662));
  jnot g03640(.din(n21662), .dout(n21663));
  jor  g03641(.dina(n21663), .dinb(n21661), .dout(n21664));
  jand g03642(.dina(n21664), .dinb(n21439), .dout(n21665));
  jxor g03643(.dina(n21431), .dinb(n433), .dout(n21666));
  jnot g03644(.din(n21666), .dout(n21667));
  jor  g03645(.dina(n21667), .dinb(n21665), .dout(n21668));
  jand g03646(.dina(n21668), .dinb(n21433), .dout(n21669));
  jxor g03647(.dina(n21425), .dinb(n421), .dout(n21670));
  jnot g03648(.din(n21670), .dout(n21671));
  jor  g03649(.dina(n21671), .dinb(n21669), .dout(n21672));
  jand g03650(.dina(n21672), .dinb(n21427), .dout(n21673));
  jxor g03651(.dina(n21419), .dinb(n422), .dout(n21674));
  jnot g03652(.din(n21674), .dout(n21675));
  jor  g03653(.dina(n21675), .dinb(n21673), .dout(n21676));
  jand g03654(.dina(n21676), .dinb(n21421), .dout(n21677));
  jxor g03655(.dina(n21413), .dinb(n416), .dout(n21678));
  jnot g03656(.din(n21678), .dout(n21679));
  jor  g03657(.dina(n21679), .dinb(n21677), .dout(n21680));
  jand g03658(.dina(n21680), .dinb(n21415), .dout(n21681));
  jxor g03659(.dina(n21407), .dinb(n417), .dout(n21682));
  jnot g03660(.din(n21682), .dout(n21683));
  jor  g03661(.dina(n21683), .dinb(n21681), .dout(n21684));
  jand g03662(.dina(n21684), .dinb(n21409), .dout(n21685));
  jxor g03663(.dina(n21401), .dinb(n2547), .dout(n21686));
  jnot g03664(.din(n21686), .dout(n21687));
  jor  g03665(.dina(n21687), .dinb(n21685), .dout(n21688));
  jand g03666(.dina(n21688), .dinb(n21403), .dout(n21689));
  jnot g03667(.din(n21395), .dout(n21690));
  jand g03668(.dina(n21690), .dinb(b22 ), .dout(n21691));
  jor  g03669(.dina(n21691), .dinb(n21689), .dout(n21692));
  jand g03670(.dina(n21692), .dinb(n21397), .dout(n21693));
  jor  g03671(.dina(n21693), .dinb(n2718), .dout(n21694));
  jand g03672(.dina(n21694), .dinb(n21395), .dout(n21695));
  jnot g03673(.din(n21512), .dout(n21696));
  jnot g03674(.din(n21518), .dout(n21697));
  jnot g03675(.din(n2852), .dout(n21698));
  jor  g03676(.dina(n21604), .dinb(n21698), .dout(n21699));
  jand g03677(.dina(n21699), .dinb(a42 ), .dout(n21700));
  jnot g03678(.din(n21605), .dout(n21701));
  jor  g03679(.dina(n21701), .dinb(n21700), .dout(n21702));
  jand g03680(.dina(n21702), .dinb(n258), .dout(n21703));
  jxor g03681(.dina(n21606), .dinb(b1 ), .dout(n21704));
  jand g03682(.dina(n21704), .dinb(n2953), .dout(n21705));
  jor  g03683(.dina(n21705), .dinb(n21703), .dout(n21706));
  jxor g03684(.dina(n21517), .dinb(b2 ), .dout(n21707));
  jand g03685(.dina(n21707), .dinb(n21706), .dout(n21708));
  jor  g03686(.dina(n21708), .dinb(n21697), .dout(n21709));
  jand g03687(.dina(n21614), .dinb(n21709), .dout(n21710));
  jor  g03688(.dina(n21710), .dinb(n21696), .dout(n21711));
  jand g03689(.dina(n21618), .dinb(n21711), .dout(n21712));
  jor  g03690(.dina(n21712), .dinb(n21504), .dout(n21713));
  jand g03691(.dina(n21622), .dinb(n21713), .dout(n21714));
  jor  g03692(.dina(n21714), .dinb(n21498), .dout(n21715));
  jand g03693(.dina(n21626), .dinb(n21715), .dout(n21716));
  jor  g03694(.dina(n21716), .dinb(n21492), .dout(n21717));
  jand g03695(.dina(n21630), .dinb(n21717), .dout(n21718));
  jor  g03696(.dina(n21718), .dinb(n21486), .dout(n21719));
  jand g03697(.dina(n21634), .dinb(n21719), .dout(n21720));
  jor  g03698(.dina(n21720), .dinb(n21480), .dout(n21721));
  jand g03699(.dina(n21638), .dinb(n21721), .dout(n21722));
  jor  g03700(.dina(n21722), .dinb(n21474), .dout(n21723));
  jand g03701(.dina(n21642), .dinb(n21723), .dout(n21724));
  jor  g03702(.dina(n21724), .dinb(n21468), .dout(n21725));
  jand g03703(.dina(n21646), .dinb(n21725), .dout(n21726));
  jor  g03704(.dina(n21726), .dinb(n21462), .dout(n21727));
  jand g03705(.dina(n21650), .dinb(n21727), .dout(n21728));
  jor  g03706(.dina(n21728), .dinb(n21456), .dout(n21729));
  jand g03707(.dina(n21654), .dinb(n21729), .dout(n21730));
  jor  g03708(.dina(n21730), .dinb(n21450), .dout(n21731));
  jand g03709(.dina(n21658), .dinb(n21731), .dout(n21732));
  jor  g03710(.dina(n21732), .dinb(n21444), .dout(n21733));
  jand g03711(.dina(n21662), .dinb(n21733), .dout(n21734));
  jor  g03712(.dina(n21734), .dinb(n21438), .dout(n21735));
  jand g03713(.dina(n21666), .dinb(n21735), .dout(n21736));
  jor  g03714(.dina(n21736), .dinb(n21432), .dout(n21737));
  jand g03715(.dina(n21670), .dinb(n21737), .dout(n21738));
  jor  g03716(.dina(n21738), .dinb(n21426), .dout(n21739));
  jand g03717(.dina(n21674), .dinb(n21739), .dout(n21740));
  jor  g03718(.dina(n21740), .dinb(n21420), .dout(n21741));
  jand g03719(.dina(n21678), .dinb(n21741), .dout(n21742));
  jor  g03720(.dina(n21742), .dinb(n21414), .dout(n21743));
  jand g03721(.dina(n21682), .dinb(n21743), .dout(n21744));
  jor  g03722(.dina(n21744), .dinb(n21408), .dout(n21745));
  jand g03723(.dina(n21686), .dinb(n21745), .dout(n21746));
  jor  g03724(.dina(n21746), .dinb(n21402), .dout(n21747));
  jand g03725(.dina(n21396), .dinb(n2719), .dout(n21748));
  jand g03726(.dina(n21748), .dinb(n21747), .dout(n21749));
  jor  g03727(.dina(n21749), .dinb(n21695), .dout(n21750));
  jand g03728(.dina(n21750), .dinb(n2719), .dout(n21751));
  jnot g03729(.din(n21751), .dout(n21752));
  jand g03730(.dina(n21694), .dinb(n21401), .dout(n21753));
  jnot g03731(.din(n21691), .dout(n21754));
  jand g03732(.dina(n21754), .dinb(n21747), .dout(n21755));
  jor  g03733(.dina(n21755), .dinb(n21396), .dout(n21756));
  jand g03734(.dina(n21756), .dinb(n2719), .dout(n21757));
  jxor g03735(.dina(n21686), .dinb(n21745), .dout(n21758));
  jand g03736(.dina(n21758), .dinb(n21757), .dout(n21759));
  jor  g03737(.dina(n21759), .dinb(n21753), .dout(n21760));
  jand g03738(.dina(n21760), .dinb(n2714), .dout(n21761));
  jnot g03739(.din(n21761), .dout(n21762));
  jand g03740(.dina(n21694), .dinb(n21407), .dout(n21763));
  jxor g03741(.dina(n21682), .dinb(n21743), .dout(n21764));
  jand g03742(.dina(n21764), .dinb(n21757), .dout(n21765));
  jor  g03743(.dina(n21765), .dinb(n21763), .dout(n21766));
  jand g03744(.dina(n21766), .dinb(n2547), .dout(n21767));
  jnot g03745(.din(n21767), .dout(n21768));
  jand g03746(.dina(n21694), .dinb(n21413), .dout(n21769));
  jxor g03747(.dina(n21678), .dinb(n21741), .dout(n21770));
  jand g03748(.dina(n21770), .dinb(n21757), .dout(n21771));
  jor  g03749(.dina(n21771), .dinb(n21769), .dout(n21772));
  jand g03750(.dina(n21772), .dinb(n417), .dout(n21773));
  jnot g03751(.din(n21773), .dout(n21774));
  jand g03752(.dina(n21694), .dinb(n21419), .dout(n21775));
  jxor g03753(.dina(n21674), .dinb(n21739), .dout(n21776));
  jand g03754(.dina(n21776), .dinb(n21757), .dout(n21777));
  jor  g03755(.dina(n21777), .dinb(n21775), .dout(n21778));
  jand g03756(.dina(n21778), .dinb(n416), .dout(n21779));
  jnot g03757(.din(n21779), .dout(n21780));
  jand g03758(.dina(n21694), .dinb(n21425), .dout(n21781));
  jxor g03759(.dina(n21670), .dinb(n21737), .dout(n21782));
  jand g03760(.dina(n21782), .dinb(n21757), .dout(n21783));
  jor  g03761(.dina(n21783), .dinb(n21781), .dout(n21784));
  jand g03762(.dina(n21784), .dinb(n422), .dout(n21785));
  jnot g03763(.din(n21785), .dout(n21786));
  jand g03764(.dina(n21694), .dinb(n21431), .dout(n21787));
  jxor g03765(.dina(n21666), .dinb(n21735), .dout(n21788));
  jand g03766(.dina(n21788), .dinb(n21757), .dout(n21789));
  jor  g03767(.dina(n21789), .dinb(n21787), .dout(n21790));
  jand g03768(.dina(n21790), .dinb(n421), .dout(n21791));
  jnot g03769(.din(n21791), .dout(n21792));
  jand g03770(.dina(n21694), .dinb(n21437), .dout(n21793));
  jxor g03771(.dina(n21662), .dinb(n21733), .dout(n21794));
  jand g03772(.dina(n21794), .dinb(n21757), .dout(n21795));
  jor  g03773(.dina(n21795), .dinb(n21793), .dout(n21796));
  jand g03774(.dina(n21796), .dinb(n433), .dout(n21797));
  jnot g03775(.din(n21797), .dout(n21798));
  jand g03776(.dina(n21694), .dinb(n21443), .dout(n21799));
  jxor g03777(.dina(n21658), .dinb(n21731), .dout(n21800));
  jand g03778(.dina(n21800), .dinb(n21757), .dout(n21801));
  jor  g03779(.dina(n21801), .dinb(n21799), .dout(n21802));
  jand g03780(.dina(n21802), .dinb(n432), .dout(n21803));
  jnot g03781(.din(n21803), .dout(n21804));
  jand g03782(.dina(n21694), .dinb(n21449), .dout(n21805));
  jxor g03783(.dina(n21654), .dinb(n21729), .dout(n21806));
  jand g03784(.dina(n21806), .dinb(n21757), .dout(n21807));
  jor  g03785(.dina(n21807), .dinb(n21805), .dout(n21808));
  jand g03786(.dina(n21808), .dinb(n436), .dout(n21809));
  jnot g03787(.din(n21809), .dout(n21810));
  jand g03788(.dina(n21694), .dinb(n21455), .dout(n21811));
  jxor g03789(.dina(n21650), .dinb(n21727), .dout(n21812));
  jand g03790(.dina(n21812), .dinb(n21757), .dout(n21813));
  jor  g03791(.dina(n21813), .dinb(n21811), .dout(n21814));
  jand g03792(.dina(n21814), .dinb(n435), .dout(n21815));
  jnot g03793(.din(n21815), .dout(n21816));
  jand g03794(.dina(n21694), .dinb(n21461), .dout(n21817));
  jxor g03795(.dina(n21646), .dinb(n21725), .dout(n21818));
  jand g03796(.dina(n21818), .dinb(n21757), .dout(n21819));
  jor  g03797(.dina(n21819), .dinb(n21817), .dout(n21820));
  jand g03798(.dina(n21820), .dinb(n440), .dout(n21821));
  jnot g03799(.din(n21821), .dout(n21822));
  jand g03800(.dina(n21694), .dinb(n21467), .dout(n21823));
  jxor g03801(.dina(n21642), .dinb(n21723), .dout(n21824));
  jand g03802(.dina(n21824), .dinb(n21757), .dout(n21825));
  jor  g03803(.dina(n21825), .dinb(n21823), .dout(n21826));
  jand g03804(.dina(n21826), .dinb(n439), .dout(n21827));
  jnot g03805(.din(n21827), .dout(n21828));
  jand g03806(.dina(n21694), .dinb(n21473), .dout(n21829));
  jxor g03807(.dina(n21638), .dinb(n21721), .dout(n21830));
  jand g03808(.dina(n21830), .dinb(n21757), .dout(n21831));
  jor  g03809(.dina(n21831), .dinb(n21829), .dout(n21832));
  jand g03810(.dina(n21832), .dinb(n325), .dout(n21833));
  jnot g03811(.din(n21833), .dout(n21834));
  jand g03812(.dina(n21694), .dinb(n21479), .dout(n21835));
  jxor g03813(.dina(n21634), .dinb(n21719), .dout(n21836));
  jand g03814(.dina(n21836), .dinb(n21757), .dout(n21837));
  jor  g03815(.dina(n21837), .dinb(n21835), .dout(n21838));
  jand g03816(.dina(n21838), .dinb(n324), .dout(n21839));
  jnot g03817(.din(n21839), .dout(n21840));
  jand g03818(.dina(n21694), .dinb(n21485), .dout(n21841));
  jxor g03819(.dina(n21630), .dinb(n21717), .dout(n21842));
  jand g03820(.dina(n21842), .dinb(n21757), .dout(n21843));
  jor  g03821(.dina(n21843), .dinb(n21841), .dout(n21844));
  jand g03822(.dina(n21844), .dinb(n323), .dout(n21845));
  jnot g03823(.din(n21845), .dout(n21846));
  jand g03824(.dina(n21694), .dinb(n21491), .dout(n21847));
  jxor g03825(.dina(n21626), .dinb(n21715), .dout(n21848));
  jand g03826(.dina(n21848), .dinb(n21757), .dout(n21849));
  jor  g03827(.dina(n21849), .dinb(n21847), .dout(n21850));
  jand g03828(.dina(n21850), .dinb(n335), .dout(n21851));
  jnot g03829(.din(n21851), .dout(n21852));
  jand g03830(.dina(n21694), .dinb(n21497), .dout(n21853));
  jxor g03831(.dina(n21622), .dinb(n21713), .dout(n21854));
  jand g03832(.dina(n21854), .dinb(n21757), .dout(n21855));
  jor  g03833(.dina(n21855), .dinb(n21853), .dout(n21856));
  jand g03834(.dina(n21856), .dinb(n334), .dout(n21857));
  jnot g03835(.din(n21857), .dout(n21858));
  jand g03836(.dina(n21694), .dinb(n21503), .dout(n21859));
  jxor g03837(.dina(n21618), .dinb(n21711), .dout(n21860));
  jand g03838(.dina(n21860), .dinb(n21757), .dout(n21861));
  jor  g03839(.dina(n21861), .dinb(n21859), .dout(n21862));
  jand g03840(.dina(n21862), .dinb(n338), .dout(n21863));
  jnot g03841(.din(n21863), .dout(n21864));
  jor  g03842(.dina(n21757), .dinb(n21511), .dout(n21865));
  jxor g03843(.dina(n21614), .dinb(n21709), .dout(n21866));
  jand g03844(.dina(n21866), .dinb(n21757), .dout(n21867));
  jnot g03845(.din(n21867), .dout(n21868));
  jand g03846(.dina(n21868), .dinb(n21865), .dout(n21869));
  jnot g03847(.din(n21869), .dout(n21870));
  jand g03848(.dina(n21870), .dinb(n337), .dout(n21871));
  jnot g03849(.din(n21871), .dout(n21872));
  jor  g03850(.dina(n21757), .dinb(n21517), .dout(n21873));
  jxor g03851(.dina(n21707), .dinb(n21706), .dout(n21874));
  jnot g03852(.din(n21874), .dout(n21875));
  jor  g03853(.dina(n21875), .dinb(n21694), .dout(n21876));
  jand g03854(.dina(n21876), .dinb(n21873), .dout(n21877));
  jnot g03855(.din(n21877), .dout(n21878));
  jand g03856(.dina(n21878), .dinb(n344), .dout(n21879));
  jnot g03857(.din(n21879), .dout(n21880));
  jand g03858(.dina(n21694), .dinb(n21702), .dout(n21881));
  jxor g03859(.dina(n21704), .dinb(n2953), .dout(n21882));
  jand g03860(.dina(n21882), .dinb(n21757), .dout(n21883));
  jor  g03861(.dina(n21883), .dinb(n21881), .dout(n21884));
  jand g03862(.dina(n21884), .dinb(n348), .dout(n21885));
  jnot g03863(.din(n21885), .dout(n21886));
  jnot g03864(.din(n3111), .dout(n21887));
  jor  g03865(.dina(n21693), .dinb(n21887), .dout(n21888));
  jand g03866(.dina(n21888), .dinb(a41 ), .dout(n21889));
  jand g03867(.dina(n21757), .dinb(n2861), .dout(n21890));
  jor  g03868(.dina(n21890), .dinb(n21889), .dout(n21891));
  jand g03869(.dina(n21891), .dinb(n258), .dout(n21892));
  jnot g03870(.din(n21892), .dout(n21893));
  jand g03871(.dina(n21756), .dinb(n3111), .dout(n21894));
  jor  g03872(.dina(n21894), .dinb(n2860), .dout(n21895));
  jor  g03873(.dina(n21694), .dinb(n2953), .dout(n21896));
  jand g03874(.dina(n21896), .dinb(n21895), .dout(n21897));
  jxor g03875(.dina(n21897), .dinb(n258), .dout(n21898));
  jor  g03876(.dina(n21898), .dinb(n3119), .dout(n21899));
  jand g03877(.dina(n21899), .dinb(n21893), .dout(n21900));
  jxor g03878(.dina(n21884), .dinb(n348), .dout(n21901));
  jnot g03879(.din(n21901), .dout(n21902));
  jor  g03880(.dina(n21902), .dinb(n21900), .dout(n21903));
  jand g03881(.dina(n21903), .dinb(n21886), .dout(n21904));
  jxor g03882(.dina(n21877), .dinb(b3 ), .dout(n21905));
  jnot g03883(.din(n21905), .dout(n21906));
  jor  g03884(.dina(n21906), .dinb(n21904), .dout(n21907));
  jand g03885(.dina(n21907), .dinb(n21880), .dout(n21908));
  jxor g03886(.dina(n21869), .dinb(b4 ), .dout(n21909));
  jnot g03887(.din(n21909), .dout(n21910));
  jor  g03888(.dina(n21910), .dinb(n21908), .dout(n21911));
  jand g03889(.dina(n21911), .dinb(n21872), .dout(n21912));
  jxor g03890(.dina(n21862), .dinb(n338), .dout(n21913));
  jnot g03891(.din(n21913), .dout(n21914));
  jor  g03892(.dina(n21914), .dinb(n21912), .dout(n21915));
  jand g03893(.dina(n21915), .dinb(n21864), .dout(n21916));
  jxor g03894(.dina(n21856), .dinb(n334), .dout(n21917));
  jnot g03895(.din(n21917), .dout(n21918));
  jor  g03896(.dina(n21918), .dinb(n21916), .dout(n21919));
  jand g03897(.dina(n21919), .dinb(n21858), .dout(n21920));
  jxor g03898(.dina(n21850), .dinb(n335), .dout(n21921));
  jnot g03899(.din(n21921), .dout(n21922));
  jor  g03900(.dina(n21922), .dinb(n21920), .dout(n21923));
  jand g03901(.dina(n21923), .dinb(n21852), .dout(n21924));
  jxor g03902(.dina(n21844), .dinb(n323), .dout(n21925));
  jnot g03903(.din(n21925), .dout(n21926));
  jor  g03904(.dina(n21926), .dinb(n21924), .dout(n21927));
  jand g03905(.dina(n21927), .dinb(n21846), .dout(n21928));
  jxor g03906(.dina(n21838), .dinb(n324), .dout(n21929));
  jnot g03907(.din(n21929), .dout(n21930));
  jor  g03908(.dina(n21930), .dinb(n21928), .dout(n21931));
  jand g03909(.dina(n21931), .dinb(n21840), .dout(n21932));
  jxor g03910(.dina(n21832), .dinb(n325), .dout(n21933));
  jnot g03911(.din(n21933), .dout(n21934));
  jor  g03912(.dina(n21934), .dinb(n21932), .dout(n21935));
  jand g03913(.dina(n21935), .dinb(n21834), .dout(n21936));
  jxor g03914(.dina(n21826), .dinb(n439), .dout(n21937));
  jnot g03915(.din(n21937), .dout(n21938));
  jor  g03916(.dina(n21938), .dinb(n21936), .dout(n21939));
  jand g03917(.dina(n21939), .dinb(n21828), .dout(n21940));
  jxor g03918(.dina(n21820), .dinb(n440), .dout(n21941));
  jnot g03919(.din(n21941), .dout(n21942));
  jor  g03920(.dina(n21942), .dinb(n21940), .dout(n21943));
  jand g03921(.dina(n21943), .dinb(n21822), .dout(n21944));
  jxor g03922(.dina(n21814), .dinb(n435), .dout(n21945));
  jnot g03923(.din(n21945), .dout(n21946));
  jor  g03924(.dina(n21946), .dinb(n21944), .dout(n21947));
  jand g03925(.dina(n21947), .dinb(n21816), .dout(n21948));
  jxor g03926(.dina(n21808), .dinb(n436), .dout(n21949));
  jnot g03927(.din(n21949), .dout(n21950));
  jor  g03928(.dina(n21950), .dinb(n21948), .dout(n21951));
  jand g03929(.dina(n21951), .dinb(n21810), .dout(n21952));
  jxor g03930(.dina(n21802), .dinb(n432), .dout(n21953));
  jnot g03931(.din(n21953), .dout(n21954));
  jor  g03932(.dina(n21954), .dinb(n21952), .dout(n21955));
  jand g03933(.dina(n21955), .dinb(n21804), .dout(n21956));
  jxor g03934(.dina(n21796), .dinb(n433), .dout(n21957));
  jnot g03935(.din(n21957), .dout(n21958));
  jor  g03936(.dina(n21958), .dinb(n21956), .dout(n21959));
  jand g03937(.dina(n21959), .dinb(n21798), .dout(n21960));
  jxor g03938(.dina(n21790), .dinb(n421), .dout(n21961));
  jnot g03939(.din(n21961), .dout(n21962));
  jor  g03940(.dina(n21962), .dinb(n21960), .dout(n21963));
  jand g03941(.dina(n21963), .dinb(n21792), .dout(n21964));
  jxor g03942(.dina(n21784), .dinb(n422), .dout(n21965));
  jnot g03943(.din(n21965), .dout(n21966));
  jor  g03944(.dina(n21966), .dinb(n21964), .dout(n21967));
  jand g03945(.dina(n21967), .dinb(n21786), .dout(n21968));
  jxor g03946(.dina(n21778), .dinb(n416), .dout(n21969));
  jnot g03947(.din(n21969), .dout(n21970));
  jor  g03948(.dina(n21970), .dinb(n21968), .dout(n21971));
  jand g03949(.dina(n21971), .dinb(n21780), .dout(n21972));
  jxor g03950(.dina(n21772), .dinb(n417), .dout(n21973));
  jnot g03951(.din(n21973), .dout(n21974));
  jor  g03952(.dina(n21974), .dinb(n21972), .dout(n21975));
  jand g03953(.dina(n21975), .dinb(n21774), .dout(n21976));
  jxor g03954(.dina(n21766), .dinb(n2547), .dout(n21977));
  jnot g03955(.din(n21977), .dout(n21978));
  jor  g03956(.dina(n21978), .dinb(n21976), .dout(n21979));
  jand g03957(.dina(n21979), .dinb(n21768), .dout(n21980));
  jxor g03958(.dina(n21760), .dinb(n2714), .dout(n21981));
  jnot g03959(.din(n21981), .dout(n21982));
  jor  g03960(.dina(n21982), .dinb(n21980), .dout(n21983));
  jand g03961(.dina(n21983), .dinb(n21762), .dout(n21984));
  jxor g03962(.dina(n21750), .dinb(b23 ), .dout(n21985));
  jor  g03963(.dina(n21985), .dinb(n21984), .dout(n21986));
  jor  g03964(.dina(n21986), .dinb(n455), .dout(n21987));
  jand g03965(.dina(n21987), .dinb(n21752), .dout(n21988));
  jand g03966(.dina(n21988), .dinb(n21750), .dout(n21989));
  jnot g03967(.din(n21989), .dout(n21990));
  jxor g03968(.dina(n21897), .dinb(b1 ), .dout(n21991));
  jand g03969(.dina(n21991), .dinb(n3120), .dout(n21992));
  jor  g03970(.dina(n21992), .dinb(n21892), .dout(n21993));
  jand g03971(.dina(n21901), .dinb(n21993), .dout(n21994));
  jor  g03972(.dina(n21994), .dinb(n21885), .dout(n21995));
  jand g03973(.dina(n21905), .dinb(n21995), .dout(n21996));
  jor  g03974(.dina(n21996), .dinb(n21879), .dout(n21997));
  jand g03975(.dina(n21909), .dinb(n21997), .dout(n21998));
  jor  g03976(.dina(n21998), .dinb(n21871), .dout(n21999));
  jand g03977(.dina(n21913), .dinb(n21999), .dout(n22000));
  jor  g03978(.dina(n22000), .dinb(n21863), .dout(n22001));
  jand g03979(.dina(n21917), .dinb(n22001), .dout(n22002));
  jor  g03980(.dina(n22002), .dinb(n21857), .dout(n22003));
  jand g03981(.dina(n21921), .dinb(n22003), .dout(n22004));
  jor  g03982(.dina(n22004), .dinb(n21851), .dout(n22005));
  jand g03983(.dina(n21925), .dinb(n22005), .dout(n22006));
  jor  g03984(.dina(n22006), .dinb(n21845), .dout(n22007));
  jand g03985(.dina(n21929), .dinb(n22007), .dout(n22008));
  jor  g03986(.dina(n22008), .dinb(n21839), .dout(n22009));
  jand g03987(.dina(n21933), .dinb(n22009), .dout(n22010));
  jor  g03988(.dina(n22010), .dinb(n21833), .dout(n22011));
  jand g03989(.dina(n21937), .dinb(n22011), .dout(n22012));
  jor  g03990(.dina(n22012), .dinb(n21827), .dout(n22013));
  jand g03991(.dina(n21941), .dinb(n22013), .dout(n22014));
  jor  g03992(.dina(n22014), .dinb(n21821), .dout(n22015));
  jand g03993(.dina(n21945), .dinb(n22015), .dout(n22016));
  jor  g03994(.dina(n22016), .dinb(n21815), .dout(n22017));
  jand g03995(.dina(n21949), .dinb(n22017), .dout(n22018));
  jor  g03996(.dina(n22018), .dinb(n21809), .dout(n22019));
  jand g03997(.dina(n21953), .dinb(n22019), .dout(n22020));
  jor  g03998(.dina(n22020), .dinb(n21803), .dout(n22021));
  jand g03999(.dina(n21957), .dinb(n22021), .dout(n22022));
  jor  g04000(.dina(n22022), .dinb(n21797), .dout(n22023));
  jand g04001(.dina(n21961), .dinb(n22023), .dout(n22024));
  jor  g04002(.dina(n22024), .dinb(n21791), .dout(n22025));
  jand g04003(.dina(n21965), .dinb(n22025), .dout(n22026));
  jor  g04004(.dina(n22026), .dinb(n21785), .dout(n22027));
  jand g04005(.dina(n21969), .dinb(n22027), .dout(n22028));
  jor  g04006(.dina(n22028), .dinb(n21779), .dout(n22029));
  jand g04007(.dina(n21973), .dinb(n22029), .dout(n22030));
  jor  g04008(.dina(n22030), .dinb(n21773), .dout(n22031));
  jand g04009(.dina(n21977), .dinb(n22031), .dout(n22032));
  jor  g04010(.dina(n22032), .dinb(n21767), .dout(n22033));
  jand g04011(.dina(n21981), .dinb(n22033), .dout(n22034));
  jor  g04012(.dina(n22034), .dinb(n21761), .dout(n22035));
  jnot g04013(.din(n21985), .dout(n22036));
  jand g04014(.dina(n22036), .dinb(n22035), .dout(n22037));
  jand g04015(.dina(n21984), .dinb(n405), .dout(n22038));
  jor  g04016(.dina(n22038), .dinb(n21752), .dout(n22039));
  jor  g04017(.dina(n22039), .dinb(n22037), .dout(n22040));
  jand g04018(.dina(n22040), .dinb(n21990), .dout(n22041));
  jnot g04019(.din(n22041), .dout(n22042));
  jand g04020(.dina(n22042), .dinb(n406), .dout(n22043));
  jand g04021(.dina(n21988), .dinb(n21760), .dout(n22044));
  jand g04022(.dina(n22037), .dinb(n592), .dout(n22045));
  jor  g04023(.dina(n22045), .dinb(n21751), .dout(n22046));
  jxor g04024(.dina(n21981), .dinb(n22033), .dout(n22047));
  jand g04025(.dina(n22047), .dinb(n22046), .dout(n22048));
  jor  g04026(.dina(n22048), .dinb(n22044), .dout(n22049));
  jand g04027(.dina(n22049), .dinb(n405), .dout(n22050));
  jand g04028(.dina(n21988), .dinb(n21766), .dout(n22051));
  jxor g04029(.dina(n21977), .dinb(n22031), .dout(n22052));
  jand g04030(.dina(n22052), .dinb(n22046), .dout(n22053));
  jor  g04031(.dina(n22053), .dinb(n22051), .dout(n22054));
  jand g04032(.dina(n22054), .dinb(n2714), .dout(n22055));
  jand g04033(.dina(n21988), .dinb(n21772), .dout(n22056));
  jxor g04034(.dina(n21973), .dinb(n22029), .dout(n22057));
  jand g04035(.dina(n22057), .dinb(n22046), .dout(n22058));
  jor  g04036(.dina(n22058), .dinb(n22056), .dout(n22059));
  jand g04037(.dina(n22059), .dinb(n2547), .dout(n22060));
  jand g04038(.dina(n21988), .dinb(n21778), .dout(n22061));
  jxor g04039(.dina(n21969), .dinb(n22027), .dout(n22062));
  jand g04040(.dina(n22062), .dinb(n22046), .dout(n22063));
  jor  g04041(.dina(n22063), .dinb(n22061), .dout(n22064));
  jand g04042(.dina(n22064), .dinb(n417), .dout(n22065));
  jand g04043(.dina(n21988), .dinb(n21784), .dout(n22066));
  jxor g04044(.dina(n21965), .dinb(n22025), .dout(n22067));
  jand g04045(.dina(n22067), .dinb(n22046), .dout(n22068));
  jor  g04046(.dina(n22068), .dinb(n22066), .dout(n22069));
  jand g04047(.dina(n22069), .dinb(n416), .dout(n22070));
  jand g04048(.dina(n21988), .dinb(n21790), .dout(n22071));
  jxor g04049(.dina(n21961), .dinb(n22023), .dout(n22072));
  jand g04050(.dina(n22072), .dinb(n22046), .dout(n22073));
  jor  g04051(.dina(n22073), .dinb(n22071), .dout(n22074));
  jand g04052(.dina(n22074), .dinb(n422), .dout(n22075));
  jand g04053(.dina(n21988), .dinb(n21796), .dout(n22076));
  jxor g04054(.dina(n21957), .dinb(n22021), .dout(n22077));
  jand g04055(.dina(n22077), .dinb(n22046), .dout(n22078));
  jor  g04056(.dina(n22078), .dinb(n22076), .dout(n22079));
  jand g04057(.dina(n22079), .dinb(n421), .dout(n22080));
  jand g04058(.dina(n21988), .dinb(n21802), .dout(n22081));
  jxor g04059(.dina(n21953), .dinb(n22019), .dout(n22082));
  jand g04060(.dina(n22082), .dinb(n22046), .dout(n22083));
  jor  g04061(.dina(n22083), .dinb(n22081), .dout(n22084));
  jand g04062(.dina(n22084), .dinb(n433), .dout(n22085));
  jand g04063(.dina(n21988), .dinb(n21808), .dout(n22086));
  jxor g04064(.dina(n21949), .dinb(n22017), .dout(n22087));
  jand g04065(.dina(n22087), .dinb(n22046), .dout(n22088));
  jor  g04066(.dina(n22088), .dinb(n22086), .dout(n22089));
  jand g04067(.dina(n22089), .dinb(n432), .dout(n22090));
  jand g04068(.dina(n21988), .dinb(n21814), .dout(n22091));
  jxor g04069(.dina(n21945), .dinb(n22015), .dout(n22092));
  jand g04070(.dina(n22092), .dinb(n22046), .dout(n22093));
  jor  g04071(.dina(n22093), .dinb(n22091), .dout(n22094));
  jand g04072(.dina(n22094), .dinb(n436), .dout(n22095));
  jand g04073(.dina(n21988), .dinb(n21820), .dout(n22096));
  jxor g04074(.dina(n21941), .dinb(n22013), .dout(n22097));
  jand g04075(.dina(n22097), .dinb(n22046), .dout(n22098));
  jor  g04076(.dina(n22098), .dinb(n22096), .dout(n22099));
  jand g04077(.dina(n22099), .dinb(n435), .dout(n22100));
  jand g04078(.dina(n21988), .dinb(n21826), .dout(n22101));
  jxor g04079(.dina(n21937), .dinb(n22011), .dout(n22102));
  jand g04080(.dina(n22102), .dinb(n22046), .dout(n22103));
  jor  g04081(.dina(n22103), .dinb(n22101), .dout(n22104));
  jand g04082(.dina(n22104), .dinb(n440), .dout(n22105));
  jand g04083(.dina(n21988), .dinb(n21832), .dout(n22106));
  jxor g04084(.dina(n21933), .dinb(n22009), .dout(n22107));
  jand g04085(.dina(n22107), .dinb(n22046), .dout(n22108));
  jor  g04086(.dina(n22108), .dinb(n22106), .dout(n22109));
  jand g04087(.dina(n22109), .dinb(n439), .dout(n22110));
  jand g04088(.dina(n21988), .dinb(n21838), .dout(n22111));
  jxor g04089(.dina(n21929), .dinb(n22007), .dout(n22112));
  jand g04090(.dina(n22112), .dinb(n22046), .dout(n22113));
  jor  g04091(.dina(n22113), .dinb(n22111), .dout(n22114));
  jand g04092(.dina(n22114), .dinb(n325), .dout(n22115));
  jand g04093(.dina(n21988), .dinb(n21844), .dout(n22116));
  jxor g04094(.dina(n21925), .dinb(n22005), .dout(n22117));
  jand g04095(.dina(n22117), .dinb(n22046), .dout(n22118));
  jor  g04096(.dina(n22118), .dinb(n22116), .dout(n22119));
  jand g04097(.dina(n22119), .dinb(n324), .dout(n22120));
  jand g04098(.dina(n21988), .dinb(n21850), .dout(n22121));
  jxor g04099(.dina(n21921), .dinb(n22003), .dout(n22122));
  jand g04100(.dina(n22122), .dinb(n22046), .dout(n22123));
  jor  g04101(.dina(n22123), .dinb(n22121), .dout(n22124));
  jand g04102(.dina(n22124), .dinb(n323), .dout(n22125));
  jand g04103(.dina(n21988), .dinb(n21856), .dout(n22126));
  jxor g04104(.dina(n21917), .dinb(n22001), .dout(n22127));
  jand g04105(.dina(n22127), .dinb(n22046), .dout(n22128));
  jor  g04106(.dina(n22128), .dinb(n22126), .dout(n22129));
  jand g04107(.dina(n22129), .dinb(n335), .dout(n22130));
  jand g04108(.dina(n21988), .dinb(n21862), .dout(n22131));
  jxor g04109(.dina(n21913), .dinb(n21999), .dout(n22132));
  jand g04110(.dina(n22132), .dinb(n22046), .dout(n22133));
  jor  g04111(.dina(n22133), .dinb(n22131), .dout(n22134));
  jand g04112(.dina(n22134), .dinb(n334), .dout(n22135));
  jand g04113(.dina(n21988), .dinb(n21870), .dout(n22136));
  jxor g04114(.dina(n21909), .dinb(n21997), .dout(n22137));
  jand g04115(.dina(n22137), .dinb(n22046), .dout(n22138));
  jor  g04116(.dina(n22138), .dinb(n22136), .dout(n22139));
  jand g04117(.dina(n22139), .dinb(n338), .dout(n22140));
  jand g04118(.dina(n21988), .dinb(n21878), .dout(n22141));
  jxor g04119(.dina(n21905), .dinb(n21995), .dout(n22142));
  jand g04120(.dina(n22142), .dinb(n22046), .dout(n22143));
  jor  g04121(.dina(n22143), .dinb(n22141), .dout(n22144));
  jand g04122(.dina(n22144), .dinb(n337), .dout(n22145));
  jand g04123(.dina(n21988), .dinb(n21884), .dout(n22146));
  jxor g04124(.dina(n21901), .dinb(n21993), .dout(n22147));
  jand g04125(.dina(n22147), .dinb(n22046), .dout(n22148));
  jor  g04126(.dina(n22148), .dinb(n22146), .dout(n22149));
  jand g04127(.dina(n22149), .dinb(n344), .dout(n22150));
  jand g04128(.dina(n21988), .dinb(n21891), .dout(n22151));
  jxor g04129(.dina(n21991), .dinb(n3120), .dout(n22152));
  jand g04130(.dina(n22152), .dinb(n22046), .dout(n22153));
  jor  g04131(.dina(n22153), .dinb(n22151), .dout(n22154));
  jand g04132(.dina(n22154), .dinb(n348), .dout(n22155));
  jor  g04133(.dina(n21988), .dinb(n18364), .dout(n22156));
  jand g04134(.dina(n22156), .dinb(a40 ), .dout(n22157));
  jor  g04135(.dina(n21988), .dinb(n3120), .dout(n22158));
  jnot g04136(.din(n22158), .dout(n22159));
  jor  g04137(.dina(n22159), .dinb(n22157), .dout(n22160));
  jand g04138(.dina(n22160), .dinb(n258), .dout(n22161));
  jand g04139(.dina(n22046), .dinb(b0 ), .dout(n22162));
  jor  g04140(.dina(n22162), .dinb(n3118), .dout(n22163));
  jand g04141(.dina(n22158), .dinb(n22163), .dout(n22164));
  jxor g04142(.dina(n22164), .dinb(b1 ), .dout(n22165));
  jand g04143(.dina(n22165), .dinb(n3322), .dout(n22166));
  jor  g04144(.dina(n22166), .dinb(n22161), .dout(n22167));
  jxor g04145(.dina(n22154), .dinb(n348), .dout(n22168));
  jand g04146(.dina(n22168), .dinb(n22167), .dout(n22169));
  jor  g04147(.dina(n22169), .dinb(n22155), .dout(n22170));
  jxor g04148(.dina(n22149), .dinb(n344), .dout(n22171));
  jand g04149(.dina(n22171), .dinb(n22170), .dout(n22172));
  jor  g04150(.dina(n22172), .dinb(n22150), .dout(n22173));
  jxor g04151(.dina(n22144), .dinb(n337), .dout(n22174));
  jand g04152(.dina(n22174), .dinb(n22173), .dout(n22175));
  jor  g04153(.dina(n22175), .dinb(n22145), .dout(n22176));
  jxor g04154(.dina(n22139), .dinb(n338), .dout(n22177));
  jand g04155(.dina(n22177), .dinb(n22176), .dout(n22178));
  jor  g04156(.dina(n22178), .dinb(n22140), .dout(n22179));
  jxor g04157(.dina(n22134), .dinb(n334), .dout(n22180));
  jand g04158(.dina(n22180), .dinb(n22179), .dout(n22181));
  jor  g04159(.dina(n22181), .dinb(n22135), .dout(n22182));
  jxor g04160(.dina(n22129), .dinb(n335), .dout(n22183));
  jand g04161(.dina(n22183), .dinb(n22182), .dout(n22184));
  jor  g04162(.dina(n22184), .dinb(n22130), .dout(n22185));
  jxor g04163(.dina(n22124), .dinb(n323), .dout(n22186));
  jand g04164(.dina(n22186), .dinb(n22185), .dout(n22187));
  jor  g04165(.dina(n22187), .dinb(n22125), .dout(n22188));
  jxor g04166(.dina(n22119), .dinb(n324), .dout(n22189));
  jand g04167(.dina(n22189), .dinb(n22188), .dout(n22190));
  jor  g04168(.dina(n22190), .dinb(n22120), .dout(n22191));
  jxor g04169(.dina(n22114), .dinb(n325), .dout(n22192));
  jand g04170(.dina(n22192), .dinb(n22191), .dout(n22193));
  jor  g04171(.dina(n22193), .dinb(n22115), .dout(n22194));
  jxor g04172(.dina(n22109), .dinb(n439), .dout(n22195));
  jand g04173(.dina(n22195), .dinb(n22194), .dout(n22196));
  jor  g04174(.dina(n22196), .dinb(n22110), .dout(n22197));
  jxor g04175(.dina(n22104), .dinb(n440), .dout(n22198));
  jand g04176(.dina(n22198), .dinb(n22197), .dout(n22199));
  jor  g04177(.dina(n22199), .dinb(n22105), .dout(n22200));
  jxor g04178(.dina(n22099), .dinb(n435), .dout(n22201));
  jand g04179(.dina(n22201), .dinb(n22200), .dout(n22202));
  jor  g04180(.dina(n22202), .dinb(n22100), .dout(n22203));
  jxor g04181(.dina(n22094), .dinb(n436), .dout(n22204));
  jand g04182(.dina(n22204), .dinb(n22203), .dout(n22205));
  jor  g04183(.dina(n22205), .dinb(n22095), .dout(n22206));
  jxor g04184(.dina(n22089), .dinb(n432), .dout(n22207));
  jand g04185(.dina(n22207), .dinb(n22206), .dout(n22208));
  jor  g04186(.dina(n22208), .dinb(n22090), .dout(n22209));
  jxor g04187(.dina(n22084), .dinb(n433), .dout(n22210));
  jand g04188(.dina(n22210), .dinb(n22209), .dout(n22211));
  jor  g04189(.dina(n22211), .dinb(n22085), .dout(n22212));
  jxor g04190(.dina(n22079), .dinb(n421), .dout(n22213));
  jand g04191(.dina(n22213), .dinb(n22212), .dout(n22214));
  jor  g04192(.dina(n22214), .dinb(n22080), .dout(n22215));
  jxor g04193(.dina(n22074), .dinb(n422), .dout(n22216));
  jand g04194(.dina(n22216), .dinb(n22215), .dout(n22217));
  jor  g04195(.dina(n22217), .dinb(n22075), .dout(n22218));
  jxor g04196(.dina(n22069), .dinb(n416), .dout(n22219));
  jand g04197(.dina(n22219), .dinb(n22218), .dout(n22220));
  jor  g04198(.dina(n22220), .dinb(n22070), .dout(n22221));
  jxor g04199(.dina(n22064), .dinb(n417), .dout(n22222));
  jand g04200(.dina(n22222), .dinb(n22221), .dout(n22223));
  jor  g04201(.dina(n22223), .dinb(n22065), .dout(n22224));
  jxor g04202(.dina(n22059), .dinb(n2547), .dout(n22225));
  jand g04203(.dina(n22225), .dinb(n22224), .dout(n22226));
  jor  g04204(.dina(n22226), .dinb(n22060), .dout(n22227));
  jxor g04205(.dina(n22054), .dinb(n2714), .dout(n22228));
  jand g04206(.dina(n22228), .dinb(n22227), .dout(n22229));
  jor  g04207(.dina(n22229), .dinb(n22055), .dout(n22230));
  jxor g04208(.dina(n22049), .dinb(n405), .dout(n22231));
  jand g04209(.dina(n22231), .dinb(n22230), .dout(n22232));
  jor  g04210(.dina(n22232), .dinb(n22050), .dout(n22233));
  jand g04211(.dina(n22041), .dinb(b24 ), .dout(n22234));
  jnot g04212(.din(n22234), .dout(n22235));
  jand g04213(.dina(n22235), .dinb(n22233), .dout(n22236));
  jor  g04214(.dina(n22236), .dinb(n22043), .dout(n22237));
  jand g04215(.dina(n22237), .dinb(n2457), .dout(n22238));
  jnot g04216(.din(n22238), .dout(n22239));
  jand g04217(.dina(n22239), .dinb(n22042), .dout(n22240));
  jand g04218(.dina(n22043), .dinb(n2457), .dout(n22241));
  jand g04219(.dina(n22241), .dinb(n22233), .dout(n22242));
  jor  g04220(.dina(n22242), .dinb(n22240), .dout(n22243));
  jand g04221(.dina(n22243), .dinb(n412), .dout(n22244));
  jnot g04222(.din(n22244), .dout(n22245));
  jand g04223(.dina(n22239), .dinb(n22049), .dout(n22246));
  jxor g04224(.dina(n22231), .dinb(n22230), .dout(n22247));
  jand g04225(.dina(n22247), .dinb(n22238), .dout(n22248));
  jor  g04226(.dina(n22248), .dinb(n22246), .dout(n22249));
  jand g04227(.dina(n22249), .dinb(n406), .dout(n22250));
  jnot g04228(.din(n22250), .dout(n22251));
  jand g04229(.dina(n22239), .dinb(n22054), .dout(n22252));
  jxor g04230(.dina(n22228), .dinb(n22227), .dout(n22253));
  jand g04231(.dina(n22253), .dinb(n22238), .dout(n22254));
  jor  g04232(.dina(n22254), .dinb(n22252), .dout(n22255));
  jand g04233(.dina(n22255), .dinb(n405), .dout(n22256));
  jnot g04234(.din(n22256), .dout(n22257));
  jand g04235(.dina(n22239), .dinb(n22059), .dout(n22258));
  jxor g04236(.dina(n22225), .dinb(n22224), .dout(n22259));
  jand g04237(.dina(n22259), .dinb(n22238), .dout(n22260));
  jor  g04238(.dina(n22260), .dinb(n22258), .dout(n22261));
  jand g04239(.dina(n22261), .dinb(n2714), .dout(n22262));
  jnot g04240(.din(n22262), .dout(n22263));
  jand g04241(.dina(n22239), .dinb(n22064), .dout(n22264));
  jxor g04242(.dina(n22222), .dinb(n22221), .dout(n22265));
  jand g04243(.dina(n22265), .dinb(n22238), .dout(n22266));
  jor  g04244(.dina(n22266), .dinb(n22264), .dout(n22267));
  jand g04245(.dina(n22267), .dinb(n2547), .dout(n22268));
  jnot g04246(.din(n22268), .dout(n22269));
  jand g04247(.dina(n22239), .dinb(n22069), .dout(n22270));
  jxor g04248(.dina(n22219), .dinb(n22218), .dout(n22271));
  jand g04249(.dina(n22271), .dinb(n22238), .dout(n22272));
  jor  g04250(.dina(n22272), .dinb(n22270), .dout(n22273));
  jand g04251(.dina(n22273), .dinb(n417), .dout(n22274));
  jnot g04252(.din(n22274), .dout(n22275));
  jand g04253(.dina(n22239), .dinb(n22074), .dout(n22276));
  jxor g04254(.dina(n22216), .dinb(n22215), .dout(n22277));
  jand g04255(.dina(n22277), .dinb(n22238), .dout(n22278));
  jor  g04256(.dina(n22278), .dinb(n22276), .dout(n22279));
  jand g04257(.dina(n22279), .dinb(n416), .dout(n22280));
  jnot g04258(.din(n22280), .dout(n22281));
  jand g04259(.dina(n22239), .dinb(n22079), .dout(n22282));
  jxor g04260(.dina(n22213), .dinb(n22212), .dout(n22283));
  jand g04261(.dina(n22283), .dinb(n22238), .dout(n22284));
  jor  g04262(.dina(n22284), .dinb(n22282), .dout(n22285));
  jand g04263(.dina(n22285), .dinb(n422), .dout(n22286));
  jnot g04264(.din(n22286), .dout(n22287));
  jand g04265(.dina(n22239), .dinb(n22084), .dout(n22288));
  jxor g04266(.dina(n22210), .dinb(n22209), .dout(n22289));
  jand g04267(.dina(n22289), .dinb(n22238), .dout(n22290));
  jor  g04268(.dina(n22290), .dinb(n22288), .dout(n22291));
  jand g04269(.dina(n22291), .dinb(n421), .dout(n22292));
  jnot g04270(.din(n22292), .dout(n22293));
  jand g04271(.dina(n22239), .dinb(n22089), .dout(n22294));
  jxor g04272(.dina(n22207), .dinb(n22206), .dout(n22295));
  jand g04273(.dina(n22295), .dinb(n22238), .dout(n22296));
  jor  g04274(.dina(n22296), .dinb(n22294), .dout(n22297));
  jand g04275(.dina(n22297), .dinb(n433), .dout(n22298));
  jnot g04276(.din(n22298), .dout(n22299));
  jand g04277(.dina(n22239), .dinb(n22094), .dout(n22300));
  jxor g04278(.dina(n22204), .dinb(n22203), .dout(n22301));
  jand g04279(.dina(n22301), .dinb(n22238), .dout(n22302));
  jor  g04280(.dina(n22302), .dinb(n22300), .dout(n22303));
  jand g04281(.dina(n22303), .dinb(n432), .dout(n22304));
  jnot g04282(.din(n22304), .dout(n22305));
  jand g04283(.dina(n22239), .dinb(n22099), .dout(n22306));
  jxor g04284(.dina(n22201), .dinb(n22200), .dout(n22307));
  jand g04285(.dina(n22307), .dinb(n22238), .dout(n22308));
  jor  g04286(.dina(n22308), .dinb(n22306), .dout(n22309));
  jand g04287(.dina(n22309), .dinb(n436), .dout(n22310));
  jnot g04288(.din(n22310), .dout(n22311));
  jand g04289(.dina(n22239), .dinb(n22104), .dout(n22312));
  jxor g04290(.dina(n22198), .dinb(n22197), .dout(n22313));
  jand g04291(.dina(n22313), .dinb(n22238), .dout(n22314));
  jor  g04292(.dina(n22314), .dinb(n22312), .dout(n22315));
  jand g04293(.dina(n22315), .dinb(n435), .dout(n22316));
  jnot g04294(.din(n22316), .dout(n22317));
  jand g04295(.dina(n22239), .dinb(n22109), .dout(n22318));
  jxor g04296(.dina(n22195), .dinb(n22194), .dout(n22319));
  jand g04297(.dina(n22319), .dinb(n22238), .dout(n22320));
  jor  g04298(.dina(n22320), .dinb(n22318), .dout(n22321));
  jand g04299(.dina(n22321), .dinb(n440), .dout(n22322));
  jnot g04300(.din(n22322), .dout(n22323));
  jand g04301(.dina(n22239), .dinb(n22114), .dout(n22324));
  jxor g04302(.dina(n22192), .dinb(n22191), .dout(n22325));
  jand g04303(.dina(n22325), .dinb(n22238), .dout(n22326));
  jor  g04304(.dina(n22326), .dinb(n22324), .dout(n22327));
  jand g04305(.dina(n22327), .dinb(n439), .dout(n22328));
  jnot g04306(.din(n22328), .dout(n22329));
  jand g04307(.dina(n22239), .dinb(n22119), .dout(n22330));
  jxor g04308(.dina(n22189), .dinb(n22188), .dout(n22331));
  jand g04309(.dina(n22331), .dinb(n22238), .dout(n22332));
  jor  g04310(.dina(n22332), .dinb(n22330), .dout(n22333));
  jand g04311(.dina(n22333), .dinb(n325), .dout(n22334));
  jnot g04312(.din(n22334), .dout(n22335));
  jand g04313(.dina(n22239), .dinb(n22124), .dout(n22336));
  jxor g04314(.dina(n22186), .dinb(n22185), .dout(n22337));
  jand g04315(.dina(n22337), .dinb(n22238), .dout(n22338));
  jor  g04316(.dina(n22338), .dinb(n22336), .dout(n22339));
  jand g04317(.dina(n22339), .dinb(n324), .dout(n22340));
  jnot g04318(.din(n22340), .dout(n22341));
  jand g04319(.dina(n22239), .dinb(n22129), .dout(n22342));
  jxor g04320(.dina(n22183), .dinb(n22182), .dout(n22343));
  jand g04321(.dina(n22343), .dinb(n22238), .dout(n22344));
  jor  g04322(.dina(n22344), .dinb(n22342), .dout(n22345));
  jand g04323(.dina(n22345), .dinb(n323), .dout(n22346));
  jnot g04324(.din(n22346), .dout(n22347));
  jand g04325(.dina(n22239), .dinb(n22134), .dout(n22348));
  jxor g04326(.dina(n22180), .dinb(n22179), .dout(n22349));
  jand g04327(.dina(n22349), .dinb(n22238), .dout(n22350));
  jor  g04328(.dina(n22350), .dinb(n22348), .dout(n22351));
  jand g04329(.dina(n22351), .dinb(n335), .dout(n22352));
  jnot g04330(.din(n22352), .dout(n22353));
  jand g04331(.dina(n22239), .dinb(n22139), .dout(n22354));
  jxor g04332(.dina(n22177), .dinb(n22176), .dout(n22355));
  jand g04333(.dina(n22355), .dinb(n22238), .dout(n22356));
  jor  g04334(.dina(n22356), .dinb(n22354), .dout(n22357));
  jand g04335(.dina(n22357), .dinb(n334), .dout(n22358));
  jnot g04336(.din(n22358), .dout(n22359));
  jand g04337(.dina(n22239), .dinb(n22144), .dout(n22360));
  jxor g04338(.dina(n22174), .dinb(n22173), .dout(n22361));
  jand g04339(.dina(n22361), .dinb(n22238), .dout(n22362));
  jor  g04340(.dina(n22362), .dinb(n22360), .dout(n22363));
  jand g04341(.dina(n22363), .dinb(n338), .dout(n22364));
  jnot g04342(.din(n22364), .dout(n22365));
  jand g04343(.dina(n22239), .dinb(n22149), .dout(n22366));
  jxor g04344(.dina(n22171), .dinb(n22170), .dout(n22367));
  jand g04345(.dina(n22367), .dinb(n22238), .dout(n22368));
  jor  g04346(.dina(n22368), .dinb(n22366), .dout(n22369));
  jand g04347(.dina(n22369), .dinb(n337), .dout(n22370));
  jnot g04348(.din(n22370), .dout(n22371));
  jnot g04349(.din(n22154), .dout(n22372));
  jor  g04350(.dina(n22238), .dinb(n22372), .dout(n22373));
  jxor g04351(.dina(n22168), .dinb(n22167), .dout(n22374));
  jnot g04352(.din(n22374), .dout(n22375));
  jor  g04353(.dina(n22375), .dinb(n22239), .dout(n22376));
  jand g04354(.dina(n22376), .dinb(n22373), .dout(n22377));
  jor  g04355(.dina(n22377), .dinb(b3 ), .dout(n22378));
  jor  g04356(.dina(n22238), .dinb(n22164), .dout(n22379));
  jxor g04357(.dina(n22165), .dinb(n3322), .dout(n22380));
  jand g04358(.dina(n22380), .dinb(n22238), .dout(n22381));
  jnot g04359(.din(n22381), .dout(n22382));
  jand g04360(.dina(n22382), .dinb(n22379), .dout(n22383));
  jor  g04361(.dina(n22383), .dinb(b2 ), .dout(n22384));
  jand g04362(.dina(n22237), .dinb(n3545), .dout(n22385));
  jor  g04363(.dina(n22385), .dinb(n3320), .dout(n22386));
  jnot g04364(.din(n3548), .dout(n22387));
  jnot g04365(.din(n22043), .dout(n22388));
  jnot g04366(.din(n22050), .dout(n22389));
  jnot g04367(.din(n22055), .dout(n22390));
  jnot g04368(.din(n22060), .dout(n22391));
  jnot g04369(.din(n22065), .dout(n22392));
  jnot g04370(.din(n22070), .dout(n22393));
  jnot g04371(.din(n22075), .dout(n22394));
  jnot g04372(.din(n22080), .dout(n22395));
  jnot g04373(.din(n22085), .dout(n22396));
  jnot g04374(.din(n22090), .dout(n22397));
  jnot g04375(.din(n22095), .dout(n22398));
  jnot g04376(.din(n22100), .dout(n22399));
  jnot g04377(.din(n22105), .dout(n22400));
  jnot g04378(.din(n22110), .dout(n22401));
  jnot g04379(.din(n22115), .dout(n22402));
  jnot g04380(.din(n22120), .dout(n22403));
  jnot g04381(.din(n22125), .dout(n22404));
  jnot g04382(.din(n22130), .dout(n22405));
  jnot g04383(.din(n22135), .dout(n22406));
  jnot g04384(.din(n22140), .dout(n22407));
  jnot g04385(.din(n22145), .dout(n22408));
  jnot g04386(.din(n22150), .dout(n22409));
  jnot g04387(.din(n22155), .dout(n22410));
  jnot g04388(.din(n22161), .dout(n22411));
  jxor g04389(.dina(n22164), .dinb(n258), .dout(n22412));
  jor  g04390(.dina(n22412), .dinb(n3321), .dout(n22413));
  jand g04391(.dina(n22413), .dinb(n22411), .dout(n22414));
  jnot g04392(.din(n22168), .dout(n22415));
  jor  g04393(.dina(n22415), .dinb(n22414), .dout(n22416));
  jand g04394(.dina(n22416), .dinb(n22410), .dout(n22417));
  jnot g04395(.din(n22171), .dout(n22418));
  jor  g04396(.dina(n22418), .dinb(n22417), .dout(n22419));
  jand g04397(.dina(n22419), .dinb(n22409), .dout(n22420));
  jnot g04398(.din(n22174), .dout(n22421));
  jor  g04399(.dina(n22421), .dinb(n22420), .dout(n22422));
  jand g04400(.dina(n22422), .dinb(n22408), .dout(n22423));
  jnot g04401(.din(n22177), .dout(n22424));
  jor  g04402(.dina(n22424), .dinb(n22423), .dout(n22425));
  jand g04403(.dina(n22425), .dinb(n22407), .dout(n22426));
  jnot g04404(.din(n22180), .dout(n22427));
  jor  g04405(.dina(n22427), .dinb(n22426), .dout(n22428));
  jand g04406(.dina(n22428), .dinb(n22406), .dout(n22429));
  jnot g04407(.din(n22183), .dout(n22430));
  jor  g04408(.dina(n22430), .dinb(n22429), .dout(n22431));
  jand g04409(.dina(n22431), .dinb(n22405), .dout(n22432));
  jnot g04410(.din(n22186), .dout(n22433));
  jor  g04411(.dina(n22433), .dinb(n22432), .dout(n22434));
  jand g04412(.dina(n22434), .dinb(n22404), .dout(n22435));
  jnot g04413(.din(n22189), .dout(n22436));
  jor  g04414(.dina(n22436), .dinb(n22435), .dout(n22437));
  jand g04415(.dina(n22437), .dinb(n22403), .dout(n22438));
  jnot g04416(.din(n22192), .dout(n22439));
  jor  g04417(.dina(n22439), .dinb(n22438), .dout(n22440));
  jand g04418(.dina(n22440), .dinb(n22402), .dout(n22441));
  jnot g04419(.din(n22195), .dout(n22442));
  jor  g04420(.dina(n22442), .dinb(n22441), .dout(n22443));
  jand g04421(.dina(n22443), .dinb(n22401), .dout(n22444));
  jnot g04422(.din(n22198), .dout(n22445));
  jor  g04423(.dina(n22445), .dinb(n22444), .dout(n22446));
  jand g04424(.dina(n22446), .dinb(n22400), .dout(n22447));
  jnot g04425(.din(n22201), .dout(n22448));
  jor  g04426(.dina(n22448), .dinb(n22447), .dout(n22449));
  jand g04427(.dina(n22449), .dinb(n22399), .dout(n22450));
  jnot g04428(.din(n22204), .dout(n22451));
  jor  g04429(.dina(n22451), .dinb(n22450), .dout(n22452));
  jand g04430(.dina(n22452), .dinb(n22398), .dout(n22453));
  jnot g04431(.din(n22207), .dout(n22454));
  jor  g04432(.dina(n22454), .dinb(n22453), .dout(n22455));
  jand g04433(.dina(n22455), .dinb(n22397), .dout(n22456));
  jnot g04434(.din(n22210), .dout(n22457));
  jor  g04435(.dina(n22457), .dinb(n22456), .dout(n22458));
  jand g04436(.dina(n22458), .dinb(n22396), .dout(n22459));
  jnot g04437(.din(n22213), .dout(n22460));
  jor  g04438(.dina(n22460), .dinb(n22459), .dout(n22461));
  jand g04439(.dina(n22461), .dinb(n22395), .dout(n22462));
  jnot g04440(.din(n22216), .dout(n22463));
  jor  g04441(.dina(n22463), .dinb(n22462), .dout(n22464));
  jand g04442(.dina(n22464), .dinb(n22394), .dout(n22465));
  jnot g04443(.din(n22219), .dout(n22466));
  jor  g04444(.dina(n22466), .dinb(n22465), .dout(n22467));
  jand g04445(.dina(n22467), .dinb(n22393), .dout(n22468));
  jnot g04446(.din(n22222), .dout(n22469));
  jor  g04447(.dina(n22469), .dinb(n22468), .dout(n22470));
  jand g04448(.dina(n22470), .dinb(n22392), .dout(n22471));
  jnot g04449(.din(n22225), .dout(n22472));
  jor  g04450(.dina(n22472), .dinb(n22471), .dout(n22473));
  jand g04451(.dina(n22473), .dinb(n22391), .dout(n22474));
  jnot g04452(.din(n22228), .dout(n22475));
  jor  g04453(.dina(n22475), .dinb(n22474), .dout(n22476));
  jand g04454(.dina(n22476), .dinb(n22390), .dout(n22477));
  jnot g04455(.din(n22231), .dout(n22478));
  jor  g04456(.dina(n22478), .dinb(n22477), .dout(n22479));
  jand g04457(.dina(n22479), .dinb(n22389), .dout(n22480));
  jor  g04458(.dina(n22234), .dinb(n22480), .dout(n22481));
  jand g04459(.dina(n22481), .dinb(n22388), .dout(n22482));
  jor  g04460(.dina(n22482), .dinb(n22387), .dout(n22483));
  jand g04461(.dina(n22483), .dinb(n22386), .dout(n22484));
  jor  g04462(.dina(n22484), .dinb(b1 ), .dout(n22485));
  jxor g04463(.dina(n22484), .dinb(n258), .dout(n22486));
  jor  g04464(.dina(n22486), .dinb(n3554), .dout(n22487));
  jand g04465(.dina(n22487), .dinb(n22485), .dout(n22488));
  jxor g04466(.dina(n22383), .dinb(n348), .dout(n22489));
  jor  g04467(.dina(n22489), .dinb(n22488), .dout(n22490));
  jand g04468(.dina(n22490), .dinb(n22384), .dout(n22491));
  jxor g04469(.dina(n22377), .dinb(b3 ), .dout(n22492));
  jnot g04470(.din(n22492), .dout(n22493));
  jor  g04471(.dina(n22493), .dinb(n22491), .dout(n22494));
  jand g04472(.dina(n22494), .dinb(n22378), .dout(n22495));
  jxor g04473(.dina(n22369), .dinb(n337), .dout(n22496));
  jnot g04474(.din(n22496), .dout(n22497));
  jor  g04475(.dina(n22497), .dinb(n22495), .dout(n22498));
  jand g04476(.dina(n22498), .dinb(n22371), .dout(n22499));
  jxor g04477(.dina(n22363), .dinb(n338), .dout(n22500));
  jnot g04478(.din(n22500), .dout(n22501));
  jor  g04479(.dina(n22501), .dinb(n22499), .dout(n22502));
  jand g04480(.dina(n22502), .dinb(n22365), .dout(n22503));
  jxor g04481(.dina(n22357), .dinb(n334), .dout(n22504));
  jnot g04482(.din(n22504), .dout(n22505));
  jor  g04483(.dina(n22505), .dinb(n22503), .dout(n22506));
  jand g04484(.dina(n22506), .dinb(n22359), .dout(n22507));
  jxor g04485(.dina(n22351), .dinb(n335), .dout(n22508));
  jnot g04486(.din(n22508), .dout(n22509));
  jor  g04487(.dina(n22509), .dinb(n22507), .dout(n22510));
  jand g04488(.dina(n22510), .dinb(n22353), .dout(n22511));
  jxor g04489(.dina(n22345), .dinb(n323), .dout(n22512));
  jnot g04490(.din(n22512), .dout(n22513));
  jor  g04491(.dina(n22513), .dinb(n22511), .dout(n22514));
  jand g04492(.dina(n22514), .dinb(n22347), .dout(n22515));
  jxor g04493(.dina(n22339), .dinb(n324), .dout(n22516));
  jnot g04494(.din(n22516), .dout(n22517));
  jor  g04495(.dina(n22517), .dinb(n22515), .dout(n22518));
  jand g04496(.dina(n22518), .dinb(n22341), .dout(n22519));
  jxor g04497(.dina(n22333), .dinb(n325), .dout(n22520));
  jnot g04498(.din(n22520), .dout(n22521));
  jor  g04499(.dina(n22521), .dinb(n22519), .dout(n22522));
  jand g04500(.dina(n22522), .dinb(n22335), .dout(n22523));
  jxor g04501(.dina(n22327), .dinb(n439), .dout(n22524));
  jnot g04502(.din(n22524), .dout(n22525));
  jor  g04503(.dina(n22525), .dinb(n22523), .dout(n22526));
  jand g04504(.dina(n22526), .dinb(n22329), .dout(n22527));
  jxor g04505(.dina(n22321), .dinb(n440), .dout(n22528));
  jnot g04506(.din(n22528), .dout(n22529));
  jor  g04507(.dina(n22529), .dinb(n22527), .dout(n22530));
  jand g04508(.dina(n22530), .dinb(n22323), .dout(n22531));
  jxor g04509(.dina(n22315), .dinb(n435), .dout(n22532));
  jnot g04510(.din(n22532), .dout(n22533));
  jor  g04511(.dina(n22533), .dinb(n22531), .dout(n22534));
  jand g04512(.dina(n22534), .dinb(n22317), .dout(n22535));
  jxor g04513(.dina(n22309), .dinb(n436), .dout(n22536));
  jnot g04514(.din(n22536), .dout(n22537));
  jor  g04515(.dina(n22537), .dinb(n22535), .dout(n22538));
  jand g04516(.dina(n22538), .dinb(n22311), .dout(n22539));
  jxor g04517(.dina(n22303), .dinb(n432), .dout(n22540));
  jnot g04518(.din(n22540), .dout(n22541));
  jor  g04519(.dina(n22541), .dinb(n22539), .dout(n22542));
  jand g04520(.dina(n22542), .dinb(n22305), .dout(n22543));
  jxor g04521(.dina(n22297), .dinb(n433), .dout(n22544));
  jnot g04522(.din(n22544), .dout(n22545));
  jor  g04523(.dina(n22545), .dinb(n22543), .dout(n22546));
  jand g04524(.dina(n22546), .dinb(n22299), .dout(n22547));
  jxor g04525(.dina(n22291), .dinb(n421), .dout(n22548));
  jnot g04526(.din(n22548), .dout(n22549));
  jor  g04527(.dina(n22549), .dinb(n22547), .dout(n22550));
  jand g04528(.dina(n22550), .dinb(n22293), .dout(n22551));
  jxor g04529(.dina(n22285), .dinb(n422), .dout(n22552));
  jnot g04530(.din(n22552), .dout(n22553));
  jor  g04531(.dina(n22553), .dinb(n22551), .dout(n22554));
  jand g04532(.dina(n22554), .dinb(n22287), .dout(n22555));
  jxor g04533(.dina(n22279), .dinb(n416), .dout(n22556));
  jnot g04534(.din(n22556), .dout(n22557));
  jor  g04535(.dina(n22557), .dinb(n22555), .dout(n22558));
  jand g04536(.dina(n22558), .dinb(n22281), .dout(n22559));
  jxor g04537(.dina(n22273), .dinb(n417), .dout(n22560));
  jnot g04538(.din(n22560), .dout(n22561));
  jor  g04539(.dina(n22561), .dinb(n22559), .dout(n22562));
  jand g04540(.dina(n22562), .dinb(n22275), .dout(n22563));
  jxor g04541(.dina(n22267), .dinb(n2547), .dout(n22564));
  jnot g04542(.din(n22564), .dout(n22565));
  jor  g04543(.dina(n22565), .dinb(n22563), .dout(n22566));
  jand g04544(.dina(n22566), .dinb(n22269), .dout(n22567));
  jxor g04545(.dina(n22261), .dinb(n2714), .dout(n22568));
  jnot g04546(.din(n22568), .dout(n22569));
  jor  g04547(.dina(n22569), .dinb(n22567), .dout(n22570));
  jand g04548(.dina(n22570), .dinb(n22263), .dout(n22571));
  jxor g04549(.dina(n22255), .dinb(n405), .dout(n22572));
  jnot g04550(.din(n22572), .dout(n22573));
  jor  g04551(.dina(n22573), .dinb(n22571), .dout(n22574));
  jand g04552(.dina(n22574), .dinb(n22257), .dout(n22575));
  jxor g04553(.dina(n22249), .dinb(n406), .dout(n22576));
  jnot g04554(.din(n22576), .dout(n22577));
  jor  g04555(.dina(n22577), .dinb(n22575), .dout(n22578));
  jand g04556(.dina(n22578), .dinb(n22251), .dout(n22579));
  jnot g04557(.din(n22243), .dout(n22580));
  jand g04558(.dina(n22580), .dinb(b25 ), .dout(n22581));
  jor  g04559(.dina(n22581), .dinb(n22579), .dout(n22582));
  jand g04560(.dina(n22582), .dinb(n22245), .dout(n22583));
  jor  g04561(.dina(n22583), .dinb(n3403), .dout(n22584));
  jand g04562(.dina(n22584), .dinb(n22243), .dout(n22585));
  jnot g04563(.din(n22378), .dout(n22586));
  jnot g04564(.din(n22384), .dout(n22587));
  jnot g04565(.din(n3545), .dout(n22588));
  jor  g04566(.dina(n22482), .dinb(n22588), .dout(n22589));
  jand g04567(.dina(n22589), .dinb(a39 ), .dout(n22590));
  jnot g04568(.din(n22483), .dout(n22591));
  jor  g04569(.dina(n22591), .dinb(n22590), .dout(n22592));
  jand g04570(.dina(n22592), .dinb(n258), .dout(n22593));
  jxor g04571(.dina(n22484), .dinb(b1 ), .dout(n22594));
  jand g04572(.dina(n22594), .dinb(n3658), .dout(n22595));
  jor  g04573(.dina(n22595), .dinb(n22593), .dout(n22596));
  jxor g04574(.dina(n22383), .dinb(b2 ), .dout(n22597));
  jand g04575(.dina(n22597), .dinb(n22596), .dout(n22598));
  jor  g04576(.dina(n22598), .dinb(n22587), .dout(n22599));
  jand g04577(.dina(n22492), .dinb(n22599), .dout(n22600));
  jor  g04578(.dina(n22600), .dinb(n22586), .dout(n22601));
  jand g04579(.dina(n22496), .dinb(n22601), .dout(n22602));
  jor  g04580(.dina(n22602), .dinb(n22370), .dout(n22603));
  jand g04581(.dina(n22500), .dinb(n22603), .dout(n22604));
  jor  g04582(.dina(n22604), .dinb(n22364), .dout(n22605));
  jand g04583(.dina(n22504), .dinb(n22605), .dout(n22606));
  jor  g04584(.dina(n22606), .dinb(n22358), .dout(n22607));
  jand g04585(.dina(n22508), .dinb(n22607), .dout(n22608));
  jor  g04586(.dina(n22608), .dinb(n22352), .dout(n22609));
  jand g04587(.dina(n22512), .dinb(n22609), .dout(n22610));
  jor  g04588(.dina(n22610), .dinb(n22346), .dout(n22611));
  jand g04589(.dina(n22516), .dinb(n22611), .dout(n22612));
  jor  g04590(.dina(n22612), .dinb(n22340), .dout(n22613));
  jand g04591(.dina(n22520), .dinb(n22613), .dout(n22614));
  jor  g04592(.dina(n22614), .dinb(n22334), .dout(n22615));
  jand g04593(.dina(n22524), .dinb(n22615), .dout(n22616));
  jor  g04594(.dina(n22616), .dinb(n22328), .dout(n22617));
  jand g04595(.dina(n22528), .dinb(n22617), .dout(n22618));
  jor  g04596(.dina(n22618), .dinb(n22322), .dout(n22619));
  jand g04597(.dina(n22532), .dinb(n22619), .dout(n22620));
  jor  g04598(.dina(n22620), .dinb(n22316), .dout(n22621));
  jand g04599(.dina(n22536), .dinb(n22621), .dout(n22622));
  jor  g04600(.dina(n22622), .dinb(n22310), .dout(n22623));
  jand g04601(.dina(n22540), .dinb(n22623), .dout(n22624));
  jor  g04602(.dina(n22624), .dinb(n22304), .dout(n22625));
  jand g04603(.dina(n22544), .dinb(n22625), .dout(n22626));
  jor  g04604(.dina(n22626), .dinb(n22298), .dout(n22627));
  jand g04605(.dina(n22548), .dinb(n22627), .dout(n22628));
  jor  g04606(.dina(n22628), .dinb(n22292), .dout(n22629));
  jand g04607(.dina(n22552), .dinb(n22629), .dout(n22630));
  jor  g04608(.dina(n22630), .dinb(n22286), .dout(n22631));
  jand g04609(.dina(n22556), .dinb(n22631), .dout(n22632));
  jor  g04610(.dina(n22632), .dinb(n22280), .dout(n22633));
  jand g04611(.dina(n22560), .dinb(n22633), .dout(n22634));
  jor  g04612(.dina(n22634), .dinb(n22274), .dout(n22635));
  jand g04613(.dina(n22564), .dinb(n22635), .dout(n22636));
  jor  g04614(.dina(n22636), .dinb(n22268), .dout(n22637));
  jand g04615(.dina(n22568), .dinb(n22637), .dout(n22638));
  jor  g04616(.dina(n22638), .dinb(n22262), .dout(n22639));
  jand g04617(.dina(n22572), .dinb(n22639), .dout(n22640));
  jor  g04618(.dina(n22640), .dinb(n22256), .dout(n22641));
  jand g04619(.dina(n22576), .dinb(n22641), .dout(n22642));
  jor  g04620(.dina(n22642), .dinb(n22250), .dout(n22643));
  jand g04621(.dina(n22244), .dinb(n3402), .dout(n22644));
  jand g04622(.dina(n22644), .dinb(n22643), .dout(n22645));
  jor  g04623(.dina(n22645), .dinb(n22585), .dout(n22646));
  jnot g04624(.din(n22646), .dout(n22647));
  jand g04625(.dina(n22584), .dinb(n22249), .dout(n22648));
  jnot g04626(.din(n22581), .dout(n22649));
  jand g04627(.dina(n22649), .dinb(n22643), .dout(n22650));
  jor  g04628(.dina(n22650), .dinb(n22244), .dout(n22651));
  jand g04629(.dina(n22651), .dinb(n3402), .dout(n22652));
  jxor g04630(.dina(n22576), .dinb(n22641), .dout(n22653));
  jand g04631(.dina(n22653), .dinb(n22652), .dout(n22654));
  jor  g04632(.dina(n22654), .dinb(n22648), .dout(n22655));
  jand g04633(.dina(n22655), .dinb(n412), .dout(n22656));
  jnot g04634(.din(n22656), .dout(n22657));
  jand g04635(.dina(n22584), .dinb(n22255), .dout(n22658));
  jxor g04636(.dina(n22572), .dinb(n22639), .dout(n22659));
  jand g04637(.dina(n22659), .dinb(n22652), .dout(n22660));
  jor  g04638(.dina(n22660), .dinb(n22658), .dout(n22661));
  jand g04639(.dina(n22661), .dinb(n406), .dout(n22662));
  jnot g04640(.din(n22662), .dout(n22663));
  jand g04641(.dina(n22584), .dinb(n22261), .dout(n22664));
  jxor g04642(.dina(n22568), .dinb(n22637), .dout(n22665));
  jand g04643(.dina(n22665), .dinb(n22652), .dout(n22666));
  jor  g04644(.dina(n22666), .dinb(n22664), .dout(n22667));
  jand g04645(.dina(n22667), .dinb(n405), .dout(n22668));
  jnot g04646(.din(n22668), .dout(n22669));
  jand g04647(.dina(n22584), .dinb(n22267), .dout(n22670));
  jxor g04648(.dina(n22564), .dinb(n22635), .dout(n22671));
  jand g04649(.dina(n22671), .dinb(n22652), .dout(n22672));
  jor  g04650(.dina(n22672), .dinb(n22670), .dout(n22673));
  jand g04651(.dina(n22673), .dinb(n2714), .dout(n22674));
  jnot g04652(.din(n22674), .dout(n22675));
  jand g04653(.dina(n22584), .dinb(n22273), .dout(n22676));
  jxor g04654(.dina(n22560), .dinb(n22633), .dout(n22677));
  jand g04655(.dina(n22677), .dinb(n22652), .dout(n22678));
  jor  g04656(.dina(n22678), .dinb(n22676), .dout(n22679));
  jand g04657(.dina(n22679), .dinb(n2547), .dout(n22680));
  jnot g04658(.din(n22680), .dout(n22681));
  jand g04659(.dina(n22584), .dinb(n22279), .dout(n22682));
  jxor g04660(.dina(n22556), .dinb(n22631), .dout(n22683));
  jand g04661(.dina(n22683), .dinb(n22652), .dout(n22684));
  jor  g04662(.dina(n22684), .dinb(n22682), .dout(n22685));
  jand g04663(.dina(n22685), .dinb(n417), .dout(n22686));
  jnot g04664(.din(n22686), .dout(n22687));
  jand g04665(.dina(n22584), .dinb(n22285), .dout(n22688));
  jxor g04666(.dina(n22552), .dinb(n22629), .dout(n22689));
  jand g04667(.dina(n22689), .dinb(n22652), .dout(n22690));
  jor  g04668(.dina(n22690), .dinb(n22688), .dout(n22691));
  jand g04669(.dina(n22691), .dinb(n416), .dout(n22692));
  jnot g04670(.din(n22692), .dout(n22693));
  jand g04671(.dina(n22584), .dinb(n22291), .dout(n22694));
  jxor g04672(.dina(n22548), .dinb(n22627), .dout(n22695));
  jand g04673(.dina(n22695), .dinb(n22652), .dout(n22696));
  jor  g04674(.dina(n22696), .dinb(n22694), .dout(n22697));
  jand g04675(.dina(n22697), .dinb(n422), .dout(n22698));
  jnot g04676(.din(n22698), .dout(n22699));
  jand g04677(.dina(n22584), .dinb(n22297), .dout(n22700));
  jxor g04678(.dina(n22544), .dinb(n22625), .dout(n22701));
  jand g04679(.dina(n22701), .dinb(n22652), .dout(n22702));
  jor  g04680(.dina(n22702), .dinb(n22700), .dout(n22703));
  jand g04681(.dina(n22703), .dinb(n421), .dout(n22704));
  jnot g04682(.din(n22704), .dout(n22705));
  jand g04683(.dina(n22584), .dinb(n22303), .dout(n22706));
  jxor g04684(.dina(n22540), .dinb(n22623), .dout(n22707));
  jand g04685(.dina(n22707), .dinb(n22652), .dout(n22708));
  jor  g04686(.dina(n22708), .dinb(n22706), .dout(n22709));
  jand g04687(.dina(n22709), .dinb(n433), .dout(n22710));
  jnot g04688(.din(n22710), .dout(n22711));
  jand g04689(.dina(n22584), .dinb(n22309), .dout(n22712));
  jxor g04690(.dina(n22536), .dinb(n22621), .dout(n22713));
  jand g04691(.dina(n22713), .dinb(n22652), .dout(n22714));
  jor  g04692(.dina(n22714), .dinb(n22712), .dout(n22715));
  jand g04693(.dina(n22715), .dinb(n432), .dout(n22716));
  jnot g04694(.din(n22716), .dout(n22717));
  jand g04695(.dina(n22584), .dinb(n22315), .dout(n22718));
  jxor g04696(.dina(n22532), .dinb(n22619), .dout(n22719));
  jand g04697(.dina(n22719), .dinb(n22652), .dout(n22720));
  jor  g04698(.dina(n22720), .dinb(n22718), .dout(n22721));
  jand g04699(.dina(n22721), .dinb(n436), .dout(n22722));
  jnot g04700(.din(n22722), .dout(n22723));
  jand g04701(.dina(n22584), .dinb(n22321), .dout(n22724));
  jxor g04702(.dina(n22528), .dinb(n22617), .dout(n22725));
  jand g04703(.dina(n22725), .dinb(n22652), .dout(n22726));
  jor  g04704(.dina(n22726), .dinb(n22724), .dout(n22727));
  jand g04705(.dina(n22727), .dinb(n435), .dout(n22728));
  jnot g04706(.din(n22728), .dout(n22729));
  jand g04707(.dina(n22584), .dinb(n22327), .dout(n22730));
  jxor g04708(.dina(n22524), .dinb(n22615), .dout(n22731));
  jand g04709(.dina(n22731), .dinb(n22652), .dout(n22732));
  jor  g04710(.dina(n22732), .dinb(n22730), .dout(n22733));
  jand g04711(.dina(n22733), .dinb(n440), .dout(n22734));
  jnot g04712(.din(n22734), .dout(n22735));
  jand g04713(.dina(n22584), .dinb(n22333), .dout(n22736));
  jxor g04714(.dina(n22520), .dinb(n22613), .dout(n22737));
  jand g04715(.dina(n22737), .dinb(n22652), .dout(n22738));
  jor  g04716(.dina(n22738), .dinb(n22736), .dout(n22739));
  jand g04717(.dina(n22739), .dinb(n439), .dout(n22740));
  jnot g04718(.din(n22740), .dout(n22741));
  jand g04719(.dina(n22584), .dinb(n22339), .dout(n22742));
  jxor g04720(.dina(n22516), .dinb(n22611), .dout(n22743));
  jand g04721(.dina(n22743), .dinb(n22652), .dout(n22744));
  jor  g04722(.dina(n22744), .dinb(n22742), .dout(n22745));
  jand g04723(.dina(n22745), .dinb(n325), .dout(n22746));
  jnot g04724(.din(n22746), .dout(n22747));
  jand g04725(.dina(n22584), .dinb(n22345), .dout(n22748));
  jxor g04726(.dina(n22512), .dinb(n22609), .dout(n22749));
  jand g04727(.dina(n22749), .dinb(n22652), .dout(n22750));
  jor  g04728(.dina(n22750), .dinb(n22748), .dout(n22751));
  jand g04729(.dina(n22751), .dinb(n324), .dout(n22752));
  jnot g04730(.din(n22752), .dout(n22753));
  jand g04731(.dina(n22584), .dinb(n22351), .dout(n22754));
  jxor g04732(.dina(n22508), .dinb(n22607), .dout(n22755));
  jand g04733(.dina(n22755), .dinb(n22652), .dout(n22756));
  jor  g04734(.dina(n22756), .dinb(n22754), .dout(n22757));
  jand g04735(.dina(n22757), .dinb(n323), .dout(n22758));
  jnot g04736(.din(n22758), .dout(n22759));
  jand g04737(.dina(n22584), .dinb(n22357), .dout(n22760));
  jxor g04738(.dina(n22504), .dinb(n22605), .dout(n22761));
  jand g04739(.dina(n22761), .dinb(n22652), .dout(n22762));
  jor  g04740(.dina(n22762), .dinb(n22760), .dout(n22763));
  jand g04741(.dina(n22763), .dinb(n335), .dout(n22764));
  jnot g04742(.din(n22764), .dout(n22765));
  jand g04743(.dina(n22584), .dinb(n22363), .dout(n22766));
  jxor g04744(.dina(n22500), .dinb(n22603), .dout(n22767));
  jand g04745(.dina(n22767), .dinb(n22652), .dout(n22768));
  jor  g04746(.dina(n22768), .dinb(n22766), .dout(n22769));
  jand g04747(.dina(n22769), .dinb(n334), .dout(n22770));
  jnot g04748(.din(n22770), .dout(n22771));
  jand g04749(.dina(n22584), .dinb(n22369), .dout(n22772));
  jxor g04750(.dina(n22496), .dinb(n22601), .dout(n22773));
  jand g04751(.dina(n22773), .dinb(n22652), .dout(n22774));
  jor  g04752(.dina(n22774), .dinb(n22772), .dout(n22775));
  jand g04753(.dina(n22775), .dinb(n338), .dout(n22776));
  jnot g04754(.din(n22776), .dout(n22777));
  jor  g04755(.dina(n22652), .dinb(n22377), .dout(n22778));
  jxor g04756(.dina(n22492), .dinb(n22599), .dout(n22779));
  jand g04757(.dina(n22779), .dinb(n22652), .dout(n22780));
  jnot g04758(.din(n22780), .dout(n22781));
  jand g04759(.dina(n22781), .dinb(n22778), .dout(n22782));
  jnot g04760(.din(n22782), .dout(n22783));
  jand g04761(.dina(n22783), .dinb(n337), .dout(n22784));
  jnot g04762(.din(n22784), .dout(n22785));
  jor  g04763(.dina(n22652), .dinb(n22383), .dout(n22786));
  jxor g04764(.dina(n22597), .dinb(n22596), .dout(n22787));
  jnot g04765(.din(n22787), .dout(n22788));
  jor  g04766(.dina(n22788), .dinb(n22584), .dout(n22789));
  jand g04767(.dina(n22789), .dinb(n22786), .dout(n22790));
  jnot g04768(.din(n22790), .dout(n22791));
  jand g04769(.dina(n22791), .dinb(n344), .dout(n22792));
  jnot g04770(.din(n22792), .dout(n22793));
  jand g04771(.dina(n22584), .dinb(n22592), .dout(n22794));
  jxor g04772(.dina(n22594), .dinb(n3658), .dout(n22795));
  jand g04773(.dina(n22795), .dinb(n22652), .dout(n22796));
  jor  g04774(.dina(n22796), .dinb(n22794), .dout(n22797));
  jand g04775(.dina(n22797), .dinb(n348), .dout(n22798));
  jnot g04776(.din(n22798), .dout(n22799));
  jnot g04777(.din(n3840), .dout(n22800));
  jor  g04778(.dina(n22583), .dinb(n22800), .dout(n22801));
  jand g04779(.dina(n22801), .dinb(a38 ), .dout(n22802));
  jand g04780(.dina(n22652), .dinb(n3554), .dout(n22803));
  jor  g04781(.dina(n22803), .dinb(n22802), .dout(n22804));
  jand g04782(.dina(n22804), .dinb(n258), .dout(n22805));
  jnot g04783(.din(n22805), .dout(n22806));
  jand g04784(.dina(n22651), .dinb(n3840), .dout(n22807));
  jor  g04785(.dina(n22807), .dinb(n3553), .dout(n22808));
  jor  g04786(.dina(n22584), .dinb(n3658), .dout(n22809));
  jand g04787(.dina(n22809), .dinb(n22808), .dout(n22810));
  jxor g04788(.dina(n22810), .dinb(n258), .dout(n22811));
  jor  g04789(.dina(n22811), .dinb(n3848), .dout(n22812));
  jand g04790(.dina(n22812), .dinb(n22806), .dout(n22813));
  jxor g04791(.dina(n22797), .dinb(n348), .dout(n22814));
  jnot g04792(.din(n22814), .dout(n22815));
  jor  g04793(.dina(n22815), .dinb(n22813), .dout(n22816));
  jand g04794(.dina(n22816), .dinb(n22799), .dout(n22817));
  jxor g04795(.dina(n22790), .dinb(b3 ), .dout(n22818));
  jnot g04796(.din(n22818), .dout(n22819));
  jor  g04797(.dina(n22819), .dinb(n22817), .dout(n22820));
  jand g04798(.dina(n22820), .dinb(n22793), .dout(n22821));
  jxor g04799(.dina(n22782), .dinb(b4 ), .dout(n22822));
  jnot g04800(.din(n22822), .dout(n22823));
  jor  g04801(.dina(n22823), .dinb(n22821), .dout(n22824));
  jand g04802(.dina(n22824), .dinb(n22785), .dout(n22825));
  jxor g04803(.dina(n22775), .dinb(n338), .dout(n22826));
  jnot g04804(.din(n22826), .dout(n22827));
  jor  g04805(.dina(n22827), .dinb(n22825), .dout(n22828));
  jand g04806(.dina(n22828), .dinb(n22777), .dout(n22829));
  jxor g04807(.dina(n22769), .dinb(n334), .dout(n22830));
  jnot g04808(.din(n22830), .dout(n22831));
  jor  g04809(.dina(n22831), .dinb(n22829), .dout(n22832));
  jand g04810(.dina(n22832), .dinb(n22771), .dout(n22833));
  jxor g04811(.dina(n22763), .dinb(n335), .dout(n22834));
  jnot g04812(.din(n22834), .dout(n22835));
  jor  g04813(.dina(n22835), .dinb(n22833), .dout(n22836));
  jand g04814(.dina(n22836), .dinb(n22765), .dout(n22837));
  jxor g04815(.dina(n22757), .dinb(n323), .dout(n22838));
  jnot g04816(.din(n22838), .dout(n22839));
  jor  g04817(.dina(n22839), .dinb(n22837), .dout(n22840));
  jand g04818(.dina(n22840), .dinb(n22759), .dout(n22841));
  jxor g04819(.dina(n22751), .dinb(n324), .dout(n22842));
  jnot g04820(.din(n22842), .dout(n22843));
  jor  g04821(.dina(n22843), .dinb(n22841), .dout(n22844));
  jand g04822(.dina(n22844), .dinb(n22753), .dout(n22845));
  jxor g04823(.dina(n22745), .dinb(n325), .dout(n22846));
  jnot g04824(.din(n22846), .dout(n22847));
  jor  g04825(.dina(n22847), .dinb(n22845), .dout(n22848));
  jand g04826(.dina(n22848), .dinb(n22747), .dout(n22849));
  jxor g04827(.dina(n22739), .dinb(n439), .dout(n22850));
  jnot g04828(.din(n22850), .dout(n22851));
  jor  g04829(.dina(n22851), .dinb(n22849), .dout(n22852));
  jand g04830(.dina(n22852), .dinb(n22741), .dout(n22853));
  jxor g04831(.dina(n22733), .dinb(n440), .dout(n22854));
  jnot g04832(.din(n22854), .dout(n22855));
  jor  g04833(.dina(n22855), .dinb(n22853), .dout(n22856));
  jand g04834(.dina(n22856), .dinb(n22735), .dout(n22857));
  jxor g04835(.dina(n22727), .dinb(n435), .dout(n22858));
  jnot g04836(.din(n22858), .dout(n22859));
  jor  g04837(.dina(n22859), .dinb(n22857), .dout(n22860));
  jand g04838(.dina(n22860), .dinb(n22729), .dout(n22861));
  jxor g04839(.dina(n22721), .dinb(n436), .dout(n22862));
  jnot g04840(.din(n22862), .dout(n22863));
  jor  g04841(.dina(n22863), .dinb(n22861), .dout(n22864));
  jand g04842(.dina(n22864), .dinb(n22723), .dout(n22865));
  jxor g04843(.dina(n22715), .dinb(n432), .dout(n22866));
  jnot g04844(.din(n22866), .dout(n22867));
  jor  g04845(.dina(n22867), .dinb(n22865), .dout(n22868));
  jand g04846(.dina(n22868), .dinb(n22717), .dout(n22869));
  jxor g04847(.dina(n22709), .dinb(n433), .dout(n22870));
  jnot g04848(.din(n22870), .dout(n22871));
  jor  g04849(.dina(n22871), .dinb(n22869), .dout(n22872));
  jand g04850(.dina(n22872), .dinb(n22711), .dout(n22873));
  jxor g04851(.dina(n22703), .dinb(n421), .dout(n22874));
  jnot g04852(.din(n22874), .dout(n22875));
  jor  g04853(.dina(n22875), .dinb(n22873), .dout(n22876));
  jand g04854(.dina(n22876), .dinb(n22705), .dout(n22877));
  jxor g04855(.dina(n22697), .dinb(n422), .dout(n22878));
  jnot g04856(.din(n22878), .dout(n22879));
  jor  g04857(.dina(n22879), .dinb(n22877), .dout(n22880));
  jand g04858(.dina(n22880), .dinb(n22699), .dout(n22881));
  jxor g04859(.dina(n22691), .dinb(n416), .dout(n22882));
  jnot g04860(.din(n22882), .dout(n22883));
  jor  g04861(.dina(n22883), .dinb(n22881), .dout(n22884));
  jand g04862(.dina(n22884), .dinb(n22693), .dout(n22885));
  jxor g04863(.dina(n22685), .dinb(n417), .dout(n22886));
  jnot g04864(.din(n22886), .dout(n22887));
  jor  g04865(.dina(n22887), .dinb(n22885), .dout(n22888));
  jand g04866(.dina(n22888), .dinb(n22687), .dout(n22889));
  jxor g04867(.dina(n22679), .dinb(n2547), .dout(n22890));
  jnot g04868(.din(n22890), .dout(n22891));
  jor  g04869(.dina(n22891), .dinb(n22889), .dout(n22892));
  jand g04870(.dina(n22892), .dinb(n22681), .dout(n22893));
  jxor g04871(.dina(n22673), .dinb(n2714), .dout(n22894));
  jnot g04872(.din(n22894), .dout(n22895));
  jor  g04873(.dina(n22895), .dinb(n22893), .dout(n22896));
  jand g04874(.dina(n22896), .dinb(n22675), .dout(n22897));
  jxor g04875(.dina(n22667), .dinb(n405), .dout(n22898));
  jnot g04876(.din(n22898), .dout(n22899));
  jor  g04877(.dina(n22899), .dinb(n22897), .dout(n22900));
  jand g04878(.dina(n22900), .dinb(n22669), .dout(n22901));
  jxor g04879(.dina(n22661), .dinb(n406), .dout(n22902));
  jnot g04880(.din(n22902), .dout(n22903));
  jor  g04881(.dina(n22903), .dinb(n22901), .dout(n22904));
  jand g04882(.dina(n22904), .dinb(n22663), .dout(n22905));
  jxor g04883(.dina(n22655), .dinb(n412), .dout(n22906));
  jnot g04884(.din(n22906), .dout(n22907));
  jor  g04885(.dina(n22907), .dinb(n22905), .dout(n22908));
  jand g04886(.dina(n22908), .dinb(n22657), .dout(n22909));
  jnot g04887(.din(n3716), .dout(n22910));
  jxor g04888(.dina(n22646), .dinb(b26 ), .dout(n22911));
  jor  g04889(.dina(n22911), .dinb(n22910), .dout(n22912));
  jor  g04890(.dina(n22912), .dinb(n22909), .dout(n22913));
  jand g04891(.dina(n22913), .dinb(n22647), .dout(n22914));
  jxor g04892(.dina(n22810), .dinb(b1 ), .dout(n22915));
  jand g04893(.dina(n22915), .dinb(n3849), .dout(n22916));
  jor  g04894(.dina(n22916), .dinb(n22805), .dout(n22917));
  jand g04895(.dina(n22814), .dinb(n22917), .dout(n22918));
  jor  g04896(.dina(n22918), .dinb(n22798), .dout(n22919));
  jand g04897(.dina(n22818), .dinb(n22919), .dout(n22920));
  jor  g04898(.dina(n22920), .dinb(n22792), .dout(n22921));
  jand g04899(.dina(n22822), .dinb(n22921), .dout(n22922));
  jor  g04900(.dina(n22922), .dinb(n22784), .dout(n22923));
  jand g04901(.dina(n22826), .dinb(n22923), .dout(n22924));
  jor  g04902(.dina(n22924), .dinb(n22776), .dout(n22925));
  jand g04903(.dina(n22830), .dinb(n22925), .dout(n22926));
  jor  g04904(.dina(n22926), .dinb(n22770), .dout(n22927));
  jand g04905(.dina(n22834), .dinb(n22927), .dout(n22928));
  jor  g04906(.dina(n22928), .dinb(n22764), .dout(n22929));
  jand g04907(.dina(n22838), .dinb(n22929), .dout(n22930));
  jor  g04908(.dina(n22930), .dinb(n22758), .dout(n22931));
  jand g04909(.dina(n22842), .dinb(n22931), .dout(n22932));
  jor  g04910(.dina(n22932), .dinb(n22752), .dout(n22933));
  jand g04911(.dina(n22846), .dinb(n22933), .dout(n22934));
  jor  g04912(.dina(n22934), .dinb(n22746), .dout(n22935));
  jand g04913(.dina(n22850), .dinb(n22935), .dout(n22936));
  jor  g04914(.dina(n22936), .dinb(n22740), .dout(n22937));
  jand g04915(.dina(n22854), .dinb(n22937), .dout(n22938));
  jor  g04916(.dina(n22938), .dinb(n22734), .dout(n22939));
  jand g04917(.dina(n22858), .dinb(n22939), .dout(n22940));
  jor  g04918(.dina(n22940), .dinb(n22728), .dout(n22941));
  jand g04919(.dina(n22862), .dinb(n22941), .dout(n22942));
  jor  g04920(.dina(n22942), .dinb(n22722), .dout(n22943));
  jand g04921(.dina(n22866), .dinb(n22943), .dout(n22944));
  jor  g04922(.dina(n22944), .dinb(n22716), .dout(n22945));
  jand g04923(.dina(n22870), .dinb(n22945), .dout(n22946));
  jor  g04924(.dina(n22946), .dinb(n22710), .dout(n22947));
  jand g04925(.dina(n22874), .dinb(n22947), .dout(n22948));
  jor  g04926(.dina(n22948), .dinb(n22704), .dout(n22949));
  jand g04927(.dina(n22878), .dinb(n22949), .dout(n22950));
  jor  g04928(.dina(n22950), .dinb(n22698), .dout(n22951));
  jand g04929(.dina(n22882), .dinb(n22951), .dout(n22952));
  jor  g04930(.dina(n22952), .dinb(n22692), .dout(n22953));
  jand g04931(.dina(n22886), .dinb(n22953), .dout(n22954));
  jor  g04932(.dina(n22954), .dinb(n22686), .dout(n22955));
  jand g04933(.dina(n22890), .dinb(n22955), .dout(n22956));
  jor  g04934(.dina(n22956), .dinb(n22680), .dout(n22957));
  jand g04935(.dina(n22894), .dinb(n22957), .dout(n22958));
  jor  g04936(.dina(n22958), .dinb(n22674), .dout(n22959));
  jand g04937(.dina(n22898), .dinb(n22959), .dout(n22960));
  jor  g04938(.dina(n22960), .dinb(n22668), .dout(n22961));
  jand g04939(.dina(n22902), .dinb(n22961), .dout(n22962));
  jor  g04940(.dina(n22962), .dinb(n22662), .dout(n22963));
  jand g04941(.dina(n22906), .dinb(n22963), .dout(n22964));
  jor  g04942(.dina(n22964), .dinb(n22656), .dout(n22965));
  jnot g04943(.din(n22912), .dout(n22966));
  jand g04944(.dina(n22966), .dinb(n22965), .dout(n22967));
  jand g04945(.dina(n22646), .dinb(n3402), .dout(n22968));
  jor  g04946(.dina(n22968), .dinb(n22967), .dout(n22969));
  jxor g04947(.dina(n22911), .dinb(n22965), .dout(n22970));
  jand g04948(.dina(n22970), .dinb(n22969), .dout(n22971));
  jor  g04949(.dina(n22971), .dinb(n22914), .dout(n22972));
  jnot g04950(.din(n22972), .dout(n22973));
  jand g04951(.dina(n22972), .dinb(b27 ), .dout(n22974));
  jnot g04952(.din(n22974), .dout(n22975));
  jand g04953(.dina(n22973), .dinb(n409), .dout(n22976));
  jnot g04954(.din(n22968), .dout(n22977));
  jand g04955(.dina(n22977), .dinb(n22913), .dout(n22978));
  jand g04956(.dina(n22978), .dinb(n22655), .dout(n22979));
  jxor g04957(.dina(n22906), .dinb(n22963), .dout(n22980));
  jand g04958(.dina(n22980), .dinb(n22969), .dout(n22981));
  jor  g04959(.dina(n22981), .dinb(n22979), .dout(n22982));
  jand g04960(.dina(n22982), .dinb(n413), .dout(n22983));
  jand g04961(.dina(n22978), .dinb(n22661), .dout(n22984));
  jxor g04962(.dina(n22902), .dinb(n22961), .dout(n22985));
  jand g04963(.dina(n22985), .dinb(n22969), .dout(n22986));
  jor  g04964(.dina(n22986), .dinb(n22984), .dout(n22987));
  jand g04965(.dina(n22987), .dinb(n412), .dout(n22988));
  jand g04966(.dina(n22978), .dinb(n22667), .dout(n22989));
  jxor g04967(.dina(n22898), .dinb(n22959), .dout(n22990));
  jand g04968(.dina(n22990), .dinb(n22969), .dout(n22991));
  jor  g04969(.dina(n22991), .dinb(n22989), .dout(n22992));
  jand g04970(.dina(n22992), .dinb(n406), .dout(n22993));
  jand g04971(.dina(n22978), .dinb(n22673), .dout(n22994));
  jxor g04972(.dina(n22894), .dinb(n22957), .dout(n22995));
  jand g04973(.dina(n22995), .dinb(n22969), .dout(n22996));
  jor  g04974(.dina(n22996), .dinb(n22994), .dout(n22997));
  jand g04975(.dina(n22997), .dinb(n405), .dout(n22998));
  jand g04976(.dina(n22978), .dinb(n22679), .dout(n22999));
  jxor g04977(.dina(n22890), .dinb(n22955), .dout(n23000));
  jand g04978(.dina(n23000), .dinb(n22969), .dout(n23001));
  jor  g04979(.dina(n23001), .dinb(n22999), .dout(n23002));
  jand g04980(.dina(n23002), .dinb(n2714), .dout(n23003));
  jand g04981(.dina(n22978), .dinb(n22685), .dout(n23004));
  jxor g04982(.dina(n22886), .dinb(n22953), .dout(n23005));
  jand g04983(.dina(n23005), .dinb(n22969), .dout(n23006));
  jor  g04984(.dina(n23006), .dinb(n23004), .dout(n23007));
  jand g04985(.dina(n23007), .dinb(n2547), .dout(n23008));
  jand g04986(.dina(n22978), .dinb(n22691), .dout(n23009));
  jxor g04987(.dina(n22882), .dinb(n22951), .dout(n23010));
  jand g04988(.dina(n23010), .dinb(n22969), .dout(n23011));
  jor  g04989(.dina(n23011), .dinb(n23009), .dout(n23012));
  jand g04990(.dina(n23012), .dinb(n417), .dout(n23013));
  jand g04991(.dina(n22978), .dinb(n22697), .dout(n23014));
  jxor g04992(.dina(n22878), .dinb(n22949), .dout(n23015));
  jand g04993(.dina(n23015), .dinb(n22969), .dout(n23016));
  jor  g04994(.dina(n23016), .dinb(n23014), .dout(n23017));
  jand g04995(.dina(n23017), .dinb(n416), .dout(n23018));
  jand g04996(.dina(n22978), .dinb(n22703), .dout(n23019));
  jxor g04997(.dina(n22874), .dinb(n22947), .dout(n23020));
  jand g04998(.dina(n23020), .dinb(n22969), .dout(n23021));
  jor  g04999(.dina(n23021), .dinb(n23019), .dout(n23022));
  jand g05000(.dina(n23022), .dinb(n422), .dout(n23023));
  jand g05001(.dina(n22978), .dinb(n22709), .dout(n23024));
  jxor g05002(.dina(n22870), .dinb(n22945), .dout(n23025));
  jand g05003(.dina(n23025), .dinb(n22969), .dout(n23026));
  jor  g05004(.dina(n23026), .dinb(n23024), .dout(n23027));
  jand g05005(.dina(n23027), .dinb(n421), .dout(n23028));
  jand g05006(.dina(n22978), .dinb(n22715), .dout(n23029));
  jxor g05007(.dina(n22866), .dinb(n22943), .dout(n23030));
  jand g05008(.dina(n23030), .dinb(n22969), .dout(n23031));
  jor  g05009(.dina(n23031), .dinb(n23029), .dout(n23032));
  jand g05010(.dina(n23032), .dinb(n433), .dout(n23033));
  jand g05011(.dina(n22978), .dinb(n22721), .dout(n23034));
  jxor g05012(.dina(n22862), .dinb(n22941), .dout(n23035));
  jand g05013(.dina(n23035), .dinb(n22969), .dout(n23036));
  jor  g05014(.dina(n23036), .dinb(n23034), .dout(n23037));
  jand g05015(.dina(n23037), .dinb(n432), .dout(n23038));
  jand g05016(.dina(n22978), .dinb(n22727), .dout(n23039));
  jxor g05017(.dina(n22858), .dinb(n22939), .dout(n23040));
  jand g05018(.dina(n23040), .dinb(n22969), .dout(n23041));
  jor  g05019(.dina(n23041), .dinb(n23039), .dout(n23042));
  jand g05020(.dina(n23042), .dinb(n436), .dout(n23043));
  jand g05021(.dina(n22978), .dinb(n22733), .dout(n23044));
  jxor g05022(.dina(n22854), .dinb(n22937), .dout(n23045));
  jand g05023(.dina(n23045), .dinb(n22969), .dout(n23046));
  jor  g05024(.dina(n23046), .dinb(n23044), .dout(n23047));
  jand g05025(.dina(n23047), .dinb(n435), .dout(n23048));
  jand g05026(.dina(n22978), .dinb(n22739), .dout(n23049));
  jxor g05027(.dina(n22850), .dinb(n22935), .dout(n23050));
  jand g05028(.dina(n23050), .dinb(n22969), .dout(n23051));
  jor  g05029(.dina(n23051), .dinb(n23049), .dout(n23052));
  jand g05030(.dina(n23052), .dinb(n440), .dout(n23053));
  jand g05031(.dina(n22978), .dinb(n22745), .dout(n23054));
  jxor g05032(.dina(n22846), .dinb(n22933), .dout(n23055));
  jand g05033(.dina(n23055), .dinb(n22969), .dout(n23056));
  jor  g05034(.dina(n23056), .dinb(n23054), .dout(n23057));
  jand g05035(.dina(n23057), .dinb(n439), .dout(n23058));
  jand g05036(.dina(n22978), .dinb(n22751), .dout(n23059));
  jxor g05037(.dina(n22842), .dinb(n22931), .dout(n23060));
  jand g05038(.dina(n23060), .dinb(n22969), .dout(n23061));
  jor  g05039(.dina(n23061), .dinb(n23059), .dout(n23062));
  jand g05040(.dina(n23062), .dinb(n325), .dout(n23063));
  jand g05041(.dina(n22978), .dinb(n22757), .dout(n23064));
  jxor g05042(.dina(n22838), .dinb(n22929), .dout(n23065));
  jand g05043(.dina(n23065), .dinb(n22969), .dout(n23066));
  jor  g05044(.dina(n23066), .dinb(n23064), .dout(n23067));
  jand g05045(.dina(n23067), .dinb(n324), .dout(n23068));
  jand g05046(.dina(n22978), .dinb(n22763), .dout(n23069));
  jxor g05047(.dina(n22834), .dinb(n22927), .dout(n23070));
  jand g05048(.dina(n23070), .dinb(n22969), .dout(n23071));
  jor  g05049(.dina(n23071), .dinb(n23069), .dout(n23072));
  jand g05050(.dina(n23072), .dinb(n323), .dout(n23073));
  jand g05051(.dina(n22978), .dinb(n22769), .dout(n23074));
  jxor g05052(.dina(n22830), .dinb(n22925), .dout(n23075));
  jand g05053(.dina(n23075), .dinb(n22969), .dout(n23076));
  jor  g05054(.dina(n23076), .dinb(n23074), .dout(n23077));
  jand g05055(.dina(n23077), .dinb(n335), .dout(n23078));
  jand g05056(.dina(n22978), .dinb(n22775), .dout(n23079));
  jxor g05057(.dina(n22826), .dinb(n22923), .dout(n23080));
  jand g05058(.dina(n23080), .dinb(n22969), .dout(n23081));
  jor  g05059(.dina(n23081), .dinb(n23079), .dout(n23082));
  jand g05060(.dina(n23082), .dinb(n334), .dout(n23083));
  jand g05061(.dina(n22978), .dinb(n22783), .dout(n23084));
  jxor g05062(.dina(n22822), .dinb(n22921), .dout(n23085));
  jand g05063(.dina(n23085), .dinb(n22969), .dout(n23086));
  jor  g05064(.dina(n23086), .dinb(n23084), .dout(n23087));
  jand g05065(.dina(n23087), .dinb(n338), .dout(n23088));
  jand g05066(.dina(n22978), .dinb(n22791), .dout(n23089));
  jxor g05067(.dina(n22818), .dinb(n22919), .dout(n23090));
  jand g05068(.dina(n23090), .dinb(n22969), .dout(n23091));
  jor  g05069(.dina(n23091), .dinb(n23089), .dout(n23092));
  jand g05070(.dina(n23092), .dinb(n337), .dout(n23093));
  jand g05071(.dina(n22978), .dinb(n22797), .dout(n23094));
  jxor g05072(.dina(n22814), .dinb(n22917), .dout(n23095));
  jand g05073(.dina(n23095), .dinb(n22969), .dout(n23096));
  jor  g05074(.dina(n23096), .dinb(n23094), .dout(n23097));
  jand g05075(.dina(n23097), .dinb(n344), .dout(n23098));
  jand g05076(.dina(n22978), .dinb(n22804), .dout(n23099));
  jxor g05077(.dina(n22915), .dinb(n3849), .dout(n23100));
  jand g05078(.dina(n23100), .dinb(n22969), .dout(n23101));
  jor  g05079(.dina(n23101), .dinb(n23099), .dout(n23102));
  jand g05080(.dina(n23102), .dinb(n348), .dout(n23103));
  jor  g05081(.dina(n22978), .dinb(n18364), .dout(n23104));
  jand g05082(.dina(n23104), .dinb(a37 ), .dout(n23105));
  jor  g05083(.dina(n22978), .dinb(n3849), .dout(n23106));
  jnot g05084(.din(n23106), .dout(n23107));
  jor  g05085(.dina(n23107), .dinb(n23105), .dout(n23108));
  jand g05086(.dina(n23108), .dinb(n258), .dout(n23109));
  jand g05087(.dina(n22969), .dinb(b0 ), .dout(n23110));
  jor  g05088(.dina(n23110), .dinb(n3847), .dout(n23111));
  jand g05089(.dina(n23106), .dinb(n23111), .dout(n23112));
  jxor g05090(.dina(n23112), .dinb(b1 ), .dout(n23113));
  jand g05091(.dina(n23113), .dinb(n4075), .dout(n23114));
  jor  g05092(.dina(n23114), .dinb(n23109), .dout(n23115));
  jxor g05093(.dina(n23102), .dinb(n348), .dout(n23116));
  jand g05094(.dina(n23116), .dinb(n23115), .dout(n23117));
  jor  g05095(.dina(n23117), .dinb(n23103), .dout(n23118));
  jxor g05096(.dina(n23097), .dinb(n344), .dout(n23119));
  jand g05097(.dina(n23119), .dinb(n23118), .dout(n23120));
  jor  g05098(.dina(n23120), .dinb(n23098), .dout(n23121));
  jxor g05099(.dina(n23092), .dinb(n337), .dout(n23122));
  jand g05100(.dina(n23122), .dinb(n23121), .dout(n23123));
  jor  g05101(.dina(n23123), .dinb(n23093), .dout(n23124));
  jxor g05102(.dina(n23087), .dinb(n338), .dout(n23125));
  jand g05103(.dina(n23125), .dinb(n23124), .dout(n23126));
  jor  g05104(.dina(n23126), .dinb(n23088), .dout(n23127));
  jxor g05105(.dina(n23082), .dinb(n334), .dout(n23128));
  jand g05106(.dina(n23128), .dinb(n23127), .dout(n23129));
  jor  g05107(.dina(n23129), .dinb(n23083), .dout(n23130));
  jxor g05108(.dina(n23077), .dinb(n335), .dout(n23131));
  jand g05109(.dina(n23131), .dinb(n23130), .dout(n23132));
  jor  g05110(.dina(n23132), .dinb(n23078), .dout(n23133));
  jxor g05111(.dina(n23072), .dinb(n323), .dout(n23134));
  jand g05112(.dina(n23134), .dinb(n23133), .dout(n23135));
  jor  g05113(.dina(n23135), .dinb(n23073), .dout(n23136));
  jxor g05114(.dina(n23067), .dinb(n324), .dout(n23137));
  jand g05115(.dina(n23137), .dinb(n23136), .dout(n23138));
  jor  g05116(.dina(n23138), .dinb(n23068), .dout(n23139));
  jxor g05117(.dina(n23062), .dinb(n325), .dout(n23140));
  jand g05118(.dina(n23140), .dinb(n23139), .dout(n23141));
  jor  g05119(.dina(n23141), .dinb(n23063), .dout(n23142));
  jxor g05120(.dina(n23057), .dinb(n439), .dout(n23143));
  jand g05121(.dina(n23143), .dinb(n23142), .dout(n23144));
  jor  g05122(.dina(n23144), .dinb(n23058), .dout(n23145));
  jxor g05123(.dina(n23052), .dinb(n440), .dout(n23146));
  jand g05124(.dina(n23146), .dinb(n23145), .dout(n23147));
  jor  g05125(.dina(n23147), .dinb(n23053), .dout(n23148));
  jxor g05126(.dina(n23047), .dinb(n435), .dout(n23149));
  jand g05127(.dina(n23149), .dinb(n23148), .dout(n23150));
  jor  g05128(.dina(n23150), .dinb(n23048), .dout(n23151));
  jxor g05129(.dina(n23042), .dinb(n436), .dout(n23152));
  jand g05130(.dina(n23152), .dinb(n23151), .dout(n23153));
  jor  g05131(.dina(n23153), .dinb(n23043), .dout(n23154));
  jxor g05132(.dina(n23037), .dinb(n432), .dout(n23155));
  jand g05133(.dina(n23155), .dinb(n23154), .dout(n23156));
  jor  g05134(.dina(n23156), .dinb(n23038), .dout(n23157));
  jxor g05135(.dina(n23032), .dinb(n433), .dout(n23158));
  jand g05136(.dina(n23158), .dinb(n23157), .dout(n23159));
  jor  g05137(.dina(n23159), .dinb(n23033), .dout(n23160));
  jxor g05138(.dina(n23027), .dinb(n421), .dout(n23161));
  jand g05139(.dina(n23161), .dinb(n23160), .dout(n23162));
  jor  g05140(.dina(n23162), .dinb(n23028), .dout(n23163));
  jxor g05141(.dina(n23022), .dinb(n422), .dout(n23164));
  jand g05142(.dina(n23164), .dinb(n23163), .dout(n23165));
  jor  g05143(.dina(n23165), .dinb(n23023), .dout(n23166));
  jxor g05144(.dina(n23017), .dinb(n416), .dout(n23167));
  jand g05145(.dina(n23167), .dinb(n23166), .dout(n23168));
  jor  g05146(.dina(n23168), .dinb(n23018), .dout(n23169));
  jxor g05147(.dina(n23012), .dinb(n417), .dout(n23170));
  jand g05148(.dina(n23170), .dinb(n23169), .dout(n23171));
  jor  g05149(.dina(n23171), .dinb(n23013), .dout(n23172));
  jxor g05150(.dina(n23007), .dinb(n2547), .dout(n23173));
  jand g05151(.dina(n23173), .dinb(n23172), .dout(n23174));
  jor  g05152(.dina(n23174), .dinb(n23008), .dout(n23175));
  jxor g05153(.dina(n23002), .dinb(n2714), .dout(n23176));
  jand g05154(.dina(n23176), .dinb(n23175), .dout(n23177));
  jor  g05155(.dina(n23177), .dinb(n23003), .dout(n23178));
  jxor g05156(.dina(n22997), .dinb(n405), .dout(n23179));
  jand g05157(.dina(n23179), .dinb(n23178), .dout(n23180));
  jor  g05158(.dina(n23180), .dinb(n22998), .dout(n23181));
  jxor g05159(.dina(n22992), .dinb(n406), .dout(n23182));
  jand g05160(.dina(n23182), .dinb(n23181), .dout(n23183));
  jor  g05161(.dina(n23183), .dinb(n22993), .dout(n23184));
  jxor g05162(.dina(n22987), .dinb(n412), .dout(n23185));
  jand g05163(.dina(n23185), .dinb(n23184), .dout(n23186));
  jor  g05164(.dina(n23186), .dinb(n22988), .dout(n23187));
  jxor g05165(.dina(n22982), .dinb(n413), .dout(n23188));
  jand g05166(.dina(n23188), .dinb(n23187), .dout(n23189));
  jor  g05167(.dina(n23189), .dinb(n22983), .dout(n23190));
  jor  g05168(.dina(n23190), .dinb(n22976), .dout(n23191));
  jand g05169(.dina(n23191), .dinb(n22975), .dout(n23192));
  jand g05170(.dina(n23192), .dinb(n3401), .dout(n23193));
  jnot g05171(.din(n23193), .dout(n23194));
  jand g05172(.dina(n23194), .dinb(n22973), .dout(n23195));
  jand g05173(.dina(n22976), .dinb(n3401), .dout(n23196));
  jand g05174(.dina(n23196), .dinb(n23190), .dout(n23197));
  jor  g05175(.dina(n23197), .dinb(n23195), .dout(n23198));
  jand g05176(.dina(n23198), .dinb(n410), .dout(n23199));
  jand g05177(.dina(n23194), .dinb(n22982), .dout(n23200));
  jxor g05178(.dina(n23188), .dinb(n23187), .dout(n23201));
  jand g05179(.dina(n23201), .dinb(n23193), .dout(n23202));
  jor  g05180(.dina(n23202), .dinb(n23200), .dout(n23203));
  jand g05181(.dina(n23203), .dinb(n409), .dout(n23204));
  jand g05182(.dina(n23194), .dinb(n22987), .dout(n23205));
  jxor g05183(.dina(n23185), .dinb(n23184), .dout(n23206));
  jand g05184(.dina(n23206), .dinb(n23193), .dout(n23207));
  jor  g05185(.dina(n23207), .dinb(n23205), .dout(n23208));
  jand g05186(.dina(n23208), .dinb(n413), .dout(n23209));
  jand g05187(.dina(n23194), .dinb(n22992), .dout(n23210));
  jxor g05188(.dina(n23182), .dinb(n23181), .dout(n23211));
  jand g05189(.dina(n23211), .dinb(n23193), .dout(n23212));
  jor  g05190(.dina(n23212), .dinb(n23210), .dout(n23213));
  jand g05191(.dina(n23213), .dinb(n412), .dout(n23214));
  jand g05192(.dina(n23194), .dinb(n22997), .dout(n23215));
  jxor g05193(.dina(n23179), .dinb(n23178), .dout(n23216));
  jand g05194(.dina(n23216), .dinb(n23193), .dout(n23217));
  jor  g05195(.dina(n23217), .dinb(n23215), .dout(n23218));
  jand g05196(.dina(n23218), .dinb(n406), .dout(n23219));
  jand g05197(.dina(n23194), .dinb(n23002), .dout(n23220));
  jxor g05198(.dina(n23176), .dinb(n23175), .dout(n23221));
  jand g05199(.dina(n23221), .dinb(n23193), .dout(n23222));
  jor  g05200(.dina(n23222), .dinb(n23220), .dout(n23223));
  jand g05201(.dina(n23223), .dinb(n405), .dout(n23224));
  jand g05202(.dina(n23194), .dinb(n23007), .dout(n23225));
  jxor g05203(.dina(n23173), .dinb(n23172), .dout(n23226));
  jand g05204(.dina(n23226), .dinb(n23193), .dout(n23227));
  jor  g05205(.dina(n23227), .dinb(n23225), .dout(n23228));
  jand g05206(.dina(n23228), .dinb(n2714), .dout(n23229));
  jand g05207(.dina(n23194), .dinb(n23012), .dout(n23230));
  jxor g05208(.dina(n23170), .dinb(n23169), .dout(n23231));
  jand g05209(.dina(n23231), .dinb(n23193), .dout(n23232));
  jor  g05210(.dina(n23232), .dinb(n23230), .dout(n23233));
  jand g05211(.dina(n23233), .dinb(n2547), .dout(n23234));
  jand g05212(.dina(n23194), .dinb(n23017), .dout(n23235));
  jxor g05213(.dina(n23167), .dinb(n23166), .dout(n23236));
  jand g05214(.dina(n23236), .dinb(n23193), .dout(n23237));
  jor  g05215(.dina(n23237), .dinb(n23235), .dout(n23238));
  jand g05216(.dina(n23238), .dinb(n417), .dout(n23239));
  jand g05217(.dina(n23194), .dinb(n23022), .dout(n23240));
  jxor g05218(.dina(n23164), .dinb(n23163), .dout(n23241));
  jand g05219(.dina(n23241), .dinb(n23193), .dout(n23242));
  jor  g05220(.dina(n23242), .dinb(n23240), .dout(n23243));
  jand g05221(.dina(n23243), .dinb(n416), .dout(n23244));
  jand g05222(.dina(n23194), .dinb(n23027), .dout(n23245));
  jxor g05223(.dina(n23161), .dinb(n23160), .dout(n23246));
  jand g05224(.dina(n23246), .dinb(n23193), .dout(n23247));
  jor  g05225(.dina(n23247), .dinb(n23245), .dout(n23248));
  jand g05226(.dina(n23248), .dinb(n422), .dout(n23249));
  jand g05227(.dina(n23194), .dinb(n23032), .dout(n23250));
  jxor g05228(.dina(n23158), .dinb(n23157), .dout(n23251));
  jand g05229(.dina(n23251), .dinb(n23193), .dout(n23252));
  jor  g05230(.dina(n23252), .dinb(n23250), .dout(n23253));
  jand g05231(.dina(n23253), .dinb(n421), .dout(n23254));
  jand g05232(.dina(n23194), .dinb(n23037), .dout(n23255));
  jxor g05233(.dina(n23155), .dinb(n23154), .dout(n23256));
  jand g05234(.dina(n23256), .dinb(n23193), .dout(n23257));
  jor  g05235(.dina(n23257), .dinb(n23255), .dout(n23258));
  jand g05236(.dina(n23258), .dinb(n433), .dout(n23259));
  jand g05237(.dina(n23194), .dinb(n23042), .dout(n23260));
  jxor g05238(.dina(n23152), .dinb(n23151), .dout(n23261));
  jand g05239(.dina(n23261), .dinb(n23193), .dout(n23262));
  jor  g05240(.dina(n23262), .dinb(n23260), .dout(n23263));
  jand g05241(.dina(n23263), .dinb(n432), .dout(n23264));
  jand g05242(.dina(n23194), .dinb(n23047), .dout(n23265));
  jxor g05243(.dina(n23149), .dinb(n23148), .dout(n23266));
  jand g05244(.dina(n23266), .dinb(n23193), .dout(n23267));
  jor  g05245(.dina(n23267), .dinb(n23265), .dout(n23268));
  jand g05246(.dina(n23268), .dinb(n436), .dout(n23269));
  jand g05247(.dina(n23194), .dinb(n23052), .dout(n23270));
  jxor g05248(.dina(n23146), .dinb(n23145), .dout(n23271));
  jand g05249(.dina(n23271), .dinb(n23193), .dout(n23272));
  jor  g05250(.dina(n23272), .dinb(n23270), .dout(n23273));
  jand g05251(.dina(n23273), .dinb(n435), .dout(n23274));
  jand g05252(.dina(n23194), .dinb(n23057), .dout(n23275));
  jxor g05253(.dina(n23143), .dinb(n23142), .dout(n23276));
  jand g05254(.dina(n23276), .dinb(n23193), .dout(n23277));
  jor  g05255(.dina(n23277), .dinb(n23275), .dout(n23278));
  jand g05256(.dina(n23278), .dinb(n440), .dout(n23279));
  jand g05257(.dina(n23194), .dinb(n23062), .dout(n23280));
  jxor g05258(.dina(n23140), .dinb(n23139), .dout(n23281));
  jand g05259(.dina(n23281), .dinb(n23193), .dout(n23282));
  jor  g05260(.dina(n23282), .dinb(n23280), .dout(n23283));
  jand g05261(.dina(n23283), .dinb(n439), .dout(n23284));
  jand g05262(.dina(n23194), .dinb(n23067), .dout(n23285));
  jxor g05263(.dina(n23137), .dinb(n23136), .dout(n23286));
  jand g05264(.dina(n23286), .dinb(n23193), .dout(n23287));
  jor  g05265(.dina(n23287), .dinb(n23285), .dout(n23288));
  jand g05266(.dina(n23288), .dinb(n325), .dout(n23289));
  jand g05267(.dina(n23194), .dinb(n23072), .dout(n23290));
  jxor g05268(.dina(n23134), .dinb(n23133), .dout(n23291));
  jand g05269(.dina(n23291), .dinb(n23193), .dout(n23292));
  jor  g05270(.dina(n23292), .dinb(n23290), .dout(n23293));
  jand g05271(.dina(n23293), .dinb(n324), .dout(n23294));
  jand g05272(.dina(n23194), .dinb(n23077), .dout(n23295));
  jxor g05273(.dina(n23131), .dinb(n23130), .dout(n23296));
  jand g05274(.dina(n23296), .dinb(n23193), .dout(n23297));
  jor  g05275(.dina(n23297), .dinb(n23295), .dout(n23298));
  jand g05276(.dina(n23298), .dinb(n323), .dout(n23299));
  jand g05277(.dina(n23194), .dinb(n23082), .dout(n23300));
  jxor g05278(.dina(n23128), .dinb(n23127), .dout(n23301));
  jand g05279(.dina(n23301), .dinb(n23193), .dout(n23302));
  jor  g05280(.dina(n23302), .dinb(n23300), .dout(n23303));
  jand g05281(.dina(n23303), .dinb(n335), .dout(n23304));
  jand g05282(.dina(n23194), .dinb(n23087), .dout(n23305));
  jxor g05283(.dina(n23125), .dinb(n23124), .dout(n23306));
  jand g05284(.dina(n23306), .dinb(n23193), .dout(n23307));
  jor  g05285(.dina(n23307), .dinb(n23305), .dout(n23308));
  jand g05286(.dina(n23308), .dinb(n334), .dout(n23309));
  jand g05287(.dina(n23194), .dinb(n23092), .dout(n23310));
  jxor g05288(.dina(n23122), .dinb(n23121), .dout(n23311));
  jand g05289(.dina(n23311), .dinb(n23193), .dout(n23312));
  jor  g05290(.dina(n23312), .dinb(n23310), .dout(n23313));
  jand g05291(.dina(n23313), .dinb(n338), .dout(n23314));
  jand g05292(.dina(n23194), .dinb(n23097), .dout(n23315));
  jxor g05293(.dina(n23119), .dinb(n23118), .dout(n23316));
  jand g05294(.dina(n23316), .dinb(n23193), .dout(n23317));
  jor  g05295(.dina(n23317), .dinb(n23315), .dout(n23318));
  jand g05296(.dina(n23318), .dinb(n337), .dout(n23319));
  jnot g05297(.din(n23102), .dout(n23320));
  jor  g05298(.dina(n23193), .dinb(n23320), .dout(n23321));
  jxor g05299(.dina(n23116), .dinb(n23115), .dout(n23322));
  jnot g05300(.din(n23322), .dout(n23323));
  jor  g05301(.dina(n23323), .dinb(n23194), .dout(n23324));
  jand g05302(.dina(n23324), .dinb(n23321), .dout(n23325));
  jnot g05303(.din(n23325), .dout(n23326));
  jand g05304(.dina(n23326), .dinb(n344), .dout(n23327));
  jor  g05305(.dina(n23193), .dinb(n23112), .dout(n23328));
  jxor g05306(.dina(n23113), .dinb(n4075), .dout(n23329));
  jand g05307(.dina(n23329), .dinb(n23193), .dout(n23330));
  jnot g05308(.din(n23330), .dout(n23331));
  jand g05309(.dina(n23331), .dinb(n23328), .dout(n23332));
  jor  g05310(.dina(n23332), .dinb(b2 ), .dout(n23333));
  jnot g05311(.din(n23333), .dout(n23334));
  jnot g05312(.din(n3839), .dout(n23335));
  jnot g05313(.din(n22976), .dout(n23336));
  jnot g05314(.din(n22983), .dout(n23337));
  jnot g05315(.din(n22988), .dout(n23338));
  jnot g05316(.din(n22993), .dout(n23339));
  jnot g05317(.din(n22998), .dout(n23340));
  jnot g05318(.din(n23003), .dout(n23341));
  jnot g05319(.din(n23008), .dout(n23342));
  jnot g05320(.din(n23013), .dout(n23343));
  jnot g05321(.din(n23018), .dout(n23344));
  jnot g05322(.din(n23023), .dout(n23345));
  jnot g05323(.din(n23028), .dout(n23346));
  jnot g05324(.din(n23033), .dout(n23347));
  jnot g05325(.din(n23038), .dout(n23348));
  jnot g05326(.din(n23043), .dout(n23349));
  jnot g05327(.din(n23048), .dout(n23350));
  jnot g05328(.din(n23053), .dout(n23351));
  jnot g05329(.din(n23058), .dout(n23352));
  jnot g05330(.din(n23063), .dout(n23353));
  jnot g05331(.din(n23068), .dout(n23354));
  jnot g05332(.din(n23073), .dout(n23355));
  jnot g05333(.din(n23078), .dout(n23356));
  jnot g05334(.din(n23083), .dout(n23357));
  jnot g05335(.din(n23088), .dout(n23358));
  jnot g05336(.din(n23093), .dout(n23359));
  jnot g05337(.din(n23098), .dout(n23360));
  jnot g05338(.din(n23103), .dout(n23361));
  jnot g05339(.din(n23109), .dout(n23362));
  jxor g05340(.dina(n23112), .dinb(n258), .dout(n23363));
  jor  g05341(.dina(n23363), .dinb(n4074), .dout(n23364));
  jand g05342(.dina(n23364), .dinb(n23362), .dout(n23365));
  jnot g05343(.din(n23116), .dout(n23366));
  jor  g05344(.dina(n23366), .dinb(n23365), .dout(n23367));
  jand g05345(.dina(n23367), .dinb(n23361), .dout(n23368));
  jnot g05346(.din(n23119), .dout(n23369));
  jor  g05347(.dina(n23369), .dinb(n23368), .dout(n23370));
  jand g05348(.dina(n23370), .dinb(n23360), .dout(n23371));
  jnot g05349(.din(n23122), .dout(n23372));
  jor  g05350(.dina(n23372), .dinb(n23371), .dout(n23373));
  jand g05351(.dina(n23373), .dinb(n23359), .dout(n23374));
  jnot g05352(.din(n23125), .dout(n23375));
  jor  g05353(.dina(n23375), .dinb(n23374), .dout(n23376));
  jand g05354(.dina(n23376), .dinb(n23358), .dout(n23377));
  jnot g05355(.din(n23128), .dout(n23378));
  jor  g05356(.dina(n23378), .dinb(n23377), .dout(n23379));
  jand g05357(.dina(n23379), .dinb(n23357), .dout(n23380));
  jnot g05358(.din(n23131), .dout(n23381));
  jor  g05359(.dina(n23381), .dinb(n23380), .dout(n23382));
  jand g05360(.dina(n23382), .dinb(n23356), .dout(n23383));
  jnot g05361(.din(n23134), .dout(n23384));
  jor  g05362(.dina(n23384), .dinb(n23383), .dout(n23385));
  jand g05363(.dina(n23385), .dinb(n23355), .dout(n23386));
  jnot g05364(.din(n23137), .dout(n23387));
  jor  g05365(.dina(n23387), .dinb(n23386), .dout(n23388));
  jand g05366(.dina(n23388), .dinb(n23354), .dout(n23389));
  jnot g05367(.din(n23140), .dout(n23390));
  jor  g05368(.dina(n23390), .dinb(n23389), .dout(n23391));
  jand g05369(.dina(n23391), .dinb(n23353), .dout(n23392));
  jnot g05370(.din(n23143), .dout(n23393));
  jor  g05371(.dina(n23393), .dinb(n23392), .dout(n23394));
  jand g05372(.dina(n23394), .dinb(n23352), .dout(n23395));
  jnot g05373(.din(n23146), .dout(n23396));
  jor  g05374(.dina(n23396), .dinb(n23395), .dout(n23397));
  jand g05375(.dina(n23397), .dinb(n23351), .dout(n23398));
  jnot g05376(.din(n23149), .dout(n23399));
  jor  g05377(.dina(n23399), .dinb(n23398), .dout(n23400));
  jand g05378(.dina(n23400), .dinb(n23350), .dout(n23401));
  jnot g05379(.din(n23152), .dout(n23402));
  jor  g05380(.dina(n23402), .dinb(n23401), .dout(n23403));
  jand g05381(.dina(n23403), .dinb(n23349), .dout(n23404));
  jnot g05382(.din(n23155), .dout(n23405));
  jor  g05383(.dina(n23405), .dinb(n23404), .dout(n23406));
  jand g05384(.dina(n23406), .dinb(n23348), .dout(n23407));
  jnot g05385(.din(n23158), .dout(n23408));
  jor  g05386(.dina(n23408), .dinb(n23407), .dout(n23409));
  jand g05387(.dina(n23409), .dinb(n23347), .dout(n23410));
  jnot g05388(.din(n23161), .dout(n23411));
  jor  g05389(.dina(n23411), .dinb(n23410), .dout(n23412));
  jand g05390(.dina(n23412), .dinb(n23346), .dout(n23413));
  jnot g05391(.din(n23164), .dout(n23414));
  jor  g05392(.dina(n23414), .dinb(n23413), .dout(n23415));
  jand g05393(.dina(n23415), .dinb(n23345), .dout(n23416));
  jnot g05394(.din(n23167), .dout(n23417));
  jor  g05395(.dina(n23417), .dinb(n23416), .dout(n23418));
  jand g05396(.dina(n23418), .dinb(n23344), .dout(n23419));
  jnot g05397(.din(n23170), .dout(n23420));
  jor  g05398(.dina(n23420), .dinb(n23419), .dout(n23421));
  jand g05399(.dina(n23421), .dinb(n23343), .dout(n23422));
  jnot g05400(.din(n23173), .dout(n23423));
  jor  g05401(.dina(n23423), .dinb(n23422), .dout(n23424));
  jand g05402(.dina(n23424), .dinb(n23342), .dout(n23425));
  jnot g05403(.din(n23176), .dout(n23426));
  jor  g05404(.dina(n23426), .dinb(n23425), .dout(n23427));
  jand g05405(.dina(n23427), .dinb(n23341), .dout(n23428));
  jnot g05406(.din(n23179), .dout(n23429));
  jor  g05407(.dina(n23429), .dinb(n23428), .dout(n23430));
  jand g05408(.dina(n23430), .dinb(n23340), .dout(n23431));
  jnot g05409(.din(n23182), .dout(n23432));
  jor  g05410(.dina(n23432), .dinb(n23431), .dout(n23433));
  jand g05411(.dina(n23433), .dinb(n23339), .dout(n23434));
  jnot g05412(.din(n23185), .dout(n23435));
  jor  g05413(.dina(n23435), .dinb(n23434), .dout(n23436));
  jand g05414(.dina(n23436), .dinb(n23338), .dout(n23437));
  jnot g05415(.din(n23188), .dout(n23438));
  jor  g05416(.dina(n23438), .dinb(n23437), .dout(n23439));
  jand g05417(.dina(n23439), .dinb(n23337), .dout(n23440));
  jand g05418(.dina(n23440), .dinb(n23336), .dout(n23441));
  jor  g05419(.dina(n23441), .dinb(n22974), .dout(n23442));
  jor  g05420(.dina(n23442), .dinb(n23335), .dout(n23443));
  jand g05421(.dina(n23443), .dinb(a36 ), .dout(n23444));
  jnot g05422(.din(n4295), .dout(n23445));
  jor  g05423(.dina(n23442), .dinb(n23445), .dout(n23446));
  jnot g05424(.din(n23446), .dout(n23447));
  jor  g05425(.dina(n23447), .dinb(n23444), .dout(n23448));
  jand g05426(.dina(n23448), .dinb(n258), .dout(n23449));
  jand g05427(.dina(n23192), .dinb(n3839), .dout(n23450));
  jor  g05428(.dina(n23450), .dinb(n4073), .dout(n23451));
  jand g05429(.dina(n23446), .dinb(n23451), .dout(n23452));
  jxor g05430(.dina(n23452), .dinb(b1 ), .dout(n23453));
  jand g05431(.dina(n23453), .dinb(n4303), .dout(n23454));
  jor  g05432(.dina(n23454), .dinb(n23449), .dout(n23455));
  jxor g05433(.dina(n23332), .dinb(b2 ), .dout(n23456));
  jand g05434(.dina(n23456), .dinb(n23455), .dout(n23457));
  jor  g05435(.dina(n23457), .dinb(n23334), .dout(n23458));
  jxor g05436(.dina(n23325), .dinb(b3 ), .dout(n23459));
  jand g05437(.dina(n23459), .dinb(n23458), .dout(n23460));
  jor  g05438(.dina(n23460), .dinb(n23327), .dout(n23461));
  jxor g05439(.dina(n23318), .dinb(n337), .dout(n23462));
  jand g05440(.dina(n23462), .dinb(n23461), .dout(n23463));
  jor  g05441(.dina(n23463), .dinb(n23319), .dout(n23464));
  jxor g05442(.dina(n23313), .dinb(n338), .dout(n23465));
  jand g05443(.dina(n23465), .dinb(n23464), .dout(n23466));
  jor  g05444(.dina(n23466), .dinb(n23314), .dout(n23467));
  jxor g05445(.dina(n23308), .dinb(n334), .dout(n23468));
  jand g05446(.dina(n23468), .dinb(n23467), .dout(n23469));
  jor  g05447(.dina(n23469), .dinb(n23309), .dout(n23470));
  jxor g05448(.dina(n23303), .dinb(n335), .dout(n23471));
  jand g05449(.dina(n23471), .dinb(n23470), .dout(n23472));
  jor  g05450(.dina(n23472), .dinb(n23304), .dout(n23473));
  jxor g05451(.dina(n23298), .dinb(n323), .dout(n23474));
  jand g05452(.dina(n23474), .dinb(n23473), .dout(n23475));
  jor  g05453(.dina(n23475), .dinb(n23299), .dout(n23476));
  jxor g05454(.dina(n23293), .dinb(n324), .dout(n23477));
  jand g05455(.dina(n23477), .dinb(n23476), .dout(n23478));
  jor  g05456(.dina(n23478), .dinb(n23294), .dout(n23479));
  jxor g05457(.dina(n23288), .dinb(n325), .dout(n23480));
  jand g05458(.dina(n23480), .dinb(n23479), .dout(n23481));
  jor  g05459(.dina(n23481), .dinb(n23289), .dout(n23482));
  jxor g05460(.dina(n23283), .dinb(n439), .dout(n23483));
  jand g05461(.dina(n23483), .dinb(n23482), .dout(n23484));
  jor  g05462(.dina(n23484), .dinb(n23284), .dout(n23485));
  jxor g05463(.dina(n23278), .dinb(n440), .dout(n23486));
  jand g05464(.dina(n23486), .dinb(n23485), .dout(n23487));
  jor  g05465(.dina(n23487), .dinb(n23279), .dout(n23488));
  jxor g05466(.dina(n23273), .dinb(n435), .dout(n23489));
  jand g05467(.dina(n23489), .dinb(n23488), .dout(n23490));
  jor  g05468(.dina(n23490), .dinb(n23274), .dout(n23491));
  jxor g05469(.dina(n23268), .dinb(n436), .dout(n23492));
  jand g05470(.dina(n23492), .dinb(n23491), .dout(n23493));
  jor  g05471(.dina(n23493), .dinb(n23269), .dout(n23494));
  jxor g05472(.dina(n23263), .dinb(n432), .dout(n23495));
  jand g05473(.dina(n23495), .dinb(n23494), .dout(n23496));
  jor  g05474(.dina(n23496), .dinb(n23264), .dout(n23497));
  jxor g05475(.dina(n23258), .dinb(n433), .dout(n23498));
  jand g05476(.dina(n23498), .dinb(n23497), .dout(n23499));
  jor  g05477(.dina(n23499), .dinb(n23259), .dout(n23500));
  jxor g05478(.dina(n23253), .dinb(n421), .dout(n23501));
  jand g05479(.dina(n23501), .dinb(n23500), .dout(n23502));
  jor  g05480(.dina(n23502), .dinb(n23254), .dout(n23503));
  jxor g05481(.dina(n23248), .dinb(n422), .dout(n23504));
  jand g05482(.dina(n23504), .dinb(n23503), .dout(n23505));
  jor  g05483(.dina(n23505), .dinb(n23249), .dout(n23506));
  jxor g05484(.dina(n23243), .dinb(n416), .dout(n23507));
  jand g05485(.dina(n23507), .dinb(n23506), .dout(n23508));
  jor  g05486(.dina(n23508), .dinb(n23244), .dout(n23509));
  jxor g05487(.dina(n23238), .dinb(n417), .dout(n23510));
  jand g05488(.dina(n23510), .dinb(n23509), .dout(n23511));
  jor  g05489(.dina(n23511), .dinb(n23239), .dout(n23512));
  jxor g05490(.dina(n23233), .dinb(n2547), .dout(n23513));
  jand g05491(.dina(n23513), .dinb(n23512), .dout(n23514));
  jor  g05492(.dina(n23514), .dinb(n23234), .dout(n23515));
  jxor g05493(.dina(n23228), .dinb(n2714), .dout(n23516));
  jand g05494(.dina(n23516), .dinb(n23515), .dout(n23517));
  jor  g05495(.dina(n23517), .dinb(n23229), .dout(n23518));
  jxor g05496(.dina(n23223), .dinb(n405), .dout(n23519));
  jand g05497(.dina(n23519), .dinb(n23518), .dout(n23520));
  jor  g05498(.dina(n23520), .dinb(n23224), .dout(n23521));
  jxor g05499(.dina(n23218), .dinb(n406), .dout(n23522));
  jand g05500(.dina(n23522), .dinb(n23521), .dout(n23523));
  jor  g05501(.dina(n23523), .dinb(n23219), .dout(n23524));
  jxor g05502(.dina(n23213), .dinb(n412), .dout(n23525));
  jand g05503(.dina(n23525), .dinb(n23524), .dout(n23526));
  jor  g05504(.dina(n23526), .dinb(n23214), .dout(n23527));
  jxor g05505(.dina(n23208), .dinb(n413), .dout(n23528));
  jand g05506(.dina(n23528), .dinb(n23527), .dout(n23529));
  jor  g05507(.dina(n23529), .dinb(n23209), .dout(n23530));
  jxor g05508(.dina(n23203), .dinb(n409), .dout(n23531));
  jand g05509(.dina(n23531), .dinb(n23530), .dout(n23532));
  jor  g05510(.dina(n23532), .dinb(n23204), .dout(n23533));
  jnot g05511(.din(n23198), .dout(n23534));
  jand g05512(.dina(n23534), .dinb(b28 ), .dout(n23535));
  jnot g05513(.din(n23535), .dout(n23536));
  jand g05514(.dina(n23536), .dinb(n23533), .dout(n23537));
  jor  g05515(.dina(n23537), .dinb(n23199), .dout(n23538));
  jand g05516(.dina(n23538), .dinb(n2196), .dout(n23539));
  jnot g05517(.din(n23539), .dout(n23540));
  jand g05518(.dina(n23540), .dinb(n23198), .dout(n23541));
  jand g05519(.dina(n23199), .dinb(n2196), .dout(n23542));
  jand g05520(.dina(n23542), .dinb(n23533), .dout(n23543));
  jor  g05521(.dina(n23543), .dinb(n23541), .dout(n23544));
  jnot g05522(.din(n23544), .dout(n23545));
  jand g05523(.dina(n23540), .dinb(n23203), .dout(n23546));
  jxor g05524(.dina(n23531), .dinb(n23530), .dout(n23547));
  jand g05525(.dina(n23547), .dinb(n23539), .dout(n23548));
  jor  g05526(.dina(n23548), .dinb(n23546), .dout(n23549));
  jand g05527(.dina(n23549), .dinb(n410), .dout(n23550));
  jnot g05528(.din(n23550), .dout(n23551));
  jand g05529(.dina(n23540), .dinb(n23208), .dout(n23552));
  jxor g05530(.dina(n23528), .dinb(n23527), .dout(n23553));
  jand g05531(.dina(n23553), .dinb(n23539), .dout(n23554));
  jor  g05532(.dina(n23554), .dinb(n23552), .dout(n23555));
  jand g05533(.dina(n23555), .dinb(n409), .dout(n23556));
  jnot g05534(.din(n23556), .dout(n23557));
  jand g05535(.dina(n23540), .dinb(n23213), .dout(n23558));
  jxor g05536(.dina(n23525), .dinb(n23524), .dout(n23559));
  jand g05537(.dina(n23559), .dinb(n23539), .dout(n23560));
  jor  g05538(.dina(n23560), .dinb(n23558), .dout(n23561));
  jand g05539(.dina(n23561), .dinb(n413), .dout(n23562));
  jnot g05540(.din(n23562), .dout(n23563));
  jand g05541(.dina(n23540), .dinb(n23218), .dout(n23564));
  jxor g05542(.dina(n23522), .dinb(n23521), .dout(n23565));
  jand g05543(.dina(n23565), .dinb(n23539), .dout(n23566));
  jor  g05544(.dina(n23566), .dinb(n23564), .dout(n23567));
  jand g05545(.dina(n23567), .dinb(n412), .dout(n23568));
  jnot g05546(.din(n23568), .dout(n23569));
  jand g05547(.dina(n23540), .dinb(n23223), .dout(n23570));
  jxor g05548(.dina(n23519), .dinb(n23518), .dout(n23571));
  jand g05549(.dina(n23571), .dinb(n23539), .dout(n23572));
  jor  g05550(.dina(n23572), .dinb(n23570), .dout(n23573));
  jand g05551(.dina(n23573), .dinb(n406), .dout(n23574));
  jnot g05552(.din(n23574), .dout(n23575));
  jand g05553(.dina(n23540), .dinb(n23228), .dout(n23576));
  jxor g05554(.dina(n23516), .dinb(n23515), .dout(n23577));
  jand g05555(.dina(n23577), .dinb(n23539), .dout(n23578));
  jor  g05556(.dina(n23578), .dinb(n23576), .dout(n23579));
  jand g05557(.dina(n23579), .dinb(n405), .dout(n23580));
  jnot g05558(.din(n23580), .dout(n23581));
  jand g05559(.dina(n23540), .dinb(n23233), .dout(n23582));
  jxor g05560(.dina(n23513), .dinb(n23512), .dout(n23583));
  jand g05561(.dina(n23583), .dinb(n23539), .dout(n23584));
  jor  g05562(.dina(n23584), .dinb(n23582), .dout(n23585));
  jand g05563(.dina(n23585), .dinb(n2714), .dout(n23586));
  jnot g05564(.din(n23586), .dout(n23587));
  jand g05565(.dina(n23540), .dinb(n23238), .dout(n23588));
  jxor g05566(.dina(n23510), .dinb(n23509), .dout(n23589));
  jand g05567(.dina(n23589), .dinb(n23539), .dout(n23590));
  jor  g05568(.dina(n23590), .dinb(n23588), .dout(n23591));
  jand g05569(.dina(n23591), .dinb(n2547), .dout(n23592));
  jnot g05570(.din(n23592), .dout(n23593));
  jand g05571(.dina(n23540), .dinb(n23243), .dout(n23594));
  jxor g05572(.dina(n23507), .dinb(n23506), .dout(n23595));
  jand g05573(.dina(n23595), .dinb(n23539), .dout(n23596));
  jor  g05574(.dina(n23596), .dinb(n23594), .dout(n23597));
  jand g05575(.dina(n23597), .dinb(n417), .dout(n23598));
  jnot g05576(.din(n23598), .dout(n23599));
  jand g05577(.dina(n23540), .dinb(n23248), .dout(n23600));
  jxor g05578(.dina(n23504), .dinb(n23503), .dout(n23601));
  jand g05579(.dina(n23601), .dinb(n23539), .dout(n23602));
  jor  g05580(.dina(n23602), .dinb(n23600), .dout(n23603));
  jand g05581(.dina(n23603), .dinb(n416), .dout(n23604));
  jnot g05582(.din(n23604), .dout(n23605));
  jand g05583(.dina(n23540), .dinb(n23253), .dout(n23606));
  jxor g05584(.dina(n23501), .dinb(n23500), .dout(n23607));
  jand g05585(.dina(n23607), .dinb(n23539), .dout(n23608));
  jor  g05586(.dina(n23608), .dinb(n23606), .dout(n23609));
  jand g05587(.dina(n23609), .dinb(n422), .dout(n23610));
  jnot g05588(.din(n23610), .dout(n23611));
  jand g05589(.dina(n23540), .dinb(n23258), .dout(n23612));
  jxor g05590(.dina(n23498), .dinb(n23497), .dout(n23613));
  jand g05591(.dina(n23613), .dinb(n23539), .dout(n23614));
  jor  g05592(.dina(n23614), .dinb(n23612), .dout(n23615));
  jand g05593(.dina(n23615), .dinb(n421), .dout(n23616));
  jnot g05594(.din(n23616), .dout(n23617));
  jand g05595(.dina(n23540), .dinb(n23263), .dout(n23618));
  jxor g05596(.dina(n23495), .dinb(n23494), .dout(n23619));
  jand g05597(.dina(n23619), .dinb(n23539), .dout(n23620));
  jor  g05598(.dina(n23620), .dinb(n23618), .dout(n23621));
  jand g05599(.dina(n23621), .dinb(n433), .dout(n23622));
  jnot g05600(.din(n23622), .dout(n23623));
  jand g05601(.dina(n23540), .dinb(n23268), .dout(n23624));
  jxor g05602(.dina(n23492), .dinb(n23491), .dout(n23625));
  jand g05603(.dina(n23625), .dinb(n23539), .dout(n23626));
  jor  g05604(.dina(n23626), .dinb(n23624), .dout(n23627));
  jand g05605(.dina(n23627), .dinb(n432), .dout(n23628));
  jnot g05606(.din(n23628), .dout(n23629));
  jand g05607(.dina(n23540), .dinb(n23273), .dout(n23630));
  jxor g05608(.dina(n23489), .dinb(n23488), .dout(n23631));
  jand g05609(.dina(n23631), .dinb(n23539), .dout(n23632));
  jor  g05610(.dina(n23632), .dinb(n23630), .dout(n23633));
  jand g05611(.dina(n23633), .dinb(n436), .dout(n23634));
  jnot g05612(.din(n23634), .dout(n23635));
  jand g05613(.dina(n23540), .dinb(n23278), .dout(n23636));
  jxor g05614(.dina(n23486), .dinb(n23485), .dout(n23637));
  jand g05615(.dina(n23637), .dinb(n23539), .dout(n23638));
  jor  g05616(.dina(n23638), .dinb(n23636), .dout(n23639));
  jand g05617(.dina(n23639), .dinb(n435), .dout(n23640));
  jnot g05618(.din(n23640), .dout(n23641));
  jand g05619(.dina(n23540), .dinb(n23283), .dout(n23642));
  jxor g05620(.dina(n23483), .dinb(n23482), .dout(n23643));
  jand g05621(.dina(n23643), .dinb(n23539), .dout(n23644));
  jor  g05622(.dina(n23644), .dinb(n23642), .dout(n23645));
  jand g05623(.dina(n23645), .dinb(n440), .dout(n23646));
  jnot g05624(.din(n23646), .dout(n23647));
  jand g05625(.dina(n23540), .dinb(n23288), .dout(n23648));
  jxor g05626(.dina(n23480), .dinb(n23479), .dout(n23649));
  jand g05627(.dina(n23649), .dinb(n23539), .dout(n23650));
  jor  g05628(.dina(n23650), .dinb(n23648), .dout(n23651));
  jand g05629(.dina(n23651), .dinb(n439), .dout(n23652));
  jnot g05630(.din(n23652), .dout(n23653));
  jand g05631(.dina(n23540), .dinb(n23293), .dout(n23654));
  jxor g05632(.dina(n23477), .dinb(n23476), .dout(n23655));
  jand g05633(.dina(n23655), .dinb(n23539), .dout(n23656));
  jor  g05634(.dina(n23656), .dinb(n23654), .dout(n23657));
  jand g05635(.dina(n23657), .dinb(n325), .dout(n23658));
  jnot g05636(.din(n23658), .dout(n23659));
  jand g05637(.dina(n23540), .dinb(n23298), .dout(n23660));
  jxor g05638(.dina(n23474), .dinb(n23473), .dout(n23661));
  jand g05639(.dina(n23661), .dinb(n23539), .dout(n23662));
  jor  g05640(.dina(n23662), .dinb(n23660), .dout(n23663));
  jand g05641(.dina(n23663), .dinb(n324), .dout(n23664));
  jnot g05642(.din(n23664), .dout(n23665));
  jand g05643(.dina(n23540), .dinb(n23303), .dout(n23666));
  jxor g05644(.dina(n23471), .dinb(n23470), .dout(n23667));
  jand g05645(.dina(n23667), .dinb(n23539), .dout(n23668));
  jor  g05646(.dina(n23668), .dinb(n23666), .dout(n23669));
  jand g05647(.dina(n23669), .dinb(n323), .dout(n23670));
  jnot g05648(.din(n23670), .dout(n23671));
  jand g05649(.dina(n23540), .dinb(n23308), .dout(n23672));
  jxor g05650(.dina(n23468), .dinb(n23467), .dout(n23673));
  jand g05651(.dina(n23673), .dinb(n23539), .dout(n23674));
  jor  g05652(.dina(n23674), .dinb(n23672), .dout(n23675));
  jand g05653(.dina(n23675), .dinb(n335), .dout(n23676));
  jnot g05654(.din(n23676), .dout(n23677));
  jand g05655(.dina(n23540), .dinb(n23313), .dout(n23678));
  jxor g05656(.dina(n23465), .dinb(n23464), .dout(n23679));
  jand g05657(.dina(n23679), .dinb(n23539), .dout(n23680));
  jor  g05658(.dina(n23680), .dinb(n23678), .dout(n23681));
  jand g05659(.dina(n23681), .dinb(n334), .dout(n23682));
  jnot g05660(.din(n23682), .dout(n23683));
  jand g05661(.dina(n23540), .dinb(n23318), .dout(n23684));
  jxor g05662(.dina(n23462), .dinb(n23461), .dout(n23685));
  jand g05663(.dina(n23685), .dinb(n23539), .dout(n23686));
  jor  g05664(.dina(n23686), .dinb(n23684), .dout(n23687));
  jand g05665(.dina(n23687), .dinb(n338), .dout(n23688));
  jnot g05666(.din(n23688), .dout(n23689));
  jand g05667(.dina(n23540), .dinb(n23326), .dout(n23690));
  jxor g05668(.dina(n23459), .dinb(n23458), .dout(n23691));
  jand g05669(.dina(n23691), .dinb(n23539), .dout(n23692));
  jor  g05670(.dina(n23692), .dinb(n23690), .dout(n23693));
  jand g05671(.dina(n23693), .dinb(n337), .dout(n23694));
  jnot g05672(.din(n23694), .dout(n23695));
  jor  g05673(.dina(n23539), .dinb(n23332), .dout(n23696));
  jxor g05674(.dina(n23456), .dinb(n23455), .dout(n23697));
  jnot g05675(.din(n23697), .dout(n23698));
  jor  g05676(.dina(n23698), .dinb(n23540), .dout(n23699));
  jand g05677(.dina(n23699), .dinb(n23696), .dout(n23700));
  jnot g05678(.din(n23700), .dout(n23701));
  jand g05679(.dina(n23701), .dinb(n344), .dout(n23702));
  jnot g05680(.din(n23702), .dout(n23703));
  jor  g05681(.dina(n23539), .dinb(n23452), .dout(n23704));
  jxor g05682(.dina(n23453), .dinb(n4303), .dout(n23705));
  jand g05683(.dina(n23705), .dinb(n23539), .dout(n23706));
  jnot g05684(.din(n23706), .dout(n23707));
  jand g05685(.dina(n23707), .dinb(n23704), .dout(n23708));
  jnot g05686(.din(n23708), .dout(n23709));
  jand g05687(.dina(n23709), .dinb(n348), .dout(n23710));
  jnot g05688(.din(n23710), .dout(n23711));
  jnot g05689(.din(n4536), .dout(n23712));
  jnot g05690(.din(n23199), .dout(n23713));
  jnot g05691(.din(n23204), .dout(n23714));
  jnot g05692(.din(n23209), .dout(n23715));
  jnot g05693(.din(n23214), .dout(n23716));
  jnot g05694(.din(n23219), .dout(n23717));
  jnot g05695(.din(n23224), .dout(n23718));
  jnot g05696(.din(n23229), .dout(n23719));
  jnot g05697(.din(n23234), .dout(n23720));
  jnot g05698(.din(n23239), .dout(n23721));
  jnot g05699(.din(n23244), .dout(n23722));
  jnot g05700(.din(n23249), .dout(n23723));
  jnot g05701(.din(n23254), .dout(n23724));
  jnot g05702(.din(n23259), .dout(n23725));
  jnot g05703(.din(n23264), .dout(n23726));
  jnot g05704(.din(n23269), .dout(n23727));
  jnot g05705(.din(n23274), .dout(n23728));
  jnot g05706(.din(n23279), .dout(n23729));
  jnot g05707(.din(n23284), .dout(n23730));
  jnot g05708(.din(n23289), .dout(n23731));
  jnot g05709(.din(n23294), .dout(n23732));
  jnot g05710(.din(n23299), .dout(n23733));
  jnot g05711(.din(n23304), .dout(n23734));
  jnot g05712(.din(n23309), .dout(n23735));
  jnot g05713(.din(n23314), .dout(n23736));
  jnot g05714(.din(n23319), .dout(n23737));
  jnot g05715(.din(n23327), .dout(n23738));
  jnot g05716(.din(n23449), .dout(n23739));
  jxor g05717(.dina(n23452), .dinb(n258), .dout(n23740));
  jor  g05718(.dina(n23740), .dinb(n4302), .dout(n23741));
  jand g05719(.dina(n23741), .dinb(n23739), .dout(n23742));
  jnot g05720(.din(n23456), .dout(n23743));
  jor  g05721(.dina(n23743), .dinb(n23742), .dout(n23744));
  jand g05722(.dina(n23744), .dinb(n23333), .dout(n23745));
  jnot g05723(.din(n23459), .dout(n23746));
  jor  g05724(.dina(n23746), .dinb(n23745), .dout(n23747));
  jand g05725(.dina(n23747), .dinb(n23738), .dout(n23748));
  jnot g05726(.din(n23462), .dout(n23749));
  jor  g05727(.dina(n23749), .dinb(n23748), .dout(n23750));
  jand g05728(.dina(n23750), .dinb(n23737), .dout(n23751));
  jnot g05729(.din(n23465), .dout(n23752));
  jor  g05730(.dina(n23752), .dinb(n23751), .dout(n23753));
  jand g05731(.dina(n23753), .dinb(n23736), .dout(n23754));
  jnot g05732(.din(n23468), .dout(n23755));
  jor  g05733(.dina(n23755), .dinb(n23754), .dout(n23756));
  jand g05734(.dina(n23756), .dinb(n23735), .dout(n23757));
  jnot g05735(.din(n23471), .dout(n23758));
  jor  g05736(.dina(n23758), .dinb(n23757), .dout(n23759));
  jand g05737(.dina(n23759), .dinb(n23734), .dout(n23760));
  jnot g05738(.din(n23474), .dout(n23761));
  jor  g05739(.dina(n23761), .dinb(n23760), .dout(n23762));
  jand g05740(.dina(n23762), .dinb(n23733), .dout(n23763));
  jnot g05741(.din(n23477), .dout(n23764));
  jor  g05742(.dina(n23764), .dinb(n23763), .dout(n23765));
  jand g05743(.dina(n23765), .dinb(n23732), .dout(n23766));
  jnot g05744(.din(n23480), .dout(n23767));
  jor  g05745(.dina(n23767), .dinb(n23766), .dout(n23768));
  jand g05746(.dina(n23768), .dinb(n23731), .dout(n23769));
  jnot g05747(.din(n23483), .dout(n23770));
  jor  g05748(.dina(n23770), .dinb(n23769), .dout(n23771));
  jand g05749(.dina(n23771), .dinb(n23730), .dout(n23772));
  jnot g05750(.din(n23486), .dout(n23773));
  jor  g05751(.dina(n23773), .dinb(n23772), .dout(n23774));
  jand g05752(.dina(n23774), .dinb(n23729), .dout(n23775));
  jnot g05753(.din(n23489), .dout(n23776));
  jor  g05754(.dina(n23776), .dinb(n23775), .dout(n23777));
  jand g05755(.dina(n23777), .dinb(n23728), .dout(n23778));
  jnot g05756(.din(n23492), .dout(n23779));
  jor  g05757(.dina(n23779), .dinb(n23778), .dout(n23780));
  jand g05758(.dina(n23780), .dinb(n23727), .dout(n23781));
  jnot g05759(.din(n23495), .dout(n23782));
  jor  g05760(.dina(n23782), .dinb(n23781), .dout(n23783));
  jand g05761(.dina(n23783), .dinb(n23726), .dout(n23784));
  jnot g05762(.din(n23498), .dout(n23785));
  jor  g05763(.dina(n23785), .dinb(n23784), .dout(n23786));
  jand g05764(.dina(n23786), .dinb(n23725), .dout(n23787));
  jnot g05765(.din(n23501), .dout(n23788));
  jor  g05766(.dina(n23788), .dinb(n23787), .dout(n23789));
  jand g05767(.dina(n23789), .dinb(n23724), .dout(n23790));
  jnot g05768(.din(n23504), .dout(n23791));
  jor  g05769(.dina(n23791), .dinb(n23790), .dout(n23792));
  jand g05770(.dina(n23792), .dinb(n23723), .dout(n23793));
  jnot g05771(.din(n23507), .dout(n23794));
  jor  g05772(.dina(n23794), .dinb(n23793), .dout(n23795));
  jand g05773(.dina(n23795), .dinb(n23722), .dout(n23796));
  jnot g05774(.din(n23510), .dout(n23797));
  jor  g05775(.dina(n23797), .dinb(n23796), .dout(n23798));
  jand g05776(.dina(n23798), .dinb(n23721), .dout(n23799));
  jnot g05777(.din(n23513), .dout(n23800));
  jor  g05778(.dina(n23800), .dinb(n23799), .dout(n23801));
  jand g05779(.dina(n23801), .dinb(n23720), .dout(n23802));
  jnot g05780(.din(n23516), .dout(n23803));
  jor  g05781(.dina(n23803), .dinb(n23802), .dout(n23804));
  jand g05782(.dina(n23804), .dinb(n23719), .dout(n23805));
  jnot g05783(.din(n23519), .dout(n23806));
  jor  g05784(.dina(n23806), .dinb(n23805), .dout(n23807));
  jand g05785(.dina(n23807), .dinb(n23718), .dout(n23808));
  jnot g05786(.din(n23522), .dout(n23809));
  jor  g05787(.dina(n23809), .dinb(n23808), .dout(n23810));
  jand g05788(.dina(n23810), .dinb(n23717), .dout(n23811));
  jnot g05789(.din(n23525), .dout(n23812));
  jor  g05790(.dina(n23812), .dinb(n23811), .dout(n23813));
  jand g05791(.dina(n23813), .dinb(n23716), .dout(n23814));
  jnot g05792(.din(n23528), .dout(n23815));
  jor  g05793(.dina(n23815), .dinb(n23814), .dout(n23816));
  jand g05794(.dina(n23816), .dinb(n23715), .dout(n23817));
  jnot g05795(.din(n23531), .dout(n23818));
  jor  g05796(.dina(n23818), .dinb(n23817), .dout(n23819));
  jand g05797(.dina(n23819), .dinb(n23714), .dout(n23820));
  jor  g05798(.dina(n23535), .dinb(n23820), .dout(n23821));
  jand g05799(.dina(n23821), .dinb(n23713), .dout(n23822));
  jor  g05800(.dina(n23822), .dinb(n23712), .dout(n23823));
  jand g05801(.dina(n23823), .dinb(a35 ), .dout(n23824));
  jnot g05802(.din(n4539), .dout(n23825));
  jor  g05803(.dina(n23822), .dinb(n23825), .dout(n23826));
  jnot g05804(.din(n23826), .dout(n23827));
  jor  g05805(.dina(n23827), .dinb(n23824), .dout(n23828));
  jand g05806(.dina(n23828), .dinb(n258), .dout(n23829));
  jnot g05807(.din(n23829), .dout(n23830));
  jand g05808(.dina(n23538), .dinb(n4536), .dout(n23831));
  jor  g05809(.dina(n23831), .dinb(n4301), .dout(n23832));
  jand g05810(.dina(n23826), .dinb(n23832), .dout(n23833));
  jxor g05811(.dina(n23833), .dinb(n258), .dout(n23834));
  jor  g05812(.dina(n23834), .dinb(n4546), .dout(n23835));
  jand g05813(.dina(n23835), .dinb(n23830), .dout(n23836));
  jxor g05814(.dina(n23708), .dinb(b2 ), .dout(n23837));
  jnot g05815(.din(n23837), .dout(n23838));
  jor  g05816(.dina(n23838), .dinb(n23836), .dout(n23839));
  jand g05817(.dina(n23839), .dinb(n23711), .dout(n23840));
  jxor g05818(.dina(n23700), .dinb(b3 ), .dout(n23841));
  jnot g05819(.din(n23841), .dout(n23842));
  jor  g05820(.dina(n23842), .dinb(n23840), .dout(n23843));
  jand g05821(.dina(n23843), .dinb(n23703), .dout(n23844));
  jxor g05822(.dina(n23693), .dinb(n337), .dout(n23845));
  jnot g05823(.din(n23845), .dout(n23846));
  jor  g05824(.dina(n23846), .dinb(n23844), .dout(n23847));
  jand g05825(.dina(n23847), .dinb(n23695), .dout(n23848));
  jxor g05826(.dina(n23687), .dinb(n338), .dout(n23849));
  jnot g05827(.din(n23849), .dout(n23850));
  jor  g05828(.dina(n23850), .dinb(n23848), .dout(n23851));
  jand g05829(.dina(n23851), .dinb(n23689), .dout(n23852));
  jxor g05830(.dina(n23681), .dinb(n334), .dout(n23853));
  jnot g05831(.din(n23853), .dout(n23854));
  jor  g05832(.dina(n23854), .dinb(n23852), .dout(n23855));
  jand g05833(.dina(n23855), .dinb(n23683), .dout(n23856));
  jxor g05834(.dina(n23675), .dinb(n335), .dout(n23857));
  jnot g05835(.din(n23857), .dout(n23858));
  jor  g05836(.dina(n23858), .dinb(n23856), .dout(n23859));
  jand g05837(.dina(n23859), .dinb(n23677), .dout(n23860));
  jxor g05838(.dina(n23669), .dinb(n323), .dout(n23861));
  jnot g05839(.din(n23861), .dout(n23862));
  jor  g05840(.dina(n23862), .dinb(n23860), .dout(n23863));
  jand g05841(.dina(n23863), .dinb(n23671), .dout(n23864));
  jxor g05842(.dina(n23663), .dinb(n324), .dout(n23865));
  jnot g05843(.din(n23865), .dout(n23866));
  jor  g05844(.dina(n23866), .dinb(n23864), .dout(n23867));
  jand g05845(.dina(n23867), .dinb(n23665), .dout(n23868));
  jxor g05846(.dina(n23657), .dinb(n325), .dout(n23869));
  jnot g05847(.din(n23869), .dout(n23870));
  jor  g05848(.dina(n23870), .dinb(n23868), .dout(n23871));
  jand g05849(.dina(n23871), .dinb(n23659), .dout(n23872));
  jxor g05850(.dina(n23651), .dinb(n439), .dout(n23873));
  jnot g05851(.din(n23873), .dout(n23874));
  jor  g05852(.dina(n23874), .dinb(n23872), .dout(n23875));
  jand g05853(.dina(n23875), .dinb(n23653), .dout(n23876));
  jxor g05854(.dina(n23645), .dinb(n440), .dout(n23877));
  jnot g05855(.din(n23877), .dout(n23878));
  jor  g05856(.dina(n23878), .dinb(n23876), .dout(n23879));
  jand g05857(.dina(n23879), .dinb(n23647), .dout(n23880));
  jxor g05858(.dina(n23639), .dinb(n435), .dout(n23881));
  jnot g05859(.din(n23881), .dout(n23882));
  jor  g05860(.dina(n23882), .dinb(n23880), .dout(n23883));
  jand g05861(.dina(n23883), .dinb(n23641), .dout(n23884));
  jxor g05862(.dina(n23633), .dinb(n436), .dout(n23885));
  jnot g05863(.din(n23885), .dout(n23886));
  jor  g05864(.dina(n23886), .dinb(n23884), .dout(n23887));
  jand g05865(.dina(n23887), .dinb(n23635), .dout(n23888));
  jxor g05866(.dina(n23627), .dinb(n432), .dout(n23889));
  jnot g05867(.din(n23889), .dout(n23890));
  jor  g05868(.dina(n23890), .dinb(n23888), .dout(n23891));
  jand g05869(.dina(n23891), .dinb(n23629), .dout(n23892));
  jxor g05870(.dina(n23621), .dinb(n433), .dout(n23893));
  jnot g05871(.din(n23893), .dout(n23894));
  jor  g05872(.dina(n23894), .dinb(n23892), .dout(n23895));
  jand g05873(.dina(n23895), .dinb(n23623), .dout(n23896));
  jxor g05874(.dina(n23615), .dinb(n421), .dout(n23897));
  jnot g05875(.din(n23897), .dout(n23898));
  jor  g05876(.dina(n23898), .dinb(n23896), .dout(n23899));
  jand g05877(.dina(n23899), .dinb(n23617), .dout(n23900));
  jxor g05878(.dina(n23609), .dinb(n422), .dout(n23901));
  jnot g05879(.din(n23901), .dout(n23902));
  jor  g05880(.dina(n23902), .dinb(n23900), .dout(n23903));
  jand g05881(.dina(n23903), .dinb(n23611), .dout(n23904));
  jxor g05882(.dina(n23603), .dinb(n416), .dout(n23905));
  jnot g05883(.din(n23905), .dout(n23906));
  jor  g05884(.dina(n23906), .dinb(n23904), .dout(n23907));
  jand g05885(.dina(n23907), .dinb(n23605), .dout(n23908));
  jxor g05886(.dina(n23597), .dinb(n417), .dout(n23909));
  jnot g05887(.din(n23909), .dout(n23910));
  jor  g05888(.dina(n23910), .dinb(n23908), .dout(n23911));
  jand g05889(.dina(n23911), .dinb(n23599), .dout(n23912));
  jxor g05890(.dina(n23591), .dinb(n2547), .dout(n23913));
  jnot g05891(.din(n23913), .dout(n23914));
  jor  g05892(.dina(n23914), .dinb(n23912), .dout(n23915));
  jand g05893(.dina(n23915), .dinb(n23593), .dout(n23916));
  jxor g05894(.dina(n23585), .dinb(n2714), .dout(n23917));
  jnot g05895(.din(n23917), .dout(n23918));
  jor  g05896(.dina(n23918), .dinb(n23916), .dout(n23919));
  jand g05897(.dina(n23919), .dinb(n23587), .dout(n23920));
  jxor g05898(.dina(n23579), .dinb(n405), .dout(n23921));
  jnot g05899(.din(n23921), .dout(n23922));
  jor  g05900(.dina(n23922), .dinb(n23920), .dout(n23923));
  jand g05901(.dina(n23923), .dinb(n23581), .dout(n23924));
  jxor g05902(.dina(n23573), .dinb(n406), .dout(n23925));
  jnot g05903(.din(n23925), .dout(n23926));
  jor  g05904(.dina(n23926), .dinb(n23924), .dout(n23927));
  jand g05905(.dina(n23927), .dinb(n23575), .dout(n23928));
  jxor g05906(.dina(n23567), .dinb(n412), .dout(n23929));
  jnot g05907(.din(n23929), .dout(n23930));
  jor  g05908(.dina(n23930), .dinb(n23928), .dout(n23931));
  jand g05909(.dina(n23931), .dinb(n23569), .dout(n23932));
  jxor g05910(.dina(n23561), .dinb(n413), .dout(n23933));
  jnot g05911(.din(n23933), .dout(n23934));
  jor  g05912(.dina(n23934), .dinb(n23932), .dout(n23935));
  jand g05913(.dina(n23935), .dinb(n23563), .dout(n23936));
  jxor g05914(.dina(n23555), .dinb(n409), .dout(n23937));
  jnot g05915(.din(n23937), .dout(n23938));
  jor  g05916(.dina(n23938), .dinb(n23936), .dout(n23939));
  jand g05917(.dina(n23939), .dinb(n23557), .dout(n23940));
  jxor g05918(.dina(n23549), .dinb(n410), .dout(n23941));
  jnot g05919(.din(n23941), .dout(n23942));
  jor  g05920(.dina(n23942), .dinb(n23940), .dout(n23943));
  jand g05921(.dina(n23943), .dinb(n23551), .dout(n23944));
  jxor g05922(.dina(n23544), .dinb(b29 ), .dout(n23945));
  jor  g05923(.dina(n23945), .dinb(n2715), .dout(n23946));
  jor  g05924(.dina(n23946), .dinb(n23944), .dout(n23947));
  jand g05925(.dina(n23947), .dinb(n23545), .dout(n23948));
  jxor g05926(.dina(n23833), .dinb(b1 ), .dout(n23949));
  jand g05927(.dina(n23949), .dinb(n4547), .dout(n23950));
  jor  g05928(.dina(n23950), .dinb(n23829), .dout(n23951));
  jand g05929(.dina(n23837), .dinb(n23951), .dout(n23952));
  jor  g05930(.dina(n23952), .dinb(n23710), .dout(n23953));
  jand g05931(.dina(n23841), .dinb(n23953), .dout(n23954));
  jor  g05932(.dina(n23954), .dinb(n23702), .dout(n23955));
  jand g05933(.dina(n23845), .dinb(n23955), .dout(n23956));
  jor  g05934(.dina(n23956), .dinb(n23694), .dout(n23957));
  jand g05935(.dina(n23849), .dinb(n23957), .dout(n23958));
  jor  g05936(.dina(n23958), .dinb(n23688), .dout(n23959));
  jand g05937(.dina(n23853), .dinb(n23959), .dout(n23960));
  jor  g05938(.dina(n23960), .dinb(n23682), .dout(n23961));
  jand g05939(.dina(n23857), .dinb(n23961), .dout(n23962));
  jor  g05940(.dina(n23962), .dinb(n23676), .dout(n23963));
  jand g05941(.dina(n23861), .dinb(n23963), .dout(n23964));
  jor  g05942(.dina(n23964), .dinb(n23670), .dout(n23965));
  jand g05943(.dina(n23865), .dinb(n23965), .dout(n23966));
  jor  g05944(.dina(n23966), .dinb(n23664), .dout(n23967));
  jand g05945(.dina(n23869), .dinb(n23967), .dout(n23968));
  jor  g05946(.dina(n23968), .dinb(n23658), .dout(n23969));
  jand g05947(.dina(n23873), .dinb(n23969), .dout(n23970));
  jor  g05948(.dina(n23970), .dinb(n23652), .dout(n23971));
  jand g05949(.dina(n23877), .dinb(n23971), .dout(n23972));
  jor  g05950(.dina(n23972), .dinb(n23646), .dout(n23973));
  jand g05951(.dina(n23881), .dinb(n23973), .dout(n23974));
  jor  g05952(.dina(n23974), .dinb(n23640), .dout(n23975));
  jand g05953(.dina(n23885), .dinb(n23975), .dout(n23976));
  jor  g05954(.dina(n23976), .dinb(n23634), .dout(n23977));
  jand g05955(.dina(n23889), .dinb(n23977), .dout(n23978));
  jor  g05956(.dina(n23978), .dinb(n23628), .dout(n23979));
  jand g05957(.dina(n23893), .dinb(n23979), .dout(n23980));
  jor  g05958(.dina(n23980), .dinb(n23622), .dout(n23981));
  jand g05959(.dina(n23897), .dinb(n23981), .dout(n23982));
  jor  g05960(.dina(n23982), .dinb(n23616), .dout(n23983));
  jand g05961(.dina(n23901), .dinb(n23983), .dout(n23984));
  jor  g05962(.dina(n23984), .dinb(n23610), .dout(n23985));
  jand g05963(.dina(n23905), .dinb(n23985), .dout(n23986));
  jor  g05964(.dina(n23986), .dinb(n23604), .dout(n23987));
  jand g05965(.dina(n23909), .dinb(n23987), .dout(n23988));
  jor  g05966(.dina(n23988), .dinb(n23598), .dout(n23989));
  jand g05967(.dina(n23913), .dinb(n23989), .dout(n23990));
  jor  g05968(.dina(n23990), .dinb(n23592), .dout(n23991));
  jand g05969(.dina(n23917), .dinb(n23991), .dout(n23992));
  jor  g05970(.dina(n23992), .dinb(n23586), .dout(n23993));
  jand g05971(.dina(n23921), .dinb(n23993), .dout(n23994));
  jor  g05972(.dina(n23994), .dinb(n23580), .dout(n23995));
  jand g05973(.dina(n23925), .dinb(n23995), .dout(n23996));
  jor  g05974(.dina(n23996), .dinb(n23574), .dout(n23997));
  jand g05975(.dina(n23929), .dinb(n23997), .dout(n23998));
  jor  g05976(.dina(n23998), .dinb(n23568), .dout(n23999));
  jand g05977(.dina(n23933), .dinb(n23999), .dout(n24000));
  jor  g05978(.dina(n24000), .dinb(n23562), .dout(n24001));
  jand g05979(.dina(n23937), .dinb(n24001), .dout(n24002));
  jor  g05980(.dina(n24002), .dinb(n23556), .dout(n24003));
  jand g05981(.dina(n23941), .dinb(n24003), .dout(n24004));
  jor  g05982(.dina(n24004), .dinb(n23550), .dout(n24005));
  jnot g05983(.din(n23946), .dout(n24006));
  jand g05984(.dina(n24006), .dinb(n24005), .dout(n24007));
  jand g05985(.dina(n23544), .dinb(n2196), .dout(n24008));
  jor  g05986(.dina(n24008), .dinb(n24007), .dout(n24009));
  jxor g05987(.dina(n23945), .dinb(n24005), .dout(n24010));
  jand g05988(.dina(n24010), .dinb(n24009), .dout(n24011));
  jor  g05989(.dina(n24011), .dinb(n23948), .dout(n24012));
  jnot g05990(.din(n24012), .dout(n24013));
  jand g05991(.dina(n24012), .dinb(b30 ), .dout(n24014));
  jnot g05992(.din(n24014), .dout(n24015));
  jand g05993(.dina(n24013), .dinb(n427), .dout(n24016));
  jnot g05994(.din(n24008), .dout(n24017));
  jand g05995(.dina(n24017), .dinb(n23947), .dout(n24018));
  jand g05996(.dina(n24018), .dinb(n23549), .dout(n24019));
  jxor g05997(.dina(n23941), .dinb(n24003), .dout(n24020));
  jand g05998(.dina(n24020), .dinb(n24009), .dout(n24021));
  jor  g05999(.dina(n24021), .dinb(n24019), .dout(n24022));
  jand g06000(.dina(n24022), .dinb(n426), .dout(n24023));
  jand g06001(.dina(n24018), .dinb(n23555), .dout(n24024));
  jxor g06002(.dina(n23937), .dinb(n24001), .dout(n24025));
  jand g06003(.dina(n24025), .dinb(n24009), .dout(n24026));
  jor  g06004(.dina(n24026), .dinb(n24024), .dout(n24027));
  jand g06005(.dina(n24027), .dinb(n410), .dout(n24028));
  jand g06006(.dina(n24018), .dinb(n23561), .dout(n24029));
  jxor g06007(.dina(n23933), .dinb(n23999), .dout(n24030));
  jand g06008(.dina(n24030), .dinb(n24009), .dout(n24031));
  jor  g06009(.dina(n24031), .dinb(n24029), .dout(n24032));
  jand g06010(.dina(n24032), .dinb(n409), .dout(n24033));
  jand g06011(.dina(n24018), .dinb(n23567), .dout(n24034));
  jxor g06012(.dina(n23929), .dinb(n23997), .dout(n24035));
  jand g06013(.dina(n24035), .dinb(n24009), .dout(n24036));
  jor  g06014(.dina(n24036), .dinb(n24034), .dout(n24037));
  jand g06015(.dina(n24037), .dinb(n413), .dout(n24038));
  jand g06016(.dina(n24018), .dinb(n23573), .dout(n24039));
  jxor g06017(.dina(n23925), .dinb(n23995), .dout(n24040));
  jand g06018(.dina(n24040), .dinb(n24009), .dout(n24041));
  jor  g06019(.dina(n24041), .dinb(n24039), .dout(n24042));
  jand g06020(.dina(n24042), .dinb(n412), .dout(n24043));
  jand g06021(.dina(n24018), .dinb(n23579), .dout(n24044));
  jxor g06022(.dina(n23921), .dinb(n23993), .dout(n24045));
  jand g06023(.dina(n24045), .dinb(n24009), .dout(n24046));
  jor  g06024(.dina(n24046), .dinb(n24044), .dout(n24047));
  jand g06025(.dina(n24047), .dinb(n406), .dout(n24048));
  jand g06026(.dina(n24018), .dinb(n23585), .dout(n24049));
  jxor g06027(.dina(n23917), .dinb(n23991), .dout(n24050));
  jand g06028(.dina(n24050), .dinb(n24009), .dout(n24051));
  jor  g06029(.dina(n24051), .dinb(n24049), .dout(n24052));
  jand g06030(.dina(n24052), .dinb(n405), .dout(n24053));
  jand g06031(.dina(n24018), .dinb(n23591), .dout(n24054));
  jxor g06032(.dina(n23913), .dinb(n23989), .dout(n24055));
  jand g06033(.dina(n24055), .dinb(n24009), .dout(n24056));
  jor  g06034(.dina(n24056), .dinb(n24054), .dout(n24057));
  jand g06035(.dina(n24057), .dinb(n2714), .dout(n24058));
  jand g06036(.dina(n24018), .dinb(n23597), .dout(n24059));
  jxor g06037(.dina(n23909), .dinb(n23987), .dout(n24060));
  jand g06038(.dina(n24060), .dinb(n24009), .dout(n24061));
  jor  g06039(.dina(n24061), .dinb(n24059), .dout(n24062));
  jand g06040(.dina(n24062), .dinb(n2547), .dout(n24063));
  jand g06041(.dina(n24018), .dinb(n23603), .dout(n24064));
  jxor g06042(.dina(n23905), .dinb(n23985), .dout(n24065));
  jand g06043(.dina(n24065), .dinb(n24009), .dout(n24066));
  jor  g06044(.dina(n24066), .dinb(n24064), .dout(n24067));
  jand g06045(.dina(n24067), .dinb(n417), .dout(n24068));
  jand g06046(.dina(n24018), .dinb(n23609), .dout(n24069));
  jxor g06047(.dina(n23901), .dinb(n23983), .dout(n24070));
  jand g06048(.dina(n24070), .dinb(n24009), .dout(n24071));
  jor  g06049(.dina(n24071), .dinb(n24069), .dout(n24072));
  jand g06050(.dina(n24072), .dinb(n416), .dout(n24073));
  jand g06051(.dina(n24018), .dinb(n23615), .dout(n24074));
  jxor g06052(.dina(n23897), .dinb(n23981), .dout(n24075));
  jand g06053(.dina(n24075), .dinb(n24009), .dout(n24076));
  jor  g06054(.dina(n24076), .dinb(n24074), .dout(n24077));
  jand g06055(.dina(n24077), .dinb(n422), .dout(n24078));
  jand g06056(.dina(n24018), .dinb(n23621), .dout(n24079));
  jxor g06057(.dina(n23893), .dinb(n23979), .dout(n24080));
  jand g06058(.dina(n24080), .dinb(n24009), .dout(n24081));
  jor  g06059(.dina(n24081), .dinb(n24079), .dout(n24082));
  jand g06060(.dina(n24082), .dinb(n421), .dout(n24083));
  jand g06061(.dina(n24018), .dinb(n23627), .dout(n24084));
  jxor g06062(.dina(n23889), .dinb(n23977), .dout(n24085));
  jand g06063(.dina(n24085), .dinb(n24009), .dout(n24086));
  jor  g06064(.dina(n24086), .dinb(n24084), .dout(n24087));
  jand g06065(.dina(n24087), .dinb(n433), .dout(n24088));
  jand g06066(.dina(n24018), .dinb(n23633), .dout(n24089));
  jxor g06067(.dina(n23885), .dinb(n23975), .dout(n24090));
  jand g06068(.dina(n24090), .dinb(n24009), .dout(n24091));
  jor  g06069(.dina(n24091), .dinb(n24089), .dout(n24092));
  jand g06070(.dina(n24092), .dinb(n432), .dout(n24093));
  jand g06071(.dina(n24018), .dinb(n23639), .dout(n24094));
  jxor g06072(.dina(n23881), .dinb(n23973), .dout(n24095));
  jand g06073(.dina(n24095), .dinb(n24009), .dout(n24096));
  jor  g06074(.dina(n24096), .dinb(n24094), .dout(n24097));
  jand g06075(.dina(n24097), .dinb(n436), .dout(n24098));
  jand g06076(.dina(n24018), .dinb(n23645), .dout(n24099));
  jxor g06077(.dina(n23877), .dinb(n23971), .dout(n24100));
  jand g06078(.dina(n24100), .dinb(n24009), .dout(n24101));
  jor  g06079(.dina(n24101), .dinb(n24099), .dout(n24102));
  jand g06080(.dina(n24102), .dinb(n435), .dout(n24103));
  jand g06081(.dina(n24018), .dinb(n23651), .dout(n24104));
  jxor g06082(.dina(n23873), .dinb(n23969), .dout(n24105));
  jand g06083(.dina(n24105), .dinb(n24009), .dout(n24106));
  jor  g06084(.dina(n24106), .dinb(n24104), .dout(n24107));
  jand g06085(.dina(n24107), .dinb(n440), .dout(n24108));
  jand g06086(.dina(n24018), .dinb(n23657), .dout(n24109));
  jxor g06087(.dina(n23869), .dinb(n23967), .dout(n24110));
  jand g06088(.dina(n24110), .dinb(n24009), .dout(n24111));
  jor  g06089(.dina(n24111), .dinb(n24109), .dout(n24112));
  jand g06090(.dina(n24112), .dinb(n439), .dout(n24113));
  jand g06091(.dina(n24018), .dinb(n23663), .dout(n24114));
  jxor g06092(.dina(n23865), .dinb(n23965), .dout(n24115));
  jand g06093(.dina(n24115), .dinb(n24009), .dout(n24116));
  jor  g06094(.dina(n24116), .dinb(n24114), .dout(n24117));
  jand g06095(.dina(n24117), .dinb(n325), .dout(n24118));
  jand g06096(.dina(n24018), .dinb(n23669), .dout(n24119));
  jxor g06097(.dina(n23861), .dinb(n23963), .dout(n24120));
  jand g06098(.dina(n24120), .dinb(n24009), .dout(n24121));
  jor  g06099(.dina(n24121), .dinb(n24119), .dout(n24122));
  jand g06100(.dina(n24122), .dinb(n324), .dout(n24123));
  jand g06101(.dina(n24018), .dinb(n23675), .dout(n24124));
  jxor g06102(.dina(n23857), .dinb(n23961), .dout(n24125));
  jand g06103(.dina(n24125), .dinb(n24009), .dout(n24126));
  jor  g06104(.dina(n24126), .dinb(n24124), .dout(n24127));
  jand g06105(.dina(n24127), .dinb(n323), .dout(n24128));
  jand g06106(.dina(n24018), .dinb(n23681), .dout(n24129));
  jxor g06107(.dina(n23853), .dinb(n23959), .dout(n24130));
  jand g06108(.dina(n24130), .dinb(n24009), .dout(n24131));
  jor  g06109(.dina(n24131), .dinb(n24129), .dout(n24132));
  jand g06110(.dina(n24132), .dinb(n335), .dout(n24133));
  jand g06111(.dina(n24018), .dinb(n23687), .dout(n24134));
  jxor g06112(.dina(n23849), .dinb(n23957), .dout(n24135));
  jand g06113(.dina(n24135), .dinb(n24009), .dout(n24136));
  jor  g06114(.dina(n24136), .dinb(n24134), .dout(n24137));
  jand g06115(.dina(n24137), .dinb(n334), .dout(n24138));
  jand g06116(.dina(n24018), .dinb(n23693), .dout(n24139));
  jxor g06117(.dina(n23845), .dinb(n23955), .dout(n24140));
  jand g06118(.dina(n24140), .dinb(n24009), .dout(n24141));
  jor  g06119(.dina(n24141), .dinb(n24139), .dout(n24142));
  jand g06120(.dina(n24142), .dinb(n338), .dout(n24143));
  jand g06121(.dina(n24018), .dinb(n23701), .dout(n24144));
  jxor g06122(.dina(n23841), .dinb(n23953), .dout(n24145));
  jand g06123(.dina(n24145), .dinb(n24009), .dout(n24146));
  jor  g06124(.dina(n24146), .dinb(n24144), .dout(n24147));
  jand g06125(.dina(n24147), .dinb(n337), .dout(n24148));
  jand g06126(.dina(n24018), .dinb(n23709), .dout(n24149));
  jxor g06127(.dina(n23837), .dinb(n23951), .dout(n24150));
  jand g06128(.dina(n24150), .dinb(n24009), .dout(n24151));
  jor  g06129(.dina(n24151), .dinb(n24149), .dout(n24152));
  jand g06130(.dina(n24152), .dinb(n344), .dout(n24153));
  jand g06131(.dina(n24018), .dinb(n23828), .dout(n24154));
  jxor g06132(.dina(n23949), .dinb(n4547), .dout(n24155));
  jand g06133(.dina(n24155), .dinb(n24009), .dout(n24156));
  jor  g06134(.dina(n24156), .dinb(n24154), .dout(n24157));
  jand g06135(.dina(n24157), .dinb(n348), .dout(n24158));
  jor  g06136(.dina(n24018), .dinb(n18364), .dout(n24159));
  jand g06137(.dina(n24159), .dinb(a34 ), .dout(n24160));
  jor  g06138(.dina(n24018), .dinb(n4547), .dout(n24161));
  jnot g06139(.din(n24161), .dout(n24162));
  jor  g06140(.dina(n24162), .dinb(n24160), .dout(n24163));
  jand g06141(.dina(n24163), .dinb(n258), .dout(n24164));
  jand g06142(.dina(n24009), .dinb(b0 ), .dout(n24165));
  jor  g06143(.dina(n24165), .dinb(n4545), .dout(n24166));
  jand g06144(.dina(n24161), .dinb(n24166), .dout(n24167));
  jxor g06145(.dina(n24167), .dinb(b1 ), .dout(n24168));
  jand g06146(.dina(n24168), .dinb(n4800), .dout(n24169));
  jor  g06147(.dina(n24169), .dinb(n24164), .dout(n24170));
  jxor g06148(.dina(n24157), .dinb(n348), .dout(n24171));
  jand g06149(.dina(n24171), .dinb(n24170), .dout(n24172));
  jor  g06150(.dina(n24172), .dinb(n24158), .dout(n24173));
  jxor g06151(.dina(n24152), .dinb(n344), .dout(n24174));
  jand g06152(.dina(n24174), .dinb(n24173), .dout(n24175));
  jor  g06153(.dina(n24175), .dinb(n24153), .dout(n24176));
  jxor g06154(.dina(n24147), .dinb(n337), .dout(n24177));
  jand g06155(.dina(n24177), .dinb(n24176), .dout(n24178));
  jor  g06156(.dina(n24178), .dinb(n24148), .dout(n24179));
  jxor g06157(.dina(n24142), .dinb(n338), .dout(n24180));
  jand g06158(.dina(n24180), .dinb(n24179), .dout(n24181));
  jor  g06159(.dina(n24181), .dinb(n24143), .dout(n24182));
  jxor g06160(.dina(n24137), .dinb(n334), .dout(n24183));
  jand g06161(.dina(n24183), .dinb(n24182), .dout(n24184));
  jor  g06162(.dina(n24184), .dinb(n24138), .dout(n24185));
  jxor g06163(.dina(n24132), .dinb(n335), .dout(n24186));
  jand g06164(.dina(n24186), .dinb(n24185), .dout(n24187));
  jor  g06165(.dina(n24187), .dinb(n24133), .dout(n24188));
  jxor g06166(.dina(n24127), .dinb(n323), .dout(n24189));
  jand g06167(.dina(n24189), .dinb(n24188), .dout(n24190));
  jor  g06168(.dina(n24190), .dinb(n24128), .dout(n24191));
  jxor g06169(.dina(n24122), .dinb(n324), .dout(n24192));
  jand g06170(.dina(n24192), .dinb(n24191), .dout(n24193));
  jor  g06171(.dina(n24193), .dinb(n24123), .dout(n24194));
  jxor g06172(.dina(n24117), .dinb(n325), .dout(n24195));
  jand g06173(.dina(n24195), .dinb(n24194), .dout(n24196));
  jor  g06174(.dina(n24196), .dinb(n24118), .dout(n24197));
  jxor g06175(.dina(n24112), .dinb(n439), .dout(n24198));
  jand g06176(.dina(n24198), .dinb(n24197), .dout(n24199));
  jor  g06177(.dina(n24199), .dinb(n24113), .dout(n24200));
  jxor g06178(.dina(n24107), .dinb(n440), .dout(n24201));
  jand g06179(.dina(n24201), .dinb(n24200), .dout(n24202));
  jor  g06180(.dina(n24202), .dinb(n24108), .dout(n24203));
  jxor g06181(.dina(n24102), .dinb(n435), .dout(n24204));
  jand g06182(.dina(n24204), .dinb(n24203), .dout(n24205));
  jor  g06183(.dina(n24205), .dinb(n24103), .dout(n24206));
  jxor g06184(.dina(n24097), .dinb(n436), .dout(n24207));
  jand g06185(.dina(n24207), .dinb(n24206), .dout(n24208));
  jor  g06186(.dina(n24208), .dinb(n24098), .dout(n24209));
  jxor g06187(.dina(n24092), .dinb(n432), .dout(n24210));
  jand g06188(.dina(n24210), .dinb(n24209), .dout(n24211));
  jor  g06189(.dina(n24211), .dinb(n24093), .dout(n24212));
  jxor g06190(.dina(n24087), .dinb(n433), .dout(n24213));
  jand g06191(.dina(n24213), .dinb(n24212), .dout(n24214));
  jor  g06192(.dina(n24214), .dinb(n24088), .dout(n24215));
  jxor g06193(.dina(n24082), .dinb(n421), .dout(n24216));
  jand g06194(.dina(n24216), .dinb(n24215), .dout(n24217));
  jor  g06195(.dina(n24217), .dinb(n24083), .dout(n24218));
  jxor g06196(.dina(n24077), .dinb(n422), .dout(n24219));
  jand g06197(.dina(n24219), .dinb(n24218), .dout(n24220));
  jor  g06198(.dina(n24220), .dinb(n24078), .dout(n24221));
  jxor g06199(.dina(n24072), .dinb(n416), .dout(n24222));
  jand g06200(.dina(n24222), .dinb(n24221), .dout(n24223));
  jor  g06201(.dina(n24223), .dinb(n24073), .dout(n24224));
  jxor g06202(.dina(n24067), .dinb(n417), .dout(n24225));
  jand g06203(.dina(n24225), .dinb(n24224), .dout(n24226));
  jor  g06204(.dina(n24226), .dinb(n24068), .dout(n24227));
  jxor g06205(.dina(n24062), .dinb(n2547), .dout(n24228));
  jand g06206(.dina(n24228), .dinb(n24227), .dout(n24229));
  jor  g06207(.dina(n24229), .dinb(n24063), .dout(n24230));
  jxor g06208(.dina(n24057), .dinb(n2714), .dout(n24231));
  jand g06209(.dina(n24231), .dinb(n24230), .dout(n24232));
  jor  g06210(.dina(n24232), .dinb(n24058), .dout(n24233));
  jxor g06211(.dina(n24052), .dinb(n405), .dout(n24234));
  jand g06212(.dina(n24234), .dinb(n24233), .dout(n24235));
  jor  g06213(.dina(n24235), .dinb(n24053), .dout(n24236));
  jxor g06214(.dina(n24047), .dinb(n406), .dout(n24237));
  jand g06215(.dina(n24237), .dinb(n24236), .dout(n24238));
  jor  g06216(.dina(n24238), .dinb(n24048), .dout(n24239));
  jxor g06217(.dina(n24042), .dinb(n412), .dout(n24240));
  jand g06218(.dina(n24240), .dinb(n24239), .dout(n24241));
  jor  g06219(.dina(n24241), .dinb(n24043), .dout(n24242));
  jxor g06220(.dina(n24037), .dinb(n413), .dout(n24243));
  jand g06221(.dina(n24243), .dinb(n24242), .dout(n24244));
  jor  g06222(.dina(n24244), .dinb(n24038), .dout(n24245));
  jxor g06223(.dina(n24032), .dinb(n409), .dout(n24246));
  jand g06224(.dina(n24246), .dinb(n24245), .dout(n24247));
  jor  g06225(.dina(n24247), .dinb(n24033), .dout(n24248));
  jxor g06226(.dina(n24027), .dinb(n410), .dout(n24249));
  jand g06227(.dina(n24249), .dinb(n24248), .dout(n24250));
  jor  g06228(.dina(n24250), .dinb(n24028), .dout(n24251));
  jxor g06229(.dina(n24022), .dinb(n426), .dout(n24252));
  jand g06230(.dina(n24252), .dinb(n24251), .dout(n24253));
  jor  g06231(.dina(n24253), .dinb(n24023), .dout(n24254));
  jor  g06232(.dina(n24254), .dinb(n24016), .dout(n24255));
  jand g06233(.dina(n24255), .dinb(n24015), .dout(n24256));
  jand g06234(.dina(n24256), .dinb(n4642), .dout(n24257));
  jnot g06235(.din(n24257), .dout(n24258));
  jand g06236(.dina(n24258), .dinb(n24013), .dout(n24259));
  jand g06237(.dina(n24016), .dinb(n4642), .dout(n24260));
  jand g06238(.dina(n24260), .dinb(n24254), .dout(n24261));
  jor  g06239(.dina(n24261), .dinb(n24259), .dout(n24262));
  jand g06240(.dina(n24262), .dinb(n424), .dout(n24263));
  jand g06241(.dina(n24258), .dinb(n24022), .dout(n24264));
  jxor g06242(.dina(n24252), .dinb(n24251), .dout(n24265));
  jand g06243(.dina(n24265), .dinb(n24257), .dout(n24266));
  jor  g06244(.dina(n24266), .dinb(n24264), .dout(n24267));
  jand g06245(.dina(n24267), .dinb(n427), .dout(n24268));
  jand g06246(.dina(n24258), .dinb(n24027), .dout(n24269));
  jxor g06247(.dina(n24249), .dinb(n24248), .dout(n24270));
  jand g06248(.dina(n24270), .dinb(n24257), .dout(n24271));
  jor  g06249(.dina(n24271), .dinb(n24269), .dout(n24272));
  jand g06250(.dina(n24272), .dinb(n426), .dout(n24273));
  jand g06251(.dina(n24258), .dinb(n24032), .dout(n24274));
  jxor g06252(.dina(n24246), .dinb(n24245), .dout(n24275));
  jand g06253(.dina(n24275), .dinb(n24257), .dout(n24276));
  jor  g06254(.dina(n24276), .dinb(n24274), .dout(n24277));
  jand g06255(.dina(n24277), .dinb(n410), .dout(n24278));
  jand g06256(.dina(n24258), .dinb(n24037), .dout(n24279));
  jxor g06257(.dina(n24243), .dinb(n24242), .dout(n24280));
  jand g06258(.dina(n24280), .dinb(n24257), .dout(n24281));
  jor  g06259(.dina(n24281), .dinb(n24279), .dout(n24282));
  jand g06260(.dina(n24282), .dinb(n409), .dout(n24283));
  jand g06261(.dina(n24258), .dinb(n24042), .dout(n24284));
  jxor g06262(.dina(n24240), .dinb(n24239), .dout(n24285));
  jand g06263(.dina(n24285), .dinb(n24257), .dout(n24286));
  jor  g06264(.dina(n24286), .dinb(n24284), .dout(n24287));
  jand g06265(.dina(n24287), .dinb(n413), .dout(n24288));
  jand g06266(.dina(n24258), .dinb(n24047), .dout(n24289));
  jxor g06267(.dina(n24237), .dinb(n24236), .dout(n24290));
  jand g06268(.dina(n24290), .dinb(n24257), .dout(n24291));
  jor  g06269(.dina(n24291), .dinb(n24289), .dout(n24292));
  jand g06270(.dina(n24292), .dinb(n412), .dout(n24293));
  jand g06271(.dina(n24258), .dinb(n24052), .dout(n24294));
  jxor g06272(.dina(n24234), .dinb(n24233), .dout(n24295));
  jand g06273(.dina(n24295), .dinb(n24257), .dout(n24296));
  jor  g06274(.dina(n24296), .dinb(n24294), .dout(n24297));
  jand g06275(.dina(n24297), .dinb(n406), .dout(n24298));
  jand g06276(.dina(n24258), .dinb(n24057), .dout(n24299));
  jxor g06277(.dina(n24231), .dinb(n24230), .dout(n24300));
  jand g06278(.dina(n24300), .dinb(n24257), .dout(n24301));
  jor  g06279(.dina(n24301), .dinb(n24299), .dout(n24302));
  jand g06280(.dina(n24302), .dinb(n405), .dout(n24303));
  jand g06281(.dina(n24258), .dinb(n24062), .dout(n24304));
  jxor g06282(.dina(n24228), .dinb(n24227), .dout(n24305));
  jand g06283(.dina(n24305), .dinb(n24257), .dout(n24306));
  jor  g06284(.dina(n24306), .dinb(n24304), .dout(n24307));
  jand g06285(.dina(n24307), .dinb(n2714), .dout(n24308));
  jand g06286(.dina(n24258), .dinb(n24067), .dout(n24309));
  jxor g06287(.dina(n24225), .dinb(n24224), .dout(n24310));
  jand g06288(.dina(n24310), .dinb(n24257), .dout(n24311));
  jor  g06289(.dina(n24311), .dinb(n24309), .dout(n24312));
  jand g06290(.dina(n24312), .dinb(n2547), .dout(n24313));
  jand g06291(.dina(n24258), .dinb(n24072), .dout(n24314));
  jxor g06292(.dina(n24222), .dinb(n24221), .dout(n24315));
  jand g06293(.dina(n24315), .dinb(n24257), .dout(n24316));
  jor  g06294(.dina(n24316), .dinb(n24314), .dout(n24317));
  jand g06295(.dina(n24317), .dinb(n417), .dout(n24318));
  jand g06296(.dina(n24258), .dinb(n24077), .dout(n24319));
  jxor g06297(.dina(n24219), .dinb(n24218), .dout(n24320));
  jand g06298(.dina(n24320), .dinb(n24257), .dout(n24321));
  jor  g06299(.dina(n24321), .dinb(n24319), .dout(n24322));
  jand g06300(.dina(n24322), .dinb(n416), .dout(n24323));
  jand g06301(.dina(n24258), .dinb(n24082), .dout(n24324));
  jxor g06302(.dina(n24216), .dinb(n24215), .dout(n24325));
  jand g06303(.dina(n24325), .dinb(n24257), .dout(n24326));
  jor  g06304(.dina(n24326), .dinb(n24324), .dout(n24327));
  jand g06305(.dina(n24327), .dinb(n422), .dout(n24328));
  jand g06306(.dina(n24258), .dinb(n24087), .dout(n24329));
  jxor g06307(.dina(n24213), .dinb(n24212), .dout(n24330));
  jand g06308(.dina(n24330), .dinb(n24257), .dout(n24331));
  jor  g06309(.dina(n24331), .dinb(n24329), .dout(n24332));
  jand g06310(.dina(n24332), .dinb(n421), .dout(n24333));
  jand g06311(.dina(n24258), .dinb(n24092), .dout(n24334));
  jxor g06312(.dina(n24210), .dinb(n24209), .dout(n24335));
  jand g06313(.dina(n24335), .dinb(n24257), .dout(n24336));
  jor  g06314(.dina(n24336), .dinb(n24334), .dout(n24337));
  jand g06315(.dina(n24337), .dinb(n433), .dout(n24338));
  jand g06316(.dina(n24258), .dinb(n24097), .dout(n24339));
  jxor g06317(.dina(n24207), .dinb(n24206), .dout(n24340));
  jand g06318(.dina(n24340), .dinb(n24257), .dout(n24341));
  jor  g06319(.dina(n24341), .dinb(n24339), .dout(n24342));
  jand g06320(.dina(n24342), .dinb(n432), .dout(n24343));
  jand g06321(.dina(n24258), .dinb(n24102), .dout(n24344));
  jxor g06322(.dina(n24204), .dinb(n24203), .dout(n24345));
  jand g06323(.dina(n24345), .dinb(n24257), .dout(n24346));
  jor  g06324(.dina(n24346), .dinb(n24344), .dout(n24347));
  jand g06325(.dina(n24347), .dinb(n436), .dout(n24348));
  jand g06326(.dina(n24258), .dinb(n24107), .dout(n24349));
  jxor g06327(.dina(n24201), .dinb(n24200), .dout(n24350));
  jand g06328(.dina(n24350), .dinb(n24257), .dout(n24351));
  jor  g06329(.dina(n24351), .dinb(n24349), .dout(n24352));
  jand g06330(.dina(n24352), .dinb(n435), .dout(n24353));
  jand g06331(.dina(n24258), .dinb(n24112), .dout(n24354));
  jxor g06332(.dina(n24198), .dinb(n24197), .dout(n24355));
  jand g06333(.dina(n24355), .dinb(n24257), .dout(n24356));
  jor  g06334(.dina(n24356), .dinb(n24354), .dout(n24357));
  jand g06335(.dina(n24357), .dinb(n440), .dout(n24358));
  jand g06336(.dina(n24258), .dinb(n24117), .dout(n24359));
  jxor g06337(.dina(n24195), .dinb(n24194), .dout(n24360));
  jand g06338(.dina(n24360), .dinb(n24257), .dout(n24361));
  jor  g06339(.dina(n24361), .dinb(n24359), .dout(n24362));
  jand g06340(.dina(n24362), .dinb(n439), .dout(n24363));
  jand g06341(.dina(n24258), .dinb(n24122), .dout(n24364));
  jxor g06342(.dina(n24192), .dinb(n24191), .dout(n24365));
  jand g06343(.dina(n24365), .dinb(n24257), .dout(n24366));
  jor  g06344(.dina(n24366), .dinb(n24364), .dout(n24367));
  jand g06345(.dina(n24367), .dinb(n325), .dout(n24368));
  jand g06346(.dina(n24258), .dinb(n24127), .dout(n24369));
  jxor g06347(.dina(n24189), .dinb(n24188), .dout(n24370));
  jand g06348(.dina(n24370), .dinb(n24257), .dout(n24371));
  jor  g06349(.dina(n24371), .dinb(n24369), .dout(n24372));
  jand g06350(.dina(n24372), .dinb(n324), .dout(n24373));
  jand g06351(.dina(n24258), .dinb(n24132), .dout(n24374));
  jxor g06352(.dina(n24186), .dinb(n24185), .dout(n24375));
  jand g06353(.dina(n24375), .dinb(n24257), .dout(n24376));
  jor  g06354(.dina(n24376), .dinb(n24374), .dout(n24377));
  jand g06355(.dina(n24377), .dinb(n323), .dout(n24378));
  jand g06356(.dina(n24258), .dinb(n24137), .dout(n24379));
  jxor g06357(.dina(n24183), .dinb(n24182), .dout(n24380));
  jand g06358(.dina(n24380), .dinb(n24257), .dout(n24381));
  jor  g06359(.dina(n24381), .dinb(n24379), .dout(n24382));
  jand g06360(.dina(n24382), .dinb(n335), .dout(n24383));
  jand g06361(.dina(n24258), .dinb(n24142), .dout(n24384));
  jxor g06362(.dina(n24180), .dinb(n24179), .dout(n24385));
  jand g06363(.dina(n24385), .dinb(n24257), .dout(n24386));
  jor  g06364(.dina(n24386), .dinb(n24384), .dout(n24387));
  jand g06365(.dina(n24387), .dinb(n334), .dout(n24388));
  jand g06366(.dina(n24258), .dinb(n24147), .dout(n24389));
  jxor g06367(.dina(n24177), .dinb(n24176), .dout(n24390));
  jand g06368(.dina(n24390), .dinb(n24257), .dout(n24391));
  jor  g06369(.dina(n24391), .dinb(n24389), .dout(n24392));
  jand g06370(.dina(n24392), .dinb(n338), .dout(n24393));
  jand g06371(.dina(n24258), .dinb(n24152), .dout(n24394));
  jxor g06372(.dina(n24174), .dinb(n24173), .dout(n24395));
  jand g06373(.dina(n24395), .dinb(n24257), .dout(n24396));
  jor  g06374(.dina(n24396), .dinb(n24394), .dout(n24397));
  jand g06375(.dina(n24397), .dinb(n337), .dout(n24398));
  jnot g06376(.din(n24157), .dout(n24399));
  jor  g06377(.dina(n24257), .dinb(n24399), .dout(n24400));
  jxor g06378(.dina(n24171), .dinb(n24170), .dout(n24401));
  jnot g06379(.din(n24401), .dout(n24402));
  jor  g06380(.dina(n24402), .dinb(n24258), .dout(n24403));
  jand g06381(.dina(n24403), .dinb(n24400), .dout(n24404));
  jnot g06382(.din(n24404), .dout(n24405));
  jand g06383(.dina(n24405), .dinb(n344), .dout(n24406));
  jor  g06384(.dina(n24257), .dinb(n24167), .dout(n24407));
  jxor g06385(.dina(n24168), .dinb(n4800), .dout(n24408));
  jand g06386(.dina(n24408), .dinb(n24257), .dout(n24409));
  jnot g06387(.din(n24409), .dout(n24410));
  jand g06388(.dina(n24410), .dinb(n24407), .dout(n24411));
  jor  g06389(.dina(n24411), .dinb(b2 ), .dout(n24412));
  jnot g06390(.din(n24412), .dout(n24413));
  jnot g06391(.din(n4535), .dout(n24414));
  jnot g06392(.din(n24016), .dout(n24415));
  jnot g06393(.din(n24023), .dout(n24416));
  jnot g06394(.din(n24028), .dout(n24417));
  jnot g06395(.din(n24033), .dout(n24418));
  jnot g06396(.din(n24038), .dout(n24419));
  jnot g06397(.din(n24043), .dout(n24420));
  jnot g06398(.din(n24048), .dout(n24421));
  jnot g06399(.din(n24053), .dout(n24422));
  jnot g06400(.din(n24058), .dout(n24423));
  jnot g06401(.din(n24063), .dout(n24424));
  jnot g06402(.din(n24068), .dout(n24425));
  jnot g06403(.din(n24073), .dout(n24426));
  jnot g06404(.din(n24078), .dout(n24427));
  jnot g06405(.din(n24083), .dout(n24428));
  jnot g06406(.din(n24088), .dout(n24429));
  jnot g06407(.din(n24093), .dout(n24430));
  jnot g06408(.din(n24098), .dout(n24431));
  jnot g06409(.din(n24103), .dout(n24432));
  jnot g06410(.din(n24108), .dout(n24433));
  jnot g06411(.din(n24113), .dout(n24434));
  jnot g06412(.din(n24118), .dout(n24435));
  jnot g06413(.din(n24123), .dout(n24436));
  jnot g06414(.din(n24128), .dout(n24437));
  jnot g06415(.din(n24133), .dout(n24438));
  jnot g06416(.din(n24138), .dout(n24439));
  jnot g06417(.din(n24143), .dout(n24440));
  jnot g06418(.din(n24148), .dout(n24441));
  jnot g06419(.din(n24153), .dout(n24442));
  jnot g06420(.din(n24158), .dout(n24443));
  jnot g06421(.din(n24164), .dout(n24444));
  jxor g06422(.dina(n24167), .dinb(n258), .dout(n24445));
  jor  g06423(.dina(n24445), .dinb(n4799), .dout(n24446));
  jand g06424(.dina(n24446), .dinb(n24444), .dout(n24447));
  jnot g06425(.din(n24171), .dout(n24448));
  jor  g06426(.dina(n24448), .dinb(n24447), .dout(n24449));
  jand g06427(.dina(n24449), .dinb(n24443), .dout(n24450));
  jnot g06428(.din(n24174), .dout(n24451));
  jor  g06429(.dina(n24451), .dinb(n24450), .dout(n24452));
  jand g06430(.dina(n24452), .dinb(n24442), .dout(n24453));
  jnot g06431(.din(n24177), .dout(n24454));
  jor  g06432(.dina(n24454), .dinb(n24453), .dout(n24455));
  jand g06433(.dina(n24455), .dinb(n24441), .dout(n24456));
  jnot g06434(.din(n24180), .dout(n24457));
  jor  g06435(.dina(n24457), .dinb(n24456), .dout(n24458));
  jand g06436(.dina(n24458), .dinb(n24440), .dout(n24459));
  jnot g06437(.din(n24183), .dout(n24460));
  jor  g06438(.dina(n24460), .dinb(n24459), .dout(n24461));
  jand g06439(.dina(n24461), .dinb(n24439), .dout(n24462));
  jnot g06440(.din(n24186), .dout(n24463));
  jor  g06441(.dina(n24463), .dinb(n24462), .dout(n24464));
  jand g06442(.dina(n24464), .dinb(n24438), .dout(n24465));
  jnot g06443(.din(n24189), .dout(n24466));
  jor  g06444(.dina(n24466), .dinb(n24465), .dout(n24467));
  jand g06445(.dina(n24467), .dinb(n24437), .dout(n24468));
  jnot g06446(.din(n24192), .dout(n24469));
  jor  g06447(.dina(n24469), .dinb(n24468), .dout(n24470));
  jand g06448(.dina(n24470), .dinb(n24436), .dout(n24471));
  jnot g06449(.din(n24195), .dout(n24472));
  jor  g06450(.dina(n24472), .dinb(n24471), .dout(n24473));
  jand g06451(.dina(n24473), .dinb(n24435), .dout(n24474));
  jnot g06452(.din(n24198), .dout(n24475));
  jor  g06453(.dina(n24475), .dinb(n24474), .dout(n24476));
  jand g06454(.dina(n24476), .dinb(n24434), .dout(n24477));
  jnot g06455(.din(n24201), .dout(n24478));
  jor  g06456(.dina(n24478), .dinb(n24477), .dout(n24479));
  jand g06457(.dina(n24479), .dinb(n24433), .dout(n24480));
  jnot g06458(.din(n24204), .dout(n24481));
  jor  g06459(.dina(n24481), .dinb(n24480), .dout(n24482));
  jand g06460(.dina(n24482), .dinb(n24432), .dout(n24483));
  jnot g06461(.din(n24207), .dout(n24484));
  jor  g06462(.dina(n24484), .dinb(n24483), .dout(n24485));
  jand g06463(.dina(n24485), .dinb(n24431), .dout(n24486));
  jnot g06464(.din(n24210), .dout(n24487));
  jor  g06465(.dina(n24487), .dinb(n24486), .dout(n24488));
  jand g06466(.dina(n24488), .dinb(n24430), .dout(n24489));
  jnot g06467(.din(n24213), .dout(n24490));
  jor  g06468(.dina(n24490), .dinb(n24489), .dout(n24491));
  jand g06469(.dina(n24491), .dinb(n24429), .dout(n24492));
  jnot g06470(.din(n24216), .dout(n24493));
  jor  g06471(.dina(n24493), .dinb(n24492), .dout(n24494));
  jand g06472(.dina(n24494), .dinb(n24428), .dout(n24495));
  jnot g06473(.din(n24219), .dout(n24496));
  jor  g06474(.dina(n24496), .dinb(n24495), .dout(n24497));
  jand g06475(.dina(n24497), .dinb(n24427), .dout(n24498));
  jnot g06476(.din(n24222), .dout(n24499));
  jor  g06477(.dina(n24499), .dinb(n24498), .dout(n24500));
  jand g06478(.dina(n24500), .dinb(n24426), .dout(n24501));
  jnot g06479(.din(n24225), .dout(n24502));
  jor  g06480(.dina(n24502), .dinb(n24501), .dout(n24503));
  jand g06481(.dina(n24503), .dinb(n24425), .dout(n24504));
  jnot g06482(.din(n24228), .dout(n24505));
  jor  g06483(.dina(n24505), .dinb(n24504), .dout(n24506));
  jand g06484(.dina(n24506), .dinb(n24424), .dout(n24507));
  jnot g06485(.din(n24231), .dout(n24508));
  jor  g06486(.dina(n24508), .dinb(n24507), .dout(n24509));
  jand g06487(.dina(n24509), .dinb(n24423), .dout(n24510));
  jnot g06488(.din(n24234), .dout(n24511));
  jor  g06489(.dina(n24511), .dinb(n24510), .dout(n24512));
  jand g06490(.dina(n24512), .dinb(n24422), .dout(n24513));
  jnot g06491(.din(n24237), .dout(n24514));
  jor  g06492(.dina(n24514), .dinb(n24513), .dout(n24515));
  jand g06493(.dina(n24515), .dinb(n24421), .dout(n24516));
  jnot g06494(.din(n24240), .dout(n24517));
  jor  g06495(.dina(n24517), .dinb(n24516), .dout(n24518));
  jand g06496(.dina(n24518), .dinb(n24420), .dout(n24519));
  jnot g06497(.din(n24243), .dout(n24520));
  jor  g06498(.dina(n24520), .dinb(n24519), .dout(n24521));
  jand g06499(.dina(n24521), .dinb(n24419), .dout(n24522));
  jnot g06500(.din(n24246), .dout(n24523));
  jor  g06501(.dina(n24523), .dinb(n24522), .dout(n24524));
  jand g06502(.dina(n24524), .dinb(n24418), .dout(n24525));
  jnot g06503(.din(n24249), .dout(n24526));
  jor  g06504(.dina(n24526), .dinb(n24525), .dout(n24527));
  jand g06505(.dina(n24527), .dinb(n24417), .dout(n24528));
  jnot g06506(.din(n24252), .dout(n24529));
  jor  g06507(.dina(n24529), .dinb(n24528), .dout(n24530));
  jand g06508(.dina(n24530), .dinb(n24416), .dout(n24531));
  jand g06509(.dina(n24531), .dinb(n24415), .dout(n24532));
  jor  g06510(.dina(n24532), .dinb(n24014), .dout(n24533));
  jor  g06511(.dina(n24533), .dinb(n24414), .dout(n24534));
  jand g06512(.dina(n24534), .dinb(a33 ), .dout(n24535));
  jnot g06513(.din(n5046), .dout(n24536));
  jor  g06514(.dina(n24533), .dinb(n24536), .dout(n24537));
  jnot g06515(.din(n24537), .dout(n24538));
  jor  g06516(.dina(n24538), .dinb(n24535), .dout(n24539));
  jand g06517(.dina(n24539), .dinb(n258), .dout(n24540));
  jand g06518(.dina(n24256), .dinb(n4535), .dout(n24541));
  jor  g06519(.dina(n24541), .dinb(n4798), .dout(n24542));
  jand g06520(.dina(n24537), .dinb(n24542), .dout(n24543));
  jxor g06521(.dina(n24543), .dinb(b1 ), .dout(n24544));
  jand g06522(.dina(n24544), .dinb(n5054), .dout(n24545));
  jor  g06523(.dina(n24545), .dinb(n24540), .dout(n24546));
  jxor g06524(.dina(n24411), .dinb(b2 ), .dout(n24547));
  jand g06525(.dina(n24547), .dinb(n24546), .dout(n24548));
  jor  g06526(.dina(n24548), .dinb(n24413), .dout(n24549));
  jxor g06527(.dina(n24404), .dinb(b3 ), .dout(n24550));
  jand g06528(.dina(n24550), .dinb(n24549), .dout(n24551));
  jor  g06529(.dina(n24551), .dinb(n24406), .dout(n24552));
  jxor g06530(.dina(n24397), .dinb(n337), .dout(n24553));
  jand g06531(.dina(n24553), .dinb(n24552), .dout(n24554));
  jor  g06532(.dina(n24554), .dinb(n24398), .dout(n24555));
  jxor g06533(.dina(n24392), .dinb(n338), .dout(n24556));
  jand g06534(.dina(n24556), .dinb(n24555), .dout(n24557));
  jor  g06535(.dina(n24557), .dinb(n24393), .dout(n24558));
  jxor g06536(.dina(n24387), .dinb(n334), .dout(n24559));
  jand g06537(.dina(n24559), .dinb(n24558), .dout(n24560));
  jor  g06538(.dina(n24560), .dinb(n24388), .dout(n24561));
  jxor g06539(.dina(n24382), .dinb(n335), .dout(n24562));
  jand g06540(.dina(n24562), .dinb(n24561), .dout(n24563));
  jor  g06541(.dina(n24563), .dinb(n24383), .dout(n24564));
  jxor g06542(.dina(n24377), .dinb(n323), .dout(n24565));
  jand g06543(.dina(n24565), .dinb(n24564), .dout(n24566));
  jor  g06544(.dina(n24566), .dinb(n24378), .dout(n24567));
  jxor g06545(.dina(n24372), .dinb(n324), .dout(n24568));
  jand g06546(.dina(n24568), .dinb(n24567), .dout(n24569));
  jor  g06547(.dina(n24569), .dinb(n24373), .dout(n24570));
  jxor g06548(.dina(n24367), .dinb(n325), .dout(n24571));
  jand g06549(.dina(n24571), .dinb(n24570), .dout(n24572));
  jor  g06550(.dina(n24572), .dinb(n24368), .dout(n24573));
  jxor g06551(.dina(n24362), .dinb(n439), .dout(n24574));
  jand g06552(.dina(n24574), .dinb(n24573), .dout(n24575));
  jor  g06553(.dina(n24575), .dinb(n24363), .dout(n24576));
  jxor g06554(.dina(n24357), .dinb(n440), .dout(n24577));
  jand g06555(.dina(n24577), .dinb(n24576), .dout(n24578));
  jor  g06556(.dina(n24578), .dinb(n24358), .dout(n24579));
  jxor g06557(.dina(n24352), .dinb(n435), .dout(n24580));
  jand g06558(.dina(n24580), .dinb(n24579), .dout(n24581));
  jor  g06559(.dina(n24581), .dinb(n24353), .dout(n24582));
  jxor g06560(.dina(n24347), .dinb(n436), .dout(n24583));
  jand g06561(.dina(n24583), .dinb(n24582), .dout(n24584));
  jor  g06562(.dina(n24584), .dinb(n24348), .dout(n24585));
  jxor g06563(.dina(n24342), .dinb(n432), .dout(n24586));
  jand g06564(.dina(n24586), .dinb(n24585), .dout(n24587));
  jor  g06565(.dina(n24587), .dinb(n24343), .dout(n24588));
  jxor g06566(.dina(n24337), .dinb(n433), .dout(n24589));
  jand g06567(.dina(n24589), .dinb(n24588), .dout(n24590));
  jor  g06568(.dina(n24590), .dinb(n24338), .dout(n24591));
  jxor g06569(.dina(n24332), .dinb(n421), .dout(n24592));
  jand g06570(.dina(n24592), .dinb(n24591), .dout(n24593));
  jor  g06571(.dina(n24593), .dinb(n24333), .dout(n24594));
  jxor g06572(.dina(n24327), .dinb(n422), .dout(n24595));
  jand g06573(.dina(n24595), .dinb(n24594), .dout(n24596));
  jor  g06574(.dina(n24596), .dinb(n24328), .dout(n24597));
  jxor g06575(.dina(n24322), .dinb(n416), .dout(n24598));
  jand g06576(.dina(n24598), .dinb(n24597), .dout(n24599));
  jor  g06577(.dina(n24599), .dinb(n24323), .dout(n24600));
  jxor g06578(.dina(n24317), .dinb(n417), .dout(n24601));
  jand g06579(.dina(n24601), .dinb(n24600), .dout(n24602));
  jor  g06580(.dina(n24602), .dinb(n24318), .dout(n24603));
  jxor g06581(.dina(n24312), .dinb(n2547), .dout(n24604));
  jand g06582(.dina(n24604), .dinb(n24603), .dout(n24605));
  jor  g06583(.dina(n24605), .dinb(n24313), .dout(n24606));
  jxor g06584(.dina(n24307), .dinb(n2714), .dout(n24607));
  jand g06585(.dina(n24607), .dinb(n24606), .dout(n24608));
  jor  g06586(.dina(n24608), .dinb(n24308), .dout(n24609));
  jxor g06587(.dina(n24302), .dinb(n405), .dout(n24610));
  jand g06588(.dina(n24610), .dinb(n24609), .dout(n24611));
  jor  g06589(.dina(n24611), .dinb(n24303), .dout(n24612));
  jxor g06590(.dina(n24297), .dinb(n406), .dout(n24613));
  jand g06591(.dina(n24613), .dinb(n24612), .dout(n24614));
  jor  g06592(.dina(n24614), .dinb(n24298), .dout(n24615));
  jxor g06593(.dina(n24292), .dinb(n412), .dout(n24616));
  jand g06594(.dina(n24616), .dinb(n24615), .dout(n24617));
  jor  g06595(.dina(n24617), .dinb(n24293), .dout(n24618));
  jxor g06596(.dina(n24287), .dinb(n413), .dout(n24619));
  jand g06597(.dina(n24619), .dinb(n24618), .dout(n24620));
  jor  g06598(.dina(n24620), .dinb(n24288), .dout(n24621));
  jxor g06599(.dina(n24282), .dinb(n409), .dout(n24622));
  jand g06600(.dina(n24622), .dinb(n24621), .dout(n24623));
  jor  g06601(.dina(n24623), .dinb(n24283), .dout(n24624));
  jxor g06602(.dina(n24277), .dinb(n410), .dout(n24625));
  jand g06603(.dina(n24625), .dinb(n24624), .dout(n24626));
  jor  g06604(.dina(n24626), .dinb(n24278), .dout(n24627));
  jxor g06605(.dina(n24272), .dinb(n426), .dout(n24628));
  jand g06606(.dina(n24628), .dinb(n24627), .dout(n24629));
  jor  g06607(.dina(n24629), .dinb(n24273), .dout(n24630));
  jxor g06608(.dina(n24267), .dinb(n427), .dout(n24631));
  jand g06609(.dina(n24631), .dinb(n24630), .dout(n24632));
  jor  g06610(.dina(n24632), .dinb(n24268), .dout(n24633));
  jnot g06611(.din(n24262), .dout(n24634));
  jand g06612(.dina(n24634), .dinb(b31 ), .dout(n24635));
  jnot g06613(.din(n24635), .dout(n24636));
  jand g06614(.dina(n24636), .dinb(n24633), .dout(n24637));
  jor  g06615(.dina(n24637), .dinb(n24263), .dout(n24638));
  jand g06616(.dina(n24638), .dinb(n590), .dout(n24639));
  jnot g06617(.din(n24639), .dout(n24640));
  jand g06618(.dina(n24640), .dinb(n24262), .dout(n24641));
  jand g06619(.dina(n24263), .dinb(n590), .dout(n24642));
  jand g06620(.dina(n24642), .dinb(n24633), .dout(n24643));
  jor  g06621(.dina(n24643), .dinb(n24641), .dout(n24644));
  jand g06622(.dina(n24644), .dinb(n590), .dout(n24645));
  jnot g06623(.din(n24645), .dout(n24646));
  jnot g06624(.din(n403), .dout(n24647));
  jand g06625(.dina(n24640), .dinb(n24267), .dout(n24648));
  jxor g06626(.dina(n24631), .dinb(n24630), .dout(n24649));
  jand g06627(.dina(n24649), .dinb(n24639), .dout(n24650));
  jor  g06628(.dina(n24650), .dinb(n24648), .dout(n24651));
  jand g06629(.dina(n24651), .dinb(n424), .dout(n24652));
  jnot g06630(.din(n24652), .dout(n24653));
  jand g06631(.dina(n24640), .dinb(n24272), .dout(n24654));
  jxor g06632(.dina(n24628), .dinb(n24627), .dout(n24655));
  jand g06633(.dina(n24655), .dinb(n24639), .dout(n24656));
  jor  g06634(.dina(n24656), .dinb(n24654), .dout(n24657));
  jand g06635(.dina(n24657), .dinb(n427), .dout(n24658));
  jnot g06636(.din(n24658), .dout(n24659));
  jand g06637(.dina(n24640), .dinb(n24277), .dout(n24660));
  jxor g06638(.dina(n24625), .dinb(n24624), .dout(n24661));
  jand g06639(.dina(n24661), .dinb(n24639), .dout(n24662));
  jor  g06640(.dina(n24662), .dinb(n24660), .dout(n24663));
  jand g06641(.dina(n24663), .dinb(n426), .dout(n24664));
  jnot g06642(.din(n24664), .dout(n24665));
  jand g06643(.dina(n24640), .dinb(n24282), .dout(n24666));
  jxor g06644(.dina(n24622), .dinb(n24621), .dout(n24667));
  jand g06645(.dina(n24667), .dinb(n24639), .dout(n24668));
  jor  g06646(.dina(n24668), .dinb(n24666), .dout(n24669));
  jand g06647(.dina(n24669), .dinb(n410), .dout(n24670));
  jnot g06648(.din(n24670), .dout(n24671));
  jand g06649(.dina(n24640), .dinb(n24287), .dout(n24672));
  jxor g06650(.dina(n24619), .dinb(n24618), .dout(n24673));
  jand g06651(.dina(n24673), .dinb(n24639), .dout(n24674));
  jor  g06652(.dina(n24674), .dinb(n24672), .dout(n24675));
  jand g06653(.dina(n24675), .dinb(n409), .dout(n24676));
  jnot g06654(.din(n24676), .dout(n24677));
  jand g06655(.dina(n24640), .dinb(n24292), .dout(n24678));
  jxor g06656(.dina(n24616), .dinb(n24615), .dout(n24679));
  jand g06657(.dina(n24679), .dinb(n24639), .dout(n24680));
  jor  g06658(.dina(n24680), .dinb(n24678), .dout(n24681));
  jand g06659(.dina(n24681), .dinb(n413), .dout(n24682));
  jnot g06660(.din(n24682), .dout(n24683));
  jand g06661(.dina(n24640), .dinb(n24297), .dout(n24684));
  jxor g06662(.dina(n24613), .dinb(n24612), .dout(n24685));
  jand g06663(.dina(n24685), .dinb(n24639), .dout(n24686));
  jor  g06664(.dina(n24686), .dinb(n24684), .dout(n24687));
  jand g06665(.dina(n24687), .dinb(n412), .dout(n24688));
  jnot g06666(.din(n24688), .dout(n24689));
  jand g06667(.dina(n24640), .dinb(n24302), .dout(n24690));
  jxor g06668(.dina(n24610), .dinb(n24609), .dout(n24691));
  jand g06669(.dina(n24691), .dinb(n24639), .dout(n24692));
  jor  g06670(.dina(n24692), .dinb(n24690), .dout(n24693));
  jand g06671(.dina(n24693), .dinb(n406), .dout(n24694));
  jnot g06672(.din(n24694), .dout(n24695));
  jand g06673(.dina(n24640), .dinb(n24307), .dout(n24696));
  jxor g06674(.dina(n24607), .dinb(n24606), .dout(n24697));
  jand g06675(.dina(n24697), .dinb(n24639), .dout(n24698));
  jor  g06676(.dina(n24698), .dinb(n24696), .dout(n24699));
  jand g06677(.dina(n24699), .dinb(n405), .dout(n24700));
  jnot g06678(.din(n24700), .dout(n24701));
  jand g06679(.dina(n24640), .dinb(n24312), .dout(n24702));
  jxor g06680(.dina(n24604), .dinb(n24603), .dout(n24703));
  jand g06681(.dina(n24703), .dinb(n24639), .dout(n24704));
  jor  g06682(.dina(n24704), .dinb(n24702), .dout(n24705));
  jand g06683(.dina(n24705), .dinb(n2714), .dout(n24706));
  jnot g06684(.din(n24706), .dout(n24707));
  jand g06685(.dina(n24640), .dinb(n24317), .dout(n24708));
  jxor g06686(.dina(n24601), .dinb(n24600), .dout(n24709));
  jand g06687(.dina(n24709), .dinb(n24639), .dout(n24710));
  jor  g06688(.dina(n24710), .dinb(n24708), .dout(n24711));
  jand g06689(.dina(n24711), .dinb(n2547), .dout(n24712));
  jnot g06690(.din(n24712), .dout(n24713));
  jand g06691(.dina(n24640), .dinb(n24322), .dout(n24714));
  jxor g06692(.dina(n24598), .dinb(n24597), .dout(n24715));
  jand g06693(.dina(n24715), .dinb(n24639), .dout(n24716));
  jor  g06694(.dina(n24716), .dinb(n24714), .dout(n24717));
  jand g06695(.dina(n24717), .dinb(n417), .dout(n24718));
  jnot g06696(.din(n24718), .dout(n24719));
  jand g06697(.dina(n24640), .dinb(n24327), .dout(n24720));
  jxor g06698(.dina(n24595), .dinb(n24594), .dout(n24721));
  jand g06699(.dina(n24721), .dinb(n24639), .dout(n24722));
  jor  g06700(.dina(n24722), .dinb(n24720), .dout(n24723));
  jand g06701(.dina(n24723), .dinb(n416), .dout(n24724));
  jnot g06702(.din(n24724), .dout(n24725));
  jand g06703(.dina(n24640), .dinb(n24332), .dout(n24726));
  jxor g06704(.dina(n24592), .dinb(n24591), .dout(n24727));
  jand g06705(.dina(n24727), .dinb(n24639), .dout(n24728));
  jor  g06706(.dina(n24728), .dinb(n24726), .dout(n24729));
  jand g06707(.dina(n24729), .dinb(n422), .dout(n24730));
  jnot g06708(.din(n24730), .dout(n24731));
  jand g06709(.dina(n24640), .dinb(n24337), .dout(n24732));
  jxor g06710(.dina(n24589), .dinb(n24588), .dout(n24733));
  jand g06711(.dina(n24733), .dinb(n24639), .dout(n24734));
  jor  g06712(.dina(n24734), .dinb(n24732), .dout(n24735));
  jand g06713(.dina(n24735), .dinb(n421), .dout(n24736));
  jnot g06714(.din(n24736), .dout(n24737));
  jand g06715(.dina(n24640), .dinb(n24342), .dout(n24738));
  jxor g06716(.dina(n24586), .dinb(n24585), .dout(n24739));
  jand g06717(.dina(n24739), .dinb(n24639), .dout(n24740));
  jor  g06718(.dina(n24740), .dinb(n24738), .dout(n24741));
  jand g06719(.dina(n24741), .dinb(n433), .dout(n24742));
  jnot g06720(.din(n24742), .dout(n24743));
  jand g06721(.dina(n24640), .dinb(n24347), .dout(n24744));
  jxor g06722(.dina(n24583), .dinb(n24582), .dout(n24745));
  jand g06723(.dina(n24745), .dinb(n24639), .dout(n24746));
  jor  g06724(.dina(n24746), .dinb(n24744), .dout(n24747));
  jand g06725(.dina(n24747), .dinb(n432), .dout(n24748));
  jnot g06726(.din(n24748), .dout(n24749));
  jand g06727(.dina(n24640), .dinb(n24352), .dout(n24750));
  jxor g06728(.dina(n24580), .dinb(n24579), .dout(n24751));
  jand g06729(.dina(n24751), .dinb(n24639), .dout(n24752));
  jor  g06730(.dina(n24752), .dinb(n24750), .dout(n24753));
  jand g06731(.dina(n24753), .dinb(n436), .dout(n24754));
  jnot g06732(.din(n24754), .dout(n24755));
  jand g06733(.dina(n24640), .dinb(n24357), .dout(n24756));
  jxor g06734(.dina(n24577), .dinb(n24576), .dout(n24757));
  jand g06735(.dina(n24757), .dinb(n24639), .dout(n24758));
  jor  g06736(.dina(n24758), .dinb(n24756), .dout(n24759));
  jand g06737(.dina(n24759), .dinb(n435), .dout(n24760));
  jnot g06738(.din(n24760), .dout(n24761));
  jand g06739(.dina(n24640), .dinb(n24362), .dout(n24762));
  jxor g06740(.dina(n24574), .dinb(n24573), .dout(n24763));
  jand g06741(.dina(n24763), .dinb(n24639), .dout(n24764));
  jor  g06742(.dina(n24764), .dinb(n24762), .dout(n24765));
  jand g06743(.dina(n24765), .dinb(n440), .dout(n24766));
  jnot g06744(.din(n24766), .dout(n24767));
  jand g06745(.dina(n24640), .dinb(n24367), .dout(n24768));
  jxor g06746(.dina(n24571), .dinb(n24570), .dout(n24769));
  jand g06747(.dina(n24769), .dinb(n24639), .dout(n24770));
  jor  g06748(.dina(n24770), .dinb(n24768), .dout(n24771));
  jand g06749(.dina(n24771), .dinb(n439), .dout(n24772));
  jnot g06750(.din(n24772), .dout(n24773));
  jand g06751(.dina(n24640), .dinb(n24372), .dout(n24774));
  jxor g06752(.dina(n24568), .dinb(n24567), .dout(n24775));
  jand g06753(.dina(n24775), .dinb(n24639), .dout(n24776));
  jor  g06754(.dina(n24776), .dinb(n24774), .dout(n24777));
  jand g06755(.dina(n24777), .dinb(n325), .dout(n24778));
  jnot g06756(.din(n24778), .dout(n24779));
  jand g06757(.dina(n24640), .dinb(n24377), .dout(n24780));
  jxor g06758(.dina(n24565), .dinb(n24564), .dout(n24781));
  jand g06759(.dina(n24781), .dinb(n24639), .dout(n24782));
  jor  g06760(.dina(n24782), .dinb(n24780), .dout(n24783));
  jand g06761(.dina(n24783), .dinb(n324), .dout(n24784));
  jnot g06762(.din(n24784), .dout(n24785));
  jand g06763(.dina(n24640), .dinb(n24382), .dout(n24786));
  jxor g06764(.dina(n24562), .dinb(n24561), .dout(n24787));
  jand g06765(.dina(n24787), .dinb(n24639), .dout(n24788));
  jor  g06766(.dina(n24788), .dinb(n24786), .dout(n24789));
  jand g06767(.dina(n24789), .dinb(n323), .dout(n24790));
  jnot g06768(.din(n24790), .dout(n24791));
  jand g06769(.dina(n24640), .dinb(n24387), .dout(n24792));
  jxor g06770(.dina(n24559), .dinb(n24558), .dout(n24793));
  jand g06771(.dina(n24793), .dinb(n24639), .dout(n24794));
  jor  g06772(.dina(n24794), .dinb(n24792), .dout(n24795));
  jand g06773(.dina(n24795), .dinb(n335), .dout(n24796));
  jnot g06774(.din(n24796), .dout(n24797));
  jand g06775(.dina(n24640), .dinb(n24392), .dout(n24798));
  jxor g06776(.dina(n24556), .dinb(n24555), .dout(n24799));
  jand g06777(.dina(n24799), .dinb(n24639), .dout(n24800));
  jor  g06778(.dina(n24800), .dinb(n24798), .dout(n24801));
  jand g06779(.dina(n24801), .dinb(n334), .dout(n24802));
  jnot g06780(.din(n24802), .dout(n24803));
  jand g06781(.dina(n24640), .dinb(n24397), .dout(n24804));
  jxor g06782(.dina(n24553), .dinb(n24552), .dout(n24805));
  jand g06783(.dina(n24805), .dinb(n24639), .dout(n24806));
  jor  g06784(.dina(n24806), .dinb(n24804), .dout(n24807));
  jand g06785(.dina(n24807), .dinb(n338), .dout(n24808));
  jnot g06786(.din(n24808), .dout(n24809));
  jand g06787(.dina(n24640), .dinb(n24405), .dout(n24810));
  jxor g06788(.dina(n24550), .dinb(n24549), .dout(n24811));
  jand g06789(.dina(n24811), .dinb(n24639), .dout(n24812));
  jor  g06790(.dina(n24812), .dinb(n24810), .dout(n24813));
  jand g06791(.dina(n24813), .dinb(n337), .dout(n24814));
  jnot g06792(.din(n24814), .dout(n24815));
  jor  g06793(.dina(n24639), .dinb(n24411), .dout(n24816));
  jxor g06794(.dina(n24547), .dinb(n24546), .dout(n24817));
  jnot g06795(.din(n24817), .dout(n24818));
  jor  g06796(.dina(n24818), .dinb(n24640), .dout(n24819));
  jand g06797(.dina(n24819), .dinb(n24816), .dout(n24820));
  jnot g06798(.din(n24820), .dout(n24821));
  jand g06799(.dina(n24821), .dinb(n344), .dout(n24822));
  jnot g06800(.din(n24822), .dout(n24823));
  jor  g06801(.dina(n24639), .dinb(n24543), .dout(n24824));
  jxor g06802(.dina(n24544), .dinb(n5054), .dout(n24825));
  jand g06803(.dina(n24825), .dinb(n24639), .dout(n24826));
  jnot g06804(.din(n24826), .dout(n24827));
  jand g06805(.dina(n24827), .dinb(n24824), .dout(n24828));
  jnot g06806(.din(n24828), .dout(n24829));
  jand g06807(.dina(n24829), .dinb(n348), .dout(n24830));
  jnot g06808(.din(n24830), .dout(n24831));
  jnot g06809(.din(n5308), .dout(n24832));
  jnot g06810(.din(n24263), .dout(n24833));
  jnot g06811(.din(n24268), .dout(n24834));
  jnot g06812(.din(n24273), .dout(n24835));
  jnot g06813(.din(n24278), .dout(n24836));
  jnot g06814(.din(n24283), .dout(n24837));
  jnot g06815(.din(n24288), .dout(n24838));
  jnot g06816(.din(n24293), .dout(n24839));
  jnot g06817(.din(n24298), .dout(n24840));
  jnot g06818(.din(n24303), .dout(n24841));
  jnot g06819(.din(n24308), .dout(n24842));
  jnot g06820(.din(n24313), .dout(n24843));
  jnot g06821(.din(n24318), .dout(n24844));
  jnot g06822(.din(n24323), .dout(n24845));
  jnot g06823(.din(n24328), .dout(n24846));
  jnot g06824(.din(n24333), .dout(n24847));
  jnot g06825(.din(n24338), .dout(n24848));
  jnot g06826(.din(n24343), .dout(n24849));
  jnot g06827(.din(n24348), .dout(n24850));
  jnot g06828(.din(n24353), .dout(n24851));
  jnot g06829(.din(n24358), .dout(n24852));
  jnot g06830(.din(n24363), .dout(n24853));
  jnot g06831(.din(n24368), .dout(n24854));
  jnot g06832(.din(n24373), .dout(n24855));
  jnot g06833(.din(n24378), .dout(n24856));
  jnot g06834(.din(n24383), .dout(n24857));
  jnot g06835(.din(n24388), .dout(n24858));
  jnot g06836(.din(n24393), .dout(n24859));
  jnot g06837(.din(n24398), .dout(n24860));
  jnot g06838(.din(n24406), .dout(n24861));
  jnot g06839(.din(n24540), .dout(n24862));
  jxor g06840(.dina(n24543), .dinb(n258), .dout(n24863));
  jor  g06841(.dina(n24863), .dinb(n5053), .dout(n24864));
  jand g06842(.dina(n24864), .dinb(n24862), .dout(n24865));
  jnot g06843(.din(n24547), .dout(n24866));
  jor  g06844(.dina(n24866), .dinb(n24865), .dout(n24867));
  jand g06845(.dina(n24867), .dinb(n24412), .dout(n24868));
  jnot g06846(.din(n24550), .dout(n24869));
  jor  g06847(.dina(n24869), .dinb(n24868), .dout(n24870));
  jand g06848(.dina(n24870), .dinb(n24861), .dout(n24871));
  jnot g06849(.din(n24553), .dout(n24872));
  jor  g06850(.dina(n24872), .dinb(n24871), .dout(n24873));
  jand g06851(.dina(n24873), .dinb(n24860), .dout(n24874));
  jnot g06852(.din(n24556), .dout(n24875));
  jor  g06853(.dina(n24875), .dinb(n24874), .dout(n24876));
  jand g06854(.dina(n24876), .dinb(n24859), .dout(n24877));
  jnot g06855(.din(n24559), .dout(n24878));
  jor  g06856(.dina(n24878), .dinb(n24877), .dout(n24879));
  jand g06857(.dina(n24879), .dinb(n24858), .dout(n24880));
  jnot g06858(.din(n24562), .dout(n24881));
  jor  g06859(.dina(n24881), .dinb(n24880), .dout(n24882));
  jand g06860(.dina(n24882), .dinb(n24857), .dout(n24883));
  jnot g06861(.din(n24565), .dout(n24884));
  jor  g06862(.dina(n24884), .dinb(n24883), .dout(n24885));
  jand g06863(.dina(n24885), .dinb(n24856), .dout(n24886));
  jnot g06864(.din(n24568), .dout(n24887));
  jor  g06865(.dina(n24887), .dinb(n24886), .dout(n24888));
  jand g06866(.dina(n24888), .dinb(n24855), .dout(n24889));
  jnot g06867(.din(n24571), .dout(n24890));
  jor  g06868(.dina(n24890), .dinb(n24889), .dout(n24891));
  jand g06869(.dina(n24891), .dinb(n24854), .dout(n24892));
  jnot g06870(.din(n24574), .dout(n24893));
  jor  g06871(.dina(n24893), .dinb(n24892), .dout(n24894));
  jand g06872(.dina(n24894), .dinb(n24853), .dout(n24895));
  jnot g06873(.din(n24577), .dout(n24896));
  jor  g06874(.dina(n24896), .dinb(n24895), .dout(n24897));
  jand g06875(.dina(n24897), .dinb(n24852), .dout(n24898));
  jnot g06876(.din(n24580), .dout(n24899));
  jor  g06877(.dina(n24899), .dinb(n24898), .dout(n24900));
  jand g06878(.dina(n24900), .dinb(n24851), .dout(n24901));
  jnot g06879(.din(n24583), .dout(n24902));
  jor  g06880(.dina(n24902), .dinb(n24901), .dout(n24903));
  jand g06881(.dina(n24903), .dinb(n24850), .dout(n24904));
  jnot g06882(.din(n24586), .dout(n24905));
  jor  g06883(.dina(n24905), .dinb(n24904), .dout(n24906));
  jand g06884(.dina(n24906), .dinb(n24849), .dout(n24907));
  jnot g06885(.din(n24589), .dout(n24908));
  jor  g06886(.dina(n24908), .dinb(n24907), .dout(n24909));
  jand g06887(.dina(n24909), .dinb(n24848), .dout(n24910));
  jnot g06888(.din(n24592), .dout(n24911));
  jor  g06889(.dina(n24911), .dinb(n24910), .dout(n24912));
  jand g06890(.dina(n24912), .dinb(n24847), .dout(n24913));
  jnot g06891(.din(n24595), .dout(n24914));
  jor  g06892(.dina(n24914), .dinb(n24913), .dout(n24915));
  jand g06893(.dina(n24915), .dinb(n24846), .dout(n24916));
  jnot g06894(.din(n24598), .dout(n24917));
  jor  g06895(.dina(n24917), .dinb(n24916), .dout(n24918));
  jand g06896(.dina(n24918), .dinb(n24845), .dout(n24919));
  jnot g06897(.din(n24601), .dout(n24920));
  jor  g06898(.dina(n24920), .dinb(n24919), .dout(n24921));
  jand g06899(.dina(n24921), .dinb(n24844), .dout(n24922));
  jnot g06900(.din(n24604), .dout(n24923));
  jor  g06901(.dina(n24923), .dinb(n24922), .dout(n24924));
  jand g06902(.dina(n24924), .dinb(n24843), .dout(n24925));
  jnot g06903(.din(n24607), .dout(n24926));
  jor  g06904(.dina(n24926), .dinb(n24925), .dout(n24927));
  jand g06905(.dina(n24927), .dinb(n24842), .dout(n24928));
  jnot g06906(.din(n24610), .dout(n24929));
  jor  g06907(.dina(n24929), .dinb(n24928), .dout(n24930));
  jand g06908(.dina(n24930), .dinb(n24841), .dout(n24931));
  jnot g06909(.din(n24613), .dout(n24932));
  jor  g06910(.dina(n24932), .dinb(n24931), .dout(n24933));
  jand g06911(.dina(n24933), .dinb(n24840), .dout(n24934));
  jnot g06912(.din(n24616), .dout(n24935));
  jor  g06913(.dina(n24935), .dinb(n24934), .dout(n24936));
  jand g06914(.dina(n24936), .dinb(n24839), .dout(n24937));
  jnot g06915(.din(n24619), .dout(n24938));
  jor  g06916(.dina(n24938), .dinb(n24937), .dout(n24939));
  jand g06917(.dina(n24939), .dinb(n24838), .dout(n24940));
  jnot g06918(.din(n24622), .dout(n24941));
  jor  g06919(.dina(n24941), .dinb(n24940), .dout(n24942));
  jand g06920(.dina(n24942), .dinb(n24837), .dout(n24943));
  jnot g06921(.din(n24625), .dout(n24944));
  jor  g06922(.dina(n24944), .dinb(n24943), .dout(n24945));
  jand g06923(.dina(n24945), .dinb(n24836), .dout(n24946));
  jnot g06924(.din(n24628), .dout(n24947));
  jor  g06925(.dina(n24947), .dinb(n24946), .dout(n24948));
  jand g06926(.dina(n24948), .dinb(n24835), .dout(n24949));
  jnot g06927(.din(n24631), .dout(n24950));
  jor  g06928(.dina(n24950), .dinb(n24949), .dout(n24951));
  jand g06929(.dina(n24951), .dinb(n24834), .dout(n24952));
  jor  g06930(.dina(n24635), .dinb(n24952), .dout(n24953));
  jand g06931(.dina(n24953), .dinb(n24833), .dout(n24954));
  jor  g06932(.dina(n24954), .dinb(n24832), .dout(n24955));
  jand g06933(.dina(n24955), .dinb(a32 ), .dout(n24956));
  jnot g06934(.din(n5311), .dout(n24957));
  jor  g06935(.dina(n24954), .dinb(n24957), .dout(n24958));
  jnot g06936(.din(n24958), .dout(n24959));
  jor  g06937(.dina(n24959), .dinb(n24956), .dout(n24960));
  jand g06938(.dina(n24960), .dinb(n258), .dout(n24961));
  jnot g06939(.din(n24961), .dout(n24962));
  jand g06940(.dina(n24638), .dinb(n5308), .dout(n24963));
  jor  g06941(.dina(n24963), .dinb(n5052), .dout(n24964));
  jand g06942(.dina(n24958), .dinb(n24964), .dout(n24965));
  jxor g06943(.dina(n24965), .dinb(n258), .dout(n24966));
  jor  g06944(.dina(n24966), .dinb(n5318), .dout(n24967));
  jand g06945(.dina(n24967), .dinb(n24962), .dout(n24968));
  jxor g06946(.dina(n24828), .dinb(b2 ), .dout(n24969));
  jnot g06947(.din(n24969), .dout(n24970));
  jor  g06948(.dina(n24970), .dinb(n24968), .dout(n24971));
  jand g06949(.dina(n24971), .dinb(n24831), .dout(n24972));
  jxor g06950(.dina(n24820), .dinb(b3 ), .dout(n24973));
  jnot g06951(.din(n24973), .dout(n24974));
  jor  g06952(.dina(n24974), .dinb(n24972), .dout(n24975));
  jand g06953(.dina(n24975), .dinb(n24823), .dout(n24976));
  jxor g06954(.dina(n24813), .dinb(n337), .dout(n24977));
  jnot g06955(.din(n24977), .dout(n24978));
  jor  g06956(.dina(n24978), .dinb(n24976), .dout(n24979));
  jand g06957(.dina(n24979), .dinb(n24815), .dout(n24980));
  jxor g06958(.dina(n24807), .dinb(n338), .dout(n24981));
  jnot g06959(.din(n24981), .dout(n24982));
  jor  g06960(.dina(n24982), .dinb(n24980), .dout(n24983));
  jand g06961(.dina(n24983), .dinb(n24809), .dout(n24984));
  jxor g06962(.dina(n24801), .dinb(n334), .dout(n24985));
  jnot g06963(.din(n24985), .dout(n24986));
  jor  g06964(.dina(n24986), .dinb(n24984), .dout(n24987));
  jand g06965(.dina(n24987), .dinb(n24803), .dout(n24988));
  jxor g06966(.dina(n24795), .dinb(n335), .dout(n24989));
  jnot g06967(.din(n24989), .dout(n24990));
  jor  g06968(.dina(n24990), .dinb(n24988), .dout(n24991));
  jand g06969(.dina(n24991), .dinb(n24797), .dout(n24992));
  jxor g06970(.dina(n24789), .dinb(n323), .dout(n24993));
  jnot g06971(.din(n24993), .dout(n24994));
  jor  g06972(.dina(n24994), .dinb(n24992), .dout(n24995));
  jand g06973(.dina(n24995), .dinb(n24791), .dout(n24996));
  jxor g06974(.dina(n24783), .dinb(n324), .dout(n24997));
  jnot g06975(.din(n24997), .dout(n24998));
  jor  g06976(.dina(n24998), .dinb(n24996), .dout(n24999));
  jand g06977(.dina(n24999), .dinb(n24785), .dout(n25000));
  jxor g06978(.dina(n24777), .dinb(n325), .dout(n25001));
  jnot g06979(.din(n25001), .dout(n25002));
  jor  g06980(.dina(n25002), .dinb(n25000), .dout(n25003));
  jand g06981(.dina(n25003), .dinb(n24779), .dout(n25004));
  jxor g06982(.dina(n24771), .dinb(n439), .dout(n25005));
  jnot g06983(.din(n25005), .dout(n25006));
  jor  g06984(.dina(n25006), .dinb(n25004), .dout(n25007));
  jand g06985(.dina(n25007), .dinb(n24773), .dout(n25008));
  jxor g06986(.dina(n24765), .dinb(n440), .dout(n25009));
  jnot g06987(.din(n25009), .dout(n25010));
  jor  g06988(.dina(n25010), .dinb(n25008), .dout(n25011));
  jand g06989(.dina(n25011), .dinb(n24767), .dout(n25012));
  jxor g06990(.dina(n24759), .dinb(n435), .dout(n25013));
  jnot g06991(.din(n25013), .dout(n25014));
  jor  g06992(.dina(n25014), .dinb(n25012), .dout(n25015));
  jand g06993(.dina(n25015), .dinb(n24761), .dout(n25016));
  jxor g06994(.dina(n24753), .dinb(n436), .dout(n25017));
  jnot g06995(.din(n25017), .dout(n25018));
  jor  g06996(.dina(n25018), .dinb(n25016), .dout(n25019));
  jand g06997(.dina(n25019), .dinb(n24755), .dout(n25020));
  jxor g06998(.dina(n24747), .dinb(n432), .dout(n25021));
  jnot g06999(.din(n25021), .dout(n25022));
  jor  g07000(.dina(n25022), .dinb(n25020), .dout(n25023));
  jand g07001(.dina(n25023), .dinb(n24749), .dout(n25024));
  jxor g07002(.dina(n24741), .dinb(n433), .dout(n25025));
  jnot g07003(.din(n25025), .dout(n25026));
  jor  g07004(.dina(n25026), .dinb(n25024), .dout(n25027));
  jand g07005(.dina(n25027), .dinb(n24743), .dout(n25028));
  jxor g07006(.dina(n24735), .dinb(n421), .dout(n25029));
  jnot g07007(.din(n25029), .dout(n25030));
  jor  g07008(.dina(n25030), .dinb(n25028), .dout(n25031));
  jand g07009(.dina(n25031), .dinb(n24737), .dout(n25032));
  jxor g07010(.dina(n24729), .dinb(n422), .dout(n25033));
  jnot g07011(.din(n25033), .dout(n25034));
  jor  g07012(.dina(n25034), .dinb(n25032), .dout(n25035));
  jand g07013(.dina(n25035), .dinb(n24731), .dout(n25036));
  jxor g07014(.dina(n24723), .dinb(n416), .dout(n25037));
  jnot g07015(.din(n25037), .dout(n25038));
  jor  g07016(.dina(n25038), .dinb(n25036), .dout(n25039));
  jand g07017(.dina(n25039), .dinb(n24725), .dout(n25040));
  jxor g07018(.dina(n24717), .dinb(n417), .dout(n25041));
  jnot g07019(.din(n25041), .dout(n25042));
  jor  g07020(.dina(n25042), .dinb(n25040), .dout(n25043));
  jand g07021(.dina(n25043), .dinb(n24719), .dout(n25044));
  jxor g07022(.dina(n24711), .dinb(n2547), .dout(n25045));
  jnot g07023(.din(n25045), .dout(n25046));
  jor  g07024(.dina(n25046), .dinb(n25044), .dout(n25047));
  jand g07025(.dina(n25047), .dinb(n24713), .dout(n25048));
  jxor g07026(.dina(n24705), .dinb(n2714), .dout(n25049));
  jnot g07027(.din(n25049), .dout(n25050));
  jor  g07028(.dina(n25050), .dinb(n25048), .dout(n25051));
  jand g07029(.dina(n25051), .dinb(n24707), .dout(n25052));
  jxor g07030(.dina(n24699), .dinb(n405), .dout(n25053));
  jnot g07031(.din(n25053), .dout(n25054));
  jor  g07032(.dina(n25054), .dinb(n25052), .dout(n25055));
  jand g07033(.dina(n25055), .dinb(n24701), .dout(n25056));
  jxor g07034(.dina(n24693), .dinb(n406), .dout(n25057));
  jnot g07035(.din(n25057), .dout(n25058));
  jor  g07036(.dina(n25058), .dinb(n25056), .dout(n25059));
  jand g07037(.dina(n25059), .dinb(n24695), .dout(n25060));
  jxor g07038(.dina(n24687), .dinb(n412), .dout(n25061));
  jnot g07039(.din(n25061), .dout(n25062));
  jor  g07040(.dina(n25062), .dinb(n25060), .dout(n25063));
  jand g07041(.dina(n25063), .dinb(n24689), .dout(n25064));
  jxor g07042(.dina(n24681), .dinb(n413), .dout(n25065));
  jnot g07043(.din(n25065), .dout(n25066));
  jor  g07044(.dina(n25066), .dinb(n25064), .dout(n25067));
  jand g07045(.dina(n25067), .dinb(n24683), .dout(n25068));
  jxor g07046(.dina(n24675), .dinb(n409), .dout(n25069));
  jnot g07047(.din(n25069), .dout(n25070));
  jor  g07048(.dina(n25070), .dinb(n25068), .dout(n25071));
  jand g07049(.dina(n25071), .dinb(n24677), .dout(n25072));
  jxor g07050(.dina(n24669), .dinb(n410), .dout(n25073));
  jnot g07051(.din(n25073), .dout(n25074));
  jor  g07052(.dina(n25074), .dinb(n25072), .dout(n25075));
  jand g07053(.dina(n25075), .dinb(n24671), .dout(n25076));
  jxor g07054(.dina(n24663), .dinb(n426), .dout(n25077));
  jnot g07055(.din(n25077), .dout(n25078));
  jor  g07056(.dina(n25078), .dinb(n25076), .dout(n25079));
  jand g07057(.dina(n25079), .dinb(n24665), .dout(n25080));
  jxor g07058(.dina(n24657), .dinb(n427), .dout(n25081));
  jnot g07059(.din(n25081), .dout(n25082));
  jor  g07060(.dina(n25082), .dinb(n25080), .dout(n25083));
  jand g07061(.dina(n25083), .dinb(n24659), .dout(n25084));
  jxor g07062(.dina(n24651), .dinb(n424), .dout(n25085));
  jnot g07063(.din(n25085), .dout(n25086));
  jor  g07064(.dina(n25086), .dinb(n25084), .dout(n25087));
  jand g07065(.dina(n25087), .dinb(n24653), .dout(n25088));
  jxor g07066(.dina(n24644), .dinb(b32 ), .dout(n25089));
  jor  g07067(.dina(n25089), .dinb(n25088), .dout(n25090));
  jor  g07068(.dina(n25090), .dinb(n24647), .dout(n25091));
  jand g07069(.dina(n25091), .dinb(n24646), .dout(n25092));
  jand g07070(.dina(n25092), .dinb(n24644), .dout(n25093));
  jnot g07071(.din(n25093), .dout(n25094));
  jxor g07072(.dina(n24965), .dinb(b1 ), .dout(n25095));
  jand g07073(.dina(n25095), .dinb(n5319), .dout(n25096));
  jor  g07074(.dina(n25096), .dinb(n24961), .dout(n25097));
  jand g07075(.dina(n24969), .dinb(n25097), .dout(n25098));
  jor  g07076(.dina(n25098), .dinb(n24830), .dout(n25099));
  jand g07077(.dina(n24973), .dinb(n25099), .dout(n25100));
  jor  g07078(.dina(n25100), .dinb(n24822), .dout(n25101));
  jand g07079(.dina(n24977), .dinb(n25101), .dout(n25102));
  jor  g07080(.dina(n25102), .dinb(n24814), .dout(n25103));
  jand g07081(.dina(n24981), .dinb(n25103), .dout(n25104));
  jor  g07082(.dina(n25104), .dinb(n24808), .dout(n25105));
  jand g07083(.dina(n24985), .dinb(n25105), .dout(n25106));
  jor  g07084(.dina(n25106), .dinb(n24802), .dout(n25107));
  jand g07085(.dina(n24989), .dinb(n25107), .dout(n25108));
  jor  g07086(.dina(n25108), .dinb(n24796), .dout(n25109));
  jand g07087(.dina(n24993), .dinb(n25109), .dout(n25110));
  jor  g07088(.dina(n25110), .dinb(n24790), .dout(n25111));
  jand g07089(.dina(n24997), .dinb(n25111), .dout(n25112));
  jor  g07090(.dina(n25112), .dinb(n24784), .dout(n25113));
  jand g07091(.dina(n25001), .dinb(n25113), .dout(n25114));
  jor  g07092(.dina(n25114), .dinb(n24778), .dout(n25115));
  jand g07093(.dina(n25005), .dinb(n25115), .dout(n25116));
  jor  g07094(.dina(n25116), .dinb(n24772), .dout(n25117));
  jand g07095(.dina(n25009), .dinb(n25117), .dout(n25118));
  jor  g07096(.dina(n25118), .dinb(n24766), .dout(n25119));
  jand g07097(.dina(n25013), .dinb(n25119), .dout(n25120));
  jor  g07098(.dina(n25120), .dinb(n24760), .dout(n25121));
  jand g07099(.dina(n25017), .dinb(n25121), .dout(n25122));
  jor  g07100(.dina(n25122), .dinb(n24754), .dout(n25123));
  jand g07101(.dina(n25021), .dinb(n25123), .dout(n25124));
  jor  g07102(.dina(n25124), .dinb(n24748), .dout(n25125));
  jand g07103(.dina(n25025), .dinb(n25125), .dout(n25126));
  jor  g07104(.dina(n25126), .dinb(n24742), .dout(n25127));
  jand g07105(.dina(n25029), .dinb(n25127), .dout(n25128));
  jor  g07106(.dina(n25128), .dinb(n24736), .dout(n25129));
  jand g07107(.dina(n25033), .dinb(n25129), .dout(n25130));
  jor  g07108(.dina(n25130), .dinb(n24730), .dout(n25131));
  jand g07109(.dina(n25037), .dinb(n25131), .dout(n25132));
  jor  g07110(.dina(n25132), .dinb(n24724), .dout(n25133));
  jand g07111(.dina(n25041), .dinb(n25133), .dout(n25134));
  jor  g07112(.dina(n25134), .dinb(n24718), .dout(n25135));
  jand g07113(.dina(n25045), .dinb(n25135), .dout(n25136));
  jor  g07114(.dina(n25136), .dinb(n24712), .dout(n25137));
  jand g07115(.dina(n25049), .dinb(n25137), .dout(n25138));
  jor  g07116(.dina(n25138), .dinb(n24706), .dout(n25139));
  jand g07117(.dina(n25053), .dinb(n25139), .dout(n25140));
  jor  g07118(.dina(n25140), .dinb(n24700), .dout(n25141));
  jand g07119(.dina(n25057), .dinb(n25141), .dout(n25142));
  jor  g07120(.dina(n25142), .dinb(n24694), .dout(n25143));
  jand g07121(.dina(n25061), .dinb(n25143), .dout(n25144));
  jor  g07122(.dina(n25144), .dinb(n24688), .dout(n25145));
  jand g07123(.dina(n25065), .dinb(n25145), .dout(n25146));
  jor  g07124(.dina(n25146), .dinb(n24682), .dout(n25147));
  jand g07125(.dina(n25069), .dinb(n25147), .dout(n25148));
  jor  g07126(.dina(n25148), .dinb(n24676), .dout(n25149));
  jand g07127(.dina(n25073), .dinb(n25149), .dout(n25150));
  jor  g07128(.dina(n25150), .dinb(n24670), .dout(n25151));
  jand g07129(.dina(n25077), .dinb(n25151), .dout(n25152));
  jor  g07130(.dina(n25152), .dinb(n24664), .dout(n25153));
  jand g07131(.dina(n25081), .dinb(n25153), .dout(n25154));
  jor  g07132(.dina(n25154), .dinb(n24658), .dout(n25155));
  jand g07133(.dina(n25085), .dinb(n25155), .dout(n25156));
  jor  g07134(.dina(n25156), .dinb(n24652), .dout(n25157));
  jnot g07135(.din(n25089), .dout(n25158));
  jand g07136(.dina(n25158), .dinb(n25157), .dout(n25159));
  jand g07137(.dina(n25088), .dinb(n300), .dout(n25160));
  jor  g07138(.dina(n25160), .dinb(n24646), .dout(n25161));
  jor  g07139(.dina(n25161), .dinb(n25159), .dout(n25162));
  jand g07140(.dina(n25162), .dinb(n25094), .dout(n25163));
  jnot g07141(.din(n25163), .dout(n25164));
  jand g07142(.dina(n25164), .dinb(n297), .dout(n25165));
  jand g07143(.dina(n25092), .dinb(n24651), .dout(n25166));
  jand g07144(.dina(n25159), .dinb(n403), .dout(n25167));
  jor  g07145(.dina(n25167), .dinb(n24645), .dout(n25168));
  jxor g07146(.dina(n25085), .dinb(n25155), .dout(n25169));
  jand g07147(.dina(n25169), .dinb(n25168), .dout(n25170));
  jor  g07148(.dina(n25170), .dinb(n25166), .dout(n25171));
  jand g07149(.dina(n25171), .dinb(n300), .dout(n25172));
  jand g07150(.dina(n25092), .dinb(n24657), .dout(n25173));
  jxor g07151(.dina(n25081), .dinb(n25153), .dout(n25174));
  jand g07152(.dina(n25174), .dinb(n25168), .dout(n25175));
  jor  g07153(.dina(n25175), .dinb(n25173), .dout(n25176));
  jand g07154(.dina(n25176), .dinb(n424), .dout(n25177));
  jand g07155(.dina(n25092), .dinb(n24663), .dout(n25178));
  jxor g07156(.dina(n25077), .dinb(n25151), .dout(n25179));
  jand g07157(.dina(n25179), .dinb(n25168), .dout(n25180));
  jor  g07158(.dina(n25180), .dinb(n25178), .dout(n25181));
  jand g07159(.dina(n25181), .dinb(n427), .dout(n25182));
  jand g07160(.dina(n25092), .dinb(n24669), .dout(n25183));
  jxor g07161(.dina(n25073), .dinb(n25149), .dout(n25184));
  jand g07162(.dina(n25184), .dinb(n25168), .dout(n25185));
  jor  g07163(.dina(n25185), .dinb(n25183), .dout(n25186));
  jand g07164(.dina(n25186), .dinb(n426), .dout(n25187));
  jand g07165(.dina(n25092), .dinb(n24675), .dout(n25188));
  jxor g07166(.dina(n25069), .dinb(n25147), .dout(n25189));
  jand g07167(.dina(n25189), .dinb(n25168), .dout(n25190));
  jor  g07168(.dina(n25190), .dinb(n25188), .dout(n25191));
  jand g07169(.dina(n25191), .dinb(n410), .dout(n25192));
  jand g07170(.dina(n25092), .dinb(n24681), .dout(n25193));
  jxor g07171(.dina(n25065), .dinb(n25145), .dout(n25194));
  jand g07172(.dina(n25194), .dinb(n25168), .dout(n25195));
  jor  g07173(.dina(n25195), .dinb(n25193), .dout(n25196));
  jand g07174(.dina(n25196), .dinb(n409), .dout(n25197));
  jand g07175(.dina(n25092), .dinb(n24687), .dout(n25198));
  jxor g07176(.dina(n25061), .dinb(n25143), .dout(n25199));
  jand g07177(.dina(n25199), .dinb(n25168), .dout(n25200));
  jor  g07178(.dina(n25200), .dinb(n25198), .dout(n25201));
  jand g07179(.dina(n25201), .dinb(n413), .dout(n25202));
  jand g07180(.dina(n25092), .dinb(n24693), .dout(n25203));
  jxor g07181(.dina(n25057), .dinb(n25141), .dout(n25204));
  jand g07182(.dina(n25204), .dinb(n25168), .dout(n25205));
  jor  g07183(.dina(n25205), .dinb(n25203), .dout(n25206));
  jand g07184(.dina(n25206), .dinb(n412), .dout(n25207));
  jand g07185(.dina(n25092), .dinb(n24699), .dout(n25208));
  jxor g07186(.dina(n25053), .dinb(n25139), .dout(n25209));
  jand g07187(.dina(n25209), .dinb(n25168), .dout(n25210));
  jor  g07188(.dina(n25210), .dinb(n25208), .dout(n25211));
  jand g07189(.dina(n25211), .dinb(n406), .dout(n25212));
  jand g07190(.dina(n25092), .dinb(n24705), .dout(n25213));
  jxor g07191(.dina(n25049), .dinb(n25137), .dout(n25214));
  jand g07192(.dina(n25214), .dinb(n25168), .dout(n25215));
  jor  g07193(.dina(n25215), .dinb(n25213), .dout(n25216));
  jand g07194(.dina(n25216), .dinb(n405), .dout(n25217));
  jand g07195(.dina(n25092), .dinb(n24711), .dout(n25218));
  jxor g07196(.dina(n25045), .dinb(n25135), .dout(n25219));
  jand g07197(.dina(n25219), .dinb(n25168), .dout(n25220));
  jor  g07198(.dina(n25220), .dinb(n25218), .dout(n25221));
  jand g07199(.dina(n25221), .dinb(n2714), .dout(n25222));
  jand g07200(.dina(n25092), .dinb(n24717), .dout(n25223));
  jxor g07201(.dina(n25041), .dinb(n25133), .dout(n25224));
  jand g07202(.dina(n25224), .dinb(n25168), .dout(n25225));
  jor  g07203(.dina(n25225), .dinb(n25223), .dout(n25226));
  jand g07204(.dina(n25226), .dinb(n2547), .dout(n25227));
  jand g07205(.dina(n25092), .dinb(n24723), .dout(n25228));
  jxor g07206(.dina(n25037), .dinb(n25131), .dout(n25229));
  jand g07207(.dina(n25229), .dinb(n25168), .dout(n25230));
  jor  g07208(.dina(n25230), .dinb(n25228), .dout(n25231));
  jand g07209(.dina(n25231), .dinb(n417), .dout(n25232));
  jand g07210(.dina(n25092), .dinb(n24729), .dout(n25233));
  jxor g07211(.dina(n25033), .dinb(n25129), .dout(n25234));
  jand g07212(.dina(n25234), .dinb(n25168), .dout(n25235));
  jor  g07213(.dina(n25235), .dinb(n25233), .dout(n25236));
  jand g07214(.dina(n25236), .dinb(n416), .dout(n25237));
  jand g07215(.dina(n25092), .dinb(n24735), .dout(n25238));
  jxor g07216(.dina(n25029), .dinb(n25127), .dout(n25239));
  jand g07217(.dina(n25239), .dinb(n25168), .dout(n25240));
  jor  g07218(.dina(n25240), .dinb(n25238), .dout(n25241));
  jand g07219(.dina(n25241), .dinb(n422), .dout(n25242));
  jand g07220(.dina(n25092), .dinb(n24741), .dout(n25243));
  jxor g07221(.dina(n25025), .dinb(n25125), .dout(n25244));
  jand g07222(.dina(n25244), .dinb(n25168), .dout(n25245));
  jor  g07223(.dina(n25245), .dinb(n25243), .dout(n25246));
  jand g07224(.dina(n25246), .dinb(n421), .dout(n25247));
  jand g07225(.dina(n25092), .dinb(n24747), .dout(n25248));
  jxor g07226(.dina(n25021), .dinb(n25123), .dout(n25249));
  jand g07227(.dina(n25249), .dinb(n25168), .dout(n25250));
  jor  g07228(.dina(n25250), .dinb(n25248), .dout(n25251));
  jand g07229(.dina(n25251), .dinb(n433), .dout(n25252));
  jand g07230(.dina(n25092), .dinb(n24753), .dout(n25253));
  jxor g07231(.dina(n25017), .dinb(n25121), .dout(n25254));
  jand g07232(.dina(n25254), .dinb(n25168), .dout(n25255));
  jor  g07233(.dina(n25255), .dinb(n25253), .dout(n25256));
  jand g07234(.dina(n25256), .dinb(n432), .dout(n25257));
  jand g07235(.dina(n25092), .dinb(n24759), .dout(n25258));
  jxor g07236(.dina(n25013), .dinb(n25119), .dout(n25259));
  jand g07237(.dina(n25259), .dinb(n25168), .dout(n25260));
  jor  g07238(.dina(n25260), .dinb(n25258), .dout(n25261));
  jand g07239(.dina(n25261), .dinb(n436), .dout(n25262));
  jand g07240(.dina(n25092), .dinb(n24765), .dout(n25263));
  jxor g07241(.dina(n25009), .dinb(n25117), .dout(n25264));
  jand g07242(.dina(n25264), .dinb(n25168), .dout(n25265));
  jor  g07243(.dina(n25265), .dinb(n25263), .dout(n25266));
  jand g07244(.dina(n25266), .dinb(n435), .dout(n25267));
  jand g07245(.dina(n25092), .dinb(n24771), .dout(n25268));
  jxor g07246(.dina(n25005), .dinb(n25115), .dout(n25269));
  jand g07247(.dina(n25269), .dinb(n25168), .dout(n25270));
  jor  g07248(.dina(n25270), .dinb(n25268), .dout(n25271));
  jand g07249(.dina(n25271), .dinb(n440), .dout(n25272));
  jand g07250(.dina(n25092), .dinb(n24777), .dout(n25273));
  jxor g07251(.dina(n25001), .dinb(n25113), .dout(n25274));
  jand g07252(.dina(n25274), .dinb(n25168), .dout(n25275));
  jor  g07253(.dina(n25275), .dinb(n25273), .dout(n25276));
  jand g07254(.dina(n25276), .dinb(n439), .dout(n25277));
  jand g07255(.dina(n25092), .dinb(n24783), .dout(n25278));
  jxor g07256(.dina(n24997), .dinb(n25111), .dout(n25279));
  jand g07257(.dina(n25279), .dinb(n25168), .dout(n25280));
  jor  g07258(.dina(n25280), .dinb(n25278), .dout(n25281));
  jand g07259(.dina(n25281), .dinb(n325), .dout(n25282));
  jand g07260(.dina(n25092), .dinb(n24789), .dout(n25283));
  jxor g07261(.dina(n24993), .dinb(n25109), .dout(n25284));
  jand g07262(.dina(n25284), .dinb(n25168), .dout(n25285));
  jor  g07263(.dina(n25285), .dinb(n25283), .dout(n25286));
  jand g07264(.dina(n25286), .dinb(n324), .dout(n25287));
  jand g07265(.dina(n25092), .dinb(n24795), .dout(n25288));
  jxor g07266(.dina(n24989), .dinb(n25107), .dout(n25289));
  jand g07267(.dina(n25289), .dinb(n25168), .dout(n25290));
  jor  g07268(.dina(n25290), .dinb(n25288), .dout(n25291));
  jand g07269(.dina(n25291), .dinb(n323), .dout(n25292));
  jand g07270(.dina(n25092), .dinb(n24801), .dout(n25293));
  jxor g07271(.dina(n24985), .dinb(n25105), .dout(n25294));
  jand g07272(.dina(n25294), .dinb(n25168), .dout(n25295));
  jor  g07273(.dina(n25295), .dinb(n25293), .dout(n25296));
  jand g07274(.dina(n25296), .dinb(n335), .dout(n25297));
  jand g07275(.dina(n25092), .dinb(n24807), .dout(n25298));
  jxor g07276(.dina(n24981), .dinb(n25103), .dout(n25299));
  jand g07277(.dina(n25299), .dinb(n25168), .dout(n25300));
  jor  g07278(.dina(n25300), .dinb(n25298), .dout(n25301));
  jand g07279(.dina(n25301), .dinb(n334), .dout(n25302));
  jand g07280(.dina(n25092), .dinb(n24813), .dout(n25303));
  jxor g07281(.dina(n24977), .dinb(n25101), .dout(n25304));
  jand g07282(.dina(n25304), .dinb(n25168), .dout(n25305));
  jor  g07283(.dina(n25305), .dinb(n25303), .dout(n25306));
  jand g07284(.dina(n25306), .dinb(n338), .dout(n25307));
  jand g07285(.dina(n25092), .dinb(n24821), .dout(n25308));
  jxor g07286(.dina(n24973), .dinb(n25099), .dout(n25309));
  jand g07287(.dina(n25309), .dinb(n25168), .dout(n25310));
  jor  g07288(.dina(n25310), .dinb(n25308), .dout(n25311));
  jand g07289(.dina(n25311), .dinb(n337), .dout(n25312));
  jand g07290(.dina(n25092), .dinb(n24829), .dout(n25313));
  jxor g07291(.dina(n24969), .dinb(n25097), .dout(n25314));
  jand g07292(.dina(n25314), .dinb(n25168), .dout(n25315));
  jor  g07293(.dina(n25315), .dinb(n25313), .dout(n25316));
  jand g07294(.dina(n25316), .dinb(n344), .dout(n25317));
  jand g07295(.dina(n25092), .dinb(n24960), .dout(n25318));
  jxor g07296(.dina(n25095), .dinb(n5319), .dout(n25319));
  jand g07297(.dina(n25319), .dinb(n25168), .dout(n25320));
  jor  g07298(.dina(n25320), .dinb(n25318), .dout(n25321));
  jand g07299(.dina(n25321), .dinb(n348), .dout(n25322));
  jor  g07300(.dina(n25092), .dinb(n18364), .dout(n25323));
  jand g07301(.dina(n25323), .dinb(a31 ), .dout(n25324));
  jor  g07302(.dina(n25092), .dinb(n5319), .dout(n25325));
  jnot g07303(.din(n25325), .dout(n25326));
  jor  g07304(.dina(n25326), .dinb(n25324), .dout(n25327));
  jand g07305(.dina(n25327), .dinb(n258), .dout(n25328));
  jand g07306(.dina(n25168), .dinb(b0 ), .dout(n25329));
  jor  g07307(.dina(n25329), .dinb(n5317), .dout(n25330));
  jand g07308(.dina(n25325), .dinb(n25330), .dout(n25331));
  jxor g07309(.dina(n25331), .dinb(b1 ), .dout(n25332));
  jand g07310(.dina(n25332), .dinb(n5593), .dout(n25333));
  jor  g07311(.dina(n25333), .dinb(n25328), .dout(n25334));
  jxor g07312(.dina(n25321), .dinb(n348), .dout(n25335));
  jand g07313(.dina(n25335), .dinb(n25334), .dout(n25336));
  jor  g07314(.dina(n25336), .dinb(n25322), .dout(n25337));
  jxor g07315(.dina(n25316), .dinb(n344), .dout(n25338));
  jand g07316(.dina(n25338), .dinb(n25337), .dout(n25339));
  jor  g07317(.dina(n25339), .dinb(n25317), .dout(n25340));
  jxor g07318(.dina(n25311), .dinb(n337), .dout(n25341));
  jand g07319(.dina(n25341), .dinb(n25340), .dout(n25342));
  jor  g07320(.dina(n25342), .dinb(n25312), .dout(n25343));
  jxor g07321(.dina(n25306), .dinb(n338), .dout(n25344));
  jand g07322(.dina(n25344), .dinb(n25343), .dout(n25345));
  jor  g07323(.dina(n25345), .dinb(n25307), .dout(n25346));
  jxor g07324(.dina(n25301), .dinb(n334), .dout(n25347));
  jand g07325(.dina(n25347), .dinb(n25346), .dout(n25348));
  jor  g07326(.dina(n25348), .dinb(n25302), .dout(n25349));
  jxor g07327(.dina(n25296), .dinb(n335), .dout(n25350));
  jand g07328(.dina(n25350), .dinb(n25349), .dout(n25351));
  jor  g07329(.dina(n25351), .dinb(n25297), .dout(n25352));
  jxor g07330(.dina(n25291), .dinb(n323), .dout(n25353));
  jand g07331(.dina(n25353), .dinb(n25352), .dout(n25354));
  jor  g07332(.dina(n25354), .dinb(n25292), .dout(n25355));
  jxor g07333(.dina(n25286), .dinb(n324), .dout(n25356));
  jand g07334(.dina(n25356), .dinb(n25355), .dout(n25357));
  jor  g07335(.dina(n25357), .dinb(n25287), .dout(n25358));
  jxor g07336(.dina(n25281), .dinb(n325), .dout(n25359));
  jand g07337(.dina(n25359), .dinb(n25358), .dout(n25360));
  jor  g07338(.dina(n25360), .dinb(n25282), .dout(n25361));
  jxor g07339(.dina(n25276), .dinb(n439), .dout(n25362));
  jand g07340(.dina(n25362), .dinb(n25361), .dout(n25363));
  jor  g07341(.dina(n25363), .dinb(n25277), .dout(n25364));
  jxor g07342(.dina(n25271), .dinb(n440), .dout(n25365));
  jand g07343(.dina(n25365), .dinb(n25364), .dout(n25366));
  jor  g07344(.dina(n25366), .dinb(n25272), .dout(n25367));
  jxor g07345(.dina(n25266), .dinb(n435), .dout(n25368));
  jand g07346(.dina(n25368), .dinb(n25367), .dout(n25369));
  jor  g07347(.dina(n25369), .dinb(n25267), .dout(n25370));
  jxor g07348(.dina(n25261), .dinb(n436), .dout(n25371));
  jand g07349(.dina(n25371), .dinb(n25370), .dout(n25372));
  jor  g07350(.dina(n25372), .dinb(n25262), .dout(n25373));
  jxor g07351(.dina(n25256), .dinb(n432), .dout(n25374));
  jand g07352(.dina(n25374), .dinb(n25373), .dout(n25375));
  jor  g07353(.dina(n25375), .dinb(n25257), .dout(n25376));
  jxor g07354(.dina(n25251), .dinb(n433), .dout(n25377));
  jand g07355(.dina(n25377), .dinb(n25376), .dout(n25378));
  jor  g07356(.dina(n25378), .dinb(n25252), .dout(n25379));
  jxor g07357(.dina(n25246), .dinb(n421), .dout(n25380));
  jand g07358(.dina(n25380), .dinb(n25379), .dout(n25381));
  jor  g07359(.dina(n25381), .dinb(n25247), .dout(n25382));
  jxor g07360(.dina(n25241), .dinb(n422), .dout(n25383));
  jand g07361(.dina(n25383), .dinb(n25382), .dout(n25384));
  jor  g07362(.dina(n25384), .dinb(n25242), .dout(n25385));
  jxor g07363(.dina(n25236), .dinb(n416), .dout(n25386));
  jand g07364(.dina(n25386), .dinb(n25385), .dout(n25387));
  jor  g07365(.dina(n25387), .dinb(n25237), .dout(n25388));
  jxor g07366(.dina(n25231), .dinb(n417), .dout(n25389));
  jand g07367(.dina(n25389), .dinb(n25388), .dout(n25390));
  jor  g07368(.dina(n25390), .dinb(n25232), .dout(n25391));
  jxor g07369(.dina(n25226), .dinb(n2547), .dout(n25392));
  jand g07370(.dina(n25392), .dinb(n25391), .dout(n25393));
  jor  g07371(.dina(n25393), .dinb(n25227), .dout(n25394));
  jxor g07372(.dina(n25221), .dinb(n2714), .dout(n25395));
  jand g07373(.dina(n25395), .dinb(n25394), .dout(n25396));
  jor  g07374(.dina(n25396), .dinb(n25222), .dout(n25397));
  jxor g07375(.dina(n25216), .dinb(n405), .dout(n25398));
  jand g07376(.dina(n25398), .dinb(n25397), .dout(n25399));
  jor  g07377(.dina(n25399), .dinb(n25217), .dout(n25400));
  jxor g07378(.dina(n25211), .dinb(n406), .dout(n25401));
  jand g07379(.dina(n25401), .dinb(n25400), .dout(n25402));
  jor  g07380(.dina(n25402), .dinb(n25212), .dout(n25403));
  jxor g07381(.dina(n25206), .dinb(n412), .dout(n25404));
  jand g07382(.dina(n25404), .dinb(n25403), .dout(n25405));
  jor  g07383(.dina(n25405), .dinb(n25207), .dout(n25406));
  jxor g07384(.dina(n25201), .dinb(n413), .dout(n25407));
  jand g07385(.dina(n25407), .dinb(n25406), .dout(n25408));
  jor  g07386(.dina(n25408), .dinb(n25202), .dout(n25409));
  jxor g07387(.dina(n25196), .dinb(n409), .dout(n25410));
  jand g07388(.dina(n25410), .dinb(n25409), .dout(n25411));
  jor  g07389(.dina(n25411), .dinb(n25197), .dout(n25412));
  jxor g07390(.dina(n25191), .dinb(n410), .dout(n25413));
  jand g07391(.dina(n25413), .dinb(n25412), .dout(n25414));
  jor  g07392(.dina(n25414), .dinb(n25192), .dout(n25415));
  jxor g07393(.dina(n25186), .dinb(n426), .dout(n25416));
  jand g07394(.dina(n25416), .dinb(n25415), .dout(n25417));
  jor  g07395(.dina(n25417), .dinb(n25187), .dout(n25418));
  jxor g07396(.dina(n25181), .dinb(n427), .dout(n25419));
  jand g07397(.dina(n25419), .dinb(n25418), .dout(n25420));
  jor  g07398(.dina(n25420), .dinb(n25182), .dout(n25421));
  jxor g07399(.dina(n25176), .dinb(n424), .dout(n25422));
  jand g07400(.dina(n25422), .dinb(n25421), .dout(n25423));
  jor  g07401(.dina(n25423), .dinb(n25177), .dout(n25424));
  jxor g07402(.dina(n25171), .dinb(n300), .dout(n25425));
  jand g07403(.dina(n25425), .dinb(n25424), .dout(n25426));
  jor  g07404(.dina(n25426), .dinb(n25172), .dout(n25427));
  jand g07405(.dina(n25163), .dinb(b33 ), .dout(n25428));
  jnot g07406(.din(n25428), .dout(n25429));
  jand g07407(.dina(n25429), .dinb(n25427), .dout(n25430));
  jor  g07408(.dina(n25430), .dinb(n25165), .dout(n25431));
  jand g07409(.dina(n25431), .dinb(n5694), .dout(n25432));
  jnot g07410(.din(n25432), .dout(n25433));
  jand g07411(.dina(n25433), .dinb(n25164), .dout(n25434));
  jand g07412(.dina(n25165), .dinb(n5694), .dout(n25435));
  jand g07413(.dina(n25435), .dinb(n25427), .dout(n25436));
  jor  g07414(.dina(n25436), .dinb(n25434), .dout(n25437));
  jand g07415(.dina(n25437), .dinb(n298), .dout(n25438));
  jnot g07416(.din(n25438), .dout(n25439));
  jand g07417(.dina(n25433), .dinb(n25171), .dout(n25440));
  jxor g07418(.dina(n25425), .dinb(n25424), .dout(n25441));
  jand g07419(.dina(n25441), .dinb(n25432), .dout(n25442));
  jor  g07420(.dina(n25442), .dinb(n25440), .dout(n25443));
  jand g07421(.dina(n25443), .dinb(n297), .dout(n25444));
  jnot g07422(.din(n25444), .dout(n25445));
  jand g07423(.dina(n25433), .dinb(n25176), .dout(n25446));
  jxor g07424(.dina(n25422), .dinb(n25421), .dout(n25447));
  jand g07425(.dina(n25447), .dinb(n25432), .dout(n25448));
  jor  g07426(.dina(n25448), .dinb(n25446), .dout(n25449));
  jand g07427(.dina(n25449), .dinb(n300), .dout(n25450));
  jnot g07428(.din(n25450), .dout(n25451));
  jand g07429(.dina(n25433), .dinb(n25181), .dout(n25452));
  jxor g07430(.dina(n25419), .dinb(n25418), .dout(n25453));
  jand g07431(.dina(n25453), .dinb(n25432), .dout(n25454));
  jor  g07432(.dina(n25454), .dinb(n25452), .dout(n25455));
  jand g07433(.dina(n25455), .dinb(n424), .dout(n25456));
  jnot g07434(.din(n25456), .dout(n25457));
  jand g07435(.dina(n25433), .dinb(n25186), .dout(n25458));
  jxor g07436(.dina(n25416), .dinb(n25415), .dout(n25459));
  jand g07437(.dina(n25459), .dinb(n25432), .dout(n25460));
  jor  g07438(.dina(n25460), .dinb(n25458), .dout(n25461));
  jand g07439(.dina(n25461), .dinb(n427), .dout(n25462));
  jnot g07440(.din(n25462), .dout(n25463));
  jand g07441(.dina(n25433), .dinb(n25191), .dout(n25464));
  jxor g07442(.dina(n25413), .dinb(n25412), .dout(n25465));
  jand g07443(.dina(n25465), .dinb(n25432), .dout(n25466));
  jor  g07444(.dina(n25466), .dinb(n25464), .dout(n25467));
  jand g07445(.dina(n25467), .dinb(n426), .dout(n25468));
  jnot g07446(.din(n25468), .dout(n25469));
  jand g07447(.dina(n25433), .dinb(n25196), .dout(n25470));
  jxor g07448(.dina(n25410), .dinb(n25409), .dout(n25471));
  jand g07449(.dina(n25471), .dinb(n25432), .dout(n25472));
  jor  g07450(.dina(n25472), .dinb(n25470), .dout(n25473));
  jand g07451(.dina(n25473), .dinb(n410), .dout(n25474));
  jnot g07452(.din(n25474), .dout(n25475));
  jand g07453(.dina(n25433), .dinb(n25201), .dout(n25476));
  jxor g07454(.dina(n25407), .dinb(n25406), .dout(n25477));
  jand g07455(.dina(n25477), .dinb(n25432), .dout(n25478));
  jor  g07456(.dina(n25478), .dinb(n25476), .dout(n25479));
  jand g07457(.dina(n25479), .dinb(n409), .dout(n25480));
  jnot g07458(.din(n25480), .dout(n25481));
  jand g07459(.dina(n25433), .dinb(n25206), .dout(n25482));
  jxor g07460(.dina(n25404), .dinb(n25403), .dout(n25483));
  jand g07461(.dina(n25483), .dinb(n25432), .dout(n25484));
  jor  g07462(.dina(n25484), .dinb(n25482), .dout(n25485));
  jand g07463(.dina(n25485), .dinb(n413), .dout(n25486));
  jnot g07464(.din(n25486), .dout(n25487));
  jand g07465(.dina(n25433), .dinb(n25211), .dout(n25488));
  jxor g07466(.dina(n25401), .dinb(n25400), .dout(n25489));
  jand g07467(.dina(n25489), .dinb(n25432), .dout(n25490));
  jor  g07468(.dina(n25490), .dinb(n25488), .dout(n25491));
  jand g07469(.dina(n25491), .dinb(n412), .dout(n25492));
  jnot g07470(.din(n25492), .dout(n25493));
  jand g07471(.dina(n25433), .dinb(n25216), .dout(n25494));
  jxor g07472(.dina(n25398), .dinb(n25397), .dout(n25495));
  jand g07473(.dina(n25495), .dinb(n25432), .dout(n25496));
  jor  g07474(.dina(n25496), .dinb(n25494), .dout(n25497));
  jand g07475(.dina(n25497), .dinb(n406), .dout(n25498));
  jnot g07476(.din(n25498), .dout(n25499));
  jand g07477(.dina(n25433), .dinb(n25221), .dout(n25500));
  jxor g07478(.dina(n25395), .dinb(n25394), .dout(n25501));
  jand g07479(.dina(n25501), .dinb(n25432), .dout(n25502));
  jor  g07480(.dina(n25502), .dinb(n25500), .dout(n25503));
  jand g07481(.dina(n25503), .dinb(n405), .dout(n25504));
  jnot g07482(.din(n25504), .dout(n25505));
  jand g07483(.dina(n25433), .dinb(n25226), .dout(n25506));
  jxor g07484(.dina(n25392), .dinb(n25391), .dout(n25507));
  jand g07485(.dina(n25507), .dinb(n25432), .dout(n25508));
  jor  g07486(.dina(n25508), .dinb(n25506), .dout(n25509));
  jand g07487(.dina(n25509), .dinb(n2714), .dout(n25510));
  jnot g07488(.din(n25510), .dout(n25511));
  jand g07489(.dina(n25433), .dinb(n25231), .dout(n25512));
  jxor g07490(.dina(n25389), .dinb(n25388), .dout(n25513));
  jand g07491(.dina(n25513), .dinb(n25432), .dout(n25514));
  jor  g07492(.dina(n25514), .dinb(n25512), .dout(n25515));
  jand g07493(.dina(n25515), .dinb(n2547), .dout(n25516));
  jnot g07494(.din(n25516), .dout(n25517));
  jand g07495(.dina(n25433), .dinb(n25236), .dout(n25518));
  jxor g07496(.dina(n25386), .dinb(n25385), .dout(n25519));
  jand g07497(.dina(n25519), .dinb(n25432), .dout(n25520));
  jor  g07498(.dina(n25520), .dinb(n25518), .dout(n25521));
  jand g07499(.dina(n25521), .dinb(n417), .dout(n25522));
  jnot g07500(.din(n25522), .dout(n25523));
  jand g07501(.dina(n25433), .dinb(n25241), .dout(n25524));
  jxor g07502(.dina(n25383), .dinb(n25382), .dout(n25525));
  jand g07503(.dina(n25525), .dinb(n25432), .dout(n25526));
  jor  g07504(.dina(n25526), .dinb(n25524), .dout(n25527));
  jand g07505(.dina(n25527), .dinb(n416), .dout(n25528));
  jnot g07506(.din(n25528), .dout(n25529));
  jand g07507(.dina(n25433), .dinb(n25246), .dout(n25530));
  jxor g07508(.dina(n25380), .dinb(n25379), .dout(n25531));
  jand g07509(.dina(n25531), .dinb(n25432), .dout(n25532));
  jor  g07510(.dina(n25532), .dinb(n25530), .dout(n25533));
  jand g07511(.dina(n25533), .dinb(n422), .dout(n25534));
  jnot g07512(.din(n25534), .dout(n25535));
  jand g07513(.dina(n25433), .dinb(n25251), .dout(n25536));
  jxor g07514(.dina(n25377), .dinb(n25376), .dout(n25537));
  jand g07515(.dina(n25537), .dinb(n25432), .dout(n25538));
  jor  g07516(.dina(n25538), .dinb(n25536), .dout(n25539));
  jand g07517(.dina(n25539), .dinb(n421), .dout(n25540));
  jnot g07518(.din(n25540), .dout(n25541));
  jand g07519(.dina(n25433), .dinb(n25256), .dout(n25542));
  jxor g07520(.dina(n25374), .dinb(n25373), .dout(n25543));
  jand g07521(.dina(n25543), .dinb(n25432), .dout(n25544));
  jor  g07522(.dina(n25544), .dinb(n25542), .dout(n25545));
  jand g07523(.dina(n25545), .dinb(n433), .dout(n25546));
  jnot g07524(.din(n25546), .dout(n25547));
  jand g07525(.dina(n25433), .dinb(n25261), .dout(n25548));
  jxor g07526(.dina(n25371), .dinb(n25370), .dout(n25549));
  jand g07527(.dina(n25549), .dinb(n25432), .dout(n25550));
  jor  g07528(.dina(n25550), .dinb(n25548), .dout(n25551));
  jand g07529(.dina(n25551), .dinb(n432), .dout(n25552));
  jnot g07530(.din(n25552), .dout(n25553));
  jand g07531(.dina(n25433), .dinb(n25266), .dout(n25554));
  jxor g07532(.dina(n25368), .dinb(n25367), .dout(n25555));
  jand g07533(.dina(n25555), .dinb(n25432), .dout(n25556));
  jor  g07534(.dina(n25556), .dinb(n25554), .dout(n25557));
  jand g07535(.dina(n25557), .dinb(n436), .dout(n25558));
  jnot g07536(.din(n25558), .dout(n25559));
  jand g07537(.dina(n25433), .dinb(n25271), .dout(n25560));
  jxor g07538(.dina(n25365), .dinb(n25364), .dout(n25561));
  jand g07539(.dina(n25561), .dinb(n25432), .dout(n25562));
  jor  g07540(.dina(n25562), .dinb(n25560), .dout(n25563));
  jand g07541(.dina(n25563), .dinb(n435), .dout(n25564));
  jnot g07542(.din(n25564), .dout(n25565));
  jand g07543(.dina(n25433), .dinb(n25276), .dout(n25566));
  jxor g07544(.dina(n25362), .dinb(n25361), .dout(n25567));
  jand g07545(.dina(n25567), .dinb(n25432), .dout(n25568));
  jor  g07546(.dina(n25568), .dinb(n25566), .dout(n25569));
  jand g07547(.dina(n25569), .dinb(n440), .dout(n25570));
  jnot g07548(.din(n25570), .dout(n25571));
  jand g07549(.dina(n25433), .dinb(n25281), .dout(n25572));
  jxor g07550(.dina(n25359), .dinb(n25358), .dout(n25573));
  jand g07551(.dina(n25573), .dinb(n25432), .dout(n25574));
  jor  g07552(.dina(n25574), .dinb(n25572), .dout(n25575));
  jand g07553(.dina(n25575), .dinb(n439), .dout(n25576));
  jnot g07554(.din(n25576), .dout(n25577));
  jand g07555(.dina(n25433), .dinb(n25286), .dout(n25578));
  jxor g07556(.dina(n25356), .dinb(n25355), .dout(n25579));
  jand g07557(.dina(n25579), .dinb(n25432), .dout(n25580));
  jor  g07558(.dina(n25580), .dinb(n25578), .dout(n25581));
  jand g07559(.dina(n25581), .dinb(n325), .dout(n25582));
  jnot g07560(.din(n25582), .dout(n25583));
  jand g07561(.dina(n25433), .dinb(n25291), .dout(n25584));
  jxor g07562(.dina(n25353), .dinb(n25352), .dout(n25585));
  jand g07563(.dina(n25585), .dinb(n25432), .dout(n25586));
  jor  g07564(.dina(n25586), .dinb(n25584), .dout(n25587));
  jand g07565(.dina(n25587), .dinb(n324), .dout(n25588));
  jnot g07566(.din(n25588), .dout(n25589));
  jand g07567(.dina(n25433), .dinb(n25296), .dout(n25590));
  jxor g07568(.dina(n25350), .dinb(n25349), .dout(n25591));
  jand g07569(.dina(n25591), .dinb(n25432), .dout(n25592));
  jor  g07570(.dina(n25592), .dinb(n25590), .dout(n25593));
  jand g07571(.dina(n25593), .dinb(n323), .dout(n25594));
  jnot g07572(.din(n25594), .dout(n25595));
  jand g07573(.dina(n25433), .dinb(n25301), .dout(n25596));
  jxor g07574(.dina(n25347), .dinb(n25346), .dout(n25597));
  jand g07575(.dina(n25597), .dinb(n25432), .dout(n25598));
  jor  g07576(.dina(n25598), .dinb(n25596), .dout(n25599));
  jand g07577(.dina(n25599), .dinb(n335), .dout(n25600));
  jnot g07578(.din(n25600), .dout(n25601));
  jand g07579(.dina(n25433), .dinb(n25306), .dout(n25602));
  jxor g07580(.dina(n25344), .dinb(n25343), .dout(n25603));
  jand g07581(.dina(n25603), .dinb(n25432), .dout(n25604));
  jor  g07582(.dina(n25604), .dinb(n25602), .dout(n25605));
  jand g07583(.dina(n25605), .dinb(n334), .dout(n25606));
  jnot g07584(.din(n25606), .dout(n25607));
  jand g07585(.dina(n25433), .dinb(n25311), .dout(n25608));
  jxor g07586(.dina(n25341), .dinb(n25340), .dout(n25609));
  jand g07587(.dina(n25609), .dinb(n25432), .dout(n25610));
  jor  g07588(.dina(n25610), .dinb(n25608), .dout(n25611));
  jand g07589(.dina(n25611), .dinb(n338), .dout(n25612));
  jnot g07590(.din(n25612), .dout(n25613));
  jand g07591(.dina(n25433), .dinb(n25316), .dout(n25614));
  jxor g07592(.dina(n25338), .dinb(n25337), .dout(n25615));
  jand g07593(.dina(n25615), .dinb(n25432), .dout(n25616));
  jor  g07594(.dina(n25616), .dinb(n25614), .dout(n25617));
  jand g07595(.dina(n25617), .dinb(n337), .dout(n25618));
  jnot g07596(.din(n25618), .dout(n25619));
  jnot g07597(.din(n25321), .dout(n25620));
  jor  g07598(.dina(n25432), .dinb(n25620), .dout(n25621));
  jxor g07599(.dina(n25335), .dinb(n25334), .dout(n25622));
  jnot g07600(.din(n25622), .dout(n25623));
  jor  g07601(.dina(n25623), .dinb(n25433), .dout(n25624));
  jand g07602(.dina(n25624), .dinb(n25621), .dout(n25625));
  jor  g07603(.dina(n25625), .dinb(b3 ), .dout(n25626));
  jor  g07604(.dina(n25432), .dinb(n25331), .dout(n25627));
  jxor g07605(.dina(n25332), .dinb(n5593), .dout(n25628));
  jand g07606(.dina(n25628), .dinb(n25432), .dout(n25629));
  jnot g07607(.din(n25629), .dout(n25630));
  jand g07608(.dina(n25630), .dinb(n25627), .dout(n25631));
  jor  g07609(.dina(n25631), .dinb(b2 ), .dout(n25632));
  jand g07610(.dina(n25431), .dinb(n5900), .dout(n25633));
  jor  g07611(.dina(n25633), .dinb(n5591), .dout(n25634));
  jnot g07612(.din(n5903), .dout(n25635));
  jnot g07613(.din(n25165), .dout(n25636));
  jnot g07614(.din(n25172), .dout(n25637));
  jnot g07615(.din(n25177), .dout(n25638));
  jnot g07616(.din(n25182), .dout(n25639));
  jnot g07617(.din(n25187), .dout(n25640));
  jnot g07618(.din(n25192), .dout(n25641));
  jnot g07619(.din(n25197), .dout(n25642));
  jnot g07620(.din(n25202), .dout(n25643));
  jnot g07621(.din(n25207), .dout(n25644));
  jnot g07622(.din(n25212), .dout(n25645));
  jnot g07623(.din(n25217), .dout(n25646));
  jnot g07624(.din(n25222), .dout(n25647));
  jnot g07625(.din(n25227), .dout(n25648));
  jnot g07626(.din(n25232), .dout(n25649));
  jnot g07627(.din(n25237), .dout(n25650));
  jnot g07628(.din(n25242), .dout(n25651));
  jnot g07629(.din(n25247), .dout(n25652));
  jnot g07630(.din(n25252), .dout(n25653));
  jnot g07631(.din(n25257), .dout(n25654));
  jnot g07632(.din(n25262), .dout(n25655));
  jnot g07633(.din(n25267), .dout(n25656));
  jnot g07634(.din(n25272), .dout(n25657));
  jnot g07635(.din(n25277), .dout(n25658));
  jnot g07636(.din(n25282), .dout(n25659));
  jnot g07637(.din(n25287), .dout(n25660));
  jnot g07638(.din(n25292), .dout(n25661));
  jnot g07639(.din(n25297), .dout(n25662));
  jnot g07640(.din(n25302), .dout(n25663));
  jnot g07641(.din(n25307), .dout(n25664));
  jnot g07642(.din(n25312), .dout(n25665));
  jnot g07643(.din(n25317), .dout(n25666));
  jnot g07644(.din(n25322), .dout(n25667));
  jnot g07645(.din(n25328), .dout(n25668));
  jxor g07646(.dina(n25331), .dinb(n258), .dout(n25669));
  jor  g07647(.dina(n25669), .dinb(n5592), .dout(n25670));
  jand g07648(.dina(n25670), .dinb(n25668), .dout(n25671));
  jnot g07649(.din(n25335), .dout(n25672));
  jor  g07650(.dina(n25672), .dinb(n25671), .dout(n25673));
  jand g07651(.dina(n25673), .dinb(n25667), .dout(n25674));
  jnot g07652(.din(n25338), .dout(n25675));
  jor  g07653(.dina(n25675), .dinb(n25674), .dout(n25676));
  jand g07654(.dina(n25676), .dinb(n25666), .dout(n25677));
  jnot g07655(.din(n25341), .dout(n25678));
  jor  g07656(.dina(n25678), .dinb(n25677), .dout(n25679));
  jand g07657(.dina(n25679), .dinb(n25665), .dout(n25680));
  jnot g07658(.din(n25344), .dout(n25681));
  jor  g07659(.dina(n25681), .dinb(n25680), .dout(n25682));
  jand g07660(.dina(n25682), .dinb(n25664), .dout(n25683));
  jnot g07661(.din(n25347), .dout(n25684));
  jor  g07662(.dina(n25684), .dinb(n25683), .dout(n25685));
  jand g07663(.dina(n25685), .dinb(n25663), .dout(n25686));
  jnot g07664(.din(n25350), .dout(n25687));
  jor  g07665(.dina(n25687), .dinb(n25686), .dout(n25688));
  jand g07666(.dina(n25688), .dinb(n25662), .dout(n25689));
  jnot g07667(.din(n25353), .dout(n25690));
  jor  g07668(.dina(n25690), .dinb(n25689), .dout(n25691));
  jand g07669(.dina(n25691), .dinb(n25661), .dout(n25692));
  jnot g07670(.din(n25356), .dout(n25693));
  jor  g07671(.dina(n25693), .dinb(n25692), .dout(n25694));
  jand g07672(.dina(n25694), .dinb(n25660), .dout(n25695));
  jnot g07673(.din(n25359), .dout(n25696));
  jor  g07674(.dina(n25696), .dinb(n25695), .dout(n25697));
  jand g07675(.dina(n25697), .dinb(n25659), .dout(n25698));
  jnot g07676(.din(n25362), .dout(n25699));
  jor  g07677(.dina(n25699), .dinb(n25698), .dout(n25700));
  jand g07678(.dina(n25700), .dinb(n25658), .dout(n25701));
  jnot g07679(.din(n25365), .dout(n25702));
  jor  g07680(.dina(n25702), .dinb(n25701), .dout(n25703));
  jand g07681(.dina(n25703), .dinb(n25657), .dout(n25704));
  jnot g07682(.din(n25368), .dout(n25705));
  jor  g07683(.dina(n25705), .dinb(n25704), .dout(n25706));
  jand g07684(.dina(n25706), .dinb(n25656), .dout(n25707));
  jnot g07685(.din(n25371), .dout(n25708));
  jor  g07686(.dina(n25708), .dinb(n25707), .dout(n25709));
  jand g07687(.dina(n25709), .dinb(n25655), .dout(n25710));
  jnot g07688(.din(n25374), .dout(n25711));
  jor  g07689(.dina(n25711), .dinb(n25710), .dout(n25712));
  jand g07690(.dina(n25712), .dinb(n25654), .dout(n25713));
  jnot g07691(.din(n25377), .dout(n25714));
  jor  g07692(.dina(n25714), .dinb(n25713), .dout(n25715));
  jand g07693(.dina(n25715), .dinb(n25653), .dout(n25716));
  jnot g07694(.din(n25380), .dout(n25717));
  jor  g07695(.dina(n25717), .dinb(n25716), .dout(n25718));
  jand g07696(.dina(n25718), .dinb(n25652), .dout(n25719));
  jnot g07697(.din(n25383), .dout(n25720));
  jor  g07698(.dina(n25720), .dinb(n25719), .dout(n25721));
  jand g07699(.dina(n25721), .dinb(n25651), .dout(n25722));
  jnot g07700(.din(n25386), .dout(n25723));
  jor  g07701(.dina(n25723), .dinb(n25722), .dout(n25724));
  jand g07702(.dina(n25724), .dinb(n25650), .dout(n25725));
  jnot g07703(.din(n25389), .dout(n25726));
  jor  g07704(.dina(n25726), .dinb(n25725), .dout(n25727));
  jand g07705(.dina(n25727), .dinb(n25649), .dout(n25728));
  jnot g07706(.din(n25392), .dout(n25729));
  jor  g07707(.dina(n25729), .dinb(n25728), .dout(n25730));
  jand g07708(.dina(n25730), .dinb(n25648), .dout(n25731));
  jnot g07709(.din(n25395), .dout(n25732));
  jor  g07710(.dina(n25732), .dinb(n25731), .dout(n25733));
  jand g07711(.dina(n25733), .dinb(n25647), .dout(n25734));
  jnot g07712(.din(n25398), .dout(n25735));
  jor  g07713(.dina(n25735), .dinb(n25734), .dout(n25736));
  jand g07714(.dina(n25736), .dinb(n25646), .dout(n25737));
  jnot g07715(.din(n25401), .dout(n25738));
  jor  g07716(.dina(n25738), .dinb(n25737), .dout(n25739));
  jand g07717(.dina(n25739), .dinb(n25645), .dout(n25740));
  jnot g07718(.din(n25404), .dout(n25741));
  jor  g07719(.dina(n25741), .dinb(n25740), .dout(n25742));
  jand g07720(.dina(n25742), .dinb(n25644), .dout(n25743));
  jnot g07721(.din(n25407), .dout(n25744));
  jor  g07722(.dina(n25744), .dinb(n25743), .dout(n25745));
  jand g07723(.dina(n25745), .dinb(n25643), .dout(n25746));
  jnot g07724(.din(n25410), .dout(n25747));
  jor  g07725(.dina(n25747), .dinb(n25746), .dout(n25748));
  jand g07726(.dina(n25748), .dinb(n25642), .dout(n25749));
  jnot g07727(.din(n25413), .dout(n25750));
  jor  g07728(.dina(n25750), .dinb(n25749), .dout(n25751));
  jand g07729(.dina(n25751), .dinb(n25641), .dout(n25752));
  jnot g07730(.din(n25416), .dout(n25753));
  jor  g07731(.dina(n25753), .dinb(n25752), .dout(n25754));
  jand g07732(.dina(n25754), .dinb(n25640), .dout(n25755));
  jnot g07733(.din(n25419), .dout(n25756));
  jor  g07734(.dina(n25756), .dinb(n25755), .dout(n25757));
  jand g07735(.dina(n25757), .dinb(n25639), .dout(n25758));
  jnot g07736(.din(n25422), .dout(n25759));
  jor  g07737(.dina(n25759), .dinb(n25758), .dout(n25760));
  jand g07738(.dina(n25760), .dinb(n25638), .dout(n25761));
  jnot g07739(.din(n25425), .dout(n25762));
  jor  g07740(.dina(n25762), .dinb(n25761), .dout(n25763));
  jand g07741(.dina(n25763), .dinb(n25637), .dout(n25764));
  jor  g07742(.dina(n25428), .dinb(n25764), .dout(n25765));
  jand g07743(.dina(n25765), .dinb(n25636), .dout(n25766));
  jor  g07744(.dina(n25766), .dinb(n25635), .dout(n25767));
  jand g07745(.dina(n25767), .dinb(n25634), .dout(n25768));
  jor  g07746(.dina(n25768), .dinb(b1 ), .dout(n25769));
  jxor g07747(.dina(n25768), .dinb(n258), .dout(n25770));
  jor  g07748(.dina(n25770), .dinb(n5909), .dout(n25771));
  jand g07749(.dina(n25771), .dinb(n25769), .dout(n25772));
  jxor g07750(.dina(n25631), .dinb(n348), .dout(n25773));
  jor  g07751(.dina(n25773), .dinb(n25772), .dout(n25774));
  jand g07752(.dina(n25774), .dinb(n25632), .dout(n25775));
  jxor g07753(.dina(n25625), .dinb(b3 ), .dout(n25776));
  jnot g07754(.din(n25776), .dout(n25777));
  jor  g07755(.dina(n25777), .dinb(n25775), .dout(n25778));
  jand g07756(.dina(n25778), .dinb(n25626), .dout(n25779));
  jxor g07757(.dina(n25617), .dinb(n337), .dout(n25780));
  jnot g07758(.din(n25780), .dout(n25781));
  jor  g07759(.dina(n25781), .dinb(n25779), .dout(n25782));
  jand g07760(.dina(n25782), .dinb(n25619), .dout(n25783));
  jxor g07761(.dina(n25611), .dinb(n338), .dout(n25784));
  jnot g07762(.din(n25784), .dout(n25785));
  jor  g07763(.dina(n25785), .dinb(n25783), .dout(n25786));
  jand g07764(.dina(n25786), .dinb(n25613), .dout(n25787));
  jxor g07765(.dina(n25605), .dinb(n334), .dout(n25788));
  jnot g07766(.din(n25788), .dout(n25789));
  jor  g07767(.dina(n25789), .dinb(n25787), .dout(n25790));
  jand g07768(.dina(n25790), .dinb(n25607), .dout(n25791));
  jxor g07769(.dina(n25599), .dinb(n335), .dout(n25792));
  jnot g07770(.din(n25792), .dout(n25793));
  jor  g07771(.dina(n25793), .dinb(n25791), .dout(n25794));
  jand g07772(.dina(n25794), .dinb(n25601), .dout(n25795));
  jxor g07773(.dina(n25593), .dinb(n323), .dout(n25796));
  jnot g07774(.din(n25796), .dout(n25797));
  jor  g07775(.dina(n25797), .dinb(n25795), .dout(n25798));
  jand g07776(.dina(n25798), .dinb(n25595), .dout(n25799));
  jxor g07777(.dina(n25587), .dinb(n324), .dout(n25800));
  jnot g07778(.din(n25800), .dout(n25801));
  jor  g07779(.dina(n25801), .dinb(n25799), .dout(n25802));
  jand g07780(.dina(n25802), .dinb(n25589), .dout(n25803));
  jxor g07781(.dina(n25581), .dinb(n325), .dout(n25804));
  jnot g07782(.din(n25804), .dout(n25805));
  jor  g07783(.dina(n25805), .dinb(n25803), .dout(n25806));
  jand g07784(.dina(n25806), .dinb(n25583), .dout(n25807));
  jxor g07785(.dina(n25575), .dinb(n439), .dout(n25808));
  jnot g07786(.din(n25808), .dout(n25809));
  jor  g07787(.dina(n25809), .dinb(n25807), .dout(n25810));
  jand g07788(.dina(n25810), .dinb(n25577), .dout(n25811));
  jxor g07789(.dina(n25569), .dinb(n440), .dout(n25812));
  jnot g07790(.din(n25812), .dout(n25813));
  jor  g07791(.dina(n25813), .dinb(n25811), .dout(n25814));
  jand g07792(.dina(n25814), .dinb(n25571), .dout(n25815));
  jxor g07793(.dina(n25563), .dinb(n435), .dout(n25816));
  jnot g07794(.din(n25816), .dout(n25817));
  jor  g07795(.dina(n25817), .dinb(n25815), .dout(n25818));
  jand g07796(.dina(n25818), .dinb(n25565), .dout(n25819));
  jxor g07797(.dina(n25557), .dinb(n436), .dout(n25820));
  jnot g07798(.din(n25820), .dout(n25821));
  jor  g07799(.dina(n25821), .dinb(n25819), .dout(n25822));
  jand g07800(.dina(n25822), .dinb(n25559), .dout(n25823));
  jxor g07801(.dina(n25551), .dinb(n432), .dout(n25824));
  jnot g07802(.din(n25824), .dout(n25825));
  jor  g07803(.dina(n25825), .dinb(n25823), .dout(n25826));
  jand g07804(.dina(n25826), .dinb(n25553), .dout(n25827));
  jxor g07805(.dina(n25545), .dinb(n433), .dout(n25828));
  jnot g07806(.din(n25828), .dout(n25829));
  jor  g07807(.dina(n25829), .dinb(n25827), .dout(n25830));
  jand g07808(.dina(n25830), .dinb(n25547), .dout(n25831));
  jxor g07809(.dina(n25539), .dinb(n421), .dout(n25832));
  jnot g07810(.din(n25832), .dout(n25833));
  jor  g07811(.dina(n25833), .dinb(n25831), .dout(n25834));
  jand g07812(.dina(n25834), .dinb(n25541), .dout(n25835));
  jxor g07813(.dina(n25533), .dinb(n422), .dout(n25836));
  jnot g07814(.din(n25836), .dout(n25837));
  jor  g07815(.dina(n25837), .dinb(n25835), .dout(n25838));
  jand g07816(.dina(n25838), .dinb(n25535), .dout(n25839));
  jxor g07817(.dina(n25527), .dinb(n416), .dout(n25840));
  jnot g07818(.din(n25840), .dout(n25841));
  jor  g07819(.dina(n25841), .dinb(n25839), .dout(n25842));
  jand g07820(.dina(n25842), .dinb(n25529), .dout(n25843));
  jxor g07821(.dina(n25521), .dinb(n417), .dout(n25844));
  jnot g07822(.din(n25844), .dout(n25845));
  jor  g07823(.dina(n25845), .dinb(n25843), .dout(n25846));
  jand g07824(.dina(n25846), .dinb(n25523), .dout(n25847));
  jxor g07825(.dina(n25515), .dinb(n2547), .dout(n25848));
  jnot g07826(.din(n25848), .dout(n25849));
  jor  g07827(.dina(n25849), .dinb(n25847), .dout(n25850));
  jand g07828(.dina(n25850), .dinb(n25517), .dout(n25851));
  jxor g07829(.dina(n25509), .dinb(n2714), .dout(n25852));
  jnot g07830(.din(n25852), .dout(n25853));
  jor  g07831(.dina(n25853), .dinb(n25851), .dout(n25854));
  jand g07832(.dina(n25854), .dinb(n25511), .dout(n25855));
  jxor g07833(.dina(n25503), .dinb(n405), .dout(n25856));
  jnot g07834(.din(n25856), .dout(n25857));
  jor  g07835(.dina(n25857), .dinb(n25855), .dout(n25858));
  jand g07836(.dina(n25858), .dinb(n25505), .dout(n25859));
  jxor g07837(.dina(n25497), .dinb(n406), .dout(n25860));
  jnot g07838(.din(n25860), .dout(n25861));
  jor  g07839(.dina(n25861), .dinb(n25859), .dout(n25862));
  jand g07840(.dina(n25862), .dinb(n25499), .dout(n25863));
  jxor g07841(.dina(n25491), .dinb(n412), .dout(n25864));
  jnot g07842(.din(n25864), .dout(n25865));
  jor  g07843(.dina(n25865), .dinb(n25863), .dout(n25866));
  jand g07844(.dina(n25866), .dinb(n25493), .dout(n25867));
  jxor g07845(.dina(n25485), .dinb(n413), .dout(n25868));
  jnot g07846(.din(n25868), .dout(n25869));
  jor  g07847(.dina(n25869), .dinb(n25867), .dout(n25870));
  jand g07848(.dina(n25870), .dinb(n25487), .dout(n25871));
  jxor g07849(.dina(n25479), .dinb(n409), .dout(n25872));
  jnot g07850(.din(n25872), .dout(n25873));
  jor  g07851(.dina(n25873), .dinb(n25871), .dout(n25874));
  jand g07852(.dina(n25874), .dinb(n25481), .dout(n25875));
  jxor g07853(.dina(n25473), .dinb(n410), .dout(n25876));
  jnot g07854(.din(n25876), .dout(n25877));
  jor  g07855(.dina(n25877), .dinb(n25875), .dout(n25878));
  jand g07856(.dina(n25878), .dinb(n25475), .dout(n25879));
  jxor g07857(.dina(n25467), .dinb(n426), .dout(n25880));
  jnot g07858(.din(n25880), .dout(n25881));
  jor  g07859(.dina(n25881), .dinb(n25879), .dout(n25882));
  jand g07860(.dina(n25882), .dinb(n25469), .dout(n25883));
  jxor g07861(.dina(n25461), .dinb(n427), .dout(n25884));
  jnot g07862(.din(n25884), .dout(n25885));
  jor  g07863(.dina(n25885), .dinb(n25883), .dout(n25886));
  jand g07864(.dina(n25886), .dinb(n25463), .dout(n25887));
  jxor g07865(.dina(n25455), .dinb(n424), .dout(n25888));
  jnot g07866(.din(n25888), .dout(n25889));
  jor  g07867(.dina(n25889), .dinb(n25887), .dout(n25890));
  jand g07868(.dina(n25890), .dinb(n25457), .dout(n25891));
  jxor g07869(.dina(n25449), .dinb(n300), .dout(n25892));
  jnot g07870(.din(n25892), .dout(n25893));
  jor  g07871(.dina(n25893), .dinb(n25891), .dout(n25894));
  jand g07872(.dina(n25894), .dinb(n25451), .dout(n25895));
  jxor g07873(.dina(n25443), .dinb(n297), .dout(n25896));
  jnot g07874(.din(n25896), .dout(n25897));
  jor  g07875(.dina(n25897), .dinb(n25895), .dout(n25898));
  jand g07876(.dina(n25898), .dinb(n25445), .dout(n25899));
  jnot g07877(.din(n25437), .dout(n25900));
  jand g07878(.dina(n25900), .dinb(b34 ), .dout(n25901));
  jor  g07879(.dina(n25901), .dinb(n25899), .dout(n25902));
  jand g07880(.dina(n25902), .dinb(n25439), .dout(n25903));
  jor  g07881(.dina(n25903), .dinb(n5704), .dout(n25904));
  jand g07882(.dina(n25904), .dinb(n25437), .dout(n25905));
  jnot g07883(.din(n25626), .dout(n25906));
  jnot g07884(.din(n25632), .dout(n25907));
  jnot g07885(.din(n5900), .dout(n25908));
  jor  g07886(.dina(n25766), .dinb(n25908), .dout(n25909));
  jand g07887(.dina(n25909), .dinb(a30 ), .dout(n25910));
  jnot g07888(.din(n25767), .dout(n25911));
  jor  g07889(.dina(n25911), .dinb(n25910), .dout(n25912));
  jand g07890(.dina(n25912), .dinb(n258), .dout(n25913));
  jxor g07891(.dina(n25768), .dinb(b1 ), .dout(n25914));
  jand g07892(.dina(n25914), .dinb(n6049), .dout(n25915));
  jor  g07893(.dina(n25915), .dinb(n25913), .dout(n25916));
  jxor g07894(.dina(n25631), .dinb(b2 ), .dout(n25917));
  jand g07895(.dina(n25917), .dinb(n25916), .dout(n25918));
  jor  g07896(.dina(n25918), .dinb(n25907), .dout(n25919));
  jand g07897(.dina(n25776), .dinb(n25919), .dout(n25920));
  jor  g07898(.dina(n25920), .dinb(n25906), .dout(n25921));
  jand g07899(.dina(n25780), .dinb(n25921), .dout(n25922));
  jor  g07900(.dina(n25922), .dinb(n25618), .dout(n25923));
  jand g07901(.dina(n25784), .dinb(n25923), .dout(n25924));
  jor  g07902(.dina(n25924), .dinb(n25612), .dout(n25925));
  jand g07903(.dina(n25788), .dinb(n25925), .dout(n25926));
  jor  g07904(.dina(n25926), .dinb(n25606), .dout(n25927));
  jand g07905(.dina(n25792), .dinb(n25927), .dout(n25928));
  jor  g07906(.dina(n25928), .dinb(n25600), .dout(n25929));
  jand g07907(.dina(n25796), .dinb(n25929), .dout(n25930));
  jor  g07908(.dina(n25930), .dinb(n25594), .dout(n25931));
  jand g07909(.dina(n25800), .dinb(n25931), .dout(n25932));
  jor  g07910(.dina(n25932), .dinb(n25588), .dout(n25933));
  jand g07911(.dina(n25804), .dinb(n25933), .dout(n25934));
  jor  g07912(.dina(n25934), .dinb(n25582), .dout(n25935));
  jand g07913(.dina(n25808), .dinb(n25935), .dout(n25936));
  jor  g07914(.dina(n25936), .dinb(n25576), .dout(n25937));
  jand g07915(.dina(n25812), .dinb(n25937), .dout(n25938));
  jor  g07916(.dina(n25938), .dinb(n25570), .dout(n25939));
  jand g07917(.dina(n25816), .dinb(n25939), .dout(n25940));
  jor  g07918(.dina(n25940), .dinb(n25564), .dout(n25941));
  jand g07919(.dina(n25820), .dinb(n25941), .dout(n25942));
  jor  g07920(.dina(n25942), .dinb(n25558), .dout(n25943));
  jand g07921(.dina(n25824), .dinb(n25943), .dout(n25944));
  jor  g07922(.dina(n25944), .dinb(n25552), .dout(n25945));
  jand g07923(.dina(n25828), .dinb(n25945), .dout(n25946));
  jor  g07924(.dina(n25946), .dinb(n25546), .dout(n25947));
  jand g07925(.dina(n25832), .dinb(n25947), .dout(n25948));
  jor  g07926(.dina(n25948), .dinb(n25540), .dout(n25949));
  jand g07927(.dina(n25836), .dinb(n25949), .dout(n25950));
  jor  g07928(.dina(n25950), .dinb(n25534), .dout(n25951));
  jand g07929(.dina(n25840), .dinb(n25951), .dout(n25952));
  jor  g07930(.dina(n25952), .dinb(n25528), .dout(n25953));
  jand g07931(.dina(n25844), .dinb(n25953), .dout(n25954));
  jor  g07932(.dina(n25954), .dinb(n25522), .dout(n25955));
  jand g07933(.dina(n25848), .dinb(n25955), .dout(n25956));
  jor  g07934(.dina(n25956), .dinb(n25516), .dout(n25957));
  jand g07935(.dina(n25852), .dinb(n25957), .dout(n25958));
  jor  g07936(.dina(n25958), .dinb(n25510), .dout(n25959));
  jand g07937(.dina(n25856), .dinb(n25959), .dout(n25960));
  jor  g07938(.dina(n25960), .dinb(n25504), .dout(n25961));
  jand g07939(.dina(n25860), .dinb(n25961), .dout(n25962));
  jor  g07940(.dina(n25962), .dinb(n25498), .dout(n25963));
  jand g07941(.dina(n25864), .dinb(n25963), .dout(n25964));
  jor  g07942(.dina(n25964), .dinb(n25492), .dout(n25965));
  jand g07943(.dina(n25868), .dinb(n25965), .dout(n25966));
  jor  g07944(.dina(n25966), .dinb(n25486), .dout(n25967));
  jand g07945(.dina(n25872), .dinb(n25967), .dout(n25968));
  jor  g07946(.dina(n25968), .dinb(n25480), .dout(n25969));
  jand g07947(.dina(n25876), .dinb(n25969), .dout(n25970));
  jor  g07948(.dina(n25970), .dinb(n25474), .dout(n25971));
  jand g07949(.dina(n25880), .dinb(n25971), .dout(n25972));
  jor  g07950(.dina(n25972), .dinb(n25468), .dout(n25973));
  jand g07951(.dina(n25884), .dinb(n25973), .dout(n25974));
  jor  g07952(.dina(n25974), .dinb(n25462), .dout(n25975));
  jand g07953(.dina(n25888), .dinb(n25975), .dout(n25976));
  jor  g07954(.dina(n25976), .dinb(n25456), .dout(n25977));
  jand g07955(.dina(n25892), .dinb(n25977), .dout(n25978));
  jor  g07956(.dina(n25978), .dinb(n25450), .dout(n25979));
  jand g07957(.dina(n25896), .dinb(n25979), .dout(n25980));
  jor  g07958(.dina(n25980), .dinb(n25444), .dout(n25981));
  jand g07959(.dina(n25438), .dinb(n5703), .dout(n25982));
  jand g07960(.dina(n25982), .dinb(n25981), .dout(n25983));
  jor  g07961(.dina(n25983), .dinb(n25905), .dout(n25984));
  jnot g07962(.din(n25984), .dout(n25985));
  jand g07963(.dina(n25904), .dinb(n25443), .dout(n25986));
  jnot g07964(.din(n25901), .dout(n25987));
  jand g07965(.dina(n25987), .dinb(n25981), .dout(n25988));
  jor  g07966(.dina(n25988), .dinb(n25438), .dout(n25989));
  jand g07967(.dina(n25989), .dinb(n5703), .dout(n25990));
  jxor g07968(.dina(n25896), .dinb(n25979), .dout(n25991));
  jand g07969(.dina(n25991), .dinb(n25990), .dout(n25992));
  jor  g07970(.dina(n25992), .dinb(n25986), .dout(n25993));
  jand g07971(.dina(n25993), .dinb(n298), .dout(n25994));
  jnot g07972(.din(n25994), .dout(n25995));
  jand g07973(.dina(n25904), .dinb(n25449), .dout(n25996));
  jxor g07974(.dina(n25892), .dinb(n25977), .dout(n25997));
  jand g07975(.dina(n25997), .dinb(n25990), .dout(n25998));
  jor  g07976(.dina(n25998), .dinb(n25996), .dout(n25999));
  jand g07977(.dina(n25999), .dinb(n297), .dout(n26000));
  jnot g07978(.din(n26000), .dout(n26001));
  jand g07979(.dina(n25904), .dinb(n25455), .dout(n26002));
  jxor g07980(.dina(n25888), .dinb(n25975), .dout(n26003));
  jand g07981(.dina(n26003), .dinb(n25990), .dout(n26004));
  jor  g07982(.dina(n26004), .dinb(n26002), .dout(n26005));
  jand g07983(.dina(n26005), .dinb(n300), .dout(n26006));
  jnot g07984(.din(n26006), .dout(n26007));
  jand g07985(.dina(n25904), .dinb(n25461), .dout(n26008));
  jxor g07986(.dina(n25884), .dinb(n25973), .dout(n26009));
  jand g07987(.dina(n26009), .dinb(n25990), .dout(n26010));
  jor  g07988(.dina(n26010), .dinb(n26008), .dout(n26011));
  jand g07989(.dina(n26011), .dinb(n424), .dout(n26012));
  jnot g07990(.din(n26012), .dout(n26013));
  jand g07991(.dina(n25904), .dinb(n25467), .dout(n26014));
  jxor g07992(.dina(n25880), .dinb(n25971), .dout(n26015));
  jand g07993(.dina(n26015), .dinb(n25990), .dout(n26016));
  jor  g07994(.dina(n26016), .dinb(n26014), .dout(n26017));
  jand g07995(.dina(n26017), .dinb(n427), .dout(n26018));
  jnot g07996(.din(n26018), .dout(n26019));
  jand g07997(.dina(n25904), .dinb(n25473), .dout(n26020));
  jxor g07998(.dina(n25876), .dinb(n25969), .dout(n26021));
  jand g07999(.dina(n26021), .dinb(n25990), .dout(n26022));
  jor  g08000(.dina(n26022), .dinb(n26020), .dout(n26023));
  jand g08001(.dina(n26023), .dinb(n426), .dout(n26024));
  jnot g08002(.din(n26024), .dout(n26025));
  jand g08003(.dina(n25904), .dinb(n25479), .dout(n26026));
  jxor g08004(.dina(n25872), .dinb(n25967), .dout(n26027));
  jand g08005(.dina(n26027), .dinb(n25990), .dout(n26028));
  jor  g08006(.dina(n26028), .dinb(n26026), .dout(n26029));
  jand g08007(.dina(n26029), .dinb(n410), .dout(n26030));
  jnot g08008(.din(n26030), .dout(n26031));
  jand g08009(.dina(n25904), .dinb(n25485), .dout(n26032));
  jxor g08010(.dina(n25868), .dinb(n25965), .dout(n26033));
  jand g08011(.dina(n26033), .dinb(n25990), .dout(n26034));
  jor  g08012(.dina(n26034), .dinb(n26032), .dout(n26035));
  jand g08013(.dina(n26035), .dinb(n409), .dout(n26036));
  jnot g08014(.din(n26036), .dout(n26037));
  jand g08015(.dina(n25904), .dinb(n25491), .dout(n26038));
  jxor g08016(.dina(n25864), .dinb(n25963), .dout(n26039));
  jand g08017(.dina(n26039), .dinb(n25990), .dout(n26040));
  jor  g08018(.dina(n26040), .dinb(n26038), .dout(n26041));
  jand g08019(.dina(n26041), .dinb(n413), .dout(n26042));
  jnot g08020(.din(n26042), .dout(n26043));
  jand g08021(.dina(n25904), .dinb(n25497), .dout(n26044));
  jxor g08022(.dina(n25860), .dinb(n25961), .dout(n26045));
  jand g08023(.dina(n26045), .dinb(n25990), .dout(n26046));
  jor  g08024(.dina(n26046), .dinb(n26044), .dout(n26047));
  jand g08025(.dina(n26047), .dinb(n412), .dout(n26048));
  jnot g08026(.din(n26048), .dout(n26049));
  jand g08027(.dina(n25904), .dinb(n25503), .dout(n26050));
  jxor g08028(.dina(n25856), .dinb(n25959), .dout(n26051));
  jand g08029(.dina(n26051), .dinb(n25990), .dout(n26052));
  jor  g08030(.dina(n26052), .dinb(n26050), .dout(n26053));
  jand g08031(.dina(n26053), .dinb(n406), .dout(n26054));
  jnot g08032(.din(n26054), .dout(n26055));
  jand g08033(.dina(n25904), .dinb(n25509), .dout(n26056));
  jxor g08034(.dina(n25852), .dinb(n25957), .dout(n26057));
  jand g08035(.dina(n26057), .dinb(n25990), .dout(n26058));
  jor  g08036(.dina(n26058), .dinb(n26056), .dout(n26059));
  jand g08037(.dina(n26059), .dinb(n405), .dout(n26060));
  jnot g08038(.din(n26060), .dout(n26061));
  jand g08039(.dina(n25904), .dinb(n25515), .dout(n26062));
  jxor g08040(.dina(n25848), .dinb(n25955), .dout(n26063));
  jand g08041(.dina(n26063), .dinb(n25990), .dout(n26064));
  jor  g08042(.dina(n26064), .dinb(n26062), .dout(n26065));
  jand g08043(.dina(n26065), .dinb(n2714), .dout(n26066));
  jnot g08044(.din(n26066), .dout(n26067));
  jand g08045(.dina(n25904), .dinb(n25521), .dout(n26068));
  jxor g08046(.dina(n25844), .dinb(n25953), .dout(n26069));
  jand g08047(.dina(n26069), .dinb(n25990), .dout(n26070));
  jor  g08048(.dina(n26070), .dinb(n26068), .dout(n26071));
  jand g08049(.dina(n26071), .dinb(n2547), .dout(n26072));
  jnot g08050(.din(n26072), .dout(n26073));
  jand g08051(.dina(n25904), .dinb(n25527), .dout(n26074));
  jxor g08052(.dina(n25840), .dinb(n25951), .dout(n26075));
  jand g08053(.dina(n26075), .dinb(n25990), .dout(n26076));
  jor  g08054(.dina(n26076), .dinb(n26074), .dout(n26077));
  jand g08055(.dina(n26077), .dinb(n417), .dout(n26078));
  jnot g08056(.din(n26078), .dout(n26079));
  jand g08057(.dina(n25904), .dinb(n25533), .dout(n26080));
  jxor g08058(.dina(n25836), .dinb(n25949), .dout(n26081));
  jand g08059(.dina(n26081), .dinb(n25990), .dout(n26082));
  jor  g08060(.dina(n26082), .dinb(n26080), .dout(n26083));
  jand g08061(.dina(n26083), .dinb(n416), .dout(n26084));
  jnot g08062(.din(n26084), .dout(n26085));
  jand g08063(.dina(n25904), .dinb(n25539), .dout(n26086));
  jxor g08064(.dina(n25832), .dinb(n25947), .dout(n26087));
  jand g08065(.dina(n26087), .dinb(n25990), .dout(n26088));
  jor  g08066(.dina(n26088), .dinb(n26086), .dout(n26089));
  jand g08067(.dina(n26089), .dinb(n422), .dout(n26090));
  jnot g08068(.din(n26090), .dout(n26091));
  jand g08069(.dina(n25904), .dinb(n25545), .dout(n26092));
  jxor g08070(.dina(n25828), .dinb(n25945), .dout(n26093));
  jand g08071(.dina(n26093), .dinb(n25990), .dout(n26094));
  jor  g08072(.dina(n26094), .dinb(n26092), .dout(n26095));
  jand g08073(.dina(n26095), .dinb(n421), .dout(n26096));
  jnot g08074(.din(n26096), .dout(n26097));
  jand g08075(.dina(n25904), .dinb(n25551), .dout(n26098));
  jxor g08076(.dina(n25824), .dinb(n25943), .dout(n26099));
  jand g08077(.dina(n26099), .dinb(n25990), .dout(n26100));
  jor  g08078(.dina(n26100), .dinb(n26098), .dout(n26101));
  jand g08079(.dina(n26101), .dinb(n433), .dout(n26102));
  jnot g08080(.din(n26102), .dout(n26103));
  jand g08081(.dina(n25904), .dinb(n25557), .dout(n26104));
  jxor g08082(.dina(n25820), .dinb(n25941), .dout(n26105));
  jand g08083(.dina(n26105), .dinb(n25990), .dout(n26106));
  jor  g08084(.dina(n26106), .dinb(n26104), .dout(n26107));
  jand g08085(.dina(n26107), .dinb(n432), .dout(n26108));
  jnot g08086(.din(n26108), .dout(n26109));
  jand g08087(.dina(n25904), .dinb(n25563), .dout(n26110));
  jxor g08088(.dina(n25816), .dinb(n25939), .dout(n26111));
  jand g08089(.dina(n26111), .dinb(n25990), .dout(n26112));
  jor  g08090(.dina(n26112), .dinb(n26110), .dout(n26113));
  jand g08091(.dina(n26113), .dinb(n436), .dout(n26114));
  jnot g08092(.din(n26114), .dout(n26115));
  jand g08093(.dina(n25904), .dinb(n25569), .dout(n26116));
  jxor g08094(.dina(n25812), .dinb(n25937), .dout(n26117));
  jand g08095(.dina(n26117), .dinb(n25990), .dout(n26118));
  jor  g08096(.dina(n26118), .dinb(n26116), .dout(n26119));
  jand g08097(.dina(n26119), .dinb(n435), .dout(n26120));
  jnot g08098(.din(n26120), .dout(n26121));
  jand g08099(.dina(n25904), .dinb(n25575), .dout(n26122));
  jxor g08100(.dina(n25808), .dinb(n25935), .dout(n26123));
  jand g08101(.dina(n26123), .dinb(n25990), .dout(n26124));
  jor  g08102(.dina(n26124), .dinb(n26122), .dout(n26125));
  jand g08103(.dina(n26125), .dinb(n440), .dout(n26126));
  jnot g08104(.din(n26126), .dout(n26127));
  jand g08105(.dina(n25904), .dinb(n25581), .dout(n26128));
  jxor g08106(.dina(n25804), .dinb(n25933), .dout(n26129));
  jand g08107(.dina(n26129), .dinb(n25990), .dout(n26130));
  jor  g08108(.dina(n26130), .dinb(n26128), .dout(n26131));
  jand g08109(.dina(n26131), .dinb(n439), .dout(n26132));
  jnot g08110(.din(n26132), .dout(n26133));
  jand g08111(.dina(n25904), .dinb(n25587), .dout(n26134));
  jxor g08112(.dina(n25800), .dinb(n25931), .dout(n26135));
  jand g08113(.dina(n26135), .dinb(n25990), .dout(n26136));
  jor  g08114(.dina(n26136), .dinb(n26134), .dout(n26137));
  jand g08115(.dina(n26137), .dinb(n325), .dout(n26138));
  jnot g08116(.din(n26138), .dout(n26139));
  jand g08117(.dina(n25904), .dinb(n25593), .dout(n26140));
  jxor g08118(.dina(n25796), .dinb(n25929), .dout(n26141));
  jand g08119(.dina(n26141), .dinb(n25990), .dout(n26142));
  jor  g08120(.dina(n26142), .dinb(n26140), .dout(n26143));
  jand g08121(.dina(n26143), .dinb(n324), .dout(n26144));
  jnot g08122(.din(n26144), .dout(n26145));
  jand g08123(.dina(n25904), .dinb(n25599), .dout(n26146));
  jxor g08124(.dina(n25792), .dinb(n25927), .dout(n26147));
  jand g08125(.dina(n26147), .dinb(n25990), .dout(n26148));
  jor  g08126(.dina(n26148), .dinb(n26146), .dout(n26149));
  jand g08127(.dina(n26149), .dinb(n323), .dout(n26150));
  jnot g08128(.din(n26150), .dout(n26151));
  jand g08129(.dina(n25904), .dinb(n25605), .dout(n26152));
  jxor g08130(.dina(n25788), .dinb(n25925), .dout(n26153));
  jand g08131(.dina(n26153), .dinb(n25990), .dout(n26154));
  jor  g08132(.dina(n26154), .dinb(n26152), .dout(n26155));
  jand g08133(.dina(n26155), .dinb(n335), .dout(n26156));
  jnot g08134(.din(n26156), .dout(n26157));
  jand g08135(.dina(n25904), .dinb(n25611), .dout(n26158));
  jxor g08136(.dina(n25784), .dinb(n25923), .dout(n26159));
  jand g08137(.dina(n26159), .dinb(n25990), .dout(n26160));
  jor  g08138(.dina(n26160), .dinb(n26158), .dout(n26161));
  jand g08139(.dina(n26161), .dinb(n334), .dout(n26162));
  jnot g08140(.din(n26162), .dout(n26163));
  jand g08141(.dina(n25904), .dinb(n25617), .dout(n26164));
  jxor g08142(.dina(n25780), .dinb(n25921), .dout(n26165));
  jand g08143(.dina(n26165), .dinb(n25990), .dout(n26166));
  jor  g08144(.dina(n26166), .dinb(n26164), .dout(n26167));
  jand g08145(.dina(n26167), .dinb(n338), .dout(n26168));
  jnot g08146(.din(n26168), .dout(n26169));
  jor  g08147(.dina(n25990), .dinb(n25625), .dout(n26170));
  jxor g08148(.dina(n25776), .dinb(n25919), .dout(n26171));
  jand g08149(.dina(n26171), .dinb(n25990), .dout(n26172));
  jnot g08150(.din(n26172), .dout(n26173));
  jand g08151(.dina(n26173), .dinb(n26170), .dout(n26174));
  jnot g08152(.din(n26174), .dout(n26175));
  jand g08153(.dina(n26175), .dinb(n337), .dout(n26176));
  jnot g08154(.din(n26176), .dout(n26177));
  jor  g08155(.dina(n25990), .dinb(n25631), .dout(n26178));
  jxor g08156(.dina(n25917), .dinb(n25916), .dout(n26179));
  jnot g08157(.din(n26179), .dout(n26180));
  jor  g08158(.dina(n26180), .dinb(n25904), .dout(n26181));
  jand g08159(.dina(n26181), .dinb(n26178), .dout(n26182));
  jnot g08160(.din(n26182), .dout(n26183));
  jand g08161(.dina(n26183), .dinb(n344), .dout(n26184));
  jnot g08162(.din(n26184), .dout(n26185));
  jand g08163(.dina(n25904), .dinb(n25912), .dout(n26186));
  jxor g08164(.dina(n25914), .dinb(n6049), .dout(n26187));
  jand g08165(.dina(n26187), .dinb(n25990), .dout(n26188));
  jor  g08166(.dina(n26188), .dinb(n26186), .dout(n26189));
  jand g08167(.dina(n26189), .dinb(n348), .dout(n26190));
  jnot g08168(.din(n26190), .dout(n26191));
  jnot g08169(.din(n6286), .dout(n26192));
  jor  g08170(.dina(n25903), .dinb(n26192), .dout(n26193));
  jand g08171(.dina(n26193), .dinb(a29 ), .dout(n26194));
  jand g08172(.dina(n25990), .dinb(n5909), .dout(n26195));
  jor  g08173(.dina(n26195), .dinb(n26194), .dout(n26196));
  jand g08174(.dina(n26196), .dinb(n258), .dout(n26197));
  jnot g08175(.din(n26197), .dout(n26198));
  jand g08176(.dina(n25989), .dinb(n6286), .dout(n26199));
  jor  g08177(.dina(n26199), .dinb(n5908), .dout(n26200));
  jor  g08178(.dina(n25904), .dinb(n6049), .dout(n26201));
  jand g08179(.dina(n26201), .dinb(n26200), .dout(n26202));
  jxor g08180(.dina(n26202), .dinb(n258), .dout(n26203));
  jor  g08181(.dina(n26203), .dinb(n6294), .dout(n26204));
  jand g08182(.dina(n26204), .dinb(n26198), .dout(n26205));
  jxor g08183(.dina(n26189), .dinb(n348), .dout(n26206));
  jnot g08184(.din(n26206), .dout(n26207));
  jor  g08185(.dina(n26207), .dinb(n26205), .dout(n26208));
  jand g08186(.dina(n26208), .dinb(n26191), .dout(n26209));
  jxor g08187(.dina(n26182), .dinb(b3 ), .dout(n26210));
  jnot g08188(.din(n26210), .dout(n26211));
  jor  g08189(.dina(n26211), .dinb(n26209), .dout(n26212));
  jand g08190(.dina(n26212), .dinb(n26185), .dout(n26213));
  jxor g08191(.dina(n26174), .dinb(b4 ), .dout(n26214));
  jnot g08192(.din(n26214), .dout(n26215));
  jor  g08193(.dina(n26215), .dinb(n26213), .dout(n26216));
  jand g08194(.dina(n26216), .dinb(n26177), .dout(n26217));
  jxor g08195(.dina(n26167), .dinb(n338), .dout(n26218));
  jnot g08196(.din(n26218), .dout(n26219));
  jor  g08197(.dina(n26219), .dinb(n26217), .dout(n26220));
  jand g08198(.dina(n26220), .dinb(n26169), .dout(n26221));
  jxor g08199(.dina(n26161), .dinb(n334), .dout(n26222));
  jnot g08200(.din(n26222), .dout(n26223));
  jor  g08201(.dina(n26223), .dinb(n26221), .dout(n26224));
  jand g08202(.dina(n26224), .dinb(n26163), .dout(n26225));
  jxor g08203(.dina(n26155), .dinb(n335), .dout(n26226));
  jnot g08204(.din(n26226), .dout(n26227));
  jor  g08205(.dina(n26227), .dinb(n26225), .dout(n26228));
  jand g08206(.dina(n26228), .dinb(n26157), .dout(n26229));
  jxor g08207(.dina(n26149), .dinb(n323), .dout(n26230));
  jnot g08208(.din(n26230), .dout(n26231));
  jor  g08209(.dina(n26231), .dinb(n26229), .dout(n26232));
  jand g08210(.dina(n26232), .dinb(n26151), .dout(n26233));
  jxor g08211(.dina(n26143), .dinb(n324), .dout(n26234));
  jnot g08212(.din(n26234), .dout(n26235));
  jor  g08213(.dina(n26235), .dinb(n26233), .dout(n26236));
  jand g08214(.dina(n26236), .dinb(n26145), .dout(n26237));
  jxor g08215(.dina(n26137), .dinb(n325), .dout(n26238));
  jnot g08216(.din(n26238), .dout(n26239));
  jor  g08217(.dina(n26239), .dinb(n26237), .dout(n26240));
  jand g08218(.dina(n26240), .dinb(n26139), .dout(n26241));
  jxor g08219(.dina(n26131), .dinb(n439), .dout(n26242));
  jnot g08220(.din(n26242), .dout(n26243));
  jor  g08221(.dina(n26243), .dinb(n26241), .dout(n26244));
  jand g08222(.dina(n26244), .dinb(n26133), .dout(n26245));
  jxor g08223(.dina(n26125), .dinb(n440), .dout(n26246));
  jnot g08224(.din(n26246), .dout(n26247));
  jor  g08225(.dina(n26247), .dinb(n26245), .dout(n26248));
  jand g08226(.dina(n26248), .dinb(n26127), .dout(n26249));
  jxor g08227(.dina(n26119), .dinb(n435), .dout(n26250));
  jnot g08228(.din(n26250), .dout(n26251));
  jor  g08229(.dina(n26251), .dinb(n26249), .dout(n26252));
  jand g08230(.dina(n26252), .dinb(n26121), .dout(n26253));
  jxor g08231(.dina(n26113), .dinb(n436), .dout(n26254));
  jnot g08232(.din(n26254), .dout(n26255));
  jor  g08233(.dina(n26255), .dinb(n26253), .dout(n26256));
  jand g08234(.dina(n26256), .dinb(n26115), .dout(n26257));
  jxor g08235(.dina(n26107), .dinb(n432), .dout(n26258));
  jnot g08236(.din(n26258), .dout(n26259));
  jor  g08237(.dina(n26259), .dinb(n26257), .dout(n26260));
  jand g08238(.dina(n26260), .dinb(n26109), .dout(n26261));
  jxor g08239(.dina(n26101), .dinb(n433), .dout(n26262));
  jnot g08240(.din(n26262), .dout(n26263));
  jor  g08241(.dina(n26263), .dinb(n26261), .dout(n26264));
  jand g08242(.dina(n26264), .dinb(n26103), .dout(n26265));
  jxor g08243(.dina(n26095), .dinb(n421), .dout(n26266));
  jnot g08244(.din(n26266), .dout(n26267));
  jor  g08245(.dina(n26267), .dinb(n26265), .dout(n26268));
  jand g08246(.dina(n26268), .dinb(n26097), .dout(n26269));
  jxor g08247(.dina(n26089), .dinb(n422), .dout(n26270));
  jnot g08248(.din(n26270), .dout(n26271));
  jor  g08249(.dina(n26271), .dinb(n26269), .dout(n26272));
  jand g08250(.dina(n26272), .dinb(n26091), .dout(n26273));
  jxor g08251(.dina(n26083), .dinb(n416), .dout(n26274));
  jnot g08252(.din(n26274), .dout(n26275));
  jor  g08253(.dina(n26275), .dinb(n26273), .dout(n26276));
  jand g08254(.dina(n26276), .dinb(n26085), .dout(n26277));
  jxor g08255(.dina(n26077), .dinb(n417), .dout(n26278));
  jnot g08256(.din(n26278), .dout(n26279));
  jor  g08257(.dina(n26279), .dinb(n26277), .dout(n26280));
  jand g08258(.dina(n26280), .dinb(n26079), .dout(n26281));
  jxor g08259(.dina(n26071), .dinb(n2547), .dout(n26282));
  jnot g08260(.din(n26282), .dout(n26283));
  jor  g08261(.dina(n26283), .dinb(n26281), .dout(n26284));
  jand g08262(.dina(n26284), .dinb(n26073), .dout(n26285));
  jxor g08263(.dina(n26065), .dinb(n2714), .dout(n26286));
  jnot g08264(.din(n26286), .dout(n26287));
  jor  g08265(.dina(n26287), .dinb(n26285), .dout(n26288));
  jand g08266(.dina(n26288), .dinb(n26067), .dout(n26289));
  jxor g08267(.dina(n26059), .dinb(n405), .dout(n26290));
  jnot g08268(.din(n26290), .dout(n26291));
  jor  g08269(.dina(n26291), .dinb(n26289), .dout(n26292));
  jand g08270(.dina(n26292), .dinb(n26061), .dout(n26293));
  jxor g08271(.dina(n26053), .dinb(n406), .dout(n26294));
  jnot g08272(.din(n26294), .dout(n26295));
  jor  g08273(.dina(n26295), .dinb(n26293), .dout(n26296));
  jand g08274(.dina(n26296), .dinb(n26055), .dout(n26297));
  jxor g08275(.dina(n26047), .dinb(n412), .dout(n26298));
  jnot g08276(.din(n26298), .dout(n26299));
  jor  g08277(.dina(n26299), .dinb(n26297), .dout(n26300));
  jand g08278(.dina(n26300), .dinb(n26049), .dout(n26301));
  jxor g08279(.dina(n26041), .dinb(n413), .dout(n26302));
  jnot g08280(.din(n26302), .dout(n26303));
  jor  g08281(.dina(n26303), .dinb(n26301), .dout(n26304));
  jand g08282(.dina(n26304), .dinb(n26043), .dout(n26305));
  jxor g08283(.dina(n26035), .dinb(n409), .dout(n26306));
  jnot g08284(.din(n26306), .dout(n26307));
  jor  g08285(.dina(n26307), .dinb(n26305), .dout(n26308));
  jand g08286(.dina(n26308), .dinb(n26037), .dout(n26309));
  jxor g08287(.dina(n26029), .dinb(n410), .dout(n26310));
  jnot g08288(.din(n26310), .dout(n26311));
  jor  g08289(.dina(n26311), .dinb(n26309), .dout(n26312));
  jand g08290(.dina(n26312), .dinb(n26031), .dout(n26313));
  jxor g08291(.dina(n26023), .dinb(n426), .dout(n26314));
  jnot g08292(.din(n26314), .dout(n26315));
  jor  g08293(.dina(n26315), .dinb(n26313), .dout(n26316));
  jand g08294(.dina(n26316), .dinb(n26025), .dout(n26317));
  jxor g08295(.dina(n26017), .dinb(n427), .dout(n26318));
  jnot g08296(.din(n26318), .dout(n26319));
  jor  g08297(.dina(n26319), .dinb(n26317), .dout(n26320));
  jand g08298(.dina(n26320), .dinb(n26019), .dout(n26321));
  jxor g08299(.dina(n26011), .dinb(n424), .dout(n26322));
  jnot g08300(.din(n26322), .dout(n26323));
  jor  g08301(.dina(n26323), .dinb(n26321), .dout(n26324));
  jand g08302(.dina(n26324), .dinb(n26013), .dout(n26325));
  jxor g08303(.dina(n26005), .dinb(n300), .dout(n26326));
  jnot g08304(.din(n26326), .dout(n26327));
  jor  g08305(.dina(n26327), .dinb(n26325), .dout(n26328));
  jand g08306(.dina(n26328), .dinb(n26007), .dout(n26329));
  jxor g08307(.dina(n25999), .dinb(n297), .dout(n26330));
  jnot g08308(.din(n26330), .dout(n26331));
  jor  g08309(.dina(n26331), .dinb(n26329), .dout(n26332));
  jand g08310(.dina(n26332), .dinb(n26001), .dout(n26333));
  jxor g08311(.dina(n25993), .dinb(n298), .dout(n26334));
  jnot g08312(.din(n26334), .dout(n26335));
  jor  g08313(.dina(n26335), .dinb(n26333), .dout(n26336));
  jand g08314(.dina(n26336), .dinb(n25995), .dout(n26337));
  jxor g08315(.dina(n25984), .dinb(b35 ), .dout(n26338));
  jor  g08316(.dina(n26338), .dinb(n6404), .dout(n26339));
  jor  g08317(.dina(n26339), .dinb(n26337), .dout(n26340));
  jand g08318(.dina(n26340), .dinb(n25985), .dout(n26341));
  jxor g08319(.dina(n26202), .dinb(b1 ), .dout(n26342));
  jand g08320(.dina(n26342), .dinb(n6295), .dout(n26343));
  jor  g08321(.dina(n26343), .dinb(n26197), .dout(n26344));
  jand g08322(.dina(n26206), .dinb(n26344), .dout(n26345));
  jor  g08323(.dina(n26345), .dinb(n26190), .dout(n26346));
  jand g08324(.dina(n26210), .dinb(n26346), .dout(n26347));
  jor  g08325(.dina(n26347), .dinb(n26184), .dout(n26348));
  jand g08326(.dina(n26214), .dinb(n26348), .dout(n26349));
  jor  g08327(.dina(n26349), .dinb(n26176), .dout(n26350));
  jand g08328(.dina(n26218), .dinb(n26350), .dout(n26351));
  jor  g08329(.dina(n26351), .dinb(n26168), .dout(n26352));
  jand g08330(.dina(n26222), .dinb(n26352), .dout(n26353));
  jor  g08331(.dina(n26353), .dinb(n26162), .dout(n26354));
  jand g08332(.dina(n26226), .dinb(n26354), .dout(n26355));
  jor  g08333(.dina(n26355), .dinb(n26156), .dout(n26356));
  jand g08334(.dina(n26230), .dinb(n26356), .dout(n26357));
  jor  g08335(.dina(n26357), .dinb(n26150), .dout(n26358));
  jand g08336(.dina(n26234), .dinb(n26358), .dout(n26359));
  jor  g08337(.dina(n26359), .dinb(n26144), .dout(n26360));
  jand g08338(.dina(n26238), .dinb(n26360), .dout(n26361));
  jor  g08339(.dina(n26361), .dinb(n26138), .dout(n26362));
  jand g08340(.dina(n26242), .dinb(n26362), .dout(n26363));
  jor  g08341(.dina(n26363), .dinb(n26132), .dout(n26364));
  jand g08342(.dina(n26246), .dinb(n26364), .dout(n26365));
  jor  g08343(.dina(n26365), .dinb(n26126), .dout(n26366));
  jand g08344(.dina(n26250), .dinb(n26366), .dout(n26367));
  jor  g08345(.dina(n26367), .dinb(n26120), .dout(n26368));
  jand g08346(.dina(n26254), .dinb(n26368), .dout(n26369));
  jor  g08347(.dina(n26369), .dinb(n26114), .dout(n26370));
  jand g08348(.dina(n26258), .dinb(n26370), .dout(n26371));
  jor  g08349(.dina(n26371), .dinb(n26108), .dout(n26372));
  jand g08350(.dina(n26262), .dinb(n26372), .dout(n26373));
  jor  g08351(.dina(n26373), .dinb(n26102), .dout(n26374));
  jand g08352(.dina(n26266), .dinb(n26374), .dout(n26375));
  jor  g08353(.dina(n26375), .dinb(n26096), .dout(n26376));
  jand g08354(.dina(n26270), .dinb(n26376), .dout(n26377));
  jor  g08355(.dina(n26377), .dinb(n26090), .dout(n26378));
  jand g08356(.dina(n26274), .dinb(n26378), .dout(n26379));
  jor  g08357(.dina(n26379), .dinb(n26084), .dout(n26380));
  jand g08358(.dina(n26278), .dinb(n26380), .dout(n26381));
  jor  g08359(.dina(n26381), .dinb(n26078), .dout(n26382));
  jand g08360(.dina(n26282), .dinb(n26382), .dout(n26383));
  jor  g08361(.dina(n26383), .dinb(n26072), .dout(n26384));
  jand g08362(.dina(n26286), .dinb(n26384), .dout(n26385));
  jor  g08363(.dina(n26385), .dinb(n26066), .dout(n26386));
  jand g08364(.dina(n26290), .dinb(n26386), .dout(n26387));
  jor  g08365(.dina(n26387), .dinb(n26060), .dout(n26388));
  jand g08366(.dina(n26294), .dinb(n26388), .dout(n26389));
  jor  g08367(.dina(n26389), .dinb(n26054), .dout(n26390));
  jand g08368(.dina(n26298), .dinb(n26390), .dout(n26391));
  jor  g08369(.dina(n26391), .dinb(n26048), .dout(n26392));
  jand g08370(.dina(n26302), .dinb(n26392), .dout(n26393));
  jor  g08371(.dina(n26393), .dinb(n26042), .dout(n26394));
  jand g08372(.dina(n26306), .dinb(n26394), .dout(n26395));
  jor  g08373(.dina(n26395), .dinb(n26036), .dout(n26396));
  jand g08374(.dina(n26310), .dinb(n26396), .dout(n26397));
  jor  g08375(.dina(n26397), .dinb(n26030), .dout(n26398));
  jand g08376(.dina(n26314), .dinb(n26398), .dout(n26399));
  jor  g08377(.dina(n26399), .dinb(n26024), .dout(n26400));
  jand g08378(.dina(n26318), .dinb(n26400), .dout(n26401));
  jor  g08379(.dina(n26401), .dinb(n26018), .dout(n26402));
  jand g08380(.dina(n26322), .dinb(n26402), .dout(n26403));
  jor  g08381(.dina(n26403), .dinb(n26012), .dout(n26404));
  jand g08382(.dina(n26326), .dinb(n26404), .dout(n26405));
  jor  g08383(.dina(n26405), .dinb(n26006), .dout(n26406));
  jand g08384(.dina(n26330), .dinb(n26406), .dout(n26407));
  jor  g08385(.dina(n26407), .dinb(n26000), .dout(n26408));
  jand g08386(.dina(n26334), .dinb(n26408), .dout(n26409));
  jor  g08387(.dina(n26409), .dinb(n25994), .dout(n26410));
  jnot g08388(.din(n26339), .dout(n26411));
  jand g08389(.dina(n26411), .dinb(n26410), .dout(n26412));
  jand g08390(.dina(n25984), .dinb(n5703), .dout(n26413));
  jor  g08391(.dina(n26413), .dinb(n26412), .dout(n26414));
  jxor g08392(.dina(n26338), .dinb(n26410), .dout(n26415));
  jand g08393(.dina(n26415), .dinb(n26414), .dout(n26416));
  jor  g08394(.dina(n26416), .dinb(n26341), .dout(n26417));
  jnot g08395(.din(n26417), .dout(n26418));
  jand g08396(.dina(n26417), .dinb(b36 ), .dout(n26419));
  jnot g08397(.din(n26419), .dout(n26420));
  jand g08398(.dina(n26418), .dinb(n293), .dout(n26421));
  jnot g08399(.din(n26413), .dout(n26422));
  jand g08400(.dina(n26422), .dinb(n26340), .dout(n26423));
  jand g08401(.dina(n26423), .dinb(n25993), .dout(n26424));
  jxor g08402(.dina(n26334), .dinb(n26408), .dout(n26425));
  jand g08403(.dina(n26425), .dinb(n26414), .dout(n26426));
  jor  g08404(.dina(n26426), .dinb(n26424), .dout(n26427));
  jand g08405(.dina(n26427), .dinb(n301), .dout(n26428));
  jand g08406(.dina(n26423), .dinb(n25999), .dout(n26429));
  jxor g08407(.dina(n26330), .dinb(n26406), .dout(n26430));
  jand g08408(.dina(n26430), .dinb(n26414), .dout(n26431));
  jor  g08409(.dina(n26431), .dinb(n26429), .dout(n26432));
  jand g08410(.dina(n26432), .dinb(n298), .dout(n26433));
  jand g08411(.dina(n26423), .dinb(n26005), .dout(n26434));
  jxor g08412(.dina(n26326), .dinb(n26404), .dout(n26435));
  jand g08413(.dina(n26435), .dinb(n26414), .dout(n26436));
  jor  g08414(.dina(n26436), .dinb(n26434), .dout(n26437));
  jand g08415(.dina(n26437), .dinb(n297), .dout(n26438));
  jand g08416(.dina(n26423), .dinb(n26011), .dout(n26439));
  jxor g08417(.dina(n26322), .dinb(n26402), .dout(n26440));
  jand g08418(.dina(n26440), .dinb(n26414), .dout(n26441));
  jor  g08419(.dina(n26441), .dinb(n26439), .dout(n26442));
  jand g08420(.dina(n26442), .dinb(n300), .dout(n26443));
  jand g08421(.dina(n26423), .dinb(n26017), .dout(n26444));
  jxor g08422(.dina(n26318), .dinb(n26400), .dout(n26445));
  jand g08423(.dina(n26445), .dinb(n26414), .dout(n26446));
  jor  g08424(.dina(n26446), .dinb(n26444), .dout(n26447));
  jand g08425(.dina(n26447), .dinb(n424), .dout(n26448));
  jand g08426(.dina(n26423), .dinb(n26023), .dout(n26449));
  jxor g08427(.dina(n26314), .dinb(n26398), .dout(n26450));
  jand g08428(.dina(n26450), .dinb(n26414), .dout(n26451));
  jor  g08429(.dina(n26451), .dinb(n26449), .dout(n26452));
  jand g08430(.dina(n26452), .dinb(n427), .dout(n26453));
  jand g08431(.dina(n26423), .dinb(n26029), .dout(n26454));
  jxor g08432(.dina(n26310), .dinb(n26396), .dout(n26455));
  jand g08433(.dina(n26455), .dinb(n26414), .dout(n26456));
  jor  g08434(.dina(n26456), .dinb(n26454), .dout(n26457));
  jand g08435(.dina(n26457), .dinb(n426), .dout(n26458));
  jand g08436(.dina(n26423), .dinb(n26035), .dout(n26459));
  jxor g08437(.dina(n26306), .dinb(n26394), .dout(n26460));
  jand g08438(.dina(n26460), .dinb(n26414), .dout(n26461));
  jor  g08439(.dina(n26461), .dinb(n26459), .dout(n26462));
  jand g08440(.dina(n26462), .dinb(n410), .dout(n26463));
  jand g08441(.dina(n26423), .dinb(n26041), .dout(n26464));
  jxor g08442(.dina(n26302), .dinb(n26392), .dout(n26465));
  jand g08443(.dina(n26465), .dinb(n26414), .dout(n26466));
  jor  g08444(.dina(n26466), .dinb(n26464), .dout(n26467));
  jand g08445(.dina(n26467), .dinb(n409), .dout(n26468));
  jand g08446(.dina(n26423), .dinb(n26047), .dout(n26469));
  jxor g08447(.dina(n26298), .dinb(n26390), .dout(n26470));
  jand g08448(.dina(n26470), .dinb(n26414), .dout(n26471));
  jor  g08449(.dina(n26471), .dinb(n26469), .dout(n26472));
  jand g08450(.dina(n26472), .dinb(n413), .dout(n26473));
  jand g08451(.dina(n26423), .dinb(n26053), .dout(n26474));
  jxor g08452(.dina(n26294), .dinb(n26388), .dout(n26475));
  jand g08453(.dina(n26475), .dinb(n26414), .dout(n26476));
  jor  g08454(.dina(n26476), .dinb(n26474), .dout(n26477));
  jand g08455(.dina(n26477), .dinb(n412), .dout(n26478));
  jand g08456(.dina(n26423), .dinb(n26059), .dout(n26479));
  jxor g08457(.dina(n26290), .dinb(n26386), .dout(n26480));
  jand g08458(.dina(n26480), .dinb(n26414), .dout(n26481));
  jor  g08459(.dina(n26481), .dinb(n26479), .dout(n26482));
  jand g08460(.dina(n26482), .dinb(n406), .dout(n26483));
  jand g08461(.dina(n26423), .dinb(n26065), .dout(n26484));
  jxor g08462(.dina(n26286), .dinb(n26384), .dout(n26485));
  jand g08463(.dina(n26485), .dinb(n26414), .dout(n26486));
  jor  g08464(.dina(n26486), .dinb(n26484), .dout(n26487));
  jand g08465(.dina(n26487), .dinb(n405), .dout(n26488));
  jand g08466(.dina(n26423), .dinb(n26071), .dout(n26489));
  jxor g08467(.dina(n26282), .dinb(n26382), .dout(n26490));
  jand g08468(.dina(n26490), .dinb(n26414), .dout(n26491));
  jor  g08469(.dina(n26491), .dinb(n26489), .dout(n26492));
  jand g08470(.dina(n26492), .dinb(n2714), .dout(n26493));
  jand g08471(.dina(n26423), .dinb(n26077), .dout(n26494));
  jxor g08472(.dina(n26278), .dinb(n26380), .dout(n26495));
  jand g08473(.dina(n26495), .dinb(n26414), .dout(n26496));
  jor  g08474(.dina(n26496), .dinb(n26494), .dout(n26497));
  jand g08475(.dina(n26497), .dinb(n2547), .dout(n26498));
  jand g08476(.dina(n26423), .dinb(n26083), .dout(n26499));
  jxor g08477(.dina(n26274), .dinb(n26378), .dout(n26500));
  jand g08478(.dina(n26500), .dinb(n26414), .dout(n26501));
  jor  g08479(.dina(n26501), .dinb(n26499), .dout(n26502));
  jand g08480(.dina(n26502), .dinb(n417), .dout(n26503));
  jand g08481(.dina(n26423), .dinb(n26089), .dout(n26504));
  jxor g08482(.dina(n26270), .dinb(n26376), .dout(n26505));
  jand g08483(.dina(n26505), .dinb(n26414), .dout(n26506));
  jor  g08484(.dina(n26506), .dinb(n26504), .dout(n26507));
  jand g08485(.dina(n26507), .dinb(n416), .dout(n26508));
  jand g08486(.dina(n26423), .dinb(n26095), .dout(n26509));
  jxor g08487(.dina(n26266), .dinb(n26374), .dout(n26510));
  jand g08488(.dina(n26510), .dinb(n26414), .dout(n26511));
  jor  g08489(.dina(n26511), .dinb(n26509), .dout(n26512));
  jand g08490(.dina(n26512), .dinb(n422), .dout(n26513));
  jand g08491(.dina(n26423), .dinb(n26101), .dout(n26514));
  jxor g08492(.dina(n26262), .dinb(n26372), .dout(n26515));
  jand g08493(.dina(n26515), .dinb(n26414), .dout(n26516));
  jor  g08494(.dina(n26516), .dinb(n26514), .dout(n26517));
  jand g08495(.dina(n26517), .dinb(n421), .dout(n26518));
  jand g08496(.dina(n26423), .dinb(n26107), .dout(n26519));
  jxor g08497(.dina(n26258), .dinb(n26370), .dout(n26520));
  jand g08498(.dina(n26520), .dinb(n26414), .dout(n26521));
  jor  g08499(.dina(n26521), .dinb(n26519), .dout(n26522));
  jand g08500(.dina(n26522), .dinb(n433), .dout(n26523));
  jand g08501(.dina(n26423), .dinb(n26113), .dout(n26524));
  jxor g08502(.dina(n26254), .dinb(n26368), .dout(n26525));
  jand g08503(.dina(n26525), .dinb(n26414), .dout(n26526));
  jor  g08504(.dina(n26526), .dinb(n26524), .dout(n26527));
  jand g08505(.dina(n26527), .dinb(n432), .dout(n26528));
  jand g08506(.dina(n26423), .dinb(n26119), .dout(n26529));
  jxor g08507(.dina(n26250), .dinb(n26366), .dout(n26530));
  jand g08508(.dina(n26530), .dinb(n26414), .dout(n26531));
  jor  g08509(.dina(n26531), .dinb(n26529), .dout(n26532));
  jand g08510(.dina(n26532), .dinb(n436), .dout(n26533));
  jand g08511(.dina(n26423), .dinb(n26125), .dout(n26534));
  jxor g08512(.dina(n26246), .dinb(n26364), .dout(n26535));
  jand g08513(.dina(n26535), .dinb(n26414), .dout(n26536));
  jor  g08514(.dina(n26536), .dinb(n26534), .dout(n26537));
  jand g08515(.dina(n26537), .dinb(n435), .dout(n26538));
  jand g08516(.dina(n26423), .dinb(n26131), .dout(n26539));
  jxor g08517(.dina(n26242), .dinb(n26362), .dout(n26540));
  jand g08518(.dina(n26540), .dinb(n26414), .dout(n26541));
  jor  g08519(.dina(n26541), .dinb(n26539), .dout(n26542));
  jand g08520(.dina(n26542), .dinb(n440), .dout(n26543));
  jand g08521(.dina(n26423), .dinb(n26137), .dout(n26544));
  jxor g08522(.dina(n26238), .dinb(n26360), .dout(n26545));
  jand g08523(.dina(n26545), .dinb(n26414), .dout(n26546));
  jor  g08524(.dina(n26546), .dinb(n26544), .dout(n26547));
  jand g08525(.dina(n26547), .dinb(n439), .dout(n26548));
  jand g08526(.dina(n26423), .dinb(n26143), .dout(n26549));
  jxor g08527(.dina(n26234), .dinb(n26358), .dout(n26550));
  jand g08528(.dina(n26550), .dinb(n26414), .dout(n26551));
  jor  g08529(.dina(n26551), .dinb(n26549), .dout(n26552));
  jand g08530(.dina(n26552), .dinb(n325), .dout(n26553));
  jand g08531(.dina(n26423), .dinb(n26149), .dout(n26554));
  jxor g08532(.dina(n26230), .dinb(n26356), .dout(n26555));
  jand g08533(.dina(n26555), .dinb(n26414), .dout(n26556));
  jor  g08534(.dina(n26556), .dinb(n26554), .dout(n26557));
  jand g08535(.dina(n26557), .dinb(n324), .dout(n26558));
  jand g08536(.dina(n26423), .dinb(n26155), .dout(n26559));
  jxor g08537(.dina(n26226), .dinb(n26354), .dout(n26560));
  jand g08538(.dina(n26560), .dinb(n26414), .dout(n26561));
  jor  g08539(.dina(n26561), .dinb(n26559), .dout(n26562));
  jand g08540(.dina(n26562), .dinb(n323), .dout(n26563));
  jand g08541(.dina(n26423), .dinb(n26161), .dout(n26564));
  jxor g08542(.dina(n26222), .dinb(n26352), .dout(n26565));
  jand g08543(.dina(n26565), .dinb(n26414), .dout(n26566));
  jor  g08544(.dina(n26566), .dinb(n26564), .dout(n26567));
  jand g08545(.dina(n26567), .dinb(n335), .dout(n26568));
  jand g08546(.dina(n26423), .dinb(n26167), .dout(n26569));
  jxor g08547(.dina(n26218), .dinb(n26350), .dout(n26570));
  jand g08548(.dina(n26570), .dinb(n26414), .dout(n26571));
  jor  g08549(.dina(n26571), .dinb(n26569), .dout(n26572));
  jand g08550(.dina(n26572), .dinb(n334), .dout(n26573));
  jand g08551(.dina(n26423), .dinb(n26175), .dout(n26574));
  jxor g08552(.dina(n26214), .dinb(n26348), .dout(n26575));
  jand g08553(.dina(n26575), .dinb(n26414), .dout(n26576));
  jor  g08554(.dina(n26576), .dinb(n26574), .dout(n26577));
  jand g08555(.dina(n26577), .dinb(n338), .dout(n26578));
  jand g08556(.dina(n26423), .dinb(n26183), .dout(n26579));
  jxor g08557(.dina(n26210), .dinb(n26346), .dout(n26580));
  jand g08558(.dina(n26580), .dinb(n26414), .dout(n26581));
  jor  g08559(.dina(n26581), .dinb(n26579), .dout(n26582));
  jand g08560(.dina(n26582), .dinb(n337), .dout(n26583));
  jand g08561(.dina(n26423), .dinb(n26189), .dout(n26584));
  jxor g08562(.dina(n26206), .dinb(n26344), .dout(n26585));
  jand g08563(.dina(n26585), .dinb(n26414), .dout(n26586));
  jor  g08564(.dina(n26586), .dinb(n26584), .dout(n26587));
  jand g08565(.dina(n26587), .dinb(n344), .dout(n26588));
  jand g08566(.dina(n26423), .dinb(n26196), .dout(n26589));
  jxor g08567(.dina(n26342), .dinb(n6295), .dout(n26590));
  jand g08568(.dina(n26590), .dinb(n26414), .dout(n26591));
  jor  g08569(.dina(n26591), .dinb(n26589), .dout(n26592));
  jand g08570(.dina(n26592), .dinb(n348), .dout(n26593));
  jor  g08571(.dina(n26423), .dinb(n18364), .dout(n26594));
  jand g08572(.dina(n26594), .dinb(a28 ), .dout(n26595));
  jor  g08573(.dina(n26423), .dinb(n6295), .dout(n26596));
  jnot g08574(.din(n26596), .dout(n26597));
  jor  g08575(.dina(n26597), .dinb(n26595), .dout(n26598));
  jand g08576(.dina(n26598), .dinb(n258), .dout(n26599));
  jand g08577(.dina(n26414), .dinb(b0 ), .dout(n26600));
  jor  g08578(.dina(n26600), .dinb(n6293), .dout(n26601));
  jand g08579(.dina(n26596), .dinb(n26601), .dout(n26602));
  jxor g08580(.dina(n26602), .dinb(b1 ), .dout(n26603));
  jand g08581(.dina(n26603), .dinb(n6601), .dout(n26604));
  jor  g08582(.dina(n26604), .dinb(n26599), .dout(n26605));
  jxor g08583(.dina(n26592), .dinb(n348), .dout(n26606));
  jand g08584(.dina(n26606), .dinb(n26605), .dout(n26607));
  jor  g08585(.dina(n26607), .dinb(n26593), .dout(n26608));
  jxor g08586(.dina(n26587), .dinb(n344), .dout(n26609));
  jand g08587(.dina(n26609), .dinb(n26608), .dout(n26610));
  jor  g08588(.dina(n26610), .dinb(n26588), .dout(n26611));
  jxor g08589(.dina(n26582), .dinb(n337), .dout(n26612));
  jand g08590(.dina(n26612), .dinb(n26611), .dout(n26613));
  jor  g08591(.dina(n26613), .dinb(n26583), .dout(n26614));
  jxor g08592(.dina(n26577), .dinb(n338), .dout(n26615));
  jand g08593(.dina(n26615), .dinb(n26614), .dout(n26616));
  jor  g08594(.dina(n26616), .dinb(n26578), .dout(n26617));
  jxor g08595(.dina(n26572), .dinb(n334), .dout(n26618));
  jand g08596(.dina(n26618), .dinb(n26617), .dout(n26619));
  jor  g08597(.dina(n26619), .dinb(n26573), .dout(n26620));
  jxor g08598(.dina(n26567), .dinb(n335), .dout(n26621));
  jand g08599(.dina(n26621), .dinb(n26620), .dout(n26622));
  jor  g08600(.dina(n26622), .dinb(n26568), .dout(n26623));
  jxor g08601(.dina(n26562), .dinb(n323), .dout(n26624));
  jand g08602(.dina(n26624), .dinb(n26623), .dout(n26625));
  jor  g08603(.dina(n26625), .dinb(n26563), .dout(n26626));
  jxor g08604(.dina(n26557), .dinb(n324), .dout(n26627));
  jand g08605(.dina(n26627), .dinb(n26626), .dout(n26628));
  jor  g08606(.dina(n26628), .dinb(n26558), .dout(n26629));
  jxor g08607(.dina(n26552), .dinb(n325), .dout(n26630));
  jand g08608(.dina(n26630), .dinb(n26629), .dout(n26631));
  jor  g08609(.dina(n26631), .dinb(n26553), .dout(n26632));
  jxor g08610(.dina(n26547), .dinb(n439), .dout(n26633));
  jand g08611(.dina(n26633), .dinb(n26632), .dout(n26634));
  jor  g08612(.dina(n26634), .dinb(n26548), .dout(n26635));
  jxor g08613(.dina(n26542), .dinb(n440), .dout(n26636));
  jand g08614(.dina(n26636), .dinb(n26635), .dout(n26637));
  jor  g08615(.dina(n26637), .dinb(n26543), .dout(n26638));
  jxor g08616(.dina(n26537), .dinb(n435), .dout(n26639));
  jand g08617(.dina(n26639), .dinb(n26638), .dout(n26640));
  jor  g08618(.dina(n26640), .dinb(n26538), .dout(n26641));
  jxor g08619(.dina(n26532), .dinb(n436), .dout(n26642));
  jand g08620(.dina(n26642), .dinb(n26641), .dout(n26643));
  jor  g08621(.dina(n26643), .dinb(n26533), .dout(n26644));
  jxor g08622(.dina(n26527), .dinb(n432), .dout(n26645));
  jand g08623(.dina(n26645), .dinb(n26644), .dout(n26646));
  jor  g08624(.dina(n26646), .dinb(n26528), .dout(n26647));
  jxor g08625(.dina(n26522), .dinb(n433), .dout(n26648));
  jand g08626(.dina(n26648), .dinb(n26647), .dout(n26649));
  jor  g08627(.dina(n26649), .dinb(n26523), .dout(n26650));
  jxor g08628(.dina(n26517), .dinb(n421), .dout(n26651));
  jand g08629(.dina(n26651), .dinb(n26650), .dout(n26652));
  jor  g08630(.dina(n26652), .dinb(n26518), .dout(n26653));
  jxor g08631(.dina(n26512), .dinb(n422), .dout(n26654));
  jand g08632(.dina(n26654), .dinb(n26653), .dout(n26655));
  jor  g08633(.dina(n26655), .dinb(n26513), .dout(n26656));
  jxor g08634(.dina(n26507), .dinb(n416), .dout(n26657));
  jand g08635(.dina(n26657), .dinb(n26656), .dout(n26658));
  jor  g08636(.dina(n26658), .dinb(n26508), .dout(n26659));
  jxor g08637(.dina(n26502), .dinb(n417), .dout(n26660));
  jand g08638(.dina(n26660), .dinb(n26659), .dout(n26661));
  jor  g08639(.dina(n26661), .dinb(n26503), .dout(n26662));
  jxor g08640(.dina(n26497), .dinb(n2547), .dout(n26663));
  jand g08641(.dina(n26663), .dinb(n26662), .dout(n26664));
  jor  g08642(.dina(n26664), .dinb(n26498), .dout(n26665));
  jxor g08643(.dina(n26492), .dinb(n2714), .dout(n26666));
  jand g08644(.dina(n26666), .dinb(n26665), .dout(n26667));
  jor  g08645(.dina(n26667), .dinb(n26493), .dout(n26668));
  jxor g08646(.dina(n26487), .dinb(n405), .dout(n26669));
  jand g08647(.dina(n26669), .dinb(n26668), .dout(n26670));
  jor  g08648(.dina(n26670), .dinb(n26488), .dout(n26671));
  jxor g08649(.dina(n26482), .dinb(n406), .dout(n26672));
  jand g08650(.dina(n26672), .dinb(n26671), .dout(n26673));
  jor  g08651(.dina(n26673), .dinb(n26483), .dout(n26674));
  jxor g08652(.dina(n26477), .dinb(n412), .dout(n26675));
  jand g08653(.dina(n26675), .dinb(n26674), .dout(n26676));
  jor  g08654(.dina(n26676), .dinb(n26478), .dout(n26677));
  jxor g08655(.dina(n26472), .dinb(n413), .dout(n26678));
  jand g08656(.dina(n26678), .dinb(n26677), .dout(n26679));
  jor  g08657(.dina(n26679), .dinb(n26473), .dout(n26680));
  jxor g08658(.dina(n26467), .dinb(n409), .dout(n26681));
  jand g08659(.dina(n26681), .dinb(n26680), .dout(n26682));
  jor  g08660(.dina(n26682), .dinb(n26468), .dout(n26683));
  jxor g08661(.dina(n26462), .dinb(n410), .dout(n26684));
  jand g08662(.dina(n26684), .dinb(n26683), .dout(n26685));
  jor  g08663(.dina(n26685), .dinb(n26463), .dout(n26686));
  jxor g08664(.dina(n26457), .dinb(n426), .dout(n26687));
  jand g08665(.dina(n26687), .dinb(n26686), .dout(n26688));
  jor  g08666(.dina(n26688), .dinb(n26458), .dout(n26689));
  jxor g08667(.dina(n26452), .dinb(n427), .dout(n26690));
  jand g08668(.dina(n26690), .dinb(n26689), .dout(n26691));
  jor  g08669(.dina(n26691), .dinb(n26453), .dout(n26692));
  jxor g08670(.dina(n26447), .dinb(n424), .dout(n26693));
  jand g08671(.dina(n26693), .dinb(n26692), .dout(n26694));
  jor  g08672(.dina(n26694), .dinb(n26448), .dout(n26695));
  jxor g08673(.dina(n26442), .dinb(n300), .dout(n26696));
  jand g08674(.dina(n26696), .dinb(n26695), .dout(n26697));
  jor  g08675(.dina(n26697), .dinb(n26443), .dout(n26698));
  jxor g08676(.dina(n26437), .dinb(n297), .dout(n26699));
  jand g08677(.dina(n26699), .dinb(n26698), .dout(n26700));
  jor  g08678(.dina(n26700), .dinb(n26438), .dout(n26701));
  jxor g08679(.dina(n26432), .dinb(n298), .dout(n26702));
  jand g08680(.dina(n26702), .dinb(n26701), .dout(n26703));
  jor  g08681(.dina(n26703), .dinb(n26433), .dout(n26704));
  jxor g08682(.dina(n26427), .dinb(n301), .dout(n26705));
  jand g08683(.dina(n26705), .dinb(n26704), .dout(n26706));
  jor  g08684(.dina(n26706), .dinb(n26428), .dout(n26707));
  jor  g08685(.dina(n26707), .dinb(n26421), .dout(n26708));
  jand g08686(.dina(n26708), .dinb(n26420), .dout(n26709));
  jand g08687(.dina(n26709), .dinb(n5702), .dout(n26710));
  jnot g08688(.din(n26710), .dout(n26711));
  jand g08689(.dina(n26711), .dinb(n26418), .dout(n26712));
  jand g08690(.dina(n26421), .dinb(n5702), .dout(n26713));
  jand g08691(.dina(n26713), .dinb(n26707), .dout(n26714));
  jor  g08692(.dina(n26714), .dinb(n26712), .dout(n26715));
  jand g08693(.dina(n26715), .dinb(n294), .dout(n26716));
  jnot g08694(.din(n26716), .dout(n26717));
  jand g08695(.dina(n26711), .dinb(n26427), .dout(n26718));
  jxor g08696(.dina(n26705), .dinb(n26704), .dout(n26719));
  jand g08697(.dina(n26719), .dinb(n26710), .dout(n26720));
  jor  g08698(.dina(n26720), .dinb(n26718), .dout(n26721));
  jand g08699(.dina(n26721), .dinb(n293), .dout(n26722));
  jnot g08700(.din(n26722), .dout(n26723));
  jand g08701(.dina(n26711), .dinb(n26432), .dout(n26724));
  jxor g08702(.dina(n26702), .dinb(n26701), .dout(n26725));
  jand g08703(.dina(n26725), .dinb(n26710), .dout(n26726));
  jor  g08704(.dina(n26726), .dinb(n26724), .dout(n26727));
  jand g08705(.dina(n26727), .dinb(n301), .dout(n26728));
  jnot g08706(.din(n26728), .dout(n26729));
  jand g08707(.dina(n26711), .dinb(n26437), .dout(n26730));
  jxor g08708(.dina(n26699), .dinb(n26698), .dout(n26731));
  jand g08709(.dina(n26731), .dinb(n26710), .dout(n26732));
  jor  g08710(.dina(n26732), .dinb(n26730), .dout(n26733));
  jand g08711(.dina(n26733), .dinb(n298), .dout(n26734));
  jnot g08712(.din(n26734), .dout(n26735));
  jand g08713(.dina(n26711), .dinb(n26442), .dout(n26736));
  jxor g08714(.dina(n26696), .dinb(n26695), .dout(n26737));
  jand g08715(.dina(n26737), .dinb(n26710), .dout(n26738));
  jor  g08716(.dina(n26738), .dinb(n26736), .dout(n26739));
  jand g08717(.dina(n26739), .dinb(n297), .dout(n26740));
  jnot g08718(.din(n26740), .dout(n26741));
  jand g08719(.dina(n26711), .dinb(n26447), .dout(n26742));
  jxor g08720(.dina(n26693), .dinb(n26692), .dout(n26743));
  jand g08721(.dina(n26743), .dinb(n26710), .dout(n26744));
  jor  g08722(.dina(n26744), .dinb(n26742), .dout(n26745));
  jand g08723(.dina(n26745), .dinb(n300), .dout(n26746));
  jnot g08724(.din(n26746), .dout(n26747));
  jand g08725(.dina(n26711), .dinb(n26452), .dout(n26748));
  jxor g08726(.dina(n26690), .dinb(n26689), .dout(n26749));
  jand g08727(.dina(n26749), .dinb(n26710), .dout(n26750));
  jor  g08728(.dina(n26750), .dinb(n26748), .dout(n26751));
  jand g08729(.dina(n26751), .dinb(n424), .dout(n26752));
  jnot g08730(.din(n26752), .dout(n26753));
  jand g08731(.dina(n26711), .dinb(n26457), .dout(n26754));
  jxor g08732(.dina(n26687), .dinb(n26686), .dout(n26755));
  jand g08733(.dina(n26755), .dinb(n26710), .dout(n26756));
  jor  g08734(.dina(n26756), .dinb(n26754), .dout(n26757));
  jand g08735(.dina(n26757), .dinb(n427), .dout(n26758));
  jnot g08736(.din(n26758), .dout(n26759));
  jand g08737(.dina(n26711), .dinb(n26462), .dout(n26760));
  jxor g08738(.dina(n26684), .dinb(n26683), .dout(n26761));
  jand g08739(.dina(n26761), .dinb(n26710), .dout(n26762));
  jor  g08740(.dina(n26762), .dinb(n26760), .dout(n26763));
  jand g08741(.dina(n26763), .dinb(n426), .dout(n26764));
  jnot g08742(.din(n26764), .dout(n26765));
  jand g08743(.dina(n26711), .dinb(n26467), .dout(n26766));
  jxor g08744(.dina(n26681), .dinb(n26680), .dout(n26767));
  jand g08745(.dina(n26767), .dinb(n26710), .dout(n26768));
  jor  g08746(.dina(n26768), .dinb(n26766), .dout(n26769));
  jand g08747(.dina(n26769), .dinb(n410), .dout(n26770));
  jnot g08748(.din(n26770), .dout(n26771));
  jand g08749(.dina(n26711), .dinb(n26472), .dout(n26772));
  jxor g08750(.dina(n26678), .dinb(n26677), .dout(n26773));
  jand g08751(.dina(n26773), .dinb(n26710), .dout(n26774));
  jor  g08752(.dina(n26774), .dinb(n26772), .dout(n26775));
  jand g08753(.dina(n26775), .dinb(n409), .dout(n26776));
  jnot g08754(.din(n26776), .dout(n26777));
  jand g08755(.dina(n26711), .dinb(n26477), .dout(n26778));
  jxor g08756(.dina(n26675), .dinb(n26674), .dout(n26779));
  jand g08757(.dina(n26779), .dinb(n26710), .dout(n26780));
  jor  g08758(.dina(n26780), .dinb(n26778), .dout(n26781));
  jand g08759(.dina(n26781), .dinb(n413), .dout(n26782));
  jnot g08760(.din(n26782), .dout(n26783));
  jand g08761(.dina(n26711), .dinb(n26482), .dout(n26784));
  jxor g08762(.dina(n26672), .dinb(n26671), .dout(n26785));
  jand g08763(.dina(n26785), .dinb(n26710), .dout(n26786));
  jor  g08764(.dina(n26786), .dinb(n26784), .dout(n26787));
  jand g08765(.dina(n26787), .dinb(n412), .dout(n26788));
  jnot g08766(.din(n26788), .dout(n26789));
  jand g08767(.dina(n26711), .dinb(n26487), .dout(n26790));
  jxor g08768(.dina(n26669), .dinb(n26668), .dout(n26791));
  jand g08769(.dina(n26791), .dinb(n26710), .dout(n26792));
  jor  g08770(.dina(n26792), .dinb(n26790), .dout(n26793));
  jand g08771(.dina(n26793), .dinb(n406), .dout(n26794));
  jnot g08772(.din(n26794), .dout(n26795));
  jand g08773(.dina(n26711), .dinb(n26492), .dout(n26796));
  jxor g08774(.dina(n26666), .dinb(n26665), .dout(n26797));
  jand g08775(.dina(n26797), .dinb(n26710), .dout(n26798));
  jor  g08776(.dina(n26798), .dinb(n26796), .dout(n26799));
  jand g08777(.dina(n26799), .dinb(n405), .dout(n26800));
  jnot g08778(.din(n26800), .dout(n26801));
  jand g08779(.dina(n26711), .dinb(n26497), .dout(n26802));
  jxor g08780(.dina(n26663), .dinb(n26662), .dout(n26803));
  jand g08781(.dina(n26803), .dinb(n26710), .dout(n26804));
  jor  g08782(.dina(n26804), .dinb(n26802), .dout(n26805));
  jand g08783(.dina(n26805), .dinb(n2714), .dout(n26806));
  jnot g08784(.din(n26806), .dout(n26807));
  jand g08785(.dina(n26711), .dinb(n26502), .dout(n26808));
  jxor g08786(.dina(n26660), .dinb(n26659), .dout(n26809));
  jand g08787(.dina(n26809), .dinb(n26710), .dout(n26810));
  jor  g08788(.dina(n26810), .dinb(n26808), .dout(n26811));
  jand g08789(.dina(n26811), .dinb(n2547), .dout(n26812));
  jnot g08790(.din(n26812), .dout(n26813));
  jand g08791(.dina(n26711), .dinb(n26507), .dout(n26814));
  jxor g08792(.dina(n26657), .dinb(n26656), .dout(n26815));
  jand g08793(.dina(n26815), .dinb(n26710), .dout(n26816));
  jor  g08794(.dina(n26816), .dinb(n26814), .dout(n26817));
  jand g08795(.dina(n26817), .dinb(n417), .dout(n26818));
  jnot g08796(.din(n26818), .dout(n26819));
  jand g08797(.dina(n26711), .dinb(n26512), .dout(n26820));
  jxor g08798(.dina(n26654), .dinb(n26653), .dout(n26821));
  jand g08799(.dina(n26821), .dinb(n26710), .dout(n26822));
  jor  g08800(.dina(n26822), .dinb(n26820), .dout(n26823));
  jand g08801(.dina(n26823), .dinb(n416), .dout(n26824));
  jnot g08802(.din(n26824), .dout(n26825));
  jand g08803(.dina(n26711), .dinb(n26517), .dout(n26826));
  jxor g08804(.dina(n26651), .dinb(n26650), .dout(n26827));
  jand g08805(.dina(n26827), .dinb(n26710), .dout(n26828));
  jor  g08806(.dina(n26828), .dinb(n26826), .dout(n26829));
  jand g08807(.dina(n26829), .dinb(n422), .dout(n26830));
  jnot g08808(.din(n26830), .dout(n26831));
  jand g08809(.dina(n26711), .dinb(n26522), .dout(n26832));
  jxor g08810(.dina(n26648), .dinb(n26647), .dout(n26833));
  jand g08811(.dina(n26833), .dinb(n26710), .dout(n26834));
  jor  g08812(.dina(n26834), .dinb(n26832), .dout(n26835));
  jand g08813(.dina(n26835), .dinb(n421), .dout(n26836));
  jnot g08814(.din(n26836), .dout(n26837));
  jand g08815(.dina(n26711), .dinb(n26527), .dout(n26838));
  jxor g08816(.dina(n26645), .dinb(n26644), .dout(n26839));
  jand g08817(.dina(n26839), .dinb(n26710), .dout(n26840));
  jor  g08818(.dina(n26840), .dinb(n26838), .dout(n26841));
  jand g08819(.dina(n26841), .dinb(n433), .dout(n26842));
  jnot g08820(.din(n26842), .dout(n26843));
  jand g08821(.dina(n26711), .dinb(n26532), .dout(n26844));
  jxor g08822(.dina(n26642), .dinb(n26641), .dout(n26845));
  jand g08823(.dina(n26845), .dinb(n26710), .dout(n26846));
  jor  g08824(.dina(n26846), .dinb(n26844), .dout(n26847));
  jand g08825(.dina(n26847), .dinb(n432), .dout(n26848));
  jnot g08826(.din(n26848), .dout(n26849));
  jand g08827(.dina(n26711), .dinb(n26537), .dout(n26850));
  jxor g08828(.dina(n26639), .dinb(n26638), .dout(n26851));
  jand g08829(.dina(n26851), .dinb(n26710), .dout(n26852));
  jor  g08830(.dina(n26852), .dinb(n26850), .dout(n26853));
  jand g08831(.dina(n26853), .dinb(n436), .dout(n26854));
  jnot g08832(.din(n26854), .dout(n26855));
  jand g08833(.dina(n26711), .dinb(n26542), .dout(n26856));
  jxor g08834(.dina(n26636), .dinb(n26635), .dout(n26857));
  jand g08835(.dina(n26857), .dinb(n26710), .dout(n26858));
  jor  g08836(.dina(n26858), .dinb(n26856), .dout(n26859));
  jand g08837(.dina(n26859), .dinb(n435), .dout(n26860));
  jnot g08838(.din(n26860), .dout(n26861));
  jand g08839(.dina(n26711), .dinb(n26547), .dout(n26862));
  jxor g08840(.dina(n26633), .dinb(n26632), .dout(n26863));
  jand g08841(.dina(n26863), .dinb(n26710), .dout(n26864));
  jor  g08842(.dina(n26864), .dinb(n26862), .dout(n26865));
  jand g08843(.dina(n26865), .dinb(n440), .dout(n26866));
  jnot g08844(.din(n26866), .dout(n26867));
  jand g08845(.dina(n26711), .dinb(n26552), .dout(n26868));
  jxor g08846(.dina(n26630), .dinb(n26629), .dout(n26869));
  jand g08847(.dina(n26869), .dinb(n26710), .dout(n26870));
  jor  g08848(.dina(n26870), .dinb(n26868), .dout(n26871));
  jand g08849(.dina(n26871), .dinb(n439), .dout(n26872));
  jnot g08850(.din(n26872), .dout(n26873));
  jand g08851(.dina(n26711), .dinb(n26557), .dout(n26874));
  jxor g08852(.dina(n26627), .dinb(n26626), .dout(n26875));
  jand g08853(.dina(n26875), .dinb(n26710), .dout(n26876));
  jor  g08854(.dina(n26876), .dinb(n26874), .dout(n26877));
  jand g08855(.dina(n26877), .dinb(n325), .dout(n26878));
  jnot g08856(.din(n26878), .dout(n26879));
  jand g08857(.dina(n26711), .dinb(n26562), .dout(n26880));
  jxor g08858(.dina(n26624), .dinb(n26623), .dout(n26881));
  jand g08859(.dina(n26881), .dinb(n26710), .dout(n26882));
  jor  g08860(.dina(n26882), .dinb(n26880), .dout(n26883));
  jand g08861(.dina(n26883), .dinb(n324), .dout(n26884));
  jnot g08862(.din(n26884), .dout(n26885));
  jand g08863(.dina(n26711), .dinb(n26567), .dout(n26886));
  jxor g08864(.dina(n26621), .dinb(n26620), .dout(n26887));
  jand g08865(.dina(n26887), .dinb(n26710), .dout(n26888));
  jor  g08866(.dina(n26888), .dinb(n26886), .dout(n26889));
  jand g08867(.dina(n26889), .dinb(n323), .dout(n26890));
  jnot g08868(.din(n26890), .dout(n26891));
  jand g08869(.dina(n26711), .dinb(n26572), .dout(n26892));
  jxor g08870(.dina(n26618), .dinb(n26617), .dout(n26893));
  jand g08871(.dina(n26893), .dinb(n26710), .dout(n26894));
  jor  g08872(.dina(n26894), .dinb(n26892), .dout(n26895));
  jand g08873(.dina(n26895), .dinb(n335), .dout(n26896));
  jnot g08874(.din(n26896), .dout(n26897));
  jand g08875(.dina(n26711), .dinb(n26577), .dout(n26898));
  jxor g08876(.dina(n26615), .dinb(n26614), .dout(n26899));
  jand g08877(.dina(n26899), .dinb(n26710), .dout(n26900));
  jor  g08878(.dina(n26900), .dinb(n26898), .dout(n26901));
  jand g08879(.dina(n26901), .dinb(n334), .dout(n26902));
  jnot g08880(.din(n26902), .dout(n26903));
  jand g08881(.dina(n26711), .dinb(n26582), .dout(n26904));
  jxor g08882(.dina(n26612), .dinb(n26611), .dout(n26905));
  jand g08883(.dina(n26905), .dinb(n26710), .dout(n26906));
  jor  g08884(.dina(n26906), .dinb(n26904), .dout(n26907));
  jand g08885(.dina(n26907), .dinb(n338), .dout(n26908));
  jnot g08886(.din(n26908), .dout(n26909));
  jand g08887(.dina(n26711), .dinb(n26587), .dout(n26910));
  jxor g08888(.dina(n26609), .dinb(n26608), .dout(n26911));
  jand g08889(.dina(n26911), .dinb(n26710), .dout(n26912));
  jor  g08890(.dina(n26912), .dinb(n26910), .dout(n26913));
  jand g08891(.dina(n26913), .dinb(n337), .dout(n26914));
  jnot g08892(.din(n26914), .dout(n26915));
  jnot g08893(.din(n26592), .dout(n26916));
  jor  g08894(.dina(n26710), .dinb(n26916), .dout(n26917));
  jxor g08895(.dina(n26606), .dinb(n26605), .dout(n26918));
  jnot g08896(.din(n26918), .dout(n26919));
  jor  g08897(.dina(n26919), .dinb(n26711), .dout(n26920));
  jand g08898(.dina(n26920), .dinb(n26917), .dout(n26921));
  jor  g08899(.dina(n26921), .dinb(b3 ), .dout(n26922));
  jor  g08900(.dina(n26710), .dinb(n26602), .dout(n26923));
  jxor g08901(.dina(n26603), .dinb(n6601), .dout(n26924));
  jand g08902(.dina(n26924), .dinb(n26710), .dout(n26925));
  jnot g08903(.din(n26925), .dout(n26926));
  jand g08904(.dina(n26926), .dinb(n26923), .dout(n26927));
  jor  g08905(.dina(n26927), .dinb(b2 ), .dout(n26928));
  jand g08906(.dina(n26709), .dinb(n6930), .dout(n26929));
  jor  g08907(.dina(n26929), .dinb(n6599), .dout(n26930));
  jnot g08908(.din(n6933), .dout(n26931));
  jnot g08909(.din(n26421), .dout(n26932));
  jnot g08910(.din(n26428), .dout(n26933));
  jnot g08911(.din(n26433), .dout(n26934));
  jnot g08912(.din(n26438), .dout(n26935));
  jnot g08913(.din(n26443), .dout(n26936));
  jnot g08914(.din(n26448), .dout(n26937));
  jnot g08915(.din(n26453), .dout(n26938));
  jnot g08916(.din(n26458), .dout(n26939));
  jnot g08917(.din(n26463), .dout(n26940));
  jnot g08918(.din(n26468), .dout(n26941));
  jnot g08919(.din(n26473), .dout(n26942));
  jnot g08920(.din(n26478), .dout(n26943));
  jnot g08921(.din(n26483), .dout(n26944));
  jnot g08922(.din(n26488), .dout(n26945));
  jnot g08923(.din(n26493), .dout(n26946));
  jnot g08924(.din(n26498), .dout(n26947));
  jnot g08925(.din(n26503), .dout(n26948));
  jnot g08926(.din(n26508), .dout(n26949));
  jnot g08927(.din(n26513), .dout(n26950));
  jnot g08928(.din(n26518), .dout(n26951));
  jnot g08929(.din(n26523), .dout(n26952));
  jnot g08930(.din(n26528), .dout(n26953));
  jnot g08931(.din(n26533), .dout(n26954));
  jnot g08932(.din(n26538), .dout(n26955));
  jnot g08933(.din(n26543), .dout(n26956));
  jnot g08934(.din(n26548), .dout(n26957));
  jnot g08935(.din(n26553), .dout(n26958));
  jnot g08936(.din(n26558), .dout(n26959));
  jnot g08937(.din(n26563), .dout(n26960));
  jnot g08938(.din(n26568), .dout(n26961));
  jnot g08939(.din(n26573), .dout(n26962));
  jnot g08940(.din(n26578), .dout(n26963));
  jnot g08941(.din(n26583), .dout(n26964));
  jnot g08942(.din(n26588), .dout(n26965));
  jnot g08943(.din(n26593), .dout(n26966));
  jnot g08944(.din(n26599), .dout(n26967));
  jxor g08945(.dina(n26602), .dinb(n258), .dout(n26968));
  jor  g08946(.dina(n26968), .dinb(n6600), .dout(n26969));
  jand g08947(.dina(n26969), .dinb(n26967), .dout(n26970));
  jnot g08948(.din(n26606), .dout(n26971));
  jor  g08949(.dina(n26971), .dinb(n26970), .dout(n26972));
  jand g08950(.dina(n26972), .dinb(n26966), .dout(n26973));
  jnot g08951(.din(n26609), .dout(n26974));
  jor  g08952(.dina(n26974), .dinb(n26973), .dout(n26975));
  jand g08953(.dina(n26975), .dinb(n26965), .dout(n26976));
  jnot g08954(.din(n26612), .dout(n26977));
  jor  g08955(.dina(n26977), .dinb(n26976), .dout(n26978));
  jand g08956(.dina(n26978), .dinb(n26964), .dout(n26979));
  jnot g08957(.din(n26615), .dout(n26980));
  jor  g08958(.dina(n26980), .dinb(n26979), .dout(n26981));
  jand g08959(.dina(n26981), .dinb(n26963), .dout(n26982));
  jnot g08960(.din(n26618), .dout(n26983));
  jor  g08961(.dina(n26983), .dinb(n26982), .dout(n26984));
  jand g08962(.dina(n26984), .dinb(n26962), .dout(n26985));
  jnot g08963(.din(n26621), .dout(n26986));
  jor  g08964(.dina(n26986), .dinb(n26985), .dout(n26987));
  jand g08965(.dina(n26987), .dinb(n26961), .dout(n26988));
  jnot g08966(.din(n26624), .dout(n26989));
  jor  g08967(.dina(n26989), .dinb(n26988), .dout(n26990));
  jand g08968(.dina(n26990), .dinb(n26960), .dout(n26991));
  jnot g08969(.din(n26627), .dout(n26992));
  jor  g08970(.dina(n26992), .dinb(n26991), .dout(n26993));
  jand g08971(.dina(n26993), .dinb(n26959), .dout(n26994));
  jnot g08972(.din(n26630), .dout(n26995));
  jor  g08973(.dina(n26995), .dinb(n26994), .dout(n26996));
  jand g08974(.dina(n26996), .dinb(n26958), .dout(n26997));
  jnot g08975(.din(n26633), .dout(n26998));
  jor  g08976(.dina(n26998), .dinb(n26997), .dout(n26999));
  jand g08977(.dina(n26999), .dinb(n26957), .dout(n27000));
  jnot g08978(.din(n26636), .dout(n27001));
  jor  g08979(.dina(n27001), .dinb(n27000), .dout(n27002));
  jand g08980(.dina(n27002), .dinb(n26956), .dout(n27003));
  jnot g08981(.din(n26639), .dout(n27004));
  jor  g08982(.dina(n27004), .dinb(n27003), .dout(n27005));
  jand g08983(.dina(n27005), .dinb(n26955), .dout(n27006));
  jnot g08984(.din(n26642), .dout(n27007));
  jor  g08985(.dina(n27007), .dinb(n27006), .dout(n27008));
  jand g08986(.dina(n27008), .dinb(n26954), .dout(n27009));
  jnot g08987(.din(n26645), .dout(n27010));
  jor  g08988(.dina(n27010), .dinb(n27009), .dout(n27011));
  jand g08989(.dina(n27011), .dinb(n26953), .dout(n27012));
  jnot g08990(.din(n26648), .dout(n27013));
  jor  g08991(.dina(n27013), .dinb(n27012), .dout(n27014));
  jand g08992(.dina(n27014), .dinb(n26952), .dout(n27015));
  jnot g08993(.din(n26651), .dout(n27016));
  jor  g08994(.dina(n27016), .dinb(n27015), .dout(n27017));
  jand g08995(.dina(n27017), .dinb(n26951), .dout(n27018));
  jnot g08996(.din(n26654), .dout(n27019));
  jor  g08997(.dina(n27019), .dinb(n27018), .dout(n27020));
  jand g08998(.dina(n27020), .dinb(n26950), .dout(n27021));
  jnot g08999(.din(n26657), .dout(n27022));
  jor  g09000(.dina(n27022), .dinb(n27021), .dout(n27023));
  jand g09001(.dina(n27023), .dinb(n26949), .dout(n27024));
  jnot g09002(.din(n26660), .dout(n27025));
  jor  g09003(.dina(n27025), .dinb(n27024), .dout(n27026));
  jand g09004(.dina(n27026), .dinb(n26948), .dout(n27027));
  jnot g09005(.din(n26663), .dout(n27028));
  jor  g09006(.dina(n27028), .dinb(n27027), .dout(n27029));
  jand g09007(.dina(n27029), .dinb(n26947), .dout(n27030));
  jnot g09008(.din(n26666), .dout(n27031));
  jor  g09009(.dina(n27031), .dinb(n27030), .dout(n27032));
  jand g09010(.dina(n27032), .dinb(n26946), .dout(n27033));
  jnot g09011(.din(n26669), .dout(n27034));
  jor  g09012(.dina(n27034), .dinb(n27033), .dout(n27035));
  jand g09013(.dina(n27035), .dinb(n26945), .dout(n27036));
  jnot g09014(.din(n26672), .dout(n27037));
  jor  g09015(.dina(n27037), .dinb(n27036), .dout(n27038));
  jand g09016(.dina(n27038), .dinb(n26944), .dout(n27039));
  jnot g09017(.din(n26675), .dout(n27040));
  jor  g09018(.dina(n27040), .dinb(n27039), .dout(n27041));
  jand g09019(.dina(n27041), .dinb(n26943), .dout(n27042));
  jnot g09020(.din(n26678), .dout(n27043));
  jor  g09021(.dina(n27043), .dinb(n27042), .dout(n27044));
  jand g09022(.dina(n27044), .dinb(n26942), .dout(n27045));
  jnot g09023(.din(n26681), .dout(n27046));
  jor  g09024(.dina(n27046), .dinb(n27045), .dout(n27047));
  jand g09025(.dina(n27047), .dinb(n26941), .dout(n27048));
  jnot g09026(.din(n26684), .dout(n27049));
  jor  g09027(.dina(n27049), .dinb(n27048), .dout(n27050));
  jand g09028(.dina(n27050), .dinb(n26940), .dout(n27051));
  jnot g09029(.din(n26687), .dout(n27052));
  jor  g09030(.dina(n27052), .dinb(n27051), .dout(n27053));
  jand g09031(.dina(n27053), .dinb(n26939), .dout(n27054));
  jnot g09032(.din(n26690), .dout(n27055));
  jor  g09033(.dina(n27055), .dinb(n27054), .dout(n27056));
  jand g09034(.dina(n27056), .dinb(n26938), .dout(n27057));
  jnot g09035(.din(n26693), .dout(n27058));
  jor  g09036(.dina(n27058), .dinb(n27057), .dout(n27059));
  jand g09037(.dina(n27059), .dinb(n26937), .dout(n27060));
  jnot g09038(.din(n26696), .dout(n27061));
  jor  g09039(.dina(n27061), .dinb(n27060), .dout(n27062));
  jand g09040(.dina(n27062), .dinb(n26936), .dout(n27063));
  jnot g09041(.din(n26699), .dout(n27064));
  jor  g09042(.dina(n27064), .dinb(n27063), .dout(n27065));
  jand g09043(.dina(n27065), .dinb(n26935), .dout(n27066));
  jnot g09044(.din(n26702), .dout(n27067));
  jor  g09045(.dina(n27067), .dinb(n27066), .dout(n27068));
  jand g09046(.dina(n27068), .dinb(n26934), .dout(n27069));
  jnot g09047(.din(n26705), .dout(n27070));
  jor  g09048(.dina(n27070), .dinb(n27069), .dout(n27071));
  jand g09049(.dina(n27071), .dinb(n26933), .dout(n27072));
  jand g09050(.dina(n27072), .dinb(n26932), .dout(n27073));
  jor  g09051(.dina(n27073), .dinb(n26419), .dout(n27074));
  jor  g09052(.dina(n27074), .dinb(n26931), .dout(n27075));
  jand g09053(.dina(n27075), .dinb(n26930), .dout(n27076));
  jor  g09054(.dina(n27076), .dinb(b1 ), .dout(n27077));
  jxor g09055(.dina(n27076), .dinb(n258), .dout(n27078));
  jor  g09056(.dina(n27078), .dinb(n6939), .dout(n27079));
  jand g09057(.dina(n27079), .dinb(n27077), .dout(n27080));
  jxor g09058(.dina(n26927), .dinb(n348), .dout(n27081));
  jor  g09059(.dina(n27081), .dinb(n27080), .dout(n27082));
  jand g09060(.dina(n27082), .dinb(n26928), .dout(n27083));
  jxor g09061(.dina(n26921), .dinb(b3 ), .dout(n27084));
  jnot g09062(.din(n27084), .dout(n27085));
  jor  g09063(.dina(n27085), .dinb(n27083), .dout(n27086));
  jand g09064(.dina(n27086), .dinb(n26922), .dout(n27087));
  jxor g09065(.dina(n26913), .dinb(n337), .dout(n27088));
  jnot g09066(.din(n27088), .dout(n27089));
  jor  g09067(.dina(n27089), .dinb(n27087), .dout(n27090));
  jand g09068(.dina(n27090), .dinb(n26915), .dout(n27091));
  jxor g09069(.dina(n26907), .dinb(n338), .dout(n27092));
  jnot g09070(.din(n27092), .dout(n27093));
  jor  g09071(.dina(n27093), .dinb(n27091), .dout(n27094));
  jand g09072(.dina(n27094), .dinb(n26909), .dout(n27095));
  jxor g09073(.dina(n26901), .dinb(n334), .dout(n27096));
  jnot g09074(.din(n27096), .dout(n27097));
  jor  g09075(.dina(n27097), .dinb(n27095), .dout(n27098));
  jand g09076(.dina(n27098), .dinb(n26903), .dout(n27099));
  jxor g09077(.dina(n26895), .dinb(n335), .dout(n27100));
  jnot g09078(.din(n27100), .dout(n27101));
  jor  g09079(.dina(n27101), .dinb(n27099), .dout(n27102));
  jand g09080(.dina(n27102), .dinb(n26897), .dout(n27103));
  jxor g09081(.dina(n26889), .dinb(n323), .dout(n27104));
  jnot g09082(.din(n27104), .dout(n27105));
  jor  g09083(.dina(n27105), .dinb(n27103), .dout(n27106));
  jand g09084(.dina(n27106), .dinb(n26891), .dout(n27107));
  jxor g09085(.dina(n26883), .dinb(n324), .dout(n27108));
  jnot g09086(.din(n27108), .dout(n27109));
  jor  g09087(.dina(n27109), .dinb(n27107), .dout(n27110));
  jand g09088(.dina(n27110), .dinb(n26885), .dout(n27111));
  jxor g09089(.dina(n26877), .dinb(n325), .dout(n27112));
  jnot g09090(.din(n27112), .dout(n27113));
  jor  g09091(.dina(n27113), .dinb(n27111), .dout(n27114));
  jand g09092(.dina(n27114), .dinb(n26879), .dout(n27115));
  jxor g09093(.dina(n26871), .dinb(n439), .dout(n27116));
  jnot g09094(.din(n27116), .dout(n27117));
  jor  g09095(.dina(n27117), .dinb(n27115), .dout(n27118));
  jand g09096(.dina(n27118), .dinb(n26873), .dout(n27119));
  jxor g09097(.dina(n26865), .dinb(n440), .dout(n27120));
  jnot g09098(.din(n27120), .dout(n27121));
  jor  g09099(.dina(n27121), .dinb(n27119), .dout(n27122));
  jand g09100(.dina(n27122), .dinb(n26867), .dout(n27123));
  jxor g09101(.dina(n26859), .dinb(n435), .dout(n27124));
  jnot g09102(.din(n27124), .dout(n27125));
  jor  g09103(.dina(n27125), .dinb(n27123), .dout(n27126));
  jand g09104(.dina(n27126), .dinb(n26861), .dout(n27127));
  jxor g09105(.dina(n26853), .dinb(n436), .dout(n27128));
  jnot g09106(.din(n27128), .dout(n27129));
  jor  g09107(.dina(n27129), .dinb(n27127), .dout(n27130));
  jand g09108(.dina(n27130), .dinb(n26855), .dout(n27131));
  jxor g09109(.dina(n26847), .dinb(n432), .dout(n27132));
  jnot g09110(.din(n27132), .dout(n27133));
  jor  g09111(.dina(n27133), .dinb(n27131), .dout(n27134));
  jand g09112(.dina(n27134), .dinb(n26849), .dout(n27135));
  jxor g09113(.dina(n26841), .dinb(n433), .dout(n27136));
  jnot g09114(.din(n27136), .dout(n27137));
  jor  g09115(.dina(n27137), .dinb(n27135), .dout(n27138));
  jand g09116(.dina(n27138), .dinb(n26843), .dout(n27139));
  jxor g09117(.dina(n26835), .dinb(n421), .dout(n27140));
  jnot g09118(.din(n27140), .dout(n27141));
  jor  g09119(.dina(n27141), .dinb(n27139), .dout(n27142));
  jand g09120(.dina(n27142), .dinb(n26837), .dout(n27143));
  jxor g09121(.dina(n26829), .dinb(n422), .dout(n27144));
  jnot g09122(.din(n27144), .dout(n27145));
  jor  g09123(.dina(n27145), .dinb(n27143), .dout(n27146));
  jand g09124(.dina(n27146), .dinb(n26831), .dout(n27147));
  jxor g09125(.dina(n26823), .dinb(n416), .dout(n27148));
  jnot g09126(.din(n27148), .dout(n27149));
  jor  g09127(.dina(n27149), .dinb(n27147), .dout(n27150));
  jand g09128(.dina(n27150), .dinb(n26825), .dout(n27151));
  jxor g09129(.dina(n26817), .dinb(n417), .dout(n27152));
  jnot g09130(.din(n27152), .dout(n27153));
  jor  g09131(.dina(n27153), .dinb(n27151), .dout(n27154));
  jand g09132(.dina(n27154), .dinb(n26819), .dout(n27155));
  jxor g09133(.dina(n26811), .dinb(n2547), .dout(n27156));
  jnot g09134(.din(n27156), .dout(n27157));
  jor  g09135(.dina(n27157), .dinb(n27155), .dout(n27158));
  jand g09136(.dina(n27158), .dinb(n26813), .dout(n27159));
  jxor g09137(.dina(n26805), .dinb(n2714), .dout(n27160));
  jnot g09138(.din(n27160), .dout(n27161));
  jor  g09139(.dina(n27161), .dinb(n27159), .dout(n27162));
  jand g09140(.dina(n27162), .dinb(n26807), .dout(n27163));
  jxor g09141(.dina(n26799), .dinb(n405), .dout(n27164));
  jnot g09142(.din(n27164), .dout(n27165));
  jor  g09143(.dina(n27165), .dinb(n27163), .dout(n27166));
  jand g09144(.dina(n27166), .dinb(n26801), .dout(n27167));
  jxor g09145(.dina(n26793), .dinb(n406), .dout(n27168));
  jnot g09146(.din(n27168), .dout(n27169));
  jor  g09147(.dina(n27169), .dinb(n27167), .dout(n27170));
  jand g09148(.dina(n27170), .dinb(n26795), .dout(n27171));
  jxor g09149(.dina(n26787), .dinb(n412), .dout(n27172));
  jnot g09150(.din(n27172), .dout(n27173));
  jor  g09151(.dina(n27173), .dinb(n27171), .dout(n27174));
  jand g09152(.dina(n27174), .dinb(n26789), .dout(n27175));
  jxor g09153(.dina(n26781), .dinb(n413), .dout(n27176));
  jnot g09154(.din(n27176), .dout(n27177));
  jor  g09155(.dina(n27177), .dinb(n27175), .dout(n27178));
  jand g09156(.dina(n27178), .dinb(n26783), .dout(n27179));
  jxor g09157(.dina(n26775), .dinb(n409), .dout(n27180));
  jnot g09158(.din(n27180), .dout(n27181));
  jor  g09159(.dina(n27181), .dinb(n27179), .dout(n27182));
  jand g09160(.dina(n27182), .dinb(n26777), .dout(n27183));
  jxor g09161(.dina(n26769), .dinb(n410), .dout(n27184));
  jnot g09162(.din(n27184), .dout(n27185));
  jor  g09163(.dina(n27185), .dinb(n27183), .dout(n27186));
  jand g09164(.dina(n27186), .dinb(n26771), .dout(n27187));
  jxor g09165(.dina(n26763), .dinb(n426), .dout(n27188));
  jnot g09166(.din(n27188), .dout(n27189));
  jor  g09167(.dina(n27189), .dinb(n27187), .dout(n27190));
  jand g09168(.dina(n27190), .dinb(n26765), .dout(n27191));
  jxor g09169(.dina(n26757), .dinb(n427), .dout(n27192));
  jnot g09170(.din(n27192), .dout(n27193));
  jor  g09171(.dina(n27193), .dinb(n27191), .dout(n27194));
  jand g09172(.dina(n27194), .dinb(n26759), .dout(n27195));
  jxor g09173(.dina(n26751), .dinb(n424), .dout(n27196));
  jnot g09174(.din(n27196), .dout(n27197));
  jor  g09175(.dina(n27197), .dinb(n27195), .dout(n27198));
  jand g09176(.dina(n27198), .dinb(n26753), .dout(n27199));
  jxor g09177(.dina(n26745), .dinb(n300), .dout(n27200));
  jnot g09178(.din(n27200), .dout(n27201));
  jor  g09179(.dina(n27201), .dinb(n27199), .dout(n27202));
  jand g09180(.dina(n27202), .dinb(n26747), .dout(n27203));
  jxor g09181(.dina(n26739), .dinb(n297), .dout(n27204));
  jnot g09182(.din(n27204), .dout(n27205));
  jor  g09183(.dina(n27205), .dinb(n27203), .dout(n27206));
  jand g09184(.dina(n27206), .dinb(n26741), .dout(n27207));
  jxor g09185(.dina(n26733), .dinb(n298), .dout(n27208));
  jnot g09186(.din(n27208), .dout(n27209));
  jor  g09187(.dina(n27209), .dinb(n27207), .dout(n27210));
  jand g09188(.dina(n27210), .dinb(n26735), .dout(n27211));
  jxor g09189(.dina(n26727), .dinb(n301), .dout(n27212));
  jnot g09190(.din(n27212), .dout(n27213));
  jor  g09191(.dina(n27213), .dinb(n27211), .dout(n27214));
  jand g09192(.dina(n27214), .dinb(n26729), .dout(n27215));
  jxor g09193(.dina(n26721), .dinb(n293), .dout(n27216));
  jnot g09194(.din(n27216), .dout(n27217));
  jor  g09195(.dina(n27217), .dinb(n27215), .dout(n27218));
  jand g09196(.dina(n27218), .dinb(n26723), .dout(n27219));
  jnot g09197(.din(n26715), .dout(n27220));
  jand g09198(.dina(n27220), .dinb(b37 ), .dout(n27221));
  jor  g09199(.dina(n27221), .dinb(n27219), .dout(n27222));
  jand g09200(.dina(n27222), .dinb(n26717), .dout(n27223));
  jor  g09201(.dina(n27223), .dinb(n6716), .dout(n27224));
  jand g09202(.dina(n27224), .dinb(n26715), .dout(n27225));
  jnot g09203(.din(n26922), .dout(n27226));
  jnot g09204(.din(n26928), .dout(n27227));
  jnot g09205(.din(n6930), .dout(n27228));
  jor  g09206(.dina(n27074), .dinb(n27228), .dout(n27229));
  jand g09207(.dina(n27229), .dinb(a27 ), .dout(n27230));
  jnot g09208(.din(n27075), .dout(n27231));
  jor  g09209(.dina(n27231), .dinb(n27230), .dout(n27232));
  jand g09210(.dina(n27232), .dinb(n258), .dout(n27233));
  jxor g09211(.dina(n27076), .dinb(b1 ), .dout(n27234));
  jand g09212(.dina(n27234), .dinb(n7091), .dout(n27235));
  jor  g09213(.dina(n27235), .dinb(n27233), .dout(n27236));
  jxor g09214(.dina(n26927), .dinb(b2 ), .dout(n27237));
  jand g09215(.dina(n27237), .dinb(n27236), .dout(n27238));
  jor  g09216(.dina(n27238), .dinb(n27227), .dout(n27239));
  jand g09217(.dina(n27084), .dinb(n27239), .dout(n27240));
  jor  g09218(.dina(n27240), .dinb(n27226), .dout(n27241));
  jand g09219(.dina(n27088), .dinb(n27241), .dout(n27242));
  jor  g09220(.dina(n27242), .dinb(n26914), .dout(n27243));
  jand g09221(.dina(n27092), .dinb(n27243), .dout(n27244));
  jor  g09222(.dina(n27244), .dinb(n26908), .dout(n27245));
  jand g09223(.dina(n27096), .dinb(n27245), .dout(n27246));
  jor  g09224(.dina(n27246), .dinb(n26902), .dout(n27247));
  jand g09225(.dina(n27100), .dinb(n27247), .dout(n27248));
  jor  g09226(.dina(n27248), .dinb(n26896), .dout(n27249));
  jand g09227(.dina(n27104), .dinb(n27249), .dout(n27250));
  jor  g09228(.dina(n27250), .dinb(n26890), .dout(n27251));
  jand g09229(.dina(n27108), .dinb(n27251), .dout(n27252));
  jor  g09230(.dina(n27252), .dinb(n26884), .dout(n27253));
  jand g09231(.dina(n27112), .dinb(n27253), .dout(n27254));
  jor  g09232(.dina(n27254), .dinb(n26878), .dout(n27255));
  jand g09233(.dina(n27116), .dinb(n27255), .dout(n27256));
  jor  g09234(.dina(n27256), .dinb(n26872), .dout(n27257));
  jand g09235(.dina(n27120), .dinb(n27257), .dout(n27258));
  jor  g09236(.dina(n27258), .dinb(n26866), .dout(n27259));
  jand g09237(.dina(n27124), .dinb(n27259), .dout(n27260));
  jor  g09238(.dina(n27260), .dinb(n26860), .dout(n27261));
  jand g09239(.dina(n27128), .dinb(n27261), .dout(n27262));
  jor  g09240(.dina(n27262), .dinb(n26854), .dout(n27263));
  jand g09241(.dina(n27132), .dinb(n27263), .dout(n27264));
  jor  g09242(.dina(n27264), .dinb(n26848), .dout(n27265));
  jand g09243(.dina(n27136), .dinb(n27265), .dout(n27266));
  jor  g09244(.dina(n27266), .dinb(n26842), .dout(n27267));
  jand g09245(.dina(n27140), .dinb(n27267), .dout(n27268));
  jor  g09246(.dina(n27268), .dinb(n26836), .dout(n27269));
  jand g09247(.dina(n27144), .dinb(n27269), .dout(n27270));
  jor  g09248(.dina(n27270), .dinb(n26830), .dout(n27271));
  jand g09249(.dina(n27148), .dinb(n27271), .dout(n27272));
  jor  g09250(.dina(n27272), .dinb(n26824), .dout(n27273));
  jand g09251(.dina(n27152), .dinb(n27273), .dout(n27274));
  jor  g09252(.dina(n27274), .dinb(n26818), .dout(n27275));
  jand g09253(.dina(n27156), .dinb(n27275), .dout(n27276));
  jor  g09254(.dina(n27276), .dinb(n26812), .dout(n27277));
  jand g09255(.dina(n27160), .dinb(n27277), .dout(n27278));
  jor  g09256(.dina(n27278), .dinb(n26806), .dout(n27279));
  jand g09257(.dina(n27164), .dinb(n27279), .dout(n27280));
  jor  g09258(.dina(n27280), .dinb(n26800), .dout(n27281));
  jand g09259(.dina(n27168), .dinb(n27281), .dout(n27282));
  jor  g09260(.dina(n27282), .dinb(n26794), .dout(n27283));
  jand g09261(.dina(n27172), .dinb(n27283), .dout(n27284));
  jor  g09262(.dina(n27284), .dinb(n26788), .dout(n27285));
  jand g09263(.dina(n27176), .dinb(n27285), .dout(n27286));
  jor  g09264(.dina(n27286), .dinb(n26782), .dout(n27287));
  jand g09265(.dina(n27180), .dinb(n27287), .dout(n27288));
  jor  g09266(.dina(n27288), .dinb(n26776), .dout(n27289));
  jand g09267(.dina(n27184), .dinb(n27289), .dout(n27290));
  jor  g09268(.dina(n27290), .dinb(n26770), .dout(n27291));
  jand g09269(.dina(n27188), .dinb(n27291), .dout(n27292));
  jor  g09270(.dina(n27292), .dinb(n26764), .dout(n27293));
  jand g09271(.dina(n27192), .dinb(n27293), .dout(n27294));
  jor  g09272(.dina(n27294), .dinb(n26758), .dout(n27295));
  jand g09273(.dina(n27196), .dinb(n27295), .dout(n27296));
  jor  g09274(.dina(n27296), .dinb(n26752), .dout(n27297));
  jand g09275(.dina(n27200), .dinb(n27297), .dout(n27298));
  jor  g09276(.dina(n27298), .dinb(n26746), .dout(n27299));
  jand g09277(.dina(n27204), .dinb(n27299), .dout(n27300));
  jor  g09278(.dina(n27300), .dinb(n26740), .dout(n27301));
  jand g09279(.dina(n27208), .dinb(n27301), .dout(n27302));
  jor  g09280(.dina(n27302), .dinb(n26734), .dout(n27303));
  jand g09281(.dina(n27212), .dinb(n27303), .dout(n27304));
  jor  g09282(.dina(n27304), .dinb(n26728), .dout(n27305));
  jand g09283(.dina(n27216), .dinb(n27305), .dout(n27306));
  jor  g09284(.dina(n27306), .dinb(n26722), .dout(n27307));
  jand g09285(.dina(n26716), .dinb(n6715), .dout(n27308));
  jand g09286(.dina(n27308), .dinb(n27307), .dout(n27309));
  jor  g09287(.dina(n27309), .dinb(n27225), .dout(n27310));
  jnot g09288(.din(n27310), .dout(n27311));
  jand g09289(.dina(n27224), .dinb(n26721), .dout(n27312));
  jnot g09290(.din(n27221), .dout(n27313));
  jand g09291(.dina(n27313), .dinb(n27307), .dout(n27314));
  jor  g09292(.dina(n27314), .dinb(n26716), .dout(n27315));
  jand g09293(.dina(n27315), .dinb(n6715), .dout(n27316));
  jxor g09294(.dina(n27216), .dinb(n27305), .dout(n27317));
  jand g09295(.dina(n27317), .dinb(n27316), .dout(n27318));
  jor  g09296(.dina(n27318), .dinb(n27312), .dout(n27319));
  jand g09297(.dina(n27319), .dinb(n294), .dout(n27320));
  jnot g09298(.din(n27320), .dout(n27321));
  jand g09299(.dina(n27224), .dinb(n26727), .dout(n27322));
  jxor g09300(.dina(n27212), .dinb(n27303), .dout(n27323));
  jand g09301(.dina(n27323), .dinb(n27316), .dout(n27324));
  jor  g09302(.dina(n27324), .dinb(n27322), .dout(n27325));
  jand g09303(.dina(n27325), .dinb(n293), .dout(n27326));
  jnot g09304(.din(n27326), .dout(n27327));
  jand g09305(.dina(n27224), .dinb(n26733), .dout(n27328));
  jxor g09306(.dina(n27208), .dinb(n27301), .dout(n27329));
  jand g09307(.dina(n27329), .dinb(n27316), .dout(n27330));
  jor  g09308(.dina(n27330), .dinb(n27328), .dout(n27331));
  jand g09309(.dina(n27331), .dinb(n301), .dout(n27332));
  jnot g09310(.din(n27332), .dout(n27333));
  jand g09311(.dina(n27224), .dinb(n26739), .dout(n27334));
  jxor g09312(.dina(n27204), .dinb(n27299), .dout(n27335));
  jand g09313(.dina(n27335), .dinb(n27316), .dout(n27336));
  jor  g09314(.dina(n27336), .dinb(n27334), .dout(n27337));
  jand g09315(.dina(n27337), .dinb(n298), .dout(n27338));
  jnot g09316(.din(n27338), .dout(n27339));
  jand g09317(.dina(n27224), .dinb(n26745), .dout(n27340));
  jxor g09318(.dina(n27200), .dinb(n27297), .dout(n27341));
  jand g09319(.dina(n27341), .dinb(n27316), .dout(n27342));
  jor  g09320(.dina(n27342), .dinb(n27340), .dout(n27343));
  jand g09321(.dina(n27343), .dinb(n297), .dout(n27344));
  jnot g09322(.din(n27344), .dout(n27345));
  jand g09323(.dina(n27224), .dinb(n26751), .dout(n27346));
  jxor g09324(.dina(n27196), .dinb(n27295), .dout(n27347));
  jand g09325(.dina(n27347), .dinb(n27316), .dout(n27348));
  jor  g09326(.dina(n27348), .dinb(n27346), .dout(n27349));
  jand g09327(.dina(n27349), .dinb(n300), .dout(n27350));
  jnot g09328(.din(n27350), .dout(n27351));
  jand g09329(.dina(n27224), .dinb(n26757), .dout(n27352));
  jxor g09330(.dina(n27192), .dinb(n27293), .dout(n27353));
  jand g09331(.dina(n27353), .dinb(n27316), .dout(n27354));
  jor  g09332(.dina(n27354), .dinb(n27352), .dout(n27355));
  jand g09333(.dina(n27355), .dinb(n424), .dout(n27356));
  jnot g09334(.din(n27356), .dout(n27357));
  jand g09335(.dina(n27224), .dinb(n26763), .dout(n27358));
  jxor g09336(.dina(n27188), .dinb(n27291), .dout(n27359));
  jand g09337(.dina(n27359), .dinb(n27316), .dout(n27360));
  jor  g09338(.dina(n27360), .dinb(n27358), .dout(n27361));
  jand g09339(.dina(n27361), .dinb(n427), .dout(n27362));
  jnot g09340(.din(n27362), .dout(n27363));
  jand g09341(.dina(n27224), .dinb(n26769), .dout(n27364));
  jxor g09342(.dina(n27184), .dinb(n27289), .dout(n27365));
  jand g09343(.dina(n27365), .dinb(n27316), .dout(n27366));
  jor  g09344(.dina(n27366), .dinb(n27364), .dout(n27367));
  jand g09345(.dina(n27367), .dinb(n426), .dout(n27368));
  jnot g09346(.din(n27368), .dout(n27369));
  jand g09347(.dina(n27224), .dinb(n26775), .dout(n27370));
  jxor g09348(.dina(n27180), .dinb(n27287), .dout(n27371));
  jand g09349(.dina(n27371), .dinb(n27316), .dout(n27372));
  jor  g09350(.dina(n27372), .dinb(n27370), .dout(n27373));
  jand g09351(.dina(n27373), .dinb(n410), .dout(n27374));
  jnot g09352(.din(n27374), .dout(n27375));
  jand g09353(.dina(n27224), .dinb(n26781), .dout(n27376));
  jxor g09354(.dina(n27176), .dinb(n27285), .dout(n27377));
  jand g09355(.dina(n27377), .dinb(n27316), .dout(n27378));
  jor  g09356(.dina(n27378), .dinb(n27376), .dout(n27379));
  jand g09357(.dina(n27379), .dinb(n409), .dout(n27380));
  jnot g09358(.din(n27380), .dout(n27381));
  jand g09359(.dina(n27224), .dinb(n26787), .dout(n27382));
  jxor g09360(.dina(n27172), .dinb(n27283), .dout(n27383));
  jand g09361(.dina(n27383), .dinb(n27316), .dout(n27384));
  jor  g09362(.dina(n27384), .dinb(n27382), .dout(n27385));
  jand g09363(.dina(n27385), .dinb(n413), .dout(n27386));
  jnot g09364(.din(n27386), .dout(n27387));
  jand g09365(.dina(n27224), .dinb(n26793), .dout(n27388));
  jxor g09366(.dina(n27168), .dinb(n27281), .dout(n27389));
  jand g09367(.dina(n27389), .dinb(n27316), .dout(n27390));
  jor  g09368(.dina(n27390), .dinb(n27388), .dout(n27391));
  jand g09369(.dina(n27391), .dinb(n412), .dout(n27392));
  jnot g09370(.din(n27392), .dout(n27393));
  jand g09371(.dina(n27224), .dinb(n26799), .dout(n27394));
  jxor g09372(.dina(n27164), .dinb(n27279), .dout(n27395));
  jand g09373(.dina(n27395), .dinb(n27316), .dout(n27396));
  jor  g09374(.dina(n27396), .dinb(n27394), .dout(n27397));
  jand g09375(.dina(n27397), .dinb(n406), .dout(n27398));
  jnot g09376(.din(n27398), .dout(n27399));
  jand g09377(.dina(n27224), .dinb(n26805), .dout(n27400));
  jxor g09378(.dina(n27160), .dinb(n27277), .dout(n27401));
  jand g09379(.dina(n27401), .dinb(n27316), .dout(n27402));
  jor  g09380(.dina(n27402), .dinb(n27400), .dout(n27403));
  jand g09381(.dina(n27403), .dinb(n405), .dout(n27404));
  jnot g09382(.din(n27404), .dout(n27405));
  jand g09383(.dina(n27224), .dinb(n26811), .dout(n27406));
  jxor g09384(.dina(n27156), .dinb(n27275), .dout(n27407));
  jand g09385(.dina(n27407), .dinb(n27316), .dout(n27408));
  jor  g09386(.dina(n27408), .dinb(n27406), .dout(n27409));
  jand g09387(.dina(n27409), .dinb(n2714), .dout(n27410));
  jnot g09388(.din(n27410), .dout(n27411));
  jand g09389(.dina(n27224), .dinb(n26817), .dout(n27412));
  jxor g09390(.dina(n27152), .dinb(n27273), .dout(n27413));
  jand g09391(.dina(n27413), .dinb(n27316), .dout(n27414));
  jor  g09392(.dina(n27414), .dinb(n27412), .dout(n27415));
  jand g09393(.dina(n27415), .dinb(n2547), .dout(n27416));
  jnot g09394(.din(n27416), .dout(n27417));
  jand g09395(.dina(n27224), .dinb(n26823), .dout(n27418));
  jxor g09396(.dina(n27148), .dinb(n27271), .dout(n27419));
  jand g09397(.dina(n27419), .dinb(n27316), .dout(n27420));
  jor  g09398(.dina(n27420), .dinb(n27418), .dout(n27421));
  jand g09399(.dina(n27421), .dinb(n417), .dout(n27422));
  jnot g09400(.din(n27422), .dout(n27423));
  jand g09401(.dina(n27224), .dinb(n26829), .dout(n27424));
  jxor g09402(.dina(n27144), .dinb(n27269), .dout(n27425));
  jand g09403(.dina(n27425), .dinb(n27316), .dout(n27426));
  jor  g09404(.dina(n27426), .dinb(n27424), .dout(n27427));
  jand g09405(.dina(n27427), .dinb(n416), .dout(n27428));
  jnot g09406(.din(n27428), .dout(n27429));
  jand g09407(.dina(n27224), .dinb(n26835), .dout(n27430));
  jxor g09408(.dina(n27140), .dinb(n27267), .dout(n27431));
  jand g09409(.dina(n27431), .dinb(n27316), .dout(n27432));
  jor  g09410(.dina(n27432), .dinb(n27430), .dout(n27433));
  jand g09411(.dina(n27433), .dinb(n422), .dout(n27434));
  jnot g09412(.din(n27434), .dout(n27435));
  jand g09413(.dina(n27224), .dinb(n26841), .dout(n27436));
  jxor g09414(.dina(n27136), .dinb(n27265), .dout(n27437));
  jand g09415(.dina(n27437), .dinb(n27316), .dout(n27438));
  jor  g09416(.dina(n27438), .dinb(n27436), .dout(n27439));
  jand g09417(.dina(n27439), .dinb(n421), .dout(n27440));
  jnot g09418(.din(n27440), .dout(n27441));
  jand g09419(.dina(n27224), .dinb(n26847), .dout(n27442));
  jxor g09420(.dina(n27132), .dinb(n27263), .dout(n27443));
  jand g09421(.dina(n27443), .dinb(n27316), .dout(n27444));
  jor  g09422(.dina(n27444), .dinb(n27442), .dout(n27445));
  jand g09423(.dina(n27445), .dinb(n433), .dout(n27446));
  jnot g09424(.din(n27446), .dout(n27447));
  jand g09425(.dina(n27224), .dinb(n26853), .dout(n27448));
  jxor g09426(.dina(n27128), .dinb(n27261), .dout(n27449));
  jand g09427(.dina(n27449), .dinb(n27316), .dout(n27450));
  jor  g09428(.dina(n27450), .dinb(n27448), .dout(n27451));
  jand g09429(.dina(n27451), .dinb(n432), .dout(n27452));
  jnot g09430(.din(n27452), .dout(n27453));
  jand g09431(.dina(n27224), .dinb(n26859), .dout(n27454));
  jxor g09432(.dina(n27124), .dinb(n27259), .dout(n27455));
  jand g09433(.dina(n27455), .dinb(n27316), .dout(n27456));
  jor  g09434(.dina(n27456), .dinb(n27454), .dout(n27457));
  jand g09435(.dina(n27457), .dinb(n436), .dout(n27458));
  jnot g09436(.din(n27458), .dout(n27459));
  jand g09437(.dina(n27224), .dinb(n26865), .dout(n27460));
  jxor g09438(.dina(n27120), .dinb(n27257), .dout(n27461));
  jand g09439(.dina(n27461), .dinb(n27316), .dout(n27462));
  jor  g09440(.dina(n27462), .dinb(n27460), .dout(n27463));
  jand g09441(.dina(n27463), .dinb(n435), .dout(n27464));
  jnot g09442(.din(n27464), .dout(n27465));
  jand g09443(.dina(n27224), .dinb(n26871), .dout(n27466));
  jxor g09444(.dina(n27116), .dinb(n27255), .dout(n27467));
  jand g09445(.dina(n27467), .dinb(n27316), .dout(n27468));
  jor  g09446(.dina(n27468), .dinb(n27466), .dout(n27469));
  jand g09447(.dina(n27469), .dinb(n440), .dout(n27470));
  jnot g09448(.din(n27470), .dout(n27471));
  jand g09449(.dina(n27224), .dinb(n26877), .dout(n27472));
  jxor g09450(.dina(n27112), .dinb(n27253), .dout(n27473));
  jand g09451(.dina(n27473), .dinb(n27316), .dout(n27474));
  jor  g09452(.dina(n27474), .dinb(n27472), .dout(n27475));
  jand g09453(.dina(n27475), .dinb(n439), .dout(n27476));
  jnot g09454(.din(n27476), .dout(n27477));
  jand g09455(.dina(n27224), .dinb(n26883), .dout(n27478));
  jxor g09456(.dina(n27108), .dinb(n27251), .dout(n27479));
  jand g09457(.dina(n27479), .dinb(n27316), .dout(n27480));
  jor  g09458(.dina(n27480), .dinb(n27478), .dout(n27481));
  jand g09459(.dina(n27481), .dinb(n325), .dout(n27482));
  jnot g09460(.din(n27482), .dout(n27483));
  jand g09461(.dina(n27224), .dinb(n26889), .dout(n27484));
  jxor g09462(.dina(n27104), .dinb(n27249), .dout(n27485));
  jand g09463(.dina(n27485), .dinb(n27316), .dout(n27486));
  jor  g09464(.dina(n27486), .dinb(n27484), .dout(n27487));
  jand g09465(.dina(n27487), .dinb(n324), .dout(n27488));
  jnot g09466(.din(n27488), .dout(n27489));
  jand g09467(.dina(n27224), .dinb(n26895), .dout(n27490));
  jxor g09468(.dina(n27100), .dinb(n27247), .dout(n27491));
  jand g09469(.dina(n27491), .dinb(n27316), .dout(n27492));
  jor  g09470(.dina(n27492), .dinb(n27490), .dout(n27493));
  jand g09471(.dina(n27493), .dinb(n323), .dout(n27494));
  jnot g09472(.din(n27494), .dout(n27495));
  jand g09473(.dina(n27224), .dinb(n26901), .dout(n27496));
  jxor g09474(.dina(n27096), .dinb(n27245), .dout(n27497));
  jand g09475(.dina(n27497), .dinb(n27316), .dout(n27498));
  jor  g09476(.dina(n27498), .dinb(n27496), .dout(n27499));
  jand g09477(.dina(n27499), .dinb(n335), .dout(n27500));
  jnot g09478(.din(n27500), .dout(n27501));
  jand g09479(.dina(n27224), .dinb(n26907), .dout(n27502));
  jxor g09480(.dina(n27092), .dinb(n27243), .dout(n27503));
  jand g09481(.dina(n27503), .dinb(n27316), .dout(n27504));
  jor  g09482(.dina(n27504), .dinb(n27502), .dout(n27505));
  jand g09483(.dina(n27505), .dinb(n334), .dout(n27506));
  jnot g09484(.din(n27506), .dout(n27507));
  jand g09485(.dina(n27224), .dinb(n26913), .dout(n27508));
  jxor g09486(.dina(n27088), .dinb(n27241), .dout(n27509));
  jand g09487(.dina(n27509), .dinb(n27316), .dout(n27510));
  jor  g09488(.dina(n27510), .dinb(n27508), .dout(n27511));
  jand g09489(.dina(n27511), .dinb(n338), .dout(n27512));
  jnot g09490(.din(n27512), .dout(n27513));
  jor  g09491(.dina(n27316), .dinb(n26921), .dout(n27514));
  jxor g09492(.dina(n27084), .dinb(n27239), .dout(n27515));
  jand g09493(.dina(n27515), .dinb(n27316), .dout(n27516));
  jnot g09494(.din(n27516), .dout(n27517));
  jand g09495(.dina(n27517), .dinb(n27514), .dout(n27518));
  jnot g09496(.din(n27518), .dout(n27519));
  jand g09497(.dina(n27519), .dinb(n337), .dout(n27520));
  jnot g09498(.din(n27520), .dout(n27521));
  jor  g09499(.dina(n27316), .dinb(n26927), .dout(n27522));
  jxor g09500(.dina(n27237), .dinb(n27236), .dout(n27523));
  jnot g09501(.din(n27523), .dout(n27524));
  jor  g09502(.dina(n27524), .dinb(n27224), .dout(n27525));
  jand g09503(.dina(n27525), .dinb(n27522), .dout(n27526));
  jnot g09504(.din(n27526), .dout(n27527));
  jand g09505(.dina(n27527), .dinb(n344), .dout(n27528));
  jnot g09506(.din(n27528), .dout(n27529));
  jand g09507(.dina(n27224), .dinb(n27232), .dout(n27530));
  jxor g09508(.dina(n27234), .dinb(n7091), .dout(n27531));
  jand g09509(.dina(n27531), .dinb(n27316), .dout(n27532));
  jor  g09510(.dina(n27532), .dinb(n27530), .dout(n27533));
  jand g09511(.dina(n27533), .dinb(n348), .dout(n27534));
  jnot g09512(.din(n27534), .dout(n27535));
  jnot g09513(.din(n7356), .dout(n27536));
  jor  g09514(.dina(n27223), .dinb(n27536), .dout(n27537));
  jand g09515(.dina(n27537), .dinb(a26 ), .dout(n27538));
  jand g09516(.dina(n27316), .dinb(n6939), .dout(n27539));
  jor  g09517(.dina(n27539), .dinb(n27538), .dout(n27540));
  jand g09518(.dina(n27540), .dinb(n258), .dout(n27541));
  jnot g09519(.din(n27541), .dout(n27542));
  jand g09520(.dina(n27315), .dinb(n7356), .dout(n27543));
  jor  g09521(.dina(n27543), .dinb(n6938), .dout(n27544));
  jor  g09522(.dina(n27224), .dinb(n7091), .dout(n27545));
  jand g09523(.dina(n27545), .dinb(n27544), .dout(n27546));
  jxor g09524(.dina(n27546), .dinb(n258), .dout(n27547));
  jor  g09525(.dina(n27547), .dinb(n7364), .dout(n27548));
  jand g09526(.dina(n27548), .dinb(n27542), .dout(n27549));
  jxor g09527(.dina(n27533), .dinb(n348), .dout(n27550));
  jnot g09528(.din(n27550), .dout(n27551));
  jor  g09529(.dina(n27551), .dinb(n27549), .dout(n27552));
  jand g09530(.dina(n27552), .dinb(n27535), .dout(n27553));
  jxor g09531(.dina(n27526), .dinb(b3 ), .dout(n27554));
  jnot g09532(.din(n27554), .dout(n27555));
  jor  g09533(.dina(n27555), .dinb(n27553), .dout(n27556));
  jand g09534(.dina(n27556), .dinb(n27529), .dout(n27557));
  jxor g09535(.dina(n27518), .dinb(b4 ), .dout(n27558));
  jnot g09536(.din(n27558), .dout(n27559));
  jor  g09537(.dina(n27559), .dinb(n27557), .dout(n27560));
  jand g09538(.dina(n27560), .dinb(n27521), .dout(n27561));
  jxor g09539(.dina(n27511), .dinb(n338), .dout(n27562));
  jnot g09540(.din(n27562), .dout(n27563));
  jor  g09541(.dina(n27563), .dinb(n27561), .dout(n27564));
  jand g09542(.dina(n27564), .dinb(n27513), .dout(n27565));
  jxor g09543(.dina(n27505), .dinb(n334), .dout(n27566));
  jnot g09544(.din(n27566), .dout(n27567));
  jor  g09545(.dina(n27567), .dinb(n27565), .dout(n27568));
  jand g09546(.dina(n27568), .dinb(n27507), .dout(n27569));
  jxor g09547(.dina(n27499), .dinb(n335), .dout(n27570));
  jnot g09548(.din(n27570), .dout(n27571));
  jor  g09549(.dina(n27571), .dinb(n27569), .dout(n27572));
  jand g09550(.dina(n27572), .dinb(n27501), .dout(n27573));
  jxor g09551(.dina(n27493), .dinb(n323), .dout(n27574));
  jnot g09552(.din(n27574), .dout(n27575));
  jor  g09553(.dina(n27575), .dinb(n27573), .dout(n27576));
  jand g09554(.dina(n27576), .dinb(n27495), .dout(n27577));
  jxor g09555(.dina(n27487), .dinb(n324), .dout(n27578));
  jnot g09556(.din(n27578), .dout(n27579));
  jor  g09557(.dina(n27579), .dinb(n27577), .dout(n27580));
  jand g09558(.dina(n27580), .dinb(n27489), .dout(n27581));
  jxor g09559(.dina(n27481), .dinb(n325), .dout(n27582));
  jnot g09560(.din(n27582), .dout(n27583));
  jor  g09561(.dina(n27583), .dinb(n27581), .dout(n27584));
  jand g09562(.dina(n27584), .dinb(n27483), .dout(n27585));
  jxor g09563(.dina(n27475), .dinb(n439), .dout(n27586));
  jnot g09564(.din(n27586), .dout(n27587));
  jor  g09565(.dina(n27587), .dinb(n27585), .dout(n27588));
  jand g09566(.dina(n27588), .dinb(n27477), .dout(n27589));
  jxor g09567(.dina(n27469), .dinb(n440), .dout(n27590));
  jnot g09568(.din(n27590), .dout(n27591));
  jor  g09569(.dina(n27591), .dinb(n27589), .dout(n27592));
  jand g09570(.dina(n27592), .dinb(n27471), .dout(n27593));
  jxor g09571(.dina(n27463), .dinb(n435), .dout(n27594));
  jnot g09572(.din(n27594), .dout(n27595));
  jor  g09573(.dina(n27595), .dinb(n27593), .dout(n27596));
  jand g09574(.dina(n27596), .dinb(n27465), .dout(n27597));
  jxor g09575(.dina(n27457), .dinb(n436), .dout(n27598));
  jnot g09576(.din(n27598), .dout(n27599));
  jor  g09577(.dina(n27599), .dinb(n27597), .dout(n27600));
  jand g09578(.dina(n27600), .dinb(n27459), .dout(n27601));
  jxor g09579(.dina(n27451), .dinb(n432), .dout(n27602));
  jnot g09580(.din(n27602), .dout(n27603));
  jor  g09581(.dina(n27603), .dinb(n27601), .dout(n27604));
  jand g09582(.dina(n27604), .dinb(n27453), .dout(n27605));
  jxor g09583(.dina(n27445), .dinb(n433), .dout(n27606));
  jnot g09584(.din(n27606), .dout(n27607));
  jor  g09585(.dina(n27607), .dinb(n27605), .dout(n27608));
  jand g09586(.dina(n27608), .dinb(n27447), .dout(n27609));
  jxor g09587(.dina(n27439), .dinb(n421), .dout(n27610));
  jnot g09588(.din(n27610), .dout(n27611));
  jor  g09589(.dina(n27611), .dinb(n27609), .dout(n27612));
  jand g09590(.dina(n27612), .dinb(n27441), .dout(n27613));
  jxor g09591(.dina(n27433), .dinb(n422), .dout(n27614));
  jnot g09592(.din(n27614), .dout(n27615));
  jor  g09593(.dina(n27615), .dinb(n27613), .dout(n27616));
  jand g09594(.dina(n27616), .dinb(n27435), .dout(n27617));
  jxor g09595(.dina(n27427), .dinb(n416), .dout(n27618));
  jnot g09596(.din(n27618), .dout(n27619));
  jor  g09597(.dina(n27619), .dinb(n27617), .dout(n27620));
  jand g09598(.dina(n27620), .dinb(n27429), .dout(n27621));
  jxor g09599(.dina(n27421), .dinb(n417), .dout(n27622));
  jnot g09600(.din(n27622), .dout(n27623));
  jor  g09601(.dina(n27623), .dinb(n27621), .dout(n27624));
  jand g09602(.dina(n27624), .dinb(n27423), .dout(n27625));
  jxor g09603(.dina(n27415), .dinb(n2547), .dout(n27626));
  jnot g09604(.din(n27626), .dout(n27627));
  jor  g09605(.dina(n27627), .dinb(n27625), .dout(n27628));
  jand g09606(.dina(n27628), .dinb(n27417), .dout(n27629));
  jxor g09607(.dina(n27409), .dinb(n2714), .dout(n27630));
  jnot g09608(.din(n27630), .dout(n27631));
  jor  g09609(.dina(n27631), .dinb(n27629), .dout(n27632));
  jand g09610(.dina(n27632), .dinb(n27411), .dout(n27633));
  jxor g09611(.dina(n27403), .dinb(n405), .dout(n27634));
  jnot g09612(.din(n27634), .dout(n27635));
  jor  g09613(.dina(n27635), .dinb(n27633), .dout(n27636));
  jand g09614(.dina(n27636), .dinb(n27405), .dout(n27637));
  jxor g09615(.dina(n27397), .dinb(n406), .dout(n27638));
  jnot g09616(.din(n27638), .dout(n27639));
  jor  g09617(.dina(n27639), .dinb(n27637), .dout(n27640));
  jand g09618(.dina(n27640), .dinb(n27399), .dout(n27641));
  jxor g09619(.dina(n27391), .dinb(n412), .dout(n27642));
  jnot g09620(.din(n27642), .dout(n27643));
  jor  g09621(.dina(n27643), .dinb(n27641), .dout(n27644));
  jand g09622(.dina(n27644), .dinb(n27393), .dout(n27645));
  jxor g09623(.dina(n27385), .dinb(n413), .dout(n27646));
  jnot g09624(.din(n27646), .dout(n27647));
  jor  g09625(.dina(n27647), .dinb(n27645), .dout(n27648));
  jand g09626(.dina(n27648), .dinb(n27387), .dout(n27649));
  jxor g09627(.dina(n27379), .dinb(n409), .dout(n27650));
  jnot g09628(.din(n27650), .dout(n27651));
  jor  g09629(.dina(n27651), .dinb(n27649), .dout(n27652));
  jand g09630(.dina(n27652), .dinb(n27381), .dout(n27653));
  jxor g09631(.dina(n27373), .dinb(n410), .dout(n27654));
  jnot g09632(.din(n27654), .dout(n27655));
  jor  g09633(.dina(n27655), .dinb(n27653), .dout(n27656));
  jand g09634(.dina(n27656), .dinb(n27375), .dout(n27657));
  jxor g09635(.dina(n27367), .dinb(n426), .dout(n27658));
  jnot g09636(.din(n27658), .dout(n27659));
  jor  g09637(.dina(n27659), .dinb(n27657), .dout(n27660));
  jand g09638(.dina(n27660), .dinb(n27369), .dout(n27661));
  jxor g09639(.dina(n27361), .dinb(n427), .dout(n27662));
  jnot g09640(.din(n27662), .dout(n27663));
  jor  g09641(.dina(n27663), .dinb(n27661), .dout(n27664));
  jand g09642(.dina(n27664), .dinb(n27363), .dout(n27665));
  jxor g09643(.dina(n27355), .dinb(n424), .dout(n27666));
  jnot g09644(.din(n27666), .dout(n27667));
  jor  g09645(.dina(n27667), .dinb(n27665), .dout(n27668));
  jand g09646(.dina(n27668), .dinb(n27357), .dout(n27669));
  jxor g09647(.dina(n27349), .dinb(n300), .dout(n27670));
  jnot g09648(.din(n27670), .dout(n27671));
  jor  g09649(.dina(n27671), .dinb(n27669), .dout(n27672));
  jand g09650(.dina(n27672), .dinb(n27351), .dout(n27673));
  jxor g09651(.dina(n27343), .dinb(n297), .dout(n27674));
  jnot g09652(.din(n27674), .dout(n27675));
  jor  g09653(.dina(n27675), .dinb(n27673), .dout(n27676));
  jand g09654(.dina(n27676), .dinb(n27345), .dout(n27677));
  jxor g09655(.dina(n27337), .dinb(n298), .dout(n27678));
  jnot g09656(.din(n27678), .dout(n27679));
  jor  g09657(.dina(n27679), .dinb(n27677), .dout(n27680));
  jand g09658(.dina(n27680), .dinb(n27339), .dout(n27681));
  jxor g09659(.dina(n27331), .dinb(n301), .dout(n27682));
  jnot g09660(.din(n27682), .dout(n27683));
  jor  g09661(.dina(n27683), .dinb(n27681), .dout(n27684));
  jand g09662(.dina(n27684), .dinb(n27333), .dout(n27685));
  jxor g09663(.dina(n27325), .dinb(n293), .dout(n27686));
  jnot g09664(.din(n27686), .dout(n27687));
  jor  g09665(.dina(n27687), .dinb(n27685), .dout(n27688));
  jand g09666(.dina(n27688), .dinb(n27327), .dout(n27689));
  jxor g09667(.dina(n27319), .dinb(n294), .dout(n27690));
  jnot g09668(.din(n27690), .dout(n27691));
  jor  g09669(.dina(n27691), .dinb(n27689), .dout(n27692));
  jand g09670(.dina(n27692), .dinb(n27321), .dout(n27693));
  jnot g09671(.din(n5701), .dout(n27694));
  jxor g09672(.dina(n27310), .dinb(b38 ), .dout(n27695));
  jor  g09673(.dina(n27695), .dinb(n27694), .dout(n27696));
  jor  g09674(.dina(n27696), .dinb(n27693), .dout(n27697));
  jand g09675(.dina(n27697), .dinb(n27311), .dout(n27698));
  jxor g09676(.dina(n27546), .dinb(b1 ), .dout(n27699));
  jand g09677(.dina(n27699), .dinb(n7365), .dout(n27700));
  jor  g09678(.dina(n27700), .dinb(n27541), .dout(n27701));
  jand g09679(.dina(n27550), .dinb(n27701), .dout(n27702));
  jor  g09680(.dina(n27702), .dinb(n27534), .dout(n27703));
  jand g09681(.dina(n27554), .dinb(n27703), .dout(n27704));
  jor  g09682(.dina(n27704), .dinb(n27528), .dout(n27705));
  jand g09683(.dina(n27558), .dinb(n27705), .dout(n27706));
  jor  g09684(.dina(n27706), .dinb(n27520), .dout(n27707));
  jand g09685(.dina(n27562), .dinb(n27707), .dout(n27708));
  jor  g09686(.dina(n27708), .dinb(n27512), .dout(n27709));
  jand g09687(.dina(n27566), .dinb(n27709), .dout(n27710));
  jor  g09688(.dina(n27710), .dinb(n27506), .dout(n27711));
  jand g09689(.dina(n27570), .dinb(n27711), .dout(n27712));
  jor  g09690(.dina(n27712), .dinb(n27500), .dout(n27713));
  jand g09691(.dina(n27574), .dinb(n27713), .dout(n27714));
  jor  g09692(.dina(n27714), .dinb(n27494), .dout(n27715));
  jand g09693(.dina(n27578), .dinb(n27715), .dout(n27716));
  jor  g09694(.dina(n27716), .dinb(n27488), .dout(n27717));
  jand g09695(.dina(n27582), .dinb(n27717), .dout(n27718));
  jor  g09696(.dina(n27718), .dinb(n27482), .dout(n27719));
  jand g09697(.dina(n27586), .dinb(n27719), .dout(n27720));
  jor  g09698(.dina(n27720), .dinb(n27476), .dout(n27721));
  jand g09699(.dina(n27590), .dinb(n27721), .dout(n27722));
  jor  g09700(.dina(n27722), .dinb(n27470), .dout(n27723));
  jand g09701(.dina(n27594), .dinb(n27723), .dout(n27724));
  jor  g09702(.dina(n27724), .dinb(n27464), .dout(n27725));
  jand g09703(.dina(n27598), .dinb(n27725), .dout(n27726));
  jor  g09704(.dina(n27726), .dinb(n27458), .dout(n27727));
  jand g09705(.dina(n27602), .dinb(n27727), .dout(n27728));
  jor  g09706(.dina(n27728), .dinb(n27452), .dout(n27729));
  jand g09707(.dina(n27606), .dinb(n27729), .dout(n27730));
  jor  g09708(.dina(n27730), .dinb(n27446), .dout(n27731));
  jand g09709(.dina(n27610), .dinb(n27731), .dout(n27732));
  jor  g09710(.dina(n27732), .dinb(n27440), .dout(n27733));
  jand g09711(.dina(n27614), .dinb(n27733), .dout(n27734));
  jor  g09712(.dina(n27734), .dinb(n27434), .dout(n27735));
  jand g09713(.dina(n27618), .dinb(n27735), .dout(n27736));
  jor  g09714(.dina(n27736), .dinb(n27428), .dout(n27737));
  jand g09715(.dina(n27622), .dinb(n27737), .dout(n27738));
  jor  g09716(.dina(n27738), .dinb(n27422), .dout(n27739));
  jand g09717(.dina(n27626), .dinb(n27739), .dout(n27740));
  jor  g09718(.dina(n27740), .dinb(n27416), .dout(n27741));
  jand g09719(.dina(n27630), .dinb(n27741), .dout(n27742));
  jor  g09720(.dina(n27742), .dinb(n27410), .dout(n27743));
  jand g09721(.dina(n27634), .dinb(n27743), .dout(n27744));
  jor  g09722(.dina(n27744), .dinb(n27404), .dout(n27745));
  jand g09723(.dina(n27638), .dinb(n27745), .dout(n27746));
  jor  g09724(.dina(n27746), .dinb(n27398), .dout(n27747));
  jand g09725(.dina(n27642), .dinb(n27747), .dout(n27748));
  jor  g09726(.dina(n27748), .dinb(n27392), .dout(n27749));
  jand g09727(.dina(n27646), .dinb(n27749), .dout(n27750));
  jor  g09728(.dina(n27750), .dinb(n27386), .dout(n27751));
  jand g09729(.dina(n27650), .dinb(n27751), .dout(n27752));
  jor  g09730(.dina(n27752), .dinb(n27380), .dout(n27753));
  jand g09731(.dina(n27654), .dinb(n27753), .dout(n27754));
  jor  g09732(.dina(n27754), .dinb(n27374), .dout(n27755));
  jand g09733(.dina(n27658), .dinb(n27755), .dout(n27756));
  jor  g09734(.dina(n27756), .dinb(n27368), .dout(n27757));
  jand g09735(.dina(n27662), .dinb(n27757), .dout(n27758));
  jor  g09736(.dina(n27758), .dinb(n27362), .dout(n27759));
  jand g09737(.dina(n27666), .dinb(n27759), .dout(n27760));
  jor  g09738(.dina(n27760), .dinb(n27356), .dout(n27761));
  jand g09739(.dina(n27670), .dinb(n27761), .dout(n27762));
  jor  g09740(.dina(n27762), .dinb(n27350), .dout(n27763));
  jand g09741(.dina(n27674), .dinb(n27763), .dout(n27764));
  jor  g09742(.dina(n27764), .dinb(n27344), .dout(n27765));
  jand g09743(.dina(n27678), .dinb(n27765), .dout(n27766));
  jor  g09744(.dina(n27766), .dinb(n27338), .dout(n27767));
  jand g09745(.dina(n27682), .dinb(n27767), .dout(n27768));
  jor  g09746(.dina(n27768), .dinb(n27332), .dout(n27769));
  jand g09747(.dina(n27686), .dinb(n27769), .dout(n27770));
  jor  g09748(.dina(n27770), .dinb(n27326), .dout(n27771));
  jand g09749(.dina(n27690), .dinb(n27771), .dout(n27772));
  jor  g09750(.dina(n27772), .dinb(n27320), .dout(n27773));
  jnot g09751(.din(n27696), .dout(n27774));
  jand g09752(.dina(n27774), .dinb(n27773), .dout(n27775));
  jand g09753(.dina(n27310), .dinb(n6715), .dout(n27776));
  jor  g09754(.dina(n27776), .dinb(n27775), .dout(n27777));
  jxor g09755(.dina(n27695), .dinb(n27773), .dout(n27778));
  jand g09756(.dina(n27778), .dinb(n27777), .dout(n27779));
  jor  g09757(.dina(n27779), .dinb(n27698), .dout(n27780));
  jnot g09758(.din(n27780), .dout(n27781));
  jand g09759(.dina(n27780), .dinb(b39 ), .dout(n27782));
  jand g09760(.dina(n27781), .dinb(n291), .dout(n27783));
  jnot g09761(.din(n27783), .dout(n27784));
  jnot g09762(.din(n27776), .dout(n27785));
  jand g09763(.dina(n27785), .dinb(n27697), .dout(n27786));
  jand g09764(.dina(n27786), .dinb(n27319), .dout(n27787));
  jxor g09765(.dina(n27690), .dinb(n27771), .dout(n27788));
  jand g09766(.dina(n27788), .dinb(n27777), .dout(n27789));
  jor  g09767(.dina(n27789), .dinb(n27787), .dout(n27790));
  jand g09768(.dina(n27790), .dinb(n290), .dout(n27791));
  jnot g09769(.din(n27791), .dout(n27792));
  jand g09770(.dina(n27786), .dinb(n27325), .dout(n27793));
  jxor g09771(.dina(n27686), .dinb(n27769), .dout(n27794));
  jand g09772(.dina(n27794), .dinb(n27777), .dout(n27795));
  jor  g09773(.dina(n27795), .dinb(n27793), .dout(n27796));
  jand g09774(.dina(n27796), .dinb(n294), .dout(n27797));
  jnot g09775(.din(n27797), .dout(n27798));
  jand g09776(.dina(n27786), .dinb(n27331), .dout(n27799));
  jxor g09777(.dina(n27682), .dinb(n27767), .dout(n27800));
  jand g09778(.dina(n27800), .dinb(n27777), .dout(n27801));
  jor  g09779(.dina(n27801), .dinb(n27799), .dout(n27802));
  jand g09780(.dina(n27802), .dinb(n293), .dout(n27803));
  jnot g09781(.din(n27803), .dout(n27804));
  jand g09782(.dina(n27786), .dinb(n27337), .dout(n27805));
  jxor g09783(.dina(n27678), .dinb(n27765), .dout(n27806));
  jand g09784(.dina(n27806), .dinb(n27777), .dout(n27807));
  jor  g09785(.dina(n27807), .dinb(n27805), .dout(n27808));
  jand g09786(.dina(n27808), .dinb(n301), .dout(n27809));
  jnot g09787(.din(n27809), .dout(n27810));
  jand g09788(.dina(n27786), .dinb(n27343), .dout(n27811));
  jxor g09789(.dina(n27674), .dinb(n27763), .dout(n27812));
  jand g09790(.dina(n27812), .dinb(n27777), .dout(n27813));
  jor  g09791(.dina(n27813), .dinb(n27811), .dout(n27814));
  jand g09792(.dina(n27814), .dinb(n298), .dout(n27815));
  jnot g09793(.din(n27815), .dout(n27816));
  jand g09794(.dina(n27786), .dinb(n27349), .dout(n27817));
  jxor g09795(.dina(n27670), .dinb(n27761), .dout(n27818));
  jand g09796(.dina(n27818), .dinb(n27777), .dout(n27819));
  jor  g09797(.dina(n27819), .dinb(n27817), .dout(n27820));
  jand g09798(.dina(n27820), .dinb(n297), .dout(n27821));
  jnot g09799(.din(n27821), .dout(n27822));
  jand g09800(.dina(n27786), .dinb(n27355), .dout(n27823));
  jxor g09801(.dina(n27666), .dinb(n27759), .dout(n27824));
  jand g09802(.dina(n27824), .dinb(n27777), .dout(n27825));
  jor  g09803(.dina(n27825), .dinb(n27823), .dout(n27826));
  jand g09804(.dina(n27826), .dinb(n300), .dout(n27827));
  jnot g09805(.din(n27827), .dout(n27828));
  jand g09806(.dina(n27786), .dinb(n27361), .dout(n27829));
  jxor g09807(.dina(n27662), .dinb(n27757), .dout(n27830));
  jand g09808(.dina(n27830), .dinb(n27777), .dout(n27831));
  jor  g09809(.dina(n27831), .dinb(n27829), .dout(n27832));
  jand g09810(.dina(n27832), .dinb(n424), .dout(n27833));
  jnot g09811(.din(n27833), .dout(n27834));
  jand g09812(.dina(n27786), .dinb(n27367), .dout(n27835));
  jxor g09813(.dina(n27658), .dinb(n27755), .dout(n27836));
  jand g09814(.dina(n27836), .dinb(n27777), .dout(n27837));
  jor  g09815(.dina(n27837), .dinb(n27835), .dout(n27838));
  jand g09816(.dina(n27838), .dinb(n427), .dout(n27839));
  jnot g09817(.din(n27839), .dout(n27840));
  jand g09818(.dina(n27786), .dinb(n27373), .dout(n27841));
  jxor g09819(.dina(n27654), .dinb(n27753), .dout(n27842));
  jand g09820(.dina(n27842), .dinb(n27777), .dout(n27843));
  jor  g09821(.dina(n27843), .dinb(n27841), .dout(n27844));
  jand g09822(.dina(n27844), .dinb(n426), .dout(n27845));
  jnot g09823(.din(n27845), .dout(n27846));
  jand g09824(.dina(n27786), .dinb(n27379), .dout(n27847));
  jxor g09825(.dina(n27650), .dinb(n27751), .dout(n27848));
  jand g09826(.dina(n27848), .dinb(n27777), .dout(n27849));
  jor  g09827(.dina(n27849), .dinb(n27847), .dout(n27850));
  jand g09828(.dina(n27850), .dinb(n410), .dout(n27851));
  jnot g09829(.din(n27851), .dout(n27852));
  jand g09830(.dina(n27786), .dinb(n27385), .dout(n27853));
  jxor g09831(.dina(n27646), .dinb(n27749), .dout(n27854));
  jand g09832(.dina(n27854), .dinb(n27777), .dout(n27855));
  jor  g09833(.dina(n27855), .dinb(n27853), .dout(n27856));
  jand g09834(.dina(n27856), .dinb(n409), .dout(n27857));
  jnot g09835(.din(n27857), .dout(n27858));
  jand g09836(.dina(n27786), .dinb(n27391), .dout(n27859));
  jxor g09837(.dina(n27642), .dinb(n27747), .dout(n27860));
  jand g09838(.dina(n27860), .dinb(n27777), .dout(n27861));
  jor  g09839(.dina(n27861), .dinb(n27859), .dout(n27862));
  jand g09840(.dina(n27862), .dinb(n413), .dout(n27863));
  jnot g09841(.din(n27863), .dout(n27864));
  jand g09842(.dina(n27786), .dinb(n27397), .dout(n27865));
  jxor g09843(.dina(n27638), .dinb(n27745), .dout(n27866));
  jand g09844(.dina(n27866), .dinb(n27777), .dout(n27867));
  jor  g09845(.dina(n27867), .dinb(n27865), .dout(n27868));
  jand g09846(.dina(n27868), .dinb(n412), .dout(n27869));
  jnot g09847(.din(n27869), .dout(n27870));
  jand g09848(.dina(n27786), .dinb(n27403), .dout(n27871));
  jxor g09849(.dina(n27634), .dinb(n27743), .dout(n27872));
  jand g09850(.dina(n27872), .dinb(n27777), .dout(n27873));
  jor  g09851(.dina(n27873), .dinb(n27871), .dout(n27874));
  jand g09852(.dina(n27874), .dinb(n406), .dout(n27875));
  jnot g09853(.din(n27875), .dout(n27876));
  jand g09854(.dina(n27786), .dinb(n27409), .dout(n27877));
  jxor g09855(.dina(n27630), .dinb(n27741), .dout(n27878));
  jand g09856(.dina(n27878), .dinb(n27777), .dout(n27879));
  jor  g09857(.dina(n27879), .dinb(n27877), .dout(n27880));
  jand g09858(.dina(n27880), .dinb(n405), .dout(n27881));
  jnot g09859(.din(n27881), .dout(n27882));
  jand g09860(.dina(n27786), .dinb(n27415), .dout(n27883));
  jxor g09861(.dina(n27626), .dinb(n27739), .dout(n27884));
  jand g09862(.dina(n27884), .dinb(n27777), .dout(n27885));
  jor  g09863(.dina(n27885), .dinb(n27883), .dout(n27886));
  jand g09864(.dina(n27886), .dinb(n2714), .dout(n27887));
  jnot g09865(.din(n27887), .dout(n27888));
  jand g09866(.dina(n27786), .dinb(n27421), .dout(n27889));
  jxor g09867(.dina(n27622), .dinb(n27737), .dout(n27890));
  jand g09868(.dina(n27890), .dinb(n27777), .dout(n27891));
  jor  g09869(.dina(n27891), .dinb(n27889), .dout(n27892));
  jand g09870(.dina(n27892), .dinb(n2547), .dout(n27893));
  jnot g09871(.din(n27893), .dout(n27894));
  jand g09872(.dina(n27786), .dinb(n27427), .dout(n27895));
  jxor g09873(.dina(n27618), .dinb(n27735), .dout(n27896));
  jand g09874(.dina(n27896), .dinb(n27777), .dout(n27897));
  jor  g09875(.dina(n27897), .dinb(n27895), .dout(n27898));
  jand g09876(.dina(n27898), .dinb(n417), .dout(n27899));
  jnot g09877(.din(n27899), .dout(n27900));
  jand g09878(.dina(n27786), .dinb(n27433), .dout(n27901));
  jxor g09879(.dina(n27614), .dinb(n27733), .dout(n27902));
  jand g09880(.dina(n27902), .dinb(n27777), .dout(n27903));
  jor  g09881(.dina(n27903), .dinb(n27901), .dout(n27904));
  jand g09882(.dina(n27904), .dinb(n416), .dout(n27905));
  jnot g09883(.din(n27905), .dout(n27906));
  jand g09884(.dina(n27786), .dinb(n27439), .dout(n27907));
  jxor g09885(.dina(n27610), .dinb(n27731), .dout(n27908));
  jand g09886(.dina(n27908), .dinb(n27777), .dout(n27909));
  jor  g09887(.dina(n27909), .dinb(n27907), .dout(n27910));
  jand g09888(.dina(n27910), .dinb(n422), .dout(n27911));
  jnot g09889(.din(n27911), .dout(n27912));
  jand g09890(.dina(n27786), .dinb(n27445), .dout(n27913));
  jxor g09891(.dina(n27606), .dinb(n27729), .dout(n27914));
  jand g09892(.dina(n27914), .dinb(n27777), .dout(n27915));
  jor  g09893(.dina(n27915), .dinb(n27913), .dout(n27916));
  jand g09894(.dina(n27916), .dinb(n421), .dout(n27917));
  jnot g09895(.din(n27917), .dout(n27918));
  jand g09896(.dina(n27786), .dinb(n27451), .dout(n27919));
  jxor g09897(.dina(n27602), .dinb(n27727), .dout(n27920));
  jand g09898(.dina(n27920), .dinb(n27777), .dout(n27921));
  jor  g09899(.dina(n27921), .dinb(n27919), .dout(n27922));
  jand g09900(.dina(n27922), .dinb(n433), .dout(n27923));
  jnot g09901(.din(n27923), .dout(n27924));
  jand g09902(.dina(n27786), .dinb(n27457), .dout(n27925));
  jxor g09903(.dina(n27598), .dinb(n27725), .dout(n27926));
  jand g09904(.dina(n27926), .dinb(n27777), .dout(n27927));
  jor  g09905(.dina(n27927), .dinb(n27925), .dout(n27928));
  jand g09906(.dina(n27928), .dinb(n432), .dout(n27929));
  jnot g09907(.din(n27929), .dout(n27930));
  jand g09908(.dina(n27786), .dinb(n27463), .dout(n27931));
  jxor g09909(.dina(n27594), .dinb(n27723), .dout(n27932));
  jand g09910(.dina(n27932), .dinb(n27777), .dout(n27933));
  jor  g09911(.dina(n27933), .dinb(n27931), .dout(n27934));
  jand g09912(.dina(n27934), .dinb(n436), .dout(n27935));
  jnot g09913(.din(n27935), .dout(n27936));
  jand g09914(.dina(n27786), .dinb(n27469), .dout(n27937));
  jxor g09915(.dina(n27590), .dinb(n27721), .dout(n27938));
  jand g09916(.dina(n27938), .dinb(n27777), .dout(n27939));
  jor  g09917(.dina(n27939), .dinb(n27937), .dout(n27940));
  jand g09918(.dina(n27940), .dinb(n435), .dout(n27941));
  jnot g09919(.din(n27941), .dout(n27942));
  jand g09920(.dina(n27786), .dinb(n27475), .dout(n27943));
  jxor g09921(.dina(n27586), .dinb(n27719), .dout(n27944));
  jand g09922(.dina(n27944), .dinb(n27777), .dout(n27945));
  jor  g09923(.dina(n27945), .dinb(n27943), .dout(n27946));
  jand g09924(.dina(n27946), .dinb(n440), .dout(n27947));
  jnot g09925(.din(n27947), .dout(n27948));
  jand g09926(.dina(n27786), .dinb(n27481), .dout(n27949));
  jxor g09927(.dina(n27582), .dinb(n27717), .dout(n27950));
  jand g09928(.dina(n27950), .dinb(n27777), .dout(n27951));
  jor  g09929(.dina(n27951), .dinb(n27949), .dout(n27952));
  jand g09930(.dina(n27952), .dinb(n439), .dout(n27953));
  jnot g09931(.din(n27953), .dout(n27954));
  jand g09932(.dina(n27786), .dinb(n27487), .dout(n27955));
  jxor g09933(.dina(n27578), .dinb(n27715), .dout(n27956));
  jand g09934(.dina(n27956), .dinb(n27777), .dout(n27957));
  jor  g09935(.dina(n27957), .dinb(n27955), .dout(n27958));
  jand g09936(.dina(n27958), .dinb(n325), .dout(n27959));
  jnot g09937(.din(n27959), .dout(n27960));
  jand g09938(.dina(n27786), .dinb(n27493), .dout(n27961));
  jxor g09939(.dina(n27574), .dinb(n27713), .dout(n27962));
  jand g09940(.dina(n27962), .dinb(n27777), .dout(n27963));
  jor  g09941(.dina(n27963), .dinb(n27961), .dout(n27964));
  jand g09942(.dina(n27964), .dinb(n324), .dout(n27965));
  jnot g09943(.din(n27965), .dout(n27966));
  jand g09944(.dina(n27786), .dinb(n27499), .dout(n27967));
  jxor g09945(.dina(n27570), .dinb(n27711), .dout(n27968));
  jand g09946(.dina(n27968), .dinb(n27777), .dout(n27969));
  jor  g09947(.dina(n27969), .dinb(n27967), .dout(n27970));
  jand g09948(.dina(n27970), .dinb(n323), .dout(n27971));
  jnot g09949(.din(n27971), .dout(n27972));
  jand g09950(.dina(n27786), .dinb(n27505), .dout(n27973));
  jxor g09951(.dina(n27566), .dinb(n27709), .dout(n27974));
  jand g09952(.dina(n27974), .dinb(n27777), .dout(n27975));
  jor  g09953(.dina(n27975), .dinb(n27973), .dout(n27976));
  jand g09954(.dina(n27976), .dinb(n335), .dout(n27977));
  jnot g09955(.din(n27977), .dout(n27978));
  jand g09956(.dina(n27786), .dinb(n27511), .dout(n27979));
  jxor g09957(.dina(n27562), .dinb(n27707), .dout(n27980));
  jand g09958(.dina(n27980), .dinb(n27777), .dout(n27981));
  jor  g09959(.dina(n27981), .dinb(n27979), .dout(n27982));
  jand g09960(.dina(n27982), .dinb(n334), .dout(n27983));
  jnot g09961(.din(n27983), .dout(n27984));
  jand g09962(.dina(n27786), .dinb(n27519), .dout(n27985));
  jxor g09963(.dina(n27558), .dinb(n27705), .dout(n27986));
  jand g09964(.dina(n27986), .dinb(n27777), .dout(n27987));
  jor  g09965(.dina(n27987), .dinb(n27985), .dout(n27988));
  jand g09966(.dina(n27988), .dinb(n338), .dout(n27989));
  jnot g09967(.din(n27989), .dout(n27990));
  jand g09968(.dina(n27786), .dinb(n27527), .dout(n27991));
  jxor g09969(.dina(n27554), .dinb(n27703), .dout(n27992));
  jand g09970(.dina(n27992), .dinb(n27777), .dout(n27993));
  jor  g09971(.dina(n27993), .dinb(n27991), .dout(n27994));
  jand g09972(.dina(n27994), .dinb(n337), .dout(n27995));
  jnot g09973(.din(n27995), .dout(n27996));
  jand g09974(.dina(n27786), .dinb(n27533), .dout(n27997));
  jxor g09975(.dina(n27550), .dinb(n27701), .dout(n27998));
  jand g09976(.dina(n27998), .dinb(n27777), .dout(n27999));
  jor  g09977(.dina(n27999), .dinb(n27997), .dout(n28000));
  jand g09978(.dina(n28000), .dinb(n344), .dout(n28001));
  jnot g09979(.din(n28001), .dout(n28002));
  jand g09980(.dina(n27786), .dinb(n27540), .dout(n28003));
  jxor g09981(.dina(n27699), .dinb(n7365), .dout(n28004));
  jand g09982(.dina(n28004), .dinb(n27777), .dout(n28005));
  jor  g09983(.dina(n28005), .dinb(n28003), .dout(n28006));
  jand g09984(.dina(n28006), .dinb(n348), .dout(n28007));
  jnot g09985(.din(n28007), .dout(n28008));
  jand g09986(.dina(n27777), .dinb(b0 ), .dout(n28009));
  jor  g09987(.dina(n28009), .dinb(n7363), .dout(n28010));
  jor  g09988(.dina(n27786), .dinb(n7365), .dout(n28011));
  jand g09989(.dina(n28011), .dinb(n28010), .dout(n28012));
  jor  g09990(.dina(n28012), .dinb(b1 ), .dout(n28013));
  jxor g09991(.dina(n28012), .dinb(n258), .dout(n28014));
  jor  g09992(.dina(n28014), .dinb(n7723), .dout(n28015));
  jand g09993(.dina(n28015), .dinb(n28013), .dout(n28016));
  jxor g09994(.dina(n28006), .dinb(n348), .dout(n28017));
  jnot g09995(.din(n28017), .dout(n28018));
  jor  g09996(.dina(n28018), .dinb(n28016), .dout(n28019));
  jand g09997(.dina(n28019), .dinb(n28008), .dout(n28020));
  jxor g09998(.dina(n28000), .dinb(n344), .dout(n28021));
  jnot g09999(.din(n28021), .dout(n28022));
  jor  g10000(.dina(n28022), .dinb(n28020), .dout(n28023));
  jand g10001(.dina(n28023), .dinb(n28002), .dout(n28024));
  jxor g10002(.dina(n27994), .dinb(n337), .dout(n28025));
  jnot g10003(.din(n28025), .dout(n28026));
  jor  g10004(.dina(n28026), .dinb(n28024), .dout(n28027));
  jand g10005(.dina(n28027), .dinb(n27996), .dout(n28028));
  jxor g10006(.dina(n27988), .dinb(n338), .dout(n28029));
  jnot g10007(.din(n28029), .dout(n28030));
  jor  g10008(.dina(n28030), .dinb(n28028), .dout(n28031));
  jand g10009(.dina(n28031), .dinb(n27990), .dout(n28032));
  jxor g10010(.dina(n27982), .dinb(n334), .dout(n28033));
  jnot g10011(.din(n28033), .dout(n28034));
  jor  g10012(.dina(n28034), .dinb(n28032), .dout(n28035));
  jand g10013(.dina(n28035), .dinb(n27984), .dout(n28036));
  jxor g10014(.dina(n27976), .dinb(n335), .dout(n28037));
  jnot g10015(.din(n28037), .dout(n28038));
  jor  g10016(.dina(n28038), .dinb(n28036), .dout(n28039));
  jand g10017(.dina(n28039), .dinb(n27978), .dout(n28040));
  jxor g10018(.dina(n27970), .dinb(n323), .dout(n28041));
  jnot g10019(.din(n28041), .dout(n28042));
  jor  g10020(.dina(n28042), .dinb(n28040), .dout(n28043));
  jand g10021(.dina(n28043), .dinb(n27972), .dout(n28044));
  jxor g10022(.dina(n27964), .dinb(n324), .dout(n28045));
  jnot g10023(.din(n28045), .dout(n28046));
  jor  g10024(.dina(n28046), .dinb(n28044), .dout(n28047));
  jand g10025(.dina(n28047), .dinb(n27966), .dout(n28048));
  jxor g10026(.dina(n27958), .dinb(n325), .dout(n28049));
  jnot g10027(.din(n28049), .dout(n28050));
  jor  g10028(.dina(n28050), .dinb(n28048), .dout(n28051));
  jand g10029(.dina(n28051), .dinb(n27960), .dout(n28052));
  jxor g10030(.dina(n27952), .dinb(n439), .dout(n28053));
  jnot g10031(.din(n28053), .dout(n28054));
  jor  g10032(.dina(n28054), .dinb(n28052), .dout(n28055));
  jand g10033(.dina(n28055), .dinb(n27954), .dout(n28056));
  jxor g10034(.dina(n27946), .dinb(n440), .dout(n28057));
  jnot g10035(.din(n28057), .dout(n28058));
  jor  g10036(.dina(n28058), .dinb(n28056), .dout(n28059));
  jand g10037(.dina(n28059), .dinb(n27948), .dout(n28060));
  jxor g10038(.dina(n27940), .dinb(n435), .dout(n28061));
  jnot g10039(.din(n28061), .dout(n28062));
  jor  g10040(.dina(n28062), .dinb(n28060), .dout(n28063));
  jand g10041(.dina(n28063), .dinb(n27942), .dout(n28064));
  jxor g10042(.dina(n27934), .dinb(n436), .dout(n28065));
  jnot g10043(.din(n28065), .dout(n28066));
  jor  g10044(.dina(n28066), .dinb(n28064), .dout(n28067));
  jand g10045(.dina(n28067), .dinb(n27936), .dout(n28068));
  jxor g10046(.dina(n27928), .dinb(n432), .dout(n28069));
  jnot g10047(.din(n28069), .dout(n28070));
  jor  g10048(.dina(n28070), .dinb(n28068), .dout(n28071));
  jand g10049(.dina(n28071), .dinb(n27930), .dout(n28072));
  jxor g10050(.dina(n27922), .dinb(n433), .dout(n28073));
  jnot g10051(.din(n28073), .dout(n28074));
  jor  g10052(.dina(n28074), .dinb(n28072), .dout(n28075));
  jand g10053(.dina(n28075), .dinb(n27924), .dout(n28076));
  jxor g10054(.dina(n27916), .dinb(n421), .dout(n28077));
  jnot g10055(.din(n28077), .dout(n28078));
  jor  g10056(.dina(n28078), .dinb(n28076), .dout(n28079));
  jand g10057(.dina(n28079), .dinb(n27918), .dout(n28080));
  jxor g10058(.dina(n27910), .dinb(n422), .dout(n28081));
  jnot g10059(.din(n28081), .dout(n28082));
  jor  g10060(.dina(n28082), .dinb(n28080), .dout(n28083));
  jand g10061(.dina(n28083), .dinb(n27912), .dout(n28084));
  jxor g10062(.dina(n27904), .dinb(n416), .dout(n28085));
  jnot g10063(.din(n28085), .dout(n28086));
  jor  g10064(.dina(n28086), .dinb(n28084), .dout(n28087));
  jand g10065(.dina(n28087), .dinb(n27906), .dout(n28088));
  jxor g10066(.dina(n27898), .dinb(n417), .dout(n28089));
  jnot g10067(.din(n28089), .dout(n28090));
  jor  g10068(.dina(n28090), .dinb(n28088), .dout(n28091));
  jand g10069(.dina(n28091), .dinb(n27900), .dout(n28092));
  jxor g10070(.dina(n27892), .dinb(n2547), .dout(n28093));
  jnot g10071(.din(n28093), .dout(n28094));
  jor  g10072(.dina(n28094), .dinb(n28092), .dout(n28095));
  jand g10073(.dina(n28095), .dinb(n27894), .dout(n28096));
  jxor g10074(.dina(n27886), .dinb(n2714), .dout(n28097));
  jnot g10075(.din(n28097), .dout(n28098));
  jor  g10076(.dina(n28098), .dinb(n28096), .dout(n28099));
  jand g10077(.dina(n28099), .dinb(n27888), .dout(n28100));
  jxor g10078(.dina(n27880), .dinb(n405), .dout(n28101));
  jnot g10079(.din(n28101), .dout(n28102));
  jor  g10080(.dina(n28102), .dinb(n28100), .dout(n28103));
  jand g10081(.dina(n28103), .dinb(n27882), .dout(n28104));
  jxor g10082(.dina(n27874), .dinb(n406), .dout(n28105));
  jnot g10083(.din(n28105), .dout(n28106));
  jor  g10084(.dina(n28106), .dinb(n28104), .dout(n28107));
  jand g10085(.dina(n28107), .dinb(n27876), .dout(n28108));
  jxor g10086(.dina(n27868), .dinb(n412), .dout(n28109));
  jnot g10087(.din(n28109), .dout(n28110));
  jor  g10088(.dina(n28110), .dinb(n28108), .dout(n28111));
  jand g10089(.dina(n28111), .dinb(n27870), .dout(n28112));
  jxor g10090(.dina(n27862), .dinb(n413), .dout(n28113));
  jnot g10091(.din(n28113), .dout(n28114));
  jor  g10092(.dina(n28114), .dinb(n28112), .dout(n28115));
  jand g10093(.dina(n28115), .dinb(n27864), .dout(n28116));
  jxor g10094(.dina(n27856), .dinb(n409), .dout(n28117));
  jnot g10095(.din(n28117), .dout(n28118));
  jor  g10096(.dina(n28118), .dinb(n28116), .dout(n28119));
  jand g10097(.dina(n28119), .dinb(n27858), .dout(n28120));
  jxor g10098(.dina(n27850), .dinb(n410), .dout(n28121));
  jnot g10099(.din(n28121), .dout(n28122));
  jor  g10100(.dina(n28122), .dinb(n28120), .dout(n28123));
  jand g10101(.dina(n28123), .dinb(n27852), .dout(n28124));
  jxor g10102(.dina(n27844), .dinb(n426), .dout(n28125));
  jnot g10103(.din(n28125), .dout(n28126));
  jor  g10104(.dina(n28126), .dinb(n28124), .dout(n28127));
  jand g10105(.dina(n28127), .dinb(n27846), .dout(n28128));
  jxor g10106(.dina(n27838), .dinb(n427), .dout(n28129));
  jnot g10107(.din(n28129), .dout(n28130));
  jor  g10108(.dina(n28130), .dinb(n28128), .dout(n28131));
  jand g10109(.dina(n28131), .dinb(n27840), .dout(n28132));
  jxor g10110(.dina(n27832), .dinb(n424), .dout(n28133));
  jnot g10111(.din(n28133), .dout(n28134));
  jor  g10112(.dina(n28134), .dinb(n28132), .dout(n28135));
  jand g10113(.dina(n28135), .dinb(n27834), .dout(n28136));
  jxor g10114(.dina(n27826), .dinb(n300), .dout(n28137));
  jnot g10115(.din(n28137), .dout(n28138));
  jor  g10116(.dina(n28138), .dinb(n28136), .dout(n28139));
  jand g10117(.dina(n28139), .dinb(n27828), .dout(n28140));
  jxor g10118(.dina(n27820), .dinb(n297), .dout(n28141));
  jnot g10119(.din(n28141), .dout(n28142));
  jor  g10120(.dina(n28142), .dinb(n28140), .dout(n28143));
  jand g10121(.dina(n28143), .dinb(n27822), .dout(n28144));
  jxor g10122(.dina(n27814), .dinb(n298), .dout(n28145));
  jnot g10123(.din(n28145), .dout(n28146));
  jor  g10124(.dina(n28146), .dinb(n28144), .dout(n28147));
  jand g10125(.dina(n28147), .dinb(n27816), .dout(n28148));
  jxor g10126(.dina(n27808), .dinb(n301), .dout(n28149));
  jnot g10127(.din(n28149), .dout(n28150));
  jor  g10128(.dina(n28150), .dinb(n28148), .dout(n28151));
  jand g10129(.dina(n28151), .dinb(n27810), .dout(n28152));
  jxor g10130(.dina(n27802), .dinb(n293), .dout(n28153));
  jnot g10131(.din(n28153), .dout(n28154));
  jor  g10132(.dina(n28154), .dinb(n28152), .dout(n28155));
  jand g10133(.dina(n28155), .dinb(n27804), .dout(n28156));
  jxor g10134(.dina(n27796), .dinb(n294), .dout(n28157));
  jnot g10135(.din(n28157), .dout(n28158));
  jor  g10136(.dina(n28158), .dinb(n28156), .dout(n28159));
  jand g10137(.dina(n28159), .dinb(n27798), .dout(n28160));
  jxor g10138(.dina(n27790), .dinb(n290), .dout(n28161));
  jnot g10139(.din(n28161), .dout(n28162));
  jor  g10140(.dina(n28162), .dinb(n28160), .dout(n28163));
  jand g10141(.dina(n28163), .dinb(n27792), .dout(n28164));
  jand g10142(.dina(n28164), .dinb(n27784), .dout(n28165));
  jor  g10143(.dina(n28165), .dinb(n27782), .dout(n28166));
  jor  g10144(.dina(n28166), .dinb(n289), .dout(n28167));
  jand g10145(.dina(n28167), .dinb(n27781), .dout(n28168));
  jor  g10146(.dina(n27786), .dinb(n18364), .dout(n28169));
  jand g10147(.dina(n28169), .dinb(a25 ), .dout(n28170));
  jnot g10148(.din(n28011), .dout(n28171));
  jor  g10149(.dina(n28171), .dinb(n28170), .dout(n28172));
  jand g10150(.dina(n28172), .dinb(n258), .dout(n28173));
  jxor g10151(.dina(n28012), .dinb(b1 ), .dout(n28174));
  jand g10152(.dina(n28174), .dinb(n7883), .dout(n28175));
  jor  g10153(.dina(n28175), .dinb(n28173), .dout(n28176));
  jand g10154(.dina(n28017), .dinb(n28176), .dout(n28177));
  jor  g10155(.dina(n28177), .dinb(n28007), .dout(n28178));
  jand g10156(.dina(n28021), .dinb(n28178), .dout(n28179));
  jor  g10157(.dina(n28179), .dinb(n28001), .dout(n28180));
  jand g10158(.dina(n28025), .dinb(n28180), .dout(n28181));
  jor  g10159(.dina(n28181), .dinb(n27995), .dout(n28182));
  jand g10160(.dina(n28029), .dinb(n28182), .dout(n28183));
  jor  g10161(.dina(n28183), .dinb(n27989), .dout(n28184));
  jand g10162(.dina(n28033), .dinb(n28184), .dout(n28185));
  jor  g10163(.dina(n28185), .dinb(n27983), .dout(n28186));
  jand g10164(.dina(n28037), .dinb(n28186), .dout(n28187));
  jor  g10165(.dina(n28187), .dinb(n27977), .dout(n28188));
  jand g10166(.dina(n28041), .dinb(n28188), .dout(n28189));
  jor  g10167(.dina(n28189), .dinb(n27971), .dout(n28190));
  jand g10168(.dina(n28045), .dinb(n28190), .dout(n28191));
  jor  g10169(.dina(n28191), .dinb(n27965), .dout(n28192));
  jand g10170(.dina(n28049), .dinb(n28192), .dout(n28193));
  jor  g10171(.dina(n28193), .dinb(n27959), .dout(n28194));
  jand g10172(.dina(n28053), .dinb(n28194), .dout(n28195));
  jor  g10173(.dina(n28195), .dinb(n27953), .dout(n28196));
  jand g10174(.dina(n28057), .dinb(n28196), .dout(n28197));
  jor  g10175(.dina(n28197), .dinb(n27947), .dout(n28198));
  jand g10176(.dina(n28061), .dinb(n28198), .dout(n28199));
  jor  g10177(.dina(n28199), .dinb(n27941), .dout(n28200));
  jand g10178(.dina(n28065), .dinb(n28200), .dout(n28201));
  jor  g10179(.dina(n28201), .dinb(n27935), .dout(n28202));
  jand g10180(.dina(n28069), .dinb(n28202), .dout(n28203));
  jor  g10181(.dina(n28203), .dinb(n27929), .dout(n28204));
  jand g10182(.dina(n28073), .dinb(n28204), .dout(n28205));
  jor  g10183(.dina(n28205), .dinb(n27923), .dout(n28206));
  jand g10184(.dina(n28077), .dinb(n28206), .dout(n28207));
  jor  g10185(.dina(n28207), .dinb(n27917), .dout(n28208));
  jand g10186(.dina(n28081), .dinb(n28208), .dout(n28209));
  jor  g10187(.dina(n28209), .dinb(n27911), .dout(n28210));
  jand g10188(.dina(n28085), .dinb(n28210), .dout(n28211));
  jor  g10189(.dina(n28211), .dinb(n27905), .dout(n28212));
  jand g10190(.dina(n28089), .dinb(n28212), .dout(n28213));
  jor  g10191(.dina(n28213), .dinb(n27899), .dout(n28214));
  jand g10192(.dina(n28093), .dinb(n28214), .dout(n28215));
  jor  g10193(.dina(n28215), .dinb(n27893), .dout(n28216));
  jand g10194(.dina(n28097), .dinb(n28216), .dout(n28217));
  jor  g10195(.dina(n28217), .dinb(n27887), .dout(n28218));
  jand g10196(.dina(n28101), .dinb(n28218), .dout(n28219));
  jor  g10197(.dina(n28219), .dinb(n27881), .dout(n28220));
  jand g10198(.dina(n28105), .dinb(n28220), .dout(n28221));
  jor  g10199(.dina(n28221), .dinb(n27875), .dout(n28222));
  jand g10200(.dina(n28109), .dinb(n28222), .dout(n28223));
  jor  g10201(.dina(n28223), .dinb(n27869), .dout(n28224));
  jand g10202(.dina(n28113), .dinb(n28224), .dout(n28225));
  jor  g10203(.dina(n28225), .dinb(n27863), .dout(n28226));
  jand g10204(.dina(n28117), .dinb(n28226), .dout(n28227));
  jor  g10205(.dina(n28227), .dinb(n27857), .dout(n28228));
  jand g10206(.dina(n28121), .dinb(n28228), .dout(n28229));
  jor  g10207(.dina(n28229), .dinb(n27851), .dout(n28230));
  jand g10208(.dina(n28125), .dinb(n28230), .dout(n28231));
  jor  g10209(.dina(n28231), .dinb(n27845), .dout(n28232));
  jand g10210(.dina(n28129), .dinb(n28232), .dout(n28233));
  jor  g10211(.dina(n28233), .dinb(n27839), .dout(n28234));
  jand g10212(.dina(n28133), .dinb(n28234), .dout(n28235));
  jor  g10213(.dina(n28235), .dinb(n27833), .dout(n28236));
  jand g10214(.dina(n28137), .dinb(n28236), .dout(n28237));
  jor  g10215(.dina(n28237), .dinb(n27827), .dout(n28238));
  jand g10216(.dina(n28141), .dinb(n28238), .dout(n28239));
  jor  g10217(.dina(n28239), .dinb(n27821), .dout(n28240));
  jand g10218(.dina(n28145), .dinb(n28240), .dout(n28241));
  jor  g10219(.dina(n28241), .dinb(n27815), .dout(n28242));
  jand g10220(.dina(n28149), .dinb(n28242), .dout(n28243));
  jor  g10221(.dina(n28243), .dinb(n27809), .dout(n28244));
  jand g10222(.dina(n28153), .dinb(n28244), .dout(n28245));
  jor  g10223(.dina(n28245), .dinb(n27803), .dout(n28246));
  jand g10224(.dina(n28157), .dinb(n28246), .dout(n28247));
  jor  g10225(.dina(n28247), .dinb(n27797), .dout(n28248));
  jand g10226(.dina(n28161), .dinb(n28248), .dout(n28249));
  jor  g10227(.dina(n28249), .dinb(n27791), .dout(n28250));
  jand g10228(.dina(n27783), .dinb(n589), .dout(n28251));
  jand g10229(.dina(n28251), .dinb(n28250), .dout(n28252));
  jor  g10230(.dina(n28252), .dinb(n28168), .dout(n28253));
  jand g10231(.dina(n28253), .dinb(n284), .dout(n28254));
  jnot g10232(.din(n28254), .dout(n28255));
  jand g10233(.dina(n28167), .dinb(n27790), .dout(n28256));
  jnot g10234(.din(n27782), .dout(n28257));
  jor  g10235(.dina(n28250), .dinb(n27783), .dout(n28258));
  jand g10236(.dina(n28258), .dinb(n28257), .dout(n28259));
  jand g10237(.dina(n28259), .dinb(n589), .dout(n28260));
  jxor g10238(.dina(n28161), .dinb(n28248), .dout(n28261));
  jand g10239(.dina(n28261), .dinb(n28260), .dout(n28262));
  jor  g10240(.dina(n28262), .dinb(n28256), .dout(n28263));
  jand g10241(.dina(n28263), .dinb(n291), .dout(n28264));
  jnot g10242(.din(n28264), .dout(n28265));
  jand g10243(.dina(n28167), .dinb(n27796), .dout(n28266));
  jxor g10244(.dina(n28157), .dinb(n28246), .dout(n28267));
  jand g10245(.dina(n28267), .dinb(n28260), .dout(n28268));
  jor  g10246(.dina(n28268), .dinb(n28266), .dout(n28269));
  jand g10247(.dina(n28269), .dinb(n290), .dout(n28270));
  jnot g10248(.din(n28270), .dout(n28271));
  jand g10249(.dina(n28167), .dinb(n27802), .dout(n28272));
  jxor g10250(.dina(n28153), .dinb(n28244), .dout(n28273));
  jand g10251(.dina(n28273), .dinb(n28260), .dout(n28274));
  jor  g10252(.dina(n28274), .dinb(n28272), .dout(n28275));
  jand g10253(.dina(n28275), .dinb(n294), .dout(n28276));
  jnot g10254(.din(n28276), .dout(n28277));
  jand g10255(.dina(n28167), .dinb(n27808), .dout(n28278));
  jxor g10256(.dina(n28149), .dinb(n28242), .dout(n28279));
  jand g10257(.dina(n28279), .dinb(n28260), .dout(n28280));
  jor  g10258(.dina(n28280), .dinb(n28278), .dout(n28281));
  jand g10259(.dina(n28281), .dinb(n293), .dout(n28282));
  jnot g10260(.din(n28282), .dout(n28283));
  jand g10261(.dina(n28167), .dinb(n27814), .dout(n28284));
  jxor g10262(.dina(n28145), .dinb(n28240), .dout(n28285));
  jand g10263(.dina(n28285), .dinb(n28260), .dout(n28286));
  jor  g10264(.dina(n28286), .dinb(n28284), .dout(n28287));
  jand g10265(.dina(n28287), .dinb(n301), .dout(n28288));
  jnot g10266(.din(n28288), .dout(n28289));
  jand g10267(.dina(n28167), .dinb(n27820), .dout(n28290));
  jxor g10268(.dina(n28141), .dinb(n28238), .dout(n28291));
  jand g10269(.dina(n28291), .dinb(n28260), .dout(n28292));
  jor  g10270(.dina(n28292), .dinb(n28290), .dout(n28293));
  jand g10271(.dina(n28293), .dinb(n298), .dout(n28294));
  jnot g10272(.din(n28294), .dout(n28295));
  jand g10273(.dina(n28167), .dinb(n27826), .dout(n28296));
  jxor g10274(.dina(n28137), .dinb(n28236), .dout(n28297));
  jand g10275(.dina(n28297), .dinb(n28260), .dout(n28298));
  jor  g10276(.dina(n28298), .dinb(n28296), .dout(n28299));
  jand g10277(.dina(n28299), .dinb(n297), .dout(n28300));
  jnot g10278(.din(n28300), .dout(n28301));
  jand g10279(.dina(n28167), .dinb(n27832), .dout(n28302));
  jxor g10280(.dina(n28133), .dinb(n28234), .dout(n28303));
  jand g10281(.dina(n28303), .dinb(n28260), .dout(n28304));
  jor  g10282(.dina(n28304), .dinb(n28302), .dout(n28305));
  jand g10283(.dina(n28305), .dinb(n300), .dout(n28306));
  jnot g10284(.din(n28306), .dout(n28307));
  jand g10285(.dina(n28167), .dinb(n27838), .dout(n28308));
  jxor g10286(.dina(n28129), .dinb(n28232), .dout(n28309));
  jand g10287(.dina(n28309), .dinb(n28260), .dout(n28310));
  jor  g10288(.dina(n28310), .dinb(n28308), .dout(n28311));
  jand g10289(.dina(n28311), .dinb(n424), .dout(n28312));
  jnot g10290(.din(n28312), .dout(n28313));
  jand g10291(.dina(n28167), .dinb(n27844), .dout(n28314));
  jxor g10292(.dina(n28125), .dinb(n28230), .dout(n28315));
  jand g10293(.dina(n28315), .dinb(n28260), .dout(n28316));
  jor  g10294(.dina(n28316), .dinb(n28314), .dout(n28317));
  jand g10295(.dina(n28317), .dinb(n427), .dout(n28318));
  jnot g10296(.din(n28318), .dout(n28319));
  jand g10297(.dina(n28167), .dinb(n27850), .dout(n28320));
  jxor g10298(.dina(n28121), .dinb(n28228), .dout(n28321));
  jand g10299(.dina(n28321), .dinb(n28260), .dout(n28322));
  jor  g10300(.dina(n28322), .dinb(n28320), .dout(n28323));
  jand g10301(.dina(n28323), .dinb(n426), .dout(n28324));
  jnot g10302(.din(n28324), .dout(n28325));
  jand g10303(.dina(n28167), .dinb(n27856), .dout(n28326));
  jxor g10304(.dina(n28117), .dinb(n28226), .dout(n28327));
  jand g10305(.dina(n28327), .dinb(n28260), .dout(n28328));
  jor  g10306(.dina(n28328), .dinb(n28326), .dout(n28329));
  jand g10307(.dina(n28329), .dinb(n410), .dout(n28330));
  jnot g10308(.din(n28330), .dout(n28331));
  jand g10309(.dina(n28167), .dinb(n27862), .dout(n28332));
  jxor g10310(.dina(n28113), .dinb(n28224), .dout(n28333));
  jand g10311(.dina(n28333), .dinb(n28260), .dout(n28334));
  jor  g10312(.dina(n28334), .dinb(n28332), .dout(n28335));
  jand g10313(.dina(n28335), .dinb(n409), .dout(n28336));
  jnot g10314(.din(n28336), .dout(n28337));
  jand g10315(.dina(n28167), .dinb(n27868), .dout(n28338));
  jxor g10316(.dina(n28109), .dinb(n28222), .dout(n28339));
  jand g10317(.dina(n28339), .dinb(n28260), .dout(n28340));
  jor  g10318(.dina(n28340), .dinb(n28338), .dout(n28341));
  jand g10319(.dina(n28341), .dinb(n413), .dout(n28342));
  jnot g10320(.din(n28342), .dout(n28343));
  jand g10321(.dina(n28167), .dinb(n27874), .dout(n28344));
  jxor g10322(.dina(n28105), .dinb(n28220), .dout(n28345));
  jand g10323(.dina(n28345), .dinb(n28260), .dout(n28346));
  jor  g10324(.dina(n28346), .dinb(n28344), .dout(n28347));
  jand g10325(.dina(n28347), .dinb(n412), .dout(n28348));
  jnot g10326(.din(n28348), .dout(n28349));
  jand g10327(.dina(n28167), .dinb(n27880), .dout(n28350));
  jxor g10328(.dina(n28101), .dinb(n28218), .dout(n28351));
  jand g10329(.dina(n28351), .dinb(n28260), .dout(n28352));
  jor  g10330(.dina(n28352), .dinb(n28350), .dout(n28353));
  jand g10331(.dina(n28353), .dinb(n406), .dout(n28354));
  jnot g10332(.din(n28354), .dout(n28355));
  jand g10333(.dina(n28167), .dinb(n27886), .dout(n28356));
  jxor g10334(.dina(n28097), .dinb(n28216), .dout(n28357));
  jand g10335(.dina(n28357), .dinb(n28260), .dout(n28358));
  jor  g10336(.dina(n28358), .dinb(n28356), .dout(n28359));
  jand g10337(.dina(n28359), .dinb(n405), .dout(n28360));
  jnot g10338(.din(n28360), .dout(n28361));
  jand g10339(.dina(n28167), .dinb(n27892), .dout(n28362));
  jxor g10340(.dina(n28093), .dinb(n28214), .dout(n28363));
  jand g10341(.dina(n28363), .dinb(n28260), .dout(n28364));
  jor  g10342(.dina(n28364), .dinb(n28362), .dout(n28365));
  jand g10343(.dina(n28365), .dinb(n2714), .dout(n28366));
  jnot g10344(.din(n28366), .dout(n28367));
  jand g10345(.dina(n28167), .dinb(n27898), .dout(n28368));
  jxor g10346(.dina(n28089), .dinb(n28212), .dout(n28369));
  jand g10347(.dina(n28369), .dinb(n28260), .dout(n28370));
  jor  g10348(.dina(n28370), .dinb(n28368), .dout(n28371));
  jand g10349(.dina(n28371), .dinb(n2547), .dout(n28372));
  jnot g10350(.din(n28372), .dout(n28373));
  jand g10351(.dina(n28167), .dinb(n27904), .dout(n28374));
  jxor g10352(.dina(n28085), .dinb(n28210), .dout(n28375));
  jand g10353(.dina(n28375), .dinb(n28260), .dout(n28376));
  jor  g10354(.dina(n28376), .dinb(n28374), .dout(n28377));
  jand g10355(.dina(n28377), .dinb(n417), .dout(n28378));
  jnot g10356(.din(n28378), .dout(n28379));
  jand g10357(.dina(n28167), .dinb(n27910), .dout(n28380));
  jxor g10358(.dina(n28081), .dinb(n28208), .dout(n28381));
  jand g10359(.dina(n28381), .dinb(n28260), .dout(n28382));
  jor  g10360(.dina(n28382), .dinb(n28380), .dout(n28383));
  jand g10361(.dina(n28383), .dinb(n416), .dout(n28384));
  jnot g10362(.din(n28384), .dout(n28385));
  jand g10363(.dina(n28167), .dinb(n27916), .dout(n28386));
  jxor g10364(.dina(n28077), .dinb(n28206), .dout(n28387));
  jand g10365(.dina(n28387), .dinb(n28260), .dout(n28388));
  jor  g10366(.dina(n28388), .dinb(n28386), .dout(n28389));
  jand g10367(.dina(n28389), .dinb(n422), .dout(n28390));
  jnot g10368(.din(n28390), .dout(n28391));
  jand g10369(.dina(n28167), .dinb(n27922), .dout(n28392));
  jxor g10370(.dina(n28073), .dinb(n28204), .dout(n28393));
  jand g10371(.dina(n28393), .dinb(n28260), .dout(n28394));
  jor  g10372(.dina(n28394), .dinb(n28392), .dout(n28395));
  jand g10373(.dina(n28395), .dinb(n421), .dout(n28396));
  jnot g10374(.din(n28396), .dout(n28397));
  jand g10375(.dina(n28167), .dinb(n27928), .dout(n28398));
  jxor g10376(.dina(n28069), .dinb(n28202), .dout(n28399));
  jand g10377(.dina(n28399), .dinb(n28260), .dout(n28400));
  jor  g10378(.dina(n28400), .dinb(n28398), .dout(n28401));
  jand g10379(.dina(n28401), .dinb(n433), .dout(n28402));
  jnot g10380(.din(n28402), .dout(n28403));
  jand g10381(.dina(n28167), .dinb(n27934), .dout(n28404));
  jxor g10382(.dina(n28065), .dinb(n28200), .dout(n28405));
  jand g10383(.dina(n28405), .dinb(n28260), .dout(n28406));
  jor  g10384(.dina(n28406), .dinb(n28404), .dout(n28407));
  jand g10385(.dina(n28407), .dinb(n432), .dout(n28408));
  jnot g10386(.din(n28408), .dout(n28409));
  jand g10387(.dina(n28167), .dinb(n27940), .dout(n28410));
  jxor g10388(.dina(n28061), .dinb(n28198), .dout(n28411));
  jand g10389(.dina(n28411), .dinb(n28260), .dout(n28412));
  jor  g10390(.dina(n28412), .dinb(n28410), .dout(n28413));
  jand g10391(.dina(n28413), .dinb(n436), .dout(n28414));
  jnot g10392(.din(n28414), .dout(n28415));
  jand g10393(.dina(n28167), .dinb(n27946), .dout(n28416));
  jxor g10394(.dina(n28057), .dinb(n28196), .dout(n28417));
  jand g10395(.dina(n28417), .dinb(n28260), .dout(n28418));
  jor  g10396(.dina(n28418), .dinb(n28416), .dout(n28419));
  jand g10397(.dina(n28419), .dinb(n435), .dout(n28420));
  jnot g10398(.din(n28420), .dout(n28421));
  jand g10399(.dina(n28167), .dinb(n27952), .dout(n28422));
  jxor g10400(.dina(n28053), .dinb(n28194), .dout(n28423));
  jand g10401(.dina(n28423), .dinb(n28260), .dout(n28424));
  jor  g10402(.dina(n28424), .dinb(n28422), .dout(n28425));
  jand g10403(.dina(n28425), .dinb(n440), .dout(n28426));
  jnot g10404(.din(n28426), .dout(n28427));
  jand g10405(.dina(n28167), .dinb(n27958), .dout(n28428));
  jxor g10406(.dina(n28049), .dinb(n28192), .dout(n28429));
  jand g10407(.dina(n28429), .dinb(n28260), .dout(n28430));
  jor  g10408(.dina(n28430), .dinb(n28428), .dout(n28431));
  jand g10409(.dina(n28431), .dinb(n439), .dout(n28432));
  jnot g10410(.din(n28432), .dout(n28433));
  jand g10411(.dina(n28167), .dinb(n27964), .dout(n28434));
  jxor g10412(.dina(n28045), .dinb(n28190), .dout(n28435));
  jand g10413(.dina(n28435), .dinb(n28260), .dout(n28436));
  jor  g10414(.dina(n28436), .dinb(n28434), .dout(n28437));
  jand g10415(.dina(n28437), .dinb(n325), .dout(n28438));
  jnot g10416(.din(n28438), .dout(n28439));
  jand g10417(.dina(n28167), .dinb(n27970), .dout(n28440));
  jxor g10418(.dina(n28041), .dinb(n28188), .dout(n28441));
  jand g10419(.dina(n28441), .dinb(n28260), .dout(n28442));
  jor  g10420(.dina(n28442), .dinb(n28440), .dout(n28443));
  jand g10421(.dina(n28443), .dinb(n324), .dout(n28444));
  jnot g10422(.din(n28444), .dout(n28445));
  jand g10423(.dina(n28167), .dinb(n27976), .dout(n28446));
  jxor g10424(.dina(n28037), .dinb(n28186), .dout(n28447));
  jand g10425(.dina(n28447), .dinb(n28260), .dout(n28448));
  jor  g10426(.dina(n28448), .dinb(n28446), .dout(n28449));
  jand g10427(.dina(n28449), .dinb(n323), .dout(n28450));
  jnot g10428(.din(n28450), .dout(n28451));
  jand g10429(.dina(n28167), .dinb(n27982), .dout(n28452));
  jxor g10430(.dina(n28033), .dinb(n28184), .dout(n28453));
  jand g10431(.dina(n28453), .dinb(n28260), .dout(n28454));
  jor  g10432(.dina(n28454), .dinb(n28452), .dout(n28455));
  jand g10433(.dina(n28455), .dinb(n335), .dout(n28456));
  jnot g10434(.din(n28456), .dout(n28457));
  jand g10435(.dina(n28167), .dinb(n27988), .dout(n28458));
  jxor g10436(.dina(n28029), .dinb(n28182), .dout(n28459));
  jand g10437(.dina(n28459), .dinb(n28260), .dout(n28460));
  jor  g10438(.dina(n28460), .dinb(n28458), .dout(n28461));
  jand g10439(.dina(n28461), .dinb(n334), .dout(n28462));
  jnot g10440(.din(n28462), .dout(n28463));
  jand g10441(.dina(n28167), .dinb(n27994), .dout(n28464));
  jxor g10442(.dina(n28025), .dinb(n28180), .dout(n28465));
  jand g10443(.dina(n28465), .dinb(n28260), .dout(n28466));
  jor  g10444(.dina(n28466), .dinb(n28464), .dout(n28467));
  jand g10445(.dina(n28467), .dinb(n338), .dout(n28468));
  jnot g10446(.din(n28468), .dout(n28469));
  jand g10447(.dina(n28167), .dinb(n28000), .dout(n28470));
  jxor g10448(.dina(n28021), .dinb(n28178), .dout(n28471));
  jand g10449(.dina(n28471), .dinb(n28260), .dout(n28472));
  jor  g10450(.dina(n28472), .dinb(n28470), .dout(n28473));
  jand g10451(.dina(n28473), .dinb(n337), .dout(n28474));
  jnot g10452(.din(n28474), .dout(n28475));
  jnot g10453(.din(n28006), .dout(n28476));
  jor  g10454(.dina(n28260), .dinb(n28476), .dout(n28477));
  jxor g10455(.dina(n28017), .dinb(n28176), .dout(n28478));
  jnot g10456(.din(n28478), .dout(n28479));
  jor  g10457(.dina(n28479), .dinb(n28167), .dout(n28480));
  jand g10458(.dina(n28480), .dinb(n28477), .dout(n28481));
  jor  g10459(.dina(n28481), .dinb(b3 ), .dout(n28482));
  jand g10460(.dina(n28167), .dinb(n28172), .dout(n28483));
  jxor g10461(.dina(n28174), .dinb(n7883), .dout(n28484));
  jand g10462(.dina(n28484), .dinb(n28260), .dout(n28485));
  jor  g10463(.dina(n28485), .dinb(n28483), .dout(n28486));
  jand g10464(.dina(n28486), .dinb(n348), .dout(n28487));
  jnot g10465(.din(n28487), .dout(n28488));
  jand g10466(.dina(n28259), .dinb(n7355), .dout(n28489));
  jor  g10467(.dina(n28489), .dinb(n7722), .dout(n28490));
  jor  g10468(.dina(n28167), .dinb(n7883), .dout(n28491));
  jand g10469(.dina(n28491), .dinb(n28490), .dout(n28492));
  jor  g10470(.dina(n28492), .dinb(b1 ), .dout(n28493));
  jxor g10471(.dina(n28492), .dinb(n258), .dout(n28494));
  jor  g10472(.dina(n28494), .dinb(n8204), .dout(n28495));
  jand g10473(.dina(n28495), .dinb(n28493), .dout(n28496));
  jxor g10474(.dina(n28486), .dinb(n348), .dout(n28497));
  jnot g10475(.din(n28497), .dout(n28498));
  jor  g10476(.dina(n28498), .dinb(n28496), .dout(n28499));
  jand g10477(.dina(n28499), .dinb(n28488), .dout(n28500));
  jxor g10478(.dina(n28481), .dinb(b3 ), .dout(n28501));
  jnot g10479(.din(n28501), .dout(n28502));
  jor  g10480(.dina(n28502), .dinb(n28500), .dout(n28503));
  jand g10481(.dina(n28503), .dinb(n28482), .dout(n28504));
  jxor g10482(.dina(n28473), .dinb(n337), .dout(n28505));
  jnot g10483(.din(n28505), .dout(n28506));
  jor  g10484(.dina(n28506), .dinb(n28504), .dout(n28507));
  jand g10485(.dina(n28507), .dinb(n28475), .dout(n28508));
  jxor g10486(.dina(n28467), .dinb(n338), .dout(n28509));
  jnot g10487(.din(n28509), .dout(n28510));
  jor  g10488(.dina(n28510), .dinb(n28508), .dout(n28511));
  jand g10489(.dina(n28511), .dinb(n28469), .dout(n28512));
  jxor g10490(.dina(n28461), .dinb(n334), .dout(n28513));
  jnot g10491(.din(n28513), .dout(n28514));
  jor  g10492(.dina(n28514), .dinb(n28512), .dout(n28515));
  jand g10493(.dina(n28515), .dinb(n28463), .dout(n28516));
  jxor g10494(.dina(n28455), .dinb(n335), .dout(n28517));
  jnot g10495(.din(n28517), .dout(n28518));
  jor  g10496(.dina(n28518), .dinb(n28516), .dout(n28519));
  jand g10497(.dina(n28519), .dinb(n28457), .dout(n28520));
  jxor g10498(.dina(n28449), .dinb(n323), .dout(n28521));
  jnot g10499(.din(n28521), .dout(n28522));
  jor  g10500(.dina(n28522), .dinb(n28520), .dout(n28523));
  jand g10501(.dina(n28523), .dinb(n28451), .dout(n28524));
  jxor g10502(.dina(n28443), .dinb(n324), .dout(n28525));
  jnot g10503(.din(n28525), .dout(n28526));
  jor  g10504(.dina(n28526), .dinb(n28524), .dout(n28527));
  jand g10505(.dina(n28527), .dinb(n28445), .dout(n28528));
  jxor g10506(.dina(n28437), .dinb(n325), .dout(n28529));
  jnot g10507(.din(n28529), .dout(n28530));
  jor  g10508(.dina(n28530), .dinb(n28528), .dout(n28531));
  jand g10509(.dina(n28531), .dinb(n28439), .dout(n28532));
  jxor g10510(.dina(n28431), .dinb(n439), .dout(n28533));
  jnot g10511(.din(n28533), .dout(n28534));
  jor  g10512(.dina(n28534), .dinb(n28532), .dout(n28535));
  jand g10513(.dina(n28535), .dinb(n28433), .dout(n28536));
  jxor g10514(.dina(n28425), .dinb(n440), .dout(n28537));
  jnot g10515(.din(n28537), .dout(n28538));
  jor  g10516(.dina(n28538), .dinb(n28536), .dout(n28539));
  jand g10517(.dina(n28539), .dinb(n28427), .dout(n28540));
  jxor g10518(.dina(n28419), .dinb(n435), .dout(n28541));
  jnot g10519(.din(n28541), .dout(n28542));
  jor  g10520(.dina(n28542), .dinb(n28540), .dout(n28543));
  jand g10521(.dina(n28543), .dinb(n28421), .dout(n28544));
  jxor g10522(.dina(n28413), .dinb(n436), .dout(n28545));
  jnot g10523(.din(n28545), .dout(n28546));
  jor  g10524(.dina(n28546), .dinb(n28544), .dout(n28547));
  jand g10525(.dina(n28547), .dinb(n28415), .dout(n28548));
  jxor g10526(.dina(n28407), .dinb(n432), .dout(n28549));
  jnot g10527(.din(n28549), .dout(n28550));
  jor  g10528(.dina(n28550), .dinb(n28548), .dout(n28551));
  jand g10529(.dina(n28551), .dinb(n28409), .dout(n28552));
  jxor g10530(.dina(n28401), .dinb(n433), .dout(n28553));
  jnot g10531(.din(n28553), .dout(n28554));
  jor  g10532(.dina(n28554), .dinb(n28552), .dout(n28555));
  jand g10533(.dina(n28555), .dinb(n28403), .dout(n28556));
  jxor g10534(.dina(n28395), .dinb(n421), .dout(n28557));
  jnot g10535(.din(n28557), .dout(n28558));
  jor  g10536(.dina(n28558), .dinb(n28556), .dout(n28559));
  jand g10537(.dina(n28559), .dinb(n28397), .dout(n28560));
  jxor g10538(.dina(n28389), .dinb(n422), .dout(n28561));
  jnot g10539(.din(n28561), .dout(n28562));
  jor  g10540(.dina(n28562), .dinb(n28560), .dout(n28563));
  jand g10541(.dina(n28563), .dinb(n28391), .dout(n28564));
  jxor g10542(.dina(n28383), .dinb(n416), .dout(n28565));
  jnot g10543(.din(n28565), .dout(n28566));
  jor  g10544(.dina(n28566), .dinb(n28564), .dout(n28567));
  jand g10545(.dina(n28567), .dinb(n28385), .dout(n28568));
  jxor g10546(.dina(n28377), .dinb(n417), .dout(n28569));
  jnot g10547(.din(n28569), .dout(n28570));
  jor  g10548(.dina(n28570), .dinb(n28568), .dout(n28571));
  jand g10549(.dina(n28571), .dinb(n28379), .dout(n28572));
  jxor g10550(.dina(n28371), .dinb(n2547), .dout(n28573));
  jnot g10551(.din(n28573), .dout(n28574));
  jor  g10552(.dina(n28574), .dinb(n28572), .dout(n28575));
  jand g10553(.dina(n28575), .dinb(n28373), .dout(n28576));
  jxor g10554(.dina(n28365), .dinb(n2714), .dout(n28577));
  jnot g10555(.din(n28577), .dout(n28578));
  jor  g10556(.dina(n28578), .dinb(n28576), .dout(n28579));
  jand g10557(.dina(n28579), .dinb(n28367), .dout(n28580));
  jxor g10558(.dina(n28359), .dinb(n405), .dout(n28581));
  jnot g10559(.din(n28581), .dout(n28582));
  jor  g10560(.dina(n28582), .dinb(n28580), .dout(n28583));
  jand g10561(.dina(n28583), .dinb(n28361), .dout(n28584));
  jxor g10562(.dina(n28353), .dinb(n406), .dout(n28585));
  jnot g10563(.din(n28585), .dout(n28586));
  jor  g10564(.dina(n28586), .dinb(n28584), .dout(n28587));
  jand g10565(.dina(n28587), .dinb(n28355), .dout(n28588));
  jxor g10566(.dina(n28347), .dinb(n412), .dout(n28589));
  jnot g10567(.din(n28589), .dout(n28590));
  jor  g10568(.dina(n28590), .dinb(n28588), .dout(n28591));
  jand g10569(.dina(n28591), .dinb(n28349), .dout(n28592));
  jxor g10570(.dina(n28341), .dinb(n413), .dout(n28593));
  jnot g10571(.din(n28593), .dout(n28594));
  jor  g10572(.dina(n28594), .dinb(n28592), .dout(n28595));
  jand g10573(.dina(n28595), .dinb(n28343), .dout(n28596));
  jxor g10574(.dina(n28335), .dinb(n409), .dout(n28597));
  jnot g10575(.din(n28597), .dout(n28598));
  jor  g10576(.dina(n28598), .dinb(n28596), .dout(n28599));
  jand g10577(.dina(n28599), .dinb(n28337), .dout(n28600));
  jxor g10578(.dina(n28329), .dinb(n410), .dout(n28601));
  jnot g10579(.din(n28601), .dout(n28602));
  jor  g10580(.dina(n28602), .dinb(n28600), .dout(n28603));
  jand g10581(.dina(n28603), .dinb(n28331), .dout(n28604));
  jxor g10582(.dina(n28323), .dinb(n426), .dout(n28605));
  jnot g10583(.din(n28605), .dout(n28606));
  jor  g10584(.dina(n28606), .dinb(n28604), .dout(n28607));
  jand g10585(.dina(n28607), .dinb(n28325), .dout(n28608));
  jxor g10586(.dina(n28317), .dinb(n427), .dout(n28609));
  jnot g10587(.din(n28609), .dout(n28610));
  jor  g10588(.dina(n28610), .dinb(n28608), .dout(n28611));
  jand g10589(.dina(n28611), .dinb(n28319), .dout(n28612));
  jxor g10590(.dina(n28311), .dinb(n424), .dout(n28613));
  jnot g10591(.din(n28613), .dout(n28614));
  jor  g10592(.dina(n28614), .dinb(n28612), .dout(n28615));
  jand g10593(.dina(n28615), .dinb(n28313), .dout(n28616));
  jxor g10594(.dina(n28305), .dinb(n300), .dout(n28617));
  jnot g10595(.din(n28617), .dout(n28618));
  jor  g10596(.dina(n28618), .dinb(n28616), .dout(n28619));
  jand g10597(.dina(n28619), .dinb(n28307), .dout(n28620));
  jxor g10598(.dina(n28299), .dinb(n297), .dout(n28621));
  jnot g10599(.din(n28621), .dout(n28622));
  jor  g10600(.dina(n28622), .dinb(n28620), .dout(n28623));
  jand g10601(.dina(n28623), .dinb(n28301), .dout(n28624));
  jxor g10602(.dina(n28293), .dinb(n298), .dout(n28625));
  jnot g10603(.din(n28625), .dout(n28626));
  jor  g10604(.dina(n28626), .dinb(n28624), .dout(n28627));
  jand g10605(.dina(n28627), .dinb(n28295), .dout(n28628));
  jxor g10606(.dina(n28287), .dinb(n301), .dout(n28629));
  jnot g10607(.din(n28629), .dout(n28630));
  jor  g10608(.dina(n28630), .dinb(n28628), .dout(n28631));
  jand g10609(.dina(n28631), .dinb(n28289), .dout(n28632));
  jxor g10610(.dina(n28281), .dinb(n293), .dout(n28633));
  jnot g10611(.din(n28633), .dout(n28634));
  jor  g10612(.dina(n28634), .dinb(n28632), .dout(n28635));
  jand g10613(.dina(n28635), .dinb(n28283), .dout(n28636));
  jxor g10614(.dina(n28275), .dinb(n294), .dout(n28637));
  jnot g10615(.din(n28637), .dout(n28638));
  jor  g10616(.dina(n28638), .dinb(n28636), .dout(n28639));
  jand g10617(.dina(n28639), .dinb(n28277), .dout(n28640));
  jxor g10618(.dina(n28269), .dinb(n290), .dout(n28641));
  jnot g10619(.din(n28641), .dout(n28642));
  jor  g10620(.dina(n28642), .dinb(n28640), .dout(n28643));
  jand g10621(.dina(n28643), .dinb(n28271), .dout(n28644));
  jxor g10622(.dina(n28263), .dinb(n291), .dout(n28645));
  jnot g10623(.din(n28645), .dout(n28646));
  jor  g10624(.dina(n28646), .dinb(n28644), .dout(n28647));
  jand g10625(.dina(n28647), .dinb(n28265), .dout(n28648));
  jnot g10626(.din(n28253), .dout(n28649));
  jand g10627(.dina(n28649), .dinb(b40 ), .dout(n28650));
  jor  g10628(.dina(n28650), .dinb(n28648), .dout(n28651));
  jand g10629(.dina(n28651), .dinb(n28255), .dout(n28652));
  jor  g10630(.dina(n28652), .dinb(n7960), .dout(n28653));
  jand g10631(.dina(n28653), .dinb(n28253), .dout(n28654));
  jnot g10632(.din(n28482), .dout(n28655));
  jnot g10633(.din(n7355), .dout(n28656));
  jor  g10634(.dina(n28166), .dinb(n28656), .dout(n28657));
  jand g10635(.dina(n28657), .dinb(a24 ), .dout(n28658));
  jand g10636(.dina(n28260), .dinb(n7723), .dout(n28659));
  jor  g10637(.dina(n28659), .dinb(n28658), .dout(n28660));
  jand g10638(.dina(n28660), .dinb(n258), .dout(n28661));
  jxor g10639(.dina(n28492), .dinb(b1 ), .dout(n28662));
  jand g10640(.dina(n28662), .dinb(n8369), .dout(n28663));
  jor  g10641(.dina(n28663), .dinb(n28661), .dout(n28664));
  jand g10642(.dina(n28497), .dinb(n28664), .dout(n28665));
  jor  g10643(.dina(n28665), .dinb(n28487), .dout(n28666));
  jand g10644(.dina(n28501), .dinb(n28666), .dout(n28667));
  jor  g10645(.dina(n28667), .dinb(n28655), .dout(n28668));
  jand g10646(.dina(n28505), .dinb(n28668), .dout(n28669));
  jor  g10647(.dina(n28669), .dinb(n28474), .dout(n28670));
  jand g10648(.dina(n28509), .dinb(n28670), .dout(n28671));
  jor  g10649(.dina(n28671), .dinb(n28468), .dout(n28672));
  jand g10650(.dina(n28513), .dinb(n28672), .dout(n28673));
  jor  g10651(.dina(n28673), .dinb(n28462), .dout(n28674));
  jand g10652(.dina(n28517), .dinb(n28674), .dout(n28675));
  jor  g10653(.dina(n28675), .dinb(n28456), .dout(n28676));
  jand g10654(.dina(n28521), .dinb(n28676), .dout(n28677));
  jor  g10655(.dina(n28677), .dinb(n28450), .dout(n28678));
  jand g10656(.dina(n28525), .dinb(n28678), .dout(n28679));
  jor  g10657(.dina(n28679), .dinb(n28444), .dout(n28680));
  jand g10658(.dina(n28529), .dinb(n28680), .dout(n28681));
  jor  g10659(.dina(n28681), .dinb(n28438), .dout(n28682));
  jand g10660(.dina(n28533), .dinb(n28682), .dout(n28683));
  jor  g10661(.dina(n28683), .dinb(n28432), .dout(n28684));
  jand g10662(.dina(n28537), .dinb(n28684), .dout(n28685));
  jor  g10663(.dina(n28685), .dinb(n28426), .dout(n28686));
  jand g10664(.dina(n28541), .dinb(n28686), .dout(n28687));
  jor  g10665(.dina(n28687), .dinb(n28420), .dout(n28688));
  jand g10666(.dina(n28545), .dinb(n28688), .dout(n28689));
  jor  g10667(.dina(n28689), .dinb(n28414), .dout(n28690));
  jand g10668(.dina(n28549), .dinb(n28690), .dout(n28691));
  jor  g10669(.dina(n28691), .dinb(n28408), .dout(n28692));
  jand g10670(.dina(n28553), .dinb(n28692), .dout(n28693));
  jor  g10671(.dina(n28693), .dinb(n28402), .dout(n28694));
  jand g10672(.dina(n28557), .dinb(n28694), .dout(n28695));
  jor  g10673(.dina(n28695), .dinb(n28396), .dout(n28696));
  jand g10674(.dina(n28561), .dinb(n28696), .dout(n28697));
  jor  g10675(.dina(n28697), .dinb(n28390), .dout(n28698));
  jand g10676(.dina(n28565), .dinb(n28698), .dout(n28699));
  jor  g10677(.dina(n28699), .dinb(n28384), .dout(n28700));
  jand g10678(.dina(n28569), .dinb(n28700), .dout(n28701));
  jor  g10679(.dina(n28701), .dinb(n28378), .dout(n28702));
  jand g10680(.dina(n28573), .dinb(n28702), .dout(n28703));
  jor  g10681(.dina(n28703), .dinb(n28372), .dout(n28704));
  jand g10682(.dina(n28577), .dinb(n28704), .dout(n28705));
  jor  g10683(.dina(n28705), .dinb(n28366), .dout(n28706));
  jand g10684(.dina(n28581), .dinb(n28706), .dout(n28707));
  jor  g10685(.dina(n28707), .dinb(n28360), .dout(n28708));
  jand g10686(.dina(n28585), .dinb(n28708), .dout(n28709));
  jor  g10687(.dina(n28709), .dinb(n28354), .dout(n28710));
  jand g10688(.dina(n28589), .dinb(n28710), .dout(n28711));
  jor  g10689(.dina(n28711), .dinb(n28348), .dout(n28712));
  jand g10690(.dina(n28593), .dinb(n28712), .dout(n28713));
  jor  g10691(.dina(n28713), .dinb(n28342), .dout(n28714));
  jand g10692(.dina(n28597), .dinb(n28714), .dout(n28715));
  jor  g10693(.dina(n28715), .dinb(n28336), .dout(n28716));
  jand g10694(.dina(n28601), .dinb(n28716), .dout(n28717));
  jor  g10695(.dina(n28717), .dinb(n28330), .dout(n28718));
  jand g10696(.dina(n28605), .dinb(n28718), .dout(n28719));
  jor  g10697(.dina(n28719), .dinb(n28324), .dout(n28720));
  jand g10698(.dina(n28609), .dinb(n28720), .dout(n28721));
  jor  g10699(.dina(n28721), .dinb(n28318), .dout(n28722));
  jand g10700(.dina(n28613), .dinb(n28722), .dout(n28723));
  jor  g10701(.dina(n28723), .dinb(n28312), .dout(n28724));
  jand g10702(.dina(n28617), .dinb(n28724), .dout(n28725));
  jor  g10703(.dina(n28725), .dinb(n28306), .dout(n28726));
  jand g10704(.dina(n28621), .dinb(n28726), .dout(n28727));
  jor  g10705(.dina(n28727), .dinb(n28300), .dout(n28728));
  jand g10706(.dina(n28625), .dinb(n28728), .dout(n28729));
  jor  g10707(.dina(n28729), .dinb(n28294), .dout(n28730));
  jand g10708(.dina(n28629), .dinb(n28730), .dout(n28731));
  jor  g10709(.dina(n28731), .dinb(n28288), .dout(n28732));
  jand g10710(.dina(n28633), .dinb(n28732), .dout(n28733));
  jor  g10711(.dina(n28733), .dinb(n28282), .dout(n28734));
  jand g10712(.dina(n28637), .dinb(n28734), .dout(n28735));
  jor  g10713(.dina(n28735), .dinb(n28276), .dout(n28736));
  jand g10714(.dina(n28641), .dinb(n28736), .dout(n28737));
  jor  g10715(.dina(n28737), .dinb(n28270), .dout(n28738));
  jand g10716(.dina(n28645), .dinb(n28738), .dout(n28739));
  jor  g10717(.dina(n28739), .dinb(n28264), .dout(n28740));
  jand g10718(.dina(n28254), .dinb(n518), .dout(n28741));
  jand g10719(.dina(n28741), .dinb(n28740), .dout(n28742));
  jor  g10720(.dina(n28742), .dinb(n28654), .dout(n28743));
  jnot g10721(.din(n28743), .dout(n28744));
  jand g10722(.dina(n28653), .dinb(n28263), .dout(n28745));
  jnot g10723(.din(n28650), .dout(n28746));
  jand g10724(.dina(n28746), .dinb(n28740), .dout(n28747));
  jor  g10725(.dina(n28747), .dinb(n28254), .dout(n28748));
  jand g10726(.dina(n28748), .dinb(n518), .dout(n28749));
  jxor g10727(.dina(n28645), .dinb(n28738), .dout(n28750));
  jand g10728(.dina(n28750), .dinb(n28749), .dout(n28751));
  jor  g10729(.dina(n28751), .dinb(n28745), .dout(n28752));
  jand g10730(.dina(n28752), .dinb(n284), .dout(n28753));
  jnot g10731(.din(n28753), .dout(n28754));
  jand g10732(.dina(n28653), .dinb(n28269), .dout(n28755));
  jxor g10733(.dina(n28641), .dinb(n28736), .dout(n28756));
  jand g10734(.dina(n28756), .dinb(n28749), .dout(n28757));
  jor  g10735(.dina(n28757), .dinb(n28755), .dout(n28758));
  jand g10736(.dina(n28758), .dinb(n291), .dout(n28759));
  jnot g10737(.din(n28759), .dout(n28760));
  jand g10738(.dina(n28653), .dinb(n28275), .dout(n28761));
  jxor g10739(.dina(n28637), .dinb(n28734), .dout(n28762));
  jand g10740(.dina(n28762), .dinb(n28749), .dout(n28763));
  jor  g10741(.dina(n28763), .dinb(n28761), .dout(n28764));
  jand g10742(.dina(n28764), .dinb(n290), .dout(n28765));
  jnot g10743(.din(n28765), .dout(n28766));
  jand g10744(.dina(n28653), .dinb(n28281), .dout(n28767));
  jxor g10745(.dina(n28633), .dinb(n28732), .dout(n28768));
  jand g10746(.dina(n28768), .dinb(n28749), .dout(n28769));
  jor  g10747(.dina(n28769), .dinb(n28767), .dout(n28770));
  jand g10748(.dina(n28770), .dinb(n294), .dout(n28771));
  jnot g10749(.din(n28771), .dout(n28772));
  jand g10750(.dina(n28653), .dinb(n28287), .dout(n28773));
  jxor g10751(.dina(n28629), .dinb(n28730), .dout(n28774));
  jand g10752(.dina(n28774), .dinb(n28749), .dout(n28775));
  jor  g10753(.dina(n28775), .dinb(n28773), .dout(n28776));
  jand g10754(.dina(n28776), .dinb(n293), .dout(n28777));
  jnot g10755(.din(n28777), .dout(n28778));
  jand g10756(.dina(n28653), .dinb(n28293), .dout(n28779));
  jxor g10757(.dina(n28625), .dinb(n28728), .dout(n28780));
  jand g10758(.dina(n28780), .dinb(n28749), .dout(n28781));
  jor  g10759(.dina(n28781), .dinb(n28779), .dout(n28782));
  jand g10760(.dina(n28782), .dinb(n301), .dout(n28783));
  jnot g10761(.din(n28783), .dout(n28784));
  jand g10762(.dina(n28653), .dinb(n28299), .dout(n28785));
  jxor g10763(.dina(n28621), .dinb(n28726), .dout(n28786));
  jand g10764(.dina(n28786), .dinb(n28749), .dout(n28787));
  jor  g10765(.dina(n28787), .dinb(n28785), .dout(n28788));
  jand g10766(.dina(n28788), .dinb(n298), .dout(n28789));
  jnot g10767(.din(n28789), .dout(n28790));
  jand g10768(.dina(n28653), .dinb(n28305), .dout(n28791));
  jxor g10769(.dina(n28617), .dinb(n28724), .dout(n28792));
  jand g10770(.dina(n28792), .dinb(n28749), .dout(n28793));
  jor  g10771(.dina(n28793), .dinb(n28791), .dout(n28794));
  jand g10772(.dina(n28794), .dinb(n297), .dout(n28795));
  jnot g10773(.din(n28795), .dout(n28796));
  jand g10774(.dina(n28653), .dinb(n28311), .dout(n28797));
  jxor g10775(.dina(n28613), .dinb(n28722), .dout(n28798));
  jand g10776(.dina(n28798), .dinb(n28749), .dout(n28799));
  jor  g10777(.dina(n28799), .dinb(n28797), .dout(n28800));
  jand g10778(.dina(n28800), .dinb(n300), .dout(n28801));
  jnot g10779(.din(n28801), .dout(n28802));
  jand g10780(.dina(n28653), .dinb(n28317), .dout(n28803));
  jxor g10781(.dina(n28609), .dinb(n28720), .dout(n28804));
  jand g10782(.dina(n28804), .dinb(n28749), .dout(n28805));
  jor  g10783(.dina(n28805), .dinb(n28803), .dout(n28806));
  jand g10784(.dina(n28806), .dinb(n424), .dout(n28807));
  jnot g10785(.din(n28807), .dout(n28808));
  jand g10786(.dina(n28653), .dinb(n28323), .dout(n28809));
  jxor g10787(.dina(n28605), .dinb(n28718), .dout(n28810));
  jand g10788(.dina(n28810), .dinb(n28749), .dout(n28811));
  jor  g10789(.dina(n28811), .dinb(n28809), .dout(n28812));
  jand g10790(.dina(n28812), .dinb(n427), .dout(n28813));
  jnot g10791(.din(n28813), .dout(n28814));
  jand g10792(.dina(n28653), .dinb(n28329), .dout(n28815));
  jxor g10793(.dina(n28601), .dinb(n28716), .dout(n28816));
  jand g10794(.dina(n28816), .dinb(n28749), .dout(n28817));
  jor  g10795(.dina(n28817), .dinb(n28815), .dout(n28818));
  jand g10796(.dina(n28818), .dinb(n426), .dout(n28819));
  jnot g10797(.din(n28819), .dout(n28820));
  jand g10798(.dina(n28653), .dinb(n28335), .dout(n28821));
  jxor g10799(.dina(n28597), .dinb(n28714), .dout(n28822));
  jand g10800(.dina(n28822), .dinb(n28749), .dout(n28823));
  jor  g10801(.dina(n28823), .dinb(n28821), .dout(n28824));
  jand g10802(.dina(n28824), .dinb(n410), .dout(n28825));
  jnot g10803(.din(n28825), .dout(n28826));
  jand g10804(.dina(n28653), .dinb(n28341), .dout(n28827));
  jxor g10805(.dina(n28593), .dinb(n28712), .dout(n28828));
  jand g10806(.dina(n28828), .dinb(n28749), .dout(n28829));
  jor  g10807(.dina(n28829), .dinb(n28827), .dout(n28830));
  jand g10808(.dina(n28830), .dinb(n409), .dout(n28831));
  jnot g10809(.din(n28831), .dout(n28832));
  jand g10810(.dina(n28653), .dinb(n28347), .dout(n28833));
  jxor g10811(.dina(n28589), .dinb(n28710), .dout(n28834));
  jand g10812(.dina(n28834), .dinb(n28749), .dout(n28835));
  jor  g10813(.dina(n28835), .dinb(n28833), .dout(n28836));
  jand g10814(.dina(n28836), .dinb(n413), .dout(n28837));
  jnot g10815(.din(n28837), .dout(n28838));
  jand g10816(.dina(n28653), .dinb(n28353), .dout(n28839));
  jxor g10817(.dina(n28585), .dinb(n28708), .dout(n28840));
  jand g10818(.dina(n28840), .dinb(n28749), .dout(n28841));
  jor  g10819(.dina(n28841), .dinb(n28839), .dout(n28842));
  jand g10820(.dina(n28842), .dinb(n412), .dout(n28843));
  jnot g10821(.din(n28843), .dout(n28844));
  jand g10822(.dina(n28653), .dinb(n28359), .dout(n28845));
  jxor g10823(.dina(n28581), .dinb(n28706), .dout(n28846));
  jand g10824(.dina(n28846), .dinb(n28749), .dout(n28847));
  jor  g10825(.dina(n28847), .dinb(n28845), .dout(n28848));
  jand g10826(.dina(n28848), .dinb(n406), .dout(n28849));
  jnot g10827(.din(n28849), .dout(n28850));
  jand g10828(.dina(n28653), .dinb(n28365), .dout(n28851));
  jxor g10829(.dina(n28577), .dinb(n28704), .dout(n28852));
  jand g10830(.dina(n28852), .dinb(n28749), .dout(n28853));
  jor  g10831(.dina(n28853), .dinb(n28851), .dout(n28854));
  jand g10832(.dina(n28854), .dinb(n405), .dout(n28855));
  jnot g10833(.din(n28855), .dout(n28856));
  jand g10834(.dina(n28653), .dinb(n28371), .dout(n28857));
  jxor g10835(.dina(n28573), .dinb(n28702), .dout(n28858));
  jand g10836(.dina(n28858), .dinb(n28749), .dout(n28859));
  jor  g10837(.dina(n28859), .dinb(n28857), .dout(n28860));
  jand g10838(.dina(n28860), .dinb(n2714), .dout(n28861));
  jnot g10839(.din(n28861), .dout(n28862));
  jand g10840(.dina(n28653), .dinb(n28377), .dout(n28863));
  jxor g10841(.dina(n28569), .dinb(n28700), .dout(n28864));
  jand g10842(.dina(n28864), .dinb(n28749), .dout(n28865));
  jor  g10843(.dina(n28865), .dinb(n28863), .dout(n28866));
  jand g10844(.dina(n28866), .dinb(n2547), .dout(n28867));
  jnot g10845(.din(n28867), .dout(n28868));
  jand g10846(.dina(n28653), .dinb(n28383), .dout(n28869));
  jxor g10847(.dina(n28565), .dinb(n28698), .dout(n28870));
  jand g10848(.dina(n28870), .dinb(n28749), .dout(n28871));
  jor  g10849(.dina(n28871), .dinb(n28869), .dout(n28872));
  jand g10850(.dina(n28872), .dinb(n417), .dout(n28873));
  jnot g10851(.din(n28873), .dout(n28874));
  jand g10852(.dina(n28653), .dinb(n28389), .dout(n28875));
  jxor g10853(.dina(n28561), .dinb(n28696), .dout(n28876));
  jand g10854(.dina(n28876), .dinb(n28749), .dout(n28877));
  jor  g10855(.dina(n28877), .dinb(n28875), .dout(n28878));
  jand g10856(.dina(n28878), .dinb(n416), .dout(n28879));
  jnot g10857(.din(n28879), .dout(n28880));
  jand g10858(.dina(n28653), .dinb(n28395), .dout(n28881));
  jxor g10859(.dina(n28557), .dinb(n28694), .dout(n28882));
  jand g10860(.dina(n28882), .dinb(n28749), .dout(n28883));
  jor  g10861(.dina(n28883), .dinb(n28881), .dout(n28884));
  jand g10862(.dina(n28884), .dinb(n422), .dout(n28885));
  jnot g10863(.din(n28885), .dout(n28886));
  jand g10864(.dina(n28653), .dinb(n28401), .dout(n28887));
  jxor g10865(.dina(n28553), .dinb(n28692), .dout(n28888));
  jand g10866(.dina(n28888), .dinb(n28749), .dout(n28889));
  jor  g10867(.dina(n28889), .dinb(n28887), .dout(n28890));
  jand g10868(.dina(n28890), .dinb(n421), .dout(n28891));
  jnot g10869(.din(n28891), .dout(n28892));
  jand g10870(.dina(n28653), .dinb(n28407), .dout(n28893));
  jxor g10871(.dina(n28549), .dinb(n28690), .dout(n28894));
  jand g10872(.dina(n28894), .dinb(n28749), .dout(n28895));
  jor  g10873(.dina(n28895), .dinb(n28893), .dout(n28896));
  jand g10874(.dina(n28896), .dinb(n433), .dout(n28897));
  jnot g10875(.din(n28897), .dout(n28898));
  jand g10876(.dina(n28653), .dinb(n28413), .dout(n28899));
  jxor g10877(.dina(n28545), .dinb(n28688), .dout(n28900));
  jand g10878(.dina(n28900), .dinb(n28749), .dout(n28901));
  jor  g10879(.dina(n28901), .dinb(n28899), .dout(n28902));
  jand g10880(.dina(n28902), .dinb(n432), .dout(n28903));
  jnot g10881(.din(n28903), .dout(n28904));
  jand g10882(.dina(n28653), .dinb(n28419), .dout(n28905));
  jxor g10883(.dina(n28541), .dinb(n28686), .dout(n28906));
  jand g10884(.dina(n28906), .dinb(n28749), .dout(n28907));
  jor  g10885(.dina(n28907), .dinb(n28905), .dout(n28908));
  jand g10886(.dina(n28908), .dinb(n436), .dout(n28909));
  jnot g10887(.din(n28909), .dout(n28910));
  jand g10888(.dina(n28653), .dinb(n28425), .dout(n28911));
  jxor g10889(.dina(n28537), .dinb(n28684), .dout(n28912));
  jand g10890(.dina(n28912), .dinb(n28749), .dout(n28913));
  jor  g10891(.dina(n28913), .dinb(n28911), .dout(n28914));
  jand g10892(.dina(n28914), .dinb(n435), .dout(n28915));
  jnot g10893(.din(n28915), .dout(n28916));
  jand g10894(.dina(n28653), .dinb(n28431), .dout(n28917));
  jxor g10895(.dina(n28533), .dinb(n28682), .dout(n28918));
  jand g10896(.dina(n28918), .dinb(n28749), .dout(n28919));
  jor  g10897(.dina(n28919), .dinb(n28917), .dout(n28920));
  jand g10898(.dina(n28920), .dinb(n440), .dout(n28921));
  jnot g10899(.din(n28921), .dout(n28922));
  jand g10900(.dina(n28653), .dinb(n28437), .dout(n28923));
  jxor g10901(.dina(n28529), .dinb(n28680), .dout(n28924));
  jand g10902(.dina(n28924), .dinb(n28749), .dout(n28925));
  jor  g10903(.dina(n28925), .dinb(n28923), .dout(n28926));
  jand g10904(.dina(n28926), .dinb(n439), .dout(n28927));
  jnot g10905(.din(n28927), .dout(n28928));
  jand g10906(.dina(n28653), .dinb(n28443), .dout(n28929));
  jxor g10907(.dina(n28525), .dinb(n28678), .dout(n28930));
  jand g10908(.dina(n28930), .dinb(n28749), .dout(n28931));
  jor  g10909(.dina(n28931), .dinb(n28929), .dout(n28932));
  jand g10910(.dina(n28932), .dinb(n325), .dout(n28933));
  jnot g10911(.din(n28933), .dout(n28934));
  jand g10912(.dina(n28653), .dinb(n28449), .dout(n28935));
  jxor g10913(.dina(n28521), .dinb(n28676), .dout(n28936));
  jand g10914(.dina(n28936), .dinb(n28749), .dout(n28937));
  jor  g10915(.dina(n28937), .dinb(n28935), .dout(n28938));
  jand g10916(.dina(n28938), .dinb(n324), .dout(n28939));
  jnot g10917(.din(n28939), .dout(n28940));
  jand g10918(.dina(n28653), .dinb(n28455), .dout(n28941));
  jxor g10919(.dina(n28517), .dinb(n28674), .dout(n28942));
  jand g10920(.dina(n28942), .dinb(n28749), .dout(n28943));
  jor  g10921(.dina(n28943), .dinb(n28941), .dout(n28944));
  jand g10922(.dina(n28944), .dinb(n323), .dout(n28945));
  jnot g10923(.din(n28945), .dout(n28946));
  jand g10924(.dina(n28653), .dinb(n28461), .dout(n28947));
  jxor g10925(.dina(n28513), .dinb(n28672), .dout(n28948));
  jand g10926(.dina(n28948), .dinb(n28749), .dout(n28949));
  jor  g10927(.dina(n28949), .dinb(n28947), .dout(n28950));
  jand g10928(.dina(n28950), .dinb(n335), .dout(n28951));
  jnot g10929(.din(n28951), .dout(n28952));
  jand g10930(.dina(n28653), .dinb(n28467), .dout(n28953));
  jxor g10931(.dina(n28509), .dinb(n28670), .dout(n28954));
  jand g10932(.dina(n28954), .dinb(n28749), .dout(n28955));
  jor  g10933(.dina(n28955), .dinb(n28953), .dout(n28956));
  jand g10934(.dina(n28956), .dinb(n334), .dout(n28957));
  jnot g10935(.din(n28957), .dout(n28958));
  jand g10936(.dina(n28653), .dinb(n28473), .dout(n28959));
  jxor g10937(.dina(n28505), .dinb(n28668), .dout(n28960));
  jand g10938(.dina(n28960), .dinb(n28749), .dout(n28961));
  jor  g10939(.dina(n28961), .dinb(n28959), .dout(n28962));
  jand g10940(.dina(n28962), .dinb(n338), .dout(n28963));
  jnot g10941(.din(n28963), .dout(n28964));
  jor  g10942(.dina(n28749), .dinb(n28481), .dout(n28965));
  jxor g10943(.dina(n28501), .dinb(n28666), .dout(n28966));
  jand g10944(.dina(n28966), .dinb(n28749), .dout(n28967));
  jnot g10945(.din(n28967), .dout(n28968));
  jand g10946(.dina(n28968), .dinb(n28965), .dout(n28969));
  jnot g10947(.din(n28969), .dout(n28970));
  jand g10948(.dina(n28970), .dinb(n337), .dout(n28971));
  jnot g10949(.din(n28971), .dout(n28972));
  jnot g10950(.din(n28486), .dout(n28973));
  jor  g10951(.dina(n28749), .dinb(n28973), .dout(n28974));
  jxor g10952(.dina(n28497), .dinb(n28664), .dout(n28975));
  jnot g10953(.din(n28975), .dout(n28976));
  jor  g10954(.dina(n28976), .dinb(n28653), .dout(n28977));
  jand g10955(.dina(n28977), .dinb(n28974), .dout(n28978));
  jnot g10956(.din(n28978), .dout(n28979));
  jand g10957(.dina(n28979), .dinb(n344), .dout(n28980));
  jnot g10958(.din(n28980), .dout(n28981));
  jand g10959(.dina(n28653), .dinb(n28660), .dout(n28982));
  jxor g10960(.dina(n28662), .dinb(n8369), .dout(n28983));
  jand g10961(.dina(n28983), .dinb(n28749), .dout(n28984));
  jor  g10962(.dina(n28984), .dinb(n28982), .dout(n28985));
  jand g10963(.dina(n28985), .dinb(n348), .dout(n28986));
  jnot g10964(.din(n28986), .dout(n28987));
  jnot g10965(.din(n8660), .dout(n28988));
  jor  g10966(.dina(n28652), .dinb(n28988), .dout(n28989));
  jand g10967(.dina(n28989), .dinb(a23 ), .dout(n28990));
  jand g10968(.dina(n28749), .dinb(n8204), .dout(n28991));
  jor  g10969(.dina(n28991), .dinb(n28990), .dout(n28992));
  jand g10970(.dina(n28992), .dinb(n258), .dout(n28993));
  jnot g10971(.din(n28993), .dout(n28994));
  jand g10972(.dina(n28748), .dinb(n8660), .dout(n28995));
  jor  g10973(.dina(n28995), .dinb(n8203), .dout(n28996));
  jor  g10974(.dina(n28653), .dinb(n8369), .dout(n28997));
  jand g10975(.dina(n28997), .dinb(n28996), .dout(n28998));
  jxor g10976(.dina(n28998), .dinb(n258), .dout(n28999));
  jor  g10977(.dina(n28999), .dinb(n8668), .dout(n29000));
  jand g10978(.dina(n29000), .dinb(n28994), .dout(n29001));
  jxor g10979(.dina(n28985), .dinb(n348), .dout(n29002));
  jnot g10980(.din(n29002), .dout(n29003));
  jor  g10981(.dina(n29003), .dinb(n29001), .dout(n29004));
  jand g10982(.dina(n29004), .dinb(n28987), .dout(n29005));
  jxor g10983(.dina(n28978), .dinb(b3 ), .dout(n29006));
  jnot g10984(.din(n29006), .dout(n29007));
  jor  g10985(.dina(n29007), .dinb(n29005), .dout(n29008));
  jand g10986(.dina(n29008), .dinb(n28981), .dout(n29009));
  jxor g10987(.dina(n28969), .dinb(b4 ), .dout(n29010));
  jnot g10988(.din(n29010), .dout(n29011));
  jor  g10989(.dina(n29011), .dinb(n29009), .dout(n29012));
  jand g10990(.dina(n29012), .dinb(n28972), .dout(n29013));
  jxor g10991(.dina(n28962), .dinb(n338), .dout(n29014));
  jnot g10992(.din(n29014), .dout(n29015));
  jor  g10993(.dina(n29015), .dinb(n29013), .dout(n29016));
  jand g10994(.dina(n29016), .dinb(n28964), .dout(n29017));
  jxor g10995(.dina(n28956), .dinb(n334), .dout(n29018));
  jnot g10996(.din(n29018), .dout(n29019));
  jor  g10997(.dina(n29019), .dinb(n29017), .dout(n29020));
  jand g10998(.dina(n29020), .dinb(n28958), .dout(n29021));
  jxor g10999(.dina(n28950), .dinb(n335), .dout(n29022));
  jnot g11000(.din(n29022), .dout(n29023));
  jor  g11001(.dina(n29023), .dinb(n29021), .dout(n29024));
  jand g11002(.dina(n29024), .dinb(n28952), .dout(n29025));
  jxor g11003(.dina(n28944), .dinb(n323), .dout(n29026));
  jnot g11004(.din(n29026), .dout(n29027));
  jor  g11005(.dina(n29027), .dinb(n29025), .dout(n29028));
  jand g11006(.dina(n29028), .dinb(n28946), .dout(n29029));
  jxor g11007(.dina(n28938), .dinb(n324), .dout(n29030));
  jnot g11008(.din(n29030), .dout(n29031));
  jor  g11009(.dina(n29031), .dinb(n29029), .dout(n29032));
  jand g11010(.dina(n29032), .dinb(n28940), .dout(n29033));
  jxor g11011(.dina(n28932), .dinb(n325), .dout(n29034));
  jnot g11012(.din(n29034), .dout(n29035));
  jor  g11013(.dina(n29035), .dinb(n29033), .dout(n29036));
  jand g11014(.dina(n29036), .dinb(n28934), .dout(n29037));
  jxor g11015(.dina(n28926), .dinb(n439), .dout(n29038));
  jnot g11016(.din(n29038), .dout(n29039));
  jor  g11017(.dina(n29039), .dinb(n29037), .dout(n29040));
  jand g11018(.dina(n29040), .dinb(n28928), .dout(n29041));
  jxor g11019(.dina(n28920), .dinb(n440), .dout(n29042));
  jnot g11020(.din(n29042), .dout(n29043));
  jor  g11021(.dina(n29043), .dinb(n29041), .dout(n29044));
  jand g11022(.dina(n29044), .dinb(n28922), .dout(n29045));
  jxor g11023(.dina(n28914), .dinb(n435), .dout(n29046));
  jnot g11024(.din(n29046), .dout(n29047));
  jor  g11025(.dina(n29047), .dinb(n29045), .dout(n29048));
  jand g11026(.dina(n29048), .dinb(n28916), .dout(n29049));
  jxor g11027(.dina(n28908), .dinb(n436), .dout(n29050));
  jnot g11028(.din(n29050), .dout(n29051));
  jor  g11029(.dina(n29051), .dinb(n29049), .dout(n29052));
  jand g11030(.dina(n29052), .dinb(n28910), .dout(n29053));
  jxor g11031(.dina(n28902), .dinb(n432), .dout(n29054));
  jnot g11032(.din(n29054), .dout(n29055));
  jor  g11033(.dina(n29055), .dinb(n29053), .dout(n29056));
  jand g11034(.dina(n29056), .dinb(n28904), .dout(n29057));
  jxor g11035(.dina(n28896), .dinb(n433), .dout(n29058));
  jnot g11036(.din(n29058), .dout(n29059));
  jor  g11037(.dina(n29059), .dinb(n29057), .dout(n29060));
  jand g11038(.dina(n29060), .dinb(n28898), .dout(n29061));
  jxor g11039(.dina(n28890), .dinb(n421), .dout(n29062));
  jnot g11040(.din(n29062), .dout(n29063));
  jor  g11041(.dina(n29063), .dinb(n29061), .dout(n29064));
  jand g11042(.dina(n29064), .dinb(n28892), .dout(n29065));
  jxor g11043(.dina(n28884), .dinb(n422), .dout(n29066));
  jnot g11044(.din(n29066), .dout(n29067));
  jor  g11045(.dina(n29067), .dinb(n29065), .dout(n29068));
  jand g11046(.dina(n29068), .dinb(n28886), .dout(n29069));
  jxor g11047(.dina(n28878), .dinb(n416), .dout(n29070));
  jnot g11048(.din(n29070), .dout(n29071));
  jor  g11049(.dina(n29071), .dinb(n29069), .dout(n29072));
  jand g11050(.dina(n29072), .dinb(n28880), .dout(n29073));
  jxor g11051(.dina(n28872), .dinb(n417), .dout(n29074));
  jnot g11052(.din(n29074), .dout(n29075));
  jor  g11053(.dina(n29075), .dinb(n29073), .dout(n29076));
  jand g11054(.dina(n29076), .dinb(n28874), .dout(n29077));
  jxor g11055(.dina(n28866), .dinb(n2547), .dout(n29078));
  jnot g11056(.din(n29078), .dout(n29079));
  jor  g11057(.dina(n29079), .dinb(n29077), .dout(n29080));
  jand g11058(.dina(n29080), .dinb(n28868), .dout(n29081));
  jxor g11059(.dina(n28860), .dinb(n2714), .dout(n29082));
  jnot g11060(.din(n29082), .dout(n29083));
  jor  g11061(.dina(n29083), .dinb(n29081), .dout(n29084));
  jand g11062(.dina(n29084), .dinb(n28862), .dout(n29085));
  jxor g11063(.dina(n28854), .dinb(n405), .dout(n29086));
  jnot g11064(.din(n29086), .dout(n29087));
  jor  g11065(.dina(n29087), .dinb(n29085), .dout(n29088));
  jand g11066(.dina(n29088), .dinb(n28856), .dout(n29089));
  jxor g11067(.dina(n28848), .dinb(n406), .dout(n29090));
  jnot g11068(.din(n29090), .dout(n29091));
  jor  g11069(.dina(n29091), .dinb(n29089), .dout(n29092));
  jand g11070(.dina(n29092), .dinb(n28850), .dout(n29093));
  jxor g11071(.dina(n28842), .dinb(n412), .dout(n29094));
  jnot g11072(.din(n29094), .dout(n29095));
  jor  g11073(.dina(n29095), .dinb(n29093), .dout(n29096));
  jand g11074(.dina(n29096), .dinb(n28844), .dout(n29097));
  jxor g11075(.dina(n28836), .dinb(n413), .dout(n29098));
  jnot g11076(.din(n29098), .dout(n29099));
  jor  g11077(.dina(n29099), .dinb(n29097), .dout(n29100));
  jand g11078(.dina(n29100), .dinb(n28838), .dout(n29101));
  jxor g11079(.dina(n28830), .dinb(n409), .dout(n29102));
  jnot g11080(.din(n29102), .dout(n29103));
  jor  g11081(.dina(n29103), .dinb(n29101), .dout(n29104));
  jand g11082(.dina(n29104), .dinb(n28832), .dout(n29105));
  jxor g11083(.dina(n28824), .dinb(n410), .dout(n29106));
  jnot g11084(.din(n29106), .dout(n29107));
  jor  g11085(.dina(n29107), .dinb(n29105), .dout(n29108));
  jand g11086(.dina(n29108), .dinb(n28826), .dout(n29109));
  jxor g11087(.dina(n28818), .dinb(n426), .dout(n29110));
  jnot g11088(.din(n29110), .dout(n29111));
  jor  g11089(.dina(n29111), .dinb(n29109), .dout(n29112));
  jand g11090(.dina(n29112), .dinb(n28820), .dout(n29113));
  jxor g11091(.dina(n28812), .dinb(n427), .dout(n29114));
  jnot g11092(.din(n29114), .dout(n29115));
  jor  g11093(.dina(n29115), .dinb(n29113), .dout(n29116));
  jand g11094(.dina(n29116), .dinb(n28814), .dout(n29117));
  jxor g11095(.dina(n28806), .dinb(n424), .dout(n29118));
  jnot g11096(.din(n29118), .dout(n29119));
  jor  g11097(.dina(n29119), .dinb(n29117), .dout(n29120));
  jand g11098(.dina(n29120), .dinb(n28808), .dout(n29121));
  jxor g11099(.dina(n28800), .dinb(n300), .dout(n29122));
  jnot g11100(.din(n29122), .dout(n29123));
  jor  g11101(.dina(n29123), .dinb(n29121), .dout(n29124));
  jand g11102(.dina(n29124), .dinb(n28802), .dout(n29125));
  jxor g11103(.dina(n28794), .dinb(n297), .dout(n29126));
  jnot g11104(.din(n29126), .dout(n29127));
  jor  g11105(.dina(n29127), .dinb(n29125), .dout(n29128));
  jand g11106(.dina(n29128), .dinb(n28796), .dout(n29129));
  jxor g11107(.dina(n28788), .dinb(n298), .dout(n29130));
  jnot g11108(.din(n29130), .dout(n29131));
  jor  g11109(.dina(n29131), .dinb(n29129), .dout(n29132));
  jand g11110(.dina(n29132), .dinb(n28790), .dout(n29133));
  jxor g11111(.dina(n28782), .dinb(n301), .dout(n29134));
  jnot g11112(.din(n29134), .dout(n29135));
  jor  g11113(.dina(n29135), .dinb(n29133), .dout(n29136));
  jand g11114(.dina(n29136), .dinb(n28784), .dout(n29137));
  jxor g11115(.dina(n28776), .dinb(n293), .dout(n29138));
  jnot g11116(.din(n29138), .dout(n29139));
  jor  g11117(.dina(n29139), .dinb(n29137), .dout(n29140));
  jand g11118(.dina(n29140), .dinb(n28778), .dout(n29141));
  jxor g11119(.dina(n28770), .dinb(n294), .dout(n29142));
  jnot g11120(.din(n29142), .dout(n29143));
  jor  g11121(.dina(n29143), .dinb(n29141), .dout(n29144));
  jand g11122(.dina(n29144), .dinb(n28772), .dout(n29145));
  jxor g11123(.dina(n28764), .dinb(n290), .dout(n29146));
  jnot g11124(.din(n29146), .dout(n29147));
  jor  g11125(.dina(n29147), .dinb(n29145), .dout(n29148));
  jand g11126(.dina(n29148), .dinb(n28766), .dout(n29149));
  jxor g11127(.dina(n28758), .dinb(n291), .dout(n29150));
  jnot g11128(.din(n29150), .dout(n29151));
  jor  g11129(.dina(n29151), .dinb(n29149), .dout(n29152));
  jand g11130(.dina(n29152), .dinb(n28760), .dout(n29153));
  jxor g11131(.dina(n28752), .dinb(n284), .dout(n29154));
  jnot g11132(.din(n29154), .dout(n29155));
  jor  g11133(.dina(n29155), .dinb(n29153), .dout(n29156));
  jand g11134(.dina(n29156), .dinb(n28754), .dout(n29157));
  jnot g11135(.din(n8458), .dout(n29158));
  jxor g11136(.dina(n28743), .dinb(b41 ), .dout(n29159));
  jor  g11137(.dina(n29159), .dinb(n29158), .dout(n29160));
  jor  g11138(.dina(n29160), .dinb(n29157), .dout(n29161));
  jand g11139(.dina(n29161), .dinb(n28744), .dout(n29162));
  jxor g11140(.dina(n28998), .dinb(b1 ), .dout(n29163));
  jand g11141(.dina(n29163), .dinb(n8669), .dout(n29164));
  jor  g11142(.dina(n29164), .dinb(n28993), .dout(n29165));
  jand g11143(.dina(n29002), .dinb(n29165), .dout(n29166));
  jor  g11144(.dina(n29166), .dinb(n28986), .dout(n29167));
  jand g11145(.dina(n29006), .dinb(n29167), .dout(n29168));
  jor  g11146(.dina(n29168), .dinb(n28980), .dout(n29169));
  jand g11147(.dina(n29010), .dinb(n29169), .dout(n29170));
  jor  g11148(.dina(n29170), .dinb(n28971), .dout(n29171));
  jand g11149(.dina(n29014), .dinb(n29171), .dout(n29172));
  jor  g11150(.dina(n29172), .dinb(n28963), .dout(n29173));
  jand g11151(.dina(n29018), .dinb(n29173), .dout(n29174));
  jor  g11152(.dina(n29174), .dinb(n28957), .dout(n29175));
  jand g11153(.dina(n29022), .dinb(n29175), .dout(n29176));
  jor  g11154(.dina(n29176), .dinb(n28951), .dout(n29177));
  jand g11155(.dina(n29026), .dinb(n29177), .dout(n29178));
  jor  g11156(.dina(n29178), .dinb(n28945), .dout(n29179));
  jand g11157(.dina(n29030), .dinb(n29179), .dout(n29180));
  jor  g11158(.dina(n29180), .dinb(n28939), .dout(n29181));
  jand g11159(.dina(n29034), .dinb(n29181), .dout(n29182));
  jor  g11160(.dina(n29182), .dinb(n28933), .dout(n29183));
  jand g11161(.dina(n29038), .dinb(n29183), .dout(n29184));
  jor  g11162(.dina(n29184), .dinb(n28927), .dout(n29185));
  jand g11163(.dina(n29042), .dinb(n29185), .dout(n29186));
  jor  g11164(.dina(n29186), .dinb(n28921), .dout(n29187));
  jand g11165(.dina(n29046), .dinb(n29187), .dout(n29188));
  jor  g11166(.dina(n29188), .dinb(n28915), .dout(n29189));
  jand g11167(.dina(n29050), .dinb(n29189), .dout(n29190));
  jor  g11168(.dina(n29190), .dinb(n28909), .dout(n29191));
  jand g11169(.dina(n29054), .dinb(n29191), .dout(n29192));
  jor  g11170(.dina(n29192), .dinb(n28903), .dout(n29193));
  jand g11171(.dina(n29058), .dinb(n29193), .dout(n29194));
  jor  g11172(.dina(n29194), .dinb(n28897), .dout(n29195));
  jand g11173(.dina(n29062), .dinb(n29195), .dout(n29196));
  jor  g11174(.dina(n29196), .dinb(n28891), .dout(n29197));
  jand g11175(.dina(n29066), .dinb(n29197), .dout(n29198));
  jor  g11176(.dina(n29198), .dinb(n28885), .dout(n29199));
  jand g11177(.dina(n29070), .dinb(n29199), .dout(n29200));
  jor  g11178(.dina(n29200), .dinb(n28879), .dout(n29201));
  jand g11179(.dina(n29074), .dinb(n29201), .dout(n29202));
  jor  g11180(.dina(n29202), .dinb(n28873), .dout(n29203));
  jand g11181(.dina(n29078), .dinb(n29203), .dout(n29204));
  jor  g11182(.dina(n29204), .dinb(n28867), .dout(n29205));
  jand g11183(.dina(n29082), .dinb(n29205), .dout(n29206));
  jor  g11184(.dina(n29206), .dinb(n28861), .dout(n29207));
  jand g11185(.dina(n29086), .dinb(n29207), .dout(n29208));
  jor  g11186(.dina(n29208), .dinb(n28855), .dout(n29209));
  jand g11187(.dina(n29090), .dinb(n29209), .dout(n29210));
  jor  g11188(.dina(n29210), .dinb(n28849), .dout(n29211));
  jand g11189(.dina(n29094), .dinb(n29211), .dout(n29212));
  jor  g11190(.dina(n29212), .dinb(n28843), .dout(n29213));
  jand g11191(.dina(n29098), .dinb(n29213), .dout(n29214));
  jor  g11192(.dina(n29214), .dinb(n28837), .dout(n29215));
  jand g11193(.dina(n29102), .dinb(n29215), .dout(n29216));
  jor  g11194(.dina(n29216), .dinb(n28831), .dout(n29217));
  jand g11195(.dina(n29106), .dinb(n29217), .dout(n29218));
  jor  g11196(.dina(n29218), .dinb(n28825), .dout(n29219));
  jand g11197(.dina(n29110), .dinb(n29219), .dout(n29220));
  jor  g11198(.dina(n29220), .dinb(n28819), .dout(n29221));
  jand g11199(.dina(n29114), .dinb(n29221), .dout(n29222));
  jor  g11200(.dina(n29222), .dinb(n28813), .dout(n29223));
  jand g11201(.dina(n29118), .dinb(n29223), .dout(n29224));
  jor  g11202(.dina(n29224), .dinb(n28807), .dout(n29225));
  jand g11203(.dina(n29122), .dinb(n29225), .dout(n29226));
  jor  g11204(.dina(n29226), .dinb(n28801), .dout(n29227));
  jand g11205(.dina(n29126), .dinb(n29227), .dout(n29228));
  jor  g11206(.dina(n29228), .dinb(n28795), .dout(n29229));
  jand g11207(.dina(n29130), .dinb(n29229), .dout(n29230));
  jor  g11208(.dina(n29230), .dinb(n28789), .dout(n29231));
  jand g11209(.dina(n29134), .dinb(n29231), .dout(n29232));
  jor  g11210(.dina(n29232), .dinb(n28783), .dout(n29233));
  jand g11211(.dina(n29138), .dinb(n29233), .dout(n29234));
  jor  g11212(.dina(n29234), .dinb(n28777), .dout(n29235));
  jand g11213(.dina(n29142), .dinb(n29235), .dout(n29236));
  jor  g11214(.dina(n29236), .dinb(n28771), .dout(n29237));
  jand g11215(.dina(n29146), .dinb(n29237), .dout(n29238));
  jor  g11216(.dina(n29238), .dinb(n28765), .dout(n29239));
  jand g11217(.dina(n29150), .dinb(n29239), .dout(n29240));
  jor  g11218(.dina(n29240), .dinb(n28759), .dout(n29241));
  jand g11219(.dina(n29154), .dinb(n29241), .dout(n29242));
  jor  g11220(.dina(n29242), .dinb(n28753), .dout(n29243));
  jnot g11221(.din(n29160), .dout(n29244));
  jand g11222(.dina(n29244), .dinb(n29243), .dout(n29245));
  jand g11223(.dina(n28743), .dinb(n518), .dout(n29246));
  jor  g11224(.dina(n29246), .dinb(n29245), .dout(n29247));
  jxor g11225(.dina(n29159), .dinb(n29243), .dout(n29248));
  jand g11226(.dina(n29248), .dinb(n29247), .dout(n29249));
  jor  g11227(.dina(n29249), .dinb(n29162), .dout(n29250));
  jnot g11228(.din(n29250), .dout(n29251));
  jand g11229(.dina(n29250), .dinb(b42 ), .dout(n29252));
  jnot g11230(.din(n29252), .dout(n29253));
  jand g11231(.dina(n29251), .dinb(n281), .dout(n29254));
  jnot g11232(.din(n29246), .dout(n29255));
  jand g11233(.dina(n29255), .dinb(n29161), .dout(n29256));
  jand g11234(.dina(n29256), .dinb(n28752), .dout(n29257));
  jxor g11235(.dina(n29154), .dinb(n29241), .dout(n29258));
  jand g11236(.dina(n29258), .dinb(n29247), .dout(n29259));
  jor  g11237(.dina(n29259), .dinb(n29257), .dout(n29260));
  jand g11238(.dina(n29260), .dinb(n285), .dout(n29261));
  jand g11239(.dina(n29256), .dinb(n28758), .dout(n29262));
  jxor g11240(.dina(n29150), .dinb(n29239), .dout(n29263));
  jand g11241(.dina(n29263), .dinb(n29247), .dout(n29264));
  jor  g11242(.dina(n29264), .dinb(n29262), .dout(n29265));
  jand g11243(.dina(n29265), .dinb(n284), .dout(n29266));
  jand g11244(.dina(n29256), .dinb(n28764), .dout(n29267));
  jxor g11245(.dina(n29146), .dinb(n29237), .dout(n29268));
  jand g11246(.dina(n29268), .dinb(n29247), .dout(n29269));
  jor  g11247(.dina(n29269), .dinb(n29267), .dout(n29270));
  jand g11248(.dina(n29270), .dinb(n291), .dout(n29271));
  jand g11249(.dina(n29256), .dinb(n28770), .dout(n29272));
  jxor g11250(.dina(n29142), .dinb(n29235), .dout(n29273));
  jand g11251(.dina(n29273), .dinb(n29247), .dout(n29274));
  jor  g11252(.dina(n29274), .dinb(n29272), .dout(n29275));
  jand g11253(.dina(n29275), .dinb(n290), .dout(n29276));
  jand g11254(.dina(n29256), .dinb(n28776), .dout(n29277));
  jxor g11255(.dina(n29138), .dinb(n29233), .dout(n29278));
  jand g11256(.dina(n29278), .dinb(n29247), .dout(n29279));
  jor  g11257(.dina(n29279), .dinb(n29277), .dout(n29280));
  jand g11258(.dina(n29280), .dinb(n294), .dout(n29281));
  jand g11259(.dina(n29256), .dinb(n28782), .dout(n29282));
  jxor g11260(.dina(n29134), .dinb(n29231), .dout(n29283));
  jand g11261(.dina(n29283), .dinb(n29247), .dout(n29284));
  jor  g11262(.dina(n29284), .dinb(n29282), .dout(n29285));
  jand g11263(.dina(n29285), .dinb(n293), .dout(n29286));
  jand g11264(.dina(n29256), .dinb(n28788), .dout(n29287));
  jxor g11265(.dina(n29130), .dinb(n29229), .dout(n29288));
  jand g11266(.dina(n29288), .dinb(n29247), .dout(n29289));
  jor  g11267(.dina(n29289), .dinb(n29287), .dout(n29290));
  jand g11268(.dina(n29290), .dinb(n301), .dout(n29291));
  jand g11269(.dina(n29256), .dinb(n28794), .dout(n29292));
  jxor g11270(.dina(n29126), .dinb(n29227), .dout(n29293));
  jand g11271(.dina(n29293), .dinb(n29247), .dout(n29294));
  jor  g11272(.dina(n29294), .dinb(n29292), .dout(n29295));
  jand g11273(.dina(n29295), .dinb(n298), .dout(n29296));
  jand g11274(.dina(n29256), .dinb(n28800), .dout(n29297));
  jxor g11275(.dina(n29122), .dinb(n29225), .dout(n29298));
  jand g11276(.dina(n29298), .dinb(n29247), .dout(n29299));
  jor  g11277(.dina(n29299), .dinb(n29297), .dout(n29300));
  jand g11278(.dina(n29300), .dinb(n297), .dout(n29301));
  jand g11279(.dina(n29256), .dinb(n28806), .dout(n29302));
  jxor g11280(.dina(n29118), .dinb(n29223), .dout(n29303));
  jand g11281(.dina(n29303), .dinb(n29247), .dout(n29304));
  jor  g11282(.dina(n29304), .dinb(n29302), .dout(n29305));
  jand g11283(.dina(n29305), .dinb(n300), .dout(n29306));
  jand g11284(.dina(n29256), .dinb(n28812), .dout(n29307));
  jxor g11285(.dina(n29114), .dinb(n29221), .dout(n29308));
  jand g11286(.dina(n29308), .dinb(n29247), .dout(n29309));
  jor  g11287(.dina(n29309), .dinb(n29307), .dout(n29310));
  jand g11288(.dina(n29310), .dinb(n424), .dout(n29311));
  jand g11289(.dina(n29256), .dinb(n28818), .dout(n29312));
  jxor g11290(.dina(n29110), .dinb(n29219), .dout(n29313));
  jand g11291(.dina(n29313), .dinb(n29247), .dout(n29314));
  jor  g11292(.dina(n29314), .dinb(n29312), .dout(n29315));
  jand g11293(.dina(n29315), .dinb(n427), .dout(n29316));
  jand g11294(.dina(n29256), .dinb(n28824), .dout(n29317));
  jxor g11295(.dina(n29106), .dinb(n29217), .dout(n29318));
  jand g11296(.dina(n29318), .dinb(n29247), .dout(n29319));
  jor  g11297(.dina(n29319), .dinb(n29317), .dout(n29320));
  jand g11298(.dina(n29320), .dinb(n426), .dout(n29321));
  jand g11299(.dina(n29256), .dinb(n28830), .dout(n29322));
  jxor g11300(.dina(n29102), .dinb(n29215), .dout(n29323));
  jand g11301(.dina(n29323), .dinb(n29247), .dout(n29324));
  jor  g11302(.dina(n29324), .dinb(n29322), .dout(n29325));
  jand g11303(.dina(n29325), .dinb(n410), .dout(n29326));
  jand g11304(.dina(n29256), .dinb(n28836), .dout(n29327));
  jxor g11305(.dina(n29098), .dinb(n29213), .dout(n29328));
  jand g11306(.dina(n29328), .dinb(n29247), .dout(n29329));
  jor  g11307(.dina(n29329), .dinb(n29327), .dout(n29330));
  jand g11308(.dina(n29330), .dinb(n409), .dout(n29331));
  jand g11309(.dina(n29256), .dinb(n28842), .dout(n29332));
  jxor g11310(.dina(n29094), .dinb(n29211), .dout(n29333));
  jand g11311(.dina(n29333), .dinb(n29247), .dout(n29334));
  jor  g11312(.dina(n29334), .dinb(n29332), .dout(n29335));
  jand g11313(.dina(n29335), .dinb(n413), .dout(n29336));
  jand g11314(.dina(n29256), .dinb(n28848), .dout(n29337));
  jxor g11315(.dina(n29090), .dinb(n29209), .dout(n29338));
  jand g11316(.dina(n29338), .dinb(n29247), .dout(n29339));
  jor  g11317(.dina(n29339), .dinb(n29337), .dout(n29340));
  jand g11318(.dina(n29340), .dinb(n412), .dout(n29341));
  jand g11319(.dina(n29256), .dinb(n28854), .dout(n29342));
  jxor g11320(.dina(n29086), .dinb(n29207), .dout(n29343));
  jand g11321(.dina(n29343), .dinb(n29247), .dout(n29344));
  jor  g11322(.dina(n29344), .dinb(n29342), .dout(n29345));
  jand g11323(.dina(n29345), .dinb(n406), .dout(n29346));
  jand g11324(.dina(n29256), .dinb(n28860), .dout(n29347));
  jxor g11325(.dina(n29082), .dinb(n29205), .dout(n29348));
  jand g11326(.dina(n29348), .dinb(n29247), .dout(n29349));
  jor  g11327(.dina(n29349), .dinb(n29347), .dout(n29350));
  jand g11328(.dina(n29350), .dinb(n405), .dout(n29351));
  jand g11329(.dina(n29256), .dinb(n28866), .dout(n29352));
  jxor g11330(.dina(n29078), .dinb(n29203), .dout(n29353));
  jand g11331(.dina(n29353), .dinb(n29247), .dout(n29354));
  jor  g11332(.dina(n29354), .dinb(n29352), .dout(n29355));
  jand g11333(.dina(n29355), .dinb(n2714), .dout(n29356));
  jand g11334(.dina(n29256), .dinb(n28872), .dout(n29357));
  jxor g11335(.dina(n29074), .dinb(n29201), .dout(n29358));
  jand g11336(.dina(n29358), .dinb(n29247), .dout(n29359));
  jor  g11337(.dina(n29359), .dinb(n29357), .dout(n29360));
  jand g11338(.dina(n29360), .dinb(n2547), .dout(n29361));
  jand g11339(.dina(n29256), .dinb(n28878), .dout(n29362));
  jxor g11340(.dina(n29070), .dinb(n29199), .dout(n29363));
  jand g11341(.dina(n29363), .dinb(n29247), .dout(n29364));
  jor  g11342(.dina(n29364), .dinb(n29362), .dout(n29365));
  jand g11343(.dina(n29365), .dinb(n417), .dout(n29366));
  jand g11344(.dina(n29256), .dinb(n28884), .dout(n29367));
  jxor g11345(.dina(n29066), .dinb(n29197), .dout(n29368));
  jand g11346(.dina(n29368), .dinb(n29247), .dout(n29369));
  jor  g11347(.dina(n29369), .dinb(n29367), .dout(n29370));
  jand g11348(.dina(n29370), .dinb(n416), .dout(n29371));
  jand g11349(.dina(n29256), .dinb(n28890), .dout(n29372));
  jxor g11350(.dina(n29062), .dinb(n29195), .dout(n29373));
  jand g11351(.dina(n29373), .dinb(n29247), .dout(n29374));
  jor  g11352(.dina(n29374), .dinb(n29372), .dout(n29375));
  jand g11353(.dina(n29375), .dinb(n422), .dout(n29376));
  jand g11354(.dina(n29256), .dinb(n28896), .dout(n29377));
  jxor g11355(.dina(n29058), .dinb(n29193), .dout(n29378));
  jand g11356(.dina(n29378), .dinb(n29247), .dout(n29379));
  jor  g11357(.dina(n29379), .dinb(n29377), .dout(n29380));
  jand g11358(.dina(n29380), .dinb(n421), .dout(n29381));
  jand g11359(.dina(n29256), .dinb(n28902), .dout(n29382));
  jxor g11360(.dina(n29054), .dinb(n29191), .dout(n29383));
  jand g11361(.dina(n29383), .dinb(n29247), .dout(n29384));
  jor  g11362(.dina(n29384), .dinb(n29382), .dout(n29385));
  jand g11363(.dina(n29385), .dinb(n433), .dout(n29386));
  jand g11364(.dina(n29256), .dinb(n28908), .dout(n29387));
  jxor g11365(.dina(n29050), .dinb(n29189), .dout(n29388));
  jand g11366(.dina(n29388), .dinb(n29247), .dout(n29389));
  jor  g11367(.dina(n29389), .dinb(n29387), .dout(n29390));
  jand g11368(.dina(n29390), .dinb(n432), .dout(n29391));
  jand g11369(.dina(n29256), .dinb(n28914), .dout(n29392));
  jxor g11370(.dina(n29046), .dinb(n29187), .dout(n29393));
  jand g11371(.dina(n29393), .dinb(n29247), .dout(n29394));
  jor  g11372(.dina(n29394), .dinb(n29392), .dout(n29395));
  jand g11373(.dina(n29395), .dinb(n436), .dout(n29396));
  jand g11374(.dina(n29256), .dinb(n28920), .dout(n29397));
  jxor g11375(.dina(n29042), .dinb(n29185), .dout(n29398));
  jand g11376(.dina(n29398), .dinb(n29247), .dout(n29399));
  jor  g11377(.dina(n29399), .dinb(n29397), .dout(n29400));
  jand g11378(.dina(n29400), .dinb(n435), .dout(n29401));
  jand g11379(.dina(n29256), .dinb(n28926), .dout(n29402));
  jxor g11380(.dina(n29038), .dinb(n29183), .dout(n29403));
  jand g11381(.dina(n29403), .dinb(n29247), .dout(n29404));
  jor  g11382(.dina(n29404), .dinb(n29402), .dout(n29405));
  jand g11383(.dina(n29405), .dinb(n440), .dout(n29406));
  jand g11384(.dina(n29256), .dinb(n28932), .dout(n29407));
  jxor g11385(.dina(n29034), .dinb(n29181), .dout(n29408));
  jand g11386(.dina(n29408), .dinb(n29247), .dout(n29409));
  jor  g11387(.dina(n29409), .dinb(n29407), .dout(n29410));
  jand g11388(.dina(n29410), .dinb(n439), .dout(n29411));
  jand g11389(.dina(n29256), .dinb(n28938), .dout(n29412));
  jxor g11390(.dina(n29030), .dinb(n29179), .dout(n29413));
  jand g11391(.dina(n29413), .dinb(n29247), .dout(n29414));
  jor  g11392(.dina(n29414), .dinb(n29412), .dout(n29415));
  jand g11393(.dina(n29415), .dinb(n325), .dout(n29416));
  jand g11394(.dina(n29256), .dinb(n28944), .dout(n29417));
  jxor g11395(.dina(n29026), .dinb(n29177), .dout(n29418));
  jand g11396(.dina(n29418), .dinb(n29247), .dout(n29419));
  jor  g11397(.dina(n29419), .dinb(n29417), .dout(n29420));
  jand g11398(.dina(n29420), .dinb(n324), .dout(n29421));
  jand g11399(.dina(n29256), .dinb(n28950), .dout(n29422));
  jxor g11400(.dina(n29022), .dinb(n29175), .dout(n29423));
  jand g11401(.dina(n29423), .dinb(n29247), .dout(n29424));
  jor  g11402(.dina(n29424), .dinb(n29422), .dout(n29425));
  jand g11403(.dina(n29425), .dinb(n323), .dout(n29426));
  jand g11404(.dina(n29256), .dinb(n28956), .dout(n29427));
  jxor g11405(.dina(n29018), .dinb(n29173), .dout(n29428));
  jand g11406(.dina(n29428), .dinb(n29247), .dout(n29429));
  jor  g11407(.dina(n29429), .dinb(n29427), .dout(n29430));
  jand g11408(.dina(n29430), .dinb(n335), .dout(n29431));
  jand g11409(.dina(n29256), .dinb(n28962), .dout(n29432));
  jxor g11410(.dina(n29014), .dinb(n29171), .dout(n29433));
  jand g11411(.dina(n29433), .dinb(n29247), .dout(n29434));
  jor  g11412(.dina(n29434), .dinb(n29432), .dout(n29435));
  jand g11413(.dina(n29435), .dinb(n334), .dout(n29436));
  jand g11414(.dina(n29256), .dinb(n28970), .dout(n29437));
  jxor g11415(.dina(n29010), .dinb(n29169), .dout(n29438));
  jand g11416(.dina(n29438), .dinb(n29247), .dout(n29439));
  jor  g11417(.dina(n29439), .dinb(n29437), .dout(n29440));
  jand g11418(.dina(n29440), .dinb(n338), .dout(n29441));
  jand g11419(.dina(n29256), .dinb(n28979), .dout(n29442));
  jxor g11420(.dina(n29006), .dinb(n29167), .dout(n29443));
  jand g11421(.dina(n29443), .dinb(n29247), .dout(n29444));
  jor  g11422(.dina(n29444), .dinb(n29442), .dout(n29445));
  jand g11423(.dina(n29445), .dinb(n337), .dout(n29446));
  jand g11424(.dina(n29256), .dinb(n28985), .dout(n29447));
  jxor g11425(.dina(n29002), .dinb(n29165), .dout(n29448));
  jand g11426(.dina(n29448), .dinb(n29247), .dout(n29449));
  jor  g11427(.dina(n29449), .dinb(n29447), .dout(n29450));
  jand g11428(.dina(n29450), .dinb(n344), .dout(n29451));
  jand g11429(.dina(n29256), .dinb(n28992), .dout(n29452));
  jxor g11430(.dina(n29163), .dinb(n8669), .dout(n29453));
  jand g11431(.dina(n29453), .dinb(n29247), .dout(n29454));
  jor  g11432(.dina(n29454), .dinb(n29452), .dout(n29455));
  jand g11433(.dina(n29455), .dinb(n348), .dout(n29456));
  jor  g11434(.dina(n29256), .dinb(n18364), .dout(n29457));
  jand g11435(.dina(n29457), .dinb(a22 ), .dout(n29458));
  jor  g11436(.dina(n29256), .dinb(n8669), .dout(n29459));
  jnot g11437(.din(n29459), .dout(n29460));
  jor  g11438(.dina(n29460), .dinb(n29458), .dout(n29461));
  jand g11439(.dina(n29461), .dinb(n258), .dout(n29462));
  jand g11440(.dina(n29247), .dinb(b0 ), .dout(n29463));
  jor  g11441(.dina(n29463), .dinb(n8667), .dout(n29464));
  jand g11442(.dina(n29459), .dinb(n29464), .dout(n29465));
  jxor g11443(.dina(n29465), .dinb(b1 ), .dout(n29466));
  jand g11444(.dina(n29466), .dinb(n9017), .dout(n29467));
  jor  g11445(.dina(n29467), .dinb(n29462), .dout(n29468));
  jxor g11446(.dina(n29455), .dinb(n348), .dout(n29469));
  jand g11447(.dina(n29469), .dinb(n29468), .dout(n29470));
  jor  g11448(.dina(n29470), .dinb(n29456), .dout(n29471));
  jxor g11449(.dina(n29450), .dinb(n344), .dout(n29472));
  jand g11450(.dina(n29472), .dinb(n29471), .dout(n29473));
  jor  g11451(.dina(n29473), .dinb(n29451), .dout(n29474));
  jxor g11452(.dina(n29445), .dinb(n337), .dout(n29475));
  jand g11453(.dina(n29475), .dinb(n29474), .dout(n29476));
  jor  g11454(.dina(n29476), .dinb(n29446), .dout(n29477));
  jxor g11455(.dina(n29440), .dinb(n338), .dout(n29478));
  jand g11456(.dina(n29478), .dinb(n29477), .dout(n29479));
  jor  g11457(.dina(n29479), .dinb(n29441), .dout(n29480));
  jxor g11458(.dina(n29435), .dinb(n334), .dout(n29481));
  jand g11459(.dina(n29481), .dinb(n29480), .dout(n29482));
  jor  g11460(.dina(n29482), .dinb(n29436), .dout(n29483));
  jxor g11461(.dina(n29430), .dinb(n335), .dout(n29484));
  jand g11462(.dina(n29484), .dinb(n29483), .dout(n29485));
  jor  g11463(.dina(n29485), .dinb(n29431), .dout(n29486));
  jxor g11464(.dina(n29425), .dinb(n323), .dout(n29487));
  jand g11465(.dina(n29487), .dinb(n29486), .dout(n29488));
  jor  g11466(.dina(n29488), .dinb(n29426), .dout(n29489));
  jxor g11467(.dina(n29420), .dinb(n324), .dout(n29490));
  jand g11468(.dina(n29490), .dinb(n29489), .dout(n29491));
  jor  g11469(.dina(n29491), .dinb(n29421), .dout(n29492));
  jxor g11470(.dina(n29415), .dinb(n325), .dout(n29493));
  jand g11471(.dina(n29493), .dinb(n29492), .dout(n29494));
  jor  g11472(.dina(n29494), .dinb(n29416), .dout(n29495));
  jxor g11473(.dina(n29410), .dinb(n439), .dout(n29496));
  jand g11474(.dina(n29496), .dinb(n29495), .dout(n29497));
  jor  g11475(.dina(n29497), .dinb(n29411), .dout(n29498));
  jxor g11476(.dina(n29405), .dinb(n440), .dout(n29499));
  jand g11477(.dina(n29499), .dinb(n29498), .dout(n29500));
  jor  g11478(.dina(n29500), .dinb(n29406), .dout(n29501));
  jxor g11479(.dina(n29400), .dinb(n435), .dout(n29502));
  jand g11480(.dina(n29502), .dinb(n29501), .dout(n29503));
  jor  g11481(.dina(n29503), .dinb(n29401), .dout(n29504));
  jxor g11482(.dina(n29395), .dinb(n436), .dout(n29505));
  jand g11483(.dina(n29505), .dinb(n29504), .dout(n29506));
  jor  g11484(.dina(n29506), .dinb(n29396), .dout(n29507));
  jxor g11485(.dina(n29390), .dinb(n432), .dout(n29508));
  jand g11486(.dina(n29508), .dinb(n29507), .dout(n29509));
  jor  g11487(.dina(n29509), .dinb(n29391), .dout(n29510));
  jxor g11488(.dina(n29385), .dinb(n433), .dout(n29511));
  jand g11489(.dina(n29511), .dinb(n29510), .dout(n29512));
  jor  g11490(.dina(n29512), .dinb(n29386), .dout(n29513));
  jxor g11491(.dina(n29380), .dinb(n421), .dout(n29514));
  jand g11492(.dina(n29514), .dinb(n29513), .dout(n29515));
  jor  g11493(.dina(n29515), .dinb(n29381), .dout(n29516));
  jxor g11494(.dina(n29375), .dinb(n422), .dout(n29517));
  jand g11495(.dina(n29517), .dinb(n29516), .dout(n29518));
  jor  g11496(.dina(n29518), .dinb(n29376), .dout(n29519));
  jxor g11497(.dina(n29370), .dinb(n416), .dout(n29520));
  jand g11498(.dina(n29520), .dinb(n29519), .dout(n29521));
  jor  g11499(.dina(n29521), .dinb(n29371), .dout(n29522));
  jxor g11500(.dina(n29365), .dinb(n417), .dout(n29523));
  jand g11501(.dina(n29523), .dinb(n29522), .dout(n29524));
  jor  g11502(.dina(n29524), .dinb(n29366), .dout(n29525));
  jxor g11503(.dina(n29360), .dinb(n2547), .dout(n29526));
  jand g11504(.dina(n29526), .dinb(n29525), .dout(n29527));
  jor  g11505(.dina(n29527), .dinb(n29361), .dout(n29528));
  jxor g11506(.dina(n29355), .dinb(n2714), .dout(n29529));
  jand g11507(.dina(n29529), .dinb(n29528), .dout(n29530));
  jor  g11508(.dina(n29530), .dinb(n29356), .dout(n29531));
  jxor g11509(.dina(n29350), .dinb(n405), .dout(n29532));
  jand g11510(.dina(n29532), .dinb(n29531), .dout(n29533));
  jor  g11511(.dina(n29533), .dinb(n29351), .dout(n29534));
  jxor g11512(.dina(n29345), .dinb(n406), .dout(n29535));
  jand g11513(.dina(n29535), .dinb(n29534), .dout(n29536));
  jor  g11514(.dina(n29536), .dinb(n29346), .dout(n29537));
  jxor g11515(.dina(n29340), .dinb(n412), .dout(n29538));
  jand g11516(.dina(n29538), .dinb(n29537), .dout(n29539));
  jor  g11517(.dina(n29539), .dinb(n29341), .dout(n29540));
  jxor g11518(.dina(n29335), .dinb(n413), .dout(n29541));
  jand g11519(.dina(n29541), .dinb(n29540), .dout(n29542));
  jor  g11520(.dina(n29542), .dinb(n29336), .dout(n29543));
  jxor g11521(.dina(n29330), .dinb(n409), .dout(n29544));
  jand g11522(.dina(n29544), .dinb(n29543), .dout(n29545));
  jor  g11523(.dina(n29545), .dinb(n29331), .dout(n29546));
  jxor g11524(.dina(n29325), .dinb(n410), .dout(n29547));
  jand g11525(.dina(n29547), .dinb(n29546), .dout(n29548));
  jor  g11526(.dina(n29548), .dinb(n29326), .dout(n29549));
  jxor g11527(.dina(n29320), .dinb(n426), .dout(n29550));
  jand g11528(.dina(n29550), .dinb(n29549), .dout(n29551));
  jor  g11529(.dina(n29551), .dinb(n29321), .dout(n29552));
  jxor g11530(.dina(n29315), .dinb(n427), .dout(n29553));
  jand g11531(.dina(n29553), .dinb(n29552), .dout(n29554));
  jor  g11532(.dina(n29554), .dinb(n29316), .dout(n29555));
  jxor g11533(.dina(n29310), .dinb(n424), .dout(n29556));
  jand g11534(.dina(n29556), .dinb(n29555), .dout(n29557));
  jor  g11535(.dina(n29557), .dinb(n29311), .dout(n29558));
  jxor g11536(.dina(n29305), .dinb(n300), .dout(n29559));
  jand g11537(.dina(n29559), .dinb(n29558), .dout(n29560));
  jor  g11538(.dina(n29560), .dinb(n29306), .dout(n29561));
  jxor g11539(.dina(n29300), .dinb(n297), .dout(n29562));
  jand g11540(.dina(n29562), .dinb(n29561), .dout(n29563));
  jor  g11541(.dina(n29563), .dinb(n29301), .dout(n29564));
  jxor g11542(.dina(n29295), .dinb(n298), .dout(n29565));
  jand g11543(.dina(n29565), .dinb(n29564), .dout(n29566));
  jor  g11544(.dina(n29566), .dinb(n29296), .dout(n29567));
  jxor g11545(.dina(n29290), .dinb(n301), .dout(n29568));
  jand g11546(.dina(n29568), .dinb(n29567), .dout(n29569));
  jor  g11547(.dina(n29569), .dinb(n29291), .dout(n29570));
  jxor g11548(.dina(n29285), .dinb(n293), .dout(n29571));
  jand g11549(.dina(n29571), .dinb(n29570), .dout(n29572));
  jor  g11550(.dina(n29572), .dinb(n29286), .dout(n29573));
  jxor g11551(.dina(n29280), .dinb(n294), .dout(n29574));
  jand g11552(.dina(n29574), .dinb(n29573), .dout(n29575));
  jor  g11553(.dina(n29575), .dinb(n29281), .dout(n29576));
  jxor g11554(.dina(n29275), .dinb(n290), .dout(n29577));
  jand g11555(.dina(n29577), .dinb(n29576), .dout(n29578));
  jor  g11556(.dina(n29578), .dinb(n29276), .dout(n29579));
  jxor g11557(.dina(n29270), .dinb(n291), .dout(n29580));
  jand g11558(.dina(n29580), .dinb(n29579), .dout(n29581));
  jor  g11559(.dina(n29581), .dinb(n29271), .dout(n29582));
  jxor g11560(.dina(n29265), .dinb(n284), .dout(n29583));
  jand g11561(.dina(n29583), .dinb(n29582), .dout(n29584));
  jor  g11562(.dina(n29584), .dinb(n29266), .dout(n29585));
  jxor g11563(.dina(n29260), .dinb(n285), .dout(n29586));
  jand g11564(.dina(n29586), .dinb(n29585), .dout(n29587));
  jor  g11565(.dina(n29587), .dinb(n29261), .dout(n29588));
  jor  g11566(.dina(n29588), .dinb(n29254), .dout(n29589));
  jand g11567(.dina(n29589), .dinb(n29253), .dout(n29590));
  jand g11568(.dina(n29590), .dinb(n517), .dout(n29591));
  jnot g11569(.din(n29591), .dout(n29592));
  jand g11570(.dina(n29592), .dinb(n29251), .dout(n29593));
  jand g11571(.dina(n29254), .dinb(n517), .dout(n29594));
  jand g11572(.dina(n29594), .dinb(n29588), .dout(n29595));
  jor  g11573(.dina(n29595), .dinb(n29593), .dout(n29596));
  jand g11574(.dina(n29596), .dinb(n517), .dout(n29597));
  jnot g11575(.din(n29597), .dout(n29598));
  jand g11576(.dina(n29592), .dinb(n29260), .dout(n29599));
  jxor g11577(.dina(n29586), .dinb(n29585), .dout(n29600));
  jand g11578(.dina(n29600), .dinb(n29591), .dout(n29601));
  jor  g11579(.dina(n29601), .dinb(n29599), .dout(n29602));
  jand g11580(.dina(n29602), .dinb(n281), .dout(n29603));
  jnot g11581(.din(n29603), .dout(n29604));
  jand g11582(.dina(n29592), .dinb(n29265), .dout(n29605));
  jxor g11583(.dina(n29583), .dinb(n29582), .dout(n29606));
  jand g11584(.dina(n29606), .dinb(n29591), .dout(n29607));
  jor  g11585(.dina(n29607), .dinb(n29605), .dout(n29608));
  jand g11586(.dina(n29608), .dinb(n285), .dout(n29609));
  jnot g11587(.din(n29609), .dout(n29610));
  jand g11588(.dina(n29592), .dinb(n29270), .dout(n29611));
  jxor g11589(.dina(n29580), .dinb(n29579), .dout(n29612));
  jand g11590(.dina(n29612), .dinb(n29591), .dout(n29613));
  jor  g11591(.dina(n29613), .dinb(n29611), .dout(n29614));
  jand g11592(.dina(n29614), .dinb(n284), .dout(n29615));
  jnot g11593(.din(n29615), .dout(n29616));
  jand g11594(.dina(n29592), .dinb(n29275), .dout(n29617));
  jxor g11595(.dina(n29577), .dinb(n29576), .dout(n29618));
  jand g11596(.dina(n29618), .dinb(n29591), .dout(n29619));
  jor  g11597(.dina(n29619), .dinb(n29617), .dout(n29620));
  jand g11598(.dina(n29620), .dinb(n291), .dout(n29621));
  jnot g11599(.din(n29621), .dout(n29622));
  jand g11600(.dina(n29592), .dinb(n29280), .dout(n29623));
  jxor g11601(.dina(n29574), .dinb(n29573), .dout(n29624));
  jand g11602(.dina(n29624), .dinb(n29591), .dout(n29625));
  jor  g11603(.dina(n29625), .dinb(n29623), .dout(n29626));
  jand g11604(.dina(n29626), .dinb(n290), .dout(n29627));
  jnot g11605(.din(n29627), .dout(n29628));
  jand g11606(.dina(n29592), .dinb(n29285), .dout(n29629));
  jxor g11607(.dina(n29571), .dinb(n29570), .dout(n29630));
  jand g11608(.dina(n29630), .dinb(n29591), .dout(n29631));
  jor  g11609(.dina(n29631), .dinb(n29629), .dout(n29632));
  jand g11610(.dina(n29632), .dinb(n294), .dout(n29633));
  jnot g11611(.din(n29633), .dout(n29634));
  jand g11612(.dina(n29592), .dinb(n29290), .dout(n29635));
  jxor g11613(.dina(n29568), .dinb(n29567), .dout(n29636));
  jand g11614(.dina(n29636), .dinb(n29591), .dout(n29637));
  jor  g11615(.dina(n29637), .dinb(n29635), .dout(n29638));
  jand g11616(.dina(n29638), .dinb(n293), .dout(n29639));
  jnot g11617(.din(n29639), .dout(n29640));
  jand g11618(.dina(n29592), .dinb(n29295), .dout(n29641));
  jxor g11619(.dina(n29565), .dinb(n29564), .dout(n29642));
  jand g11620(.dina(n29642), .dinb(n29591), .dout(n29643));
  jor  g11621(.dina(n29643), .dinb(n29641), .dout(n29644));
  jand g11622(.dina(n29644), .dinb(n301), .dout(n29645));
  jnot g11623(.din(n29645), .dout(n29646));
  jand g11624(.dina(n29592), .dinb(n29300), .dout(n29647));
  jxor g11625(.dina(n29562), .dinb(n29561), .dout(n29648));
  jand g11626(.dina(n29648), .dinb(n29591), .dout(n29649));
  jor  g11627(.dina(n29649), .dinb(n29647), .dout(n29650));
  jand g11628(.dina(n29650), .dinb(n298), .dout(n29651));
  jnot g11629(.din(n29651), .dout(n29652));
  jand g11630(.dina(n29592), .dinb(n29305), .dout(n29653));
  jxor g11631(.dina(n29559), .dinb(n29558), .dout(n29654));
  jand g11632(.dina(n29654), .dinb(n29591), .dout(n29655));
  jor  g11633(.dina(n29655), .dinb(n29653), .dout(n29656));
  jand g11634(.dina(n29656), .dinb(n297), .dout(n29657));
  jnot g11635(.din(n29657), .dout(n29658));
  jand g11636(.dina(n29592), .dinb(n29310), .dout(n29659));
  jxor g11637(.dina(n29556), .dinb(n29555), .dout(n29660));
  jand g11638(.dina(n29660), .dinb(n29591), .dout(n29661));
  jor  g11639(.dina(n29661), .dinb(n29659), .dout(n29662));
  jand g11640(.dina(n29662), .dinb(n300), .dout(n29663));
  jnot g11641(.din(n29663), .dout(n29664));
  jand g11642(.dina(n29592), .dinb(n29315), .dout(n29665));
  jxor g11643(.dina(n29553), .dinb(n29552), .dout(n29666));
  jand g11644(.dina(n29666), .dinb(n29591), .dout(n29667));
  jor  g11645(.dina(n29667), .dinb(n29665), .dout(n29668));
  jand g11646(.dina(n29668), .dinb(n424), .dout(n29669));
  jnot g11647(.din(n29669), .dout(n29670));
  jand g11648(.dina(n29592), .dinb(n29320), .dout(n29671));
  jxor g11649(.dina(n29550), .dinb(n29549), .dout(n29672));
  jand g11650(.dina(n29672), .dinb(n29591), .dout(n29673));
  jor  g11651(.dina(n29673), .dinb(n29671), .dout(n29674));
  jand g11652(.dina(n29674), .dinb(n427), .dout(n29675));
  jnot g11653(.din(n29675), .dout(n29676));
  jand g11654(.dina(n29592), .dinb(n29325), .dout(n29677));
  jxor g11655(.dina(n29547), .dinb(n29546), .dout(n29678));
  jand g11656(.dina(n29678), .dinb(n29591), .dout(n29679));
  jor  g11657(.dina(n29679), .dinb(n29677), .dout(n29680));
  jand g11658(.dina(n29680), .dinb(n426), .dout(n29681));
  jnot g11659(.din(n29681), .dout(n29682));
  jand g11660(.dina(n29592), .dinb(n29330), .dout(n29683));
  jxor g11661(.dina(n29544), .dinb(n29543), .dout(n29684));
  jand g11662(.dina(n29684), .dinb(n29591), .dout(n29685));
  jor  g11663(.dina(n29685), .dinb(n29683), .dout(n29686));
  jand g11664(.dina(n29686), .dinb(n410), .dout(n29687));
  jnot g11665(.din(n29687), .dout(n29688));
  jand g11666(.dina(n29592), .dinb(n29335), .dout(n29689));
  jxor g11667(.dina(n29541), .dinb(n29540), .dout(n29690));
  jand g11668(.dina(n29690), .dinb(n29591), .dout(n29691));
  jor  g11669(.dina(n29691), .dinb(n29689), .dout(n29692));
  jand g11670(.dina(n29692), .dinb(n409), .dout(n29693));
  jnot g11671(.din(n29693), .dout(n29694));
  jand g11672(.dina(n29592), .dinb(n29340), .dout(n29695));
  jxor g11673(.dina(n29538), .dinb(n29537), .dout(n29696));
  jand g11674(.dina(n29696), .dinb(n29591), .dout(n29697));
  jor  g11675(.dina(n29697), .dinb(n29695), .dout(n29698));
  jand g11676(.dina(n29698), .dinb(n413), .dout(n29699));
  jnot g11677(.din(n29699), .dout(n29700));
  jand g11678(.dina(n29592), .dinb(n29345), .dout(n29701));
  jxor g11679(.dina(n29535), .dinb(n29534), .dout(n29702));
  jand g11680(.dina(n29702), .dinb(n29591), .dout(n29703));
  jor  g11681(.dina(n29703), .dinb(n29701), .dout(n29704));
  jand g11682(.dina(n29704), .dinb(n412), .dout(n29705));
  jnot g11683(.din(n29705), .dout(n29706));
  jand g11684(.dina(n29592), .dinb(n29350), .dout(n29707));
  jxor g11685(.dina(n29532), .dinb(n29531), .dout(n29708));
  jand g11686(.dina(n29708), .dinb(n29591), .dout(n29709));
  jor  g11687(.dina(n29709), .dinb(n29707), .dout(n29710));
  jand g11688(.dina(n29710), .dinb(n406), .dout(n29711));
  jnot g11689(.din(n29711), .dout(n29712));
  jand g11690(.dina(n29592), .dinb(n29355), .dout(n29713));
  jxor g11691(.dina(n29529), .dinb(n29528), .dout(n29714));
  jand g11692(.dina(n29714), .dinb(n29591), .dout(n29715));
  jor  g11693(.dina(n29715), .dinb(n29713), .dout(n29716));
  jand g11694(.dina(n29716), .dinb(n405), .dout(n29717));
  jnot g11695(.din(n29717), .dout(n29718));
  jand g11696(.dina(n29592), .dinb(n29360), .dout(n29719));
  jxor g11697(.dina(n29526), .dinb(n29525), .dout(n29720));
  jand g11698(.dina(n29720), .dinb(n29591), .dout(n29721));
  jor  g11699(.dina(n29721), .dinb(n29719), .dout(n29722));
  jand g11700(.dina(n29722), .dinb(n2714), .dout(n29723));
  jnot g11701(.din(n29723), .dout(n29724));
  jand g11702(.dina(n29592), .dinb(n29365), .dout(n29725));
  jxor g11703(.dina(n29523), .dinb(n29522), .dout(n29726));
  jand g11704(.dina(n29726), .dinb(n29591), .dout(n29727));
  jor  g11705(.dina(n29727), .dinb(n29725), .dout(n29728));
  jand g11706(.dina(n29728), .dinb(n2547), .dout(n29729));
  jnot g11707(.din(n29729), .dout(n29730));
  jand g11708(.dina(n29592), .dinb(n29370), .dout(n29731));
  jxor g11709(.dina(n29520), .dinb(n29519), .dout(n29732));
  jand g11710(.dina(n29732), .dinb(n29591), .dout(n29733));
  jor  g11711(.dina(n29733), .dinb(n29731), .dout(n29734));
  jand g11712(.dina(n29734), .dinb(n417), .dout(n29735));
  jnot g11713(.din(n29735), .dout(n29736));
  jand g11714(.dina(n29592), .dinb(n29375), .dout(n29737));
  jxor g11715(.dina(n29517), .dinb(n29516), .dout(n29738));
  jand g11716(.dina(n29738), .dinb(n29591), .dout(n29739));
  jor  g11717(.dina(n29739), .dinb(n29737), .dout(n29740));
  jand g11718(.dina(n29740), .dinb(n416), .dout(n29741));
  jnot g11719(.din(n29741), .dout(n29742));
  jand g11720(.dina(n29592), .dinb(n29380), .dout(n29743));
  jxor g11721(.dina(n29514), .dinb(n29513), .dout(n29744));
  jand g11722(.dina(n29744), .dinb(n29591), .dout(n29745));
  jor  g11723(.dina(n29745), .dinb(n29743), .dout(n29746));
  jand g11724(.dina(n29746), .dinb(n422), .dout(n29747));
  jnot g11725(.din(n29747), .dout(n29748));
  jand g11726(.dina(n29592), .dinb(n29385), .dout(n29749));
  jxor g11727(.dina(n29511), .dinb(n29510), .dout(n29750));
  jand g11728(.dina(n29750), .dinb(n29591), .dout(n29751));
  jor  g11729(.dina(n29751), .dinb(n29749), .dout(n29752));
  jand g11730(.dina(n29752), .dinb(n421), .dout(n29753));
  jnot g11731(.din(n29753), .dout(n29754));
  jand g11732(.dina(n29592), .dinb(n29390), .dout(n29755));
  jxor g11733(.dina(n29508), .dinb(n29507), .dout(n29756));
  jand g11734(.dina(n29756), .dinb(n29591), .dout(n29757));
  jor  g11735(.dina(n29757), .dinb(n29755), .dout(n29758));
  jand g11736(.dina(n29758), .dinb(n433), .dout(n29759));
  jnot g11737(.din(n29759), .dout(n29760));
  jand g11738(.dina(n29592), .dinb(n29395), .dout(n29761));
  jxor g11739(.dina(n29505), .dinb(n29504), .dout(n29762));
  jand g11740(.dina(n29762), .dinb(n29591), .dout(n29763));
  jor  g11741(.dina(n29763), .dinb(n29761), .dout(n29764));
  jand g11742(.dina(n29764), .dinb(n432), .dout(n29765));
  jnot g11743(.din(n29765), .dout(n29766));
  jand g11744(.dina(n29592), .dinb(n29400), .dout(n29767));
  jxor g11745(.dina(n29502), .dinb(n29501), .dout(n29768));
  jand g11746(.dina(n29768), .dinb(n29591), .dout(n29769));
  jor  g11747(.dina(n29769), .dinb(n29767), .dout(n29770));
  jand g11748(.dina(n29770), .dinb(n436), .dout(n29771));
  jnot g11749(.din(n29771), .dout(n29772));
  jand g11750(.dina(n29592), .dinb(n29405), .dout(n29773));
  jxor g11751(.dina(n29499), .dinb(n29498), .dout(n29774));
  jand g11752(.dina(n29774), .dinb(n29591), .dout(n29775));
  jor  g11753(.dina(n29775), .dinb(n29773), .dout(n29776));
  jand g11754(.dina(n29776), .dinb(n435), .dout(n29777));
  jnot g11755(.din(n29777), .dout(n29778));
  jand g11756(.dina(n29592), .dinb(n29410), .dout(n29779));
  jxor g11757(.dina(n29496), .dinb(n29495), .dout(n29780));
  jand g11758(.dina(n29780), .dinb(n29591), .dout(n29781));
  jor  g11759(.dina(n29781), .dinb(n29779), .dout(n29782));
  jand g11760(.dina(n29782), .dinb(n440), .dout(n29783));
  jnot g11761(.din(n29783), .dout(n29784));
  jand g11762(.dina(n29592), .dinb(n29415), .dout(n29785));
  jxor g11763(.dina(n29493), .dinb(n29492), .dout(n29786));
  jand g11764(.dina(n29786), .dinb(n29591), .dout(n29787));
  jor  g11765(.dina(n29787), .dinb(n29785), .dout(n29788));
  jand g11766(.dina(n29788), .dinb(n439), .dout(n29789));
  jnot g11767(.din(n29789), .dout(n29790));
  jand g11768(.dina(n29592), .dinb(n29420), .dout(n29791));
  jxor g11769(.dina(n29490), .dinb(n29489), .dout(n29792));
  jand g11770(.dina(n29792), .dinb(n29591), .dout(n29793));
  jor  g11771(.dina(n29793), .dinb(n29791), .dout(n29794));
  jand g11772(.dina(n29794), .dinb(n325), .dout(n29795));
  jnot g11773(.din(n29795), .dout(n29796));
  jand g11774(.dina(n29592), .dinb(n29425), .dout(n29797));
  jxor g11775(.dina(n29487), .dinb(n29486), .dout(n29798));
  jand g11776(.dina(n29798), .dinb(n29591), .dout(n29799));
  jor  g11777(.dina(n29799), .dinb(n29797), .dout(n29800));
  jand g11778(.dina(n29800), .dinb(n324), .dout(n29801));
  jnot g11779(.din(n29801), .dout(n29802));
  jand g11780(.dina(n29592), .dinb(n29430), .dout(n29803));
  jxor g11781(.dina(n29484), .dinb(n29483), .dout(n29804));
  jand g11782(.dina(n29804), .dinb(n29591), .dout(n29805));
  jor  g11783(.dina(n29805), .dinb(n29803), .dout(n29806));
  jand g11784(.dina(n29806), .dinb(n323), .dout(n29807));
  jnot g11785(.din(n29807), .dout(n29808));
  jand g11786(.dina(n29592), .dinb(n29435), .dout(n29809));
  jxor g11787(.dina(n29481), .dinb(n29480), .dout(n29810));
  jand g11788(.dina(n29810), .dinb(n29591), .dout(n29811));
  jor  g11789(.dina(n29811), .dinb(n29809), .dout(n29812));
  jand g11790(.dina(n29812), .dinb(n335), .dout(n29813));
  jnot g11791(.din(n29813), .dout(n29814));
  jand g11792(.dina(n29592), .dinb(n29440), .dout(n29815));
  jxor g11793(.dina(n29478), .dinb(n29477), .dout(n29816));
  jand g11794(.dina(n29816), .dinb(n29591), .dout(n29817));
  jor  g11795(.dina(n29817), .dinb(n29815), .dout(n29818));
  jand g11796(.dina(n29818), .dinb(n334), .dout(n29819));
  jnot g11797(.din(n29819), .dout(n29820));
  jand g11798(.dina(n29592), .dinb(n29445), .dout(n29821));
  jxor g11799(.dina(n29475), .dinb(n29474), .dout(n29822));
  jand g11800(.dina(n29822), .dinb(n29591), .dout(n29823));
  jor  g11801(.dina(n29823), .dinb(n29821), .dout(n29824));
  jand g11802(.dina(n29824), .dinb(n338), .dout(n29825));
  jnot g11803(.din(n29825), .dout(n29826));
  jand g11804(.dina(n29592), .dinb(n29450), .dout(n29827));
  jxor g11805(.dina(n29472), .dinb(n29471), .dout(n29828));
  jand g11806(.dina(n29828), .dinb(n29591), .dout(n29829));
  jor  g11807(.dina(n29829), .dinb(n29827), .dout(n29830));
  jand g11808(.dina(n29830), .dinb(n337), .dout(n29831));
  jnot g11809(.din(n29831), .dout(n29832));
  jnot g11810(.din(n29455), .dout(n29833));
  jor  g11811(.dina(n29591), .dinb(n29833), .dout(n29834));
  jxor g11812(.dina(n29469), .dinb(n29468), .dout(n29835));
  jnot g11813(.din(n29835), .dout(n29836));
  jor  g11814(.dina(n29836), .dinb(n29592), .dout(n29837));
  jand g11815(.dina(n29837), .dinb(n29834), .dout(n29838));
  jnot g11816(.din(n29838), .dout(n29839));
  jand g11817(.dina(n29839), .dinb(n344), .dout(n29840));
  jnot g11818(.din(n29840), .dout(n29841));
  jor  g11819(.dina(n29591), .dinb(n29465), .dout(n29842));
  jxor g11820(.dina(n29466), .dinb(n9017), .dout(n29843));
  jand g11821(.dina(n29843), .dinb(n29591), .dout(n29844));
  jnot g11822(.din(n29844), .dout(n29845));
  jand g11823(.dina(n29845), .dinb(n29842), .dout(n29846));
  jnot g11824(.din(n29846), .dout(n29847));
  jand g11825(.dina(n29847), .dinb(n348), .dout(n29848));
  jnot g11826(.din(n29848), .dout(n29849));
  jnot g11827(.din(n8659), .dout(n29850));
  jnot g11828(.din(n29254), .dout(n29851));
  jnot g11829(.din(n29261), .dout(n29852));
  jnot g11830(.din(n29266), .dout(n29853));
  jnot g11831(.din(n29271), .dout(n29854));
  jnot g11832(.din(n29276), .dout(n29855));
  jnot g11833(.din(n29281), .dout(n29856));
  jnot g11834(.din(n29286), .dout(n29857));
  jnot g11835(.din(n29291), .dout(n29858));
  jnot g11836(.din(n29296), .dout(n29859));
  jnot g11837(.din(n29301), .dout(n29860));
  jnot g11838(.din(n29306), .dout(n29861));
  jnot g11839(.din(n29311), .dout(n29862));
  jnot g11840(.din(n29316), .dout(n29863));
  jnot g11841(.din(n29321), .dout(n29864));
  jnot g11842(.din(n29326), .dout(n29865));
  jnot g11843(.din(n29331), .dout(n29866));
  jnot g11844(.din(n29336), .dout(n29867));
  jnot g11845(.din(n29341), .dout(n29868));
  jnot g11846(.din(n29346), .dout(n29869));
  jnot g11847(.din(n29351), .dout(n29870));
  jnot g11848(.din(n29356), .dout(n29871));
  jnot g11849(.din(n29361), .dout(n29872));
  jnot g11850(.din(n29366), .dout(n29873));
  jnot g11851(.din(n29371), .dout(n29874));
  jnot g11852(.din(n29376), .dout(n29875));
  jnot g11853(.din(n29381), .dout(n29876));
  jnot g11854(.din(n29386), .dout(n29877));
  jnot g11855(.din(n29391), .dout(n29878));
  jnot g11856(.din(n29396), .dout(n29879));
  jnot g11857(.din(n29401), .dout(n29880));
  jnot g11858(.din(n29406), .dout(n29881));
  jnot g11859(.din(n29411), .dout(n29882));
  jnot g11860(.din(n29416), .dout(n29883));
  jnot g11861(.din(n29421), .dout(n29884));
  jnot g11862(.din(n29426), .dout(n29885));
  jnot g11863(.din(n29431), .dout(n29886));
  jnot g11864(.din(n29436), .dout(n29887));
  jnot g11865(.din(n29441), .dout(n29888));
  jnot g11866(.din(n29446), .dout(n29889));
  jnot g11867(.din(n29451), .dout(n29890));
  jnot g11868(.din(n29456), .dout(n29891));
  jnot g11869(.din(n29462), .dout(n29892));
  jxor g11870(.dina(n29465), .dinb(n258), .dout(n29893));
  jor  g11871(.dina(n29893), .dinb(n9016), .dout(n29894));
  jand g11872(.dina(n29894), .dinb(n29892), .dout(n29895));
  jnot g11873(.din(n29469), .dout(n29896));
  jor  g11874(.dina(n29896), .dinb(n29895), .dout(n29897));
  jand g11875(.dina(n29897), .dinb(n29891), .dout(n29898));
  jnot g11876(.din(n29472), .dout(n29899));
  jor  g11877(.dina(n29899), .dinb(n29898), .dout(n29900));
  jand g11878(.dina(n29900), .dinb(n29890), .dout(n29901));
  jnot g11879(.din(n29475), .dout(n29902));
  jor  g11880(.dina(n29902), .dinb(n29901), .dout(n29903));
  jand g11881(.dina(n29903), .dinb(n29889), .dout(n29904));
  jnot g11882(.din(n29478), .dout(n29905));
  jor  g11883(.dina(n29905), .dinb(n29904), .dout(n29906));
  jand g11884(.dina(n29906), .dinb(n29888), .dout(n29907));
  jnot g11885(.din(n29481), .dout(n29908));
  jor  g11886(.dina(n29908), .dinb(n29907), .dout(n29909));
  jand g11887(.dina(n29909), .dinb(n29887), .dout(n29910));
  jnot g11888(.din(n29484), .dout(n29911));
  jor  g11889(.dina(n29911), .dinb(n29910), .dout(n29912));
  jand g11890(.dina(n29912), .dinb(n29886), .dout(n29913));
  jnot g11891(.din(n29487), .dout(n29914));
  jor  g11892(.dina(n29914), .dinb(n29913), .dout(n29915));
  jand g11893(.dina(n29915), .dinb(n29885), .dout(n29916));
  jnot g11894(.din(n29490), .dout(n29917));
  jor  g11895(.dina(n29917), .dinb(n29916), .dout(n29918));
  jand g11896(.dina(n29918), .dinb(n29884), .dout(n29919));
  jnot g11897(.din(n29493), .dout(n29920));
  jor  g11898(.dina(n29920), .dinb(n29919), .dout(n29921));
  jand g11899(.dina(n29921), .dinb(n29883), .dout(n29922));
  jnot g11900(.din(n29496), .dout(n29923));
  jor  g11901(.dina(n29923), .dinb(n29922), .dout(n29924));
  jand g11902(.dina(n29924), .dinb(n29882), .dout(n29925));
  jnot g11903(.din(n29499), .dout(n29926));
  jor  g11904(.dina(n29926), .dinb(n29925), .dout(n29927));
  jand g11905(.dina(n29927), .dinb(n29881), .dout(n29928));
  jnot g11906(.din(n29502), .dout(n29929));
  jor  g11907(.dina(n29929), .dinb(n29928), .dout(n29930));
  jand g11908(.dina(n29930), .dinb(n29880), .dout(n29931));
  jnot g11909(.din(n29505), .dout(n29932));
  jor  g11910(.dina(n29932), .dinb(n29931), .dout(n29933));
  jand g11911(.dina(n29933), .dinb(n29879), .dout(n29934));
  jnot g11912(.din(n29508), .dout(n29935));
  jor  g11913(.dina(n29935), .dinb(n29934), .dout(n29936));
  jand g11914(.dina(n29936), .dinb(n29878), .dout(n29937));
  jnot g11915(.din(n29511), .dout(n29938));
  jor  g11916(.dina(n29938), .dinb(n29937), .dout(n29939));
  jand g11917(.dina(n29939), .dinb(n29877), .dout(n29940));
  jnot g11918(.din(n29514), .dout(n29941));
  jor  g11919(.dina(n29941), .dinb(n29940), .dout(n29942));
  jand g11920(.dina(n29942), .dinb(n29876), .dout(n29943));
  jnot g11921(.din(n29517), .dout(n29944));
  jor  g11922(.dina(n29944), .dinb(n29943), .dout(n29945));
  jand g11923(.dina(n29945), .dinb(n29875), .dout(n29946));
  jnot g11924(.din(n29520), .dout(n29947));
  jor  g11925(.dina(n29947), .dinb(n29946), .dout(n29948));
  jand g11926(.dina(n29948), .dinb(n29874), .dout(n29949));
  jnot g11927(.din(n29523), .dout(n29950));
  jor  g11928(.dina(n29950), .dinb(n29949), .dout(n29951));
  jand g11929(.dina(n29951), .dinb(n29873), .dout(n29952));
  jnot g11930(.din(n29526), .dout(n29953));
  jor  g11931(.dina(n29953), .dinb(n29952), .dout(n29954));
  jand g11932(.dina(n29954), .dinb(n29872), .dout(n29955));
  jnot g11933(.din(n29529), .dout(n29956));
  jor  g11934(.dina(n29956), .dinb(n29955), .dout(n29957));
  jand g11935(.dina(n29957), .dinb(n29871), .dout(n29958));
  jnot g11936(.din(n29532), .dout(n29959));
  jor  g11937(.dina(n29959), .dinb(n29958), .dout(n29960));
  jand g11938(.dina(n29960), .dinb(n29870), .dout(n29961));
  jnot g11939(.din(n29535), .dout(n29962));
  jor  g11940(.dina(n29962), .dinb(n29961), .dout(n29963));
  jand g11941(.dina(n29963), .dinb(n29869), .dout(n29964));
  jnot g11942(.din(n29538), .dout(n29965));
  jor  g11943(.dina(n29965), .dinb(n29964), .dout(n29966));
  jand g11944(.dina(n29966), .dinb(n29868), .dout(n29967));
  jnot g11945(.din(n29541), .dout(n29968));
  jor  g11946(.dina(n29968), .dinb(n29967), .dout(n29969));
  jand g11947(.dina(n29969), .dinb(n29867), .dout(n29970));
  jnot g11948(.din(n29544), .dout(n29971));
  jor  g11949(.dina(n29971), .dinb(n29970), .dout(n29972));
  jand g11950(.dina(n29972), .dinb(n29866), .dout(n29973));
  jnot g11951(.din(n29547), .dout(n29974));
  jor  g11952(.dina(n29974), .dinb(n29973), .dout(n29975));
  jand g11953(.dina(n29975), .dinb(n29865), .dout(n29976));
  jnot g11954(.din(n29550), .dout(n29977));
  jor  g11955(.dina(n29977), .dinb(n29976), .dout(n29978));
  jand g11956(.dina(n29978), .dinb(n29864), .dout(n29979));
  jnot g11957(.din(n29553), .dout(n29980));
  jor  g11958(.dina(n29980), .dinb(n29979), .dout(n29981));
  jand g11959(.dina(n29981), .dinb(n29863), .dout(n29982));
  jnot g11960(.din(n29556), .dout(n29983));
  jor  g11961(.dina(n29983), .dinb(n29982), .dout(n29984));
  jand g11962(.dina(n29984), .dinb(n29862), .dout(n29985));
  jnot g11963(.din(n29559), .dout(n29986));
  jor  g11964(.dina(n29986), .dinb(n29985), .dout(n29987));
  jand g11965(.dina(n29987), .dinb(n29861), .dout(n29988));
  jnot g11966(.din(n29562), .dout(n29989));
  jor  g11967(.dina(n29989), .dinb(n29988), .dout(n29990));
  jand g11968(.dina(n29990), .dinb(n29860), .dout(n29991));
  jnot g11969(.din(n29565), .dout(n29992));
  jor  g11970(.dina(n29992), .dinb(n29991), .dout(n29993));
  jand g11971(.dina(n29993), .dinb(n29859), .dout(n29994));
  jnot g11972(.din(n29568), .dout(n29995));
  jor  g11973(.dina(n29995), .dinb(n29994), .dout(n29996));
  jand g11974(.dina(n29996), .dinb(n29858), .dout(n29997));
  jnot g11975(.din(n29571), .dout(n29998));
  jor  g11976(.dina(n29998), .dinb(n29997), .dout(n29999));
  jand g11977(.dina(n29999), .dinb(n29857), .dout(n30000));
  jnot g11978(.din(n29574), .dout(n30001));
  jor  g11979(.dina(n30001), .dinb(n30000), .dout(n30002));
  jand g11980(.dina(n30002), .dinb(n29856), .dout(n30003));
  jnot g11981(.din(n29577), .dout(n30004));
  jor  g11982(.dina(n30004), .dinb(n30003), .dout(n30005));
  jand g11983(.dina(n30005), .dinb(n29855), .dout(n30006));
  jnot g11984(.din(n29580), .dout(n30007));
  jor  g11985(.dina(n30007), .dinb(n30006), .dout(n30008));
  jand g11986(.dina(n30008), .dinb(n29854), .dout(n30009));
  jnot g11987(.din(n29583), .dout(n30010));
  jor  g11988(.dina(n30010), .dinb(n30009), .dout(n30011));
  jand g11989(.dina(n30011), .dinb(n29853), .dout(n30012));
  jnot g11990(.din(n29586), .dout(n30013));
  jor  g11991(.dina(n30013), .dinb(n30012), .dout(n30014));
  jand g11992(.dina(n30014), .dinb(n29852), .dout(n30015));
  jand g11993(.dina(n30015), .dinb(n29851), .dout(n30016));
  jor  g11994(.dina(n30016), .dinb(n29252), .dout(n30017));
  jor  g11995(.dina(n30017), .dinb(n29850), .dout(n30018));
  jand g11996(.dina(n30018), .dinb(a21 ), .dout(n30019));
  jnot g11997(.din(n9354), .dout(n30020));
  jor  g11998(.dina(n30017), .dinb(n30020), .dout(n30021));
  jnot g11999(.din(n30021), .dout(n30022));
  jor  g12000(.dina(n30022), .dinb(n30019), .dout(n30023));
  jand g12001(.dina(n30023), .dinb(n258), .dout(n30024));
  jnot g12002(.din(n30024), .dout(n30025));
  jand g12003(.dina(n29590), .dinb(n8659), .dout(n30026));
  jor  g12004(.dina(n30026), .dinb(n9015), .dout(n30027));
  jand g12005(.dina(n30021), .dinb(n30027), .dout(n30028));
  jxor g12006(.dina(n30028), .dinb(n258), .dout(n30029));
  jor  g12007(.dina(n30029), .dinb(n9361), .dout(n30030));
  jand g12008(.dina(n30030), .dinb(n30025), .dout(n30031));
  jxor g12009(.dina(n29846), .dinb(b2 ), .dout(n30032));
  jnot g12010(.din(n30032), .dout(n30033));
  jor  g12011(.dina(n30033), .dinb(n30031), .dout(n30034));
  jand g12012(.dina(n30034), .dinb(n29849), .dout(n30035));
  jxor g12013(.dina(n29838), .dinb(b3 ), .dout(n30036));
  jnot g12014(.din(n30036), .dout(n30037));
  jor  g12015(.dina(n30037), .dinb(n30035), .dout(n30038));
  jand g12016(.dina(n30038), .dinb(n29841), .dout(n30039));
  jxor g12017(.dina(n29830), .dinb(n337), .dout(n30040));
  jnot g12018(.din(n30040), .dout(n30041));
  jor  g12019(.dina(n30041), .dinb(n30039), .dout(n30042));
  jand g12020(.dina(n30042), .dinb(n29832), .dout(n30043));
  jxor g12021(.dina(n29824), .dinb(n338), .dout(n30044));
  jnot g12022(.din(n30044), .dout(n30045));
  jor  g12023(.dina(n30045), .dinb(n30043), .dout(n30046));
  jand g12024(.dina(n30046), .dinb(n29826), .dout(n30047));
  jxor g12025(.dina(n29818), .dinb(n334), .dout(n30048));
  jnot g12026(.din(n30048), .dout(n30049));
  jor  g12027(.dina(n30049), .dinb(n30047), .dout(n30050));
  jand g12028(.dina(n30050), .dinb(n29820), .dout(n30051));
  jxor g12029(.dina(n29812), .dinb(n335), .dout(n30052));
  jnot g12030(.din(n30052), .dout(n30053));
  jor  g12031(.dina(n30053), .dinb(n30051), .dout(n30054));
  jand g12032(.dina(n30054), .dinb(n29814), .dout(n30055));
  jxor g12033(.dina(n29806), .dinb(n323), .dout(n30056));
  jnot g12034(.din(n30056), .dout(n30057));
  jor  g12035(.dina(n30057), .dinb(n30055), .dout(n30058));
  jand g12036(.dina(n30058), .dinb(n29808), .dout(n30059));
  jxor g12037(.dina(n29800), .dinb(n324), .dout(n30060));
  jnot g12038(.din(n30060), .dout(n30061));
  jor  g12039(.dina(n30061), .dinb(n30059), .dout(n30062));
  jand g12040(.dina(n30062), .dinb(n29802), .dout(n30063));
  jxor g12041(.dina(n29794), .dinb(n325), .dout(n30064));
  jnot g12042(.din(n30064), .dout(n30065));
  jor  g12043(.dina(n30065), .dinb(n30063), .dout(n30066));
  jand g12044(.dina(n30066), .dinb(n29796), .dout(n30067));
  jxor g12045(.dina(n29788), .dinb(n439), .dout(n30068));
  jnot g12046(.din(n30068), .dout(n30069));
  jor  g12047(.dina(n30069), .dinb(n30067), .dout(n30070));
  jand g12048(.dina(n30070), .dinb(n29790), .dout(n30071));
  jxor g12049(.dina(n29782), .dinb(n440), .dout(n30072));
  jnot g12050(.din(n30072), .dout(n30073));
  jor  g12051(.dina(n30073), .dinb(n30071), .dout(n30074));
  jand g12052(.dina(n30074), .dinb(n29784), .dout(n30075));
  jxor g12053(.dina(n29776), .dinb(n435), .dout(n30076));
  jnot g12054(.din(n30076), .dout(n30077));
  jor  g12055(.dina(n30077), .dinb(n30075), .dout(n30078));
  jand g12056(.dina(n30078), .dinb(n29778), .dout(n30079));
  jxor g12057(.dina(n29770), .dinb(n436), .dout(n30080));
  jnot g12058(.din(n30080), .dout(n30081));
  jor  g12059(.dina(n30081), .dinb(n30079), .dout(n30082));
  jand g12060(.dina(n30082), .dinb(n29772), .dout(n30083));
  jxor g12061(.dina(n29764), .dinb(n432), .dout(n30084));
  jnot g12062(.din(n30084), .dout(n30085));
  jor  g12063(.dina(n30085), .dinb(n30083), .dout(n30086));
  jand g12064(.dina(n30086), .dinb(n29766), .dout(n30087));
  jxor g12065(.dina(n29758), .dinb(n433), .dout(n30088));
  jnot g12066(.din(n30088), .dout(n30089));
  jor  g12067(.dina(n30089), .dinb(n30087), .dout(n30090));
  jand g12068(.dina(n30090), .dinb(n29760), .dout(n30091));
  jxor g12069(.dina(n29752), .dinb(n421), .dout(n30092));
  jnot g12070(.din(n30092), .dout(n30093));
  jor  g12071(.dina(n30093), .dinb(n30091), .dout(n30094));
  jand g12072(.dina(n30094), .dinb(n29754), .dout(n30095));
  jxor g12073(.dina(n29746), .dinb(n422), .dout(n30096));
  jnot g12074(.din(n30096), .dout(n30097));
  jor  g12075(.dina(n30097), .dinb(n30095), .dout(n30098));
  jand g12076(.dina(n30098), .dinb(n29748), .dout(n30099));
  jxor g12077(.dina(n29740), .dinb(n416), .dout(n30100));
  jnot g12078(.din(n30100), .dout(n30101));
  jor  g12079(.dina(n30101), .dinb(n30099), .dout(n30102));
  jand g12080(.dina(n30102), .dinb(n29742), .dout(n30103));
  jxor g12081(.dina(n29734), .dinb(n417), .dout(n30104));
  jnot g12082(.din(n30104), .dout(n30105));
  jor  g12083(.dina(n30105), .dinb(n30103), .dout(n30106));
  jand g12084(.dina(n30106), .dinb(n29736), .dout(n30107));
  jxor g12085(.dina(n29728), .dinb(n2547), .dout(n30108));
  jnot g12086(.din(n30108), .dout(n30109));
  jor  g12087(.dina(n30109), .dinb(n30107), .dout(n30110));
  jand g12088(.dina(n30110), .dinb(n29730), .dout(n30111));
  jxor g12089(.dina(n29722), .dinb(n2714), .dout(n30112));
  jnot g12090(.din(n30112), .dout(n30113));
  jor  g12091(.dina(n30113), .dinb(n30111), .dout(n30114));
  jand g12092(.dina(n30114), .dinb(n29724), .dout(n30115));
  jxor g12093(.dina(n29716), .dinb(n405), .dout(n30116));
  jnot g12094(.din(n30116), .dout(n30117));
  jor  g12095(.dina(n30117), .dinb(n30115), .dout(n30118));
  jand g12096(.dina(n30118), .dinb(n29718), .dout(n30119));
  jxor g12097(.dina(n29710), .dinb(n406), .dout(n30120));
  jnot g12098(.din(n30120), .dout(n30121));
  jor  g12099(.dina(n30121), .dinb(n30119), .dout(n30122));
  jand g12100(.dina(n30122), .dinb(n29712), .dout(n30123));
  jxor g12101(.dina(n29704), .dinb(n412), .dout(n30124));
  jnot g12102(.din(n30124), .dout(n30125));
  jor  g12103(.dina(n30125), .dinb(n30123), .dout(n30126));
  jand g12104(.dina(n30126), .dinb(n29706), .dout(n30127));
  jxor g12105(.dina(n29698), .dinb(n413), .dout(n30128));
  jnot g12106(.din(n30128), .dout(n30129));
  jor  g12107(.dina(n30129), .dinb(n30127), .dout(n30130));
  jand g12108(.dina(n30130), .dinb(n29700), .dout(n30131));
  jxor g12109(.dina(n29692), .dinb(n409), .dout(n30132));
  jnot g12110(.din(n30132), .dout(n30133));
  jor  g12111(.dina(n30133), .dinb(n30131), .dout(n30134));
  jand g12112(.dina(n30134), .dinb(n29694), .dout(n30135));
  jxor g12113(.dina(n29686), .dinb(n410), .dout(n30136));
  jnot g12114(.din(n30136), .dout(n30137));
  jor  g12115(.dina(n30137), .dinb(n30135), .dout(n30138));
  jand g12116(.dina(n30138), .dinb(n29688), .dout(n30139));
  jxor g12117(.dina(n29680), .dinb(n426), .dout(n30140));
  jnot g12118(.din(n30140), .dout(n30141));
  jor  g12119(.dina(n30141), .dinb(n30139), .dout(n30142));
  jand g12120(.dina(n30142), .dinb(n29682), .dout(n30143));
  jxor g12121(.dina(n29674), .dinb(n427), .dout(n30144));
  jnot g12122(.din(n30144), .dout(n30145));
  jor  g12123(.dina(n30145), .dinb(n30143), .dout(n30146));
  jand g12124(.dina(n30146), .dinb(n29676), .dout(n30147));
  jxor g12125(.dina(n29668), .dinb(n424), .dout(n30148));
  jnot g12126(.din(n30148), .dout(n30149));
  jor  g12127(.dina(n30149), .dinb(n30147), .dout(n30150));
  jand g12128(.dina(n30150), .dinb(n29670), .dout(n30151));
  jxor g12129(.dina(n29662), .dinb(n300), .dout(n30152));
  jnot g12130(.din(n30152), .dout(n30153));
  jor  g12131(.dina(n30153), .dinb(n30151), .dout(n30154));
  jand g12132(.dina(n30154), .dinb(n29664), .dout(n30155));
  jxor g12133(.dina(n29656), .dinb(n297), .dout(n30156));
  jnot g12134(.din(n30156), .dout(n30157));
  jor  g12135(.dina(n30157), .dinb(n30155), .dout(n30158));
  jand g12136(.dina(n30158), .dinb(n29658), .dout(n30159));
  jxor g12137(.dina(n29650), .dinb(n298), .dout(n30160));
  jnot g12138(.din(n30160), .dout(n30161));
  jor  g12139(.dina(n30161), .dinb(n30159), .dout(n30162));
  jand g12140(.dina(n30162), .dinb(n29652), .dout(n30163));
  jxor g12141(.dina(n29644), .dinb(n301), .dout(n30164));
  jnot g12142(.din(n30164), .dout(n30165));
  jor  g12143(.dina(n30165), .dinb(n30163), .dout(n30166));
  jand g12144(.dina(n30166), .dinb(n29646), .dout(n30167));
  jxor g12145(.dina(n29638), .dinb(n293), .dout(n30168));
  jnot g12146(.din(n30168), .dout(n30169));
  jor  g12147(.dina(n30169), .dinb(n30167), .dout(n30170));
  jand g12148(.dina(n30170), .dinb(n29640), .dout(n30171));
  jxor g12149(.dina(n29632), .dinb(n294), .dout(n30172));
  jnot g12150(.din(n30172), .dout(n30173));
  jor  g12151(.dina(n30173), .dinb(n30171), .dout(n30174));
  jand g12152(.dina(n30174), .dinb(n29634), .dout(n30175));
  jxor g12153(.dina(n29626), .dinb(n290), .dout(n30176));
  jnot g12154(.din(n30176), .dout(n30177));
  jor  g12155(.dina(n30177), .dinb(n30175), .dout(n30178));
  jand g12156(.dina(n30178), .dinb(n29628), .dout(n30179));
  jxor g12157(.dina(n29620), .dinb(n291), .dout(n30180));
  jnot g12158(.din(n30180), .dout(n30181));
  jor  g12159(.dina(n30181), .dinb(n30179), .dout(n30182));
  jand g12160(.dina(n30182), .dinb(n29622), .dout(n30183));
  jxor g12161(.dina(n29614), .dinb(n284), .dout(n30184));
  jnot g12162(.din(n30184), .dout(n30185));
  jor  g12163(.dina(n30185), .dinb(n30183), .dout(n30186));
  jand g12164(.dina(n30186), .dinb(n29616), .dout(n30187));
  jxor g12165(.dina(n29608), .dinb(n285), .dout(n30188));
  jnot g12166(.din(n30188), .dout(n30189));
  jor  g12167(.dina(n30189), .dinb(n30187), .dout(n30190));
  jand g12168(.dina(n30190), .dinb(n29610), .dout(n30191));
  jxor g12169(.dina(n29602), .dinb(n281), .dout(n30192));
  jnot g12170(.din(n30192), .dout(n30193));
  jor  g12171(.dina(n30193), .dinb(n30191), .dout(n30194));
  jand g12172(.dina(n30194), .dinb(n29604), .dout(n30195));
  jxor g12173(.dina(n29596), .dinb(b43 ), .dout(n30196));
  jor  g12174(.dina(n30196), .dinb(n30195), .dout(n30197));
  jor  g12175(.dina(n30197), .dinb(n280), .dout(n30198));
  jand g12176(.dina(n30198), .dinb(n29598), .dout(n30199));
  jand g12177(.dina(n30199), .dinb(n29596), .dout(n30200));
  jnot g12178(.din(n30200), .dout(n30201));
  jxor g12179(.dina(n30028), .dinb(b1 ), .dout(n30202));
  jand g12180(.dina(n30202), .dinb(n9362), .dout(n30203));
  jor  g12181(.dina(n30203), .dinb(n30024), .dout(n30204));
  jand g12182(.dina(n30032), .dinb(n30204), .dout(n30205));
  jor  g12183(.dina(n30205), .dinb(n29848), .dout(n30206));
  jand g12184(.dina(n30036), .dinb(n30206), .dout(n30207));
  jor  g12185(.dina(n30207), .dinb(n29840), .dout(n30208));
  jand g12186(.dina(n30040), .dinb(n30208), .dout(n30209));
  jor  g12187(.dina(n30209), .dinb(n29831), .dout(n30210));
  jand g12188(.dina(n30044), .dinb(n30210), .dout(n30211));
  jor  g12189(.dina(n30211), .dinb(n29825), .dout(n30212));
  jand g12190(.dina(n30048), .dinb(n30212), .dout(n30213));
  jor  g12191(.dina(n30213), .dinb(n29819), .dout(n30214));
  jand g12192(.dina(n30052), .dinb(n30214), .dout(n30215));
  jor  g12193(.dina(n30215), .dinb(n29813), .dout(n30216));
  jand g12194(.dina(n30056), .dinb(n30216), .dout(n30217));
  jor  g12195(.dina(n30217), .dinb(n29807), .dout(n30218));
  jand g12196(.dina(n30060), .dinb(n30218), .dout(n30219));
  jor  g12197(.dina(n30219), .dinb(n29801), .dout(n30220));
  jand g12198(.dina(n30064), .dinb(n30220), .dout(n30221));
  jor  g12199(.dina(n30221), .dinb(n29795), .dout(n30222));
  jand g12200(.dina(n30068), .dinb(n30222), .dout(n30223));
  jor  g12201(.dina(n30223), .dinb(n29789), .dout(n30224));
  jand g12202(.dina(n30072), .dinb(n30224), .dout(n30225));
  jor  g12203(.dina(n30225), .dinb(n29783), .dout(n30226));
  jand g12204(.dina(n30076), .dinb(n30226), .dout(n30227));
  jor  g12205(.dina(n30227), .dinb(n29777), .dout(n30228));
  jand g12206(.dina(n30080), .dinb(n30228), .dout(n30229));
  jor  g12207(.dina(n30229), .dinb(n29771), .dout(n30230));
  jand g12208(.dina(n30084), .dinb(n30230), .dout(n30231));
  jor  g12209(.dina(n30231), .dinb(n29765), .dout(n30232));
  jand g12210(.dina(n30088), .dinb(n30232), .dout(n30233));
  jor  g12211(.dina(n30233), .dinb(n29759), .dout(n30234));
  jand g12212(.dina(n30092), .dinb(n30234), .dout(n30235));
  jor  g12213(.dina(n30235), .dinb(n29753), .dout(n30236));
  jand g12214(.dina(n30096), .dinb(n30236), .dout(n30237));
  jor  g12215(.dina(n30237), .dinb(n29747), .dout(n30238));
  jand g12216(.dina(n30100), .dinb(n30238), .dout(n30239));
  jor  g12217(.dina(n30239), .dinb(n29741), .dout(n30240));
  jand g12218(.dina(n30104), .dinb(n30240), .dout(n30241));
  jor  g12219(.dina(n30241), .dinb(n29735), .dout(n30242));
  jand g12220(.dina(n30108), .dinb(n30242), .dout(n30243));
  jor  g12221(.dina(n30243), .dinb(n29729), .dout(n30244));
  jand g12222(.dina(n30112), .dinb(n30244), .dout(n30245));
  jor  g12223(.dina(n30245), .dinb(n29723), .dout(n30246));
  jand g12224(.dina(n30116), .dinb(n30246), .dout(n30247));
  jor  g12225(.dina(n30247), .dinb(n29717), .dout(n30248));
  jand g12226(.dina(n30120), .dinb(n30248), .dout(n30249));
  jor  g12227(.dina(n30249), .dinb(n29711), .dout(n30250));
  jand g12228(.dina(n30124), .dinb(n30250), .dout(n30251));
  jor  g12229(.dina(n30251), .dinb(n29705), .dout(n30252));
  jand g12230(.dina(n30128), .dinb(n30252), .dout(n30253));
  jor  g12231(.dina(n30253), .dinb(n29699), .dout(n30254));
  jand g12232(.dina(n30132), .dinb(n30254), .dout(n30255));
  jor  g12233(.dina(n30255), .dinb(n29693), .dout(n30256));
  jand g12234(.dina(n30136), .dinb(n30256), .dout(n30257));
  jor  g12235(.dina(n30257), .dinb(n29687), .dout(n30258));
  jand g12236(.dina(n30140), .dinb(n30258), .dout(n30259));
  jor  g12237(.dina(n30259), .dinb(n29681), .dout(n30260));
  jand g12238(.dina(n30144), .dinb(n30260), .dout(n30261));
  jor  g12239(.dina(n30261), .dinb(n29675), .dout(n30262));
  jand g12240(.dina(n30148), .dinb(n30262), .dout(n30263));
  jor  g12241(.dina(n30263), .dinb(n29669), .dout(n30264));
  jand g12242(.dina(n30152), .dinb(n30264), .dout(n30265));
  jor  g12243(.dina(n30265), .dinb(n29663), .dout(n30266));
  jand g12244(.dina(n30156), .dinb(n30266), .dout(n30267));
  jor  g12245(.dina(n30267), .dinb(n29657), .dout(n30268));
  jand g12246(.dina(n30160), .dinb(n30268), .dout(n30269));
  jor  g12247(.dina(n30269), .dinb(n29651), .dout(n30270));
  jand g12248(.dina(n30164), .dinb(n30270), .dout(n30271));
  jor  g12249(.dina(n30271), .dinb(n29645), .dout(n30272));
  jand g12250(.dina(n30168), .dinb(n30272), .dout(n30273));
  jor  g12251(.dina(n30273), .dinb(n29639), .dout(n30274));
  jand g12252(.dina(n30172), .dinb(n30274), .dout(n30275));
  jor  g12253(.dina(n30275), .dinb(n29633), .dout(n30276));
  jand g12254(.dina(n30176), .dinb(n30276), .dout(n30277));
  jor  g12255(.dina(n30277), .dinb(n29627), .dout(n30278));
  jand g12256(.dina(n30180), .dinb(n30278), .dout(n30279));
  jor  g12257(.dina(n30279), .dinb(n29621), .dout(n30280));
  jand g12258(.dina(n30184), .dinb(n30280), .dout(n30281));
  jor  g12259(.dina(n30281), .dinb(n29615), .dout(n30282));
  jand g12260(.dina(n30188), .dinb(n30282), .dout(n30283));
  jor  g12261(.dina(n30283), .dinb(n29609), .dout(n30284));
  jand g12262(.dina(n30192), .dinb(n30284), .dout(n30285));
  jor  g12263(.dina(n30285), .dinb(n29603), .dout(n30286));
  jnot g12264(.din(n30196), .dout(n30287));
  jand g12265(.dina(n30287), .dinb(n30286), .dout(n30288));
  jand g12266(.dina(n30195), .dinb(n282), .dout(n30289));
  jor  g12267(.dina(n30289), .dinb(n29598), .dout(n30290));
  jor  g12268(.dina(n30290), .dinb(n30288), .dout(n30291));
  jand g12269(.dina(n30291), .dinb(n30201), .dout(n30292));
  jand g12270(.dina(n30199), .dinb(n29602), .dout(n30293));
  jand g12271(.dina(n30288), .dinb(n588), .dout(n30294));
  jor  g12272(.dina(n30294), .dinb(n29597), .dout(n30295));
  jxor g12273(.dina(n30192), .dinb(n30284), .dout(n30296));
  jand g12274(.dina(n30296), .dinb(n30295), .dout(n30297));
  jor  g12275(.dina(n30297), .dinb(n30293), .dout(n30298));
  jand g12276(.dina(n30298), .dinb(n282), .dout(n30299));
  jnot g12277(.din(n30299), .dout(n30300));
  jand g12278(.dina(n30199), .dinb(n29608), .dout(n30301));
  jxor g12279(.dina(n30188), .dinb(n30282), .dout(n30302));
  jand g12280(.dina(n30302), .dinb(n30295), .dout(n30303));
  jor  g12281(.dina(n30303), .dinb(n30301), .dout(n30304));
  jand g12282(.dina(n30304), .dinb(n281), .dout(n30305));
  jnot g12283(.din(n30305), .dout(n30306));
  jand g12284(.dina(n30199), .dinb(n29614), .dout(n30307));
  jxor g12285(.dina(n30184), .dinb(n30280), .dout(n30308));
  jand g12286(.dina(n30308), .dinb(n30295), .dout(n30309));
  jor  g12287(.dina(n30309), .dinb(n30307), .dout(n30310));
  jand g12288(.dina(n30310), .dinb(n285), .dout(n30311));
  jnot g12289(.din(n30311), .dout(n30312));
  jand g12290(.dina(n30199), .dinb(n29620), .dout(n30313));
  jxor g12291(.dina(n30180), .dinb(n30278), .dout(n30314));
  jand g12292(.dina(n30314), .dinb(n30295), .dout(n30315));
  jor  g12293(.dina(n30315), .dinb(n30313), .dout(n30316));
  jand g12294(.dina(n30316), .dinb(n284), .dout(n30317));
  jnot g12295(.din(n30317), .dout(n30318));
  jand g12296(.dina(n30199), .dinb(n29626), .dout(n30319));
  jxor g12297(.dina(n30176), .dinb(n30276), .dout(n30320));
  jand g12298(.dina(n30320), .dinb(n30295), .dout(n30321));
  jor  g12299(.dina(n30321), .dinb(n30319), .dout(n30322));
  jand g12300(.dina(n30322), .dinb(n291), .dout(n30323));
  jnot g12301(.din(n30323), .dout(n30324));
  jand g12302(.dina(n30199), .dinb(n29632), .dout(n30325));
  jxor g12303(.dina(n30172), .dinb(n30274), .dout(n30326));
  jand g12304(.dina(n30326), .dinb(n30295), .dout(n30327));
  jor  g12305(.dina(n30327), .dinb(n30325), .dout(n30328));
  jand g12306(.dina(n30328), .dinb(n290), .dout(n30329));
  jnot g12307(.din(n30329), .dout(n30330));
  jand g12308(.dina(n30199), .dinb(n29638), .dout(n30331));
  jxor g12309(.dina(n30168), .dinb(n30272), .dout(n30332));
  jand g12310(.dina(n30332), .dinb(n30295), .dout(n30333));
  jor  g12311(.dina(n30333), .dinb(n30331), .dout(n30334));
  jand g12312(.dina(n30334), .dinb(n294), .dout(n30335));
  jnot g12313(.din(n30335), .dout(n30336));
  jand g12314(.dina(n30199), .dinb(n29644), .dout(n30337));
  jxor g12315(.dina(n30164), .dinb(n30270), .dout(n30338));
  jand g12316(.dina(n30338), .dinb(n30295), .dout(n30339));
  jor  g12317(.dina(n30339), .dinb(n30337), .dout(n30340));
  jand g12318(.dina(n30340), .dinb(n293), .dout(n30341));
  jnot g12319(.din(n30341), .dout(n30342));
  jand g12320(.dina(n30199), .dinb(n29650), .dout(n30343));
  jxor g12321(.dina(n30160), .dinb(n30268), .dout(n30344));
  jand g12322(.dina(n30344), .dinb(n30295), .dout(n30345));
  jor  g12323(.dina(n30345), .dinb(n30343), .dout(n30346));
  jand g12324(.dina(n30346), .dinb(n301), .dout(n30347));
  jnot g12325(.din(n30347), .dout(n30348));
  jand g12326(.dina(n30199), .dinb(n29656), .dout(n30349));
  jxor g12327(.dina(n30156), .dinb(n30266), .dout(n30350));
  jand g12328(.dina(n30350), .dinb(n30295), .dout(n30351));
  jor  g12329(.dina(n30351), .dinb(n30349), .dout(n30352));
  jand g12330(.dina(n30352), .dinb(n298), .dout(n30353));
  jnot g12331(.din(n30353), .dout(n30354));
  jand g12332(.dina(n30199), .dinb(n29662), .dout(n30355));
  jxor g12333(.dina(n30152), .dinb(n30264), .dout(n30356));
  jand g12334(.dina(n30356), .dinb(n30295), .dout(n30357));
  jor  g12335(.dina(n30357), .dinb(n30355), .dout(n30358));
  jand g12336(.dina(n30358), .dinb(n297), .dout(n30359));
  jnot g12337(.din(n30359), .dout(n30360));
  jand g12338(.dina(n30199), .dinb(n29668), .dout(n30361));
  jxor g12339(.dina(n30148), .dinb(n30262), .dout(n30362));
  jand g12340(.dina(n30362), .dinb(n30295), .dout(n30363));
  jor  g12341(.dina(n30363), .dinb(n30361), .dout(n30364));
  jand g12342(.dina(n30364), .dinb(n300), .dout(n30365));
  jnot g12343(.din(n30365), .dout(n30366));
  jand g12344(.dina(n30199), .dinb(n29674), .dout(n30367));
  jxor g12345(.dina(n30144), .dinb(n30260), .dout(n30368));
  jand g12346(.dina(n30368), .dinb(n30295), .dout(n30369));
  jor  g12347(.dina(n30369), .dinb(n30367), .dout(n30370));
  jand g12348(.dina(n30370), .dinb(n424), .dout(n30371));
  jnot g12349(.din(n30371), .dout(n30372));
  jand g12350(.dina(n30199), .dinb(n29680), .dout(n30373));
  jxor g12351(.dina(n30140), .dinb(n30258), .dout(n30374));
  jand g12352(.dina(n30374), .dinb(n30295), .dout(n30375));
  jor  g12353(.dina(n30375), .dinb(n30373), .dout(n30376));
  jand g12354(.dina(n30376), .dinb(n427), .dout(n30377));
  jnot g12355(.din(n30377), .dout(n30378));
  jand g12356(.dina(n30199), .dinb(n29686), .dout(n30379));
  jxor g12357(.dina(n30136), .dinb(n30256), .dout(n30380));
  jand g12358(.dina(n30380), .dinb(n30295), .dout(n30381));
  jor  g12359(.dina(n30381), .dinb(n30379), .dout(n30382));
  jand g12360(.dina(n30382), .dinb(n426), .dout(n30383));
  jnot g12361(.din(n30383), .dout(n30384));
  jand g12362(.dina(n30199), .dinb(n29692), .dout(n30385));
  jxor g12363(.dina(n30132), .dinb(n30254), .dout(n30386));
  jand g12364(.dina(n30386), .dinb(n30295), .dout(n30387));
  jor  g12365(.dina(n30387), .dinb(n30385), .dout(n30388));
  jand g12366(.dina(n30388), .dinb(n410), .dout(n30389));
  jnot g12367(.din(n30389), .dout(n30390));
  jand g12368(.dina(n30199), .dinb(n29698), .dout(n30391));
  jxor g12369(.dina(n30128), .dinb(n30252), .dout(n30392));
  jand g12370(.dina(n30392), .dinb(n30295), .dout(n30393));
  jor  g12371(.dina(n30393), .dinb(n30391), .dout(n30394));
  jand g12372(.dina(n30394), .dinb(n409), .dout(n30395));
  jnot g12373(.din(n30395), .dout(n30396));
  jand g12374(.dina(n30199), .dinb(n29704), .dout(n30397));
  jxor g12375(.dina(n30124), .dinb(n30250), .dout(n30398));
  jand g12376(.dina(n30398), .dinb(n30295), .dout(n30399));
  jor  g12377(.dina(n30399), .dinb(n30397), .dout(n30400));
  jand g12378(.dina(n30400), .dinb(n413), .dout(n30401));
  jnot g12379(.din(n30401), .dout(n30402));
  jand g12380(.dina(n30199), .dinb(n29710), .dout(n30403));
  jxor g12381(.dina(n30120), .dinb(n30248), .dout(n30404));
  jand g12382(.dina(n30404), .dinb(n30295), .dout(n30405));
  jor  g12383(.dina(n30405), .dinb(n30403), .dout(n30406));
  jand g12384(.dina(n30406), .dinb(n412), .dout(n30407));
  jnot g12385(.din(n30407), .dout(n30408));
  jand g12386(.dina(n30199), .dinb(n29716), .dout(n30409));
  jxor g12387(.dina(n30116), .dinb(n30246), .dout(n30410));
  jand g12388(.dina(n30410), .dinb(n30295), .dout(n30411));
  jor  g12389(.dina(n30411), .dinb(n30409), .dout(n30412));
  jand g12390(.dina(n30412), .dinb(n406), .dout(n30413));
  jnot g12391(.din(n30413), .dout(n30414));
  jand g12392(.dina(n30199), .dinb(n29722), .dout(n30415));
  jxor g12393(.dina(n30112), .dinb(n30244), .dout(n30416));
  jand g12394(.dina(n30416), .dinb(n30295), .dout(n30417));
  jor  g12395(.dina(n30417), .dinb(n30415), .dout(n30418));
  jand g12396(.dina(n30418), .dinb(n405), .dout(n30419));
  jnot g12397(.din(n30419), .dout(n30420));
  jand g12398(.dina(n30199), .dinb(n29728), .dout(n30421));
  jxor g12399(.dina(n30108), .dinb(n30242), .dout(n30422));
  jand g12400(.dina(n30422), .dinb(n30295), .dout(n30423));
  jor  g12401(.dina(n30423), .dinb(n30421), .dout(n30424));
  jand g12402(.dina(n30424), .dinb(n2714), .dout(n30425));
  jnot g12403(.din(n30425), .dout(n30426));
  jand g12404(.dina(n30199), .dinb(n29734), .dout(n30427));
  jxor g12405(.dina(n30104), .dinb(n30240), .dout(n30428));
  jand g12406(.dina(n30428), .dinb(n30295), .dout(n30429));
  jor  g12407(.dina(n30429), .dinb(n30427), .dout(n30430));
  jand g12408(.dina(n30430), .dinb(n2547), .dout(n30431));
  jnot g12409(.din(n30431), .dout(n30432));
  jand g12410(.dina(n30199), .dinb(n29740), .dout(n30433));
  jxor g12411(.dina(n30100), .dinb(n30238), .dout(n30434));
  jand g12412(.dina(n30434), .dinb(n30295), .dout(n30435));
  jor  g12413(.dina(n30435), .dinb(n30433), .dout(n30436));
  jand g12414(.dina(n30436), .dinb(n417), .dout(n30437));
  jnot g12415(.din(n30437), .dout(n30438));
  jand g12416(.dina(n30199), .dinb(n29746), .dout(n30439));
  jxor g12417(.dina(n30096), .dinb(n30236), .dout(n30440));
  jand g12418(.dina(n30440), .dinb(n30295), .dout(n30441));
  jor  g12419(.dina(n30441), .dinb(n30439), .dout(n30442));
  jand g12420(.dina(n30442), .dinb(n416), .dout(n30443));
  jnot g12421(.din(n30443), .dout(n30444));
  jand g12422(.dina(n30199), .dinb(n29752), .dout(n30445));
  jxor g12423(.dina(n30092), .dinb(n30234), .dout(n30446));
  jand g12424(.dina(n30446), .dinb(n30295), .dout(n30447));
  jor  g12425(.dina(n30447), .dinb(n30445), .dout(n30448));
  jand g12426(.dina(n30448), .dinb(n422), .dout(n30449));
  jnot g12427(.din(n30449), .dout(n30450));
  jand g12428(.dina(n30199), .dinb(n29758), .dout(n30451));
  jxor g12429(.dina(n30088), .dinb(n30232), .dout(n30452));
  jand g12430(.dina(n30452), .dinb(n30295), .dout(n30453));
  jor  g12431(.dina(n30453), .dinb(n30451), .dout(n30454));
  jand g12432(.dina(n30454), .dinb(n421), .dout(n30455));
  jnot g12433(.din(n30455), .dout(n30456));
  jand g12434(.dina(n30199), .dinb(n29764), .dout(n30457));
  jxor g12435(.dina(n30084), .dinb(n30230), .dout(n30458));
  jand g12436(.dina(n30458), .dinb(n30295), .dout(n30459));
  jor  g12437(.dina(n30459), .dinb(n30457), .dout(n30460));
  jand g12438(.dina(n30460), .dinb(n433), .dout(n30461));
  jnot g12439(.din(n30461), .dout(n30462));
  jand g12440(.dina(n30199), .dinb(n29770), .dout(n30463));
  jxor g12441(.dina(n30080), .dinb(n30228), .dout(n30464));
  jand g12442(.dina(n30464), .dinb(n30295), .dout(n30465));
  jor  g12443(.dina(n30465), .dinb(n30463), .dout(n30466));
  jand g12444(.dina(n30466), .dinb(n432), .dout(n30467));
  jnot g12445(.din(n30467), .dout(n30468));
  jand g12446(.dina(n30199), .dinb(n29776), .dout(n30469));
  jxor g12447(.dina(n30076), .dinb(n30226), .dout(n30470));
  jand g12448(.dina(n30470), .dinb(n30295), .dout(n30471));
  jor  g12449(.dina(n30471), .dinb(n30469), .dout(n30472));
  jand g12450(.dina(n30472), .dinb(n436), .dout(n30473));
  jnot g12451(.din(n30473), .dout(n30474));
  jand g12452(.dina(n30199), .dinb(n29782), .dout(n30475));
  jxor g12453(.dina(n30072), .dinb(n30224), .dout(n30476));
  jand g12454(.dina(n30476), .dinb(n30295), .dout(n30477));
  jor  g12455(.dina(n30477), .dinb(n30475), .dout(n30478));
  jand g12456(.dina(n30478), .dinb(n435), .dout(n30479));
  jnot g12457(.din(n30479), .dout(n30480));
  jand g12458(.dina(n30199), .dinb(n29788), .dout(n30481));
  jxor g12459(.dina(n30068), .dinb(n30222), .dout(n30482));
  jand g12460(.dina(n30482), .dinb(n30295), .dout(n30483));
  jor  g12461(.dina(n30483), .dinb(n30481), .dout(n30484));
  jand g12462(.dina(n30484), .dinb(n440), .dout(n30485));
  jnot g12463(.din(n30485), .dout(n30486));
  jand g12464(.dina(n30199), .dinb(n29794), .dout(n30487));
  jxor g12465(.dina(n30064), .dinb(n30220), .dout(n30488));
  jand g12466(.dina(n30488), .dinb(n30295), .dout(n30489));
  jor  g12467(.dina(n30489), .dinb(n30487), .dout(n30490));
  jand g12468(.dina(n30490), .dinb(n439), .dout(n30491));
  jnot g12469(.din(n30491), .dout(n30492));
  jand g12470(.dina(n30199), .dinb(n29800), .dout(n30493));
  jxor g12471(.dina(n30060), .dinb(n30218), .dout(n30494));
  jand g12472(.dina(n30494), .dinb(n30295), .dout(n30495));
  jor  g12473(.dina(n30495), .dinb(n30493), .dout(n30496));
  jand g12474(.dina(n30496), .dinb(n325), .dout(n30497));
  jnot g12475(.din(n30497), .dout(n30498));
  jand g12476(.dina(n30199), .dinb(n29806), .dout(n30499));
  jxor g12477(.dina(n30056), .dinb(n30216), .dout(n30500));
  jand g12478(.dina(n30500), .dinb(n30295), .dout(n30501));
  jor  g12479(.dina(n30501), .dinb(n30499), .dout(n30502));
  jand g12480(.dina(n30502), .dinb(n324), .dout(n30503));
  jnot g12481(.din(n30503), .dout(n30504));
  jand g12482(.dina(n30199), .dinb(n29812), .dout(n30505));
  jxor g12483(.dina(n30052), .dinb(n30214), .dout(n30506));
  jand g12484(.dina(n30506), .dinb(n30295), .dout(n30507));
  jor  g12485(.dina(n30507), .dinb(n30505), .dout(n30508));
  jand g12486(.dina(n30508), .dinb(n323), .dout(n30509));
  jnot g12487(.din(n30509), .dout(n30510));
  jand g12488(.dina(n30199), .dinb(n29818), .dout(n30511));
  jxor g12489(.dina(n30048), .dinb(n30212), .dout(n30512));
  jand g12490(.dina(n30512), .dinb(n30295), .dout(n30513));
  jor  g12491(.dina(n30513), .dinb(n30511), .dout(n30514));
  jand g12492(.dina(n30514), .dinb(n335), .dout(n30515));
  jnot g12493(.din(n30515), .dout(n30516));
  jand g12494(.dina(n30199), .dinb(n29824), .dout(n30517));
  jxor g12495(.dina(n30044), .dinb(n30210), .dout(n30518));
  jand g12496(.dina(n30518), .dinb(n30295), .dout(n30519));
  jor  g12497(.dina(n30519), .dinb(n30517), .dout(n30520));
  jand g12498(.dina(n30520), .dinb(n334), .dout(n30521));
  jnot g12499(.din(n30521), .dout(n30522));
  jand g12500(.dina(n30199), .dinb(n29830), .dout(n30523));
  jxor g12501(.dina(n30040), .dinb(n30208), .dout(n30524));
  jand g12502(.dina(n30524), .dinb(n30295), .dout(n30525));
  jor  g12503(.dina(n30525), .dinb(n30523), .dout(n30526));
  jand g12504(.dina(n30526), .dinb(n338), .dout(n30527));
  jnot g12505(.din(n30527), .dout(n30528));
  jand g12506(.dina(n30199), .dinb(n29839), .dout(n30529));
  jxor g12507(.dina(n30036), .dinb(n30206), .dout(n30530));
  jand g12508(.dina(n30530), .dinb(n30295), .dout(n30531));
  jor  g12509(.dina(n30531), .dinb(n30529), .dout(n30532));
  jand g12510(.dina(n30532), .dinb(n337), .dout(n30533));
  jnot g12511(.din(n30533), .dout(n30534));
  jand g12512(.dina(n30199), .dinb(n29847), .dout(n30535));
  jxor g12513(.dina(n30032), .dinb(n30204), .dout(n30536));
  jand g12514(.dina(n30536), .dinb(n30295), .dout(n30537));
  jor  g12515(.dina(n30537), .dinb(n30535), .dout(n30538));
  jand g12516(.dina(n30538), .dinb(n344), .dout(n30539));
  jnot g12517(.din(n30539), .dout(n30540));
  jand g12518(.dina(n30199), .dinb(n30023), .dout(n30541));
  jxor g12519(.dina(n30202), .dinb(n9362), .dout(n30542));
  jand g12520(.dina(n30542), .dinb(n30295), .dout(n30543));
  jor  g12521(.dina(n30543), .dinb(n30541), .dout(n30544));
  jand g12522(.dina(n30544), .dinb(n348), .dout(n30545));
  jnot g12523(.din(n30545), .dout(n30546));
  jor  g12524(.dina(n30199), .dinb(n18364), .dout(n30547));
  jand g12525(.dina(n30547), .dinb(a20 ), .dout(n30548));
  jor  g12526(.dina(n30199), .dinb(n9362), .dout(n30549));
  jnot g12527(.din(n30549), .dout(n30550));
  jor  g12528(.dina(n30550), .dinb(n30548), .dout(n30551));
  jand g12529(.dina(n30551), .dinb(n258), .dout(n30552));
  jnot g12530(.din(n30552), .dout(n30553));
  jand g12531(.dina(n30295), .dinb(b0 ), .dout(n30554));
  jor  g12532(.dina(n30554), .dinb(n9360), .dout(n30555));
  jand g12533(.dina(n30549), .dinb(n30555), .dout(n30556));
  jxor g12534(.dina(n30556), .dinb(n258), .dout(n30557));
  jor  g12535(.dina(n30557), .dinb(n9720), .dout(n30558));
  jand g12536(.dina(n30558), .dinb(n30553), .dout(n30559));
  jxor g12537(.dina(n30544), .dinb(n348), .dout(n30560));
  jnot g12538(.din(n30560), .dout(n30561));
  jor  g12539(.dina(n30561), .dinb(n30559), .dout(n30562));
  jand g12540(.dina(n30562), .dinb(n30546), .dout(n30563));
  jxor g12541(.dina(n30538), .dinb(n344), .dout(n30564));
  jnot g12542(.din(n30564), .dout(n30565));
  jor  g12543(.dina(n30565), .dinb(n30563), .dout(n30566));
  jand g12544(.dina(n30566), .dinb(n30540), .dout(n30567));
  jxor g12545(.dina(n30532), .dinb(n337), .dout(n30568));
  jnot g12546(.din(n30568), .dout(n30569));
  jor  g12547(.dina(n30569), .dinb(n30567), .dout(n30570));
  jand g12548(.dina(n30570), .dinb(n30534), .dout(n30571));
  jxor g12549(.dina(n30526), .dinb(n338), .dout(n30572));
  jnot g12550(.din(n30572), .dout(n30573));
  jor  g12551(.dina(n30573), .dinb(n30571), .dout(n30574));
  jand g12552(.dina(n30574), .dinb(n30528), .dout(n30575));
  jxor g12553(.dina(n30520), .dinb(n334), .dout(n30576));
  jnot g12554(.din(n30576), .dout(n30577));
  jor  g12555(.dina(n30577), .dinb(n30575), .dout(n30578));
  jand g12556(.dina(n30578), .dinb(n30522), .dout(n30579));
  jxor g12557(.dina(n30514), .dinb(n335), .dout(n30580));
  jnot g12558(.din(n30580), .dout(n30581));
  jor  g12559(.dina(n30581), .dinb(n30579), .dout(n30582));
  jand g12560(.dina(n30582), .dinb(n30516), .dout(n30583));
  jxor g12561(.dina(n30508), .dinb(n323), .dout(n30584));
  jnot g12562(.din(n30584), .dout(n30585));
  jor  g12563(.dina(n30585), .dinb(n30583), .dout(n30586));
  jand g12564(.dina(n30586), .dinb(n30510), .dout(n30587));
  jxor g12565(.dina(n30502), .dinb(n324), .dout(n30588));
  jnot g12566(.din(n30588), .dout(n30589));
  jor  g12567(.dina(n30589), .dinb(n30587), .dout(n30590));
  jand g12568(.dina(n30590), .dinb(n30504), .dout(n30591));
  jxor g12569(.dina(n30496), .dinb(n325), .dout(n30592));
  jnot g12570(.din(n30592), .dout(n30593));
  jor  g12571(.dina(n30593), .dinb(n30591), .dout(n30594));
  jand g12572(.dina(n30594), .dinb(n30498), .dout(n30595));
  jxor g12573(.dina(n30490), .dinb(n439), .dout(n30596));
  jnot g12574(.din(n30596), .dout(n30597));
  jor  g12575(.dina(n30597), .dinb(n30595), .dout(n30598));
  jand g12576(.dina(n30598), .dinb(n30492), .dout(n30599));
  jxor g12577(.dina(n30484), .dinb(n440), .dout(n30600));
  jnot g12578(.din(n30600), .dout(n30601));
  jor  g12579(.dina(n30601), .dinb(n30599), .dout(n30602));
  jand g12580(.dina(n30602), .dinb(n30486), .dout(n30603));
  jxor g12581(.dina(n30478), .dinb(n435), .dout(n30604));
  jnot g12582(.din(n30604), .dout(n30605));
  jor  g12583(.dina(n30605), .dinb(n30603), .dout(n30606));
  jand g12584(.dina(n30606), .dinb(n30480), .dout(n30607));
  jxor g12585(.dina(n30472), .dinb(n436), .dout(n30608));
  jnot g12586(.din(n30608), .dout(n30609));
  jor  g12587(.dina(n30609), .dinb(n30607), .dout(n30610));
  jand g12588(.dina(n30610), .dinb(n30474), .dout(n30611));
  jxor g12589(.dina(n30466), .dinb(n432), .dout(n30612));
  jnot g12590(.din(n30612), .dout(n30613));
  jor  g12591(.dina(n30613), .dinb(n30611), .dout(n30614));
  jand g12592(.dina(n30614), .dinb(n30468), .dout(n30615));
  jxor g12593(.dina(n30460), .dinb(n433), .dout(n30616));
  jnot g12594(.din(n30616), .dout(n30617));
  jor  g12595(.dina(n30617), .dinb(n30615), .dout(n30618));
  jand g12596(.dina(n30618), .dinb(n30462), .dout(n30619));
  jxor g12597(.dina(n30454), .dinb(n421), .dout(n30620));
  jnot g12598(.din(n30620), .dout(n30621));
  jor  g12599(.dina(n30621), .dinb(n30619), .dout(n30622));
  jand g12600(.dina(n30622), .dinb(n30456), .dout(n30623));
  jxor g12601(.dina(n30448), .dinb(n422), .dout(n30624));
  jnot g12602(.din(n30624), .dout(n30625));
  jor  g12603(.dina(n30625), .dinb(n30623), .dout(n30626));
  jand g12604(.dina(n30626), .dinb(n30450), .dout(n30627));
  jxor g12605(.dina(n30442), .dinb(n416), .dout(n30628));
  jnot g12606(.din(n30628), .dout(n30629));
  jor  g12607(.dina(n30629), .dinb(n30627), .dout(n30630));
  jand g12608(.dina(n30630), .dinb(n30444), .dout(n30631));
  jxor g12609(.dina(n30436), .dinb(n417), .dout(n30632));
  jnot g12610(.din(n30632), .dout(n30633));
  jor  g12611(.dina(n30633), .dinb(n30631), .dout(n30634));
  jand g12612(.dina(n30634), .dinb(n30438), .dout(n30635));
  jxor g12613(.dina(n30430), .dinb(n2547), .dout(n30636));
  jnot g12614(.din(n30636), .dout(n30637));
  jor  g12615(.dina(n30637), .dinb(n30635), .dout(n30638));
  jand g12616(.dina(n30638), .dinb(n30432), .dout(n30639));
  jxor g12617(.dina(n30424), .dinb(n2714), .dout(n30640));
  jnot g12618(.din(n30640), .dout(n30641));
  jor  g12619(.dina(n30641), .dinb(n30639), .dout(n30642));
  jand g12620(.dina(n30642), .dinb(n30426), .dout(n30643));
  jxor g12621(.dina(n30418), .dinb(n405), .dout(n30644));
  jnot g12622(.din(n30644), .dout(n30645));
  jor  g12623(.dina(n30645), .dinb(n30643), .dout(n30646));
  jand g12624(.dina(n30646), .dinb(n30420), .dout(n30647));
  jxor g12625(.dina(n30412), .dinb(n406), .dout(n30648));
  jnot g12626(.din(n30648), .dout(n30649));
  jor  g12627(.dina(n30649), .dinb(n30647), .dout(n30650));
  jand g12628(.dina(n30650), .dinb(n30414), .dout(n30651));
  jxor g12629(.dina(n30406), .dinb(n412), .dout(n30652));
  jnot g12630(.din(n30652), .dout(n30653));
  jor  g12631(.dina(n30653), .dinb(n30651), .dout(n30654));
  jand g12632(.dina(n30654), .dinb(n30408), .dout(n30655));
  jxor g12633(.dina(n30400), .dinb(n413), .dout(n30656));
  jnot g12634(.din(n30656), .dout(n30657));
  jor  g12635(.dina(n30657), .dinb(n30655), .dout(n30658));
  jand g12636(.dina(n30658), .dinb(n30402), .dout(n30659));
  jxor g12637(.dina(n30394), .dinb(n409), .dout(n30660));
  jnot g12638(.din(n30660), .dout(n30661));
  jor  g12639(.dina(n30661), .dinb(n30659), .dout(n30662));
  jand g12640(.dina(n30662), .dinb(n30396), .dout(n30663));
  jxor g12641(.dina(n30388), .dinb(n410), .dout(n30664));
  jnot g12642(.din(n30664), .dout(n30665));
  jor  g12643(.dina(n30665), .dinb(n30663), .dout(n30666));
  jand g12644(.dina(n30666), .dinb(n30390), .dout(n30667));
  jxor g12645(.dina(n30382), .dinb(n426), .dout(n30668));
  jnot g12646(.din(n30668), .dout(n30669));
  jor  g12647(.dina(n30669), .dinb(n30667), .dout(n30670));
  jand g12648(.dina(n30670), .dinb(n30384), .dout(n30671));
  jxor g12649(.dina(n30376), .dinb(n427), .dout(n30672));
  jnot g12650(.din(n30672), .dout(n30673));
  jor  g12651(.dina(n30673), .dinb(n30671), .dout(n30674));
  jand g12652(.dina(n30674), .dinb(n30378), .dout(n30675));
  jxor g12653(.dina(n30370), .dinb(n424), .dout(n30676));
  jnot g12654(.din(n30676), .dout(n30677));
  jor  g12655(.dina(n30677), .dinb(n30675), .dout(n30678));
  jand g12656(.dina(n30678), .dinb(n30372), .dout(n30679));
  jxor g12657(.dina(n30364), .dinb(n300), .dout(n30680));
  jnot g12658(.din(n30680), .dout(n30681));
  jor  g12659(.dina(n30681), .dinb(n30679), .dout(n30682));
  jand g12660(.dina(n30682), .dinb(n30366), .dout(n30683));
  jxor g12661(.dina(n30358), .dinb(n297), .dout(n30684));
  jnot g12662(.din(n30684), .dout(n30685));
  jor  g12663(.dina(n30685), .dinb(n30683), .dout(n30686));
  jand g12664(.dina(n30686), .dinb(n30360), .dout(n30687));
  jxor g12665(.dina(n30352), .dinb(n298), .dout(n30688));
  jnot g12666(.din(n30688), .dout(n30689));
  jor  g12667(.dina(n30689), .dinb(n30687), .dout(n30690));
  jand g12668(.dina(n30690), .dinb(n30354), .dout(n30691));
  jxor g12669(.dina(n30346), .dinb(n301), .dout(n30692));
  jnot g12670(.din(n30692), .dout(n30693));
  jor  g12671(.dina(n30693), .dinb(n30691), .dout(n30694));
  jand g12672(.dina(n30694), .dinb(n30348), .dout(n30695));
  jxor g12673(.dina(n30340), .dinb(n293), .dout(n30696));
  jnot g12674(.din(n30696), .dout(n30697));
  jor  g12675(.dina(n30697), .dinb(n30695), .dout(n30698));
  jand g12676(.dina(n30698), .dinb(n30342), .dout(n30699));
  jxor g12677(.dina(n30334), .dinb(n294), .dout(n30700));
  jnot g12678(.din(n30700), .dout(n30701));
  jor  g12679(.dina(n30701), .dinb(n30699), .dout(n30702));
  jand g12680(.dina(n30702), .dinb(n30336), .dout(n30703));
  jxor g12681(.dina(n30328), .dinb(n290), .dout(n30704));
  jnot g12682(.din(n30704), .dout(n30705));
  jor  g12683(.dina(n30705), .dinb(n30703), .dout(n30706));
  jand g12684(.dina(n30706), .dinb(n30330), .dout(n30707));
  jxor g12685(.dina(n30322), .dinb(n291), .dout(n30708));
  jnot g12686(.din(n30708), .dout(n30709));
  jor  g12687(.dina(n30709), .dinb(n30707), .dout(n30710));
  jand g12688(.dina(n30710), .dinb(n30324), .dout(n30711));
  jxor g12689(.dina(n30316), .dinb(n284), .dout(n30712));
  jnot g12690(.din(n30712), .dout(n30713));
  jor  g12691(.dina(n30713), .dinb(n30711), .dout(n30714));
  jand g12692(.dina(n30714), .dinb(n30318), .dout(n30715));
  jxor g12693(.dina(n30310), .dinb(n285), .dout(n30716));
  jnot g12694(.din(n30716), .dout(n30717));
  jor  g12695(.dina(n30717), .dinb(n30715), .dout(n30718));
  jand g12696(.dina(n30718), .dinb(n30312), .dout(n30719));
  jxor g12697(.dina(n30304), .dinb(n281), .dout(n30720));
  jnot g12698(.din(n30720), .dout(n30721));
  jor  g12699(.dina(n30721), .dinb(n30719), .dout(n30722));
  jand g12700(.dina(n30722), .dinb(n30306), .dout(n30723));
  jxor g12701(.dina(n30298), .dinb(n282), .dout(n30724));
  jnot g12702(.din(n30724), .dout(n30725));
  jor  g12703(.dina(n30725), .dinb(n30723), .dout(n30726));
  jand g12704(.dina(n30726), .dinb(n30300), .dout(n30727));
  jxor g12705(.dina(n30292), .dinb(n397), .dout(n30728));
  jnot g12706(.din(n30728), .dout(n30729));
  jand g12707(.dina(n30729), .dinb(n516), .dout(n30730));
  jnot g12708(.din(n30730), .dout(n30731));
  jor  g12709(.dina(n30731), .dinb(n30727), .dout(n30732));
  jand g12710(.dina(n30732), .dinb(n30292), .dout(n30733));
  jxor g12711(.dina(n30556), .dinb(b1 ), .dout(n30734));
  jand g12712(.dina(n30734), .dinb(n9721), .dout(n30735));
  jor  g12713(.dina(n30735), .dinb(n30552), .dout(n30736));
  jand g12714(.dina(n30560), .dinb(n30736), .dout(n30737));
  jor  g12715(.dina(n30737), .dinb(n30545), .dout(n30738));
  jand g12716(.dina(n30564), .dinb(n30738), .dout(n30739));
  jor  g12717(.dina(n30739), .dinb(n30539), .dout(n30740));
  jand g12718(.dina(n30568), .dinb(n30740), .dout(n30741));
  jor  g12719(.dina(n30741), .dinb(n30533), .dout(n30742));
  jand g12720(.dina(n30572), .dinb(n30742), .dout(n30743));
  jor  g12721(.dina(n30743), .dinb(n30527), .dout(n30744));
  jand g12722(.dina(n30576), .dinb(n30744), .dout(n30745));
  jor  g12723(.dina(n30745), .dinb(n30521), .dout(n30746));
  jand g12724(.dina(n30580), .dinb(n30746), .dout(n30747));
  jor  g12725(.dina(n30747), .dinb(n30515), .dout(n30748));
  jand g12726(.dina(n30584), .dinb(n30748), .dout(n30749));
  jor  g12727(.dina(n30749), .dinb(n30509), .dout(n30750));
  jand g12728(.dina(n30588), .dinb(n30750), .dout(n30751));
  jor  g12729(.dina(n30751), .dinb(n30503), .dout(n30752));
  jand g12730(.dina(n30592), .dinb(n30752), .dout(n30753));
  jor  g12731(.dina(n30753), .dinb(n30497), .dout(n30754));
  jand g12732(.dina(n30596), .dinb(n30754), .dout(n30755));
  jor  g12733(.dina(n30755), .dinb(n30491), .dout(n30756));
  jand g12734(.dina(n30600), .dinb(n30756), .dout(n30757));
  jor  g12735(.dina(n30757), .dinb(n30485), .dout(n30758));
  jand g12736(.dina(n30604), .dinb(n30758), .dout(n30759));
  jor  g12737(.dina(n30759), .dinb(n30479), .dout(n30760));
  jand g12738(.dina(n30608), .dinb(n30760), .dout(n30761));
  jor  g12739(.dina(n30761), .dinb(n30473), .dout(n30762));
  jand g12740(.dina(n30612), .dinb(n30762), .dout(n30763));
  jor  g12741(.dina(n30763), .dinb(n30467), .dout(n30764));
  jand g12742(.dina(n30616), .dinb(n30764), .dout(n30765));
  jor  g12743(.dina(n30765), .dinb(n30461), .dout(n30766));
  jand g12744(.dina(n30620), .dinb(n30766), .dout(n30767));
  jor  g12745(.dina(n30767), .dinb(n30455), .dout(n30768));
  jand g12746(.dina(n30624), .dinb(n30768), .dout(n30769));
  jor  g12747(.dina(n30769), .dinb(n30449), .dout(n30770));
  jand g12748(.dina(n30628), .dinb(n30770), .dout(n30771));
  jor  g12749(.dina(n30771), .dinb(n30443), .dout(n30772));
  jand g12750(.dina(n30632), .dinb(n30772), .dout(n30773));
  jor  g12751(.dina(n30773), .dinb(n30437), .dout(n30774));
  jand g12752(.dina(n30636), .dinb(n30774), .dout(n30775));
  jor  g12753(.dina(n30775), .dinb(n30431), .dout(n30776));
  jand g12754(.dina(n30640), .dinb(n30776), .dout(n30777));
  jor  g12755(.dina(n30777), .dinb(n30425), .dout(n30778));
  jand g12756(.dina(n30644), .dinb(n30778), .dout(n30779));
  jor  g12757(.dina(n30779), .dinb(n30419), .dout(n30780));
  jand g12758(.dina(n30648), .dinb(n30780), .dout(n30781));
  jor  g12759(.dina(n30781), .dinb(n30413), .dout(n30782));
  jand g12760(.dina(n30652), .dinb(n30782), .dout(n30783));
  jor  g12761(.dina(n30783), .dinb(n30407), .dout(n30784));
  jand g12762(.dina(n30656), .dinb(n30784), .dout(n30785));
  jor  g12763(.dina(n30785), .dinb(n30401), .dout(n30786));
  jand g12764(.dina(n30660), .dinb(n30786), .dout(n30787));
  jor  g12765(.dina(n30787), .dinb(n30395), .dout(n30788));
  jand g12766(.dina(n30664), .dinb(n30788), .dout(n30789));
  jor  g12767(.dina(n30789), .dinb(n30389), .dout(n30790));
  jand g12768(.dina(n30668), .dinb(n30790), .dout(n30791));
  jor  g12769(.dina(n30791), .dinb(n30383), .dout(n30792));
  jand g12770(.dina(n30672), .dinb(n30792), .dout(n30793));
  jor  g12771(.dina(n30793), .dinb(n30377), .dout(n30794));
  jand g12772(.dina(n30676), .dinb(n30794), .dout(n30795));
  jor  g12773(.dina(n30795), .dinb(n30371), .dout(n30796));
  jand g12774(.dina(n30680), .dinb(n30796), .dout(n30797));
  jor  g12775(.dina(n30797), .dinb(n30365), .dout(n30798));
  jand g12776(.dina(n30684), .dinb(n30798), .dout(n30799));
  jor  g12777(.dina(n30799), .dinb(n30359), .dout(n30800));
  jand g12778(.dina(n30688), .dinb(n30800), .dout(n30801));
  jor  g12779(.dina(n30801), .dinb(n30353), .dout(n30802));
  jand g12780(.dina(n30692), .dinb(n30802), .dout(n30803));
  jor  g12781(.dina(n30803), .dinb(n30347), .dout(n30804));
  jand g12782(.dina(n30696), .dinb(n30804), .dout(n30805));
  jor  g12783(.dina(n30805), .dinb(n30341), .dout(n30806));
  jand g12784(.dina(n30700), .dinb(n30806), .dout(n30807));
  jor  g12785(.dina(n30807), .dinb(n30335), .dout(n30808));
  jand g12786(.dina(n30704), .dinb(n30808), .dout(n30809));
  jor  g12787(.dina(n30809), .dinb(n30329), .dout(n30810));
  jand g12788(.dina(n30708), .dinb(n30810), .dout(n30811));
  jor  g12789(.dina(n30811), .dinb(n30323), .dout(n30812));
  jand g12790(.dina(n30712), .dinb(n30812), .dout(n30813));
  jor  g12791(.dina(n30813), .dinb(n30317), .dout(n30814));
  jand g12792(.dina(n30716), .dinb(n30814), .dout(n30815));
  jor  g12793(.dina(n30815), .dinb(n30311), .dout(n30816));
  jand g12794(.dina(n30720), .dinb(n30816), .dout(n30817));
  jor  g12795(.dina(n30817), .dinb(n30305), .dout(n30818));
  jand g12796(.dina(n30724), .dinb(n30818), .dout(n30819));
  jor  g12797(.dina(n30819), .dinb(n30299), .dout(n30820));
  jand g12798(.dina(n30730), .dinb(n30820), .dout(n30821));
  jor  g12799(.dina(n30292), .dinb(n280), .dout(n30822));
  jnot g12800(.din(n30822), .dout(n30823));
  jor  g12801(.dina(n30823), .dinb(n30821), .dout(n30824));
  jxor g12802(.dina(n30728), .dinb(n30820), .dout(n30825));
  jand g12803(.dina(n30825), .dinb(n30824), .dout(n30826));
  jor  g12804(.dina(n30826), .dinb(n30733), .dout(n30827));
  jnot g12805(.din(n30827), .dout(n30828));
  jand g12806(.dina(n30827), .dinb(b45 ), .dout(n30829));
  jnot g12807(.din(n30829), .dout(n30830));
  jand g12808(.dina(n30828), .dinb(n513), .dout(n30831));
  jand g12809(.dina(n30822), .dinb(n30732), .dout(n30832));
  jand g12810(.dina(n30832), .dinb(n30298), .dout(n30833));
  jxor g12811(.dina(n30724), .dinb(n30818), .dout(n30834));
  jand g12812(.dina(n30834), .dinb(n30824), .dout(n30835));
  jor  g12813(.dina(n30835), .dinb(n30833), .dout(n30836));
  jand g12814(.dina(n30836), .dinb(n397), .dout(n30837));
  jand g12815(.dina(n30832), .dinb(n30304), .dout(n30838));
  jxor g12816(.dina(n30720), .dinb(n30816), .dout(n30839));
  jand g12817(.dina(n30839), .dinb(n30824), .dout(n30840));
  jor  g12818(.dina(n30840), .dinb(n30838), .dout(n30841));
  jand g12819(.dina(n30841), .dinb(n282), .dout(n30842));
  jand g12820(.dina(n30832), .dinb(n30310), .dout(n30843));
  jxor g12821(.dina(n30716), .dinb(n30814), .dout(n30844));
  jand g12822(.dina(n30844), .dinb(n30824), .dout(n30845));
  jor  g12823(.dina(n30845), .dinb(n30843), .dout(n30846));
  jand g12824(.dina(n30846), .dinb(n281), .dout(n30847));
  jand g12825(.dina(n30832), .dinb(n30316), .dout(n30848));
  jxor g12826(.dina(n30712), .dinb(n30812), .dout(n30849));
  jand g12827(.dina(n30849), .dinb(n30824), .dout(n30850));
  jor  g12828(.dina(n30850), .dinb(n30848), .dout(n30851));
  jand g12829(.dina(n30851), .dinb(n285), .dout(n30852));
  jand g12830(.dina(n30832), .dinb(n30322), .dout(n30853));
  jxor g12831(.dina(n30708), .dinb(n30810), .dout(n30854));
  jand g12832(.dina(n30854), .dinb(n30824), .dout(n30855));
  jor  g12833(.dina(n30855), .dinb(n30853), .dout(n30856));
  jand g12834(.dina(n30856), .dinb(n284), .dout(n30857));
  jand g12835(.dina(n30832), .dinb(n30328), .dout(n30858));
  jxor g12836(.dina(n30704), .dinb(n30808), .dout(n30859));
  jand g12837(.dina(n30859), .dinb(n30824), .dout(n30860));
  jor  g12838(.dina(n30860), .dinb(n30858), .dout(n30861));
  jand g12839(.dina(n30861), .dinb(n291), .dout(n30862));
  jand g12840(.dina(n30832), .dinb(n30334), .dout(n30863));
  jxor g12841(.dina(n30700), .dinb(n30806), .dout(n30864));
  jand g12842(.dina(n30864), .dinb(n30824), .dout(n30865));
  jor  g12843(.dina(n30865), .dinb(n30863), .dout(n30866));
  jand g12844(.dina(n30866), .dinb(n290), .dout(n30867));
  jand g12845(.dina(n30832), .dinb(n30340), .dout(n30868));
  jxor g12846(.dina(n30696), .dinb(n30804), .dout(n30869));
  jand g12847(.dina(n30869), .dinb(n30824), .dout(n30870));
  jor  g12848(.dina(n30870), .dinb(n30868), .dout(n30871));
  jand g12849(.dina(n30871), .dinb(n294), .dout(n30872));
  jand g12850(.dina(n30832), .dinb(n30346), .dout(n30873));
  jxor g12851(.dina(n30692), .dinb(n30802), .dout(n30874));
  jand g12852(.dina(n30874), .dinb(n30824), .dout(n30875));
  jor  g12853(.dina(n30875), .dinb(n30873), .dout(n30876));
  jand g12854(.dina(n30876), .dinb(n293), .dout(n30877));
  jand g12855(.dina(n30832), .dinb(n30352), .dout(n30878));
  jxor g12856(.dina(n30688), .dinb(n30800), .dout(n30879));
  jand g12857(.dina(n30879), .dinb(n30824), .dout(n30880));
  jor  g12858(.dina(n30880), .dinb(n30878), .dout(n30881));
  jand g12859(.dina(n30881), .dinb(n301), .dout(n30882));
  jand g12860(.dina(n30832), .dinb(n30358), .dout(n30883));
  jxor g12861(.dina(n30684), .dinb(n30798), .dout(n30884));
  jand g12862(.dina(n30884), .dinb(n30824), .dout(n30885));
  jor  g12863(.dina(n30885), .dinb(n30883), .dout(n30886));
  jand g12864(.dina(n30886), .dinb(n298), .dout(n30887));
  jand g12865(.dina(n30832), .dinb(n30364), .dout(n30888));
  jxor g12866(.dina(n30680), .dinb(n30796), .dout(n30889));
  jand g12867(.dina(n30889), .dinb(n30824), .dout(n30890));
  jor  g12868(.dina(n30890), .dinb(n30888), .dout(n30891));
  jand g12869(.dina(n30891), .dinb(n297), .dout(n30892));
  jand g12870(.dina(n30832), .dinb(n30370), .dout(n30893));
  jxor g12871(.dina(n30676), .dinb(n30794), .dout(n30894));
  jand g12872(.dina(n30894), .dinb(n30824), .dout(n30895));
  jor  g12873(.dina(n30895), .dinb(n30893), .dout(n30896));
  jand g12874(.dina(n30896), .dinb(n300), .dout(n30897));
  jand g12875(.dina(n30832), .dinb(n30376), .dout(n30898));
  jxor g12876(.dina(n30672), .dinb(n30792), .dout(n30899));
  jand g12877(.dina(n30899), .dinb(n30824), .dout(n30900));
  jor  g12878(.dina(n30900), .dinb(n30898), .dout(n30901));
  jand g12879(.dina(n30901), .dinb(n424), .dout(n30902));
  jand g12880(.dina(n30832), .dinb(n30382), .dout(n30903));
  jxor g12881(.dina(n30668), .dinb(n30790), .dout(n30904));
  jand g12882(.dina(n30904), .dinb(n30824), .dout(n30905));
  jor  g12883(.dina(n30905), .dinb(n30903), .dout(n30906));
  jand g12884(.dina(n30906), .dinb(n427), .dout(n30907));
  jand g12885(.dina(n30832), .dinb(n30388), .dout(n30908));
  jxor g12886(.dina(n30664), .dinb(n30788), .dout(n30909));
  jand g12887(.dina(n30909), .dinb(n30824), .dout(n30910));
  jor  g12888(.dina(n30910), .dinb(n30908), .dout(n30911));
  jand g12889(.dina(n30911), .dinb(n426), .dout(n30912));
  jand g12890(.dina(n30832), .dinb(n30394), .dout(n30913));
  jxor g12891(.dina(n30660), .dinb(n30786), .dout(n30914));
  jand g12892(.dina(n30914), .dinb(n30824), .dout(n30915));
  jor  g12893(.dina(n30915), .dinb(n30913), .dout(n30916));
  jand g12894(.dina(n30916), .dinb(n410), .dout(n30917));
  jand g12895(.dina(n30832), .dinb(n30400), .dout(n30918));
  jxor g12896(.dina(n30656), .dinb(n30784), .dout(n30919));
  jand g12897(.dina(n30919), .dinb(n30824), .dout(n30920));
  jor  g12898(.dina(n30920), .dinb(n30918), .dout(n30921));
  jand g12899(.dina(n30921), .dinb(n409), .dout(n30922));
  jand g12900(.dina(n30832), .dinb(n30406), .dout(n30923));
  jxor g12901(.dina(n30652), .dinb(n30782), .dout(n30924));
  jand g12902(.dina(n30924), .dinb(n30824), .dout(n30925));
  jor  g12903(.dina(n30925), .dinb(n30923), .dout(n30926));
  jand g12904(.dina(n30926), .dinb(n413), .dout(n30927));
  jand g12905(.dina(n30832), .dinb(n30412), .dout(n30928));
  jxor g12906(.dina(n30648), .dinb(n30780), .dout(n30929));
  jand g12907(.dina(n30929), .dinb(n30824), .dout(n30930));
  jor  g12908(.dina(n30930), .dinb(n30928), .dout(n30931));
  jand g12909(.dina(n30931), .dinb(n412), .dout(n30932));
  jand g12910(.dina(n30832), .dinb(n30418), .dout(n30933));
  jxor g12911(.dina(n30644), .dinb(n30778), .dout(n30934));
  jand g12912(.dina(n30934), .dinb(n30824), .dout(n30935));
  jor  g12913(.dina(n30935), .dinb(n30933), .dout(n30936));
  jand g12914(.dina(n30936), .dinb(n406), .dout(n30937));
  jand g12915(.dina(n30832), .dinb(n30424), .dout(n30938));
  jxor g12916(.dina(n30640), .dinb(n30776), .dout(n30939));
  jand g12917(.dina(n30939), .dinb(n30824), .dout(n30940));
  jor  g12918(.dina(n30940), .dinb(n30938), .dout(n30941));
  jand g12919(.dina(n30941), .dinb(n405), .dout(n30942));
  jand g12920(.dina(n30832), .dinb(n30430), .dout(n30943));
  jxor g12921(.dina(n30636), .dinb(n30774), .dout(n30944));
  jand g12922(.dina(n30944), .dinb(n30824), .dout(n30945));
  jor  g12923(.dina(n30945), .dinb(n30943), .dout(n30946));
  jand g12924(.dina(n30946), .dinb(n2714), .dout(n30947));
  jand g12925(.dina(n30832), .dinb(n30436), .dout(n30948));
  jxor g12926(.dina(n30632), .dinb(n30772), .dout(n30949));
  jand g12927(.dina(n30949), .dinb(n30824), .dout(n30950));
  jor  g12928(.dina(n30950), .dinb(n30948), .dout(n30951));
  jand g12929(.dina(n30951), .dinb(n2547), .dout(n30952));
  jand g12930(.dina(n30832), .dinb(n30442), .dout(n30953));
  jxor g12931(.dina(n30628), .dinb(n30770), .dout(n30954));
  jand g12932(.dina(n30954), .dinb(n30824), .dout(n30955));
  jor  g12933(.dina(n30955), .dinb(n30953), .dout(n30956));
  jand g12934(.dina(n30956), .dinb(n417), .dout(n30957));
  jand g12935(.dina(n30832), .dinb(n30448), .dout(n30958));
  jxor g12936(.dina(n30624), .dinb(n30768), .dout(n30959));
  jand g12937(.dina(n30959), .dinb(n30824), .dout(n30960));
  jor  g12938(.dina(n30960), .dinb(n30958), .dout(n30961));
  jand g12939(.dina(n30961), .dinb(n416), .dout(n30962));
  jand g12940(.dina(n30832), .dinb(n30454), .dout(n30963));
  jxor g12941(.dina(n30620), .dinb(n30766), .dout(n30964));
  jand g12942(.dina(n30964), .dinb(n30824), .dout(n30965));
  jor  g12943(.dina(n30965), .dinb(n30963), .dout(n30966));
  jand g12944(.dina(n30966), .dinb(n422), .dout(n30967));
  jand g12945(.dina(n30832), .dinb(n30460), .dout(n30968));
  jxor g12946(.dina(n30616), .dinb(n30764), .dout(n30969));
  jand g12947(.dina(n30969), .dinb(n30824), .dout(n30970));
  jor  g12948(.dina(n30970), .dinb(n30968), .dout(n30971));
  jand g12949(.dina(n30971), .dinb(n421), .dout(n30972));
  jand g12950(.dina(n30832), .dinb(n30466), .dout(n30973));
  jxor g12951(.dina(n30612), .dinb(n30762), .dout(n30974));
  jand g12952(.dina(n30974), .dinb(n30824), .dout(n30975));
  jor  g12953(.dina(n30975), .dinb(n30973), .dout(n30976));
  jand g12954(.dina(n30976), .dinb(n433), .dout(n30977));
  jand g12955(.dina(n30832), .dinb(n30472), .dout(n30978));
  jxor g12956(.dina(n30608), .dinb(n30760), .dout(n30979));
  jand g12957(.dina(n30979), .dinb(n30824), .dout(n30980));
  jor  g12958(.dina(n30980), .dinb(n30978), .dout(n30981));
  jand g12959(.dina(n30981), .dinb(n432), .dout(n30982));
  jand g12960(.dina(n30832), .dinb(n30478), .dout(n30983));
  jxor g12961(.dina(n30604), .dinb(n30758), .dout(n30984));
  jand g12962(.dina(n30984), .dinb(n30824), .dout(n30985));
  jor  g12963(.dina(n30985), .dinb(n30983), .dout(n30986));
  jand g12964(.dina(n30986), .dinb(n436), .dout(n30987));
  jand g12965(.dina(n30832), .dinb(n30484), .dout(n30988));
  jxor g12966(.dina(n30600), .dinb(n30756), .dout(n30989));
  jand g12967(.dina(n30989), .dinb(n30824), .dout(n30990));
  jor  g12968(.dina(n30990), .dinb(n30988), .dout(n30991));
  jand g12969(.dina(n30991), .dinb(n435), .dout(n30992));
  jand g12970(.dina(n30832), .dinb(n30490), .dout(n30993));
  jxor g12971(.dina(n30596), .dinb(n30754), .dout(n30994));
  jand g12972(.dina(n30994), .dinb(n30824), .dout(n30995));
  jor  g12973(.dina(n30995), .dinb(n30993), .dout(n30996));
  jand g12974(.dina(n30996), .dinb(n440), .dout(n30997));
  jand g12975(.dina(n30832), .dinb(n30496), .dout(n30998));
  jxor g12976(.dina(n30592), .dinb(n30752), .dout(n30999));
  jand g12977(.dina(n30999), .dinb(n30824), .dout(n31000));
  jor  g12978(.dina(n31000), .dinb(n30998), .dout(n31001));
  jand g12979(.dina(n31001), .dinb(n439), .dout(n31002));
  jand g12980(.dina(n30832), .dinb(n30502), .dout(n31003));
  jxor g12981(.dina(n30588), .dinb(n30750), .dout(n31004));
  jand g12982(.dina(n31004), .dinb(n30824), .dout(n31005));
  jor  g12983(.dina(n31005), .dinb(n31003), .dout(n31006));
  jand g12984(.dina(n31006), .dinb(n325), .dout(n31007));
  jand g12985(.dina(n30832), .dinb(n30508), .dout(n31008));
  jxor g12986(.dina(n30584), .dinb(n30748), .dout(n31009));
  jand g12987(.dina(n31009), .dinb(n30824), .dout(n31010));
  jor  g12988(.dina(n31010), .dinb(n31008), .dout(n31011));
  jand g12989(.dina(n31011), .dinb(n324), .dout(n31012));
  jand g12990(.dina(n30832), .dinb(n30514), .dout(n31013));
  jxor g12991(.dina(n30580), .dinb(n30746), .dout(n31014));
  jand g12992(.dina(n31014), .dinb(n30824), .dout(n31015));
  jor  g12993(.dina(n31015), .dinb(n31013), .dout(n31016));
  jand g12994(.dina(n31016), .dinb(n323), .dout(n31017));
  jand g12995(.dina(n30832), .dinb(n30520), .dout(n31018));
  jxor g12996(.dina(n30576), .dinb(n30744), .dout(n31019));
  jand g12997(.dina(n31019), .dinb(n30824), .dout(n31020));
  jor  g12998(.dina(n31020), .dinb(n31018), .dout(n31021));
  jand g12999(.dina(n31021), .dinb(n335), .dout(n31022));
  jand g13000(.dina(n30832), .dinb(n30526), .dout(n31023));
  jxor g13001(.dina(n30572), .dinb(n30742), .dout(n31024));
  jand g13002(.dina(n31024), .dinb(n30824), .dout(n31025));
  jor  g13003(.dina(n31025), .dinb(n31023), .dout(n31026));
  jand g13004(.dina(n31026), .dinb(n334), .dout(n31027));
  jand g13005(.dina(n30832), .dinb(n30532), .dout(n31028));
  jxor g13006(.dina(n30568), .dinb(n30740), .dout(n31029));
  jand g13007(.dina(n31029), .dinb(n30824), .dout(n31030));
  jor  g13008(.dina(n31030), .dinb(n31028), .dout(n31031));
  jand g13009(.dina(n31031), .dinb(n338), .dout(n31032));
  jand g13010(.dina(n30832), .dinb(n30538), .dout(n31033));
  jxor g13011(.dina(n30564), .dinb(n30738), .dout(n31034));
  jand g13012(.dina(n31034), .dinb(n30824), .dout(n31035));
  jor  g13013(.dina(n31035), .dinb(n31033), .dout(n31036));
  jand g13014(.dina(n31036), .dinb(n337), .dout(n31037));
  jand g13015(.dina(n30832), .dinb(n30544), .dout(n31038));
  jxor g13016(.dina(n30560), .dinb(n30736), .dout(n31039));
  jand g13017(.dina(n31039), .dinb(n30824), .dout(n31040));
  jor  g13018(.dina(n31040), .dinb(n31038), .dout(n31041));
  jand g13019(.dina(n31041), .dinb(n344), .dout(n31042));
  jand g13020(.dina(n30832), .dinb(n30551), .dout(n31043));
  jxor g13021(.dina(n30734), .dinb(n9721), .dout(n31044));
  jand g13022(.dina(n31044), .dinb(n30824), .dout(n31045));
  jor  g13023(.dina(n31045), .dinb(n31043), .dout(n31046));
  jand g13024(.dina(n31046), .dinb(n348), .dout(n31047));
  jor  g13025(.dina(n30832), .dinb(n18364), .dout(n31048));
  jand g13026(.dina(n31048), .dinb(a19 ), .dout(n31049));
  jor  g13027(.dina(n30832), .dinb(n9721), .dout(n31050));
  jnot g13028(.din(n31050), .dout(n31051));
  jor  g13029(.dina(n31051), .dinb(n31049), .dout(n31052));
  jand g13030(.dina(n31052), .dinb(n258), .dout(n31053));
  jand g13031(.dina(n30824), .dinb(b0 ), .dout(n31054));
  jor  g13032(.dina(n31054), .dinb(n9719), .dout(n31055));
  jand g13033(.dina(n31050), .dinb(n31055), .dout(n31056));
  jxor g13034(.dina(n31056), .dinb(b1 ), .dout(n31057));
  jand g13035(.dina(n31057), .dinb(n10102), .dout(n31058));
  jor  g13036(.dina(n31058), .dinb(n31053), .dout(n31059));
  jxor g13037(.dina(n31046), .dinb(n348), .dout(n31060));
  jand g13038(.dina(n31060), .dinb(n31059), .dout(n31061));
  jor  g13039(.dina(n31061), .dinb(n31047), .dout(n31062));
  jxor g13040(.dina(n31041), .dinb(n344), .dout(n31063));
  jand g13041(.dina(n31063), .dinb(n31062), .dout(n31064));
  jor  g13042(.dina(n31064), .dinb(n31042), .dout(n31065));
  jxor g13043(.dina(n31036), .dinb(n337), .dout(n31066));
  jand g13044(.dina(n31066), .dinb(n31065), .dout(n31067));
  jor  g13045(.dina(n31067), .dinb(n31037), .dout(n31068));
  jxor g13046(.dina(n31031), .dinb(n338), .dout(n31069));
  jand g13047(.dina(n31069), .dinb(n31068), .dout(n31070));
  jor  g13048(.dina(n31070), .dinb(n31032), .dout(n31071));
  jxor g13049(.dina(n31026), .dinb(n334), .dout(n31072));
  jand g13050(.dina(n31072), .dinb(n31071), .dout(n31073));
  jor  g13051(.dina(n31073), .dinb(n31027), .dout(n31074));
  jxor g13052(.dina(n31021), .dinb(n335), .dout(n31075));
  jand g13053(.dina(n31075), .dinb(n31074), .dout(n31076));
  jor  g13054(.dina(n31076), .dinb(n31022), .dout(n31077));
  jxor g13055(.dina(n31016), .dinb(n323), .dout(n31078));
  jand g13056(.dina(n31078), .dinb(n31077), .dout(n31079));
  jor  g13057(.dina(n31079), .dinb(n31017), .dout(n31080));
  jxor g13058(.dina(n31011), .dinb(n324), .dout(n31081));
  jand g13059(.dina(n31081), .dinb(n31080), .dout(n31082));
  jor  g13060(.dina(n31082), .dinb(n31012), .dout(n31083));
  jxor g13061(.dina(n31006), .dinb(n325), .dout(n31084));
  jand g13062(.dina(n31084), .dinb(n31083), .dout(n31085));
  jor  g13063(.dina(n31085), .dinb(n31007), .dout(n31086));
  jxor g13064(.dina(n31001), .dinb(n439), .dout(n31087));
  jand g13065(.dina(n31087), .dinb(n31086), .dout(n31088));
  jor  g13066(.dina(n31088), .dinb(n31002), .dout(n31089));
  jxor g13067(.dina(n30996), .dinb(n440), .dout(n31090));
  jand g13068(.dina(n31090), .dinb(n31089), .dout(n31091));
  jor  g13069(.dina(n31091), .dinb(n30997), .dout(n31092));
  jxor g13070(.dina(n30991), .dinb(n435), .dout(n31093));
  jand g13071(.dina(n31093), .dinb(n31092), .dout(n31094));
  jor  g13072(.dina(n31094), .dinb(n30992), .dout(n31095));
  jxor g13073(.dina(n30986), .dinb(n436), .dout(n31096));
  jand g13074(.dina(n31096), .dinb(n31095), .dout(n31097));
  jor  g13075(.dina(n31097), .dinb(n30987), .dout(n31098));
  jxor g13076(.dina(n30981), .dinb(n432), .dout(n31099));
  jand g13077(.dina(n31099), .dinb(n31098), .dout(n31100));
  jor  g13078(.dina(n31100), .dinb(n30982), .dout(n31101));
  jxor g13079(.dina(n30976), .dinb(n433), .dout(n31102));
  jand g13080(.dina(n31102), .dinb(n31101), .dout(n31103));
  jor  g13081(.dina(n31103), .dinb(n30977), .dout(n31104));
  jxor g13082(.dina(n30971), .dinb(n421), .dout(n31105));
  jand g13083(.dina(n31105), .dinb(n31104), .dout(n31106));
  jor  g13084(.dina(n31106), .dinb(n30972), .dout(n31107));
  jxor g13085(.dina(n30966), .dinb(n422), .dout(n31108));
  jand g13086(.dina(n31108), .dinb(n31107), .dout(n31109));
  jor  g13087(.dina(n31109), .dinb(n30967), .dout(n31110));
  jxor g13088(.dina(n30961), .dinb(n416), .dout(n31111));
  jand g13089(.dina(n31111), .dinb(n31110), .dout(n31112));
  jor  g13090(.dina(n31112), .dinb(n30962), .dout(n31113));
  jxor g13091(.dina(n30956), .dinb(n417), .dout(n31114));
  jand g13092(.dina(n31114), .dinb(n31113), .dout(n31115));
  jor  g13093(.dina(n31115), .dinb(n30957), .dout(n31116));
  jxor g13094(.dina(n30951), .dinb(n2547), .dout(n31117));
  jand g13095(.dina(n31117), .dinb(n31116), .dout(n31118));
  jor  g13096(.dina(n31118), .dinb(n30952), .dout(n31119));
  jxor g13097(.dina(n30946), .dinb(n2714), .dout(n31120));
  jand g13098(.dina(n31120), .dinb(n31119), .dout(n31121));
  jor  g13099(.dina(n31121), .dinb(n30947), .dout(n31122));
  jxor g13100(.dina(n30941), .dinb(n405), .dout(n31123));
  jand g13101(.dina(n31123), .dinb(n31122), .dout(n31124));
  jor  g13102(.dina(n31124), .dinb(n30942), .dout(n31125));
  jxor g13103(.dina(n30936), .dinb(n406), .dout(n31126));
  jand g13104(.dina(n31126), .dinb(n31125), .dout(n31127));
  jor  g13105(.dina(n31127), .dinb(n30937), .dout(n31128));
  jxor g13106(.dina(n30931), .dinb(n412), .dout(n31129));
  jand g13107(.dina(n31129), .dinb(n31128), .dout(n31130));
  jor  g13108(.dina(n31130), .dinb(n30932), .dout(n31131));
  jxor g13109(.dina(n30926), .dinb(n413), .dout(n31132));
  jand g13110(.dina(n31132), .dinb(n31131), .dout(n31133));
  jor  g13111(.dina(n31133), .dinb(n30927), .dout(n31134));
  jxor g13112(.dina(n30921), .dinb(n409), .dout(n31135));
  jand g13113(.dina(n31135), .dinb(n31134), .dout(n31136));
  jor  g13114(.dina(n31136), .dinb(n30922), .dout(n31137));
  jxor g13115(.dina(n30916), .dinb(n410), .dout(n31138));
  jand g13116(.dina(n31138), .dinb(n31137), .dout(n31139));
  jor  g13117(.dina(n31139), .dinb(n30917), .dout(n31140));
  jxor g13118(.dina(n30911), .dinb(n426), .dout(n31141));
  jand g13119(.dina(n31141), .dinb(n31140), .dout(n31142));
  jor  g13120(.dina(n31142), .dinb(n30912), .dout(n31143));
  jxor g13121(.dina(n30906), .dinb(n427), .dout(n31144));
  jand g13122(.dina(n31144), .dinb(n31143), .dout(n31145));
  jor  g13123(.dina(n31145), .dinb(n30907), .dout(n31146));
  jxor g13124(.dina(n30901), .dinb(n424), .dout(n31147));
  jand g13125(.dina(n31147), .dinb(n31146), .dout(n31148));
  jor  g13126(.dina(n31148), .dinb(n30902), .dout(n31149));
  jxor g13127(.dina(n30896), .dinb(n300), .dout(n31150));
  jand g13128(.dina(n31150), .dinb(n31149), .dout(n31151));
  jor  g13129(.dina(n31151), .dinb(n30897), .dout(n31152));
  jxor g13130(.dina(n30891), .dinb(n297), .dout(n31153));
  jand g13131(.dina(n31153), .dinb(n31152), .dout(n31154));
  jor  g13132(.dina(n31154), .dinb(n30892), .dout(n31155));
  jxor g13133(.dina(n30886), .dinb(n298), .dout(n31156));
  jand g13134(.dina(n31156), .dinb(n31155), .dout(n31157));
  jor  g13135(.dina(n31157), .dinb(n30887), .dout(n31158));
  jxor g13136(.dina(n30881), .dinb(n301), .dout(n31159));
  jand g13137(.dina(n31159), .dinb(n31158), .dout(n31160));
  jor  g13138(.dina(n31160), .dinb(n30882), .dout(n31161));
  jxor g13139(.dina(n30876), .dinb(n293), .dout(n31162));
  jand g13140(.dina(n31162), .dinb(n31161), .dout(n31163));
  jor  g13141(.dina(n31163), .dinb(n30877), .dout(n31164));
  jxor g13142(.dina(n30871), .dinb(n294), .dout(n31165));
  jand g13143(.dina(n31165), .dinb(n31164), .dout(n31166));
  jor  g13144(.dina(n31166), .dinb(n30872), .dout(n31167));
  jxor g13145(.dina(n30866), .dinb(n290), .dout(n31168));
  jand g13146(.dina(n31168), .dinb(n31167), .dout(n31169));
  jor  g13147(.dina(n31169), .dinb(n30867), .dout(n31170));
  jxor g13148(.dina(n30861), .dinb(n291), .dout(n31171));
  jand g13149(.dina(n31171), .dinb(n31170), .dout(n31172));
  jor  g13150(.dina(n31172), .dinb(n30862), .dout(n31173));
  jxor g13151(.dina(n30856), .dinb(n284), .dout(n31174));
  jand g13152(.dina(n31174), .dinb(n31173), .dout(n31175));
  jor  g13153(.dina(n31175), .dinb(n30857), .dout(n31176));
  jxor g13154(.dina(n30851), .dinb(n285), .dout(n31177));
  jand g13155(.dina(n31177), .dinb(n31176), .dout(n31178));
  jor  g13156(.dina(n31178), .dinb(n30852), .dout(n31179));
  jxor g13157(.dina(n30846), .dinb(n281), .dout(n31180));
  jand g13158(.dina(n31180), .dinb(n31179), .dout(n31181));
  jor  g13159(.dina(n31181), .dinb(n30847), .dout(n31182));
  jxor g13160(.dina(n30841), .dinb(n282), .dout(n31183));
  jand g13161(.dina(n31183), .dinb(n31182), .dout(n31184));
  jor  g13162(.dina(n31184), .dinb(n30842), .dout(n31185));
  jxor g13163(.dina(n30836), .dinb(n397), .dout(n31186));
  jand g13164(.dina(n31186), .dinb(n31185), .dout(n31187));
  jor  g13165(.dina(n31187), .dinb(n30837), .dout(n31188));
  jor  g13166(.dina(n31188), .dinb(n30831), .dout(n31189));
  jand g13167(.dina(n31189), .dinb(n30830), .dout(n31190));
  jand g13168(.dina(n31190), .dinb(n9869), .dout(n31191));
  jnot g13169(.din(n31191), .dout(n31192));
  jand g13170(.dina(n31192), .dinb(n30828), .dout(n31193));
  jand g13171(.dina(n30831), .dinb(n9869), .dout(n31194));
  jand g13172(.dina(n31194), .dinb(n31188), .dout(n31195));
  jor  g13173(.dina(n31195), .dinb(n31193), .dout(n31196));
  jand g13174(.dina(n31196), .dinb(n9869), .dout(n31197));
  jnot g13175(.din(n31197), .dout(n31198));
  jand g13176(.dina(n31192), .dinb(n30836), .dout(n31199));
  jxor g13177(.dina(n31186), .dinb(n31185), .dout(n31200));
  jand g13178(.dina(n31200), .dinb(n31191), .dout(n31201));
  jor  g13179(.dina(n31201), .dinb(n31199), .dout(n31202));
  jand g13180(.dina(n31202), .dinb(n513), .dout(n31203));
  jnot g13181(.din(n31203), .dout(n31204));
  jand g13182(.dina(n31192), .dinb(n30841), .dout(n31205));
  jxor g13183(.dina(n31183), .dinb(n31182), .dout(n31206));
  jand g13184(.dina(n31206), .dinb(n31191), .dout(n31207));
  jor  g13185(.dina(n31207), .dinb(n31205), .dout(n31208));
  jand g13186(.dina(n31208), .dinb(n397), .dout(n31209));
  jnot g13187(.din(n31209), .dout(n31210));
  jand g13188(.dina(n31192), .dinb(n30846), .dout(n31211));
  jxor g13189(.dina(n31180), .dinb(n31179), .dout(n31212));
  jand g13190(.dina(n31212), .dinb(n31191), .dout(n31213));
  jor  g13191(.dina(n31213), .dinb(n31211), .dout(n31214));
  jand g13192(.dina(n31214), .dinb(n282), .dout(n31215));
  jnot g13193(.din(n31215), .dout(n31216));
  jand g13194(.dina(n31192), .dinb(n30851), .dout(n31217));
  jxor g13195(.dina(n31177), .dinb(n31176), .dout(n31218));
  jand g13196(.dina(n31218), .dinb(n31191), .dout(n31219));
  jor  g13197(.dina(n31219), .dinb(n31217), .dout(n31220));
  jand g13198(.dina(n31220), .dinb(n281), .dout(n31221));
  jnot g13199(.din(n31221), .dout(n31222));
  jand g13200(.dina(n31192), .dinb(n30856), .dout(n31223));
  jxor g13201(.dina(n31174), .dinb(n31173), .dout(n31224));
  jand g13202(.dina(n31224), .dinb(n31191), .dout(n31225));
  jor  g13203(.dina(n31225), .dinb(n31223), .dout(n31226));
  jand g13204(.dina(n31226), .dinb(n285), .dout(n31227));
  jnot g13205(.din(n31227), .dout(n31228));
  jand g13206(.dina(n31192), .dinb(n30861), .dout(n31229));
  jxor g13207(.dina(n31171), .dinb(n31170), .dout(n31230));
  jand g13208(.dina(n31230), .dinb(n31191), .dout(n31231));
  jor  g13209(.dina(n31231), .dinb(n31229), .dout(n31232));
  jand g13210(.dina(n31232), .dinb(n284), .dout(n31233));
  jnot g13211(.din(n31233), .dout(n31234));
  jand g13212(.dina(n31192), .dinb(n30866), .dout(n31235));
  jxor g13213(.dina(n31168), .dinb(n31167), .dout(n31236));
  jand g13214(.dina(n31236), .dinb(n31191), .dout(n31237));
  jor  g13215(.dina(n31237), .dinb(n31235), .dout(n31238));
  jand g13216(.dina(n31238), .dinb(n291), .dout(n31239));
  jnot g13217(.din(n31239), .dout(n31240));
  jand g13218(.dina(n31192), .dinb(n30871), .dout(n31241));
  jxor g13219(.dina(n31165), .dinb(n31164), .dout(n31242));
  jand g13220(.dina(n31242), .dinb(n31191), .dout(n31243));
  jor  g13221(.dina(n31243), .dinb(n31241), .dout(n31244));
  jand g13222(.dina(n31244), .dinb(n290), .dout(n31245));
  jnot g13223(.din(n31245), .dout(n31246));
  jand g13224(.dina(n31192), .dinb(n30876), .dout(n31247));
  jxor g13225(.dina(n31162), .dinb(n31161), .dout(n31248));
  jand g13226(.dina(n31248), .dinb(n31191), .dout(n31249));
  jor  g13227(.dina(n31249), .dinb(n31247), .dout(n31250));
  jand g13228(.dina(n31250), .dinb(n294), .dout(n31251));
  jnot g13229(.din(n31251), .dout(n31252));
  jand g13230(.dina(n31192), .dinb(n30881), .dout(n31253));
  jxor g13231(.dina(n31159), .dinb(n31158), .dout(n31254));
  jand g13232(.dina(n31254), .dinb(n31191), .dout(n31255));
  jor  g13233(.dina(n31255), .dinb(n31253), .dout(n31256));
  jand g13234(.dina(n31256), .dinb(n293), .dout(n31257));
  jnot g13235(.din(n31257), .dout(n31258));
  jand g13236(.dina(n31192), .dinb(n30886), .dout(n31259));
  jxor g13237(.dina(n31156), .dinb(n31155), .dout(n31260));
  jand g13238(.dina(n31260), .dinb(n31191), .dout(n31261));
  jor  g13239(.dina(n31261), .dinb(n31259), .dout(n31262));
  jand g13240(.dina(n31262), .dinb(n301), .dout(n31263));
  jnot g13241(.din(n31263), .dout(n31264));
  jand g13242(.dina(n31192), .dinb(n30891), .dout(n31265));
  jxor g13243(.dina(n31153), .dinb(n31152), .dout(n31266));
  jand g13244(.dina(n31266), .dinb(n31191), .dout(n31267));
  jor  g13245(.dina(n31267), .dinb(n31265), .dout(n31268));
  jand g13246(.dina(n31268), .dinb(n298), .dout(n31269));
  jnot g13247(.din(n31269), .dout(n31270));
  jand g13248(.dina(n31192), .dinb(n30896), .dout(n31271));
  jxor g13249(.dina(n31150), .dinb(n31149), .dout(n31272));
  jand g13250(.dina(n31272), .dinb(n31191), .dout(n31273));
  jor  g13251(.dina(n31273), .dinb(n31271), .dout(n31274));
  jand g13252(.dina(n31274), .dinb(n297), .dout(n31275));
  jnot g13253(.din(n31275), .dout(n31276));
  jand g13254(.dina(n31192), .dinb(n30901), .dout(n31277));
  jxor g13255(.dina(n31147), .dinb(n31146), .dout(n31278));
  jand g13256(.dina(n31278), .dinb(n31191), .dout(n31279));
  jor  g13257(.dina(n31279), .dinb(n31277), .dout(n31280));
  jand g13258(.dina(n31280), .dinb(n300), .dout(n31281));
  jnot g13259(.din(n31281), .dout(n31282));
  jand g13260(.dina(n31192), .dinb(n30906), .dout(n31283));
  jxor g13261(.dina(n31144), .dinb(n31143), .dout(n31284));
  jand g13262(.dina(n31284), .dinb(n31191), .dout(n31285));
  jor  g13263(.dina(n31285), .dinb(n31283), .dout(n31286));
  jand g13264(.dina(n31286), .dinb(n424), .dout(n31287));
  jnot g13265(.din(n31287), .dout(n31288));
  jand g13266(.dina(n31192), .dinb(n30911), .dout(n31289));
  jxor g13267(.dina(n31141), .dinb(n31140), .dout(n31290));
  jand g13268(.dina(n31290), .dinb(n31191), .dout(n31291));
  jor  g13269(.dina(n31291), .dinb(n31289), .dout(n31292));
  jand g13270(.dina(n31292), .dinb(n427), .dout(n31293));
  jnot g13271(.din(n31293), .dout(n31294));
  jand g13272(.dina(n31192), .dinb(n30916), .dout(n31295));
  jxor g13273(.dina(n31138), .dinb(n31137), .dout(n31296));
  jand g13274(.dina(n31296), .dinb(n31191), .dout(n31297));
  jor  g13275(.dina(n31297), .dinb(n31295), .dout(n31298));
  jand g13276(.dina(n31298), .dinb(n426), .dout(n31299));
  jnot g13277(.din(n31299), .dout(n31300));
  jand g13278(.dina(n31192), .dinb(n30921), .dout(n31301));
  jxor g13279(.dina(n31135), .dinb(n31134), .dout(n31302));
  jand g13280(.dina(n31302), .dinb(n31191), .dout(n31303));
  jor  g13281(.dina(n31303), .dinb(n31301), .dout(n31304));
  jand g13282(.dina(n31304), .dinb(n410), .dout(n31305));
  jnot g13283(.din(n31305), .dout(n31306));
  jand g13284(.dina(n31192), .dinb(n30926), .dout(n31307));
  jxor g13285(.dina(n31132), .dinb(n31131), .dout(n31308));
  jand g13286(.dina(n31308), .dinb(n31191), .dout(n31309));
  jor  g13287(.dina(n31309), .dinb(n31307), .dout(n31310));
  jand g13288(.dina(n31310), .dinb(n409), .dout(n31311));
  jnot g13289(.din(n31311), .dout(n31312));
  jand g13290(.dina(n31192), .dinb(n30931), .dout(n31313));
  jxor g13291(.dina(n31129), .dinb(n31128), .dout(n31314));
  jand g13292(.dina(n31314), .dinb(n31191), .dout(n31315));
  jor  g13293(.dina(n31315), .dinb(n31313), .dout(n31316));
  jand g13294(.dina(n31316), .dinb(n413), .dout(n31317));
  jnot g13295(.din(n31317), .dout(n31318));
  jand g13296(.dina(n31192), .dinb(n30936), .dout(n31319));
  jxor g13297(.dina(n31126), .dinb(n31125), .dout(n31320));
  jand g13298(.dina(n31320), .dinb(n31191), .dout(n31321));
  jor  g13299(.dina(n31321), .dinb(n31319), .dout(n31322));
  jand g13300(.dina(n31322), .dinb(n412), .dout(n31323));
  jnot g13301(.din(n31323), .dout(n31324));
  jand g13302(.dina(n31192), .dinb(n30941), .dout(n31325));
  jxor g13303(.dina(n31123), .dinb(n31122), .dout(n31326));
  jand g13304(.dina(n31326), .dinb(n31191), .dout(n31327));
  jor  g13305(.dina(n31327), .dinb(n31325), .dout(n31328));
  jand g13306(.dina(n31328), .dinb(n406), .dout(n31329));
  jnot g13307(.din(n31329), .dout(n31330));
  jand g13308(.dina(n31192), .dinb(n30946), .dout(n31331));
  jxor g13309(.dina(n31120), .dinb(n31119), .dout(n31332));
  jand g13310(.dina(n31332), .dinb(n31191), .dout(n31333));
  jor  g13311(.dina(n31333), .dinb(n31331), .dout(n31334));
  jand g13312(.dina(n31334), .dinb(n405), .dout(n31335));
  jnot g13313(.din(n31335), .dout(n31336));
  jand g13314(.dina(n31192), .dinb(n30951), .dout(n31337));
  jxor g13315(.dina(n31117), .dinb(n31116), .dout(n31338));
  jand g13316(.dina(n31338), .dinb(n31191), .dout(n31339));
  jor  g13317(.dina(n31339), .dinb(n31337), .dout(n31340));
  jand g13318(.dina(n31340), .dinb(n2714), .dout(n31341));
  jnot g13319(.din(n31341), .dout(n31342));
  jand g13320(.dina(n31192), .dinb(n30956), .dout(n31343));
  jxor g13321(.dina(n31114), .dinb(n31113), .dout(n31344));
  jand g13322(.dina(n31344), .dinb(n31191), .dout(n31345));
  jor  g13323(.dina(n31345), .dinb(n31343), .dout(n31346));
  jand g13324(.dina(n31346), .dinb(n2547), .dout(n31347));
  jnot g13325(.din(n31347), .dout(n31348));
  jand g13326(.dina(n31192), .dinb(n30961), .dout(n31349));
  jxor g13327(.dina(n31111), .dinb(n31110), .dout(n31350));
  jand g13328(.dina(n31350), .dinb(n31191), .dout(n31351));
  jor  g13329(.dina(n31351), .dinb(n31349), .dout(n31352));
  jand g13330(.dina(n31352), .dinb(n417), .dout(n31353));
  jnot g13331(.din(n31353), .dout(n31354));
  jand g13332(.dina(n31192), .dinb(n30966), .dout(n31355));
  jxor g13333(.dina(n31108), .dinb(n31107), .dout(n31356));
  jand g13334(.dina(n31356), .dinb(n31191), .dout(n31357));
  jor  g13335(.dina(n31357), .dinb(n31355), .dout(n31358));
  jand g13336(.dina(n31358), .dinb(n416), .dout(n31359));
  jnot g13337(.din(n31359), .dout(n31360));
  jand g13338(.dina(n31192), .dinb(n30971), .dout(n31361));
  jxor g13339(.dina(n31105), .dinb(n31104), .dout(n31362));
  jand g13340(.dina(n31362), .dinb(n31191), .dout(n31363));
  jor  g13341(.dina(n31363), .dinb(n31361), .dout(n31364));
  jand g13342(.dina(n31364), .dinb(n422), .dout(n31365));
  jnot g13343(.din(n31365), .dout(n31366));
  jand g13344(.dina(n31192), .dinb(n30976), .dout(n31367));
  jxor g13345(.dina(n31102), .dinb(n31101), .dout(n31368));
  jand g13346(.dina(n31368), .dinb(n31191), .dout(n31369));
  jor  g13347(.dina(n31369), .dinb(n31367), .dout(n31370));
  jand g13348(.dina(n31370), .dinb(n421), .dout(n31371));
  jnot g13349(.din(n31371), .dout(n31372));
  jand g13350(.dina(n31192), .dinb(n30981), .dout(n31373));
  jxor g13351(.dina(n31099), .dinb(n31098), .dout(n31374));
  jand g13352(.dina(n31374), .dinb(n31191), .dout(n31375));
  jor  g13353(.dina(n31375), .dinb(n31373), .dout(n31376));
  jand g13354(.dina(n31376), .dinb(n433), .dout(n31377));
  jnot g13355(.din(n31377), .dout(n31378));
  jand g13356(.dina(n31192), .dinb(n30986), .dout(n31379));
  jxor g13357(.dina(n31096), .dinb(n31095), .dout(n31380));
  jand g13358(.dina(n31380), .dinb(n31191), .dout(n31381));
  jor  g13359(.dina(n31381), .dinb(n31379), .dout(n31382));
  jand g13360(.dina(n31382), .dinb(n432), .dout(n31383));
  jnot g13361(.din(n31383), .dout(n31384));
  jand g13362(.dina(n31192), .dinb(n30991), .dout(n31385));
  jxor g13363(.dina(n31093), .dinb(n31092), .dout(n31386));
  jand g13364(.dina(n31386), .dinb(n31191), .dout(n31387));
  jor  g13365(.dina(n31387), .dinb(n31385), .dout(n31388));
  jand g13366(.dina(n31388), .dinb(n436), .dout(n31389));
  jnot g13367(.din(n31389), .dout(n31390));
  jand g13368(.dina(n31192), .dinb(n30996), .dout(n31391));
  jxor g13369(.dina(n31090), .dinb(n31089), .dout(n31392));
  jand g13370(.dina(n31392), .dinb(n31191), .dout(n31393));
  jor  g13371(.dina(n31393), .dinb(n31391), .dout(n31394));
  jand g13372(.dina(n31394), .dinb(n435), .dout(n31395));
  jnot g13373(.din(n31395), .dout(n31396));
  jand g13374(.dina(n31192), .dinb(n31001), .dout(n31397));
  jxor g13375(.dina(n31087), .dinb(n31086), .dout(n31398));
  jand g13376(.dina(n31398), .dinb(n31191), .dout(n31399));
  jor  g13377(.dina(n31399), .dinb(n31397), .dout(n31400));
  jand g13378(.dina(n31400), .dinb(n440), .dout(n31401));
  jnot g13379(.din(n31401), .dout(n31402));
  jand g13380(.dina(n31192), .dinb(n31006), .dout(n31403));
  jxor g13381(.dina(n31084), .dinb(n31083), .dout(n31404));
  jand g13382(.dina(n31404), .dinb(n31191), .dout(n31405));
  jor  g13383(.dina(n31405), .dinb(n31403), .dout(n31406));
  jand g13384(.dina(n31406), .dinb(n439), .dout(n31407));
  jnot g13385(.din(n31407), .dout(n31408));
  jand g13386(.dina(n31192), .dinb(n31011), .dout(n31409));
  jxor g13387(.dina(n31081), .dinb(n31080), .dout(n31410));
  jand g13388(.dina(n31410), .dinb(n31191), .dout(n31411));
  jor  g13389(.dina(n31411), .dinb(n31409), .dout(n31412));
  jand g13390(.dina(n31412), .dinb(n325), .dout(n31413));
  jnot g13391(.din(n31413), .dout(n31414));
  jand g13392(.dina(n31192), .dinb(n31016), .dout(n31415));
  jxor g13393(.dina(n31078), .dinb(n31077), .dout(n31416));
  jand g13394(.dina(n31416), .dinb(n31191), .dout(n31417));
  jor  g13395(.dina(n31417), .dinb(n31415), .dout(n31418));
  jand g13396(.dina(n31418), .dinb(n324), .dout(n31419));
  jnot g13397(.din(n31419), .dout(n31420));
  jand g13398(.dina(n31192), .dinb(n31021), .dout(n31421));
  jxor g13399(.dina(n31075), .dinb(n31074), .dout(n31422));
  jand g13400(.dina(n31422), .dinb(n31191), .dout(n31423));
  jor  g13401(.dina(n31423), .dinb(n31421), .dout(n31424));
  jand g13402(.dina(n31424), .dinb(n323), .dout(n31425));
  jnot g13403(.din(n31425), .dout(n31426));
  jand g13404(.dina(n31192), .dinb(n31026), .dout(n31427));
  jxor g13405(.dina(n31072), .dinb(n31071), .dout(n31428));
  jand g13406(.dina(n31428), .dinb(n31191), .dout(n31429));
  jor  g13407(.dina(n31429), .dinb(n31427), .dout(n31430));
  jand g13408(.dina(n31430), .dinb(n335), .dout(n31431));
  jnot g13409(.din(n31431), .dout(n31432));
  jand g13410(.dina(n31192), .dinb(n31031), .dout(n31433));
  jxor g13411(.dina(n31069), .dinb(n31068), .dout(n31434));
  jand g13412(.dina(n31434), .dinb(n31191), .dout(n31435));
  jor  g13413(.dina(n31435), .dinb(n31433), .dout(n31436));
  jand g13414(.dina(n31436), .dinb(n334), .dout(n31437));
  jnot g13415(.din(n31437), .dout(n31438));
  jand g13416(.dina(n31192), .dinb(n31036), .dout(n31439));
  jxor g13417(.dina(n31066), .dinb(n31065), .dout(n31440));
  jand g13418(.dina(n31440), .dinb(n31191), .dout(n31441));
  jor  g13419(.dina(n31441), .dinb(n31439), .dout(n31442));
  jand g13420(.dina(n31442), .dinb(n338), .dout(n31443));
  jnot g13421(.din(n31443), .dout(n31444));
  jand g13422(.dina(n31192), .dinb(n31041), .dout(n31445));
  jxor g13423(.dina(n31063), .dinb(n31062), .dout(n31446));
  jand g13424(.dina(n31446), .dinb(n31191), .dout(n31447));
  jor  g13425(.dina(n31447), .dinb(n31445), .dout(n31448));
  jand g13426(.dina(n31448), .dinb(n337), .dout(n31449));
  jnot g13427(.din(n31449), .dout(n31450));
  jnot g13428(.din(n31046), .dout(n31451));
  jor  g13429(.dina(n31191), .dinb(n31451), .dout(n31452));
  jxor g13430(.dina(n31060), .dinb(n31059), .dout(n31453));
  jnot g13431(.din(n31453), .dout(n31454));
  jor  g13432(.dina(n31454), .dinb(n31192), .dout(n31455));
  jand g13433(.dina(n31455), .dinb(n31452), .dout(n31456));
  jnot g13434(.din(n31456), .dout(n31457));
  jand g13435(.dina(n31457), .dinb(n344), .dout(n31458));
  jnot g13436(.din(n31458), .dout(n31459));
  jor  g13437(.dina(n31191), .dinb(n31056), .dout(n31460));
  jxor g13438(.dina(n31057), .dinb(n10102), .dout(n31461));
  jand g13439(.dina(n31461), .dinb(n31191), .dout(n31462));
  jnot g13440(.din(n31462), .dout(n31463));
  jand g13441(.dina(n31463), .dinb(n31460), .dout(n31464));
  jnot g13442(.din(n31464), .dout(n31465));
  jand g13443(.dina(n31465), .dinb(n348), .dout(n31466));
  jnot g13444(.din(n31466), .dout(n31467));
  jnot g13445(.din(n10460), .dout(n31468));
  jnot g13446(.din(n30831), .dout(n31469));
  jnot g13447(.din(n30837), .dout(n31470));
  jnot g13448(.din(n30842), .dout(n31471));
  jnot g13449(.din(n30847), .dout(n31472));
  jnot g13450(.din(n30852), .dout(n31473));
  jnot g13451(.din(n30857), .dout(n31474));
  jnot g13452(.din(n30862), .dout(n31475));
  jnot g13453(.din(n30867), .dout(n31476));
  jnot g13454(.din(n30872), .dout(n31477));
  jnot g13455(.din(n30877), .dout(n31478));
  jnot g13456(.din(n30882), .dout(n31479));
  jnot g13457(.din(n30887), .dout(n31480));
  jnot g13458(.din(n30892), .dout(n31481));
  jnot g13459(.din(n30897), .dout(n31482));
  jnot g13460(.din(n30902), .dout(n31483));
  jnot g13461(.din(n30907), .dout(n31484));
  jnot g13462(.din(n30912), .dout(n31485));
  jnot g13463(.din(n30917), .dout(n31486));
  jnot g13464(.din(n30922), .dout(n31487));
  jnot g13465(.din(n30927), .dout(n31488));
  jnot g13466(.din(n30932), .dout(n31489));
  jnot g13467(.din(n30937), .dout(n31490));
  jnot g13468(.din(n30942), .dout(n31491));
  jnot g13469(.din(n30947), .dout(n31492));
  jnot g13470(.din(n30952), .dout(n31493));
  jnot g13471(.din(n30957), .dout(n31494));
  jnot g13472(.din(n30962), .dout(n31495));
  jnot g13473(.din(n30967), .dout(n31496));
  jnot g13474(.din(n30972), .dout(n31497));
  jnot g13475(.din(n30977), .dout(n31498));
  jnot g13476(.din(n30982), .dout(n31499));
  jnot g13477(.din(n30987), .dout(n31500));
  jnot g13478(.din(n30992), .dout(n31501));
  jnot g13479(.din(n30997), .dout(n31502));
  jnot g13480(.din(n31002), .dout(n31503));
  jnot g13481(.din(n31007), .dout(n31504));
  jnot g13482(.din(n31012), .dout(n31505));
  jnot g13483(.din(n31017), .dout(n31506));
  jnot g13484(.din(n31022), .dout(n31507));
  jnot g13485(.din(n31027), .dout(n31508));
  jnot g13486(.din(n31032), .dout(n31509));
  jnot g13487(.din(n31037), .dout(n31510));
  jnot g13488(.din(n31042), .dout(n31511));
  jnot g13489(.din(n31047), .dout(n31512));
  jnot g13490(.din(n31053), .dout(n31513));
  jxor g13491(.dina(n31056), .dinb(n258), .dout(n31514));
  jor  g13492(.dina(n31514), .dinb(n10101), .dout(n31515));
  jand g13493(.dina(n31515), .dinb(n31513), .dout(n31516));
  jnot g13494(.din(n31060), .dout(n31517));
  jor  g13495(.dina(n31517), .dinb(n31516), .dout(n31518));
  jand g13496(.dina(n31518), .dinb(n31512), .dout(n31519));
  jnot g13497(.din(n31063), .dout(n31520));
  jor  g13498(.dina(n31520), .dinb(n31519), .dout(n31521));
  jand g13499(.dina(n31521), .dinb(n31511), .dout(n31522));
  jnot g13500(.din(n31066), .dout(n31523));
  jor  g13501(.dina(n31523), .dinb(n31522), .dout(n31524));
  jand g13502(.dina(n31524), .dinb(n31510), .dout(n31525));
  jnot g13503(.din(n31069), .dout(n31526));
  jor  g13504(.dina(n31526), .dinb(n31525), .dout(n31527));
  jand g13505(.dina(n31527), .dinb(n31509), .dout(n31528));
  jnot g13506(.din(n31072), .dout(n31529));
  jor  g13507(.dina(n31529), .dinb(n31528), .dout(n31530));
  jand g13508(.dina(n31530), .dinb(n31508), .dout(n31531));
  jnot g13509(.din(n31075), .dout(n31532));
  jor  g13510(.dina(n31532), .dinb(n31531), .dout(n31533));
  jand g13511(.dina(n31533), .dinb(n31507), .dout(n31534));
  jnot g13512(.din(n31078), .dout(n31535));
  jor  g13513(.dina(n31535), .dinb(n31534), .dout(n31536));
  jand g13514(.dina(n31536), .dinb(n31506), .dout(n31537));
  jnot g13515(.din(n31081), .dout(n31538));
  jor  g13516(.dina(n31538), .dinb(n31537), .dout(n31539));
  jand g13517(.dina(n31539), .dinb(n31505), .dout(n31540));
  jnot g13518(.din(n31084), .dout(n31541));
  jor  g13519(.dina(n31541), .dinb(n31540), .dout(n31542));
  jand g13520(.dina(n31542), .dinb(n31504), .dout(n31543));
  jnot g13521(.din(n31087), .dout(n31544));
  jor  g13522(.dina(n31544), .dinb(n31543), .dout(n31545));
  jand g13523(.dina(n31545), .dinb(n31503), .dout(n31546));
  jnot g13524(.din(n31090), .dout(n31547));
  jor  g13525(.dina(n31547), .dinb(n31546), .dout(n31548));
  jand g13526(.dina(n31548), .dinb(n31502), .dout(n31549));
  jnot g13527(.din(n31093), .dout(n31550));
  jor  g13528(.dina(n31550), .dinb(n31549), .dout(n31551));
  jand g13529(.dina(n31551), .dinb(n31501), .dout(n31552));
  jnot g13530(.din(n31096), .dout(n31553));
  jor  g13531(.dina(n31553), .dinb(n31552), .dout(n31554));
  jand g13532(.dina(n31554), .dinb(n31500), .dout(n31555));
  jnot g13533(.din(n31099), .dout(n31556));
  jor  g13534(.dina(n31556), .dinb(n31555), .dout(n31557));
  jand g13535(.dina(n31557), .dinb(n31499), .dout(n31558));
  jnot g13536(.din(n31102), .dout(n31559));
  jor  g13537(.dina(n31559), .dinb(n31558), .dout(n31560));
  jand g13538(.dina(n31560), .dinb(n31498), .dout(n31561));
  jnot g13539(.din(n31105), .dout(n31562));
  jor  g13540(.dina(n31562), .dinb(n31561), .dout(n31563));
  jand g13541(.dina(n31563), .dinb(n31497), .dout(n31564));
  jnot g13542(.din(n31108), .dout(n31565));
  jor  g13543(.dina(n31565), .dinb(n31564), .dout(n31566));
  jand g13544(.dina(n31566), .dinb(n31496), .dout(n31567));
  jnot g13545(.din(n31111), .dout(n31568));
  jor  g13546(.dina(n31568), .dinb(n31567), .dout(n31569));
  jand g13547(.dina(n31569), .dinb(n31495), .dout(n31570));
  jnot g13548(.din(n31114), .dout(n31571));
  jor  g13549(.dina(n31571), .dinb(n31570), .dout(n31572));
  jand g13550(.dina(n31572), .dinb(n31494), .dout(n31573));
  jnot g13551(.din(n31117), .dout(n31574));
  jor  g13552(.dina(n31574), .dinb(n31573), .dout(n31575));
  jand g13553(.dina(n31575), .dinb(n31493), .dout(n31576));
  jnot g13554(.din(n31120), .dout(n31577));
  jor  g13555(.dina(n31577), .dinb(n31576), .dout(n31578));
  jand g13556(.dina(n31578), .dinb(n31492), .dout(n31579));
  jnot g13557(.din(n31123), .dout(n31580));
  jor  g13558(.dina(n31580), .dinb(n31579), .dout(n31581));
  jand g13559(.dina(n31581), .dinb(n31491), .dout(n31582));
  jnot g13560(.din(n31126), .dout(n31583));
  jor  g13561(.dina(n31583), .dinb(n31582), .dout(n31584));
  jand g13562(.dina(n31584), .dinb(n31490), .dout(n31585));
  jnot g13563(.din(n31129), .dout(n31586));
  jor  g13564(.dina(n31586), .dinb(n31585), .dout(n31587));
  jand g13565(.dina(n31587), .dinb(n31489), .dout(n31588));
  jnot g13566(.din(n31132), .dout(n31589));
  jor  g13567(.dina(n31589), .dinb(n31588), .dout(n31590));
  jand g13568(.dina(n31590), .dinb(n31488), .dout(n31591));
  jnot g13569(.din(n31135), .dout(n31592));
  jor  g13570(.dina(n31592), .dinb(n31591), .dout(n31593));
  jand g13571(.dina(n31593), .dinb(n31487), .dout(n31594));
  jnot g13572(.din(n31138), .dout(n31595));
  jor  g13573(.dina(n31595), .dinb(n31594), .dout(n31596));
  jand g13574(.dina(n31596), .dinb(n31486), .dout(n31597));
  jnot g13575(.din(n31141), .dout(n31598));
  jor  g13576(.dina(n31598), .dinb(n31597), .dout(n31599));
  jand g13577(.dina(n31599), .dinb(n31485), .dout(n31600));
  jnot g13578(.din(n31144), .dout(n31601));
  jor  g13579(.dina(n31601), .dinb(n31600), .dout(n31602));
  jand g13580(.dina(n31602), .dinb(n31484), .dout(n31603));
  jnot g13581(.din(n31147), .dout(n31604));
  jor  g13582(.dina(n31604), .dinb(n31603), .dout(n31605));
  jand g13583(.dina(n31605), .dinb(n31483), .dout(n31606));
  jnot g13584(.din(n31150), .dout(n31607));
  jor  g13585(.dina(n31607), .dinb(n31606), .dout(n31608));
  jand g13586(.dina(n31608), .dinb(n31482), .dout(n31609));
  jnot g13587(.din(n31153), .dout(n31610));
  jor  g13588(.dina(n31610), .dinb(n31609), .dout(n31611));
  jand g13589(.dina(n31611), .dinb(n31481), .dout(n31612));
  jnot g13590(.din(n31156), .dout(n31613));
  jor  g13591(.dina(n31613), .dinb(n31612), .dout(n31614));
  jand g13592(.dina(n31614), .dinb(n31480), .dout(n31615));
  jnot g13593(.din(n31159), .dout(n31616));
  jor  g13594(.dina(n31616), .dinb(n31615), .dout(n31617));
  jand g13595(.dina(n31617), .dinb(n31479), .dout(n31618));
  jnot g13596(.din(n31162), .dout(n31619));
  jor  g13597(.dina(n31619), .dinb(n31618), .dout(n31620));
  jand g13598(.dina(n31620), .dinb(n31478), .dout(n31621));
  jnot g13599(.din(n31165), .dout(n31622));
  jor  g13600(.dina(n31622), .dinb(n31621), .dout(n31623));
  jand g13601(.dina(n31623), .dinb(n31477), .dout(n31624));
  jnot g13602(.din(n31168), .dout(n31625));
  jor  g13603(.dina(n31625), .dinb(n31624), .dout(n31626));
  jand g13604(.dina(n31626), .dinb(n31476), .dout(n31627));
  jnot g13605(.din(n31171), .dout(n31628));
  jor  g13606(.dina(n31628), .dinb(n31627), .dout(n31629));
  jand g13607(.dina(n31629), .dinb(n31475), .dout(n31630));
  jnot g13608(.din(n31174), .dout(n31631));
  jor  g13609(.dina(n31631), .dinb(n31630), .dout(n31632));
  jand g13610(.dina(n31632), .dinb(n31474), .dout(n31633));
  jnot g13611(.din(n31177), .dout(n31634));
  jor  g13612(.dina(n31634), .dinb(n31633), .dout(n31635));
  jand g13613(.dina(n31635), .dinb(n31473), .dout(n31636));
  jnot g13614(.din(n31180), .dout(n31637));
  jor  g13615(.dina(n31637), .dinb(n31636), .dout(n31638));
  jand g13616(.dina(n31638), .dinb(n31472), .dout(n31639));
  jnot g13617(.din(n31183), .dout(n31640));
  jor  g13618(.dina(n31640), .dinb(n31639), .dout(n31641));
  jand g13619(.dina(n31641), .dinb(n31471), .dout(n31642));
  jnot g13620(.din(n31186), .dout(n31643));
  jor  g13621(.dina(n31643), .dinb(n31642), .dout(n31644));
  jand g13622(.dina(n31644), .dinb(n31470), .dout(n31645));
  jand g13623(.dina(n31645), .dinb(n31469), .dout(n31646));
  jor  g13624(.dina(n31646), .dinb(n30829), .dout(n31647));
  jor  g13625(.dina(n31647), .dinb(n31468), .dout(n31648));
  jand g13626(.dina(n31648), .dinb(a18 ), .dout(n31649));
  jnot g13627(.din(n10463), .dout(n31650));
  jor  g13628(.dina(n31647), .dinb(n31650), .dout(n31651));
  jnot g13629(.din(n31651), .dout(n31652));
  jor  g13630(.dina(n31652), .dinb(n31649), .dout(n31653));
  jand g13631(.dina(n31653), .dinb(n258), .dout(n31654));
  jnot g13632(.din(n31654), .dout(n31655));
  jand g13633(.dina(n31190), .dinb(n10460), .dout(n31656));
  jor  g13634(.dina(n31656), .dinb(n10100), .dout(n31657));
  jand g13635(.dina(n31651), .dinb(n31657), .dout(n31658));
  jxor g13636(.dina(n31658), .dinb(n258), .dout(n31659));
  jor  g13637(.dina(n31659), .dinb(n10470), .dout(n31660));
  jand g13638(.dina(n31660), .dinb(n31655), .dout(n31661));
  jxor g13639(.dina(n31464), .dinb(b2 ), .dout(n31662));
  jnot g13640(.din(n31662), .dout(n31663));
  jor  g13641(.dina(n31663), .dinb(n31661), .dout(n31664));
  jand g13642(.dina(n31664), .dinb(n31467), .dout(n31665));
  jxor g13643(.dina(n31456), .dinb(b3 ), .dout(n31666));
  jnot g13644(.din(n31666), .dout(n31667));
  jor  g13645(.dina(n31667), .dinb(n31665), .dout(n31668));
  jand g13646(.dina(n31668), .dinb(n31459), .dout(n31669));
  jxor g13647(.dina(n31448), .dinb(n337), .dout(n31670));
  jnot g13648(.din(n31670), .dout(n31671));
  jor  g13649(.dina(n31671), .dinb(n31669), .dout(n31672));
  jand g13650(.dina(n31672), .dinb(n31450), .dout(n31673));
  jxor g13651(.dina(n31442), .dinb(n338), .dout(n31674));
  jnot g13652(.din(n31674), .dout(n31675));
  jor  g13653(.dina(n31675), .dinb(n31673), .dout(n31676));
  jand g13654(.dina(n31676), .dinb(n31444), .dout(n31677));
  jxor g13655(.dina(n31436), .dinb(n334), .dout(n31678));
  jnot g13656(.din(n31678), .dout(n31679));
  jor  g13657(.dina(n31679), .dinb(n31677), .dout(n31680));
  jand g13658(.dina(n31680), .dinb(n31438), .dout(n31681));
  jxor g13659(.dina(n31430), .dinb(n335), .dout(n31682));
  jnot g13660(.din(n31682), .dout(n31683));
  jor  g13661(.dina(n31683), .dinb(n31681), .dout(n31684));
  jand g13662(.dina(n31684), .dinb(n31432), .dout(n31685));
  jxor g13663(.dina(n31424), .dinb(n323), .dout(n31686));
  jnot g13664(.din(n31686), .dout(n31687));
  jor  g13665(.dina(n31687), .dinb(n31685), .dout(n31688));
  jand g13666(.dina(n31688), .dinb(n31426), .dout(n31689));
  jxor g13667(.dina(n31418), .dinb(n324), .dout(n31690));
  jnot g13668(.din(n31690), .dout(n31691));
  jor  g13669(.dina(n31691), .dinb(n31689), .dout(n31692));
  jand g13670(.dina(n31692), .dinb(n31420), .dout(n31693));
  jxor g13671(.dina(n31412), .dinb(n325), .dout(n31694));
  jnot g13672(.din(n31694), .dout(n31695));
  jor  g13673(.dina(n31695), .dinb(n31693), .dout(n31696));
  jand g13674(.dina(n31696), .dinb(n31414), .dout(n31697));
  jxor g13675(.dina(n31406), .dinb(n439), .dout(n31698));
  jnot g13676(.din(n31698), .dout(n31699));
  jor  g13677(.dina(n31699), .dinb(n31697), .dout(n31700));
  jand g13678(.dina(n31700), .dinb(n31408), .dout(n31701));
  jxor g13679(.dina(n31400), .dinb(n440), .dout(n31702));
  jnot g13680(.din(n31702), .dout(n31703));
  jor  g13681(.dina(n31703), .dinb(n31701), .dout(n31704));
  jand g13682(.dina(n31704), .dinb(n31402), .dout(n31705));
  jxor g13683(.dina(n31394), .dinb(n435), .dout(n31706));
  jnot g13684(.din(n31706), .dout(n31707));
  jor  g13685(.dina(n31707), .dinb(n31705), .dout(n31708));
  jand g13686(.dina(n31708), .dinb(n31396), .dout(n31709));
  jxor g13687(.dina(n31388), .dinb(n436), .dout(n31710));
  jnot g13688(.din(n31710), .dout(n31711));
  jor  g13689(.dina(n31711), .dinb(n31709), .dout(n31712));
  jand g13690(.dina(n31712), .dinb(n31390), .dout(n31713));
  jxor g13691(.dina(n31382), .dinb(n432), .dout(n31714));
  jnot g13692(.din(n31714), .dout(n31715));
  jor  g13693(.dina(n31715), .dinb(n31713), .dout(n31716));
  jand g13694(.dina(n31716), .dinb(n31384), .dout(n31717));
  jxor g13695(.dina(n31376), .dinb(n433), .dout(n31718));
  jnot g13696(.din(n31718), .dout(n31719));
  jor  g13697(.dina(n31719), .dinb(n31717), .dout(n31720));
  jand g13698(.dina(n31720), .dinb(n31378), .dout(n31721));
  jxor g13699(.dina(n31370), .dinb(n421), .dout(n31722));
  jnot g13700(.din(n31722), .dout(n31723));
  jor  g13701(.dina(n31723), .dinb(n31721), .dout(n31724));
  jand g13702(.dina(n31724), .dinb(n31372), .dout(n31725));
  jxor g13703(.dina(n31364), .dinb(n422), .dout(n31726));
  jnot g13704(.din(n31726), .dout(n31727));
  jor  g13705(.dina(n31727), .dinb(n31725), .dout(n31728));
  jand g13706(.dina(n31728), .dinb(n31366), .dout(n31729));
  jxor g13707(.dina(n31358), .dinb(n416), .dout(n31730));
  jnot g13708(.din(n31730), .dout(n31731));
  jor  g13709(.dina(n31731), .dinb(n31729), .dout(n31732));
  jand g13710(.dina(n31732), .dinb(n31360), .dout(n31733));
  jxor g13711(.dina(n31352), .dinb(n417), .dout(n31734));
  jnot g13712(.din(n31734), .dout(n31735));
  jor  g13713(.dina(n31735), .dinb(n31733), .dout(n31736));
  jand g13714(.dina(n31736), .dinb(n31354), .dout(n31737));
  jxor g13715(.dina(n31346), .dinb(n2547), .dout(n31738));
  jnot g13716(.din(n31738), .dout(n31739));
  jor  g13717(.dina(n31739), .dinb(n31737), .dout(n31740));
  jand g13718(.dina(n31740), .dinb(n31348), .dout(n31741));
  jxor g13719(.dina(n31340), .dinb(n2714), .dout(n31742));
  jnot g13720(.din(n31742), .dout(n31743));
  jor  g13721(.dina(n31743), .dinb(n31741), .dout(n31744));
  jand g13722(.dina(n31744), .dinb(n31342), .dout(n31745));
  jxor g13723(.dina(n31334), .dinb(n405), .dout(n31746));
  jnot g13724(.din(n31746), .dout(n31747));
  jor  g13725(.dina(n31747), .dinb(n31745), .dout(n31748));
  jand g13726(.dina(n31748), .dinb(n31336), .dout(n31749));
  jxor g13727(.dina(n31328), .dinb(n406), .dout(n31750));
  jnot g13728(.din(n31750), .dout(n31751));
  jor  g13729(.dina(n31751), .dinb(n31749), .dout(n31752));
  jand g13730(.dina(n31752), .dinb(n31330), .dout(n31753));
  jxor g13731(.dina(n31322), .dinb(n412), .dout(n31754));
  jnot g13732(.din(n31754), .dout(n31755));
  jor  g13733(.dina(n31755), .dinb(n31753), .dout(n31756));
  jand g13734(.dina(n31756), .dinb(n31324), .dout(n31757));
  jxor g13735(.dina(n31316), .dinb(n413), .dout(n31758));
  jnot g13736(.din(n31758), .dout(n31759));
  jor  g13737(.dina(n31759), .dinb(n31757), .dout(n31760));
  jand g13738(.dina(n31760), .dinb(n31318), .dout(n31761));
  jxor g13739(.dina(n31310), .dinb(n409), .dout(n31762));
  jnot g13740(.din(n31762), .dout(n31763));
  jor  g13741(.dina(n31763), .dinb(n31761), .dout(n31764));
  jand g13742(.dina(n31764), .dinb(n31312), .dout(n31765));
  jxor g13743(.dina(n31304), .dinb(n410), .dout(n31766));
  jnot g13744(.din(n31766), .dout(n31767));
  jor  g13745(.dina(n31767), .dinb(n31765), .dout(n31768));
  jand g13746(.dina(n31768), .dinb(n31306), .dout(n31769));
  jxor g13747(.dina(n31298), .dinb(n426), .dout(n31770));
  jnot g13748(.din(n31770), .dout(n31771));
  jor  g13749(.dina(n31771), .dinb(n31769), .dout(n31772));
  jand g13750(.dina(n31772), .dinb(n31300), .dout(n31773));
  jxor g13751(.dina(n31292), .dinb(n427), .dout(n31774));
  jnot g13752(.din(n31774), .dout(n31775));
  jor  g13753(.dina(n31775), .dinb(n31773), .dout(n31776));
  jand g13754(.dina(n31776), .dinb(n31294), .dout(n31777));
  jxor g13755(.dina(n31286), .dinb(n424), .dout(n31778));
  jnot g13756(.din(n31778), .dout(n31779));
  jor  g13757(.dina(n31779), .dinb(n31777), .dout(n31780));
  jand g13758(.dina(n31780), .dinb(n31288), .dout(n31781));
  jxor g13759(.dina(n31280), .dinb(n300), .dout(n31782));
  jnot g13760(.din(n31782), .dout(n31783));
  jor  g13761(.dina(n31783), .dinb(n31781), .dout(n31784));
  jand g13762(.dina(n31784), .dinb(n31282), .dout(n31785));
  jxor g13763(.dina(n31274), .dinb(n297), .dout(n31786));
  jnot g13764(.din(n31786), .dout(n31787));
  jor  g13765(.dina(n31787), .dinb(n31785), .dout(n31788));
  jand g13766(.dina(n31788), .dinb(n31276), .dout(n31789));
  jxor g13767(.dina(n31268), .dinb(n298), .dout(n31790));
  jnot g13768(.din(n31790), .dout(n31791));
  jor  g13769(.dina(n31791), .dinb(n31789), .dout(n31792));
  jand g13770(.dina(n31792), .dinb(n31270), .dout(n31793));
  jxor g13771(.dina(n31262), .dinb(n301), .dout(n31794));
  jnot g13772(.din(n31794), .dout(n31795));
  jor  g13773(.dina(n31795), .dinb(n31793), .dout(n31796));
  jand g13774(.dina(n31796), .dinb(n31264), .dout(n31797));
  jxor g13775(.dina(n31256), .dinb(n293), .dout(n31798));
  jnot g13776(.din(n31798), .dout(n31799));
  jor  g13777(.dina(n31799), .dinb(n31797), .dout(n31800));
  jand g13778(.dina(n31800), .dinb(n31258), .dout(n31801));
  jxor g13779(.dina(n31250), .dinb(n294), .dout(n31802));
  jnot g13780(.din(n31802), .dout(n31803));
  jor  g13781(.dina(n31803), .dinb(n31801), .dout(n31804));
  jand g13782(.dina(n31804), .dinb(n31252), .dout(n31805));
  jxor g13783(.dina(n31244), .dinb(n290), .dout(n31806));
  jnot g13784(.din(n31806), .dout(n31807));
  jor  g13785(.dina(n31807), .dinb(n31805), .dout(n31808));
  jand g13786(.dina(n31808), .dinb(n31246), .dout(n31809));
  jxor g13787(.dina(n31238), .dinb(n291), .dout(n31810));
  jnot g13788(.din(n31810), .dout(n31811));
  jor  g13789(.dina(n31811), .dinb(n31809), .dout(n31812));
  jand g13790(.dina(n31812), .dinb(n31240), .dout(n31813));
  jxor g13791(.dina(n31232), .dinb(n284), .dout(n31814));
  jnot g13792(.din(n31814), .dout(n31815));
  jor  g13793(.dina(n31815), .dinb(n31813), .dout(n31816));
  jand g13794(.dina(n31816), .dinb(n31234), .dout(n31817));
  jxor g13795(.dina(n31226), .dinb(n285), .dout(n31818));
  jnot g13796(.din(n31818), .dout(n31819));
  jor  g13797(.dina(n31819), .dinb(n31817), .dout(n31820));
  jand g13798(.dina(n31820), .dinb(n31228), .dout(n31821));
  jxor g13799(.dina(n31220), .dinb(n281), .dout(n31822));
  jnot g13800(.din(n31822), .dout(n31823));
  jor  g13801(.dina(n31823), .dinb(n31821), .dout(n31824));
  jand g13802(.dina(n31824), .dinb(n31222), .dout(n31825));
  jxor g13803(.dina(n31214), .dinb(n282), .dout(n31826));
  jnot g13804(.din(n31826), .dout(n31827));
  jor  g13805(.dina(n31827), .dinb(n31825), .dout(n31828));
  jand g13806(.dina(n31828), .dinb(n31216), .dout(n31829));
  jxor g13807(.dina(n31208), .dinb(n397), .dout(n31830));
  jnot g13808(.din(n31830), .dout(n31831));
  jor  g13809(.dina(n31831), .dinb(n31829), .dout(n31832));
  jand g13810(.dina(n31832), .dinb(n31210), .dout(n31833));
  jxor g13811(.dina(n31202), .dinb(n513), .dout(n31834));
  jnot g13812(.din(n31834), .dout(n31835));
  jor  g13813(.dina(n31835), .dinb(n31833), .dout(n31836));
  jand g13814(.dina(n31836), .dinb(n31204), .dout(n31837));
  jxor g13815(.dina(n31196), .dinb(b46 ), .dout(n31838));
  jor  g13816(.dina(n31838), .dinb(n31837), .dout(n31839));
  jor  g13817(.dina(n31839), .dinb(n10607), .dout(n31840));
  jand g13818(.dina(n31840), .dinb(n31198), .dout(n31841));
  jand g13819(.dina(n31841), .dinb(n31196), .dout(n31842));
  jnot g13820(.din(n31842), .dout(n31843));
  jxor g13821(.dina(n31658), .dinb(b1 ), .dout(n31844));
  jand g13822(.dina(n31844), .dinb(n10471), .dout(n31845));
  jor  g13823(.dina(n31845), .dinb(n31654), .dout(n31846));
  jand g13824(.dina(n31662), .dinb(n31846), .dout(n31847));
  jor  g13825(.dina(n31847), .dinb(n31466), .dout(n31848));
  jand g13826(.dina(n31666), .dinb(n31848), .dout(n31849));
  jor  g13827(.dina(n31849), .dinb(n31458), .dout(n31850));
  jand g13828(.dina(n31670), .dinb(n31850), .dout(n31851));
  jor  g13829(.dina(n31851), .dinb(n31449), .dout(n31852));
  jand g13830(.dina(n31674), .dinb(n31852), .dout(n31853));
  jor  g13831(.dina(n31853), .dinb(n31443), .dout(n31854));
  jand g13832(.dina(n31678), .dinb(n31854), .dout(n31855));
  jor  g13833(.dina(n31855), .dinb(n31437), .dout(n31856));
  jand g13834(.dina(n31682), .dinb(n31856), .dout(n31857));
  jor  g13835(.dina(n31857), .dinb(n31431), .dout(n31858));
  jand g13836(.dina(n31686), .dinb(n31858), .dout(n31859));
  jor  g13837(.dina(n31859), .dinb(n31425), .dout(n31860));
  jand g13838(.dina(n31690), .dinb(n31860), .dout(n31861));
  jor  g13839(.dina(n31861), .dinb(n31419), .dout(n31862));
  jand g13840(.dina(n31694), .dinb(n31862), .dout(n31863));
  jor  g13841(.dina(n31863), .dinb(n31413), .dout(n31864));
  jand g13842(.dina(n31698), .dinb(n31864), .dout(n31865));
  jor  g13843(.dina(n31865), .dinb(n31407), .dout(n31866));
  jand g13844(.dina(n31702), .dinb(n31866), .dout(n31867));
  jor  g13845(.dina(n31867), .dinb(n31401), .dout(n31868));
  jand g13846(.dina(n31706), .dinb(n31868), .dout(n31869));
  jor  g13847(.dina(n31869), .dinb(n31395), .dout(n31870));
  jand g13848(.dina(n31710), .dinb(n31870), .dout(n31871));
  jor  g13849(.dina(n31871), .dinb(n31389), .dout(n31872));
  jand g13850(.dina(n31714), .dinb(n31872), .dout(n31873));
  jor  g13851(.dina(n31873), .dinb(n31383), .dout(n31874));
  jand g13852(.dina(n31718), .dinb(n31874), .dout(n31875));
  jor  g13853(.dina(n31875), .dinb(n31377), .dout(n31876));
  jand g13854(.dina(n31722), .dinb(n31876), .dout(n31877));
  jor  g13855(.dina(n31877), .dinb(n31371), .dout(n31878));
  jand g13856(.dina(n31726), .dinb(n31878), .dout(n31879));
  jor  g13857(.dina(n31879), .dinb(n31365), .dout(n31880));
  jand g13858(.dina(n31730), .dinb(n31880), .dout(n31881));
  jor  g13859(.dina(n31881), .dinb(n31359), .dout(n31882));
  jand g13860(.dina(n31734), .dinb(n31882), .dout(n31883));
  jor  g13861(.dina(n31883), .dinb(n31353), .dout(n31884));
  jand g13862(.dina(n31738), .dinb(n31884), .dout(n31885));
  jor  g13863(.dina(n31885), .dinb(n31347), .dout(n31886));
  jand g13864(.dina(n31742), .dinb(n31886), .dout(n31887));
  jor  g13865(.dina(n31887), .dinb(n31341), .dout(n31888));
  jand g13866(.dina(n31746), .dinb(n31888), .dout(n31889));
  jor  g13867(.dina(n31889), .dinb(n31335), .dout(n31890));
  jand g13868(.dina(n31750), .dinb(n31890), .dout(n31891));
  jor  g13869(.dina(n31891), .dinb(n31329), .dout(n31892));
  jand g13870(.dina(n31754), .dinb(n31892), .dout(n31893));
  jor  g13871(.dina(n31893), .dinb(n31323), .dout(n31894));
  jand g13872(.dina(n31758), .dinb(n31894), .dout(n31895));
  jor  g13873(.dina(n31895), .dinb(n31317), .dout(n31896));
  jand g13874(.dina(n31762), .dinb(n31896), .dout(n31897));
  jor  g13875(.dina(n31897), .dinb(n31311), .dout(n31898));
  jand g13876(.dina(n31766), .dinb(n31898), .dout(n31899));
  jor  g13877(.dina(n31899), .dinb(n31305), .dout(n31900));
  jand g13878(.dina(n31770), .dinb(n31900), .dout(n31901));
  jor  g13879(.dina(n31901), .dinb(n31299), .dout(n31902));
  jand g13880(.dina(n31774), .dinb(n31902), .dout(n31903));
  jor  g13881(.dina(n31903), .dinb(n31293), .dout(n31904));
  jand g13882(.dina(n31778), .dinb(n31904), .dout(n31905));
  jor  g13883(.dina(n31905), .dinb(n31287), .dout(n31906));
  jand g13884(.dina(n31782), .dinb(n31906), .dout(n31907));
  jor  g13885(.dina(n31907), .dinb(n31281), .dout(n31908));
  jand g13886(.dina(n31786), .dinb(n31908), .dout(n31909));
  jor  g13887(.dina(n31909), .dinb(n31275), .dout(n31910));
  jand g13888(.dina(n31790), .dinb(n31910), .dout(n31911));
  jor  g13889(.dina(n31911), .dinb(n31269), .dout(n31912));
  jand g13890(.dina(n31794), .dinb(n31912), .dout(n31913));
  jor  g13891(.dina(n31913), .dinb(n31263), .dout(n31914));
  jand g13892(.dina(n31798), .dinb(n31914), .dout(n31915));
  jor  g13893(.dina(n31915), .dinb(n31257), .dout(n31916));
  jand g13894(.dina(n31802), .dinb(n31916), .dout(n31917));
  jor  g13895(.dina(n31917), .dinb(n31251), .dout(n31918));
  jand g13896(.dina(n31806), .dinb(n31918), .dout(n31919));
  jor  g13897(.dina(n31919), .dinb(n31245), .dout(n31920));
  jand g13898(.dina(n31810), .dinb(n31920), .dout(n31921));
  jor  g13899(.dina(n31921), .dinb(n31239), .dout(n31922));
  jand g13900(.dina(n31814), .dinb(n31922), .dout(n31923));
  jor  g13901(.dina(n31923), .dinb(n31233), .dout(n31924));
  jand g13902(.dina(n31818), .dinb(n31924), .dout(n31925));
  jor  g13903(.dina(n31925), .dinb(n31227), .dout(n31926));
  jand g13904(.dina(n31822), .dinb(n31926), .dout(n31927));
  jor  g13905(.dina(n31927), .dinb(n31221), .dout(n31928));
  jand g13906(.dina(n31826), .dinb(n31928), .dout(n31929));
  jor  g13907(.dina(n31929), .dinb(n31215), .dout(n31930));
  jand g13908(.dina(n31830), .dinb(n31930), .dout(n31931));
  jor  g13909(.dina(n31931), .dinb(n31209), .dout(n31932));
  jand g13910(.dina(n31834), .dinb(n31932), .dout(n31933));
  jor  g13911(.dina(n31933), .dinb(n31203), .dout(n31934));
  jnot g13912(.din(n31838), .dout(n31935));
  jand g13913(.dina(n31935), .dinb(n31934), .dout(n31936));
  jand g13914(.dina(n31837), .dinb(n514), .dout(n31937));
  jor  g13915(.dina(n31937), .dinb(n31198), .dout(n31938));
  jor  g13916(.dina(n31938), .dinb(n31936), .dout(n31939));
  jand g13917(.dina(n31939), .dinb(n31843), .dout(n31940));
  jnot g13918(.din(n31940), .dout(n31941));
  jand g13919(.dina(n31941), .dinb(n512), .dout(n31942));
  jnot g13920(.din(n31942), .dout(n31943));
  jnot g13921(.din(n9868), .dout(n31944));
  jand g13922(.dina(n31841), .dinb(n31202), .dout(n31945));
  jand g13923(.dina(n31936), .dinb(n512), .dout(n31946));
  jor  g13924(.dina(n31946), .dinb(n31197), .dout(n31947));
  jxor g13925(.dina(n31834), .dinb(n31932), .dout(n31948));
  jand g13926(.dina(n31948), .dinb(n31947), .dout(n31949));
  jor  g13927(.dina(n31949), .dinb(n31945), .dout(n31950));
  jand g13928(.dina(n31950), .dinb(n514), .dout(n31951));
  jnot g13929(.din(n31951), .dout(n31952));
  jand g13930(.dina(n31841), .dinb(n31208), .dout(n31953));
  jxor g13931(.dina(n31830), .dinb(n31930), .dout(n31954));
  jand g13932(.dina(n31954), .dinb(n31947), .dout(n31955));
  jor  g13933(.dina(n31955), .dinb(n31953), .dout(n31956));
  jand g13934(.dina(n31956), .dinb(n513), .dout(n31957));
  jnot g13935(.din(n31957), .dout(n31958));
  jand g13936(.dina(n31841), .dinb(n31214), .dout(n31959));
  jxor g13937(.dina(n31826), .dinb(n31928), .dout(n31960));
  jand g13938(.dina(n31960), .dinb(n31947), .dout(n31961));
  jor  g13939(.dina(n31961), .dinb(n31959), .dout(n31962));
  jand g13940(.dina(n31962), .dinb(n397), .dout(n31963));
  jnot g13941(.din(n31963), .dout(n31964));
  jand g13942(.dina(n31841), .dinb(n31220), .dout(n31965));
  jxor g13943(.dina(n31822), .dinb(n31926), .dout(n31966));
  jand g13944(.dina(n31966), .dinb(n31947), .dout(n31967));
  jor  g13945(.dina(n31967), .dinb(n31965), .dout(n31968));
  jand g13946(.dina(n31968), .dinb(n282), .dout(n31969));
  jnot g13947(.din(n31969), .dout(n31970));
  jand g13948(.dina(n31841), .dinb(n31226), .dout(n31971));
  jxor g13949(.dina(n31818), .dinb(n31924), .dout(n31972));
  jand g13950(.dina(n31972), .dinb(n31947), .dout(n31973));
  jor  g13951(.dina(n31973), .dinb(n31971), .dout(n31974));
  jand g13952(.dina(n31974), .dinb(n281), .dout(n31975));
  jnot g13953(.din(n31975), .dout(n31976));
  jand g13954(.dina(n31841), .dinb(n31232), .dout(n31977));
  jxor g13955(.dina(n31814), .dinb(n31922), .dout(n31978));
  jand g13956(.dina(n31978), .dinb(n31947), .dout(n31979));
  jor  g13957(.dina(n31979), .dinb(n31977), .dout(n31980));
  jand g13958(.dina(n31980), .dinb(n285), .dout(n31981));
  jnot g13959(.din(n31981), .dout(n31982));
  jand g13960(.dina(n31841), .dinb(n31238), .dout(n31983));
  jxor g13961(.dina(n31810), .dinb(n31920), .dout(n31984));
  jand g13962(.dina(n31984), .dinb(n31947), .dout(n31985));
  jor  g13963(.dina(n31985), .dinb(n31983), .dout(n31986));
  jand g13964(.dina(n31986), .dinb(n284), .dout(n31987));
  jnot g13965(.din(n31987), .dout(n31988));
  jand g13966(.dina(n31841), .dinb(n31244), .dout(n31989));
  jxor g13967(.dina(n31806), .dinb(n31918), .dout(n31990));
  jand g13968(.dina(n31990), .dinb(n31947), .dout(n31991));
  jor  g13969(.dina(n31991), .dinb(n31989), .dout(n31992));
  jand g13970(.dina(n31992), .dinb(n291), .dout(n31993));
  jnot g13971(.din(n31993), .dout(n31994));
  jand g13972(.dina(n31841), .dinb(n31250), .dout(n31995));
  jxor g13973(.dina(n31802), .dinb(n31916), .dout(n31996));
  jand g13974(.dina(n31996), .dinb(n31947), .dout(n31997));
  jor  g13975(.dina(n31997), .dinb(n31995), .dout(n31998));
  jand g13976(.dina(n31998), .dinb(n290), .dout(n31999));
  jnot g13977(.din(n31999), .dout(n32000));
  jand g13978(.dina(n31841), .dinb(n31256), .dout(n32001));
  jxor g13979(.dina(n31798), .dinb(n31914), .dout(n32002));
  jand g13980(.dina(n32002), .dinb(n31947), .dout(n32003));
  jor  g13981(.dina(n32003), .dinb(n32001), .dout(n32004));
  jand g13982(.dina(n32004), .dinb(n294), .dout(n32005));
  jnot g13983(.din(n32005), .dout(n32006));
  jand g13984(.dina(n31841), .dinb(n31262), .dout(n32007));
  jxor g13985(.dina(n31794), .dinb(n31912), .dout(n32008));
  jand g13986(.dina(n32008), .dinb(n31947), .dout(n32009));
  jor  g13987(.dina(n32009), .dinb(n32007), .dout(n32010));
  jand g13988(.dina(n32010), .dinb(n293), .dout(n32011));
  jnot g13989(.din(n32011), .dout(n32012));
  jand g13990(.dina(n31841), .dinb(n31268), .dout(n32013));
  jxor g13991(.dina(n31790), .dinb(n31910), .dout(n32014));
  jand g13992(.dina(n32014), .dinb(n31947), .dout(n32015));
  jor  g13993(.dina(n32015), .dinb(n32013), .dout(n32016));
  jand g13994(.dina(n32016), .dinb(n301), .dout(n32017));
  jnot g13995(.din(n32017), .dout(n32018));
  jand g13996(.dina(n31841), .dinb(n31274), .dout(n32019));
  jxor g13997(.dina(n31786), .dinb(n31908), .dout(n32020));
  jand g13998(.dina(n32020), .dinb(n31947), .dout(n32021));
  jor  g13999(.dina(n32021), .dinb(n32019), .dout(n32022));
  jand g14000(.dina(n32022), .dinb(n298), .dout(n32023));
  jnot g14001(.din(n32023), .dout(n32024));
  jand g14002(.dina(n31841), .dinb(n31280), .dout(n32025));
  jxor g14003(.dina(n31782), .dinb(n31906), .dout(n32026));
  jand g14004(.dina(n32026), .dinb(n31947), .dout(n32027));
  jor  g14005(.dina(n32027), .dinb(n32025), .dout(n32028));
  jand g14006(.dina(n32028), .dinb(n297), .dout(n32029));
  jnot g14007(.din(n32029), .dout(n32030));
  jand g14008(.dina(n31841), .dinb(n31286), .dout(n32031));
  jxor g14009(.dina(n31778), .dinb(n31904), .dout(n32032));
  jand g14010(.dina(n32032), .dinb(n31947), .dout(n32033));
  jor  g14011(.dina(n32033), .dinb(n32031), .dout(n32034));
  jand g14012(.dina(n32034), .dinb(n300), .dout(n32035));
  jnot g14013(.din(n32035), .dout(n32036));
  jand g14014(.dina(n31841), .dinb(n31292), .dout(n32037));
  jxor g14015(.dina(n31774), .dinb(n31902), .dout(n32038));
  jand g14016(.dina(n32038), .dinb(n31947), .dout(n32039));
  jor  g14017(.dina(n32039), .dinb(n32037), .dout(n32040));
  jand g14018(.dina(n32040), .dinb(n424), .dout(n32041));
  jnot g14019(.din(n32041), .dout(n32042));
  jand g14020(.dina(n31841), .dinb(n31298), .dout(n32043));
  jxor g14021(.dina(n31770), .dinb(n31900), .dout(n32044));
  jand g14022(.dina(n32044), .dinb(n31947), .dout(n32045));
  jor  g14023(.dina(n32045), .dinb(n32043), .dout(n32046));
  jand g14024(.dina(n32046), .dinb(n427), .dout(n32047));
  jnot g14025(.din(n32047), .dout(n32048));
  jand g14026(.dina(n31841), .dinb(n31304), .dout(n32049));
  jxor g14027(.dina(n31766), .dinb(n31898), .dout(n32050));
  jand g14028(.dina(n32050), .dinb(n31947), .dout(n32051));
  jor  g14029(.dina(n32051), .dinb(n32049), .dout(n32052));
  jand g14030(.dina(n32052), .dinb(n426), .dout(n32053));
  jnot g14031(.din(n32053), .dout(n32054));
  jand g14032(.dina(n31841), .dinb(n31310), .dout(n32055));
  jxor g14033(.dina(n31762), .dinb(n31896), .dout(n32056));
  jand g14034(.dina(n32056), .dinb(n31947), .dout(n32057));
  jor  g14035(.dina(n32057), .dinb(n32055), .dout(n32058));
  jand g14036(.dina(n32058), .dinb(n410), .dout(n32059));
  jnot g14037(.din(n32059), .dout(n32060));
  jand g14038(.dina(n31841), .dinb(n31316), .dout(n32061));
  jxor g14039(.dina(n31758), .dinb(n31894), .dout(n32062));
  jand g14040(.dina(n32062), .dinb(n31947), .dout(n32063));
  jor  g14041(.dina(n32063), .dinb(n32061), .dout(n32064));
  jand g14042(.dina(n32064), .dinb(n409), .dout(n32065));
  jnot g14043(.din(n32065), .dout(n32066));
  jand g14044(.dina(n31841), .dinb(n31322), .dout(n32067));
  jxor g14045(.dina(n31754), .dinb(n31892), .dout(n32068));
  jand g14046(.dina(n32068), .dinb(n31947), .dout(n32069));
  jor  g14047(.dina(n32069), .dinb(n32067), .dout(n32070));
  jand g14048(.dina(n32070), .dinb(n413), .dout(n32071));
  jnot g14049(.din(n32071), .dout(n32072));
  jand g14050(.dina(n31841), .dinb(n31328), .dout(n32073));
  jxor g14051(.dina(n31750), .dinb(n31890), .dout(n32074));
  jand g14052(.dina(n32074), .dinb(n31947), .dout(n32075));
  jor  g14053(.dina(n32075), .dinb(n32073), .dout(n32076));
  jand g14054(.dina(n32076), .dinb(n412), .dout(n32077));
  jnot g14055(.din(n32077), .dout(n32078));
  jand g14056(.dina(n31841), .dinb(n31334), .dout(n32079));
  jxor g14057(.dina(n31746), .dinb(n31888), .dout(n32080));
  jand g14058(.dina(n32080), .dinb(n31947), .dout(n32081));
  jor  g14059(.dina(n32081), .dinb(n32079), .dout(n32082));
  jand g14060(.dina(n32082), .dinb(n406), .dout(n32083));
  jnot g14061(.din(n32083), .dout(n32084));
  jand g14062(.dina(n31841), .dinb(n31340), .dout(n32085));
  jxor g14063(.dina(n31742), .dinb(n31886), .dout(n32086));
  jand g14064(.dina(n32086), .dinb(n31947), .dout(n32087));
  jor  g14065(.dina(n32087), .dinb(n32085), .dout(n32088));
  jand g14066(.dina(n32088), .dinb(n405), .dout(n32089));
  jnot g14067(.din(n32089), .dout(n32090));
  jand g14068(.dina(n31841), .dinb(n31346), .dout(n32091));
  jxor g14069(.dina(n31738), .dinb(n31884), .dout(n32092));
  jand g14070(.dina(n32092), .dinb(n31947), .dout(n32093));
  jor  g14071(.dina(n32093), .dinb(n32091), .dout(n32094));
  jand g14072(.dina(n32094), .dinb(n2714), .dout(n32095));
  jnot g14073(.din(n32095), .dout(n32096));
  jand g14074(.dina(n31841), .dinb(n31352), .dout(n32097));
  jxor g14075(.dina(n31734), .dinb(n31882), .dout(n32098));
  jand g14076(.dina(n32098), .dinb(n31947), .dout(n32099));
  jor  g14077(.dina(n32099), .dinb(n32097), .dout(n32100));
  jand g14078(.dina(n32100), .dinb(n2547), .dout(n32101));
  jnot g14079(.din(n32101), .dout(n32102));
  jand g14080(.dina(n31841), .dinb(n31358), .dout(n32103));
  jxor g14081(.dina(n31730), .dinb(n31880), .dout(n32104));
  jand g14082(.dina(n32104), .dinb(n31947), .dout(n32105));
  jor  g14083(.dina(n32105), .dinb(n32103), .dout(n32106));
  jand g14084(.dina(n32106), .dinb(n417), .dout(n32107));
  jnot g14085(.din(n32107), .dout(n32108));
  jand g14086(.dina(n31841), .dinb(n31364), .dout(n32109));
  jxor g14087(.dina(n31726), .dinb(n31878), .dout(n32110));
  jand g14088(.dina(n32110), .dinb(n31947), .dout(n32111));
  jor  g14089(.dina(n32111), .dinb(n32109), .dout(n32112));
  jand g14090(.dina(n32112), .dinb(n416), .dout(n32113));
  jnot g14091(.din(n32113), .dout(n32114));
  jand g14092(.dina(n31841), .dinb(n31370), .dout(n32115));
  jxor g14093(.dina(n31722), .dinb(n31876), .dout(n32116));
  jand g14094(.dina(n32116), .dinb(n31947), .dout(n32117));
  jor  g14095(.dina(n32117), .dinb(n32115), .dout(n32118));
  jand g14096(.dina(n32118), .dinb(n422), .dout(n32119));
  jnot g14097(.din(n32119), .dout(n32120));
  jand g14098(.dina(n31841), .dinb(n31376), .dout(n32121));
  jxor g14099(.dina(n31718), .dinb(n31874), .dout(n32122));
  jand g14100(.dina(n32122), .dinb(n31947), .dout(n32123));
  jor  g14101(.dina(n32123), .dinb(n32121), .dout(n32124));
  jand g14102(.dina(n32124), .dinb(n421), .dout(n32125));
  jnot g14103(.din(n32125), .dout(n32126));
  jand g14104(.dina(n31841), .dinb(n31382), .dout(n32127));
  jxor g14105(.dina(n31714), .dinb(n31872), .dout(n32128));
  jand g14106(.dina(n32128), .dinb(n31947), .dout(n32129));
  jor  g14107(.dina(n32129), .dinb(n32127), .dout(n32130));
  jand g14108(.dina(n32130), .dinb(n433), .dout(n32131));
  jnot g14109(.din(n32131), .dout(n32132));
  jand g14110(.dina(n31841), .dinb(n31388), .dout(n32133));
  jxor g14111(.dina(n31710), .dinb(n31870), .dout(n32134));
  jand g14112(.dina(n32134), .dinb(n31947), .dout(n32135));
  jor  g14113(.dina(n32135), .dinb(n32133), .dout(n32136));
  jand g14114(.dina(n32136), .dinb(n432), .dout(n32137));
  jnot g14115(.din(n32137), .dout(n32138));
  jand g14116(.dina(n31841), .dinb(n31394), .dout(n32139));
  jxor g14117(.dina(n31706), .dinb(n31868), .dout(n32140));
  jand g14118(.dina(n32140), .dinb(n31947), .dout(n32141));
  jor  g14119(.dina(n32141), .dinb(n32139), .dout(n32142));
  jand g14120(.dina(n32142), .dinb(n436), .dout(n32143));
  jnot g14121(.din(n32143), .dout(n32144));
  jand g14122(.dina(n31841), .dinb(n31400), .dout(n32145));
  jxor g14123(.dina(n31702), .dinb(n31866), .dout(n32146));
  jand g14124(.dina(n32146), .dinb(n31947), .dout(n32147));
  jor  g14125(.dina(n32147), .dinb(n32145), .dout(n32148));
  jand g14126(.dina(n32148), .dinb(n435), .dout(n32149));
  jnot g14127(.din(n32149), .dout(n32150));
  jand g14128(.dina(n31841), .dinb(n31406), .dout(n32151));
  jxor g14129(.dina(n31698), .dinb(n31864), .dout(n32152));
  jand g14130(.dina(n32152), .dinb(n31947), .dout(n32153));
  jor  g14131(.dina(n32153), .dinb(n32151), .dout(n32154));
  jand g14132(.dina(n32154), .dinb(n440), .dout(n32155));
  jnot g14133(.din(n32155), .dout(n32156));
  jand g14134(.dina(n31841), .dinb(n31412), .dout(n32157));
  jxor g14135(.dina(n31694), .dinb(n31862), .dout(n32158));
  jand g14136(.dina(n32158), .dinb(n31947), .dout(n32159));
  jor  g14137(.dina(n32159), .dinb(n32157), .dout(n32160));
  jand g14138(.dina(n32160), .dinb(n439), .dout(n32161));
  jnot g14139(.din(n32161), .dout(n32162));
  jand g14140(.dina(n31841), .dinb(n31418), .dout(n32163));
  jxor g14141(.dina(n31690), .dinb(n31860), .dout(n32164));
  jand g14142(.dina(n32164), .dinb(n31947), .dout(n32165));
  jor  g14143(.dina(n32165), .dinb(n32163), .dout(n32166));
  jand g14144(.dina(n32166), .dinb(n325), .dout(n32167));
  jnot g14145(.din(n32167), .dout(n32168));
  jand g14146(.dina(n31841), .dinb(n31424), .dout(n32169));
  jxor g14147(.dina(n31686), .dinb(n31858), .dout(n32170));
  jand g14148(.dina(n32170), .dinb(n31947), .dout(n32171));
  jor  g14149(.dina(n32171), .dinb(n32169), .dout(n32172));
  jand g14150(.dina(n32172), .dinb(n324), .dout(n32173));
  jnot g14151(.din(n32173), .dout(n32174));
  jand g14152(.dina(n31841), .dinb(n31430), .dout(n32175));
  jxor g14153(.dina(n31682), .dinb(n31856), .dout(n32176));
  jand g14154(.dina(n32176), .dinb(n31947), .dout(n32177));
  jor  g14155(.dina(n32177), .dinb(n32175), .dout(n32178));
  jand g14156(.dina(n32178), .dinb(n323), .dout(n32179));
  jnot g14157(.din(n32179), .dout(n32180));
  jand g14158(.dina(n31841), .dinb(n31436), .dout(n32181));
  jxor g14159(.dina(n31678), .dinb(n31854), .dout(n32182));
  jand g14160(.dina(n32182), .dinb(n31947), .dout(n32183));
  jor  g14161(.dina(n32183), .dinb(n32181), .dout(n32184));
  jand g14162(.dina(n32184), .dinb(n335), .dout(n32185));
  jnot g14163(.din(n32185), .dout(n32186));
  jand g14164(.dina(n31841), .dinb(n31442), .dout(n32187));
  jxor g14165(.dina(n31674), .dinb(n31852), .dout(n32188));
  jand g14166(.dina(n32188), .dinb(n31947), .dout(n32189));
  jor  g14167(.dina(n32189), .dinb(n32187), .dout(n32190));
  jand g14168(.dina(n32190), .dinb(n334), .dout(n32191));
  jnot g14169(.din(n32191), .dout(n32192));
  jand g14170(.dina(n31841), .dinb(n31448), .dout(n32193));
  jxor g14171(.dina(n31670), .dinb(n31850), .dout(n32194));
  jand g14172(.dina(n32194), .dinb(n31947), .dout(n32195));
  jor  g14173(.dina(n32195), .dinb(n32193), .dout(n32196));
  jand g14174(.dina(n32196), .dinb(n338), .dout(n32197));
  jnot g14175(.din(n32197), .dout(n32198));
  jand g14176(.dina(n31841), .dinb(n31457), .dout(n32199));
  jxor g14177(.dina(n31666), .dinb(n31848), .dout(n32200));
  jand g14178(.dina(n32200), .dinb(n31947), .dout(n32201));
  jor  g14179(.dina(n32201), .dinb(n32199), .dout(n32202));
  jand g14180(.dina(n32202), .dinb(n337), .dout(n32203));
  jnot g14181(.din(n32203), .dout(n32204));
  jand g14182(.dina(n31841), .dinb(n31465), .dout(n32205));
  jxor g14183(.dina(n31662), .dinb(n31846), .dout(n32206));
  jand g14184(.dina(n32206), .dinb(n31947), .dout(n32207));
  jor  g14185(.dina(n32207), .dinb(n32205), .dout(n32208));
  jand g14186(.dina(n32208), .dinb(n344), .dout(n32209));
  jnot g14187(.din(n32209), .dout(n32210));
  jand g14188(.dina(n31841), .dinb(n31653), .dout(n32211));
  jxor g14189(.dina(n31844), .dinb(n10471), .dout(n32212));
  jand g14190(.dina(n32212), .dinb(n31947), .dout(n32213));
  jor  g14191(.dina(n32213), .dinb(n32211), .dout(n32214));
  jand g14192(.dina(n32214), .dinb(n348), .dout(n32215));
  jnot g14193(.din(n32215), .dout(n32216));
  jor  g14194(.dina(n31841), .dinb(n18364), .dout(n32217));
  jand g14195(.dina(n32217), .dinb(a17 ), .dout(n32218));
  jor  g14196(.dina(n31841), .dinb(n10471), .dout(n32219));
  jnot g14197(.din(n32219), .dout(n32220));
  jor  g14198(.dina(n32220), .dinb(n32218), .dout(n32221));
  jand g14199(.dina(n32221), .dinb(n258), .dout(n32222));
  jnot g14200(.din(n32222), .dout(n32223));
  jand g14201(.dina(n31947), .dinb(b0 ), .dout(n32224));
  jor  g14202(.dina(n32224), .dinb(n10469), .dout(n32225));
  jand g14203(.dina(n32219), .dinb(n32225), .dout(n32226));
  jxor g14204(.dina(n32226), .dinb(n258), .dout(n32227));
  jor  g14205(.dina(n32227), .dinb(n10854), .dout(n32228));
  jand g14206(.dina(n32228), .dinb(n32223), .dout(n32229));
  jxor g14207(.dina(n32214), .dinb(n348), .dout(n32230));
  jnot g14208(.din(n32230), .dout(n32231));
  jor  g14209(.dina(n32231), .dinb(n32229), .dout(n32232));
  jand g14210(.dina(n32232), .dinb(n32216), .dout(n32233));
  jxor g14211(.dina(n32208), .dinb(n344), .dout(n32234));
  jnot g14212(.din(n32234), .dout(n32235));
  jor  g14213(.dina(n32235), .dinb(n32233), .dout(n32236));
  jand g14214(.dina(n32236), .dinb(n32210), .dout(n32237));
  jxor g14215(.dina(n32202), .dinb(n337), .dout(n32238));
  jnot g14216(.din(n32238), .dout(n32239));
  jor  g14217(.dina(n32239), .dinb(n32237), .dout(n32240));
  jand g14218(.dina(n32240), .dinb(n32204), .dout(n32241));
  jxor g14219(.dina(n32196), .dinb(n338), .dout(n32242));
  jnot g14220(.din(n32242), .dout(n32243));
  jor  g14221(.dina(n32243), .dinb(n32241), .dout(n32244));
  jand g14222(.dina(n32244), .dinb(n32198), .dout(n32245));
  jxor g14223(.dina(n32190), .dinb(n334), .dout(n32246));
  jnot g14224(.din(n32246), .dout(n32247));
  jor  g14225(.dina(n32247), .dinb(n32245), .dout(n32248));
  jand g14226(.dina(n32248), .dinb(n32192), .dout(n32249));
  jxor g14227(.dina(n32184), .dinb(n335), .dout(n32250));
  jnot g14228(.din(n32250), .dout(n32251));
  jor  g14229(.dina(n32251), .dinb(n32249), .dout(n32252));
  jand g14230(.dina(n32252), .dinb(n32186), .dout(n32253));
  jxor g14231(.dina(n32178), .dinb(n323), .dout(n32254));
  jnot g14232(.din(n32254), .dout(n32255));
  jor  g14233(.dina(n32255), .dinb(n32253), .dout(n32256));
  jand g14234(.dina(n32256), .dinb(n32180), .dout(n32257));
  jxor g14235(.dina(n32172), .dinb(n324), .dout(n32258));
  jnot g14236(.din(n32258), .dout(n32259));
  jor  g14237(.dina(n32259), .dinb(n32257), .dout(n32260));
  jand g14238(.dina(n32260), .dinb(n32174), .dout(n32261));
  jxor g14239(.dina(n32166), .dinb(n325), .dout(n32262));
  jnot g14240(.din(n32262), .dout(n32263));
  jor  g14241(.dina(n32263), .dinb(n32261), .dout(n32264));
  jand g14242(.dina(n32264), .dinb(n32168), .dout(n32265));
  jxor g14243(.dina(n32160), .dinb(n439), .dout(n32266));
  jnot g14244(.din(n32266), .dout(n32267));
  jor  g14245(.dina(n32267), .dinb(n32265), .dout(n32268));
  jand g14246(.dina(n32268), .dinb(n32162), .dout(n32269));
  jxor g14247(.dina(n32154), .dinb(n440), .dout(n32270));
  jnot g14248(.din(n32270), .dout(n32271));
  jor  g14249(.dina(n32271), .dinb(n32269), .dout(n32272));
  jand g14250(.dina(n32272), .dinb(n32156), .dout(n32273));
  jxor g14251(.dina(n32148), .dinb(n435), .dout(n32274));
  jnot g14252(.din(n32274), .dout(n32275));
  jor  g14253(.dina(n32275), .dinb(n32273), .dout(n32276));
  jand g14254(.dina(n32276), .dinb(n32150), .dout(n32277));
  jxor g14255(.dina(n32142), .dinb(n436), .dout(n32278));
  jnot g14256(.din(n32278), .dout(n32279));
  jor  g14257(.dina(n32279), .dinb(n32277), .dout(n32280));
  jand g14258(.dina(n32280), .dinb(n32144), .dout(n32281));
  jxor g14259(.dina(n32136), .dinb(n432), .dout(n32282));
  jnot g14260(.din(n32282), .dout(n32283));
  jor  g14261(.dina(n32283), .dinb(n32281), .dout(n32284));
  jand g14262(.dina(n32284), .dinb(n32138), .dout(n32285));
  jxor g14263(.dina(n32130), .dinb(n433), .dout(n32286));
  jnot g14264(.din(n32286), .dout(n32287));
  jor  g14265(.dina(n32287), .dinb(n32285), .dout(n32288));
  jand g14266(.dina(n32288), .dinb(n32132), .dout(n32289));
  jxor g14267(.dina(n32124), .dinb(n421), .dout(n32290));
  jnot g14268(.din(n32290), .dout(n32291));
  jor  g14269(.dina(n32291), .dinb(n32289), .dout(n32292));
  jand g14270(.dina(n32292), .dinb(n32126), .dout(n32293));
  jxor g14271(.dina(n32118), .dinb(n422), .dout(n32294));
  jnot g14272(.din(n32294), .dout(n32295));
  jor  g14273(.dina(n32295), .dinb(n32293), .dout(n32296));
  jand g14274(.dina(n32296), .dinb(n32120), .dout(n32297));
  jxor g14275(.dina(n32112), .dinb(n416), .dout(n32298));
  jnot g14276(.din(n32298), .dout(n32299));
  jor  g14277(.dina(n32299), .dinb(n32297), .dout(n32300));
  jand g14278(.dina(n32300), .dinb(n32114), .dout(n32301));
  jxor g14279(.dina(n32106), .dinb(n417), .dout(n32302));
  jnot g14280(.din(n32302), .dout(n32303));
  jor  g14281(.dina(n32303), .dinb(n32301), .dout(n32304));
  jand g14282(.dina(n32304), .dinb(n32108), .dout(n32305));
  jxor g14283(.dina(n32100), .dinb(n2547), .dout(n32306));
  jnot g14284(.din(n32306), .dout(n32307));
  jor  g14285(.dina(n32307), .dinb(n32305), .dout(n32308));
  jand g14286(.dina(n32308), .dinb(n32102), .dout(n32309));
  jxor g14287(.dina(n32094), .dinb(n2714), .dout(n32310));
  jnot g14288(.din(n32310), .dout(n32311));
  jor  g14289(.dina(n32311), .dinb(n32309), .dout(n32312));
  jand g14290(.dina(n32312), .dinb(n32096), .dout(n32313));
  jxor g14291(.dina(n32088), .dinb(n405), .dout(n32314));
  jnot g14292(.din(n32314), .dout(n32315));
  jor  g14293(.dina(n32315), .dinb(n32313), .dout(n32316));
  jand g14294(.dina(n32316), .dinb(n32090), .dout(n32317));
  jxor g14295(.dina(n32082), .dinb(n406), .dout(n32318));
  jnot g14296(.din(n32318), .dout(n32319));
  jor  g14297(.dina(n32319), .dinb(n32317), .dout(n32320));
  jand g14298(.dina(n32320), .dinb(n32084), .dout(n32321));
  jxor g14299(.dina(n32076), .dinb(n412), .dout(n32322));
  jnot g14300(.din(n32322), .dout(n32323));
  jor  g14301(.dina(n32323), .dinb(n32321), .dout(n32324));
  jand g14302(.dina(n32324), .dinb(n32078), .dout(n32325));
  jxor g14303(.dina(n32070), .dinb(n413), .dout(n32326));
  jnot g14304(.din(n32326), .dout(n32327));
  jor  g14305(.dina(n32327), .dinb(n32325), .dout(n32328));
  jand g14306(.dina(n32328), .dinb(n32072), .dout(n32329));
  jxor g14307(.dina(n32064), .dinb(n409), .dout(n32330));
  jnot g14308(.din(n32330), .dout(n32331));
  jor  g14309(.dina(n32331), .dinb(n32329), .dout(n32332));
  jand g14310(.dina(n32332), .dinb(n32066), .dout(n32333));
  jxor g14311(.dina(n32058), .dinb(n410), .dout(n32334));
  jnot g14312(.din(n32334), .dout(n32335));
  jor  g14313(.dina(n32335), .dinb(n32333), .dout(n32336));
  jand g14314(.dina(n32336), .dinb(n32060), .dout(n32337));
  jxor g14315(.dina(n32052), .dinb(n426), .dout(n32338));
  jnot g14316(.din(n32338), .dout(n32339));
  jor  g14317(.dina(n32339), .dinb(n32337), .dout(n32340));
  jand g14318(.dina(n32340), .dinb(n32054), .dout(n32341));
  jxor g14319(.dina(n32046), .dinb(n427), .dout(n32342));
  jnot g14320(.din(n32342), .dout(n32343));
  jor  g14321(.dina(n32343), .dinb(n32341), .dout(n32344));
  jand g14322(.dina(n32344), .dinb(n32048), .dout(n32345));
  jxor g14323(.dina(n32040), .dinb(n424), .dout(n32346));
  jnot g14324(.din(n32346), .dout(n32347));
  jor  g14325(.dina(n32347), .dinb(n32345), .dout(n32348));
  jand g14326(.dina(n32348), .dinb(n32042), .dout(n32349));
  jxor g14327(.dina(n32034), .dinb(n300), .dout(n32350));
  jnot g14328(.din(n32350), .dout(n32351));
  jor  g14329(.dina(n32351), .dinb(n32349), .dout(n32352));
  jand g14330(.dina(n32352), .dinb(n32036), .dout(n32353));
  jxor g14331(.dina(n32028), .dinb(n297), .dout(n32354));
  jnot g14332(.din(n32354), .dout(n32355));
  jor  g14333(.dina(n32355), .dinb(n32353), .dout(n32356));
  jand g14334(.dina(n32356), .dinb(n32030), .dout(n32357));
  jxor g14335(.dina(n32022), .dinb(n298), .dout(n32358));
  jnot g14336(.din(n32358), .dout(n32359));
  jor  g14337(.dina(n32359), .dinb(n32357), .dout(n32360));
  jand g14338(.dina(n32360), .dinb(n32024), .dout(n32361));
  jxor g14339(.dina(n32016), .dinb(n301), .dout(n32362));
  jnot g14340(.din(n32362), .dout(n32363));
  jor  g14341(.dina(n32363), .dinb(n32361), .dout(n32364));
  jand g14342(.dina(n32364), .dinb(n32018), .dout(n32365));
  jxor g14343(.dina(n32010), .dinb(n293), .dout(n32366));
  jnot g14344(.din(n32366), .dout(n32367));
  jor  g14345(.dina(n32367), .dinb(n32365), .dout(n32368));
  jand g14346(.dina(n32368), .dinb(n32012), .dout(n32369));
  jxor g14347(.dina(n32004), .dinb(n294), .dout(n32370));
  jnot g14348(.din(n32370), .dout(n32371));
  jor  g14349(.dina(n32371), .dinb(n32369), .dout(n32372));
  jand g14350(.dina(n32372), .dinb(n32006), .dout(n32373));
  jxor g14351(.dina(n31998), .dinb(n290), .dout(n32374));
  jnot g14352(.din(n32374), .dout(n32375));
  jor  g14353(.dina(n32375), .dinb(n32373), .dout(n32376));
  jand g14354(.dina(n32376), .dinb(n32000), .dout(n32377));
  jxor g14355(.dina(n31992), .dinb(n291), .dout(n32378));
  jnot g14356(.din(n32378), .dout(n32379));
  jor  g14357(.dina(n32379), .dinb(n32377), .dout(n32380));
  jand g14358(.dina(n32380), .dinb(n31994), .dout(n32381));
  jxor g14359(.dina(n31986), .dinb(n284), .dout(n32382));
  jnot g14360(.din(n32382), .dout(n32383));
  jor  g14361(.dina(n32383), .dinb(n32381), .dout(n32384));
  jand g14362(.dina(n32384), .dinb(n31988), .dout(n32385));
  jxor g14363(.dina(n31980), .dinb(n285), .dout(n32386));
  jnot g14364(.din(n32386), .dout(n32387));
  jor  g14365(.dina(n32387), .dinb(n32385), .dout(n32388));
  jand g14366(.dina(n32388), .dinb(n31982), .dout(n32389));
  jxor g14367(.dina(n31974), .dinb(n281), .dout(n32390));
  jnot g14368(.din(n32390), .dout(n32391));
  jor  g14369(.dina(n32391), .dinb(n32389), .dout(n32392));
  jand g14370(.dina(n32392), .dinb(n31976), .dout(n32393));
  jxor g14371(.dina(n31968), .dinb(n282), .dout(n32394));
  jnot g14372(.din(n32394), .dout(n32395));
  jor  g14373(.dina(n32395), .dinb(n32393), .dout(n32396));
  jand g14374(.dina(n32396), .dinb(n31970), .dout(n32397));
  jxor g14375(.dina(n31962), .dinb(n397), .dout(n32398));
  jnot g14376(.din(n32398), .dout(n32399));
  jor  g14377(.dina(n32399), .dinb(n32397), .dout(n32400));
  jand g14378(.dina(n32400), .dinb(n31964), .dout(n32401));
  jxor g14379(.dina(n31956), .dinb(n513), .dout(n32402));
  jnot g14380(.din(n32402), .dout(n32403));
  jor  g14381(.dina(n32403), .dinb(n32401), .dout(n32404));
  jand g14382(.dina(n32404), .dinb(n31958), .dout(n32405));
  jxor g14383(.dina(n31950), .dinb(n514), .dout(n32406));
  jnot g14384(.din(n32406), .dout(n32407));
  jor  g14385(.dina(n32407), .dinb(n32405), .dout(n32408));
  jand g14386(.dina(n32408), .dinb(n31952), .dout(n32409));
  jxor g14387(.dina(n31940), .dinb(n510), .dout(n32410));
  jor  g14388(.dina(n32410), .dinb(n32409), .dout(n32411));
  jor  g14389(.dina(n32411), .dinb(n31944), .dout(n32412));
  jand g14390(.dina(n32412), .dinb(n31943), .dout(n32413));
  jand g14391(.dina(n32413), .dinb(n31941), .dout(n32414));
  jnot g14392(.din(n32414), .dout(n32415));
  jxor g14393(.dina(n32226), .dinb(b1 ), .dout(n32416));
  jand g14394(.dina(n32416), .dinb(n10855), .dout(n32417));
  jor  g14395(.dina(n32417), .dinb(n32222), .dout(n32418));
  jand g14396(.dina(n32230), .dinb(n32418), .dout(n32419));
  jor  g14397(.dina(n32419), .dinb(n32215), .dout(n32420));
  jand g14398(.dina(n32234), .dinb(n32420), .dout(n32421));
  jor  g14399(.dina(n32421), .dinb(n32209), .dout(n32422));
  jand g14400(.dina(n32238), .dinb(n32422), .dout(n32423));
  jor  g14401(.dina(n32423), .dinb(n32203), .dout(n32424));
  jand g14402(.dina(n32242), .dinb(n32424), .dout(n32425));
  jor  g14403(.dina(n32425), .dinb(n32197), .dout(n32426));
  jand g14404(.dina(n32246), .dinb(n32426), .dout(n32427));
  jor  g14405(.dina(n32427), .dinb(n32191), .dout(n32428));
  jand g14406(.dina(n32250), .dinb(n32428), .dout(n32429));
  jor  g14407(.dina(n32429), .dinb(n32185), .dout(n32430));
  jand g14408(.dina(n32254), .dinb(n32430), .dout(n32431));
  jor  g14409(.dina(n32431), .dinb(n32179), .dout(n32432));
  jand g14410(.dina(n32258), .dinb(n32432), .dout(n32433));
  jor  g14411(.dina(n32433), .dinb(n32173), .dout(n32434));
  jand g14412(.dina(n32262), .dinb(n32434), .dout(n32435));
  jor  g14413(.dina(n32435), .dinb(n32167), .dout(n32436));
  jand g14414(.dina(n32266), .dinb(n32436), .dout(n32437));
  jor  g14415(.dina(n32437), .dinb(n32161), .dout(n32438));
  jand g14416(.dina(n32270), .dinb(n32438), .dout(n32439));
  jor  g14417(.dina(n32439), .dinb(n32155), .dout(n32440));
  jand g14418(.dina(n32274), .dinb(n32440), .dout(n32441));
  jor  g14419(.dina(n32441), .dinb(n32149), .dout(n32442));
  jand g14420(.dina(n32278), .dinb(n32442), .dout(n32443));
  jor  g14421(.dina(n32443), .dinb(n32143), .dout(n32444));
  jand g14422(.dina(n32282), .dinb(n32444), .dout(n32445));
  jor  g14423(.dina(n32445), .dinb(n32137), .dout(n32446));
  jand g14424(.dina(n32286), .dinb(n32446), .dout(n32447));
  jor  g14425(.dina(n32447), .dinb(n32131), .dout(n32448));
  jand g14426(.dina(n32290), .dinb(n32448), .dout(n32449));
  jor  g14427(.dina(n32449), .dinb(n32125), .dout(n32450));
  jand g14428(.dina(n32294), .dinb(n32450), .dout(n32451));
  jor  g14429(.dina(n32451), .dinb(n32119), .dout(n32452));
  jand g14430(.dina(n32298), .dinb(n32452), .dout(n32453));
  jor  g14431(.dina(n32453), .dinb(n32113), .dout(n32454));
  jand g14432(.dina(n32302), .dinb(n32454), .dout(n32455));
  jor  g14433(.dina(n32455), .dinb(n32107), .dout(n32456));
  jand g14434(.dina(n32306), .dinb(n32456), .dout(n32457));
  jor  g14435(.dina(n32457), .dinb(n32101), .dout(n32458));
  jand g14436(.dina(n32310), .dinb(n32458), .dout(n32459));
  jor  g14437(.dina(n32459), .dinb(n32095), .dout(n32460));
  jand g14438(.dina(n32314), .dinb(n32460), .dout(n32461));
  jor  g14439(.dina(n32461), .dinb(n32089), .dout(n32462));
  jand g14440(.dina(n32318), .dinb(n32462), .dout(n32463));
  jor  g14441(.dina(n32463), .dinb(n32083), .dout(n32464));
  jand g14442(.dina(n32322), .dinb(n32464), .dout(n32465));
  jor  g14443(.dina(n32465), .dinb(n32077), .dout(n32466));
  jand g14444(.dina(n32326), .dinb(n32466), .dout(n32467));
  jor  g14445(.dina(n32467), .dinb(n32071), .dout(n32468));
  jand g14446(.dina(n32330), .dinb(n32468), .dout(n32469));
  jor  g14447(.dina(n32469), .dinb(n32065), .dout(n32470));
  jand g14448(.dina(n32334), .dinb(n32470), .dout(n32471));
  jor  g14449(.dina(n32471), .dinb(n32059), .dout(n32472));
  jand g14450(.dina(n32338), .dinb(n32472), .dout(n32473));
  jor  g14451(.dina(n32473), .dinb(n32053), .dout(n32474));
  jand g14452(.dina(n32342), .dinb(n32474), .dout(n32475));
  jor  g14453(.dina(n32475), .dinb(n32047), .dout(n32476));
  jand g14454(.dina(n32346), .dinb(n32476), .dout(n32477));
  jor  g14455(.dina(n32477), .dinb(n32041), .dout(n32478));
  jand g14456(.dina(n32350), .dinb(n32478), .dout(n32479));
  jor  g14457(.dina(n32479), .dinb(n32035), .dout(n32480));
  jand g14458(.dina(n32354), .dinb(n32480), .dout(n32481));
  jor  g14459(.dina(n32481), .dinb(n32029), .dout(n32482));
  jand g14460(.dina(n32358), .dinb(n32482), .dout(n32483));
  jor  g14461(.dina(n32483), .dinb(n32023), .dout(n32484));
  jand g14462(.dina(n32362), .dinb(n32484), .dout(n32485));
  jor  g14463(.dina(n32485), .dinb(n32017), .dout(n32486));
  jand g14464(.dina(n32366), .dinb(n32486), .dout(n32487));
  jor  g14465(.dina(n32487), .dinb(n32011), .dout(n32488));
  jand g14466(.dina(n32370), .dinb(n32488), .dout(n32489));
  jor  g14467(.dina(n32489), .dinb(n32005), .dout(n32490));
  jand g14468(.dina(n32374), .dinb(n32490), .dout(n32491));
  jor  g14469(.dina(n32491), .dinb(n31999), .dout(n32492));
  jand g14470(.dina(n32378), .dinb(n32492), .dout(n32493));
  jor  g14471(.dina(n32493), .dinb(n31993), .dout(n32494));
  jand g14472(.dina(n32382), .dinb(n32494), .dout(n32495));
  jor  g14473(.dina(n32495), .dinb(n31987), .dout(n32496));
  jand g14474(.dina(n32386), .dinb(n32496), .dout(n32497));
  jor  g14475(.dina(n32497), .dinb(n31981), .dout(n32498));
  jand g14476(.dina(n32390), .dinb(n32498), .dout(n32499));
  jor  g14477(.dina(n32499), .dinb(n31975), .dout(n32500));
  jand g14478(.dina(n32394), .dinb(n32500), .dout(n32501));
  jor  g14479(.dina(n32501), .dinb(n31969), .dout(n32502));
  jand g14480(.dina(n32398), .dinb(n32502), .dout(n32503));
  jor  g14481(.dina(n32503), .dinb(n31963), .dout(n32504));
  jand g14482(.dina(n32402), .dinb(n32504), .dout(n32505));
  jor  g14483(.dina(n32505), .dinb(n31957), .dout(n32506));
  jand g14484(.dina(n32406), .dinb(n32506), .dout(n32507));
  jor  g14485(.dina(n32507), .dinb(n31951), .dout(n32508));
  jnot g14486(.din(n32410), .dout(n32509));
  jand g14487(.dina(n32509), .dinb(n32508), .dout(n32510));
  jand g14488(.dina(n32409), .dinb(n510), .dout(n32511));
  jor  g14489(.dina(n32511), .dinb(n31943), .dout(n32512));
  jor  g14490(.dina(n32512), .dinb(n32510), .dout(n32513));
  jand g14491(.dina(n32513), .dinb(n32415), .dout(n32514));
  jnot g14492(.din(n32514), .dout(n32515));
  jand g14493(.dina(n32515), .dinb(n396), .dout(n32516));
  jand g14494(.dina(n32413), .dinb(n31950), .dout(n32517));
  jand g14495(.dina(n32510), .dinb(n9868), .dout(n32518));
  jor  g14496(.dina(n32518), .dinb(n31942), .dout(n32519));
  jxor g14497(.dina(n32406), .dinb(n32506), .dout(n32520));
  jand g14498(.dina(n32520), .dinb(n32519), .dout(n32521));
  jor  g14499(.dina(n32521), .dinb(n32517), .dout(n32522));
  jand g14500(.dina(n32522), .dinb(n510), .dout(n32523));
  jand g14501(.dina(n32413), .dinb(n31956), .dout(n32524));
  jxor g14502(.dina(n32402), .dinb(n32504), .dout(n32525));
  jand g14503(.dina(n32525), .dinb(n32519), .dout(n32526));
  jor  g14504(.dina(n32526), .dinb(n32524), .dout(n32527));
  jand g14505(.dina(n32527), .dinb(n514), .dout(n32528));
  jand g14506(.dina(n32413), .dinb(n31962), .dout(n32529));
  jxor g14507(.dina(n32398), .dinb(n32502), .dout(n32530));
  jand g14508(.dina(n32530), .dinb(n32519), .dout(n32531));
  jor  g14509(.dina(n32531), .dinb(n32529), .dout(n32532));
  jand g14510(.dina(n32532), .dinb(n513), .dout(n32533));
  jand g14511(.dina(n32413), .dinb(n31968), .dout(n32534));
  jxor g14512(.dina(n32394), .dinb(n32500), .dout(n32535));
  jand g14513(.dina(n32535), .dinb(n32519), .dout(n32536));
  jor  g14514(.dina(n32536), .dinb(n32534), .dout(n32537));
  jand g14515(.dina(n32537), .dinb(n397), .dout(n32538));
  jand g14516(.dina(n32413), .dinb(n31974), .dout(n32539));
  jxor g14517(.dina(n32390), .dinb(n32498), .dout(n32540));
  jand g14518(.dina(n32540), .dinb(n32519), .dout(n32541));
  jor  g14519(.dina(n32541), .dinb(n32539), .dout(n32542));
  jand g14520(.dina(n32542), .dinb(n282), .dout(n32543));
  jand g14521(.dina(n32413), .dinb(n31980), .dout(n32544));
  jxor g14522(.dina(n32386), .dinb(n32496), .dout(n32545));
  jand g14523(.dina(n32545), .dinb(n32519), .dout(n32546));
  jor  g14524(.dina(n32546), .dinb(n32544), .dout(n32547));
  jand g14525(.dina(n32547), .dinb(n281), .dout(n32548));
  jand g14526(.dina(n32413), .dinb(n31986), .dout(n32549));
  jxor g14527(.dina(n32382), .dinb(n32494), .dout(n32550));
  jand g14528(.dina(n32550), .dinb(n32519), .dout(n32551));
  jor  g14529(.dina(n32551), .dinb(n32549), .dout(n32552));
  jand g14530(.dina(n32552), .dinb(n285), .dout(n32553));
  jand g14531(.dina(n32413), .dinb(n31992), .dout(n32554));
  jxor g14532(.dina(n32378), .dinb(n32492), .dout(n32555));
  jand g14533(.dina(n32555), .dinb(n32519), .dout(n32556));
  jor  g14534(.dina(n32556), .dinb(n32554), .dout(n32557));
  jand g14535(.dina(n32557), .dinb(n284), .dout(n32558));
  jand g14536(.dina(n32413), .dinb(n31998), .dout(n32559));
  jxor g14537(.dina(n32374), .dinb(n32490), .dout(n32560));
  jand g14538(.dina(n32560), .dinb(n32519), .dout(n32561));
  jor  g14539(.dina(n32561), .dinb(n32559), .dout(n32562));
  jand g14540(.dina(n32562), .dinb(n291), .dout(n32563));
  jand g14541(.dina(n32413), .dinb(n32004), .dout(n32564));
  jxor g14542(.dina(n32370), .dinb(n32488), .dout(n32565));
  jand g14543(.dina(n32565), .dinb(n32519), .dout(n32566));
  jor  g14544(.dina(n32566), .dinb(n32564), .dout(n32567));
  jand g14545(.dina(n32567), .dinb(n290), .dout(n32568));
  jand g14546(.dina(n32413), .dinb(n32010), .dout(n32569));
  jxor g14547(.dina(n32366), .dinb(n32486), .dout(n32570));
  jand g14548(.dina(n32570), .dinb(n32519), .dout(n32571));
  jor  g14549(.dina(n32571), .dinb(n32569), .dout(n32572));
  jand g14550(.dina(n32572), .dinb(n294), .dout(n32573));
  jand g14551(.dina(n32413), .dinb(n32016), .dout(n32574));
  jxor g14552(.dina(n32362), .dinb(n32484), .dout(n32575));
  jand g14553(.dina(n32575), .dinb(n32519), .dout(n32576));
  jor  g14554(.dina(n32576), .dinb(n32574), .dout(n32577));
  jand g14555(.dina(n32577), .dinb(n293), .dout(n32578));
  jand g14556(.dina(n32413), .dinb(n32022), .dout(n32579));
  jxor g14557(.dina(n32358), .dinb(n32482), .dout(n32580));
  jand g14558(.dina(n32580), .dinb(n32519), .dout(n32581));
  jor  g14559(.dina(n32581), .dinb(n32579), .dout(n32582));
  jand g14560(.dina(n32582), .dinb(n301), .dout(n32583));
  jand g14561(.dina(n32413), .dinb(n32028), .dout(n32584));
  jxor g14562(.dina(n32354), .dinb(n32480), .dout(n32585));
  jand g14563(.dina(n32585), .dinb(n32519), .dout(n32586));
  jor  g14564(.dina(n32586), .dinb(n32584), .dout(n32587));
  jand g14565(.dina(n32587), .dinb(n298), .dout(n32588));
  jand g14566(.dina(n32413), .dinb(n32034), .dout(n32589));
  jxor g14567(.dina(n32350), .dinb(n32478), .dout(n32590));
  jand g14568(.dina(n32590), .dinb(n32519), .dout(n32591));
  jor  g14569(.dina(n32591), .dinb(n32589), .dout(n32592));
  jand g14570(.dina(n32592), .dinb(n297), .dout(n32593));
  jand g14571(.dina(n32413), .dinb(n32040), .dout(n32594));
  jxor g14572(.dina(n32346), .dinb(n32476), .dout(n32595));
  jand g14573(.dina(n32595), .dinb(n32519), .dout(n32596));
  jor  g14574(.dina(n32596), .dinb(n32594), .dout(n32597));
  jand g14575(.dina(n32597), .dinb(n300), .dout(n32598));
  jand g14576(.dina(n32413), .dinb(n32046), .dout(n32599));
  jxor g14577(.dina(n32342), .dinb(n32474), .dout(n32600));
  jand g14578(.dina(n32600), .dinb(n32519), .dout(n32601));
  jor  g14579(.dina(n32601), .dinb(n32599), .dout(n32602));
  jand g14580(.dina(n32602), .dinb(n424), .dout(n32603));
  jand g14581(.dina(n32413), .dinb(n32052), .dout(n32604));
  jxor g14582(.dina(n32338), .dinb(n32472), .dout(n32605));
  jand g14583(.dina(n32605), .dinb(n32519), .dout(n32606));
  jor  g14584(.dina(n32606), .dinb(n32604), .dout(n32607));
  jand g14585(.dina(n32607), .dinb(n427), .dout(n32608));
  jand g14586(.dina(n32413), .dinb(n32058), .dout(n32609));
  jxor g14587(.dina(n32334), .dinb(n32470), .dout(n32610));
  jand g14588(.dina(n32610), .dinb(n32519), .dout(n32611));
  jor  g14589(.dina(n32611), .dinb(n32609), .dout(n32612));
  jand g14590(.dina(n32612), .dinb(n426), .dout(n32613));
  jand g14591(.dina(n32413), .dinb(n32064), .dout(n32614));
  jxor g14592(.dina(n32330), .dinb(n32468), .dout(n32615));
  jand g14593(.dina(n32615), .dinb(n32519), .dout(n32616));
  jor  g14594(.dina(n32616), .dinb(n32614), .dout(n32617));
  jand g14595(.dina(n32617), .dinb(n410), .dout(n32618));
  jand g14596(.dina(n32413), .dinb(n32070), .dout(n32619));
  jxor g14597(.dina(n32326), .dinb(n32466), .dout(n32620));
  jand g14598(.dina(n32620), .dinb(n32519), .dout(n32621));
  jor  g14599(.dina(n32621), .dinb(n32619), .dout(n32622));
  jand g14600(.dina(n32622), .dinb(n409), .dout(n32623));
  jand g14601(.dina(n32413), .dinb(n32076), .dout(n32624));
  jxor g14602(.dina(n32322), .dinb(n32464), .dout(n32625));
  jand g14603(.dina(n32625), .dinb(n32519), .dout(n32626));
  jor  g14604(.dina(n32626), .dinb(n32624), .dout(n32627));
  jand g14605(.dina(n32627), .dinb(n413), .dout(n32628));
  jand g14606(.dina(n32413), .dinb(n32082), .dout(n32629));
  jxor g14607(.dina(n32318), .dinb(n32462), .dout(n32630));
  jand g14608(.dina(n32630), .dinb(n32519), .dout(n32631));
  jor  g14609(.dina(n32631), .dinb(n32629), .dout(n32632));
  jand g14610(.dina(n32632), .dinb(n412), .dout(n32633));
  jand g14611(.dina(n32413), .dinb(n32088), .dout(n32634));
  jxor g14612(.dina(n32314), .dinb(n32460), .dout(n32635));
  jand g14613(.dina(n32635), .dinb(n32519), .dout(n32636));
  jor  g14614(.dina(n32636), .dinb(n32634), .dout(n32637));
  jand g14615(.dina(n32637), .dinb(n406), .dout(n32638));
  jand g14616(.dina(n32413), .dinb(n32094), .dout(n32639));
  jxor g14617(.dina(n32310), .dinb(n32458), .dout(n32640));
  jand g14618(.dina(n32640), .dinb(n32519), .dout(n32641));
  jor  g14619(.dina(n32641), .dinb(n32639), .dout(n32642));
  jand g14620(.dina(n32642), .dinb(n405), .dout(n32643));
  jand g14621(.dina(n32413), .dinb(n32100), .dout(n32644));
  jxor g14622(.dina(n32306), .dinb(n32456), .dout(n32645));
  jand g14623(.dina(n32645), .dinb(n32519), .dout(n32646));
  jor  g14624(.dina(n32646), .dinb(n32644), .dout(n32647));
  jand g14625(.dina(n32647), .dinb(n2714), .dout(n32648));
  jand g14626(.dina(n32413), .dinb(n32106), .dout(n32649));
  jxor g14627(.dina(n32302), .dinb(n32454), .dout(n32650));
  jand g14628(.dina(n32650), .dinb(n32519), .dout(n32651));
  jor  g14629(.dina(n32651), .dinb(n32649), .dout(n32652));
  jand g14630(.dina(n32652), .dinb(n2547), .dout(n32653));
  jand g14631(.dina(n32413), .dinb(n32112), .dout(n32654));
  jxor g14632(.dina(n32298), .dinb(n32452), .dout(n32655));
  jand g14633(.dina(n32655), .dinb(n32519), .dout(n32656));
  jor  g14634(.dina(n32656), .dinb(n32654), .dout(n32657));
  jand g14635(.dina(n32657), .dinb(n417), .dout(n32658));
  jand g14636(.dina(n32413), .dinb(n32118), .dout(n32659));
  jxor g14637(.dina(n32294), .dinb(n32450), .dout(n32660));
  jand g14638(.dina(n32660), .dinb(n32519), .dout(n32661));
  jor  g14639(.dina(n32661), .dinb(n32659), .dout(n32662));
  jand g14640(.dina(n32662), .dinb(n416), .dout(n32663));
  jand g14641(.dina(n32413), .dinb(n32124), .dout(n32664));
  jxor g14642(.dina(n32290), .dinb(n32448), .dout(n32665));
  jand g14643(.dina(n32665), .dinb(n32519), .dout(n32666));
  jor  g14644(.dina(n32666), .dinb(n32664), .dout(n32667));
  jand g14645(.dina(n32667), .dinb(n422), .dout(n32668));
  jand g14646(.dina(n32413), .dinb(n32130), .dout(n32669));
  jxor g14647(.dina(n32286), .dinb(n32446), .dout(n32670));
  jand g14648(.dina(n32670), .dinb(n32519), .dout(n32671));
  jor  g14649(.dina(n32671), .dinb(n32669), .dout(n32672));
  jand g14650(.dina(n32672), .dinb(n421), .dout(n32673));
  jand g14651(.dina(n32413), .dinb(n32136), .dout(n32674));
  jxor g14652(.dina(n32282), .dinb(n32444), .dout(n32675));
  jand g14653(.dina(n32675), .dinb(n32519), .dout(n32676));
  jor  g14654(.dina(n32676), .dinb(n32674), .dout(n32677));
  jand g14655(.dina(n32677), .dinb(n433), .dout(n32678));
  jand g14656(.dina(n32413), .dinb(n32142), .dout(n32679));
  jxor g14657(.dina(n32278), .dinb(n32442), .dout(n32680));
  jand g14658(.dina(n32680), .dinb(n32519), .dout(n32681));
  jor  g14659(.dina(n32681), .dinb(n32679), .dout(n32682));
  jand g14660(.dina(n32682), .dinb(n432), .dout(n32683));
  jand g14661(.dina(n32413), .dinb(n32148), .dout(n32684));
  jxor g14662(.dina(n32274), .dinb(n32440), .dout(n32685));
  jand g14663(.dina(n32685), .dinb(n32519), .dout(n32686));
  jor  g14664(.dina(n32686), .dinb(n32684), .dout(n32687));
  jand g14665(.dina(n32687), .dinb(n436), .dout(n32688));
  jand g14666(.dina(n32413), .dinb(n32154), .dout(n32689));
  jxor g14667(.dina(n32270), .dinb(n32438), .dout(n32690));
  jand g14668(.dina(n32690), .dinb(n32519), .dout(n32691));
  jor  g14669(.dina(n32691), .dinb(n32689), .dout(n32692));
  jand g14670(.dina(n32692), .dinb(n435), .dout(n32693));
  jand g14671(.dina(n32413), .dinb(n32160), .dout(n32694));
  jxor g14672(.dina(n32266), .dinb(n32436), .dout(n32695));
  jand g14673(.dina(n32695), .dinb(n32519), .dout(n32696));
  jor  g14674(.dina(n32696), .dinb(n32694), .dout(n32697));
  jand g14675(.dina(n32697), .dinb(n440), .dout(n32698));
  jand g14676(.dina(n32413), .dinb(n32166), .dout(n32699));
  jxor g14677(.dina(n32262), .dinb(n32434), .dout(n32700));
  jand g14678(.dina(n32700), .dinb(n32519), .dout(n32701));
  jor  g14679(.dina(n32701), .dinb(n32699), .dout(n32702));
  jand g14680(.dina(n32702), .dinb(n439), .dout(n32703));
  jand g14681(.dina(n32413), .dinb(n32172), .dout(n32704));
  jxor g14682(.dina(n32258), .dinb(n32432), .dout(n32705));
  jand g14683(.dina(n32705), .dinb(n32519), .dout(n32706));
  jor  g14684(.dina(n32706), .dinb(n32704), .dout(n32707));
  jand g14685(.dina(n32707), .dinb(n325), .dout(n32708));
  jand g14686(.dina(n32413), .dinb(n32178), .dout(n32709));
  jxor g14687(.dina(n32254), .dinb(n32430), .dout(n32710));
  jand g14688(.dina(n32710), .dinb(n32519), .dout(n32711));
  jor  g14689(.dina(n32711), .dinb(n32709), .dout(n32712));
  jand g14690(.dina(n32712), .dinb(n324), .dout(n32713));
  jand g14691(.dina(n32413), .dinb(n32184), .dout(n32714));
  jxor g14692(.dina(n32250), .dinb(n32428), .dout(n32715));
  jand g14693(.dina(n32715), .dinb(n32519), .dout(n32716));
  jor  g14694(.dina(n32716), .dinb(n32714), .dout(n32717));
  jand g14695(.dina(n32717), .dinb(n323), .dout(n32718));
  jand g14696(.dina(n32413), .dinb(n32190), .dout(n32719));
  jxor g14697(.dina(n32246), .dinb(n32426), .dout(n32720));
  jand g14698(.dina(n32720), .dinb(n32519), .dout(n32721));
  jor  g14699(.dina(n32721), .dinb(n32719), .dout(n32722));
  jand g14700(.dina(n32722), .dinb(n335), .dout(n32723));
  jand g14701(.dina(n32413), .dinb(n32196), .dout(n32724));
  jxor g14702(.dina(n32242), .dinb(n32424), .dout(n32725));
  jand g14703(.dina(n32725), .dinb(n32519), .dout(n32726));
  jor  g14704(.dina(n32726), .dinb(n32724), .dout(n32727));
  jand g14705(.dina(n32727), .dinb(n334), .dout(n32728));
  jand g14706(.dina(n32413), .dinb(n32202), .dout(n32729));
  jxor g14707(.dina(n32238), .dinb(n32422), .dout(n32730));
  jand g14708(.dina(n32730), .dinb(n32519), .dout(n32731));
  jor  g14709(.dina(n32731), .dinb(n32729), .dout(n32732));
  jand g14710(.dina(n32732), .dinb(n338), .dout(n32733));
  jand g14711(.dina(n32413), .dinb(n32208), .dout(n32734));
  jxor g14712(.dina(n32234), .dinb(n32420), .dout(n32735));
  jand g14713(.dina(n32735), .dinb(n32519), .dout(n32736));
  jor  g14714(.dina(n32736), .dinb(n32734), .dout(n32737));
  jand g14715(.dina(n32737), .dinb(n337), .dout(n32738));
  jand g14716(.dina(n32413), .dinb(n32214), .dout(n32739));
  jxor g14717(.dina(n32230), .dinb(n32418), .dout(n32740));
  jand g14718(.dina(n32740), .dinb(n32519), .dout(n32741));
  jor  g14719(.dina(n32741), .dinb(n32739), .dout(n32742));
  jand g14720(.dina(n32742), .dinb(n344), .dout(n32743));
  jand g14721(.dina(n32413), .dinb(n32221), .dout(n32744));
  jxor g14722(.dina(n32416), .dinb(n10855), .dout(n32745));
  jand g14723(.dina(n32745), .dinb(n32519), .dout(n32746));
  jor  g14724(.dina(n32746), .dinb(n32744), .dout(n32747));
  jand g14725(.dina(n32747), .dinb(n348), .dout(n32748));
  jor  g14726(.dina(n32413), .dinb(n18364), .dout(n32749));
  jand g14727(.dina(n32749), .dinb(a16 ), .dout(n32750));
  jor  g14728(.dina(n32413), .dinb(n10855), .dout(n32751));
  jnot g14729(.din(n32751), .dout(n32752));
  jor  g14730(.dina(n32752), .dinb(n32750), .dout(n32753));
  jand g14731(.dina(n32753), .dinb(n258), .dout(n32754));
  jand g14732(.dina(n32519), .dinb(b0 ), .dout(n32755));
  jor  g14733(.dina(n32755), .dinb(n10853), .dout(n32756));
  jand g14734(.dina(n32751), .dinb(n32756), .dout(n32757));
  jxor g14735(.dina(n32757), .dinb(b1 ), .dout(n32758));
  jand g14736(.dina(n32758), .dinb(n11256), .dout(n32759));
  jor  g14737(.dina(n32759), .dinb(n32754), .dout(n32760));
  jxor g14738(.dina(n32747), .dinb(n348), .dout(n32761));
  jand g14739(.dina(n32761), .dinb(n32760), .dout(n32762));
  jor  g14740(.dina(n32762), .dinb(n32748), .dout(n32763));
  jxor g14741(.dina(n32742), .dinb(n344), .dout(n32764));
  jand g14742(.dina(n32764), .dinb(n32763), .dout(n32765));
  jor  g14743(.dina(n32765), .dinb(n32743), .dout(n32766));
  jxor g14744(.dina(n32737), .dinb(n337), .dout(n32767));
  jand g14745(.dina(n32767), .dinb(n32766), .dout(n32768));
  jor  g14746(.dina(n32768), .dinb(n32738), .dout(n32769));
  jxor g14747(.dina(n32732), .dinb(n338), .dout(n32770));
  jand g14748(.dina(n32770), .dinb(n32769), .dout(n32771));
  jor  g14749(.dina(n32771), .dinb(n32733), .dout(n32772));
  jxor g14750(.dina(n32727), .dinb(n334), .dout(n32773));
  jand g14751(.dina(n32773), .dinb(n32772), .dout(n32774));
  jor  g14752(.dina(n32774), .dinb(n32728), .dout(n32775));
  jxor g14753(.dina(n32722), .dinb(n335), .dout(n32776));
  jand g14754(.dina(n32776), .dinb(n32775), .dout(n32777));
  jor  g14755(.dina(n32777), .dinb(n32723), .dout(n32778));
  jxor g14756(.dina(n32717), .dinb(n323), .dout(n32779));
  jand g14757(.dina(n32779), .dinb(n32778), .dout(n32780));
  jor  g14758(.dina(n32780), .dinb(n32718), .dout(n32781));
  jxor g14759(.dina(n32712), .dinb(n324), .dout(n32782));
  jand g14760(.dina(n32782), .dinb(n32781), .dout(n32783));
  jor  g14761(.dina(n32783), .dinb(n32713), .dout(n32784));
  jxor g14762(.dina(n32707), .dinb(n325), .dout(n32785));
  jand g14763(.dina(n32785), .dinb(n32784), .dout(n32786));
  jor  g14764(.dina(n32786), .dinb(n32708), .dout(n32787));
  jxor g14765(.dina(n32702), .dinb(n439), .dout(n32788));
  jand g14766(.dina(n32788), .dinb(n32787), .dout(n32789));
  jor  g14767(.dina(n32789), .dinb(n32703), .dout(n32790));
  jxor g14768(.dina(n32697), .dinb(n440), .dout(n32791));
  jand g14769(.dina(n32791), .dinb(n32790), .dout(n32792));
  jor  g14770(.dina(n32792), .dinb(n32698), .dout(n32793));
  jxor g14771(.dina(n32692), .dinb(n435), .dout(n32794));
  jand g14772(.dina(n32794), .dinb(n32793), .dout(n32795));
  jor  g14773(.dina(n32795), .dinb(n32693), .dout(n32796));
  jxor g14774(.dina(n32687), .dinb(n436), .dout(n32797));
  jand g14775(.dina(n32797), .dinb(n32796), .dout(n32798));
  jor  g14776(.dina(n32798), .dinb(n32688), .dout(n32799));
  jxor g14777(.dina(n32682), .dinb(n432), .dout(n32800));
  jand g14778(.dina(n32800), .dinb(n32799), .dout(n32801));
  jor  g14779(.dina(n32801), .dinb(n32683), .dout(n32802));
  jxor g14780(.dina(n32677), .dinb(n433), .dout(n32803));
  jand g14781(.dina(n32803), .dinb(n32802), .dout(n32804));
  jor  g14782(.dina(n32804), .dinb(n32678), .dout(n32805));
  jxor g14783(.dina(n32672), .dinb(n421), .dout(n32806));
  jand g14784(.dina(n32806), .dinb(n32805), .dout(n32807));
  jor  g14785(.dina(n32807), .dinb(n32673), .dout(n32808));
  jxor g14786(.dina(n32667), .dinb(n422), .dout(n32809));
  jand g14787(.dina(n32809), .dinb(n32808), .dout(n32810));
  jor  g14788(.dina(n32810), .dinb(n32668), .dout(n32811));
  jxor g14789(.dina(n32662), .dinb(n416), .dout(n32812));
  jand g14790(.dina(n32812), .dinb(n32811), .dout(n32813));
  jor  g14791(.dina(n32813), .dinb(n32663), .dout(n32814));
  jxor g14792(.dina(n32657), .dinb(n417), .dout(n32815));
  jand g14793(.dina(n32815), .dinb(n32814), .dout(n32816));
  jor  g14794(.dina(n32816), .dinb(n32658), .dout(n32817));
  jxor g14795(.dina(n32652), .dinb(n2547), .dout(n32818));
  jand g14796(.dina(n32818), .dinb(n32817), .dout(n32819));
  jor  g14797(.dina(n32819), .dinb(n32653), .dout(n32820));
  jxor g14798(.dina(n32647), .dinb(n2714), .dout(n32821));
  jand g14799(.dina(n32821), .dinb(n32820), .dout(n32822));
  jor  g14800(.dina(n32822), .dinb(n32648), .dout(n32823));
  jxor g14801(.dina(n32642), .dinb(n405), .dout(n32824));
  jand g14802(.dina(n32824), .dinb(n32823), .dout(n32825));
  jor  g14803(.dina(n32825), .dinb(n32643), .dout(n32826));
  jxor g14804(.dina(n32637), .dinb(n406), .dout(n32827));
  jand g14805(.dina(n32827), .dinb(n32826), .dout(n32828));
  jor  g14806(.dina(n32828), .dinb(n32638), .dout(n32829));
  jxor g14807(.dina(n32632), .dinb(n412), .dout(n32830));
  jand g14808(.dina(n32830), .dinb(n32829), .dout(n32831));
  jor  g14809(.dina(n32831), .dinb(n32633), .dout(n32832));
  jxor g14810(.dina(n32627), .dinb(n413), .dout(n32833));
  jand g14811(.dina(n32833), .dinb(n32832), .dout(n32834));
  jor  g14812(.dina(n32834), .dinb(n32628), .dout(n32835));
  jxor g14813(.dina(n32622), .dinb(n409), .dout(n32836));
  jand g14814(.dina(n32836), .dinb(n32835), .dout(n32837));
  jor  g14815(.dina(n32837), .dinb(n32623), .dout(n32838));
  jxor g14816(.dina(n32617), .dinb(n410), .dout(n32839));
  jand g14817(.dina(n32839), .dinb(n32838), .dout(n32840));
  jor  g14818(.dina(n32840), .dinb(n32618), .dout(n32841));
  jxor g14819(.dina(n32612), .dinb(n426), .dout(n32842));
  jand g14820(.dina(n32842), .dinb(n32841), .dout(n32843));
  jor  g14821(.dina(n32843), .dinb(n32613), .dout(n32844));
  jxor g14822(.dina(n32607), .dinb(n427), .dout(n32845));
  jand g14823(.dina(n32845), .dinb(n32844), .dout(n32846));
  jor  g14824(.dina(n32846), .dinb(n32608), .dout(n32847));
  jxor g14825(.dina(n32602), .dinb(n424), .dout(n32848));
  jand g14826(.dina(n32848), .dinb(n32847), .dout(n32849));
  jor  g14827(.dina(n32849), .dinb(n32603), .dout(n32850));
  jxor g14828(.dina(n32597), .dinb(n300), .dout(n32851));
  jand g14829(.dina(n32851), .dinb(n32850), .dout(n32852));
  jor  g14830(.dina(n32852), .dinb(n32598), .dout(n32853));
  jxor g14831(.dina(n32592), .dinb(n297), .dout(n32854));
  jand g14832(.dina(n32854), .dinb(n32853), .dout(n32855));
  jor  g14833(.dina(n32855), .dinb(n32593), .dout(n32856));
  jxor g14834(.dina(n32587), .dinb(n298), .dout(n32857));
  jand g14835(.dina(n32857), .dinb(n32856), .dout(n32858));
  jor  g14836(.dina(n32858), .dinb(n32588), .dout(n32859));
  jxor g14837(.dina(n32582), .dinb(n301), .dout(n32860));
  jand g14838(.dina(n32860), .dinb(n32859), .dout(n32861));
  jor  g14839(.dina(n32861), .dinb(n32583), .dout(n32862));
  jxor g14840(.dina(n32577), .dinb(n293), .dout(n32863));
  jand g14841(.dina(n32863), .dinb(n32862), .dout(n32864));
  jor  g14842(.dina(n32864), .dinb(n32578), .dout(n32865));
  jxor g14843(.dina(n32572), .dinb(n294), .dout(n32866));
  jand g14844(.dina(n32866), .dinb(n32865), .dout(n32867));
  jor  g14845(.dina(n32867), .dinb(n32573), .dout(n32868));
  jxor g14846(.dina(n32567), .dinb(n290), .dout(n32869));
  jand g14847(.dina(n32869), .dinb(n32868), .dout(n32870));
  jor  g14848(.dina(n32870), .dinb(n32568), .dout(n32871));
  jxor g14849(.dina(n32562), .dinb(n291), .dout(n32872));
  jand g14850(.dina(n32872), .dinb(n32871), .dout(n32873));
  jor  g14851(.dina(n32873), .dinb(n32563), .dout(n32874));
  jxor g14852(.dina(n32557), .dinb(n284), .dout(n32875));
  jand g14853(.dina(n32875), .dinb(n32874), .dout(n32876));
  jor  g14854(.dina(n32876), .dinb(n32558), .dout(n32877));
  jxor g14855(.dina(n32552), .dinb(n285), .dout(n32878));
  jand g14856(.dina(n32878), .dinb(n32877), .dout(n32879));
  jor  g14857(.dina(n32879), .dinb(n32553), .dout(n32880));
  jxor g14858(.dina(n32547), .dinb(n281), .dout(n32881));
  jand g14859(.dina(n32881), .dinb(n32880), .dout(n32882));
  jor  g14860(.dina(n32882), .dinb(n32548), .dout(n32883));
  jxor g14861(.dina(n32542), .dinb(n282), .dout(n32884));
  jand g14862(.dina(n32884), .dinb(n32883), .dout(n32885));
  jor  g14863(.dina(n32885), .dinb(n32543), .dout(n32886));
  jxor g14864(.dina(n32537), .dinb(n397), .dout(n32887));
  jand g14865(.dina(n32887), .dinb(n32886), .dout(n32888));
  jor  g14866(.dina(n32888), .dinb(n32538), .dout(n32889));
  jxor g14867(.dina(n32532), .dinb(n513), .dout(n32890));
  jand g14868(.dina(n32890), .dinb(n32889), .dout(n32891));
  jor  g14869(.dina(n32891), .dinb(n32533), .dout(n32892));
  jxor g14870(.dina(n32527), .dinb(n514), .dout(n32893));
  jand g14871(.dina(n32893), .dinb(n32892), .dout(n32894));
  jor  g14872(.dina(n32894), .dinb(n32528), .dout(n32895));
  jxor g14873(.dina(n32522), .dinb(n510), .dout(n32896));
  jand g14874(.dina(n32896), .dinb(n32895), .dout(n32897));
  jor  g14875(.dina(n32897), .dinb(n32523), .dout(n32898));
  jand g14876(.dina(n32514), .dinb(b48 ), .dout(n32899));
  jnot g14877(.din(n32899), .dout(n32900));
  jand g14878(.dina(n32900), .dinb(n32898), .dout(n32901));
  jor  g14879(.dina(n32901), .dinb(n32516), .dout(n32902));
  jand g14880(.dina(n32902), .dinb(n387), .dout(n32903));
  jnot g14881(.din(n32903), .dout(n32904));
  jand g14882(.dina(n32904), .dinb(n32515), .dout(n32905));
  jand g14883(.dina(n32516), .dinb(n387), .dout(n32906));
  jand g14884(.dina(n32906), .dinb(n32898), .dout(n32907));
  jor  g14885(.dina(n32907), .dinb(n32905), .dout(n32908));
  jnot g14886(.din(n32908), .dout(n32909));
  jand g14887(.dina(n32904), .dinb(n32522), .dout(n32910));
  jxor g14888(.dina(n32896), .dinb(n32895), .dout(n32911));
  jand g14889(.dina(n32911), .dinb(n32903), .dout(n32912));
  jor  g14890(.dina(n32912), .dinb(n32910), .dout(n32913));
  jand g14891(.dina(n32913), .dinb(n396), .dout(n32914));
  jnot g14892(.din(n32914), .dout(n32915));
  jand g14893(.dina(n32904), .dinb(n32527), .dout(n32916));
  jxor g14894(.dina(n32893), .dinb(n32892), .dout(n32917));
  jand g14895(.dina(n32917), .dinb(n32903), .dout(n32918));
  jor  g14896(.dina(n32918), .dinb(n32916), .dout(n32919));
  jand g14897(.dina(n32919), .dinb(n510), .dout(n32920));
  jnot g14898(.din(n32920), .dout(n32921));
  jand g14899(.dina(n32904), .dinb(n32532), .dout(n32922));
  jxor g14900(.dina(n32890), .dinb(n32889), .dout(n32923));
  jand g14901(.dina(n32923), .dinb(n32903), .dout(n32924));
  jor  g14902(.dina(n32924), .dinb(n32922), .dout(n32925));
  jand g14903(.dina(n32925), .dinb(n514), .dout(n32926));
  jnot g14904(.din(n32926), .dout(n32927));
  jand g14905(.dina(n32904), .dinb(n32537), .dout(n32928));
  jxor g14906(.dina(n32887), .dinb(n32886), .dout(n32929));
  jand g14907(.dina(n32929), .dinb(n32903), .dout(n32930));
  jor  g14908(.dina(n32930), .dinb(n32928), .dout(n32931));
  jand g14909(.dina(n32931), .dinb(n513), .dout(n32932));
  jnot g14910(.din(n32932), .dout(n32933));
  jand g14911(.dina(n32904), .dinb(n32542), .dout(n32934));
  jxor g14912(.dina(n32884), .dinb(n32883), .dout(n32935));
  jand g14913(.dina(n32935), .dinb(n32903), .dout(n32936));
  jor  g14914(.dina(n32936), .dinb(n32934), .dout(n32937));
  jand g14915(.dina(n32937), .dinb(n397), .dout(n32938));
  jnot g14916(.din(n32938), .dout(n32939));
  jand g14917(.dina(n32904), .dinb(n32547), .dout(n32940));
  jxor g14918(.dina(n32881), .dinb(n32880), .dout(n32941));
  jand g14919(.dina(n32941), .dinb(n32903), .dout(n32942));
  jor  g14920(.dina(n32942), .dinb(n32940), .dout(n32943));
  jand g14921(.dina(n32943), .dinb(n282), .dout(n32944));
  jnot g14922(.din(n32944), .dout(n32945));
  jand g14923(.dina(n32904), .dinb(n32552), .dout(n32946));
  jxor g14924(.dina(n32878), .dinb(n32877), .dout(n32947));
  jand g14925(.dina(n32947), .dinb(n32903), .dout(n32948));
  jor  g14926(.dina(n32948), .dinb(n32946), .dout(n32949));
  jand g14927(.dina(n32949), .dinb(n281), .dout(n32950));
  jnot g14928(.din(n32950), .dout(n32951));
  jand g14929(.dina(n32904), .dinb(n32557), .dout(n32952));
  jxor g14930(.dina(n32875), .dinb(n32874), .dout(n32953));
  jand g14931(.dina(n32953), .dinb(n32903), .dout(n32954));
  jor  g14932(.dina(n32954), .dinb(n32952), .dout(n32955));
  jand g14933(.dina(n32955), .dinb(n285), .dout(n32956));
  jnot g14934(.din(n32956), .dout(n32957));
  jand g14935(.dina(n32904), .dinb(n32562), .dout(n32958));
  jxor g14936(.dina(n32872), .dinb(n32871), .dout(n32959));
  jand g14937(.dina(n32959), .dinb(n32903), .dout(n32960));
  jor  g14938(.dina(n32960), .dinb(n32958), .dout(n32961));
  jand g14939(.dina(n32961), .dinb(n284), .dout(n32962));
  jnot g14940(.din(n32962), .dout(n32963));
  jand g14941(.dina(n32904), .dinb(n32567), .dout(n32964));
  jxor g14942(.dina(n32869), .dinb(n32868), .dout(n32965));
  jand g14943(.dina(n32965), .dinb(n32903), .dout(n32966));
  jor  g14944(.dina(n32966), .dinb(n32964), .dout(n32967));
  jand g14945(.dina(n32967), .dinb(n291), .dout(n32968));
  jnot g14946(.din(n32968), .dout(n32969));
  jand g14947(.dina(n32904), .dinb(n32572), .dout(n32970));
  jxor g14948(.dina(n32866), .dinb(n32865), .dout(n32971));
  jand g14949(.dina(n32971), .dinb(n32903), .dout(n32972));
  jor  g14950(.dina(n32972), .dinb(n32970), .dout(n32973));
  jand g14951(.dina(n32973), .dinb(n290), .dout(n32974));
  jnot g14952(.din(n32974), .dout(n32975));
  jand g14953(.dina(n32904), .dinb(n32577), .dout(n32976));
  jxor g14954(.dina(n32863), .dinb(n32862), .dout(n32977));
  jand g14955(.dina(n32977), .dinb(n32903), .dout(n32978));
  jor  g14956(.dina(n32978), .dinb(n32976), .dout(n32979));
  jand g14957(.dina(n32979), .dinb(n294), .dout(n32980));
  jnot g14958(.din(n32980), .dout(n32981));
  jand g14959(.dina(n32904), .dinb(n32582), .dout(n32982));
  jxor g14960(.dina(n32860), .dinb(n32859), .dout(n32983));
  jand g14961(.dina(n32983), .dinb(n32903), .dout(n32984));
  jor  g14962(.dina(n32984), .dinb(n32982), .dout(n32985));
  jand g14963(.dina(n32985), .dinb(n293), .dout(n32986));
  jnot g14964(.din(n32986), .dout(n32987));
  jand g14965(.dina(n32904), .dinb(n32587), .dout(n32988));
  jxor g14966(.dina(n32857), .dinb(n32856), .dout(n32989));
  jand g14967(.dina(n32989), .dinb(n32903), .dout(n32990));
  jor  g14968(.dina(n32990), .dinb(n32988), .dout(n32991));
  jand g14969(.dina(n32991), .dinb(n301), .dout(n32992));
  jnot g14970(.din(n32992), .dout(n32993));
  jand g14971(.dina(n32904), .dinb(n32592), .dout(n32994));
  jxor g14972(.dina(n32854), .dinb(n32853), .dout(n32995));
  jand g14973(.dina(n32995), .dinb(n32903), .dout(n32996));
  jor  g14974(.dina(n32996), .dinb(n32994), .dout(n32997));
  jand g14975(.dina(n32997), .dinb(n298), .dout(n32998));
  jnot g14976(.din(n32998), .dout(n32999));
  jand g14977(.dina(n32904), .dinb(n32597), .dout(n33000));
  jxor g14978(.dina(n32851), .dinb(n32850), .dout(n33001));
  jand g14979(.dina(n33001), .dinb(n32903), .dout(n33002));
  jor  g14980(.dina(n33002), .dinb(n33000), .dout(n33003));
  jand g14981(.dina(n33003), .dinb(n297), .dout(n33004));
  jnot g14982(.din(n33004), .dout(n33005));
  jand g14983(.dina(n32904), .dinb(n32602), .dout(n33006));
  jxor g14984(.dina(n32848), .dinb(n32847), .dout(n33007));
  jand g14985(.dina(n33007), .dinb(n32903), .dout(n33008));
  jor  g14986(.dina(n33008), .dinb(n33006), .dout(n33009));
  jand g14987(.dina(n33009), .dinb(n300), .dout(n33010));
  jnot g14988(.din(n33010), .dout(n33011));
  jand g14989(.dina(n32904), .dinb(n32607), .dout(n33012));
  jxor g14990(.dina(n32845), .dinb(n32844), .dout(n33013));
  jand g14991(.dina(n33013), .dinb(n32903), .dout(n33014));
  jor  g14992(.dina(n33014), .dinb(n33012), .dout(n33015));
  jand g14993(.dina(n33015), .dinb(n424), .dout(n33016));
  jnot g14994(.din(n33016), .dout(n33017));
  jand g14995(.dina(n32904), .dinb(n32612), .dout(n33018));
  jxor g14996(.dina(n32842), .dinb(n32841), .dout(n33019));
  jand g14997(.dina(n33019), .dinb(n32903), .dout(n33020));
  jor  g14998(.dina(n33020), .dinb(n33018), .dout(n33021));
  jand g14999(.dina(n33021), .dinb(n427), .dout(n33022));
  jnot g15000(.din(n33022), .dout(n33023));
  jand g15001(.dina(n32904), .dinb(n32617), .dout(n33024));
  jxor g15002(.dina(n32839), .dinb(n32838), .dout(n33025));
  jand g15003(.dina(n33025), .dinb(n32903), .dout(n33026));
  jor  g15004(.dina(n33026), .dinb(n33024), .dout(n33027));
  jand g15005(.dina(n33027), .dinb(n426), .dout(n33028));
  jnot g15006(.din(n33028), .dout(n33029));
  jand g15007(.dina(n32904), .dinb(n32622), .dout(n33030));
  jxor g15008(.dina(n32836), .dinb(n32835), .dout(n33031));
  jand g15009(.dina(n33031), .dinb(n32903), .dout(n33032));
  jor  g15010(.dina(n33032), .dinb(n33030), .dout(n33033));
  jand g15011(.dina(n33033), .dinb(n410), .dout(n33034));
  jnot g15012(.din(n33034), .dout(n33035));
  jand g15013(.dina(n32904), .dinb(n32627), .dout(n33036));
  jxor g15014(.dina(n32833), .dinb(n32832), .dout(n33037));
  jand g15015(.dina(n33037), .dinb(n32903), .dout(n33038));
  jor  g15016(.dina(n33038), .dinb(n33036), .dout(n33039));
  jand g15017(.dina(n33039), .dinb(n409), .dout(n33040));
  jnot g15018(.din(n33040), .dout(n33041));
  jand g15019(.dina(n32904), .dinb(n32632), .dout(n33042));
  jxor g15020(.dina(n32830), .dinb(n32829), .dout(n33043));
  jand g15021(.dina(n33043), .dinb(n32903), .dout(n33044));
  jor  g15022(.dina(n33044), .dinb(n33042), .dout(n33045));
  jand g15023(.dina(n33045), .dinb(n413), .dout(n33046));
  jnot g15024(.din(n33046), .dout(n33047));
  jand g15025(.dina(n32904), .dinb(n32637), .dout(n33048));
  jxor g15026(.dina(n32827), .dinb(n32826), .dout(n33049));
  jand g15027(.dina(n33049), .dinb(n32903), .dout(n33050));
  jor  g15028(.dina(n33050), .dinb(n33048), .dout(n33051));
  jand g15029(.dina(n33051), .dinb(n412), .dout(n33052));
  jnot g15030(.din(n33052), .dout(n33053));
  jand g15031(.dina(n32904), .dinb(n32642), .dout(n33054));
  jxor g15032(.dina(n32824), .dinb(n32823), .dout(n33055));
  jand g15033(.dina(n33055), .dinb(n32903), .dout(n33056));
  jor  g15034(.dina(n33056), .dinb(n33054), .dout(n33057));
  jand g15035(.dina(n33057), .dinb(n406), .dout(n33058));
  jnot g15036(.din(n33058), .dout(n33059));
  jand g15037(.dina(n32904), .dinb(n32647), .dout(n33060));
  jxor g15038(.dina(n32821), .dinb(n32820), .dout(n33061));
  jand g15039(.dina(n33061), .dinb(n32903), .dout(n33062));
  jor  g15040(.dina(n33062), .dinb(n33060), .dout(n33063));
  jand g15041(.dina(n33063), .dinb(n405), .dout(n33064));
  jnot g15042(.din(n33064), .dout(n33065));
  jand g15043(.dina(n32904), .dinb(n32652), .dout(n33066));
  jxor g15044(.dina(n32818), .dinb(n32817), .dout(n33067));
  jand g15045(.dina(n33067), .dinb(n32903), .dout(n33068));
  jor  g15046(.dina(n33068), .dinb(n33066), .dout(n33069));
  jand g15047(.dina(n33069), .dinb(n2714), .dout(n33070));
  jnot g15048(.din(n33070), .dout(n33071));
  jand g15049(.dina(n32904), .dinb(n32657), .dout(n33072));
  jxor g15050(.dina(n32815), .dinb(n32814), .dout(n33073));
  jand g15051(.dina(n33073), .dinb(n32903), .dout(n33074));
  jor  g15052(.dina(n33074), .dinb(n33072), .dout(n33075));
  jand g15053(.dina(n33075), .dinb(n2547), .dout(n33076));
  jnot g15054(.din(n33076), .dout(n33077));
  jand g15055(.dina(n32904), .dinb(n32662), .dout(n33078));
  jxor g15056(.dina(n32812), .dinb(n32811), .dout(n33079));
  jand g15057(.dina(n33079), .dinb(n32903), .dout(n33080));
  jor  g15058(.dina(n33080), .dinb(n33078), .dout(n33081));
  jand g15059(.dina(n33081), .dinb(n417), .dout(n33082));
  jnot g15060(.din(n33082), .dout(n33083));
  jand g15061(.dina(n32904), .dinb(n32667), .dout(n33084));
  jxor g15062(.dina(n32809), .dinb(n32808), .dout(n33085));
  jand g15063(.dina(n33085), .dinb(n32903), .dout(n33086));
  jor  g15064(.dina(n33086), .dinb(n33084), .dout(n33087));
  jand g15065(.dina(n33087), .dinb(n416), .dout(n33088));
  jnot g15066(.din(n33088), .dout(n33089));
  jand g15067(.dina(n32904), .dinb(n32672), .dout(n33090));
  jxor g15068(.dina(n32806), .dinb(n32805), .dout(n33091));
  jand g15069(.dina(n33091), .dinb(n32903), .dout(n33092));
  jor  g15070(.dina(n33092), .dinb(n33090), .dout(n33093));
  jand g15071(.dina(n33093), .dinb(n422), .dout(n33094));
  jnot g15072(.din(n33094), .dout(n33095));
  jand g15073(.dina(n32904), .dinb(n32677), .dout(n33096));
  jxor g15074(.dina(n32803), .dinb(n32802), .dout(n33097));
  jand g15075(.dina(n33097), .dinb(n32903), .dout(n33098));
  jor  g15076(.dina(n33098), .dinb(n33096), .dout(n33099));
  jand g15077(.dina(n33099), .dinb(n421), .dout(n33100));
  jnot g15078(.din(n33100), .dout(n33101));
  jand g15079(.dina(n32904), .dinb(n32682), .dout(n33102));
  jxor g15080(.dina(n32800), .dinb(n32799), .dout(n33103));
  jand g15081(.dina(n33103), .dinb(n32903), .dout(n33104));
  jor  g15082(.dina(n33104), .dinb(n33102), .dout(n33105));
  jand g15083(.dina(n33105), .dinb(n433), .dout(n33106));
  jnot g15084(.din(n33106), .dout(n33107));
  jand g15085(.dina(n32904), .dinb(n32687), .dout(n33108));
  jxor g15086(.dina(n32797), .dinb(n32796), .dout(n33109));
  jand g15087(.dina(n33109), .dinb(n32903), .dout(n33110));
  jor  g15088(.dina(n33110), .dinb(n33108), .dout(n33111));
  jand g15089(.dina(n33111), .dinb(n432), .dout(n33112));
  jnot g15090(.din(n33112), .dout(n33113));
  jand g15091(.dina(n32904), .dinb(n32692), .dout(n33114));
  jxor g15092(.dina(n32794), .dinb(n32793), .dout(n33115));
  jand g15093(.dina(n33115), .dinb(n32903), .dout(n33116));
  jor  g15094(.dina(n33116), .dinb(n33114), .dout(n33117));
  jand g15095(.dina(n33117), .dinb(n436), .dout(n33118));
  jnot g15096(.din(n33118), .dout(n33119));
  jand g15097(.dina(n32904), .dinb(n32697), .dout(n33120));
  jxor g15098(.dina(n32791), .dinb(n32790), .dout(n33121));
  jand g15099(.dina(n33121), .dinb(n32903), .dout(n33122));
  jor  g15100(.dina(n33122), .dinb(n33120), .dout(n33123));
  jand g15101(.dina(n33123), .dinb(n435), .dout(n33124));
  jnot g15102(.din(n33124), .dout(n33125));
  jand g15103(.dina(n32904), .dinb(n32702), .dout(n33126));
  jxor g15104(.dina(n32788), .dinb(n32787), .dout(n33127));
  jand g15105(.dina(n33127), .dinb(n32903), .dout(n33128));
  jor  g15106(.dina(n33128), .dinb(n33126), .dout(n33129));
  jand g15107(.dina(n33129), .dinb(n440), .dout(n33130));
  jnot g15108(.din(n33130), .dout(n33131));
  jand g15109(.dina(n32904), .dinb(n32707), .dout(n33132));
  jxor g15110(.dina(n32785), .dinb(n32784), .dout(n33133));
  jand g15111(.dina(n33133), .dinb(n32903), .dout(n33134));
  jor  g15112(.dina(n33134), .dinb(n33132), .dout(n33135));
  jand g15113(.dina(n33135), .dinb(n439), .dout(n33136));
  jnot g15114(.din(n33136), .dout(n33137));
  jand g15115(.dina(n32904), .dinb(n32712), .dout(n33138));
  jxor g15116(.dina(n32782), .dinb(n32781), .dout(n33139));
  jand g15117(.dina(n33139), .dinb(n32903), .dout(n33140));
  jor  g15118(.dina(n33140), .dinb(n33138), .dout(n33141));
  jand g15119(.dina(n33141), .dinb(n325), .dout(n33142));
  jnot g15120(.din(n33142), .dout(n33143));
  jand g15121(.dina(n32904), .dinb(n32717), .dout(n33144));
  jxor g15122(.dina(n32779), .dinb(n32778), .dout(n33145));
  jand g15123(.dina(n33145), .dinb(n32903), .dout(n33146));
  jor  g15124(.dina(n33146), .dinb(n33144), .dout(n33147));
  jand g15125(.dina(n33147), .dinb(n324), .dout(n33148));
  jnot g15126(.din(n33148), .dout(n33149));
  jand g15127(.dina(n32904), .dinb(n32722), .dout(n33150));
  jxor g15128(.dina(n32776), .dinb(n32775), .dout(n33151));
  jand g15129(.dina(n33151), .dinb(n32903), .dout(n33152));
  jor  g15130(.dina(n33152), .dinb(n33150), .dout(n33153));
  jand g15131(.dina(n33153), .dinb(n323), .dout(n33154));
  jnot g15132(.din(n33154), .dout(n33155));
  jand g15133(.dina(n32904), .dinb(n32727), .dout(n33156));
  jxor g15134(.dina(n32773), .dinb(n32772), .dout(n33157));
  jand g15135(.dina(n33157), .dinb(n32903), .dout(n33158));
  jor  g15136(.dina(n33158), .dinb(n33156), .dout(n33159));
  jand g15137(.dina(n33159), .dinb(n335), .dout(n33160));
  jnot g15138(.din(n33160), .dout(n33161));
  jand g15139(.dina(n32904), .dinb(n32732), .dout(n33162));
  jxor g15140(.dina(n32770), .dinb(n32769), .dout(n33163));
  jand g15141(.dina(n33163), .dinb(n32903), .dout(n33164));
  jor  g15142(.dina(n33164), .dinb(n33162), .dout(n33165));
  jand g15143(.dina(n33165), .dinb(n334), .dout(n33166));
  jnot g15144(.din(n33166), .dout(n33167));
  jand g15145(.dina(n32904), .dinb(n32737), .dout(n33168));
  jxor g15146(.dina(n32767), .dinb(n32766), .dout(n33169));
  jand g15147(.dina(n33169), .dinb(n32903), .dout(n33170));
  jor  g15148(.dina(n33170), .dinb(n33168), .dout(n33171));
  jand g15149(.dina(n33171), .dinb(n338), .dout(n33172));
  jnot g15150(.din(n33172), .dout(n33173));
  jand g15151(.dina(n32904), .dinb(n32742), .dout(n33174));
  jxor g15152(.dina(n32764), .dinb(n32763), .dout(n33175));
  jand g15153(.dina(n33175), .dinb(n32903), .dout(n33176));
  jor  g15154(.dina(n33176), .dinb(n33174), .dout(n33177));
  jand g15155(.dina(n33177), .dinb(n337), .dout(n33178));
  jnot g15156(.din(n33178), .dout(n33179));
  jnot g15157(.din(n32747), .dout(n33180));
  jor  g15158(.dina(n32903), .dinb(n33180), .dout(n33181));
  jxor g15159(.dina(n32761), .dinb(n32760), .dout(n33182));
  jnot g15160(.din(n33182), .dout(n33183));
  jor  g15161(.dina(n33183), .dinb(n32904), .dout(n33184));
  jand g15162(.dina(n33184), .dinb(n33181), .dout(n33185));
  jnot g15163(.din(n33185), .dout(n33186));
  jand g15164(.dina(n33186), .dinb(n344), .dout(n33187));
  jnot g15165(.din(n33187), .dout(n33188));
  jor  g15166(.dina(n32903), .dinb(n32757), .dout(n33189));
  jxor g15167(.dina(n32758), .dinb(n11256), .dout(n33190));
  jand g15168(.dina(n33190), .dinb(n32903), .dout(n33191));
  jnot g15169(.din(n33191), .dout(n33192));
  jand g15170(.dina(n33192), .dinb(n33189), .dout(n33193));
  jnot g15171(.din(n33193), .dout(n33194));
  jand g15172(.dina(n33194), .dinb(n348), .dout(n33195));
  jnot g15173(.din(n33195), .dout(n33196));
  jnot g15174(.din(n11638), .dout(n33197));
  jnot g15175(.din(n32516), .dout(n33198));
  jnot g15176(.din(n32523), .dout(n33199));
  jnot g15177(.din(n32528), .dout(n33200));
  jnot g15178(.din(n32533), .dout(n33201));
  jnot g15179(.din(n32538), .dout(n33202));
  jnot g15180(.din(n32543), .dout(n33203));
  jnot g15181(.din(n32548), .dout(n33204));
  jnot g15182(.din(n32553), .dout(n33205));
  jnot g15183(.din(n32558), .dout(n33206));
  jnot g15184(.din(n32563), .dout(n33207));
  jnot g15185(.din(n32568), .dout(n33208));
  jnot g15186(.din(n32573), .dout(n33209));
  jnot g15187(.din(n32578), .dout(n33210));
  jnot g15188(.din(n32583), .dout(n33211));
  jnot g15189(.din(n32588), .dout(n33212));
  jnot g15190(.din(n32593), .dout(n33213));
  jnot g15191(.din(n32598), .dout(n33214));
  jnot g15192(.din(n32603), .dout(n33215));
  jnot g15193(.din(n32608), .dout(n33216));
  jnot g15194(.din(n32613), .dout(n33217));
  jnot g15195(.din(n32618), .dout(n33218));
  jnot g15196(.din(n32623), .dout(n33219));
  jnot g15197(.din(n32628), .dout(n33220));
  jnot g15198(.din(n32633), .dout(n33221));
  jnot g15199(.din(n32638), .dout(n33222));
  jnot g15200(.din(n32643), .dout(n33223));
  jnot g15201(.din(n32648), .dout(n33224));
  jnot g15202(.din(n32653), .dout(n33225));
  jnot g15203(.din(n32658), .dout(n33226));
  jnot g15204(.din(n32663), .dout(n33227));
  jnot g15205(.din(n32668), .dout(n33228));
  jnot g15206(.din(n32673), .dout(n33229));
  jnot g15207(.din(n32678), .dout(n33230));
  jnot g15208(.din(n32683), .dout(n33231));
  jnot g15209(.din(n32688), .dout(n33232));
  jnot g15210(.din(n32693), .dout(n33233));
  jnot g15211(.din(n32698), .dout(n33234));
  jnot g15212(.din(n32703), .dout(n33235));
  jnot g15213(.din(n32708), .dout(n33236));
  jnot g15214(.din(n32713), .dout(n33237));
  jnot g15215(.din(n32718), .dout(n33238));
  jnot g15216(.din(n32723), .dout(n33239));
  jnot g15217(.din(n32728), .dout(n33240));
  jnot g15218(.din(n32733), .dout(n33241));
  jnot g15219(.din(n32738), .dout(n33242));
  jnot g15220(.din(n32743), .dout(n33243));
  jnot g15221(.din(n32748), .dout(n33244));
  jnot g15222(.din(n32754), .dout(n33245));
  jxor g15223(.dina(n32757), .dinb(n258), .dout(n33246));
  jor  g15224(.dina(n33246), .dinb(n11255), .dout(n33247));
  jand g15225(.dina(n33247), .dinb(n33245), .dout(n33248));
  jnot g15226(.din(n32761), .dout(n33249));
  jor  g15227(.dina(n33249), .dinb(n33248), .dout(n33250));
  jand g15228(.dina(n33250), .dinb(n33244), .dout(n33251));
  jnot g15229(.din(n32764), .dout(n33252));
  jor  g15230(.dina(n33252), .dinb(n33251), .dout(n33253));
  jand g15231(.dina(n33253), .dinb(n33243), .dout(n33254));
  jnot g15232(.din(n32767), .dout(n33255));
  jor  g15233(.dina(n33255), .dinb(n33254), .dout(n33256));
  jand g15234(.dina(n33256), .dinb(n33242), .dout(n33257));
  jnot g15235(.din(n32770), .dout(n33258));
  jor  g15236(.dina(n33258), .dinb(n33257), .dout(n33259));
  jand g15237(.dina(n33259), .dinb(n33241), .dout(n33260));
  jnot g15238(.din(n32773), .dout(n33261));
  jor  g15239(.dina(n33261), .dinb(n33260), .dout(n33262));
  jand g15240(.dina(n33262), .dinb(n33240), .dout(n33263));
  jnot g15241(.din(n32776), .dout(n33264));
  jor  g15242(.dina(n33264), .dinb(n33263), .dout(n33265));
  jand g15243(.dina(n33265), .dinb(n33239), .dout(n33266));
  jnot g15244(.din(n32779), .dout(n33267));
  jor  g15245(.dina(n33267), .dinb(n33266), .dout(n33268));
  jand g15246(.dina(n33268), .dinb(n33238), .dout(n33269));
  jnot g15247(.din(n32782), .dout(n33270));
  jor  g15248(.dina(n33270), .dinb(n33269), .dout(n33271));
  jand g15249(.dina(n33271), .dinb(n33237), .dout(n33272));
  jnot g15250(.din(n32785), .dout(n33273));
  jor  g15251(.dina(n33273), .dinb(n33272), .dout(n33274));
  jand g15252(.dina(n33274), .dinb(n33236), .dout(n33275));
  jnot g15253(.din(n32788), .dout(n33276));
  jor  g15254(.dina(n33276), .dinb(n33275), .dout(n33277));
  jand g15255(.dina(n33277), .dinb(n33235), .dout(n33278));
  jnot g15256(.din(n32791), .dout(n33279));
  jor  g15257(.dina(n33279), .dinb(n33278), .dout(n33280));
  jand g15258(.dina(n33280), .dinb(n33234), .dout(n33281));
  jnot g15259(.din(n32794), .dout(n33282));
  jor  g15260(.dina(n33282), .dinb(n33281), .dout(n33283));
  jand g15261(.dina(n33283), .dinb(n33233), .dout(n33284));
  jnot g15262(.din(n32797), .dout(n33285));
  jor  g15263(.dina(n33285), .dinb(n33284), .dout(n33286));
  jand g15264(.dina(n33286), .dinb(n33232), .dout(n33287));
  jnot g15265(.din(n32800), .dout(n33288));
  jor  g15266(.dina(n33288), .dinb(n33287), .dout(n33289));
  jand g15267(.dina(n33289), .dinb(n33231), .dout(n33290));
  jnot g15268(.din(n32803), .dout(n33291));
  jor  g15269(.dina(n33291), .dinb(n33290), .dout(n33292));
  jand g15270(.dina(n33292), .dinb(n33230), .dout(n33293));
  jnot g15271(.din(n32806), .dout(n33294));
  jor  g15272(.dina(n33294), .dinb(n33293), .dout(n33295));
  jand g15273(.dina(n33295), .dinb(n33229), .dout(n33296));
  jnot g15274(.din(n32809), .dout(n33297));
  jor  g15275(.dina(n33297), .dinb(n33296), .dout(n33298));
  jand g15276(.dina(n33298), .dinb(n33228), .dout(n33299));
  jnot g15277(.din(n32812), .dout(n33300));
  jor  g15278(.dina(n33300), .dinb(n33299), .dout(n33301));
  jand g15279(.dina(n33301), .dinb(n33227), .dout(n33302));
  jnot g15280(.din(n32815), .dout(n33303));
  jor  g15281(.dina(n33303), .dinb(n33302), .dout(n33304));
  jand g15282(.dina(n33304), .dinb(n33226), .dout(n33305));
  jnot g15283(.din(n32818), .dout(n33306));
  jor  g15284(.dina(n33306), .dinb(n33305), .dout(n33307));
  jand g15285(.dina(n33307), .dinb(n33225), .dout(n33308));
  jnot g15286(.din(n32821), .dout(n33309));
  jor  g15287(.dina(n33309), .dinb(n33308), .dout(n33310));
  jand g15288(.dina(n33310), .dinb(n33224), .dout(n33311));
  jnot g15289(.din(n32824), .dout(n33312));
  jor  g15290(.dina(n33312), .dinb(n33311), .dout(n33313));
  jand g15291(.dina(n33313), .dinb(n33223), .dout(n33314));
  jnot g15292(.din(n32827), .dout(n33315));
  jor  g15293(.dina(n33315), .dinb(n33314), .dout(n33316));
  jand g15294(.dina(n33316), .dinb(n33222), .dout(n33317));
  jnot g15295(.din(n32830), .dout(n33318));
  jor  g15296(.dina(n33318), .dinb(n33317), .dout(n33319));
  jand g15297(.dina(n33319), .dinb(n33221), .dout(n33320));
  jnot g15298(.din(n32833), .dout(n33321));
  jor  g15299(.dina(n33321), .dinb(n33320), .dout(n33322));
  jand g15300(.dina(n33322), .dinb(n33220), .dout(n33323));
  jnot g15301(.din(n32836), .dout(n33324));
  jor  g15302(.dina(n33324), .dinb(n33323), .dout(n33325));
  jand g15303(.dina(n33325), .dinb(n33219), .dout(n33326));
  jnot g15304(.din(n32839), .dout(n33327));
  jor  g15305(.dina(n33327), .dinb(n33326), .dout(n33328));
  jand g15306(.dina(n33328), .dinb(n33218), .dout(n33329));
  jnot g15307(.din(n32842), .dout(n33330));
  jor  g15308(.dina(n33330), .dinb(n33329), .dout(n33331));
  jand g15309(.dina(n33331), .dinb(n33217), .dout(n33332));
  jnot g15310(.din(n32845), .dout(n33333));
  jor  g15311(.dina(n33333), .dinb(n33332), .dout(n33334));
  jand g15312(.dina(n33334), .dinb(n33216), .dout(n33335));
  jnot g15313(.din(n32848), .dout(n33336));
  jor  g15314(.dina(n33336), .dinb(n33335), .dout(n33337));
  jand g15315(.dina(n33337), .dinb(n33215), .dout(n33338));
  jnot g15316(.din(n32851), .dout(n33339));
  jor  g15317(.dina(n33339), .dinb(n33338), .dout(n33340));
  jand g15318(.dina(n33340), .dinb(n33214), .dout(n33341));
  jnot g15319(.din(n32854), .dout(n33342));
  jor  g15320(.dina(n33342), .dinb(n33341), .dout(n33343));
  jand g15321(.dina(n33343), .dinb(n33213), .dout(n33344));
  jnot g15322(.din(n32857), .dout(n33345));
  jor  g15323(.dina(n33345), .dinb(n33344), .dout(n33346));
  jand g15324(.dina(n33346), .dinb(n33212), .dout(n33347));
  jnot g15325(.din(n32860), .dout(n33348));
  jor  g15326(.dina(n33348), .dinb(n33347), .dout(n33349));
  jand g15327(.dina(n33349), .dinb(n33211), .dout(n33350));
  jnot g15328(.din(n32863), .dout(n33351));
  jor  g15329(.dina(n33351), .dinb(n33350), .dout(n33352));
  jand g15330(.dina(n33352), .dinb(n33210), .dout(n33353));
  jnot g15331(.din(n32866), .dout(n33354));
  jor  g15332(.dina(n33354), .dinb(n33353), .dout(n33355));
  jand g15333(.dina(n33355), .dinb(n33209), .dout(n33356));
  jnot g15334(.din(n32869), .dout(n33357));
  jor  g15335(.dina(n33357), .dinb(n33356), .dout(n33358));
  jand g15336(.dina(n33358), .dinb(n33208), .dout(n33359));
  jnot g15337(.din(n32872), .dout(n33360));
  jor  g15338(.dina(n33360), .dinb(n33359), .dout(n33361));
  jand g15339(.dina(n33361), .dinb(n33207), .dout(n33362));
  jnot g15340(.din(n32875), .dout(n33363));
  jor  g15341(.dina(n33363), .dinb(n33362), .dout(n33364));
  jand g15342(.dina(n33364), .dinb(n33206), .dout(n33365));
  jnot g15343(.din(n32878), .dout(n33366));
  jor  g15344(.dina(n33366), .dinb(n33365), .dout(n33367));
  jand g15345(.dina(n33367), .dinb(n33205), .dout(n33368));
  jnot g15346(.din(n32881), .dout(n33369));
  jor  g15347(.dina(n33369), .dinb(n33368), .dout(n33370));
  jand g15348(.dina(n33370), .dinb(n33204), .dout(n33371));
  jnot g15349(.din(n32884), .dout(n33372));
  jor  g15350(.dina(n33372), .dinb(n33371), .dout(n33373));
  jand g15351(.dina(n33373), .dinb(n33203), .dout(n33374));
  jnot g15352(.din(n32887), .dout(n33375));
  jor  g15353(.dina(n33375), .dinb(n33374), .dout(n33376));
  jand g15354(.dina(n33376), .dinb(n33202), .dout(n33377));
  jnot g15355(.din(n32890), .dout(n33378));
  jor  g15356(.dina(n33378), .dinb(n33377), .dout(n33379));
  jand g15357(.dina(n33379), .dinb(n33201), .dout(n33380));
  jnot g15358(.din(n32893), .dout(n33381));
  jor  g15359(.dina(n33381), .dinb(n33380), .dout(n33382));
  jand g15360(.dina(n33382), .dinb(n33200), .dout(n33383));
  jnot g15361(.din(n32896), .dout(n33384));
  jor  g15362(.dina(n33384), .dinb(n33383), .dout(n33385));
  jand g15363(.dina(n33385), .dinb(n33199), .dout(n33386));
  jor  g15364(.dina(n32899), .dinb(n33386), .dout(n33387));
  jand g15365(.dina(n33387), .dinb(n33198), .dout(n33388));
  jor  g15366(.dina(n33388), .dinb(n33197), .dout(n33389));
  jand g15367(.dina(n33389), .dinb(a15 ), .dout(n33390));
  jnot g15368(.din(n11641), .dout(n33391));
  jor  g15369(.dina(n33388), .dinb(n33391), .dout(n33392));
  jnot g15370(.din(n33392), .dout(n33393));
  jor  g15371(.dina(n33393), .dinb(n33390), .dout(n33394));
  jand g15372(.dina(n33394), .dinb(n258), .dout(n33395));
  jnot g15373(.din(n33395), .dout(n33396));
  jand g15374(.dina(n32902), .dinb(n11638), .dout(n33397));
  jor  g15375(.dina(n33397), .dinb(n11254), .dout(n33398));
  jand g15376(.dina(n33392), .dinb(n33398), .dout(n33399));
  jxor g15377(.dina(n33399), .dinb(n258), .dout(n33400));
  jor  g15378(.dina(n33400), .dinb(n11648), .dout(n33401));
  jand g15379(.dina(n33401), .dinb(n33396), .dout(n33402));
  jxor g15380(.dina(n33193), .dinb(b2 ), .dout(n33403));
  jnot g15381(.din(n33403), .dout(n33404));
  jor  g15382(.dina(n33404), .dinb(n33402), .dout(n33405));
  jand g15383(.dina(n33405), .dinb(n33196), .dout(n33406));
  jxor g15384(.dina(n33185), .dinb(b3 ), .dout(n33407));
  jnot g15385(.din(n33407), .dout(n33408));
  jor  g15386(.dina(n33408), .dinb(n33406), .dout(n33409));
  jand g15387(.dina(n33409), .dinb(n33188), .dout(n33410));
  jxor g15388(.dina(n33177), .dinb(n337), .dout(n33411));
  jnot g15389(.din(n33411), .dout(n33412));
  jor  g15390(.dina(n33412), .dinb(n33410), .dout(n33413));
  jand g15391(.dina(n33413), .dinb(n33179), .dout(n33414));
  jxor g15392(.dina(n33171), .dinb(n338), .dout(n33415));
  jnot g15393(.din(n33415), .dout(n33416));
  jor  g15394(.dina(n33416), .dinb(n33414), .dout(n33417));
  jand g15395(.dina(n33417), .dinb(n33173), .dout(n33418));
  jxor g15396(.dina(n33165), .dinb(n334), .dout(n33419));
  jnot g15397(.din(n33419), .dout(n33420));
  jor  g15398(.dina(n33420), .dinb(n33418), .dout(n33421));
  jand g15399(.dina(n33421), .dinb(n33167), .dout(n33422));
  jxor g15400(.dina(n33159), .dinb(n335), .dout(n33423));
  jnot g15401(.din(n33423), .dout(n33424));
  jor  g15402(.dina(n33424), .dinb(n33422), .dout(n33425));
  jand g15403(.dina(n33425), .dinb(n33161), .dout(n33426));
  jxor g15404(.dina(n33153), .dinb(n323), .dout(n33427));
  jnot g15405(.din(n33427), .dout(n33428));
  jor  g15406(.dina(n33428), .dinb(n33426), .dout(n33429));
  jand g15407(.dina(n33429), .dinb(n33155), .dout(n33430));
  jxor g15408(.dina(n33147), .dinb(n324), .dout(n33431));
  jnot g15409(.din(n33431), .dout(n33432));
  jor  g15410(.dina(n33432), .dinb(n33430), .dout(n33433));
  jand g15411(.dina(n33433), .dinb(n33149), .dout(n33434));
  jxor g15412(.dina(n33141), .dinb(n325), .dout(n33435));
  jnot g15413(.din(n33435), .dout(n33436));
  jor  g15414(.dina(n33436), .dinb(n33434), .dout(n33437));
  jand g15415(.dina(n33437), .dinb(n33143), .dout(n33438));
  jxor g15416(.dina(n33135), .dinb(n439), .dout(n33439));
  jnot g15417(.din(n33439), .dout(n33440));
  jor  g15418(.dina(n33440), .dinb(n33438), .dout(n33441));
  jand g15419(.dina(n33441), .dinb(n33137), .dout(n33442));
  jxor g15420(.dina(n33129), .dinb(n440), .dout(n33443));
  jnot g15421(.din(n33443), .dout(n33444));
  jor  g15422(.dina(n33444), .dinb(n33442), .dout(n33445));
  jand g15423(.dina(n33445), .dinb(n33131), .dout(n33446));
  jxor g15424(.dina(n33123), .dinb(n435), .dout(n33447));
  jnot g15425(.din(n33447), .dout(n33448));
  jor  g15426(.dina(n33448), .dinb(n33446), .dout(n33449));
  jand g15427(.dina(n33449), .dinb(n33125), .dout(n33450));
  jxor g15428(.dina(n33117), .dinb(n436), .dout(n33451));
  jnot g15429(.din(n33451), .dout(n33452));
  jor  g15430(.dina(n33452), .dinb(n33450), .dout(n33453));
  jand g15431(.dina(n33453), .dinb(n33119), .dout(n33454));
  jxor g15432(.dina(n33111), .dinb(n432), .dout(n33455));
  jnot g15433(.din(n33455), .dout(n33456));
  jor  g15434(.dina(n33456), .dinb(n33454), .dout(n33457));
  jand g15435(.dina(n33457), .dinb(n33113), .dout(n33458));
  jxor g15436(.dina(n33105), .dinb(n433), .dout(n33459));
  jnot g15437(.din(n33459), .dout(n33460));
  jor  g15438(.dina(n33460), .dinb(n33458), .dout(n33461));
  jand g15439(.dina(n33461), .dinb(n33107), .dout(n33462));
  jxor g15440(.dina(n33099), .dinb(n421), .dout(n33463));
  jnot g15441(.din(n33463), .dout(n33464));
  jor  g15442(.dina(n33464), .dinb(n33462), .dout(n33465));
  jand g15443(.dina(n33465), .dinb(n33101), .dout(n33466));
  jxor g15444(.dina(n33093), .dinb(n422), .dout(n33467));
  jnot g15445(.din(n33467), .dout(n33468));
  jor  g15446(.dina(n33468), .dinb(n33466), .dout(n33469));
  jand g15447(.dina(n33469), .dinb(n33095), .dout(n33470));
  jxor g15448(.dina(n33087), .dinb(n416), .dout(n33471));
  jnot g15449(.din(n33471), .dout(n33472));
  jor  g15450(.dina(n33472), .dinb(n33470), .dout(n33473));
  jand g15451(.dina(n33473), .dinb(n33089), .dout(n33474));
  jxor g15452(.dina(n33081), .dinb(n417), .dout(n33475));
  jnot g15453(.din(n33475), .dout(n33476));
  jor  g15454(.dina(n33476), .dinb(n33474), .dout(n33477));
  jand g15455(.dina(n33477), .dinb(n33083), .dout(n33478));
  jxor g15456(.dina(n33075), .dinb(n2547), .dout(n33479));
  jnot g15457(.din(n33479), .dout(n33480));
  jor  g15458(.dina(n33480), .dinb(n33478), .dout(n33481));
  jand g15459(.dina(n33481), .dinb(n33077), .dout(n33482));
  jxor g15460(.dina(n33069), .dinb(n2714), .dout(n33483));
  jnot g15461(.din(n33483), .dout(n33484));
  jor  g15462(.dina(n33484), .dinb(n33482), .dout(n33485));
  jand g15463(.dina(n33485), .dinb(n33071), .dout(n33486));
  jxor g15464(.dina(n33063), .dinb(n405), .dout(n33487));
  jnot g15465(.din(n33487), .dout(n33488));
  jor  g15466(.dina(n33488), .dinb(n33486), .dout(n33489));
  jand g15467(.dina(n33489), .dinb(n33065), .dout(n33490));
  jxor g15468(.dina(n33057), .dinb(n406), .dout(n33491));
  jnot g15469(.din(n33491), .dout(n33492));
  jor  g15470(.dina(n33492), .dinb(n33490), .dout(n33493));
  jand g15471(.dina(n33493), .dinb(n33059), .dout(n33494));
  jxor g15472(.dina(n33051), .dinb(n412), .dout(n33495));
  jnot g15473(.din(n33495), .dout(n33496));
  jor  g15474(.dina(n33496), .dinb(n33494), .dout(n33497));
  jand g15475(.dina(n33497), .dinb(n33053), .dout(n33498));
  jxor g15476(.dina(n33045), .dinb(n413), .dout(n33499));
  jnot g15477(.din(n33499), .dout(n33500));
  jor  g15478(.dina(n33500), .dinb(n33498), .dout(n33501));
  jand g15479(.dina(n33501), .dinb(n33047), .dout(n33502));
  jxor g15480(.dina(n33039), .dinb(n409), .dout(n33503));
  jnot g15481(.din(n33503), .dout(n33504));
  jor  g15482(.dina(n33504), .dinb(n33502), .dout(n33505));
  jand g15483(.dina(n33505), .dinb(n33041), .dout(n33506));
  jxor g15484(.dina(n33033), .dinb(n410), .dout(n33507));
  jnot g15485(.din(n33507), .dout(n33508));
  jor  g15486(.dina(n33508), .dinb(n33506), .dout(n33509));
  jand g15487(.dina(n33509), .dinb(n33035), .dout(n33510));
  jxor g15488(.dina(n33027), .dinb(n426), .dout(n33511));
  jnot g15489(.din(n33511), .dout(n33512));
  jor  g15490(.dina(n33512), .dinb(n33510), .dout(n33513));
  jand g15491(.dina(n33513), .dinb(n33029), .dout(n33514));
  jxor g15492(.dina(n33021), .dinb(n427), .dout(n33515));
  jnot g15493(.din(n33515), .dout(n33516));
  jor  g15494(.dina(n33516), .dinb(n33514), .dout(n33517));
  jand g15495(.dina(n33517), .dinb(n33023), .dout(n33518));
  jxor g15496(.dina(n33015), .dinb(n424), .dout(n33519));
  jnot g15497(.din(n33519), .dout(n33520));
  jor  g15498(.dina(n33520), .dinb(n33518), .dout(n33521));
  jand g15499(.dina(n33521), .dinb(n33017), .dout(n33522));
  jxor g15500(.dina(n33009), .dinb(n300), .dout(n33523));
  jnot g15501(.din(n33523), .dout(n33524));
  jor  g15502(.dina(n33524), .dinb(n33522), .dout(n33525));
  jand g15503(.dina(n33525), .dinb(n33011), .dout(n33526));
  jxor g15504(.dina(n33003), .dinb(n297), .dout(n33527));
  jnot g15505(.din(n33527), .dout(n33528));
  jor  g15506(.dina(n33528), .dinb(n33526), .dout(n33529));
  jand g15507(.dina(n33529), .dinb(n33005), .dout(n33530));
  jxor g15508(.dina(n32997), .dinb(n298), .dout(n33531));
  jnot g15509(.din(n33531), .dout(n33532));
  jor  g15510(.dina(n33532), .dinb(n33530), .dout(n33533));
  jand g15511(.dina(n33533), .dinb(n32999), .dout(n33534));
  jxor g15512(.dina(n32991), .dinb(n301), .dout(n33535));
  jnot g15513(.din(n33535), .dout(n33536));
  jor  g15514(.dina(n33536), .dinb(n33534), .dout(n33537));
  jand g15515(.dina(n33537), .dinb(n32993), .dout(n33538));
  jxor g15516(.dina(n32985), .dinb(n293), .dout(n33539));
  jnot g15517(.din(n33539), .dout(n33540));
  jor  g15518(.dina(n33540), .dinb(n33538), .dout(n33541));
  jand g15519(.dina(n33541), .dinb(n32987), .dout(n33542));
  jxor g15520(.dina(n32979), .dinb(n294), .dout(n33543));
  jnot g15521(.din(n33543), .dout(n33544));
  jor  g15522(.dina(n33544), .dinb(n33542), .dout(n33545));
  jand g15523(.dina(n33545), .dinb(n32981), .dout(n33546));
  jxor g15524(.dina(n32973), .dinb(n290), .dout(n33547));
  jnot g15525(.din(n33547), .dout(n33548));
  jor  g15526(.dina(n33548), .dinb(n33546), .dout(n33549));
  jand g15527(.dina(n33549), .dinb(n32975), .dout(n33550));
  jxor g15528(.dina(n32967), .dinb(n291), .dout(n33551));
  jnot g15529(.din(n33551), .dout(n33552));
  jor  g15530(.dina(n33552), .dinb(n33550), .dout(n33553));
  jand g15531(.dina(n33553), .dinb(n32969), .dout(n33554));
  jxor g15532(.dina(n32961), .dinb(n284), .dout(n33555));
  jnot g15533(.din(n33555), .dout(n33556));
  jor  g15534(.dina(n33556), .dinb(n33554), .dout(n33557));
  jand g15535(.dina(n33557), .dinb(n32963), .dout(n33558));
  jxor g15536(.dina(n32955), .dinb(n285), .dout(n33559));
  jnot g15537(.din(n33559), .dout(n33560));
  jor  g15538(.dina(n33560), .dinb(n33558), .dout(n33561));
  jand g15539(.dina(n33561), .dinb(n32957), .dout(n33562));
  jxor g15540(.dina(n32949), .dinb(n281), .dout(n33563));
  jnot g15541(.din(n33563), .dout(n33564));
  jor  g15542(.dina(n33564), .dinb(n33562), .dout(n33565));
  jand g15543(.dina(n33565), .dinb(n32951), .dout(n33566));
  jxor g15544(.dina(n32943), .dinb(n282), .dout(n33567));
  jnot g15545(.din(n33567), .dout(n33568));
  jor  g15546(.dina(n33568), .dinb(n33566), .dout(n33569));
  jand g15547(.dina(n33569), .dinb(n32945), .dout(n33570));
  jxor g15548(.dina(n32937), .dinb(n397), .dout(n33571));
  jnot g15549(.din(n33571), .dout(n33572));
  jor  g15550(.dina(n33572), .dinb(n33570), .dout(n33573));
  jand g15551(.dina(n33573), .dinb(n32939), .dout(n33574));
  jxor g15552(.dina(n32931), .dinb(n513), .dout(n33575));
  jnot g15553(.din(n33575), .dout(n33576));
  jor  g15554(.dina(n33576), .dinb(n33574), .dout(n33577));
  jand g15555(.dina(n33577), .dinb(n32933), .dout(n33578));
  jxor g15556(.dina(n32925), .dinb(n514), .dout(n33579));
  jnot g15557(.din(n33579), .dout(n33580));
  jor  g15558(.dina(n33580), .dinb(n33578), .dout(n33581));
  jand g15559(.dina(n33581), .dinb(n32927), .dout(n33582));
  jxor g15560(.dina(n32919), .dinb(n510), .dout(n33583));
  jnot g15561(.din(n33583), .dout(n33584));
  jor  g15562(.dina(n33584), .dinb(n33582), .dout(n33585));
  jand g15563(.dina(n33585), .dinb(n32921), .dout(n33586));
  jxor g15564(.dina(n32913), .dinb(n396), .dout(n33587));
  jnot g15565(.din(n33587), .dout(n33588));
  jor  g15566(.dina(n33588), .dinb(n33586), .dout(n33589));
  jand g15567(.dina(n33589), .dinb(n32915), .dout(n33590));
  jxor g15568(.dina(n32908), .dinb(b49 ), .dout(n33591));
  jor  g15569(.dina(n33591), .dinb(n11794), .dout(n33592));
  jor  g15570(.dina(n33592), .dinb(n33590), .dout(n33593));
  jand g15571(.dina(n33593), .dinb(n32909), .dout(n33594));
  jxor g15572(.dina(n33399), .dinb(b1 ), .dout(n33595));
  jand g15573(.dina(n33595), .dinb(n11649), .dout(n33596));
  jor  g15574(.dina(n33596), .dinb(n33395), .dout(n33597));
  jand g15575(.dina(n33403), .dinb(n33597), .dout(n33598));
  jor  g15576(.dina(n33598), .dinb(n33195), .dout(n33599));
  jand g15577(.dina(n33407), .dinb(n33599), .dout(n33600));
  jor  g15578(.dina(n33600), .dinb(n33187), .dout(n33601));
  jand g15579(.dina(n33411), .dinb(n33601), .dout(n33602));
  jor  g15580(.dina(n33602), .dinb(n33178), .dout(n33603));
  jand g15581(.dina(n33415), .dinb(n33603), .dout(n33604));
  jor  g15582(.dina(n33604), .dinb(n33172), .dout(n33605));
  jand g15583(.dina(n33419), .dinb(n33605), .dout(n33606));
  jor  g15584(.dina(n33606), .dinb(n33166), .dout(n33607));
  jand g15585(.dina(n33423), .dinb(n33607), .dout(n33608));
  jor  g15586(.dina(n33608), .dinb(n33160), .dout(n33609));
  jand g15587(.dina(n33427), .dinb(n33609), .dout(n33610));
  jor  g15588(.dina(n33610), .dinb(n33154), .dout(n33611));
  jand g15589(.dina(n33431), .dinb(n33611), .dout(n33612));
  jor  g15590(.dina(n33612), .dinb(n33148), .dout(n33613));
  jand g15591(.dina(n33435), .dinb(n33613), .dout(n33614));
  jor  g15592(.dina(n33614), .dinb(n33142), .dout(n33615));
  jand g15593(.dina(n33439), .dinb(n33615), .dout(n33616));
  jor  g15594(.dina(n33616), .dinb(n33136), .dout(n33617));
  jand g15595(.dina(n33443), .dinb(n33617), .dout(n33618));
  jor  g15596(.dina(n33618), .dinb(n33130), .dout(n33619));
  jand g15597(.dina(n33447), .dinb(n33619), .dout(n33620));
  jor  g15598(.dina(n33620), .dinb(n33124), .dout(n33621));
  jand g15599(.dina(n33451), .dinb(n33621), .dout(n33622));
  jor  g15600(.dina(n33622), .dinb(n33118), .dout(n33623));
  jand g15601(.dina(n33455), .dinb(n33623), .dout(n33624));
  jor  g15602(.dina(n33624), .dinb(n33112), .dout(n33625));
  jand g15603(.dina(n33459), .dinb(n33625), .dout(n33626));
  jor  g15604(.dina(n33626), .dinb(n33106), .dout(n33627));
  jand g15605(.dina(n33463), .dinb(n33627), .dout(n33628));
  jor  g15606(.dina(n33628), .dinb(n33100), .dout(n33629));
  jand g15607(.dina(n33467), .dinb(n33629), .dout(n33630));
  jor  g15608(.dina(n33630), .dinb(n33094), .dout(n33631));
  jand g15609(.dina(n33471), .dinb(n33631), .dout(n33632));
  jor  g15610(.dina(n33632), .dinb(n33088), .dout(n33633));
  jand g15611(.dina(n33475), .dinb(n33633), .dout(n33634));
  jor  g15612(.dina(n33634), .dinb(n33082), .dout(n33635));
  jand g15613(.dina(n33479), .dinb(n33635), .dout(n33636));
  jor  g15614(.dina(n33636), .dinb(n33076), .dout(n33637));
  jand g15615(.dina(n33483), .dinb(n33637), .dout(n33638));
  jor  g15616(.dina(n33638), .dinb(n33070), .dout(n33639));
  jand g15617(.dina(n33487), .dinb(n33639), .dout(n33640));
  jor  g15618(.dina(n33640), .dinb(n33064), .dout(n33641));
  jand g15619(.dina(n33491), .dinb(n33641), .dout(n33642));
  jor  g15620(.dina(n33642), .dinb(n33058), .dout(n33643));
  jand g15621(.dina(n33495), .dinb(n33643), .dout(n33644));
  jor  g15622(.dina(n33644), .dinb(n33052), .dout(n33645));
  jand g15623(.dina(n33499), .dinb(n33645), .dout(n33646));
  jor  g15624(.dina(n33646), .dinb(n33046), .dout(n33647));
  jand g15625(.dina(n33503), .dinb(n33647), .dout(n33648));
  jor  g15626(.dina(n33648), .dinb(n33040), .dout(n33649));
  jand g15627(.dina(n33507), .dinb(n33649), .dout(n33650));
  jor  g15628(.dina(n33650), .dinb(n33034), .dout(n33651));
  jand g15629(.dina(n33511), .dinb(n33651), .dout(n33652));
  jor  g15630(.dina(n33652), .dinb(n33028), .dout(n33653));
  jand g15631(.dina(n33515), .dinb(n33653), .dout(n33654));
  jor  g15632(.dina(n33654), .dinb(n33022), .dout(n33655));
  jand g15633(.dina(n33519), .dinb(n33655), .dout(n33656));
  jor  g15634(.dina(n33656), .dinb(n33016), .dout(n33657));
  jand g15635(.dina(n33523), .dinb(n33657), .dout(n33658));
  jor  g15636(.dina(n33658), .dinb(n33010), .dout(n33659));
  jand g15637(.dina(n33527), .dinb(n33659), .dout(n33660));
  jor  g15638(.dina(n33660), .dinb(n33004), .dout(n33661));
  jand g15639(.dina(n33531), .dinb(n33661), .dout(n33662));
  jor  g15640(.dina(n33662), .dinb(n32998), .dout(n33663));
  jand g15641(.dina(n33535), .dinb(n33663), .dout(n33664));
  jor  g15642(.dina(n33664), .dinb(n32992), .dout(n33665));
  jand g15643(.dina(n33539), .dinb(n33665), .dout(n33666));
  jor  g15644(.dina(n33666), .dinb(n32986), .dout(n33667));
  jand g15645(.dina(n33543), .dinb(n33667), .dout(n33668));
  jor  g15646(.dina(n33668), .dinb(n32980), .dout(n33669));
  jand g15647(.dina(n33547), .dinb(n33669), .dout(n33670));
  jor  g15648(.dina(n33670), .dinb(n32974), .dout(n33671));
  jand g15649(.dina(n33551), .dinb(n33671), .dout(n33672));
  jor  g15650(.dina(n33672), .dinb(n32968), .dout(n33673));
  jand g15651(.dina(n33555), .dinb(n33673), .dout(n33674));
  jor  g15652(.dina(n33674), .dinb(n32962), .dout(n33675));
  jand g15653(.dina(n33559), .dinb(n33675), .dout(n33676));
  jor  g15654(.dina(n33676), .dinb(n32956), .dout(n33677));
  jand g15655(.dina(n33563), .dinb(n33677), .dout(n33678));
  jor  g15656(.dina(n33678), .dinb(n32950), .dout(n33679));
  jand g15657(.dina(n33567), .dinb(n33679), .dout(n33680));
  jor  g15658(.dina(n33680), .dinb(n32944), .dout(n33681));
  jand g15659(.dina(n33571), .dinb(n33681), .dout(n33682));
  jor  g15660(.dina(n33682), .dinb(n32938), .dout(n33683));
  jand g15661(.dina(n33575), .dinb(n33683), .dout(n33684));
  jor  g15662(.dina(n33684), .dinb(n32932), .dout(n33685));
  jand g15663(.dina(n33579), .dinb(n33685), .dout(n33686));
  jor  g15664(.dina(n33686), .dinb(n32926), .dout(n33687));
  jand g15665(.dina(n33583), .dinb(n33687), .dout(n33688));
  jor  g15666(.dina(n33688), .dinb(n32920), .dout(n33689));
  jand g15667(.dina(n33587), .dinb(n33689), .dout(n33690));
  jor  g15668(.dina(n33690), .dinb(n32914), .dout(n33691));
  jnot g15669(.din(n33592), .dout(n33692));
  jand g15670(.dina(n33692), .dinb(n33691), .dout(n33693));
  jand g15671(.dina(n32908), .dinb(n387), .dout(n33694));
  jor  g15672(.dina(n33694), .dinb(n33693), .dout(n33695));
  jxor g15673(.dina(n33591), .dinb(n33691), .dout(n33696));
  jand g15674(.dina(n33696), .dinb(n33695), .dout(n33697));
  jor  g15675(.dina(n33697), .dinb(n33594), .dout(n33698));
  jnot g15676(.din(n33694), .dout(n33699));
  jand g15677(.dina(n33699), .dinb(n33593), .dout(n33700));
  jand g15678(.dina(n33700), .dinb(n32913), .dout(n33701));
  jxor g15679(.dina(n33587), .dinb(n33689), .dout(n33702));
  jand g15680(.dina(n33702), .dinb(n33695), .dout(n33703));
  jor  g15681(.dina(n33703), .dinb(n33701), .dout(n33704));
  jand g15682(.dina(n33704), .dinb(n383), .dout(n33705));
  jnot g15683(.din(n33705), .dout(n33706));
  jand g15684(.dina(n33700), .dinb(n32919), .dout(n33707));
  jxor g15685(.dina(n33583), .dinb(n33687), .dout(n33708));
  jand g15686(.dina(n33708), .dinb(n33695), .dout(n33709));
  jor  g15687(.dina(n33709), .dinb(n33707), .dout(n33710));
  jand g15688(.dina(n33710), .dinb(n396), .dout(n33711));
  jnot g15689(.din(n33711), .dout(n33712));
  jand g15690(.dina(n33700), .dinb(n32925), .dout(n33713));
  jxor g15691(.dina(n33579), .dinb(n33685), .dout(n33714));
  jand g15692(.dina(n33714), .dinb(n33695), .dout(n33715));
  jor  g15693(.dina(n33715), .dinb(n33713), .dout(n33716));
  jand g15694(.dina(n33716), .dinb(n510), .dout(n33717));
  jnot g15695(.din(n33717), .dout(n33718));
  jand g15696(.dina(n33700), .dinb(n32931), .dout(n33719));
  jxor g15697(.dina(n33575), .dinb(n33683), .dout(n33720));
  jand g15698(.dina(n33720), .dinb(n33695), .dout(n33721));
  jor  g15699(.dina(n33721), .dinb(n33719), .dout(n33722));
  jand g15700(.dina(n33722), .dinb(n514), .dout(n33723));
  jnot g15701(.din(n33723), .dout(n33724));
  jand g15702(.dina(n33700), .dinb(n32937), .dout(n33725));
  jxor g15703(.dina(n33571), .dinb(n33681), .dout(n33726));
  jand g15704(.dina(n33726), .dinb(n33695), .dout(n33727));
  jor  g15705(.dina(n33727), .dinb(n33725), .dout(n33728));
  jand g15706(.dina(n33728), .dinb(n513), .dout(n33729));
  jnot g15707(.din(n33729), .dout(n33730));
  jand g15708(.dina(n33700), .dinb(n32943), .dout(n33731));
  jxor g15709(.dina(n33567), .dinb(n33679), .dout(n33732));
  jand g15710(.dina(n33732), .dinb(n33695), .dout(n33733));
  jor  g15711(.dina(n33733), .dinb(n33731), .dout(n33734));
  jand g15712(.dina(n33734), .dinb(n397), .dout(n33735));
  jnot g15713(.din(n33735), .dout(n33736));
  jand g15714(.dina(n33700), .dinb(n32949), .dout(n33737));
  jxor g15715(.dina(n33563), .dinb(n33677), .dout(n33738));
  jand g15716(.dina(n33738), .dinb(n33695), .dout(n33739));
  jor  g15717(.dina(n33739), .dinb(n33737), .dout(n33740));
  jand g15718(.dina(n33740), .dinb(n282), .dout(n33741));
  jnot g15719(.din(n33741), .dout(n33742));
  jand g15720(.dina(n33700), .dinb(n32955), .dout(n33743));
  jxor g15721(.dina(n33559), .dinb(n33675), .dout(n33744));
  jand g15722(.dina(n33744), .dinb(n33695), .dout(n33745));
  jor  g15723(.dina(n33745), .dinb(n33743), .dout(n33746));
  jand g15724(.dina(n33746), .dinb(n281), .dout(n33747));
  jnot g15725(.din(n33747), .dout(n33748));
  jand g15726(.dina(n33700), .dinb(n32961), .dout(n33749));
  jxor g15727(.dina(n33555), .dinb(n33673), .dout(n33750));
  jand g15728(.dina(n33750), .dinb(n33695), .dout(n33751));
  jor  g15729(.dina(n33751), .dinb(n33749), .dout(n33752));
  jand g15730(.dina(n33752), .dinb(n285), .dout(n33753));
  jnot g15731(.din(n33753), .dout(n33754));
  jand g15732(.dina(n33700), .dinb(n32967), .dout(n33755));
  jxor g15733(.dina(n33551), .dinb(n33671), .dout(n33756));
  jand g15734(.dina(n33756), .dinb(n33695), .dout(n33757));
  jor  g15735(.dina(n33757), .dinb(n33755), .dout(n33758));
  jand g15736(.dina(n33758), .dinb(n284), .dout(n33759));
  jnot g15737(.din(n33759), .dout(n33760));
  jand g15738(.dina(n33700), .dinb(n32973), .dout(n33761));
  jxor g15739(.dina(n33547), .dinb(n33669), .dout(n33762));
  jand g15740(.dina(n33762), .dinb(n33695), .dout(n33763));
  jor  g15741(.dina(n33763), .dinb(n33761), .dout(n33764));
  jand g15742(.dina(n33764), .dinb(n291), .dout(n33765));
  jnot g15743(.din(n33765), .dout(n33766));
  jand g15744(.dina(n33700), .dinb(n32979), .dout(n33767));
  jxor g15745(.dina(n33543), .dinb(n33667), .dout(n33768));
  jand g15746(.dina(n33768), .dinb(n33695), .dout(n33769));
  jor  g15747(.dina(n33769), .dinb(n33767), .dout(n33770));
  jand g15748(.dina(n33770), .dinb(n290), .dout(n33771));
  jnot g15749(.din(n33771), .dout(n33772));
  jand g15750(.dina(n33700), .dinb(n32985), .dout(n33773));
  jxor g15751(.dina(n33539), .dinb(n33665), .dout(n33774));
  jand g15752(.dina(n33774), .dinb(n33695), .dout(n33775));
  jor  g15753(.dina(n33775), .dinb(n33773), .dout(n33776));
  jand g15754(.dina(n33776), .dinb(n294), .dout(n33777));
  jnot g15755(.din(n33777), .dout(n33778));
  jand g15756(.dina(n33700), .dinb(n32991), .dout(n33779));
  jxor g15757(.dina(n33535), .dinb(n33663), .dout(n33780));
  jand g15758(.dina(n33780), .dinb(n33695), .dout(n33781));
  jor  g15759(.dina(n33781), .dinb(n33779), .dout(n33782));
  jand g15760(.dina(n33782), .dinb(n293), .dout(n33783));
  jnot g15761(.din(n33783), .dout(n33784));
  jand g15762(.dina(n33700), .dinb(n32997), .dout(n33785));
  jxor g15763(.dina(n33531), .dinb(n33661), .dout(n33786));
  jand g15764(.dina(n33786), .dinb(n33695), .dout(n33787));
  jor  g15765(.dina(n33787), .dinb(n33785), .dout(n33788));
  jand g15766(.dina(n33788), .dinb(n301), .dout(n33789));
  jnot g15767(.din(n33789), .dout(n33790));
  jand g15768(.dina(n33700), .dinb(n33003), .dout(n33791));
  jxor g15769(.dina(n33527), .dinb(n33659), .dout(n33792));
  jand g15770(.dina(n33792), .dinb(n33695), .dout(n33793));
  jor  g15771(.dina(n33793), .dinb(n33791), .dout(n33794));
  jand g15772(.dina(n33794), .dinb(n298), .dout(n33795));
  jnot g15773(.din(n33795), .dout(n33796));
  jand g15774(.dina(n33700), .dinb(n33009), .dout(n33797));
  jxor g15775(.dina(n33523), .dinb(n33657), .dout(n33798));
  jand g15776(.dina(n33798), .dinb(n33695), .dout(n33799));
  jor  g15777(.dina(n33799), .dinb(n33797), .dout(n33800));
  jand g15778(.dina(n33800), .dinb(n297), .dout(n33801));
  jnot g15779(.din(n33801), .dout(n33802));
  jand g15780(.dina(n33700), .dinb(n33015), .dout(n33803));
  jxor g15781(.dina(n33519), .dinb(n33655), .dout(n33804));
  jand g15782(.dina(n33804), .dinb(n33695), .dout(n33805));
  jor  g15783(.dina(n33805), .dinb(n33803), .dout(n33806));
  jand g15784(.dina(n33806), .dinb(n300), .dout(n33807));
  jnot g15785(.din(n33807), .dout(n33808));
  jand g15786(.dina(n33700), .dinb(n33021), .dout(n33809));
  jxor g15787(.dina(n33515), .dinb(n33653), .dout(n33810));
  jand g15788(.dina(n33810), .dinb(n33695), .dout(n33811));
  jor  g15789(.dina(n33811), .dinb(n33809), .dout(n33812));
  jand g15790(.dina(n33812), .dinb(n424), .dout(n33813));
  jnot g15791(.din(n33813), .dout(n33814));
  jand g15792(.dina(n33700), .dinb(n33027), .dout(n33815));
  jxor g15793(.dina(n33511), .dinb(n33651), .dout(n33816));
  jand g15794(.dina(n33816), .dinb(n33695), .dout(n33817));
  jor  g15795(.dina(n33817), .dinb(n33815), .dout(n33818));
  jand g15796(.dina(n33818), .dinb(n427), .dout(n33819));
  jnot g15797(.din(n33819), .dout(n33820));
  jand g15798(.dina(n33700), .dinb(n33033), .dout(n33821));
  jxor g15799(.dina(n33507), .dinb(n33649), .dout(n33822));
  jand g15800(.dina(n33822), .dinb(n33695), .dout(n33823));
  jor  g15801(.dina(n33823), .dinb(n33821), .dout(n33824));
  jand g15802(.dina(n33824), .dinb(n426), .dout(n33825));
  jnot g15803(.din(n33825), .dout(n33826));
  jand g15804(.dina(n33700), .dinb(n33039), .dout(n33827));
  jxor g15805(.dina(n33503), .dinb(n33647), .dout(n33828));
  jand g15806(.dina(n33828), .dinb(n33695), .dout(n33829));
  jor  g15807(.dina(n33829), .dinb(n33827), .dout(n33830));
  jand g15808(.dina(n33830), .dinb(n410), .dout(n33831));
  jnot g15809(.din(n33831), .dout(n33832));
  jand g15810(.dina(n33700), .dinb(n33045), .dout(n33833));
  jxor g15811(.dina(n33499), .dinb(n33645), .dout(n33834));
  jand g15812(.dina(n33834), .dinb(n33695), .dout(n33835));
  jor  g15813(.dina(n33835), .dinb(n33833), .dout(n33836));
  jand g15814(.dina(n33836), .dinb(n409), .dout(n33837));
  jnot g15815(.din(n33837), .dout(n33838));
  jand g15816(.dina(n33700), .dinb(n33051), .dout(n33839));
  jxor g15817(.dina(n33495), .dinb(n33643), .dout(n33840));
  jand g15818(.dina(n33840), .dinb(n33695), .dout(n33841));
  jor  g15819(.dina(n33841), .dinb(n33839), .dout(n33842));
  jand g15820(.dina(n33842), .dinb(n413), .dout(n33843));
  jnot g15821(.din(n33843), .dout(n33844));
  jand g15822(.dina(n33700), .dinb(n33057), .dout(n33845));
  jxor g15823(.dina(n33491), .dinb(n33641), .dout(n33846));
  jand g15824(.dina(n33846), .dinb(n33695), .dout(n33847));
  jor  g15825(.dina(n33847), .dinb(n33845), .dout(n33848));
  jand g15826(.dina(n33848), .dinb(n412), .dout(n33849));
  jnot g15827(.din(n33849), .dout(n33850));
  jand g15828(.dina(n33700), .dinb(n33063), .dout(n33851));
  jxor g15829(.dina(n33487), .dinb(n33639), .dout(n33852));
  jand g15830(.dina(n33852), .dinb(n33695), .dout(n33853));
  jor  g15831(.dina(n33853), .dinb(n33851), .dout(n33854));
  jand g15832(.dina(n33854), .dinb(n406), .dout(n33855));
  jnot g15833(.din(n33855), .dout(n33856));
  jand g15834(.dina(n33700), .dinb(n33069), .dout(n33857));
  jxor g15835(.dina(n33483), .dinb(n33637), .dout(n33858));
  jand g15836(.dina(n33858), .dinb(n33695), .dout(n33859));
  jor  g15837(.dina(n33859), .dinb(n33857), .dout(n33860));
  jand g15838(.dina(n33860), .dinb(n405), .dout(n33861));
  jnot g15839(.din(n33861), .dout(n33862));
  jand g15840(.dina(n33700), .dinb(n33075), .dout(n33863));
  jxor g15841(.dina(n33479), .dinb(n33635), .dout(n33864));
  jand g15842(.dina(n33864), .dinb(n33695), .dout(n33865));
  jor  g15843(.dina(n33865), .dinb(n33863), .dout(n33866));
  jand g15844(.dina(n33866), .dinb(n2714), .dout(n33867));
  jnot g15845(.din(n33867), .dout(n33868));
  jand g15846(.dina(n33700), .dinb(n33081), .dout(n33869));
  jxor g15847(.dina(n33475), .dinb(n33633), .dout(n33870));
  jand g15848(.dina(n33870), .dinb(n33695), .dout(n33871));
  jor  g15849(.dina(n33871), .dinb(n33869), .dout(n33872));
  jand g15850(.dina(n33872), .dinb(n2547), .dout(n33873));
  jnot g15851(.din(n33873), .dout(n33874));
  jand g15852(.dina(n33700), .dinb(n33087), .dout(n33875));
  jxor g15853(.dina(n33471), .dinb(n33631), .dout(n33876));
  jand g15854(.dina(n33876), .dinb(n33695), .dout(n33877));
  jor  g15855(.dina(n33877), .dinb(n33875), .dout(n33878));
  jand g15856(.dina(n33878), .dinb(n417), .dout(n33879));
  jnot g15857(.din(n33879), .dout(n33880));
  jand g15858(.dina(n33700), .dinb(n33093), .dout(n33881));
  jxor g15859(.dina(n33467), .dinb(n33629), .dout(n33882));
  jand g15860(.dina(n33882), .dinb(n33695), .dout(n33883));
  jor  g15861(.dina(n33883), .dinb(n33881), .dout(n33884));
  jand g15862(.dina(n33884), .dinb(n416), .dout(n33885));
  jnot g15863(.din(n33885), .dout(n33886));
  jand g15864(.dina(n33700), .dinb(n33099), .dout(n33887));
  jxor g15865(.dina(n33463), .dinb(n33627), .dout(n33888));
  jand g15866(.dina(n33888), .dinb(n33695), .dout(n33889));
  jor  g15867(.dina(n33889), .dinb(n33887), .dout(n33890));
  jand g15868(.dina(n33890), .dinb(n422), .dout(n33891));
  jnot g15869(.din(n33891), .dout(n33892));
  jand g15870(.dina(n33700), .dinb(n33105), .dout(n33893));
  jxor g15871(.dina(n33459), .dinb(n33625), .dout(n33894));
  jand g15872(.dina(n33894), .dinb(n33695), .dout(n33895));
  jor  g15873(.dina(n33895), .dinb(n33893), .dout(n33896));
  jand g15874(.dina(n33896), .dinb(n421), .dout(n33897));
  jnot g15875(.din(n33897), .dout(n33898));
  jand g15876(.dina(n33700), .dinb(n33111), .dout(n33899));
  jxor g15877(.dina(n33455), .dinb(n33623), .dout(n33900));
  jand g15878(.dina(n33900), .dinb(n33695), .dout(n33901));
  jor  g15879(.dina(n33901), .dinb(n33899), .dout(n33902));
  jand g15880(.dina(n33902), .dinb(n433), .dout(n33903));
  jnot g15881(.din(n33903), .dout(n33904));
  jand g15882(.dina(n33700), .dinb(n33117), .dout(n33905));
  jxor g15883(.dina(n33451), .dinb(n33621), .dout(n33906));
  jand g15884(.dina(n33906), .dinb(n33695), .dout(n33907));
  jor  g15885(.dina(n33907), .dinb(n33905), .dout(n33908));
  jand g15886(.dina(n33908), .dinb(n432), .dout(n33909));
  jnot g15887(.din(n33909), .dout(n33910));
  jand g15888(.dina(n33700), .dinb(n33123), .dout(n33911));
  jxor g15889(.dina(n33447), .dinb(n33619), .dout(n33912));
  jand g15890(.dina(n33912), .dinb(n33695), .dout(n33913));
  jor  g15891(.dina(n33913), .dinb(n33911), .dout(n33914));
  jand g15892(.dina(n33914), .dinb(n436), .dout(n33915));
  jnot g15893(.din(n33915), .dout(n33916));
  jand g15894(.dina(n33700), .dinb(n33129), .dout(n33917));
  jxor g15895(.dina(n33443), .dinb(n33617), .dout(n33918));
  jand g15896(.dina(n33918), .dinb(n33695), .dout(n33919));
  jor  g15897(.dina(n33919), .dinb(n33917), .dout(n33920));
  jand g15898(.dina(n33920), .dinb(n435), .dout(n33921));
  jnot g15899(.din(n33921), .dout(n33922));
  jand g15900(.dina(n33700), .dinb(n33135), .dout(n33923));
  jxor g15901(.dina(n33439), .dinb(n33615), .dout(n33924));
  jand g15902(.dina(n33924), .dinb(n33695), .dout(n33925));
  jor  g15903(.dina(n33925), .dinb(n33923), .dout(n33926));
  jand g15904(.dina(n33926), .dinb(n440), .dout(n33927));
  jnot g15905(.din(n33927), .dout(n33928));
  jand g15906(.dina(n33700), .dinb(n33141), .dout(n33929));
  jxor g15907(.dina(n33435), .dinb(n33613), .dout(n33930));
  jand g15908(.dina(n33930), .dinb(n33695), .dout(n33931));
  jor  g15909(.dina(n33931), .dinb(n33929), .dout(n33932));
  jand g15910(.dina(n33932), .dinb(n439), .dout(n33933));
  jnot g15911(.din(n33933), .dout(n33934));
  jand g15912(.dina(n33700), .dinb(n33147), .dout(n33935));
  jxor g15913(.dina(n33431), .dinb(n33611), .dout(n33936));
  jand g15914(.dina(n33936), .dinb(n33695), .dout(n33937));
  jor  g15915(.dina(n33937), .dinb(n33935), .dout(n33938));
  jand g15916(.dina(n33938), .dinb(n325), .dout(n33939));
  jnot g15917(.din(n33939), .dout(n33940));
  jand g15918(.dina(n33700), .dinb(n33153), .dout(n33941));
  jxor g15919(.dina(n33427), .dinb(n33609), .dout(n33942));
  jand g15920(.dina(n33942), .dinb(n33695), .dout(n33943));
  jor  g15921(.dina(n33943), .dinb(n33941), .dout(n33944));
  jand g15922(.dina(n33944), .dinb(n324), .dout(n33945));
  jnot g15923(.din(n33945), .dout(n33946));
  jand g15924(.dina(n33700), .dinb(n33159), .dout(n33947));
  jxor g15925(.dina(n33423), .dinb(n33607), .dout(n33948));
  jand g15926(.dina(n33948), .dinb(n33695), .dout(n33949));
  jor  g15927(.dina(n33949), .dinb(n33947), .dout(n33950));
  jand g15928(.dina(n33950), .dinb(n323), .dout(n33951));
  jnot g15929(.din(n33951), .dout(n33952));
  jand g15930(.dina(n33700), .dinb(n33165), .dout(n33953));
  jxor g15931(.dina(n33419), .dinb(n33605), .dout(n33954));
  jand g15932(.dina(n33954), .dinb(n33695), .dout(n33955));
  jor  g15933(.dina(n33955), .dinb(n33953), .dout(n33956));
  jand g15934(.dina(n33956), .dinb(n335), .dout(n33957));
  jnot g15935(.din(n33957), .dout(n33958));
  jand g15936(.dina(n33700), .dinb(n33171), .dout(n33959));
  jxor g15937(.dina(n33415), .dinb(n33603), .dout(n33960));
  jand g15938(.dina(n33960), .dinb(n33695), .dout(n33961));
  jor  g15939(.dina(n33961), .dinb(n33959), .dout(n33962));
  jand g15940(.dina(n33962), .dinb(n334), .dout(n33963));
  jnot g15941(.din(n33963), .dout(n33964));
  jand g15942(.dina(n33700), .dinb(n33177), .dout(n33965));
  jxor g15943(.dina(n33411), .dinb(n33601), .dout(n33966));
  jand g15944(.dina(n33966), .dinb(n33695), .dout(n33967));
  jor  g15945(.dina(n33967), .dinb(n33965), .dout(n33968));
  jand g15946(.dina(n33968), .dinb(n338), .dout(n33969));
  jnot g15947(.din(n33969), .dout(n33970));
  jand g15948(.dina(n33700), .dinb(n33186), .dout(n33971));
  jxor g15949(.dina(n33407), .dinb(n33599), .dout(n33972));
  jand g15950(.dina(n33972), .dinb(n33695), .dout(n33973));
  jor  g15951(.dina(n33973), .dinb(n33971), .dout(n33974));
  jand g15952(.dina(n33974), .dinb(n337), .dout(n33975));
  jnot g15953(.din(n33975), .dout(n33976));
  jand g15954(.dina(n33700), .dinb(n33194), .dout(n33977));
  jxor g15955(.dina(n33403), .dinb(n33597), .dout(n33978));
  jand g15956(.dina(n33978), .dinb(n33695), .dout(n33979));
  jor  g15957(.dina(n33979), .dinb(n33977), .dout(n33980));
  jand g15958(.dina(n33980), .dinb(n344), .dout(n33981));
  jnot g15959(.din(n33981), .dout(n33982));
  jand g15960(.dina(n33700), .dinb(n33394), .dout(n33983));
  jxor g15961(.dina(n33595), .dinb(n11649), .dout(n33984));
  jand g15962(.dina(n33984), .dinb(n33695), .dout(n33985));
  jor  g15963(.dina(n33985), .dinb(n33983), .dout(n33986));
  jand g15964(.dina(n33986), .dinb(n348), .dout(n33987));
  jnot g15965(.din(n33987), .dout(n33988));
  jor  g15966(.dina(n33700), .dinb(n18364), .dout(n33989));
  jand g15967(.dina(n33989), .dinb(a14 ), .dout(n33990));
  jor  g15968(.dina(n33700), .dinb(n11649), .dout(n33991));
  jnot g15969(.din(n33991), .dout(n33992));
  jor  g15970(.dina(n33992), .dinb(n33990), .dout(n33993));
  jand g15971(.dina(n33993), .dinb(n258), .dout(n33994));
  jnot g15972(.din(n33994), .dout(n33995));
  jand g15973(.dina(n33695), .dinb(b0 ), .dout(n33996));
  jor  g15974(.dina(n33996), .dinb(n11647), .dout(n33997));
  jand g15975(.dina(n33991), .dinb(n33997), .dout(n33998));
  jxor g15976(.dina(n33998), .dinb(n258), .dout(n33999));
  jor  g15977(.dina(n33999), .dinb(n12062), .dout(n34000));
  jand g15978(.dina(n34000), .dinb(n33995), .dout(n34001));
  jxor g15979(.dina(n33986), .dinb(n348), .dout(n34002));
  jnot g15980(.din(n34002), .dout(n34003));
  jor  g15981(.dina(n34003), .dinb(n34001), .dout(n34004));
  jand g15982(.dina(n34004), .dinb(n33988), .dout(n34005));
  jxor g15983(.dina(n33980), .dinb(n344), .dout(n34006));
  jnot g15984(.din(n34006), .dout(n34007));
  jor  g15985(.dina(n34007), .dinb(n34005), .dout(n34008));
  jand g15986(.dina(n34008), .dinb(n33982), .dout(n34009));
  jxor g15987(.dina(n33974), .dinb(n337), .dout(n34010));
  jnot g15988(.din(n34010), .dout(n34011));
  jor  g15989(.dina(n34011), .dinb(n34009), .dout(n34012));
  jand g15990(.dina(n34012), .dinb(n33976), .dout(n34013));
  jxor g15991(.dina(n33968), .dinb(n338), .dout(n34014));
  jnot g15992(.din(n34014), .dout(n34015));
  jor  g15993(.dina(n34015), .dinb(n34013), .dout(n34016));
  jand g15994(.dina(n34016), .dinb(n33970), .dout(n34017));
  jxor g15995(.dina(n33962), .dinb(n334), .dout(n34018));
  jnot g15996(.din(n34018), .dout(n34019));
  jor  g15997(.dina(n34019), .dinb(n34017), .dout(n34020));
  jand g15998(.dina(n34020), .dinb(n33964), .dout(n34021));
  jxor g15999(.dina(n33956), .dinb(n335), .dout(n34022));
  jnot g16000(.din(n34022), .dout(n34023));
  jor  g16001(.dina(n34023), .dinb(n34021), .dout(n34024));
  jand g16002(.dina(n34024), .dinb(n33958), .dout(n34025));
  jxor g16003(.dina(n33950), .dinb(n323), .dout(n34026));
  jnot g16004(.din(n34026), .dout(n34027));
  jor  g16005(.dina(n34027), .dinb(n34025), .dout(n34028));
  jand g16006(.dina(n34028), .dinb(n33952), .dout(n34029));
  jxor g16007(.dina(n33944), .dinb(n324), .dout(n34030));
  jnot g16008(.din(n34030), .dout(n34031));
  jor  g16009(.dina(n34031), .dinb(n34029), .dout(n34032));
  jand g16010(.dina(n34032), .dinb(n33946), .dout(n34033));
  jxor g16011(.dina(n33938), .dinb(n325), .dout(n34034));
  jnot g16012(.din(n34034), .dout(n34035));
  jor  g16013(.dina(n34035), .dinb(n34033), .dout(n34036));
  jand g16014(.dina(n34036), .dinb(n33940), .dout(n34037));
  jxor g16015(.dina(n33932), .dinb(n439), .dout(n34038));
  jnot g16016(.din(n34038), .dout(n34039));
  jor  g16017(.dina(n34039), .dinb(n34037), .dout(n34040));
  jand g16018(.dina(n34040), .dinb(n33934), .dout(n34041));
  jxor g16019(.dina(n33926), .dinb(n440), .dout(n34042));
  jnot g16020(.din(n34042), .dout(n34043));
  jor  g16021(.dina(n34043), .dinb(n34041), .dout(n34044));
  jand g16022(.dina(n34044), .dinb(n33928), .dout(n34045));
  jxor g16023(.dina(n33920), .dinb(n435), .dout(n34046));
  jnot g16024(.din(n34046), .dout(n34047));
  jor  g16025(.dina(n34047), .dinb(n34045), .dout(n34048));
  jand g16026(.dina(n34048), .dinb(n33922), .dout(n34049));
  jxor g16027(.dina(n33914), .dinb(n436), .dout(n34050));
  jnot g16028(.din(n34050), .dout(n34051));
  jor  g16029(.dina(n34051), .dinb(n34049), .dout(n34052));
  jand g16030(.dina(n34052), .dinb(n33916), .dout(n34053));
  jxor g16031(.dina(n33908), .dinb(n432), .dout(n34054));
  jnot g16032(.din(n34054), .dout(n34055));
  jor  g16033(.dina(n34055), .dinb(n34053), .dout(n34056));
  jand g16034(.dina(n34056), .dinb(n33910), .dout(n34057));
  jxor g16035(.dina(n33902), .dinb(n433), .dout(n34058));
  jnot g16036(.din(n34058), .dout(n34059));
  jor  g16037(.dina(n34059), .dinb(n34057), .dout(n34060));
  jand g16038(.dina(n34060), .dinb(n33904), .dout(n34061));
  jxor g16039(.dina(n33896), .dinb(n421), .dout(n34062));
  jnot g16040(.din(n34062), .dout(n34063));
  jor  g16041(.dina(n34063), .dinb(n34061), .dout(n34064));
  jand g16042(.dina(n34064), .dinb(n33898), .dout(n34065));
  jxor g16043(.dina(n33890), .dinb(n422), .dout(n34066));
  jnot g16044(.din(n34066), .dout(n34067));
  jor  g16045(.dina(n34067), .dinb(n34065), .dout(n34068));
  jand g16046(.dina(n34068), .dinb(n33892), .dout(n34069));
  jxor g16047(.dina(n33884), .dinb(n416), .dout(n34070));
  jnot g16048(.din(n34070), .dout(n34071));
  jor  g16049(.dina(n34071), .dinb(n34069), .dout(n34072));
  jand g16050(.dina(n34072), .dinb(n33886), .dout(n34073));
  jxor g16051(.dina(n33878), .dinb(n417), .dout(n34074));
  jnot g16052(.din(n34074), .dout(n34075));
  jor  g16053(.dina(n34075), .dinb(n34073), .dout(n34076));
  jand g16054(.dina(n34076), .dinb(n33880), .dout(n34077));
  jxor g16055(.dina(n33872), .dinb(n2547), .dout(n34078));
  jnot g16056(.din(n34078), .dout(n34079));
  jor  g16057(.dina(n34079), .dinb(n34077), .dout(n34080));
  jand g16058(.dina(n34080), .dinb(n33874), .dout(n34081));
  jxor g16059(.dina(n33866), .dinb(n2714), .dout(n34082));
  jnot g16060(.din(n34082), .dout(n34083));
  jor  g16061(.dina(n34083), .dinb(n34081), .dout(n34084));
  jand g16062(.dina(n34084), .dinb(n33868), .dout(n34085));
  jxor g16063(.dina(n33860), .dinb(n405), .dout(n34086));
  jnot g16064(.din(n34086), .dout(n34087));
  jor  g16065(.dina(n34087), .dinb(n34085), .dout(n34088));
  jand g16066(.dina(n34088), .dinb(n33862), .dout(n34089));
  jxor g16067(.dina(n33854), .dinb(n406), .dout(n34090));
  jnot g16068(.din(n34090), .dout(n34091));
  jor  g16069(.dina(n34091), .dinb(n34089), .dout(n34092));
  jand g16070(.dina(n34092), .dinb(n33856), .dout(n34093));
  jxor g16071(.dina(n33848), .dinb(n412), .dout(n34094));
  jnot g16072(.din(n34094), .dout(n34095));
  jor  g16073(.dina(n34095), .dinb(n34093), .dout(n34096));
  jand g16074(.dina(n34096), .dinb(n33850), .dout(n34097));
  jxor g16075(.dina(n33842), .dinb(n413), .dout(n34098));
  jnot g16076(.din(n34098), .dout(n34099));
  jor  g16077(.dina(n34099), .dinb(n34097), .dout(n34100));
  jand g16078(.dina(n34100), .dinb(n33844), .dout(n34101));
  jxor g16079(.dina(n33836), .dinb(n409), .dout(n34102));
  jnot g16080(.din(n34102), .dout(n34103));
  jor  g16081(.dina(n34103), .dinb(n34101), .dout(n34104));
  jand g16082(.dina(n34104), .dinb(n33838), .dout(n34105));
  jxor g16083(.dina(n33830), .dinb(n410), .dout(n34106));
  jnot g16084(.din(n34106), .dout(n34107));
  jor  g16085(.dina(n34107), .dinb(n34105), .dout(n34108));
  jand g16086(.dina(n34108), .dinb(n33832), .dout(n34109));
  jxor g16087(.dina(n33824), .dinb(n426), .dout(n34110));
  jnot g16088(.din(n34110), .dout(n34111));
  jor  g16089(.dina(n34111), .dinb(n34109), .dout(n34112));
  jand g16090(.dina(n34112), .dinb(n33826), .dout(n34113));
  jxor g16091(.dina(n33818), .dinb(n427), .dout(n34114));
  jnot g16092(.din(n34114), .dout(n34115));
  jor  g16093(.dina(n34115), .dinb(n34113), .dout(n34116));
  jand g16094(.dina(n34116), .dinb(n33820), .dout(n34117));
  jxor g16095(.dina(n33812), .dinb(n424), .dout(n34118));
  jnot g16096(.din(n34118), .dout(n34119));
  jor  g16097(.dina(n34119), .dinb(n34117), .dout(n34120));
  jand g16098(.dina(n34120), .dinb(n33814), .dout(n34121));
  jxor g16099(.dina(n33806), .dinb(n300), .dout(n34122));
  jnot g16100(.din(n34122), .dout(n34123));
  jor  g16101(.dina(n34123), .dinb(n34121), .dout(n34124));
  jand g16102(.dina(n34124), .dinb(n33808), .dout(n34125));
  jxor g16103(.dina(n33800), .dinb(n297), .dout(n34126));
  jnot g16104(.din(n34126), .dout(n34127));
  jor  g16105(.dina(n34127), .dinb(n34125), .dout(n34128));
  jand g16106(.dina(n34128), .dinb(n33802), .dout(n34129));
  jxor g16107(.dina(n33794), .dinb(n298), .dout(n34130));
  jnot g16108(.din(n34130), .dout(n34131));
  jor  g16109(.dina(n34131), .dinb(n34129), .dout(n34132));
  jand g16110(.dina(n34132), .dinb(n33796), .dout(n34133));
  jxor g16111(.dina(n33788), .dinb(n301), .dout(n34134));
  jnot g16112(.din(n34134), .dout(n34135));
  jor  g16113(.dina(n34135), .dinb(n34133), .dout(n34136));
  jand g16114(.dina(n34136), .dinb(n33790), .dout(n34137));
  jxor g16115(.dina(n33782), .dinb(n293), .dout(n34138));
  jnot g16116(.din(n34138), .dout(n34139));
  jor  g16117(.dina(n34139), .dinb(n34137), .dout(n34140));
  jand g16118(.dina(n34140), .dinb(n33784), .dout(n34141));
  jxor g16119(.dina(n33776), .dinb(n294), .dout(n34142));
  jnot g16120(.din(n34142), .dout(n34143));
  jor  g16121(.dina(n34143), .dinb(n34141), .dout(n34144));
  jand g16122(.dina(n34144), .dinb(n33778), .dout(n34145));
  jxor g16123(.dina(n33770), .dinb(n290), .dout(n34146));
  jnot g16124(.din(n34146), .dout(n34147));
  jor  g16125(.dina(n34147), .dinb(n34145), .dout(n34148));
  jand g16126(.dina(n34148), .dinb(n33772), .dout(n34149));
  jxor g16127(.dina(n33764), .dinb(n291), .dout(n34150));
  jnot g16128(.din(n34150), .dout(n34151));
  jor  g16129(.dina(n34151), .dinb(n34149), .dout(n34152));
  jand g16130(.dina(n34152), .dinb(n33766), .dout(n34153));
  jxor g16131(.dina(n33758), .dinb(n284), .dout(n34154));
  jnot g16132(.din(n34154), .dout(n34155));
  jor  g16133(.dina(n34155), .dinb(n34153), .dout(n34156));
  jand g16134(.dina(n34156), .dinb(n33760), .dout(n34157));
  jxor g16135(.dina(n33752), .dinb(n285), .dout(n34158));
  jnot g16136(.din(n34158), .dout(n34159));
  jor  g16137(.dina(n34159), .dinb(n34157), .dout(n34160));
  jand g16138(.dina(n34160), .dinb(n33754), .dout(n34161));
  jxor g16139(.dina(n33746), .dinb(n281), .dout(n34162));
  jnot g16140(.din(n34162), .dout(n34163));
  jor  g16141(.dina(n34163), .dinb(n34161), .dout(n34164));
  jand g16142(.dina(n34164), .dinb(n33748), .dout(n34165));
  jxor g16143(.dina(n33740), .dinb(n282), .dout(n34166));
  jnot g16144(.din(n34166), .dout(n34167));
  jor  g16145(.dina(n34167), .dinb(n34165), .dout(n34168));
  jand g16146(.dina(n34168), .dinb(n33742), .dout(n34169));
  jxor g16147(.dina(n33734), .dinb(n397), .dout(n34170));
  jnot g16148(.din(n34170), .dout(n34171));
  jor  g16149(.dina(n34171), .dinb(n34169), .dout(n34172));
  jand g16150(.dina(n34172), .dinb(n33736), .dout(n34173));
  jxor g16151(.dina(n33728), .dinb(n513), .dout(n34174));
  jnot g16152(.din(n34174), .dout(n34175));
  jor  g16153(.dina(n34175), .dinb(n34173), .dout(n34176));
  jand g16154(.dina(n34176), .dinb(n33730), .dout(n34177));
  jxor g16155(.dina(n33722), .dinb(n514), .dout(n34178));
  jnot g16156(.din(n34178), .dout(n34179));
  jor  g16157(.dina(n34179), .dinb(n34177), .dout(n34180));
  jand g16158(.dina(n34180), .dinb(n33724), .dout(n34181));
  jxor g16159(.dina(n33716), .dinb(n510), .dout(n34182));
  jnot g16160(.din(n34182), .dout(n34183));
  jor  g16161(.dina(n34183), .dinb(n34181), .dout(n34184));
  jand g16162(.dina(n34184), .dinb(n33718), .dout(n34185));
  jxor g16163(.dina(n33710), .dinb(n396), .dout(n34186));
  jnot g16164(.din(n34186), .dout(n34187));
  jor  g16165(.dina(n34187), .dinb(n34185), .dout(n34188));
  jand g16166(.dina(n34188), .dinb(n33712), .dout(n34189));
  jxor g16167(.dina(n33704), .dinb(n383), .dout(n34190));
  jnot g16168(.din(n34190), .dout(n34191));
  jor  g16169(.dina(n34191), .dinb(n34189), .dout(n34192));
  jand g16170(.dina(n34192), .dinb(n33706), .dout(n34193));
  jxor g16171(.dina(n33698), .dinb(b50 ), .dout(n34194));
  jand g16172(.dina(n34194), .dinb(n12216), .dout(n34195));
  jnot g16173(.din(n34195), .dout(n34196));
  jor  g16174(.dina(n34196), .dinb(n34193), .dout(n34197));
  jand g16175(.dina(n34197), .dinb(n33698), .dout(n34198));
  jxor g16176(.dina(n33998), .dinb(b1 ), .dout(n34199));
  jand g16177(.dina(n34199), .dinb(n12063), .dout(n34200));
  jor  g16178(.dina(n34200), .dinb(n33994), .dout(n34201));
  jand g16179(.dina(n34002), .dinb(n34201), .dout(n34202));
  jor  g16180(.dina(n34202), .dinb(n33987), .dout(n34203));
  jand g16181(.dina(n34006), .dinb(n34203), .dout(n34204));
  jor  g16182(.dina(n34204), .dinb(n33981), .dout(n34205));
  jand g16183(.dina(n34010), .dinb(n34205), .dout(n34206));
  jor  g16184(.dina(n34206), .dinb(n33975), .dout(n34207));
  jand g16185(.dina(n34014), .dinb(n34207), .dout(n34208));
  jor  g16186(.dina(n34208), .dinb(n33969), .dout(n34209));
  jand g16187(.dina(n34018), .dinb(n34209), .dout(n34210));
  jor  g16188(.dina(n34210), .dinb(n33963), .dout(n34211));
  jand g16189(.dina(n34022), .dinb(n34211), .dout(n34212));
  jor  g16190(.dina(n34212), .dinb(n33957), .dout(n34213));
  jand g16191(.dina(n34026), .dinb(n34213), .dout(n34214));
  jor  g16192(.dina(n34214), .dinb(n33951), .dout(n34215));
  jand g16193(.dina(n34030), .dinb(n34215), .dout(n34216));
  jor  g16194(.dina(n34216), .dinb(n33945), .dout(n34217));
  jand g16195(.dina(n34034), .dinb(n34217), .dout(n34218));
  jor  g16196(.dina(n34218), .dinb(n33939), .dout(n34219));
  jand g16197(.dina(n34038), .dinb(n34219), .dout(n34220));
  jor  g16198(.dina(n34220), .dinb(n33933), .dout(n34221));
  jand g16199(.dina(n34042), .dinb(n34221), .dout(n34222));
  jor  g16200(.dina(n34222), .dinb(n33927), .dout(n34223));
  jand g16201(.dina(n34046), .dinb(n34223), .dout(n34224));
  jor  g16202(.dina(n34224), .dinb(n33921), .dout(n34225));
  jand g16203(.dina(n34050), .dinb(n34225), .dout(n34226));
  jor  g16204(.dina(n34226), .dinb(n33915), .dout(n34227));
  jand g16205(.dina(n34054), .dinb(n34227), .dout(n34228));
  jor  g16206(.dina(n34228), .dinb(n33909), .dout(n34229));
  jand g16207(.dina(n34058), .dinb(n34229), .dout(n34230));
  jor  g16208(.dina(n34230), .dinb(n33903), .dout(n34231));
  jand g16209(.dina(n34062), .dinb(n34231), .dout(n34232));
  jor  g16210(.dina(n34232), .dinb(n33897), .dout(n34233));
  jand g16211(.dina(n34066), .dinb(n34233), .dout(n34234));
  jor  g16212(.dina(n34234), .dinb(n33891), .dout(n34235));
  jand g16213(.dina(n34070), .dinb(n34235), .dout(n34236));
  jor  g16214(.dina(n34236), .dinb(n33885), .dout(n34237));
  jand g16215(.dina(n34074), .dinb(n34237), .dout(n34238));
  jor  g16216(.dina(n34238), .dinb(n33879), .dout(n34239));
  jand g16217(.dina(n34078), .dinb(n34239), .dout(n34240));
  jor  g16218(.dina(n34240), .dinb(n33873), .dout(n34241));
  jand g16219(.dina(n34082), .dinb(n34241), .dout(n34242));
  jor  g16220(.dina(n34242), .dinb(n33867), .dout(n34243));
  jand g16221(.dina(n34086), .dinb(n34243), .dout(n34244));
  jor  g16222(.dina(n34244), .dinb(n33861), .dout(n34245));
  jand g16223(.dina(n34090), .dinb(n34245), .dout(n34246));
  jor  g16224(.dina(n34246), .dinb(n33855), .dout(n34247));
  jand g16225(.dina(n34094), .dinb(n34247), .dout(n34248));
  jor  g16226(.dina(n34248), .dinb(n33849), .dout(n34249));
  jand g16227(.dina(n34098), .dinb(n34249), .dout(n34250));
  jor  g16228(.dina(n34250), .dinb(n33843), .dout(n34251));
  jand g16229(.dina(n34102), .dinb(n34251), .dout(n34252));
  jor  g16230(.dina(n34252), .dinb(n33837), .dout(n34253));
  jand g16231(.dina(n34106), .dinb(n34253), .dout(n34254));
  jor  g16232(.dina(n34254), .dinb(n33831), .dout(n34255));
  jand g16233(.dina(n34110), .dinb(n34255), .dout(n34256));
  jor  g16234(.dina(n34256), .dinb(n33825), .dout(n34257));
  jand g16235(.dina(n34114), .dinb(n34257), .dout(n34258));
  jor  g16236(.dina(n34258), .dinb(n33819), .dout(n34259));
  jand g16237(.dina(n34118), .dinb(n34259), .dout(n34260));
  jor  g16238(.dina(n34260), .dinb(n33813), .dout(n34261));
  jand g16239(.dina(n34122), .dinb(n34261), .dout(n34262));
  jor  g16240(.dina(n34262), .dinb(n33807), .dout(n34263));
  jand g16241(.dina(n34126), .dinb(n34263), .dout(n34264));
  jor  g16242(.dina(n34264), .dinb(n33801), .dout(n34265));
  jand g16243(.dina(n34130), .dinb(n34265), .dout(n34266));
  jor  g16244(.dina(n34266), .dinb(n33795), .dout(n34267));
  jand g16245(.dina(n34134), .dinb(n34267), .dout(n34268));
  jor  g16246(.dina(n34268), .dinb(n33789), .dout(n34269));
  jand g16247(.dina(n34138), .dinb(n34269), .dout(n34270));
  jor  g16248(.dina(n34270), .dinb(n33783), .dout(n34271));
  jand g16249(.dina(n34142), .dinb(n34271), .dout(n34272));
  jor  g16250(.dina(n34272), .dinb(n33777), .dout(n34273));
  jand g16251(.dina(n34146), .dinb(n34273), .dout(n34274));
  jor  g16252(.dina(n34274), .dinb(n33771), .dout(n34275));
  jand g16253(.dina(n34150), .dinb(n34275), .dout(n34276));
  jor  g16254(.dina(n34276), .dinb(n33765), .dout(n34277));
  jand g16255(.dina(n34154), .dinb(n34277), .dout(n34278));
  jor  g16256(.dina(n34278), .dinb(n33759), .dout(n34279));
  jand g16257(.dina(n34158), .dinb(n34279), .dout(n34280));
  jor  g16258(.dina(n34280), .dinb(n33753), .dout(n34281));
  jand g16259(.dina(n34162), .dinb(n34281), .dout(n34282));
  jor  g16260(.dina(n34282), .dinb(n33747), .dout(n34283));
  jand g16261(.dina(n34166), .dinb(n34283), .dout(n34284));
  jor  g16262(.dina(n34284), .dinb(n33741), .dout(n34285));
  jand g16263(.dina(n34170), .dinb(n34285), .dout(n34286));
  jor  g16264(.dina(n34286), .dinb(n33735), .dout(n34287));
  jand g16265(.dina(n34174), .dinb(n34287), .dout(n34288));
  jor  g16266(.dina(n34288), .dinb(n33729), .dout(n34289));
  jand g16267(.dina(n34178), .dinb(n34289), .dout(n34290));
  jor  g16268(.dina(n34290), .dinb(n33723), .dout(n34291));
  jand g16269(.dina(n34182), .dinb(n34291), .dout(n34292));
  jor  g16270(.dina(n34292), .dinb(n33717), .dout(n34293));
  jand g16271(.dina(n34186), .dinb(n34293), .dout(n34294));
  jor  g16272(.dina(n34294), .dinb(n33711), .dout(n34295));
  jand g16273(.dina(n34190), .dinb(n34295), .dout(n34296));
  jor  g16274(.dina(n34296), .dinb(n33705), .dout(n34297));
  jand g16275(.dina(n34195), .dinb(n34297), .dout(n34298));
  jor  g16276(.dina(n33698), .dinb(n11794), .dout(n34299));
  jnot g16277(.din(n34299), .dout(n34300));
  jor  g16278(.dina(n34300), .dinb(n34298), .dout(n34301));
  jxor g16279(.dina(n34194), .dinb(n34193), .dout(n34302));
  jand g16280(.dina(n34302), .dinb(n34301), .dout(n34303));
  jor  g16281(.dina(n34303), .dinb(n34198), .dout(n34304));
  jnot g16282(.din(n34304), .dout(n34305));
  jand g16283(.dina(n34304), .dinb(b51 ), .dout(n34306));
  jnot g16284(.din(n34306), .dout(n34307));
  jand g16285(.dina(n34305), .dinb(n12214), .dout(n34308));
  jand g16286(.dina(n34299), .dinb(n34197), .dout(n34309));
  jand g16287(.dina(n34309), .dinb(n33704), .dout(n34310));
  jxor g16288(.dina(n34190), .dinb(n34295), .dout(n34311));
  jand g16289(.dina(n34311), .dinb(n34301), .dout(n34312));
  jor  g16290(.dina(n34312), .dinb(n34310), .dout(n34313));
  jand g16291(.dina(n34313), .dinb(n12211), .dout(n34314));
  jand g16292(.dina(n34309), .dinb(n33710), .dout(n34315));
  jxor g16293(.dina(n34186), .dinb(n34293), .dout(n34316));
  jand g16294(.dina(n34316), .dinb(n34301), .dout(n34317));
  jor  g16295(.dina(n34317), .dinb(n34315), .dout(n34318));
  jand g16296(.dina(n34318), .dinb(n383), .dout(n34319));
  jand g16297(.dina(n34309), .dinb(n33716), .dout(n34320));
  jxor g16298(.dina(n34182), .dinb(n34291), .dout(n34321));
  jand g16299(.dina(n34321), .dinb(n34301), .dout(n34322));
  jor  g16300(.dina(n34322), .dinb(n34320), .dout(n34323));
  jand g16301(.dina(n34323), .dinb(n396), .dout(n34324));
  jand g16302(.dina(n34309), .dinb(n33722), .dout(n34325));
  jxor g16303(.dina(n34178), .dinb(n34289), .dout(n34326));
  jand g16304(.dina(n34326), .dinb(n34301), .dout(n34327));
  jor  g16305(.dina(n34327), .dinb(n34325), .dout(n34328));
  jand g16306(.dina(n34328), .dinb(n510), .dout(n34329));
  jand g16307(.dina(n34309), .dinb(n33728), .dout(n34330));
  jxor g16308(.dina(n34174), .dinb(n34287), .dout(n34331));
  jand g16309(.dina(n34331), .dinb(n34301), .dout(n34332));
  jor  g16310(.dina(n34332), .dinb(n34330), .dout(n34333));
  jand g16311(.dina(n34333), .dinb(n514), .dout(n34334));
  jand g16312(.dina(n34309), .dinb(n33734), .dout(n34335));
  jxor g16313(.dina(n34170), .dinb(n34285), .dout(n34336));
  jand g16314(.dina(n34336), .dinb(n34301), .dout(n34337));
  jor  g16315(.dina(n34337), .dinb(n34335), .dout(n34338));
  jand g16316(.dina(n34338), .dinb(n513), .dout(n34339));
  jand g16317(.dina(n34309), .dinb(n33740), .dout(n34340));
  jxor g16318(.dina(n34166), .dinb(n34283), .dout(n34341));
  jand g16319(.dina(n34341), .dinb(n34301), .dout(n34342));
  jor  g16320(.dina(n34342), .dinb(n34340), .dout(n34343));
  jand g16321(.dina(n34343), .dinb(n397), .dout(n34344));
  jand g16322(.dina(n34309), .dinb(n33746), .dout(n34345));
  jxor g16323(.dina(n34162), .dinb(n34281), .dout(n34346));
  jand g16324(.dina(n34346), .dinb(n34301), .dout(n34347));
  jor  g16325(.dina(n34347), .dinb(n34345), .dout(n34348));
  jand g16326(.dina(n34348), .dinb(n282), .dout(n34349));
  jand g16327(.dina(n34309), .dinb(n33752), .dout(n34350));
  jxor g16328(.dina(n34158), .dinb(n34279), .dout(n34351));
  jand g16329(.dina(n34351), .dinb(n34301), .dout(n34352));
  jor  g16330(.dina(n34352), .dinb(n34350), .dout(n34353));
  jand g16331(.dina(n34353), .dinb(n281), .dout(n34354));
  jand g16332(.dina(n34309), .dinb(n33758), .dout(n34355));
  jxor g16333(.dina(n34154), .dinb(n34277), .dout(n34356));
  jand g16334(.dina(n34356), .dinb(n34301), .dout(n34357));
  jor  g16335(.dina(n34357), .dinb(n34355), .dout(n34358));
  jand g16336(.dina(n34358), .dinb(n285), .dout(n34359));
  jand g16337(.dina(n34309), .dinb(n33764), .dout(n34360));
  jxor g16338(.dina(n34150), .dinb(n34275), .dout(n34361));
  jand g16339(.dina(n34361), .dinb(n34301), .dout(n34362));
  jor  g16340(.dina(n34362), .dinb(n34360), .dout(n34363));
  jand g16341(.dina(n34363), .dinb(n284), .dout(n34364));
  jand g16342(.dina(n34309), .dinb(n33770), .dout(n34365));
  jxor g16343(.dina(n34146), .dinb(n34273), .dout(n34366));
  jand g16344(.dina(n34366), .dinb(n34301), .dout(n34367));
  jor  g16345(.dina(n34367), .dinb(n34365), .dout(n34368));
  jand g16346(.dina(n34368), .dinb(n291), .dout(n34369));
  jand g16347(.dina(n34309), .dinb(n33776), .dout(n34370));
  jxor g16348(.dina(n34142), .dinb(n34271), .dout(n34371));
  jand g16349(.dina(n34371), .dinb(n34301), .dout(n34372));
  jor  g16350(.dina(n34372), .dinb(n34370), .dout(n34373));
  jand g16351(.dina(n34373), .dinb(n290), .dout(n34374));
  jand g16352(.dina(n34309), .dinb(n33782), .dout(n34375));
  jxor g16353(.dina(n34138), .dinb(n34269), .dout(n34376));
  jand g16354(.dina(n34376), .dinb(n34301), .dout(n34377));
  jor  g16355(.dina(n34377), .dinb(n34375), .dout(n34378));
  jand g16356(.dina(n34378), .dinb(n294), .dout(n34379));
  jand g16357(.dina(n34309), .dinb(n33788), .dout(n34380));
  jxor g16358(.dina(n34134), .dinb(n34267), .dout(n34381));
  jand g16359(.dina(n34381), .dinb(n34301), .dout(n34382));
  jor  g16360(.dina(n34382), .dinb(n34380), .dout(n34383));
  jand g16361(.dina(n34383), .dinb(n293), .dout(n34384));
  jand g16362(.dina(n34309), .dinb(n33794), .dout(n34385));
  jxor g16363(.dina(n34130), .dinb(n34265), .dout(n34386));
  jand g16364(.dina(n34386), .dinb(n34301), .dout(n34387));
  jor  g16365(.dina(n34387), .dinb(n34385), .dout(n34388));
  jand g16366(.dina(n34388), .dinb(n301), .dout(n34389));
  jand g16367(.dina(n34309), .dinb(n33800), .dout(n34390));
  jxor g16368(.dina(n34126), .dinb(n34263), .dout(n34391));
  jand g16369(.dina(n34391), .dinb(n34301), .dout(n34392));
  jor  g16370(.dina(n34392), .dinb(n34390), .dout(n34393));
  jand g16371(.dina(n34393), .dinb(n298), .dout(n34394));
  jand g16372(.dina(n34309), .dinb(n33806), .dout(n34395));
  jxor g16373(.dina(n34122), .dinb(n34261), .dout(n34396));
  jand g16374(.dina(n34396), .dinb(n34301), .dout(n34397));
  jor  g16375(.dina(n34397), .dinb(n34395), .dout(n34398));
  jand g16376(.dina(n34398), .dinb(n297), .dout(n34399));
  jand g16377(.dina(n34309), .dinb(n33812), .dout(n34400));
  jxor g16378(.dina(n34118), .dinb(n34259), .dout(n34401));
  jand g16379(.dina(n34401), .dinb(n34301), .dout(n34402));
  jor  g16380(.dina(n34402), .dinb(n34400), .dout(n34403));
  jand g16381(.dina(n34403), .dinb(n300), .dout(n34404));
  jand g16382(.dina(n34309), .dinb(n33818), .dout(n34405));
  jxor g16383(.dina(n34114), .dinb(n34257), .dout(n34406));
  jand g16384(.dina(n34406), .dinb(n34301), .dout(n34407));
  jor  g16385(.dina(n34407), .dinb(n34405), .dout(n34408));
  jand g16386(.dina(n34408), .dinb(n424), .dout(n34409));
  jand g16387(.dina(n34309), .dinb(n33824), .dout(n34410));
  jxor g16388(.dina(n34110), .dinb(n34255), .dout(n34411));
  jand g16389(.dina(n34411), .dinb(n34301), .dout(n34412));
  jor  g16390(.dina(n34412), .dinb(n34410), .dout(n34413));
  jand g16391(.dina(n34413), .dinb(n427), .dout(n34414));
  jand g16392(.dina(n34309), .dinb(n33830), .dout(n34415));
  jxor g16393(.dina(n34106), .dinb(n34253), .dout(n34416));
  jand g16394(.dina(n34416), .dinb(n34301), .dout(n34417));
  jor  g16395(.dina(n34417), .dinb(n34415), .dout(n34418));
  jand g16396(.dina(n34418), .dinb(n426), .dout(n34419));
  jand g16397(.dina(n34309), .dinb(n33836), .dout(n34420));
  jxor g16398(.dina(n34102), .dinb(n34251), .dout(n34421));
  jand g16399(.dina(n34421), .dinb(n34301), .dout(n34422));
  jor  g16400(.dina(n34422), .dinb(n34420), .dout(n34423));
  jand g16401(.dina(n34423), .dinb(n410), .dout(n34424));
  jand g16402(.dina(n34309), .dinb(n33842), .dout(n34425));
  jxor g16403(.dina(n34098), .dinb(n34249), .dout(n34426));
  jand g16404(.dina(n34426), .dinb(n34301), .dout(n34427));
  jor  g16405(.dina(n34427), .dinb(n34425), .dout(n34428));
  jand g16406(.dina(n34428), .dinb(n409), .dout(n34429));
  jand g16407(.dina(n34309), .dinb(n33848), .dout(n34430));
  jxor g16408(.dina(n34094), .dinb(n34247), .dout(n34431));
  jand g16409(.dina(n34431), .dinb(n34301), .dout(n34432));
  jor  g16410(.dina(n34432), .dinb(n34430), .dout(n34433));
  jand g16411(.dina(n34433), .dinb(n413), .dout(n34434));
  jand g16412(.dina(n34309), .dinb(n33854), .dout(n34435));
  jxor g16413(.dina(n34090), .dinb(n34245), .dout(n34436));
  jand g16414(.dina(n34436), .dinb(n34301), .dout(n34437));
  jor  g16415(.dina(n34437), .dinb(n34435), .dout(n34438));
  jand g16416(.dina(n34438), .dinb(n412), .dout(n34439));
  jand g16417(.dina(n34309), .dinb(n33860), .dout(n34440));
  jxor g16418(.dina(n34086), .dinb(n34243), .dout(n34441));
  jand g16419(.dina(n34441), .dinb(n34301), .dout(n34442));
  jor  g16420(.dina(n34442), .dinb(n34440), .dout(n34443));
  jand g16421(.dina(n34443), .dinb(n406), .dout(n34444));
  jand g16422(.dina(n34309), .dinb(n33866), .dout(n34445));
  jxor g16423(.dina(n34082), .dinb(n34241), .dout(n34446));
  jand g16424(.dina(n34446), .dinb(n34301), .dout(n34447));
  jor  g16425(.dina(n34447), .dinb(n34445), .dout(n34448));
  jand g16426(.dina(n34448), .dinb(n405), .dout(n34449));
  jand g16427(.dina(n34309), .dinb(n33872), .dout(n34450));
  jxor g16428(.dina(n34078), .dinb(n34239), .dout(n34451));
  jand g16429(.dina(n34451), .dinb(n34301), .dout(n34452));
  jor  g16430(.dina(n34452), .dinb(n34450), .dout(n34453));
  jand g16431(.dina(n34453), .dinb(n2714), .dout(n34454));
  jand g16432(.dina(n34309), .dinb(n33878), .dout(n34455));
  jxor g16433(.dina(n34074), .dinb(n34237), .dout(n34456));
  jand g16434(.dina(n34456), .dinb(n34301), .dout(n34457));
  jor  g16435(.dina(n34457), .dinb(n34455), .dout(n34458));
  jand g16436(.dina(n34458), .dinb(n2547), .dout(n34459));
  jand g16437(.dina(n34309), .dinb(n33884), .dout(n34460));
  jxor g16438(.dina(n34070), .dinb(n34235), .dout(n34461));
  jand g16439(.dina(n34461), .dinb(n34301), .dout(n34462));
  jor  g16440(.dina(n34462), .dinb(n34460), .dout(n34463));
  jand g16441(.dina(n34463), .dinb(n417), .dout(n34464));
  jand g16442(.dina(n34309), .dinb(n33890), .dout(n34465));
  jxor g16443(.dina(n34066), .dinb(n34233), .dout(n34466));
  jand g16444(.dina(n34466), .dinb(n34301), .dout(n34467));
  jor  g16445(.dina(n34467), .dinb(n34465), .dout(n34468));
  jand g16446(.dina(n34468), .dinb(n416), .dout(n34469));
  jand g16447(.dina(n34309), .dinb(n33896), .dout(n34470));
  jxor g16448(.dina(n34062), .dinb(n34231), .dout(n34471));
  jand g16449(.dina(n34471), .dinb(n34301), .dout(n34472));
  jor  g16450(.dina(n34472), .dinb(n34470), .dout(n34473));
  jand g16451(.dina(n34473), .dinb(n422), .dout(n34474));
  jand g16452(.dina(n34309), .dinb(n33902), .dout(n34475));
  jxor g16453(.dina(n34058), .dinb(n34229), .dout(n34476));
  jand g16454(.dina(n34476), .dinb(n34301), .dout(n34477));
  jor  g16455(.dina(n34477), .dinb(n34475), .dout(n34478));
  jand g16456(.dina(n34478), .dinb(n421), .dout(n34479));
  jand g16457(.dina(n34309), .dinb(n33908), .dout(n34480));
  jxor g16458(.dina(n34054), .dinb(n34227), .dout(n34481));
  jand g16459(.dina(n34481), .dinb(n34301), .dout(n34482));
  jor  g16460(.dina(n34482), .dinb(n34480), .dout(n34483));
  jand g16461(.dina(n34483), .dinb(n433), .dout(n34484));
  jand g16462(.dina(n34309), .dinb(n33914), .dout(n34485));
  jxor g16463(.dina(n34050), .dinb(n34225), .dout(n34486));
  jand g16464(.dina(n34486), .dinb(n34301), .dout(n34487));
  jor  g16465(.dina(n34487), .dinb(n34485), .dout(n34488));
  jand g16466(.dina(n34488), .dinb(n432), .dout(n34489));
  jand g16467(.dina(n34309), .dinb(n33920), .dout(n34490));
  jxor g16468(.dina(n34046), .dinb(n34223), .dout(n34491));
  jand g16469(.dina(n34491), .dinb(n34301), .dout(n34492));
  jor  g16470(.dina(n34492), .dinb(n34490), .dout(n34493));
  jand g16471(.dina(n34493), .dinb(n436), .dout(n34494));
  jand g16472(.dina(n34309), .dinb(n33926), .dout(n34495));
  jxor g16473(.dina(n34042), .dinb(n34221), .dout(n34496));
  jand g16474(.dina(n34496), .dinb(n34301), .dout(n34497));
  jor  g16475(.dina(n34497), .dinb(n34495), .dout(n34498));
  jand g16476(.dina(n34498), .dinb(n435), .dout(n34499));
  jand g16477(.dina(n34309), .dinb(n33932), .dout(n34500));
  jxor g16478(.dina(n34038), .dinb(n34219), .dout(n34501));
  jand g16479(.dina(n34501), .dinb(n34301), .dout(n34502));
  jor  g16480(.dina(n34502), .dinb(n34500), .dout(n34503));
  jand g16481(.dina(n34503), .dinb(n440), .dout(n34504));
  jand g16482(.dina(n34309), .dinb(n33938), .dout(n34505));
  jxor g16483(.dina(n34034), .dinb(n34217), .dout(n34506));
  jand g16484(.dina(n34506), .dinb(n34301), .dout(n34507));
  jor  g16485(.dina(n34507), .dinb(n34505), .dout(n34508));
  jand g16486(.dina(n34508), .dinb(n439), .dout(n34509));
  jand g16487(.dina(n34309), .dinb(n33944), .dout(n34510));
  jxor g16488(.dina(n34030), .dinb(n34215), .dout(n34511));
  jand g16489(.dina(n34511), .dinb(n34301), .dout(n34512));
  jor  g16490(.dina(n34512), .dinb(n34510), .dout(n34513));
  jand g16491(.dina(n34513), .dinb(n325), .dout(n34514));
  jand g16492(.dina(n34309), .dinb(n33950), .dout(n34515));
  jxor g16493(.dina(n34026), .dinb(n34213), .dout(n34516));
  jand g16494(.dina(n34516), .dinb(n34301), .dout(n34517));
  jor  g16495(.dina(n34517), .dinb(n34515), .dout(n34518));
  jand g16496(.dina(n34518), .dinb(n324), .dout(n34519));
  jand g16497(.dina(n34309), .dinb(n33956), .dout(n34520));
  jxor g16498(.dina(n34022), .dinb(n34211), .dout(n34521));
  jand g16499(.dina(n34521), .dinb(n34301), .dout(n34522));
  jor  g16500(.dina(n34522), .dinb(n34520), .dout(n34523));
  jand g16501(.dina(n34523), .dinb(n323), .dout(n34524));
  jand g16502(.dina(n34309), .dinb(n33962), .dout(n34525));
  jxor g16503(.dina(n34018), .dinb(n34209), .dout(n34526));
  jand g16504(.dina(n34526), .dinb(n34301), .dout(n34527));
  jor  g16505(.dina(n34527), .dinb(n34525), .dout(n34528));
  jand g16506(.dina(n34528), .dinb(n335), .dout(n34529));
  jand g16507(.dina(n34309), .dinb(n33968), .dout(n34530));
  jxor g16508(.dina(n34014), .dinb(n34207), .dout(n34531));
  jand g16509(.dina(n34531), .dinb(n34301), .dout(n34532));
  jor  g16510(.dina(n34532), .dinb(n34530), .dout(n34533));
  jand g16511(.dina(n34533), .dinb(n334), .dout(n34534));
  jand g16512(.dina(n34309), .dinb(n33974), .dout(n34535));
  jxor g16513(.dina(n34010), .dinb(n34205), .dout(n34536));
  jand g16514(.dina(n34536), .dinb(n34301), .dout(n34537));
  jor  g16515(.dina(n34537), .dinb(n34535), .dout(n34538));
  jand g16516(.dina(n34538), .dinb(n338), .dout(n34539));
  jand g16517(.dina(n34309), .dinb(n33980), .dout(n34540));
  jxor g16518(.dina(n34006), .dinb(n34203), .dout(n34541));
  jand g16519(.dina(n34541), .dinb(n34301), .dout(n34542));
  jor  g16520(.dina(n34542), .dinb(n34540), .dout(n34543));
  jand g16521(.dina(n34543), .dinb(n337), .dout(n34544));
  jand g16522(.dina(n34309), .dinb(n33986), .dout(n34545));
  jxor g16523(.dina(n34002), .dinb(n34201), .dout(n34546));
  jand g16524(.dina(n34546), .dinb(n34301), .dout(n34547));
  jor  g16525(.dina(n34547), .dinb(n34545), .dout(n34548));
  jand g16526(.dina(n34548), .dinb(n344), .dout(n34549));
  jand g16527(.dina(n34309), .dinb(n33993), .dout(n34550));
  jxor g16528(.dina(n34199), .dinb(n12063), .dout(n34551));
  jand g16529(.dina(n34551), .dinb(n34301), .dout(n34552));
  jor  g16530(.dina(n34552), .dinb(n34550), .dout(n34553));
  jand g16531(.dina(n34553), .dinb(n348), .dout(n34554));
  jor  g16532(.dina(n34309), .dinb(n18364), .dout(n34555));
  jand g16533(.dina(n34555), .dinb(a13 ), .dout(n34556));
  jor  g16534(.dina(n34309), .dinb(n12063), .dout(n34557));
  jnot g16535(.din(n34557), .dout(n34558));
  jor  g16536(.dina(n34558), .dinb(n34556), .dout(n34559));
  jand g16537(.dina(n34559), .dinb(n258), .dout(n34560));
  jand g16538(.dina(n34301), .dinb(b0 ), .dout(n34561));
  jor  g16539(.dina(n34561), .dinb(n12061), .dout(n34562));
  jand g16540(.dina(n34557), .dinb(n34562), .dout(n34563));
  jxor g16541(.dina(n34563), .dinb(b1 ), .dout(n34564));
  jand g16542(.dina(n34564), .dinb(n12487), .dout(n34565));
  jor  g16543(.dina(n34565), .dinb(n34560), .dout(n34566));
  jxor g16544(.dina(n34553), .dinb(n348), .dout(n34567));
  jand g16545(.dina(n34567), .dinb(n34566), .dout(n34568));
  jor  g16546(.dina(n34568), .dinb(n34554), .dout(n34569));
  jxor g16547(.dina(n34548), .dinb(n344), .dout(n34570));
  jand g16548(.dina(n34570), .dinb(n34569), .dout(n34571));
  jor  g16549(.dina(n34571), .dinb(n34549), .dout(n34572));
  jxor g16550(.dina(n34543), .dinb(n337), .dout(n34573));
  jand g16551(.dina(n34573), .dinb(n34572), .dout(n34574));
  jor  g16552(.dina(n34574), .dinb(n34544), .dout(n34575));
  jxor g16553(.dina(n34538), .dinb(n338), .dout(n34576));
  jand g16554(.dina(n34576), .dinb(n34575), .dout(n34577));
  jor  g16555(.dina(n34577), .dinb(n34539), .dout(n34578));
  jxor g16556(.dina(n34533), .dinb(n334), .dout(n34579));
  jand g16557(.dina(n34579), .dinb(n34578), .dout(n34580));
  jor  g16558(.dina(n34580), .dinb(n34534), .dout(n34581));
  jxor g16559(.dina(n34528), .dinb(n335), .dout(n34582));
  jand g16560(.dina(n34582), .dinb(n34581), .dout(n34583));
  jor  g16561(.dina(n34583), .dinb(n34529), .dout(n34584));
  jxor g16562(.dina(n34523), .dinb(n323), .dout(n34585));
  jand g16563(.dina(n34585), .dinb(n34584), .dout(n34586));
  jor  g16564(.dina(n34586), .dinb(n34524), .dout(n34587));
  jxor g16565(.dina(n34518), .dinb(n324), .dout(n34588));
  jand g16566(.dina(n34588), .dinb(n34587), .dout(n34589));
  jor  g16567(.dina(n34589), .dinb(n34519), .dout(n34590));
  jxor g16568(.dina(n34513), .dinb(n325), .dout(n34591));
  jand g16569(.dina(n34591), .dinb(n34590), .dout(n34592));
  jor  g16570(.dina(n34592), .dinb(n34514), .dout(n34593));
  jxor g16571(.dina(n34508), .dinb(n439), .dout(n34594));
  jand g16572(.dina(n34594), .dinb(n34593), .dout(n34595));
  jor  g16573(.dina(n34595), .dinb(n34509), .dout(n34596));
  jxor g16574(.dina(n34503), .dinb(n440), .dout(n34597));
  jand g16575(.dina(n34597), .dinb(n34596), .dout(n34598));
  jor  g16576(.dina(n34598), .dinb(n34504), .dout(n34599));
  jxor g16577(.dina(n34498), .dinb(n435), .dout(n34600));
  jand g16578(.dina(n34600), .dinb(n34599), .dout(n34601));
  jor  g16579(.dina(n34601), .dinb(n34499), .dout(n34602));
  jxor g16580(.dina(n34493), .dinb(n436), .dout(n34603));
  jand g16581(.dina(n34603), .dinb(n34602), .dout(n34604));
  jor  g16582(.dina(n34604), .dinb(n34494), .dout(n34605));
  jxor g16583(.dina(n34488), .dinb(n432), .dout(n34606));
  jand g16584(.dina(n34606), .dinb(n34605), .dout(n34607));
  jor  g16585(.dina(n34607), .dinb(n34489), .dout(n34608));
  jxor g16586(.dina(n34483), .dinb(n433), .dout(n34609));
  jand g16587(.dina(n34609), .dinb(n34608), .dout(n34610));
  jor  g16588(.dina(n34610), .dinb(n34484), .dout(n34611));
  jxor g16589(.dina(n34478), .dinb(n421), .dout(n34612));
  jand g16590(.dina(n34612), .dinb(n34611), .dout(n34613));
  jor  g16591(.dina(n34613), .dinb(n34479), .dout(n34614));
  jxor g16592(.dina(n34473), .dinb(n422), .dout(n34615));
  jand g16593(.dina(n34615), .dinb(n34614), .dout(n34616));
  jor  g16594(.dina(n34616), .dinb(n34474), .dout(n34617));
  jxor g16595(.dina(n34468), .dinb(n416), .dout(n34618));
  jand g16596(.dina(n34618), .dinb(n34617), .dout(n34619));
  jor  g16597(.dina(n34619), .dinb(n34469), .dout(n34620));
  jxor g16598(.dina(n34463), .dinb(n417), .dout(n34621));
  jand g16599(.dina(n34621), .dinb(n34620), .dout(n34622));
  jor  g16600(.dina(n34622), .dinb(n34464), .dout(n34623));
  jxor g16601(.dina(n34458), .dinb(n2547), .dout(n34624));
  jand g16602(.dina(n34624), .dinb(n34623), .dout(n34625));
  jor  g16603(.dina(n34625), .dinb(n34459), .dout(n34626));
  jxor g16604(.dina(n34453), .dinb(n2714), .dout(n34627));
  jand g16605(.dina(n34627), .dinb(n34626), .dout(n34628));
  jor  g16606(.dina(n34628), .dinb(n34454), .dout(n34629));
  jxor g16607(.dina(n34448), .dinb(n405), .dout(n34630));
  jand g16608(.dina(n34630), .dinb(n34629), .dout(n34631));
  jor  g16609(.dina(n34631), .dinb(n34449), .dout(n34632));
  jxor g16610(.dina(n34443), .dinb(n406), .dout(n34633));
  jand g16611(.dina(n34633), .dinb(n34632), .dout(n34634));
  jor  g16612(.dina(n34634), .dinb(n34444), .dout(n34635));
  jxor g16613(.dina(n34438), .dinb(n412), .dout(n34636));
  jand g16614(.dina(n34636), .dinb(n34635), .dout(n34637));
  jor  g16615(.dina(n34637), .dinb(n34439), .dout(n34638));
  jxor g16616(.dina(n34433), .dinb(n413), .dout(n34639));
  jand g16617(.dina(n34639), .dinb(n34638), .dout(n34640));
  jor  g16618(.dina(n34640), .dinb(n34434), .dout(n34641));
  jxor g16619(.dina(n34428), .dinb(n409), .dout(n34642));
  jand g16620(.dina(n34642), .dinb(n34641), .dout(n34643));
  jor  g16621(.dina(n34643), .dinb(n34429), .dout(n34644));
  jxor g16622(.dina(n34423), .dinb(n410), .dout(n34645));
  jand g16623(.dina(n34645), .dinb(n34644), .dout(n34646));
  jor  g16624(.dina(n34646), .dinb(n34424), .dout(n34647));
  jxor g16625(.dina(n34418), .dinb(n426), .dout(n34648));
  jand g16626(.dina(n34648), .dinb(n34647), .dout(n34649));
  jor  g16627(.dina(n34649), .dinb(n34419), .dout(n34650));
  jxor g16628(.dina(n34413), .dinb(n427), .dout(n34651));
  jand g16629(.dina(n34651), .dinb(n34650), .dout(n34652));
  jor  g16630(.dina(n34652), .dinb(n34414), .dout(n34653));
  jxor g16631(.dina(n34408), .dinb(n424), .dout(n34654));
  jand g16632(.dina(n34654), .dinb(n34653), .dout(n34655));
  jor  g16633(.dina(n34655), .dinb(n34409), .dout(n34656));
  jxor g16634(.dina(n34403), .dinb(n300), .dout(n34657));
  jand g16635(.dina(n34657), .dinb(n34656), .dout(n34658));
  jor  g16636(.dina(n34658), .dinb(n34404), .dout(n34659));
  jxor g16637(.dina(n34398), .dinb(n297), .dout(n34660));
  jand g16638(.dina(n34660), .dinb(n34659), .dout(n34661));
  jor  g16639(.dina(n34661), .dinb(n34399), .dout(n34662));
  jxor g16640(.dina(n34393), .dinb(n298), .dout(n34663));
  jand g16641(.dina(n34663), .dinb(n34662), .dout(n34664));
  jor  g16642(.dina(n34664), .dinb(n34394), .dout(n34665));
  jxor g16643(.dina(n34388), .dinb(n301), .dout(n34666));
  jand g16644(.dina(n34666), .dinb(n34665), .dout(n34667));
  jor  g16645(.dina(n34667), .dinb(n34389), .dout(n34668));
  jxor g16646(.dina(n34383), .dinb(n293), .dout(n34669));
  jand g16647(.dina(n34669), .dinb(n34668), .dout(n34670));
  jor  g16648(.dina(n34670), .dinb(n34384), .dout(n34671));
  jxor g16649(.dina(n34378), .dinb(n294), .dout(n34672));
  jand g16650(.dina(n34672), .dinb(n34671), .dout(n34673));
  jor  g16651(.dina(n34673), .dinb(n34379), .dout(n34674));
  jxor g16652(.dina(n34373), .dinb(n290), .dout(n34675));
  jand g16653(.dina(n34675), .dinb(n34674), .dout(n34676));
  jor  g16654(.dina(n34676), .dinb(n34374), .dout(n34677));
  jxor g16655(.dina(n34368), .dinb(n291), .dout(n34678));
  jand g16656(.dina(n34678), .dinb(n34677), .dout(n34679));
  jor  g16657(.dina(n34679), .dinb(n34369), .dout(n34680));
  jxor g16658(.dina(n34363), .dinb(n284), .dout(n34681));
  jand g16659(.dina(n34681), .dinb(n34680), .dout(n34682));
  jor  g16660(.dina(n34682), .dinb(n34364), .dout(n34683));
  jxor g16661(.dina(n34358), .dinb(n285), .dout(n34684));
  jand g16662(.dina(n34684), .dinb(n34683), .dout(n34685));
  jor  g16663(.dina(n34685), .dinb(n34359), .dout(n34686));
  jxor g16664(.dina(n34353), .dinb(n281), .dout(n34687));
  jand g16665(.dina(n34687), .dinb(n34686), .dout(n34688));
  jor  g16666(.dina(n34688), .dinb(n34354), .dout(n34689));
  jxor g16667(.dina(n34348), .dinb(n282), .dout(n34690));
  jand g16668(.dina(n34690), .dinb(n34689), .dout(n34691));
  jor  g16669(.dina(n34691), .dinb(n34349), .dout(n34692));
  jxor g16670(.dina(n34343), .dinb(n397), .dout(n34693));
  jand g16671(.dina(n34693), .dinb(n34692), .dout(n34694));
  jor  g16672(.dina(n34694), .dinb(n34344), .dout(n34695));
  jxor g16673(.dina(n34338), .dinb(n513), .dout(n34696));
  jand g16674(.dina(n34696), .dinb(n34695), .dout(n34697));
  jor  g16675(.dina(n34697), .dinb(n34339), .dout(n34698));
  jxor g16676(.dina(n34333), .dinb(n514), .dout(n34699));
  jand g16677(.dina(n34699), .dinb(n34698), .dout(n34700));
  jor  g16678(.dina(n34700), .dinb(n34334), .dout(n34701));
  jxor g16679(.dina(n34328), .dinb(n510), .dout(n34702));
  jand g16680(.dina(n34702), .dinb(n34701), .dout(n34703));
  jor  g16681(.dina(n34703), .dinb(n34329), .dout(n34704));
  jxor g16682(.dina(n34323), .dinb(n396), .dout(n34705));
  jand g16683(.dina(n34705), .dinb(n34704), .dout(n34706));
  jor  g16684(.dina(n34706), .dinb(n34324), .dout(n34707));
  jxor g16685(.dina(n34318), .dinb(n383), .dout(n34708));
  jand g16686(.dina(n34708), .dinb(n34707), .dout(n34709));
  jor  g16687(.dina(n34709), .dinb(n34319), .dout(n34710));
  jxor g16688(.dina(n34313), .dinb(n12211), .dout(n34711));
  jand g16689(.dina(n34711), .dinb(n34710), .dout(n34712));
  jor  g16690(.dina(n34712), .dinb(n34314), .dout(n34713));
  jor  g16691(.dina(n34713), .dinb(n34308), .dout(n34714));
  jand g16692(.dina(n34714), .dinb(n34307), .dout(n34715));
  jand g16693(.dina(n34715), .dinb(n583), .dout(n34716));
  jnot g16694(.din(n34716), .dout(n34717));
  jand g16695(.dina(n34717), .dinb(n34305), .dout(n34718));
  jand g16696(.dina(n34308), .dinb(n583), .dout(n34719));
  jand g16697(.dina(n34719), .dinb(n34713), .dout(n34720));
  jor  g16698(.dina(n34720), .dinb(n34718), .dout(n34721));
  jnot g16699(.din(n34721), .dout(n34722));
  jand g16700(.dina(n34717), .dinb(n34313), .dout(n34723));
  jxor g16701(.dina(n34711), .dinb(n34710), .dout(n34724));
  jand g16702(.dina(n34724), .dinb(n34716), .dout(n34725));
  jor  g16703(.dina(n34725), .dinb(n34723), .dout(n34726));
  jand g16704(.dina(n34726), .dinb(n12214), .dout(n34727));
  jnot g16705(.din(n34727), .dout(n34728));
  jand g16706(.dina(n34717), .dinb(n34318), .dout(n34729));
  jxor g16707(.dina(n34708), .dinb(n34707), .dout(n34730));
  jand g16708(.dina(n34730), .dinb(n34716), .dout(n34731));
  jor  g16709(.dina(n34731), .dinb(n34729), .dout(n34732));
  jand g16710(.dina(n34732), .dinb(n12211), .dout(n34733));
  jnot g16711(.din(n34733), .dout(n34734));
  jand g16712(.dina(n34717), .dinb(n34323), .dout(n34735));
  jxor g16713(.dina(n34705), .dinb(n34704), .dout(n34736));
  jand g16714(.dina(n34736), .dinb(n34716), .dout(n34737));
  jor  g16715(.dina(n34737), .dinb(n34735), .dout(n34738));
  jand g16716(.dina(n34738), .dinb(n383), .dout(n34739));
  jnot g16717(.din(n34739), .dout(n34740));
  jand g16718(.dina(n34717), .dinb(n34328), .dout(n34741));
  jxor g16719(.dina(n34702), .dinb(n34701), .dout(n34742));
  jand g16720(.dina(n34742), .dinb(n34716), .dout(n34743));
  jor  g16721(.dina(n34743), .dinb(n34741), .dout(n34744));
  jand g16722(.dina(n34744), .dinb(n396), .dout(n34745));
  jnot g16723(.din(n34745), .dout(n34746));
  jand g16724(.dina(n34717), .dinb(n34333), .dout(n34747));
  jxor g16725(.dina(n34699), .dinb(n34698), .dout(n34748));
  jand g16726(.dina(n34748), .dinb(n34716), .dout(n34749));
  jor  g16727(.dina(n34749), .dinb(n34747), .dout(n34750));
  jand g16728(.dina(n34750), .dinb(n510), .dout(n34751));
  jnot g16729(.din(n34751), .dout(n34752));
  jand g16730(.dina(n34717), .dinb(n34338), .dout(n34753));
  jxor g16731(.dina(n34696), .dinb(n34695), .dout(n34754));
  jand g16732(.dina(n34754), .dinb(n34716), .dout(n34755));
  jor  g16733(.dina(n34755), .dinb(n34753), .dout(n34756));
  jand g16734(.dina(n34756), .dinb(n514), .dout(n34757));
  jnot g16735(.din(n34757), .dout(n34758));
  jand g16736(.dina(n34717), .dinb(n34343), .dout(n34759));
  jxor g16737(.dina(n34693), .dinb(n34692), .dout(n34760));
  jand g16738(.dina(n34760), .dinb(n34716), .dout(n34761));
  jor  g16739(.dina(n34761), .dinb(n34759), .dout(n34762));
  jand g16740(.dina(n34762), .dinb(n513), .dout(n34763));
  jnot g16741(.din(n34763), .dout(n34764));
  jand g16742(.dina(n34717), .dinb(n34348), .dout(n34765));
  jxor g16743(.dina(n34690), .dinb(n34689), .dout(n34766));
  jand g16744(.dina(n34766), .dinb(n34716), .dout(n34767));
  jor  g16745(.dina(n34767), .dinb(n34765), .dout(n34768));
  jand g16746(.dina(n34768), .dinb(n397), .dout(n34769));
  jnot g16747(.din(n34769), .dout(n34770));
  jand g16748(.dina(n34717), .dinb(n34353), .dout(n34771));
  jxor g16749(.dina(n34687), .dinb(n34686), .dout(n34772));
  jand g16750(.dina(n34772), .dinb(n34716), .dout(n34773));
  jor  g16751(.dina(n34773), .dinb(n34771), .dout(n34774));
  jand g16752(.dina(n34774), .dinb(n282), .dout(n34775));
  jnot g16753(.din(n34775), .dout(n34776));
  jand g16754(.dina(n34717), .dinb(n34358), .dout(n34777));
  jxor g16755(.dina(n34684), .dinb(n34683), .dout(n34778));
  jand g16756(.dina(n34778), .dinb(n34716), .dout(n34779));
  jor  g16757(.dina(n34779), .dinb(n34777), .dout(n34780));
  jand g16758(.dina(n34780), .dinb(n281), .dout(n34781));
  jnot g16759(.din(n34781), .dout(n34782));
  jand g16760(.dina(n34717), .dinb(n34363), .dout(n34783));
  jxor g16761(.dina(n34681), .dinb(n34680), .dout(n34784));
  jand g16762(.dina(n34784), .dinb(n34716), .dout(n34785));
  jor  g16763(.dina(n34785), .dinb(n34783), .dout(n34786));
  jand g16764(.dina(n34786), .dinb(n285), .dout(n34787));
  jnot g16765(.din(n34787), .dout(n34788));
  jand g16766(.dina(n34717), .dinb(n34368), .dout(n34789));
  jxor g16767(.dina(n34678), .dinb(n34677), .dout(n34790));
  jand g16768(.dina(n34790), .dinb(n34716), .dout(n34791));
  jor  g16769(.dina(n34791), .dinb(n34789), .dout(n34792));
  jand g16770(.dina(n34792), .dinb(n284), .dout(n34793));
  jnot g16771(.din(n34793), .dout(n34794));
  jand g16772(.dina(n34717), .dinb(n34373), .dout(n34795));
  jxor g16773(.dina(n34675), .dinb(n34674), .dout(n34796));
  jand g16774(.dina(n34796), .dinb(n34716), .dout(n34797));
  jor  g16775(.dina(n34797), .dinb(n34795), .dout(n34798));
  jand g16776(.dina(n34798), .dinb(n291), .dout(n34799));
  jnot g16777(.din(n34799), .dout(n34800));
  jand g16778(.dina(n34717), .dinb(n34378), .dout(n34801));
  jxor g16779(.dina(n34672), .dinb(n34671), .dout(n34802));
  jand g16780(.dina(n34802), .dinb(n34716), .dout(n34803));
  jor  g16781(.dina(n34803), .dinb(n34801), .dout(n34804));
  jand g16782(.dina(n34804), .dinb(n290), .dout(n34805));
  jnot g16783(.din(n34805), .dout(n34806));
  jand g16784(.dina(n34717), .dinb(n34383), .dout(n34807));
  jxor g16785(.dina(n34669), .dinb(n34668), .dout(n34808));
  jand g16786(.dina(n34808), .dinb(n34716), .dout(n34809));
  jor  g16787(.dina(n34809), .dinb(n34807), .dout(n34810));
  jand g16788(.dina(n34810), .dinb(n294), .dout(n34811));
  jnot g16789(.din(n34811), .dout(n34812));
  jand g16790(.dina(n34717), .dinb(n34388), .dout(n34813));
  jxor g16791(.dina(n34666), .dinb(n34665), .dout(n34814));
  jand g16792(.dina(n34814), .dinb(n34716), .dout(n34815));
  jor  g16793(.dina(n34815), .dinb(n34813), .dout(n34816));
  jand g16794(.dina(n34816), .dinb(n293), .dout(n34817));
  jnot g16795(.din(n34817), .dout(n34818));
  jand g16796(.dina(n34717), .dinb(n34393), .dout(n34819));
  jxor g16797(.dina(n34663), .dinb(n34662), .dout(n34820));
  jand g16798(.dina(n34820), .dinb(n34716), .dout(n34821));
  jor  g16799(.dina(n34821), .dinb(n34819), .dout(n34822));
  jand g16800(.dina(n34822), .dinb(n301), .dout(n34823));
  jnot g16801(.din(n34823), .dout(n34824));
  jand g16802(.dina(n34717), .dinb(n34398), .dout(n34825));
  jxor g16803(.dina(n34660), .dinb(n34659), .dout(n34826));
  jand g16804(.dina(n34826), .dinb(n34716), .dout(n34827));
  jor  g16805(.dina(n34827), .dinb(n34825), .dout(n34828));
  jand g16806(.dina(n34828), .dinb(n298), .dout(n34829));
  jnot g16807(.din(n34829), .dout(n34830));
  jand g16808(.dina(n34717), .dinb(n34403), .dout(n34831));
  jxor g16809(.dina(n34657), .dinb(n34656), .dout(n34832));
  jand g16810(.dina(n34832), .dinb(n34716), .dout(n34833));
  jor  g16811(.dina(n34833), .dinb(n34831), .dout(n34834));
  jand g16812(.dina(n34834), .dinb(n297), .dout(n34835));
  jnot g16813(.din(n34835), .dout(n34836));
  jand g16814(.dina(n34717), .dinb(n34408), .dout(n34837));
  jxor g16815(.dina(n34654), .dinb(n34653), .dout(n34838));
  jand g16816(.dina(n34838), .dinb(n34716), .dout(n34839));
  jor  g16817(.dina(n34839), .dinb(n34837), .dout(n34840));
  jand g16818(.dina(n34840), .dinb(n300), .dout(n34841));
  jnot g16819(.din(n34841), .dout(n34842));
  jand g16820(.dina(n34717), .dinb(n34413), .dout(n34843));
  jxor g16821(.dina(n34651), .dinb(n34650), .dout(n34844));
  jand g16822(.dina(n34844), .dinb(n34716), .dout(n34845));
  jor  g16823(.dina(n34845), .dinb(n34843), .dout(n34846));
  jand g16824(.dina(n34846), .dinb(n424), .dout(n34847));
  jnot g16825(.din(n34847), .dout(n34848));
  jand g16826(.dina(n34717), .dinb(n34418), .dout(n34849));
  jxor g16827(.dina(n34648), .dinb(n34647), .dout(n34850));
  jand g16828(.dina(n34850), .dinb(n34716), .dout(n34851));
  jor  g16829(.dina(n34851), .dinb(n34849), .dout(n34852));
  jand g16830(.dina(n34852), .dinb(n427), .dout(n34853));
  jnot g16831(.din(n34853), .dout(n34854));
  jand g16832(.dina(n34717), .dinb(n34423), .dout(n34855));
  jxor g16833(.dina(n34645), .dinb(n34644), .dout(n34856));
  jand g16834(.dina(n34856), .dinb(n34716), .dout(n34857));
  jor  g16835(.dina(n34857), .dinb(n34855), .dout(n34858));
  jand g16836(.dina(n34858), .dinb(n426), .dout(n34859));
  jnot g16837(.din(n34859), .dout(n34860));
  jand g16838(.dina(n34717), .dinb(n34428), .dout(n34861));
  jxor g16839(.dina(n34642), .dinb(n34641), .dout(n34862));
  jand g16840(.dina(n34862), .dinb(n34716), .dout(n34863));
  jor  g16841(.dina(n34863), .dinb(n34861), .dout(n34864));
  jand g16842(.dina(n34864), .dinb(n410), .dout(n34865));
  jnot g16843(.din(n34865), .dout(n34866));
  jand g16844(.dina(n34717), .dinb(n34433), .dout(n34867));
  jxor g16845(.dina(n34639), .dinb(n34638), .dout(n34868));
  jand g16846(.dina(n34868), .dinb(n34716), .dout(n34869));
  jor  g16847(.dina(n34869), .dinb(n34867), .dout(n34870));
  jand g16848(.dina(n34870), .dinb(n409), .dout(n34871));
  jnot g16849(.din(n34871), .dout(n34872));
  jand g16850(.dina(n34717), .dinb(n34438), .dout(n34873));
  jxor g16851(.dina(n34636), .dinb(n34635), .dout(n34874));
  jand g16852(.dina(n34874), .dinb(n34716), .dout(n34875));
  jor  g16853(.dina(n34875), .dinb(n34873), .dout(n34876));
  jand g16854(.dina(n34876), .dinb(n413), .dout(n34877));
  jnot g16855(.din(n34877), .dout(n34878));
  jand g16856(.dina(n34717), .dinb(n34443), .dout(n34879));
  jxor g16857(.dina(n34633), .dinb(n34632), .dout(n34880));
  jand g16858(.dina(n34880), .dinb(n34716), .dout(n34881));
  jor  g16859(.dina(n34881), .dinb(n34879), .dout(n34882));
  jand g16860(.dina(n34882), .dinb(n412), .dout(n34883));
  jnot g16861(.din(n34883), .dout(n34884));
  jand g16862(.dina(n34717), .dinb(n34448), .dout(n34885));
  jxor g16863(.dina(n34630), .dinb(n34629), .dout(n34886));
  jand g16864(.dina(n34886), .dinb(n34716), .dout(n34887));
  jor  g16865(.dina(n34887), .dinb(n34885), .dout(n34888));
  jand g16866(.dina(n34888), .dinb(n406), .dout(n34889));
  jnot g16867(.din(n34889), .dout(n34890));
  jand g16868(.dina(n34717), .dinb(n34453), .dout(n34891));
  jxor g16869(.dina(n34627), .dinb(n34626), .dout(n34892));
  jand g16870(.dina(n34892), .dinb(n34716), .dout(n34893));
  jor  g16871(.dina(n34893), .dinb(n34891), .dout(n34894));
  jand g16872(.dina(n34894), .dinb(n405), .dout(n34895));
  jnot g16873(.din(n34895), .dout(n34896));
  jand g16874(.dina(n34717), .dinb(n34458), .dout(n34897));
  jxor g16875(.dina(n34624), .dinb(n34623), .dout(n34898));
  jand g16876(.dina(n34898), .dinb(n34716), .dout(n34899));
  jor  g16877(.dina(n34899), .dinb(n34897), .dout(n34900));
  jand g16878(.dina(n34900), .dinb(n2714), .dout(n34901));
  jnot g16879(.din(n34901), .dout(n34902));
  jand g16880(.dina(n34717), .dinb(n34463), .dout(n34903));
  jxor g16881(.dina(n34621), .dinb(n34620), .dout(n34904));
  jand g16882(.dina(n34904), .dinb(n34716), .dout(n34905));
  jor  g16883(.dina(n34905), .dinb(n34903), .dout(n34906));
  jand g16884(.dina(n34906), .dinb(n2547), .dout(n34907));
  jnot g16885(.din(n34907), .dout(n34908));
  jand g16886(.dina(n34717), .dinb(n34468), .dout(n34909));
  jxor g16887(.dina(n34618), .dinb(n34617), .dout(n34910));
  jand g16888(.dina(n34910), .dinb(n34716), .dout(n34911));
  jor  g16889(.dina(n34911), .dinb(n34909), .dout(n34912));
  jand g16890(.dina(n34912), .dinb(n417), .dout(n34913));
  jnot g16891(.din(n34913), .dout(n34914));
  jand g16892(.dina(n34717), .dinb(n34473), .dout(n34915));
  jxor g16893(.dina(n34615), .dinb(n34614), .dout(n34916));
  jand g16894(.dina(n34916), .dinb(n34716), .dout(n34917));
  jor  g16895(.dina(n34917), .dinb(n34915), .dout(n34918));
  jand g16896(.dina(n34918), .dinb(n416), .dout(n34919));
  jnot g16897(.din(n34919), .dout(n34920));
  jand g16898(.dina(n34717), .dinb(n34478), .dout(n34921));
  jxor g16899(.dina(n34612), .dinb(n34611), .dout(n34922));
  jand g16900(.dina(n34922), .dinb(n34716), .dout(n34923));
  jor  g16901(.dina(n34923), .dinb(n34921), .dout(n34924));
  jand g16902(.dina(n34924), .dinb(n422), .dout(n34925));
  jnot g16903(.din(n34925), .dout(n34926));
  jand g16904(.dina(n34717), .dinb(n34483), .dout(n34927));
  jxor g16905(.dina(n34609), .dinb(n34608), .dout(n34928));
  jand g16906(.dina(n34928), .dinb(n34716), .dout(n34929));
  jor  g16907(.dina(n34929), .dinb(n34927), .dout(n34930));
  jand g16908(.dina(n34930), .dinb(n421), .dout(n34931));
  jnot g16909(.din(n34931), .dout(n34932));
  jand g16910(.dina(n34717), .dinb(n34488), .dout(n34933));
  jxor g16911(.dina(n34606), .dinb(n34605), .dout(n34934));
  jand g16912(.dina(n34934), .dinb(n34716), .dout(n34935));
  jor  g16913(.dina(n34935), .dinb(n34933), .dout(n34936));
  jand g16914(.dina(n34936), .dinb(n433), .dout(n34937));
  jnot g16915(.din(n34937), .dout(n34938));
  jand g16916(.dina(n34717), .dinb(n34493), .dout(n34939));
  jxor g16917(.dina(n34603), .dinb(n34602), .dout(n34940));
  jand g16918(.dina(n34940), .dinb(n34716), .dout(n34941));
  jor  g16919(.dina(n34941), .dinb(n34939), .dout(n34942));
  jand g16920(.dina(n34942), .dinb(n432), .dout(n34943));
  jnot g16921(.din(n34943), .dout(n34944));
  jand g16922(.dina(n34717), .dinb(n34498), .dout(n34945));
  jxor g16923(.dina(n34600), .dinb(n34599), .dout(n34946));
  jand g16924(.dina(n34946), .dinb(n34716), .dout(n34947));
  jor  g16925(.dina(n34947), .dinb(n34945), .dout(n34948));
  jand g16926(.dina(n34948), .dinb(n436), .dout(n34949));
  jnot g16927(.din(n34949), .dout(n34950));
  jand g16928(.dina(n34717), .dinb(n34503), .dout(n34951));
  jxor g16929(.dina(n34597), .dinb(n34596), .dout(n34952));
  jand g16930(.dina(n34952), .dinb(n34716), .dout(n34953));
  jor  g16931(.dina(n34953), .dinb(n34951), .dout(n34954));
  jand g16932(.dina(n34954), .dinb(n435), .dout(n34955));
  jnot g16933(.din(n34955), .dout(n34956));
  jand g16934(.dina(n34717), .dinb(n34508), .dout(n34957));
  jxor g16935(.dina(n34594), .dinb(n34593), .dout(n34958));
  jand g16936(.dina(n34958), .dinb(n34716), .dout(n34959));
  jor  g16937(.dina(n34959), .dinb(n34957), .dout(n34960));
  jand g16938(.dina(n34960), .dinb(n440), .dout(n34961));
  jnot g16939(.din(n34961), .dout(n34962));
  jand g16940(.dina(n34717), .dinb(n34513), .dout(n34963));
  jxor g16941(.dina(n34591), .dinb(n34590), .dout(n34964));
  jand g16942(.dina(n34964), .dinb(n34716), .dout(n34965));
  jor  g16943(.dina(n34965), .dinb(n34963), .dout(n34966));
  jand g16944(.dina(n34966), .dinb(n439), .dout(n34967));
  jnot g16945(.din(n34967), .dout(n34968));
  jand g16946(.dina(n34717), .dinb(n34518), .dout(n34969));
  jxor g16947(.dina(n34588), .dinb(n34587), .dout(n34970));
  jand g16948(.dina(n34970), .dinb(n34716), .dout(n34971));
  jor  g16949(.dina(n34971), .dinb(n34969), .dout(n34972));
  jand g16950(.dina(n34972), .dinb(n325), .dout(n34973));
  jnot g16951(.din(n34973), .dout(n34974));
  jand g16952(.dina(n34717), .dinb(n34523), .dout(n34975));
  jxor g16953(.dina(n34585), .dinb(n34584), .dout(n34976));
  jand g16954(.dina(n34976), .dinb(n34716), .dout(n34977));
  jor  g16955(.dina(n34977), .dinb(n34975), .dout(n34978));
  jand g16956(.dina(n34978), .dinb(n324), .dout(n34979));
  jnot g16957(.din(n34979), .dout(n34980));
  jand g16958(.dina(n34717), .dinb(n34528), .dout(n34981));
  jxor g16959(.dina(n34582), .dinb(n34581), .dout(n34982));
  jand g16960(.dina(n34982), .dinb(n34716), .dout(n34983));
  jor  g16961(.dina(n34983), .dinb(n34981), .dout(n34984));
  jand g16962(.dina(n34984), .dinb(n323), .dout(n34985));
  jnot g16963(.din(n34985), .dout(n34986));
  jand g16964(.dina(n34717), .dinb(n34533), .dout(n34987));
  jxor g16965(.dina(n34579), .dinb(n34578), .dout(n34988));
  jand g16966(.dina(n34988), .dinb(n34716), .dout(n34989));
  jor  g16967(.dina(n34989), .dinb(n34987), .dout(n34990));
  jand g16968(.dina(n34990), .dinb(n335), .dout(n34991));
  jnot g16969(.din(n34991), .dout(n34992));
  jand g16970(.dina(n34717), .dinb(n34538), .dout(n34993));
  jxor g16971(.dina(n34576), .dinb(n34575), .dout(n34994));
  jand g16972(.dina(n34994), .dinb(n34716), .dout(n34995));
  jor  g16973(.dina(n34995), .dinb(n34993), .dout(n34996));
  jand g16974(.dina(n34996), .dinb(n334), .dout(n34997));
  jnot g16975(.din(n34997), .dout(n34998));
  jand g16976(.dina(n34717), .dinb(n34543), .dout(n34999));
  jxor g16977(.dina(n34573), .dinb(n34572), .dout(n35000));
  jand g16978(.dina(n35000), .dinb(n34716), .dout(n35001));
  jor  g16979(.dina(n35001), .dinb(n34999), .dout(n35002));
  jand g16980(.dina(n35002), .dinb(n338), .dout(n35003));
  jnot g16981(.din(n35003), .dout(n35004));
  jand g16982(.dina(n34717), .dinb(n34548), .dout(n35005));
  jxor g16983(.dina(n34570), .dinb(n34569), .dout(n35006));
  jand g16984(.dina(n35006), .dinb(n34716), .dout(n35007));
  jor  g16985(.dina(n35007), .dinb(n35005), .dout(n35008));
  jand g16986(.dina(n35008), .dinb(n337), .dout(n35009));
  jnot g16987(.din(n35009), .dout(n35010));
  jnot g16988(.din(n34553), .dout(n35011));
  jor  g16989(.dina(n34716), .dinb(n35011), .dout(n35012));
  jxor g16990(.dina(n34567), .dinb(n34566), .dout(n35013));
  jnot g16991(.din(n35013), .dout(n35014));
  jor  g16992(.dina(n35014), .dinb(n34717), .dout(n35015));
  jand g16993(.dina(n35015), .dinb(n35012), .dout(n35016));
  jnot g16994(.din(n35016), .dout(n35017));
  jand g16995(.dina(n35017), .dinb(n344), .dout(n35018));
  jnot g16996(.din(n35018), .dout(n35019));
  jor  g16997(.dina(n34716), .dinb(n34563), .dout(n35020));
  jxor g16998(.dina(n34564), .dinb(n12487), .dout(n35021));
  jand g16999(.dina(n35021), .dinb(n34716), .dout(n35022));
  jnot g17000(.din(n35022), .dout(n35023));
  jand g17001(.dina(n35023), .dinb(n35020), .dout(n35024));
  jnot g17002(.din(n35024), .dout(n35025));
  jand g17003(.dina(n35025), .dinb(n348), .dout(n35026));
  jnot g17004(.din(n35026), .dout(n35027));
  jnot g17005(.din(n12895), .dout(n35028));
  jnot g17006(.din(n34308), .dout(n35029));
  jnot g17007(.din(n34314), .dout(n35030));
  jnot g17008(.din(n34319), .dout(n35031));
  jnot g17009(.din(n34324), .dout(n35032));
  jnot g17010(.din(n34329), .dout(n35033));
  jnot g17011(.din(n34334), .dout(n35034));
  jnot g17012(.din(n34339), .dout(n35035));
  jnot g17013(.din(n34344), .dout(n35036));
  jnot g17014(.din(n34349), .dout(n35037));
  jnot g17015(.din(n34354), .dout(n35038));
  jnot g17016(.din(n34359), .dout(n35039));
  jnot g17017(.din(n34364), .dout(n35040));
  jnot g17018(.din(n34369), .dout(n35041));
  jnot g17019(.din(n34374), .dout(n35042));
  jnot g17020(.din(n34379), .dout(n35043));
  jnot g17021(.din(n34384), .dout(n35044));
  jnot g17022(.din(n34389), .dout(n35045));
  jnot g17023(.din(n34394), .dout(n35046));
  jnot g17024(.din(n34399), .dout(n35047));
  jnot g17025(.din(n34404), .dout(n35048));
  jnot g17026(.din(n34409), .dout(n35049));
  jnot g17027(.din(n34414), .dout(n35050));
  jnot g17028(.din(n34419), .dout(n35051));
  jnot g17029(.din(n34424), .dout(n35052));
  jnot g17030(.din(n34429), .dout(n35053));
  jnot g17031(.din(n34434), .dout(n35054));
  jnot g17032(.din(n34439), .dout(n35055));
  jnot g17033(.din(n34444), .dout(n35056));
  jnot g17034(.din(n34449), .dout(n35057));
  jnot g17035(.din(n34454), .dout(n35058));
  jnot g17036(.din(n34459), .dout(n35059));
  jnot g17037(.din(n34464), .dout(n35060));
  jnot g17038(.din(n34469), .dout(n35061));
  jnot g17039(.din(n34474), .dout(n35062));
  jnot g17040(.din(n34479), .dout(n35063));
  jnot g17041(.din(n34484), .dout(n35064));
  jnot g17042(.din(n34489), .dout(n35065));
  jnot g17043(.din(n34494), .dout(n35066));
  jnot g17044(.din(n34499), .dout(n35067));
  jnot g17045(.din(n34504), .dout(n35068));
  jnot g17046(.din(n34509), .dout(n35069));
  jnot g17047(.din(n34514), .dout(n35070));
  jnot g17048(.din(n34519), .dout(n35071));
  jnot g17049(.din(n34524), .dout(n35072));
  jnot g17050(.din(n34529), .dout(n35073));
  jnot g17051(.din(n34534), .dout(n35074));
  jnot g17052(.din(n34539), .dout(n35075));
  jnot g17053(.din(n34544), .dout(n35076));
  jnot g17054(.din(n34549), .dout(n35077));
  jnot g17055(.din(n34554), .dout(n35078));
  jnot g17056(.din(n34560), .dout(n35079));
  jxor g17057(.dina(n34563), .dinb(n258), .dout(n35080));
  jor  g17058(.dina(n35080), .dinb(n12486), .dout(n35081));
  jand g17059(.dina(n35081), .dinb(n35079), .dout(n35082));
  jnot g17060(.din(n34567), .dout(n35083));
  jor  g17061(.dina(n35083), .dinb(n35082), .dout(n35084));
  jand g17062(.dina(n35084), .dinb(n35078), .dout(n35085));
  jnot g17063(.din(n34570), .dout(n35086));
  jor  g17064(.dina(n35086), .dinb(n35085), .dout(n35087));
  jand g17065(.dina(n35087), .dinb(n35077), .dout(n35088));
  jnot g17066(.din(n34573), .dout(n35089));
  jor  g17067(.dina(n35089), .dinb(n35088), .dout(n35090));
  jand g17068(.dina(n35090), .dinb(n35076), .dout(n35091));
  jnot g17069(.din(n34576), .dout(n35092));
  jor  g17070(.dina(n35092), .dinb(n35091), .dout(n35093));
  jand g17071(.dina(n35093), .dinb(n35075), .dout(n35094));
  jnot g17072(.din(n34579), .dout(n35095));
  jor  g17073(.dina(n35095), .dinb(n35094), .dout(n35096));
  jand g17074(.dina(n35096), .dinb(n35074), .dout(n35097));
  jnot g17075(.din(n34582), .dout(n35098));
  jor  g17076(.dina(n35098), .dinb(n35097), .dout(n35099));
  jand g17077(.dina(n35099), .dinb(n35073), .dout(n35100));
  jnot g17078(.din(n34585), .dout(n35101));
  jor  g17079(.dina(n35101), .dinb(n35100), .dout(n35102));
  jand g17080(.dina(n35102), .dinb(n35072), .dout(n35103));
  jnot g17081(.din(n34588), .dout(n35104));
  jor  g17082(.dina(n35104), .dinb(n35103), .dout(n35105));
  jand g17083(.dina(n35105), .dinb(n35071), .dout(n35106));
  jnot g17084(.din(n34591), .dout(n35107));
  jor  g17085(.dina(n35107), .dinb(n35106), .dout(n35108));
  jand g17086(.dina(n35108), .dinb(n35070), .dout(n35109));
  jnot g17087(.din(n34594), .dout(n35110));
  jor  g17088(.dina(n35110), .dinb(n35109), .dout(n35111));
  jand g17089(.dina(n35111), .dinb(n35069), .dout(n35112));
  jnot g17090(.din(n34597), .dout(n35113));
  jor  g17091(.dina(n35113), .dinb(n35112), .dout(n35114));
  jand g17092(.dina(n35114), .dinb(n35068), .dout(n35115));
  jnot g17093(.din(n34600), .dout(n35116));
  jor  g17094(.dina(n35116), .dinb(n35115), .dout(n35117));
  jand g17095(.dina(n35117), .dinb(n35067), .dout(n35118));
  jnot g17096(.din(n34603), .dout(n35119));
  jor  g17097(.dina(n35119), .dinb(n35118), .dout(n35120));
  jand g17098(.dina(n35120), .dinb(n35066), .dout(n35121));
  jnot g17099(.din(n34606), .dout(n35122));
  jor  g17100(.dina(n35122), .dinb(n35121), .dout(n35123));
  jand g17101(.dina(n35123), .dinb(n35065), .dout(n35124));
  jnot g17102(.din(n34609), .dout(n35125));
  jor  g17103(.dina(n35125), .dinb(n35124), .dout(n35126));
  jand g17104(.dina(n35126), .dinb(n35064), .dout(n35127));
  jnot g17105(.din(n34612), .dout(n35128));
  jor  g17106(.dina(n35128), .dinb(n35127), .dout(n35129));
  jand g17107(.dina(n35129), .dinb(n35063), .dout(n35130));
  jnot g17108(.din(n34615), .dout(n35131));
  jor  g17109(.dina(n35131), .dinb(n35130), .dout(n35132));
  jand g17110(.dina(n35132), .dinb(n35062), .dout(n35133));
  jnot g17111(.din(n34618), .dout(n35134));
  jor  g17112(.dina(n35134), .dinb(n35133), .dout(n35135));
  jand g17113(.dina(n35135), .dinb(n35061), .dout(n35136));
  jnot g17114(.din(n34621), .dout(n35137));
  jor  g17115(.dina(n35137), .dinb(n35136), .dout(n35138));
  jand g17116(.dina(n35138), .dinb(n35060), .dout(n35139));
  jnot g17117(.din(n34624), .dout(n35140));
  jor  g17118(.dina(n35140), .dinb(n35139), .dout(n35141));
  jand g17119(.dina(n35141), .dinb(n35059), .dout(n35142));
  jnot g17120(.din(n34627), .dout(n35143));
  jor  g17121(.dina(n35143), .dinb(n35142), .dout(n35144));
  jand g17122(.dina(n35144), .dinb(n35058), .dout(n35145));
  jnot g17123(.din(n34630), .dout(n35146));
  jor  g17124(.dina(n35146), .dinb(n35145), .dout(n35147));
  jand g17125(.dina(n35147), .dinb(n35057), .dout(n35148));
  jnot g17126(.din(n34633), .dout(n35149));
  jor  g17127(.dina(n35149), .dinb(n35148), .dout(n35150));
  jand g17128(.dina(n35150), .dinb(n35056), .dout(n35151));
  jnot g17129(.din(n34636), .dout(n35152));
  jor  g17130(.dina(n35152), .dinb(n35151), .dout(n35153));
  jand g17131(.dina(n35153), .dinb(n35055), .dout(n35154));
  jnot g17132(.din(n34639), .dout(n35155));
  jor  g17133(.dina(n35155), .dinb(n35154), .dout(n35156));
  jand g17134(.dina(n35156), .dinb(n35054), .dout(n35157));
  jnot g17135(.din(n34642), .dout(n35158));
  jor  g17136(.dina(n35158), .dinb(n35157), .dout(n35159));
  jand g17137(.dina(n35159), .dinb(n35053), .dout(n35160));
  jnot g17138(.din(n34645), .dout(n35161));
  jor  g17139(.dina(n35161), .dinb(n35160), .dout(n35162));
  jand g17140(.dina(n35162), .dinb(n35052), .dout(n35163));
  jnot g17141(.din(n34648), .dout(n35164));
  jor  g17142(.dina(n35164), .dinb(n35163), .dout(n35165));
  jand g17143(.dina(n35165), .dinb(n35051), .dout(n35166));
  jnot g17144(.din(n34651), .dout(n35167));
  jor  g17145(.dina(n35167), .dinb(n35166), .dout(n35168));
  jand g17146(.dina(n35168), .dinb(n35050), .dout(n35169));
  jnot g17147(.din(n34654), .dout(n35170));
  jor  g17148(.dina(n35170), .dinb(n35169), .dout(n35171));
  jand g17149(.dina(n35171), .dinb(n35049), .dout(n35172));
  jnot g17150(.din(n34657), .dout(n35173));
  jor  g17151(.dina(n35173), .dinb(n35172), .dout(n35174));
  jand g17152(.dina(n35174), .dinb(n35048), .dout(n35175));
  jnot g17153(.din(n34660), .dout(n35176));
  jor  g17154(.dina(n35176), .dinb(n35175), .dout(n35177));
  jand g17155(.dina(n35177), .dinb(n35047), .dout(n35178));
  jnot g17156(.din(n34663), .dout(n35179));
  jor  g17157(.dina(n35179), .dinb(n35178), .dout(n35180));
  jand g17158(.dina(n35180), .dinb(n35046), .dout(n35181));
  jnot g17159(.din(n34666), .dout(n35182));
  jor  g17160(.dina(n35182), .dinb(n35181), .dout(n35183));
  jand g17161(.dina(n35183), .dinb(n35045), .dout(n35184));
  jnot g17162(.din(n34669), .dout(n35185));
  jor  g17163(.dina(n35185), .dinb(n35184), .dout(n35186));
  jand g17164(.dina(n35186), .dinb(n35044), .dout(n35187));
  jnot g17165(.din(n34672), .dout(n35188));
  jor  g17166(.dina(n35188), .dinb(n35187), .dout(n35189));
  jand g17167(.dina(n35189), .dinb(n35043), .dout(n35190));
  jnot g17168(.din(n34675), .dout(n35191));
  jor  g17169(.dina(n35191), .dinb(n35190), .dout(n35192));
  jand g17170(.dina(n35192), .dinb(n35042), .dout(n35193));
  jnot g17171(.din(n34678), .dout(n35194));
  jor  g17172(.dina(n35194), .dinb(n35193), .dout(n35195));
  jand g17173(.dina(n35195), .dinb(n35041), .dout(n35196));
  jnot g17174(.din(n34681), .dout(n35197));
  jor  g17175(.dina(n35197), .dinb(n35196), .dout(n35198));
  jand g17176(.dina(n35198), .dinb(n35040), .dout(n35199));
  jnot g17177(.din(n34684), .dout(n35200));
  jor  g17178(.dina(n35200), .dinb(n35199), .dout(n35201));
  jand g17179(.dina(n35201), .dinb(n35039), .dout(n35202));
  jnot g17180(.din(n34687), .dout(n35203));
  jor  g17181(.dina(n35203), .dinb(n35202), .dout(n35204));
  jand g17182(.dina(n35204), .dinb(n35038), .dout(n35205));
  jnot g17183(.din(n34690), .dout(n35206));
  jor  g17184(.dina(n35206), .dinb(n35205), .dout(n35207));
  jand g17185(.dina(n35207), .dinb(n35037), .dout(n35208));
  jnot g17186(.din(n34693), .dout(n35209));
  jor  g17187(.dina(n35209), .dinb(n35208), .dout(n35210));
  jand g17188(.dina(n35210), .dinb(n35036), .dout(n35211));
  jnot g17189(.din(n34696), .dout(n35212));
  jor  g17190(.dina(n35212), .dinb(n35211), .dout(n35213));
  jand g17191(.dina(n35213), .dinb(n35035), .dout(n35214));
  jnot g17192(.din(n34699), .dout(n35215));
  jor  g17193(.dina(n35215), .dinb(n35214), .dout(n35216));
  jand g17194(.dina(n35216), .dinb(n35034), .dout(n35217));
  jnot g17195(.din(n34702), .dout(n35218));
  jor  g17196(.dina(n35218), .dinb(n35217), .dout(n35219));
  jand g17197(.dina(n35219), .dinb(n35033), .dout(n35220));
  jnot g17198(.din(n34705), .dout(n35221));
  jor  g17199(.dina(n35221), .dinb(n35220), .dout(n35222));
  jand g17200(.dina(n35222), .dinb(n35032), .dout(n35223));
  jnot g17201(.din(n34708), .dout(n35224));
  jor  g17202(.dina(n35224), .dinb(n35223), .dout(n35225));
  jand g17203(.dina(n35225), .dinb(n35031), .dout(n35226));
  jnot g17204(.din(n34711), .dout(n35227));
  jor  g17205(.dina(n35227), .dinb(n35226), .dout(n35228));
  jand g17206(.dina(n35228), .dinb(n35030), .dout(n35229));
  jand g17207(.dina(n35229), .dinb(n35029), .dout(n35230));
  jor  g17208(.dina(n35230), .dinb(n34306), .dout(n35231));
  jor  g17209(.dina(n35231), .dinb(n35028), .dout(n35232));
  jand g17210(.dina(n35232), .dinb(a12 ), .dout(n35233));
  jnot g17211(.din(n12898), .dout(n35234));
  jor  g17212(.dina(n35231), .dinb(n35234), .dout(n35235));
  jnot g17213(.din(n35235), .dout(n35236));
  jor  g17214(.dina(n35236), .dinb(n35233), .dout(n35237));
  jand g17215(.dina(n35237), .dinb(n258), .dout(n35238));
  jnot g17216(.din(n35238), .dout(n35239));
  jand g17217(.dina(n34715), .dinb(n12895), .dout(n35240));
  jor  g17218(.dina(n35240), .dinb(n12485), .dout(n35241));
  jand g17219(.dina(n35235), .dinb(n35241), .dout(n35242));
  jxor g17220(.dina(n35242), .dinb(n258), .dout(n35243));
  jor  g17221(.dina(n35243), .dinb(n12905), .dout(n35244));
  jand g17222(.dina(n35244), .dinb(n35239), .dout(n35245));
  jxor g17223(.dina(n35024), .dinb(b2 ), .dout(n35246));
  jnot g17224(.din(n35246), .dout(n35247));
  jor  g17225(.dina(n35247), .dinb(n35245), .dout(n35248));
  jand g17226(.dina(n35248), .dinb(n35027), .dout(n35249));
  jxor g17227(.dina(n35016), .dinb(b3 ), .dout(n35250));
  jnot g17228(.din(n35250), .dout(n35251));
  jor  g17229(.dina(n35251), .dinb(n35249), .dout(n35252));
  jand g17230(.dina(n35252), .dinb(n35019), .dout(n35253));
  jxor g17231(.dina(n35008), .dinb(n337), .dout(n35254));
  jnot g17232(.din(n35254), .dout(n35255));
  jor  g17233(.dina(n35255), .dinb(n35253), .dout(n35256));
  jand g17234(.dina(n35256), .dinb(n35010), .dout(n35257));
  jxor g17235(.dina(n35002), .dinb(n338), .dout(n35258));
  jnot g17236(.din(n35258), .dout(n35259));
  jor  g17237(.dina(n35259), .dinb(n35257), .dout(n35260));
  jand g17238(.dina(n35260), .dinb(n35004), .dout(n35261));
  jxor g17239(.dina(n34996), .dinb(n334), .dout(n35262));
  jnot g17240(.din(n35262), .dout(n35263));
  jor  g17241(.dina(n35263), .dinb(n35261), .dout(n35264));
  jand g17242(.dina(n35264), .dinb(n34998), .dout(n35265));
  jxor g17243(.dina(n34990), .dinb(n335), .dout(n35266));
  jnot g17244(.din(n35266), .dout(n35267));
  jor  g17245(.dina(n35267), .dinb(n35265), .dout(n35268));
  jand g17246(.dina(n35268), .dinb(n34992), .dout(n35269));
  jxor g17247(.dina(n34984), .dinb(n323), .dout(n35270));
  jnot g17248(.din(n35270), .dout(n35271));
  jor  g17249(.dina(n35271), .dinb(n35269), .dout(n35272));
  jand g17250(.dina(n35272), .dinb(n34986), .dout(n35273));
  jxor g17251(.dina(n34978), .dinb(n324), .dout(n35274));
  jnot g17252(.din(n35274), .dout(n35275));
  jor  g17253(.dina(n35275), .dinb(n35273), .dout(n35276));
  jand g17254(.dina(n35276), .dinb(n34980), .dout(n35277));
  jxor g17255(.dina(n34972), .dinb(n325), .dout(n35278));
  jnot g17256(.din(n35278), .dout(n35279));
  jor  g17257(.dina(n35279), .dinb(n35277), .dout(n35280));
  jand g17258(.dina(n35280), .dinb(n34974), .dout(n35281));
  jxor g17259(.dina(n34966), .dinb(n439), .dout(n35282));
  jnot g17260(.din(n35282), .dout(n35283));
  jor  g17261(.dina(n35283), .dinb(n35281), .dout(n35284));
  jand g17262(.dina(n35284), .dinb(n34968), .dout(n35285));
  jxor g17263(.dina(n34960), .dinb(n440), .dout(n35286));
  jnot g17264(.din(n35286), .dout(n35287));
  jor  g17265(.dina(n35287), .dinb(n35285), .dout(n35288));
  jand g17266(.dina(n35288), .dinb(n34962), .dout(n35289));
  jxor g17267(.dina(n34954), .dinb(n435), .dout(n35290));
  jnot g17268(.din(n35290), .dout(n35291));
  jor  g17269(.dina(n35291), .dinb(n35289), .dout(n35292));
  jand g17270(.dina(n35292), .dinb(n34956), .dout(n35293));
  jxor g17271(.dina(n34948), .dinb(n436), .dout(n35294));
  jnot g17272(.din(n35294), .dout(n35295));
  jor  g17273(.dina(n35295), .dinb(n35293), .dout(n35296));
  jand g17274(.dina(n35296), .dinb(n34950), .dout(n35297));
  jxor g17275(.dina(n34942), .dinb(n432), .dout(n35298));
  jnot g17276(.din(n35298), .dout(n35299));
  jor  g17277(.dina(n35299), .dinb(n35297), .dout(n35300));
  jand g17278(.dina(n35300), .dinb(n34944), .dout(n35301));
  jxor g17279(.dina(n34936), .dinb(n433), .dout(n35302));
  jnot g17280(.din(n35302), .dout(n35303));
  jor  g17281(.dina(n35303), .dinb(n35301), .dout(n35304));
  jand g17282(.dina(n35304), .dinb(n34938), .dout(n35305));
  jxor g17283(.dina(n34930), .dinb(n421), .dout(n35306));
  jnot g17284(.din(n35306), .dout(n35307));
  jor  g17285(.dina(n35307), .dinb(n35305), .dout(n35308));
  jand g17286(.dina(n35308), .dinb(n34932), .dout(n35309));
  jxor g17287(.dina(n34924), .dinb(n422), .dout(n35310));
  jnot g17288(.din(n35310), .dout(n35311));
  jor  g17289(.dina(n35311), .dinb(n35309), .dout(n35312));
  jand g17290(.dina(n35312), .dinb(n34926), .dout(n35313));
  jxor g17291(.dina(n34918), .dinb(n416), .dout(n35314));
  jnot g17292(.din(n35314), .dout(n35315));
  jor  g17293(.dina(n35315), .dinb(n35313), .dout(n35316));
  jand g17294(.dina(n35316), .dinb(n34920), .dout(n35317));
  jxor g17295(.dina(n34912), .dinb(n417), .dout(n35318));
  jnot g17296(.din(n35318), .dout(n35319));
  jor  g17297(.dina(n35319), .dinb(n35317), .dout(n35320));
  jand g17298(.dina(n35320), .dinb(n34914), .dout(n35321));
  jxor g17299(.dina(n34906), .dinb(n2547), .dout(n35322));
  jnot g17300(.din(n35322), .dout(n35323));
  jor  g17301(.dina(n35323), .dinb(n35321), .dout(n35324));
  jand g17302(.dina(n35324), .dinb(n34908), .dout(n35325));
  jxor g17303(.dina(n34900), .dinb(n2714), .dout(n35326));
  jnot g17304(.din(n35326), .dout(n35327));
  jor  g17305(.dina(n35327), .dinb(n35325), .dout(n35328));
  jand g17306(.dina(n35328), .dinb(n34902), .dout(n35329));
  jxor g17307(.dina(n34894), .dinb(n405), .dout(n35330));
  jnot g17308(.din(n35330), .dout(n35331));
  jor  g17309(.dina(n35331), .dinb(n35329), .dout(n35332));
  jand g17310(.dina(n35332), .dinb(n34896), .dout(n35333));
  jxor g17311(.dina(n34888), .dinb(n406), .dout(n35334));
  jnot g17312(.din(n35334), .dout(n35335));
  jor  g17313(.dina(n35335), .dinb(n35333), .dout(n35336));
  jand g17314(.dina(n35336), .dinb(n34890), .dout(n35337));
  jxor g17315(.dina(n34882), .dinb(n412), .dout(n35338));
  jnot g17316(.din(n35338), .dout(n35339));
  jor  g17317(.dina(n35339), .dinb(n35337), .dout(n35340));
  jand g17318(.dina(n35340), .dinb(n34884), .dout(n35341));
  jxor g17319(.dina(n34876), .dinb(n413), .dout(n35342));
  jnot g17320(.din(n35342), .dout(n35343));
  jor  g17321(.dina(n35343), .dinb(n35341), .dout(n35344));
  jand g17322(.dina(n35344), .dinb(n34878), .dout(n35345));
  jxor g17323(.dina(n34870), .dinb(n409), .dout(n35346));
  jnot g17324(.din(n35346), .dout(n35347));
  jor  g17325(.dina(n35347), .dinb(n35345), .dout(n35348));
  jand g17326(.dina(n35348), .dinb(n34872), .dout(n35349));
  jxor g17327(.dina(n34864), .dinb(n410), .dout(n35350));
  jnot g17328(.din(n35350), .dout(n35351));
  jor  g17329(.dina(n35351), .dinb(n35349), .dout(n35352));
  jand g17330(.dina(n35352), .dinb(n34866), .dout(n35353));
  jxor g17331(.dina(n34858), .dinb(n426), .dout(n35354));
  jnot g17332(.din(n35354), .dout(n35355));
  jor  g17333(.dina(n35355), .dinb(n35353), .dout(n35356));
  jand g17334(.dina(n35356), .dinb(n34860), .dout(n35357));
  jxor g17335(.dina(n34852), .dinb(n427), .dout(n35358));
  jnot g17336(.din(n35358), .dout(n35359));
  jor  g17337(.dina(n35359), .dinb(n35357), .dout(n35360));
  jand g17338(.dina(n35360), .dinb(n34854), .dout(n35361));
  jxor g17339(.dina(n34846), .dinb(n424), .dout(n35362));
  jnot g17340(.din(n35362), .dout(n35363));
  jor  g17341(.dina(n35363), .dinb(n35361), .dout(n35364));
  jand g17342(.dina(n35364), .dinb(n34848), .dout(n35365));
  jxor g17343(.dina(n34840), .dinb(n300), .dout(n35366));
  jnot g17344(.din(n35366), .dout(n35367));
  jor  g17345(.dina(n35367), .dinb(n35365), .dout(n35368));
  jand g17346(.dina(n35368), .dinb(n34842), .dout(n35369));
  jxor g17347(.dina(n34834), .dinb(n297), .dout(n35370));
  jnot g17348(.din(n35370), .dout(n35371));
  jor  g17349(.dina(n35371), .dinb(n35369), .dout(n35372));
  jand g17350(.dina(n35372), .dinb(n34836), .dout(n35373));
  jxor g17351(.dina(n34828), .dinb(n298), .dout(n35374));
  jnot g17352(.din(n35374), .dout(n35375));
  jor  g17353(.dina(n35375), .dinb(n35373), .dout(n35376));
  jand g17354(.dina(n35376), .dinb(n34830), .dout(n35377));
  jxor g17355(.dina(n34822), .dinb(n301), .dout(n35378));
  jnot g17356(.din(n35378), .dout(n35379));
  jor  g17357(.dina(n35379), .dinb(n35377), .dout(n35380));
  jand g17358(.dina(n35380), .dinb(n34824), .dout(n35381));
  jxor g17359(.dina(n34816), .dinb(n293), .dout(n35382));
  jnot g17360(.din(n35382), .dout(n35383));
  jor  g17361(.dina(n35383), .dinb(n35381), .dout(n35384));
  jand g17362(.dina(n35384), .dinb(n34818), .dout(n35385));
  jxor g17363(.dina(n34810), .dinb(n294), .dout(n35386));
  jnot g17364(.din(n35386), .dout(n35387));
  jor  g17365(.dina(n35387), .dinb(n35385), .dout(n35388));
  jand g17366(.dina(n35388), .dinb(n34812), .dout(n35389));
  jxor g17367(.dina(n34804), .dinb(n290), .dout(n35390));
  jnot g17368(.din(n35390), .dout(n35391));
  jor  g17369(.dina(n35391), .dinb(n35389), .dout(n35392));
  jand g17370(.dina(n35392), .dinb(n34806), .dout(n35393));
  jxor g17371(.dina(n34798), .dinb(n291), .dout(n35394));
  jnot g17372(.din(n35394), .dout(n35395));
  jor  g17373(.dina(n35395), .dinb(n35393), .dout(n35396));
  jand g17374(.dina(n35396), .dinb(n34800), .dout(n35397));
  jxor g17375(.dina(n34792), .dinb(n284), .dout(n35398));
  jnot g17376(.din(n35398), .dout(n35399));
  jor  g17377(.dina(n35399), .dinb(n35397), .dout(n35400));
  jand g17378(.dina(n35400), .dinb(n34794), .dout(n35401));
  jxor g17379(.dina(n34786), .dinb(n285), .dout(n35402));
  jnot g17380(.din(n35402), .dout(n35403));
  jor  g17381(.dina(n35403), .dinb(n35401), .dout(n35404));
  jand g17382(.dina(n35404), .dinb(n34788), .dout(n35405));
  jxor g17383(.dina(n34780), .dinb(n281), .dout(n35406));
  jnot g17384(.din(n35406), .dout(n35407));
  jor  g17385(.dina(n35407), .dinb(n35405), .dout(n35408));
  jand g17386(.dina(n35408), .dinb(n34782), .dout(n35409));
  jxor g17387(.dina(n34774), .dinb(n282), .dout(n35410));
  jnot g17388(.din(n35410), .dout(n35411));
  jor  g17389(.dina(n35411), .dinb(n35409), .dout(n35412));
  jand g17390(.dina(n35412), .dinb(n34776), .dout(n35413));
  jxor g17391(.dina(n34768), .dinb(n397), .dout(n35414));
  jnot g17392(.din(n35414), .dout(n35415));
  jor  g17393(.dina(n35415), .dinb(n35413), .dout(n35416));
  jand g17394(.dina(n35416), .dinb(n34770), .dout(n35417));
  jxor g17395(.dina(n34762), .dinb(n513), .dout(n35418));
  jnot g17396(.din(n35418), .dout(n35419));
  jor  g17397(.dina(n35419), .dinb(n35417), .dout(n35420));
  jand g17398(.dina(n35420), .dinb(n34764), .dout(n35421));
  jxor g17399(.dina(n34756), .dinb(n514), .dout(n35422));
  jnot g17400(.din(n35422), .dout(n35423));
  jor  g17401(.dina(n35423), .dinb(n35421), .dout(n35424));
  jand g17402(.dina(n35424), .dinb(n34758), .dout(n35425));
  jxor g17403(.dina(n34750), .dinb(n510), .dout(n35426));
  jnot g17404(.din(n35426), .dout(n35427));
  jor  g17405(.dina(n35427), .dinb(n35425), .dout(n35428));
  jand g17406(.dina(n35428), .dinb(n34752), .dout(n35429));
  jxor g17407(.dina(n34744), .dinb(n396), .dout(n35430));
  jnot g17408(.din(n35430), .dout(n35431));
  jor  g17409(.dina(n35431), .dinb(n35429), .dout(n35432));
  jand g17410(.dina(n35432), .dinb(n34746), .dout(n35433));
  jxor g17411(.dina(n34738), .dinb(n383), .dout(n35434));
  jnot g17412(.din(n35434), .dout(n35435));
  jor  g17413(.dina(n35435), .dinb(n35433), .dout(n35436));
  jand g17414(.dina(n35436), .dinb(n34740), .dout(n35437));
  jxor g17415(.dina(n34732), .dinb(n12211), .dout(n35438));
  jnot g17416(.din(n35438), .dout(n35439));
  jor  g17417(.dina(n35439), .dinb(n35437), .dout(n35440));
  jand g17418(.dina(n35440), .dinb(n34734), .dout(n35441));
  jxor g17419(.dina(n34726), .dinb(n12214), .dout(n35442));
  jnot g17420(.din(n35442), .dout(n35443));
  jor  g17421(.dina(n35443), .dinb(n35441), .dout(n35444));
  jand g17422(.dina(n35444), .dinb(n34728), .dout(n35445));
  jxor g17423(.dina(n34721), .dinb(b52 ), .dout(n35446));
  jor  g17424(.dina(n35446), .dinb(n13060), .dout(n35447));
  jor  g17425(.dina(n35447), .dinb(n35445), .dout(n35448));
  jand g17426(.dina(n35448), .dinb(n34722), .dout(n35449));
  jxor g17427(.dina(n35242), .dinb(b1 ), .dout(n35450));
  jand g17428(.dina(n35450), .dinb(n12906), .dout(n35451));
  jor  g17429(.dina(n35451), .dinb(n35238), .dout(n35452));
  jand g17430(.dina(n35246), .dinb(n35452), .dout(n35453));
  jor  g17431(.dina(n35453), .dinb(n35026), .dout(n35454));
  jand g17432(.dina(n35250), .dinb(n35454), .dout(n35455));
  jor  g17433(.dina(n35455), .dinb(n35018), .dout(n35456));
  jand g17434(.dina(n35254), .dinb(n35456), .dout(n35457));
  jor  g17435(.dina(n35457), .dinb(n35009), .dout(n35458));
  jand g17436(.dina(n35258), .dinb(n35458), .dout(n35459));
  jor  g17437(.dina(n35459), .dinb(n35003), .dout(n35460));
  jand g17438(.dina(n35262), .dinb(n35460), .dout(n35461));
  jor  g17439(.dina(n35461), .dinb(n34997), .dout(n35462));
  jand g17440(.dina(n35266), .dinb(n35462), .dout(n35463));
  jor  g17441(.dina(n35463), .dinb(n34991), .dout(n35464));
  jand g17442(.dina(n35270), .dinb(n35464), .dout(n35465));
  jor  g17443(.dina(n35465), .dinb(n34985), .dout(n35466));
  jand g17444(.dina(n35274), .dinb(n35466), .dout(n35467));
  jor  g17445(.dina(n35467), .dinb(n34979), .dout(n35468));
  jand g17446(.dina(n35278), .dinb(n35468), .dout(n35469));
  jor  g17447(.dina(n35469), .dinb(n34973), .dout(n35470));
  jand g17448(.dina(n35282), .dinb(n35470), .dout(n35471));
  jor  g17449(.dina(n35471), .dinb(n34967), .dout(n35472));
  jand g17450(.dina(n35286), .dinb(n35472), .dout(n35473));
  jor  g17451(.dina(n35473), .dinb(n34961), .dout(n35474));
  jand g17452(.dina(n35290), .dinb(n35474), .dout(n35475));
  jor  g17453(.dina(n35475), .dinb(n34955), .dout(n35476));
  jand g17454(.dina(n35294), .dinb(n35476), .dout(n35477));
  jor  g17455(.dina(n35477), .dinb(n34949), .dout(n35478));
  jand g17456(.dina(n35298), .dinb(n35478), .dout(n35479));
  jor  g17457(.dina(n35479), .dinb(n34943), .dout(n35480));
  jand g17458(.dina(n35302), .dinb(n35480), .dout(n35481));
  jor  g17459(.dina(n35481), .dinb(n34937), .dout(n35482));
  jand g17460(.dina(n35306), .dinb(n35482), .dout(n35483));
  jor  g17461(.dina(n35483), .dinb(n34931), .dout(n35484));
  jand g17462(.dina(n35310), .dinb(n35484), .dout(n35485));
  jor  g17463(.dina(n35485), .dinb(n34925), .dout(n35486));
  jand g17464(.dina(n35314), .dinb(n35486), .dout(n35487));
  jor  g17465(.dina(n35487), .dinb(n34919), .dout(n35488));
  jand g17466(.dina(n35318), .dinb(n35488), .dout(n35489));
  jor  g17467(.dina(n35489), .dinb(n34913), .dout(n35490));
  jand g17468(.dina(n35322), .dinb(n35490), .dout(n35491));
  jor  g17469(.dina(n35491), .dinb(n34907), .dout(n35492));
  jand g17470(.dina(n35326), .dinb(n35492), .dout(n35493));
  jor  g17471(.dina(n35493), .dinb(n34901), .dout(n35494));
  jand g17472(.dina(n35330), .dinb(n35494), .dout(n35495));
  jor  g17473(.dina(n35495), .dinb(n34895), .dout(n35496));
  jand g17474(.dina(n35334), .dinb(n35496), .dout(n35497));
  jor  g17475(.dina(n35497), .dinb(n34889), .dout(n35498));
  jand g17476(.dina(n35338), .dinb(n35498), .dout(n35499));
  jor  g17477(.dina(n35499), .dinb(n34883), .dout(n35500));
  jand g17478(.dina(n35342), .dinb(n35500), .dout(n35501));
  jor  g17479(.dina(n35501), .dinb(n34877), .dout(n35502));
  jand g17480(.dina(n35346), .dinb(n35502), .dout(n35503));
  jor  g17481(.dina(n35503), .dinb(n34871), .dout(n35504));
  jand g17482(.dina(n35350), .dinb(n35504), .dout(n35505));
  jor  g17483(.dina(n35505), .dinb(n34865), .dout(n35506));
  jand g17484(.dina(n35354), .dinb(n35506), .dout(n35507));
  jor  g17485(.dina(n35507), .dinb(n34859), .dout(n35508));
  jand g17486(.dina(n35358), .dinb(n35508), .dout(n35509));
  jor  g17487(.dina(n35509), .dinb(n34853), .dout(n35510));
  jand g17488(.dina(n35362), .dinb(n35510), .dout(n35511));
  jor  g17489(.dina(n35511), .dinb(n34847), .dout(n35512));
  jand g17490(.dina(n35366), .dinb(n35512), .dout(n35513));
  jor  g17491(.dina(n35513), .dinb(n34841), .dout(n35514));
  jand g17492(.dina(n35370), .dinb(n35514), .dout(n35515));
  jor  g17493(.dina(n35515), .dinb(n34835), .dout(n35516));
  jand g17494(.dina(n35374), .dinb(n35516), .dout(n35517));
  jor  g17495(.dina(n35517), .dinb(n34829), .dout(n35518));
  jand g17496(.dina(n35378), .dinb(n35518), .dout(n35519));
  jor  g17497(.dina(n35519), .dinb(n34823), .dout(n35520));
  jand g17498(.dina(n35382), .dinb(n35520), .dout(n35521));
  jor  g17499(.dina(n35521), .dinb(n34817), .dout(n35522));
  jand g17500(.dina(n35386), .dinb(n35522), .dout(n35523));
  jor  g17501(.dina(n35523), .dinb(n34811), .dout(n35524));
  jand g17502(.dina(n35390), .dinb(n35524), .dout(n35525));
  jor  g17503(.dina(n35525), .dinb(n34805), .dout(n35526));
  jand g17504(.dina(n35394), .dinb(n35526), .dout(n35527));
  jor  g17505(.dina(n35527), .dinb(n34799), .dout(n35528));
  jand g17506(.dina(n35398), .dinb(n35528), .dout(n35529));
  jor  g17507(.dina(n35529), .dinb(n34793), .dout(n35530));
  jand g17508(.dina(n35402), .dinb(n35530), .dout(n35531));
  jor  g17509(.dina(n35531), .dinb(n34787), .dout(n35532));
  jand g17510(.dina(n35406), .dinb(n35532), .dout(n35533));
  jor  g17511(.dina(n35533), .dinb(n34781), .dout(n35534));
  jand g17512(.dina(n35410), .dinb(n35534), .dout(n35535));
  jor  g17513(.dina(n35535), .dinb(n34775), .dout(n35536));
  jand g17514(.dina(n35414), .dinb(n35536), .dout(n35537));
  jor  g17515(.dina(n35537), .dinb(n34769), .dout(n35538));
  jand g17516(.dina(n35418), .dinb(n35538), .dout(n35539));
  jor  g17517(.dina(n35539), .dinb(n34763), .dout(n35540));
  jand g17518(.dina(n35422), .dinb(n35540), .dout(n35541));
  jor  g17519(.dina(n35541), .dinb(n34757), .dout(n35542));
  jand g17520(.dina(n35426), .dinb(n35542), .dout(n35543));
  jor  g17521(.dina(n35543), .dinb(n34751), .dout(n35544));
  jand g17522(.dina(n35430), .dinb(n35544), .dout(n35545));
  jor  g17523(.dina(n35545), .dinb(n34745), .dout(n35546));
  jand g17524(.dina(n35434), .dinb(n35546), .dout(n35547));
  jor  g17525(.dina(n35547), .dinb(n34739), .dout(n35548));
  jand g17526(.dina(n35438), .dinb(n35548), .dout(n35549));
  jor  g17527(.dina(n35549), .dinb(n34733), .dout(n35550));
  jand g17528(.dina(n35442), .dinb(n35550), .dout(n35551));
  jor  g17529(.dina(n35551), .dinb(n34727), .dout(n35552));
  jnot g17530(.din(n35447), .dout(n35553));
  jand g17531(.dina(n35553), .dinb(n35552), .dout(n35554));
  jand g17532(.dina(n34721), .dinb(n583), .dout(n35555));
  jor  g17533(.dina(n35555), .dinb(n35554), .dout(n35556));
  jxor g17534(.dina(n35446), .dinb(n35552), .dout(n35557));
  jand g17535(.dina(n35557), .dinb(n35556), .dout(n35558));
  jor  g17536(.dina(n35558), .dinb(n35449), .dout(n35559));
  jnot g17537(.din(n35559), .dout(n35560));
  jnot g17538(.din(n35555), .dout(n35561));
  jand g17539(.dina(n35561), .dinb(n35448), .dout(n35562));
  jand g17540(.dina(n35562), .dinb(n34726), .dout(n35563));
  jxor g17541(.dina(n35442), .dinb(n35550), .dout(n35564));
  jand g17542(.dina(n35564), .dinb(n35556), .dout(n35565));
  jor  g17543(.dina(n35565), .dinb(n35563), .dout(n35566));
  jand g17544(.dina(n35566), .dinb(n384), .dout(n35567));
  jand g17545(.dina(n35562), .dinb(n34732), .dout(n35568));
  jxor g17546(.dina(n35438), .dinb(n35548), .dout(n35569));
  jand g17547(.dina(n35569), .dinb(n35556), .dout(n35570));
  jor  g17548(.dina(n35570), .dinb(n35568), .dout(n35571));
  jand g17549(.dina(n35571), .dinb(n12214), .dout(n35572));
  jand g17550(.dina(n35562), .dinb(n34738), .dout(n35573));
  jxor g17551(.dina(n35434), .dinb(n35546), .dout(n35574));
  jand g17552(.dina(n35574), .dinb(n35556), .dout(n35575));
  jor  g17553(.dina(n35575), .dinb(n35573), .dout(n35576));
  jand g17554(.dina(n35576), .dinb(n12211), .dout(n35577));
  jand g17555(.dina(n35562), .dinb(n34744), .dout(n35578));
  jxor g17556(.dina(n35430), .dinb(n35544), .dout(n35579));
  jand g17557(.dina(n35579), .dinb(n35556), .dout(n35580));
  jor  g17558(.dina(n35580), .dinb(n35578), .dout(n35581));
  jand g17559(.dina(n35581), .dinb(n383), .dout(n35582));
  jand g17560(.dina(n35562), .dinb(n34750), .dout(n35583));
  jxor g17561(.dina(n35426), .dinb(n35542), .dout(n35584));
  jand g17562(.dina(n35584), .dinb(n35556), .dout(n35585));
  jor  g17563(.dina(n35585), .dinb(n35583), .dout(n35586));
  jand g17564(.dina(n35586), .dinb(n396), .dout(n35587));
  jand g17565(.dina(n35562), .dinb(n34756), .dout(n35588));
  jxor g17566(.dina(n35422), .dinb(n35540), .dout(n35589));
  jand g17567(.dina(n35589), .dinb(n35556), .dout(n35590));
  jor  g17568(.dina(n35590), .dinb(n35588), .dout(n35591));
  jand g17569(.dina(n35591), .dinb(n510), .dout(n35592));
  jand g17570(.dina(n35562), .dinb(n34762), .dout(n35593));
  jxor g17571(.dina(n35418), .dinb(n35538), .dout(n35594));
  jand g17572(.dina(n35594), .dinb(n35556), .dout(n35595));
  jor  g17573(.dina(n35595), .dinb(n35593), .dout(n35596));
  jand g17574(.dina(n35596), .dinb(n514), .dout(n35597));
  jand g17575(.dina(n35562), .dinb(n34768), .dout(n35598));
  jxor g17576(.dina(n35414), .dinb(n35536), .dout(n35599));
  jand g17577(.dina(n35599), .dinb(n35556), .dout(n35600));
  jor  g17578(.dina(n35600), .dinb(n35598), .dout(n35601));
  jand g17579(.dina(n35601), .dinb(n513), .dout(n35602));
  jand g17580(.dina(n35562), .dinb(n34774), .dout(n35603));
  jxor g17581(.dina(n35410), .dinb(n35534), .dout(n35604));
  jand g17582(.dina(n35604), .dinb(n35556), .dout(n35605));
  jor  g17583(.dina(n35605), .dinb(n35603), .dout(n35606));
  jand g17584(.dina(n35606), .dinb(n397), .dout(n35607));
  jand g17585(.dina(n35562), .dinb(n34780), .dout(n35608));
  jxor g17586(.dina(n35406), .dinb(n35532), .dout(n35609));
  jand g17587(.dina(n35609), .dinb(n35556), .dout(n35610));
  jor  g17588(.dina(n35610), .dinb(n35608), .dout(n35611));
  jand g17589(.dina(n35611), .dinb(n282), .dout(n35612));
  jand g17590(.dina(n35562), .dinb(n34786), .dout(n35613));
  jxor g17591(.dina(n35402), .dinb(n35530), .dout(n35614));
  jand g17592(.dina(n35614), .dinb(n35556), .dout(n35615));
  jor  g17593(.dina(n35615), .dinb(n35613), .dout(n35616));
  jand g17594(.dina(n35616), .dinb(n281), .dout(n35617));
  jand g17595(.dina(n35562), .dinb(n34792), .dout(n35618));
  jxor g17596(.dina(n35398), .dinb(n35528), .dout(n35619));
  jand g17597(.dina(n35619), .dinb(n35556), .dout(n35620));
  jor  g17598(.dina(n35620), .dinb(n35618), .dout(n35621));
  jand g17599(.dina(n35621), .dinb(n285), .dout(n35622));
  jand g17600(.dina(n35562), .dinb(n34798), .dout(n35623));
  jxor g17601(.dina(n35394), .dinb(n35526), .dout(n35624));
  jand g17602(.dina(n35624), .dinb(n35556), .dout(n35625));
  jor  g17603(.dina(n35625), .dinb(n35623), .dout(n35626));
  jand g17604(.dina(n35626), .dinb(n284), .dout(n35627));
  jand g17605(.dina(n35562), .dinb(n34804), .dout(n35628));
  jxor g17606(.dina(n35390), .dinb(n35524), .dout(n35629));
  jand g17607(.dina(n35629), .dinb(n35556), .dout(n35630));
  jor  g17608(.dina(n35630), .dinb(n35628), .dout(n35631));
  jand g17609(.dina(n35631), .dinb(n291), .dout(n35632));
  jand g17610(.dina(n35562), .dinb(n34810), .dout(n35633));
  jxor g17611(.dina(n35386), .dinb(n35522), .dout(n35634));
  jand g17612(.dina(n35634), .dinb(n35556), .dout(n35635));
  jor  g17613(.dina(n35635), .dinb(n35633), .dout(n35636));
  jand g17614(.dina(n35636), .dinb(n290), .dout(n35637));
  jand g17615(.dina(n35562), .dinb(n34816), .dout(n35638));
  jxor g17616(.dina(n35382), .dinb(n35520), .dout(n35639));
  jand g17617(.dina(n35639), .dinb(n35556), .dout(n35640));
  jor  g17618(.dina(n35640), .dinb(n35638), .dout(n35641));
  jand g17619(.dina(n35641), .dinb(n294), .dout(n35642));
  jand g17620(.dina(n35562), .dinb(n34822), .dout(n35643));
  jxor g17621(.dina(n35378), .dinb(n35518), .dout(n35644));
  jand g17622(.dina(n35644), .dinb(n35556), .dout(n35645));
  jor  g17623(.dina(n35645), .dinb(n35643), .dout(n35646));
  jand g17624(.dina(n35646), .dinb(n293), .dout(n35647));
  jand g17625(.dina(n35562), .dinb(n34828), .dout(n35648));
  jxor g17626(.dina(n35374), .dinb(n35516), .dout(n35649));
  jand g17627(.dina(n35649), .dinb(n35556), .dout(n35650));
  jor  g17628(.dina(n35650), .dinb(n35648), .dout(n35651));
  jand g17629(.dina(n35651), .dinb(n301), .dout(n35652));
  jand g17630(.dina(n35562), .dinb(n34834), .dout(n35653));
  jxor g17631(.dina(n35370), .dinb(n35514), .dout(n35654));
  jand g17632(.dina(n35654), .dinb(n35556), .dout(n35655));
  jor  g17633(.dina(n35655), .dinb(n35653), .dout(n35656));
  jand g17634(.dina(n35656), .dinb(n298), .dout(n35657));
  jand g17635(.dina(n35562), .dinb(n34840), .dout(n35658));
  jxor g17636(.dina(n35366), .dinb(n35512), .dout(n35659));
  jand g17637(.dina(n35659), .dinb(n35556), .dout(n35660));
  jor  g17638(.dina(n35660), .dinb(n35658), .dout(n35661));
  jand g17639(.dina(n35661), .dinb(n297), .dout(n35662));
  jand g17640(.dina(n35562), .dinb(n34846), .dout(n35663));
  jxor g17641(.dina(n35362), .dinb(n35510), .dout(n35664));
  jand g17642(.dina(n35664), .dinb(n35556), .dout(n35665));
  jor  g17643(.dina(n35665), .dinb(n35663), .dout(n35666));
  jand g17644(.dina(n35666), .dinb(n300), .dout(n35667));
  jand g17645(.dina(n35562), .dinb(n34852), .dout(n35668));
  jxor g17646(.dina(n35358), .dinb(n35508), .dout(n35669));
  jand g17647(.dina(n35669), .dinb(n35556), .dout(n35670));
  jor  g17648(.dina(n35670), .dinb(n35668), .dout(n35671));
  jand g17649(.dina(n35671), .dinb(n424), .dout(n35672));
  jand g17650(.dina(n35562), .dinb(n34858), .dout(n35673));
  jxor g17651(.dina(n35354), .dinb(n35506), .dout(n35674));
  jand g17652(.dina(n35674), .dinb(n35556), .dout(n35675));
  jor  g17653(.dina(n35675), .dinb(n35673), .dout(n35676));
  jand g17654(.dina(n35676), .dinb(n427), .dout(n35677));
  jand g17655(.dina(n35562), .dinb(n34864), .dout(n35678));
  jxor g17656(.dina(n35350), .dinb(n35504), .dout(n35679));
  jand g17657(.dina(n35679), .dinb(n35556), .dout(n35680));
  jor  g17658(.dina(n35680), .dinb(n35678), .dout(n35681));
  jand g17659(.dina(n35681), .dinb(n426), .dout(n35682));
  jand g17660(.dina(n35562), .dinb(n34870), .dout(n35683));
  jxor g17661(.dina(n35346), .dinb(n35502), .dout(n35684));
  jand g17662(.dina(n35684), .dinb(n35556), .dout(n35685));
  jor  g17663(.dina(n35685), .dinb(n35683), .dout(n35686));
  jand g17664(.dina(n35686), .dinb(n410), .dout(n35687));
  jand g17665(.dina(n35562), .dinb(n34876), .dout(n35688));
  jxor g17666(.dina(n35342), .dinb(n35500), .dout(n35689));
  jand g17667(.dina(n35689), .dinb(n35556), .dout(n35690));
  jor  g17668(.dina(n35690), .dinb(n35688), .dout(n35691));
  jand g17669(.dina(n35691), .dinb(n409), .dout(n35692));
  jand g17670(.dina(n35562), .dinb(n34882), .dout(n35693));
  jxor g17671(.dina(n35338), .dinb(n35498), .dout(n35694));
  jand g17672(.dina(n35694), .dinb(n35556), .dout(n35695));
  jor  g17673(.dina(n35695), .dinb(n35693), .dout(n35696));
  jand g17674(.dina(n35696), .dinb(n413), .dout(n35697));
  jand g17675(.dina(n35562), .dinb(n34888), .dout(n35698));
  jxor g17676(.dina(n35334), .dinb(n35496), .dout(n35699));
  jand g17677(.dina(n35699), .dinb(n35556), .dout(n35700));
  jor  g17678(.dina(n35700), .dinb(n35698), .dout(n35701));
  jand g17679(.dina(n35701), .dinb(n412), .dout(n35702));
  jand g17680(.dina(n35562), .dinb(n34894), .dout(n35703));
  jxor g17681(.dina(n35330), .dinb(n35494), .dout(n35704));
  jand g17682(.dina(n35704), .dinb(n35556), .dout(n35705));
  jor  g17683(.dina(n35705), .dinb(n35703), .dout(n35706));
  jand g17684(.dina(n35706), .dinb(n406), .dout(n35707));
  jand g17685(.dina(n35562), .dinb(n34900), .dout(n35708));
  jxor g17686(.dina(n35326), .dinb(n35492), .dout(n35709));
  jand g17687(.dina(n35709), .dinb(n35556), .dout(n35710));
  jor  g17688(.dina(n35710), .dinb(n35708), .dout(n35711));
  jand g17689(.dina(n35711), .dinb(n405), .dout(n35712));
  jand g17690(.dina(n35562), .dinb(n34906), .dout(n35713));
  jxor g17691(.dina(n35322), .dinb(n35490), .dout(n35714));
  jand g17692(.dina(n35714), .dinb(n35556), .dout(n35715));
  jor  g17693(.dina(n35715), .dinb(n35713), .dout(n35716));
  jand g17694(.dina(n35716), .dinb(n2714), .dout(n35717));
  jand g17695(.dina(n35562), .dinb(n34912), .dout(n35718));
  jxor g17696(.dina(n35318), .dinb(n35488), .dout(n35719));
  jand g17697(.dina(n35719), .dinb(n35556), .dout(n35720));
  jor  g17698(.dina(n35720), .dinb(n35718), .dout(n35721));
  jand g17699(.dina(n35721), .dinb(n2547), .dout(n35722));
  jand g17700(.dina(n35562), .dinb(n34918), .dout(n35723));
  jxor g17701(.dina(n35314), .dinb(n35486), .dout(n35724));
  jand g17702(.dina(n35724), .dinb(n35556), .dout(n35725));
  jor  g17703(.dina(n35725), .dinb(n35723), .dout(n35726));
  jand g17704(.dina(n35726), .dinb(n417), .dout(n35727));
  jand g17705(.dina(n35562), .dinb(n34924), .dout(n35728));
  jxor g17706(.dina(n35310), .dinb(n35484), .dout(n35729));
  jand g17707(.dina(n35729), .dinb(n35556), .dout(n35730));
  jor  g17708(.dina(n35730), .dinb(n35728), .dout(n35731));
  jand g17709(.dina(n35731), .dinb(n416), .dout(n35732));
  jand g17710(.dina(n35562), .dinb(n34930), .dout(n35733));
  jxor g17711(.dina(n35306), .dinb(n35482), .dout(n35734));
  jand g17712(.dina(n35734), .dinb(n35556), .dout(n35735));
  jor  g17713(.dina(n35735), .dinb(n35733), .dout(n35736));
  jand g17714(.dina(n35736), .dinb(n422), .dout(n35737));
  jand g17715(.dina(n35562), .dinb(n34936), .dout(n35738));
  jxor g17716(.dina(n35302), .dinb(n35480), .dout(n35739));
  jand g17717(.dina(n35739), .dinb(n35556), .dout(n35740));
  jor  g17718(.dina(n35740), .dinb(n35738), .dout(n35741));
  jand g17719(.dina(n35741), .dinb(n421), .dout(n35742));
  jand g17720(.dina(n35562), .dinb(n34942), .dout(n35743));
  jxor g17721(.dina(n35298), .dinb(n35478), .dout(n35744));
  jand g17722(.dina(n35744), .dinb(n35556), .dout(n35745));
  jor  g17723(.dina(n35745), .dinb(n35743), .dout(n35746));
  jand g17724(.dina(n35746), .dinb(n433), .dout(n35747));
  jand g17725(.dina(n35562), .dinb(n34948), .dout(n35748));
  jxor g17726(.dina(n35294), .dinb(n35476), .dout(n35749));
  jand g17727(.dina(n35749), .dinb(n35556), .dout(n35750));
  jor  g17728(.dina(n35750), .dinb(n35748), .dout(n35751));
  jand g17729(.dina(n35751), .dinb(n432), .dout(n35752));
  jand g17730(.dina(n35562), .dinb(n34954), .dout(n35753));
  jxor g17731(.dina(n35290), .dinb(n35474), .dout(n35754));
  jand g17732(.dina(n35754), .dinb(n35556), .dout(n35755));
  jor  g17733(.dina(n35755), .dinb(n35753), .dout(n35756));
  jand g17734(.dina(n35756), .dinb(n436), .dout(n35757));
  jand g17735(.dina(n35562), .dinb(n34960), .dout(n35758));
  jxor g17736(.dina(n35286), .dinb(n35472), .dout(n35759));
  jand g17737(.dina(n35759), .dinb(n35556), .dout(n35760));
  jor  g17738(.dina(n35760), .dinb(n35758), .dout(n35761));
  jand g17739(.dina(n35761), .dinb(n435), .dout(n35762));
  jand g17740(.dina(n35562), .dinb(n34966), .dout(n35763));
  jxor g17741(.dina(n35282), .dinb(n35470), .dout(n35764));
  jand g17742(.dina(n35764), .dinb(n35556), .dout(n35765));
  jor  g17743(.dina(n35765), .dinb(n35763), .dout(n35766));
  jand g17744(.dina(n35766), .dinb(n440), .dout(n35767));
  jand g17745(.dina(n35562), .dinb(n34972), .dout(n35768));
  jxor g17746(.dina(n35278), .dinb(n35468), .dout(n35769));
  jand g17747(.dina(n35769), .dinb(n35556), .dout(n35770));
  jor  g17748(.dina(n35770), .dinb(n35768), .dout(n35771));
  jand g17749(.dina(n35771), .dinb(n439), .dout(n35772));
  jand g17750(.dina(n35562), .dinb(n34978), .dout(n35773));
  jxor g17751(.dina(n35274), .dinb(n35466), .dout(n35774));
  jand g17752(.dina(n35774), .dinb(n35556), .dout(n35775));
  jor  g17753(.dina(n35775), .dinb(n35773), .dout(n35776));
  jand g17754(.dina(n35776), .dinb(n325), .dout(n35777));
  jand g17755(.dina(n35562), .dinb(n34984), .dout(n35778));
  jxor g17756(.dina(n35270), .dinb(n35464), .dout(n35779));
  jand g17757(.dina(n35779), .dinb(n35556), .dout(n35780));
  jor  g17758(.dina(n35780), .dinb(n35778), .dout(n35781));
  jand g17759(.dina(n35781), .dinb(n324), .dout(n35782));
  jand g17760(.dina(n35562), .dinb(n34990), .dout(n35783));
  jxor g17761(.dina(n35266), .dinb(n35462), .dout(n35784));
  jand g17762(.dina(n35784), .dinb(n35556), .dout(n35785));
  jor  g17763(.dina(n35785), .dinb(n35783), .dout(n35786));
  jand g17764(.dina(n35786), .dinb(n323), .dout(n35787));
  jand g17765(.dina(n35562), .dinb(n34996), .dout(n35788));
  jxor g17766(.dina(n35262), .dinb(n35460), .dout(n35789));
  jand g17767(.dina(n35789), .dinb(n35556), .dout(n35790));
  jor  g17768(.dina(n35790), .dinb(n35788), .dout(n35791));
  jand g17769(.dina(n35791), .dinb(n335), .dout(n35792));
  jand g17770(.dina(n35562), .dinb(n35002), .dout(n35793));
  jxor g17771(.dina(n35258), .dinb(n35458), .dout(n35794));
  jand g17772(.dina(n35794), .dinb(n35556), .dout(n35795));
  jor  g17773(.dina(n35795), .dinb(n35793), .dout(n35796));
  jand g17774(.dina(n35796), .dinb(n334), .dout(n35797));
  jand g17775(.dina(n35562), .dinb(n35008), .dout(n35798));
  jxor g17776(.dina(n35254), .dinb(n35456), .dout(n35799));
  jand g17777(.dina(n35799), .dinb(n35556), .dout(n35800));
  jor  g17778(.dina(n35800), .dinb(n35798), .dout(n35801));
  jand g17779(.dina(n35801), .dinb(n338), .dout(n35802));
  jand g17780(.dina(n35562), .dinb(n35017), .dout(n35803));
  jxor g17781(.dina(n35250), .dinb(n35454), .dout(n35804));
  jand g17782(.dina(n35804), .dinb(n35556), .dout(n35805));
  jor  g17783(.dina(n35805), .dinb(n35803), .dout(n35806));
  jand g17784(.dina(n35806), .dinb(n337), .dout(n35807));
  jand g17785(.dina(n35562), .dinb(n35025), .dout(n35808));
  jxor g17786(.dina(n35246), .dinb(n35452), .dout(n35809));
  jand g17787(.dina(n35809), .dinb(n35556), .dout(n35810));
  jor  g17788(.dina(n35810), .dinb(n35808), .dout(n35811));
  jand g17789(.dina(n35811), .dinb(n344), .dout(n35812));
  jand g17790(.dina(n35562), .dinb(n35237), .dout(n35813));
  jxor g17791(.dina(n35450), .dinb(n12906), .dout(n35814));
  jand g17792(.dina(n35814), .dinb(n35556), .dout(n35815));
  jor  g17793(.dina(n35815), .dinb(n35813), .dout(n35816));
  jand g17794(.dina(n35816), .dinb(n348), .dout(n35817));
  jor  g17795(.dina(n35562), .dinb(n18364), .dout(n35818));
  jand g17796(.dina(n35818), .dinb(a11 ), .dout(n35819));
  jor  g17797(.dina(n35562), .dinb(n12906), .dout(n35820));
  jnot g17798(.din(n35820), .dout(n35821));
  jor  g17799(.dina(n35821), .dinb(n35819), .dout(n35822));
  jand g17800(.dina(n35822), .dinb(n258), .dout(n35823));
  jand g17801(.dina(n35556), .dinb(b0 ), .dout(n35824));
  jor  g17802(.dina(n35824), .dinb(n12904), .dout(n35825));
  jand g17803(.dina(n35820), .dinb(n35825), .dout(n35826));
  jxor g17804(.dina(n35826), .dinb(b1 ), .dout(n35827));
  jand g17805(.dina(n35827), .dinb(n13344), .dout(n35828));
  jor  g17806(.dina(n35828), .dinb(n35823), .dout(n35829));
  jxor g17807(.dina(n35816), .dinb(n348), .dout(n35830));
  jand g17808(.dina(n35830), .dinb(n35829), .dout(n35831));
  jor  g17809(.dina(n35831), .dinb(n35817), .dout(n35832));
  jxor g17810(.dina(n35811), .dinb(n344), .dout(n35833));
  jand g17811(.dina(n35833), .dinb(n35832), .dout(n35834));
  jor  g17812(.dina(n35834), .dinb(n35812), .dout(n35835));
  jxor g17813(.dina(n35806), .dinb(n337), .dout(n35836));
  jand g17814(.dina(n35836), .dinb(n35835), .dout(n35837));
  jor  g17815(.dina(n35837), .dinb(n35807), .dout(n35838));
  jxor g17816(.dina(n35801), .dinb(n338), .dout(n35839));
  jand g17817(.dina(n35839), .dinb(n35838), .dout(n35840));
  jor  g17818(.dina(n35840), .dinb(n35802), .dout(n35841));
  jxor g17819(.dina(n35796), .dinb(n334), .dout(n35842));
  jand g17820(.dina(n35842), .dinb(n35841), .dout(n35843));
  jor  g17821(.dina(n35843), .dinb(n35797), .dout(n35844));
  jxor g17822(.dina(n35791), .dinb(n335), .dout(n35845));
  jand g17823(.dina(n35845), .dinb(n35844), .dout(n35846));
  jor  g17824(.dina(n35846), .dinb(n35792), .dout(n35847));
  jxor g17825(.dina(n35786), .dinb(n323), .dout(n35848));
  jand g17826(.dina(n35848), .dinb(n35847), .dout(n35849));
  jor  g17827(.dina(n35849), .dinb(n35787), .dout(n35850));
  jxor g17828(.dina(n35781), .dinb(n324), .dout(n35851));
  jand g17829(.dina(n35851), .dinb(n35850), .dout(n35852));
  jor  g17830(.dina(n35852), .dinb(n35782), .dout(n35853));
  jxor g17831(.dina(n35776), .dinb(n325), .dout(n35854));
  jand g17832(.dina(n35854), .dinb(n35853), .dout(n35855));
  jor  g17833(.dina(n35855), .dinb(n35777), .dout(n35856));
  jxor g17834(.dina(n35771), .dinb(n439), .dout(n35857));
  jand g17835(.dina(n35857), .dinb(n35856), .dout(n35858));
  jor  g17836(.dina(n35858), .dinb(n35772), .dout(n35859));
  jxor g17837(.dina(n35766), .dinb(n440), .dout(n35860));
  jand g17838(.dina(n35860), .dinb(n35859), .dout(n35861));
  jor  g17839(.dina(n35861), .dinb(n35767), .dout(n35862));
  jxor g17840(.dina(n35761), .dinb(n435), .dout(n35863));
  jand g17841(.dina(n35863), .dinb(n35862), .dout(n35864));
  jor  g17842(.dina(n35864), .dinb(n35762), .dout(n35865));
  jxor g17843(.dina(n35756), .dinb(n436), .dout(n35866));
  jand g17844(.dina(n35866), .dinb(n35865), .dout(n35867));
  jor  g17845(.dina(n35867), .dinb(n35757), .dout(n35868));
  jxor g17846(.dina(n35751), .dinb(n432), .dout(n35869));
  jand g17847(.dina(n35869), .dinb(n35868), .dout(n35870));
  jor  g17848(.dina(n35870), .dinb(n35752), .dout(n35871));
  jxor g17849(.dina(n35746), .dinb(n433), .dout(n35872));
  jand g17850(.dina(n35872), .dinb(n35871), .dout(n35873));
  jor  g17851(.dina(n35873), .dinb(n35747), .dout(n35874));
  jxor g17852(.dina(n35741), .dinb(n421), .dout(n35875));
  jand g17853(.dina(n35875), .dinb(n35874), .dout(n35876));
  jor  g17854(.dina(n35876), .dinb(n35742), .dout(n35877));
  jxor g17855(.dina(n35736), .dinb(n422), .dout(n35878));
  jand g17856(.dina(n35878), .dinb(n35877), .dout(n35879));
  jor  g17857(.dina(n35879), .dinb(n35737), .dout(n35880));
  jxor g17858(.dina(n35731), .dinb(n416), .dout(n35881));
  jand g17859(.dina(n35881), .dinb(n35880), .dout(n35882));
  jor  g17860(.dina(n35882), .dinb(n35732), .dout(n35883));
  jxor g17861(.dina(n35726), .dinb(n417), .dout(n35884));
  jand g17862(.dina(n35884), .dinb(n35883), .dout(n35885));
  jor  g17863(.dina(n35885), .dinb(n35727), .dout(n35886));
  jxor g17864(.dina(n35721), .dinb(n2547), .dout(n35887));
  jand g17865(.dina(n35887), .dinb(n35886), .dout(n35888));
  jor  g17866(.dina(n35888), .dinb(n35722), .dout(n35889));
  jxor g17867(.dina(n35716), .dinb(n2714), .dout(n35890));
  jand g17868(.dina(n35890), .dinb(n35889), .dout(n35891));
  jor  g17869(.dina(n35891), .dinb(n35717), .dout(n35892));
  jxor g17870(.dina(n35711), .dinb(n405), .dout(n35893));
  jand g17871(.dina(n35893), .dinb(n35892), .dout(n35894));
  jor  g17872(.dina(n35894), .dinb(n35712), .dout(n35895));
  jxor g17873(.dina(n35706), .dinb(n406), .dout(n35896));
  jand g17874(.dina(n35896), .dinb(n35895), .dout(n35897));
  jor  g17875(.dina(n35897), .dinb(n35707), .dout(n35898));
  jxor g17876(.dina(n35701), .dinb(n412), .dout(n35899));
  jand g17877(.dina(n35899), .dinb(n35898), .dout(n35900));
  jor  g17878(.dina(n35900), .dinb(n35702), .dout(n35901));
  jxor g17879(.dina(n35696), .dinb(n413), .dout(n35902));
  jand g17880(.dina(n35902), .dinb(n35901), .dout(n35903));
  jor  g17881(.dina(n35903), .dinb(n35697), .dout(n35904));
  jxor g17882(.dina(n35691), .dinb(n409), .dout(n35905));
  jand g17883(.dina(n35905), .dinb(n35904), .dout(n35906));
  jor  g17884(.dina(n35906), .dinb(n35692), .dout(n35907));
  jxor g17885(.dina(n35686), .dinb(n410), .dout(n35908));
  jand g17886(.dina(n35908), .dinb(n35907), .dout(n35909));
  jor  g17887(.dina(n35909), .dinb(n35687), .dout(n35910));
  jxor g17888(.dina(n35681), .dinb(n426), .dout(n35911));
  jand g17889(.dina(n35911), .dinb(n35910), .dout(n35912));
  jor  g17890(.dina(n35912), .dinb(n35682), .dout(n35913));
  jxor g17891(.dina(n35676), .dinb(n427), .dout(n35914));
  jand g17892(.dina(n35914), .dinb(n35913), .dout(n35915));
  jor  g17893(.dina(n35915), .dinb(n35677), .dout(n35916));
  jxor g17894(.dina(n35671), .dinb(n424), .dout(n35917));
  jand g17895(.dina(n35917), .dinb(n35916), .dout(n35918));
  jor  g17896(.dina(n35918), .dinb(n35672), .dout(n35919));
  jxor g17897(.dina(n35666), .dinb(n300), .dout(n35920));
  jand g17898(.dina(n35920), .dinb(n35919), .dout(n35921));
  jor  g17899(.dina(n35921), .dinb(n35667), .dout(n35922));
  jxor g17900(.dina(n35661), .dinb(n297), .dout(n35923));
  jand g17901(.dina(n35923), .dinb(n35922), .dout(n35924));
  jor  g17902(.dina(n35924), .dinb(n35662), .dout(n35925));
  jxor g17903(.dina(n35656), .dinb(n298), .dout(n35926));
  jand g17904(.dina(n35926), .dinb(n35925), .dout(n35927));
  jor  g17905(.dina(n35927), .dinb(n35657), .dout(n35928));
  jxor g17906(.dina(n35651), .dinb(n301), .dout(n35929));
  jand g17907(.dina(n35929), .dinb(n35928), .dout(n35930));
  jor  g17908(.dina(n35930), .dinb(n35652), .dout(n35931));
  jxor g17909(.dina(n35646), .dinb(n293), .dout(n35932));
  jand g17910(.dina(n35932), .dinb(n35931), .dout(n35933));
  jor  g17911(.dina(n35933), .dinb(n35647), .dout(n35934));
  jxor g17912(.dina(n35641), .dinb(n294), .dout(n35935));
  jand g17913(.dina(n35935), .dinb(n35934), .dout(n35936));
  jor  g17914(.dina(n35936), .dinb(n35642), .dout(n35937));
  jxor g17915(.dina(n35636), .dinb(n290), .dout(n35938));
  jand g17916(.dina(n35938), .dinb(n35937), .dout(n35939));
  jor  g17917(.dina(n35939), .dinb(n35637), .dout(n35940));
  jxor g17918(.dina(n35631), .dinb(n291), .dout(n35941));
  jand g17919(.dina(n35941), .dinb(n35940), .dout(n35942));
  jor  g17920(.dina(n35942), .dinb(n35632), .dout(n35943));
  jxor g17921(.dina(n35626), .dinb(n284), .dout(n35944));
  jand g17922(.dina(n35944), .dinb(n35943), .dout(n35945));
  jor  g17923(.dina(n35945), .dinb(n35627), .dout(n35946));
  jxor g17924(.dina(n35621), .dinb(n285), .dout(n35947));
  jand g17925(.dina(n35947), .dinb(n35946), .dout(n35948));
  jor  g17926(.dina(n35948), .dinb(n35622), .dout(n35949));
  jxor g17927(.dina(n35616), .dinb(n281), .dout(n35950));
  jand g17928(.dina(n35950), .dinb(n35949), .dout(n35951));
  jor  g17929(.dina(n35951), .dinb(n35617), .dout(n35952));
  jxor g17930(.dina(n35611), .dinb(n282), .dout(n35953));
  jand g17931(.dina(n35953), .dinb(n35952), .dout(n35954));
  jor  g17932(.dina(n35954), .dinb(n35612), .dout(n35955));
  jxor g17933(.dina(n35606), .dinb(n397), .dout(n35956));
  jand g17934(.dina(n35956), .dinb(n35955), .dout(n35957));
  jor  g17935(.dina(n35957), .dinb(n35607), .dout(n35958));
  jxor g17936(.dina(n35601), .dinb(n513), .dout(n35959));
  jand g17937(.dina(n35959), .dinb(n35958), .dout(n35960));
  jor  g17938(.dina(n35960), .dinb(n35602), .dout(n35961));
  jxor g17939(.dina(n35596), .dinb(n514), .dout(n35962));
  jand g17940(.dina(n35962), .dinb(n35961), .dout(n35963));
  jor  g17941(.dina(n35963), .dinb(n35597), .dout(n35964));
  jxor g17942(.dina(n35591), .dinb(n510), .dout(n35965));
  jand g17943(.dina(n35965), .dinb(n35964), .dout(n35966));
  jor  g17944(.dina(n35966), .dinb(n35592), .dout(n35967));
  jxor g17945(.dina(n35586), .dinb(n396), .dout(n35968));
  jand g17946(.dina(n35968), .dinb(n35967), .dout(n35969));
  jor  g17947(.dina(n35969), .dinb(n35587), .dout(n35970));
  jxor g17948(.dina(n35581), .dinb(n383), .dout(n35971));
  jand g17949(.dina(n35971), .dinb(n35970), .dout(n35972));
  jor  g17950(.dina(n35972), .dinb(n35582), .dout(n35973));
  jxor g17951(.dina(n35576), .dinb(n12211), .dout(n35974));
  jand g17952(.dina(n35974), .dinb(n35973), .dout(n35975));
  jor  g17953(.dina(n35975), .dinb(n35577), .dout(n35976));
  jxor g17954(.dina(n35571), .dinb(n12214), .dout(n35977));
  jand g17955(.dina(n35977), .dinb(n35976), .dout(n35978));
  jor  g17956(.dina(n35978), .dinb(n35572), .dout(n35979));
  jxor g17957(.dina(n35566), .dinb(n384), .dout(n35980));
  jand g17958(.dina(n35980), .dinb(n35979), .dout(n35981));
  jor  g17959(.dina(n35981), .dinb(n35567), .dout(n35982));
  jand g17960(.dina(n35982), .dinb(n374), .dout(n35983));
  jnot g17961(.din(n13503), .dout(n35984));
  jnot g17962(.din(n35567), .dout(n35985));
  jnot g17963(.din(n35572), .dout(n35986));
  jnot g17964(.din(n35577), .dout(n35987));
  jnot g17965(.din(n35582), .dout(n35988));
  jnot g17966(.din(n35587), .dout(n35989));
  jnot g17967(.din(n35592), .dout(n35990));
  jnot g17968(.din(n35597), .dout(n35991));
  jnot g17969(.din(n35602), .dout(n35992));
  jnot g17970(.din(n35607), .dout(n35993));
  jnot g17971(.din(n35612), .dout(n35994));
  jnot g17972(.din(n35617), .dout(n35995));
  jnot g17973(.din(n35622), .dout(n35996));
  jnot g17974(.din(n35627), .dout(n35997));
  jnot g17975(.din(n35632), .dout(n35998));
  jnot g17976(.din(n35637), .dout(n35999));
  jnot g17977(.din(n35642), .dout(n36000));
  jnot g17978(.din(n35647), .dout(n36001));
  jnot g17979(.din(n35652), .dout(n36002));
  jnot g17980(.din(n35657), .dout(n36003));
  jnot g17981(.din(n35662), .dout(n36004));
  jnot g17982(.din(n35667), .dout(n36005));
  jnot g17983(.din(n35672), .dout(n36006));
  jnot g17984(.din(n35677), .dout(n36007));
  jnot g17985(.din(n35682), .dout(n36008));
  jnot g17986(.din(n35687), .dout(n36009));
  jnot g17987(.din(n35692), .dout(n36010));
  jnot g17988(.din(n35697), .dout(n36011));
  jnot g17989(.din(n35702), .dout(n36012));
  jnot g17990(.din(n35707), .dout(n36013));
  jnot g17991(.din(n35712), .dout(n36014));
  jnot g17992(.din(n35717), .dout(n36015));
  jnot g17993(.din(n35722), .dout(n36016));
  jnot g17994(.din(n35727), .dout(n36017));
  jnot g17995(.din(n35732), .dout(n36018));
  jnot g17996(.din(n35737), .dout(n36019));
  jnot g17997(.din(n35742), .dout(n36020));
  jnot g17998(.din(n35747), .dout(n36021));
  jnot g17999(.din(n35752), .dout(n36022));
  jnot g18000(.din(n35757), .dout(n36023));
  jnot g18001(.din(n35762), .dout(n36024));
  jnot g18002(.din(n35767), .dout(n36025));
  jnot g18003(.din(n35772), .dout(n36026));
  jnot g18004(.din(n35777), .dout(n36027));
  jnot g18005(.din(n35782), .dout(n36028));
  jnot g18006(.din(n35787), .dout(n36029));
  jnot g18007(.din(n35792), .dout(n36030));
  jnot g18008(.din(n35797), .dout(n36031));
  jnot g18009(.din(n35802), .dout(n36032));
  jnot g18010(.din(n35807), .dout(n36033));
  jnot g18011(.din(n35812), .dout(n36034));
  jnot g18012(.din(n35817), .dout(n36035));
  jnot g18013(.din(n35823), .dout(n36036));
  jxor g18014(.dina(n35826), .dinb(n258), .dout(n36037));
  jor  g18015(.dina(n36037), .dinb(n13343), .dout(n36038));
  jand g18016(.dina(n36038), .dinb(n36036), .dout(n36039));
  jnot g18017(.din(n35830), .dout(n36040));
  jor  g18018(.dina(n36040), .dinb(n36039), .dout(n36041));
  jand g18019(.dina(n36041), .dinb(n36035), .dout(n36042));
  jnot g18020(.din(n35833), .dout(n36043));
  jor  g18021(.dina(n36043), .dinb(n36042), .dout(n36044));
  jand g18022(.dina(n36044), .dinb(n36034), .dout(n36045));
  jnot g18023(.din(n35836), .dout(n36046));
  jor  g18024(.dina(n36046), .dinb(n36045), .dout(n36047));
  jand g18025(.dina(n36047), .dinb(n36033), .dout(n36048));
  jnot g18026(.din(n35839), .dout(n36049));
  jor  g18027(.dina(n36049), .dinb(n36048), .dout(n36050));
  jand g18028(.dina(n36050), .dinb(n36032), .dout(n36051));
  jnot g18029(.din(n35842), .dout(n36052));
  jor  g18030(.dina(n36052), .dinb(n36051), .dout(n36053));
  jand g18031(.dina(n36053), .dinb(n36031), .dout(n36054));
  jnot g18032(.din(n35845), .dout(n36055));
  jor  g18033(.dina(n36055), .dinb(n36054), .dout(n36056));
  jand g18034(.dina(n36056), .dinb(n36030), .dout(n36057));
  jnot g18035(.din(n35848), .dout(n36058));
  jor  g18036(.dina(n36058), .dinb(n36057), .dout(n36059));
  jand g18037(.dina(n36059), .dinb(n36029), .dout(n36060));
  jnot g18038(.din(n35851), .dout(n36061));
  jor  g18039(.dina(n36061), .dinb(n36060), .dout(n36062));
  jand g18040(.dina(n36062), .dinb(n36028), .dout(n36063));
  jnot g18041(.din(n35854), .dout(n36064));
  jor  g18042(.dina(n36064), .dinb(n36063), .dout(n36065));
  jand g18043(.dina(n36065), .dinb(n36027), .dout(n36066));
  jnot g18044(.din(n35857), .dout(n36067));
  jor  g18045(.dina(n36067), .dinb(n36066), .dout(n36068));
  jand g18046(.dina(n36068), .dinb(n36026), .dout(n36069));
  jnot g18047(.din(n35860), .dout(n36070));
  jor  g18048(.dina(n36070), .dinb(n36069), .dout(n36071));
  jand g18049(.dina(n36071), .dinb(n36025), .dout(n36072));
  jnot g18050(.din(n35863), .dout(n36073));
  jor  g18051(.dina(n36073), .dinb(n36072), .dout(n36074));
  jand g18052(.dina(n36074), .dinb(n36024), .dout(n36075));
  jnot g18053(.din(n35866), .dout(n36076));
  jor  g18054(.dina(n36076), .dinb(n36075), .dout(n36077));
  jand g18055(.dina(n36077), .dinb(n36023), .dout(n36078));
  jnot g18056(.din(n35869), .dout(n36079));
  jor  g18057(.dina(n36079), .dinb(n36078), .dout(n36080));
  jand g18058(.dina(n36080), .dinb(n36022), .dout(n36081));
  jnot g18059(.din(n35872), .dout(n36082));
  jor  g18060(.dina(n36082), .dinb(n36081), .dout(n36083));
  jand g18061(.dina(n36083), .dinb(n36021), .dout(n36084));
  jnot g18062(.din(n35875), .dout(n36085));
  jor  g18063(.dina(n36085), .dinb(n36084), .dout(n36086));
  jand g18064(.dina(n36086), .dinb(n36020), .dout(n36087));
  jnot g18065(.din(n35878), .dout(n36088));
  jor  g18066(.dina(n36088), .dinb(n36087), .dout(n36089));
  jand g18067(.dina(n36089), .dinb(n36019), .dout(n36090));
  jnot g18068(.din(n35881), .dout(n36091));
  jor  g18069(.dina(n36091), .dinb(n36090), .dout(n36092));
  jand g18070(.dina(n36092), .dinb(n36018), .dout(n36093));
  jnot g18071(.din(n35884), .dout(n36094));
  jor  g18072(.dina(n36094), .dinb(n36093), .dout(n36095));
  jand g18073(.dina(n36095), .dinb(n36017), .dout(n36096));
  jnot g18074(.din(n35887), .dout(n36097));
  jor  g18075(.dina(n36097), .dinb(n36096), .dout(n36098));
  jand g18076(.dina(n36098), .dinb(n36016), .dout(n36099));
  jnot g18077(.din(n35890), .dout(n36100));
  jor  g18078(.dina(n36100), .dinb(n36099), .dout(n36101));
  jand g18079(.dina(n36101), .dinb(n36015), .dout(n36102));
  jnot g18080(.din(n35893), .dout(n36103));
  jor  g18081(.dina(n36103), .dinb(n36102), .dout(n36104));
  jand g18082(.dina(n36104), .dinb(n36014), .dout(n36105));
  jnot g18083(.din(n35896), .dout(n36106));
  jor  g18084(.dina(n36106), .dinb(n36105), .dout(n36107));
  jand g18085(.dina(n36107), .dinb(n36013), .dout(n36108));
  jnot g18086(.din(n35899), .dout(n36109));
  jor  g18087(.dina(n36109), .dinb(n36108), .dout(n36110));
  jand g18088(.dina(n36110), .dinb(n36012), .dout(n36111));
  jnot g18089(.din(n35902), .dout(n36112));
  jor  g18090(.dina(n36112), .dinb(n36111), .dout(n36113));
  jand g18091(.dina(n36113), .dinb(n36011), .dout(n36114));
  jnot g18092(.din(n35905), .dout(n36115));
  jor  g18093(.dina(n36115), .dinb(n36114), .dout(n36116));
  jand g18094(.dina(n36116), .dinb(n36010), .dout(n36117));
  jnot g18095(.din(n35908), .dout(n36118));
  jor  g18096(.dina(n36118), .dinb(n36117), .dout(n36119));
  jand g18097(.dina(n36119), .dinb(n36009), .dout(n36120));
  jnot g18098(.din(n35911), .dout(n36121));
  jor  g18099(.dina(n36121), .dinb(n36120), .dout(n36122));
  jand g18100(.dina(n36122), .dinb(n36008), .dout(n36123));
  jnot g18101(.din(n35914), .dout(n36124));
  jor  g18102(.dina(n36124), .dinb(n36123), .dout(n36125));
  jand g18103(.dina(n36125), .dinb(n36007), .dout(n36126));
  jnot g18104(.din(n35917), .dout(n36127));
  jor  g18105(.dina(n36127), .dinb(n36126), .dout(n36128));
  jand g18106(.dina(n36128), .dinb(n36006), .dout(n36129));
  jnot g18107(.din(n35920), .dout(n36130));
  jor  g18108(.dina(n36130), .dinb(n36129), .dout(n36131));
  jand g18109(.dina(n36131), .dinb(n36005), .dout(n36132));
  jnot g18110(.din(n35923), .dout(n36133));
  jor  g18111(.dina(n36133), .dinb(n36132), .dout(n36134));
  jand g18112(.dina(n36134), .dinb(n36004), .dout(n36135));
  jnot g18113(.din(n35926), .dout(n36136));
  jor  g18114(.dina(n36136), .dinb(n36135), .dout(n36137));
  jand g18115(.dina(n36137), .dinb(n36003), .dout(n36138));
  jnot g18116(.din(n35929), .dout(n36139));
  jor  g18117(.dina(n36139), .dinb(n36138), .dout(n36140));
  jand g18118(.dina(n36140), .dinb(n36002), .dout(n36141));
  jnot g18119(.din(n35932), .dout(n36142));
  jor  g18120(.dina(n36142), .dinb(n36141), .dout(n36143));
  jand g18121(.dina(n36143), .dinb(n36001), .dout(n36144));
  jnot g18122(.din(n35935), .dout(n36145));
  jor  g18123(.dina(n36145), .dinb(n36144), .dout(n36146));
  jand g18124(.dina(n36146), .dinb(n36000), .dout(n36147));
  jnot g18125(.din(n35938), .dout(n36148));
  jor  g18126(.dina(n36148), .dinb(n36147), .dout(n36149));
  jand g18127(.dina(n36149), .dinb(n35999), .dout(n36150));
  jnot g18128(.din(n35941), .dout(n36151));
  jor  g18129(.dina(n36151), .dinb(n36150), .dout(n36152));
  jand g18130(.dina(n36152), .dinb(n35998), .dout(n36153));
  jnot g18131(.din(n35944), .dout(n36154));
  jor  g18132(.dina(n36154), .dinb(n36153), .dout(n36155));
  jand g18133(.dina(n36155), .dinb(n35997), .dout(n36156));
  jnot g18134(.din(n35947), .dout(n36157));
  jor  g18135(.dina(n36157), .dinb(n36156), .dout(n36158));
  jand g18136(.dina(n36158), .dinb(n35996), .dout(n36159));
  jnot g18137(.din(n35950), .dout(n36160));
  jor  g18138(.dina(n36160), .dinb(n36159), .dout(n36161));
  jand g18139(.dina(n36161), .dinb(n35995), .dout(n36162));
  jnot g18140(.din(n35953), .dout(n36163));
  jor  g18141(.dina(n36163), .dinb(n36162), .dout(n36164));
  jand g18142(.dina(n36164), .dinb(n35994), .dout(n36165));
  jnot g18143(.din(n35956), .dout(n36166));
  jor  g18144(.dina(n36166), .dinb(n36165), .dout(n36167));
  jand g18145(.dina(n36167), .dinb(n35993), .dout(n36168));
  jnot g18146(.din(n35959), .dout(n36169));
  jor  g18147(.dina(n36169), .dinb(n36168), .dout(n36170));
  jand g18148(.dina(n36170), .dinb(n35992), .dout(n36171));
  jnot g18149(.din(n35962), .dout(n36172));
  jor  g18150(.dina(n36172), .dinb(n36171), .dout(n36173));
  jand g18151(.dina(n36173), .dinb(n35991), .dout(n36174));
  jnot g18152(.din(n35965), .dout(n36175));
  jor  g18153(.dina(n36175), .dinb(n36174), .dout(n36176));
  jand g18154(.dina(n36176), .dinb(n35990), .dout(n36177));
  jnot g18155(.din(n35968), .dout(n36178));
  jor  g18156(.dina(n36178), .dinb(n36177), .dout(n36179));
  jand g18157(.dina(n36179), .dinb(n35989), .dout(n36180));
  jnot g18158(.din(n35971), .dout(n36181));
  jor  g18159(.dina(n36181), .dinb(n36180), .dout(n36182));
  jand g18160(.dina(n36182), .dinb(n35988), .dout(n36183));
  jnot g18161(.din(n35974), .dout(n36184));
  jor  g18162(.dina(n36184), .dinb(n36183), .dout(n36185));
  jand g18163(.dina(n36185), .dinb(n35987), .dout(n36186));
  jnot g18164(.din(n35977), .dout(n36187));
  jor  g18165(.dina(n36187), .dinb(n36186), .dout(n36188));
  jand g18166(.dina(n36188), .dinb(n35986), .dout(n36189));
  jnot g18167(.din(n35980), .dout(n36190));
  jor  g18168(.dina(n36190), .dinb(n36189), .dout(n36191));
  jand g18169(.dina(n36191), .dinb(n35985), .dout(n36192));
  jand g18170(.dina(n36192), .dinb(b53 ), .dout(n36193));
  jor  g18171(.dina(n36193), .dinb(n35984), .dout(n36194));
  jor  g18172(.dina(n36194), .dinb(n35983), .dout(n36195));
  jand g18173(.dina(n36195), .dinb(n35560), .dout(n36196));
  jnot g18174(.din(n36196), .dout(n36197));
  jand g18175(.dina(n36197), .dinb(b54 ), .dout(n36198));
  jand g18176(.dina(n36196), .dinb(n376), .dout(n36199));
  jnot g18177(.din(n36199), .dout(n36200));
  jand g18178(.dina(n35560), .dinb(n374), .dout(n36201));
  jnot g18179(.din(n36201), .dout(n36202));
  jand g18180(.dina(n36202), .dinb(n36192), .dout(n36203));
  jand g18181(.dina(n35559), .dinb(b53 ), .dout(n36204));
  jor  g18182(.dina(n36204), .dinb(n35984), .dout(n36205));
  jor  g18183(.dina(n36205), .dinb(n36203), .dout(n36206));
  jand g18184(.dina(n36206), .dinb(n35566), .dout(n36207));
  jor  g18185(.dina(n36201), .dinb(n35982), .dout(n36208));
  jnot g18186(.din(n36205), .dout(n36209));
  jand g18187(.dina(n36209), .dinb(n36208), .dout(n36210));
  jxor g18188(.dina(n35980), .dinb(n35979), .dout(n36211));
  jand g18189(.dina(n36211), .dinb(n36210), .dout(n36212));
  jor  g18190(.dina(n36212), .dinb(n36207), .dout(n36213));
  jand g18191(.dina(n36213), .dinb(n374), .dout(n36214));
  jnot g18192(.din(n36214), .dout(n36215));
  jand g18193(.dina(n36206), .dinb(n35571), .dout(n36216));
  jxor g18194(.dina(n35977), .dinb(n35976), .dout(n36217));
  jand g18195(.dina(n36217), .dinb(n36210), .dout(n36218));
  jor  g18196(.dina(n36218), .dinb(n36216), .dout(n36219));
  jand g18197(.dina(n36219), .dinb(n384), .dout(n36220));
  jnot g18198(.din(n36220), .dout(n36221));
  jand g18199(.dina(n36206), .dinb(n35576), .dout(n36222));
  jxor g18200(.dina(n35974), .dinb(n35973), .dout(n36223));
  jand g18201(.dina(n36223), .dinb(n36210), .dout(n36224));
  jor  g18202(.dina(n36224), .dinb(n36222), .dout(n36225));
  jand g18203(.dina(n36225), .dinb(n12214), .dout(n36226));
  jnot g18204(.din(n36226), .dout(n36227));
  jand g18205(.dina(n36206), .dinb(n35581), .dout(n36228));
  jxor g18206(.dina(n35971), .dinb(n35970), .dout(n36229));
  jand g18207(.dina(n36229), .dinb(n36210), .dout(n36230));
  jor  g18208(.dina(n36230), .dinb(n36228), .dout(n36231));
  jand g18209(.dina(n36231), .dinb(n12211), .dout(n36232));
  jnot g18210(.din(n36232), .dout(n36233));
  jand g18211(.dina(n36206), .dinb(n35586), .dout(n36234));
  jxor g18212(.dina(n35968), .dinb(n35967), .dout(n36235));
  jand g18213(.dina(n36235), .dinb(n36210), .dout(n36236));
  jor  g18214(.dina(n36236), .dinb(n36234), .dout(n36237));
  jand g18215(.dina(n36237), .dinb(n383), .dout(n36238));
  jnot g18216(.din(n36238), .dout(n36239));
  jand g18217(.dina(n36206), .dinb(n35591), .dout(n36240));
  jxor g18218(.dina(n35965), .dinb(n35964), .dout(n36241));
  jand g18219(.dina(n36241), .dinb(n36210), .dout(n36242));
  jor  g18220(.dina(n36242), .dinb(n36240), .dout(n36243));
  jand g18221(.dina(n36243), .dinb(n396), .dout(n36244));
  jnot g18222(.din(n36244), .dout(n36245));
  jand g18223(.dina(n36206), .dinb(n35596), .dout(n36246));
  jxor g18224(.dina(n35962), .dinb(n35961), .dout(n36247));
  jand g18225(.dina(n36247), .dinb(n36210), .dout(n36248));
  jor  g18226(.dina(n36248), .dinb(n36246), .dout(n36249));
  jand g18227(.dina(n36249), .dinb(n510), .dout(n36250));
  jnot g18228(.din(n36250), .dout(n36251));
  jand g18229(.dina(n36206), .dinb(n35601), .dout(n36252));
  jxor g18230(.dina(n35959), .dinb(n35958), .dout(n36253));
  jand g18231(.dina(n36253), .dinb(n36210), .dout(n36254));
  jor  g18232(.dina(n36254), .dinb(n36252), .dout(n36255));
  jand g18233(.dina(n36255), .dinb(n514), .dout(n36256));
  jnot g18234(.din(n36256), .dout(n36257));
  jand g18235(.dina(n36206), .dinb(n35606), .dout(n36258));
  jxor g18236(.dina(n35956), .dinb(n35955), .dout(n36259));
  jand g18237(.dina(n36259), .dinb(n36210), .dout(n36260));
  jor  g18238(.dina(n36260), .dinb(n36258), .dout(n36261));
  jand g18239(.dina(n36261), .dinb(n513), .dout(n36262));
  jnot g18240(.din(n36262), .dout(n36263));
  jand g18241(.dina(n36206), .dinb(n35611), .dout(n36264));
  jxor g18242(.dina(n35953), .dinb(n35952), .dout(n36265));
  jand g18243(.dina(n36265), .dinb(n36210), .dout(n36266));
  jor  g18244(.dina(n36266), .dinb(n36264), .dout(n36267));
  jand g18245(.dina(n36267), .dinb(n397), .dout(n36268));
  jnot g18246(.din(n36268), .dout(n36269));
  jand g18247(.dina(n36206), .dinb(n35616), .dout(n36270));
  jxor g18248(.dina(n35950), .dinb(n35949), .dout(n36271));
  jand g18249(.dina(n36271), .dinb(n36210), .dout(n36272));
  jor  g18250(.dina(n36272), .dinb(n36270), .dout(n36273));
  jand g18251(.dina(n36273), .dinb(n282), .dout(n36274));
  jnot g18252(.din(n36274), .dout(n36275));
  jand g18253(.dina(n36206), .dinb(n35621), .dout(n36276));
  jxor g18254(.dina(n35947), .dinb(n35946), .dout(n36277));
  jand g18255(.dina(n36277), .dinb(n36210), .dout(n36278));
  jor  g18256(.dina(n36278), .dinb(n36276), .dout(n36279));
  jand g18257(.dina(n36279), .dinb(n281), .dout(n36280));
  jnot g18258(.din(n36280), .dout(n36281));
  jand g18259(.dina(n36206), .dinb(n35626), .dout(n36282));
  jxor g18260(.dina(n35944), .dinb(n35943), .dout(n36283));
  jand g18261(.dina(n36283), .dinb(n36210), .dout(n36284));
  jor  g18262(.dina(n36284), .dinb(n36282), .dout(n36285));
  jand g18263(.dina(n36285), .dinb(n285), .dout(n36286));
  jnot g18264(.din(n36286), .dout(n36287));
  jand g18265(.dina(n36206), .dinb(n35631), .dout(n36288));
  jxor g18266(.dina(n35941), .dinb(n35940), .dout(n36289));
  jand g18267(.dina(n36289), .dinb(n36210), .dout(n36290));
  jor  g18268(.dina(n36290), .dinb(n36288), .dout(n36291));
  jand g18269(.dina(n36291), .dinb(n284), .dout(n36292));
  jnot g18270(.din(n36292), .dout(n36293));
  jand g18271(.dina(n36206), .dinb(n35636), .dout(n36294));
  jxor g18272(.dina(n35938), .dinb(n35937), .dout(n36295));
  jand g18273(.dina(n36295), .dinb(n36210), .dout(n36296));
  jor  g18274(.dina(n36296), .dinb(n36294), .dout(n36297));
  jand g18275(.dina(n36297), .dinb(n291), .dout(n36298));
  jnot g18276(.din(n36298), .dout(n36299));
  jand g18277(.dina(n36206), .dinb(n35641), .dout(n36300));
  jxor g18278(.dina(n35935), .dinb(n35934), .dout(n36301));
  jand g18279(.dina(n36301), .dinb(n36210), .dout(n36302));
  jor  g18280(.dina(n36302), .dinb(n36300), .dout(n36303));
  jand g18281(.dina(n36303), .dinb(n290), .dout(n36304));
  jnot g18282(.din(n36304), .dout(n36305));
  jand g18283(.dina(n36206), .dinb(n35646), .dout(n36306));
  jxor g18284(.dina(n35932), .dinb(n35931), .dout(n36307));
  jand g18285(.dina(n36307), .dinb(n36210), .dout(n36308));
  jor  g18286(.dina(n36308), .dinb(n36306), .dout(n36309));
  jand g18287(.dina(n36309), .dinb(n294), .dout(n36310));
  jnot g18288(.din(n36310), .dout(n36311));
  jand g18289(.dina(n36206), .dinb(n35651), .dout(n36312));
  jxor g18290(.dina(n35929), .dinb(n35928), .dout(n36313));
  jand g18291(.dina(n36313), .dinb(n36210), .dout(n36314));
  jor  g18292(.dina(n36314), .dinb(n36312), .dout(n36315));
  jand g18293(.dina(n36315), .dinb(n293), .dout(n36316));
  jnot g18294(.din(n36316), .dout(n36317));
  jand g18295(.dina(n36206), .dinb(n35656), .dout(n36318));
  jxor g18296(.dina(n35926), .dinb(n35925), .dout(n36319));
  jand g18297(.dina(n36319), .dinb(n36210), .dout(n36320));
  jor  g18298(.dina(n36320), .dinb(n36318), .dout(n36321));
  jand g18299(.dina(n36321), .dinb(n301), .dout(n36322));
  jnot g18300(.din(n36322), .dout(n36323));
  jand g18301(.dina(n36206), .dinb(n35661), .dout(n36324));
  jxor g18302(.dina(n35923), .dinb(n35922), .dout(n36325));
  jand g18303(.dina(n36325), .dinb(n36210), .dout(n36326));
  jor  g18304(.dina(n36326), .dinb(n36324), .dout(n36327));
  jand g18305(.dina(n36327), .dinb(n298), .dout(n36328));
  jnot g18306(.din(n36328), .dout(n36329));
  jand g18307(.dina(n36206), .dinb(n35666), .dout(n36330));
  jxor g18308(.dina(n35920), .dinb(n35919), .dout(n36331));
  jand g18309(.dina(n36331), .dinb(n36210), .dout(n36332));
  jor  g18310(.dina(n36332), .dinb(n36330), .dout(n36333));
  jand g18311(.dina(n36333), .dinb(n297), .dout(n36334));
  jnot g18312(.din(n36334), .dout(n36335));
  jand g18313(.dina(n36206), .dinb(n35671), .dout(n36336));
  jxor g18314(.dina(n35917), .dinb(n35916), .dout(n36337));
  jand g18315(.dina(n36337), .dinb(n36210), .dout(n36338));
  jor  g18316(.dina(n36338), .dinb(n36336), .dout(n36339));
  jand g18317(.dina(n36339), .dinb(n300), .dout(n36340));
  jnot g18318(.din(n36340), .dout(n36341));
  jand g18319(.dina(n36206), .dinb(n35676), .dout(n36342));
  jxor g18320(.dina(n35914), .dinb(n35913), .dout(n36343));
  jand g18321(.dina(n36343), .dinb(n36210), .dout(n36344));
  jor  g18322(.dina(n36344), .dinb(n36342), .dout(n36345));
  jand g18323(.dina(n36345), .dinb(n424), .dout(n36346));
  jnot g18324(.din(n36346), .dout(n36347));
  jand g18325(.dina(n36206), .dinb(n35681), .dout(n36348));
  jxor g18326(.dina(n35911), .dinb(n35910), .dout(n36349));
  jand g18327(.dina(n36349), .dinb(n36210), .dout(n36350));
  jor  g18328(.dina(n36350), .dinb(n36348), .dout(n36351));
  jand g18329(.dina(n36351), .dinb(n427), .dout(n36352));
  jnot g18330(.din(n36352), .dout(n36353));
  jand g18331(.dina(n36206), .dinb(n35686), .dout(n36354));
  jxor g18332(.dina(n35908), .dinb(n35907), .dout(n36355));
  jand g18333(.dina(n36355), .dinb(n36210), .dout(n36356));
  jor  g18334(.dina(n36356), .dinb(n36354), .dout(n36357));
  jand g18335(.dina(n36357), .dinb(n426), .dout(n36358));
  jnot g18336(.din(n36358), .dout(n36359));
  jand g18337(.dina(n36206), .dinb(n35691), .dout(n36360));
  jxor g18338(.dina(n35905), .dinb(n35904), .dout(n36361));
  jand g18339(.dina(n36361), .dinb(n36210), .dout(n36362));
  jor  g18340(.dina(n36362), .dinb(n36360), .dout(n36363));
  jand g18341(.dina(n36363), .dinb(n410), .dout(n36364));
  jnot g18342(.din(n36364), .dout(n36365));
  jand g18343(.dina(n36206), .dinb(n35696), .dout(n36366));
  jxor g18344(.dina(n35902), .dinb(n35901), .dout(n36367));
  jand g18345(.dina(n36367), .dinb(n36210), .dout(n36368));
  jor  g18346(.dina(n36368), .dinb(n36366), .dout(n36369));
  jand g18347(.dina(n36369), .dinb(n409), .dout(n36370));
  jnot g18348(.din(n36370), .dout(n36371));
  jand g18349(.dina(n36206), .dinb(n35701), .dout(n36372));
  jxor g18350(.dina(n35899), .dinb(n35898), .dout(n36373));
  jand g18351(.dina(n36373), .dinb(n36210), .dout(n36374));
  jor  g18352(.dina(n36374), .dinb(n36372), .dout(n36375));
  jand g18353(.dina(n36375), .dinb(n413), .dout(n36376));
  jnot g18354(.din(n36376), .dout(n36377));
  jand g18355(.dina(n36206), .dinb(n35706), .dout(n36378));
  jxor g18356(.dina(n35896), .dinb(n35895), .dout(n36379));
  jand g18357(.dina(n36379), .dinb(n36210), .dout(n36380));
  jor  g18358(.dina(n36380), .dinb(n36378), .dout(n36381));
  jand g18359(.dina(n36381), .dinb(n412), .dout(n36382));
  jnot g18360(.din(n36382), .dout(n36383));
  jand g18361(.dina(n36206), .dinb(n35711), .dout(n36384));
  jxor g18362(.dina(n35893), .dinb(n35892), .dout(n36385));
  jand g18363(.dina(n36385), .dinb(n36210), .dout(n36386));
  jor  g18364(.dina(n36386), .dinb(n36384), .dout(n36387));
  jand g18365(.dina(n36387), .dinb(n406), .dout(n36388));
  jnot g18366(.din(n36388), .dout(n36389));
  jand g18367(.dina(n36206), .dinb(n35716), .dout(n36390));
  jxor g18368(.dina(n35890), .dinb(n35889), .dout(n36391));
  jand g18369(.dina(n36391), .dinb(n36210), .dout(n36392));
  jor  g18370(.dina(n36392), .dinb(n36390), .dout(n36393));
  jand g18371(.dina(n36393), .dinb(n405), .dout(n36394));
  jnot g18372(.din(n36394), .dout(n36395));
  jand g18373(.dina(n36206), .dinb(n35721), .dout(n36396));
  jxor g18374(.dina(n35887), .dinb(n35886), .dout(n36397));
  jand g18375(.dina(n36397), .dinb(n36210), .dout(n36398));
  jor  g18376(.dina(n36398), .dinb(n36396), .dout(n36399));
  jand g18377(.dina(n36399), .dinb(n2714), .dout(n36400));
  jnot g18378(.din(n36400), .dout(n36401));
  jand g18379(.dina(n36206), .dinb(n35726), .dout(n36402));
  jxor g18380(.dina(n35884), .dinb(n35883), .dout(n36403));
  jand g18381(.dina(n36403), .dinb(n36210), .dout(n36404));
  jor  g18382(.dina(n36404), .dinb(n36402), .dout(n36405));
  jand g18383(.dina(n36405), .dinb(n2547), .dout(n36406));
  jnot g18384(.din(n36406), .dout(n36407));
  jand g18385(.dina(n36206), .dinb(n35731), .dout(n36408));
  jxor g18386(.dina(n35881), .dinb(n35880), .dout(n36409));
  jand g18387(.dina(n36409), .dinb(n36210), .dout(n36410));
  jor  g18388(.dina(n36410), .dinb(n36408), .dout(n36411));
  jand g18389(.dina(n36411), .dinb(n417), .dout(n36412));
  jnot g18390(.din(n36412), .dout(n36413));
  jand g18391(.dina(n36206), .dinb(n35736), .dout(n36414));
  jxor g18392(.dina(n35878), .dinb(n35877), .dout(n36415));
  jand g18393(.dina(n36415), .dinb(n36210), .dout(n36416));
  jor  g18394(.dina(n36416), .dinb(n36414), .dout(n36417));
  jand g18395(.dina(n36417), .dinb(n416), .dout(n36418));
  jnot g18396(.din(n36418), .dout(n36419));
  jand g18397(.dina(n36206), .dinb(n35741), .dout(n36420));
  jxor g18398(.dina(n35875), .dinb(n35874), .dout(n36421));
  jand g18399(.dina(n36421), .dinb(n36210), .dout(n36422));
  jor  g18400(.dina(n36422), .dinb(n36420), .dout(n36423));
  jand g18401(.dina(n36423), .dinb(n422), .dout(n36424));
  jnot g18402(.din(n36424), .dout(n36425));
  jand g18403(.dina(n36206), .dinb(n35746), .dout(n36426));
  jxor g18404(.dina(n35872), .dinb(n35871), .dout(n36427));
  jand g18405(.dina(n36427), .dinb(n36210), .dout(n36428));
  jor  g18406(.dina(n36428), .dinb(n36426), .dout(n36429));
  jand g18407(.dina(n36429), .dinb(n421), .dout(n36430));
  jnot g18408(.din(n36430), .dout(n36431));
  jand g18409(.dina(n36206), .dinb(n35751), .dout(n36432));
  jxor g18410(.dina(n35869), .dinb(n35868), .dout(n36433));
  jand g18411(.dina(n36433), .dinb(n36210), .dout(n36434));
  jor  g18412(.dina(n36434), .dinb(n36432), .dout(n36435));
  jand g18413(.dina(n36435), .dinb(n433), .dout(n36436));
  jnot g18414(.din(n36436), .dout(n36437));
  jand g18415(.dina(n36206), .dinb(n35756), .dout(n36438));
  jxor g18416(.dina(n35866), .dinb(n35865), .dout(n36439));
  jand g18417(.dina(n36439), .dinb(n36210), .dout(n36440));
  jor  g18418(.dina(n36440), .dinb(n36438), .dout(n36441));
  jand g18419(.dina(n36441), .dinb(n432), .dout(n36442));
  jnot g18420(.din(n36442), .dout(n36443));
  jand g18421(.dina(n36206), .dinb(n35761), .dout(n36444));
  jxor g18422(.dina(n35863), .dinb(n35862), .dout(n36445));
  jand g18423(.dina(n36445), .dinb(n36210), .dout(n36446));
  jor  g18424(.dina(n36446), .dinb(n36444), .dout(n36447));
  jand g18425(.dina(n36447), .dinb(n436), .dout(n36448));
  jnot g18426(.din(n36448), .dout(n36449));
  jand g18427(.dina(n36206), .dinb(n35766), .dout(n36450));
  jxor g18428(.dina(n35860), .dinb(n35859), .dout(n36451));
  jand g18429(.dina(n36451), .dinb(n36210), .dout(n36452));
  jor  g18430(.dina(n36452), .dinb(n36450), .dout(n36453));
  jand g18431(.dina(n36453), .dinb(n435), .dout(n36454));
  jnot g18432(.din(n36454), .dout(n36455));
  jand g18433(.dina(n36206), .dinb(n35771), .dout(n36456));
  jxor g18434(.dina(n35857), .dinb(n35856), .dout(n36457));
  jand g18435(.dina(n36457), .dinb(n36210), .dout(n36458));
  jor  g18436(.dina(n36458), .dinb(n36456), .dout(n36459));
  jand g18437(.dina(n36459), .dinb(n440), .dout(n36460));
  jnot g18438(.din(n36460), .dout(n36461));
  jand g18439(.dina(n36206), .dinb(n35776), .dout(n36462));
  jxor g18440(.dina(n35854), .dinb(n35853), .dout(n36463));
  jand g18441(.dina(n36463), .dinb(n36210), .dout(n36464));
  jor  g18442(.dina(n36464), .dinb(n36462), .dout(n36465));
  jand g18443(.dina(n36465), .dinb(n439), .dout(n36466));
  jnot g18444(.din(n36466), .dout(n36467));
  jand g18445(.dina(n36206), .dinb(n35781), .dout(n36468));
  jxor g18446(.dina(n35851), .dinb(n35850), .dout(n36469));
  jand g18447(.dina(n36469), .dinb(n36210), .dout(n36470));
  jor  g18448(.dina(n36470), .dinb(n36468), .dout(n36471));
  jand g18449(.dina(n36471), .dinb(n325), .dout(n36472));
  jnot g18450(.din(n36472), .dout(n36473));
  jand g18451(.dina(n36206), .dinb(n35786), .dout(n36474));
  jxor g18452(.dina(n35848), .dinb(n35847), .dout(n36475));
  jand g18453(.dina(n36475), .dinb(n36210), .dout(n36476));
  jor  g18454(.dina(n36476), .dinb(n36474), .dout(n36477));
  jand g18455(.dina(n36477), .dinb(n324), .dout(n36478));
  jnot g18456(.din(n36478), .dout(n36479));
  jand g18457(.dina(n36206), .dinb(n35791), .dout(n36480));
  jxor g18458(.dina(n35845), .dinb(n35844), .dout(n36481));
  jand g18459(.dina(n36481), .dinb(n36210), .dout(n36482));
  jor  g18460(.dina(n36482), .dinb(n36480), .dout(n36483));
  jand g18461(.dina(n36483), .dinb(n323), .dout(n36484));
  jnot g18462(.din(n36484), .dout(n36485));
  jand g18463(.dina(n36206), .dinb(n35796), .dout(n36486));
  jxor g18464(.dina(n35842), .dinb(n35841), .dout(n36487));
  jand g18465(.dina(n36487), .dinb(n36210), .dout(n36488));
  jor  g18466(.dina(n36488), .dinb(n36486), .dout(n36489));
  jand g18467(.dina(n36489), .dinb(n335), .dout(n36490));
  jnot g18468(.din(n36490), .dout(n36491));
  jand g18469(.dina(n36206), .dinb(n35801), .dout(n36492));
  jxor g18470(.dina(n35839), .dinb(n35838), .dout(n36493));
  jand g18471(.dina(n36493), .dinb(n36210), .dout(n36494));
  jor  g18472(.dina(n36494), .dinb(n36492), .dout(n36495));
  jand g18473(.dina(n36495), .dinb(n334), .dout(n36496));
  jnot g18474(.din(n36496), .dout(n36497));
  jand g18475(.dina(n36206), .dinb(n35806), .dout(n36498));
  jxor g18476(.dina(n35836), .dinb(n35835), .dout(n36499));
  jand g18477(.dina(n36499), .dinb(n36210), .dout(n36500));
  jor  g18478(.dina(n36500), .dinb(n36498), .dout(n36501));
  jand g18479(.dina(n36501), .dinb(n338), .dout(n36502));
  jnot g18480(.din(n36502), .dout(n36503));
  jand g18481(.dina(n36206), .dinb(n35811), .dout(n36504));
  jxor g18482(.dina(n35833), .dinb(n35832), .dout(n36505));
  jand g18483(.dina(n36505), .dinb(n36210), .dout(n36506));
  jor  g18484(.dina(n36506), .dinb(n36504), .dout(n36507));
  jand g18485(.dina(n36507), .dinb(n337), .dout(n36508));
  jnot g18486(.din(n36508), .dout(n36509));
  jand g18487(.dina(n36206), .dinb(n35816), .dout(n36510));
  jxor g18488(.dina(n35830), .dinb(n35829), .dout(n36511));
  jand g18489(.dina(n36511), .dinb(n36210), .dout(n36512));
  jor  g18490(.dina(n36512), .dinb(n36510), .dout(n36513));
  jand g18491(.dina(n36513), .dinb(n344), .dout(n36514));
  jnot g18492(.din(n36514), .dout(n36515));
  jand g18493(.dina(n36206), .dinb(n35822), .dout(n36516));
  jxor g18494(.dina(n35827), .dinb(n13344), .dout(n36517));
  jand g18495(.dina(n36517), .dinb(n36210), .dout(n36518));
  jor  g18496(.dina(n36518), .dinb(n36516), .dout(n36519));
  jand g18497(.dina(n36519), .dinb(n348), .dout(n36520));
  jnot g18498(.din(n36520), .dout(n36521));
  jor  g18499(.dina(n36206), .dinb(n18364), .dout(n36522));
  jand g18500(.dina(n36522), .dinb(a10 ), .dout(n36523));
  jor  g18501(.dina(n36206), .dinb(n13344), .dout(n36524));
  jnot g18502(.din(n36524), .dout(n36525));
  jor  g18503(.dina(n36525), .dinb(n36523), .dout(n36526));
  jand g18504(.dina(n36526), .dinb(n258), .dout(n36527));
  jnot g18505(.din(n36527), .dout(n36528));
  jand g18506(.dina(n36210), .dinb(b0 ), .dout(n36529));
  jor  g18507(.dina(n36529), .dinb(n13342), .dout(n36530));
  jand g18508(.dina(n36524), .dinb(n36530), .dout(n36531));
  jxor g18509(.dina(n36531), .dinb(n258), .dout(n36532));
  jor  g18510(.dina(n36532), .dinb(n13838), .dout(n36533));
  jand g18511(.dina(n36533), .dinb(n36528), .dout(n36534));
  jxor g18512(.dina(n36519), .dinb(n348), .dout(n36535));
  jnot g18513(.din(n36535), .dout(n36536));
  jor  g18514(.dina(n36536), .dinb(n36534), .dout(n36537));
  jand g18515(.dina(n36537), .dinb(n36521), .dout(n36538));
  jxor g18516(.dina(n36513), .dinb(n344), .dout(n36539));
  jnot g18517(.din(n36539), .dout(n36540));
  jor  g18518(.dina(n36540), .dinb(n36538), .dout(n36541));
  jand g18519(.dina(n36541), .dinb(n36515), .dout(n36542));
  jxor g18520(.dina(n36507), .dinb(n337), .dout(n36543));
  jnot g18521(.din(n36543), .dout(n36544));
  jor  g18522(.dina(n36544), .dinb(n36542), .dout(n36545));
  jand g18523(.dina(n36545), .dinb(n36509), .dout(n36546));
  jxor g18524(.dina(n36501), .dinb(n338), .dout(n36547));
  jnot g18525(.din(n36547), .dout(n36548));
  jor  g18526(.dina(n36548), .dinb(n36546), .dout(n36549));
  jand g18527(.dina(n36549), .dinb(n36503), .dout(n36550));
  jxor g18528(.dina(n36495), .dinb(n334), .dout(n36551));
  jnot g18529(.din(n36551), .dout(n36552));
  jor  g18530(.dina(n36552), .dinb(n36550), .dout(n36553));
  jand g18531(.dina(n36553), .dinb(n36497), .dout(n36554));
  jxor g18532(.dina(n36489), .dinb(n335), .dout(n36555));
  jnot g18533(.din(n36555), .dout(n36556));
  jor  g18534(.dina(n36556), .dinb(n36554), .dout(n36557));
  jand g18535(.dina(n36557), .dinb(n36491), .dout(n36558));
  jxor g18536(.dina(n36483), .dinb(n323), .dout(n36559));
  jnot g18537(.din(n36559), .dout(n36560));
  jor  g18538(.dina(n36560), .dinb(n36558), .dout(n36561));
  jand g18539(.dina(n36561), .dinb(n36485), .dout(n36562));
  jxor g18540(.dina(n36477), .dinb(n324), .dout(n36563));
  jnot g18541(.din(n36563), .dout(n36564));
  jor  g18542(.dina(n36564), .dinb(n36562), .dout(n36565));
  jand g18543(.dina(n36565), .dinb(n36479), .dout(n36566));
  jxor g18544(.dina(n36471), .dinb(n325), .dout(n36567));
  jnot g18545(.din(n36567), .dout(n36568));
  jor  g18546(.dina(n36568), .dinb(n36566), .dout(n36569));
  jand g18547(.dina(n36569), .dinb(n36473), .dout(n36570));
  jxor g18548(.dina(n36465), .dinb(n439), .dout(n36571));
  jnot g18549(.din(n36571), .dout(n36572));
  jor  g18550(.dina(n36572), .dinb(n36570), .dout(n36573));
  jand g18551(.dina(n36573), .dinb(n36467), .dout(n36574));
  jxor g18552(.dina(n36459), .dinb(n440), .dout(n36575));
  jnot g18553(.din(n36575), .dout(n36576));
  jor  g18554(.dina(n36576), .dinb(n36574), .dout(n36577));
  jand g18555(.dina(n36577), .dinb(n36461), .dout(n36578));
  jxor g18556(.dina(n36453), .dinb(n435), .dout(n36579));
  jnot g18557(.din(n36579), .dout(n36580));
  jor  g18558(.dina(n36580), .dinb(n36578), .dout(n36581));
  jand g18559(.dina(n36581), .dinb(n36455), .dout(n36582));
  jxor g18560(.dina(n36447), .dinb(n436), .dout(n36583));
  jnot g18561(.din(n36583), .dout(n36584));
  jor  g18562(.dina(n36584), .dinb(n36582), .dout(n36585));
  jand g18563(.dina(n36585), .dinb(n36449), .dout(n36586));
  jxor g18564(.dina(n36441), .dinb(n432), .dout(n36587));
  jnot g18565(.din(n36587), .dout(n36588));
  jor  g18566(.dina(n36588), .dinb(n36586), .dout(n36589));
  jand g18567(.dina(n36589), .dinb(n36443), .dout(n36590));
  jxor g18568(.dina(n36435), .dinb(n433), .dout(n36591));
  jnot g18569(.din(n36591), .dout(n36592));
  jor  g18570(.dina(n36592), .dinb(n36590), .dout(n36593));
  jand g18571(.dina(n36593), .dinb(n36437), .dout(n36594));
  jxor g18572(.dina(n36429), .dinb(n421), .dout(n36595));
  jnot g18573(.din(n36595), .dout(n36596));
  jor  g18574(.dina(n36596), .dinb(n36594), .dout(n36597));
  jand g18575(.dina(n36597), .dinb(n36431), .dout(n36598));
  jxor g18576(.dina(n36423), .dinb(n422), .dout(n36599));
  jnot g18577(.din(n36599), .dout(n36600));
  jor  g18578(.dina(n36600), .dinb(n36598), .dout(n36601));
  jand g18579(.dina(n36601), .dinb(n36425), .dout(n36602));
  jxor g18580(.dina(n36417), .dinb(n416), .dout(n36603));
  jnot g18581(.din(n36603), .dout(n36604));
  jor  g18582(.dina(n36604), .dinb(n36602), .dout(n36605));
  jand g18583(.dina(n36605), .dinb(n36419), .dout(n36606));
  jxor g18584(.dina(n36411), .dinb(n417), .dout(n36607));
  jnot g18585(.din(n36607), .dout(n36608));
  jor  g18586(.dina(n36608), .dinb(n36606), .dout(n36609));
  jand g18587(.dina(n36609), .dinb(n36413), .dout(n36610));
  jxor g18588(.dina(n36405), .dinb(n2547), .dout(n36611));
  jnot g18589(.din(n36611), .dout(n36612));
  jor  g18590(.dina(n36612), .dinb(n36610), .dout(n36613));
  jand g18591(.dina(n36613), .dinb(n36407), .dout(n36614));
  jxor g18592(.dina(n36399), .dinb(n2714), .dout(n36615));
  jnot g18593(.din(n36615), .dout(n36616));
  jor  g18594(.dina(n36616), .dinb(n36614), .dout(n36617));
  jand g18595(.dina(n36617), .dinb(n36401), .dout(n36618));
  jxor g18596(.dina(n36393), .dinb(n405), .dout(n36619));
  jnot g18597(.din(n36619), .dout(n36620));
  jor  g18598(.dina(n36620), .dinb(n36618), .dout(n36621));
  jand g18599(.dina(n36621), .dinb(n36395), .dout(n36622));
  jxor g18600(.dina(n36387), .dinb(n406), .dout(n36623));
  jnot g18601(.din(n36623), .dout(n36624));
  jor  g18602(.dina(n36624), .dinb(n36622), .dout(n36625));
  jand g18603(.dina(n36625), .dinb(n36389), .dout(n36626));
  jxor g18604(.dina(n36381), .dinb(n412), .dout(n36627));
  jnot g18605(.din(n36627), .dout(n36628));
  jor  g18606(.dina(n36628), .dinb(n36626), .dout(n36629));
  jand g18607(.dina(n36629), .dinb(n36383), .dout(n36630));
  jxor g18608(.dina(n36375), .dinb(n413), .dout(n36631));
  jnot g18609(.din(n36631), .dout(n36632));
  jor  g18610(.dina(n36632), .dinb(n36630), .dout(n36633));
  jand g18611(.dina(n36633), .dinb(n36377), .dout(n36634));
  jxor g18612(.dina(n36369), .dinb(n409), .dout(n36635));
  jnot g18613(.din(n36635), .dout(n36636));
  jor  g18614(.dina(n36636), .dinb(n36634), .dout(n36637));
  jand g18615(.dina(n36637), .dinb(n36371), .dout(n36638));
  jxor g18616(.dina(n36363), .dinb(n410), .dout(n36639));
  jnot g18617(.din(n36639), .dout(n36640));
  jor  g18618(.dina(n36640), .dinb(n36638), .dout(n36641));
  jand g18619(.dina(n36641), .dinb(n36365), .dout(n36642));
  jxor g18620(.dina(n36357), .dinb(n426), .dout(n36643));
  jnot g18621(.din(n36643), .dout(n36644));
  jor  g18622(.dina(n36644), .dinb(n36642), .dout(n36645));
  jand g18623(.dina(n36645), .dinb(n36359), .dout(n36646));
  jxor g18624(.dina(n36351), .dinb(n427), .dout(n36647));
  jnot g18625(.din(n36647), .dout(n36648));
  jor  g18626(.dina(n36648), .dinb(n36646), .dout(n36649));
  jand g18627(.dina(n36649), .dinb(n36353), .dout(n36650));
  jxor g18628(.dina(n36345), .dinb(n424), .dout(n36651));
  jnot g18629(.din(n36651), .dout(n36652));
  jor  g18630(.dina(n36652), .dinb(n36650), .dout(n36653));
  jand g18631(.dina(n36653), .dinb(n36347), .dout(n36654));
  jxor g18632(.dina(n36339), .dinb(n300), .dout(n36655));
  jnot g18633(.din(n36655), .dout(n36656));
  jor  g18634(.dina(n36656), .dinb(n36654), .dout(n36657));
  jand g18635(.dina(n36657), .dinb(n36341), .dout(n36658));
  jxor g18636(.dina(n36333), .dinb(n297), .dout(n36659));
  jnot g18637(.din(n36659), .dout(n36660));
  jor  g18638(.dina(n36660), .dinb(n36658), .dout(n36661));
  jand g18639(.dina(n36661), .dinb(n36335), .dout(n36662));
  jxor g18640(.dina(n36327), .dinb(n298), .dout(n36663));
  jnot g18641(.din(n36663), .dout(n36664));
  jor  g18642(.dina(n36664), .dinb(n36662), .dout(n36665));
  jand g18643(.dina(n36665), .dinb(n36329), .dout(n36666));
  jxor g18644(.dina(n36321), .dinb(n301), .dout(n36667));
  jnot g18645(.din(n36667), .dout(n36668));
  jor  g18646(.dina(n36668), .dinb(n36666), .dout(n36669));
  jand g18647(.dina(n36669), .dinb(n36323), .dout(n36670));
  jxor g18648(.dina(n36315), .dinb(n293), .dout(n36671));
  jnot g18649(.din(n36671), .dout(n36672));
  jor  g18650(.dina(n36672), .dinb(n36670), .dout(n36673));
  jand g18651(.dina(n36673), .dinb(n36317), .dout(n36674));
  jxor g18652(.dina(n36309), .dinb(n294), .dout(n36675));
  jnot g18653(.din(n36675), .dout(n36676));
  jor  g18654(.dina(n36676), .dinb(n36674), .dout(n36677));
  jand g18655(.dina(n36677), .dinb(n36311), .dout(n36678));
  jxor g18656(.dina(n36303), .dinb(n290), .dout(n36679));
  jnot g18657(.din(n36679), .dout(n36680));
  jor  g18658(.dina(n36680), .dinb(n36678), .dout(n36681));
  jand g18659(.dina(n36681), .dinb(n36305), .dout(n36682));
  jxor g18660(.dina(n36297), .dinb(n291), .dout(n36683));
  jnot g18661(.din(n36683), .dout(n36684));
  jor  g18662(.dina(n36684), .dinb(n36682), .dout(n36685));
  jand g18663(.dina(n36685), .dinb(n36299), .dout(n36686));
  jxor g18664(.dina(n36291), .dinb(n284), .dout(n36687));
  jnot g18665(.din(n36687), .dout(n36688));
  jor  g18666(.dina(n36688), .dinb(n36686), .dout(n36689));
  jand g18667(.dina(n36689), .dinb(n36293), .dout(n36690));
  jxor g18668(.dina(n36285), .dinb(n285), .dout(n36691));
  jnot g18669(.din(n36691), .dout(n36692));
  jor  g18670(.dina(n36692), .dinb(n36690), .dout(n36693));
  jand g18671(.dina(n36693), .dinb(n36287), .dout(n36694));
  jxor g18672(.dina(n36279), .dinb(n281), .dout(n36695));
  jnot g18673(.din(n36695), .dout(n36696));
  jor  g18674(.dina(n36696), .dinb(n36694), .dout(n36697));
  jand g18675(.dina(n36697), .dinb(n36281), .dout(n36698));
  jxor g18676(.dina(n36273), .dinb(n282), .dout(n36699));
  jnot g18677(.din(n36699), .dout(n36700));
  jor  g18678(.dina(n36700), .dinb(n36698), .dout(n36701));
  jand g18679(.dina(n36701), .dinb(n36275), .dout(n36702));
  jxor g18680(.dina(n36267), .dinb(n397), .dout(n36703));
  jnot g18681(.din(n36703), .dout(n36704));
  jor  g18682(.dina(n36704), .dinb(n36702), .dout(n36705));
  jand g18683(.dina(n36705), .dinb(n36269), .dout(n36706));
  jxor g18684(.dina(n36261), .dinb(n513), .dout(n36707));
  jnot g18685(.din(n36707), .dout(n36708));
  jor  g18686(.dina(n36708), .dinb(n36706), .dout(n36709));
  jand g18687(.dina(n36709), .dinb(n36263), .dout(n36710));
  jxor g18688(.dina(n36255), .dinb(n514), .dout(n36711));
  jnot g18689(.din(n36711), .dout(n36712));
  jor  g18690(.dina(n36712), .dinb(n36710), .dout(n36713));
  jand g18691(.dina(n36713), .dinb(n36257), .dout(n36714));
  jxor g18692(.dina(n36249), .dinb(n510), .dout(n36715));
  jnot g18693(.din(n36715), .dout(n36716));
  jor  g18694(.dina(n36716), .dinb(n36714), .dout(n36717));
  jand g18695(.dina(n36717), .dinb(n36251), .dout(n36718));
  jxor g18696(.dina(n36243), .dinb(n396), .dout(n36719));
  jnot g18697(.din(n36719), .dout(n36720));
  jor  g18698(.dina(n36720), .dinb(n36718), .dout(n36721));
  jand g18699(.dina(n36721), .dinb(n36245), .dout(n36722));
  jxor g18700(.dina(n36237), .dinb(n383), .dout(n36723));
  jnot g18701(.din(n36723), .dout(n36724));
  jor  g18702(.dina(n36724), .dinb(n36722), .dout(n36725));
  jand g18703(.dina(n36725), .dinb(n36239), .dout(n36726));
  jxor g18704(.dina(n36231), .dinb(n12211), .dout(n36727));
  jnot g18705(.din(n36727), .dout(n36728));
  jor  g18706(.dina(n36728), .dinb(n36726), .dout(n36729));
  jand g18707(.dina(n36729), .dinb(n36233), .dout(n36730));
  jxor g18708(.dina(n36225), .dinb(n12214), .dout(n36731));
  jnot g18709(.din(n36731), .dout(n36732));
  jor  g18710(.dina(n36732), .dinb(n36730), .dout(n36733));
  jand g18711(.dina(n36733), .dinb(n36227), .dout(n36734));
  jxor g18712(.dina(n36219), .dinb(n384), .dout(n36735));
  jnot g18713(.din(n36735), .dout(n36736));
  jor  g18714(.dina(n36736), .dinb(n36734), .dout(n36737));
  jand g18715(.dina(n36737), .dinb(n36221), .dout(n36738));
  jxor g18716(.dina(n36213), .dinb(n374), .dout(n36739));
  jnot g18717(.din(n36739), .dout(n36740));
  jor  g18718(.dina(n36740), .dinb(n36738), .dout(n36741));
  jand g18719(.dina(n36741), .dinb(n36215), .dout(n36742));
  jand g18720(.dina(n36742), .dinb(n36200), .dout(n36743));
  jor  g18721(.dina(n36743), .dinb(n36198), .dout(n36744));
  jor  g18722(.dina(n36744), .dinb(n14055), .dout(n36745));
  jand g18723(.dina(n36745), .dinb(n36196), .dout(n36746));
  jxor g18724(.dina(n36531), .dinb(b1 ), .dout(n36747));
  jand g18725(.dina(n36747), .dinb(n14061), .dout(n36748));
  jor  g18726(.dina(n36748), .dinb(n36527), .dout(n36749));
  jand g18727(.dina(n36535), .dinb(n36749), .dout(n36750));
  jor  g18728(.dina(n36750), .dinb(n36520), .dout(n36751));
  jand g18729(.dina(n36539), .dinb(n36751), .dout(n36752));
  jor  g18730(.dina(n36752), .dinb(n36514), .dout(n36753));
  jand g18731(.dina(n36543), .dinb(n36753), .dout(n36754));
  jor  g18732(.dina(n36754), .dinb(n36508), .dout(n36755));
  jand g18733(.dina(n36547), .dinb(n36755), .dout(n36756));
  jor  g18734(.dina(n36756), .dinb(n36502), .dout(n36757));
  jand g18735(.dina(n36551), .dinb(n36757), .dout(n36758));
  jor  g18736(.dina(n36758), .dinb(n36496), .dout(n36759));
  jand g18737(.dina(n36555), .dinb(n36759), .dout(n36760));
  jor  g18738(.dina(n36760), .dinb(n36490), .dout(n36761));
  jand g18739(.dina(n36559), .dinb(n36761), .dout(n36762));
  jor  g18740(.dina(n36762), .dinb(n36484), .dout(n36763));
  jand g18741(.dina(n36563), .dinb(n36763), .dout(n36764));
  jor  g18742(.dina(n36764), .dinb(n36478), .dout(n36765));
  jand g18743(.dina(n36567), .dinb(n36765), .dout(n36766));
  jor  g18744(.dina(n36766), .dinb(n36472), .dout(n36767));
  jand g18745(.dina(n36571), .dinb(n36767), .dout(n36768));
  jor  g18746(.dina(n36768), .dinb(n36466), .dout(n36769));
  jand g18747(.dina(n36575), .dinb(n36769), .dout(n36770));
  jor  g18748(.dina(n36770), .dinb(n36460), .dout(n36771));
  jand g18749(.dina(n36579), .dinb(n36771), .dout(n36772));
  jor  g18750(.dina(n36772), .dinb(n36454), .dout(n36773));
  jand g18751(.dina(n36583), .dinb(n36773), .dout(n36774));
  jor  g18752(.dina(n36774), .dinb(n36448), .dout(n36775));
  jand g18753(.dina(n36587), .dinb(n36775), .dout(n36776));
  jor  g18754(.dina(n36776), .dinb(n36442), .dout(n36777));
  jand g18755(.dina(n36591), .dinb(n36777), .dout(n36778));
  jor  g18756(.dina(n36778), .dinb(n36436), .dout(n36779));
  jand g18757(.dina(n36595), .dinb(n36779), .dout(n36780));
  jor  g18758(.dina(n36780), .dinb(n36430), .dout(n36781));
  jand g18759(.dina(n36599), .dinb(n36781), .dout(n36782));
  jor  g18760(.dina(n36782), .dinb(n36424), .dout(n36783));
  jand g18761(.dina(n36603), .dinb(n36783), .dout(n36784));
  jor  g18762(.dina(n36784), .dinb(n36418), .dout(n36785));
  jand g18763(.dina(n36607), .dinb(n36785), .dout(n36786));
  jor  g18764(.dina(n36786), .dinb(n36412), .dout(n36787));
  jand g18765(.dina(n36611), .dinb(n36787), .dout(n36788));
  jor  g18766(.dina(n36788), .dinb(n36406), .dout(n36789));
  jand g18767(.dina(n36615), .dinb(n36789), .dout(n36790));
  jor  g18768(.dina(n36790), .dinb(n36400), .dout(n36791));
  jand g18769(.dina(n36619), .dinb(n36791), .dout(n36792));
  jor  g18770(.dina(n36792), .dinb(n36394), .dout(n36793));
  jand g18771(.dina(n36623), .dinb(n36793), .dout(n36794));
  jor  g18772(.dina(n36794), .dinb(n36388), .dout(n36795));
  jand g18773(.dina(n36627), .dinb(n36795), .dout(n36796));
  jor  g18774(.dina(n36796), .dinb(n36382), .dout(n36797));
  jand g18775(.dina(n36631), .dinb(n36797), .dout(n36798));
  jor  g18776(.dina(n36798), .dinb(n36376), .dout(n36799));
  jand g18777(.dina(n36635), .dinb(n36799), .dout(n36800));
  jor  g18778(.dina(n36800), .dinb(n36370), .dout(n36801));
  jand g18779(.dina(n36639), .dinb(n36801), .dout(n36802));
  jor  g18780(.dina(n36802), .dinb(n36364), .dout(n36803));
  jand g18781(.dina(n36643), .dinb(n36803), .dout(n36804));
  jor  g18782(.dina(n36804), .dinb(n36358), .dout(n36805));
  jand g18783(.dina(n36647), .dinb(n36805), .dout(n36806));
  jor  g18784(.dina(n36806), .dinb(n36352), .dout(n36807));
  jand g18785(.dina(n36651), .dinb(n36807), .dout(n36808));
  jor  g18786(.dina(n36808), .dinb(n36346), .dout(n36809));
  jand g18787(.dina(n36655), .dinb(n36809), .dout(n36810));
  jor  g18788(.dina(n36810), .dinb(n36340), .dout(n36811));
  jand g18789(.dina(n36659), .dinb(n36811), .dout(n36812));
  jor  g18790(.dina(n36812), .dinb(n36334), .dout(n36813));
  jand g18791(.dina(n36663), .dinb(n36813), .dout(n36814));
  jor  g18792(.dina(n36814), .dinb(n36328), .dout(n36815));
  jand g18793(.dina(n36667), .dinb(n36815), .dout(n36816));
  jor  g18794(.dina(n36816), .dinb(n36322), .dout(n36817));
  jand g18795(.dina(n36671), .dinb(n36817), .dout(n36818));
  jor  g18796(.dina(n36818), .dinb(n36316), .dout(n36819));
  jand g18797(.dina(n36675), .dinb(n36819), .dout(n36820));
  jor  g18798(.dina(n36820), .dinb(n36310), .dout(n36821));
  jand g18799(.dina(n36679), .dinb(n36821), .dout(n36822));
  jor  g18800(.dina(n36822), .dinb(n36304), .dout(n36823));
  jand g18801(.dina(n36683), .dinb(n36823), .dout(n36824));
  jor  g18802(.dina(n36824), .dinb(n36298), .dout(n36825));
  jand g18803(.dina(n36687), .dinb(n36825), .dout(n36826));
  jor  g18804(.dina(n36826), .dinb(n36292), .dout(n36827));
  jand g18805(.dina(n36691), .dinb(n36827), .dout(n36828));
  jor  g18806(.dina(n36828), .dinb(n36286), .dout(n36829));
  jand g18807(.dina(n36695), .dinb(n36829), .dout(n36830));
  jor  g18808(.dina(n36830), .dinb(n36280), .dout(n36831));
  jand g18809(.dina(n36699), .dinb(n36831), .dout(n36832));
  jor  g18810(.dina(n36832), .dinb(n36274), .dout(n36833));
  jand g18811(.dina(n36703), .dinb(n36833), .dout(n36834));
  jor  g18812(.dina(n36834), .dinb(n36268), .dout(n36835));
  jand g18813(.dina(n36707), .dinb(n36835), .dout(n36836));
  jor  g18814(.dina(n36836), .dinb(n36262), .dout(n36837));
  jand g18815(.dina(n36711), .dinb(n36837), .dout(n36838));
  jor  g18816(.dina(n36838), .dinb(n36256), .dout(n36839));
  jand g18817(.dina(n36715), .dinb(n36839), .dout(n36840));
  jor  g18818(.dina(n36840), .dinb(n36250), .dout(n36841));
  jand g18819(.dina(n36719), .dinb(n36841), .dout(n36842));
  jor  g18820(.dina(n36842), .dinb(n36244), .dout(n36843));
  jand g18821(.dina(n36723), .dinb(n36843), .dout(n36844));
  jor  g18822(.dina(n36844), .dinb(n36238), .dout(n36845));
  jand g18823(.dina(n36727), .dinb(n36845), .dout(n36846));
  jor  g18824(.dina(n36846), .dinb(n36232), .dout(n36847));
  jand g18825(.dina(n36731), .dinb(n36847), .dout(n36848));
  jor  g18826(.dina(n36848), .dinb(n36226), .dout(n36849));
  jand g18827(.dina(n36735), .dinb(n36849), .dout(n36850));
  jor  g18828(.dina(n36850), .dinb(n36220), .dout(n36851));
  jand g18829(.dina(n36739), .dinb(n36851), .dout(n36852));
  jor  g18830(.dina(n36852), .dinb(n36214), .dout(n36853));
  jand g18831(.dina(n36199), .dinb(n14054), .dout(n36854));
  jand g18832(.dina(n36854), .dinb(n36853), .dout(n36855));
  jor  g18833(.dina(n36855), .dinb(n36746), .dout(n36856));
  jand g18834(.dina(n36745), .dinb(n36213), .dout(n36857));
  jnot g18835(.din(n36198), .dout(n36858));
  jor  g18836(.dina(n36853), .dinb(n36199), .dout(n36859));
  jand g18837(.dina(n36859), .dinb(n36858), .dout(n36860));
  jand g18838(.dina(n36860), .dinb(n14054), .dout(n36861));
  jxor g18839(.dina(n36739), .dinb(n36851), .dout(n36862));
  jand g18840(.dina(n36862), .dinb(n36861), .dout(n36863));
  jor  g18841(.dina(n36863), .dinb(n36857), .dout(n36864));
  jand g18842(.dina(n36864), .dinb(n376), .dout(n36865));
  jand g18843(.dina(n36745), .dinb(n36219), .dout(n36866));
  jxor g18844(.dina(n36735), .dinb(n36849), .dout(n36867));
  jand g18845(.dina(n36867), .dinb(n36861), .dout(n36868));
  jor  g18846(.dina(n36868), .dinb(n36866), .dout(n36869));
  jand g18847(.dina(n36869), .dinb(n374), .dout(n36870));
  jand g18848(.dina(n36745), .dinb(n36225), .dout(n36871));
  jxor g18849(.dina(n36731), .dinb(n36847), .dout(n36872));
  jand g18850(.dina(n36872), .dinb(n36861), .dout(n36873));
  jor  g18851(.dina(n36873), .dinb(n36871), .dout(n36874));
  jand g18852(.dina(n36874), .dinb(n384), .dout(n36875));
  jand g18853(.dina(n36745), .dinb(n36231), .dout(n36876));
  jxor g18854(.dina(n36727), .dinb(n36845), .dout(n36877));
  jand g18855(.dina(n36877), .dinb(n36861), .dout(n36878));
  jor  g18856(.dina(n36878), .dinb(n36876), .dout(n36879));
  jand g18857(.dina(n36879), .dinb(n12214), .dout(n36880));
  jand g18858(.dina(n36745), .dinb(n36237), .dout(n36881));
  jxor g18859(.dina(n36723), .dinb(n36843), .dout(n36882));
  jand g18860(.dina(n36882), .dinb(n36861), .dout(n36883));
  jor  g18861(.dina(n36883), .dinb(n36881), .dout(n36884));
  jand g18862(.dina(n36884), .dinb(n12211), .dout(n36885));
  jand g18863(.dina(n36745), .dinb(n36243), .dout(n36886));
  jxor g18864(.dina(n36719), .dinb(n36841), .dout(n36887));
  jand g18865(.dina(n36887), .dinb(n36861), .dout(n36888));
  jor  g18866(.dina(n36888), .dinb(n36886), .dout(n36889));
  jand g18867(.dina(n36889), .dinb(n383), .dout(n36890));
  jand g18868(.dina(n36745), .dinb(n36249), .dout(n36891));
  jxor g18869(.dina(n36715), .dinb(n36839), .dout(n36892));
  jand g18870(.dina(n36892), .dinb(n36861), .dout(n36893));
  jor  g18871(.dina(n36893), .dinb(n36891), .dout(n36894));
  jand g18872(.dina(n36894), .dinb(n396), .dout(n36895));
  jand g18873(.dina(n36745), .dinb(n36255), .dout(n36896));
  jxor g18874(.dina(n36711), .dinb(n36837), .dout(n36897));
  jand g18875(.dina(n36897), .dinb(n36861), .dout(n36898));
  jor  g18876(.dina(n36898), .dinb(n36896), .dout(n36899));
  jand g18877(.dina(n36899), .dinb(n510), .dout(n36900));
  jand g18878(.dina(n36745), .dinb(n36261), .dout(n36901));
  jxor g18879(.dina(n36707), .dinb(n36835), .dout(n36902));
  jand g18880(.dina(n36902), .dinb(n36861), .dout(n36903));
  jor  g18881(.dina(n36903), .dinb(n36901), .dout(n36904));
  jand g18882(.dina(n36904), .dinb(n514), .dout(n36905));
  jand g18883(.dina(n36745), .dinb(n36267), .dout(n36906));
  jxor g18884(.dina(n36703), .dinb(n36833), .dout(n36907));
  jand g18885(.dina(n36907), .dinb(n36861), .dout(n36908));
  jor  g18886(.dina(n36908), .dinb(n36906), .dout(n36909));
  jand g18887(.dina(n36909), .dinb(n513), .dout(n36910));
  jand g18888(.dina(n36745), .dinb(n36273), .dout(n36911));
  jxor g18889(.dina(n36699), .dinb(n36831), .dout(n36912));
  jand g18890(.dina(n36912), .dinb(n36861), .dout(n36913));
  jor  g18891(.dina(n36913), .dinb(n36911), .dout(n36914));
  jand g18892(.dina(n36914), .dinb(n397), .dout(n36915));
  jand g18893(.dina(n36745), .dinb(n36279), .dout(n36916));
  jxor g18894(.dina(n36695), .dinb(n36829), .dout(n36917));
  jand g18895(.dina(n36917), .dinb(n36861), .dout(n36918));
  jor  g18896(.dina(n36918), .dinb(n36916), .dout(n36919));
  jand g18897(.dina(n36919), .dinb(n282), .dout(n36920));
  jand g18898(.dina(n36745), .dinb(n36285), .dout(n36921));
  jxor g18899(.dina(n36691), .dinb(n36827), .dout(n36922));
  jand g18900(.dina(n36922), .dinb(n36861), .dout(n36923));
  jor  g18901(.dina(n36923), .dinb(n36921), .dout(n36924));
  jand g18902(.dina(n36924), .dinb(n281), .dout(n36925));
  jand g18903(.dina(n36745), .dinb(n36291), .dout(n36926));
  jxor g18904(.dina(n36687), .dinb(n36825), .dout(n36927));
  jand g18905(.dina(n36927), .dinb(n36861), .dout(n36928));
  jor  g18906(.dina(n36928), .dinb(n36926), .dout(n36929));
  jand g18907(.dina(n36929), .dinb(n285), .dout(n36930));
  jand g18908(.dina(n36745), .dinb(n36297), .dout(n36931));
  jxor g18909(.dina(n36683), .dinb(n36823), .dout(n36932));
  jand g18910(.dina(n36932), .dinb(n36861), .dout(n36933));
  jor  g18911(.dina(n36933), .dinb(n36931), .dout(n36934));
  jand g18912(.dina(n36934), .dinb(n284), .dout(n36935));
  jand g18913(.dina(n36745), .dinb(n36303), .dout(n36936));
  jxor g18914(.dina(n36679), .dinb(n36821), .dout(n36937));
  jand g18915(.dina(n36937), .dinb(n36861), .dout(n36938));
  jor  g18916(.dina(n36938), .dinb(n36936), .dout(n36939));
  jand g18917(.dina(n36939), .dinb(n291), .dout(n36940));
  jand g18918(.dina(n36745), .dinb(n36309), .dout(n36941));
  jxor g18919(.dina(n36675), .dinb(n36819), .dout(n36942));
  jand g18920(.dina(n36942), .dinb(n36861), .dout(n36943));
  jor  g18921(.dina(n36943), .dinb(n36941), .dout(n36944));
  jand g18922(.dina(n36944), .dinb(n290), .dout(n36945));
  jand g18923(.dina(n36745), .dinb(n36315), .dout(n36946));
  jxor g18924(.dina(n36671), .dinb(n36817), .dout(n36947));
  jand g18925(.dina(n36947), .dinb(n36861), .dout(n36948));
  jor  g18926(.dina(n36948), .dinb(n36946), .dout(n36949));
  jand g18927(.dina(n36949), .dinb(n294), .dout(n36950));
  jand g18928(.dina(n36745), .dinb(n36321), .dout(n36951));
  jxor g18929(.dina(n36667), .dinb(n36815), .dout(n36952));
  jand g18930(.dina(n36952), .dinb(n36861), .dout(n36953));
  jor  g18931(.dina(n36953), .dinb(n36951), .dout(n36954));
  jand g18932(.dina(n36954), .dinb(n293), .dout(n36955));
  jand g18933(.dina(n36745), .dinb(n36327), .dout(n36956));
  jxor g18934(.dina(n36663), .dinb(n36813), .dout(n36957));
  jand g18935(.dina(n36957), .dinb(n36861), .dout(n36958));
  jor  g18936(.dina(n36958), .dinb(n36956), .dout(n36959));
  jand g18937(.dina(n36959), .dinb(n301), .dout(n36960));
  jand g18938(.dina(n36745), .dinb(n36333), .dout(n36961));
  jxor g18939(.dina(n36659), .dinb(n36811), .dout(n36962));
  jand g18940(.dina(n36962), .dinb(n36861), .dout(n36963));
  jor  g18941(.dina(n36963), .dinb(n36961), .dout(n36964));
  jand g18942(.dina(n36964), .dinb(n298), .dout(n36965));
  jand g18943(.dina(n36745), .dinb(n36339), .dout(n36966));
  jxor g18944(.dina(n36655), .dinb(n36809), .dout(n36967));
  jand g18945(.dina(n36967), .dinb(n36861), .dout(n36968));
  jor  g18946(.dina(n36968), .dinb(n36966), .dout(n36969));
  jand g18947(.dina(n36969), .dinb(n297), .dout(n36970));
  jand g18948(.dina(n36745), .dinb(n36345), .dout(n36971));
  jxor g18949(.dina(n36651), .dinb(n36807), .dout(n36972));
  jand g18950(.dina(n36972), .dinb(n36861), .dout(n36973));
  jor  g18951(.dina(n36973), .dinb(n36971), .dout(n36974));
  jand g18952(.dina(n36974), .dinb(n300), .dout(n36975));
  jand g18953(.dina(n36745), .dinb(n36351), .dout(n36976));
  jxor g18954(.dina(n36647), .dinb(n36805), .dout(n36977));
  jand g18955(.dina(n36977), .dinb(n36861), .dout(n36978));
  jor  g18956(.dina(n36978), .dinb(n36976), .dout(n36979));
  jand g18957(.dina(n36979), .dinb(n424), .dout(n36980));
  jand g18958(.dina(n36745), .dinb(n36357), .dout(n36981));
  jxor g18959(.dina(n36643), .dinb(n36803), .dout(n36982));
  jand g18960(.dina(n36982), .dinb(n36861), .dout(n36983));
  jor  g18961(.dina(n36983), .dinb(n36981), .dout(n36984));
  jand g18962(.dina(n36984), .dinb(n427), .dout(n36985));
  jand g18963(.dina(n36745), .dinb(n36363), .dout(n36986));
  jxor g18964(.dina(n36639), .dinb(n36801), .dout(n36987));
  jand g18965(.dina(n36987), .dinb(n36861), .dout(n36988));
  jor  g18966(.dina(n36988), .dinb(n36986), .dout(n36989));
  jand g18967(.dina(n36989), .dinb(n426), .dout(n36990));
  jand g18968(.dina(n36745), .dinb(n36369), .dout(n36991));
  jxor g18969(.dina(n36635), .dinb(n36799), .dout(n36992));
  jand g18970(.dina(n36992), .dinb(n36861), .dout(n36993));
  jor  g18971(.dina(n36993), .dinb(n36991), .dout(n36994));
  jand g18972(.dina(n36994), .dinb(n410), .dout(n36995));
  jand g18973(.dina(n36745), .dinb(n36375), .dout(n36996));
  jxor g18974(.dina(n36631), .dinb(n36797), .dout(n36997));
  jand g18975(.dina(n36997), .dinb(n36861), .dout(n36998));
  jor  g18976(.dina(n36998), .dinb(n36996), .dout(n36999));
  jand g18977(.dina(n36999), .dinb(n409), .dout(n37000));
  jand g18978(.dina(n36745), .dinb(n36381), .dout(n37001));
  jxor g18979(.dina(n36627), .dinb(n36795), .dout(n37002));
  jand g18980(.dina(n37002), .dinb(n36861), .dout(n37003));
  jor  g18981(.dina(n37003), .dinb(n37001), .dout(n37004));
  jand g18982(.dina(n37004), .dinb(n413), .dout(n37005));
  jand g18983(.dina(n36745), .dinb(n36387), .dout(n37006));
  jxor g18984(.dina(n36623), .dinb(n36793), .dout(n37007));
  jand g18985(.dina(n37007), .dinb(n36861), .dout(n37008));
  jor  g18986(.dina(n37008), .dinb(n37006), .dout(n37009));
  jand g18987(.dina(n37009), .dinb(n412), .dout(n37010));
  jand g18988(.dina(n36745), .dinb(n36393), .dout(n37011));
  jxor g18989(.dina(n36619), .dinb(n36791), .dout(n37012));
  jand g18990(.dina(n37012), .dinb(n36861), .dout(n37013));
  jor  g18991(.dina(n37013), .dinb(n37011), .dout(n37014));
  jand g18992(.dina(n37014), .dinb(n406), .dout(n37015));
  jand g18993(.dina(n36745), .dinb(n36399), .dout(n37016));
  jxor g18994(.dina(n36615), .dinb(n36789), .dout(n37017));
  jand g18995(.dina(n37017), .dinb(n36861), .dout(n37018));
  jor  g18996(.dina(n37018), .dinb(n37016), .dout(n37019));
  jand g18997(.dina(n37019), .dinb(n405), .dout(n37020));
  jand g18998(.dina(n36745), .dinb(n36405), .dout(n37021));
  jxor g18999(.dina(n36611), .dinb(n36787), .dout(n37022));
  jand g19000(.dina(n37022), .dinb(n36861), .dout(n37023));
  jor  g19001(.dina(n37023), .dinb(n37021), .dout(n37024));
  jand g19002(.dina(n37024), .dinb(n2714), .dout(n37025));
  jand g19003(.dina(n36745), .dinb(n36411), .dout(n37026));
  jxor g19004(.dina(n36607), .dinb(n36785), .dout(n37027));
  jand g19005(.dina(n37027), .dinb(n36861), .dout(n37028));
  jor  g19006(.dina(n37028), .dinb(n37026), .dout(n37029));
  jand g19007(.dina(n37029), .dinb(n2547), .dout(n37030));
  jand g19008(.dina(n36745), .dinb(n36417), .dout(n37031));
  jxor g19009(.dina(n36603), .dinb(n36783), .dout(n37032));
  jand g19010(.dina(n37032), .dinb(n36861), .dout(n37033));
  jor  g19011(.dina(n37033), .dinb(n37031), .dout(n37034));
  jand g19012(.dina(n37034), .dinb(n417), .dout(n37035));
  jand g19013(.dina(n36745), .dinb(n36423), .dout(n37036));
  jxor g19014(.dina(n36599), .dinb(n36781), .dout(n37037));
  jand g19015(.dina(n37037), .dinb(n36861), .dout(n37038));
  jor  g19016(.dina(n37038), .dinb(n37036), .dout(n37039));
  jand g19017(.dina(n37039), .dinb(n416), .dout(n37040));
  jand g19018(.dina(n36745), .dinb(n36429), .dout(n37041));
  jxor g19019(.dina(n36595), .dinb(n36779), .dout(n37042));
  jand g19020(.dina(n37042), .dinb(n36861), .dout(n37043));
  jor  g19021(.dina(n37043), .dinb(n37041), .dout(n37044));
  jand g19022(.dina(n37044), .dinb(n422), .dout(n37045));
  jand g19023(.dina(n36745), .dinb(n36435), .dout(n37046));
  jxor g19024(.dina(n36591), .dinb(n36777), .dout(n37047));
  jand g19025(.dina(n37047), .dinb(n36861), .dout(n37048));
  jor  g19026(.dina(n37048), .dinb(n37046), .dout(n37049));
  jand g19027(.dina(n37049), .dinb(n421), .dout(n37050));
  jand g19028(.dina(n36745), .dinb(n36441), .dout(n37051));
  jxor g19029(.dina(n36587), .dinb(n36775), .dout(n37052));
  jand g19030(.dina(n37052), .dinb(n36861), .dout(n37053));
  jor  g19031(.dina(n37053), .dinb(n37051), .dout(n37054));
  jand g19032(.dina(n37054), .dinb(n433), .dout(n37055));
  jand g19033(.dina(n36745), .dinb(n36447), .dout(n37056));
  jxor g19034(.dina(n36583), .dinb(n36773), .dout(n37057));
  jand g19035(.dina(n37057), .dinb(n36861), .dout(n37058));
  jor  g19036(.dina(n37058), .dinb(n37056), .dout(n37059));
  jand g19037(.dina(n37059), .dinb(n432), .dout(n37060));
  jand g19038(.dina(n36745), .dinb(n36453), .dout(n37061));
  jxor g19039(.dina(n36579), .dinb(n36771), .dout(n37062));
  jand g19040(.dina(n37062), .dinb(n36861), .dout(n37063));
  jor  g19041(.dina(n37063), .dinb(n37061), .dout(n37064));
  jand g19042(.dina(n37064), .dinb(n436), .dout(n37065));
  jand g19043(.dina(n36745), .dinb(n36459), .dout(n37066));
  jxor g19044(.dina(n36575), .dinb(n36769), .dout(n37067));
  jand g19045(.dina(n37067), .dinb(n36861), .dout(n37068));
  jor  g19046(.dina(n37068), .dinb(n37066), .dout(n37069));
  jand g19047(.dina(n37069), .dinb(n435), .dout(n37070));
  jand g19048(.dina(n36745), .dinb(n36465), .dout(n37071));
  jxor g19049(.dina(n36571), .dinb(n36767), .dout(n37072));
  jand g19050(.dina(n37072), .dinb(n36861), .dout(n37073));
  jor  g19051(.dina(n37073), .dinb(n37071), .dout(n37074));
  jand g19052(.dina(n37074), .dinb(n440), .dout(n37075));
  jand g19053(.dina(n36745), .dinb(n36471), .dout(n37076));
  jxor g19054(.dina(n36567), .dinb(n36765), .dout(n37077));
  jand g19055(.dina(n37077), .dinb(n36861), .dout(n37078));
  jor  g19056(.dina(n37078), .dinb(n37076), .dout(n37079));
  jand g19057(.dina(n37079), .dinb(n439), .dout(n37080));
  jand g19058(.dina(n36745), .dinb(n36477), .dout(n37081));
  jxor g19059(.dina(n36563), .dinb(n36763), .dout(n37082));
  jand g19060(.dina(n37082), .dinb(n36861), .dout(n37083));
  jor  g19061(.dina(n37083), .dinb(n37081), .dout(n37084));
  jand g19062(.dina(n37084), .dinb(n325), .dout(n37085));
  jand g19063(.dina(n36745), .dinb(n36483), .dout(n37086));
  jxor g19064(.dina(n36559), .dinb(n36761), .dout(n37087));
  jand g19065(.dina(n37087), .dinb(n36861), .dout(n37088));
  jor  g19066(.dina(n37088), .dinb(n37086), .dout(n37089));
  jand g19067(.dina(n37089), .dinb(n324), .dout(n37090));
  jand g19068(.dina(n36745), .dinb(n36489), .dout(n37091));
  jxor g19069(.dina(n36555), .dinb(n36759), .dout(n37092));
  jand g19070(.dina(n37092), .dinb(n36861), .dout(n37093));
  jor  g19071(.dina(n37093), .dinb(n37091), .dout(n37094));
  jand g19072(.dina(n37094), .dinb(n323), .dout(n37095));
  jand g19073(.dina(n36745), .dinb(n36495), .dout(n37096));
  jxor g19074(.dina(n36551), .dinb(n36757), .dout(n37097));
  jand g19075(.dina(n37097), .dinb(n36861), .dout(n37098));
  jor  g19076(.dina(n37098), .dinb(n37096), .dout(n37099));
  jand g19077(.dina(n37099), .dinb(n335), .dout(n37100));
  jand g19078(.dina(n36745), .dinb(n36501), .dout(n37101));
  jxor g19079(.dina(n36547), .dinb(n36755), .dout(n37102));
  jand g19080(.dina(n37102), .dinb(n36861), .dout(n37103));
  jor  g19081(.dina(n37103), .dinb(n37101), .dout(n37104));
  jand g19082(.dina(n37104), .dinb(n334), .dout(n37105));
  jand g19083(.dina(n36745), .dinb(n36507), .dout(n37106));
  jxor g19084(.dina(n36543), .dinb(n36753), .dout(n37107));
  jand g19085(.dina(n37107), .dinb(n36861), .dout(n37108));
  jor  g19086(.dina(n37108), .dinb(n37106), .dout(n37109));
  jand g19087(.dina(n37109), .dinb(n338), .dout(n37110));
  jand g19088(.dina(n36745), .dinb(n36513), .dout(n37111));
  jxor g19089(.dina(n36539), .dinb(n36751), .dout(n37112));
  jand g19090(.dina(n37112), .dinb(n36861), .dout(n37113));
  jor  g19091(.dina(n37113), .dinb(n37111), .dout(n37114));
  jand g19092(.dina(n37114), .dinb(n337), .dout(n37115));
  jand g19093(.dina(n36745), .dinb(n36519), .dout(n37116));
  jxor g19094(.dina(n36535), .dinb(n36749), .dout(n37117));
  jand g19095(.dina(n37117), .dinb(n36861), .dout(n37118));
  jor  g19096(.dina(n37118), .dinb(n37116), .dout(n37119));
  jand g19097(.dina(n37119), .dinb(n344), .dout(n37120));
  jor  g19098(.dina(n36861), .dinb(n36531), .dout(n37121));
  jxor g19099(.dina(n36747), .dinb(n14061), .dout(n37122));
  jnot g19100(.din(n37122), .dout(n37123));
  jor  g19101(.dina(n37123), .dinb(n36745), .dout(n37124));
  jand g19102(.dina(n37124), .dinb(n37121), .dout(n37125));
  jnot g19103(.din(n37125), .dout(n37126));
  jand g19104(.dina(n37126), .dinb(n348), .dout(n37127));
  jand g19105(.dina(n36860), .dinb(n14440), .dout(n37128));
  jxor g19106(.dina(n37128), .dinb(a9 ), .dout(n37129));
  jand g19107(.dina(n37129), .dinb(n258), .dout(n37130));
  jxor g19108(.dina(n37128), .dinb(n13837), .dout(n37131));
  jxor g19109(.dina(n37131), .dinb(b1 ), .dout(n37132));
  jand g19110(.dina(n37132), .dinb(n14449), .dout(n37133));
  jor  g19111(.dina(n37133), .dinb(n37130), .dout(n37134));
  jxor g19112(.dina(n37125), .dinb(b2 ), .dout(n37135));
  jand g19113(.dina(n37135), .dinb(n37134), .dout(n37136));
  jor  g19114(.dina(n37136), .dinb(n37127), .dout(n37137));
  jxor g19115(.dina(n37119), .dinb(n344), .dout(n37138));
  jand g19116(.dina(n37138), .dinb(n37137), .dout(n37139));
  jor  g19117(.dina(n37139), .dinb(n37120), .dout(n37140));
  jxor g19118(.dina(n37114), .dinb(n337), .dout(n37141));
  jand g19119(.dina(n37141), .dinb(n37140), .dout(n37142));
  jor  g19120(.dina(n37142), .dinb(n37115), .dout(n37143));
  jxor g19121(.dina(n37109), .dinb(n338), .dout(n37144));
  jand g19122(.dina(n37144), .dinb(n37143), .dout(n37145));
  jor  g19123(.dina(n37145), .dinb(n37110), .dout(n37146));
  jxor g19124(.dina(n37104), .dinb(n334), .dout(n37147));
  jand g19125(.dina(n37147), .dinb(n37146), .dout(n37148));
  jor  g19126(.dina(n37148), .dinb(n37105), .dout(n37149));
  jxor g19127(.dina(n37099), .dinb(n335), .dout(n37150));
  jand g19128(.dina(n37150), .dinb(n37149), .dout(n37151));
  jor  g19129(.dina(n37151), .dinb(n37100), .dout(n37152));
  jxor g19130(.dina(n37094), .dinb(n323), .dout(n37153));
  jand g19131(.dina(n37153), .dinb(n37152), .dout(n37154));
  jor  g19132(.dina(n37154), .dinb(n37095), .dout(n37155));
  jxor g19133(.dina(n37089), .dinb(n324), .dout(n37156));
  jand g19134(.dina(n37156), .dinb(n37155), .dout(n37157));
  jor  g19135(.dina(n37157), .dinb(n37090), .dout(n37158));
  jxor g19136(.dina(n37084), .dinb(n325), .dout(n37159));
  jand g19137(.dina(n37159), .dinb(n37158), .dout(n37160));
  jor  g19138(.dina(n37160), .dinb(n37085), .dout(n37161));
  jxor g19139(.dina(n37079), .dinb(n439), .dout(n37162));
  jand g19140(.dina(n37162), .dinb(n37161), .dout(n37163));
  jor  g19141(.dina(n37163), .dinb(n37080), .dout(n37164));
  jxor g19142(.dina(n37074), .dinb(n440), .dout(n37165));
  jand g19143(.dina(n37165), .dinb(n37164), .dout(n37166));
  jor  g19144(.dina(n37166), .dinb(n37075), .dout(n37167));
  jxor g19145(.dina(n37069), .dinb(n435), .dout(n37168));
  jand g19146(.dina(n37168), .dinb(n37167), .dout(n37169));
  jor  g19147(.dina(n37169), .dinb(n37070), .dout(n37170));
  jxor g19148(.dina(n37064), .dinb(n436), .dout(n37171));
  jand g19149(.dina(n37171), .dinb(n37170), .dout(n37172));
  jor  g19150(.dina(n37172), .dinb(n37065), .dout(n37173));
  jxor g19151(.dina(n37059), .dinb(n432), .dout(n37174));
  jand g19152(.dina(n37174), .dinb(n37173), .dout(n37175));
  jor  g19153(.dina(n37175), .dinb(n37060), .dout(n37176));
  jxor g19154(.dina(n37054), .dinb(n433), .dout(n37177));
  jand g19155(.dina(n37177), .dinb(n37176), .dout(n37178));
  jor  g19156(.dina(n37178), .dinb(n37055), .dout(n37179));
  jxor g19157(.dina(n37049), .dinb(n421), .dout(n37180));
  jand g19158(.dina(n37180), .dinb(n37179), .dout(n37181));
  jor  g19159(.dina(n37181), .dinb(n37050), .dout(n37182));
  jxor g19160(.dina(n37044), .dinb(n422), .dout(n37183));
  jand g19161(.dina(n37183), .dinb(n37182), .dout(n37184));
  jor  g19162(.dina(n37184), .dinb(n37045), .dout(n37185));
  jxor g19163(.dina(n37039), .dinb(n416), .dout(n37186));
  jand g19164(.dina(n37186), .dinb(n37185), .dout(n37187));
  jor  g19165(.dina(n37187), .dinb(n37040), .dout(n37188));
  jxor g19166(.dina(n37034), .dinb(n417), .dout(n37189));
  jand g19167(.dina(n37189), .dinb(n37188), .dout(n37190));
  jor  g19168(.dina(n37190), .dinb(n37035), .dout(n37191));
  jxor g19169(.dina(n37029), .dinb(n2547), .dout(n37192));
  jand g19170(.dina(n37192), .dinb(n37191), .dout(n37193));
  jor  g19171(.dina(n37193), .dinb(n37030), .dout(n37194));
  jxor g19172(.dina(n37024), .dinb(n2714), .dout(n37195));
  jand g19173(.dina(n37195), .dinb(n37194), .dout(n37196));
  jor  g19174(.dina(n37196), .dinb(n37025), .dout(n37197));
  jxor g19175(.dina(n37019), .dinb(n405), .dout(n37198));
  jand g19176(.dina(n37198), .dinb(n37197), .dout(n37199));
  jor  g19177(.dina(n37199), .dinb(n37020), .dout(n37200));
  jxor g19178(.dina(n37014), .dinb(n406), .dout(n37201));
  jand g19179(.dina(n37201), .dinb(n37200), .dout(n37202));
  jor  g19180(.dina(n37202), .dinb(n37015), .dout(n37203));
  jxor g19181(.dina(n37009), .dinb(n412), .dout(n37204));
  jand g19182(.dina(n37204), .dinb(n37203), .dout(n37205));
  jor  g19183(.dina(n37205), .dinb(n37010), .dout(n37206));
  jxor g19184(.dina(n37004), .dinb(n413), .dout(n37207));
  jand g19185(.dina(n37207), .dinb(n37206), .dout(n37208));
  jor  g19186(.dina(n37208), .dinb(n37005), .dout(n37209));
  jxor g19187(.dina(n36999), .dinb(n409), .dout(n37210));
  jand g19188(.dina(n37210), .dinb(n37209), .dout(n37211));
  jor  g19189(.dina(n37211), .dinb(n37000), .dout(n37212));
  jxor g19190(.dina(n36994), .dinb(n410), .dout(n37213));
  jand g19191(.dina(n37213), .dinb(n37212), .dout(n37214));
  jor  g19192(.dina(n37214), .dinb(n36995), .dout(n37215));
  jxor g19193(.dina(n36989), .dinb(n426), .dout(n37216));
  jand g19194(.dina(n37216), .dinb(n37215), .dout(n37217));
  jor  g19195(.dina(n37217), .dinb(n36990), .dout(n37218));
  jxor g19196(.dina(n36984), .dinb(n427), .dout(n37219));
  jand g19197(.dina(n37219), .dinb(n37218), .dout(n37220));
  jor  g19198(.dina(n37220), .dinb(n36985), .dout(n37221));
  jxor g19199(.dina(n36979), .dinb(n424), .dout(n37222));
  jand g19200(.dina(n37222), .dinb(n37221), .dout(n37223));
  jor  g19201(.dina(n37223), .dinb(n36980), .dout(n37224));
  jxor g19202(.dina(n36974), .dinb(n300), .dout(n37225));
  jand g19203(.dina(n37225), .dinb(n37224), .dout(n37226));
  jor  g19204(.dina(n37226), .dinb(n36975), .dout(n37227));
  jxor g19205(.dina(n36969), .dinb(n297), .dout(n37228));
  jand g19206(.dina(n37228), .dinb(n37227), .dout(n37229));
  jor  g19207(.dina(n37229), .dinb(n36970), .dout(n37230));
  jxor g19208(.dina(n36964), .dinb(n298), .dout(n37231));
  jand g19209(.dina(n37231), .dinb(n37230), .dout(n37232));
  jor  g19210(.dina(n37232), .dinb(n36965), .dout(n37233));
  jxor g19211(.dina(n36959), .dinb(n301), .dout(n37234));
  jand g19212(.dina(n37234), .dinb(n37233), .dout(n37235));
  jor  g19213(.dina(n37235), .dinb(n36960), .dout(n37236));
  jxor g19214(.dina(n36954), .dinb(n293), .dout(n37237));
  jand g19215(.dina(n37237), .dinb(n37236), .dout(n37238));
  jor  g19216(.dina(n37238), .dinb(n36955), .dout(n37239));
  jxor g19217(.dina(n36949), .dinb(n294), .dout(n37240));
  jand g19218(.dina(n37240), .dinb(n37239), .dout(n37241));
  jor  g19219(.dina(n37241), .dinb(n36950), .dout(n37242));
  jxor g19220(.dina(n36944), .dinb(n290), .dout(n37243));
  jand g19221(.dina(n37243), .dinb(n37242), .dout(n37244));
  jor  g19222(.dina(n37244), .dinb(n36945), .dout(n37245));
  jxor g19223(.dina(n36939), .dinb(n291), .dout(n37246));
  jand g19224(.dina(n37246), .dinb(n37245), .dout(n37247));
  jor  g19225(.dina(n37247), .dinb(n36940), .dout(n37248));
  jxor g19226(.dina(n36934), .dinb(n284), .dout(n37249));
  jand g19227(.dina(n37249), .dinb(n37248), .dout(n37250));
  jor  g19228(.dina(n37250), .dinb(n36935), .dout(n37251));
  jxor g19229(.dina(n36929), .dinb(n285), .dout(n37252));
  jand g19230(.dina(n37252), .dinb(n37251), .dout(n37253));
  jor  g19231(.dina(n37253), .dinb(n36930), .dout(n37254));
  jxor g19232(.dina(n36924), .dinb(n281), .dout(n37255));
  jand g19233(.dina(n37255), .dinb(n37254), .dout(n37256));
  jor  g19234(.dina(n37256), .dinb(n36925), .dout(n37257));
  jxor g19235(.dina(n36919), .dinb(n282), .dout(n37258));
  jand g19236(.dina(n37258), .dinb(n37257), .dout(n37259));
  jor  g19237(.dina(n37259), .dinb(n36920), .dout(n37260));
  jxor g19238(.dina(n36914), .dinb(n397), .dout(n37261));
  jand g19239(.dina(n37261), .dinb(n37260), .dout(n37262));
  jor  g19240(.dina(n37262), .dinb(n36915), .dout(n37263));
  jxor g19241(.dina(n36909), .dinb(n513), .dout(n37264));
  jand g19242(.dina(n37264), .dinb(n37263), .dout(n37265));
  jor  g19243(.dina(n37265), .dinb(n36910), .dout(n37266));
  jxor g19244(.dina(n36904), .dinb(n514), .dout(n37267));
  jand g19245(.dina(n37267), .dinb(n37266), .dout(n37268));
  jor  g19246(.dina(n37268), .dinb(n36905), .dout(n37269));
  jxor g19247(.dina(n36899), .dinb(n510), .dout(n37270));
  jand g19248(.dina(n37270), .dinb(n37269), .dout(n37271));
  jor  g19249(.dina(n37271), .dinb(n36900), .dout(n37272));
  jxor g19250(.dina(n36894), .dinb(n396), .dout(n37273));
  jand g19251(.dina(n37273), .dinb(n37272), .dout(n37274));
  jor  g19252(.dina(n37274), .dinb(n36895), .dout(n37275));
  jxor g19253(.dina(n36889), .dinb(n383), .dout(n37276));
  jand g19254(.dina(n37276), .dinb(n37275), .dout(n37277));
  jor  g19255(.dina(n37277), .dinb(n36890), .dout(n37278));
  jxor g19256(.dina(n36884), .dinb(n12211), .dout(n37279));
  jand g19257(.dina(n37279), .dinb(n37278), .dout(n37280));
  jor  g19258(.dina(n37280), .dinb(n36885), .dout(n37281));
  jxor g19259(.dina(n36879), .dinb(n12214), .dout(n37282));
  jand g19260(.dina(n37282), .dinb(n37281), .dout(n37283));
  jor  g19261(.dina(n37283), .dinb(n36880), .dout(n37284));
  jxor g19262(.dina(n36874), .dinb(n384), .dout(n37285));
  jand g19263(.dina(n37285), .dinb(n37284), .dout(n37286));
  jor  g19264(.dina(n37286), .dinb(n36875), .dout(n37287));
  jxor g19265(.dina(n36869), .dinb(n374), .dout(n37288));
  jand g19266(.dina(n37288), .dinb(n37287), .dout(n37289));
  jor  g19267(.dina(n37289), .dinb(n36870), .dout(n37290));
  jxor g19268(.dina(n36864), .dinb(n376), .dout(n37291));
  jand g19269(.dina(n37291), .dinb(n37290), .dout(n37292));
  jor  g19270(.dina(n37292), .dinb(n36865), .dout(n37293));
  jand g19271(.dina(n37293), .dinb(n377), .dout(n37294));
  jnot g19272(.din(n36865), .dout(n37295));
  jnot g19273(.din(n36870), .dout(n37296));
  jnot g19274(.din(n36875), .dout(n37297));
  jnot g19275(.din(n36880), .dout(n37298));
  jnot g19276(.din(n36885), .dout(n37299));
  jnot g19277(.din(n36890), .dout(n37300));
  jnot g19278(.din(n36895), .dout(n37301));
  jnot g19279(.din(n36900), .dout(n37302));
  jnot g19280(.din(n36905), .dout(n37303));
  jnot g19281(.din(n36910), .dout(n37304));
  jnot g19282(.din(n36915), .dout(n37305));
  jnot g19283(.din(n36920), .dout(n37306));
  jnot g19284(.din(n36925), .dout(n37307));
  jnot g19285(.din(n36930), .dout(n37308));
  jnot g19286(.din(n36935), .dout(n37309));
  jnot g19287(.din(n36940), .dout(n37310));
  jnot g19288(.din(n36945), .dout(n37311));
  jnot g19289(.din(n36950), .dout(n37312));
  jnot g19290(.din(n36955), .dout(n37313));
  jnot g19291(.din(n36960), .dout(n37314));
  jnot g19292(.din(n36965), .dout(n37315));
  jnot g19293(.din(n36970), .dout(n37316));
  jnot g19294(.din(n36975), .dout(n37317));
  jnot g19295(.din(n36980), .dout(n37318));
  jnot g19296(.din(n36985), .dout(n37319));
  jnot g19297(.din(n36990), .dout(n37320));
  jnot g19298(.din(n36995), .dout(n37321));
  jnot g19299(.din(n37000), .dout(n37322));
  jnot g19300(.din(n37005), .dout(n37323));
  jnot g19301(.din(n37010), .dout(n37324));
  jnot g19302(.din(n37015), .dout(n37325));
  jnot g19303(.din(n37020), .dout(n37326));
  jnot g19304(.din(n37025), .dout(n37327));
  jnot g19305(.din(n37030), .dout(n37328));
  jnot g19306(.din(n37035), .dout(n37329));
  jnot g19307(.din(n37040), .dout(n37330));
  jnot g19308(.din(n37045), .dout(n37331));
  jnot g19309(.din(n37050), .dout(n37332));
  jnot g19310(.din(n37055), .dout(n37333));
  jnot g19311(.din(n37060), .dout(n37334));
  jnot g19312(.din(n37065), .dout(n37335));
  jnot g19313(.din(n37070), .dout(n37336));
  jnot g19314(.din(n37075), .dout(n37337));
  jnot g19315(.din(n37080), .dout(n37338));
  jnot g19316(.din(n37085), .dout(n37339));
  jnot g19317(.din(n37090), .dout(n37340));
  jnot g19318(.din(n37095), .dout(n37341));
  jnot g19319(.din(n37100), .dout(n37342));
  jnot g19320(.din(n37105), .dout(n37343));
  jnot g19321(.din(n37110), .dout(n37344));
  jnot g19322(.din(n37115), .dout(n37345));
  jnot g19323(.din(n37120), .dout(n37346));
  jnot g19324(.din(n37127), .dout(n37347));
  jnot g19325(.din(n37130), .dout(n37348));
  jxor g19326(.dina(n37131), .dinb(n258), .dout(n37349));
  jor  g19327(.dina(n37349), .dinb(n14448), .dout(n37350));
  jand g19328(.dina(n37350), .dinb(n37348), .dout(n37351));
  jnot g19329(.din(n37135), .dout(n37352));
  jor  g19330(.dina(n37352), .dinb(n37351), .dout(n37353));
  jand g19331(.dina(n37353), .dinb(n37347), .dout(n37354));
  jnot g19332(.din(n37138), .dout(n37355));
  jor  g19333(.dina(n37355), .dinb(n37354), .dout(n37356));
  jand g19334(.dina(n37356), .dinb(n37346), .dout(n37357));
  jnot g19335(.din(n37141), .dout(n37358));
  jor  g19336(.dina(n37358), .dinb(n37357), .dout(n37359));
  jand g19337(.dina(n37359), .dinb(n37345), .dout(n37360));
  jnot g19338(.din(n37144), .dout(n37361));
  jor  g19339(.dina(n37361), .dinb(n37360), .dout(n37362));
  jand g19340(.dina(n37362), .dinb(n37344), .dout(n37363));
  jnot g19341(.din(n37147), .dout(n37364));
  jor  g19342(.dina(n37364), .dinb(n37363), .dout(n37365));
  jand g19343(.dina(n37365), .dinb(n37343), .dout(n37366));
  jnot g19344(.din(n37150), .dout(n37367));
  jor  g19345(.dina(n37367), .dinb(n37366), .dout(n37368));
  jand g19346(.dina(n37368), .dinb(n37342), .dout(n37369));
  jnot g19347(.din(n37153), .dout(n37370));
  jor  g19348(.dina(n37370), .dinb(n37369), .dout(n37371));
  jand g19349(.dina(n37371), .dinb(n37341), .dout(n37372));
  jnot g19350(.din(n37156), .dout(n37373));
  jor  g19351(.dina(n37373), .dinb(n37372), .dout(n37374));
  jand g19352(.dina(n37374), .dinb(n37340), .dout(n37375));
  jnot g19353(.din(n37159), .dout(n37376));
  jor  g19354(.dina(n37376), .dinb(n37375), .dout(n37377));
  jand g19355(.dina(n37377), .dinb(n37339), .dout(n37378));
  jnot g19356(.din(n37162), .dout(n37379));
  jor  g19357(.dina(n37379), .dinb(n37378), .dout(n37380));
  jand g19358(.dina(n37380), .dinb(n37338), .dout(n37381));
  jnot g19359(.din(n37165), .dout(n37382));
  jor  g19360(.dina(n37382), .dinb(n37381), .dout(n37383));
  jand g19361(.dina(n37383), .dinb(n37337), .dout(n37384));
  jnot g19362(.din(n37168), .dout(n37385));
  jor  g19363(.dina(n37385), .dinb(n37384), .dout(n37386));
  jand g19364(.dina(n37386), .dinb(n37336), .dout(n37387));
  jnot g19365(.din(n37171), .dout(n37388));
  jor  g19366(.dina(n37388), .dinb(n37387), .dout(n37389));
  jand g19367(.dina(n37389), .dinb(n37335), .dout(n37390));
  jnot g19368(.din(n37174), .dout(n37391));
  jor  g19369(.dina(n37391), .dinb(n37390), .dout(n37392));
  jand g19370(.dina(n37392), .dinb(n37334), .dout(n37393));
  jnot g19371(.din(n37177), .dout(n37394));
  jor  g19372(.dina(n37394), .dinb(n37393), .dout(n37395));
  jand g19373(.dina(n37395), .dinb(n37333), .dout(n37396));
  jnot g19374(.din(n37180), .dout(n37397));
  jor  g19375(.dina(n37397), .dinb(n37396), .dout(n37398));
  jand g19376(.dina(n37398), .dinb(n37332), .dout(n37399));
  jnot g19377(.din(n37183), .dout(n37400));
  jor  g19378(.dina(n37400), .dinb(n37399), .dout(n37401));
  jand g19379(.dina(n37401), .dinb(n37331), .dout(n37402));
  jnot g19380(.din(n37186), .dout(n37403));
  jor  g19381(.dina(n37403), .dinb(n37402), .dout(n37404));
  jand g19382(.dina(n37404), .dinb(n37330), .dout(n37405));
  jnot g19383(.din(n37189), .dout(n37406));
  jor  g19384(.dina(n37406), .dinb(n37405), .dout(n37407));
  jand g19385(.dina(n37407), .dinb(n37329), .dout(n37408));
  jnot g19386(.din(n37192), .dout(n37409));
  jor  g19387(.dina(n37409), .dinb(n37408), .dout(n37410));
  jand g19388(.dina(n37410), .dinb(n37328), .dout(n37411));
  jnot g19389(.din(n37195), .dout(n37412));
  jor  g19390(.dina(n37412), .dinb(n37411), .dout(n37413));
  jand g19391(.dina(n37413), .dinb(n37327), .dout(n37414));
  jnot g19392(.din(n37198), .dout(n37415));
  jor  g19393(.dina(n37415), .dinb(n37414), .dout(n37416));
  jand g19394(.dina(n37416), .dinb(n37326), .dout(n37417));
  jnot g19395(.din(n37201), .dout(n37418));
  jor  g19396(.dina(n37418), .dinb(n37417), .dout(n37419));
  jand g19397(.dina(n37419), .dinb(n37325), .dout(n37420));
  jnot g19398(.din(n37204), .dout(n37421));
  jor  g19399(.dina(n37421), .dinb(n37420), .dout(n37422));
  jand g19400(.dina(n37422), .dinb(n37324), .dout(n37423));
  jnot g19401(.din(n37207), .dout(n37424));
  jor  g19402(.dina(n37424), .dinb(n37423), .dout(n37425));
  jand g19403(.dina(n37425), .dinb(n37323), .dout(n37426));
  jnot g19404(.din(n37210), .dout(n37427));
  jor  g19405(.dina(n37427), .dinb(n37426), .dout(n37428));
  jand g19406(.dina(n37428), .dinb(n37322), .dout(n37429));
  jnot g19407(.din(n37213), .dout(n37430));
  jor  g19408(.dina(n37430), .dinb(n37429), .dout(n37431));
  jand g19409(.dina(n37431), .dinb(n37321), .dout(n37432));
  jnot g19410(.din(n37216), .dout(n37433));
  jor  g19411(.dina(n37433), .dinb(n37432), .dout(n37434));
  jand g19412(.dina(n37434), .dinb(n37320), .dout(n37435));
  jnot g19413(.din(n37219), .dout(n37436));
  jor  g19414(.dina(n37436), .dinb(n37435), .dout(n37437));
  jand g19415(.dina(n37437), .dinb(n37319), .dout(n37438));
  jnot g19416(.din(n37222), .dout(n37439));
  jor  g19417(.dina(n37439), .dinb(n37438), .dout(n37440));
  jand g19418(.dina(n37440), .dinb(n37318), .dout(n37441));
  jnot g19419(.din(n37225), .dout(n37442));
  jor  g19420(.dina(n37442), .dinb(n37441), .dout(n37443));
  jand g19421(.dina(n37443), .dinb(n37317), .dout(n37444));
  jnot g19422(.din(n37228), .dout(n37445));
  jor  g19423(.dina(n37445), .dinb(n37444), .dout(n37446));
  jand g19424(.dina(n37446), .dinb(n37316), .dout(n37447));
  jnot g19425(.din(n37231), .dout(n37448));
  jor  g19426(.dina(n37448), .dinb(n37447), .dout(n37449));
  jand g19427(.dina(n37449), .dinb(n37315), .dout(n37450));
  jnot g19428(.din(n37234), .dout(n37451));
  jor  g19429(.dina(n37451), .dinb(n37450), .dout(n37452));
  jand g19430(.dina(n37452), .dinb(n37314), .dout(n37453));
  jnot g19431(.din(n37237), .dout(n37454));
  jor  g19432(.dina(n37454), .dinb(n37453), .dout(n37455));
  jand g19433(.dina(n37455), .dinb(n37313), .dout(n37456));
  jnot g19434(.din(n37240), .dout(n37457));
  jor  g19435(.dina(n37457), .dinb(n37456), .dout(n37458));
  jand g19436(.dina(n37458), .dinb(n37312), .dout(n37459));
  jnot g19437(.din(n37243), .dout(n37460));
  jor  g19438(.dina(n37460), .dinb(n37459), .dout(n37461));
  jand g19439(.dina(n37461), .dinb(n37311), .dout(n37462));
  jnot g19440(.din(n37246), .dout(n37463));
  jor  g19441(.dina(n37463), .dinb(n37462), .dout(n37464));
  jand g19442(.dina(n37464), .dinb(n37310), .dout(n37465));
  jnot g19443(.din(n37249), .dout(n37466));
  jor  g19444(.dina(n37466), .dinb(n37465), .dout(n37467));
  jand g19445(.dina(n37467), .dinb(n37309), .dout(n37468));
  jnot g19446(.din(n37252), .dout(n37469));
  jor  g19447(.dina(n37469), .dinb(n37468), .dout(n37470));
  jand g19448(.dina(n37470), .dinb(n37308), .dout(n37471));
  jnot g19449(.din(n37255), .dout(n37472));
  jor  g19450(.dina(n37472), .dinb(n37471), .dout(n37473));
  jand g19451(.dina(n37473), .dinb(n37307), .dout(n37474));
  jnot g19452(.din(n37258), .dout(n37475));
  jor  g19453(.dina(n37475), .dinb(n37474), .dout(n37476));
  jand g19454(.dina(n37476), .dinb(n37306), .dout(n37477));
  jnot g19455(.din(n37261), .dout(n37478));
  jor  g19456(.dina(n37478), .dinb(n37477), .dout(n37479));
  jand g19457(.dina(n37479), .dinb(n37305), .dout(n37480));
  jnot g19458(.din(n37264), .dout(n37481));
  jor  g19459(.dina(n37481), .dinb(n37480), .dout(n37482));
  jand g19460(.dina(n37482), .dinb(n37304), .dout(n37483));
  jnot g19461(.din(n37267), .dout(n37484));
  jor  g19462(.dina(n37484), .dinb(n37483), .dout(n37485));
  jand g19463(.dina(n37485), .dinb(n37303), .dout(n37486));
  jnot g19464(.din(n37270), .dout(n37487));
  jor  g19465(.dina(n37487), .dinb(n37486), .dout(n37488));
  jand g19466(.dina(n37488), .dinb(n37302), .dout(n37489));
  jnot g19467(.din(n37273), .dout(n37490));
  jor  g19468(.dina(n37490), .dinb(n37489), .dout(n37491));
  jand g19469(.dina(n37491), .dinb(n37301), .dout(n37492));
  jnot g19470(.din(n37276), .dout(n37493));
  jor  g19471(.dina(n37493), .dinb(n37492), .dout(n37494));
  jand g19472(.dina(n37494), .dinb(n37300), .dout(n37495));
  jnot g19473(.din(n37279), .dout(n37496));
  jor  g19474(.dina(n37496), .dinb(n37495), .dout(n37497));
  jand g19475(.dina(n37497), .dinb(n37299), .dout(n37498));
  jnot g19476(.din(n37282), .dout(n37499));
  jor  g19477(.dina(n37499), .dinb(n37498), .dout(n37500));
  jand g19478(.dina(n37500), .dinb(n37298), .dout(n37501));
  jnot g19479(.din(n37285), .dout(n37502));
  jor  g19480(.dina(n37502), .dinb(n37501), .dout(n37503));
  jand g19481(.dina(n37503), .dinb(n37297), .dout(n37504));
  jnot g19482(.din(n37288), .dout(n37505));
  jor  g19483(.dina(n37505), .dinb(n37504), .dout(n37506));
  jand g19484(.dina(n37506), .dinb(n37296), .dout(n37507));
  jnot g19485(.din(n37291), .dout(n37508));
  jor  g19486(.dina(n37508), .dinb(n37507), .dout(n37509));
  jand g19487(.dina(n37509), .dinb(n37295), .dout(n37510));
  jand g19488(.dina(n37510), .dinb(b55 ), .dout(n37511));
  jor  g19489(.dina(n37511), .dinb(n14612), .dout(n37512));
  jor  g19490(.dina(n37512), .dinb(n37294), .dout(n37513));
  jand g19491(.dina(n37513), .dinb(n36856), .dout(n37514));
  jnot g19492(.din(n37514), .dout(n37515));
  jxor g19493(.dina(n36856), .dinb(b55 ), .dout(n37516));
  jor  g19494(.dina(n37516), .dinb(n14612), .dout(n37517));
  jor  g19495(.dina(n37517), .dinb(n37510), .dout(n37518));
  jand g19496(.dina(n36856), .dinb(n14054), .dout(n37519));
  jnot g19497(.din(n37519), .dout(n37520));
  jand g19498(.dina(n37520), .dinb(n37518), .dout(n37521));
  jand g19499(.dina(n37521), .dinb(n36864), .dout(n37522));
  jnot g19500(.din(n37517), .dout(n37523));
  jand g19501(.dina(n37523), .dinb(n37293), .dout(n37524));
  jor  g19502(.dina(n37519), .dinb(n37524), .dout(n37525));
  jxor g19503(.dina(n37291), .dinb(n37290), .dout(n37526));
  jand g19504(.dina(n37526), .dinb(n37525), .dout(n37527));
  jor  g19505(.dina(n37527), .dinb(n37522), .dout(n37528));
  jand g19506(.dina(n37528), .dinb(n377), .dout(n37529));
  jnot g19507(.din(n37529), .dout(n37530));
  jand g19508(.dina(n37521), .dinb(n36869), .dout(n37531));
  jxor g19509(.dina(n37288), .dinb(n37287), .dout(n37532));
  jand g19510(.dina(n37532), .dinb(n37525), .dout(n37533));
  jor  g19511(.dina(n37533), .dinb(n37531), .dout(n37534));
  jand g19512(.dina(n37534), .dinb(n376), .dout(n37535));
  jnot g19513(.din(n37535), .dout(n37536));
  jand g19514(.dina(n37521), .dinb(n36874), .dout(n37537));
  jxor g19515(.dina(n37285), .dinb(n37284), .dout(n37538));
  jand g19516(.dina(n37538), .dinb(n37525), .dout(n37539));
  jor  g19517(.dina(n37539), .dinb(n37537), .dout(n37540));
  jand g19518(.dina(n37540), .dinb(n374), .dout(n37541));
  jnot g19519(.din(n37541), .dout(n37542));
  jand g19520(.dina(n37521), .dinb(n36879), .dout(n37543));
  jxor g19521(.dina(n37282), .dinb(n37281), .dout(n37544));
  jand g19522(.dina(n37544), .dinb(n37525), .dout(n37545));
  jor  g19523(.dina(n37545), .dinb(n37543), .dout(n37546));
  jand g19524(.dina(n37546), .dinb(n384), .dout(n37547));
  jnot g19525(.din(n37547), .dout(n37548));
  jand g19526(.dina(n37521), .dinb(n36884), .dout(n37549));
  jxor g19527(.dina(n37279), .dinb(n37278), .dout(n37550));
  jand g19528(.dina(n37550), .dinb(n37525), .dout(n37551));
  jor  g19529(.dina(n37551), .dinb(n37549), .dout(n37552));
  jand g19530(.dina(n37552), .dinb(n12214), .dout(n37553));
  jnot g19531(.din(n37553), .dout(n37554));
  jand g19532(.dina(n37521), .dinb(n36889), .dout(n37555));
  jxor g19533(.dina(n37276), .dinb(n37275), .dout(n37556));
  jand g19534(.dina(n37556), .dinb(n37525), .dout(n37557));
  jor  g19535(.dina(n37557), .dinb(n37555), .dout(n37558));
  jand g19536(.dina(n37558), .dinb(n12211), .dout(n37559));
  jnot g19537(.din(n37559), .dout(n37560));
  jand g19538(.dina(n37521), .dinb(n36894), .dout(n37561));
  jxor g19539(.dina(n37273), .dinb(n37272), .dout(n37562));
  jand g19540(.dina(n37562), .dinb(n37525), .dout(n37563));
  jor  g19541(.dina(n37563), .dinb(n37561), .dout(n37564));
  jand g19542(.dina(n37564), .dinb(n383), .dout(n37565));
  jnot g19543(.din(n37565), .dout(n37566));
  jand g19544(.dina(n37521), .dinb(n36899), .dout(n37567));
  jxor g19545(.dina(n37270), .dinb(n37269), .dout(n37568));
  jand g19546(.dina(n37568), .dinb(n37525), .dout(n37569));
  jor  g19547(.dina(n37569), .dinb(n37567), .dout(n37570));
  jand g19548(.dina(n37570), .dinb(n396), .dout(n37571));
  jnot g19549(.din(n37571), .dout(n37572));
  jand g19550(.dina(n37521), .dinb(n36904), .dout(n37573));
  jxor g19551(.dina(n37267), .dinb(n37266), .dout(n37574));
  jand g19552(.dina(n37574), .dinb(n37525), .dout(n37575));
  jor  g19553(.dina(n37575), .dinb(n37573), .dout(n37576));
  jand g19554(.dina(n37576), .dinb(n510), .dout(n37577));
  jnot g19555(.din(n37577), .dout(n37578));
  jand g19556(.dina(n37521), .dinb(n36909), .dout(n37579));
  jxor g19557(.dina(n37264), .dinb(n37263), .dout(n37580));
  jand g19558(.dina(n37580), .dinb(n37525), .dout(n37581));
  jor  g19559(.dina(n37581), .dinb(n37579), .dout(n37582));
  jand g19560(.dina(n37582), .dinb(n514), .dout(n37583));
  jnot g19561(.din(n37583), .dout(n37584));
  jand g19562(.dina(n37521), .dinb(n36914), .dout(n37585));
  jxor g19563(.dina(n37261), .dinb(n37260), .dout(n37586));
  jand g19564(.dina(n37586), .dinb(n37525), .dout(n37587));
  jor  g19565(.dina(n37587), .dinb(n37585), .dout(n37588));
  jand g19566(.dina(n37588), .dinb(n513), .dout(n37589));
  jnot g19567(.din(n37589), .dout(n37590));
  jand g19568(.dina(n37521), .dinb(n36919), .dout(n37591));
  jxor g19569(.dina(n37258), .dinb(n37257), .dout(n37592));
  jand g19570(.dina(n37592), .dinb(n37525), .dout(n37593));
  jor  g19571(.dina(n37593), .dinb(n37591), .dout(n37594));
  jand g19572(.dina(n37594), .dinb(n397), .dout(n37595));
  jnot g19573(.din(n37595), .dout(n37596));
  jand g19574(.dina(n37521), .dinb(n36924), .dout(n37597));
  jxor g19575(.dina(n37255), .dinb(n37254), .dout(n37598));
  jand g19576(.dina(n37598), .dinb(n37525), .dout(n37599));
  jor  g19577(.dina(n37599), .dinb(n37597), .dout(n37600));
  jand g19578(.dina(n37600), .dinb(n282), .dout(n37601));
  jnot g19579(.din(n37601), .dout(n37602));
  jand g19580(.dina(n37521), .dinb(n36929), .dout(n37603));
  jxor g19581(.dina(n37252), .dinb(n37251), .dout(n37604));
  jand g19582(.dina(n37604), .dinb(n37525), .dout(n37605));
  jor  g19583(.dina(n37605), .dinb(n37603), .dout(n37606));
  jand g19584(.dina(n37606), .dinb(n281), .dout(n37607));
  jnot g19585(.din(n37607), .dout(n37608));
  jand g19586(.dina(n37521), .dinb(n36934), .dout(n37609));
  jxor g19587(.dina(n37249), .dinb(n37248), .dout(n37610));
  jand g19588(.dina(n37610), .dinb(n37525), .dout(n37611));
  jor  g19589(.dina(n37611), .dinb(n37609), .dout(n37612));
  jand g19590(.dina(n37612), .dinb(n285), .dout(n37613));
  jnot g19591(.din(n37613), .dout(n37614));
  jand g19592(.dina(n37521), .dinb(n36939), .dout(n37615));
  jxor g19593(.dina(n37246), .dinb(n37245), .dout(n37616));
  jand g19594(.dina(n37616), .dinb(n37525), .dout(n37617));
  jor  g19595(.dina(n37617), .dinb(n37615), .dout(n37618));
  jand g19596(.dina(n37618), .dinb(n284), .dout(n37619));
  jnot g19597(.din(n37619), .dout(n37620));
  jand g19598(.dina(n37521), .dinb(n36944), .dout(n37621));
  jxor g19599(.dina(n37243), .dinb(n37242), .dout(n37622));
  jand g19600(.dina(n37622), .dinb(n37525), .dout(n37623));
  jor  g19601(.dina(n37623), .dinb(n37621), .dout(n37624));
  jand g19602(.dina(n37624), .dinb(n291), .dout(n37625));
  jnot g19603(.din(n37625), .dout(n37626));
  jand g19604(.dina(n37521), .dinb(n36949), .dout(n37627));
  jxor g19605(.dina(n37240), .dinb(n37239), .dout(n37628));
  jand g19606(.dina(n37628), .dinb(n37525), .dout(n37629));
  jor  g19607(.dina(n37629), .dinb(n37627), .dout(n37630));
  jand g19608(.dina(n37630), .dinb(n290), .dout(n37631));
  jnot g19609(.din(n37631), .dout(n37632));
  jand g19610(.dina(n37521), .dinb(n36954), .dout(n37633));
  jxor g19611(.dina(n37237), .dinb(n37236), .dout(n37634));
  jand g19612(.dina(n37634), .dinb(n37525), .dout(n37635));
  jor  g19613(.dina(n37635), .dinb(n37633), .dout(n37636));
  jand g19614(.dina(n37636), .dinb(n294), .dout(n37637));
  jnot g19615(.din(n37637), .dout(n37638));
  jand g19616(.dina(n37521), .dinb(n36959), .dout(n37639));
  jxor g19617(.dina(n37234), .dinb(n37233), .dout(n37640));
  jand g19618(.dina(n37640), .dinb(n37525), .dout(n37641));
  jor  g19619(.dina(n37641), .dinb(n37639), .dout(n37642));
  jand g19620(.dina(n37642), .dinb(n293), .dout(n37643));
  jnot g19621(.din(n37643), .dout(n37644));
  jand g19622(.dina(n37521), .dinb(n36964), .dout(n37645));
  jxor g19623(.dina(n37231), .dinb(n37230), .dout(n37646));
  jand g19624(.dina(n37646), .dinb(n37525), .dout(n37647));
  jor  g19625(.dina(n37647), .dinb(n37645), .dout(n37648));
  jand g19626(.dina(n37648), .dinb(n301), .dout(n37649));
  jnot g19627(.din(n37649), .dout(n37650));
  jand g19628(.dina(n37521), .dinb(n36969), .dout(n37651));
  jxor g19629(.dina(n37228), .dinb(n37227), .dout(n37652));
  jand g19630(.dina(n37652), .dinb(n37525), .dout(n37653));
  jor  g19631(.dina(n37653), .dinb(n37651), .dout(n37654));
  jand g19632(.dina(n37654), .dinb(n298), .dout(n37655));
  jnot g19633(.din(n37655), .dout(n37656));
  jand g19634(.dina(n37521), .dinb(n36974), .dout(n37657));
  jxor g19635(.dina(n37225), .dinb(n37224), .dout(n37658));
  jand g19636(.dina(n37658), .dinb(n37525), .dout(n37659));
  jor  g19637(.dina(n37659), .dinb(n37657), .dout(n37660));
  jand g19638(.dina(n37660), .dinb(n297), .dout(n37661));
  jnot g19639(.din(n37661), .dout(n37662));
  jand g19640(.dina(n37521), .dinb(n36979), .dout(n37663));
  jxor g19641(.dina(n37222), .dinb(n37221), .dout(n37664));
  jand g19642(.dina(n37664), .dinb(n37525), .dout(n37665));
  jor  g19643(.dina(n37665), .dinb(n37663), .dout(n37666));
  jand g19644(.dina(n37666), .dinb(n300), .dout(n37667));
  jnot g19645(.din(n37667), .dout(n37668));
  jand g19646(.dina(n37521), .dinb(n36984), .dout(n37669));
  jxor g19647(.dina(n37219), .dinb(n37218), .dout(n37670));
  jand g19648(.dina(n37670), .dinb(n37525), .dout(n37671));
  jor  g19649(.dina(n37671), .dinb(n37669), .dout(n37672));
  jand g19650(.dina(n37672), .dinb(n424), .dout(n37673));
  jnot g19651(.din(n37673), .dout(n37674));
  jand g19652(.dina(n37521), .dinb(n36989), .dout(n37675));
  jxor g19653(.dina(n37216), .dinb(n37215), .dout(n37676));
  jand g19654(.dina(n37676), .dinb(n37525), .dout(n37677));
  jor  g19655(.dina(n37677), .dinb(n37675), .dout(n37678));
  jand g19656(.dina(n37678), .dinb(n427), .dout(n37679));
  jnot g19657(.din(n37679), .dout(n37680));
  jand g19658(.dina(n37521), .dinb(n36994), .dout(n37681));
  jxor g19659(.dina(n37213), .dinb(n37212), .dout(n37682));
  jand g19660(.dina(n37682), .dinb(n37525), .dout(n37683));
  jor  g19661(.dina(n37683), .dinb(n37681), .dout(n37684));
  jand g19662(.dina(n37684), .dinb(n426), .dout(n37685));
  jnot g19663(.din(n37685), .dout(n37686));
  jand g19664(.dina(n37521), .dinb(n36999), .dout(n37687));
  jxor g19665(.dina(n37210), .dinb(n37209), .dout(n37688));
  jand g19666(.dina(n37688), .dinb(n37525), .dout(n37689));
  jor  g19667(.dina(n37689), .dinb(n37687), .dout(n37690));
  jand g19668(.dina(n37690), .dinb(n410), .dout(n37691));
  jnot g19669(.din(n37691), .dout(n37692));
  jand g19670(.dina(n37521), .dinb(n37004), .dout(n37693));
  jxor g19671(.dina(n37207), .dinb(n37206), .dout(n37694));
  jand g19672(.dina(n37694), .dinb(n37525), .dout(n37695));
  jor  g19673(.dina(n37695), .dinb(n37693), .dout(n37696));
  jand g19674(.dina(n37696), .dinb(n409), .dout(n37697));
  jnot g19675(.din(n37697), .dout(n37698));
  jand g19676(.dina(n37521), .dinb(n37009), .dout(n37699));
  jxor g19677(.dina(n37204), .dinb(n37203), .dout(n37700));
  jand g19678(.dina(n37700), .dinb(n37525), .dout(n37701));
  jor  g19679(.dina(n37701), .dinb(n37699), .dout(n37702));
  jand g19680(.dina(n37702), .dinb(n413), .dout(n37703));
  jnot g19681(.din(n37703), .dout(n37704));
  jand g19682(.dina(n37521), .dinb(n37014), .dout(n37705));
  jxor g19683(.dina(n37201), .dinb(n37200), .dout(n37706));
  jand g19684(.dina(n37706), .dinb(n37525), .dout(n37707));
  jor  g19685(.dina(n37707), .dinb(n37705), .dout(n37708));
  jand g19686(.dina(n37708), .dinb(n412), .dout(n37709));
  jnot g19687(.din(n37709), .dout(n37710));
  jand g19688(.dina(n37521), .dinb(n37019), .dout(n37711));
  jxor g19689(.dina(n37198), .dinb(n37197), .dout(n37712));
  jand g19690(.dina(n37712), .dinb(n37525), .dout(n37713));
  jor  g19691(.dina(n37713), .dinb(n37711), .dout(n37714));
  jand g19692(.dina(n37714), .dinb(n406), .dout(n37715));
  jnot g19693(.din(n37715), .dout(n37716));
  jand g19694(.dina(n37521), .dinb(n37024), .dout(n37717));
  jxor g19695(.dina(n37195), .dinb(n37194), .dout(n37718));
  jand g19696(.dina(n37718), .dinb(n37525), .dout(n37719));
  jor  g19697(.dina(n37719), .dinb(n37717), .dout(n37720));
  jand g19698(.dina(n37720), .dinb(n405), .dout(n37721));
  jnot g19699(.din(n37721), .dout(n37722));
  jand g19700(.dina(n37521), .dinb(n37029), .dout(n37723));
  jxor g19701(.dina(n37192), .dinb(n37191), .dout(n37724));
  jand g19702(.dina(n37724), .dinb(n37525), .dout(n37725));
  jor  g19703(.dina(n37725), .dinb(n37723), .dout(n37726));
  jand g19704(.dina(n37726), .dinb(n2714), .dout(n37727));
  jnot g19705(.din(n37727), .dout(n37728));
  jand g19706(.dina(n37521), .dinb(n37034), .dout(n37729));
  jxor g19707(.dina(n37189), .dinb(n37188), .dout(n37730));
  jand g19708(.dina(n37730), .dinb(n37525), .dout(n37731));
  jor  g19709(.dina(n37731), .dinb(n37729), .dout(n37732));
  jand g19710(.dina(n37732), .dinb(n2547), .dout(n37733));
  jnot g19711(.din(n37733), .dout(n37734));
  jand g19712(.dina(n37521), .dinb(n37039), .dout(n37735));
  jxor g19713(.dina(n37186), .dinb(n37185), .dout(n37736));
  jand g19714(.dina(n37736), .dinb(n37525), .dout(n37737));
  jor  g19715(.dina(n37737), .dinb(n37735), .dout(n37738));
  jand g19716(.dina(n37738), .dinb(n417), .dout(n37739));
  jnot g19717(.din(n37739), .dout(n37740));
  jand g19718(.dina(n37521), .dinb(n37044), .dout(n37741));
  jxor g19719(.dina(n37183), .dinb(n37182), .dout(n37742));
  jand g19720(.dina(n37742), .dinb(n37525), .dout(n37743));
  jor  g19721(.dina(n37743), .dinb(n37741), .dout(n37744));
  jand g19722(.dina(n37744), .dinb(n416), .dout(n37745));
  jnot g19723(.din(n37745), .dout(n37746));
  jand g19724(.dina(n37521), .dinb(n37049), .dout(n37747));
  jxor g19725(.dina(n37180), .dinb(n37179), .dout(n37748));
  jand g19726(.dina(n37748), .dinb(n37525), .dout(n37749));
  jor  g19727(.dina(n37749), .dinb(n37747), .dout(n37750));
  jand g19728(.dina(n37750), .dinb(n422), .dout(n37751));
  jnot g19729(.din(n37751), .dout(n37752));
  jand g19730(.dina(n37521), .dinb(n37054), .dout(n37753));
  jxor g19731(.dina(n37177), .dinb(n37176), .dout(n37754));
  jand g19732(.dina(n37754), .dinb(n37525), .dout(n37755));
  jor  g19733(.dina(n37755), .dinb(n37753), .dout(n37756));
  jand g19734(.dina(n37756), .dinb(n421), .dout(n37757));
  jnot g19735(.din(n37757), .dout(n37758));
  jand g19736(.dina(n37521), .dinb(n37059), .dout(n37759));
  jxor g19737(.dina(n37174), .dinb(n37173), .dout(n37760));
  jand g19738(.dina(n37760), .dinb(n37525), .dout(n37761));
  jor  g19739(.dina(n37761), .dinb(n37759), .dout(n37762));
  jand g19740(.dina(n37762), .dinb(n433), .dout(n37763));
  jnot g19741(.din(n37763), .dout(n37764));
  jand g19742(.dina(n37521), .dinb(n37064), .dout(n37765));
  jxor g19743(.dina(n37171), .dinb(n37170), .dout(n37766));
  jand g19744(.dina(n37766), .dinb(n37525), .dout(n37767));
  jor  g19745(.dina(n37767), .dinb(n37765), .dout(n37768));
  jand g19746(.dina(n37768), .dinb(n432), .dout(n37769));
  jnot g19747(.din(n37769), .dout(n37770));
  jand g19748(.dina(n37521), .dinb(n37069), .dout(n37771));
  jxor g19749(.dina(n37168), .dinb(n37167), .dout(n37772));
  jand g19750(.dina(n37772), .dinb(n37525), .dout(n37773));
  jor  g19751(.dina(n37773), .dinb(n37771), .dout(n37774));
  jand g19752(.dina(n37774), .dinb(n436), .dout(n37775));
  jnot g19753(.din(n37775), .dout(n37776));
  jand g19754(.dina(n37521), .dinb(n37074), .dout(n37777));
  jxor g19755(.dina(n37165), .dinb(n37164), .dout(n37778));
  jand g19756(.dina(n37778), .dinb(n37525), .dout(n37779));
  jor  g19757(.dina(n37779), .dinb(n37777), .dout(n37780));
  jand g19758(.dina(n37780), .dinb(n435), .dout(n37781));
  jnot g19759(.din(n37781), .dout(n37782));
  jand g19760(.dina(n37521), .dinb(n37079), .dout(n37783));
  jxor g19761(.dina(n37162), .dinb(n37161), .dout(n37784));
  jand g19762(.dina(n37784), .dinb(n37525), .dout(n37785));
  jor  g19763(.dina(n37785), .dinb(n37783), .dout(n37786));
  jand g19764(.dina(n37786), .dinb(n440), .dout(n37787));
  jnot g19765(.din(n37787), .dout(n37788));
  jand g19766(.dina(n37521), .dinb(n37084), .dout(n37789));
  jxor g19767(.dina(n37159), .dinb(n37158), .dout(n37790));
  jand g19768(.dina(n37790), .dinb(n37525), .dout(n37791));
  jor  g19769(.dina(n37791), .dinb(n37789), .dout(n37792));
  jand g19770(.dina(n37792), .dinb(n439), .dout(n37793));
  jnot g19771(.din(n37793), .dout(n37794));
  jand g19772(.dina(n37521), .dinb(n37089), .dout(n37795));
  jxor g19773(.dina(n37156), .dinb(n37155), .dout(n37796));
  jand g19774(.dina(n37796), .dinb(n37525), .dout(n37797));
  jor  g19775(.dina(n37797), .dinb(n37795), .dout(n37798));
  jand g19776(.dina(n37798), .dinb(n325), .dout(n37799));
  jnot g19777(.din(n37799), .dout(n37800));
  jand g19778(.dina(n37521), .dinb(n37094), .dout(n37801));
  jxor g19779(.dina(n37153), .dinb(n37152), .dout(n37802));
  jand g19780(.dina(n37802), .dinb(n37525), .dout(n37803));
  jor  g19781(.dina(n37803), .dinb(n37801), .dout(n37804));
  jand g19782(.dina(n37804), .dinb(n324), .dout(n37805));
  jnot g19783(.din(n37805), .dout(n37806));
  jand g19784(.dina(n37521), .dinb(n37099), .dout(n37807));
  jxor g19785(.dina(n37150), .dinb(n37149), .dout(n37808));
  jand g19786(.dina(n37808), .dinb(n37525), .dout(n37809));
  jor  g19787(.dina(n37809), .dinb(n37807), .dout(n37810));
  jand g19788(.dina(n37810), .dinb(n323), .dout(n37811));
  jnot g19789(.din(n37811), .dout(n37812));
  jand g19790(.dina(n37521), .dinb(n37104), .dout(n37813));
  jxor g19791(.dina(n37147), .dinb(n37146), .dout(n37814));
  jand g19792(.dina(n37814), .dinb(n37525), .dout(n37815));
  jor  g19793(.dina(n37815), .dinb(n37813), .dout(n37816));
  jand g19794(.dina(n37816), .dinb(n335), .dout(n37817));
  jnot g19795(.din(n37817), .dout(n37818));
  jand g19796(.dina(n37521), .dinb(n37109), .dout(n37819));
  jxor g19797(.dina(n37144), .dinb(n37143), .dout(n37820));
  jand g19798(.dina(n37820), .dinb(n37525), .dout(n37821));
  jor  g19799(.dina(n37821), .dinb(n37819), .dout(n37822));
  jand g19800(.dina(n37822), .dinb(n334), .dout(n37823));
  jnot g19801(.din(n37823), .dout(n37824));
  jand g19802(.dina(n37521), .dinb(n37114), .dout(n37825));
  jxor g19803(.dina(n37141), .dinb(n37140), .dout(n37826));
  jand g19804(.dina(n37826), .dinb(n37525), .dout(n37827));
  jor  g19805(.dina(n37827), .dinb(n37825), .dout(n37828));
  jand g19806(.dina(n37828), .dinb(n338), .dout(n37829));
  jnot g19807(.din(n37829), .dout(n37830));
  jand g19808(.dina(n37521), .dinb(n37119), .dout(n37831));
  jxor g19809(.dina(n37138), .dinb(n37137), .dout(n37832));
  jand g19810(.dina(n37832), .dinb(n37525), .dout(n37833));
  jor  g19811(.dina(n37833), .dinb(n37831), .dout(n37834));
  jand g19812(.dina(n37834), .dinb(n337), .dout(n37835));
  jnot g19813(.din(n37835), .dout(n37836));
  jand g19814(.dina(n37521), .dinb(n37126), .dout(n37837));
  jxor g19815(.dina(n37135), .dinb(n37134), .dout(n37838));
  jand g19816(.dina(n37838), .dinb(n37525), .dout(n37839));
  jor  g19817(.dina(n37839), .dinb(n37837), .dout(n37840));
  jand g19818(.dina(n37840), .dinb(n344), .dout(n37841));
  jnot g19819(.din(n37841), .dout(n37842));
  jand g19820(.dina(n37521), .dinb(n37129), .dout(n37843));
  jxor g19821(.dina(n37132), .dinb(n14449), .dout(n37844));
  jand g19822(.dina(n37844), .dinb(n37525), .dout(n37845));
  jor  g19823(.dina(n37845), .dinb(n37843), .dout(n37846));
  jand g19824(.dina(n37846), .dinb(n348), .dout(n37847));
  jnot g19825(.din(n37847), .dout(n37848));
  jor  g19826(.dina(n37521), .dinb(n18364), .dout(n37849));
  jand g19827(.dina(n37849), .dinb(a8 ), .dout(n37850));
  jor  g19828(.dina(n37521), .dinb(n14449), .dout(n37851));
  jnot g19829(.din(n37851), .dout(n37852));
  jor  g19830(.dina(n37852), .dinb(n37850), .dout(n37853));
  jand g19831(.dina(n37853), .dinb(n258), .dout(n37854));
  jnot g19832(.din(n37854), .dout(n37855));
  jand g19833(.dina(n37525), .dinb(b0 ), .dout(n37856));
  jor  g19834(.dina(n37856), .dinb(n14447), .dout(n37857));
  jand g19835(.dina(n37851), .dinb(n37857), .dout(n37858));
  jxor g19836(.dina(n37858), .dinb(n258), .dout(n37859));
  jor  g19837(.dina(n37859), .dinb(n14904), .dout(n37860));
  jand g19838(.dina(n37860), .dinb(n37855), .dout(n37861));
  jxor g19839(.dina(n37846), .dinb(n348), .dout(n37862));
  jnot g19840(.din(n37862), .dout(n37863));
  jor  g19841(.dina(n37863), .dinb(n37861), .dout(n37864));
  jand g19842(.dina(n37864), .dinb(n37848), .dout(n37865));
  jxor g19843(.dina(n37840), .dinb(n344), .dout(n37866));
  jnot g19844(.din(n37866), .dout(n37867));
  jor  g19845(.dina(n37867), .dinb(n37865), .dout(n37868));
  jand g19846(.dina(n37868), .dinb(n37842), .dout(n37869));
  jxor g19847(.dina(n37834), .dinb(n337), .dout(n37870));
  jnot g19848(.din(n37870), .dout(n37871));
  jor  g19849(.dina(n37871), .dinb(n37869), .dout(n37872));
  jand g19850(.dina(n37872), .dinb(n37836), .dout(n37873));
  jxor g19851(.dina(n37828), .dinb(n338), .dout(n37874));
  jnot g19852(.din(n37874), .dout(n37875));
  jor  g19853(.dina(n37875), .dinb(n37873), .dout(n37876));
  jand g19854(.dina(n37876), .dinb(n37830), .dout(n37877));
  jxor g19855(.dina(n37822), .dinb(n334), .dout(n37878));
  jnot g19856(.din(n37878), .dout(n37879));
  jor  g19857(.dina(n37879), .dinb(n37877), .dout(n37880));
  jand g19858(.dina(n37880), .dinb(n37824), .dout(n37881));
  jxor g19859(.dina(n37816), .dinb(n335), .dout(n37882));
  jnot g19860(.din(n37882), .dout(n37883));
  jor  g19861(.dina(n37883), .dinb(n37881), .dout(n37884));
  jand g19862(.dina(n37884), .dinb(n37818), .dout(n37885));
  jxor g19863(.dina(n37810), .dinb(n323), .dout(n37886));
  jnot g19864(.din(n37886), .dout(n37887));
  jor  g19865(.dina(n37887), .dinb(n37885), .dout(n37888));
  jand g19866(.dina(n37888), .dinb(n37812), .dout(n37889));
  jxor g19867(.dina(n37804), .dinb(n324), .dout(n37890));
  jnot g19868(.din(n37890), .dout(n37891));
  jor  g19869(.dina(n37891), .dinb(n37889), .dout(n37892));
  jand g19870(.dina(n37892), .dinb(n37806), .dout(n37893));
  jxor g19871(.dina(n37798), .dinb(n325), .dout(n37894));
  jnot g19872(.din(n37894), .dout(n37895));
  jor  g19873(.dina(n37895), .dinb(n37893), .dout(n37896));
  jand g19874(.dina(n37896), .dinb(n37800), .dout(n37897));
  jxor g19875(.dina(n37792), .dinb(n439), .dout(n37898));
  jnot g19876(.din(n37898), .dout(n37899));
  jor  g19877(.dina(n37899), .dinb(n37897), .dout(n37900));
  jand g19878(.dina(n37900), .dinb(n37794), .dout(n37901));
  jxor g19879(.dina(n37786), .dinb(n440), .dout(n37902));
  jnot g19880(.din(n37902), .dout(n37903));
  jor  g19881(.dina(n37903), .dinb(n37901), .dout(n37904));
  jand g19882(.dina(n37904), .dinb(n37788), .dout(n37905));
  jxor g19883(.dina(n37780), .dinb(n435), .dout(n37906));
  jnot g19884(.din(n37906), .dout(n37907));
  jor  g19885(.dina(n37907), .dinb(n37905), .dout(n37908));
  jand g19886(.dina(n37908), .dinb(n37782), .dout(n37909));
  jxor g19887(.dina(n37774), .dinb(n436), .dout(n37910));
  jnot g19888(.din(n37910), .dout(n37911));
  jor  g19889(.dina(n37911), .dinb(n37909), .dout(n37912));
  jand g19890(.dina(n37912), .dinb(n37776), .dout(n37913));
  jxor g19891(.dina(n37768), .dinb(n432), .dout(n37914));
  jnot g19892(.din(n37914), .dout(n37915));
  jor  g19893(.dina(n37915), .dinb(n37913), .dout(n37916));
  jand g19894(.dina(n37916), .dinb(n37770), .dout(n37917));
  jxor g19895(.dina(n37762), .dinb(n433), .dout(n37918));
  jnot g19896(.din(n37918), .dout(n37919));
  jor  g19897(.dina(n37919), .dinb(n37917), .dout(n37920));
  jand g19898(.dina(n37920), .dinb(n37764), .dout(n37921));
  jxor g19899(.dina(n37756), .dinb(n421), .dout(n37922));
  jnot g19900(.din(n37922), .dout(n37923));
  jor  g19901(.dina(n37923), .dinb(n37921), .dout(n37924));
  jand g19902(.dina(n37924), .dinb(n37758), .dout(n37925));
  jxor g19903(.dina(n37750), .dinb(n422), .dout(n37926));
  jnot g19904(.din(n37926), .dout(n37927));
  jor  g19905(.dina(n37927), .dinb(n37925), .dout(n37928));
  jand g19906(.dina(n37928), .dinb(n37752), .dout(n37929));
  jxor g19907(.dina(n37744), .dinb(n416), .dout(n37930));
  jnot g19908(.din(n37930), .dout(n37931));
  jor  g19909(.dina(n37931), .dinb(n37929), .dout(n37932));
  jand g19910(.dina(n37932), .dinb(n37746), .dout(n37933));
  jxor g19911(.dina(n37738), .dinb(n417), .dout(n37934));
  jnot g19912(.din(n37934), .dout(n37935));
  jor  g19913(.dina(n37935), .dinb(n37933), .dout(n37936));
  jand g19914(.dina(n37936), .dinb(n37740), .dout(n37937));
  jxor g19915(.dina(n37732), .dinb(n2547), .dout(n37938));
  jnot g19916(.din(n37938), .dout(n37939));
  jor  g19917(.dina(n37939), .dinb(n37937), .dout(n37940));
  jand g19918(.dina(n37940), .dinb(n37734), .dout(n37941));
  jxor g19919(.dina(n37726), .dinb(n2714), .dout(n37942));
  jnot g19920(.din(n37942), .dout(n37943));
  jor  g19921(.dina(n37943), .dinb(n37941), .dout(n37944));
  jand g19922(.dina(n37944), .dinb(n37728), .dout(n37945));
  jxor g19923(.dina(n37720), .dinb(n405), .dout(n37946));
  jnot g19924(.din(n37946), .dout(n37947));
  jor  g19925(.dina(n37947), .dinb(n37945), .dout(n37948));
  jand g19926(.dina(n37948), .dinb(n37722), .dout(n37949));
  jxor g19927(.dina(n37714), .dinb(n406), .dout(n37950));
  jnot g19928(.din(n37950), .dout(n37951));
  jor  g19929(.dina(n37951), .dinb(n37949), .dout(n37952));
  jand g19930(.dina(n37952), .dinb(n37716), .dout(n37953));
  jxor g19931(.dina(n37708), .dinb(n412), .dout(n37954));
  jnot g19932(.din(n37954), .dout(n37955));
  jor  g19933(.dina(n37955), .dinb(n37953), .dout(n37956));
  jand g19934(.dina(n37956), .dinb(n37710), .dout(n37957));
  jxor g19935(.dina(n37702), .dinb(n413), .dout(n37958));
  jnot g19936(.din(n37958), .dout(n37959));
  jor  g19937(.dina(n37959), .dinb(n37957), .dout(n37960));
  jand g19938(.dina(n37960), .dinb(n37704), .dout(n37961));
  jxor g19939(.dina(n37696), .dinb(n409), .dout(n37962));
  jnot g19940(.din(n37962), .dout(n37963));
  jor  g19941(.dina(n37963), .dinb(n37961), .dout(n37964));
  jand g19942(.dina(n37964), .dinb(n37698), .dout(n37965));
  jxor g19943(.dina(n37690), .dinb(n410), .dout(n37966));
  jnot g19944(.din(n37966), .dout(n37967));
  jor  g19945(.dina(n37967), .dinb(n37965), .dout(n37968));
  jand g19946(.dina(n37968), .dinb(n37692), .dout(n37969));
  jxor g19947(.dina(n37684), .dinb(n426), .dout(n37970));
  jnot g19948(.din(n37970), .dout(n37971));
  jor  g19949(.dina(n37971), .dinb(n37969), .dout(n37972));
  jand g19950(.dina(n37972), .dinb(n37686), .dout(n37973));
  jxor g19951(.dina(n37678), .dinb(n427), .dout(n37974));
  jnot g19952(.din(n37974), .dout(n37975));
  jor  g19953(.dina(n37975), .dinb(n37973), .dout(n37976));
  jand g19954(.dina(n37976), .dinb(n37680), .dout(n37977));
  jxor g19955(.dina(n37672), .dinb(n424), .dout(n37978));
  jnot g19956(.din(n37978), .dout(n37979));
  jor  g19957(.dina(n37979), .dinb(n37977), .dout(n37980));
  jand g19958(.dina(n37980), .dinb(n37674), .dout(n37981));
  jxor g19959(.dina(n37666), .dinb(n300), .dout(n37982));
  jnot g19960(.din(n37982), .dout(n37983));
  jor  g19961(.dina(n37983), .dinb(n37981), .dout(n37984));
  jand g19962(.dina(n37984), .dinb(n37668), .dout(n37985));
  jxor g19963(.dina(n37660), .dinb(n297), .dout(n37986));
  jnot g19964(.din(n37986), .dout(n37987));
  jor  g19965(.dina(n37987), .dinb(n37985), .dout(n37988));
  jand g19966(.dina(n37988), .dinb(n37662), .dout(n37989));
  jxor g19967(.dina(n37654), .dinb(n298), .dout(n37990));
  jnot g19968(.din(n37990), .dout(n37991));
  jor  g19969(.dina(n37991), .dinb(n37989), .dout(n37992));
  jand g19970(.dina(n37992), .dinb(n37656), .dout(n37993));
  jxor g19971(.dina(n37648), .dinb(n301), .dout(n37994));
  jnot g19972(.din(n37994), .dout(n37995));
  jor  g19973(.dina(n37995), .dinb(n37993), .dout(n37996));
  jand g19974(.dina(n37996), .dinb(n37650), .dout(n37997));
  jxor g19975(.dina(n37642), .dinb(n293), .dout(n37998));
  jnot g19976(.din(n37998), .dout(n37999));
  jor  g19977(.dina(n37999), .dinb(n37997), .dout(n38000));
  jand g19978(.dina(n38000), .dinb(n37644), .dout(n38001));
  jxor g19979(.dina(n37636), .dinb(n294), .dout(n38002));
  jnot g19980(.din(n38002), .dout(n38003));
  jor  g19981(.dina(n38003), .dinb(n38001), .dout(n38004));
  jand g19982(.dina(n38004), .dinb(n37638), .dout(n38005));
  jxor g19983(.dina(n37630), .dinb(n290), .dout(n38006));
  jnot g19984(.din(n38006), .dout(n38007));
  jor  g19985(.dina(n38007), .dinb(n38005), .dout(n38008));
  jand g19986(.dina(n38008), .dinb(n37632), .dout(n38009));
  jxor g19987(.dina(n37624), .dinb(n291), .dout(n38010));
  jnot g19988(.din(n38010), .dout(n38011));
  jor  g19989(.dina(n38011), .dinb(n38009), .dout(n38012));
  jand g19990(.dina(n38012), .dinb(n37626), .dout(n38013));
  jxor g19991(.dina(n37618), .dinb(n284), .dout(n38014));
  jnot g19992(.din(n38014), .dout(n38015));
  jor  g19993(.dina(n38015), .dinb(n38013), .dout(n38016));
  jand g19994(.dina(n38016), .dinb(n37620), .dout(n38017));
  jxor g19995(.dina(n37612), .dinb(n285), .dout(n38018));
  jnot g19996(.din(n38018), .dout(n38019));
  jor  g19997(.dina(n38019), .dinb(n38017), .dout(n38020));
  jand g19998(.dina(n38020), .dinb(n37614), .dout(n38021));
  jxor g19999(.dina(n37606), .dinb(n281), .dout(n38022));
  jnot g20000(.din(n38022), .dout(n38023));
  jor  g20001(.dina(n38023), .dinb(n38021), .dout(n38024));
  jand g20002(.dina(n38024), .dinb(n37608), .dout(n38025));
  jxor g20003(.dina(n37600), .dinb(n282), .dout(n38026));
  jnot g20004(.din(n38026), .dout(n38027));
  jor  g20005(.dina(n38027), .dinb(n38025), .dout(n38028));
  jand g20006(.dina(n38028), .dinb(n37602), .dout(n38029));
  jxor g20007(.dina(n37594), .dinb(n397), .dout(n38030));
  jnot g20008(.din(n38030), .dout(n38031));
  jor  g20009(.dina(n38031), .dinb(n38029), .dout(n38032));
  jand g20010(.dina(n38032), .dinb(n37596), .dout(n38033));
  jxor g20011(.dina(n37588), .dinb(n513), .dout(n38034));
  jnot g20012(.din(n38034), .dout(n38035));
  jor  g20013(.dina(n38035), .dinb(n38033), .dout(n38036));
  jand g20014(.dina(n38036), .dinb(n37590), .dout(n38037));
  jxor g20015(.dina(n37582), .dinb(n514), .dout(n38038));
  jnot g20016(.din(n38038), .dout(n38039));
  jor  g20017(.dina(n38039), .dinb(n38037), .dout(n38040));
  jand g20018(.dina(n38040), .dinb(n37584), .dout(n38041));
  jxor g20019(.dina(n37576), .dinb(n510), .dout(n38042));
  jnot g20020(.din(n38042), .dout(n38043));
  jor  g20021(.dina(n38043), .dinb(n38041), .dout(n38044));
  jand g20022(.dina(n38044), .dinb(n37578), .dout(n38045));
  jxor g20023(.dina(n37570), .dinb(n396), .dout(n38046));
  jnot g20024(.din(n38046), .dout(n38047));
  jor  g20025(.dina(n38047), .dinb(n38045), .dout(n38048));
  jand g20026(.dina(n38048), .dinb(n37572), .dout(n38049));
  jxor g20027(.dina(n37564), .dinb(n383), .dout(n38050));
  jnot g20028(.din(n38050), .dout(n38051));
  jor  g20029(.dina(n38051), .dinb(n38049), .dout(n38052));
  jand g20030(.dina(n38052), .dinb(n37566), .dout(n38053));
  jxor g20031(.dina(n37558), .dinb(n12211), .dout(n38054));
  jnot g20032(.din(n38054), .dout(n38055));
  jor  g20033(.dina(n38055), .dinb(n38053), .dout(n38056));
  jand g20034(.dina(n38056), .dinb(n37560), .dout(n38057));
  jxor g20035(.dina(n37552), .dinb(n12214), .dout(n38058));
  jnot g20036(.din(n38058), .dout(n38059));
  jor  g20037(.dina(n38059), .dinb(n38057), .dout(n38060));
  jand g20038(.dina(n38060), .dinb(n37554), .dout(n38061));
  jxor g20039(.dina(n37546), .dinb(n384), .dout(n38062));
  jnot g20040(.din(n38062), .dout(n38063));
  jor  g20041(.dina(n38063), .dinb(n38061), .dout(n38064));
  jand g20042(.dina(n38064), .dinb(n37548), .dout(n38065));
  jxor g20043(.dina(n37540), .dinb(n374), .dout(n38066));
  jnot g20044(.din(n38066), .dout(n38067));
  jor  g20045(.dina(n38067), .dinb(n38065), .dout(n38068));
  jand g20046(.dina(n38068), .dinb(n37542), .dout(n38069));
  jxor g20047(.dina(n37534), .dinb(n376), .dout(n38070));
  jnot g20048(.din(n38070), .dout(n38071));
  jor  g20049(.dina(n38071), .dinb(n38069), .dout(n38072));
  jand g20050(.dina(n38072), .dinb(n37536), .dout(n38073));
  jxor g20051(.dina(n37528), .dinb(n377), .dout(n38074));
  jnot g20052(.din(n38074), .dout(n38075));
  jor  g20053(.dina(n38075), .dinb(n38073), .dout(n38076));
  jand g20054(.dina(n38076), .dinb(n37530), .dout(n38077));
  jand g20055(.dina(n36856), .dinb(b56 ), .dout(n38078));
  jand g20056(.dina(n37515), .dinb(n375), .dout(n38079));
  jor  g20057(.dina(n38079), .dinb(n38078), .dout(n38080));
  jand g20058(.dina(n38080), .dinb(n373), .dout(n38081));
  jnot g20059(.din(n38081), .dout(n38082));
  jor  g20060(.dina(n38082), .dinb(n38077), .dout(n38083));
  jand g20061(.dina(n38083), .dinb(n37515), .dout(n38084));
  jxor g20062(.dina(n37858), .dinb(b1 ), .dout(n38085));
  jand g20063(.dina(n38085), .dinb(n14905), .dout(n38086));
  jor  g20064(.dina(n38086), .dinb(n37854), .dout(n38087));
  jand g20065(.dina(n37862), .dinb(n38087), .dout(n38088));
  jor  g20066(.dina(n38088), .dinb(n37847), .dout(n38089));
  jand g20067(.dina(n37866), .dinb(n38089), .dout(n38090));
  jor  g20068(.dina(n38090), .dinb(n37841), .dout(n38091));
  jand g20069(.dina(n37870), .dinb(n38091), .dout(n38092));
  jor  g20070(.dina(n38092), .dinb(n37835), .dout(n38093));
  jand g20071(.dina(n37874), .dinb(n38093), .dout(n38094));
  jor  g20072(.dina(n38094), .dinb(n37829), .dout(n38095));
  jand g20073(.dina(n37878), .dinb(n38095), .dout(n38096));
  jor  g20074(.dina(n38096), .dinb(n37823), .dout(n38097));
  jand g20075(.dina(n37882), .dinb(n38097), .dout(n38098));
  jor  g20076(.dina(n38098), .dinb(n37817), .dout(n38099));
  jand g20077(.dina(n37886), .dinb(n38099), .dout(n38100));
  jor  g20078(.dina(n38100), .dinb(n37811), .dout(n38101));
  jand g20079(.dina(n37890), .dinb(n38101), .dout(n38102));
  jor  g20080(.dina(n38102), .dinb(n37805), .dout(n38103));
  jand g20081(.dina(n37894), .dinb(n38103), .dout(n38104));
  jor  g20082(.dina(n38104), .dinb(n37799), .dout(n38105));
  jand g20083(.dina(n37898), .dinb(n38105), .dout(n38106));
  jor  g20084(.dina(n38106), .dinb(n37793), .dout(n38107));
  jand g20085(.dina(n37902), .dinb(n38107), .dout(n38108));
  jor  g20086(.dina(n38108), .dinb(n37787), .dout(n38109));
  jand g20087(.dina(n37906), .dinb(n38109), .dout(n38110));
  jor  g20088(.dina(n38110), .dinb(n37781), .dout(n38111));
  jand g20089(.dina(n37910), .dinb(n38111), .dout(n38112));
  jor  g20090(.dina(n38112), .dinb(n37775), .dout(n38113));
  jand g20091(.dina(n37914), .dinb(n38113), .dout(n38114));
  jor  g20092(.dina(n38114), .dinb(n37769), .dout(n38115));
  jand g20093(.dina(n37918), .dinb(n38115), .dout(n38116));
  jor  g20094(.dina(n38116), .dinb(n37763), .dout(n38117));
  jand g20095(.dina(n37922), .dinb(n38117), .dout(n38118));
  jor  g20096(.dina(n38118), .dinb(n37757), .dout(n38119));
  jand g20097(.dina(n37926), .dinb(n38119), .dout(n38120));
  jor  g20098(.dina(n38120), .dinb(n37751), .dout(n38121));
  jand g20099(.dina(n37930), .dinb(n38121), .dout(n38122));
  jor  g20100(.dina(n38122), .dinb(n37745), .dout(n38123));
  jand g20101(.dina(n37934), .dinb(n38123), .dout(n38124));
  jor  g20102(.dina(n38124), .dinb(n37739), .dout(n38125));
  jand g20103(.dina(n37938), .dinb(n38125), .dout(n38126));
  jor  g20104(.dina(n38126), .dinb(n37733), .dout(n38127));
  jand g20105(.dina(n37942), .dinb(n38127), .dout(n38128));
  jor  g20106(.dina(n38128), .dinb(n37727), .dout(n38129));
  jand g20107(.dina(n37946), .dinb(n38129), .dout(n38130));
  jor  g20108(.dina(n38130), .dinb(n37721), .dout(n38131));
  jand g20109(.dina(n37950), .dinb(n38131), .dout(n38132));
  jor  g20110(.dina(n38132), .dinb(n37715), .dout(n38133));
  jand g20111(.dina(n37954), .dinb(n38133), .dout(n38134));
  jor  g20112(.dina(n38134), .dinb(n37709), .dout(n38135));
  jand g20113(.dina(n37958), .dinb(n38135), .dout(n38136));
  jor  g20114(.dina(n38136), .dinb(n37703), .dout(n38137));
  jand g20115(.dina(n37962), .dinb(n38137), .dout(n38138));
  jor  g20116(.dina(n38138), .dinb(n37697), .dout(n38139));
  jand g20117(.dina(n37966), .dinb(n38139), .dout(n38140));
  jor  g20118(.dina(n38140), .dinb(n37691), .dout(n38141));
  jand g20119(.dina(n37970), .dinb(n38141), .dout(n38142));
  jor  g20120(.dina(n38142), .dinb(n37685), .dout(n38143));
  jand g20121(.dina(n37974), .dinb(n38143), .dout(n38144));
  jor  g20122(.dina(n38144), .dinb(n37679), .dout(n38145));
  jand g20123(.dina(n37978), .dinb(n38145), .dout(n38146));
  jor  g20124(.dina(n38146), .dinb(n37673), .dout(n38147));
  jand g20125(.dina(n37982), .dinb(n38147), .dout(n38148));
  jor  g20126(.dina(n38148), .dinb(n37667), .dout(n38149));
  jand g20127(.dina(n37986), .dinb(n38149), .dout(n38150));
  jor  g20128(.dina(n38150), .dinb(n37661), .dout(n38151));
  jand g20129(.dina(n37990), .dinb(n38151), .dout(n38152));
  jor  g20130(.dina(n38152), .dinb(n37655), .dout(n38153));
  jand g20131(.dina(n37994), .dinb(n38153), .dout(n38154));
  jor  g20132(.dina(n38154), .dinb(n37649), .dout(n38155));
  jand g20133(.dina(n37998), .dinb(n38155), .dout(n38156));
  jor  g20134(.dina(n38156), .dinb(n37643), .dout(n38157));
  jand g20135(.dina(n38002), .dinb(n38157), .dout(n38158));
  jor  g20136(.dina(n38158), .dinb(n37637), .dout(n38159));
  jand g20137(.dina(n38006), .dinb(n38159), .dout(n38160));
  jor  g20138(.dina(n38160), .dinb(n37631), .dout(n38161));
  jand g20139(.dina(n38010), .dinb(n38161), .dout(n38162));
  jor  g20140(.dina(n38162), .dinb(n37625), .dout(n38163));
  jand g20141(.dina(n38014), .dinb(n38163), .dout(n38164));
  jor  g20142(.dina(n38164), .dinb(n37619), .dout(n38165));
  jand g20143(.dina(n38018), .dinb(n38165), .dout(n38166));
  jor  g20144(.dina(n38166), .dinb(n37613), .dout(n38167));
  jand g20145(.dina(n38022), .dinb(n38167), .dout(n38168));
  jor  g20146(.dina(n38168), .dinb(n37607), .dout(n38169));
  jand g20147(.dina(n38026), .dinb(n38169), .dout(n38170));
  jor  g20148(.dina(n38170), .dinb(n37601), .dout(n38171));
  jand g20149(.dina(n38030), .dinb(n38171), .dout(n38172));
  jor  g20150(.dina(n38172), .dinb(n37595), .dout(n38173));
  jand g20151(.dina(n38034), .dinb(n38173), .dout(n38174));
  jor  g20152(.dina(n38174), .dinb(n37589), .dout(n38175));
  jand g20153(.dina(n38038), .dinb(n38175), .dout(n38176));
  jor  g20154(.dina(n38176), .dinb(n37583), .dout(n38177));
  jand g20155(.dina(n38042), .dinb(n38177), .dout(n38178));
  jor  g20156(.dina(n38178), .dinb(n37577), .dout(n38179));
  jand g20157(.dina(n38046), .dinb(n38179), .dout(n38180));
  jor  g20158(.dina(n38180), .dinb(n37571), .dout(n38181));
  jand g20159(.dina(n38050), .dinb(n38181), .dout(n38182));
  jor  g20160(.dina(n38182), .dinb(n37565), .dout(n38183));
  jand g20161(.dina(n38054), .dinb(n38183), .dout(n38184));
  jor  g20162(.dina(n38184), .dinb(n37559), .dout(n38185));
  jand g20163(.dina(n38058), .dinb(n38185), .dout(n38186));
  jor  g20164(.dina(n38186), .dinb(n37553), .dout(n38187));
  jand g20165(.dina(n38062), .dinb(n38187), .dout(n38188));
  jor  g20166(.dina(n38188), .dinb(n37547), .dout(n38189));
  jand g20167(.dina(n38066), .dinb(n38189), .dout(n38190));
  jor  g20168(.dina(n38190), .dinb(n37541), .dout(n38191));
  jand g20169(.dina(n38070), .dinb(n38191), .dout(n38192));
  jor  g20170(.dina(n38192), .dinb(n37535), .dout(n38193));
  jand g20171(.dina(n38074), .dinb(n38193), .dout(n38194));
  jor  g20172(.dina(n38194), .dinb(n37529), .dout(n38195));
  jand g20173(.dina(n38081), .dinb(n38195), .dout(n38196));
  jand g20174(.dina(n37514), .dinb(n14053), .dout(n38197));
  jor  g20175(.dina(n38197), .dinb(n38196), .dout(n38198));
  jxor g20176(.dina(n38080), .dinb(n38077), .dout(n38199));
  jand g20177(.dina(n38199), .dinb(n38198), .dout(n38200));
  jor  g20178(.dina(n38200), .dinb(n38084), .dout(n38201));
  jnot g20179(.din(n38201), .dout(n38202));
  jnot g20180(.din(n15090), .dout(n38203));
  jand g20181(.dina(n38201), .dinb(b57 ), .dout(n38204));
  jand g20182(.dina(n38202), .dinb(n362), .dout(n38205));
  jnot g20183(.din(n38205), .dout(n38206));
  jnot g20184(.din(n38197), .dout(n38207));
  jand g20185(.dina(n38207), .dinb(n38083), .dout(n38208));
  jand g20186(.dina(n38208), .dinb(n37528), .dout(n38209));
  jxor g20187(.dina(n38074), .dinb(n38193), .dout(n38210));
  jand g20188(.dina(n38210), .dinb(n38198), .dout(n38211));
  jor  g20189(.dina(n38211), .dinb(n38209), .dout(n38212));
  jand g20190(.dina(n38212), .dinb(n375), .dout(n38213));
  jnot g20191(.din(n38213), .dout(n38214));
  jand g20192(.dina(n38208), .dinb(n37534), .dout(n38215));
  jxor g20193(.dina(n38070), .dinb(n38191), .dout(n38216));
  jand g20194(.dina(n38216), .dinb(n38198), .dout(n38217));
  jor  g20195(.dina(n38217), .dinb(n38215), .dout(n38218));
  jand g20196(.dina(n38218), .dinb(n377), .dout(n38219));
  jnot g20197(.din(n38219), .dout(n38220));
  jand g20198(.dina(n38208), .dinb(n37540), .dout(n38221));
  jxor g20199(.dina(n38066), .dinb(n38189), .dout(n38222));
  jand g20200(.dina(n38222), .dinb(n38198), .dout(n38223));
  jor  g20201(.dina(n38223), .dinb(n38221), .dout(n38224));
  jand g20202(.dina(n38224), .dinb(n376), .dout(n38225));
  jnot g20203(.din(n38225), .dout(n38226));
  jand g20204(.dina(n38208), .dinb(n37546), .dout(n38227));
  jxor g20205(.dina(n38062), .dinb(n38187), .dout(n38228));
  jand g20206(.dina(n38228), .dinb(n38198), .dout(n38229));
  jor  g20207(.dina(n38229), .dinb(n38227), .dout(n38230));
  jand g20208(.dina(n38230), .dinb(n374), .dout(n38231));
  jnot g20209(.din(n38231), .dout(n38232));
  jand g20210(.dina(n38208), .dinb(n37552), .dout(n38233));
  jxor g20211(.dina(n38058), .dinb(n38185), .dout(n38234));
  jand g20212(.dina(n38234), .dinb(n38198), .dout(n38235));
  jor  g20213(.dina(n38235), .dinb(n38233), .dout(n38236));
  jand g20214(.dina(n38236), .dinb(n384), .dout(n38237));
  jnot g20215(.din(n38237), .dout(n38238));
  jand g20216(.dina(n38208), .dinb(n37558), .dout(n38239));
  jxor g20217(.dina(n38054), .dinb(n38183), .dout(n38240));
  jand g20218(.dina(n38240), .dinb(n38198), .dout(n38241));
  jor  g20219(.dina(n38241), .dinb(n38239), .dout(n38242));
  jand g20220(.dina(n38242), .dinb(n12214), .dout(n38243));
  jnot g20221(.din(n38243), .dout(n38244));
  jand g20222(.dina(n38208), .dinb(n37564), .dout(n38245));
  jxor g20223(.dina(n38050), .dinb(n38181), .dout(n38246));
  jand g20224(.dina(n38246), .dinb(n38198), .dout(n38247));
  jor  g20225(.dina(n38247), .dinb(n38245), .dout(n38248));
  jand g20226(.dina(n38248), .dinb(n12211), .dout(n38249));
  jnot g20227(.din(n38249), .dout(n38250));
  jand g20228(.dina(n38208), .dinb(n37570), .dout(n38251));
  jxor g20229(.dina(n38046), .dinb(n38179), .dout(n38252));
  jand g20230(.dina(n38252), .dinb(n38198), .dout(n38253));
  jor  g20231(.dina(n38253), .dinb(n38251), .dout(n38254));
  jand g20232(.dina(n38254), .dinb(n383), .dout(n38255));
  jnot g20233(.din(n38255), .dout(n38256));
  jand g20234(.dina(n38208), .dinb(n37576), .dout(n38257));
  jxor g20235(.dina(n38042), .dinb(n38177), .dout(n38258));
  jand g20236(.dina(n38258), .dinb(n38198), .dout(n38259));
  jor  g20237(.dina(n38259), .dinb(n38257), .dout(n38260));
  jand g20238(.dina(n38260), .dinb(n396), .dout(n38261));
  jnot g20239(.din(n38261), .dout(n38262));
  jand g20240(.dina(n38208), .dinb(n37582), .dout(n38263));
  jxor g20241(.dina(n38038), .dinb(n38175), .dout(n38264));
  jand g20242(.dina(n38264), .dinb(n38198), .dout(n38265));
  jor  g20243(.dina(n38265), .dinb(n38263), .dout(n38266));
  jand g20244(.dina(n38266), .dinb(n510), .dout(n38267));
  jnot g20245(.din(n38267), .dout(n38268));
  jand g20246(.dina(n38208), .dinb(n37588), .dout(n38269));
  jxor g20247(.dina(n38034), .dinb(n38173), .dout(n38270));
  jand g20248(.dina(n38270), .dinb(n38198), .dout(n38271));
  jor  g20249(.dina(n38271), .dinb(n38269), .dout(n38272));
  jand g20250(.dina(n38272), .dinb(n514), .dout(n38273));
  jnot g20251(.din(n38273), .dout(n38274));
  jand g20252(.dina(n38208), .dinb(n37594), .dout(n38275));
  jxor g20253(.dina(n38030), .dinb(n38171), .dout(n38276));
  jand g20254(.dina(n38276), .dinb(n38198), .dout(n38277));
  jor  g20255(.dina(n38277), .dinb(n38275), .dout(n38278));
  jand g20256(.dina(n38278), .dinb(n513), .dout(n38279));
  jnot g20257(.din(n38279), .dout(n38280));
  jand g20258(.dina(n38208), .dinb(n37600), .dout(n38281));
  jxor g20259(.dina(n38026), .dinb(n38169), .dout(n38282));
  jand g20260(.dina(n38282), .dinb(n38198), .dout(n38283));
  jor  g20261(.dina(n38283), .dinb(n38281), .dout(n38284));
  jand g20262(.dina(n38284), .dinb(n397), .dout(n38285));
  jnot g20263(.din(n38285), .dout(n38286));
  jand g20264(.dina(n38208), .dinb(n37606), .dout(n38287));
  jxor g20265(.dina(n38022), .dinb(n38167), .dout(n38288));
  jand g20266(.dina(n38288), .dinb(n38198), .dout(n38289));
  jor  g20267(.dina(n38289), .dinb(n38287), .dout(n38290));
  jand g20268(.dina(n38290), .dinb(n282), .dout(n38291));
  jnot g20269(.din(n38291), .dout(n38292));
  jand g20270(.dina(n38208), .dinb(n37612), .dout(n38293));
  jxor g20271(.dina(n38018), .dinb(n38165), .dout(n38294));
  jand g20272(.dina(n38294), .dinb(n38198), .dout(n38295));
  jor  g20273(.dina(n38295), .dinb(n38293), .dout(n38296));
  jand g20274(.dina(n38296), .dinb(n281), .dout(n38297));
  jnot g20275(.din(n38297), .dout(n38298));
  jand g20276(.dina(n38208), .dinb(n37618), .dout(n38299));
  jxor g20277(.dina(n38014), .dinb(n38163), .dout(n38300));
  jand g20278(.dina(n38300), .dinb(n38198), .dout(n38301));
  jor  g20279(.dina(n38301), .dinb(n38299), .dout(n38302));
  jand g20280(.dina(n38302), .dinb(n285), .dout(n38303));
  jnot g20281(.din(n38303), .dout(n38304));
  jand g20282(.dina(n38208), .dinb(n37624), .dout(n38305));
  jxor g20283(.dina(n38010), .dinb(n38161), .dout(n38306));
  jand g20284(.dina(n38306), .dinb(n38198), .dout(n38307));
  jor  g20285(.dina(n38307), .dinb(n38305), .dout(n38308));
  jand g20286(.dina(n38308), .dinb(n284), .dout(n38309));
  jnot g20287(.din(n38309), .dout(n38310));
  jand g20288(.dina(n38208), .dinb(n37630), .dout(n38311));
  jxor g20289(.dina(n38006), .dinb(n38159), .dout(n38312));
  jand g20290(.dina(n38312), .dinb(n38198), .dout(n38313));
  jor  g20291(.dina(n38313), .dinb(n38311), .dout(n38314));
  jand g20292(.dina(n38314), .dinb(n291), .dout(n38315));
  jnot g20293(.din(n38315), .dout(n38316));
  jand g20294(.dina(n38208), .dinb(n37636), .dout(n38317));
  jxor g20295(.dina(n38002), .dinb(n38157), .dout(n38318));
  jand g20296(.dina(n38318), .dinb(n38198), .dout(n38319));
  jor  g20297(.dina(n38319), .dinb(n38317), .dout(n38320));
  jand g20298(.dina(n38320), .dinb(n290), .dout(n38321));
  jnot g20299(.din(n38321), .dout(n38322));
  jand g20300(.dina(n38208), .dinb(n37642), .dout(n38323));
  jxor g20301(.dina(n37998), .dinb(n38155), .dout(n38324));
  jand g20302(.dina(n38324), .dinb(n38198), .dout(n38325));
  jor  g20303(.dina(n38325), .dinb(n38323), .dout(n38326));
  jand g20304(.dina(n38326), .dinb(n294), .dout(n38327));
  jnot g20305(.din(n38327), .dout(n38328));
  jand g20306(.dina(n38208), .dinb(n37648), .dout(n38329));
  jxor g20307(.dina(n37994), .dinb(n38153), .dout(n38330));
  jand g20308(.dina(n38330), .dinb(n38198), .dout(n38331));
  jor  g20309(.dina(n38331), .dinb(n38329), .dout(n38332));
  jand g20310(.dina(n38332), .dinb(n293), .dout(n38333));
  jnot g20311(.din(n38333), .dout(n38334));
  jand g20312(.dina(n38208), .dinb(n37654), .dout(n38335));
  jxor g20313(.dina(n37990), .dinb(n38151), .dout(n38336));
  jand g20314(.dina(n38336), .dinb(n38198), .dout(n38337));
  jor  g20315(.dina(n38337), .dinb(n38335), .dout(n38338));
  jand g20316(.dina(n38338), .dinb(n301), .dout(n38339));
  jnot g20317(.din(n38339), .dout(n38340));
  jand g20318(.dina(n38208), .dinb(n37660), .dout(n38341));
  jxor g20319(.dina(n37986), .dinb(n38149), .dout(n38342));
  jand g20320(.dina(n38342), .dinb(n38198), .dout(n38343));
  jor  g20321(.dina(n38343), .dinb(n38341), .dout(n38344));
  jand g20322(.dina(n38344), .dinb(n298), .dout(n38345));
  jnot g20323(.din(n38345), .dout(n38346));
  jand g20324(.dina(n38208), .dinb(n37666), .dout(n38347));
  jxor g20325(.dina(n37982), .dinb(n38147), .dout(n38348));
  jand g20326(.dina(n38348), .dinb(n38198), .dout(n38349));
  jor  g20327(.dina(n38349), .dinb(n38347), .dout(n38350));
  jand g20328(.dina(n38350), .dinb(n297), .dout(n38351));
  jnot g20329(.din(n38351), .dout(n38352));
  jand g20330(.dina(n38208), .dinb(n37672), .dout(n38353));
  jxor g20331(.dina(n37978), .dinb(n38145), .dout(n38354));
  jand g20332(.dina(n38354), .dinb(n38198), .dout(n38355));
  jor  g20333(.dina(n38355), .dinb(n38353), .dout(n38356));
  jand g20334(.dina(n38356), .dinb(n300), .dout(n38357));
  jnot g20335(.din(n38357), .dout(n38358));
  jand g20336(.dina(n38208), .dinb(n37678), .dout(n38359));
  jxor g20337(.dina(n37974), .dinb(n38143), .dout(n38360));
  jand g20338(.dina(n38360), .dinb(n38198), .dout(n38361));
  jor  g20339(.dina(n38361), .dinb(n38359), .dout(n38362));
  jand g20340(.dina(n38362), .dinb(n424), .dout(n38363));
  jnot g20341(.din(n38363), .dout(n38364));
  jand g20342(.dina(n38208), .dinb(n37684), .dout(n38365));
  jxor g20343(.dina(n37970), .dinb(n38141), .dout(n38366));
  jand g20344(.dina(n38366), .dinb(n38198), .dout(n38367));
  jor  g20345(.dina(n38367), .dinb(n38365), .dout(n38368));
  jand g20346(.dina(n38368), .dinb(n427), .dout(n38369));
  jnot g20347(.din(n38369), .dout(n38370));
  jand g20348(.dina(n38208), .dinb(n37690), .dout(n38371));
  jxor g20349(.dina(n37966), .dinb(n38139), .dout(n38372));
  jand g20350(.dina(n38372), .dinb(n38198), .dout(n38373));
  jor  g20351(.dina(n38373), .dinb(n38371), .dout(n38374));
  jand g20352(.dina(n38374), .dinb(n426), .dout(n38375));
  jnot g20353(.din(n38375), .dout(n38376));
  jand g20354(.dina(n38208), .dinb(n37696), .dout(n38377));
  jxor g20355(.dina(n37962), .dinb(n38137), .dout(n38378));
  jand g20356(.dina(n38378), .dinb(n38198), .dout(n38379));
  jor  g20357(.dina(n38379), .dinb(n38377), .dout(n38380));
  jand g20358(.dina(n38380), .dinb(n410), .dout(n38381));
  jnot g20359(.din(n38381), .dout(n38382));
  jand g20360(.dina(n38208), .dinb(n37702), .dout(n38383));
  jxor g20361(.dina(n37958), .dinb(n38135), .dout(n38384));
  jand g20362(.dina(n38384), .dinb(n38198), .dout(n38385));
  jor  g20363(.dina(n38385), .dinb(n38383), .dout(n38386));
  jand g20364(.dina(n38386), .dinb(n409), .dout(n38387));
  jnot g20365(.din(n38387), .dout(n38388));
  jand g20366(.dina(n38208), .dinb(n37708), .dout(n38389));
  jxor g20367(.dina(n37954), .dinb(n38133), .dout(n38390));
  jand g20368(.dina(n38390), .dinb(n38198), .dout(n38391));
  jor  g20369(.dina(n38391), .dinb(n38389), .dout(n38392));
  jand g20370(.dina(n38392), .dinb(n413), .dout(n38393));
  jnot g20371(.din(n38393), .dout(n38394));
  jand g20372(.dina(n38208), .dinb(n37714), .dout(n38395));
  jxor g20373(.dina(n37950), .dinb(n38131), .dout(n38396));
  jand g20374(.dina(n38396), .dinb(n38198), .dout(n38397));
  jor  g20375(.dina(n38397), .dinb(n38395), .dout(n38398));
  jand g20376(.dina(n38398), .dinb(n412), .dout(n38399));
  jnot g20377(.din(n38399), .dout(n38400));
  jand g20378(.dina(n38208), .dinb(n37720), .dout(n38401));
  jxor g20379(.dina(n37946), .dinb(n38129), .dout(n38402));
  jand g20380(.dina(n38402), .dinb(n38198), .dout(n38403));
  jor  g20381(.dina(n38403), .dinb(n38401), .dout(n38404));
  jand g20382(.dina(n38404), .dinb(n406), .dout(n38405));
  jnot g20383(.din(n38405), .dout(n38406));
  jand g20384(.dina(n38208), .dinb(n37726), .dout(n38407));
  jxor g20385(.dina(n37942), .dinb(n38127), .dout(n38408));
  jand g20386(.dina(n38408), .dinb(n38198), .dout(n38409));
  jor  g20387(.dina(n38409), .dinb(n38407), .dout(n38410));
  jand g20388(.dina(n38410), .dinb(n405), .dout(n38411));
  jnot g20389(.din(n38411), .dout(n38412));
  jand g20390(.dina(n38208), .dinb(n37732), .dout(n38413));
  jxor g20391(.dina(n37938), .dinb(n38125), .dout(n38414));
  jand g20392(.dina(n38414), .dinb(n38198), .dout(n38415));
  jor  g20393(.dina(n38415), .dinb(n38413), .dout(n38416));
  jand g20394(.dina(n38416), .dinb(n2714), .dout(n38417));
  jnot g20395(.din(n38417), .dout(n38418));
  jand g20396(.dina(n38208), .dinb(n37738), .dout(n38419));
  jxor g20397(.dina(n37934), .dinb(n38123), .dout(n38420));
  jand g20398(.dina(n38420), .dinb(n38198), .dout(n38421));
  jor  g20399(.dina(n38421), .dinb(n38419), .dout(n38422));
  jand g20400(.dina(n38422), .dinb(n2547), .dout(n38423));
  jnot g20401(.din(n38423), .dout(n38424));
  jand g20402(.dina(n38208), .dinb(n37744), .dout(n38425));
  jxor g20403(.dina(n37930), .dinb(n38121), .dout(n38426));
  jand g20404(.dina(n38426), .dinb(n38198), .dout(n38427));
  jor  g20405(.dina(n38427), .dinb(n38425), .dout(n38428));
  jand g20406(.dina(n38428), .dinb(n417), .dout(n38429));
  jnot g20407(.din(n38429), .dout(n38430));
  jand g20408(.dina(n38208), .dinb(n37750), .dout(n38431));
  jxor g20409(.dina(n37926), .dinb(n38119), .dout(n38432));
  jand g20410(.dina(n38432), .dinb(n38198), .dout(n38433));
  jor  g20411(.dina(n38433), .dinb(n38431), .dout(n38434));
  jand g20412(.dina(n38434), .dinb(n416), .dout(n38435));
  jnot g20413(.din(n38435), .dout(n38436));
  jand g20414(.dina(n38208), .dinb(n37756), .dout(n38437));
  jxor g20415(.dina(n37922), .dinb(n38117), .dout(n38438));
  jand g20416(.dina(n38438), .dinb(n38198), .dout(n38439));
  jor  g20417(.dina(n38439), .dinb(n38437), .dout(n38440));
  jand g20418(.dina(n38440), .dinb(n422), .dout(n38441));
  jnot g20419(.din(n38441), .dout(n38442));
  jand g20420(.dina(n38208), .dinb(n37762), .dout(n38443));
  jxor g20421(.dina(n37918), .dinb(n38115), .dout(n38444));
  jand g20422(.dina(n38444), .dinb(n38198), .dout(n38445));
  jor  g20423(.dina(n38445), .dinb(n38443), .dout(n38446));
  jand g20424(.dina(n38446), .dinb(n421), .dout(n38447));
  jnot g20425(.din(n38447), .dout(n38448));
  jand g20426(.dina(n38208), .dinb(n37768), .dout(n38449));
  jxor g20427(.dina(n37914), .dinb(n38113), .dout(n38450));
  jand g20428(.dina(n38450), .dinb(n38198), .dout(n38451));
  jor  g20429(.dina(n38451), .dinb(n38449), .dout(n38452));
  jand g20430(.dina(n38452), .dinb(n433), .dout(n38453));
  jnot g20431(.din(n38453), .dout(n38454));
  jand g20432(.dina(n38208), .dinb(n37774), .dout(n38455));
  jxor g20433(.dina(n37910), .dinb(n38111), .dout(n38456));
  jand g20434(.dina(n38456), .dinb(n38198), .dout(n38457));
  jor  g20435(.dina(n38457), .dinb(n38455), .dout(n38458));
  jand g20436(.dina(n38458), .dinb(n432), .dout(n38459));
  jnot g20437(.din(n38459), .dout(n38460));
  jand g20438(.dina(n38208), .dinb(n37780), .dout(n38461));
  jxor g20439(.dina(n37906), .dinb(n38109), .dout(n38462));
  jand g20440(.dina(n38462), .dinb(n38198), .dout(n38463));
  jor  g20441(.dina(n38463), .dinb(n38461), .dout(n38464));
  jand g20442(.dina(n38464), .dinb(n436), .dout(n38465));
  jnot g20443(.din(n38465), .dout(n38466));
  jand g20444(.dina(n38208), .dinb(n37786), .dout(n38467));
  jxor g20445(.dina(n37902), .dinb(n38107), .dout(n38468));
  jand g20446(.dina(n38468), .dinb(n38198), .dout(n38469));
  jor  g20447(.dina(n38469), .dinb(n38467), .dout(n38470));
  jand g20448(.dina(n38470), .dinb(n435), .dout(n38471));
  jnot g20449(.din(n38471), .dout(n38472));
  jand g20450(.dina(n38208), .dinb(n37792), .dout(n38473));
  jxor g20451(.dina(n37898), .dinb(n38105), .dout(n38474));
  jand g20452(.dina(n38474), .dinb(n38198), .dout(n38475));
  jor  g20453(.dina(n38475), .dinb(n38473), .dout(n38476));
  jand g20454(.dina(n38476), .dinb(n440), .dout(n38477));
  jnot g20455(.din(n38477), .dout(n38478));
  jand g20456(.dina(n38208), .dinb(n37798), .dout(n38479));
  jxor g20457(.dina(n37894), .dinb(n38103), .dout(n38480));
  jand g20458(.dina(n38480), .dinb(n38198), .dout(n38481));
  jor  g20459(.dina(n38481), .dinb(n38479), .dout(n38482));
  jand g20460(.dina(n38482), .dinb(n439), .dout(n38483));
  jnot g20461(.din(n38483), .dout(n38484));
  jand g20462(.dina(n38208), .dinb(n37804), .dout(n38485));
  jxor g20463(.dina(n37890), .dinb(n38101), .dout(n38486));
  jand g20464(.dina(n38486), .dinb(n38198), .dout(n38487));
  jor  g20465(.dina(n38487), .dinb(n38485), .dout(n38488));
  jand g20466(.dina(n38488), .dinb(n325), .dout(n38489));
  jnot g20467(.din(n38489), .dout(n38490));
  jand g20468(.dina(n38208), .dinb(n37810), .dout(n38491));
  jxor g20469(.dina(n37886), .dinb(n38099), .dout(n38492));
  jand g20470(.dina(n38492), .dinb(n38198), .dout(n38493));
  jor  g20471(.dina(n38493), .dinb(n38491), .dout(n38494));
  jand g20472(.dina(n38494), .dinb(n324), .dout(n38495));
  jnot g20473(.din(n38495), .dout(n38496));
  jand g20474(.dina(n38208), .dinb(n37816), .dout(n38497));
  jxor g20475(.dina(n37882), .dinb(n38097), .dout(n38498));
  jand g20476(.dina(n38498), .dinb(n38198), .dout(n38499));
  jor  g20477(.dina(n38499), .dinb(n38497), .dout(n38500));
  jand g20478(.dina(n38500), .dinb(n323), .dout(n38501));
  jnot g20479(.din(n38501), .dout(n38502));
  jand g20480(.dina(n38208), .dinb(n37822), .dout(n38503));
  jxor g20481(.dina(n37878), .dinb(n38095), .dout(n38504));
  jand g20482(.dina(n38504), .dinb(n38198), .dout(n38505));
  jor  g20483(.dina(n38505), .dinb(n38503), .dout(n38506));
  jand g20484(.dina(n38506), .dinb(n335), .dout(n38507));
  jnot g20485(.din(n38507), .dout(n38508));
  jand g20486(.dina(n38208), .dinb(n37828), .dout(n38509));
  jxor g20487(.dina(n37874), .dinb(n38093), .dout(n38510));
  jand g20488(.dina(n38510), .dinb(n38198), .dout(n38511));
  jor  g20489(.dina(n38511), .dinb(n38509), .dout(n38512));
  jand g20490(.dina(n38512), .dinb(n334), .dout(n38513));
  jnot g20491(.din(n38513), .dout(n38514));
  jand g20492(.dina(n38208), .dinb(n37834), .dout(n38515));
  jxor g20493(.dina(n37870), .dinb(n38091), .dout(n38516));
  jand g20494(.dina(n38516), .dinb(n38198), .dout(n38517));
  jor  g20495(.dina(n38517), .dinb(n38515), .dout(n38518));
  jand g20496(.dina(n38518), .dinb(n338), .dout(n38519));
  jnot g20497(.din(n38519), .dout(n38520));
  jand g20498(.dina(n38208), .dinb(n37840), .dout(n38521));
  jxor g20499(.dina(n37866), .dinb(n38089), .dout(n38522));
  jand g20500(.dina(n38522), .dinb(n38198), .dout(n38523));
  jor  g20501(.dina(n38523), .dinb(n38521), .dout(n38524));
  jand g20502(.dina(n38524), .dinb(n337), .dout(n38525));
  jnot g20503(.din(n38525), .dout(n38526));
  jand g20504(.dina(n38208), .dinb(n37846), .dout(n38527));
  jxor g20505(.dina(n37862), .dinb(n38087), .dout(n38528));
  jand g20506(.dina(n38528), .dinb(n38198), .dout(n38529));
  jor  g20507(.dina(n38529), .dinb(n38527), .dout(n38530));
  jand g20508(.dina(n38530), .dinb(n344), .dout(n38531));
  jnot g20509(.din(n38531), .dout(n38532));
  jand g20510(.dina(n38208), .dinb(n37853), .dout(n38533));
  jxor g20511(.dina(n38085), .dinb(n14905), .dout(n38534));
  jand g20512(.dina(n38534), .dinb(n38198), .dout(n38535));
  jor  g20513(.dina(n38535), .dinb(n38533), .dout(n38536));
  jand g20514(.dina(n38536), .dinb(n348), .dout(n38537));
  jnot g20515(.din(n38537), .dout(n38538));
  jor  g20516(.dina(n38208), .dinb(n18364), .dout(n38539));
  jand g20517(.dina(n38539), .dinb(a7 ), .dout(n38540));
  jor  g20518(.dina(n38208), .dinb(n14905), .dout(n38541));
  jnot g20519(.din(n38541), .dout(n38542));
  jor  g20520(.dina(n38542), .dinb(n38540), .dout(n38543));
  jand g20521(.dina(n38543), .dinb(n258), .dout(n38544));
  jnot g20522(.din(n38544), .dout(n38545));
  jand g20523(.dina(n38198), .dinb(b0 ), .dout(n38546));
  jor  g20524(.dina(n38546), .dinb(n14903), .dout(n38547));
  jand g20525(.dina(n38541), .dinb(n38547), .dout(n38548));
  jxor g20526(.dina(n38548), .dinb(n258), .dout(n38549));
  jor  g20527(.dina(n38549), .dinb(n15382), .dout(n38550));
  jand g20528(.dina(n38550), .dinb(n38545), .dout(n38551));
  jxor g20529(.dina(n38536), .dinb(n348), .dout(n38552));
  jnot g20530(.din(n38552), .dout(n38553));
  jor  g20531(.dina(n38553), .dinb(n38551), .dout(n38554));
  jand g20532(.dina(n38554), .dinb(n38538), .dout(n38555));
  jxor g20533(.dina(n38530), .dinb(n344), .dout(n38556));
  jnot g20534(.din(n38556), .dout(n38557));
  jor  g20535(.dina(n38557), .dinb(n38555), .dout(n38558));
  jand g20536(.dina(n38558), .dinb(n38532), .dout(n38559));
  jxor g20537(.dina(n38524), .dinb(n337), .dout(n38560));
  jnot g20538(.din(n38560), .dout(n38561));
  jor  g20539(.dina(n38561), .dinb(n38559), .dout(n38562));
  jand g20540(.dina(n38562), .dinb(n38526), .dout(n38563));
  jxor g20541(.dina(n38518), .dinb(n338), .dout(n38564));
  jnot g20542(.din(n38564), .dout(n38565));
  jor  g20543(.dina(n38565), .dinb(n38563), .dout(n38566));
  jand g20544(.dina(n38566), .dinb(n38520), .dout(n38567));
  jxor g20545(.dina(n38512), .dinb(n334), .dout(n38568));
  jnot g20546(.din(n38568), .dout(n38569));
  jor  g20547(.dina(n38569), .dinb(n38567), .dout(n38570));
  jand g20548(.dina(n38570), .dinb(n38514), .dout(n38571));
  jxor g20549(.dina(n38506), .dinb(n335), .dout(n38572));
  jnot g20550(.din(n38572), .dout(n38573));
  jor  g20551(.dina(n38573), .dinb(n38571), .dout(n38574));
  jand g20552(.dina(n38574), .dinb(n38508), .dout(n38575));
  jxor g20553(.dina(n38500), .dinb(n323), .dout(n38576));
  jnot g20554(.din(n38576), .dout(n38577));
  jor  g20555(.dina(n38577), .dinb(n38575), .dout(n38578));
  jand g20556(.dina(n38578), .dinb(n38502), .dout(n38579));
  jxor g20557(.dina(n38494), .dinb(n324), .dout(n38580));
  jnot g20558(.din(n38580), .dout(n38581));
  jor  g20559(.dina(n38581), .dinb(n38579), .dout(n38582));
  jand g20560(.dina(n38582), .dinb(n38496), .dout(n38583));
  jxor g20561(.dina(n38488), .dinb(n325), .dout(n38584));
  jnot g20562(.din(n38584), .dout(n38585));
  jor  g20563(.dina(n38585), .dinb(n38583), .dout(n38586));
  jand g20564(.dina(n38586), .dinb(n38490), .dout(n38587));
  jxor g20565(.dina(n38482), .dinb(n439), .dout(n38588));
  jnot g20566(.din(n38588), .dout(n38589));
  jor  g20567(.dina(n38589), .dinb(n38587), .dout(n38590));
  jand g20568(.dina(n38590), .dinb(n38484), .dout(n38591));
  jxor g20569(.dina(n38476), .dinb(n440), .dout(n38592));
  jnot g20570(.din(n38592), .dout(n38593));
  jor  g20571(.dina(n38593), .dinb(n38591), .dout(n38594));
  jand g20572(.dina(n38594), .dinb(n38478), .dout(n38595));
  jxor g20573(.dina(n38470), .dinb(n435), .dout(n38596));
  jnot g20574(.din(n38596), .dout(n38597));
  jor  g20575(.dina(n38597), .dinb(n38595), .dout(n38598));
  jand g20576(.dina(n38598), .dinb(n38472), .dout(n38599));
  jxor g20577(.dina(n38464), .dinb(n436), .dout(n38600));
  jnot g20578(.din(n38600), .dout(n38601));
  jor  g20579(.dina(n38601), .dinb(n38599), .dout(n38602));
  jand g20580(.dina(n38602), .dinb(n38466), .dout(n38603));
  jxor g20581(.dina(n38458), .dinb(n432), .dout(n38604));
  jnot g20582(.din(n38604), .dout(n38605));
  jor  g20583(.dina(n38605), .dinb(n38603), .dout(n38606));
  jand g20584(.dina(n38606), .dinb(n38460), .dout(n38607));
  jxor g20585(.dina(n38452), .dinb(n433), .dout(n38608));
  jnot g20586(.din(n38608), .dout(n38609));
  jor  g20587(.dina(n38609), .dinb(n38607), .dout(n38610));
  jand g20588(.dina(n38610), .dinb(n38454), .dout(n38611));
  jxor g20589(.dina(n38446), .dinb(n421), .dout(n38612));
  jnot g20590(.din(n38612), .dout(n38613));
  jor  g20591(.dina(n38613), .dinb(n38611), .dout(n38614));
  jand g20592(.dina(n38614), .dinb(n38448), .dout(n38615));
  jxor g20593(.dina(n38440), .dinb(n422), .dout(n38616));
  jnot g20594(.din(n38616), .dout(n38617));
  jor  g20595(.dina(n38617), .dinb(n38615), .dout(n38618));
  jand g20596(.dina(n38618), .dinb(n38442), .dout(n38619));
  jxor g20597(.dina(n38434), .dinb(n416), .dout(n38620));
  jnot g20598(.din(n38620), .dout(n38621));
  jor  g20599(.dina(n38621), .dinb(n38619), .dout(n38622));
  jand g20600(.dina(n38622), .dinb(n38436), .dout(n38623));
  jxor g20601(.dina(n38428), .dinb(n417), .dout(n38624));
  jnot g20602(.din(n38624), .dout(n38625));
  jor  g20603(.dina(n38625), .dinb(n38623), .dout(n38626));
  jand g20604(.dina(n38626), .dinb(n38430), .dout(n38627));
  jxor g20605(.dina(n38422), .dinb(n2547), .dout(n38628));
  jnot g20606(.din(n38628), .dout(n38629));
  jor  g20607(.dina(n38629), .dinb(n38627), .dout(n38630));
  jand g20608(.dina(n38630), .dinb(n38424), .dout(n38631));
  jxor g20609(.dina(n38416), .dinb(n2714), .dout(n38632));
  jnot g20610(.din(n38632), .dout(n38633));
  jor  g20611(.dina(n38633), .dinb(n38631), .dout(n38634));
  jand g20612(.dina(n38634), .dinb(n38418), .dout(n38635));
  jxor g20613(.dina(n38410), .dinb(n405), .dout(n38636));
  jnot g20614(.din(n38636), .dout(n38637));
  jor  g20615(.dina(n38637), .dinb(n38635), .dout(n38638));
  jand g20616(.dina(n38638), .dinb(n38412), .dout(n38639));
  jxor g20617(.dina(n38404), .dinb(n406), .dout(n38640));
  jnot g20618(.din(n38640), .dout(n38641));
  jor  g20619(.dina(n38641), .dinb(n38639), .dout(n38642));
  jand g20620(.dina(n38642), .dinb(n38406), .dout(n38643));
  jxor g20621(.dina(n38398), .dinb(n412), .dout(n38644));
  jnot g20622(.din(n38644), .dout(n38645));
  jor  g20623(.dina(n38645), .dinb(n38643), .dout(n38646));
  jand g20624(.dina(n38646), .dinb(n38400), .dout(n38647));
  jxor g20625(.dina(n38392), .dinb(n413), .dout(n38648));
  jnot g20626(.din(n38648), .dout(n38649));
  jor  g20627(.dina(n38649), .dinb(n38647), .dout(n38650));
  jand g20628(.dina(n38650), .dinb(n38394), .dout(n38651));
  jxor g20629(.dina(n38386), .dinb(n409), .dout(n38652));
  jnot g20630(.din(n38652), .dout(n38653));
  jor  g20631(.dina(n38653), .dinb(n38651), .dout(n38654));
  jand g20632(.dina(n38654), .dinb(n38388), .dout(n38655));
  jxor g20633(.dina(n38380), .dinb(n410), .dout(n38656));
  jnot g20634(.din(n38656), .dout(n38657));
  jor  g20635(.dina(n38657), .dinb(n38655), .dout(n38658));
  jand g20636(.dina(n38658), .dinb(n38382), .dout(n38659));
  jxor g20637(.dina(n38374), .dinb(n426), .dout(n38660));
  jnot g20638(.din(n38660), .dout(n38661));
  jor  g20639(.dina(n38661), .dinb(n38659), .dout(n38662));
  jand g20640(.dina(n38662), .dinb(n38376), .dout(n38663));
  jxor g20641(.dina(n38368), .dinb(n427), .dout(n38664));
  jnot g20642(.din(n38664), .dout(n38665));
  jor  g20643(.dina(n38665), .dinb(n38663), .dout(n38666));
  jand g20644(.dina(n38666), .dinb(n38370), .dout(n38667));
  jxor g20645(.dina(n38362), .dinb(n424), .dout(n38668));
  jnot g20646(.din(n38668), .dout(n38669));
  jor  g20647(.dina(n38669), .dinb(n38667), .dout(n38670));
  jand g20648(.dina(n38670), .dinb(n38364), .dout(n38671));
  jxor g20649(.dina(n38356), .dinb(n300), .dout(n38672));
  jnot g20650(.din(n38672), .dout(n38673));
  jor  g20651(.dina(n38673), .dinb(n38671), .dout(n38674));
  jand g20652(.dina(n38674), .dinb(n38358), .dout(n38675));
  jxor g20653(.dina(n38350), .dinb(n297), .dout(n38676));
  jnot g20654(.din(n38676), .dout(n38677));
  jor  g20655(.dina(n38677), .dinb(n38675), .dout(n38678));
  jand g20656(.dina(n38678), .dinb(n38352), .dout(n38679));
  jxor g20657(.dina(n38344), .dinb(n298), .dout(n38680));
  jnot g20658(.din(n38680), .dout(n38681));
  jor  g20659(.dina(n38681), .dinb(n38679), .dout(n38682));
  jand g20660(.dina(n38682), .dinb(n38346), .dout(n38683));
  jxor g20661(.dina(n38338), .dinb(n301), .dout(n38684));
  jnot g20662(.din(n38684), .dout(n38685));
  jor  g20663(.dina(n38685), .dinb(n38683), .dout(n38686));
  jand g20664(.dina(n38686), .dinb(n38340), .dout(n38687));
  jxor g20665(.dina(n38332), .dinb(n293), .dout(n38688));
  jnot g20666(.din(n38688), .dout(n38689));
  jor  g20667(.dina(n38689), .dinb(n38687), .dout(n38690));
  jand g20668(.dina(n38690), .dinb(n38334), .dout(n38691));
  jxor g20669(.dina(n38326), .dinb(n294), .dout(n38692));
  jnot g20670(.din(n38692), .dout(n38693));
  jor  g20671(.dina(n38693), .dinb(n38691), .dout(n38694));
  jand g20672(.dina(n38694), .dinb(n38328), .dout(n38695));
  jxor g20673(.dina(n38320), .dinb(n290), .dout(n38696));
  jnot g20674(.din(n38696), .dout(n38697));
  jor  g20675(.dina(n38697), .dinb(n38695), .dout(n38698));
  jand g20676(.dina(n38698), .dinb(n38322), .dout(n38699));
  jxor g20677(.dina(n38314), .dinb(n291), .dout(n38700));
  jnot g20678(.din(n38700), .dout(n38701));
  jor  g20679(.dina(n38701), .dinb(n38699), .dout(n38702));
  jand g20680(.dina(n38702), .dinb(n38316), .dout(n38703));
  jxor g20681(.dina(n38308), .dinb(n284), .dout(n38704));
  jnot g20682(.din(n38704), .dout(n38705));
  jor  g20683(.dina(n38705), .dinb(n38703), .dout(n38706));
  jand g20684(.dina(n38706), .dinb(n38310), .dout(n38707));
  jxor g20685(.dina(n38302), .dinb(n285), .dout(n38708));
  jnot g20686(.din(n38708), .dout(n38709));
  jor  g20687(.dina(n38709), .dinb(n38707), .dout(n38710));
  jand g20688(.dina(n38710), .dinb(n38304), .dout(n38711));
  jxor g20689(.dina(n38296), .dinb(n281), .dout(n38712));
  jnot g20690(.din(n38712), .dout(n38713));
  jor  g20691(.dina(n38713), .dinb(n38711), .dout(n38714));
  jand g20692(.dina(n38714), .dinb(n38298), .dout(n38715));
  jxor g20693(.dina(n38290), .dinb(n282), .dout(n38716));
  jnot g20694(.din(n38716), .dout(n38717));
  jor  g20695(.dina(n38717), .dinb(n38715), .dout(n38718));
  jand g20696(.dina(n38718), .dinb(n38292), .dout(n38719));
  jxor g20697(.dina(n38284), .dinb(n397), .dout(n38720));
  jnot g20698(.din(n38720), .dout(n38721));
  jor  g20699(.dina(n38721), .dinb(n38719), .dout(n38722));
  jand g20700(.dina(n38722), .dinb(n38286), .dout(n38723));
  jxor g20701(.dina(n38278), .dinb(n513), .dout(n38724));
  jnot g20702(.din(n38724), .dout(n38725));
  jor  g20703(.dina(n38725), .dinb(n38723), .dout(n38726));
  jand g20704(.dina(n38726), .dinb(n38280), .dout(n38727));
  jxor g20705(.dina(n38272), .dinb(n514), .dout(n38728));
  jnot g20706(.din(n38728), .dout(n38729));
  jor  g20707(.dina(n38729), .dinb(n38727), .dout(n38730));
  jand g20708(.dina(n38730), .dinb(n38274), .dout(n38731));
  jxor g20709(.dina(n38266), .dinb(n510), .dout(n38732));
  jnot g20710(.din(n38732), .dout(n38733));
  jor  g20711(.dina(n38733), .dinb(n38731), .dout(n38734));
  jand g20712(.dina(n38734), .dinb(n38268), .dout(n38735));
  jxor g20713(.dina(n38260), .dinb(n396), .dout(n38736));
  jnot g20714(.din(n38736), .dout(n38737));
  jor  g20715(.dina(n38737), .dinb(n38735), .dout(n38738));
  jand g20716(.dina(n38738), .dinb(n38262), .dout(n38739));
  jxor g20717(.dina(n38254), .dinb(n383), .dout(n38740));
  jnot g20718(.din(n38740), .dout(n38741));
  jor  g20719(.dina(n38741), .dinb(n38739), .dout(n38742));
  jand g20720(.dina(n38742), .dinb(n38256), .dout(n38743));
  jxor g20721(.dina(n38248), .dinb(n12211), .dout(n38744));
  jnot g20722(.din(n38744), .dout(n38745));
  jor  g20723(.dina(n38745), .dinb(n38743), .dout(n38746));
  jand g20724(.dina(n38746), .dinb(n38250), .dout(n38747));
  jxor g20725(.dina(n38242), .dinb(n12214), .dout(n38748));
  jnot g20726(.din(n38748), .dout(n38749));
  jor  g20727(.dina(n38749), .dinb(n38747), .dout(n38750));
  jand g20728(.dina(n38750), .dinb(n38244), .dout(n38751));
  jxor g20729(.dina(n38236), .dinb(n384), .dout(n38752));
  jnot g20730(.din(n38752), .dout(n38753));
  jor  g20731(.dina(n38753), .dinb(n38751), .dout(n38754));
  jand g20732(.dina(n38754), .dinb(n38238), .dout(n38755));
  jxor g20733(.dina(n38230), .dinb(n374), .dout(n38756));
  jnot g20734(.din(n38756), .dout(n38757));
  jor  g20735(.dina(n38757), .dinb(n38755), .dout(n38758));
  jand g20736(.dina(n38758), .dinb(n38232), .dout(n38759));
  jxor g20737(.dina(n38224), .dinb(n376), .dout(n38760));
  jnot g20738(.din(n38760), .dout(n38761));
  jor  g20739(.dina(n38761), .dinb(n38759), .dout(n38762));
  jand g20740(.dina(n38762), .dinb(n38226), .dout(n38763));
  jxor g20741(.dina(n38218), .dinb(n377), .dout(n38764));
  jnot g20742(.din(n38764), .dout(n38765));
  jor  g20743(.dina(n38765), .dinb(n38763), .dout(n38766));
  jand g20744(.dina(n38766), .dinb(n38220), .dout(n38767));
  jxor g20745(.dina(n38212), .dinb(n375), .dout(n38768));
  jnot g20746(.din(n38768), .dout(n38769));
  jor  g20747(.dina(n38769), .dinb(n38767), .dout(n38770));
  jand g20748(.dina(n38770), .dinb(n38214), .dout(n38771));
  jand g20749(.dina(n38771), .dinb(n38206), .dout(n38772));
  jor  g20750(.dina(n38772), .dinb(n38204), .dout(n38773));
  jor  g20751(.dina(n38773), .dinb(n38203), .dout(n38774));
  jxor g20752(.dina(n38548), .dinb(b1 ), .dout(n38775));
  jand g20753(.dina(n38775), .dinb(n15383), .dout(n38776));
  jor  g20754(.dina(n38776), .dinb(n38544), .dout(n38777));
  jand g20755(.dina(n38552), .dinb(n38777), .dout(n38778));
  jor  g20756(.dina(n38778), .dinb(n38537), .dout(n38779));
  jand g20757(.dina(n38556), .dinb(n38779), .dout(n38780));
  jor  g20758(.dina(n38780), .dinb(n38531), .dout(n38781));
  jand g20759(.dina(n38560), .dinb(n38781), .dout(n38782));
  jor  g20760(.dina(n38782), .dinb(n38525), .dout(n38783));
  jand g20761(.dina(n38564), .dinb(n38783), .dout(n38784));
  jor  g20762(.dina(n38784), .dinb(n38519), .dout(n38785));
  jand g20763(.dina(n38568), .dinb(n38785), .dout(n38786));
  jor  g20764(.dina(n38786), .dinb(n38513), .dout(n38787));
  jand g20765(.dina(n38572), .dinb(n38787), .dout(n38788));
  jor  g20766(.dina(n38788), .dinb(n38507), .dout(n38789));
  jand g20767(.dina(n38576), .dinb(n38789), .dout(n38790));
  jor  g20768(.dina(n38790), .dinb(n38501), .dout(n38791));
  jand g20769(.dina(n38580), .dinb(n38791), .dout(n38792));
  jor  g20770(.dina(n38792), .dinb(n38495), .dout(n38793));
  jand g20771(.dina(n38584), .dinb(n38793), .dout(n38794));
  jor  g20772(.dina(n38794), .dinb(n38489), .dout(n38795));
  jand g20773(.dina(n38588), .dinb(n38795), .dout(n38796));
  jor  g20774(.dina(n38796), .dinb(n38483), .dout(n38797));
  jand g20775(.dina(n38592), .dinb(n38797), .dout(n38798));
  jor  g20776(.dina(n38798), .dinb(n38477), .dout(n38799));
  jand g20777(.dina(n38596), .dinb(n38799), .dout(n38800));
  jor  g20778(.dina(n38800), .dinb(n38471), .dout(n38801));
  jand g20779(.dina(n38600), .dinb(n38801), .dout(n38802));
  jor  g20780(.dina(n38802), .dinb(n38465), .dout(n38803));
  jand g20781(.dina(n38604), .dinb(n38803), .dout(n38804));
  jor  g20782(.dina(n38804), .dinb(n38459), .dout(n38805));
  jand g20783(.dina(n38608), .dinb(n38805), .dout(n38806));
  jor  g20784(.dina(n38806), .dinb(n38453), .dout(n38807));
  jand g20785(.dina(n38612), .dinb(n38807), .dout(n38808));
  jor  g20786(.dina(n38808), .dinb(n38447), .dout(n38809));
  jand g20787(.dina(n38616), .dinb(n38809), .dout(n38810));
  jor  g20788(.dina(n38810), .dinb(n38441), .dout(n38811));
  jand g20789(.dina(n38620), .dinb(n38811), .dout(n38812));
  jor  g20790(.dina(n38812), .dinb(n38435), .dout(n38813));
  jand g20791(.dina(n38624), .dinb(n38813), .dout(n38814));
  jor  g20792(.dina(n38814), .dinb(n38429), .dout(n38815));
  jand g20793(.dina(n38628), .dinb(n38815), .dout(n38816));
  jor  g20794(.dina(n38816), .dinb(n38423), .dout(n38817));
  jand g20795(.dina(n38632), .dinb(n38817), .dout(n38818));
  jor  g20796(.dina(n38818), .dinb(n38417), .dout(n38819));
  jand g20797(.dina(n38636), .dinb(n38819), .dout(n38820));
  jor  g20798(.dina(n38820), .dinb(n38411), .dout(n38821));
  jand g20799(.dina(n38640), .dinb(n38821), .dout(n38822));
  jor  g20800(.dina(n38822), .dinb(n38405), .dout(n38823));
  jand g20801(.dina(n38644), .dinb(n38823), .dout(n38824));
  jor  g20802(.dina(n38824), .dinb(n38399), .dout(n38825));
  jand g20803(.dina(n38648), .dinb(n38825), .dout(n38826));
  jor  g20804(.dina(n38826), .dinb(n38393), .dout(n38827));
  jand g20805(.dina(n38652), .dinb(n38827), .dout(n38828));
  jor  g20806(.dina(n38828), .dinb(n38387), .dout(n38829));
  jand g20807(.dina(n38656), .dinb(n38829), .dout(n38830));
  jor  g20808(.dina(n38830), .dinb(n38381), .dout(n38831));
  jand g20809(.dina(n38660), .dinb(n38831), .dout(n38832));
  jor  g20810(.dina(n38832), .dinb(n38375), .dout(n38833));
  jand g20811(.dina(n38664), .dinb(n38833), .dout(n38834));
  jor  g20812(.dina(n38834), .dinb(n38369), .dout(n38835));
  jand g20813(.dina(n38668), .dinb(n38835), .dout(n38836));
  jor  g20814(.dina(n38836), .dinb(n38363), .dout(n38837));
  jand g20815(.dina(n38672), .dinb(n38837), .dout(n38838));
  jor  g20816(.dina(n38838), .dinb(n38357), .dout(n38839));
  jand g20817(.dina(n38676), .dinb(n38839), .dout(n38840));
  jor  g20818(.dina(n38840), .dinb(n38351), .dout(n38841));
  jand g20819(.dina(n38680), .dinb(n38841), .dout(n38842));
  jor  g20820(.dina(n38842), .dinb(n38345), .dout(n38843));
  jand g20821(.dina(n38684), .dinb(n38843), .dout(n38844));
  jor  g20822(.dina(n38844), .dinb(n38339), .dout(n38845));
  jand g20823(.dina(n38688), .dinb(n38845), .dout(n38846));
  jor  g20824(.dina(n38846), .dinb(n38333), .dout(n38847));
  jand g20825(.dina(n38692), .dinb(n38847), .dout(n38848));
  jor  g20826(.dina(n38848), .dinb(n38327), .dout(n38849));
  jand g20827(.dina(n38696), .dinb(n38849), .dout(n38850));
  jor  g20828(.dina(n38850), .dinb(n38321), .dout(n38851));
  jand g20829(.dina(n38700), .dinb(n38851), .dout(n38852));
  jor  g20830(.dina(n38852), .dinb(n38315), .dout(n38853));
  jand g20831(.dina(n38704), .dinb(n38853), .dout(n38854));
  jor  g20832(.dina(n38854), .dinb(n38309), .dout(n38855));
  jand g20833(.dina(n38708), .dinb(n38855), .dout(n38856));
  jor  g20834(.dina(n38856), .dinb(n38303), .dout(n38857));
  jand g20835(.dina(n38712), .dinb(n38857), .dout(n38858));
  jor  g20836(.dina(n38858), .dinb(n38297), .dout(n38859));
  jand g20837(.dina(n38716), .dinb(n38859), .dout(n38860));
  jor  g20838(.dina(n38860), .dinb(n38291), .dout(n38861));
  jand g20839(.dina(n38720), .dinb(n38861), .dout(n38862));
  jor  g20840(.dina(n38862), .dinb(n38285), .dout(n38863));
  jand g20841(.dina(n38724), .dinb(n38863), .dout(n38864));
  jor  g20842(.dina(n38864), .dinb(n38279), .dout(n38865));
  jand g20843(.dina(n38728), .dinb(n38865), .dout(n38866));
  jor  g20844(.dina(n38866), .dinb(n38273), .dout(n38867));
  jand g20845(.dina(n38732), .dinb(n38867), .dout(n38868));
  jor  g20846(.dina(n38868), .dinb(n38267), .dout(n38869));
  jand g20847(.dina(n38736), .dinb(n38869), .dout(n38870));
  jor  g20848(.dina(n38870), .dinb(n38261), .dout(n38871));
  jand g20849(.dina(n38740), .dinb(n38871), .dout(n38872));
  jor  g20850(.dina(n38872), .dinb(n38255), .dout(n38873));
  jand g20851(.dina(n38744), .dinb(n38873), .dout(n38874));
  jor  g20852(.dina(n38874), .dinb(n38249), .dout(n38875));
  jand g20853(.dina(n38748), .dinb(n38875), .dout(n38876));
  jor  g20854(.dina(n38876), .dinb(n38243), .dout(n38877));
  jand g20855(.dina(n38752), .dinb(n38877), .dout(n38878));
  jor  g20856(.dina(n38878), .dinb(n38237), .dout(n38879));
  jand g20857(.dina(n38756), .dinb(n38879), .dout(n38880));
  jor  g20858(.dina(n38880), .dinb(n38231), .dout(n38881));
  jand g20859(.dina(n38760), .dinb(n38881), .dout(n38882));
  jor  g20860(.dina(n38882), .dinb(n38225), .dout(n38883));
  jand g20861(.dina(n38764), .dinb(n38883), .dout(n38884));
  jor  g20862(.dina(n38884), .dinb(n38219), .dout(n38885));
  jand g20863(.dina(n38768), .dinb(n38885), .dout(n38886));
  jor  g20864(.dina(n38886), .dinb(n38213), .dout(n38887));
  jand g20865(.dina(n38887), .dinb(n373), .dout(n38888));
  jor  g20866(.dina(n38888), .dinb(n38774), .dout(n38889));
  jand g20867(.dina(n38889), .dinb(n38202), .dout(n38890));
  jand g20868(.dina(n38774), .dinb(n38212), .dout(n38891));
  jnot g20869(.din(n38204), .dout(n38892));
  jor  g20870(.dina(n38887), .dinb(n38205), .dout(n38893));
  jand g20871(.dina(n38893), .dinb(n38892), .dout(n38894));
  jand g20872(.dina(n38894), .dinb(n15090), .dout(n38895));
  jxor g20873(.dina(n38768), .dinb(n38885), .dout(n38896));
  jand g20874(.dina(n38896), .dinb(n38895), .dout(n38897));
  jor  g20875(.dina(n38897), .dinb(n38891), .dout(n38898));
  jand g20876(.dina(n38898), .dinb(n362), .dout(n38899));
  jnot g20877(.din(n38899), .dout(n38900));
  jand g20878(.dina(n38774), .dinb(n38218), .dout(n38901));
  jxor g20879(.dina(n38764), .dinb(n38883), .dout(n38902));
  jand g20880(.dina(n38902), .dinb(n38895), .dout(n38903));
  jor  g20881(.dina(n38903), .dinb(n38901), .dout(n38904));
  jand g20882(.dina(n38904), .dinb(n375), .dout(n38905));
  jnot g20883(.din(n38905), .dout(n38906));
  jand g20884(.dina(n38774), .dinb(n38224), .dout(n38907));
  jxor g20885(.dina(n38760), .dinb(n38881), .dout(n38908));
  jand g20886(.dina(n38908), .dinb(n38895), .dout(n38909));
  jor  g20887(.dina(n38909), .dinb(n38907), .dout(n38910));
  jand g20888(.dina(n38910), .dinb(n377), .dout(n38911));
  jnot g20889(.din(n38911), .dout(n38912));
  jand g20890(.dina(n38774), .dinb(n38230), .dout(n38913));
  jxor g20891(.dina(n38756), .dinb(n38879), .dout(n38914));
  jand g20892(.dina(n38914), .dinb(n38895), .dout(n38915));
  jor  g20893(.dina(n38915), .dinb(n38913), .dout(n38916));
  jand g20894(.dina(n38916), .dinb(n376), .dout(n38917));
  jnot g20895(.din(n38917), .dout(n38918));
  jand g20896(.dina(n38774), .dinb(n38236), .dout(n38919));
  jxor g20897(.dina(n38752), .dinb(n38877), .dout(n38920));
  jand g20898(.dina(n38920), .dinb(n38895), .dout(n38921));
  jor  g20899(.dina(n38921), .dinb(n38919), .dout(n38922));
  jand g20900(.dina(n38922), .dinb(n374), .dout(n38923));
  jnot g20901(.din(n38923), .dout(n38924));
  jand g20902(.dina(n38774), .dinb(n38242), .dout(n38925));
  jxor g20903(.dina(n38748), .dinb(n38875), .dout(n38926));
  jand g20904(.dina(n38926), .dinb(n38895), .dout(n38927));
  jor  g20905(.dina(n38927), .dinb(n38925), .dout(n38928));
  jand g20906(.dina(n38928), .dinb(n384), .dout(n38929));
  jnot g20907(.din(n38929), .dout(n38930));
  jand g20908(.dina(n38774), .dinb(n38248), .dout(n38931));
  jxor g20909(.dina(n38744), .dinb(n38873), .dout(n38932));
  jand g20910(.dina(n38932), .dinb(n38895), .dout(n38933));
  jor  g20911(.dina(n38933), .dinb(n38931), .dout(n38934));
  jand g20912(.dina(n38934), .dinb(n12214), .dout(n38935));
  jnot g20913(.din(n38935), .dout(n38936));
  jand g20914(.dina(n38774), .dinb(n38254), .dout(n38937));
  jxor g20915(.dina(n38740), .dinb(n38871), .dout(n38938));
  jand g20916(.dina(n38938), .dinb(n38895), .dout(n38939));
  jor  g20917(.dina(n38939), .dinb(n38937), .dout(n38940));
  jand g20918(.dina(n38940), .dinb(n12211), .dout(n38941));
  jnot g20919(.din(n38941), .dout(n38942));
  jand g20920(.dina(n38774), .dinb(n38260), .dout(n38943));
  jxor g20921(.dina(n38736), .dinb(n38869), .dout(n38944));
  jand g20922(.dina(n38944), .dinb(n38895), .dout(n38945));
  jor  g20923(.dina(n38945), .dinb(n38943), .dout(n38946));
  jand g20924(.dina(n38946), .dinb(n383), .dout(n38947));
  jnot g20925(.din(n38947), .dout(n38948));
  jand g20926(.dina(n38774), .dinb(n38266), .dout(n38949));
  jxor g20927(.dina(n38732), .dinb(n38867), .dout(n38950));
  jand g20928(.dina(n38950), .dinb(n38895), .dout(n38951));
  jor  g20929(.dina(n38951), .dinb(n38949), .dout(n38952));
  jand g20930(.dina(n38952), .dinb(n396), .dout(n38953));
  jnot g20931(.din(n38953), .dout(n38954));
  jand g20932(.dina(n38774), .dinb(n38272), .dout(n38955));
  jxor g20933(.dina(n38728), .dinb(n38865), .dout(n38956));
  jand g20934(.dina(n38956), .dinb(n38895), .dout(n38957));
  jor  g20935(.dina(n38957), .dinb(n38955), .dout(n38958));
  jand g20936(.dina(n38958), .dinb(n510), .dout(n38959));
  jnot g20937(.din(n38959), .dout(n38960));
  jand g20938(.dina(n38774), .dinb(n38278), .dout(n38961));
  jxor g20939(.dina(n38724), .dinb(n38863), .dout(n38962));
  jand g20940(.dina(n38962), .dinb(n38895), .dout(n38963));
  jor  g20941(.dina(n38963), .dinb(n38961), .dout(n38964));
  jand g20942(.dina(n38964), .dinb(n514), .dout(n38965));
  jnot g20943(.din(n38965), .dout(n38966));
  jand g20944(.dina(n38774), .dinb(n38284), .dout(n38967));
  jxor g20945(.dina(n38720), .dinb(n38861), .dout(n38968));
  jand g20946(.dina(n38968), .dinb(n38895), .dout(n38969));
  jor  g20947(.dina(n38969), .dinb(n38967), .dout(n38970));
  jand g20948(.dina(n38970), .dinb(n513), .dout(n38971));
  jnot g20949(.din(n38971), .dout(n38972));
  jand g20950(.dina(n38774), .dinb(n38290), .dout(n38973));
  jxor g20951(.dina(n38716), .dinb(n38859), .dout(n38974));
  jand g20952(.dina(n38974), .dinb(n38895), .dout(n38975));
  jor  g20953(.dina(n38975), .dinb(n38973), .dout(n38976));
  jand g20954(.dina(n38976), .dinb(n397), .dout(n38977));
  jnot g20955(.din(n38977), .dout(n38978));
  jand g20956(.dina(n38774), .dinb(n38296), .dout(n38979));
  jxor g20957(.dina(n38712), .dinb(n38857), .dout(n38980));
  jand g20958(.dina(n38980), .dinb(n38895), .dout(n38981));
  jor  g20959(.dina(n38981), .dinb(n38979), .dout(n38982));
  jand g20960(.dina(n38982), .dinb(n282), .dout(n38983));
  jnot g20961(.din(n38983), .dout(n38984));
  jand g20962(.dina(n38774), .dinb(n38302), .dout(n38985));
  jxor g20963(.dina(n38708), .dinb(n38855), .dout(n38986));
  jand g20964(.dina(n38986), .dinb(n38895), .dout(n38987));
  jor  g20965(.dina(n38987), .dinb(n38985), .dout(n38988));
  jand g20966(.dina(n38988), .dinb(n281), .dout(n38989));
  jnot g20967(.din(n38989), .dout(n38990));
  jand g20968(.dina(n38774), .dinb(n38308), .dout(n38991));
  jxor g20969(.dina(n38704), .dinb(n38853), .dout(n38992));
  jand g20970(.dina(n38992), .dinb(n38895), .dout(n38993));
  jor  g20971(.dina(n38993), .dinb(n38991), .dout(n38994));
  jand g20972(.dina(n38994), .dinb(n285), .dout(n38995));
  jnot g20973(.din(n38995), .dout(n38996));
  jand g20974(.dina(n38774), .dinb(n38314), .dout(n38997));
  jxor g20975(.dina(n38700), .dinb(n38851), .dout(n38998));
  jand g20976(.dina(n38998), .dinb(n38895), .dout(n38999));
  jor  g20977(.dina(n38999), .dinb(n38997), .dout(n39000));
  jand g20978(.dina(n39000), .dinb(n284), .dout(n39001));
  jnot g20979(.din(n39001), .dout(n39002));
  jand g20980(.dina(n38774), .dinb(n38320), .dout(n39003));
  jxor g20981(.dina(n38696), .dinb(n38849), .dout(n39004));
  jand g20982(.dina(n39004), .dinb(n38895), .dout(n39005));
  jor  g20983(.dina(n39005), .dinb(n39003), .dout(n39006));
  jand g20984(.dina(n39006), .dinb(n291), .dout(n39007));
  jnot g20985(.din(n39007), .dout(n39008));
  jand g20986(.dina(n38774), .dinb(n38326), .dout(n39009));
  jxor g20987(.dina(n38692), .dinb(n38847), .dout(n39010));
  jand g20988(.dina(n39010), .dinb(n38895), .dout(n39011));
  jor  g20989(.dina(n39011), .dinb(n39009), .dout(n39012));
  jand g20990(.dina(n39012), .dinb(n290), .dout(n39013));
  jnot g20991(.din(n39013), .dout(n39014));
  jand g20992(.dina(n38774), .dinb(n38332), .dout(n39015));
  jxor g20993(.dina(n38688), .dinb(n38845), .dout(n39016));
  jand g20994(.dina(n39016), .dinb(n38895), .dout(n39017));
  jor  g20995(.dina(n39017), .dinb(n39015), .dout(n39018));
  jand g20996(.dina(n39018), .dinb(n294), .dout(n39019));
  jnot g20997(.din(n39019), .dout(n39020));
  jand g20998(.dina(n38774), .dinb(n38338), .dout(n39021));
  jxor g20999(.dina(n38684), .dinb(n38843), .dout(n39022));
  jand g21000(.dina(n39022), .dinb(n38895), .dout(n39023));
  jor  g21001(.dina(n39023), .dinb(n39021), .dout(n39024));
  jand g21002(.dina(n39024), .dinb(n293), .dout(n39025));
  jnot g21003(.din(n39025), .dout(n39026));
  jand g21004(.dina(n38774), .dinb(n38344), .dout(n39027));
  jxor g21005(.dina(n38680), .dinb(n38841), .dout(n39028));
  jand g21006(.dina(n39028), .dinb(n38895), .dout(n39029));
  jor  g21007(.dina(n39029), .dinb(n39027), .dout(n39030));
  jand g21008(.dina(n39030), .dinb(n301), .dout(n39031));
  jnot g21009(.din(n39031), .dout(n39032));
  jand g21010(.dina(n38774), .dinb(n38350), .dout(n39033));
  jxor g21011(.dina(n38676), .dinb(n38839), .dout(n39034));
  jand g21012(.dina(n39034), .dinb(n38895), .dout(n39035));
  jor  g21013(.dina(n39035), .dinb(n39033), .dout(n39036));
  jand g21014(.dina(n39036), .dinb(n298), .dout(n39037));
  jnot g21015(.din(n39037), .dout(n39038));
  jand g21016(.dina(n38774), .dinb(n38356), .dout(n39039));
  jxor g21017(.dina(n38672), .dinb(n38837), .dout(n39040));
  jand g21018(.dina(n39040), .dinb(n38895), .dout(n39041));
  jor  g21019(.dina(n39041), .dinb(n39039), .dout(n39042));
  jand g21020(.dina(n39042), .dinb(n297), .dout(n39043));
  jnot g21021(.din(n39043), .dout(n39044));
  jand g21022(.dina(n38774), .dinb(n38362), .dout(n39045));
  jxor g21023(.dina(n38668), .dinb(n38835), .dout(n39046));
  jand g21024(.dina(n39046), .dinb(n38895), .dout(n39047));
  jor  g21025(.dina(n39047), .dinb(n39045), .dout(n39048));
  jand g21026(.dina(n39048), .dinb(n300), .dout(n39049));
  jnot g21027(.din(n39049), .dout(n39050));
  jand g21028(.dina(n38774), .dinb(n38368), .dout(n39051));
  jxor g21029(.dina(n38664), .dinb(n38833), .dout(n39052));
  jand g21030(.dina(n39052), .dinb(n38895), .dout(n39053));
  jor  g21031(.dina(n39053), .dinb(n39051), .dout(n39054));
  jand g21032(.dina(n39054), .dinb(n424), .dout(n39055));
  jnot g21033(.din(n39055), .dout(n39056));
  jand g21034(.dina(n38774), .dinb(n38374), .dout(n39057));
  jxor g21035(.dina(n38660), .dinb(n38831), .dout(n39058));
  jand g21036(.dina(n39058), .dinb(n38895), .dout(n39059));
  jor  g21037(.dina(n39059), .dinb(n39057), .dout(n39060));
  jand g21038(.dina(n39060), .dinb(n427), .dout(n39061));
  jnot g21039(.din(n39061), .dout(n39062));
  jand g21040(.dina(n38774), .dinb(n38380), .dout(n39063));
  jxor g21041(.dina(n38656), .dinb(n38829), .dout(n39064));
  jand g21042(.dina(n39064), .dinb(n38895), .dout(n39065));
  jor  g21043(.dina(n39065), .dinb(n39063), .dout(n39066));
  jand g21044(.dina(n39066), .dinb(n426), .dout(n39067));
  jnot g21045(.din(n39067), .dout(n39068));
  jand g21046(.dina(n38774), .dinb(n38386), .dout(n39069));
  jxor g21047(.dina(n38652), .dinb(n38827), .dout(n39070));
  jand g21048(.dina(n39070), .dinb(n38895), .dout(n39071));
  jor  g21049(.dina(n39071), .dinb(n39069), .dout(n39072));
  jand g21050(.dina(n39072), .dinb(n410), .dout(n39073));
  jnot g21051(.din(n39073), .dout(n39074));
  jand g21052(.dina(n38774), .dinb(n38392), .dout(n39075));
  jxor g21053(.dina(n38648), .dinb(n38825), .dout(n39076));
  jand g21054(.dina(n39076), .dinb(n38895), .dout(n39077));
  jor  g21055(.dina(n39077), .dinb(n39075), .dout(n39078));
  jand g21056(.dina(n39078), .dinb(n409), .dout(n39079));
  jnot g21057(.din(n39079), .dout(n39080));
  jand g21058(.dina(n38774), .dinb(n38398), .dout(n39081));
  jxor g21059(.dina(n38644), .dinb(n38823), .dout(n39082));
  jand g21060(.dina(n39082), .dinb(n38895), .dout(n39083));
  jor  g21061(.dina(n39083), .dinb(n39081), .dout(n39084));
  jand g21062(.dina(n39084), .dinb(n413), .dout(n39085));
  jnot g21063(.din(n39085), .dout(n39086));
  jand g21064(.dina(n38774), .dinb(n38404), .dout(n39087));
  jxor g21065(.dina(n38640), .dinb(n38821), .dout(n39088));
  jand g21066(.dina(n39088), .dinb(n38895), .dout(n39089));
  jor  g21067(.dina(n39089), .dinb(n39087), .dout(n39090));
  jand g21068(.dina(n39090), .dinb(n412), .dout(n39091));
  jnot g21069(.din(n39091), .dout(n39092));
  jand g21070(.dina(n38774), .dinb(n38410), .dout(n39093));
  jxor g21071(.dina(n38636), .dinb(n38819), .dout(n39094));
  jand g21072(.dina(n39094), .dinb(n38895), .dout(n39095));
  jor  g21073(.dina(n39095), .dinb(n39093), .dout(n39096));
  jand g21074(.dina(n39096), .dinb(n406), .dout(n39097));
  jnot g21075(.din(n39097), .dout(n39098));
  jand g21076(.dina(n38774), .dinb(n38416), .dout(n39099));
  jxor g21077(.dina(n38632), .dinb(n38817), .dout(n39100));
  jand g21078(.dina(n39100), .dinb(n38895), .dout(n39101));
  jor  g21079(.dina(n39101), .dinb(n39099), .dout(n39102));
  jand g21080(.dina(n39102), .dinb(n405), .dout(n39103));
  jnot g21081(.din(n39103), .dout(n39104));
  jand g21082(.dina(n38774), .dinb(n38422), .dout(n39105));
  jxor g21083(.dina(n38628), .dinb(n38815), .dout(n39106));
  jand g21084(.dina(n39106), .dinb(n38895), .dout(n39107));
  jor  g21085(.dina(n39107), .dinb(n39105), .dout(n39108));
  jand g21086(.dina(n39108), .dinb(n2714), .dout(n39109));
  jnot g21087(.din(n39109), .dout(n39110));
  jand g21088(.dina(n38774), .dinb(n38428), .dout(n39111));
  jxor g21089(.dina(n38624), .dinb(n38813), .dout(n39112));
  jand g21090(.dina(n39112), .dinb(n38895), .dout(n39113));
  jor  g21091(.dina(n39113), .dinb(n39111), .dout(n39114));
  jand g21092(.dina(n39114), .dinb(n2547), .dout(n39115));
  jnot g21093(.din(n39115), .dout(n39116));
  jand g21094(.dina(n38774), .dinb(n38434), .dout(n39117));
  jxor g21095(.dina(n38620), .dinb(n38811), .dout(n39118));
  jand g21096(.dina(n39118), .dinb(n38895), .dout(n39119));
  jor  g21097(.dina(n39119), .dinb(n39117), .dout(n39120));
  jand g21098(.dina(n39120), .dinb(n417), .dout(n39121));
  jnot g21099(.din(n39121), .dout(n39122));
  jand g21100(.dina(n38774), .dinb(n38440), .dout(n39123));
  jxor g21101(.dina(n38616), .dinb(n38809), .dout(n39124));
  jand g21102(.dina(n39124), .dinb(n38895), .dout(n39125));
  jor  g21103(.dina(n39125), .dinb(n39123), .dout(n39126));
  jand g21104(.dina(n39126), .dinb(n416), .dout(n39127));
  jnot g21105(.din(n39127), .dout(n39128));
  jand g21106(.dina(n38774), .dinb(n38446), .dout(n39129));
  jxor g21107(.dina(n38612), .dinb(n38807), .dout(n39130));
  jand g21108(.dina(n39130), .dinb(n38895), .dout(n39131));
  jor  g21109(.dina(n39131), .dinb(n39129), .dout(n39132));
  jand g21110(.dina(n39132), .dinb(n422), .dout(n39133));
  jnot g21111(.din(n39133), .dout(n39134));
  jand g21112(.dina(n38774), .dinb(n38452), .dout(n39135));
  jxor g21113(.dina(n38608), .dinb(n38805), .dout(n39136));
  jand g21114(.dina(n39136), .dinb(n38895), .dout(n39137));
  jor  g21115(.dina(n39137), .dinb(n39135), .dout(n39138));
  jand g21116(.dina(n39138), .dinb(n421), .dout(n39139));
  jnot g21117(.din(n39139), .dout(n39140));
  jand g21118(.dina(n38774), .dinb(n38458), .dout(n39141));
  jxor g21119(.dina(n38604), .dinb(n38803), .dout(n39142));
  jand g21120(.dina(n39142), .dinb(n38895), .dout(n39143));
  jor  g21121(.dina(n39143), .dinb(n39141), .dout(n39144));
  jand g21122(.dina(n39144), .dinb(n433), .dout(n39145));
  jnot g21123(.din(n39145), .dout(n39146));
  jand g21124(.dina(n38774), .dinb(n38464), .dout(n39147));
  jxor g21125(.dina(n38600), .dinb(n38801), .dout(n39148));
  jand g21126(.dina(n39148), .dinb(n38895), .dout(n39149));
  jor  g21127(.dina(n39149), .dinb(n39147), .dout(n39150));
  jand g21128(.dina(n39150), .dinb(n432), .dout(n39151));
  jnot g21129(.din(n39151), .dout(n39152));
  jand g21130(.dina(n38774), .dinb(n38470), .dout(n39153));
  jxor g21131(.dina(n38596), .dinb(n38799), .dout(n39154));
  jand g21132(.dina(n39154), .dinb(n38895), .dout(n39155));
  jor  g21133(.dina(n39155), .dinb(n39153), .dout(n39156));
  jand g21134(.dina(n39156), .dinb(n436), .dout(n39157));
  jnot g21135(.din(n39157), .dout(n39158));
  jand g21136(.dina(n38774), .dinb(n38476), .dout(n39159));
  jxor g21137(.dina(n38592), .dinb(n38797), .dout(n39160));
  jand g21138(.dina(n39160), .dinb(n38895), .dout(n39161));
  jor  g21139(.dina(n39161), .dinb(n39159), .dout(n39162));
  jand g21140(.dina(n39162), .dinb(n435), .dout(n39163));
  jnot g21141(.din(n39163), .dout(n39164));
  jand g21142(.dina(n38774), .dinb(n38482), .dout(n39165));
  jxor g21143(.dina(n38588), .dinb(n38795), .dout(n39166));
  jand g21144(.dina(n39166), .dinb(n38895), .dout(n39167));
  jor  g21145(.dina(n39167), .dinb(n39165), .dout(n39168));
  jand g21146(.dina(n39168), .dinb(n440), .dout(n39169));
  jnot g21147(.din(n39169), .dout(n39170));
  jand g21148(.dina(n38774), .dinb(n38488), .dout(n39171));
  jxor g21149(.dina(n38584), .dinb(n38793), .dout(n39172));
  jand g21150(.dina(n39172), .dinb(n38895), .dout(n39173));
  jor  g21151(.dina(n39173), .dinb(n39171), .dout(n39174));
  jand g21152(.dina(n39174), .dinb(n439), .dout(n39175));
  jnot g21153(.din(n39175), .dout(n39176));
  jand g21154(.dina(n38774), .dinb(n38494), .dout(n39177));
  jxor g21155(.dina(n38580), .dinb(n38791), .dout(n39178));
  jand g21156(.dina(n39178), .dinb(n38895), .dout(n39179));
  jor  g21157(.dina(n39179), .dinb(n39177), .dout(n39180));
  jand g21158(.dina(n39180), .dinb(n325), .dout(n39181));
  jnot g21159(.din(n39181), .dout(n39182));
  jand g21160(.dina(n38774), .dinb(n38500), .dout(n39183));
  jxor g21161(.dina(n38576), .dinb(n38789), .dout(n39184));
  jand g21162(.dina(n39184), .dinb(n38895), .dout(n39185));
  jor  g21163(.dina(n39185), .dinb(n39183), .dout(n39186));
  jand g21164(.dina(n39186), .dinb(n324), .dout(n39187));
  jnot g21165(.din(n39187), .dout(n39188));
  jand g21166(.dina(n38774), .dinb(n38506), .dout(n39189));
  jxor g21167(.dina(n38572), .dinb(n38787), .dout(n39190));
  jand g21168(.dina(n39190), .dinb(n38895), .dout(n39191));
  jor  g21169(.dina(n39191), .dinb(n39189), .dout(n39192));
  jand g21170(.dina(n39192), .dinb(n323), .dout(n39193));
  jnot g21171(.din(n39193), .dout(n39194));
  jand g21172(.dina(n38774), .dinb(n38512), .dout(n39195));
  jxor g21173(.dina(n38568), .dinb(n38785), .dout(n39196));
  jand g21174(.dina(n39196), .dinb(n38895), .dout(n39197));
  jor  g21175(.dina(n39197), .dinb(n39195), .dout(n39198));
  jand g21176(.dina(n39198), .dinb(n335), .dout(n39199));
  jnot g21177(.din(n39199), .dout(n39200));
  jand g21178(.dina(n38774), .dinb(n38518), .dout(n39201));
  jxor g21179(.dina(n38564), .dinb(n38783), .dout(n39202));
  jand g21180(.dina(n39202), .dinb(n38895), .dout(n39203));
  jor  g21181(.dina(n39203), .dinb(n39201), .dout(n39204));
  jand g21182(.dina(n39204), .dinb(n334), .dout(n39205));
  jnot g21183(.din(n39205), .dout(n39206));
  jand g21184(.dina(n38774), .dinb(n38524), .dout(n39207));
  jxor g21185(.dina(n38560), .dinb(n38781), .dout(n39208));
  jand g21186(.dina(n39208), .dinb(n38895), .dout(n39209));
  jor  g21187(.dina(n39209), .dinb(n39207), .dout(n39210));
  jand g21188(.dina(n39210), .dinb(n338), .dout(n39211));
  jnot g21189(.din(n39211), .dout(n39212));
  jand g21190(.dina(n38774), .dinb(n38530), .dout(n39213));
  jxor g21191(.dina(n38556), .dinb(n38779), .dout(n39214));
  jand g21192(.dina(n39214), .dinb(n38895), .dout(n39215));
  jor  g21193(.dina(n39215), .dinb(n39213), .dout(n39216));
  jand g21194(.dina(n39216), .dinb(n337), .dout(n39217));
  jnot g21195(.din(n39217), .dout(n39218));
  jand g21196(.dina(n38774), .dinb(n38536), .dout(n39219));
  jxor g21197(.dina(n38552), .dinb(n38777), .dout(n39220));
  jand g21198(.dina(n39220), .dinb(n38895), .dout(n39221));
  jor  g21199(.dina(n39221), .dinb(n39219), .dout(n39222));
  jand g21200(.dina(n39222), .dinb(n344), .dout(n39223));
  jnot g21201(.din(n39223), .dout(n39224));
  jor  g21202(.dina(n38895), .dinb(n38548), .dout(n39225));
  jxor g21203(.dina(n38775), .dinb(n15383), .dout(n39226));
  jnot g21204(.din(n39226), .dout(n39227));
  jor  g21205(.dina(n39227), .dinb(n38774), .dout(n39228));
  jand g21206(.dina(n39228), .dinb(n39225), .dout(n39229));
  jnot g21207(.din(n39229), .dout(n39230));
  jand g21208(.dina(n39230), .dinb(n348), .dout(n39231));
  jnot g21209(.din(n39231), .dout(n39232));
  jand g21210(.dina(n38894), .dinb(n15840), .dout(n39233));
  jxor g21211(.dina(n39233), .dinb(a6 ), .dout(n39234));
  jand g21212(.dina(n39234), .dinb(n258), .dout(n39235));
  jnot g21213(.din(n39235), .dout(n39236));
  jxor g21214(.dina(n39233), .dinb(n15381), .dout(n39237));
  jxor g21215(.dina(n39237), .dinb(n258), .dout(n39238));
  jor  g21216(.dina(n39238), .dinb(n15846), .dout(n39239));
  jand g21217(.dina(n39239), .dinb(n39236), .dout(n39240));
  jxor g21218(.dina(n39229), .dinb(b2 ), .dout(n39241));
  jnot g21219(.din(n39241), .dout(n39242));
  jor  g21220(.dina(n39242), .dinb(n39240), .dout(n39243));
  jand g21221(.dina(n39243), .dinb(n39232), .dout(n39244));
  jxor g21222(.dina(n39222), .dinb(n344), .dout(n39245));
  jnot g21223(.din(n39245), .dout(n39246));
  jor  g21224(.dina(n39246), .dinb(n39244), .dout(n39247));
  jand g21225(.dina(n39247), .dinb(n39224), .dout(n39248));
  jxor g21226(.dina(n39216), .dinb(n337), .dout(n39249));
  jnot g21227(.din(n39249), .dout(n39250));
  jor  g21228(.dina(n39250), .dinb(n39248), .dout(n39251));
  jand g21229(.dina(n39251), .dinb(n39218), .dout(n39252));
  jxor g21230(.dina(n39210), .dinb(n338), .dout(n39253));
  jnot g21231(.din(n39253), .dout(n39254));
  jor  g21232(.dina(n39254), .dinb(n39252), .dout(n39255));
  jand g21233(.dina(n39255), .dinb(n39212), .dout(n39256));
  jxor g21234(.dina(n39204), .dinb(n334), .dout(n39257));
  jnot g21235(.din(n39257), .dout(n39258));
  jor  g21236(.dina(n39258), .dinb(n39256), .dout(n39259));
  jand g21237(.dina(n39259), .dinb(n39206), .dout(n39260));
  jxor g21238(.dina(n39198), .dinb(n335), .dout(n39261));
  jnot g21239(.din(n39261), .dout(n39262));
  jor  g21240(.dina(n39262), .dinb(n39260), .dout(n39263));
  jand g21241(.dina(n39263), .dinb(n39200), .dout(n39264));
  jxor g21242(.dina(n39192), .dinb(n323), .dout(n39265));
  jnot g21243(.din(n39265), .dout(n39266));
  jor  g21244(.dina(n39266), .dinb(n39264), .dout(n39267));
  jand g21245(.dina(n39267), .dinb(n39194), .dout(n39268));
  jxor g21246(.dina(n39186), .dinb(n324), .dout(n39269));
  jnot g21247(.din(n39269), .dout(n39270));
  jor  g21248(.dina(n39270), .dinb(n39268), .dout(n39271));
  jand g21249(.dina(n39271), .dinb(n39188), .dout(n39272));
  jxor g21250(.dina(n39180), .dinb(n325), .dout(n39273));
  jnot g21251(.din(n39273), .dout(n39274));
  jor  g21252(.dina(n39274), .dinb(n39272), .dout(n39275));
  jand g21253(.dina(n39275), .dinb(n39182), .dout(n39276));
  jxor g21254(.dina(n39174), .dinb(n439), .dout(n39277));
  jnot g21255(.din(n39277), .dout(n39278));
  jor  g21256(.dina(n39278), .dinb(n39276), .dout(n39279));
  jand g21257(.dina(n39279), .dinb(n39176), .dout(n39280));
  jxor g21258(.dina(n39168), .dinb(n440), .dout(n39281));
  jnot g21259(.din(n39281), .dout(n39282));
  jor  g21260(.dina(n39282), .dinb(n39280), .dout(n39283));
  jand g21261(.dina(n39283), .dinb(n39170), .dout(n39284));
  jxor g21262(.dina(n39162), .dinb(n435), .dout(n39285));
  jnot g21263(.din(n39285), .dout(n39286));
  jor  g21264(.dina(n39286), .dinb(n39284), .dout(n39287));
  jand g21265(.dina(n39287), .dinb(n39164), .dout(n39288));
  jxor g21266(.dina(n39156), .dinb(n436), .dout(n39289));
  jnot g21267(.din(n39289), .dout(n39290));
  jor  g21268(.dina(n39290), .dinb(n39288), .dout(n39291));
  jand g21269(.dina(n39291), .dinb(n39158), .dout(n39292));
  jxor g21270(.dina(n39150), .dinb(n432), .dout(n39293));
  jnot g21271(.din(n39293), .dout(n39294));
  jor  g21272(.dina(n39294), .dinb(n39292), .dout(n39295));
  jand g21273(.dina(n39295), .dinb(n39152), .dout(n39296));
  jxor g21274(.dina(n39144), .dinb(n433), .dout(n39297));
  jnot g21275(.din(n39297), .dout(n39298));
  jor  g21276(.dina(n39298), .dinb(n39296), .dout(n39299));
  jand g21277(.dina(n39299), .dinb(n39146), .dout(n39300));
  jxor g21278(.dina(n39138), .dinb(n421), .dout(n39301));
  jnot g21279(.din(n39301), .dout(n39302));
  jor  g21280(.dina(n39302), .dinb(n39300), .dout(n39303));
  jand g21281(.dina(n39303), .dinb(n39140), .dout(n39304));
  jxor g21282(.dina(n39132), .dinb(n422), .dout(n39305));
  jnot g21283(.din(n39305), .dout(n39306));
  jor  g21284(.dina(n39306), .dinb(n39304), .dout(n39307));
  jand g21285(.dina(n39307), .dinb(n39134), .dout(n39308));
  jxor g21286(.dina(n39126), .dinb(n416), .dout(n39309));
  jnot g21287(.din(n39309), .dout(n39310));
  jor  g21288(.dina(n39310), .dinb(n39308), .dout(n39311));
  jand g21289(.dina(n39311), .dinb(n39128), .dout(n39312));
  jxor g21290(.dina(n39120), .dinb(n417), .dout(n39313));
  jnot g21291(.din(n39313), .dout(n39314));
  jor  g21292(.dina(n39314), .dinb(n39312), .dout(n39315));
  jand g21293(.dina(n39315), .dinb(n39122), .dout(n39316));
  jxor g21294(.dina(n39114), .dinb(n2547), .dout(n39317));
  jnot g21295(.din(n39317), .dout(n39318));
  jor  g21296(.dina(n39318), .dinb(n39316), .dout(n39319));
  jand g21297(.dina(n39319), .dinb(n39116), .dout(n39320));
  jxor g21298(.dina(n39108), .dinb(n2714), .dout(n39321));
  jnot g21299(.din(n39321), .dout(n39322));
  jor  g21300(.dina(n39322), .dinb(n39320), .dout(n39323));
  jand g21301(.dina(n39323), .dinb(n39110), .dout(n39324));
  jxor g21302(.dina(n39102), .dinb(n405), .dout(n39325));
  jnot g21303(.din(n39325), .dout(n39326));
  jor  g21304(.dina(n39326), .dinb(n39324), .dout(n39327));
  jand g21305(.dina(n39327), .dinb(n39104), .dout(n39328));
  jxor g21306(.dina(n39096), .dinb(n406), .dout(n39329));
  jnot g21307(.din(n39329), .dout(n39330));
  jor  g21308(.dina(n39330), .dinb(n39328), .dout(n39331));
  jand g21309(.dina(n39331), .dinb(n39098), .dout(n39332));
  jxor g21310(.dina(n39090), .dinb(n412), .dout(n39333));
  jnot g21311(.din(n39333), .dout(n39334));
  jor  g21312(.dina(n39334), .dinb(n39332), .dout(n39335));
  jand g21313(.dina(n39335), .dinb(n39092), .dout(n39336));
  jxor g21314(.dina(n39084), .dinb(n413), .dout(n39337));
  jnot g21315(.din(n39337), .dout(n39338));
  jor  g21316(.dina(n39338), .dinb(n39336), .dout(n39339));
  jand g21317(.dina(n39339), .dinb(n39086), .dout(n39340));
  jxor g21318(.dina(n39078), .dinb(n409), .dout(n39341));
  jnot g21319(.din(n39341), .dout(n39342));
  jor  g21320(.dina(n39342), .dinb(n39340), .dout(n39343));
  jand g21321(.dina(n39343), .dinb(n39080), .dout(n39344));
  jxor g21322(.dina(n39072), .dinb(n410), .dout(n39345));
  jnot g21323(.din(n39345), .dout(n39346));
  jor  g21324(.dina(n39346), .dinb(n39344), .dout(n39347));
  jand g21325(.dina(n39347), .dinb(n39074), .dout(n39348));
  jxor g21326(.dina(n39066), .dinb(n426), .dout(n39349));
  jnot g21327(.din(n39349), .dout(n39350));
  jor  g21328(.dina(n39350), .dinb(n39348), .dout(n39351));
  jand g21329(.dina(n39351), .dinb(n39068), .dout(n39352));
  jxor g21330(.dina(n39060), .dinb(n427), .dout(n39353));
  jnot g21331(.din(n39353), .dout(n39354));
  jor  g21332(.dina(n39354), .dinb(n39352), .dout(n39355));
  jand g21333(.dina(n39355), .dinb(n39062), .dout(n39356));
  jxor g21334(.dina(n39054), .dinb(n424), .dout(n39357));
  jnot g21335(.din(n39357), .dout(n39358));
  jor  g21336(.dina(n39358), .dinb(n39356), .dout(n39359));
  jand g21337(.dina(n39359), .dinb(n39056), .dout(n39360));
  jxor g21338(.dina(n39048), .dinb(n300), .dout(n39361));
  jnot g21339(.din(n39361), .dout(n39362));
  jor  g21340(.dina(n39362), .dinb(n39360), .dout(n39363));
  jand g21341(.dina(n39363), .dinb(n39050), .dout(n39364));
  jxor g21342(.dina(n39042), .dinb(n297), .dout(n39365));
  jnot g21343(.din(n39365), .dout(n39366));
  jor  g21344(.dina(n39366), .dinb(n39364), .dout(n39367));
  jand g21345(.dina(n39367), .dinb(n39044), .dout(n39368));
  jxor g21346(.dina(n39036), .dinb(n298), .dout(n39369));
  jnot g21347(.din(n39369), .dout(n39370));
  jor  g21348(.dina(n39370), .dinb(n39368), .dout(n39371));
  jand g21349(.dina(n39371), .dinb(n39038), .dout(n39372));
  jxor g21350(.dina(n39030), .dinb(n301), .dout(n39373));
  jnot g21351(.din(n39373), .dout(n39374));
  jor  g21352(.dina(n39374), .dinb(n39372), .dout(n39375));
  jand g21353(.dina(n39375), .dinb(n39032), .dout(n39376));
  jxor g21354(.dina(n39024), .dinb(n293), .dout(n39377));
  jnot g21355(.din(n39377), .dout(n39378));
  jor  g21356(.dina(n39378), .dinb(n39376), .dout(n39379));
  jand g21357(.dina(n39379), .dinb(n39026), .dout(n39380));
  jxor g21358(.dina(n39018), .dinb(n294), .dout(n39381));
  jnot g21359(.din(n39381), .dout(n39382));
  jor  g21360(.dina(n39382), .dinb(n39380), .dout(n39383));
  jand g21361(.dina(n39383), .dinb(n39020), .dout(n39384));
  jxor g21362(.dina(n39012), .dinb(n290), .dout(n39385));
  jnot g21363(.din(n39385), .dout(n39386));
  jor  g21364(.dina(n39386), .dinb(n39384), .dout(n39387));
  jand g21365(.dina(n39387), .dinb(n39014), .dout(n39388));
  jxor g21366(.dina(n39006), .dinb(n291), .dout(n39389));
  jnot g21367(.din(n39389), .dout(n39390));
  jor  g21368(.dina(n39390), .dinb(n39388), .dout(n39391));
  jand g21369(.dina(n39391), .dinb(n39008), .dout(n39392));
  jxor g21370(.dina(n39000), .dinb(n284), .dout(n39393));
  jnot g21371(.din(n39393), .dout(n39394));
  jor  g21372(.dina(n39394), .dinb(n39392), .dout(n39395));
  jand g21373(.dina(n39395), .dinb(n39002), .dout(n39396));
  jxor g21374(.dina(n38994), .dinb(n285), .dout(n39397));
  jnot g21375(.din(n39397), .dout(n39398));
  jor  g21376(.dina(n39398), .dinb(n39396), .dout(n39399));
  jand g21377(.dina(n39399), .dinb(n38996), .dout(n39400));
  jxor g21378(.dina(n38988), .dinb(n281), .dout(n39401));
  jnot g21379(.din(n39401), .dout(n39402));
  jor  g21380(.dina(n39402), .dinb(n39400), .dout(n39403));
  jand g21381(.dina(n39403), .dinb(n38990), .dout(n39404));
  jxor g21382(.dina(n38982), .dinb(n282), .dout(n39405));
  jnot g21383(.din(n39405), .dout(n39406));
  jor  g21384(.dina(n39406), .dinb(n39404), .dout(n39407));
  jand g21385(.dina(n39407), .dinb(n38984), .dout(n39408));
  jxor g21386(.dina(n38976), .dinb(n397), .dout(n39409));
  jnot g21387(.din(n39409), .dout(n39410));
  jor  g21388(.dina(n39410), .dinb(n39408), .dout(n39411));
  jand g21389(.dina(n39411), .dinb(n38978), .dout(n39412));
  jxor g21390(.dina(n38970), .dinb(n513), .dout(n39413));
  jnot g21391(.din(n39413), .dout(n39414));
  jor  g21392(.dina(n39414), .dinb(n39412), .dout(n39415));
  jand g21393(.dina(n39415), .dinb(n38972), .dout(n39416));
  jxor g21394(.dina(n38964), .dinb(n514), .dout(n39417));
  jnot g21395(.din(n39417), .dout(n39418));
  jor  g21396(.dina(n39418), .dinb(n39416), .dout(n39419));
  jand g21397(.dina(n39419), .dinb(n38966), .dout(n39420));
  jxor g21398(.dina(n38958), .dinb(n510), .dout(n39421));
  jnot g21399(.din(n39421), .dout(n39422));
  jor  g21400(.dina(n39422), .dinb(n39420), .dout(n39423));
  jand g21401(.dina(n39423), .dinb(n38960), .dout(n39424));
  jxor g21402(.dina(n38952), .dinb(n396), .dout(n39425));
  jnot g21403(.din(n39425), .dout(n39426));
  jor  g21404(.dina(n39426), .dinb(n39424), .dout(n39427));
  jand g21405(.dina(n39427), .dinb(n38954), .dout(n39428));
  jxor g21406(.dina(n38946), .dinb(n383), .dout(n39429));
  jnot g21407(.din(n39429), .dout(n39430));
  jor  g21408(.dina(n39430), .dinb(n39428), .dout(n39431));
  jand g21409(.dina(n39431), .dinb(n38948), .dout(n39432));
  jxor g21410(.dina(n38940), .dinb(n12211), .dout(n39433));
  jnot g21411(.din(n39433), .dout(n39434));
  jor  g21412(.dina(n39434), .dinb(n39432), .dout(n39435));
  jand g21413(.dina(n39435), .dinb(n38942), .dout(n39436));
  jxor g21414(.dina(n38934), .dinb(n12214), .dout(n39437));
  jnot g21415(.din(n39437), .dout(n39438));
  jor  g21416(.dina(n39438), .dinb(n39436), .dout(n39439));
  jand g21417(.dina(n39439), .dinb(n38936), .dout(n39440));
  jxor g21418(.dina(n38928), .dinb(n384), .dout(n39441));
  jnot g21419(.din(n39441), .dout(n39442));
  jor  g21420(.dina(n39442), .dinb(n39440), .dout(n39443));
  jand g21421(.dina(n39443), .dinb(n38930), .dout(n39444));
  jxor g21422(.dina(n38922), .dinb(n374), .dout(n39445));
  jnot g21423(.din(n39445), .dout(n39446));
  jor  g21424(.dina(n39446), .dinb(n39444), .dout(n39447));
  jand g21425(.dina(n39447), .dinb(n38924), .dout(n39448));
  jxor g21426(.dina(n38916), .dinb(n376), .dout(n39449));
  jnot g21427(.din(n39449), .dout(n39450));
  jor  g21428(.dina(n39450), .dinb(n39448), .dout(n39451));
  jand g21429(.dina(n39451), .dinb(n38918), .dout(n39452));
  jxor g21430(.dina(n38910), .dinb(n377), .dout(n39453));
  jnot g21431(.din(n39453), .dout(n39454));
  jor  g21432(.dina(n39454), .dinb(n39452), .dout(n39455));
  jand g21433(.dina(n39455), .dinb(n38912), .dout(n39456));
  jxor g21434(.dina(n38904), .dinb(n375), .dout(n39457));
  jnot g21435(.din(n39457), .dout(n39458));
  jor  g21436(.dina(n39458), .dinb(n39456), .dout(n39459));
  jand g21437(.dina(n39459), .dinb(n38906), .dout(n39460));
  jxor g21438(.dina(n38898), .dinb(n362), .dout(n39461));
  jnot g21439(.din(n39461), .dout(n39462));
  jor  g21440(.dina(n39462), .dinb(n39460), .dout(n39463));
  jand g21441(.dina(n39463), .dinb(n38900), .dout(n39464));
  jand g21442(.dina(n38890), .dinb(n363), .dout(n39465));
  jnot g21443(.din(n39465), .dout(n39466));
  jand g21444(.dina(n39466), .dinb(n39464), .dout(n39467));
  jnot g21445(.din(n38890), .dout(n39468));
  jand g21446(.dina(n39468), .dinb(b58 ), .dout(n39469));
  jor  g21447(.dina(n39469), .dinb(n16024), .dout(n39470));
  jor  g21448(.dina(n39470), .dinb(n39467), .dout(n39471));
  jxor g21449(.dina(n39237), .dinb(b1 ), .dout(n39472));
  jand g21450(.dina(n39472), .dinb(n15847), .dout(n39473));
  jor  g21451(.dina(n39473), .dinb(n39235), .dout(n39474));
  jand g21452(.dina(n39241), .dinb(n39474), .dout(n39475));
  jor  g21453(.dina(n39475), .dinb(n39231), .dout(n39476));
  jand g21454(.dina(n39245), .dinb(n39476), .dout(n39477));
  jor  g21455(.dina(n39477), .dinb(n39223), .dout(n39478));
  jand g21456(.dina(n39249), .dinb(n39478), .dout(n39479));
  jor  g21457(.dina(n39479), .dinb(n39217), .dout(n39480));
  jand g21458(.dina(n39253), .dinb(n39480), .dout(n39481));
  jor  g21459(.dina(n39481), .dinb(n39211), .dout(n39482));
  jand g21460(.dina(n39257), .dinb(n39482), .dout(n39483));
  jor  g21461(.dina(n39483), .dinb(n39205), .dout(n39484));
  jand g21462(.dina(n39261), .dinb(n39484), .dout(n39485));
  jor  g21463(.dina(n39485), .dinb(n39199), .dout(n39486));
  jand g21464(.dina(n39265), .dinb(n39486), .dout(n39487));
  jor  g21465(.dina(n39487), .dinb(n39193), .dout(n39488));
  jand g21466(.dina(n39269), .dinb(n39488), .dout(n39489));
  jor  g21467(.dina(n39489), .dinb(n39187), .dout(n39490));
  jand g21468(.dina(n39273), .dinb(n39490), .dout(n39491));
  jor  g21469(.dina(n39491), .dinb(n39181), .dout(n39492));
  jand g21470(.dina(n39277), .dinb(n39492), .dout(n39493));
  jor  g21471(.dina(n39493), .dinb(n39175), .dout(n39494));
  jand g21472(.dina(n39281), .dinb(n39494), .dout(n39495));
  jor  g21473(.dina(n39495), .dinb(n39169), .dout(n39496));
  jand g21474(.dina(n39285), .dinb(n39496), .dout(n39497));
  jor  g21475(.dina(n39497), .dinb(n39163), .dout(n39498));
  jand g21476(.dina(n39289), .dinb(n39498), .dout(n39499));
  jor  g21477(.dina(n39499), .dinb(n39157), .dout(n39500));
  jand g21478(.dina(n39293), .dinb(n39500), .dout(n39501));
  jor  g21479(.dina(n39501), .dinb(n39151), .dout(n39502));
  jand g21480(.dina(n39297), .dinb(n39502), .dout(n39503));
  jor  g21481(.dina(n39503), .dinb(n39145), .dout(n39504));
  jand g21482(.dina(n39301), .dinb(n39504), .dout(n39505));
  jor  g21483(.dina(n39505), .dinb(n39139), .dout(n39506));
  jand g21484(.dina(n39305), .dinb(n39506), .dout(n39507));
  jor  g21485(.dina(n39507), .dinb(n39133), .dout(n39508));
  jand g21486(.dina(n39309), .dinb(n39508), .dout(n39509));
  jor  g21487(.dina(n39509), .dinb(n39127), .dout(n39510));
  jand g21488(.dina(n39313), .dinb(n39510), .dout(n39511));
  jor  g21489(.dina(n39511), .dinb(n39121), .dout(n39512));
  jand g21490(.dina(n39317), .dinb(n39512), .dout(n39513));
  jor  g21491(.dina(n39513), .dinb(n39115), .dout(n39514));
  jand g21492(.dina(n39321), .dinb(n39514), .dout(n39515));
  jor  g21493(.dina(n39515), .dinb(n39109), .dout(n39516));
  jand g21494(.dina(n39325), .dinb(n39516), .dout(n39517));
  jor  g21495(.dina(n39517), .dinb(n39103), .dout(n39518));
  jand g21496(.dina(n39329), .dinb(n39518), .dout(n39519));
  jor  g21497(.dina(n39519), .dinb(n39097), .dout(n39520));
  jand g21498(.dina(n39333), .dinb(n39520), .dout(n39521));
  jor  g21499(.dina(n39521), .dinb(n39091), .dout(n39522));
  jand g21500(.dina(n39337), .dinb(n39522), .dout(n39523));
  jor  g21501(.dina(n39523), .dinb(n39085), .dout(n39524));
  jand g21502(.dina(n39341), .dinb(n39524), .dout(n39525));
  jor  g21503(.dina(n39525), .dinb(n39079), .dout(n39526));
  jand g21504(.dina(n39345), .dinb(n39526), .dout(n39527));
  jor  g21505(.dina(n39527), .dinb(n39073), .dout(n39528));
  jand g21506(.dina(n39349), .dinb(n39528), .dout(n39529));
  jor  g21507(.dina(n39529), .dinb(n39067), .dout(n39530));
  jand g21508(.dina(n39353), .dinb(n39530), .dout(n39531));
  jor  g21509(.dina(n39531), .dinb(n39061), .dout(n39532));
  jand g21510(.dina(n39357), .dinb(n39532), .dout(n39533));
  jor  g21511(.dina(n39533), .dinb(n39055), .dout(n39534));
  jand g21512(.dina(n39361), .dinb(n39534), .dout(n39535));
  jor  g21513(.dina(n39535), .dinb(n39049), .dout(n39536));
  jand g21514(.dina(n39365), .dinb(n39536), .dout(n39537));
  jor  g21515(.dina(n39537), .dinb(n39043), .dout(n39538));
  jand g21516(.dina(n39369), .dinb(n39538), .dout(n39539));
  jor  g21517(.dina(n39539), .dinb(n39037), .dout(n39540));
  jand g21518(.dina(n39373), .dinb(n39540), .dout(n39541));
  jor  g21519(.dina(n39541), .dinb(n39031), .dout(n39542));
  jand g21520(.dina(n39377), .dinb(n39542), .dout(n39543));
  jor  g21521(.dina(n39543), .dinb(n39025), .dout(n39544));
  jand g21522(.dina(n39381), .dinb(n39544), .dout(n39545));
  jor  g21523(.dina(n39545), .dinb(n39019), .dout(n39546));
  jand g21524(.dina(n39385), .dinb(n39546), .dout(n39547));
  jor  g21525(.dina(n39547), .dinb(n39013), .dout(n39548));
  jand g21526(.dina(n39389), .dinb(n39548), .dout(n39549));
  jor  g21527(.dina(n39549), .dinb(n39007), .dout(n39550));
  jand g21528(.dina(n39393), .dinb(n39550), .dout(n39551));
  jor  g21529(.dina(n39551), .dinb(n39001), .dout(n39552));
  jand g21530(.dina(n39397), .dinb(n39552), .dout(n39553));
  jor  g21531(.dina(n39553), .dinb(n38995), .dout(n39554));
  jand g21532(.dina(n39401), .dinb(n39554), .dout(n39555));
  jor  g21533(.dina(n39555), .dinb(n38989), .dout(n39556));
  jand g21534(.dina(n39405), .dinb(n39556), .dout(n39557));
  jor  g21535(.dina(n39557), .dinb(n38983), .dout(n39558));
  jand g21536(.dina(n39409), .dinb(n39558), .dout(n39559));
  jor  g21537(.dina(n39559), .dinb(n38977), .dout(n39560));
  jand g21538(.dina(n39413), .dinb(n39560), .dout(n39561));
  jor  g21539(.dina(n39561), .dinb(n38971), .dout(n39562));
  jand g21540(.dina(n39417), .dinb(n39562), .dout(n39563));
  jor  g21541(.dina(n39563), .dinb(n38965), .dout(n39564));
  jand g21542(.dina(n39421), .dinb(n39564), .dout(n39565));
  jor  g21543(.dina(n39565), .dinb(n38959), .dout(n39566));
  jand g21544(.dina(n39425), .dinb(n39566), .dout(n39567));
  jor  g21545(.dina(n39567), .dinb(n38953), .dout(n39568));
  jand g21546(.dina(n39429), .dinb(n39568), .dout(n39569));
  jor  g21547(.dina(n39569), .dinb(n38947), .dout(n39570));
  jand g21548(.dina(n39433), .dinb(n39570), .dout(n39571));
  jor  g21549(.dina(n39571), .dinb(n38941), .dout(n39572));
  jand g21550(.dina(n39437), .dinb(n39572), .dout(n39573));
  jor  g21551(.dina(n39573), .dinb(n38935), .dout(n39574));
  jand g21552(.dina(n39441), .dinb(n39574), .dout(n39575));
  jor  g21553(.dina(n39575), .dinb(n38929), .dout(n39576));
  jand g21554(.dina(n39445), .dinb(n39576), .dout(n39577));
  jor  g21555(.dina(n39577), .dinb(n38923), .dout(n39578));
  jand g21556(.dina(n39449), .dinb(n39578), .dout(n39579));
  jor  g21557(.dina(n39579), .dinb(n38917), .dout(n39580));
  jand g21558(.dina(n39453), .dinb(n39580), .dout(n39581));
  jor  g21559(.dina(n39581), .dinb(n38911), .dout(n39582));
  jand g21560(.dina(n39457), .dinb(n39582), .dout(n39583));
  jor  g21561(.dina(n39583), .dinb(n38905), .dout(n39584));
  jand g21562(.dina(n39461), .dinb(n39584), .dout(n39585));
  jor  g21563(.dina(n39585), .dinb(n38899), .dout(n39586));
  jand g21564(.dina(n39586), .dinb(n15090), .dout(n39587));
  jor  g21565(.dina(n39587), .dinb(n39471), .dout(n39588));
  jand g21566(.dina(n39588), .dinb(n38890), .dout(n39589));
  jand g21567(.dina(n39471), .dinb(n38898), .dout(n39590));
  jor  g21568(.dina(n39465), .dinb(n39586), .dout(n39591));
  jnot g21569(.din(n39470), .dout(n39592));
  jand g21570(.dina(n39592), .dinb(n39591), .dout(n39593));
  jxor g21571(.dina(n39461), .dinb(n39584), .dout(n39594));
  jand g21572(.dina(n39594), .dinb(n39593), .dout(n39595));
  jor  g21573(.dina(n39595), .dinb(n39590), .dout(n39596));
  jand g21574(.dina(n39596), .dinb(n363), .dout(n39597));
  jnot g21575(.din(n39597), .dout(n39598));
  jand g21576(.dina(n39471), .dinb(n38904), .dout(n39599));
  jxor g21577(.dina(n39457), .dinb(n39582), .dout(n39600));
  jand g21578(.dina(n39600), .dinb(n39593), .dout(n39601));
  jor  g21579(.dina(n39601), .dinb(n39599), .dout(n39602));
  jand g21580(.dina(n39602), .dinb(n362), .dout(n39603));
  jnot g21581(.din(n39603), .dout(n39604));
  jand g21582(.dina(n39471), .dinb(n38910), .dout(n39605));
  jxor g21583(.dina(n39453), .dinb(n39580), .dout(n39606));
  jand g21584(.dina(n39606), .dinb(n39593), .dout(n39607));
  jor  g21585(.dina(n39607), .dinb(n39605), .dout(n39608));
  jand g21586(.dina(n39608), .dinb(n375), .dout(n39609));
  jnot g21587(.din(n39609), .dout(n39610));
  jand g21588(.dina(n39471), .dinb(n38916), .dout(n39611));
  jxor g21589(.dina(n39449), .dinb(n39578), .dout(n39612));
  jand g21590(.dina(n39612), .dinb(n39593), .dout(n39613));
  jor  g21591(.dina(n39613), .dinb(n39611), .dout(n39614));
  jand g21592(.dina(n39614), .dinb(n377), .dout(n39615));
  jnot g21593(.din(n39615), .dout(n39616));
  jand g21594(.dina(n39471), .dinb(n38922), .dout(n39617));
  jxor g21595(.dina(n39445), .dinb(n39576), .dout(n39618));
  jand g21596(.dina(n39618), .dinb(n39593), .dout(n39619));
  jor  g21597(.dina(n39619), .dinb(n39617), .dout(n39620));
  jand g21598(.dina(n39620), .dinb(n376), .dout(n39621));
  jnot g21599(.din(n39621), .dout(n39622));
  jand g21600(.dina(n39471), .dinb(n38928), .dout(n39623));
  jxor g21601(.dina(n39441), .dinb(n39574), .dout(n39624));
  jand g21602(.dina(n39624), .dinb(n39593), .dout(n39625));
  jor  g21603(.dina(n39625), .dinb(n39623), .dout(n39626));
  jand g21604(.dina(n39626), .dinb(n374), .dout(n39627));
  jnot g21605(.din(n39627), .dout(n39628));
  jand g21606(.dina(n39471), .dinb(n38934), .dout(n39629));
  jxor g21607(.dina(n39437), .dinb(n39572), .dout(n39630));
  jand g21608(.dina(n39630), .dinb(n39593), .dout(n39631));
  jor  g21609(.dina(n39631), .dinb(n39629), .dout(n39632));
  jand g21610(.dina(n39632), .dinb(n384), .dout(n39633));
  jnot g21611(.din(n39633), .dout(n39634));
  jand g21612(.dina(n39471), .dinb(n38940), .dout(n39635));
  jxor g21613(.dina(n39433), .dinb(n39570), .dout(n39636));
  jand g21614(.dina(n39636), .dinb(n39593), .dout(n39637));
  jor  g21615(.dina(n39637), .dinb(n39635), .dout(n39638));
  jand g21616(.dina(n39638), .dinb(n12214), .dout(n39639));
  jnot g21617(.din(n39639), .dout(n39640));
  jand g21618(.dina(n39471), .dinb(n38946), .dout(n39641));
  jxor g21619(.dina(n39429), .dinb(n39568), .dout(n39642));
  jand g21620(.dina(n39642), .dinb(n39593), .dout(n39643));
  jor  g21621(.dina(n39643), .dinb(n39641), .dout(n39644));
  jand g21622(.dina(n39644), .dinb(n12211), .dout(n39645));
  jnot g21623(.din(n39645), .dout(n39646));
  jand g21624(.dina(n39471), .dinb(n38952), .dout(n39647));
  jxor g21625(.dina(n39425), .dinb(n39566), .dout(n39648));
  jand g21626(.dina(n39648), .dinb(n39593), .dout(n39649));
  jor  g21627(.dina(n39649), .dinb(n39647), .dout(n39650));
  jand g21628(.dina(n39650), .dinb(n383), .dout(n39651));
  jnot g21629(.din(n39651), .dout(n39652));
  jand g21630(.dina(n39471), .dinb(n38958), .dout(n39653));
  jxor g21631(.dina(n39421), .dinb(n39564), .dout(n39654));
  jand g21632(.dina(n39654), .dinb(n39593), .dout(n39655));
  jor  g21633(.dina(n39655), .dinb(n39653), .dout(n39656));
  jand g21634(.dina(n39656), .dinb(n396), .dout(n39657));
  jnot g21635(.din(n39657), .dout(n39658));
  jand g21636(.dina(n39471), .dinb(n38964), .dout(n39659));
  jxor g21637(.dina(n39417), .dinb(n39562), .dout(n39660));
  jand g21638(.dina(n39660), .dinb(n39593), .dout(n39661));
  jor  g21639(.dina(n39661), .dinb(n39659), .dout(n39662));
  jand g21640(.dina(n39662), .dinb(n510), .dout(n39663));
  jnot g21641(.din(n39663), .dout(n39664));
  jand g21642(.dina(n39471), .dinb(n38970), .dout(n39665));
  jxor g21643(.dina(n39413), .dinb(n39560), .dout(n39666));
  jand g21644(.dina(n39666), .dinb(n39593), .dout(n39667));
  jor  g21645(.dina(n39667), .dinb(n39665), .dout(n39668));
  jand g21646(.dina(n39668), .dinb(n514), .dout(n39669));
  jnot g21647(.din(n39669), .dout(n39670));
  jand g21648(.dina(n39471), .dinb(n38976), .dout(n39671));
  jxor g21649(.dina(n39409), .dinb(n39558), .dout(n39672));
  jand g21650(.dina(n39672), .dinb(n39593), .dout(n39673));
  jor  g21651(.dina(n39673), .dinb(n39671), .dout(n39674));
  jand g21652(.dina(n39674), .dinb(n513), .dout(n39675));
  jnot g21653(.din(n39675), .dout(n39676));
  jand g21654(.dina(n39471), .dinb(n38982), .dout(n39677));
  jxor g21655(.dina(n39405), .dinb(n39556), .dout(n39678));
  jand g21656(.dina(n39678), .dinb(n39593), .dout(n39679));
  jor  g21657(.dina(n39679), .dinb(n39677), .dout(n39680));
  jand g21658(.dina(n39680), .dinb(n397), .dout(n39681));
  jnot g21659(.din(n39681), .dout(n39682));
  jand g21660(.dina(n39471), .dinb(n38988), .dout(n39683));
  jxor g21661(.dina(n39401), .dinb(n39554), .dout(n39684));
  jand g21662(.dina(n39684), .dinb(n39593), .dout(n39685));
  jor  g21663(.dina(n39685), .dinb(n39683), .dout(n39686));
  jand g21664(.dina(n39686), .dinb(n282), .dout(n39687));
  jnot g21665(.din(n39687), .dout(n39688));
  jand g21666(.dina(n39471), .dinb(n38994), .dout(n39689));
  jxor g21667(.dina(n39397), .dinb(n39552), .dout(n39690));
  jand g21668(.dina(n39690), .dinb(n39593), .dout(n39691));
  jor  g21669(.dina(n39691), .dinb(n39689), .dout(n39692));
  jand g21670(.dina(n39692), .dinb(n281), .dout(n39693));
  jnot g21671(.din(n39693), .dout(n39694));
  jand g21672(.dina(n39471), .dinb(n39000), .dout(n39695));
  jxor g21673(.dina(n39393), .dinb(n39550), .dout(n39696));
  jand g21674(.dina(n39696), .dinb(n39593), .dout(n39697));
  jor  g21675(.dina(n39697), .dinb(n39695), .dout(n39698));
  jand g21676(.dina(n39698), .dinb(n285), .dout(n39699));
  jnot g21677(.din(n39699), .dout(n39700));
  jand g21678(.dina(n39471), .dinb(n39006), .dout(n39701));
  jxor g21679(.dina(n39389), .dinb(n39548), .dout(n39702));
  jand g21680(.dina(n39702), .dinb(n39593), .dout(n39703));
  jor  g21681(.dina(n39703), .dinb(n39701), .dout(n39704));
  jand g21682(.dina(n39704), .dinb(n284), .dout(n39705));
  jnot g21683(.din(n39705), .dout(n39706));
  jand g21684(.dina(n39471), .dinb(n39012), .dout(n39707));
  jxor g21685(.dina(n39385), .dinb(n39546), .dout(n39708));
  jand g21686(.dina(n39708), .dinb(n39593), .dout(n39709));
  jor  g21687(.dina(n39709), .dinb(n39707), .dout(n39710));
  jand g21688(.dina(n39710), .dinb(n291), .dout(n39711));
  jnot g21689(.din(n39711), .dout(n39712));
  jand g21690(.dina(n39471), .dinb(n39018), .dout(n39713));
  jxor g21691(.dina(n39381), .dinb(n39544), .dout(n39714));
  jand g21692(.dina(n39714), .dinb(n39593), .dout(n39715));
  jor  g21693(.dina(n39715), .dinb(n39713), .dout(n39716));
  jand g21694(.dina(n39716), .dinb(n290), .dout(n39717));
  jnot g21695(.din(n39717), .dout(n39718));
  jand g21696(.dina(n39471), .dinb(n39024), .dout(n39719));
  jxor g21697(.dina(n39377), .dinb(n39542), .dout(n39720));
  jand g21698(.dina(n39720), .dinb(n39593), .dout(n39721));
  jor  g21699(.dina(n39721), .dinb(n39719), .dout(n39722));
  jand g21700(.dina(n39722), .dinb(n294), .dout(n39723));
  jnot g21701(.din(n39723), .dout(n39724));
  jand g21702(.dina(n39471), .dinb(n39030), .dout(n39725));
  jxor g21703(.dina(n39373), .dinb(n39540), .dout(n39726));
  jand g21704(.dina(n39726), .dinb(n39593), .dout(n39727));
  jor  g21705(.dina(n39727), .dinb(n39725), .dout(n39728));
  jand g21706(.dina(n39728), .dinb(n293), .dout(n39729));
  jnot g21707(.din(n39729), .dout(n39730));
  jand g21708(.dina(n39471), .dinb(n39036), .dout(n39731));
  jxor g21709(.dina(n39369), .dinb(n39538), .dout(n39732));
  jand g21710(.dina(n39732), .dinb(n39593), .dout(n39733));
  jor  g21711(.dina(n39733), .dinb(n39731), .dout(n39734));
  jand g21712(.dina(n39734), .dinb(n301), .dout(n39735));
  jnot g21713(.din(n39735), .dout(n39736));
  jand g21714(.dina(n39471), .dinb(n39042), .dout(n39737));
  jxor g21715(.dina(n39365), .dinb(n39536), .dout(n39738));
  jand g21716(.dina(n39738), .dinb(n39593), .dout(n39739));
  jor  g21717(.dina(n39739), .dinb(n39737), .dout(n39740));
  jand g21718(.dina(n39740), .dinb(n298), .dout(n39741));
  jnot g21719(.din(n39741), .dout(n39742));
  jand g21720(.dina(n39471), .dinb(n39048), .dout(n39743));
  jxor g21721(.dina(n39361), .dinb(n39534), .dout(n39744));
  jand g21722(.dina(n39744), .dinb(n39593), .dout(n39745));
  jor  g21723(.dina(n39745), .dinb(n39743), .dout(n39746));
  jand g21724(.dina(n39746), .dinb(n297), .dout(n39747));
  jnot g21725(.din(n39747), .dout(n39748));
  jand g21726(.dina(n39471), .dinb(n39054), .dout(n39749));
  jxor g21727(.dina(n39357), .dinb(n39532), .dout(n39750));
  jand g21728(.dina(n39750), .dinb(n39593), .dout(n39751));
  jor  g21729(.dina(n39751), .dinb(n39749), .dout(n39752));
  jand g21730(.dina(n39752), .dinb(n300), .dout(n39753));
  jnot g21731(.din(n39753), .dout(n39754));
  jand g21732(.dina(n39471), .dinb(n39060), .dout(n39755));
  jxor g21733(.dina(n39353), .dinb(n39530), .dout(n39756));
  jand g21734(.dina(n39756), .dinb(n39593), .dout(n39757));
  jor  g21735(.dina(n39757), .dinb(n39755), .dout(n39758));
  jand g21736(.dina(n39758), .dinb(n424), .dout(n39759));
  jnot g21737(.din(n39759), .dout(n39760));
  jand g21738(.dina(n39471), .dinb(n39066), .dout(n39761));
  jxor g21739(.dina(n39349), .dinb(n39528), .dout(n39762));
  jand g21740(.dina(n39762), .dinb(n39593), .dout(n39763));
  jor  g21741(.dina(n39763), .dinb(n39761), .dout(n39764));
  jand g21742(.dina(n39764), .dinb(n427), .dout(n39765));
  jnot g21743(.din(n39765), .dout(n39766));
  jand g21744(.dina(n39471), .dinb(n39072), .dout(n39767));
  jxor g21745(.dina(n39345), .dinb(n39526), .dout(n39768));
  jand g21746(.dina(n39768), .dinb(n39593), .dout(n39769));
  jor  g21747(.dina(n39769), .dinb(n39767), .dout(n39770));
  jand g21748(.dina(n39770), .dinb(n426), .dout(n39771));
  jnot g21749(.din(n39771), .dout(n39772));
  jand g21750(.dina(n39471), .dinb(n39078), .dout(n39773));
  jxor g21751(.dina(n39341), .dinb(n39524), .dout(n39774));
  jand g21752(.dina(n39774), .dinb(n39593), .dout(n39775));
  jor  g21753(.dina(n39775), .dinb(n39773), .dout(n39776));
  jand g21754(.dina(n39776), .dinb(n410), .dout(n39777));
  jnot g21755(.din(n39777), .dout(n39778));
  jand g21756(.dina(n39471), .dinb(n39084), .dout(n39779));
  jxor g21757(.dina(n39337), .dinb(n39522), .dout(n39780));
  jand g21758(.dina(n39780), .dinb(n39593), .dout(n39781));
  jor  g21759(.dina(n39781), .dinb(n39779), .dout(n39782));
  jand g21760(.dina(n39782), .dinb(n409), .dout(n39783));
  jnot g21761(.din(n39783), .dout(n39784));
  jand g21762(.dina(n39471), .dinb(n39090), .dout(n39785));
  jxor g21763(.dina(n39333), .dinb(n39520), .dout(n39786));
  jand g21764(.dina(n39786), .dinb(n39593), .dout(n39787));
  jor  g21765(.dina(n39787), .dinb(n39785), .dout(n39788));
  jand g21766(.dina(n39788), .dinb(n413), .dout(n39789));
  jnot g21767(.din(n39789), .dout(n39790));
  jand g21768(.dina(n39471), .dinb(n39096), .dout(n39791));
  jxor g21769(.dina(n39329), .dinb(n39518), .dout(n39792));
  jand g21770(.dina(n39792), .dinb(n39593), .dout(n39793));
  jor  g21771(.dina(n39793), .dinb(n39791), .dout(n39794));
  jand g21772(.dina(n39794), .dinb(n412), .dout(n39795));
  jnot g21773(.din(n39795), .dout(n39796));
  jand g21774(.dina(n39471), .dinb(n39102), .dout(n39797));
  jxor g21775(.dina(n39325), .dinb(n39516), .dout(n39798));
  jand g21776(.dina(n39798), .dinb(n39593), .dout(n39799));
  jor  g21777(.dina(n39799), .dinb(n39797), .dout(n39800));
  jand g21778(.dina(n39800), .dinb(n406), .dout(n39801));
  jnot g21779(.din(n39801), .dout(n39802));
  jand g21780(.dina(n39471), .dinb(n39108), .dout(n39803));
  jxor g21781(.dina(n39321), .dinb(n39514), .dout(n39804));
  jand g21782(.dina(n39804), .dinb(n39593), .dout(n39805));
  jor  g21783(.dina(n39805), .dinb(n39803), .dout(n39806));
  jand g21784(.dina(n39806), .dinb(n405), .dout(n39807));
  jnot g21785(.din(n39807), .dout(n39808));
  jand g21786(.dina(n39471), .dinb(n39114), .dout(n39809));
  jxor g21787(.dina(n39317), .dinb(n39512), .dout(n39810));
  jand g21788(.dina(n39810), .dinb(n39593), .dout(n39811));
  jor  g21789(.dina(n39811), .dinb(n39809), .dout(n39812));
  jand g21790(.dina(n39812), .dinb(n2714), .dout(n39813));
  jnot g21791(.din(n39813), .dout(n39814));
  jand g21792(.dina(n39471), .dinb(n39120), .dout(n39815));
  jxor g21793(.dina(n39313), .dinb(n39510), .dout(n39816));
  jand g21794(.dina(n39816), .dinb(n39593), .dout(n39817));
  jor  g21795(.dina(n39817), .dinb(n39815), .dout(n39818));
  jand g21796(.dina(n39818), .dinb(n2547), .dout(n39819));
  jnot g21797(.din(n39819), .dout(n39820));
  jand g21798(.dina(n39471), .dinb(n39126), .dout(n39821));
  jxor g21799(.dina(n39309), .dinb(n39508), .dout(n39822));
  jand g21800(.dina(n39822), .dinb(n39593), .dout(n39823));
  jor  g21801(.dina(n39823), .dinb(n39821), .dout(n39824));
  jand g21802(.dina(n39824), .dinb(n417), .dout(n39825));
  jnot g21803(.din(n39825), .dout(n39826));
  jand g21804(.dina(n39471), .dinb(n39132), .dout(n39827));
  jxor g21805(.dina(n39305), .dinb(n39506), .dout(n39828));
  jand g21806(.dina(n39828), .dinb(n39593), .dout(n39829));
  jor  g21807(.dina(n39829), .dinb(n39827), .dout(n39830));
  jand g21808(.dina(n39830), .dinb(n416), .dout(n39831));
  jnot g21809(.din(n39831), .dout(n39832));
  jand g21810(.dina(n39471), .dinb(n39138), .dout(n39833));
  jxor g21811(.dina(n39301), .dinb(n39504), .dout(n39834));
  jand g21812(.dina(n39834), .dinb(n39593), .dout(n39835));
  jor  g21813(.dina(n39835), .dinb(n39833), .dout(n39836));
  jand g21814(.dina(n39836), .dinb(n422), .dout(n39837));
  jnot g21815(.din(n39837), .dout(n39838));
  jand g21816(.dina(n39471), .dinb(n39144), .dout(n39839));
  jxor g21817(.dina(n39297), .dinb(n39502), .dout(n39840));
  jand g21818(.dina(n39840), .dinb(n39593), .dout(n39841));
  jor  g21819(.dina(n39841), .dinb(n39839), .dout(n39842));
  jand g21820(.dina(n39842), .dinb(n421), .dout(n39843));
  jnot g21821(.din(n39843), .dout(n39844));
  jand g21822(.dina(n39471), .dinb(n39150), .dout(n39845));
  jxor g21823(.dina(n39293), .dinb(n39500), .dout(n39846));
  jand g21824(.dina(n39846), .dinb(n39593), .dout(n39847));
  jor  g21825(.dina(n39847), .dinb(n39845), .dout(n39848));
  jand g21826(.dina(n39848), .dinb(n433), .dout(n39849));
  jnot g21827(.din(n39849), .dout(n39850));
  jand g21828(.dina(n39471), .dinb(n39156), .dout(n39851));
  jxor g21829(.dina(n39289), .dinb(n39498), .dout(n39852));
  jand g21830(.dina(n39852), .dinb(n39593), .dout(n39853));
  jor  g21831(.dina(n39853), .dinb(n39851), .dout(n39854));
  jand g21832(.dina(n39854), .dinb(n432), .dout(n39855));
  jnot g21833(.din(n39855), .dout(n39856));
  jand g21834(.dina(n39471), .dinb(n39162), .dout(n39857));
  jxor g21835(.dina(n39285), .dinb(n39496), .dout(n39858));
  jand g21836(.dina(n39858), .dinb(n39593), .dout(n39859));
  jor  g21837(.dina(n39859), .dinb(n39857), .dout(n39860));
  jand g21838(.dina(n39860), .dinb(n436), .dout(n39861));
  jnot g21839(.din(n39861), .dout(n39862));
  jand g21840(.dina(n39471), .dinb(n39168), .dout(n39863));
  jxor g21841(.dina(n39281), .dinb(n39494), .dout(n39864));
  jand g21842(.dina(n39864), .dinb(n39593), .dout(n39865));
  jor  g21843(.dina(n39865), .dinb(n39863), .dout(n39866));
  jand g21844(.dina(n39866), .dinb(n435), .dout(n39867));
  jnot g21845(.din(n39867), .dout(n39868));
  jand g21846(.dina(n39471), .dinb(n39174), .dout(n39869));
  jxor g21847(.dina(n39277), .dinb(n39492), .dout(n39870));
  jand g21848(.dina(n39870), .dinb(n39593), .dout(n39871));
  jor  g21849(.dina(n39871), .dinb(n39869), .dout(n39872));
  jand g21850(.dina(n39872), .dinb(n440), .dout(n39873));
  jnot g21851(.din(n39873), .dout(n39874));
  jand g21852(.dina(n39471), .dinb(n39180), .dout(n39875));
  jxor g21853(.dina(n39273), .dinb(n39490), .dout(n39876));
  jand g21854(.dina(n39876), .dinb(n39593), .dout(n39877));
  jor  g21855(.dina(n39877), .dinb(n39875), .dout(n39878));
  jand g21856(.dina(n39878), .dinb(n439), .dout(n39879));
  jnot g21857(.din(n39879), .dout(n39880));
  jand g21858(.dina(n39471), .dinb(n39186), .dout(n39881));
  jxor g21859(.dina(n39269), .dinb(n39488), .dout(n39882));
  jand g21860(.dina(n39882), .dinb(n39593), .dout(n39883));
  jor  g21861(.dina(n39883), .dinb(n39881), .dout(n39884));
  jand g21862(.dina(n39884), .dinb(n325), .dout(n39885));
  jnot g21863(.din(n39885), .dout(n39886));
  jand g21864(.dina(n39471), .dinb(n39192), .dout(n39887));
  jxor g21865(.dina(n39265), .dinb(n39486), .dout(n39888));
  jand g21866(.dina(n39888), .dinb(n39593), .dout(n39889));
  jor  g21867(.dina(n39889), .dinb(n39887), .dout(n39890));
  jand g21868(.dina(n39890), .dinb(n324), .dout(n39891));
  jnot g21869(.din(n39891), .dout(n39892));
  jand g21870(.dina(n39471), .dinb(n39198), .dout(n39893));
  jxor g21871(.dina(n39261), .dinb(n39484), .dout(n39894));
  jand g21872(.dina(n39894), .dinb(n39593), .dout(n39895));
  jor  g21873(.dina(n39895), .dinb(n39893), .dout(n39896));
  jand g21874(.dina(n39896), .dinb(n323), .dout(n39897));
  jnot g21875(.din(n39897), .dout(n39898));
  jand g21876(.dina(n39471), .dinb(n39204), .dout(n39899));
  jxor g21877(.dina(n39257), .dinb(n39482), .dout(n39900));
  jand g21878(.dina(n39900), .dinb(n39593), .dout(n39901));
  jor  g21879(.dina(n39901), .dinb(n39899), .dout(n39902));
  jand g21880(.dina(n39902), .dinb(n335), .dout(n39903));
  jnot g21881(.din(n39903), .dout(n39904));
  jand g21882(.dina(n39471), .dinb(n39210), .dout(n39905));
  jxor g21883(.dina(n39253), .dinb(n39480), .dout(n39906));
  jand g21884(.dina(n39906), .dinb(n39593), .dout(n39907));
  jor  g21885(.dina(n39907), .dinb(n39905), .dout(n39908));
  jand g21886(.dina(n39908), .dinb(n334), .dout(n39909));
  jnot g21887(.din(n39909), .dout(n39910));
  jand g21888(.dina(n39471), .dinb(n39216), .dout(n39911));
  jxor g21889(.dina(n39249), .dinb(n39478), .dout(n39912));
  jand g21890(.dina(n39912), .dinb(n39593), .dout(n39913));
  jor  g21891(.dina(n39913), .dinb(n39911), .dout(n39914));
  jand g21892(.dina(n39914), .dinb(n338), .dout(n39915));
  jnot g21893(.din(n39915), .dout(n39916));
  jand g21894(.dina(n39471), .dinb(n39222), .dout(n39917));
  jxor g21895(.dina(n39245), .dinb(n39476), .dout(n39918));
  jand g21896(.dina(n39918), .dinb(n39593), .dout(n39919));
  jor  g21897(.dina(n39919), .dinb(n39917), .dout(n39920));
  jand g21898(.dina(n39920), .dinb(n337), .dout(n39921));
  jnot g21899(.din(n39921), .dout(n39922));
  jand g21900(.dina(n39471), .dinb(n39230), .dout(n39923));
  jxor g21901(.dina(n39241), .dinb(n39474), .dout(n39924));
  jand g21902(.dina(n39924), .dinb(n39593), .dout(n39925));
  jor  g21903(.dina(n39925), .dinb(n39923), .dout(n39926));
  jand g21904(.dina(n39926), .dinb(n344), .dout(n39927));
  jnot g21905(.din(n39927), .dout(n39928));
  jand g21906(.dina(n39471), .dinb(n39234), .dout(n39929));
  jxor g21907(.dina(n39472), .dinb(n15847), .dout(n39930));
  jand g21908(.dina(n39930), .dinb(n39593), .dout(n39931));
  jor  g21909(.dina(n39931), .dinb(n39929), .dout(n39932));
  jand g21910(.dina(n39932), .dinb(n348), .dout(n39933));
  jnot g21911(.din(n39933), .dout(n39934));
  jor  g21912(.dina(n39471), .dinb(n18364), .dout(n39935));
  jand g21913(.dina(n39935), .dinb(a5 ), .dout(n39936));
  jor  g21914(.dina(n39471), .dinb(n15847), .dout(n39937));
  jnot g21915(.din(n39937), .dout(n39938));
  jor  g21916(.dina(n39938), .dinb(n39936), .dout(n39939));
  jand g21917(.dina(n39939), .dinb(n258), .dout(n39940));
  jnot g21918(.din(n39940), .dout(n39941));
  jand g21919(.dina(n39593), .dinb(b0 ), .dout(n39942));
  jor  g21920(.dina(n39942), .dinb(n15845), .dout(n39943));
  jand g21921(.dina(n39937), .dinb(n39943), .dout(n39944));
  jxor g21922(.dina(n39944), .dinb(n258), .dout(n39945));
  jor  g21923(.dina(n39945), .dinb(n16326), .dout(n39946));
  jand g21924(.dina(n39946), .dinb(n39941), .dout(n39947));
  jxor g21925(.dina(n39932), .dinb(n348), .dout(n39948));
  jnot g21926(.din(n39948), .dout(n39949));
  jor  g21927(.dina(n39949), .dinb(n39947), .dout(n39950));
  jand g21928(.dina(n39950), .dinb(n39934), .dout(n39951));
  jxor g21929(.dina(n39926), .dinb(n344), .dout(n39952));
  jnot g21930(.din(n39952), .dout(n39953));
  jor  g21931(.dina(n39953), .dinb(n39951), .dout(n39954));
  jand g21932(.dina(n39954), .dinb(n39928), .dout(n39955));
  jxor g21933(.dina(n39920), .dinb(n337), .dout(n39956));
  jnot g21934(.din(n39956), .dout(n39957));
  jor  g21935(.dina(n39957), .dinb(n39955), .dout(n39958));
  jand g21936(.dina(n39958), .dinb(n39922), .dout(n39959));
  jxor g21937(.dina(n39914), .dinb(n338), .dout(n39960));
  jnot g21938(.din(n39960), .dout(n39961));
  jor  g21939(.dina(n39961), .dinb(n39959), .dout(n39962));
  jand g21940(.dina(n39962), .dinb(n39916), .dout(n39963));
  jxor g21941(.dina(n39908), .dinb(n334), .dout(n39964));
  jnot g21942(.din(n39964), .dout(n39965));
  jor  g21943(.dina(n39965), .dinb(n39963), .dout(n39966));
  jand g21944(.dina(n39966), .dinb(n39910), .dout(n39967));
  jxor g21945(.dina(n39902), .dinb(n335), .dout(n39968));
  jnot g21946(.din(n39968), .dout(n39969));
  jor  g21947(.dina(n39969), .dinb(n39967), .dout(n39970));
  jand g21948(.dina(n39970), .dinb(n39904), .dout(n39971));
  jxor g21949(.dina(n39896), .dinb(n323), .dout(n39972));
  jnot g21950(.din(n39972), .dout(n39973));
  jor  g21951(.dina(n39973), .dinb(n39971), .dout(n39974));
  jand g21952(.dina(n39974), .dinb(n39898), .dout(n39975));
  jxor g21953(.dina(n39890), .dinb(n324), .dout(n39976));
  jnot g21954(.din(n39976), .dout(n39977));
  jor  g21955(.dina(n39977), .dinb(n39975), .dout(n39978));
  jand g21956(.dina(n39978), .dinb(n39892), .dout(n39979));
  jxor g21957(.dina(n39884), .dinb(n325), .dout(n39980));
  jnot g21958(.din(n39980), .dout(n39981));
  jor  g21959(.dina(n39981), .dinb(n39979), .dout(n39982));
  jand g21960(.dina(n39982), .dinb(n39886), .dout(n39983));
  jxor g21961(.dina(n39878), .dinb(n439), .dout(n39984));
  jnot g21962(.din(n39984), .dout(n39985));
  jor  g21963(.dina(n39985), .dinb(n39983), .dout(n39986));
  jand g21964(.dina(n39986), .dinb(n39880), .dout(n39987));
  jxor g21965(.dina(n39872), .dinb(n440), .dout(n39988));
  jnot g21966(.din(n39988), .dout(n39989));
  jor  g21967(.dina(n39989), .dinb(n39987), .dout(n39990));
  jand g21968(.dina(n39990), .dinb(n39874), .dout(n39991));
  jxor g21969(.dina(n39866), .dinb(n435), .dout(n39992));
  jnot g21970(.din(n39992), .dout(n39993));
  jor  g21971(.dina(n39993), .dinb(n39991), .dout(n39994));
  jand g21972(.dina(n39994), .dinb(n39868), .dout(n39995));
  jxor g21973(.dina(n39860), .dinb(n436), .dout(n39996));
  jnot g21974(.din(n39996), .dout(n39997));
  jor  g21975(.dina(n39997), .dinb(n39995), .dout(n39998));
  jand g21976(.dina(n39998), .dinb(n39862), .dout(n39999));
  jxor g21977(.dina(n39854), .dinb(n432), .dout(n40000));
  jnot g21978(.din(n40000), .dout(n40001));
  jor  g21979(.dina(n40001), .dinb(n39999), .dout(n40002));
  jand g21980(.dina(n40002), .dinb(n39856), .dout(n40003));
  jxor g21981(.dina(n39848), .dinb(n433), .dout(n40004));
  jnot g21982(.din(n40004), .dout(n40005));
  jor  g21983(.dina(n40005), .dinb(n40003), .dout(n40006));
  jand g21984(.dina(n40006), .dinb(n39850), .dout(n40007));
  jxor g21985(.dina(n39842), .dinb(n421), .dout(n40008));
  jnot g21986(.din(n40008), .dout(n40009));
  jor  g21987(.dina(n40009), .dinb(n40007), .dout(n40010));
  jand g21988(.dina(n40010), .dinb(n39844), .dout(n40011));
  jxor g21989(.dina(n39836), .dinb(n422), .dout(n40012));
  jnot g21990(.din(n40012), .dout(n40013));
  jor  g21991(.dina(n40013), .dinb(n40011), .dout(n40014));
  jand g21992(.dina(n40014), .dinb(n39838), .dout(n40015));
  jxor g21993(.dina(n39830), .dinb(n416), .dout(n40016));
  jnot g21994(.din(n40016), .dout(n40017));
  jor  g21995(.dina(n40017), .dinb(n40015), .dout(n40018));
  jand g21996(.dina(n40018), .dinb(n39832), .dout(n40019));
  jxor g21997(.dina(n39824), .dinb(n417), .dout(n40020));
  jnot g21998(.din(n40020), .dout(n40021));
  jor  g21999(.dina(n40021), .dinb(n40019), .dout(n40022));
  jand g22000(.dina(n40022), .dinb(n39826), .dout(n40023));
  jxor g22001(.dina(n39818), .dinb(n2547), .dout(n40024));
  jnot g22002(.din(n40024), .dout(n40025));
  jor  g22003(.dina(n40025), .dinb(n40023), .dout(n40026));
  jand g22004(.dina(n40026), .dinb(n39820), .dout(n40027));
  jxor g22005(.dina(n39812), .dinb(n2714), .dout(n40028));
  jnot g22006(.din(n40028), .dout(n40029));
  jor  g22007(.dina(n40029), .dinb(n40027), .dout(n40030));
  jand g22008(.dina(n40030), .dinb(n39814), .dout(n40031));
  jxor g22009(.dina(n39806), .dinb(n405), .dout(n40032));
  jnot g22010(.din(n40032), .dout(n40033));
  jor  g22011(.dina(n40033), .dinb(n40031), .dout(n40034));
  jand g22012(.dina(n40034), .dinb(n39808), .dout(n40035));
  jxor g22013(.dina(n39800), .dinb(n406), .dout(n40036));
  jnot g22014(.din(n40036), .dout(n40037));
  jor  g22015(.dina(n40037), .dinb(n40035), .dout(n40038));
  jand g22016(.dina(n40038), .dinb(n39802), .dout(n40039));
  jxor g22017(.dina(n39794), .dinb(n412), .dout(n40040));
  jnot g22018(.din(n40040), .dout(n40041));
  jor  g22019(.dina(n40041), .dinb(n40039), .dout(n40042));
  jand g22020(.dina(n40042), .dinb(n39796), .dout(n40043));
  jxor g22021(.dina(n39788), .dinb(n413), .dout(n40044));
  jnot g22022(.din(n40044), .dout(n40045));
  jor  g22023(.dina(n40045), .dinb(n40043), .dout(n40046));
  jand g22024(.dina(n40046), .dinb(n39790), .dout(n40047));
  jxor g22025(.dina(n39782), .dinb(n409), .dout(n40048));
  jnot g22026(.din(n40048), .dout(n40049));
  jor  g22027(.dina(n40049), .dinb(n40047), .dout(n40050));
  jand g22028(.dina(n40050), .dinb(n39784), .dout(n40051));
  jxor g22029(.dina(n39776), .dinb(n410), .dout(n40052));
  jnot g22030(.din(n40052), .dout(n40053));
  jor  g22031(.dina(n40053), .dinb(n40051), .dout(n40054));
  jand g22032(.dina(n40054), .dinb(n39778), .dout(n40055));
  jxor g22033(.dina(n39770), .dinb(n426), .dout(n40056));
  jnot g22034(.din(n40056), .dout(n40057));
  jor  g22035(.dina(n40057), .dinb(n40055), .dout(n40058));
  jand g22036(.dina(n40058), .dinb(n39772), .dout(n40059));
  jxor g22037(.dina(n39764), .dinb(n427), .dout(n40060));
  jnot g22038(.din(n40060), .dout(n40061));
  jor  g22039(.dina(n40061), .dinb(n40059), .dout(n40062));
  jand g22040(.dina(n40062), .dinb(n39766), .dout(n40063));
  jxor g22041(.dina(n39758), .dinb(n424), .dout(n40064));
  jnot g22042(.din(n40064), .dout(n40065));
  jor  g22043(.dina(n40065), .dinb(n40063), .dout(n40066));
  jand g22044(.dina(n40066), .dinb(n39760), .dout(n40067));
  jxor g22045(.dina(n39752), .dinb(n300), .dout(n40068));
  jnot g22046(.din(n40068), .dout(n40069));
  jor  g22047(.dina(n40069), .dinb(n40067), .dout(n40070));
  jand g22048(.dina(n40070), .dinb(n39754), .dout(n40071));
  jxor g22049(.dina(n39746), .dinb(n297), .dout(n40072));
  jnot g22050(.din(n40072), .dout(n40073));
  jor  g22051(.dina(n40073), .dinb(n40071), .dout(n40074));
  jand g22052(.dina(n40074), .dinb(n39748), .dout(n40075));
  jxor g22053(.dina(n39740), .dinb(n298), .dout(n40076));
  jnot g22054(.din(n40076), .dout(n40077));
  jor  g22055(.dina(n40077), .dinb(n40075), .dout(n40078));
  jand g22056(.dina(n40078), .dinb(n39742), .dout(n40079));
  jxor g22057(.dina(n39734), .dinb(n301), .dout(n40080));
  jnot g22058(.din(n40080), .dout(n40081));
  jor  g22059(.dina(n40081), .dinb(n40079), .dout(n40082));
  jand g22060(.dina(n40082), .dinb(n39736), .dout(n40083));
  jxor g22061(.dina(n39728), .dinb(n293), .dout(n40084));
  jnot g22062(.din(n40084), .dout(n40085));
  jor  g22063(.dina(n40085), .dinb(n40083), .dout(n40086));
  jand g22064(.dina(n40086), .dinb(n39730), .dout(n40087));
  jxor g22065(.dina(n39722), .dinb(n294), .dout(n40088));
  jnot g22066(.din(n40088), .dout(n40089));
  jor  g22067(.dina(n40089), .dinb(n40087), .dout(n40090));
  jand g22068(.dina(n40090), .dinb(n39724), .dout(n40091));
  jxor g22069(.dina(n39716), .dinb(n290), .dout(n40092));
  jnot g22070(.din(n40092), .dout(n40093));
  jor  g22071(.dina(n40093), .dinb(n40091), .dout(n40094));
  jand g22072(.dina(n40094), .dinb(n39718), .dout(n40095));
  jxor g22073(.dina(n39710), .dinb(n291), .dout(n40096));
  jnot g22074(.din(n40096), .dout(n40097));
  jor  g22075(.dina(n40097), .dinb(n40095), .dout(n40098));
  jand g22076(.dina(n40098), .dinb(n39712), .dout(n40099));
  jxor g22077(.dina(n39704), .dinb(n284), .dout(n40100));
  jnot g22078(.din(n40100), .dout(n40101));
  jor  g22079(.dina(n40101), .dinb(n40099), .dout(n40102));
  jand g22080(.dina(n40102), .dinb(n39706), .dout(n40103));
  jxor g22081(.dina(n39698), .dinb(n285), .dout(n40104));
  jnot g22082(.din(n40104), .dout(n40105));
  jor  g22083(.dina(n40105), .dinb(n40103), .dout(n40106));
  jand g22084(.dina(n40106), .dinb(n39700), .dout(n40107));
  jxor g22085(.dina(n39692), .dinb(n281), .dout(n40108));
  jnot g22086(.din(n40108), .dout(n40109));
  jor  g22087(.dina(n40109), .dinb(n40107), .dout(n40110));
  jand g22088(.dina(n40110), .dinb(n39694), .dout(n40111));
  jxor g22089(.dina(n39686), .dinb(n282), .dout(n40112));
  jnot g22090(.din(n40112), .dout(n40113));
  jor  g22091(.dina(n40113), .dinb(n40111), .dout(n40114));
  jand g22092(.dina(n40114), .dinb(n39688), .dout(n40115));
  jxor g22093(.dina(n39680), .dinb(n397), .dout(n40116));
  jnot g22094(.din(n40116), .dout(n40117));
  jor  g22095(.dina(n40117), .dinb(n40115), .dout(n40118));
  jand g22096(.dina(n40118), .dinb(n39682), .dout(n40119));
  jxor g22097(.dina(n39674), .dinb(n513), .dout(n40120));
  jnot g22098(.din(n40120), .dout(n40121));
  jor  g22099(.dina(n40121), .dinb(n40119), .dout(n40122));
  jand g22100(.dina(n40122), .dinb(n39676), .dout(n40123));
  jxor g22101(.dina(n39668), .dinb(n514), .dout(n40124));
  jnot g22102(.din(n40124), .dout(n40125));
  jor  g22103(.dina(n40125), .dinb(n40123), .dout(n40126));
  jand g22104(.dina(n40126), .dinb(n39670), .dout(n40127));
  jxor g22105(.dina(n39662), .dinb(n510), .dout(n40128));
  jnot g22106(.din(n40128), .dout(n40129));
  jor  g22107(.dina(n40129), .dinb(n40127), .dout(n40130));
  jand g22108(.dina(n40130), .dinb(n39664), .dout(n40131));
  jxor g22109(.dina(n39656), .dinb(n396), .dout(n40132));
  jnot g22110(.din(n40132), .dout(n40133));
  jor  g22111(.dina(n40133), .dinb(n40131), .dout(n40134));
  jand g22112(.dina(n40134), .dinb(n39658), .dout(n40135));
  jxor g22113(.dina(n39650), .dinb(n383), .dout(n40136));
  jnot g22114(.din(n40136), .dout(n40137));
  jor  g22115(.dina(n40137), .dinb(n40135), .dout(n40138));
  jand g22116(.dina(n40138), .dinb(n39652), .dout(n40139));
  jxor g22117(.dina(n39644), .dinb(n12211), .dout(n40140));
  jnot g22118(.din(n40140), .dout(n40141));
  jor  g22119(.dina(n40141), .dinb(n40139), .dout(n40142));
  jand g22120(.dina(n40142), .dinb(n39646), .dout(n40143));
  jxor g22121(.dina(n39638), .dinb(n12214), .dout(n40144));
  jnot g22122(.din(n40144), .dout(n40145));
  jor  g22123(.dina(n40145), .dinb(n40143), .dout(n40146));
  jand g22124(.dina(n40146), .dinb(n39640), .dout(n40147));
  jxor g22125(.dina(n39632), .dinb(n384), .dout(n40148));
  jnot g22126(.din(n40148), .dout(n40149));
  jor  g22127(.dina(n40149), .dinb(n40147), .dout(n40150));
  jand g22128(.dina(n40150), .dinb(n39634), .dout(n40151));
  jxor g22129(.dina(n39626), .dinb(n374), .dout(n40152));
  jnot g22130(.din(n40152), .dout(n40153));
  jor  g22131(.dina(n40153), .dinb(n40151), .dout(n40154));
  jand g22132(.dina(n40154), .dinb(n39628), .dout(n40155));
  jxor g22133(.dina(n39620), .dinb(n376), .dout(n40156));
  jnot g22134(.din(n40156), .dout(n40157));
  jor  g22135(.dina(n40157), .dinb(n40155), .dout(n40158));
  jand g22136(.dina(n40158), .dinb(n39622), .dout(n40159));
  jxor g22137(.dina(n39614), .dinb(n377), .dout(n40160));
  jnot g22138(.din(n40160), .dout(n40161));
  jor  g22139(.dina(n40161), .dinb(n40159), .dout(n40162));
  jand g22140(.dina(n40162), .dinb(n39616), .dout(n40163));
  jxor g22141(.dina(n39608), .dinb(n375), .dout(n40164));
  jnot g22142(.din(n40164), .dout(n40165));
  jor  g22143(.dina(n40165), .dinb(n40163), .dout(n40166));
  jand g22144(.dina(n40166), .dinb(n39610), .dout(n40167));
  jxor g22145(.dina(n39602), .dinb(n362), .dout(n40168));
  jnot g22146(.din(n40168), .dout(n40169));
  jor  g22147(.dina(n40169), .dinb(n40167), .dout(n40170));
  jand g22148(.dina(n40170), .dinb(n39604), .dout(n40171));
  jxor g22149(.dina(n39596), .dinb(n363), .dout(n40172));
  jnot g22150(.din(n40172), .dout(n40173));
  jor  g22151(.dina(n40173), .dinb(n40171), .dout(n40174));
  jand g22152(.dina(n40174), .dinb(n39598), .dout(n40175));
  jand g22153(.dina(n39589), .dinb(n365), .dout(n40176));
  jnot g22154(.din(n40176), .dout(n40177));
  jand g22155(.dina(n40177), .dinb(n40175), .dout(n40178));
  jnot g22156(.din(n39589), .dout(n40179));
  jand g22157(.dina(n40179), .dinb(b59 ), .dout(n40180));
  jor  g22158(.dina(n40180), .dinb(n264), .dout(n40181));
  jor  g22159(.dina(n40181), .dinb(n40178), .dout(n40182));
  jxor g22160(.dina(n39944), .dinb(b1 ), .dout(n40183));
  jand g22161(.dina(n40183), .dinb(n16327), .dout(n40184));
  jor  g22162(.dina(n40184), .dinb(n39940), .dout(n40185));
  jand g22163(.dina(n39948), .dinb(n40185), .dout(n40186));
  jor  g22164(.dina(n40186), .dinb(n39933), .dout(n40187));
  jand g22165(.dina(n39952), .dinb(n40187), .dout(n40188));
  jor  g22166(.dina(n40188), .dinb(n39927), .dout(n40189));
  jand g22167(.dina(n39956), .dinb(n40189), .dout(n40190));
  jor  g22168(.dina(n40190), .dinb(n39921), .dout(n40191));
  jand g22169(.dina(n39960), .dinb(n40191), .dout(n40192));
  jor  g22170(.dina(n40192), .dinb(n39915), .dout(n40193));
  jand g22171(.dina(n39964), .dinb(n40193), .dout(n40194));
  jor  g22172(.dina(n40194), .dinb(n39909), .dout(n40195));
  jand g22173(.dina(n39968), .dinb(n40195), .dout(n40196));
  jor  g22174(.dina(n40196), .dinb(n39903), .dout(n40197));
  jand g22175(.dina(n39972), .dinb(n40197), .dout(n40198));
  jor  g22176(.dina(n40198), .dinb(n39897), .dout(n40199));
  jand g22177(.dina(n39976), .dinb(n40199), .dout(n40200));
  jor  g22178(.dina(n40200), .dinb(n39891), .dout(n40201));
  jand g22179(.dina(n39980), .dinb(n40201), .dout(n40202));
  jor  g22180(.dina(n40202), .dinb(n39885), .dout(n40203));
  jand g22181(.dina(n39984), .dinb(n40203), .dout(n40204));
  jor  g22182(.dina(n40204), .dinb(n39879), .dout(n40205));
  jand g22183(.dina(n39988), .dinb(n40205), .dout(n40206));
  jor  g22184(.dina(n40206), .dinb(n39873), .dout(n40207));
  jand g22185(.dina(n39992), .dinb(n40207), .dout(n40208));
  jor  g22186(.dina(n40208), .dinb(n39867), .dout(n40209));
  jand g22187(.dina(n39996), .dinb(n40209), .dout(n40210));
  jor  g22188(.dina(n40210), .dinb(n39861), .dout(n40211));
  jand g22189(.dina(n40000), .dinb(n40211), .dout(n40212));
  jor  g22190(.dina(n40212), .dinb(n39855), .dout(n40213));
  jand g22191(.dina(n40004), .dinb(n40213), .dout(n40214));
  jor  g22192(.dina(n40214), .dinb(n39849), .dout(n40215));
  jand g22193(.dina(n40008), .dinb(n40215), .dout(n40216));
  jor  g22194(.dina(n40216), .dinb(n39843), .dout(n40217));
  jand g22195(.dina(n40012), .dinb(n40217), .dout(n40218));
  jor  g22196(.dina(n40218), .dinb(n39837), .dout(n40219));
  jand g22197(.dina(n40016), .dinb(n40219), .dout(n40220));
  jor  g22198(.dina(n40220), .dinb(n39831), .dout(n40221));
  jand g22199(.dina(n40020), .dinb(n40221), .dout(n40222));
  jor  g22200(.dina(n40222), .dinb(n39825), .dout(n40223));
  jand g22201(.dina(n40024), .dinb(n40223), .dout(n40224));
  jor  g22202(.dina(n40224), .dinb(n39819), .dout(n40225));
  jand g22203(.dina(n40028), .dinb(n40225), .dout(n40226));
  jor  g22204(.dina(n40226), .dinb(n39813), .dout(n40227));
  jand g22205(.dina(n40032), .dinb(n40227), .dout(n40228));
  jor  g22206(.dina(n40228), .dinb(n39807), .dout(n40229));
  jand g22207(.dina(n40036), .dinb(n40229), .dout(n40230));
  jor  g22208(.dina(n40230), .dinb(n39801), .dout(n40231));
  jand g22209(.dina(n40040), .dinb(n40231), .dout(n40232));
  jor  g22210(.dina(n40232), .dinb(n39795), .dout(n40233));
  jand g22211(.dina(n40044), .dinb(n40233), .dout(n40234));
  jor  g22212(.dina(n40234), .dinb(n39789), .dout(n40235));
  jand g22213(.dina(n40048), .dinb(n40235), .dout(n40236));
  jor  g22214(.dina(n40236), .dinb(n39783), .dout(n40237));
  jand g22215(.dina(n40052), .dinb(n40237), .dout(n40238));
  jor  g22216(.dina(n40238), .dinb(n39777), .dout(n40239));
  jand g22217(.dina(n40056), .dinb(n40239), .dout(n40240));
  jor  g22218(.dina(n40240), .dinb(n39771), .dout(n40241));
  jand g22219(.dina(n40060), .dinb(n40241), .dout(n40242));
  jor  g22220(.dina(n40242), .dinb(n39765), .dout(n40243));
  jand g22221(.dina(n40064), .dinb(n40243), .dout(n40244));
  jor  g22222(.dina(n40244), .dinb(n39759), .dout(n40245));
  jand g22223(.dina(n40068), .dinb(n40245), .dout(n40246));
  jor  g22224(.dina(n40246), .dinb(n39753), .dout(n40247));
  jand g22225(.dina(n40072), .dinb(n40247), .dout(n40248));
  jor  g22226(.dina(n40248), .dinb(n39747), .dout(n40249));
  jand g22227(.dina(n40076), .dinb(n40249), .dout(n40250));
  jor  g22228(.dina(n40250), .dinb(n39741), .dout(n40251));
  jand g22229(.dina(n40080), .dinb(n40251), .dout(n40252));
  jor  g22230(.dina(n40252), .dinb(n39735), .dout(n40253));
  jand g22231(.dina(n40084), .dinb(n40253), .dout(n40254));
  jor  g22232(.dina(n40254), .dinb(n39729), .dout(n40255));
  jand g22233(.dina(n40088), .dinb(n40255), .dout(n40256));
  jor  g22234(.dina(n40256), .dinb(n39723), .dout(n40257));
  jand g22235(.dina(n40092), .dinb(n40257), .dout(n40258));
  jor  g22236(.dina(n40258), .dinb(n39717), .dout(n40259));
  jand g22237(.dina(n40096), .dinb(n40259), .dout(n40260));
  jor  g22238(.dina(n40260), .dinb(n39711), .dout(n40261));
  jand g22239(.dina(n40100), .dinb(n40261), .dout(n40262));
  jor  g22240(.dina(n40262), .dinb(n39705), .dout(n40263));
  jand g22241(.dina(n40104), .dinb(n40263), .dout(n40264));
  jor  g22242(.dina(n40264), .dinb(n39699), .dout(n40265));
  jand g22243(.dina(n40108), .dinb(n40265), .dout(n40266));
  jor  g22244(.dina(n40266), .dinb(n39693), .dout(n40267));
  jand g22245(.dina(n40112), .dinb(n40267), .dout(n40268));
  jor  g22246(.dina(n40268), .dinb(n39687), .dout(n40269));
  jand g22247(.dina(n40116), .dinb(n40269), .dout(n40270));
  jor  g22248(.dina(n40270), .dinb(n39681), .dout(n40271));
  jand g22249(.dina(n40120), .dinb(n40271), .dout(n40272));
  jor  g22250(.dina(n40272), .dinb(n39675), .dout(n40273));
  jand g22251(.dina(n40124), .dinb(n40273), .dout(n40274));
  jor  g22252(.dina(n40274), .dinb(n39669), .dout(n40275));
  jand g22253(.dina(n40128), .dinb(n40275), .dout(n40276));
  jor  g22254(.dina(n40276), .dinb(n39663), .dout(n40277));
  jand g22255(.dina(n40132), .dinb(n40277), .dout(n40278));
  jor  g22256(.dina(n40278), .dinb(n39657), .dout(n40279));
  jand g22257(.dina(n40136), .dinb(n40279), .dout(n40280));
  jor  g22258(.dina(n40280), .dinb(n39651), .dout(n40281));
  jand g22259(.dina(n40140), .dinb(n40281), .dout(n40282));
  jor  g22260(.dina(n40282), .dinb(n39645), .dout(n40283));
  jand g22261(.dina(n40144), .dinb(n40283), .dout(n40284));
  jor  g22262(.dina(n40284), .dinb(n39639), .dout(n40285));
  jand g22263(.dina(n40148), .dinb(n40285), .dout(n40286));
  jor  g22264(.dina(n40286), .dinb(n39633), .dout(n40287));
  jand g22265(.dina(n40152), .dinb(n40287), .dout(n40288));
  jor  g22266(.dina(n40288), .dinb(n39627), .dout(n40289));
  jand g22267(.dina(n40156), .dinb(n40289), .dout(n40290));
  jor  g22268(.dina(n40290), .dinb(n39621), .dout(n40291));
  jand g22269(.dina(n40160), .dinb(n40291), .dout(n40292));
  jor  g22270(.dina(n40292), .dinb(n39615), .dout(n40293));
  jand g22271(.dina(n40164), .dinb(n40293), .dout(n40294));
  jor  g22272(.dina(n40294), .dinb(n39609), .dout(n40295));
  jand g22273(.dina(n40168), .dinb(n40295), .dout(n40296));
  jor  g22274(.dina(n40296), .dinb(n39603), .dout(n40297));
  jand g22275(.dina(n40172), .dinb(n40297), .dout(n40298));
  jor  g22276(.dina(n40298), .dinb(n39597), .dout(n40299));
  jand g22277(.dina(n40299), .dinb(n372), .dout(n40300));
  jor  g22278(.dina(n40300), .dinb(n40182), .dout(n40301));
  jand g22279(.dina(n40301), .dinb(n39589), .dout(n40302));
  jand g22280(.dina(n40182), .dinb(n39596), .dout(n40303));
  jor  g22281(.dina(n40176), .dinb(n40299), .dout(n40304));
  jnot g22282(.din(n40181), .dout(n40305));
  jand g22283(.dina(n40305), .dinb(n40304), .dout(n40306));
  jxor g22284(.dina(n40172), .dinb(n40297), .dout(n40307));
  jand g22285(.dina(n40307), .dinb(n40306), .dout(n40308));
  jor  g22286(.dina(n40308), .dinb(n40303), .dout(n40309));
  jand g22287(.dina(n40309), .dinb(n365), .dout(n40310));
  jnot g22288(.din(n40310), .dout(n40311));
  jand g22289(.dina(n40182), .dinb(n39602), .dout(n40312));
  jxor g22290(.dina(n40168), .dinb(n40295), .dout(n40313));
  jand g22291(.dina(n40313), .dinb(n40306), .dout(n40314));
  jor  g22292(.dina(n40314), .dinb(n40312), .dout(n40315));
  jand g22293(.dina(n40315), .dinb(n363), .dout(n40316));
  jnot g22294(.din(n40316), .dout(n40317));
  jand g22295(.dina(n40182), .dinb(n39608), .dout(n40318));
  jxor g22296(.dina(n40164), .dinb(n40293), .dout(n40319));
  jand g22297(.dina(n40319), .dinb(n40306), .dout(n40320));
  jor  g22298(.dina(n40320), .dinb(n40318), .dout(n40321));
  jand g22299(.dina(n40321), .dinb(n362), .dout(n40322));
  jnot g22300(.din(n40322), .dout(n40323));
  jand g22301(.dina(n40182), .dinb(n39614), .dout(n40324));
  jxor g22302(.dina(n40160), .dinb(n40291), .dout(n40325));
  jand g22303(.dina(n40325), .dinb(n40306), .dout(n40326));
  jor  g22304(.dina(n40326), .dinb(n40324), .dout(n40327));
  jand g22305(.dina(n40327), .dinb(n375), .dout(n40328));
  jnot g22306(.din(n40328), .dout(n40329));
  jand g22307(.dina(n40182), .dinb(n39620), .dout(n40330));
  jxor g22308(.dina(n40156), .dinb(n40289), .dout(n40331));
  jand g22309(.dina(n40331), .dinb(n40306), .dout(n40332));
  jor  g22310(.dina(n40332), .dinb(n40330), .dout(n40333));
  jand g22311(.dina(n40333), .dinb(n377), .dout(n40334));
  jnot g22312(.din(n40334), .dout(n40335));
  jand g22313(.dina(n40182), .dinb(n39626), .dout(n40336));
  jxor g22314(.dina(n40152), .dinb(n40287), .dout(n40337));
  jand g22315(.dina(n40337), .dinb(n40306), .dout(n40338));
  jor  g22316(.dina(n40338), .dinb(n40336), .dout(n40339));
  jand g22317(.dina(n40339), .dinb(n376), .dout(n40340));
  jnot g22318(.din(n40340), .dout(n40341));
  jand g22319(.dina(n40182), .dinb(n39632), .dout(n40342));
  jxor g22320(.dina(n40148), .dinb(n40285), .dout(n40343));
  jand g22321(.dina(n40343), .dinb(n40306), .dout(n40344));
  jor  g22322(.dina(n40344), .dinb(n40342), .dout(n40345));
  jand g22323(.dina(n40345), .dinb(n374), .dout(n40346));
  jnot g22324(.din(n40346), .dout(n40347));
  jand g22325(.dina(n40182), .dinb(n39638), .dout(n40348));
  jxor g22326(.dina(n40144), .dinb(n40283), .dout(n40349));
  jand g22327(.dina(n40349), .dinb(n40306), .dout(n40350));
  jor  g22328(.dina(n40350), .dinb(n40348), .dout(n40351));
  jand g22329(.dina(n40351), .dinb(n384), .dout(n40352));
  jnot g22330(.din(n40352), .dout(n40353));
  jand g22331(.dina(n40182), .dinb(n39644), .dout(n40354));
  jxor g22332(.dina(n40140), .dinb(n40281), .dout(n40355));
  jand g22333(.dina(n40355), .dinb(n40306), .dout(n40356));
  jor  g22334(.dina(n40356), .dinb(n40354), .dout(n40357));
  jand g22335(.dina(n40357), .dinb(n12214), .dout(n40358));
  jnot g22336(.din(n40358), .dout(n40359));
  jand g22337(.dina(n40182), .dinb(n39650), .dout(n40360));
  jxor g22338(.dina(n40136), .dinb(n40279), .dout(n40361));
  jand g22339(.dina(n40361), .dinb(n40306), .dout(n40362));
  jor  g22340(.dina(n40362), .dinb(n40360), .dout(n40363));
  jand g22341(.dina(n40363), .dinb(n12211), .dout(n40364));
  jnot g22342(.din(n40364), .dout(n40365));
  jand g22343(.dina(n40182), .dinb(n39656), .dout(n40366));
  jxor g22344(.dina(n40132), .dinb(n40277), .dout(n40367));
  jand g22345(.dina(n40367), .dinb(n40306), .dout(n40368));
  jor  g22346(.dina(n40368), .dinb(n40366), .dout(n40369));
  jand g22347(.dina(n40369), .dinb(n383), .dout(n40370));
  jnot g22348(.din(n40370), .dout(n40371));
  jand g22349(.dina(n40182), .dinb(n39662), .dout(n40372));
  jxor g22350(.dina(n40128), .dinb(n40275), .dout(n40373));
  jand g22351(.dina(n40373), .dinb(n40306), .dout(n40374));
  jor  g22352(.dina(n40374), .dinb(n40372), .dout(n40375));
  jand g22353(.dina(n40375), .dinb(n396), .dout(n40376));
  jnot g22354(.din(n40376), .dout(n40377));
  jand g22355(.dina(n40182), .dinb(n39668), .dout(n40378));
  jxor g22356(.dina(n40124), .dinb(n40273), .dout(n40379));
  jand g22357(.dina(n40379), .dinb(n40306), .dout(n40380));
  jor  g22358(.dina(n40380), .dinb(n40378), .dout(n40381));
  jand g22359(.dina(n40381), .dinb(n510), .dout(n40382));
  jnot g22360(.din(n40382), .dout(n40383));
  jand g22361(.dina(n40182), .dinb(n39674), .dout(n40384));
  jxor g22362(.dina(n40120), .dinb(n40271), .dout(n40385));
  jand g22363(.dina(n40385), .dinb(n40306), .dout(n40386));
  jor  g22364(.dina(n40386), .dinb(n40384), .dout(n40387));
  jand g22365(.dina(n40387), .dinb(n514), .dout(n40388));
  jnot g22366(.din(n40388), .dout(n40389));
  jand g22367(.dina(n40182), .dinb(n39680), .dout(n40390));
  jxor g22368(.dina(n40116), .dinb(n40269), .dout(n40391));
  jand g22369(.dina(n40391), .dinb(n40306), .dout(n40392));
  jor  g22370(.dina(n40392), .dinb(n40390), .dout(n40393));
  jand g22371(.dina(n40393), .dinb(n513), .dout(n40394));
  jnot g22372(.din(n40394), .dout(n40395));
  jand g22373(.dina(n40182), .dinb(n39686), .dout(n40396));
  jxor g22374(.dina(n40112), .dinb(n40267), .dout(n40397));
  jand g22375(.dina(n40397), .dinb(n40306), .dout(n40398));
  jor  g22376(.dina(n40398), .dinb(n40396), .dout(n40399));
  jand g22377(.dina(n40399), .dinb(n397), .dout(n40400));
  jnot g22378(.din(n40400), .dout(n40401));
  jand g22379(.dina(n40182), .dinb(n39692), .dout(n40402));
  jxor g22380(.dina(n40108), .dinb(n40265), .dout(n40403));
  jand g22381(.dina(n40403), .dinb(n40306), .dout(n40404));
  jor  g22382(.dina(n40404), .dinb(n40402), .dout(n40405));
  jand g22383(.dina(n40405), .dinb(n282), .dout(n40406));
  jnot g22384(.din(n40406), .dout(n40407));
  jand g22385(.dina(n40182), .dinb(n39698), .dout(n40408));
  jxor g22386(.dina(n40104), .dinb(n40263), .dout(n40409));
  jand g22387(.dina(n40409), .dinb(n40306), .dout(n40410));
  jor  g22388(.dina(n40410), .dinb(n40408), .dout(n40411));
  jand g22389(.dina(n40411), .dinb(n281), .dout(n40412));
  jnot g22390(.din(n40412), .dout(n40413));
  jand g22391(.dina(n40182), .dinb(n39704), .dout(n40414));
  jxor g22392(.dina(n40100), .dinb(n40261), .dout(n40415));
  jand g22393(.dina(n40415), .dinb(n40306), .dout(n40416));
  jor  g22394(.dina(n40416), .dinb(n40414), .dout(n40417));
  jand g22395(.dina(n40417), .dinb(n285), .dout(n40418));
  jnot g22396(.din(n40418), .dout(n40419));
  jand g22397(.dina(n40182), .dinb(n39710), .dout(n40420));
  jxor g22398(.dina(n40096), .dinb(n40259), .dout(n40421));
  jand g22399(.dina(n40421), .dinb(n40306), .dout(n40422));
  jor  g22400(.dina(n40422), .dinb(n40420), .dout(n40423));
  jand g22401(.dina(n40423), .dinb(n284), .dout(n40424));
  jnot g22402(.din(n40424), .dout(n40425));
  jand g22403(.dina(n40182), .dinb(n39716), .dout(n40426));
  jxor g22404(.dina(n40092), .dinb(n40257), .dout(n40427));
  jand g22405(.dina(n40427), .dinb(n40306), .dout(n40428));
  jor  g22406(.dina(n40428), .dinb(n40426), .dout(n40429));
  jand g22407(.dina(n40429), .dinb(n291), .dout(n40430));
  jnot g22408(.din(n40430), .dout(n40431));
  jand g22409(.dina(n40182), .dinb(n39722), .dout(n40432));
  jxor g22410(.dina(n40088), .dinb(n40255), .dout(n40433));
  jand g22411(.dina(n40433), .dinb(n40306), .dout(n40434));
  jor  g22412(.dina(n40434), .dinb(n40432), .dout(n40435));
  jand g22413(.dina(n40435), .dinb(n290), .dout(n40436));
  jnot g22414(.din(n40436), .dout(n40437));
  jand g22415(.dina(n40182), .dinb(n39728), .dout(n40438));
  jxor g22416(.dina(n40084), .dinb(n40253), .dout(n40439));
  jand g22417(.dina(n40439), .dinb(n40306), .dout(n40440));
  jor  g22418(.dina(n40440), .dinb(n40438), .dout(n40441));
  jand g22419(.dina(n40441), .dinb(n294), .dout(n40442));
  jnot g22420(.din(n40442), .dout(n40443));
  jand g22421(.dina(n40182), .dinb(n39734), .dout(n40444));
  jxor g22422(.dina(n40080), .dinb(n40251), .dout(n40445));
  jand g22423(.dina(n40445), .dinb(n40306), .dout(n40446));
  jor  g22424(.dina(n40446), .dinb(n40444), .dout(n40447));
  jand g22425(.dina(n40447), .dinb(n293), .dout(n40448));
  jnot g22426(.din(n40448), .dout(n40449));
  jand g22427(.dina(n40182), .dinb(n39740), .dout(n40450));
  jxor g22428(.dina(n40076), .dinb(n40249), .dout(n40451));
  jand g22429(.dina(n40451), .dinb(n40306), .dout(n40452));
  jor  g22430(.dina(n40452), .dinb(n40450), .dout(n40453));
  jand g22431(.dina(n40453), .dinb(n301), .dout(n40454));
  jnot g22432(.din(n40454), .dout(n40455));
  jand g22433(.dina(n40182), .dinb(n39746), .dout(n40456));
  jxor g22434(.dina(n40072), .dinb(n40247), .dout(n40457));
  jand g22435(.dina(n40457), .dinb(n40306), .dout(n40458));
  jor  g22436(.dina(n40458), .dinb(n40456), .dout(n40459));
  jand g22437(.dina(n40459), .dinb(n298), .dout(n40460));
  jnot g22438(.din(n40460), .dout(n40461));
  jand g22439(.dina(n40182), .dinb(n39752), .dout(n40462));
  jxor g22440(.dina(n40068), .dinb(n40245), .dout(n40463));
  jand g22441(.dina(n40463), .dinb(n40306), .dout(n40464));
  jor  g22442(.dina(n40464), .dinb(n40462), .dout(n40465));
  jand g22443(.dina(n40465), .dinb(n297), .dout(n40466));
  jnot g22444(.din(n40466), .dout(n40467));
  jand g22445(.dina(n40182), .dinb(n39758), .dout(n40468));
  jxor g22446(.dina(n40064), .dinb(n40243), .dout(n40469));
  jand g22447(.dina(n40469), .dinb(n40306), .dout(n40470));
  jor  g22448(.dina(n40470), .dinb(n40468), .dout(n40471));
  jand g22449(.dina(n40471), .dinb(n300), .dout(n40472));
  jnot g22450(.din(n40472), .dout(n40473));
  jand g22451(.dina(n40182), .dinb(n39764), .dout(n40474));
  jxor g22452(.dina(n40060), .dinb(n40241), .dout(n40475));
  jand g22453(.dina(n40475), .dinb(n40306), .dout(n40476));
  jor  g22454(.dina(n40476), .dinb(n40474), .dout(n40477));
  jand g22455(.dina(n40477), .dinb(n424), .dout(n40478));
  jnot g22456(.din(n40478), .dout(n40479));
  jand g22457(.dina(n40182), .dinb(n39770), .dout(n40480));
  jxor g22458(.dina(n40056), .dinb(n40239), .dout(n40481));
  jand g22459(.dina(n40481), .dinb(n40306), .dout(n40482));
  jor  g22460(.dina(n40482), .dinb(n40480), .dout(n40483));
  jand g22461(.dina(n40483), .dinb(n427), .dout(n40484));
  jnot g22462(.din(n40484), .dout(n40485));
  jand g22463(.dina(n40182), .dinb(n39776), .dout(n40486));
  jxor g22464(.dina(n40052), .dinb(n40237), .dout(n40487));
  jand g22465(.dina(n40487), .dinb(n40306), .dout(n40488));
  jor  g22466(.dina(n40488), .dinb(n40486), .dout(n40489));
  jand g22467(.dina(n40489), .dinb(n426), .dout(n40490));
  jnot g22468(.din(n40490), .dout(n40491));
  jand g22469(.dina(n40182), .dinb(n39782), .dout(n40492));
  jxor g22470(.dina(n40048), .dinb(n40235), .dout(n40493));
  jand g22471(.dina(n40493), .dinb(n40306), .dout(n40494));
  jor  g22472(.dina(n40494), .dinb(n40492), .dout(n40495));
  jand g22473(.dina(n40495), .dinb(n410), .dout(n40496));
  jnot g22474(.din(n40496), .dout(n40497));
  jand g22475(.dina(n40182), .dinb(n39788), .dout(n40498));
  jxor g22476(.dina(n40044), .dinb(n40233), .dout(n40499));
  jand g22477(.dina(n40499), .dinb(n40306), .dout(n40500));
  jor  g22478(.dina(n40500), .dinb(n40498), .dout(n40501));
  jand g22479(.dina(n40501), .dinb(n409), .dout(n40502));
  jnot g22480(.din(n40502), .dout(n40503));
  jand g22481(.dina(n40182), .dinb(n39794), .dout(n40504));
  jxor g22482(.dina(n40040), .dinb(n40231), .dout(n40505));
  jand g22483(.dina(n40505), .dinb(n40306), .dout(n40506));
  jor  g22484(.dina(n40506), .dinb(n40504), .dout(n40507));
  jand g22485(.dina(n40507), .dinb(n413), .dout(n40508));
  jnot g22486(.din(n40508), .dout(n40509));
  jand g22487(.dina(n40182), .dinb(n39800), .dout(n40510));
  jxor g22488(.dina(n40036), .dinb(n40229), .dout(n40511));
  jand g22489(.dina(n40511), .dinb(n40306), .dout(n40512));
  jor  g22490(.dina(n40512), .dinb(n40510), .dout(n40513));
  jand g22491(.dina(n40513), .dinb(n412), .dout(n40514));
  jnot g22492(.din(n40514), .dout(n40515));
  jand g22493(.dina(n40182), .dinb(n39806), .dout(n40516));
  jxor g22494(.dina(n40032), .dinb(n40227), .dout(n40517));
  jand g22495(.dina(n40517), .dinb(n40306), .dout(n40518));
  jor  g22496(.dina(n40518), .dinb(n40516), .dout(n40519));
  jand g22497(.dina(n40519), .dinb(n406), .dout(n40520));
  jnot g22498(.din(n40520), .dout(n40521));
  jand g22499(.dina(n40182), .dinb(n39812), .dout(n40522));
  jxor g22500(.dina(n40028), .dinb(n40225), .dout(n40523));
  jand g22501(.dina(n40523), .dinb(n40306), .dout(n40524));
  jor  g22502(.dina(n40524), .dinb(n40522), .dout(n40525));
  jand g22503(.dina(n40525), .dinb(n405), .dout(n40526));
  jnot g22504(.din(n40526), .dout(n40527));
  jand g22505(.dina(n40182), .dinb(n39818), .dout(n40528));
  jxor g22506(.dina(n40024), .dinb(n40223), .dout(n40529));
  jand g22507(.dina(n40529), .dinb(n40306), .dout(n40530));
  jor  g22508(.dina(n40530), .dinb(n40528), .dout(n40531));
  jand g22509(.dina(n40531), .dinb(n2714), .dout(n40532));
  jnot g22510(.din(n40532), .dout(n40533));
  jand g22511(.dina(n40182), .dinb(n39824), .dout(n40534));
  jxor g22512(.dina(n40020), .dinb(n40221), .dout(n40535));
  jand g22513(.dina(n40535), .dinb(n40306), .dout(n40536));
  jor  g22514(.dina(n40536), .dinb(n40534), .dout(n40537));
  jand g22515(.dina(n40537), .dinb(n2547), .dout(n40538));
  jnot g22516(.din(n40538), .dout(n40539));
  jand g22517(.dina(n40182), .dinb(n39830), .dout(n40540));
  jxor g22518(.dina(n40016), .dinb(n40219), .dout(n40541));
  jand g22519(.dina(n40541), .dinb(n40306), .dout(n40542));
  jor  g22520(.dina(n40542), .dinb(n40540), .dout(n40543));
  jand g22521(.dina(n40543), .dinb(n417), .dout(n40544));
  jnot g22522(.din(n40544), .dout(n40545));
  jand g22523(.dina(n40182), .dinb(n39836), .dout(n40546));
  jxor g22524(.dina(n40012), .dinb(n40217), .dout(n40547));
  jand g22525(.dina(n40547), .dinb(n40306), .dout(n40548));
  jor  g22526(.dina(n40548), .dinb(n40546), .dout(n40549));
  jand g22527(.dina(n40549), .dinb(n416), .dout(n40550));
  jnot g22528(.din(n40550), .dout(n40551));
  jand g22529(.dina(n40182), .dinb(n39842), .dout(n40552));
  jxor g22530(.dina(n40008), .dinb(n40215), .dout(n40553));
  jand g22531(.dina(n40553), .dinb(n40306), .dout(n40554));
  jor  g22532(.dina(n40554), .dinb(n40552), .dout(n40555));
  jand g22533(.dina(n40555), .dinb(n422), .dout(n40556));
  jnot g22534(.din(n40556), .dout(n40557));
  jand g22535(.dina(n40182), .dinb(n39848), .dout(n40558));
  jxor g22536(.dina(n40004), .dinb(n40213), .dout(n40559));
  jand g22537(.dina(n40559), .dinb(n40306), .dout(n40560));
  jor  g22538(.dina(n40560), .dinb(n40558), .dout(n40561));
  jand g22539(.dina(n40561), .dinb(n421), .dout(n40562));
  jnot g22540(.din(n40562), .dout(n40563));
  jand g22541(.dina(n40182), .dinb(n39854), .dout(n40564));
  jxor g22542(.dina(n40000), .dinb(n40211), .dout(n40565));
  jand g22543(.dina(n40565), .dinb(n40306), .dout(n40566));
  jor  g22544(.dina(n40566), .dinb(n40564), .dout(n40567));
  jand g22545(.dina(n40567), .dinb(n433), .dout(n40568));
  jnot g22546(.din(n40568), .dout(n40569));
  jand g22547(.dina(n40182), .dinb(n39860), .dout(n40570));
  jxor g22548(.dina(n39996), .dinb(n40209), .dout(n40571));
  jand g22549(.dina(n40571), .dinb(n40306), .dout(n40572));
  jor  g22550(.dina(n40572), .dinb(n40570), .dout(n40573));
  jand g22551(.dina(n40573), .dinb(n432), .dout(n40574));
  jnot g22552(.din(n40574), .dout(n40575));
  jand g22553(.dina(n40182), .dinb(n39866), .dout(n40576));
  jxor g22554(.dina(n39992), .dinb(n40207), .dout(n40577));
  jand g22555(.dina(n40577), .dinb(n40306), .dout(n40578));
  jor  g22556(.dina(n40578), .dinb(n40576), .dout(n40579));
  jand g22557(.dina(n40579), .dinb(n436), .dout(n40580));
  jnot g22558(.din(n40580), .dout(n40581));
  jand g22559(.dina(n40182), .dinb(n39872), .dout(n40582));
  jxor g22560(.dina(n39988), .dinb(n40205), .dout(n40583));
  jand g22561(.dina(n40583), .dinb(n40306), .dout(n40584));
  jor  g22562(.dina(n40584), .dinb(n40582), .dout(n40585));
  jand g22563(.dina(n40585), .dinb(n435), .dout(n40586));
  jnot g22564(.din(n40586), .dout(n40587));
  jand g22565(.dina(n40182), .dinb(n39878), .dout(n40588));
  jxor g22566(.dina(n39984), .dinb(n40203), .dout(n40589));
  jand g22567(.dina(n40589), .dinb(n40306), .dout(n40590));
  jor  g22568(.dina(n40590), .dinb(n40588), .dout(n40591));
  jand g22569(.dina(n40591), .dinb(n440), .dout(n40592));
  jnot g22570(.din(n40592), .dout(n40593));
  jand g22571(.dina(n40182), .dinb(n39884), .dout(n40594));
  jxor g22572(.dina(n39980), .dinb(n40201), .dout(n40595));
  jand g22573(.dina(n40595), .dinb(n40306), .dout(n40596));
  jor  g22574(.dina(n40596), .dinb(n40594), .dout(n40597));
  jand g22575(.dina(n40597), .dinb(n439), .dout(n40598));
  jnot g22576(.din(n40598), .dout(n40599));
  jand g22577(.dina(n40182), .dinb(n39890), .dout(n40600));
  jxor g22578(.dina(n39976), .dinb(n40199), .dout(n40601));
  jand g22579(.dina(n40601), .dinb(n40306), .dout(n40602));
  jor  g22580(.dina(n40602), .dinb(n40600), .dout(n40603));
  jand g22581(.dina(n40603), .dinb(n325), .dout(n40604));
  jnot g22582(.din(n40604), .dout(n40605));
  jand g22583(.dina(n40182), .dinb(n39896), .dout(n40606));
  jxor g22584(.dina(n39972), .dinb(n40197), .dout(n40607));
  jand g22585(.dina(n40607), .dinb(n40306), .dout(n40608));
  jor  g22586(.dina(n40608), .dinb(n40606), .dout(n40609));
  jand g22587(.dina(n40609), .dinb(n324), .dout(n40610));
  jnot g22588(.din(n40610), .dout(n40611));
  jand g22589(.dina(n40182), .dinb(n39902), .dout(n40612));
  jxor g22590(.dina(n39968), .dinb(n40195), .dout(n40613));
  jand g22591(.dina(n40613), .dinb(n40306), .dout(n40614));
  jor  g22592(.dina(n40614), .dinb(n40612), .dout(n40615));
  jand g22593(.dina(n40615), .dinb(n323), .dout(n40616));
  jnot g22594(.din(n40616), .dout(n40617));
  jand g22595(.dina(n40182), .dinb(n39908), .dout(n40618));
  jxor g22596(.dina(n39964), .dinb(n40193), .dout(n40619));
  jand g22597(.dina(n40619), .dinb(n40306), .dout(n40620));
  jor  g22598(.dina(n40620), .dinb(n40618), .dout(n40621));
  jand g22599(.dina(n40621), .dinb(n335), .dout(n40622));
  jnot g22600(.din(n40622), .dout(n40623));
  jand g22601(.dina(n40182), .dinb(n39914), .dout(n40624));
  jxor g22602(.dina(n39960), .dinb(n40191), .dout(n40625));
  jand g22603(.dina(n40625), .dinb(n40306), .dout(n40626));
  jor  g22604(.dina(n40626), .dinb(n40624), .dout(n40627));
  jand g22605(.dina(n40627), .dinb(n334), .dout(n40628));
  jnot g22606(.din(n40628), .dout(n40629));
  jand g22607(.dina(n40182), .dinb(n39920), .dout(n40630));
  jxor g22608(.dina(n39956), .dinb(n40189), .dout(n40631));
  jand g22609(.dina(n40631), .dinb(n40306), .dout(n40632));
  jor  g22610(.dina(n40632), .dinb(n40630), .dout(n40633));
  jand g22611(.dina(n40633), .dinb(n338), .dout(n40634));
  jnot g22612(.din(n40634), .dout(n40635));
  jand g22613(.dina(n40182), .dinb(n39926), .dout(n40636));
  jxor g22614(.dina(n39952), .dinb(n40187), .dout(n40637));
  jand g22615(.dina(n40637), .dinb(n40306), .dout(n40638));
  jor  g22616(.dina(n40638), .dinb(n40636), .dout(n40639));
  jand g22617(.dina(n40639), .dinb(n337), .dout(n40640));
  jnot g22618(.din(n40640), .dout(n40641));
  jand g22619(.dina(n40182), .dinb(n39932), .dout(n40642));
  jxor g22620(.dina(n39948), .dinb(n40185), .dout(n40643));
  jand g22621(.dina(n40643), .dinb(n40306), .dout(n40644));
  jor  g22622(.dina(n40644), .dinb(n40642), .dout(n40645));
  jand g22623(.dina(n40645), .dinb(n344), .dout(n40646));
  jnot g22624(.din(n40646), .dout(n40647));
  jand g22625(.dina(n40182), .dinb(n39939), .dout(n40648));
  jxor g22626(.dina(n40183), .dinb(n16327), .dout(n40649));
  jand g22627(.dina(n40649), .dinb(n40306), .dout(n40650));
  jor  g22628(.dina(n40650), .dinb(n40648), .dout(n40651));
  jand g22629(.dina(n40651), .dinb(n348), .dout(n40652));
  jnot g22630(.din(n40652), .dout(n40653));
  jor  g22631(.dina(n40182), .dinb(n18364), .dout(n40654));
  jand g22632(.dina(n40654), .dinb(a4 ), .dout(n40655));
  jor  g22633(.dina(n40182), .dinb(n16327), .dout(n40656));
  jnot g22634(.din(n40656), .dout(n40657));
  jor  g22635(.dina(n40657), .dinb(n40655), .dout(n40658));
  jand g22636(.dina(n40658), .dinb(n258), .dout(n40659));
  jnot g22637(.din(n40659), .dout(n40660));
  jand g22638(.dina(n40306), .dinb(b0 ), .dout(n40661));
  jor  g22639(.dina(n40661), .dinb(n16325), .dout(n40662));
  jand g22640(.dina(n40656), .dinb(n40662), .dout(n40663));
  jxor g22641(.dina(n40663), .dinb(n258), .dout(n40664));
  jor  g22642(.dina(n40664), .dinb(n16813), .dout(n40665));
  jand g22643(.dina(n40665), .dinb(n40660), .dout(n40666));
  jxor g22644(.dina(n40651), .dinb(n348), .dout(n40667));
  jnot g22645(.din(n40667), .dout(n40668));
  jor  g22646(.dina(n40668), .dinb(n40666), .dout(n40669));
  jand g22647(.dina(n40669), .dinb(n40653), .dout(n40670));
  jxor g22648(.dina(n40645), .dinb(n344), .dout(n40671));
  jnot g22649(.din(n40671), .dout(n40672));
  jor  g22650(.dina(n40672), .dinb(n40670), .dout(n40673));
  jand g22651(.dina(n40673), .dinb(n40647), .dout(n40674));
  jxor g22652(.dina(n40639), .dinb(n337), .dout(n40675));
  jnot g22653(.din(n40675), .dout(n40676));
  jor  g22654(.dina(n40676), .dinb(n40674), .dout(n40677));
  jand g22655(.dina(n40677), .dinb(n40641), .dout(n40678));
  jxor g22656(.dina(n40633), .dinb(n338), .dout(n40679));
  jnot g22657(.din(n40679), .dout(n40680));
  jor  g22658(.dina(n40680), .dinb(n40678), .dout(n40681));
  jand g22659(.dina(n40681), .dinb(n40635), .dout(n40682));
  jxor g22660(.dina(n40627), .dinb(n334), .dout(n40683));
  jnot g22661(.din(n40683), .dout(n40684));
  jor  g22662(.dina(n40684), .dinb(n40682), .dout(n40685));
  jand g22663(.dina(n40685), .dinb(n40629), .dout(n40686));
  jxor g22664(.dina(n40621), .dinb(n335), .dout(n40687));
  jnot g22665(.din(n40687), .dout(n40688));
  jor  g22666(.dina(n40688), .dinb(n40686), .dout(n40689));
  jand g22667(.dina(n40689), .dinb(n40623), .dout(n40690));
  jxor g22668(.dina(n40615), .dinb(n323), .dout(n40691));
  jnot g22669(.din(n40691), .dout(n40692));
  jor  g22670(.dina(n40692), .dinb(n40690), .dout(n40693));
  jand g22671(.dina(n40693), .dinb(n40617), .dout(n40694));
  jxor g22672(.dina(n40609), .dinb(n324), .dout(n40695));
  jnot g22673(.din(n40695), .dout(n40696));
  jor  g22674(.dina(n40696), .dinb(n40694), .dout(n40697));
  jand g22675(.dina(n40697), .dinb(n40611), .dout(n40698));
  jxor g22676(.dina(n40603), .dinb(n325), .dout(n40699));
  jnot g22677(.din(n40699), .dout(n40700));
  jor  g22678(.dina(n40700), .dinb(n40698), .dout(n40701));
  jand g22679(.dina(n40701), .dinb(n40605), .dout(n40702));
  jxor g22680(.dina(n40597), .dinb(n439), .dout(n40703));
  jnot g22681(.din(n40703), .dout(n40704));
  jor  g22682(.dina(n40704), .dinb(n40702), .dout(n40705));
  jand g22683(.dina(n40705), .dinb(n40599), .dout(n40706));
  jxor g22684(.dina(n40591), .dinb(n440), .dout(n40707));
  jnot g22685(.din(n40707), .dout(n40708));
  jor  g22686(.dina(n40708), .dinb(n40706), .dout(n40709));
  jand g22687(.dina(n40709), .dinb(n40593), .dout(n40710));
  jxor g22688(.dina(n40585), .dinb(n435), .dout(n40711));
  jnot g22689(.din(n40711), .dout(n40712));
  jor  g22690(.dina(n40712), .dinb(n40710), .dout(n40713));
  jand g22691(.dina(n40713), .dinb(n40587), .dout(n40714));
  jxor g22692(.dina(n40579), .dinb(n436), .dout(n40715));
  jnot g22693(.din(n40715), .dout(n40716));
  jor  g22694(.dina(n40716), .dinb(n40714), .dout(n40717));
  jand g22695(.dina(n40717), .dinb(n40581), .dout(n40718));
  jxor g22696(.dina(n40573), .dinb(n432), .dout(n40719));
  jnot g22697(.din(n40719), .dout(n40720));
  jor  g22698(.dina(n40720), .dinb(n40718), .dout(n40721));
  jand g22699(.dina(n40721), .dinb(n40575), .dout(n40722));
  jxor g22700(.dina(n40567), .dinb(n433), .dout(n40723));
  jnot g22701(.din(n40723), .dout(n40724));
  jor  g22702(.dina(n40724), .dinb(n40722), .dout(n40725));
  jand g22703(.dina(n40725), .dinb(n40569), .dout(n40726));
  jxor g22704(.dina(n40561), .dinb(n421), .dout(n40727));
  jnot g22705(.din(n40727), .dout(n40728));
  jor  g22706(.dina(n40728), .dinb(n40726), .dout(n40729));
  jand g22707(.dina(n40729), .dinb(n40563), .dout(n40730));
  jxor g22708(.dina(n40555), .dinb(n422), .dout(n40731));
  jnot g22709(.din(n40731), .dout(n40732));
  jor  g22710(.dina(n40732), .dinb(n40730), .dout(n40733));
  jand g22711(.dina(n40733), .dinb(n40557), .dout(n40734));
  jxor g22712(.dina(n40549), .dinb(n416), .dout(n40735));
  jnot g22713(.din(n40735), .dout(n40736));
  jor  g22714(.dina(n40736), .dinb(n40734), .dout(n40737));
  jand g22715(.dina(n40737), .dinb(n40551), .dout(n40738));
  jxor g22716(.dina(n40543), .dinb(n417), .dout(n40739));
  jnot g22717(.din(n40739), .dout(n40740));
  jor  g22718(.dina(n40740), .dinb(n40738), .dout(n40741));
  jand g22719(.dina(n40741), .dinb(n40545), .dout(n40742));
  jxor g22720(.dina(n40537), .dinb(n2547), .dout(n40743));
  jnot g22721(.din(n40743), .dout(n40744));
  jor  g22722(.dina(n40744), .dinb(n40742), .dout(n40745));
  jand g22723(.dina(n40745), .dinb(n40539), .dout(n40746));
  jxor g22724(.dina(n40531), .dinb(n2714), .dout(n40747));
  jnot g22725(.din(n40747), .dout(n40748));
  jor  g22726(.dina(n40748), .dinb(n40746), .dout(n40749));
  jand g22727(.dina(n40749), .dinb(n40533), .dout(n40750));
  jxor g22728(.dina(n40525), .dinb(n405), .dout(n40751));
  jnot g22729(.din(n40751), .dout(n40752));
  jor  g22730(.dina(n40752), .dinb(n40750), .dout(n40753));
  jand g22731(.dina(n40753), .dinb(n40527), .dout(n40754));
  jxor g22732(.dina(n40519), .dinb(n406), .dout(n40755));
  jnot g22733(.din(n40755), .dout(n40756));
  jor  g22734(.dina(n40756), .dinb(n40754), .dout(n40757));
  jand g22735(.dina(n40757), .dinb(n40521), .dout(n40758));
  jxor g22736(.dina(n40513), .dinb(n412), .dout(n40759));
  jnot g22737(.din(n40759), .dout(n40760));
  jor  g22738(.dina(n40760), .dinb(n40758), .dout(n40761));
  jand g22739(.dina(n40761), .dinb(n40515), .dout(n40762));
  jxor g22740(.dina(n40507), .dinb(n413), .dout(n40763));
  jnot g22741(.din(n40763), .dout(n40764));
  jor  g22742(.dina(n40764), .dinb(n40762), .dout(n40765));
  jand g22743(.dina(n40765), .dinb(n40509), .dout(n40766));
  jxor g22744(.dina(n40501), .dinb(n409), .dout(n40767));
  jnot g22745(.din(n40767), .dout(n40768));
  jor  g22746(.dina(n40768), .dinb(n40766), .dout(n40769));
  jand g22747(.dina(n40769), .dinb(n40503), .dout(n40770));
  jxor g22748(.dina(n40495), .dinb(n410), .dout(n40771));
  jnot g22749(.din(n40771), .dout(n40772));
  jor  g22750(.dina(n40772), .dinb(n40770), .dout(n40773));
  jand g22751(.dina(n40773), .dinb(n40497), .dout(n40774));
  jxor g22752(.dina(n40489), .dinb(n426), .dout(n40775));
  jnot g22753(.din(n40775), .dout(n40776));
  jor  g22754(.dina(n40776), .dinb(n40774), .dout(n40777));
  jand g22755(.dina(n40777), .dinb(n40491), .dout(n40778));
  jxor g22756(.dina(n40483), .dinb(n427), .dout(n40779));
  jnot g22757(.din(n40779), .dout(n40780));
  jor  g22758(.dina(n40780), .dinb(n40778), .dout(n40781));
  jand g22759(.dina(n40781), .dinb(n40485), .dout(n40782));
  jxor g22760(.dina(n40477), .dinb(n424), .dout(n40783));
  jnot g22761(.din(n40783), .dout(n40784));
  jor  g22762(.dina(n40784), .dinb(n40782), .dout(n40785));
  jand g22763(.dina(n40785), .dinb(n40479), .dout(n40786));
  jxor g22764(.dina(n40471), .dinb(n300), .dout(n40787));
  jnot g22765(.din(n40787), .dout(n40788));
  jor  g22766(.dina(n40788), .dinb(n40786), .dout(n40789));
  jand g22767(.dina(n40789), .dinb(n40473), .dout(n40790));
  jxor g22768(.dina(n40465), .dinb(n297), .dout(n40791));
  jnot g22769(.din(n40791), .dout(n40792));
  jor  g22770(.dina(n40792), .dinb(n40790), .dout(n40793));
  jand g22771(.dina(n40793), .dinb(n40467), .dout(n40794));
  jxor g22772(.dina(n40459), .dinb(n298), .dout(n40795));
  jnot g22773(.din(n40795), .dout(n40796));
  jor  g22774(.dina(n40796), .dinb(n40794), .dout(n40797));
  jand g22775(.dina(n40797), .dinb(n40461), .dout(n40798));
  jxor g22776(.dina(n40453), .dinb(n301), .dout(n40799));
  jnot g22777(.din(n40799), .dout(n40800));
  jor  g22778(.dina(n40800), .dinb(n40798), .dout(n40801));
  jand g22779(.dina(n40801), .dinb(n40455), .dout(n40802));
  jxor g22780(.dina(n40447), .dinb(n293), .dout(n40803));
  jnot g22781(.din(n40803), .dout(n40804));
  jor  g22782(.dina(n40804), .dinb(n40802), .dout(n40805));
  jand g22783(.dina(n40805), .dinb(n40449), .dout(n40806));
  jxor g22784(.dina(n40441), .dinb(n294), .dout(n40807));
  jnot g22785(.din(n40807), .dout(n40808));
  jor  g22786(.dina(n40808), .dinb(n40806), .dout(n40809));
  jand g22787(.dina(n40809), .dinb(n40443), .dout(n40810));
  jxor g22788(.dina(n40435), .dinb(n290), .dout(n40811));
  jnot g22789(.din(n40811), .dout(n40812));
  jor  g22790(.dina(n40812), .dinb(n40810), .dout(n40813));
  jand g22791(.dina(n40813), .dinb(n40437), .dout(n40814));
  jxor g22792(.dina(n40429), .dinb(n291), .dout(n40815));
  jnot g22793(.din(n40815), .dout(n40816));
  jor  g22794(.dina(n40816), .dinb(n40814), .dout(n40817));
  jand g22795(.dina(n40817), .dinb(n40431), .dout(n40818));
  jxor g22796(.dina(n40423), .dinb(n284), .dout(n40819));
  jnot g22797(.din(n40819), .dout(n40820));
  jor  g22798(.dina(n40820), .dinb(n40818), .dout(n40821));
  jand g22799(.dina(n40821), .dinb(n40425), .dout(n40822));
  jxor g22800(.dina(n40417), .dinb(n285), .dout(n40823));
  jnot g22801(.din(n40823), .dout(n40824));
  jor  g22802(.dina(n40824), .dinb(n40822), .dout(n40825));
  jand g22803(.dina(n40825), .dinb(n40419), .dout(n40826));
  jxor g22804(.dina(n40411), .dinb(n281), .dout(n40827));
  jnot g22805(.din(n40827), .dout(n40828));
  jor  g22806(.dina(n40828), .dinb(n40826), .dout(n40829));
  jand g22807(.dina(n40829), .dinb(n40413), .dout(n40830));
  jxor g22808(.dina(n40405), .dinb(n282), .dout(n40831));
  jnot g22809(.din(n40831), .dout(n40832));
  jor  g22810(.dina(n40832), .dinb(n40830), .dout(n40833));
  jand g22811(.dina(n40833), .dinb(n40407), .dout(n40834));
  jxor g22812(.dina(n40399), .dinb(n397), .dout(n40835));
  jnot g22813(.din(n40835), .dout(n40836));
  jor  g22814(.dina(n40836), .dinb(n40834), .dout(n40837));
  jand g22815(.dina(n40837), .dinb(n40401), .dout(n40838));
  jxor g22816(.dina(n40393), .dinb(n513), .dout(n40839));
  jnot g22817(.din(n40839), .dout(n40840));
  jor  g22818(.dina(n40840), .dinb(n40838), .dout(n40841));
  jand g22819(.dina(n40841), .dinb(n40395), .dout(n40842));
  jxor g22820(.dina(n40387), .dinb(n514), .dout(n40843));
  jnot g22821(.din(n40843), .dout(n40844));
  jor  g22822(.dina(n40844), .dinb(n40842), .dout(n40845));
  jand g22823(.dina(n40845), .dinb(n40389), .dout(n40846));
  jxor g22824(.dina(n40381), .dinb(n510), .dout(n40847));
  jnot g22825(.din(n40847), .dout(n40848));
  jor  g22826(.dina(n40848), .dinb(n40846), .dout(n40849));
  jand g22827(.dina(n40849), .dinb(n40383), .dout(n40850));
  jxor g22828(.dina(n40375), .dinb(n396), .dout(n40851));
  jnot g22829(.din(n40851), .dout(n40852));
  jor  g22830(.dina(n40852), .dinb(n40850), .dout(n40853));
  jand g22831(.dina(n40853), .dinb(n40377), .dout(n40854));
  jxor g22832(.dina(n40369), .dinb(n383), .dout(n40855));
  jnot g22833(.din(n40855), .dout(n40856));
  jor  g22834(.dina(n40856), .dinb(n40854), .dout(n40857));
  jand g22835(.dina(n40857), .dinb(n40371), .dout(n40858));
  jxor g22836(.dina(n40363), .dinb(n12211), .dout(n40859));
  jnot g22837(.din(n40859), .dout(n40860));
  jor  g22838(.dina(n40860), .dinb(n40858), .dout(n40861));
  jand g22839(.dina(n40861), .dinb(n40365), .dout(n40862));
  jxor g22840(.dina(n40357), .dinb(n12214), .dout(n40863));
  jnot g22841(.din(n40863), .dout(n40864));
  jor  g22842(.dina(n40864), .dinb(n40862), .dout(n40865));
  jand g22843(.dina(n40865), .dinb(n40359), .dout(n40866));
  jxor g22844(.dina(n40351), .dinb(n384), .dout(n40867));
  jnot g22845(.din(n40867), .dout(n40868));
  jor  g22846(.dina(n40868), .dinb(n40866), .dout(n40869));
  jand g22847(.dina(n40869), .dinb(n40353), .dout(n40870));
  jxor g22848(.dina(n40345), .dinb(n374), .dout(n40871));
  jnot g22849(.din(n40871), .dout(n40872));
  jor  g22850(.dina(n40872), .dinb(n40870), .dout(n40873));
  jand g22851(.dina(n40873), .dinb(n40347), .dout(n40874));
  jxor g22852(.dina(n40339), .dinb(n376), .dout(n40875));
  jnot g22853(.din(n40875), .dout(n40876));
  jor  g22854(.dina(n40876), .dinb(n40874), .dout(n40877));
  jand g22855(.dina(n40877), .dinb(n40341), .dout(n40878));
  jxor g22856(.dina(n40333), .dinb(n377), .dout(n40879));
  jnot g22857(.din(n40879), .dout(n40880));
  jor  g22858(.dina(n40880), .dinb(n40878), .dout(n40881));
  jand g22859(.dina(n40881), .dinb(n40335), .dout(n40882));
  jxor g22860(.dina(n40327), .dinb(n375), .dout(n40883));
  jnot g22861(.din(n40883), .dout(n40884));
  jor  g22862(.dina(n40884), .dinb(n40882), .dout(n40885));
  jand g22863(.dina(n40885), .dinb(n40329), .dout(n40886));
  jxor g22864(.dina(n40321), .dinb(n362), .dout(n40887));
  jnot g22865(.din(n40887), .dout(n40888));
  jor  g22866(.dina(n40888), .dinb(n40886), .dout(n40889));
  jand g22867(.dina(n40889), .dinb(n40323), .dout(n40890));
  jxor g22868(.dina(n40315), .dinb(n363), .dout(n40891));
  jnot g22869(.din(n40891), .dout(n40892));
  jor  g22870(.dina(n40892), .dinb(n40890), .dout(n40893));
  jand g22871(.dina(n40893), .dinb(n40317), .dout(n40894));
  jxor g22872(.dina(n40309), .dinb(n365), .dout(n40895));
  jnot g22873(.din(n40895), .dout(n40896));
  jor  g22874(.dina(n40896), .dinb(n40894), .dout(n40897));
  jand g22875(.dina(n40897), .dinb(n40311), .dout(n40898));
  jand g22876(.dina(n40302), .dinb(n366), .dout(n40899));
  jnot g22877(.din(n40899), .dout(n40900));
  jand g22878(.dina(n40900), .dinb(n40898), .dout(n40901));
  jnot g22879(.din(n40302), .dout(n40902));
  jand g22880(.dina(n40902), .dinb(b60 ), .dout(n40903));
  jor  g22881(.dina(n40903), .dinb(n263), .dout(n40904));
  jor  g22882(.dina(n40904), .dinb(n40901), .dout(n40905));
  jxor g22883(.dina(n40663), .dinb(b1 ), .dout(n40906));
  jand g22884(.dina(n40906), .dinb(n16814), .dout(n40907));
  jor  g22885(.dina(n40907), .dinb(n40659), .dout(n40908));
  jand g22886(.dina(n40667), .dinb(n40908), .dout(n40909));
  jor  g22887(.dina(n40909), .dinb(n40652), .dout(n40910));
  jand g22888(.dina(n40671), .dinb(n40910), .dout(n40911));
  jor  g22889(.dina(n40911), .dinb(n40646), .dout(n40912));
  jand g22890(.dina(n40675), .dinb(n40912), .dout(n40913));
  jor  g22891(.dina(n40913), .dinb(n40640), .dout(n40914));
  jand g22892(.dina(n40679), .dinb(n40914), .dout(n40915));
  jor  g22893(.dina(n40915), .dinb(n40634), .dout(n40916));
  jand g22894(.dina(n40683), .dinb(n40916), .dout(n40917));
  jor  g22895(.dina(n40917), .dinb(n40628), .dout(n40918));
  jand g22896(.dina(n40687), .dinb(n40918), .dout(n40919));
  jor  g22897(.dina(n40919), .dinb(n40622), .dout(n40920));
  jand g22898(.dina(n40691), .dinb(n40920), .dout(n40921));
  jor  g22899(.dina(n40921), .dinb(n40616), .dout(n40922));
  jand g22900(.dina(n40695), .dinb(n40922), .dout(n40923));
  jor  g22901(.dina(n40923), .dinb(n40610), .dout(n40924));
  jand g22902(.dina(n40699), .dinb(n40924), .dout(n40925));
  jor  g22903(.dina(n40925), .dinb(n40604), .dout(n40926));
  jand g22904(.dina(n40703), .dinb(n40926), .dout(n40927));
  jor  g22905(.dina(n40927), .dinb(n40598), .dout(n40928));
  jand g22906(.dina(n40707), .dinb(n40928), .dout(n40929));
  jor  g22907(.dina(n40929), .dinb(n40592), .dout(n40930));
  jand g22908(.dina(n40711), .dinb(n40930), .dout(n40931));
  jor  g22909(.dina(n40931), .dinb(n40586), .dout(n40932));
  jand g22910(.dina(n40715), .dinb(n40932), .dout(n40933));
  jor  g22911(.dina(n40933), .dinb(n40580), .dout(n40934));
  jand g22912(.dina(n40719), .dinb(n40934), .dout(n40935));
  jor  g22913(.dina(n40935), .dinb(n40574), .dout(n40936));
  jand g22914(.dina(n40723), .dinb(n40936), .dout(n40937));
  jor  g22915(.dina(n40937), .dinb(n40568), .dout(n40938));
  jand g22916(.dina(n40727), .dinb(n40938), .dout(n40939));
  jor  g22917(.dina(n40939), .dinb(n40562), .dout(n40940));
  jand g22918(.dina(n40731), .dinb(n40940), .dout(n40941));
  jor  g22919(.dina(n40941), .dinb(n40556), .dout(n40942));
  jand g22920(.dina(n40735), .dinb(n40942), .dout(n40943));
  jor  g22921(.dina(n40943), .dinb(n40550), .dout(n40944));
  jand g22922(.dina(n40739), .dinb(n40944), .dout(n40945));
  jor  g22923(.dina(n40945), .dinb(n40544), .dout(n40946));
  jand g22924(.dina(n40743), .dinb(n40946), .dout(n40947));
  jor  g22925(.dina(n40947), .dinb(n40538), .dout(n40948));
  jand g22926(.dina(n40747), .dinb(n40948), .dout(n40949));
  jor  g22927(.dina(n40949), .dinb(n40532), .dout(n40950));
  jand g22928(.dina(n40751), .dinb(n40950), .dout(n40951));
  jor  g22929(.dina(n40951), .dinb(n40526), .dout(n40952));
  jand g22930(.dina(n40755), .dinb(n40952), .dout(n40953));
  jor  g22931(.dina(n40953), .dinb(n40520), .dout(n40954));
  jand g22932(.dina(n40759), .dinb(n40954), .dout(n40955));
  jor  g22933(.dina(n40955), .dinb(n40514), .dout(n40956));
  jand g22934(.dina(n40763), .dinb(n40956), .dout(n40957));
  jor  g22935(.dina(n40957), .dinb(n40508), .dout(n40958));
  jand g22936(.dina(n40767), .dinb(n40958), .dout(n40959));
  jor  g22937(.dina(n40959), .dinb(n40502), .dout(n40960));
  jand g22938(.dina(n40771), .dinb(n40960), .dout(n40961));
  jor  g22939(.dina(n40961), .dinb(n40496), .dout(n40962));
  jand g22940(.dina(n40775), .dinb(n40962), .dout(n40963));
  jor  g22941(.dina(n40963), .dinb(n40490), .dout(n40964));
  jand g22942(.dina(n40779), .dinb(n40964), .dout(n40965));
  jor  g22943(.dina(n40965), .dinb(n40484), .dout(n40966));
  jand g22944(.dina(n40783), .dinb(n40966), .dout(n40967));
  jor  g22945(.dina(n40967), .dinb(n40478), .dout(n40968));
  jand g22946(.dina(n40787), .dinb(n40968), .dout(n40969));
  jor  g22947(.dina(n40969), .dinb(n40472), .dout(n40970));
  jand g22948(.dina(n40791), .dinb(n40970), .dout(n40971));
  jor  g22949(.dina(n40971), .dinb(n40466), .dout(n40972));
  jand g22950(.dina(n40795), .dinb(n40972), .dout(n40973));
  jor  g22951(.dina(n40973), .dinb(n40460), .dout(n40974));
  jand g22952(.dina(n40799), .dinb(n40974), .dout(n40975));
  jor  g22953(.dina(n40975), .dinb(n40454), .dout(n40976));
  jand g22954(.dina(n40803), .dinb(n40976), .dout(n40977));
  jor  g22955(.dina(n40977), .dinb(n40448), .dout(n40978));
  jand g22956(.dina(n40807), .dinb(n40978), .dout(n40979));
  jor  g22957(.dina(n40979), .dinb(n40442), .dout(n40980));
  jand g22958(.dina(n40811), .dinb(n40980), .dout(n40981));
  jor  g22959(.dina(n40981), .dinb(n40436), .dout(n40982));
  jand g22960(.dina(n40815), .dinb(n40982), .dout(n40983));
  jor  g22961(.dina(n40983), .dinb(n40430), .dout(n40984));
  jand g22962(.dina(n40819), .dinb(n40984), .dout(n40985));
  jor  g22963(.dina(n40985), .dinb(n40424), .dout(n40986));
  jand g22964(.dina(n40823), .dinb(n40986), .dout(n40987));
  jor  g22965(.dina(n40987), .dinb(n40418), .dout(n40988));
  jand g22966(.dina(n40827), .dinb(n40988), .dout(n40989));
  jor  g22967(.dina(n40989), .dinb(n40412), .dout(n40990));
  jand g22968(.dina(n40831), .dinb(n40990), .dout(n40991));
  jor  g22969(.dina(n40991), .dinb(n40406), .dout(n40992));
  jand g22970(.dina(n40835), .dinb(n40992), .dout(n40993));
  jor  g22971(.dina(n40993), .dinb(n40400), .dout(n40994));
  jand g22972(.dina(n40839), .dinb(n40994), .dout(n40995));
  jor  g22973(.dina(n40995), .dinb(n40394), .dout(n40996));
  jand g22974(.dina(n40843), .dinb(n40996), .dout(n40997));
  jor  g22975(.dina(n40997), .dinb(n40388), .dout(n40998));
  jand g22976(.dina(n40847), .dinb(n40998), .dout(n40999));
  jor  g22977(.dina(n40999), .dinb(n40382), .dout(n41000));
  jand g22978(.dina(n40851), .dinb(n41000), .dout(n41001));
  jor  g22979(.dina(n41001), .dinb(n40376), .dout(n41002));
  jand g22980(.dina(n40855), .dinb(n41002), .dout(n41003));
  jor  g22981(.dina(n41003), .dinb(n40370), .dout(n41004));
  jand g22982(.dina(n40859), .dinb(n41004), .dout(n41005));
  jor  g22983(.dina(n41005), .dinb(n40364), .dout(n41006));
  jand g22984(.dina(n40863), .dinb(n41006), .dout(n41007));
  jor  g22985(.dina(n41007), .dinb(n40358), .dout(n41008));
  jand g22986(.dina(n40867), .dinb(n41008), .dout(n41009));
  jor  g22987(.dina(n41009), .dinb(n40352), .dout(n41010));
  jand g22988(.dina(n40871), .dinb(n41010), .dout(n41011));
  jor  g22989(.dina(n41011), .dinb(n40346), .dout(n41012));
  jand g22990(.dina(n40875), .dinb(n41012), .dout(n41013));
  jor  g22991(.dina(n41013), .dinb(n40340), .dout(n41014));
  jand g22992(.dina(n40879), .dinb(n41014), .dout(n41015));
  jor  g22993(.dina(n41015), .dinb(n40334), .dout(n41016));
  jand g22994(.dina(n40883), .dinb(n41016), .dout(n41017));
  jor  g22995(.dina(n41017), .dinb(n40328), .dout(n41018));
  jand g22996(.dina(n40887), .dinb(n41018), .dout(n41019));
  jor  g22997(.dina(n41019), .dinb(n40322), .dout(n41020));
  jand g22998(.dina(n40891), .dinb(n41020), .dout(n41021));
  jor  g22999(.dina(n41021), .dinb(n40316), .dout(n41022));
  jand g23000(.dina(n40895), .dinb(n41022), .dout(n41023));
  jor  g23001(.dina(n41023), .dinb(n40310), .dout(n41024));
  jand g23002(.dina(n41024), .dinb(n371), .dout(n41025));
  jor  g23003(.dina(n41025), .dinb(n40905), .dout(n41026));
  jand g23004(.dina(n41026), .dinb(n40302), .dout(n41027));
  jand g23005(.dina(n40905), .dinb(n40309), .dout(n41028));
  jor  g23006(.dina(n40899), .dinb(n41024), .dout(n41029));
  jnot g23007(.din(n40904), .dout(n41030));
  jand g23008(.dina(n41030), .dinb(n41029), .dout(n41031));
  jxor g23009(.dina(n40895), .dinb(n41022), .dout(n41032));
  jand g23010(.dina(n41032), .dinb(n41031), .dout(n41033));
  jor  g23011(.dina(n41033), .dinb(n41028), .dout(n41034));
  jand g23012(.dina(n41034), .dinb(n366), .dout(n41035));
  jnot g23013(.din(n41035), .dout(n41036));
  jand g23014(.dina(n40905), .dinb(n40315), .dout(n41037));
  jxor g23015(.dina(n40891), .dinb(n41020), .dout(n41038));
  jand g23016(.dina(n41038), .dinb(n41031), .dout(n41039));
  jor  g23017(.dina(n41039), .dinb(n41037), .dout(n41040));
  jand g23018(.dina(n41040), .dinb(n365), .dout(n41041));
  jnot g23019(.din(n41041), .dout(n41042));
  jand g23020(.dina(n40905), .dinb(n40321), .dout(n41043));
  jxor g23021(.dina(n40887), .dinb(n41018), .dout(n41044));
  jand g23022(.dina(n41044), .dinb(n41031), .dout(n41045));
  jor  g23023(.dina(n41045), .dinb(n41043), .dout(n41046));
  jand g23024(.dina(n41046), .dinb(n363), .dout(n41047));
  jnot g23025(.din(n41047), .dout(n41048));
  jand g23026(.dina(n40905), .dinb(n40327), .dout(n41049));
  jxor g23027(.dina(n40883), .dinb(n41016), .dout(n41050));
  jand g23028(.dina(n41050), .dinb(n41031), .dout(n41051));
  jor  g23029(.dina(n41051), .dinb(n41049), .dout(n41052));
  jand g23030(.dina(n41052), .dinb(n362), .dout(n41053));
  jnot g23031(.din(n41053), .dout(n41054));
  jand g23032(.dina(n40905), .dinb(n40333), .dout(n41055));
  jxor g23033(.dina(n40879), .dinb(n41014), .dout(n41056));
  jand g23034(.dina(n41056), .dinb(n41031), .dout(n41057));
  jor  g23035(.dina(n41057), .dinb(n41055), .dout(n41058));
  jand g23036(.dina(n41058), .dinb(n375), .dout(n41059));
  jnot g23037(.din(n41059), .dout(n41060));
  jand g23038(.dina(n40905), .dinb(n40339), .dout(n41061));
  jxor g23039(.dina(n40875), .dinb(n41012), .dout(n41062));
  jand g23040(.dina(n41062), .dinb(n41031), .dout(n41063));
  jor  g23041(.dina(n41063), .dinb(n41061), .dout(n41064));
  jand g23042(.dina(n41064), .dinb(n377), .dout(n41065));
  jnot g23043(.din(n41065), .dout(n41066));
  jand g23044(.dina(n40905), .dinb(n40345), .dout(n41067));
  jxor g23045(.dina(n40871), .dinb(n41010), .dout(n41068));
  jand g23046(.dina(n41068), .dinb(n41031), .dout(n41069));
  jor  g23047(.dina(n41069), .dinb(n41067), .dout(n41070));
  jand g23048(.dina(n41070), .dinb(n376), .dout(n41071));
  jnot g23049(.din(n41071), .dout(n41072));
  jand g23050(.dina(n40905), .dinb(n40351), .dout(n41073));
  jxor g23051(.dina(n40867), .dinb(n41008), .dout(n41074));
  jand g23052(.dina(n41074), .dinb(n41031), .dout(n41075));
  jor  g23053(.dina(n41075), .dinb(n41073), .dout(n41076));
  jand g23054(.dina(n41076), .dinb(n374), .dout(n41077));
  jnot g23055(.din(n41077), .dout(n41078));
  jand g23056(.dina(n40905), .dinb(n40357), .dout(n41079));
  jxor g23057(.dina(n40863), .dinb(n41006), .dout(n41080));
  jand g23058(.dina(n41080), .dinb(n41031), .dout(n41081));
  jor  g23059(.dina(n41081), .dinb(n41079), .dout(n41082));
  jand g23060(.dina(n41082), .dinb(n384), .dout(n41083));
  jnot g23061(.din(n41083), .dout(n41084));
  jand g23062(.dina(n40905), .dinb(n40363), .dout(n41085));
  jxor g23063(.dina(n40859), .dinb(n41004), .dout(n41086));
  jand g23064(.dina(n41086), .dinb(n41031), .dout(n41087));
  jor  g23065(.dina(n41087), .dinb(n41085), .dout(n41088));
  jand g23066(.dina(n41088), .dinb(n12214), .dout(n41089));
  jnot g23067(.din(n41089), .dout(n41090));
  jand g23068(.dina(n40905), .dinb(n40369), .dout(n41091));
  jxor g23069(.dina(n40855), .dinb(n41002), .dout(n41092));
  jand g23070(.dina(n41092), .dinb(n41031), .dout(n41093));
  jor  g23071(.dina(n41093), .dinb(n41091), .dout(n41094));
  jand g23072(.dina(n41094), .dinb(n12211), .dout(n41095));
  jnot g23073(.din(n41095), .dout(n41096));
  jand g23074(.dina(n40905), .dinb(n40375), .dout(n41097));
  jxor g23075(.dina(n40851), .dinb(n41000), .dout(n41098));
  jand g23076(.dina(n41098), .dinb(n41031), .dout(n41099));
  jor  g23077(.dina(n41099), .dinb(n41097), .dout(n41100));
  jand g23078(.dina(n41100), .dinb(n383), .dout(n41101));
  jnot g23079(.din(n41101), .dout(n41102));
  jand g23080(.dina(n40905), .dinb(n40381), .dout(n41103));
  jxor g23081(.dina(n40847), .dinb(n40998), .dout(n41104));
  jand g23082(.dina(n41104), .dinb(n41031), .dout(n41105));
  jor  g23083(.dina(n41105), .dinb(n41103), .dout(n41106));
  jand g23084(.dina(n41106), .dinb(n396), .dout(n41107));
  jnot g23085(.din(n41107), .dout(n41108));
  jand g23086(.dina(n40905), .dinb(n40387), .dout(n41109));
  jxor g23087(.dina(n40843), .dinb(n40996), .dout(n41110));
  jand g23088(.dina(n41110), .dinb(n41031), .dout(n41111));
  jor  g23089(.dina(n41111), .dinb(n41109), .dout(n41112));
  jand g23090(.dina(n41112), .dinb(n510), .dout(n41113));
  jnot g23091(.din(n41113), .dout(n41114));
  jand g23092(.dina(n40905), .dinb(n40393), .dout(n41115));
  jxor g23093(.dina(n40839), .dinb(n40994), .dout(n41116));
  jand g23094(.dina(n41116), .dinb(n41031), .dout(n41117));
  jor  g23095(.dina(n41117), .dinb(n41115), .dout(n41118));
  jand g23096(.dina(n41118), .dinb(n514), .dout(n41119));
  jnot g23097(.din(n41119), .dout(n41120));
  jand g23098(.dina(n40905), .dinb(n40399), .dout(n41121));
  jxor g23099(.dina(n40835), .dinb(n40992), .dout(n41122));
  jand g23100(.dina(n41122), .dinb(n41031), .dout(n41123));
  jor  g23101(.dina(n41123), .dinb(n41121), .dout(n41124));
  jand g23102(.dina(n41124), .dinb(n513), .dout(n41125));
  jnot g23103(.din(n41125), .dout(n41126));
  jand g23104(.dina(n40905), .dinb(n40405), .dout(n41127));
  jxor g23105(.dina(n40831), .dinb(n40990), .dout(n41128));
  jand g23106(.dina(n41128), .dinb(n41031), .dout(n41129));
  jor  g23107(.dina(n41129), .dinb(n41127), .dout(n41130));
  jand g23108(.dina(n41130), .dinb(n397), .dout(n41131));
  jnot g23109(.din(n41131), .dout(n41132));
  jand g23110(.dina(n40905), .dinb(n40411), .dout(n41133));
  jxor g23111(.dina(n40827), .dinb(n40988), .dout(n41134));
  jand g23112(.dina(n41134), .dinb(n41031), .dout(n41135));
  jor  g23113(.dina(n41135), .dinb(n41133), .dout(n41136));
  jand g23114(.dina(n41136), .dinb(n282), .dout(n41137));
  jnot g23115(.din(n41137), .dout(n41138));
  jand g23116(.dina(n40905), .dinb(n40417), .dout(n41139));
  jxor g23117(.dina(n40823), .dinb(n40986), .dout(n41140));
  jand g23118(.dina(n41140), .dinb(n41031), .dout(n41141));
  jor  g23119(.dina(n41141), .dinb(n41139), .dout(n41142));
  jand g23120(.dina(n41142), .dinb(n281), .dout(n41143));
  jnot g23121(.din(n41143), .dout(n41144));
  jand g23122(.dina(n40905), .dinb(n40423), .dout(n41145));
  jxor g23123(.dina(n40819), .dinb(n40984), .dout(n41146));
  jand g23124(.dina(n41146), .dinb(n41031), .dout(n41147));
  jor  g23125(.dina(n41147), .dinb(n41145), .dout(n41148));
  jand g23126(.dina(n41148), .dinb(n285), .dout(n41149));
  jnot g23127(.din(n41149), .dout(n41150));
  jand g23128(.dina(n40905), .dinb(n40429), .dout(n41151));
  jxor g23129(.dina(n40815), .dinb(n40982), .dout(n41152));
  jand g23130(.dina(n41152), .dinb(n41031), .dout(n41153));
  jor  g23131(.dina(n41153), .dinb(n41151), .dout(n41154));
  jand g23132(.dina(n41154), .dinb(n284), .dout(n41155));
  jnot g23133(.din(n41155), .dout(n41156));
  jand g23134(.dina(n40905), .dinb(n40435), .dout(n41157));
  jxor g23135(.dina(n40811), .dinb(n40980), .dout(n41158));
  jand g23136(.dina(n41158), .dinb(n41031), .dout(n41159));
  jor  g23137(.dina(n41159), .dinb(n41157), .dout(n41160));
  jand g23138(.dina(n41160), .dinb(n291), .dout(n41161));
  jnot g23139(.din(n41161), .dout(n41162));
  jand g23140(.dina(n40905), .dinb(n40441), .dout(n41163));
  jxor g23141(.dina(n40807), .dinb(n40978), .dout(n41164));
  jand g23142(.dina(n41164), .dinb(n41031), .dout(n41165));
  jor  g23143(.dina(n41165), .dinb(n41163), .dout(n41166));
  jand g23144(.dina(n41166), .dinb(n290), .dout(n41167));
  jnot g23145(.din(n41167), .dout(n41168));
  jand g23146(.dina(n40905), .dinb(n40447), .dout(n41169));
  jxor g23147(.dina(n40803), .dinb(n40976), .dout(n41170));
  jand g23148(.dina(n41170), .dinb(n41031), .dout(n41171));
  jor  g23149(.dina(n41171), .dinb(n41169), .dout(n41172));
  jand g23150(.dina(n41172), .dinb(n294), .dout(n41173));
  jnot g23151(.din(n41173), .dout(n41174));
  jand g23152(.dina(n40905), .dinb(n40453), .dout(n41175));
  jxor g23153(.dina(n40799), .dinb(n40974), .dout(n41176));
  jand g23154(.dina(n41176), .dinb(n41031), .dout(n41177));
  jor  g23155(.dina(n41177), .dinb(n41175), .dout(n41178));
  jand g23156(.dina(n41178), .dinb(n293), .dout(n41179));
  jnot g23157(.din(n41179), .dout(n41180));
  jand g23158(.dina(n40905), .dinb(n40459), .dout(n41181));
  jxor g23159(.dina(n40795), .dinb(n40972), .dout(n41182));
  jand g23160(.dina(n41182), .dinb(n41031), .dout(n41183));
  jor  g23161(.dina(n41183), .dinb(n41181), .dout(n41184));
  jand g23162(.dina(n41184), .dinb(n301), .dout(n41185));
  jnot g23163(.din(n41185), .dout(n41186));
  jand g23164(.dina(n40905), .dinb(n40465), .dout(n41187));
  jxor g23165(.dina(n40791), .dinb(n40970), .dout(n41188));
  jand g23166(.dina(n41188), .dinb(n41031), .dout(n41189));
  jor  g23167(.dina(n41189), .dinb(n41187), .dout(n41190));
  jand g23168(.dina(n41190), .dinb(n298), .dout(n41191));
  jnot g23169(.din(n41191), .dout(n41192));
  jand g23170(.dina(n40905), .dinb(n40471), .dout(n41193));
  jxor g23171(.dina(n40787), .dinb(n40968), .dout(n41194));
  jand g23172(.dina(n41194), .dinb(n41031), .dout(n41195));
  jor  g23173(.dina(n41195), .dinb(n41193), .dout(n41196));
  jand g23174(.dina(n41196), .dinb(n297), .dout(n41197));
  jnot g23175(.din(n41197), .dout(n41198));
  jand g23176(.dina(n40905), .dinb(n40477), .dout(n41199));
  jxor g23177(.dina(n40783), .dinb(n40966), .dout(n41200));
  jand g23178(.dina(n41200), .dinb(n41031), .dout(n41201));
  jor  g23179(.dina(n41201), .dinb(n41199), .dout(n41202));
  jand g23180(.dina(n41202), .dinb(n300), .dout(n41203));
  jnot g23181(.din(n41203), .dout(n41204));
  jand g23182(.dina(n40905), .dinb(n40483), .dout(n41205));
  jxor g23183(.dina(n40779), .dinb(n40964), .dout(n41206));
  jand g23184(.dina(n41206), .dinb(n41031), .dout(n41207));
  jor  g23185(.dina(n41207), .dinb(n41205), .dout(n41208));
  jand g23186(.dina(n41208), .dinb(n424), .dout(n41209));
  jnot g23187(.din(n41209), .dout(n41210));
  jand g23188(.dina(n40905), .dinb(n40489), .dout(n41211));
  jxor g23189(.dina(n40775), .dinb(n40962), .dout(n41212));
  jand g23190(.dina(n41212), .dinb(n41031), .dout(n41213));
  jor  g23191(.dina(n41213), .dinb(n41211), .dout(n41214));
  jand g23192(.dina(n41214), .dinb(n427), .dout(n41215));
  jnot g23193(.din(n41215), .dout(n41216));
  jand g23194(.dina(n40905), .dinb(n40495), .dout(n41217));
  jxor g23195(.dina(n40771), .dinb(n40960), .dout(n41218));
  jand g23196(.dina(n41218), .dinb(n41031), .dout(n41219));
  jor  g23197(.dina(n41219), .dinb(n41217), .dout(n41220));
  jand g23198(.dina(n41220), .dinb(n426), .dout(n41221));
  jnot g23199(.din(n41221), .dout(n41222));
  jand g23200(.dina(n40905), .dinb(n40501), .dout(n41223));
  jxor g23201(.dina(n40767), .dinb(n40958), .dout(n41224));
  jand g23202(.dina(n41224), .dinb(n41031), .dout(n41225));
  jor  g23203(.dina(n41225), .dinb(n41223), .dout(n41226));
  jand g23204(.dina(n41226), .dinb(n410), .dout(n41227));
  jnot g23205(.din(n41227), .dout(n41228));
  jand g23206(.dina(n40905), .dinb(n40507), .dout(n41229));
  jxor g23207(.dina(n40763), .dinb(n40956), .dout(n41230));
  jand g23208(.dina(n41230), .dinb(n41031), .dout(n41231));
  jor  g23209(.dina(n41231), .dinb(n41229), .dout(n41232));
  jand g23210(.dina(n41232), .dinb(n409), .dout(n41233));
  jnot g23211(.din(n41233), .dout(n41234));
  jand g23212(.dina(n40905), .dinb(n40513), .dout(n41235));
  jxor g23213(.dina(n40759), .dinb(n40954), .dout(n41236));
  jand g23214(.dina(n41236), .dinb(n41031), .dout(n41237));
  jor  g23215(.dina(n41237), .dinb(n41235), .dout(n41238));
  jand g23216(.dina(n41238), .dinb(n413), .dout(n41239));
  jnot g23217(.din(n41239), .dout(n41240));
  jand g23218(.dina(n40905), .dinb(n40519), .dout(n41241));
  jxor g23219(.dina(n40755), .dinb(n40952), .dout(n41242));
  jand g23220(.dina(n41242), .dinb(n41031), .dout(n41243));
  jor  g23221(.dina(n41243), .dinb(n41241), .dout(n41244));
  jand g23222(.dina(n41244), .dinb(n412), .dout(n41245));
  jnot g23223(.din(n41245), .dout(n41246));
  jand g23224(.dina(n40905), .dinb(n40525), .dout(n41247));
  jxor g23225(.dina(n40751), .dinb(n40950), .dout(n41248));
  jand g23226(.dina(n41248), .dinb(n41031), .dout(n41249));
  jor  g23227(.dina(n41249), .dinb(n41247), .dout(n41250));
  jand g23228(.dina(n41250), .dinb(n406), .dout(n41251));
  jnot g23229(.din(n41251), .dout(n41252));
  jand g23230(.dina(n40905), .dinb(n40531), .dout(n41253));
  jxor g23231(.dina(n40747), .dinb(n40948), .dout(n41254));
  jand g23232(.dina(n41254), .dinb(n41031), .dout(n41255));
  jor  g23233(.dina(n41255), .dinb(n41253), .dout(n41256));
  jand g23234(.dina(n41256), .dinb(n405), .dout(n41257));
  jnot g23235(.din(n41257), .dout(n41258));
  jand g23236(.dina(n40905), .dinb(n40537), .dout(n41259));
  jxor g23237(.dina(n40743), .dinb(n40946), .dout(n41260));
  jand g23238(.dina(n41260), .dinb(n41031), .dout(n41261));
  jor  g23239(.dina(n41261), .dinb(n41259), .dout(n41262));
  jand g23240(.dina(n41262), .dinb(n2714), .dout(n41263));
  jnot g23241(.din(n41263), .dout(n41264));
  jand g23242(.dina(n40905), .dinb(n40543), .dout(n41265));
  jxor g23243(.dina(n40739), .dinb(n40944), .dout(n41266));
  jand g23244(.dina(n41266), .dinb(n41031), .dout(n41267));
  jor  g23245(.dina(n41267), .dinb(n41265), .dout(n41268));
  jand g23246(.dina(n41268), .dinb(n2547), .dout(n41269));
  jnot g23247(.din(n41269), .dout(n41270));
  jand g23248(.dina(n40905), .dinb(n40549), .dout(n41271));
  jxor g23249(.dina(n40735), .dinb(n40942), .dout(n41272));
  jand g23250(.dina(n41272), .dinb(n41031), .dout(n41273));
  jor  g23251(.dina(n41273), .dinb(n41271), .dout(n41274));
  jand g23252(.dina(n41274), .dinb(n417), .dout(n41275));
  jnot g23253(.din(n41275), .dout(n41276));
  jand g23254(.dina(n40905), .dinb(n40555), .dout(n41277));
  jxor g23255(.dina(n40731), .dinb(n40940), .dout(n41278));
  jand g23256(.dina(n41278), .dinb(n41031), .dout(n41279));
  jor  g23257(.dina(n41279), .dinb(n41277), .dout(n41280));
  jand g23258(.dina(n41280), .dinb(n416), .dout(n41281));
  jnot g23259(.din(n41281), .dout(n41282));
  jand g23260(.dina(n40905), .dinb(n40561), .dout(n41283));
  jxor g23261(.dina(n40727), .dinb(n40938), .dout(n41284));
  jand g23262(.dina(n41284), .dinb(n41031), .dout(n41285));
  jor  g23263(.dina(n41285), .dinb(n41283), .dout(n41286));
  jand g23264(.dina(n41286), .dinb(n422), .dout(n41287));
  jnot g23265(.din(n41287), .dout(n41288));
  jand g23266(.dina(n40905), .dinb(n40567), .dout(n41289));
  jxor g23267(.dina(n40723), .dinb(n40936), .dout(n41290));
  jand g23268(.dina(n41290), .dinb(n41031), .dout(n41291));
  jor  g23269(.dina(n41291), .dinb(n41289), .dout(n41292));
  jand g23270(.dina(n41292), .dinb(n421), .dout(n41293));
  jnot g23271(.din(n41293), .dout(n41294));
  jand g23272(.dina(n40905), .dinb(n40573), .dout(n41295));
  jxor g23273(.dina(n40719), .dinb(n40934), .dout(n41296));
  jand g23274(.dina(n41296), .dinb(n41031), .dout(n41297));
  jor  g23275(.dina(n41297), .dinb(n41295), .dout(n41298));
  jand g23276(.dina(n41298), .dinb(n433), .dout(n41299));
  jnot g23277(.din(n41299), .dout(n41300));
  jand g23278(.dina(n40905), .dinb(n40579), .dout(n41301));
  jxor g23279(.dina(n40715), .dinb(n40932), .dout(n41302));
  jand g23280(.dina(n41302), .dinb(n41031), .dout(n41303));
  jor  g23281(.dina(n41303), .dinb(n41301), .dout(n41304));
  jand g23282(.dina(n41304), .dinb(n432), .dout(n41305));
  jnot g23283(.din(n41305), .dout(n41306));
  jand g23284(.dina(n40905), .dinb(n40585), .dout(n41307));
  jxor g23285(.dina(n40711), .dinb(n40930), .dout(n41308));
  jand g23286(.dina(n41308), .dinb(n41031), .dout(n41309));
  jor  g23287(.dina(n41309), .dinb(n41307), .dout(n41310));
  jand g23288(.dina(n41310), .dinb(n436), .dout(n41311));
  jnot g23289(.din(n41311), .dout(n41312));
  jand g23290(.dina(n40905), .dinb(n40591), .dout(n41313));
  jxor g23291(.dina(n40707), .dinb(n40928), .dout(n41314));
  jand g23292(.dina(n41314), .dinb(n41031), .dout(n41315));
  jor  g23293(.dina(n41315), .dinb(n41313), .dout(n41316));
  jand g23294(.dina(n41316), .dinb(n435), .dout(n41317));
  jnot g23295(.din(n41317), .dout(n41318));
  jand g23296(.dina(n40905), .dinb(n40597), .dout(n41319));
  jxor g23297(.dina(n40703), .dinb(n40926), .dout(n41320));
  jand g23298(.dina(n41320), .dinb(n41031), .dout(n41321));
  jor  g23299(.dina(n41321), .dinb(n41319), .dout(n41322));
  jand g23300(.dina(n41322), .dinb(n440), .dout(n41323));
  jnot g23301(.din(n41323), .dout(n41324));
  jand g23302(.dina(n40905), .dinb(n40603), .dout(n41325));
  jxor g23303(.dina(n40699), .dinb(n40924), .dout(n41326));
  jand g23304(.dina(n41326), .dinb(n41031), .dout(n41327));
  jor  g23305(.dina(n41327), .dinb(n41325), .dout(n41328));
  jand g23306(.dina(n41328), .dinb(n439), .dout(n41329));
  jnot g23307(.din(n41329), .dout(n41330));
  jand g23308(.dina(n40905), .dinb(n40609), .dout(n41331));
  jxor g23309(.dina(n40695), .dinb(n40922), .dout(n41332));
  jand g23310(.dina(n41332), .dinb(n41031), .dout(n41333));
  jor  g23311(.dina(n41333), .dinb(n41331), .dout(n41334));
  jand g23312(.dina(n41334), .dinb(n325), .dout(n41335));
  jnot g23313(.din(n41335), .dout(n41336));
  jand g23314(.dina(n40905), .dinb(n40615), .dout(n41337));
  jxor g23315(.dina(n40691), .dinb(n40920), .dout(n41338));
  jand g23316(.dina(n41338), .dinb(n41031), .dout(n41339));
  jor  g23317(.dina(n41339), .dinb(n41337), .dout(n41340));
  jand g23318(.dina(n41340), .dinb(n324), .dout(n41341));
  jnot g23319(.din(n41341), .dout(n41342));
  jand g23320(.dina(n40905), .dinb(n40621), .dout(n41343));
  jxor g23321(.dina(n40687), .dinb(n40918), .dout(n41344));
  jand g23322(.dina(n41344), .dinb(n41031), .dout(n41345));
  jor  g23323(.dina(n41345), .dinb(n41343), .dout(n41346));
  jand g23324(.dina(n41346), .dinb(n323), .dout(n41347));
  jnot g23325(.din(n41347), .dout(n41348));
  jand g23326(.dina(n40905), .dinb(n40627), .dout(n41349));
  jxor g23327(.dina(n40683), .dinb(n40916), .dout(n41350));
  jand g23328(.dina(n41350), .dinb(n41031), .dout(n41351));
  jor  g23329(.dina(n41351), .dinb(n41349), .dout(n41352));
  jand g23330(.dina(n41352), .dinb(n335), .dout(n41353));
  jnot g23331(.din(n41353), .dout(n41354));
  jand g23332(.dina(n40905), .dinb(n40633), .dout(n41355));
  jxor g23333(.dina(n40679), .dinb(n40914), .dout(n41356));
  jand g23334(.dina(n41356), .dinb(n41031), .dout(n41357));
  jor  g23335(.dina(n41357), .dinb(n41355), .dout(n41358));
  jand g23336(.dina(n41358), .dinb(n334), .dout(n41359));
  jnot g23337(.din(n41359), .dout(n41360));
  jand g23338(.dina(n40905), .dinb(n40639), .dout(n41361));
  jxor g23339(.dina(n40675), .dinb(n40912), .dout(n41362));
  jand g23340(.dina(n41362), .dinb(n41031), .dout(n41363));
  jor  g23341(.dina(n41363), .dinb(n41361), .dout(n41364));
  jand g23342(.dina(n41364), .dinb(n338), .dout(n41365));
  jnot g23343(.din(n41365), .dout(n41366));
  jand g23344(.dina(n40905), .dinb(n40645), .dout(n41367));
  jxor g23345(.dina(n40671), .dinb(n40910), .dout(n41368));
  jand g23346(.dina(n41368), .dinb(n41031), .dout(n41369));
  jor  g23347(.dina(n41369), .dinb(n41367), .dout(n41370));
  jand g23348(.dina(n41370), .dinb(n337), .dout(n41371));
  jnot g23349(.din(n41371), .dout(n41372));
  jand g23350(.dina(n40905), .dinb(n40651), .dout(n41373));
  jxor g23351(.dina(n40667), .dinb(n40908), .dout(n41374));
  jand g23352(.dina(n41374), .dinb(n41031), .dout(n41375));
  jor  g23353(.dina(n41375), .dinb(n41373), .dout(n41376));
  jand g23354(.dina(n41376), .dinb(n344), .dout(n41377));
  jnot g23355(.din(n41377), .dout(n41378));
  jand g23356(.dina(n40905), .dinb(n40658), .dout(n41379));
  jxor g23357(.dina(n40906), .dinb(n16814), .dout(n41380));
  jand g23358(.dina(n41380), .dinb(n41031), .dout(n41381));
  jor  g23359(.dina(n41381), .dinb(n41379), .dout(n41382));
  jand g23360(.dina(n41382), .dinb(n348), .dout(n41383));
  jnot g23361(.din(n41383), .dout(n41384));
  jor  g23362(.dina(n40905), .dinb(n18364), .dout(n41385));
  jand g23363(.dina(n41385), .dinb(a3 ), .dout(n41386));
  jor  g23364(.dina(n40905), .dinb(n16814), .dout(n41387));
  jnot g23365(.din(n41387), .dout(n41388));
  jor  g23366(.dina(n41388), .dinb(n41386), .dout(n41389));
  jand g23367(.dina(n41389), .dinb(n258), .dout(n41390));
  jnot g23368(.din(n41390), .dout(n41391));
  jand g23369(.dina(n41031), .dinb(b0 ), .dout(n41392));
  jor  g23370(.dina(n41392), .dinb(n16812), .dout(n41393));
  jand g23371(.dina(n41387), .dinb(n41393), .dout(n41394));
  jxor g23372(.dina(n41394), .dinb(n258), .dout(n41395));
  jor  g23373(.dina(n41395), .dinb(n17308), .dout(n41396));
  jand g23374(.dina(n41396), .dinb(n41391), .dout(n41397));
  jxor g23375(.dina(n41382), .dinb(n348), .dout(n41398));
  jnot g23376(.din(n41398), .dout(n41399));
  jor  g23377(.dina(n41399), .dinb(n41397), .dout(n41400));
  jand g23378(.dina(n41400), .dinb(n41384), .dout(n41401));
  jxor g23379(.dina(n41376), .dinb(n344), .dout(n41402));
  jnot g23380(.din(n41402), .dout(n41403));
  jor  g23381(.dina(n41403), .dinb(n41401), .dout(n41404));
  jand g23382(.dina(n41404), .dinb(n41378), .dout(n41405));
  jxor g23383(.dina(n41370), .dinb(n337), .dout(n41406));
  jnot g23384(.din(n41406), .dout(n41407));
  jor  g23385(.dina(n41407), .dinb(n41405), .dout(n41408));
  jand g23386(.dina(n41408), .dinb(n41372), .dout(n41409));
  jxor g23387(.dina(n41364), .dinb(n338), .dout(n41410));
  jnot g23388(.din(n41410), .dout(n41411));
  jor  g23389(.dina(n41411), .dinb(n41409), .dout(n41412));
  jand g23390(.dina(n41412), .dinb(n41366), .dout(n41413));
  jxor g23391(.dina(n41358), .dinb(n334), .dout(n41414));
  jnot g23392(.din(n41414), .dout(n41415));
  jor  g23393(.dina(n41415), .dinb(n41413), .dout(n41416));
  jand g23394(.dina(n41416), .dinb(n41360), .dout(n41417));
  jxor g23395(.dina(n41352), .dinb(n335), .dout(n41418));
  jnot g23396(.din(n41418), .dout(n41419));
  jor  g23397(.dina(n41419), .dinb(n41417), .dout(n41420));
  jand g23398(.dina(n41420), .dinb(n41354), .dout(n41421));
  jxor g23399(.dina(n41346), .dinb(n323), .dout(n41422));
  jnot g23400(.din(n41422), .dout(n41423));
  jor  g23401(.dina(n41423), .dinb(n41421), .dout(n41424));
  jand g23402(.dina(n41424), .dinb(n41348), .dout(n41425));
  jxor g23403(.dina(n41340), .dinb(n324), .dout(n41426));
  jnot g23404(.din(n41426), .dout(n41427));
  jor  g23405(.dina(n41427), .dinb(n41425), .dout(n41428));
  jand g23406(.dina(n41428), .dinb(n41342), .dout(n41429));
  jxor g23407(.dina(n41334), .dinb(n325), .dout(n41430));
  jnot g23408(.din(n41430), .dout(n41431));
  jor  g23409(.dina(n41431), .dinb(n41429), .dout(n41432));
  jand g23410(.dina(n41432), .dinb(n41336), .dout(n41433));
  jxor g23411(.dina(n41328), .dinb(n439), .dout(n41434));
  jnot g23412(.din(n41434), .dout(n41435));
  jor  g23413(.dina(n41435), .dinb(n41433), .dout(n41436));
  jand g23414(.dina(n41436), .dinb(n41330), .dout(n41437));
  jxor g23415(.dina(n41322), .dinb(n440), .dout(n41438));
  jnot g23416(.din(n41438), .dout(n41439));
  jor  g23417(.dina(n41439), .dinb(n41437), .dout(n41440));
  jand g23418(.dina(n41440), .dinb(n41324), .dout(n41441));
  jxor g23419(.dina(n41316), .dinb(n435), .dout(n41442));
  jnot g23420(.din(n41442), .dout(n41443));
  jor  g23421(.dina(n41443), .dinb(n41441), .dout(n41444));
  jand g23422(.dina(n41444), .dinb(n41318), .dout(n41445));
  jxor g23423(.dina(n41310), .dinb(n436), .dout(n41446));
  jnot g23424(.din(n41446), .dout(n41447));
  jor  g23425(.dina(n41447), .dinb(n41445), .dout(n41448));
  jand g23426(.dina(n41448), .dinb(n41312), .dout(n41449));
  jxor g23427(.dina(n41304), .dinb(n432), .dout(n41450));
  jnot g23428(.din(n41450), .dout(n41451));
  jor  g23429(.dina(n41451), .dinb(n41449), .dout(n41452));
  jand g23430(.dina(n41452), .dinb(n41306), .dout(n41453));
  jxor g23431(.dina(n41298), .dinb(n433), .dout(n41454));
  jnot g23432(.din(n41454), .dout(n41455));
  jor  g23433(.dina(n41455), .dinb(n41453), .dout(n41456));
  jand g23434(.dina(n41456), .dinb(n41300), .dout(n41457));
  jxor g23435(.dina(n41292), .dinb(n421), .dout(n41458));
  jnot g23436(.din(n41458), .dout(n41459));
  jor  g23437(.dina(n41459), .dinb(n41457), .dout(n41460));
  jand g23438(.dina(n41460), .dinb(n41294), .dout(n41461));
  jxor g23439(.dina(n41286), .dinb(n422), .dout(n41462));
  jnot g23440(.din(n41462), .dout(n41463));
  jor  g23441(.dina(n41463), .dinb(n41461), .dout(n41464));
  jand g23442(.dina(n41464), .dinb(n41288), .dout(n41465));
  jxor g23443(.dina(n41280), .dinb(n416), .dout(n41466));
  jnot g23444(.din(n41466), .dout(n41467));
  jor  g23445(.dina(n41467), .dinb(n41465), .dout(n41468));
  jand g23446(.dina(n41468), .dinb(n41282), .dout(n41469));
  jxor g23447(.dina(n41274), .dinb(n417), .dout(n41470));
  jnot g23448(.din(n41470), .dout(n41471));
  jor  g23449(.dina(n41471), .dinb(n41469), .dout(n41472));
  jand g23450(.dina(n41472), .dinb(n41276), .dout(n41473));
  jxor g23451(.dina(n41268), .dinb(n2547), .dout(n41474));
  jnot g23452(.din(n41474), .dout(n41475));
  jor  g23453(.dina(n41475), .dinb(n41473), .dout(n41476));
  jand g23454(.dina(n41476), .dinb(n41270), .dout(n41477));
  jxor g23455(.dina(n41262), .dinb(n2714), .dout(n41478));
  jnot g23456(.din(n41478), .dout(n41479));
  jor  g23457(.dina(n41479), .dinb(n41477), .dout(n41480));
  jand g23458(.dina(n41480), .dinb(n41264), .dout(n41481));
  jxor g23459(.dina(n41256), .dinb(n405), .dout(n41482));
  jnot g23460(.din(n41482), .dout(n41483));
  jor  g23461(.dina(n41483), .dinb(n41481), .dout(n41484));
  jand g23462(.dina(n41484), .dinb(n41258), .dout(n41485));
  jxor g23463(.dina(n41250), .dinb(n406), .dout(n41486));
  jnot g23464(.din(n41486), .dout(n41487));
  jor  g23465(.dina(n41487), .dinb(n41485), .dout(n41488));
  jand g23466(.dina(n41488), .dinb(n41252), .dout(n41489));
  jxor g23467(.dina(n41244), .dinb(n412), .dout(n41490));
  jnot g23468(.din(n41490), .dout(n41491));
  jor  g23469(.dina(n41491), .dinb(n41489), .dout(n41492));
  jand g23470(.dina(n41492), .dinb(n41246), .dout(n41493));
  jxor g23471(.dina(n41238), .dinb(n413), .dout(n41494));
  jnot g23472(.din(n41494), .dout(n41495));
  jor  g23473(.dina(n41495), .dinb(n41493), .dout(n41496));
  jand g23474(.dina(n41496), .dinb(n41240), .dout(n41497));
  jxor g23475(.dina(n41232), .dinb(n409), .dout(n41498));
  jnot g23476(.din(n41498), .dout(n41499));
  jor  g23477(.dina(n41499), .dinb(n41497), .dout(n41500));
  jand g23478(.dina(n41500), .dinb(n41234), .dout(n41501));
  jxor g23479(.dina(n41226), .dinb(n410), .dout(n41502));
  jnot g23480(.din(n41502), .dout(n41503));
  jor  g23481(.dina(n41503), .dinb(n41501), .dout(n41504));
  jand g23482(.dina(n41504), .dinb(n41228), .dout(n41505));
  jxor g23483(.dina(n41220), .dinb(n426), .dout(n41506));
  jnot g23484(.din(n41506), .dout(n41507));
  jor  g23485(.dina(n41507), .dinb(n41505), .dout(n41508));
  jand g23486(.dina(n41508), .dinb(n41222), .dout(n41509));
  jxor g23487(.dina(n41214), .dinb(n427), .dout(n41510));
  jnot g23488(.din(n41510), .dout(n41511));
  jor  g23489(.dina(n41511), .dinb(n41509), .dout(n41512));
  jand g23490(.dina(n41512), .dinb(n41216), .dout(n41513));
  jxor g23491(.dina(n41208), .dinb(n424), .dout(n41514));
  jnot g23492(.din(n41514), .dout(n41515));
  jor  g23493(.dina(n41515), .dinb(n41513), .dout(n41516));
  jand g23494(.dina(n41516), .dinb(n41210), .dout(n41517));
  jxor g23495(.dina(n41202), .dinb(n300), .dout(n41518));
  jnot g23496(.din(n41518), .dout(n41519));
  jor  g23497(.dina(n41519), .dinb(n41517), .dout(n41520));
  jand g23498(.dina(n41520), .dinb(n41204), .dout(n41521));
  jxor g23499(.dina(n41196), .dinb(n297), .dout(n41522));
  jnot g23500(.din(n41522), .dout(n41523));
  jor  g23501(.dina(n41523), .dinb(n41521), .dout(n41524));
  jand g23502(.dina(n41524), .dinb(n41198), .dout(n41525));
  jxor g23503(.dina(n41190), .dinb(n298), .dout(n41526));
  jnot g23504(.din(n41526), .dout(n41527));
  jor  g23505(.dina(n41527), .dinb(n41525), .dout(n41528));
  jand g23506(.dina(n41528), .dinb(n41192), .dout(n41529));
  jxor g23507(.dina(n41184), .dinb(n301), .dout(n41530));
  jnot g23508(.din(n41530), .dout(n41531));
  jor  g23509(.dina(n41531), .dinb(n41529), .dout(n41532));
  jand g23510(.dina(n41532), .dinb(n41186), .dout(n41533));
  jxor g23511(.dina(n41178), .dinb(n293), .dout(n41534));
  jnot g23512(.din(n41534), .dout(n41535));
  jor  g23513(.dina(n41535), .dinb(n41533), .dout(n41536));
  jand g23514(.dina(n41536), .dinb(n41180), .dout(n41537));
  jxor g23515(.dina(n41172), .dinb(n294), .dout(n41538));
  jnot g23516(.din(n41538), .dout(n41539));
  jor  g23517(.dina(n41539), .dinb(n41537), .dout(n41540));
  jand g23518(.dina(n41540), .dinb(n41174), .dout(n41541));
  jxor g23519(.dina(n41166), .dinb(n290), .dout(n41542));
  jnot g23520(.din(n41542), .dout(n41543));
  jor  g23521(.dina(n41543), .dinb(n41541), .dout(n41544));
  jand g23522(.dina(n41544), .dinb(n41168), .dout(n41545));
  jxor g23523(.dina(n41160), .dinb(n291), .dout(n41546));
  jnot g23524(.din(n41546), .dout(n41547));
  jor  g23525(.dina(n41547), .dinb(n41545), .dout(n41548));
  jand g23526(.dina(n41548), .dinb(n41162), .dout(n41549));
  jxor g23527(.dina(n41154), .dinb(n284), .dout(n41550));
  jnot g23528(.din(n41550), .dout(n41551));
  jor  g23529(.dina(n41551), .dinb(n41549), .dout(n41552));
  jand g23530(.dina(n41552), .dinb(n41156), .dout(n41553));
  jxor g23531(.dina(n41148), .dinb(n285), .dout(n41554));
  jnot g23532(.din(n41554), .dout(n41555));
  jor  g23533(.dina(n41555), .dinb(n41553), .dout(n41556));
  jand g23534(.dina(n41556), .dinb(n41150), .dout(n41557));
  jxor g23535(.dina(n41142), .dinb(n281), .dout(n41558));
  jnot g23536(.din(n41558), .dout(n41559));
  jor  g23537(.dina(n41559), .dinb(n41557), .dout(n41560));
  jand g23538(.dina(n41560), .dinb(n41144), .dout(n41561));
  jxor g23539(.dina(n41136), .dinb(n282), .dout(n41562));
  jnot g23540(.din(n41562), .dout(n41563));
  jor  g23541(.dina(n41563), .dinb(n41561), .dout(n41564));
  jand g23542(.dina(n41564), .dinb(n41138), .dout(n41565));
  jxor g23543(.dina(n41130), .dinb(n397), .dout(n41566));
  jnot g23544(.din(n41566), .dout(n41567));
  jor  g23545(.dina(n41567), .dinb(n41565), .dout(n41568));
  jand g23546(.dina(n41568), .dinb(n41132), .dout(n41569));
  jxor g23547(.dina(n41124), .dinb(n513), .dout(n41570));
  jnot g23548(.din(n41570), .dout(n41571));
  jor  g23549(.dina(n41571), .dinb(n41569), .dout(n41572));
  jand g23550(.dina(n41572), .dinb(n41126), .dout(n41573));
  jxor g23551(.dina(n41118), .dinb(n514), .dout(n41574));
  jnot g23552(.din(n41574), .dout(n41575));
  jor  g23553(.dina(n41575), .dinb(n41573), .dout(n41576));
  jand g23554(.dina(n41576), .dinb(n41120), .dout(n41577));
  jxor g23555(.dina(n41112), .dinb(n510), .dout(n41578));
  jnot g23556(.din(n41578), .dout(n41579));
  jor  g23557(.dina(n41579), .dinb(n41577), .dout(n41580));
  jand g23558(.dina(n41580), .dinb(n41114), .dout(n41581));
  jxor g23559(.dina(n41106), .dinb(n396), .dout(n41582));
  jnot g23560(.din(n41582), .dout(n41583));
  jor  g23561(.dina(n41583), .dinb(n41581), .dout(n41584));
  jand g23562(.dina(n41584), .dinb(n41108), .dout(n41585));
  jxor g23563(.dina(n41100), .dinb(n383), .dout(n41586));
  jnot g23564(.din(n41586), .dout(n41587));
  jor  g23565(.dina(n41587), .dinb(n41585), .dout(n41588));
  jand g23566(.dina(n41588), .dinb(n41102), .dout(n41589));
  jxor g23567(.dina(n41094), .dinb(n12211), .dout(n41590));
  jnot g23568(.din(n41590), .dout(n41591));
  jor  g23569(.dina(n41591), .dinb(n41589), .dout(n41592));
  jand g23570(.dina(n41592), .dinb(n41096), .dout(n41593));
  jxor g23571(.dina(n41088), .dinb(n12214), .dout(n41594));
  jnot g23572(.din(n41594), .dout(n41595));
  jor  g23573(.dina(n41595), .dinb(n41593), .dout(n41596));
  jand g23574(.dina(n41596), .dinb(n41090), .dout(n41597));
  jxor g23575(.dina(n41082), .dinb(n384), .dout(n41598));
  jnot g23576(.din(n41598), .dout(n41599));
  jor  g23577(.dina(n41599), .dinb(n41597), .dout(n41600));
  jand g23578(.dina(n41600), .dinb(n41084), .dout(n41601));
  jxor g23579(.dina(n41076), .dinb(n374), .dout(n41602));
  jnot g23580(.din(n41602), .dout(n41603));
  jor  g23581(.dina(n41603), .dinb(n41601), .dout(n41604));
  jand g23582(.dina(n41604), .dinb(n41078), .dout(n41605));
  jxor g23583(.dina(n41070), .dinb(n376), .dout(n41606));
  jnot g23584(.din(n41606), .dout(n41607));
  jor  g23585(.dina(n41607), .dinb(n41605), .dout(n41608));
  jand g23586(.dina(n41608), .dinb(n41072), .dout(n41609));
  jxor g23587(.dina(n41064), .dinb(n377), .dout(n41610));
  jnot g23588(.din(n41610), .dout(n41611));
  jor  g23589(.dina(n41611), .dinb(n41609), .dout(n41612));
  jand g23590(.dina(n41612), .dinb(n41066), .dout(n41613));
  jxor g23591(.dina(n41058), .dinb(n375), .dout(n41614));
  jnot g23592(.din(n41614), .dout(n41615));
  jor  g23593(.dina(n41615), .dinb(n41613), .dout(n41616));
  jand g23594(.dina(n41616), .dinb(n41060), .dout(n41617));
  jxor g23595(.dina(n41052), .dinb(n362), .dout(n41618));
  jnot g23596(.din(n41618), .dout(n41619));
  jor  g23597(.dina(n41619), .dinb(n41617), .dout(n41620));
  jand g23598(.dina(n41620), .dinb(n41054), .dout(n41621));
  jxor g23599(.dina(n41046), .dinb(n363), .dout(n41622));
  jnot g23600(.din(n41622), .dout(n41623));
  jor  g23601(.dina(n41623), .dinb(n41621), .dout(n41624));
  jand g23602(.dina(n41624), .dinb(n41048), .dout(n41625));
  jxor g23603(.dina(n41040), .dinb(n365), .dout(n41626));
  jnot g23604(.din(n41626), .dout(n41627));
  jor  g23605(.dina(n41627), .dinb(n41625), .dout(n41628));
  jand g23606(.dina(n41628), .dinb(n41042), .dout(n41629));
  jxor g23607(.dina(n41034), .dinb(n366), .dout(n41630));
  jnot g23608(.din(n41630), .dout(n41631));
  jor  g23609(.dina(n41631), .dinb(n41629), .dout(n41632));
  jand g23610(.dina(n41632), .dinb(n41036), .dout(n41633));
  jand g23611(.dina(n41027), .dinb(n256), .dout(n41634));
  jnot g23612(.din(n41634), .dout(n41635));
  jand g23613(.dina(n41635), .dinb(n41633), .dout(n41636));
  jnot g23614(.din(n41027), .dout(n41637));
  jand g23615(.dina(n41637), .dinb(b61 ), .dout(n41638));
  jor  g23616(.dina(n41638), .dinb(n262), .dout(n41639));
  jor  g23617(.dina(n41639), .dinb(n41636), .dout(n41640));
  jxor g23618(.dina(n41394), .dinb(b1 ), .dout(n41641));
  jand g23619(.dina(n41641), .dinb(n17309), .dout(n41642));
  jor  g23620(.dina(n41642), .dinb(n41390), .dout(n41643));
  jand g23621(.dina(n41398), .dinb(n41643), .dout(n41644));
  jor  g23622(.dina(n41644), .dinb(n41383), .dout(n41645));
  jand g23623(.dina(n41402), .dinb(n41645), .dout(n41646));
  jor  g23624(.dina(n41646), .dinb(n41377), .dout(n41647));
  jand g23625(.dina(n41406), .dinb(n41647), .dout(n41648));
  jor  g23626(.dina(n41648), .dinb(n41371), .dout(n41649));
  jand g23627(.dina(n41410), .dinb(n41649), .dout(n41650));
  jor  g23628(.dina(n41650), .dinb(n41365), .dout(n41651));
  jand g23629(.dina(n41414), .dinb(n41651), .dout(n41652));
  jor  g23630(.dina(n41652), .dinb(n41359), .dout(n41653));
  jand g23631(.dina(n41418), .dinb(n41653), .dout(n41654));
  jor  g23632(.dina(n41654), .dinb(n41353), .dout(n41655));
  jand g23633(.dina(n41422), .dinb(n41655), .dout(n41656));
  jor  g23634(.dina(n41656), .dinb(n41347), .dout(n41657));
  jand g23635(.dina(n41426), .dinb(n41657), .dout(n41658));
  jor  g23636(.dina(n41658), .dinb(n41341), .dout(n41659));
  jand g23637(.dina(n41430), .dinb(n41659), .dout(n41660));
  jor  g23638(.dina(n41660), .dinb(n41335), .dout(n41661));
  jand g23639(.dina(n41434), .dinb(n41661), .dout(n41662));
  jor  g23640(.dina(n41662), .dinb(n41329), .dout(n41663));
  jand g23641(.dina(n41438), .dinb(n41663), .dout(n41664));
  jor  g23642(.dina(n41664), .dinb(n41323), .dout(n41665));
  jand g23643(.dina(n41442), .dinb(n41665), .dout(n41666));
  jor  g23644(.dina(n41666), .dinb(n41317), .dout(n41667));
  jand g23645(.dina(n41446), .dinb(n41667), .dout(n41668));
  jor  g23646(.dina(n41668), .dinb(n41311), .dout(n41669));
  jand g23647(.dina(n41450), .dinb(n41669), .dout(n41670));
  jor  g23648(.dina(n41670), .dinb(n41305), .dout(n41671));
  jand g23649(.dina(n41454), .dinb(n41671), .dout(n41672));
  jor  g23650(.dina(n41672), .dinb(n41299), .dout(n41673));
  jand g23651(.dina(n41458), .dinb(n41673), .dout(n41674));
  jor  g23652(.dina(n41674), .dinb(n41293), .dout(n41675));
  jand g23653(.dina(n41462), .dinb(n41675), .dout(n41676));
  jor  g23654(.dina(n41676), .dinb(n41287), .dout(n41677));
  jand g23655(.dina(n41466), .dinb(n41677), .dout(n41678));
  jor  g23656(.dina(n41678), .dinb(n41281), .dout(n41679));
  jand g23657(.dina(n41470), .dinb(n41679), .dout(n41680));
  jor  g23658(.dina(n41680), .dinb(n41275), .dout(n41681));
  jand g23659(.dina(n41474), .dinb(n41681), .dout(n41682));
  jor  g23660(.dina(n41682), .dinb(n41269), .dout(n41683));
  jand g23661(.dina(n41478), .dinb(n41683), .dout(n41684));
  jor  g23662(.dina(n41684), .dinb(n41263), .dout(n41685));
  jand g23663(.dina(n41482), .dinb(n41685), .dout(n41686));
  jor  g23664(.dina(n41686), .dinb(n41257), .dout(n41687));
  jand g23665(.dina(n41486), .dinb(n41687), .dout(n41688));
  jor  g23666(.dina(n41688), .dinb(n41251), .dout(n41689));
  jand g23667(.dina(n41490), .dinb(n41689), .dout(n41690));
  jor  g23668(.dina(n41690), .dinb(n41245), .dout(n41691));
  jand g23669(.dina(n41494), .dinb(n41691), .dout(n41692));
  jor  g23670(.dina(n41692), .dinb(n41239), .dout(n41693));
  jand g23671(.dina(n41498), .dinb(n41693), .dout(n41694));
  jor  g23672(.dina(n41694), .dinb(n41233), .dout(n41695));
  jand g23673(.dina(n41502), .dinb(n41695), .dout(n41696));
  jor  g23674(.dina(n41696), .dinb(n41227), .dout(n41697));
  jand g23675(.dina(n41506), .dinb(n41697), .dout(n41698));
  jor  g23676(.dina(n41698), .dinb(n41221), .dout(n41699));
  jand g23677(.dina(n41510), .dinb(n41699), .dout(n41700));
  jor  g23678(.dina(n41700), .dinb(n41215), .dout(n41701));
  jand g23679(.dina(n41514), .dinb(n41701), .dout(n41702));
  jor  g23680(.dina(n41702), .dinb(n41209), .dout(n41703));
  jand g23681(.dina(n41518), .dinb(n41703), .dout(n41704));
  jor  g23682(.dina(n41704), .dinb(n41203), .dout(n41705));
  jand g23683(.dina(n41522), .dinb(n41705), .dout(n41706));
  jor  g23684(.dina(n41706), .dinb(n41197), .dout(n41707));
  jand g23685(.dina(n41526), .dinb(n41707), .dout(n41708));
  jor  g23686(.dina(n41708), .dinb(n41191), .dout(n41709));
  jand g23687(.dina(n41530), .dinb(n41709), .dout(n41710));
  jor  g23688(.dina(n41710), .dinb(n41185), .dout(n41711));
  jand g23689(.dina(n41534), .dinb(n41711), .dout(n41712));
  jor  g23690(.dina(n41712), .dinb(n41179), .dout(n41713));
  jand g23691(.dina(n41538), .dinb(n41713), .dout(n41714));
  jor  g23692(.dina(n41714), .dinb(n41173), .dout(n41715));
  jand g23693(.dina(n41542), .dinb(n41715), .dout(n41716));
  jor  g23694(.dina(n41716), .dinb(n41167), .dout(n41717));
  jand g23695(.dina(n41546), .dinb(n41717), .dout(n41718));
  jor  g23696(.dina(n41718), .dinb(n41161), .dout(n41719));
  jand g23697(.dina(n41550), .dinb(n41719), .dout(n41720));
  jor  g23698(.dina(n41720), .dinb(n41155), .dout(n41721));
  jand g23699(.dina(n41554), .dinb(n41721), .dout(n41722));
  jor  g23700(.dina(n41722), .dinb(n41149), .dout(n41723));
  jand g23701(.dina(n41558), .dinb(n41723), .dout(n41724));
  jor  g23702(.dina(n41724), .dinb(n41143), .dout(n41725));
  jand g23703(.dina(n41562), .dinb(n41725), .dout(n41726));
  jor  g23704(.dina(n41726), .dinb(n41137), .dout(n41727));
  jand g23705(.dina(n41566), .dinb(n41727), .dout(n41728));
  jor  g23706(.dina(n41728), .dinb(n41131), .dout(n41729));
  jand g23707(.dina(n41570), .dinb(n41729), .dout(n41730));
  jor  g23708(.dina(n41730), .dinb(n41125), .dout(n41731));
  jand g23709(.dina(n41574), .dinb(n41731), .dout(n41732));
  jor  g23710(.dina(n41732), .dinb(n41119), .dout(n41733));
  jand g23711(.dina(n41578), .dinb(n41733), .dout(n41734));
  jor  g23712(.dina(n41734), .dinb(n41113), .dout(n41735));
  jand g23713(.dina(n41582), .dinb(n41735), .dout(n41736));
  jor  g23714(.dina(n41736), .dinb(n41107), .dout(n41737));
  jand g23715(.dina(n41586), .dinb(n41737), .dout(n41738));
  jor  g23716(.dina(n41738), .dinb(n41101), .dout(n41739));
  jand g23717(.dina(n41590), .dinb(n41739), .dout(n41740));
  jor  g23718(.dina(n41740), .dinb(n41095), .dout(n41741));
  jand g23719(.dina(n41594), .dinb(n41741), .dout(n41742));
  jor  g23720(.dina(n41742), .dinb(n41089), .dout(n41743));
  jand g23721(.dina(n41598), .dinb(n41743), .dout(n41744));
  jor  g23722(.dina(n41744), .dinb(n41083), .dout(n41745));
  jand g23723(.dina(n41602), .dinb(n41745), .dout(n41746));
  jor  g23724(.dina(n41746), .dinb(n41077), .dout(n41747));
  jand g23725(.dina(n41606), .dinb(n41747), .dout(n41748));
  jor  g23726(.dina(n41748), .dinb(n41071), .dout(n41749));
  jand g23727(.dina(n41610), .dinb(n41749), .dout(n41750));
  jor  g23728(.dina(n41750), .dinb(n41065), .dout(n41751));
  jand g23729(.dina(n41614), .dinb(n41751), .dout(n41752));
  jor  g23730(.dina(n41752), .dinb(n41059), .dout(n41753));
  jand g23731(.dina(n41618), .dinb(n41753), .dout(n41754));
  jor  g23732(.dina(n41754), .dinb(n41053), .dout(n41755));
  jand g23733(.dina(n41622), .dinb(n41755), .dout(n41756));
  jor  g23734(.dina(n41756), .dinb(n41047), .dout(n41757));
  jand g23735(.dina(n41626), .dinb(n41757), .dout(n41758));
  jor  g23736(.dina(n41758), .dinb(n41041), .dout(n41759));
  jand g23737(.dina(n41630), .dinb(n41759), .dout(n41760));
  jor  g23738(.dina(n41760), .dinb(n41035), .dout(n41761));
  jand g23739(.dina(n41761), .dinb(n370), .dout(n41762));
  jor  g23740(.dina(n41762), .dinb(n41640), .dout(n41763));
  jand g23741(.dina(n41763), .dinb(n41027), .dout(n41764));
  jnot g23742(.din(n41764), .dout(n41765));
  jand g23743(.dina(n41765), .dinb(b63 ), .dout(n41766));
  jand g23744(.dina(n41640), .dinb(n41034), .dout(n41767));
  jor  g23745(.dina(n41634), .dinb(n41761), .dout(n41768));
  jnot g23746(.din(n41639), .dout(n41769));
  jand g23747(.dina(n41769), .dinb(n41768), .dout(n41770));
  jxor g23748(.dina(n41630), .dinb(n41759), .dout(n41771));
  jand g23749(.dina(n41771), .dinb(n41770), .dout(n41772));
  jor  g23750(.dina(n41772), .dinb(n41767), .dout(n41773));
  jand g23751(.dina(n41773), .dinb(n256), .dout(n41774));
  jnot g23752(.din(n41774), .dout(n41775));
  jand g23753(.dina(n41640), .dinb(n41040), .dout(n41776));
  jxor g23754(.dina(n41626), .dinb(n41757), .dout(n41777));
  jand g23755(.dina(n41777), .dinb(n41770), .dout(n41778));
  jor  g23756(.dina(n41778), .dinb(n41776), .dout(n41779));
  jand g23757(.dina(n41779), .dinb(n366), .dout(n41780));
  jnot g23758(.din(n41780), .dout(n41781));
  jand g23759(.dina(n41640), .dinb(n41046), .dout(n41782));
  jxor g23760(.dina(n41622), .dinb(n41755), .dout(n41783));
  jand g23761(.dina(n41783), .dinb(n41770), .dout(n41784));
  jor  g23762(.dina(n41784), .dinb(n41782), .dout(n41785));
  jand g23763(.dina(n41785), .dinb(n365), .dout(n41786));
  jnot g23764(.din(n41786), .dout(n41787));
  jand g23765(.dina(n41640), .dinb(n41052), .dout(n41788));
  jxor g23766(.dina(n41618), .dinb(n41753), .dout(n41789));
  jand g23767(.dina(n41789), .dinb(n41770), .dout(n41790));
  jor  g23768(.dina(n41790), .dinb(n41788), .dout(n41791));
  jand g23769(.dina(n41791), .dinb(n363), .dout(n41792));
  jnot g23770(.din(n41792), .dout(n41793));
  jand g23771(.dina(n41640), .dinb(n41058), .dout(n41794));
  jxor g23772(.dina(n41614), .dinb(n41751), .dout(n41795));
  jand g23773(.dina(n41795), .dinb(n41770), .dout(n41796));
  jor  g23774(.dina(n41796), .dinb(n41794), .dout(n41797));
  jand g23775(.dina(n41797), .dinb(n362), .dout(n41798));
  jnot g23776(.din(n41798), .dout(n41799));
  jand g23777(.dina(n41640), .dinb(n41064), .dout(n41800));
  jxor g23778(.dina(n41610), .dinb(n41749), .dout(n41801));
  jand g23779(.dina(n41801), .dinb(n41770), .dout(n41802));
  jor  g23780(.dina(n41802), .dinb(n41800), .dout(n41803));
  jand g23781(.dina(n41803), .dinb(n375), .dout(n41804));
  jnot g23782(.din(n41804), .dout(n41805));
  jand g23783(.dina(n41640), .dinb(n41070), .dout(n41806));
  jxor g23784(.dina(n41606), .dinb(n41747), .dout(n41807));
  jand g23785(.dina(n41807), .dinb(n41770), .dout(n41808));
  jor  g23786(.dina(n41808), .dinb(n41806), .dout(n41809));
  jand g23787(.dina(n41809), .dinb(n377), .dout(n41810));
  jnot g23788(.din(n41810), .dout(n41811));
  jand g23789(.dina(n41640), .dinb(n41076), .dout(n41812));
  jxor g23790(.dina(n41602), .dinb(n41745), .dout(n41813));
  jand g23791(.dina(n41813), .dinb(n41770), .dout(n41814));
  jor  g23792(.dina(n41814), .dinb(n41812), .dout(n41815));
  jand g23793(.dina(n41815), .dinb(n376), .dout(n41816));
  jnot g23794(.din(n41816), .dout(n41817));
  jand g23795(.dina(n41640), .dinb(n41082), .dout(n41818));
  jxor g23796(.dina(n41598), .dinb(n41743), .dout(n41819));
  jand g23797(.dina(n41819), .dinb(n41770), .dout(n41820));
  jor  g23798(.dina(n41820), .dinb(n41818), .dout(n41821));
  jand g23799(.dina(n41821), .dinb(n374), .dout(n41822));
  jnot g23800(.din(n41822), .dout(n41823));
  jand g23801(.dina(n41640), .dinb(n41088), .dout(n41824));
  jxor g23802(.dina(n41594), .dinb(n41741), .dout(n41825));
  jand g23803(.dina(n41825), .dinb(n41770), .dout(n41826));
  jor  g23804(.dina(n41826), .dinb(n41824), .dout(n41827));
  jand g23805(.dina(n41827), .dinb(n384), .dout(n41828));
  jnot g23806(.din(n41828), .dout(n41829));
  jand g23807(.dina(n41640), .dinb(n41094), .dout(n41830));
  jxor g23808(.dina(n41590), .dinb(n41739), .dout(n41831));
  jand g23809(.dina(n41831), .dinb(n41770), .dout(n41832));
  jor  g23810(.dina(n41832), .dinb(n41830), .dout(n41833));
  jand g23811(.dina(n41833), .dinb(n12214), .dout(n41834));
  jnot g23812(.din(n41834), .dout(n41835));
  jand g23813(.dina(n41640), .dinb(n41100), .dout(n41836));
  jxor g23814(.dina(n41586), .dinb(n41737), .dout(n41837));
  jand g23815(.dina(n41837), .dinb(n41770), .dout(n41838));
  jor  g23816(.dina(n41838), .dinb(n41836), .dout(n41839));
  jand g23817(.dina(n41839), .dinb(n12211), .dout(n41840));
  jnot g23818(.din(n41840), .dout(n41841));
  jand g23819(.dina(n41640), .dinb(n41106), .dout(n41842));
  jxor g23820(.dina(n41582), .dinb(n41735), .dout(n41843));
  jand g23821(.dina(n41843), .dinb(n41770), .dout(n41844));
  jor  g23822(.dina(n41844), .dinb(n41842), .dout(n41845));
  jand g23823(.dina(n41845), .dinb(n383), .dout(n41846));
  jnot g23824(.din(n41846), .dout(n41847));
  jand g23825(.dina(n41640), .dinb(n41112), .dout(n41848));
  jxor g23826(.dina(n41578), .dinb(n41733), .dout(n41849));
  jand g23827(.dina(n41849), .dinb(n41770), .dout(n41850));
  jor  g23828(.dina(n41850), .dinb(n41848), .dout(n41851));
  jand g23829(.dina(n41851), .dinb(n396), .dout(n41852));
  jnot g23830(.din(n41852), .dout(n41853));
  jand g23831(.dina(n41640), .dinb(n41118), .dout(n41854));
  jxor g23832(.dina(n41574), .dinb(n41731), .dout(n41855));
  jand g23833(.dina(n41855), .dinb(n41770), .dout(n41856));
  jor  g23834(.dina(n41856), .dinb(n41854), .dout(n41857));
  jand g23835(.dina(n41857), .dinb(n510), .dout(n41858));
  jnot g23836(.din(n41858), .dout(n41859));
  jand g23837(.dina(n41640), .dinb(n41124), .dout(n41860));
  jxor g23838(.dina(n41570), .dinb(n41729), .dout(n41861));
  jand g23839(.dina(n41861), .dinb(n41770), .dout(n41862));
  jor  g23840(.dina(n41862), .dinb(n41860), .dout(n41863));
  jand g23841(.dina(n41863), .dinb(n514), .dout(n41864));
  jnot g23842(.din(n41864), .dout(n41865));
  jand g23843(.dina(n41640), .dinb(n41130), .dout(n41866));
  jxor g23844(.dina(n41566), .dinb(n41727), .dout(n41867));
  jand g23845(.dina(n41867), .dinb(n41770), .dout(n41868));
  jor  g23846(.dina(n41868), .dinb(n41866), .dout(n41869));
  jand g23847(.dina(n41869), .dinb(n513), .dout(n41870));
  jnot g23848(.din(n41870), .dout(n41871));
  jand g23849(.dina(n41640), .dinb(n41136), .dout(n41872));
  jxor g23850(.dina(n41562), .dinb(n41725), .dout(n41873));
  jand g23851(.dina(n41873), .dinb(n41770), .dout(n41874));
  jor  g23852(.dina(n41874), .dinb(n41872), .dout(n41875));
  jand g23853(.dina(n41875), .dinb(n397), .dout(n41876));
  jnot g23854(.din(n41876), .dout(n41877));
  jand g23855(.dina(n41640), .dinb(n41142), .dout(n41878));
  jxor g23856(.dina(n41558), .dinb(n41723), .dout(n41879));
  jand g23857(.dina(n41879), .dinb(n41770), .dout(n41880));
  jor  g23858(.dina(n41880), .dinb(n41878), .dout(n41881));
  jand g23859(.dina(n41881), .dinb(n282), .dout(n41882));
  jnot g23860(.din(n41882), .dout(n41883));
  jand g23861(.dina(n41640), .dinb(n41148), .dout(n41884));
  jxor g23862(.dina(n41554), .dinb(n41721), .dout(n41885));
  jand g23863(.dina(n41885), .dinb(n41770), .dout(n41886));
  jor  g23864(.dina(n41886), .dinb(n41884), .dout(n41887));
  jand g23865(.dina(n41887), .dinb(n281), .dout(n41888));
  jnot g23866(.din(n41888), .dout(n41889));
  jand g23867(.dina(n41640), .dinb(n41154), .dout(n41890));
  jxor g23868(.dina(n41550), .dinb(n41719), .dout(n41891));
  jand g23869(.dina(n41891), .dinb(n41770), .dout(n41892));
  jor  g23870(.dina(n41892), .dinb(n41890), .dout(n41893));
  jand g23871(.dina(n41893), .dinb(n285), .dout(n41894));
  jnot g23872(.din(n41894), .dout(n41895));
  jand g23873(.dina(n41640), .dinb(n41160), .dout(n41896));
  jxor g23874(.dina(n41546), .dinb(n41717), .dout(n41897));
  jand g23875(.dina(n41897), .dinb(n41770), .dout(n41898));
  jor  g23876(.dina(n41898), .dinb(n41896), .dout(n41899));
  jand g23877(.dina(n41899), .dinb(n284), .dout(n41900));
  jnot g23878(.din(n41900), .dout(n41901));
  jand g23879(.dina(n41640), .dinb(n41166), .dout(n41902));
  jxor g23880(.dina(n41542), .dinb(n41715), .dout(n41903));
  jand g23881(.dina(n41903), .dinb(n41770), .dout(n41904));
  jor  g23882(.dina(n41904), .dinb(n41902), .dout(n41905));
  jand g23883(.dina(n41905), .dinb(n291), .dout(n41906));
  jnot g23884(.din(n41906), .dout(n41907));
  jand g23885(.dina(n41640), .dinb(n41172), .dout(n41908));
  jxor g23886(.dina(n41538), .dinb(n41713), .dout(n41909));
  jand g23887(.dina(n41909), .dinb(n41770), .dout(n41910));
  jor  g23888(.dina(n41910), .dinb(n41908), .dout(n41911));
  jand g23889(.dina(n41911), .dinb(n290), .dout(n41912));
  jnot g23890(.din(n41912), .dout(n41913));
  jand g23891(.dina(n41640), .dinb(n41178), .dout(n41914));
  jxor g23892(.dina(n41534), .dinb(n41711), .dout(n41915));
  jand g23893(.dina(n41915), .dinb(n41770), .dout(n41916));
  jor  g23894(.dina(n41916), .dinb(n41914), .dout(n41917));
  jand g23895(.dina(n41917), .dinb(n294), .dout(n41918));
  jnot g23896(.din(n41918), .dout(n41919));
  jand g23897(.dina(n41640), .dinb(n41184), .dout(n41920));
  jxor g23898(.dina(n41530), .dinb(n41709), .dout(n41921));
  jand g23899(.dina(n41921), .dinb(n41770), .dout(n41922));
  jor  g23900(.dina(n41922), .dinb(n41920), .dout(n41923));
  jand g23901(.dina(n41923), .dinb(n293), .dout(n41924));
  jnot g23902(.din(n41924), .dout(n41925));
  jand g23903(.dina(n41640), .dinb(n41190), .dout(n41926));
  jxor g23904(.dina(n41526), .dinb(n41707), .dout(n41927));
  jand g23905(.dina(n41927), .dinb(n41770), .dout(n41928));
  jor  g23906(.dina(n41928), .dinb(n41926), .dout(n41929));
  jand g23907(.dina(n41929), .dinb(n301), .dout(n41930));
  jnot g23908(.din(n41930), .dout(n41931));
  jand g23909(.dina(n41640), .dinb(n41196), .dout(n41932));
  jxor g23910(.dina(n41522), .dinb(n41705), .dout(n41933));
  jand g23911(.dina(n41933), .dinb(n41770), .dout(n41934));
  jor  g23912(.dina(n41934), .dinb(n41932), .dout(n41935));
  jand g23913(.dina(n41935), .dinb(n298), .dout(n41936));
  jnot g23914(.din(n41936), .dout(n41937));
  jand g23915(.dina(n41640), .dinb(n41202), .dout(n41938));
  jxor g23916(.dina(n41518), .dinb(n41703), .dout(n41939));
  jand g23917(.dina(n41939), .dinb(n41770), .dout(n41940));
  jor  g23918(.dina(n41940), .dinb(n41938), .dout(n41941));
  jand g23919(.dina(n41941), .dinb(n297), .dout(n41942));
  jnot g23920(.din(n41942), .dout(n41943));
  jand g23921(.dina(n41640), .dinb(n41208), .dout(n41944));
  jxor g23922(.dina(n41514), .dinb(n41701), .dout(n41945));
  jand g23923(.dina(n41945), .dinb(n41770), .dout(n41946));
  jor  g23924(.dina(n41946), .dinb(n41944), .dout(n41947));
  jand g23925(.dina(n41947), .dinb(n300), .dout(n41948));
  jnot g23926(.din(n41948), .dout(n41949));
  jand g23927(.dina(n41640), .dinb(n41214), .dout(n41950));
  jxor g23928(.dina(n41510), .dinb(n41699), .dout(n41951));
  jand g23929(.dina(n41951), .dinb(n41770), .dout(n41952));
  jor  g23930(.dina(n41952), .dinb(n41950), .dout(n41953));
  jand g23931(.dina(n41953), .dinb(n424), .dout(n41954));
  jnot g23932(.din(n41954), .dout(n41955));
  jand g23933(.dina(n41640), .dinb(n41220), .dout(n41956));
  jxor g23934(.dina(n41506), .dinb(n41697), .dout(n41957));
  jand g23935(.dina(n41957), .dinb(n41770), .dout(n41958));
  jor  g23936(.dina(n41958), .dinb(n41956), .dout(n41959));
  jand g23937(.dina(n41959), .dinb(n427), .dout(n41960));
  jnot g23938(.din(n41960), .dout(n41961));
  jand g23939(.dina(n41640), .dinb(n41226), .dout(n41962));
  jxor g23940(.dina(n41502), .dinb(n41695), .dout(n41963));
  jand g23941(.dina(n41963), .dinb(n41770), .dout(n41964));
  jor  g23942(.dina(n41964), .dinb(n41962), .dout(n41965));
  jand g23943(.dina(n41965), .dinb(n426), .dout(n41966));
  jnot g23944(.din(n41966), .dout(n41967));
  jand g23945(.dina(n41640), .dinb(n41232), .dout(n41968));
  jxor g23946(.dina(n41498), .dinb(n41693), .dout(n41969));
  jand g23947(.dina(n41969), .dinb(n41770), .dout(n41970));
  jor  g23948(.dina(n41970), .dinb(n41968), .dout(n41971));
  jand g23949(.dina(n41971), .dinb(n410), .dout(n41972));
  jnot g23950(.din(n41972), .dout(n41973));
  jand g23951(.dina(n41640), .dinb(n41238), .dout(n41974));
  jxor g23952(.dina(n41494), .dinb(n41691), .dout(n41975));
  jand g23953(.dina(n41975), .dinb(n41770), .dout(n41976));
  jor  g23954(.dina(n41976), .dinb(n41974), .dout(n41977));
  jand g23955(.dina(n41977), .dinb(n409), .dout(n41978));
  jnot g23956(.din(n41978), .dout(n41979));
  jand g23957(.dina(n41640), .dinb(n41244), .dout(n41980));
  jxor g23958(.dina(n41490), .dinb(n41689), .dout(n41981));
  jand g23959(.dina(n41981), .dinb(n41770), .dout(n41982));
  jor  g23960(.dina(n41982), .dinb(n41980), .dout(n41983));
  jand g23961(.dina(n41983), .dinb(n413), .dout(n41984));
  jnot g23962(.din(n41984), .dout(n41985));
  jand g23963(.dina(n41640), .dinb(n41250), .dout(n41986));
  jxor g23964(.dina(n41486), .dinb(n41687), .dout(n41987));
  jand g23965(.dina(n41987), .dinb(n41770), .dout(n41988));
  jor  g23966(.dina(n41988), .dinb(n41986), .dout(n41989));
  jand g23967(.dina(n41989), .dinb(n412), .dout(n41990));
  jnot g23968(.din(n41990), .dout(n41991));
  jand g23969(.dina(n41640), .dinb(n41256), .dout(n41992));
  jxor g23970(.dina(n41482), .dinb(n41685), .dout(n41993));
  jand g23971(.dina(n41993), .dinb(n41770), .dout(n41994));
  jor  g23972(.dina(n41994), .dinb(n41992), .dout(n41995));
  jand g23973(.dina(n41995), .dinb(n406), .dout(n41996));
  jnot g23974(.din(n41996), .dout(n41997));
  jand g23975(.dina(n41640), .dinb(n41262), .dout(n41998));
  jxor g23976(.dina(n41478), .dinb(n41683), .dout(n41999));
  jand g23977(.dina(n41999), .dinb(n41770), .dout(n42000));
  jor  g23978(.dina(n42000), .dinb(n41998), .dout(n42001));
  jand g23979(.dina(n42001), .dinb(n405), .dout(n42002));
  jnot g23980(.din(n42002), .dout(n42003));
  jand g23981(.dina(n41640), .dinb(n41268), .dout(n42004));
  jxor g23982(.dina(n41474), .dinb(n41681), .dout(n42005));
  jand g23983(.dina(n42005), .dinb(n41770), .dout(n42006));
  jor  g23984(.dina(n42006), .dinb(n42004), .dout(n42007));
  jand g23985(.dina(n42007), .dinb(n2714), .dout(n42008));
  jnot g23986(.din(n42008), .dout(n42009));
  jand g23987(.dina(n41640), .dinb(n41274), .dout(n42010));
  jxor g23988(.dina(n41470), .dinb(n41679), .dout(n42011));
  jand g23989(.dina(n42011), .dinb(n41770), .dout(n42012));
  jor  g23990(.dina(n42012), .dinb(n42010), .dout(n42013));
  jand g23991(.dina(n42013), .dinb(n2547), .dout(n42014));
  jnot g23992(.din(n42014), .dout(n42015));
  jand g23993(.dina(n41640), .dinb(n41280), .dout(n42016));
  jxor g23994(.dina(n41466), .dinb(n41677), .dout(n42017));
  jand g23995(.dina(n42017), .dinb(n41770), .dout(n42018));
  jor  g23996(.dina(n42018), .dinb(n42016), .dout(n42019));
  jand g23997(.dina(n42019), .dinb(n417), .dout(n42020));
  jnot g23998(.din(n42020), .dout(n42021));
  jand g23999(.dina(n41640), .dinb(n41286), .dout(n42022));
  jxor g24000(.dina(n41462), .dinb(n41675), .dout(n42023));
  jand g24001(.dina(n42023), .dinb(n41770), .dout(n42024));
  jor  g24002(.dina(n42024), .dinb(n42022), .dout(n42025));
  jand g24003(.dina(n42025), .dinb(n416), .dout(n42026));
  jnot g24004(.din(n42026), .dout(n42027));
  jand g24005(.dina(n41640), .dinb(n41292), .dout(n42028));
  jxor g24006(.dina(n41458), .dinb(n41673), .dout(n42029));
  jand g24007(.dina(n42029), .dinb(n41770), .dout(n42030));
  jor  g24008(.dina(n42030), .dinb(n42028), .dout(n42031));
  jand g24009(.dina(n42031), .dinb(n422), .dout(n42032));
  jnot g24010(.din(n42032), .dout(n42033));
  jand g24011(.dina(n41640), .dinb(n41298), .dout(n42034));
  jxor g24012(.dina(n41454), .dinb(n41671), .dout(n42035));
  jand g24013(.dina(n42035), .dinb(n41770), .dout(n42036));
  jor  g24014(.dina(n42036), .dinb(n42034), .dout(n42037));
  jand g24015(.dina(n42037), .dinb(n421), .dout(n42038));
  jnot g24016(.din(n42038), .dout(n42039));
  jand g24017(.dina(n41640), .dinb(n41304), .dout(n42040));
  jxor g24018(.dina(n41450), .dinb(n41669), .dout(n42041));
  jand g24019(.dina(n42041), .dinb(n41770), .dout(n42042));
  jor  g24020(.dina(n42042), .dinb(n42040), .dout(n42043));
  jand g24021(.dina(n42043), .dinb(n433), .dout(n42044));
  jnot g24022(.din(n42044), .dout(n42045));
  jand g24023(.dina(n41640), .dinb(n41310), .dout(n42046));
  jxor g24024(.dina(n41446), .dinb(n41667), .dout(n42047));
  jand g24025(.dina(n42047), .dinb(n41770), .dout(n42048));
  jor  g24026(.dina(n42048), .dinb(n42046), .dout(n42049));
  jand g24027(.dina(n42049), .dinb(n432), .dout(n42050));
  jnot g24028(.din(n42050), .dout(n42051));
  jand g24029(.dina(n41640), .dinb(n41316), .dout(n42052));
  jxor g24030(.dina(n41442), .dinb(n41665), .dout(n42053));
  jand g24031(.dina(n42053), .dinb(n41770), .dout(n42054));
  jor  g24032(.dina(n42054), .dinb(n42052), .dout(n42055));
  jand g24033(.dina(n42055), .dinb(n436), .dout(n42056));
  jnot g24034(.din(n42056), .dout(n42057));
  jand g24035(.dina(n41640), .dinb(n41322), .dout(n42058));
  jxor g24036(.dina(n41438), .dinb(n41663), .dout(n42059));
  jand g24037(.dina(n42059), .dinb(n41770), .dout(n42060));
  jor  g24038(.dina(n42060), .dinb(n42058), .dout(n42061));
  jand g24039(.dina(n42061), .dinb(n435), .dout(n42062));
  jnot g24040(.din(n42062), .dout(n42063));
  jand g24041(.dina(n41640), .dinb(n41328), .dout(n42064));
  jxor g24042(.dina(n41434), .dinb(n41661), .dout(n42065));
  jand g24043(.dina(n42065), .dinb(n41770), .dout(n42066));
  jor  g24044(.dina(n42066), .dinb(n42064), .dout(n42067));
  jand g24045(.dina(n42067), .dinb(n440), .dout(n42068));
  jnot g24046(.din(n42068), .dout(n42069));
  jand g24047(.dina(n41640), .dinb(n41334), .dout(n42070));
  jxor g24048(.dina(n41430), .dinb(n41659), .dout(n42071));
  jand g24049(.dina(n42071), .dinb(n41770), .dout(n42072));
  jor  g24050(.dina(n42072), .dinb(n42070), .dout(n42073));
  jand g24051(.dina(n42073), .dinb(n439), .dout(n42074));
  jnot g24052(.din(n42074), .dout(n42075));
  jand g24053(.dina(n41640), .dinb(n41340), .dout(n42076));
  jxor g24054(.dina(n41426), .dinb(n41657), .dout(n42077));
  jand g24055(.dina(n42077), .dinb(n41770), .dout(n42078));
  jor  g24056(.dina(n42078), .dinb(n42076), .dout(n42079));
  jand g24057(.dina(n42079), .dinb(n325), .dout(n42080));
  jnot g24058(.din(n42080), .dout(n42081));
  jand g24059(.dina(n41640), .dinb(n41346), .dout(n42082));
  jxor g24060(.dina(n41422), .dinb(n41655), .dout(n42083));
  jand g24061(.dina(n42083), .dinb(n41770), .dout(n42084));
  jor  g24062(.dina(n42084), .dinb(n42082), .dout(n42085));
  jand g24063(.dina(n42085), .dinb(n324), .dout(n42086));
  jnot g24064(.din(n42086), .dout(n42087));
  jand g24065(.dina(n41640), .dinb(n41352), .dout(n42088));
  jxor g24066(.dina(n41418), .dinb(n41653), .dout(n42089));
  jand g24067(.dina(n42089), .dinb(n41770), .dout(n42090));
  jor  g24068(.dina(n42090), .dinb(n42088), .dout(n42091));
  jand g24069(.dina(n42091), .dinb(n323), .dout(n42092));
  jnot g24070(.din(n42092), .dout(n42093));
  jand g24071(.dina(n41640), .dinb(n41358), .dout(n42094));
  jxor g24072(.dina(n41414), .dinb(n41651), .dout(n42095));
  jand g24073(.dina(n42095), .dinb(n41770), .dout(n42096));
  jor  g24074(.dina(n42096), .dinb(n42094), .dout(n42097));
  jand g24075(.dina(n42097), .dinb(n335), .dout(n42098));
  jnot g24076(.din(n42098), .dout(n42099));
  jand g24077(.dina(n41640), .dinb(n41364), .dout(n42100));
  jxor g24078(.dina(n41410), .dinb(n41649), .dout(n42101));
  jand g24079(.dina(n42101), .dinb(n41770), .dout(n42102));
  jor  g24080(.dina(n42102), .dinb(n42100), .dout(n42103));
  jand g24081(.dina(n42103), .dinb(n334), .dout(n42104));
  jnot g24082(.din(n42104), .dout(n42105));
  jand g24083(.dina(n41640), .dinb(n41370), .dout(n42106));
  jxor g24084(.dina(n41406), .dinb(n41647), .dout(n42107));
  jand g24085(.dina(n42107), .dinb(n41770), .dout(n42108));
  jor  g24086(.dina(n42108), .dinb(n42106), .dout(n42109));
  jand g24087(.dina(n42109), .dinb(n338), .dout(n42110));
  jnot g24088(.din(n42110), .dout(n42111));
  jand g24089(.dina(n41640), .dinb(n41376), .dout(n42112));
  jxor g24090(.dina(n41402), .dinb(n41645), .dout(n42113));
  jand g24091(.dina(n42113), .dinb(n41770), .dout(n42114));
  jor  g24092(.dina(n42114), .dinb(n42112), .dout(n42115));
  jand g24093(.dina(n42115), .dinb(n337), .dout(n42116));
  jnot g24094(.din(n42116), .dout(n42117));
  jand g24095(.dina(n41640), .dinb(n41382), .dout(n42118));
  jxor g24096(.dina(n41398), .dinb(n41643), .dout(n42119));
  jand g24097(.dina(n42119), .dinb(n41770), .dout(n42120));
  jor  g24098(.dina(n42120), .dinb(n42118), .dout(n42121));
  jand g24099(.dina(n42121), .dinb(n344), .dout(n42122));
  jnot g24100(.din(n42122), .dout(n42123));
  jand g24101(.dina(n41640), .dinb(n41389), .dout(n42124));
  jxor g24102(.dina(n41641), .dinb(n17309), .dout(n42125));
  jand g24103(.dina(n42125), .dinb(n41770), .dout(n42126));
  jor  g24104(.dina(n42126), .dinb(n42124), .dout(n42127));
  jand g24105(.dina(n42127), .dinb(n348), .dout(n42128));
  jnot g24106(.din(n42128), .dout(n42129));
  jor  g24107(.dina(n41640), .dinb(n18364), .dout(n42130));
  jand g24108(.dina(n42130), .dinb(a2 ), .dout(n42131));
  jor  g24109(.dina(n41640), .dinb(n17309), .dout(n42132));
  jnot g24110(.din(n42132), .dout(n42133));
  jor  g24111(.dina(n42133), .dinb(n42131), .dout(n42134));
  jand g24112(.dina(n42134), .dinb(n258), .dout(n42135));
  jnot g24113(.din(n42135), .dout(n42136));
  jand g24114(.dina(n41770), .dinb(b0 ), .dout(n42137));
  jor  g24115(.dina(n42137), .dinb(n17307), .dout(n42138));
  jand g24116(.dina(n42132), .dinb(n42138), .dout(n42139));
  jxor g24117(.dina(n42139), .dinb(n258), .dout(n42140));
  jor  g24118(.dina(n42140), .dinb(n17811), .dout(n42141));
  jand g24119(.dina(n42141), .dinb(n42136), .dout(n42142));
  jxor g24120(.dina(n42127), .dinb(n348), .dout(n42143));
  jnot g24121(.din(n42143), .dout(n42144));
  jor  g24122(.dina(n42144), .dinb(n42142), .dout(n42145));
  jand g24123(.dina(n42145), .dinb(n42129), .dout(n42146));
  jxor g24124(.dina(n42121), .dinb(n344), .dout(n42147));
  jnot g24125(.din(n42147), .dout(n42148));
  jor  g24126(.dina(n42148), .dinb(n42146), .dout(n42149));
  jand g24127(.dina(n42149), .dinb(n42123), .dout(n42150));
  jxor g24128(.dina(n42115), .dinb(n337), .dout(n42151));
  jnot g24129(.din(n42151), .dout(n42152));
  jor  g24130(.dina(n42152), .dinb(n42150), .dout(n42153));
  jand g24131(.dina(n42153), .dinb(n42117), .dout(n42154));
  jxor g24132(.dina(n42109), .dinb(n338), .dout(n42155));
  jnot g24133(.din(n42155), .dout(n42156));
  jor  g24134(.dina(n42156), .dinb(n42154), .dout(n42157));
  jand g24135(.dina(n42157), .dinb(n42111), .dout(n42158));
  jxor g24136(.dina(n42103), .dinb(n334), .dout(n42159));
  jnot g24137(.din(n42159), .dout(n42160));
  jor  g24138(.dina(n42160), .dinb(n42158), .dout(n42161));
  jand g24139(.dina(n42161), .dinb(n42105), .dout(n42162));
  jxor g24140(.dina(n42097), .dinb(n335), .dout(n42163));
  jnot g24141(.din(n42163), .dout(n42164));
  jor  g24142(.dina(n42164), .dinb(n42162), .dout(n42165));
  jand g24143(.dina(n42165), .dinb(n42099), .dout(n42166));
  jxor g24144(.dina(n42091), .dinb(n323), .dout(n42167));
  jnot g24145(.din(n42167), .dout(n42168));
  jor  g24146(.dina(n42168), .dinb(n42166), .dout(n42169));
  jand g24147(.dina(n42169), .dinb(n42093), .dout(n42170));
  jxor g24148(.dina(n42085), .dinb(n324), .dout(n42171));
  jnot g24149(.din(n42171), .dout(n42172));
  jor  g24150(.dina(n42172), .dinb(n42170), .dout(n42173));
  jand g24151(.dina(n42173), .dinb(n42087), .dout(n42174));
  jxor g24152(.dina(n42079), .dinb(n325), .dout(n42175));
  jnot g24153(.din(n42175), .dout(n42176));
  jor  g24154(.dina(n42176), .dinb(n42174), .dout(n42177));
  jand g24155(.dina(n42177), .dinb(n42081), .dout(n42178));
  jxor g24156(.dina(n42073), .dinb(n439), .dout(n42179));
  jnot g24157(.din(n42179), .dout(n42180));
  jor  g24158(.dina(n42180), .dinb(n42178), .dout(n42181));
  jand g24159(.dina(n42181), .dinb(n42075), .dout(n42182));
  jxor g24160(.dina(n42067), .dinb(n440), .dout(n42183));
  jnot g24161(.din(n42183), .dout(n42184));
  jor  g24162(.dina(n42184), .dinb(n42182), .dout(n42185));
  jand g24163(.dina(n42185), .dinb(n42069), .dout(n42186));
  jxor g24164(.dina(n42061), .dinb(n435), .dout(n42187));
  jnot g24165(.din(n42187), .dout(n42188));
  jor  g24166(.dina(n42188), .dinb(n42186), .dout(n42189));
  jand g24167(.dina(n42189), .dinb(n42063), .dout(n42190));
  jxor g24168(.dina(n42055), .dinb(n436), .dout(n42191));
  jnot g24169(.din(n42191), .dout(n42192));
  jor  g24170(.dina(n42192), .dinb(n42190), .dout(n42193));
  jand g24171(.dina(n42193), .dinb(n42057), .dout(n42194));
  jxor g24172(.dina(n42049), .dinb(n432), .dout(n42195));
  jnot g24173(.din(n42195), .dout(n42196));
  jor  g24174(.dina(n42196), .dinb(n42194), .dout(n42197));
  jand g24175(.dina(n42197), .dinb(n42051), .dout(n42198));
  jxor g24176(.dina(n42043), .dinb(n433), .dout(n42199));
  jnot g24177(.din(n42199), .dout(n42200));
  jor  g24178(.dina(n42200), .dinb(n42198), .dout(n42201));
  jand g24179(.dina(n42201), .dinb(n42045), .dout(n42202));
  jxor g24180(.dina(n42037), .dinb(n421), .dout(n42203));
  jnot g24181(.din(n42203), .dout(n42204));
  jor  g24182(.dina(n42204), .dinb(n42202), .dout(n42205));
  jand g24183(.dina(n42205), .dinb(n42039), .dout(n42206));
  jxor g24184(.dina(n42031), .dinb(n422), .dout(n42207));
  jnot g24185(.din(n42207), .dout(n42208));
  jor  g24186(.dina(n42208), .dinb(n42206), .dout(n42209));
  jand g24187(.dina(n42209), .dinb(n42033), .dout(n42210));
  jxor g24188(.dina(n42025), .dinb(n416), .dout(n42211));
  jnot g24189(.din(n42211), .dout(n42212));
  jor  g24190(.dina(n42212), .dinb(n42210), .dout(n42213));
  jand g24191(.dina(n42213), .dinb(n42027), .dout(n42214));
  jxor g24192(.dina(n42019), .dinb(n417), .dout(n42215));
  jnot g24193(.din(n42215), .dout(n42216));
  jor  g24194(.dina(n42216), .dinb(n42214), .dout(n42217));
  jand g24195(.dina(n42217), .dinb(n42021), .dout(n42218));
  jxor g24196(.dina(n42013), .dinb(n2547), .dout(n42219));
  jnot g24197(.din(n42219), .dout(n42220));
  jor  g24198(.dina(n42220), .dinb(n42218), .dout(n42221));
  jand g24199(.dina(n42221), .dinb(n42015), .dout(n42222));
  jxor g24200(.dina(n42007), .dinb(n2714), .dout(n42223));
  jnot g24201(.din(n42223), .dout(n42224));
  jor  g24202(.dina(n42224), .dinb(n42222), .dout(n42225));
  jand g24203(.dina(n42225), .dinb(n42009), .dout(n42226));
  jxor g24204(.dina(n42001), .dinb(n405), .dout(n42227));
  jnot g24205(.din(n42227), .dout(n42228));
  jor  g24206(.dina(n42228), .dinb(n42226), .dout(n42229));
  jand g24207(.dina(n42229), .dinb(n42003), .dout(n42230));
  jxor g24208(.dina(n41995), .dinb(n406), .dout(n42231));
  jnot g24209(.din(n42231), .dout(n42232));
  jor  g24210(.dina(n42232), .dinb(n42230), .dout(n42233));
  jand g24211(.dina(n42233), .dinb(n41997), .dout(n42234));
  jxor g24212(.dina(n41989), .dinb(n412), .dout(n42235));
  jnot g24213(.din(n42235), .dout(n42236));
  jor  g24214(.dina(n42236), .dinb(n42234), .dout(n42237));
  jand g24215(.dina(n42237), .dinb(n41991), .dout(n42238));
  jxor g24216(.dina(n41983), .dinb(n413), .dout(n42239));
  jnot g24217(.din(n42239), .dout(n42240));
  jor  g24218(.dina(n42240), .dinb(n42238), .dout(n42241));
  jand g24219(.dina(n42241), .dinb(n41985), .dout(n42242));
  jxor g24220(.dina(n41977), .dinb(n409), .dout(n42243));
  jnot g24221(.din(n42243), .dout(n42244));
  jor  g24222(.dina(n42244), .dinb(n42242), .dout(n42245));
  jand g24223(.dina(n42245), .dinb(n41979), .dout(n42246));
  jxor g24224(.dina(n41971), .dinb(n410), .dout(n42247));
  jnot g24225(.din(n42247), .dout(n42248));
  jor  g24226(.dina(n42248), .dinb(n42246), .dout(n42249));
  jand g24227(.dina(n42249), .dinb(n41973), .dout(n42250));
  jxor g24228(.dina(n41965), .dinb(n426), .dout(n42251));
  jnot g24229(.din(n42251), .dout(n42252));
  jor  g24230(.dina(n42252), .dinb(n42250), .dout(n42253));
  jand g24231(.dina(n42253), .dinb(n41967), .dout(n42254));
  jxor g24232(.dina(n41959), .dinb(n427), .dout(n42255));
  jnot g24233(.din(n42255), .dout(n42256));
  jor  g24234(.dina(n42256), .dinb(n42254), .dout(n42257));
  jand g24235(.dina(n42257), .dinb(n41961), .dout(n42258));
  jxor g24236(.dina(n41953), .dinb(n424), .dout(n42259));
  jnot g24237(.din(n42259), .dout(n42260));
  jor  g24238(.dina(n42260), .dinb(n42258), .dout(n42261));
  jand g24239(.dina(n42261), .dinb(n41955), .dout(n42262));
  jxor g24240(.dina(n41947), .dinb(n300), .dout(n42263));
  jnot g24241(.din(n42263), .dout(n42264));
  jor  g24242(.dina(n42264), .dinb(n42262), .dout(n42265));
  jand g24243(.dina(n42265), .dinb(n41949), .dout(n42266));
  jxor g24244(.dina(n41941), .dinb(n297), .dout(n42267));
  jnot g24245(.din(n42267), .dout(n42268));
  jor  g24246(.dina(n42268), .dinb(n42266), .dout(n42269));
  jand g24247(.dina(n42269), .dinb(n41943), .dout(n42270));
  jxor g24248(.dina(n41935), .dinb(n298), .dout(n42271));
  jnot g24249(.din(n42271), .dout(n42272));
  jor  g24250(.dina(n42272), .dinb(n42270), .dout(n42273));
  jand g24251(.dina(n42273), .dinb(n41937), .dout(n42274));
  jxor g24252(.dina(n41929), .dinb(n301), .dout(n42275));
  jnot g24253(.din(n42275), .dout(n42276));
  jor  g24254(.dina(n42276), .dinb(n42274), .dout(n42277));
  jand g24255(.dina(n42277), .dinb(n41931), .dout(n42278));
  jxor g24256(.dina(n41923), .dinb(n293), .dout(n42279));
  jnot g24257(.din(n42279), .dout(n42280));
  jor  g24258(.dina(n42280), .dinb(n42278), .dout(n42281));
  jand g24259(.dina(n42281), .dinb(n41925), .dout(n42282));
  jxor g24260(.dina(n41917), .dinb(n294), .dout(n42283));
  jnot g24261(.din(n42283), .dout(n42284));
  jor  g24262(.dina(n42284), .dinb(n42282), .dout(n42285));
  jand g24263(.dina(n42285), .dinb(n41919), .dout(n42286));
  jxor g24264(.dina(n41911), .dinb(n290), .dout(n42287));
  jnot g24265(.din(n42287), .dout(n42288));
  jor  g24266(.dina(n42288), .dinb(n42286), .dout(n42289));
  jand g24267(.dina(n42289), .dinb(n41913), .dout(n42290));
  jxor g24268(.dina(n41905), .dinb(n291), .dout(n42291));
  jnot g24269(.din(n42291), .dout(n42292));
  jor  g24270(.dina(n42292), .dinb(n42290), .dout(n42293));
  jand g24271(.dina(n42293), .dinb(n41907), .dout(n42294));
  jxor g24272(.dina(n41899), .dinb(n284), .dout(n42295));
  jnot g24273(.din(n42295), .dout(n42296));
  jor  g24274(.dina(n42296), .dinb(n42294), .dout(n42297));
  jand g24275(.dina(n42297), .dinb(n41901), .dout(n42298));
  jxor g24276(.dina(n41893), .dinb(n285), .dout(n42299));
  jnot g24277(.din(n42299), .dout(n42300));
  jor  g24278(.dina(n42300), .dinb(n42298), .dout(n42301));
  jand g24279(.dina(n42301), .dinb(n41895), .dout(n42302));
  jxor g24280(.dina(n41887), .dinb(n281), .dout(n42303));
  jnot g24281(.din(n42303), .dout(n42304));
  jor  g24282(.dina(n42304), .dinb(n42302), .dout(n42305));
  jand g24283(.dina(n42305), .dinb(n41889), .dout(n42306));
  jxor g24284(.dina(n41881), .dinb(n282), .dout(n42307));
  jnot g24285(.din(n42307), .dout(n42308));
  jor  g24286(.dina(n42308), .dinb(n42306), .dout(n42309));
  jand g24287(.dina(n42309), .dinb(n41883), .dout(n42310));
  jxor g24288(.dina(n41875), .dinb(n397), .dout(n42311));
  jnot g24289(.din(n42311), .dout(n42312));
  jor  g24290(.dina(n42312), .dinb(n42310), .dout(n42313));
  jand g24291(.dina(n42313), .dinb(n41877), .dout(n42314));
  jxor g24292(.dina(n41869), .dinb(n513), .dout(n42315));
  jnot g24293(.din(n42315), .dout(n42316));
  jor  g24294(.dina(n42316), .dinb(n42314), .dout(n42317));
  jand g24295(.dina(n42317), .dinb(n41871), .dout(n42318));
  jxor g24296(.dina(n41863), .dinb(n514), .dout(n42319));
  jnot g24297(.din(n42319), .dout(n42320));
  jor  g24298(.dina(n42320), .dinb(n42318), .dout(n42321));
  jand g24299(.dina(n42321), .dinb(n41865), .dout(n42322));
  jxor g24300(.dina(n41857), .dinb(n510), .dout(n42323));
  jnot g24301(.din(n42323), .dout(n42324));
  jor  g24302(.dina(n42324), .dinb(n42322), .dout(n42325));
  jand g24303(.dina(n42325), .dinb(n41859), .dout(n42326));
  jxor g24304(.dina(n41851), .dinb(n396), .dout(n42327));
  jnot g24305(.din(n42327), .dout(n42328));
  jor  g24306(.dina(n42328), .dinb(n42326), .dout(n42329));
  jand g24307(.dina(n42329), .dinb(n41853), .dout(n42330));
  jxor g24308(.dina(n41845), .dinb(n383), .dout(n42331));
  jnot g24309(.din(n42331), .dout(n42332));
  jor  g24310(.dina(n42332), .dinb(n42330), .dout(n42333));
  jand g24311(.dina(n42333), .dinb(n41847), .dout(n42334));
  jxor g24312(.dina(n41839), .dinb(n12211), .dout(n42335));
  jnot g24313(.din(n42335), .dout(n42336));
  jor  g24314(.dina(n42336), .dinb(n42334), .dout(n42337));
  jand g24315(.dina(n42337), .dinb(n41841), .dout(n42338));
  jxor g24316(.dina(n41833), .dinb(n12214), .dout(n42339));
  jnot g24317(.din(n42339), .dout(n42340));
  jor  g24318(.dina(n42340), .dinb(n42338), .dout(n42341));
  jand g24319(.dina(n42341), .dinb(n41835), .dout(n42342));
  jxor g24320(.dina(n41827), .dinb(n384), .dout(n42343));
  jnot g24321(.din(n42343), .dout(n42344));
  jor  g24322(.dina(n42344), .dinb(n42342), .dout(n42345));
  jand g24323(.dina(n42345), .dinb(n41829), .dout(n42346));
  jxor g24324(.dina(n41821), .dinb(n374), .dout(n42347));
  jnot g24325(.din(n42347), .dout(n42348));
  jor  g24326(.dina(n42348), .dinb(n42346), .dout(n42349));
  jand g24327(.dina(n42349), .dinb(n41823), .dout(n42350));
  jxor g24328(.dina(n41815), .dinb(n376), .dout(n42351));
  jnot g24329(.din(n42351), .dout(n42352));
  jor  g24330(.dina(n42352), .dinb(n42350), .dout(n42353));
  jand g24331(.dina(n42353), .dinb(n41817), .dout(n42354));
  jxor g24332(.dina(n41809), .dinb(n377), .dout(n42355));
  jnot g24333(.din(n42355), .dout(n42356));
  jor  g24334(.dina(n42356), .dinb(n42354), .dout(n42357));
  jand g24335(.dina(n42357), .dinb(n41811), .dout(n42358));
  jxor g24336(.dina(n41803), .dinb(n375), .dout(n42359));
  jnot g24337(.din(n42359), .dout(n42360));
  jor  g24338(.dina(n42360), .dinb(n42358), .dout(n42361));
  jand g24339(.dina(n42361), .dinb(n41805), .dout(n42362));
  jxor g24340(.dina(n41797), .dinb(n362), .dout(n42363));
  jnot g24341(.din(n42363), .dout(n42364));
  jor  g24342(.dina(n42364), .dinb(n42362), .dout(n42365));
  jand g24343(.dina(n42365), .dinb(n41799), .dout(n42366));
  jxor g24344(.dina(n41791), .dinb(n363), .dout(n42367));
  jnot g24345(.din(n42367), .dout(n42368));
  jor  g24346(.dina(n42368), .dinb(n42366), .dout(n42369));
  jand g24347(.dina(n42369), .dinb(n41793), .dout(n42370));
  jxor g24348(.dina(n41785), .dinb(n365), .dout(n42371));
  jnot g24349(.din(n42371), .dout(n42372));
  jor  g24350(.dina(n42372), .dinb(n42370), .dout(n42373));
  jand g24351(.dina(n42373), .dinb(n41787), .dout(n42374));
  jxor g24352(.dina(n41779), .dinb(n366), .dout(n42375));
  jnot g24353(.din(n42375), .dout(n42376));
  jor  g24354(.dina(n42376), .dinb(n42374), .dout(n42377));
  jand g24355(.dina(n42377), .dinb(n41781), .dout(n42378));
  jxor g24356(.dina(n41773), .dinb(n256), .dout(n42379));
  jnot g24357(.din(n42379), .dout(n42380));
  jor  g24358(.dina(n42380), .dinb(n42378), .dout(n42381));
  jand g24359(.dina(n42381), .dinb(n41775), .dout(n42382));
  jand g24360(.dina(n41764), .dinb(n367), .dout(n42383));
  jnot g24361(.din(n42383), .dout(n42384));
  jand g24362(.dina(n42384), .dinb(n42382), .dout(n42385));
  jand g24363(.dina(n41765), .dinb(b62 ), .dout(n42386));
  jor  g24364(.dina(n42386), .dinb(b63 ), .dout(n42387));
  jor  g24365(.dina(n42387), .dinb(n42385), .dout(n42388));
  jxor g24366(.dina(n42139), .dinb(b1 ), .dout(n42389));
  jand g24367(.dina(n42389), .dinb(n17812), .dout(n42390));
  jor  g24368(.dina(n42390), .dinb(n42135), .dout(n42391));
  jand g24369(.dina(n42143), .dinb(n42391), .dout(n42392));
  jor  g24370(.dina(n42392), .dinb(n42128), .dout(n42393));
  jand g24371(.dina(n42147), .dinb(n42393), .dout(n42394));
  jor  g24372(.dina(n42394), .dinb(n42122), .dout(n42395));
  jand g24373(.dina(n42151), .dinb(n42395), .dout(n42396));
  jor  g24374(.dina(n42396), .dinb(n42116), .dout(n42397));
  jand g24375(.dina(n42155), .dinb(n42397), .dout(n42398));
  jor  g24376(.dina(n42398), .dinb(n42110), .dout(n42399));
  jand g24377(.dina(n42159), .dinb(n42399), .dout(n42400));
  jor  g24378(.dina(n42400), .dinb(n42104), .dout(n42401));
  jand g24379(.dina(n42163), .dinb(n42401), .dout(n42402));
  jor  g24380(.dina(n42402), .dinb(n42098), .dout(n42403));
  jand g24381(.dina(n42167), .dinb(n42403), .dout(n42404));
  jor  g24382(.dina(n42404), .dinb(n42092), .dout(n42405));
  jand g24383(.dina(n42171), .dinb(n42405), .dout(n42406));
  jor  g24384(.dina(n42406), .dinb(n42086), .dout(n42407));
  jand g24385(.dina(n42175), .dinb(n42407), .dout(n42408));
  jor  g24386(.dina(n42408), .dinb(n42080), .dout(n42409));
  jand g24387(.dina(n42179), .dinb(n42409), .dout(n42410));
  jor  g24388(.dina(n42410), .dinb(n42074), .dout(n42411));
  jand g24389(.dina(n42183), .dinb(n42411), .dout(n42412));
  jor  g24390(.dina(n42412), .dinb(n42068), .dout(n42413));
  jand g24391(.dina(n42187), .dinb(n42413), .dout(n42414));
  jor  g24392(.dina(n42414), .dinb(n42062), .dout(n42415));
  jand g24393(.dina(n42191), .dinb(n42415), .dout(n42416));
  jor  g24394(.dina(n42416), .dinb(n42056), .dout(n42417));
  jand g24395(.dina(n42195), .dinb(n42417), .dout(n42418));
  jor  g24396(.dina(n42418), .dinb(n42050), .dout(n42419));
  jand g24397(.dina(n42199), .dinb(n42419), .dout(n42420));
  jor  g24398(.dina(n42420), .dinb(n42044), .dout(n42421));
  jand g24399(.dina(n42203), .dinb(n42421), .dout(n42422));
  jor  g24400(.dina(n42422), .dinb(n42038), .dout(n42423));
  jand g24401(.dina(n42207), .dinb(n42423), .dout(n42424));
  jor  g24402(.dina(n42424), .dinb(n42032), .dout(n42425));
  jand g24403(.dina(n42211), .dinb(n42425), .dout(n42426));
  jor  g24404(.dina(n42426), .dinb(n42026), .dout(n42427));
  jand g24405(.dina(n42215), .dinb(n42427), .dout(n42428));
  jor  g24406(.dina(n42428), .dinb(n42020), .dout(n42429));
  jand g24407(.dina(n42219), .dinb(n42429), .dout(n42430));
  jor  g24408(.dina(n42430), .dinb(n42014), .dout(n42431));
  jand g24409(.dina(n42223), .dinb(n42431), .dout(n42432));
  jor  g24410(.dina(n42432), .dinb(n42008), .dout(n42433));
  jand g24411(.dina(n42227), .dinb(n42433), .dout(n42434));
  jor  g24412(.dina(n42434), .dinb(n42002), .dout(n42435));
  jand g24413(.dina(n42231), .dinb(n42435), .dout(n42436));
  jor  g24414(.dina(n42436), .dinb(n41996), .dout(n42437));
  jand g24415(.dina(n42235), .dinb(n42437), .dout(n42438));
  jor  g24416(.dina(n42438), .dinb(n41990), .dout(n42439));
  jand g24417(.dina(n42239), .dinb(n42439), .dout(n42440));
  jor  g24418(.dina(n42440), .dinb(n41984), .dout(n42441));
  jand g24419(.dina(n42243), .dinb(n42441), .dout(n42442));
  jor  g24420(.dina(n42442), .dinb(n41978), .dout(n42443));
  jand g24421(.dina(n42247), .dinb(n42443), .dout(n42444));
  jor  g24422(.dina(n42444), .dinb(n41972), .dout(n42445));
  jand g24423(.dina(n42251), .dinb(n42445), .dout(n42446));
  jor  g24424(.dina(n42446), .dinb(n41966), .dout(n42447));
  jand g24425(.dina(n42255), .dinb(n42447), .dout(n42448));
  jor  g24426(.dina(n42448), .dinb(n41960), .dout(n42449));
  jand g24427(.dina(n42259), .dinb(n42449), .dout(n42450));
  jor  g24428(.dina(n42450), .dinb(n41954), .dout(n42451));
  jand g24429(.dina(n42263), .dinb(n42451), .dout(n42452));
  jor  g24430(.dina(n42452), .dinb(n41948), .dout(n42453));
  jand g24431(.dina(n42267), .dinb(n42453), .dout(n42454));
  jor  g24432(.dina(n42454), .dinb(n41942), .dout(n42455));
  jand g24433(.dina(n42271), .dinb(n42455), .dout(n42456));
  jor  g24434(.dina(n42456), .dinb(n41936), .dout(n42457));
  jand g24435(.dina(n42275), .dinb(n42457), .dout(n42458));
  jor  g24436(.dina(n42458), .dinb(n41930), .dout(n42459));
  jand g24437(.dina(n42279), .dinb(n42459), .dout(n42460));
  jor  g24438(.dina(n42460), .dinb(n41924), .dout(n42461));
  jand g24439(.dina(n42283), .dinb(n42461), .dout(n42462));
  jor  g24440(.dina(n42462), .dinb(n41918), .dout(n42463));
  jand g24441(.dina(n42287), .dinb(n42463), .dout(n42464));
  jor  g24442(.dina(n42464), .dinb(n41912), .dout(n42465));
  jand g24443(.dina(n42291), .dinb(n42465), .dout(n42466));
  jor  g24444(.dina(n42466), .dinb(n41906), .dout(n42467));
  jand g24445(.dina(n42295), .dinb(n42467), .dout(n42468));
  jor  g24446(.dina(n42468), .dinb(n41900), .dout(n42469));
  jand g24447(.dina(n42299), .dinb(n42469), .dout(n42470));
  jor  g24448(.dina(n42470), .dinb(n41894), .dout(n42471));
  jand g24449(.dina(n42303), .dinb(n42471), .dout(n42472));
  jor  g24450(.dina(n42472), .dinb(n41888), .dout(n42473));
  jand g24451(.dina(n42307), .dinb(n42473), .dout(n42474));
  jor  g24452(.dina(n42474), .dinb(n41882), .dout(n42475));
  jand g24453(.dina(n42311), .dinb(n42475), .dout(n42476));
  jor  g24454(.dina(n42476), .dinb(n41876), .dout(n42477));
  jand g24455(.dina(n42315), .dinb(n42477), .dout(n42478));
  jor  g24456(.dina(n42478), .dinb(n41870), .dout(n42479));
  jand g24457(.dina(n42319), .dinb(n42479), .dout(n42480));
  jor  g24458(.dina(n42480), .dinb(n41864), .dout(n42481));
  jand g24459(.dina(n42323), .dinb(n42481), .dout(n42482));
  jor  g24460(.dina(n42482), .dinb(n41858), .dout(n42483));
  jand g24461(.dina(n42327), .dinb(n42483), .dout(n42484));
  jor  g24462(.dina(n42484), .dinb(n41852), .dout(n42485));
  jand g24463(.dina(n42331), .dinb(n42485), .dout(n42486));
  jor  g24464(.dina(n42486), .dinb(n41846), .dout(n42487));
  jand g24465(.dina(n42335), .dinb(n42487), .dout(n42488));
  jor  g24466(.dina(n42488), .dinb(n41840), .dout(n42489));
  jand g24467(.dina(n42339), .dinb(n42489), .dout(n42490));
  jor  g24468(.dina(n42490), .dinb(n41834), .dout(n42491));
  jand g24469(.dina(n42343), .dinb(n42491), .dout(n42492));
  jor  g24470(.dina(n42492), .dinb(n41828), .dout(n42493));
  jand g24471(.dina(n42347), .dinb(n42493), .dout(n42494));
  jor  g24472(.dina(n42494), .dinb(n41822), .dout(n42495));
  jand g24473(.dina(n42351), .dinb(n42495), .dout(n42496));
  jor  g24474(.dina(n42496), .dinb(n41816), .dout(n42497));
  jand g24475(.dina(n42355), .dinb(n42497), .dout(n42498));
  jor  g24476(.dina(n42498), .dinb(n41810), .dout(n42499));
  jand g24477(.dina(n42359), .dinb(n42499), .dout(n42500));
  jor  g24478(.dina(n42500), .dinb(n41804), .dout(n42501));
  jand g24479(.dina(n42363), .dinb(n42501), .dout(n42502));
  jor  g24480(.dina(n42502), .dinb(n41798), .dout(n42503));
  jand g24481(.dina(n42367), .dinb(n42503), .dout(n42504));
  jor  g24482(.dina(n42504), .dinb(n41792), .dout(n42505));
  jand g24483(.dina(n42371), .dinb(n42505), .dout(n42506));
  jor  g24484(.dina(n42506), .dinb(n41786), .dout(n42507));
  jand g24485(.dina(n42375), .dinb(n42507), .dout(n42508));
  jor  g24486(.dina(n42508), .dinb(n41780), .dout(n42509));
  jand g24487(.dina(n42379), .dinb(n42509), .dout(n42510));
  jor  g24488(.dina(n42510), .dinb(n41774), .dout(n42511));
  jand g24489(.dina(n42511), .dinb(n369), .dout(n42512));
  jor  g24490(.dina(n42512), .dinb(n42388), .dout(n42513));
  jand g24491(.dina(n42513), .dinb(n41764), .dout(n42514));
  jand g24492(.dina(n42514), .dinb(n368), .dout(n42515));
  jnot g24493(.din(n42515), .dout(n42516));
  jand g24494(.dina(n42388), .dinb(n41773), .dout(n42517));
  jor  g24495(.dina(n42383), .dinb(n42511), .dout(n42518));
  jnot g24496(.din(n42387), .dout(n42519));
  jand g24497(.dina(n42519), .dinb(n42518), .dout(n42520));
  jxor g24498(.dina(n42379), .dinb(n42509), .dout(n42521));
  jand g24499(.dina(n42521), .dinb(n42520), .dout(n42522));
  jor  g24500(.dina(n42522), .dinb(n42517), .dout(n42523));
  jand g24501(.dina(n42523), .dinb(n367), .dout(n42524));
  jnot g24502(.din(n42524), .dout(n42525));
  jand g24503(.dina(n42388), .dinb(n41779), .dout(n42526));
  jxor g24504(.dina(n42375), .dinb(n42507), .dout(n42527));
  jand g24505(.dina(n42527), .dinb(n42520), .dout(n42528));
  jor  g24506(.dina(n42528), .dinb(n42526), .dout(n42529));
  jand g24507(.dina(n42529), .dinb(n256), .dout(n42530));
  jnot g24508(.din(n42530), .dout(n42531));
  jand g24509(.dina(n42388), .dinb(n41785), .dout(n42532));
  jxor g24510(.dina(n42371), .dinb(n42505), .dout(n42533));
  jand g24511(.dina(n42533), .dinb(n42520), .dout(n42534));
  jor  g24512(.dina(n42534), .dinb(n42532), .dout(n42535));
  jand g24513(.dina(n42535), .dinb(n366), .dout(n42536));
  jnot g24514(.din(n42536), .dout(n42537));
  jand g24515(.dina(n42388), .dinb(n41791), .dout(n42538));
  jxor g24516(.dina(n42367), .dinb(n42503), .dout(n42539));
  jand g24517(.dina(n42539), .dinb(n42520), .dout(n42540));
  jor  g24518(.dina(n42540), .dinb(n42538), .dout(n42541));
  jand g24519(.dina(n42541), .dinb(n365), .dout(n42542));
  jnot g24520(.din(n42542), .dout(n42543));
  jand g24521(.dina(n42388), .dinb(n41797), .dout(n42544));
  jxor g24522(.dina(n42363), .dinb(n42501), .dout(n42545));
  jand g24523(.dina(n42545), .dinb(n42520), .dout(n42546));
  jor  g24524(.dina(n42546), .dinb(n42544), .dout(n42547));
  jand g24525(.dina(n42547), .dinb(n363), .dout(n42548));
  jnot g24526(.din(n42548), .dout(n42549));
  jand g24527(.dina(n42388), .dinb(n41803), .dout(n42550));
  jxor g24528(.dina(n42359), .dinb(n42499), .dout(n42551));
  jand g24529(.dina(n42551), .dinb(n42520), .dout(n42552));
  jor  g24530(.dina(n42552), .dinb(n42550), .dout(n42553));
  jand g24531(.dina(n42553), .dinb(n362), .dout(n42554));
  jnot g24532(.din(n42554), .dout(n42555));
  jand g24533(.dina(n42388), .dinb(n41809), .dout(n42556));
  jxor g24534(.dina(n42355), .dinb(n42497), .dout(n42557));
  jand g24535(.dina(n42557), .dinb(n42520), .dout(n42558));
  jor  g24536(.dina(n42558), .dinb(n42556), .dout(n42559));
  jand g24537(.dina(n42559), .dinb(n375), .dout(n42560));
  jnot g24538(.din(n42560), .dout(n42561));
  jand g24539(.dina(n42388), .dinb(n41815), .dout(n42562));
  jxor g24540(.dina(n42351), .dinb(n42495), .dout(n42563));
  jand g24541(.dina(n42563), .dinb(n42520), .dout(n42564));
  jor  g24542(.dina(n42564), .dinb(n42562), .dout(n42565));
  jand g24543(.dina(n42565), .dinb(n377), .dout(n42566));
  jnot g24544(.din(n42566), .dout(n42567));
  jand g24545(.dina(n42388), .dinb(n41821), .dout(n42568));
  jxor g24546(.dina(n42347), .dinb(n42493), .dout(n42569));
  jand g24547(.dina(n42569), .dinb(n42520), .dout(n42570));
  jor  g24548(.dina(n42570), .dinb(n42568), .dout(n42571));
  jand g24549(.dina(n42571), .dinb(n376), .dout(n42572));
  jnot g24550(.din(n42572), .dout(n42573));
  jand g24551(.dina(n42388), .dinb(n41827), .dout(n42574));
  jxor g24552(.dina(n42343), .dinb(n42491), .dout(n42575));
  jand g24553(.dina(n42575), .dinb(n42520), .dout(n42576));
  jor  g24554(.dina(n42576), .dinb(n42574), .dout(n42577));
  jand g24555(.dina(n42577), .dinb(n374), .dout(n42578));
  jnot g24556(.din(n42578), .dout(n42579));
  jand g24557(.dina(n42388), .dinb(n41833), .dout(n42580));
  jxor g24558(.dina(n42339), .dinb(n42489), .dout(n42581));
  jand g24559(.dina(n42581), .dinb(n42520), .dout(n42582));
  jor  g24560(.dina(n42582), .dinb(n42580), .dout(n42583));
  jand g24561(.dina(n42583), .dinb(n384), .dout(n42584));
  jnot g24562(.din(n42584), .dout(n42585));
  jand g24563(.dina(n42388), .dinb(n41839), .dout(n42586));
  jxor g24564(.dina(n42335), .dinb(n42487), .dout(n42587));
  jand g24565(.dina(n42587), .dinb(n42520), .dout(n42588));
  jor  g24566(.dina(n42588), .dinb(n42586), .dout(n42589));
  jand g24567(.dina(n42589), .dinb(n12214), .dout(n42590));
  jnot g24568(.din(n42590), .dout(n42591));
  jand g24569(.dina(n42388), .dinb(n41845), .dout(n42592));
  jxor g24570(.dina(n42331), .dinb(n42485), .dout(n42593));
  jand g24571(.dina(n42593), .dinb(n42520), .dout(n42594));
  jor  g24572(.dina(n42594), .dinb(n42592), .dout(n42595));
  jand g24573(.dina(n42595), .dinb(n12211), .dout(n42596));
  jnot g24574(.din(n42596), .dout(n42597));
  jand g24575(.dina(n42388), .dinb(n41851), .dout(n42598));
  jxor g24576(.dina(n42327), .dinb(n42483), .dout(n42599));
  jand g24577(.dina(n42599), .dinb(n42520), .dout(n42600));
  jor  g24578(.dina(n42600), .dinb(n42598), .dout(n42601));
  jand g24579(.dina(n42601), .dinb(n383), .dout(n42602));
  jnot g24580(.din(n42602), .dout(n42603));
  jand g24581(.dina(n42388), .dinb(n41857), .dout(n42604));
  jxor g24582(.dina(n42323), .dinb(n42481), .dout(n42605));
  jand g24583(.dina(n42605), .dinb(n42520), .dout(n42606));
  jor  g24584(.dina(n42606), .dinb(n42604), .dout(n42607));
  jand g24585(.dina(n42607), .dinb(n396), .dout(n42608));
  jnot g24586(.din(n42608), .dout(n42609));
  jand g24587(.dina(n42388), .dinb(n41863), .dout(n42610));
  jxor g24588(.dina(n42319), .dinb(n42479), .dout(n42611));
  jand g24589(.dina(n42611), .dinb(n42520), .dout(n42612));
  jor  g24590(.dina(n42612), .dinb(n42610), .dout(n42613));
  jand g24591(.dina(n42613), .dinb(n510), .dout(n42614));
  jnot g24592(.din(n42614), .dout(n42615));
  jand g24593(.dina(n42388), .dinb(n41869), .dout(n42616));
  jxor g24594(.dina(n42315), .dinb(n42477), .dout(n42617));
  jand g24595(.dina(n42617), .dinb(n42520), .dout(n42618));
  jor  g24596(.dina(n42618), .dinb(n42616), .dout(n42619));
  jand g24597(.dina(n42619), .dinb(n514), .dout(n42620));
  jnot g24598(.din(n42620), .dout(n42621));
  jand g24599(.dina(n42388), .dinb(n41875), .dout(n42622));
  jxor g24600(.dina(n42311), .dinb(n42475), .dout(n42623));
  jand g24601(.dina(n42623), .dinb(n42520), .dout(n42624));
  jor  g24602(.dina(n42624), .dinb(n42622), .dout(n42625));
  jand g24603(.dina(n42625), .dinb(n513), .dout(n42626));
  jnot g24604(.din(n42626), .dout(n42627));
  jand g24605(.dina(n42388), .dinb(n41881), .dout(n42628));
  jxor g24606(.dina(n42307), .dinb(n42473), .dout(n42629));
  jand g24607(.dina(n42629), .dinb(n42520), .dout(n42630));
  jor  g24608(.dina(n42630), .dinb(n42628), .dout(n42631));
  jand g24609(.dina(n42631), .dinb(n397), .dout(n42632));
  jnot g24610(.din(n42632), .dout(n42633));
  jand g24611(.dina(n42388), .dinb(n41887), .dout(n42634));
  jxor g24612(.dina(n42303), .dinb(n42471), .dout(n42635));
  jand g24613(.dina(n42635), .dinb(n42520), .dout(n42636));
  jor  g24614(.dina(n42636), .dinb(n42634), .dout(n42637));
  jand g24615(.dina(n42637), .dinb(n282), .dout(n42638));
  jnot g24616(.din(n42638), .dout(n42639));
  jand g24617(.dina(n42388), .dinb(n41893), .dout(n42640));
  jxor g24618(.dina(n42299), .dinb(n42469), .dout(n42641));
  jand g24619(.dina(n42641), .dinb(n42520), .dout(n42642));
  jor  g24620(.dina(n42642), .dinb(n42640), .dout(n42643));
  jand g24621(.dina(n42643), .dinb(n281), .dout(n42644));
  jnot g24622(.din(n42644), .dout(n42645));
  jand g24623(.dina(n42388), .dinb(n41899), .dout(n42646));
  jxor g24624(.dina(n42295), .dinb(n42467), .dout(n42647));
  jand g24625(.dina(n42647), .dinb(n42520), .dout(n42648));
  jor  g24626(.dina(n42648), .dinb(n42646), .dout(n42649));
  jand g24627(.dina(n42649), .dinb(n285), .dout(n42650));
  jnot g24628(.din(n42650), .dout(n42651));
  jand g24629(.dina(n42388), .dinb(n41905), .dout(n42652));
  jxor g24630(.dina(n42291), .dinb(n42465), .dout(n42653));
  jand g24631(.dina(n42653), .dinb(n42520), .dout(n42654));
  jor  g24632(.dina(n42654), .dinb(n42652), .dout(n42655));
  jand g24633(.dina(n42655), .dinb(n284), .dout(n42656));
  jnot g24634(.din(n42656), .dout(n42657));
  jand g24635(.dina(n42388), .dinb(n41911), .dout(n42658));
  jxor g24636(.dina(n42287), .dinb(n42463), .dout(n42659));
  jand g24637(.dina(n42659), .dinb(n42520), .dout(n42660));
  jor  g24638(.dina(n42660), .dinb(n42658), .dout(n42661));
  jand g24639(.dina(n42661), .dinb(n291), .dout(n42662));
  jnot g24640(.din(n42662), .dout(n42663));
  jand g24641(.dina(n42388), .dinb(n41917), .dout(n42664));
  jxor g24642(.dina(n42283), .dinb(n42461), .dout(n42665));
  jand g24643(.dina(n42665), .dinb(n42520), .dout(n42666));
  jor  g24644(.dina(n42666), .dinb(n42664), .dout(n42667));
  jand g24645(.dina(n42667), .dinb(n290), .dout(n42668));
  jnot g24646(.din(n42668), .dout(n42669));
  jand g24647(.dina(n42388), .dinb(n41923), .dout(n42670));
  jxor g24648(.dina(n42279), .dinb(n42459), .dout(n42671));
  jand g24649(.dina(n42671), .dinb(n42520), .dout(n42672));
  jor  g24650(.dina(n42672), .dinb(n42670), .dout(n42673));
  jand g24651(.dina(n42673), .dinb(n294), .dout(n42674));
  jnot g24652(.din(n42674), .dout(n42675));
  jand g24653(.dina(n42388), .dinb(n41929), .dout(n42676));
  jxor g24654(.dina(n42275), .dinb(n42457), .dout(n42677));
  jand g24655(.dina(n42677), .dinb(n42520), .dout(n42678));
  jor  g24656(.dina(n42678), .dinb(n42676), .dout(n42679));
  jand g24657(.dina(n42679), .dinb(n293), .dout(n42680));
  jnot g24658(.din(n42680), .dout(n42681));
  jand g24659(.dina(n42388), .dinb(n41935), .dout(n42682));
  jxor g24660(.dina(n42271), .dinb(n42455), .dout(n42683));
  jand g24661(.dina(n42683), .dinb(n42520), .dout(n42684));
  jor  g24662(.dina(n42684), .dinb(n42682), .dout(n42685));
  jand g24663(.dina(n42685), .dinb(n301), .dout(n42686));
  jnot g24664(.din(n42686), .dout(n42687));
  jand g24665(.dina(n42388), .dinb(n41941), .dout(n42688));
  jxor g24666(.dina(n42267), .dinb(n42453), .dout(n42689));
  jand g24667(.dina(n42689), .dinb(n42520), .dout(n42690));
  jor  g24668(.dina(n42690), .dinb(n42688), .dout(n42691));
  jand g24669(.dina(n42691), .dinb(n298), .dout(n42692));
  jnot g24670(.din(n42692), .dout(n42693));
  jand g24671(.dina(n42388), .dinb(n41947), .dout(n42694));
  jxor g24672(.dina(n42263), .dinb(n42451), .dout(n42695));
  jand g24673(.dina(n42695), .dinb(n42520), .dout(n42696));
  jor  g24674(.dina(n42696), .dinb(n42694), .dout(n42697));
  jand g24675(.dina(n42697), .dinb(n297), .dout(n42698));
  jnot g24676(.din(n42698), .dout(n42699));
  jand g24677(.dina(n42388), .dinb(n41953), .dout(n42700));
  jxor g24678(.dina(n42259), .dinb(n42449), .dout(n42701));
  jand g24679(.dina(n42701), .dinb(n42520), .dout(n42702));
  jor  g24680(.dina(n42702), .dinb(n42700), .dout(n42703));
  jand g24681(.dina(n42703), .dinb(n300), .dout(n42704));
  jnot g24682(.din(n42704), .dout(n42705));
  jand g24683(.dina(n42388), .dinb(n41959), .dout(n42706));
  jxor g24684(.dina(n42255), .dinb(n42447), .dout(n42707));
  jand g24685(.dina(n42707), .dinb(n42520), .dout(n42708));
  jor  g24686(.dina(n42708), .dinb(n42706), .dout(n42709));
  jand g24687(.dina(n42709), .dinb(n424), .dout(n42710));
  jnot g24688(.din(n42710), .dout(n42711));
  jand g24689(.dina(n42388), .dinb(n41965), .dout(n42712));
  jxor g24690(.dina(n42251), .dinb(n42445), .dout(n42713));
  jand g24691(.dina(n42713), .dinb(n42520), .dout(n42714));
  jor  g24692(.dina(n42714), .dinb(n42712), .dout(n42715));
  jand g24693(.dina(n42715), .dinb(n427), .dout(n42716));
  jnot g24694(.din(n42716), .dout(n42717));
  jand g24695(.dina(n42388), .dinb(n41971), .dout(n42718));
  jxor g24696(.dina(n42247), .dinb(n42443), .dout(n42719));
  jand g24697(.dina(n42719), .dinb(n42520), .dout(n42720));
  jor  g24698(.dina(n42720), .dinb(n42718), .dout(n42721));
  jand g24699(.dina(n42721), .dinb(n426), .dout(n42722));
  jnot g24700(.din(n42722), .dout(n42723));
  jand g24701(.dina(n42388), .dinb(n41977), .dout(n42724));
  jxor g24702(.dina(n42243), .dinb(n42441), .dout(n42725));
  jand g24703(.dina(n42725), .dinb(n42520), .dout(n42726));
  jor  g24704(.dina(n42726), .dinb(n42724), .dout(n42727));
  jand g24705(.dina(n42727), .dinb(n410), .dout(n42728));
  jnot g24706(.din(n42728), .dout(n42729));
  jand g24707(.dina(n42388), .dinb(n41983), .dout(n42730));
  jxor g24708(.dina(n42239), .dinb(n42439), .dout(n42731));
  jand g24709(.dina(n42731), .dinb(n42520), .dout(n42732));
  jor  g24710(.dina(n42732), .dinb(n42730), .dout(n42733));
  jand g24711(.dina(n42733), .dinb(n409), .dout(n42734));
  jnot g24712(.din(n42734), .dout(n42735));
  jand g24713(.dina(n42388), .dinb(n41989), .dout(n42736));
  jxor g24714(.dina(n42235), .dinb(n42437), .dout(n42737));
  jand g24715(.dina(n42737), .dinb(n42520), .dout(n42738));
  jor  g24716(.dina(n42738), .dinb(n42736), .dout(n42739));
  jand g24717(.dina(n42739), .dinb(n413), .dout(n42740));
  jnot g24718(.din(n42740), .dout(n42741));
  jand g24719(.dina(n42388), .dinb(n41995), .dout(n42742));
  jxor g24720(.dina(n42231), .dinb(n42435), .dout(n42743));
  jand g24721(.dina(n42743), .dinb(n42520), .dout(n42744));
  jor  g24722(.dina(n42744), .dinb(n42742), .dout(n42745));
  jand g24723(.dina(n42745), .dinb(n412), .dout(n42746));
  jnot g24724(.din(n42746), .dout(n42747));
  jand g24725(.dina(n42388), .dinb(n42001), .dout(n42748));
  jxor g24726(.dina(n42227), .dinb(n42433), .dout(n42749));
  jand g24727(.dina(n42749), .dinb(n42520), .dout(n42750));
  jor  g24728(.dina(n42750), .dinb(n42748), .dout(n42751));
  jand g24729(.dina(n42751), .dinb(n406), .dout(n42752));
  jnot g24730(.din(n42752), .dout(n42753));
  jand g24731(.dina(n42388), .dinb(n42007), .dout(n42754));
  jxor g24732(.dina(n42223), .dinb(n42431), .dout(n42755));
  jand g24733(.dina(n42755), .dinb(n42520), .dout(n42756));
  jor  g24734(.dina(n42756), .dinb(n42754), .dout(n42757));
  jand g24735(.dina(n42757), .dinb(n405), .dout(n42758));
  jnot g24736(.din(n42758), .dout(n42759));
  jand g24737(.dina(n42388), .dinb(n42013), .dout(n42760));
  jxor g24738(.dina(n42219), .dinb(n42429), .dout(n42761));
  jand g24739(.dina(n42761), .dinb(n42520), .dout(n42762));
  jor  g24740(.dina(n42762), .dinb(n42760), .dout(n42763));
  jand g24741(.dina(n42763), .dinb(n2714), .dout(n42764));
  jnot g24742(.din(n42764), .dout(n42765));
  jand g24743(.dina(n42388), .dinb(n42019), .dout(n42766));
  jxor g24744(.dina(n42215), .dinb(n42427), .dout(n42767));
  jand g24745(.dina(n42767), .dinb(n42520), .dout(n42768));
  jor  g24746(.dina(n42768), .dinb(n42766), .dout(n42769));
  jand g24747(.dina(n42769), .dinb(n2547), .dout(n42770));
  jnot g24748(.din(n42770), .dout(n42771));
  jand g24749(.dina(n42388), .dinb(n42025), .dout(n42772));
  jxor g24750(.dina(n42211), .dinb(n42425), .dout(n42773));
  jand g24751(.dina(n42773), .dinb(n42520), .dout(n42774));
  jor  g24752(.dina(n42774), .dinb(n42772), .dout(n42775));
  jand g24753(.dina(n42775), .dinb(n417), .dout(n42776));
  jnot g24754(.din(n42776), .dout(n42777));
  jand g24755(.dina(n42388), .dinb(n42031), .dout(n42778));
  jxor g24756(.dina(n42207), .dinb(n42423), .dout(n42779));
  jand g24757(.dina(n42779), .dinb(n42520), .dout(n42780));
  jor  g24758(.dina(n42780), .dinb(n42778), .dout(n42781));
  jand g24759(.dina(n42781), .dinb(n416), .dout(n42782));
  jnot g24760(.din(n42782), .dout(n42783));
  jand g24761(.dina(n42388), .dinb(n42037), .dout(n42784));
  jxor g24762(.dina(n42203), .dinb(n42421), .dout(n42785));
  jand g24763(.dina(n42785), .dinb(n42520), .dout(n42786));
  jor  g24764(.dina(n42786), .dinb(n42784), .dout(n42787));
  jand g24765(.dina(n42787), .dinb(n422), .dout(n42788));
  jnot g24766(.din(n42788), .dout(n42789));
  jand g24767(.dina(n42388), .dinb(n42043), .dout(n42790));
  jxor g24768(.dina(n42199), .dinb(n42419), .dout(n42791));
  jand g24769(.dina(n42791), .dinb(n42520), .dout(n42792));
  jor  g24770(.dina(n42792), .dinb(n42790), .dout(n42793));
  jand g24771(.dina(n42793), .dinb(n421), .dout(n42794));
  jnot g24772(.din(n42794), .dout(n42795));
  jand g24773(.dina(n42388), .dinb(n42049), .dout(n42796));
  jxor g24774(.dina(n42195), .dinb(n42417), .dout(n42797));
  jand g24775(.dina(n42797), .dinb(n42520), .dout(n42798));
  jor  g24776(.dina(n42798), .dinb(n42796), .dout(n42799));
  jand g24777(.dina(n42799), .dinb(n433), .dout(n42800));
  jnot g24778(.din(n42800), .dout(n42801));
  jand g24779(.dina(n42388), .dinb(n42055), .dout(n42802));
  jxor g24780(.dina(n42191), .dinb(n42415), .dout(n42803));
  jand g24781(.dina(n42803), .dinb(n42520), .dout(n42804));
  jor  g24782(.dina(n42804), .dinb(n42802), .dout(n42805));
  jand g24783(.dina(n42805), .dinb(n432), .dout(n42806));
  jnot g24784(.din(n42806), .dout(n42807));
  jand g24785(.dina(n42388), .dinb(n42061), .dout(n42808));
  jxor g24786(.dina(n42187), .dinb(n42413), .dout(n42809));
  jand g24787(.dina(n42809), .dinb(n42520), .dout(n42810));
  jor  g24788(.dina(n42810), .dinb(n42808), .dout(n42811));
  jand g24789(.dina(n42811), .dinb(n436), .dout(n42812));
  jnot g24790(.din(n42812), .dout(n42813));
  jand g24791(.dina(n42388), .dinb(n42067), .dout(n42814));
  jxor g24792(.dina(n42183), .dinb(n42411), .dout(n42815));
  jand g24793(.dina(n42815), .dinb(n42520), .dout(n42816));
  jor  g24794(.dina(n42816), .dinb(n42814), .dout(n42817));
  jand g24795(.dina(n42817), .dinb(n435), .dout(n42818));
  jnot g24796(.din(n42818), .dout(n42819));
  jand g24797(.dina(n42388), .dinb(n42073), .dout(n42820));
  jxor g24798(.dina(n42179), .dinb(n42409), .dout(n42821));
  jand g24799(.dina(n42821), .dinb(n42520), .dout(n42822));
  jor  g24800(.dina(n42822), .dinb(n42820), .dout(n42823));
  jand g24801(.dina(n42823), .dinb(n440), .dout(n42824));
  jnot g24802(.din(n42824), .dout(n42825));
  jand g24803(.dina(n42388), .dinb(n42079), .dout(n42826));
  jxor g24804(.dina(n42175), .dinb(n42407), .dout(n42827));
  jand g24805(.dina(n42827), .dinb(n42520), .dout(n42828));
  jor  g24806(.dina(n42828), .dinb(n42826), .dout(n42829));
  jand g24807(.dina(n42829), .dinb(n439), .dout(n42830));
  jnot g24808(.din(n42830), .dout(n42831));
  jand g24809(.dina(n42388), .dinb(n42085), .dout(n42832));
  jxor g24810(.dina(n42171), .dinb(n42405), .dout(n42833));
  jand g24811(.dina(n42833), .dinb(n42520), .dout(n42834));
  jor  g24812(.dina(n42834), .dinb(n42832), .dout(n42835));
  jand g24813(.dina(n42835), .dinb(n325), .dout(n42836));
  jnot g24814(.din(n42836), .dout(n42837));
  jand g24815(.dina(n42388), .dinb(n42091), .dout(n42838));
  jxor g24816(.dina(n42167), .dinb(n42403), .dout(n42839));
  jand g24817(.dina(n42839), .dinb(n42520), .dout(n42840));
  jor  g24818(.dina(n42840), .dinb(n42838), .dout(n42841));
  jand g24819(.dina(n42841), .dinb(n324), .dout(n42842));
  jnot g24820(.din(n42842), .dout(n42843));
  jand g24821(.dina(n42388), .dinb(n42097), .dout(n42844));
  jxor g24822(.dina(n42163), .dinb(n42401), .dout(n42845));
  jand g24823(.dina(n42845), .dinb(n42520), .dout(n42846));
  jor  g24824(.dina(n42846), .dinb(n42844), .dout(n42847));
  jand g24825(.dina(n42847), .dinb(n323), .dout(n42848));
  jnot g24826(.din(n42848), .dout(n42849));
  jand g24827(.dina(n42388), .dinb(n42103), .dout(n42850));
  jxor g24828(.dina(n42159), .dinb(n42399), .dout(n42851));
  jand g24829(.dina(n42851), .dinb(n42520), .dout(n42852));
  jor  g24830(.dina(n42852), .dinb(n42850), .dout(n42853));
  jand g24831(.dina(n42853), .dinb(n335), .dout(n42854));
  jnot g24832(.din(n42854), .dout(n42855));
  jand g24833(.dina(n42388), .dinb(n42109), .dout(n42856));
  jxor g24834(.dina(n42155), .dinb(n42397), .dout(n42857));
  jand g24835(.dina(n42857), .dinb(n42520), .dout(n42858));
  jor  g24836(.dina(n42858), .dinb(n42856), .dout(n42859));
  jand g24837(.dina(n42859), .dinb(n334), .dout(n42860));
  jnot g24838(.din(n42860), .dout(n42861));
  jand g24839(.dina(n42388), .dinb(n42115), .dout(n42862));
  jxor g24840(.dina(n42151), .dinb(n42395), .dout(n42863));
  jand g24841(.dina(n42863), .dinb(n42520), .dout(n42864));
  jor  g24842(.dina(n42864), .dinb(n42862), .dout(n42865));
  jand g24843(.dina(n42865), .dinb(n338), .dout(n42866));
  jnot g24844(.din(n42866), .dout(n42867));
  jand g24845(.dina(n42388), .dinb(n42121), .dout(n42868));
  jxor g24846(.dina(n42147), .dinb(n42393), .dout(n42869));
  jand g24847(.dina(n42869), .dinb(n42520), .dout(n42870));
  jor  g24848(.dina(n42870), .dinb(n42868), .dout(n42871));
  jand g24849(.dina(n42871), .dinb(n337), .dout(n42872));
  jnot g24850(.din(n42872), .dout(n42873));
  jand g24851(.dina(n42388), .dinb(n42127), .dout(n42874));
  jxor g24852(.dina(n42143), .dinb(n42391), .dout(n42875));
  jand g24853(.dina(n42875), .dinb(n42520), .dout(n42876));
  jor  g24854(.dina(n42876), .dinb(n42874), .dout(n42877));
  jand g24855(.dina(n42877), .dinb(n344), .dout(n42878));
  jnot g24856(.din(n42878), .dout(n42879));
  jor  g24857(.dina(n42520), .dinb(n42139), .dout(n42880));
  jxor g24858(.dina(n42389), .dinb(n17812), .dout(n42881));
  jnot g24859(.din(n42881), .dout(n42882));
  jor  g24860(.dina(n42882), .dinb(n42388), .dout(n42883));
  jand g24861(.dina(n42883), .dinb(n42880), .dout(n42884));
  jor  g24862(.dina(n42884), .dinb(b2 ), .dout(n42885));
  jand g24863(.dina(n42520), .dinb(b0 ), .dout(n42886));
  jor  g24864(.dina(n42886), .dinb(n17810), .dout(n42887));
  jor  g24865(.dina(n42388), .dinb(n17812), .dout(n42888));
  jand g24866(.dina(n42888), .dinb(n42887), .dout(n42889));
  jor  g24867(.dina(n42889), .dinb(b1 ), .dout(n42890));
  jnot g24868(.din(n18365), .dout(n42891));
  jxor g24869(.dina(n42889), .dinb(n258), .dout(n42892));
  jor  g24870(.dina(n42892), .dinb(n42891), .dout(n42893));
  jand g24871(.dina(n42893), .dinb(n42890), .dout(n42894));
  jxor g24872(.dina(n42884), .dinb(b2 ), .dout(n42895));
  jnot g24873(.din(n42895), .dout(n42896));
  jor  g24874(.dina(n42896), .dinb(n42894), .dout(n42897));
  jand g24875(.dina(n42897), .dinb(n42885), .dout(n42898));
  jxor g24876(.dina(n42877), .dinb(n344), .dout(n42899));
  jnot g24877(.din(n42899), .dout(n42900));
  jor  g24878(.dina(n42900), .dinb(n42898), .dout(n42901));
  jand g24879(.dina(n42901), .dinb(n42879), .dout(n42902));
  jxor g24880(.dina(n42871), .dinb(n337), .dout(n42903));
  jnot g24881(.din(n42903), .dout(n42904));
  jor  g24882(.dina(n42904), .dinb(n42902), .dout(n42905));
  jand g24883(.dina(n42905), .dinb(n42873), .dout(n42906));
  jxor g24884(.dina(n42865), .dinb(n338), .dout(n42907));
  jnot g24885(.din(n42907), .dout(n42908));
  jor  g24886(.dina(n42908), .dinb(n42906), .dout(n42909));
  jand g24887(.dina(n42909), .dinb(n42867), .dout(n42910));
  jxor g24888(.dina(n42859), .dinb(n334), .dout(n42911));
  jnot g24889(.din(n42911), .dout(n42912));
  jor  g24890(.dina(n42912), .dinb(n42910), .dout(n42913));
  jand g24891(.dina(n42913), .dinb(n42861), .dout(n42914));
  jxor g24892(.dina(n42853), .dinb(n335), .dout(n42915));
  jnot g24893(.din(n42915), .dout(n42916));
  jor  g24894(.dina(n42916), .dinb(n42914), .dout(n42917));
  jand g24895(.dina(n42917), .dinb(n42855), .dout(n42918));
  jxor g24896(.dina(n42847), .dinb(n323), .dout(n42919));
  jnot g24897(.din(n42919), .dout(n42920));
  jor  g24898(.dina(n42920), .dinb(n42918), .dout(n42921));
  jand g24899(.dina(n42921), .dinb(n42849), .dout(n42922));
  jxor g24900(.dina(n42841), .dinb(n324), .dout(n42923));
  jnot g24901(.din(n42923), .dout(n42924));
  jor  g24902(.dina(n42924), .dinb(n42922), .dout(n42925));
  jand g24903(.dina(n42925), .dinb(n42843), .dout(n42926));
  jxor g24904(.dina(n42835), .dinb(n325), .dout(n42927));
  jnot g24905(.din(n42927), .dout(n42928));
  jor  g24906(.dina(n42928), .dinb(n42926), .dout(n42929));
  jand g24907(.dina(n42929), .dinb(n42837), .dout(n42930));
  jxor g24908(.dina(n42829), .dinb(n439), .dout(n42931));
  jnot g24909(.din(n42931), .dout(n42932));
  jor  g24910(.dina(n42932), .dinb(n42930), .dout(n42933));
  jand g24911(.dina(n42933), .dinb(n42831), .dout(n42934));
  jxor g24912(.dina(n42823), .dinb(n440), .dout(n42935));
  jnot g24913(.din(n42935), .dout(n42936));
  jor  g24914(.dina(n42936), .dinb(n42934), .dout(n42937));
  jand g24915(.dina(n42937), .dinb(n42825), .dout(n42938));
  jxor g24916(.dina(n42817), .dinb(n435), .dout(n42939));
  jnot g24917(.din(n42939), .dout(n42940));
  jor  g24918(.dina(n42940), .dinb(n42938), .dout(n42941));
  jand g24919(.dina(n42941), .dinb(n42819), .dout(n42942));
  jxor g24920(.dina(n42811), .dinb(n436), .dout(n42943));
  jnot g24921(.din(n42943), .dout(n42944));
  jor  g24922(.dina(n42944), .dinb(n42942), .dout(n42945));
  jand g24923(.dina(n42945), .dinb(n42813), .dout(n42946));
  jxor g24924(.dina(n42805), .dinb(n432), .dout(n42947));
  jnot g24925(.din(n42947), .dout(n42948));
  jor  g24926(.dina(n42948), .dinb(n42946), .dout(n42949));
  jand g24927(.dina(n42949), .dinb(n42807), .dout(n42950));
  jxor g24928(.dina(n42799), .dinb(n433), .dout(n42951));
  jnot g24929(.din(n42951), .dout(n42952));
  jor  g24930(.dina(n42952), .dinb(n42950), .dout(n42953));
  jand g24931(.dina(n42953), .dinb(n42801), .dout(n42954));
  jxor g24932(.dina(n42793), .dinb(n421), .dout(n42955));
  jnot g24933(.din(n42955), .dout(n42956));
  jor  g24934(.dina(n42956), .dinb(n42954), .dout(n42957));
  jand g24935(.dina(n42957), .dinb(n42795), .dout(n42958));
  jxor g24936(.dina(n42787), .dinb(n422), .dout(n42959));
  jnot g24937(.din(n42959), .dout(n42960));
  jor  g24938(.dina(n42960), .dinb(n42958), .dout(n42961));
  jand g24939(.dina(n42961), .dinb(n42789), .dout(n42962));
  jxor g24940(.dina(n42781), .dinb(n416), .dout(n42963));
  jnot g24941(.din(n42963), .dout(n42964));
  jor  g24942(.dina(n42964), .dinb(n42962), .dout(n42965));
  jand g24943(.dina(n42965), .dinb(n42783), .dout(n42966));
  jxor g24944(.dina(n42775), .dinb(n417), .dout(n42967));
  jnot g24945(.din(n42967), .dout(n42968));
  jor  g24946(.dina(n42968), .dinb(n42966), .dout(n42969));
  jand g24947(.dina(n42969), .dinb(n42777), .dout(n42970));
  jxor g24948(.dina(n42769), .dinb(n2547), .dout(n42971));
  jnot g24949(.din(n42971), .dout(n42972));
  jor  g24950(.dina(n42972), .dinb(n42970), .dout(n42973));
  jand g24951(.dina(n42973), .dinb(n42771), .dout(n42974));
  jxor g24952(.dina(n42763), .dinb(n2714), .dout(n42975));
  jnot g24953(.din(n42975), .dout(n42976));
  jor  g24954(.dina(n42976), .dinb(n42974), .dout(n42977));
  jand g24955(.dina(n42977), .dinb(n42765), .dout(n42978));
  jxor g24956(.dina(n42757), .dinb(n405), .dout(n42979));
  jnot g24957(.din(n42979), .dout(n42980));
  jor  g24958(.dina(n42980), .dinb(n42978), .dout(n42981));
  jand g24959(.dina(n42981), .dinb(n42759), .dout(n42982));
  jxor g24960(.dina(n42751), .dinb(n406), .dout(n42983));
  jnot g24961(.din(n42983), .dout(n42984));
  jor  g24962(.dina(n42984), .dinb(n42982), .dout(n42985));
  jand g24963(.dina(n42985), .dinb(n42753), .dout(n42986));
  jxor g24964(.dina(n42745), .dinb(n412), .dout(n42987));
  jnot g24965(.din(n42987), .dout(n42988));
  jor  g24966(.dina(n42988), .dinb(n42986), .dout(n42989));
  jand g24967(.dina(n42989), .dinb(n42747), .dout(n42990));
  jxor g24968(.dina(n42739), .dinb(n413), .dout(n42991));
  jnot g24969(.din(n42991), .dout(n42992));
  jor  g24970(.dina(n42992), .dinb(n42990), .dout(n42993));
  jand g24971(.dina(n42993), .dinb(n42741), .dout(n42994));
  jxor g24972(.dina(n42733), .dinb(n409), .dout(n42995));
  jnot g24973(.din(n42995), .dout(n42996));
  jor  g24974(.dina(n42996), .dinb(n42994), .dout(n42997));
  jand g24975(.dina(n42997), .dinb(n42735), .dout(n42998));
  jxor g24976(.dina(n42727), .dinb(n410), .dout(n42999));
  jnot g24977(.din(n42999), .dout(n43000));
  jor  g24978(.dina(n43000), .dinb(n42998), .dout(n43001));
  jand g24979(.dina(n43001), .dinb(n42729), .dout(n43002));
  jxor g24980(.dina(n42721), .dinb(n426), .dout(n43003));
  jnot g24981(.din(n43003), .dout(n43004));
  jor  g24982(.dina(n43004), .dinb(n43002), .dout(n43005));
  jand g24983(.dina(n43005), .dinb(n42723), .dout(n43006));
  jxor g24984(.dina(n42715), .dinb(n427), .dout(n43007));
  jnot g24985(.din(n43007), .dout(n43008));
  jor  g24986(.dina(n43008), .dinb(n43006), .dout(n43009));
  jand g24987(.dina(n43009), .dinb(n42717), .dout(n43010));
  jxor g24988(.dina(n42709), .dinb(n424), .dout(n43011));
  jnot g24989(.din(n43011), .dout(n43012));
  jor  g24990(.dina(n43012), .dinb(n43010), .dout(n43013));
  jand g24991(.dina(n43013), .dinb(n42711), .dout(n43014));
  jxor g24992(.dina(n42703), .dinb(n300), .dout(n43015));
  jnot g24993(.din(n43015), .dout(n43016));
  jor  g24994(.dina(n43016), .dinb(n43014), .dout(n43017));
  jand g24995(.dina(n43017), .dinb(n42705), .dout(n43018));
  jxor g24996(.dina(n42697), .dinb(n297), .dout(n43019));
  jnot g24997(.din(n43019), .dout(n43020));
  jor  g24998(.dina(n43020), .dinb(n43018), .dout(n43021));
  jand g24999(.dina(n43021), .dinb(n42699), .dout(n43022));
  jxor g25000(.dina(n42691), .dinb(n298), .dout(n43023));
  jnot g25001(.din(n43023), .dout(n43024));
  jor  g25002(.dina(n43024), .dinb(n43022), .dout(n43025));
  jand g25003(.dina(n43025), .dinb(n42693), .dout(n43026));
  jxor g25004(.dina(n42685), .dinb(n301), .dout(n43027));
  jnot g25005(.din(n43027), .dout(n43028));
  jor  g25006(.dina(n43028), .dinb(n43026), .dout(n43029));
  jand g25007(.dina(n43029), .dinb(n42687), .dout(n43030));
  jxor g25008(.dina(n42679), .dinb(n293), .dout(n43031));
  jnot g25009(.din(n43031), .dout(n43032));
  jor  g25010(.dina(n43032), .dinb(n43030), .dout(n43033));
  jand g25011(.dina(n43033), .dinb(n42681), .dout(n43034));
  jxor g25012(.dina(n42673), .dinb(n294), .dout(n43035));
  jnot g25013(.din(n43035), .dout(n43036));
  jor  g25014(.dina(n43036), .dinb(n43034), .dout(n43037));
  jand g25015(.dina(n43037), .dinb(n42675), .dout(n43038));
  jxor g25016(.dina(n42667), .dinb(n290), .dout(n43039));
  jnot g25017(.din(n43039), .dout(n43040));
  jor  g25018(.dina(n43040), .dinb(n43038), .dout(n43041));
  jand g25019(.dina(n43041), .dinb(n42669), .dout(n43042));
  jxor g25020(.dina(n42661), .dinb(n291), .dout(n43043));
  jnot g25021(.din(n43043), .dout(n43044));
  jor  g25022(.dina(n43044), .dinb(n43042), .dout(n43045));
  jand g25023(.dina(n43045), .dinb(n42663), .dout(n43046));
  jxor g25024(.dina(n42655), .dinb(n284), .dout(n43047));
  jnot g25025(.din(n43047), .dout(n43048));
  jor  g25026(.dina(n43048), .dinb(n43046), .dout(n43049));
  jand g25027(.dina(n43049), .dinb(n42657), .dout(n43050));
  jxor g25028(.dina(n42649), .dinb(n285), .dout(n43051));
  jnot g25029(.din(n43051), .dout(n43052));
  jor  g25030(.dina(n43052), .dinb(n43050), .dout(n43053));
  jand g25031(.dina(n43053), .dinb(n42651), .dout(n43054));
  jxor g25032(.dina(n42643), .dinb(n281), .dout(n43055));
  jnot g25033(.din(n43055), .dout(n43056));
  jor  g25034(.dina(n43056), .dinb(n43054), .dout(n43057));
  jand g25035(.dina(n43057), .dinb(n42645), .dout(n43058));
  jxor g25036(.dina(n42637), .dinb(n282), .dout(n43059));
  jnot g25037(.din(n43059), .dout(n43060));
  jor  g25038(.dina(n43060), .dinb(n43058), .dout(n43061));
  jand g25039(.dina(n43061), .dinb(n42639), .dout(n43062));
  jxor g25040(.dina(n42631), .dinb(n397), .dout(n43063));
  jnot g25041(.din(n43063), .dout(n43064));
  jor  g25042(.dina(n43064), .dinb(n43062), .dout(n43065));
  jand g25043(.dina(n43065), .dinb(n42633), .dout(n43066));
  jxor g25044(.dina(n42625), .dinb(n513), .dout(n43067));
  jnot g25045(.din(n43067), .dout(n43068));
  jor  g25046(.dina(n43068), .dinb(n43066), .dout(n43069));
  jand g25047(.dina(n43069), .dinb(n42627), .dout(n43070));
  jxor g25048(.dina(n42619), .dinb(n514), .dout(n43071));
  jnot g25049(.din(n43071), .dout(n43072));
  jor  g25050(.dina(n43072), .dinb(n43070), .dout(n43073));
  jand g25051(.dina(n43073), .dinb(n42621), .dout(n43074));
  jxor g25052(.dina(n42613), .dinb(n510), .dout(n43075));
  jnot g25053(.din(n43075), .dout(n43076));
  jor  g25054(.dina(n43076), .dinb(n43074), .dout(n43077));
  jand g25055(.dina(n43077), .dinb(n42615), .dout(n43078));
  jxor g25056(.dina(n42607), .dinb(n396), .dout(n43079));
  jnot g25057(.din(n43079), .dout(n43080));
  jor  g25058(.dina(n43080), .dinb(n43078), .dout(n43081));
  jand g25059(.dina(n43081), .dinb(n42609), .dout(n43082));
  jxor g25060(.dina(n42601), .dinb(n383), .dout(n43083));
  jnot g25061(.din(n43083), .dout(n43084));
  jor  g25062(.dina(n43084), .dinb(n43082), .dout(n43085));
  jand g25063(.dina(n43085), .dinb(n42603), .dout(n43086));
  jxor g25064(.dina(n42595), .dinb(n12211), .dout(n43087));
  jnot g25065(.din(n43087), .dout(n43088));
  jor  g25066(.dina(n43088), .dinb(n43086), .dout(n43089));
  jand g25067(.dina(n43089), .dinb(n42597), .dout(n43090));
  jxor g25068(.dina(n42589), .dinb(n12214), .dout(n43091));
  jnot g25069(.din(n43091), .dout(n43092));
  jor  g25070(.dina(n43092), .dinb(n43090), .dout(n43093));
  jand g25071(.dina(n43093), .dinb(n42591), .dout(n43094));
  jxor g25072(.dina(n42583), .dinb(n384), .dout(n43095));
  jnot g25073(.din(n43095), .dout(n43096));
  jor  g25074(.dina(n43096), .dinb(n43094), .dout(n43097));
  jand g25075(.dina(n43097), .dinb(n42585), .dout(n43098));
  jxor g25076(.dina(n42577), .dinb(n374), .dout(n43099));
  jnot g25077(.din(n43099), .dout(n43100));
  jor  g25078(.dina(n43100), .dinb(n43098), .dout(n43101));
  jand g25079(.dina(n43101), .dinb(n42579), .dout(n43102));
  jxor g25080(.dina(n42571), .dinb(n376), .dout(n43103));
  jnot g25081(.din(n43103), .dout(n43104));
  jor  g25082(.dina(n43104), .dinb(n43102), .dout(n43105));
  jand g25083(.dina(n43105), .dinb(n42573), .dout(n43106));
  jxor g25084(.dina(n42565), .dinb(n377), .dout(n43107));
  jnot g25085(.din(n43107), .dout(n43108));
  jor  g25086(.dina(n43108), .dinb(n43106), .dout(n43109));
  jand g25087(.dina(n43109), .dinb(n42567), .dout(n43110));
  jxor g25088(.dina(n42559), .dinb(n375), .dout(n43111));
  jnot g25089(.din(n43111), .dout(n43112));
  jor  g25090(.dina(n43112), .dinb(n43110), .dout(n43113));
  jand g25091(.dina(n43113), .dinb(n42561), .dout(n43114));
  jxor g25092(.dina(n42553), .dinb(n362), .dout(n43115));
  jnot g25093(.din(n43115), .dout(n43116));
  jor  g25094(.dina(n43116), .dinb(n43114), .dout(n43117));
  jand g25095(.dina(n43117), .dinb(n42555), .dout(n43118));
  jxor g25096(.dina(n42547), .dinb(n363), .dout(n43119));
  jnot g25097(.din(n43119), .dout(n43120));
  jor  g25098(.dina(n43120), .dinb(n43118), .dout(n43121));
  jand g25099(.dina(n43121), .dinb(n42549), .dout(n43122));
  jxor g25100(.dina(n42541), .dinb(n365), .dout(n43123));
  jnot g25101(.din(n43123), .dout(n43124));
  jor  g25102(.dina(n43124), .dinb(n43122), .dout(n43125));
  jand g25103(.dina(n43125), .dinb(n42543), .dout(n43126));
  jxor g25104(.dina(n42535), .dinb(n366), .dout(n43127));
  jnot g25105(.din(n43127), .dout(n43128));
  jor  g25106(.dina(n43128), .dinb(n43126), .dout(n43129));
  jand g25107(.dina(n43129), .dinb(n42537), .dout(n43130));
  jxor g25108(.dina(n42529), .dinb(n256), .dout(n43131));
  jnot g25109(.din(n43131), .dout(n43132));
  jor  g25110(.dina(n43132), .dinb(n43130), .dout(n43133));
  jand g25111(.dina(n43133), .dinb(n42531), .dout(n43134));
  jxor g25112(.dina(n42523), .dinb(n367), .dout(n43135));
  jnot g25113(.din(n43135), .dout(n43136));
  jor  g25114(.dina(n43136), .dinb(n43134), .dout(n43137));
  jand g25115(.dina(n43137), .dinb(n42525), .dout(n43138));
  jand g25116(.dina(n43138), .dinb(n42516), .dout(n43139));
  jor  g25117(.dina(n43139), .dinb(n41766), .dout(n43140));
  jor  g25118(.dina(n43140), .dinb(n18364), .dout(n43141));
  jand g25119(.dina(n43141), .dinb(a0 ), .dout(n43142));
  jnot g25120(.din(n41766), .dout(n43143));
  jnot g25121(.din(n42885), .dout(n43144));
  jnot g25122(.din(n42890), .dout(n43145));
  jxor g25123(.dina(n42889), .dinb(b1 ), .dout(n43146));
  jand g25124(.dina(n43146), .dinb(n18365), .dout(n43147));
  jor  g25125(.dina(n43147), .dinb(n43145), .dout(n43148));
  jand g25126(.dina(n42895), .dinb(n43148), .dout(n43149));
  jor  g25127(.dina(n43149), .dinb(n43144), .dout(n43150));
  jand g25128(.dina(n42899), .dinb(n43150), .dout(n43151));
  jor  g25129(.dina(n43151), .dinb(n42878), .dout(n43152));
  jand g25130(.dina(n42903), .dinb(n43152), .dout(n43153));
  jor  g25131(.dina(n43153), .dinb(n42872), .dout(n43154));
  jand g25132(.dina(n42907), .dinb(n43154), .dout(n43155));
  jor  g25133(.dina(n43155), .dinb(n42866), .dout(n43156));
  jand g25134(.dina(n42911), .dinb(n43156), .dout(n43157));
  jor  g25135(.dina(n43157), .dinb(n42860), .dout(n43158));
  jand g25136(.dina(n42915), .dinb(n43158), .dout(n43159));
  jor  g25137(.dina(n43159), .dinb(n42854), .dout(n43160));
  jand g25138(.dina(n42919), .dinb(n43160), .dout(n43161));
  jor  g25139(.dina(n43161), .dinb(n42848), .dout(n43162));
  jand g25140(.dina(n42923), .dinb(n43162), .dout(n43163));
  jor  g25141(.dina(n43163), .dinb(n42842), .dout(n43164));
  jand g25142(.dina(n42927), .dinb(n43164), .dout(n43165));
  jor  g25143(.dina(n43165), .dinb(n42836), .dout(n43166));
  jand g25144(.dina(n42931), .dinb(n43166), .dout(n43167));
  jor  g25145(.dina(n43167), .dinb(n42830), .dout(n43168));
  jand g25146(.dina(n42935), .dinb(n43168), .dout(n43169));
  jor  g25147(.dina(n43169), .dinb(n42824), .dout(n43170));
  jand g25148(.dina(n42939), .dinb(n43170), .dout(n43171));
  jor  g25149(.dina(n43171), .dinb(n42818), .dout(n43172));
  jand g25150(.dina(n42943), .dinb(n43172), .dout(n43173));
  jor  g25151(.dina(n43173), .dinb(n42812), .dout(n43174));
  jand g25152(.dina(n42947), .dinb(n43174), .dout(n43175));
  jor  g25153(.dina(n43175), .dinb(n42806), .dout(n43176));
  jand g25154(.dina(n42951), .dinb(n43176), .dout(n43177));
  jor  g25155(.dina(n43177), .dinb(n42800), .dout(n43178));
  jand g25156(.dina(n42955), .dinb(n43178), .dout(n43179));
  jor  g25157(.dina(n43179), .dinb(n42794), .dout(n43180));
  jand g25158(.dina(n42959), .dinb(n43180), .dout(n43181));
  jor  g25159(.dina(n43181), .dinb(n42788), .dout(n43182));
  jand g25160(.dina(n42963), .dinb(n43182), .dout(n43183));
  jor  g25161(.dina(n43183), .dinb(n42782), .dout(n43184));
  jand g25162(.dina(n42967), .dinb(n43184), .dout(n43185));
  jor  g25163(.dina(n43185), .dinb(n42776), .dout(n43186));
  jand g25164(.dina(n42971), .dinb(n43186), .dout(n43187));
  jor  g25165(.dina(n43187), .dinb(n42770), .dout(n43188));
  jand g25166(.dina(n42975), .dinb(n43188), .dout(n43189));
  jor  g25167(.dina(n43189), .dinb(n42764), .dout(n43190));
  jand g25168(.dina(n42979), .dinb(n43190), .dout(n43191));
  jor  g25169(.dina(n43191), .dinb(n42758), .dout(n43192));
  jand g25170(.dina(n42983), .dinb(n43192), .dout(n43193));
  jor  g25171(.dina(n43193), .dinb(n42752), .dout(n43194));
  jand g25172(.dina(n42987), .dinb(n43194), .dout(n43195));
  jor  g25173(.dina(n43195), .dinb(n42746), .dout(n43196));
  jand g25174(.dina(n42991), .dinb(n43196), .dout(n43197));
  jor  g25175(.dina(n43197), .dinb(n42740), .dout(n43198));
  jand g25176(.dina(n42995), .dinb(n43198), .dout(n43199));
  jor  g25177(.dina(n43199), .dinb(n42734), .dout(n43200));
  jand g25178(.dina(n42999), .dinb(n43200), .dout(n43201));
  jor  g25179(.dina(n43201), .dinb(n42728), .dout(n43202));
  jand g25180(.dina(n43003), .dinb(n43202), .dout(n43203));
  jor  g25181(.dina(n43203), .dinb(n42722), .dout(n43204));
  jand g25182(.dina(n43007), .dinb(n43204), .dout(n43205));
  jor  g25183(.dina(n43205), .dinb(n42716), .dout(n43206));
  jand g25184(.dina(n43011), .dinb(n43206), .dout(n43207));
  jor  g25185(.dina(n43207), .dinb(n42710), .dout(n43208));
  jand g25186(.dina(n43015), .dinb(n43208), .dout(n43209));
  jor  g25187(.dina(n43209), .dinb(n42704), .dout(n43210));
  jand g25188(.dina(n43019), .dinb(n43210), .dout(n43211));
  jor  g25189(.dina(n43211), .dinb(n42698), .dout(n43212));
  jand g25190(.dina(n43023), .dinb(n43212), .dout(n43213));
  jor  g25191(.dina(n43213), .dinb(n42692), .dout(n43214));
  jand g25192(.dina(n43027), .dinb(n43214), .dout(n43215));
  jor  g25193(.dina(n43215), .dinb(n42686), .dout(n43216));
  jand g25194(.dina(n43031), .dinb(n43216), .dout(n43217));
  jor  g25195(.dina(n43217), .dinb(n42680), .dout(n43218));
  jand g25196(.dina(n43035), .dinb(n43218), .dout(n43219));
  jor  g25197(.dina(n43219), .dinb(n42674), .dout(n43220));
  jand g25198(.dina(n43039), .dinb(n43220), .dout(n43221));
  jor  g25199(.dina(n43221), .dinb(n42668), .dout(n43222));
  jand g25200(.dina(n43043), .dinb(n43222), .dout(n43223));
  jor  g25201(.dina(n43223), .dinb(n42662), .dout(n43224));
  jand g25202(.dina(n43047), .dinb(n43224), .dout(n43225));
  jor  g25203(.dina(n43225), .dinb(n42656), .dout(n43226));
  jand g25204(.dina(n43051), .dinb(n43226), .dout(n43227));
  jor  g25205(.dina(n43227), .dinb(n42650), .dout(n43228));
  jand g25206(.dina(n43055), .dinb(n43228), .dout(n43229));
  jor  g25207(.dina(n43229), .dinb(n42644), .dout(n43230));
  jand g25208(.dina(n43059), .dinb(n43230), .dout(n43231));
  jor  g25209(.dina(n43231), .dinb(n42638), .dout(n43232));
  jand g25210(.dina(n43063), .dinb(n43232), .dout(n43233));
  jor  g25211(.dina(n43233), .dinb(n42632), .dout(n43234));
  jand g25212(.dina(n43067), .dinb(n43234), .dout(n43235));
  jor  g25213(.dina(n43235), .dinb(n42626), .dout(n43236));
  jand g25214(.dina(n43071), .dinb(n43236), .dout(n43237));
  jor  g25215(.dina(n43237), .dinb(n42620), .dout(n43238));
  jand g25216(.dina(n43075), .dinb(n43238), .dout(n43239));
  jor  g25217(.dina(n43239), .dinb(n42614), .dout(n43240));
  jand g25218(.dina(n43079), .dinb(n43240), .dout(n43241));
  jor  g25219(.dina(n43241), .dinb(n42608), .dout(n43242));
  jand g25220(.dina(n43083), .dinb(n43242), .dout(n43243));
  jor  g25221(.dina(n43243), .dinb(n42602), .dout(n43244));
  jand g25222(.dina(n43087), .dinb(n43244), .dout(n43245));
  jor  g25223(.dina(n43245), .dinb(n42596), .dout(n43246));
  jand g25224(.dina(n43091), .dinb(n43246), .dout(n43247));
  jor  g25225(.dina(n43247), .dinb(n42590), .dout(n43248));
  jand g25226(.dina(n43095), .dinb(n43248), .dout(n43249));
  jor  g25227(.dina(n43249), .dinb(n42584), .dout(n43250));
  jand g25228(.dina(n43099), .dinb(n43250), .dout(n43251));
  jor  g25229(.dina(n43251), .dinb(n42578), .dout(n43252));
  jand g25230(.dina(n43103), .dinb(n43252), .dout(n43253));
  jor  g25231(.dina(n43253), .dinb(n42572), .dout(n43254));
  jand g25232(.dina(n43107), .dinb(n43254), .dout(n43255));
  jor  g25233(.dina(n43255), .dinb(n42566), .dout(n43256));
  jand g25234(.dina(n43111), .dinb(n43256), .dout(n43257));
  jor  g25235(.dina(n43257), .dinb(n42560), .dout(n43258));
  jand g25236(.dina(n43115), .dinb(n43258), .dout(n43259));
  jor  g25237(.dina(n43259), .dinb(n42554), .dout(n43260));
  jand g25238(.dina(n43119), .dinb(n43260), .dout(n43261));
  jor  g25239(.dina(n43261), .dinb(n42548), .dout(n43262));
  jand g25240(.dina(n43123), .dinb(n43262), .dout(n43263));
  jor  g25241(.dina(n43263), .dinb(n42542), .dout(n43264));
  jand g25242(.dina(n43127), .dinb(n43264), .dout(n43265));
  jor  g25243(.dina(n43265), .dinb(n42536), .dout(n43266));
  jand g25244(.dina(n43131), .dinb(n43266), .dout(n43267));
  jor  g25245(.dina(n43267), .dinb(n42530), .dout(n43268));
  jand g25246(.dina(n43135), .dinb(n43268), .dout(n43269));
  jor  g25247(.dina(n43269), .dinb(n42524), .dout(n43270));
  jor  g25248(.dina(n43270), .dinb(n42515), .dout(n43271));
  jand g25249(.dina(n43271), .dinb(n43143), .dout(n43272));
  jand g25250(.dina(n43272), .dinb(n42891), .dout(n43273));
  jor  g25251(.dina(n43273), .dinb(n43142), .dout(remainder0 ));
  jnot g25252(.din(n42889), .dout(n43275));
  jand g25253(.dina(n43140), .dinb(n43275), .dout(n43276));
  jxor g25254(.dina(n43146), .dinb(n18365), .dout(n43277));
  jand g25255(.dina(n43277), .dinb(n43272), .dout(n43278));
  jor  g25256(.dina(n43278), .dinb(n43276), .dout(remainder1 ));
  jnot g25257(.din(n42884), .dout(n43280));
  jand g25258(.dina(n43140), .dinb(n43280), .dout(n43281));
  jxor g25259(.dina(n42895), .dinb(n43148), .dout(n43282));
  jand g25260(.dina(n43282), .dinb(n43272), .dout(n43283));
  jor  g25261(.dina(n43283), .dinb(n43281), .dout(remainder2 ));
  jand g25262(.dina(n43140), .dinb(n42877), .dout(n43285));
  jxor g25263(.dina(n42899), .dinb(n43150), .dout(n43286));
  jand g25264(.dina(n43286), .dinb(n43272), .dout(n43287));
  jor  g25265(.dina(n43287), .dinb(n43285), .dout(remainder3 ));
  jand g25266(.dina(n43140), .dinb(n42871), .dout(n43289));
  jxor g25267(.dina(n42903), .dinb(n43152), .dout(n43290));
  jand g25268(.dina(n43290), .dinb(n43272), .dout(n43291));
  jor  g25269(.dina(n43291), .dinb(n43289), .dout(remainder4 ));
  jand g25270(.dina(n43140), .dinb(n42865), .dout(n43293));
  jxor g25271(.dina(n42907), .dinb(n43154), .dout(n43294));
  jand g25272(.dina(n43294), .dinb(n43272), .dout(n43295));
  jor  g25273(.dina(n43295), .dinb(n43293), .dout(remainder5 ));
  jand g25274(.dina(n43140), .dinb(n42859), .dout(n43297));
  jxor g25275(.dina(n42911), .dinb(n43156), .dout(n43298));
  jand g25276(.dina(n43298), .dinb(n43272), .dout(n43299));
  jor  g25277(.dina(n43299), .dinb(n43297), .dout(remainder6 ));
  jand g25278(.dina(n43140), .dinb(n42853), .dout(n43301));
  jxor g25279(.dina(n42915), .dinb(n43158), .dout(n43302));
  jand g25280(.dina(n43302), .dinb(n43272), .dout(n43303));
  jor  g25281(.dina(n43303), .dinb(n43301), .dout(remainder7 ));
  jand g25282(.dina(n43140), .dinb(n42847), .dout(n43305));
  jxor g25283(.dina(n42919), .dinb(n43160), .dout(n43306));
  jand g25284(.dina(n43306), .dinb(n43272), .dout(n43307));
  jor  g25285(.dina(n43307), .dinb(n43305), .dout(remainder8 ));
  jand g25286(.dina(n43140), .dinb(n42841), .dout(n43309));
  jxor g25287(.dina(n42923), .dinb(n43162), .dout(n43310));
  jand g25288(.dina(n43310), .dinb(n43272), .dout(n43311));
  jor  g25289(.dina(n43311), .dinb(n43309), .dout(remainder9 ));
  jand g25290(.dina(n43140), .dinb(n42835), .dout(n43313));
  jxor g25291(.dina(n42927), .dinb(n43164), .dout(n43314));
  jand g25292(.dina(n43314), .dinb(n43272), .dout(n43315));
  jor  g25293(.dina(n43315), .dinb(n43313), .dout(remainder10 ));
  jand g25294(.dina(n43140), .dinb(n42829), .dout(n43317));
  jxor g25295(.dina(n42931), .dinb(n43166), .dout(n43318));
  jand g25296(.dina(n43318), .dinb(n43272), .dout(n43319));
  jor  g25297(.dina(n43319), .dinb(n43317), .dout(remainder11 ));
  jand g25298(.dina(n43140), .dinb(n42823), .dout(n43321));
  jxor g25299(.dina(n42935), .dinb(n43168), .dout(n43322));
  jand g25300(.dina(n43322), .dinb(n43272), .dout(n43323));
  jor  g25301(.dina(n43323), .dinb(n43321), .dout(remainder12 ));
  jand g25302(.dina(n43140), .dinb(n42817), .dout(n43325));
  jxor g25303(.dina(n42939), .dinb(n43170), .dout(n43326));
  jand g25304(.dina(n43326), .dinb(n43272), .dout(n43327));
  jor  g25305(.dina(n43327), .dinb(n43325), .dout(remainder13 ));
  jand g25306(.dina(n43140), .dinb(n42811), .dout(n43329));
  jxor g25307(.dina(n42943), .dinb(n43172), .dout(n43330));
  jand g25308(.dina(n43330), .dinb(n43272), .dout(n43331));
  jor  g25309(.dina(n43331), .dinb(n43329), .dout(remainder14 ));
  jand g25310(.dina(n43140), .dinb(n42805), .dout(n43333));
  jxor g25311(.dina(n42947), .dinb(n43174), .dout(n43334));
  jand g25312(.dina(n43334), .dinb(n43272), .dout(n43335));
  jor  g25313(.dina(n43335), .dinb(n43333), .dout(remainder15 ));
  jand g25314(.dina(n43140), .dinb(n42799), .dout(n43337));
  jxor g25315(.dina(n42951), .dinb(n43176), .dout(n43338));
  jand g25316(.dina(n43338), .dinb(n43272), .dout(n43339));
  jor  g25317(.dina(n43339), .dinb(n43337), .dout(remainder16 ));
  jand g25318(.dina(n43140), .dinb(n42793), .dout(n43341));
  jxor g25319(.dina(n42955), .dinb(n43178), .dout(n43342));
  jand g25320(.dina(n43342), .dinb(n43272), .dout(n43343));
  jor  g25321(.dina(n43343), .dinb(n43341), .dout(remainder17 ));
  jand g25322(.dina(n43140), .dinb(n42787), .dout(n43345));
  jxor g25323(.dina(n42959), .dinb(n43180), .dout(n43346));
  jand g25324(.dina(n43346), .dinb(n43272), .dout(n43347));
  jor  g25325(.dina(n43347), .dinb(n43345), .dout(remainder18 ));
  jand g25326(.dina(n43140), .dinb(n42781), .dout(n43349));
  jxor g25327(.dina(n42963), .dinb(n43182), .dout(n43350));
  jand g25328(.dina(n43350), .dinb(n43272), .dout(n43351));
  jor  g25329(.dina(n43351), .dinb(n43349), .dout(remainder19 ));
  jand g25330(.dina(n43140), .dinb(n42775), .dout(n43353));
  jxor g25331(.dina(n42967), .dinb(n43184), .dout(n43354));
  jand g25332(.dina(n43354), .dinb(n43272), .dout(n43355));
  jor  g25333(.dina(n43355), .dinb(n43353), .dout(remainder20 ));
  jand g25334(.dina(n43140), .dinb(n42769), .dout(n43357));
  jxor g25335(.dina(n42971), .dinb(n43186), .dout(n43358));
  jand g25336(.dina(n43358), .dinb(n43272), .dout(n43359));
  jor  g25337(.dina(n43359), .dinb(n43357), .dout(remainder21 ));
  jand g25338(.dina(n43140), .dinb(n42763), .dout(n43361));
  jxor g25339(.dina(n42975), .dinb(n43188), .dout(n43362));
  jand g25340(.dina(n43362), .dinb(n43272), .dout(n43363));
  jor  g25341(.dina(n43363), .dinb(n43361), .dout(remainder22 ));
  jand g25342(.dina(n43140), .dinb(n42757), .dout(n43365));
  jxor g25343(.dina(n42979), .dinb(n43190), .dout(n43366));
  jand g25344(.dina(n43366), .dinb(n43272), .dout(n43367));
  jor  g25345(.dina(n43367), .dinb(n43365), .dout(remainder23 ));
  jand g25346(.dina(n43140), .dinb(n42751), .dout(n43369));
  jxor g25347(.dina(n42983), .dinb(n43192), .dout(n43370));
  jand g25348(.dina(n43370), .dinb(n43272), .dout(n43371));
  jor  g25349(.dina(n43371), .dinb(n43369), .dout(remainder24 ));
  jand g25350(.dina(n43140), .dinb(n42745), .dout(n43373));
  jxor g25351(.dina(n42987), .dinb(n43194), .dout(n43374));
  jand g25352(.dina(n43374), .dinb(n43272), .dout(n43375));
  jor  g25353(.dina(n43375), .dinb(n43373), .dout(remainder25 ));
  jand g25354(.dina(n43140), .dinb(n42739), .dout(n43377));
  jxor g25355(.dina(n42991), .dinb(n43196), .dout(n43378));
  jand g25356(.dina(n43378), .dinb(n43272), .dout(n43379));
  jor  g25357(.dina(n43379), .dinb(n43377), .dout(remainder26 ));
  jand g25358(.dina(n43140), .dinb(n42733), .dout(n43381));
  jxor g25359(.dina(n42995), .dinb(n43198), .dout(n43382));
  jand g25360(.dina(n43382), .dinb(n43272), .dout(n43383));
  jor  g25361(.dina(n43383), .dinb(n43381), .dout(remainder27 ));
  jand g25362(.dina(n43140), .dinb(n42727), .dout(n43385));
  jxor g25363(.dina(n42999), .dinb(n43200), .dout(n43386));
  jand g25364(.dina(n43386), .dinb(n43272), .dout(n43387));
  jor  g25365(.dina(n43387), .dinb(n43385), .dout(remainder28 ));
  jand g25366(.dina(n43140), .dinb(n42721), .dout(n43389));
  jxor g25367(.dina(n43003), .dinb(n43202), .dout(n43390));
  jand g25368(.dina(n43390), .dinb(n43272), .dout(n43391));
  jor  g25369(.dina(n43391), .dinb(n43389), .dout(remainder29 ));
  jand g25370(.dina(n43140), .dinb(n42715), .dout(n43393));
  jxor g25371(.dina(n43007), .dinb(n43204), .dout(n43394));
  jand g25372(.dina(n43394), .dinb(n43272), .dout(n43395));
  jor  g25373(.dina(n43395), .dinb(n43393), .dout(remainder30 ));
  jand g25374(.dina(n43140), .dinb(n42709), .dout(n43397));
  jxor g25375(.dina(n43011), .dinb(n43206), .dout(n43398));
  jand g25376(.dina(n43398), .dinb(n43272), .dout(n43399));
  jor  g25377(.dina(n43399), .dinb(n43397), .dout(remainder31 ));
  jand g25378(.dina(n43140), .dinb(n42703), .dout(n43401));
  jxor g25379(.dina(n43015), .dinb(n43208), .dout(n43402));
  jand g25380(.dina(n43402), .dinb(n43272), .dout(n43403));
  jor  g25381(.dina(n43403), .dinb(n43401), .dout(remainder32 ));
  jand g25382(.dina(n43140), .dinb(n42697), .dout(n43405));
  jxor g25383(.dina(n43019), .dinb(n43210), .dout(n43406));
  jand g25384(.dina(n43406), .dinb(n43272), .dout(n43407));
  jor  g25385(.dina(n43407), .dinb(n43405), .dout(remainder33 ));
  jand g25386(.dina(n43140), .dinb(n42691), .dout(n43409));
  jxor g25387(.dina(n43023), .dinb(n43212), .dout(n43410));
  jand g25388(.dina(n43410), .dinb(n43272), .dout(n43411));
  jor  g25389(.dina(n43411), .dinb(n43409), .dout(remainder34 ));
  jand g25390(.dina(n43140), .dinb(n42685), .dout(n43413));
  jxor g25391(.dina(n43027), .dinb(n43214), .dout(n43414));
  jand g25392(.dina(n43414), .dinb(n43272), .dout(n43415));
  jor  g25393(.dina(n43415), .dinb(n43413), .dout(remainder35 ));
  jand g25394(.dina(n43140), .dinb(n42679), .dout(n43417));
  jxor g25395(.dina(n43031), .dinb(n43216), .dout(n43418));
  jand g25396(.dina(n43418), .dinb(n43272), .dout(n43419));
  jor  g25397(.dina(n43419), .dinb(n43417), .dout(remainder36 ));
  jand g25398(.dina(n43140), .dinb(n42673), .dout(n43421));
  jxor g25399(.dina(n43035), .dinb(n43218), .dout(n43422));
  jand g25400(.dina(n43422), .dinb(n43272), .dout(n43423));
  jor  g25401(.dina(n43423), .dinb(n43421), .dout(remainder37 ));
  jand g25402(.dina(n43140), .dinb(n42667), .dout(n43425));
  jxor g25403(.dina(n43039), .dinb(n43220), .dout(n43426));
  jand g25404(.dina(n43426), .dinb(n43272), .dout(n43427));
  jor  g25405(.dina(n43427), .dinb(n43425), .dout(remainder38 ));
  jand g25406(.dina(n43140), .dinb(n42661), .dout(n43429));
  jxor g25407(.dina(n43043), .dinb(n43222), .dout(n43430));
  jand g25408(.dina(n43430), .dinb(n43272), .dout(n43431));
  jor  g25409(.dina(n43431), .dinb(n43429), .dout(remainder39 ));
  jand g25410(.dina(n43140), .dinb(n42655), .dout(n43433));
  jxor g25411(.dina(n43047), .dinb(n43224), .dout(n43434));
  jand g25412(.dina(n43434), .dinb(n43272), .dout(n43435));
  jor  g25413(.dina(n43435), .dinb(n43433), .dout(remainder40 ));
  jand g25414(.dina(n43140), .dinb(n42649), .dout(n43437));
  jxor g25415(.dina(n43051), .dinb(n43226), .dout(n43438));
  jand g25416(.dina(n43438), .dinb(n43272), .dout(n43439));
  jor  g25417(.dina(n43439), .dinb(n43437), .dout(remainder41 ));
  jand g25418(.dina(n43140), .dinb(n42643), .dout(n43441));
  jxor g25419(.dina(n43055), .dinb(n43228), .dout(n43442));
  jand g25420(.dina(n43442), .dinb(n43272), .dout(n43443));
  jor  g25421(.dina(n43443), .dinb(n43441), .dout(remainder42 ));
  jand g25422(.dina(n43140), .dinb(n42637), .dout(n43445));
  jxor g25423(.dina(n43059), .dinb(n43230), .dout(n43446));
  jand g25424(.dina(n43446), .dinb(n43272), .dout(n43447));
  jor  g25425(.dina(n43447), .dinb(n43445), .dout(remainder43 ));
  jand g25426(.dina(n43140), .dinb(n42631), .dout(n43449));
  jxor g25427(.dina(n43063), .dinb(n43232), .dout(n43450));
  jand g25428(.dina(n43450), .dinb(n43272), .dout(n43451));
  jor  g25429(.dina(n43451), .dinb(n43449), .dout(remainder44 ));
  jand g25430(.dina(n43140), .dinb(n42625), .dout(n43453));
  jxor g25431(.dina(n43067), .dinb(n43234), .dout(n43454));
  jand g25432(.dina(n43454), .dinb(n43272), .dout(n43455));
  jor  g25433(.dina(n43455), .dinb(n43453), .dout(remainder45 ));
  jand g25434(.dina(n43140), .dinb(n42619), .dout(n43457));
  jxor g25435(.dina(n43071), .dinb(n43236), .dout(n43458));
  jand g25436(.dina(n43458), .dinb(n43272), .dout(n43459));
  jor  g25437(.dina(n43459), .dinb(n43457), .dout(remainder46 ));
  jand g25438(.dina(n43140), .dinb(n42613), .dout(n43461));
  jxor g25439(.dina(n43075), .dinb(n43238), .dout(n43462));
  jand g25440(.dina(n43462), .dinb(n43272), .dout(n43463));
  jor  g25441(.dina(n43463), .dinb(n43461), .dout(remainder47 ));
  jand g25442(.dina(n43140), .dinb(n42607), .dout(n43465));
  jxor g25443(.dina(n43079), .dinb(n43240), .dout(n43466));
  jand g25444(.dina(n43466), .dinb(n43272), .dout(n43467));
  jor  g25445(.dina(n43467), .dinb(n43465), .dout(remainder48 ));
  jand g25446(.dina(n43140), .dinb(n42601), .dout(n43469));
  jxor g25447(.dina(n43083), .dinb(n43242), .dout(n43470));
  jand g25448(.dina(n43470), .dinb(n43272), .dout(n43471));
  jor  g25449(.dina(n43471), .dinb(n43469), .dout(remainder49 ));
  jand g25450(.dina(n43140), .dinb(n42595), .dout(n43473));
  jxor g25451(.dina(n43087), .dinb(n43244), .dout(n43474));
  jand g25452(.dina(n43474), .dinb(n43272), .dout(n43475));
  jor  g25453(.dina(n43475), .dinb(n43473), .dout(remainder50 ));
  jand g25454(.dina(n43140), .dinb(n42589), .dout(n43477));
  jxor g25455(.dina(n43091), .dinb(n43246), .dout(n43478));
  jand g25456(.dina(n43478), .dinb(n43272), .dout(n43479));
  jor  g25457(.dina(n43479), .dinb(n43477), .dout(remainder51 ));
  jand g25458(.dina(n43140), .dinb(n42583), .dout(n43481));
  jxor g25459(.dina(n43095), .dinb(n43248), .dout(n43482));
  jand g25460(.dina(n43482), .dinb(n43272), .dout(n43483));
  jor  g25461(.dina(n43483), .dinb(n43481), .dout(remainder52 ));
  jand g25462(.dina(n43140), .dinb(n42577), .dout(n43485));
  jxor g25463(.dina(n43099), .dinb(n43250), .dout(n43486));
  jand g25464(.dina(n43486), .dinb(n43272), .dout(n43487));
  jor  g25465(.dina(n43487), .dinb(n43485), .dout(remainder53 ));
  jand g25466(.dina(n43140), .dinb(n42571), .dout(n43489));
  jxor g25467(.dina(n43103), .dinb(n43252), .dout(n43490));
  jand g25468(.dina(n43490), .dinb(n43272), .dout(n43491));
  jor  g25469(.dina(n43491), .dinb(n43489), .dout(remainder54 ));
  jand g25470(.dina(n43140), .dinb(n42565), .dout(n43493));
  jxor g25471(.dina(n43107), .dinb(n43254), .dout(n43494));
  jand g25472(.dina(n43494), .dinb(n43272), .dout(n43495));
  jor  g25473(.dina(n43495), .dinb(n43493), .dout(remainder55 ));
  jand g25474(.dina(n43140), .dinb(n42559), .dout(n43497));
  jxor g25475(.dina(n43111), .dinb(n43256), .dout(n43498));
  jand g25476(.dina(n43498), .dinb(n43272), .dout(n43499));
  jor  g25477(.dina(n43499), .dinb(n43497), .dout(remainder56 ));
  jand g25478(.dina(n43140), .dinb(n42553), .dout(n43501));
  jxor g25479(.dina(n43115), .dinb(n43258), .dout(n43502));
  jand g25480(.dina(n43502), .dinb(n43272), .dout(n43503));
  jor  g25481(.dina(n43503), .dinb(n43501), .dout(remainder57 ));
  jand g25482(.dina(n43140), .dinb(n42547), .dout(n43505));
  jxor g25483(.dina(n43119), .dinb(n43260), .dout(n43506));
  jand g25484(.dina(n43506), .dinb(n43272), .dout(n43507));
  jor  g25485(.dina(n43507), .dinb(n43505), .dout(remainder58 ));
  jand g25486(.dina(n43140), .dinb(n42541), .dout(n43509));
  jxor g25487(.dina(n43123), .dinb(n43262), .dout(n43510));
  jand g25488(.dina(n43510), .dinb(n43272), .dout(n43511));
  jor  g25489(.dina(n43511), .dinb(n43509), .dout(remainder59 ));
  jand g25490(.dina(n43140), .dinb(n42535), .dout(n43513));
  jxor g25491(.dina(n43127), .dinb(n43264), .dout(n43514));
  jand g25492(.dina(n43514), .dinb(n43272), .dout(n43515));
  jor  g25493(.dina(n43515), .dinb(n43513), .dout(remainder60 ));
  jand g25494(.dina(n43140), .dinb(n42529), .dout(n43517));
  jxor g25495(.dina(n43131), .dinb(n43266), .dout(n43518));
  jand g25496(.dina(n43518), .dinb(n43272), .dout(n43519));
  jor  g25497(.dina(n43519), .dinb(n43517), .dout(remainder61 ));
  jand g25498(.dina(n43140), .dinb(n42523), .dout(n43521));
  jxor g25499(.dina(n43135), .dinb(n43268), .dout(n43522));
  jand g25500(.dina(n43522), .dinb(n43272), .dout(n43523));
  jor  g25501(.dina(n43523), .dinb(n43521), .dout(remainder62 ));
  jand g25502(.dina(n43270), .dinb(n42515), .dout(n43525));
  jand g25503(.dina(n43139), .dinb(n42514), .dout(n43526));
  jor  g25504(.dina(n43526), .dinb(n43525), .dout(remainder63 ));
endmodule


