/*

c1908:
	jxor: 78
	jspl: 105
	jspl3: 86
	jnot: 30
	jdff: 969
	jor: 87
	jand: 120

Summary:
	jxor: 78
	jspl: 105
	jspl3: 86
	jnot: 30
	jdff: 969
	jor: 87
	jand: 120
*/

module c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n173;
	wire n174;
	wire n175;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n201;
	wire n203;
	wire n204;
	wire n206;
	wire n207;
	wire n208;
	wire n210;
	wire n211;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n220;
	wire n222;
	wire n223;
	wire n224;
	wire n226;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n270;
	wire n271;
	wire n272;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n348;
	wire n349;
	wire n350;
	wire n352;
	wire n353;
	wire n354;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n369;
	wire n370;
	wire n371;
	wire[2:0] w_G101_0;
	wire[2:0] w_G104_0;
	wire[2:0] w_G107_0;
	wire[2:0] w_G110_0;
	wire[2:0] w_G113_0;
	wire[2:0] w_G116_0;
	wire[2:0] w_G119_0;
	wire[2:0] w_G122_0;
	wire[1:0] w_G122_1;
	wire[2:0] w_G125_0;
	wire[2:0] w_G128_0;
	wire[2:0] w_G131_0;
	wire[2:0] w_G134_0;
	wire[2:0] w_G137_0;
	wire[2:0] w_G140_0;
	wire[2:0] w_G143_0;
	wire[2:0] w_G146_0;
	wire[2:0] w_G210_0;
	wire[1:0] w_G214_0;
	wire[2:0] w_G217_0;
	wire[1:0] w_G221_0;
	wire[1:0] w_G224_0;
	wire[1:0] w_G227_0;
	wire[2:0] w_G234_0;
	wire[1:0] w_G234_1;
	wire[2:0] w_G237_0;
	wire[2:0] w_G469_0;
	wire[2:0] w_G472_0;
	wire[2:0] w_G475_0;
	wire[2:0] w_G478_0;
	wire[1:0] w_G898_0;
	wire[1:0] w_G900_0;
	wire[2:0] w_G902_0;
	wire[2:0] w_G902_1;
	wire[2:0] w_G902_2;
	wire[2:0] w_G902_3;
	wire[2:0] w_G952_0;
	wire[2:0] w_G953_0;
	wire[2:0] w_G953_1;
	wire[1:0] w_G953_2;
	wire[2:0] w_n58_0;
	wire[2:0] w_n58_1;
	wire[2:0] w_n58_2;
	wire[1:0] w_n63_0;
	wire[1:0] w_n66_0;
	wire[1:0] w_n67_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n71_0;
	wire[1:0] w_n73_0;
	wire[1:0] w_n74_0;
	wire[2:0] w_n76_0;
	wire[2:0] w_n76_1;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[2:0] w_n81_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[1:0] w_n90_0;
	wire[1:0] w_n91_0;
	wire[2:0] w_n92_0;
	wire[1:0] w_n92_1;
	wire[2:0] w_n93_0;
	wire[1:0] w_n93_1;
	wire[1:0] w_n94_0;
	wire[2:0] w_n95_0;
	wire[1:0] w_n95_1;
	wire[2:0] w_n96_0;
	wire[1:0] w_n99_0;
	wire[1:0] w_n102_0;
	wire[2:0] w_n103_0;
	wire[2:0] w_n103_1;
	wire[2:0] w_n103_2;
	wire[2:0] w_n103_3;
	wire[1:0] w_n107_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n109_0;
	wire[1:0] w_n110_0;
	wire[1:0] w_n111_0;
	wire[2:0] w_n112_0;
	wire[1:0] w_n112_1;
	wire[2:0] w_n113_0;
	wire[1:0] w_n118_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[1:0] w_n121_0;
	wire[2:0] w_n122_0;
	wire[1:0] w_n122_1;
	wire[1:0] w_n124_0;
	wire[1:0] w_n126_0;
	wire[1:0] w_n127_0;
	wire[2:0] w_n130_0;
	wire[1:0] w_n130_1;
	wire[2:0] w_n131_0;
	wire[2:0] w_n131_1;
	wire[1:0] w_n139_0;
	wire[1:0] w_n140_0;
	wire[2:0] w_n141_0;
	wire[1:0] w_n141_1;
	wire[2:0] w_n151_0;
	wire[1:0] w_n152_0;
	wire[2:0] w_n153_0;
	wire[1:0] w_n153_1;
	wire[2:0] w_n154_0;
	wire[1:0] w_n154_1;
	wire[1:0] w_n155_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n157_0;
	wire[2:0] w_n160_0;
	wire[2:0] w_n160_1;
	wire[2:0] w_n161_0;
	wire[1:0] w_n161_1;
	wire[1:0] w_n162_0;
	wire[2:0] w_n163_0;
	wire[1:0] w_n163_1;
	wire[1:0] w_n164_0;
	wire[2:0] w_n165_0;
	wire[1:0] w_n166_0;
	wire[2:0] w_n168_0;
	wire[1:0] w_n168_1;
	wire[1:0] w_n169_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n171_0;
	wire[2:0] w_n173_0;
	wire[1:0] w_n173_1;
	wire[1:0] w_n174_0;
	wire[1:0] w_n175_0;
	wire[2:0] w_n177_0;
	wire[1:0] w_n178_0;
	wire[1:0] w_n180_0;
	wire[2:0] w_n182_0;
	wire[2:0] w_n182_1;
	wire[2:0] w_n183_0;
	wire[1:0] w_n184_0;
	wire[1:0] w_n186_0;
	wire[1:0] w_n189_0;
	wire[2:0] w_n191_0;
	wire[2:0] w_n192_0;
	wire[2:0] w_n195_0;
	wire[2:0] w_n197_0;
	wire[1:0] w_n197_1;
	wire[1:0] w_n198_0;
	wire[2:0] w_n199_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n208_0;
	wire[1:0] w_n210_0;
	wire[1:0] w_n211_0;
	wire[2:0] w_n214_0;
	wire[2:0] w_n216_0;
	wire[1:0] w_n216_1;
	wire[1:0] w_n217_0;
	wire[1:0] w_n218_0;
	wire[1:0] w_n220_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n226_0;
	wire[2:0] w_n242_0;
	wire[2:0] w_n242_1;
	wire[2:0] w_n242_2;
	wire[1:0] w_n243_0;
	wire[1:0] w_n249_0;
	wire[2:0] w_n258_0;
	wire[2:0] w_n265_0;
	wire[2:0] w_n265_1;
	wire[1:0] w_n265_2;
	wire[1:0] w_n274_0;
	wire[2:0] w_n278_0;
	wire[1:0] w_n279_0;
	wire[1:0] w_n280_0;
	wire[2:0] w_n282_0;
	wire[1:0] w_n282_1;
	wire[1:0] w_n286_0;
	wire[2:0] w_n287_0;
	wire[1:0] w_n287_1;
	wire[1:0] w_n288_0;
	wire[2:0] w_n291_0;
	wire[1:0] w_n291_1;
	wire[1:0] w_n292_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n294_0;
	wire[1:0] w_n297_0;
	wire[1:0] w_n303_0;
	wire[2:0] w_n307_0;
	wire[1:0] w_n313_0;
	wire[2:0] w_n316_0;
	wire[2:0] w_n317_0;
	wire[1:0] w_n322_0;
	wire[1:0] w_n323_0;
	wire[1:0] w_n327_0;
	wire[1:0] w_n329_0;
	wire[1:0] w_n341_0;
	wire w_dff_B_CdRx2ofj8_0;
	wire w_dff_B_Jofgn1S76_0;
	wire w_dff_B_tSrBdNNg0_0;
	wire w_dff_B_uzJKMgZJ8_0;
	wire w_dff_B_mdhrHRyX3_0;
	wire w_dff_B_rKkOArAP6_0;
	wire w_dff_B_2UGfDtp09_0;
	wire w_dff_B_EjutnVrS9_0;
	wire w_dff_A_PKCFZb8h0_0;
	wire w_dff_A_dSFONKfV8_0;
	wire w_dff_B_bWLtcQoM2_0;
	wire w_dff_B_rTOt5aZC3_0;
	wire w_dff_B_P74BFHHB6_0;
	wire w_dff_B_qX0R8aqj3_0;
	wire w_dff_B_Y7JkvRCC7_0;
	wire w_dff_B_UhkGRgaT1_1;
	wire w_dff_B_gvI1qoJE5_1;
	wire w_dff_B_Ss4VEQKz8_1;
	wire w_dff_B_RoDxmlQO3_1;
	wire w_dff_B_noQphQOk8_1;
	wire w_dff_B_G6zvj8GB8_1;
	wire w_dff_B_33x2tQbN4_1;
	wire w_dff_B_kUGQb4pD9_1;
	wire w_dff_B_SkxkywiX2_1;
	wire w_dff_B_vqkQtcQR0_1;
	wire w_dff_B_GvNAzZn29_1;
	wire w_dff_B_Pdmthr8R4_1;
	wire w_dff_B_E4Ub7aYc9_0;
	wire w_dff_B_BJZXmpsT4_0;
	wire w_dff_B_Rw3IvUap5_0;
	wire w_dff_B_VQsxdqKi4_0;
	wire w_dff_B_NAPbsLZ77_0;
	wire w_dff_B_SNo6lWGV8_0;
	wire w_dff_B_s02w2U9v6_0;
	wire w_dff_B_lQ3kIVHT5_0;
	wire w_dff_B_Umxg7UHQ6_0;
	wire w_dff_B_wD9nMmlb6_0;
	wire w_dff_B_dMIT6iMI9_0;
	wire w_dff_B_P7YEjKFB7_0;
	wire w_dff_B_dEkIWPHf4_0;
	wire w_dff_B_xTtMqEP62_0;
	wire w_dff_A_01Zlvuku6_1;
	wire w_dff_A_JyQbwjjG5_1;
	wire w_dff_A_RGq2ecjx2_1;
	wire w_dff_A_BxZUUVZb4_1;
	wire w_dff_A_BAX7EPEZ4_1;
	wire w_dff_A_NiXjGfW73_1;
	wire w_dff_A_ULNlmOgF4_1;
	wire w_dff_A_IDzbWCqW0_1;
	wire w_dff_A_Fa6hmuCA7_1;
	wire w_dff_A_4FTO6hXT7_1;
	wire w_dff_A_2ccFVnGw1_1;
	wire w_dff_A_9ZosgNHH8_1;
	wire w_dff_A_W4IyJAAy8_1;
	wire w_dff_A_46gwKBMl0_1;
	wire w_dff_A_DIdKlfsT9_1;
	wire w_dff_A_Y3wGLXRM6_1;
	wire w_dff_A_JgZ3KUDw3_1;
	wire w_dff_A_g9GM441z5_1;
	wire w_dff_A_utWSeLvC1_1;
	wire w_dff_A_8e7MtCfJ0_1;
	wire w_dff_A_etSqSXhN7_1;
	wire w_dff_A_HivJmHxQ4_1;
	wire w_dff_A_scdTvfje6_1;
	wire w_dff_A_GGnSifdZ0_1;
	wire w_dff_A_iJL4TF6P3_1;
	wire w_dff_A_6c9bOjaF0_1;
	wire w_dff_A_6QuDRRlY4_1;
	wire w_dff_A_LefPmnEp8_1;
	wire w_dff_A_JNikaNm51_1;
	wire w_dff_A_jg6GCSEe1_1;
	wire w_dff_A_Xm3ei6mZ7_1;
	wire w_dff_A_VyTK4dvY7_1;
	wire w_dff_A_97odHxbd8_2;
	wire w_dff_A_1geQscUf2_2;
	wire w_dff_A_V2qqzgfI7_2;
	wire w_dff_A_IEObQtub7_2;
	wire w_dff_A_z0XG4Ye59_2;
	wire w_dff_A_M7usmQGk8_2;
	wire w_dff_A_0nY5riSl9_2;
	wire w_dff_A_krg8bAKb9_2;
	wire w_dff_A_raRC3OMP1_2;
	wire w_dff_A_6WVtgcq52_2;
	wire w_dff_A_WxVODHg12_2;
	wire w_dff_A_rkvpdkLv3_2;
	wire w_dff_A_DPq1QHOl5_2;
	wire w_dff_A_HQ7adru01_2;
	wire w_dff_A_RXlS4zgb6_2;
	wire w_dff_A_PfNa3u4S7_2;
	wire w_dff_A_WN7aDri63_2;
	wire w_dff_A_eSyyHdl70_0;
	wire w_dff_A_ClAuuYEU2_1;
	wire w_dff_B_KLwBtMBo5_1;
	wire w_dff_B_Pqzg5Onq1_1;
	wire w_dff_B_580wu7Pw4_1;
	wire w_dff_B_8MBa5YkG5_1;
	wire w_dff_B_jCJcTw8x9_1;
	wire w_dff_B_mNbCnYs29_1;
	wire w_dff_B_Iu3AWsBL9_1;
	wire w_dff_B_HhoRgETG3_1;
	wire w_dff_B_ggwC78Ie4_1;
	wire w_dff_B_kddSgT1I0_1;
	wire w_dff_B_32whL4Fq2_1;
	wire w_dff_B_mm3w6rtw5_1;
	wire w_dff_B_sZyVdW0g1_0;
	wire w_dff_B_fwm0Thr30_0;
	wire w_dff_B_WKX6vTOm1_0;
	wire w_dff_B_7jWup1Di6_0;
	wire w_dff_B_r5yi4Ilk2_0;
	wire w_dff_B_7dfcLZX26_0;
	wire w_dff_B_3vQk8ReK6_0;
	wire w_dff_B_Nf4iurPA5_0;
	wire w_dff_B_v0JEP4p01_0;
	wire w_dff_B_G059g5QF4_0;
	wire w_dff_B_OIzh3tr73_0;
	wire w_dff_B_qMy3jbYl2_0;
	wire w_dff_B_9igCQlhx5_0;
	wire w_dff_B_CT4BKni72_0;
	wire w_dff_B_H0KRGSsn2_1;
	wire w_dff_B_XYKnHp0j2_1;
	wire w_dff_B_5rQkiA8U2_1;
	wire w_dff_B_IBTGc6487_1;
	wire w_dff_B_D7S2f1cO7_2;
	wire w_dff_A_KyQhiGUQ8_1;
	wire w_dff_B_GBnHB9Zw8_2;
	wire w_dff_A_E82yDAXB3_2;
	wire w_dff_A_T9L4824r0_2;
	wire w_dff_B_ZUyHbJGO8_3;
	wire w_dff_B_642pIuUB7_3;
	wire w_dff_B_bw6JouIo8_0;
	wire w_dff_B_nrGvtlF21_0;
	wire w_dff_B_dfrEfNZa3_0;
	wire w_dff_B_85COfi2C0_0;
	wire w_dff_B_AHPfHRnc0_0;
	wire w_dff_B_3V0w02l23_0;
	wire w_dff_B_8LlYVvKp9_0;
	wire w_dff_B_Rw29LyWx0_0;
	wire w_dff_B_qr30Hv1l1_0;
	wire w_dff_B_lRvMcX6T0_0;
	wire w_dff_B_xlV9W2jf8_0;
	wire w_dff_B_pHDAhxtA7_0;
	wire w_dff_B_yr50cWre3_0;
	wire w_dff_B_aUCGbcsC7_0;
	wire w_dff_B_IcUCqYEo6_0;
	wire w_dff_B_sJs3Z4DR0_0;
	wire w_dff_B_RwsggDky2_0;
	wire w_dff_B_n4RqY0dh1_0;
	wire w_dff_B_myFuCQOt5_0;
	wire w_dff_B_O9WwE1F88_0;
	wire w_dff_B_qlIthqTp6_0;
	wire w_dff_B_G6zDwesT8_0;
	wire w_dff_B_kPJIySp34_0;
	wire w_dff_B_MWH7XePi5_0;
	wire w_dff_B_FJyLm5td2_0;
	wire w_dff_B_XgqYe2sI5_0;
	wire w_dff_B_jaVsgVn29_1;
	wire w_dff_B_favqS1wC0_1;
	wire w_dff_B_S6Ympi2H6_1;
	wire w_dff_A_DEqNbgcH4_1;
	wire w_dff_A_x6yjkDmP3_2;
	wire w_dff_A_ZODl5Moa2_1;
	wire w_dff_A_8refZzbe8_1;
	wire w_dff_A_moB27oGJ2_1;
	wire w_dff_A_MWZ48N6Z3_2;
	wire w_dff_A_Ql1RQxrt9_1;
	wire w_dff_A_U0yY5g6B5_0;
	wire w_dff_A_3bKSKJPS4_2;
	wire w_dff_A_vRssUqsX6_0;
	wire w_dff_A_WvrPjgf76_1;
	wire w_dff_B_8U3ot9Yd8_2;
	wire w_dff_A_QwYvSUKV8_0;
	wire w_dff_A_YwRCZHgK4_2;
	wire w_dff_A_LnZaJCs82_0;
	wire w_dff_A_Fxn3f38s5_2;
	wire w_dff_B_iF8xxByB5_3;
	wire w_dff_B_KSiHxSKO7_3;
	wire w_dff_A_aiYopAbc9_1;
	wire w_dff_A_4HYK9vc51_2;
	wire w_dff_B_VMwPWO1d1_0;
	wire w_dff_B_05WJY39F9_0;
	wire w_dff_B_F0oEXzHH5_0;
	wire w_dff_B_FmogL4Tr6_0;
	wire w_dff_B_PVEGtvjN1_0;
	wire w_dff_B_DLzdOQkj4_0;
	wire w_dff_B_XLT3ylCP2_0;
	wire w_dff_B_DxleLwwm5_0;
	wire w_dff_B_qnQsVxvs5_0;
	wire w_dff_B_2H44TzEw4_0;
	wire w_dff_B_E2OGXQWx4_0;
	wire w_dff_B_T60XriuG8_0;
	wire w_dff_B_dbNB63XD4_0;
	wire w_dff_B_UcTr2xLm2_0;
	wire w_dff_B_iHdfZUwO1_0;
	wire w_dff_A_QDdCYJo07_1;
	wire w_dff_A_JRGb2gXD7_1;
	wire w_dff_A_PmhDL7eN5_1;
	wire w_dff_A_Kr47xTpf5_1;
	wire w_dff_A_lKPvVncS4_1;
	wire w_dff_A_5q0iiHtL2_1;
	wire w_dff_A_rqkgNDsE1_1;
	wire w_dff_A_C7DW2jBL0_1;
	wire w_dff_A_UN8YvMYk7_1;
	wire w_dff_A_2qnLViUH1_1;
	wire w_dff_A_ZVEVOxHd0_1;
	wire w_dff_A_fzb2ey0u6_1;
	wire w_dff_A_4aRytuxL4_1;
	wire w_dff_A_ayle6BcB5_1;
	wire w_dff_A_JKobmPW97_1;
	wire w_dff_A_b4baawxQ5_1;
	wire w_dff_A_Xa2aGWVJ7_1;
	wire w_dff_A_u7xQmrzd0_2;
	wire w_dff_A_BipGxom86_2;
	wire w_dff_A_7MWomFnc0_2;
	wire w_dff_A_aySddW5V9_2;
	wire w_dff_A_QL6ZRlOf8_2;
	wire w_dff_A_07B2X1Ur5_2;
	wire w_dff_A_i60C2Ups4_2;
	wire w_dff_A_Xyp4qGUm3_2;
	wire w_dff_A_w2vnCVdz4_2;
	wire w_dff_A_7Y6mJfUR5_2;
	wire w_dff_A_BrrfhQ5v1_2;
	wire w_dff_A_ycwMGVna9_2;
	wire w_dff_A_eNZWx0B75_2;
	wire w_dff_A_jBTPX2LO1_2;
	wire w_dff_A_HFqMOeIh1_2;
	wire w_dff_A_5z7CCzzn1_2;
	wire w_dff_A_TPWjdESN3_2;
	wire w_dff_B_HfhpR8ps8_1;
	wire w_dff_B_8bRbkbHo2_1;
	wire w_dff_A_nft3XXuY3_0;
	wire w_dff_A_sdWzoRyN7_1;
	wire w_dff_A_YL2Miv7Q0_2;
	wire w_dff_A_mvYfA7ak6_0;
	wire w_dff_A_sehqTj2E5_2;
	wire w_dff_B_yc4fuzHt1_0;
	wire w_dff_B_x0dXhVj88_0;
	wire w_dff_B_9Vd1GOLh7_0;
	wire w_dff_A_t2ZLaWgT3_1;
	wire w_dff_A_6H0WDGGA8_0;
	wire w_dff_A_bCtB2c645_2;
	wire w_dff_A_QnfWgLoo0_1;
	wire w_dff_A_jGjusVUl4_0;
	wire w_dff_A_wGfFCvUd2_0;
	wire w_dff_A_WL8mdX3K8_0;
	wire w_dff_A_Gf1fOO9v0_2;
	wire w_dff_A_4Dnh2owz6_2;
	wire w_dff_A_Axm0Vv1I7_2;
	wire w_dff_A_YoKxsKfO2_2;
	wire w_dff_A_y3BIuxuQ6_0;
	wire w_dff_A_o5HX76V06_1;
	wire w_dff_A_yuQe9kTT3_1;
	wire w_dff_A_r82Pybnj4_2;
	wire w_dff_A_Eo3OP6EE2_0;
	wire w_dff_A_H2zQJU8B6_1;
	wire w_dff_B_2dksoSKa9_2;
	wire w_dff_A_ljf1Bi7P1_1;
	wire w_dff_A_yPIgSjky6_1;
	wire w_dff_A_3UBavrO18_0;
	wire w_dff_B_bAL3FZPL7_2;
	wire w_dff_A_vbbhBETj6_2;
	wire w_dff_A_YQvrdROC5_2;
	wire w_dff_A_Rn7lfHCP7_2;
	wire w_dff_A_TB3CFVc45_2;
	wire w_dff_B_raM7NCsX4_1;
	wire w_dff_B_b594Y2jO9_1;
	wire w_dff_B_ztlquN5g3_1;
	wire w_dff_B_oA9mZ8LN9_1;
	wire w_dff_B_Mxv7YFLo4_1;
	wire w_dff_A_bs9puDA28_1;
	wire w_dff_A_gt2VHgWJ4_1;
	wire w_dff_A_LhbJ3WDd8_1;
	wire w_dff_A_OsegNpXQ2_2;
	wire w_dff_A_CSeTQGlo6_0;
	wire w_dff_A_dWLe2s8Q4_1;
	wire w_dff_A_XBGQncMn4_2;
	wire w_dff_B_dIolIVmb4_1;
	wire w_dff_B_fvnInEzm1_1;
	wire w_dff_B_Yg7vPTC64_1;
	wire w_dff_B_dvmuNwsN3_1;
	wire w_dff_B_nKMMM2cI3_1;
	wire w_dff_A_BqKbgA812_1;
	wire w_dff_A_rQqc1nWU3_0;
	wire w_dff_A_D6wwbt1I7_1;
	wire w_dff_B_cYVFmp2Q2_1;
	wire w_dff_B_AAI2YqKa1_1;
	wire w_dff_B_nFzxAVfw5_1;
	wire w_dff_B_hNv2kRgM7_1;
	wire w_dff_B_EZajK4Zx4_1;
	wire w_dff_A_mWbAcvmq0_0;
	wire w_dff_A_FeUaWPZB4_0;
	wire w_dff_A_7vFu0o4n8_0;
	wire w_dff_A_MbAnB5Qd6_0;
	wire w_dff_A_MNOQRZPF0_0;
	wire w_dff_A_AUxs2JCG2_0;
	wire w_dff_A_qQ9Fba7L5_0;
	wire w_dff_A_knnKQf9j0_0;
	wire w_dff_A_AAeKoEmm2_0;
	wire w_dff_A_znJYkK2h1_0;
	wire w_dff_A_XtzpvVlA5_0;
	wire w_dff_A_CqFgFXHW0_0;
	wire w_dff_A_wqXB6xBt2_0;
	wire w_dff_A_PSy1Ef8v9_1;
	wire w_dff_A_fTujv3rS0_0;
	wire w_dff_A_W26QZD3x7_0;
	wire w_dff_A_glZCvSbV0_0;
	wire w_dff_A_LfdWhR0k2_0;
	wire w_dff_A_BIkT6B4Y6_0;
	wire w_dff_A_152QaVWZ4_0;
	wire w_dff_A_TVAszvr33_0;
	wire w_dff_A_jQwZCwyL4_0;
	wire w_dff_A_RmLCvJR08_0;
	wire w_dff_A_FsXolQU91_0;
	wire w_dff_A_USbeHMh75_0;
	wire w_dff_A_g0hz9BCR9_0;
	wire w_dff_A_jJXHTid63_0;
	wire w_dff_A_fts2igdj9_0;
	wire w_dff_A_9afLu5cr4_0;
	wire w_dff_A_Ki5uAwD32_0;
	wire w_dff_A_qTumxMiU7_2;
	wire w_dff_A_VjfWHbZr1_2;
	wire w_dff_A_4ygaUCMi0_2;
	wire w_dff_A_OeVzAPap7_2;
	wire w_dff_A_aEk61aJ43_2;
	wire w_dff_A_Ainhjsqa1_2;
	wire w_dff_A_Fao2cAqc6_1;
	wire w_dff_A_pQOq6Uh58_1;
	wire w_dff_A_37wy3utU9_2;
	wire w_dff_A_glx4b2HU7_2;
	wire w_dff_A_MyexSgyj5_1;
	wire w_dff_A_jsgNo3aG6_1;
	wire w_dff_A_szorhQwO6_1;
	wire w_dff_A_Z9JB7D5B1_2;
	wire w_dff_A_BMhIXWMj5_2;
	wire w_dff_A_4ZH5GRqy3_2;
	wire w_dff_A_wxCamwqG0_1;
	wire w_dff_A_vs0lCKW85_1;
	wire w_dff_A_PKSGSRMF5_1;
	wire w_dff_A_XXodlFnk5_1;
	wire w_dff_A_Jq81yBNG1_0;
	wire w_dff_A_mbCLDJc58_0;
	wire w_dff_A_eVJwQ8Rd6_0;
	wire w_dff_A_dlUm5GdS9_0;
	wire w_dff_A_5l6aGnp06_0;
	wire w_dff_A_6Znmh7On2_0;
	wire w_dff_A_KBIeAkO20_0;
	wire w_dff_A_7bhc17KK1_0;
	wire w_dff_A_ovrl5xYy2_0;
	wire w_dff_A_MUlJkXFG9_0;
	wire w_dff_A_koMlqWKZ0_0;
	wire w_dff_A_ohN5pEQc0_0;
	wire w_dff_A_8DSmAR8e6_0;
	wire w_dff_B_OOoXnuC15_1;
	wire w_dff_A_wdwqTUD03_1;
	wire w_dff_B_yLgtjOzk6_0;
	wire w_dff_B_tglVqJNZ7_0;
	wire w_dff_A_dYQ2sOnO3_0;
	wire w_dff_A_Jjn2Iy6I8_1;
	wire w_dff_A_kiIlB8Vh1_1;
	wire w_dff_A_PFqwSlRL6_2;
	wire w_dff_A_H8F0IXdL4_2;
	wire w_dff_B_O4s8zUHl7_3;
	wire w_dff_B_JCHEIWWr5_3;
	wire w_dff_A_5YQM2Dv99_0;
	wire w_dff_A_ufFIFDr17_0;
	wire w_dff_A_in8rgn4A9_1;
	wire w_dff_A_kvKSfVHq6_1;
	wire w_dff_A_lp5uNfOn0_1;
	wire w_dff_A_ChyF10g46_1;
	wire w_dff_A_TAIfjDqB5_1;
	wire w_dff_A_hTI2R2GC7_2;
	wire w_dff_A_O8CXT4Og7_2;
	wire w_dff_A_ECJUwDdp2_2;
	wire w_dff_A_9pp1EhMF8_2;
	wire w_dff_A_0SNZBjMI2_2;
	wire w_dff_A_4mbwf4eE1_1;
	wire w_dff_A_Yc2wWo9e0_2;
	wire w_dff_B_LUzLjp6Q9_3;
	wire w_dff_B_IbDQEo7i1_1;
	wire w_dff_B_hFX4NJtE3_1;
	wire w_dff_B_YeSQtdKL2_1;
	wire w_dff_B_373lpKxb8_1;
	wire w_dff_B_oEXkI1vY7_1;
	wire w_dff_A_IVJjGBzk6_0;
	wire w_dff_A_XpbkbB1C2_0;
	wire w_dff_A_fSRLNKkA8_0;
	wire w_dff_A_HvLa1AXe2_0;
	wire w_dff_A_uyyNAPEa2_0;
	wire w_dff_A_3jmxAeI24_0;
	wire w_dff_A_P1ifWpEv2_0;
	wire w_dff_A_Hrd8bJTN3_0;
	wire w_dff_A_eS4RkAuC2_0;
	wire w_dff_A_cVEwS4jw2_0;
	wire w_dff_A_bwh7ArJO1_0;
	wire w_dff_A_lDGQmxr08_0;
	wire w_dff_A_WaaanRHD1_0;
	wire w_dff_A_X4uqIgWo4_0;
	wire w_dff_A_MU7cEkiq8_0;
	wire w_dff_A_RMZzRwnv4_0;
	wire w_dff_A_mXfaxYyM3_0;
	wire w_dff_A_VD3Cy5BD7_0;
	wire w_dff_A_AkfgV1Eh4_0;
	wire w_dff_A_Tjz2ZwEm3_0;
	wire w_dff_A_YCF3mrwO9_0;
	wire w_dff_A_HWNHflyG8_0;
	wire w_dff_A_bDfma8U30_0;
	wire w_dff_A_Iu1zOiwH6_0;
	wire w_dff_A_TAGELWTD5_0;
	wire w_dff_A_TfkoPOzq8_0;
	wire w_dff_A_TTg2vcIa2_0;
	wire w_dff_A_Dvrpoyht9_0;
	wire w_dff_A_Fnzdoirm6_1;
	wire w_dff_A_63Xj2V504_0;
	wire w_dff_A_7ptXhgKe3_0;
	wire w_dff_A_okrlDpS29_0;
	wire w_dff_A_I8vmvHrG2_0;
	wire w_dff_A_7M5jHN025_0;
	wire w_dff_A_7gCRq0WD5_0;
	wire w_dff_A_Oo6WF2vO3_0;
	wire w_dff_A_vXHwLd4q7_0;
	wire w_dff_A_HmwdAIXL9_0;
	wire w_dff_A_2Se3tiNk8_0;
	wire w_dff_A_R8YlHE2w3_0;
	wire w_dff_A_6g28ZD0h5_2;
	wire w_dff_A_VXWWuc3X5_2;
	wire w_dff_A_DTpVIFKE5_1;
	wire w_dff_A_0W73h6m64_1;
	wire w_dff_A_1jcsAr9G2_2;
	wire w_dff_A_hVdLlbEz0_2;
	wire w_dff_A_hL5gAhwG1_2;
	wire w_dff_A_XAJyGXLt1_2;
	wire w_dff_A_4odj30ia1_2;
	wire w_dff_A_zpzRYhAj1_2;
	wire w_dff_A_ngie6Vjf5_2;
	wire w_dff_B_gdUnpY1m1_0;
	wire w_dff_A_RwYGsJCT6_0;
	wire w_dff_A_O1ecZPEC7_0;
	wire w_dff_A_hgOT9GkU1_0;
	wire w_dff_A_GXhKf2iZ7_0;
	wire w_dff_A_gZQjpllN0_0;
	wire w_dff_A_TT9wvXy35_0;
	wire w_dff_A_yrBFt94H4_0;
	wire w_dff_A_lQpPB3ZW5_0;
	wire w_dff_A_qCeLwvIR4_0;
	wire w_dff_A_0rwgrJoI1_0;
	wire w_dff_A_AXRqwrCx0_0;
	wire w_dff_A_RSaRzvei8_0;
	wire w_dff_A_QZSIMUtJ3_0;
	wire w_dff_A_xs6BUOcj4_0;
	wire w_dff_A_RtDpuMvy0_0;
	wire w_dff_B_fOfk53P32_0;
	wire w_dff_B_SezSqpel8_0;
	wire w_dff_A_pKZNHe552_0;
	wire w_dff_A_3oi60fMZ4_0;
	wire w_dff_A_mhuuLXXT6_0;
	wire w_dff_A_d1KPOBMq1_0;
	wire w_dff_A_mHAJuHcK2_0;
	wire w_dff_A_Hpte4vfu5_0;
	wire w_dff_A_TK4fxhqT6_0;
	wire w_dff_A_S0XfC0pO6_0;
	wire w_dff_A_g5sZoqxD7_0;
	wire w_dff_A_kk5aMkAw7_0;
	wire w_dff_A_QKqVNlEN5_0;
	wire w_dff_B_E2gMzbzZ7_0;
	wire w_dff_A_tNTC83n08_0;
	wire w_dff_A_ksZUfEAq9_0;
	wire w_dff_A_sJWnaMA38_0;
	wire w_dff_A_j4SrJ4Ch5_0;
	wire w_dff_A_btybmDyg1_0;
	wire w_dff_A_pDflvThv8_0;
	wire w_dff_A_sBiep1zc3_0;
	wire w_dff_A_OsVdRZSh4_0;
	wire w_dff_A_IfvaPOnB3_0;
	wire w_dff_A_uAxIQxjG2_0;
	wire w_dff_A_I5DHfcvg5_0;
	wire w_dff_A_0lugVVhC9_2;
	wire w_dff_A_5Asyo8uZ5_0;
	wire w_dff_A_9eEG8FuC2_0;
	wire w_dff_A_OwOH84eF1_0;
	wire w_dff_A_xNDl61YB7_0;
	wire w_dff_A_8acG0xR55_0;
	wire w_dff_A_rRjvU9CP0_0;
	wire w_dff_A_FV2sbfqf7_0;
	wire w_dff_A_WaBbkL3Z2_0;
	wire w_dff_A_QQGZNuYD6_0;
	wire w_dff_A_JXdWwEvB1_0;
	wire w_dff_A_sEbjAvFW8_0;
	wire w_dff_B_MYlh2hkP6_1;
	wire w_dff_A_FpyAogCZ2_0;
	wire w_dff_A_WuZeBu4y0_0;
	wire w_dff_A_WxG6asbp1_0;
	wire w_dff_A_bfGVxm1p0_0;
	wire w_dff_A_1X4jttEt0_0;
	wire w_dff_A_ks7Lw3Sr8_0;
	wire w_dff_A_PUx7N4Rs1_0;
	wire w_dff_A_rQECRfdN9_0;
	wire w_dff_A_JJUYwFe61_2;
	wire w_dff_A_o3ZTjruz8_2;
	wire w_dff_A_RPe0UhA67_2;
	wire w_dff_A_1kggSPbO3_2;
	wire w_dff_A_Z90Zwh8F3_0;
	wire w_dff_A_n8nmovg17_0;
	wire w_dff_A_I8pmQhjl7_0;
	wire w_dff_A_2GMuLE8Z3_2;
	wire w_dff_A_lJ5AhLZ90_2;
	wire w_dff_A_J4tJ1UPO0_2;
	wire w_dff_A_hgCRujL88_2;
	wire w_dff_A_BGe6APbO8_2;
	wire w_dff_A_Uv9nZhjH3_1;
	wire w_dff_A_qnLsnTcA7_1;
	wire w_dff_A_EGiaBh7U6_1;
	wire w_dff_A_yMoIAGfu6_1;
	wire w_dff_A_7XIVxcxE2_2;
	wire w_dff_A_8o5KYpZZ0_2;
	wire w_dff_A_GR1uVg2b9_2;
	wire w_dff_A_Bxamrgzn8_2;
	wire w_dff_A_VWtukREt6_2;
	wire w_dff_A_wE6cvfsv4_2;
	wire w_dff_A_35AQNABq7_2;
	wire w_dff_A_iwleWXhp5_2;
	wire w_dff_A_EfsTyA2Z4_2;
	wire w_dff_A_O9bDVYXm7_0;
	wire w_dff_A_WgfzuJgN5_1;
	wire w_dff_A_3b2YPRZZ3_0;
	wire w_dff_A_cfc6Fpsw1_0;
	wire w_dff_A_0S7blAa62_0;
	wire w_dff_A_KZ7hGh7y2_1;
	wire w_dff_A_fwasoT2e1_1;
	wire w_dff_A_RuHp7h8W7_1;
	wire w_dff_A_xt1G26Iq5_1;
	wire w_dff_A_ot761LEK5_1;
	wire w_dff_A_jucyTyvX1_1;
	wire w_dff_A_o6nx9h7l6_1;
	wire w_dff_A_0FXadMBX7_1;
	wire w_dff_A_SM2TfiJu9_1;
	wire w_dff_A_fmEMOViY1_1;
	wire w_dff_A_eDYUT59i0_1;
	wire w_dff_A_05lP8yaM7_1;
	wire w_dff_B_7UJZZigs3_1;
	wire w_dff_B_RpTxSUap7_1;
	wire w_dff_A_6abGK1HB3_0;
	wire w_dff_A_hoSnWOJF9_0;
	wire w_dff_A_M1pWkXlx1_0;
	wire w_dff_A_XEpaEkmy8_0;
	wire w_dff_A_iLf9I2Gs5_0;
	wire w_dff_A_9YUT2xh85_0;
	wire w_dff_A_6ako0U6V3_0;
	wire w_dff_A_jXzzJuGt6_0;
	wire w_dff_A_y0Az1ZHM7_0;
	wire w_dff_A_IT8zjJY29_0;
	wire w_dff_A_UCtd2EQc3_0;
	wire w_dff_A_kWJYUDkj6_2;
	wire w_dff_A_YMmS6L9s1_1;
	wire w_dff_A_smhmllAO2_1;
	wire w_dff_A_zFmTtjw79_0;
	wire w_dff_A_AuvSAvHW6_0;
	wire w_dff_A_YZJPXvwV8_0;
	wire w_dff_A_ObWUNuaj5_0;
	wire w_dff_A_jFmNtVyD2_0;
	wire w_dff_A_uVJug44B3_0;
	wire w_dff_A_O4VLiglz5_0;
	wire w_dff_A_AkCyC8ka5_0;
	wire w_dff_A_kN6ymnwt2_0;
	wire w_dff_A_MPRMm5fR2_0;
	wire w_dff_A_IKjUIpAw9_0;
	wire w_dff_A_slcVONpW6_0;
	wire w_dff_A_o9s3hDUl8_0;
	wire w_dff_A_n6GAev5Y8_0;
	wire w_dff_A_6GQaVU096_1;
	wire w_dff_A_iUAE4Xef2_0;
	wire w_dff_A_gYmzkazS2_0;
	wire w_dff_A_YiaGsrrI9_0;
	wire w_dff_A_qEcDgUcA5_0;
	wire w_dff_A_pgvuoAmg9_0;
	wire w_dff_A_sLveICmz3_0;
	wire w_dff_A_E3qJyMaQ9_0;
	wire w_dff_A_piWuwKyK9_0;
	wire w_dff_A_vIvjCqFI3_0;
	wire w_dff_A_x4Y6JPWi6_0;
	wire w_dff_A_7Z5JpQnk7_0;
	wire w_dff_A_fOjlT9f56_1;
	wire w_dff_A_L4xYoWA20_1;
	wire w_dff_A_JKeSEgmt2_0;
	wire w_dff_A_0oWuuqk64_0;
	wire w_dff_A_mwKgX20g9_0;
	wire w_dff_A_bZol1qMW1_0;
	wire w_dff_A_M7Eav1Li4_0;
	wire w_dff_A_Uiorhndm8_0;
	wire w_dff_A_vPPoHPEg1_0;
	wire w_dff_A_C0sjlLTX4_0;
	wire w_dff_A_MJ64zJmb7_0;
	wire w_dff_A_LqyqEvkk1_0;
	wire w_dff_B_tDf7LaZP8_3;
	wire w_dff_A_1ci5hxao0_0;
	wire w_dff_A_17BTM5Yb1_0;
	wire w_dff_A_cuQw0M3q5_0;
	wire w_dff_A_uoyEAyqJ2_0;
	wire w_dff_A_JpVJFe6h4_0;
	wire w_dff_A_Ho1MDuCO0_0;
	wire w_dff_A_J9OsFp8x5_0;
	wire w_dff_A_Fqq7HPkV7_0;
	wire w_dff_A_JNmo33VS1_0;
	wire w_dff_A_VTqvuAUF2_0;
	wire w_dff_A_KDlWnTBC2_0;
	wire w_dff_A_7cswBw1t9_0;
	wire w_dff_A_d5GERTO76_0;
	wire w_dff_A_eEk1WIa76_0;
	wire w_dff_A_7C97W6zW1_0;
	wire w_dff_A_DrSQHbmK8_0;
	wire w_dff_A_lErC70C12_0;
	wire w_dff_A_znjD7QcY3_0;
	wire w_dff_A_3ipr91Wf5_0;
	wire w_dff_A_TzPKrYpL1_0;
	wire w_dff_A_AXWvgzbM5_0;
	wire w_dff_A_QxyRqpiz9_0;
	wire w_dff_A_UXNkOvNP1_1;
	wire w_dff_A_eRzFMcPL9_1;
	wire w_dff_A_bfN0Q0R15_1;
	wire w_dff_A_fCpVzSGy4_1;
	wire w_dff_A_BdXfqQ4o7_1;
	wire w_dff_A_u6rrTcFq6_1;
	wire w_dff_A_UuWofEKp8_1;
	wire w_dff_A_yoCtgT8M5_0;
	wire w_dff_A_WkwsjzLT5_0;
	wire w_dff_A_kvNusFHk3_0;
	wire w_dff_A_Bi6OkHbp1_0;
	wire w_dff_A_omCrb17u3_0;
	wire w_dff_A_6ZJLDOnL9_0;
	wire w_dff_A_lQ5MsYHa4_0;
	wire w_dff_A_AoqoFddy4_0;
	wire w_dff_A_Vramqusf3_0;
	wire w_dff_A_ExHkzXRH6_0;
	wire w_dff_A_tBfZmiO65_0;
	wire w_dff_A_SfD5si6v2_0;
	wire w_dff_A_sOCpEAii1_0;
	wire w_dff_B_AaC27EVr9_1;
	wire w_dff_B_rGJeMbm67_1;
	wire w_dff_B_0KLhEgVX2_0;
	wire w_dff_A_FJcUi0DD7_1;
	wire w_dff_A_zOU00Jo50_1;
	wire w_dff_A_uFRrlYmx5_1;
	wire w_dff_A_HNWrLLCV9_1;
	wire w_dff_A_8pJLPnNb8_1;
	wire w_dff_A_lpQKkEot6_1;
	wire w_dff_A_fUfjc2Nt5_1;
	wire w_dff_A_xzjcm0HP9_1;
	wire w_dff_A_pV7U0BwU0_1;
	wire w_dff_A_1StxXajN7_1;
	wire w_dff_A_yJRJj9yl0_1;
	wire w_dff_A_uAcqtmzT1_1;
	wire w_dff_A_CGPkWkbw4_0;
	wire w_dff_A_rxo7xlto1_0;
	wire w_dff_A_VQGxGIqE0_0;
	wire w_dff_A_AMgOlEnP1_0;
	wire w_dff_A_9vKkCo9I6_0;
	wire w_dff_A_gZimZZuF4_0;
	wire w_dff_A_Ze4lYX293_0;
	wire w_dff_A_YADflOyV4_0;
	wire w_dff_A_Jje4ToyZ2_0;
	wire w_dff_A_eyyGZype4_0;
	wire w_dff_A_rvYggMYV9_0;
	wire w_dff_A_4EsmdIrz9_0;
	wire w_dff_A_Kuba5AAk3_0;
	wire w_dff_A_pE3Qa32p8_0;
	wire w_dff_A_6iiqElcM2_0;
	wire w_dff_A_Af1fojlL4_0;
	wire w_dff_A_cl0m71280_0;
	wire w_dff_A_bNj1RzFi8_0;
	wire w_dff_A_iaoM9yXH4_0;
	wire w_dff_A_QrVaYf3R7_0;
	wire w_dff_A_ZaSg8bTT6_0;
	wire w_dff_A_7X63bgxk9_0;
	wire w_dff_A_4yWwIPGb3_1;
	wire w_dff_A_LCBQVhYw9_2;
	wire w_dff_A_8Riq3MXW9_2;
	wire w_dff_A_QulWFVfe7_1;
	wire w_dff_A_LHdbYX1l4_0;
	wire w_dff_A_fgM0rRkI3_0;
	wire w_dff_A_9MRPvmYd4_0;
	wire w_dff_A_thdJSFsO7_0;
	wire w_dff_A_QCy9DNjg5_0;
	wire w_dff_A_xLKU9s3N0_0;
	wire w_dff_A_gigbAQeI1_0;
	wire w_dff_A_y6u6BAZH1_0;
	wire w_dff_A_xxpNAW7v3_0;
	wire w_dff_A_O2cWDeTR9_0;
	wire w_dff_A_qaqcQl2I7_0;
	wire w_dff_A_Hi1Blwi94_0;
	wire w_dff_A_95ypSuxk4_0;
	wire w_dff_A_MWoF7v4d9_0;
	wire w_dff_A_u45MO1NO5_2;
	wire w_dff_B_dBsVMmw73_3;
	wire w_dff_B_n2egPD6k4_3;
	wire w_dff_A_5vbmP3rN7_0;
	wire w_dff_A_r0TRfFGO6_0;
	wire w_dff_A_wwTKFn1p7_0;
	wire w_dff_A_3HY76bT19_0;
	wire w_dff_A_43RCmt4a0_0;
	wire w_dff_A_8BX39smi2_0;
	wire w_dff_A_z8q9eX0b6_0;
	wire w_dff_A_12hBlNlt8_0;
	wire w_dff_A_9CADTxuV0_0;
	wire w_dff_A_BhggG4sV1_0;
	wire w_dff_A_oEciDPoY5_0;
	wire w_dff_A_t0QOJokZ5_1;
	wire w_dff_A_Wk3nflXf8_0;
	wire w_dff_A_AcqzBmno9_0;
	wire w_dff_A_ke57k9Ly9_0;
	wire w_dff_A_JzS1N3x26_0;
	wire w_dff_A_ITmY9NBD9_0;
	wire w_dff_A_CoCJX8gk1_0;
	wire w_dff_A_XuS2VIxY7_0;
	wire w_dff_A_L2ye1Ak59_0;
	wire w_dff_A_NEO4XSwV2_0;
	wire w_dff_A_cKt2JESH7_0;
	wire w_dff_A_jj354q4q8_0;
	wire w_dff_A_wpf09Gme3_0;
	wire w_dff_A_MxM8sEm29_0;
	wire w_dff_A_pEwiFNb82_0;
	wire w_dff_A_MV6gKf3u8_0;
	wire w_dff_A_Kp4fMU0B1_0;
	wire w_dff_A_oeQf53br4_0;
	wire w_dff_A_O1R10r377_0;
	wire w_dff_A_Ux2feFDC8_0;
	wire w_dff_A_B6l5WYiX2_0;
	wire w_dff_A_OZdOeCCq2_0;
	wire w_dff_A_bDdjKQWW9_0;
	wire w_dff_A_Vr5KbPGm8_1;
	wire w_dff_A_JOXvNFby4_0;
	wire w_dff_A_b8WsRpQW0_0;
	wire w_dff_A_WxXg8hHp6_0;
	wire w_dff_A_iqkRzPY84_0;
	wire w_dff_A_CfEJDDX21_2;
	wire w_dff_A_pErA9So75_2;
	wire w_dff_A_2SsQnHsJ0_2;
	wire w_dff_A_3N0rDgif6_2;
	wire w_dff_A_thEhU3rG8_0;
	wire w_dff_A_KuNoHgdm8_0;
	wire w_dff_A_XO2NXqmB5_0;
	wire w_dff_A_YLd838JQ1_0;
	wire w_dff_A_Ejkc2pvE5_0;
	wire w_dff_A_GMhsnH2r1_0;
	wire w_dff_A_kBaZRqQp3_0;
	wire w_dff_A_bq1snYzD8_0;
	wire w_dff_A_UwmH1h3q7_0;
	wire w_dff_A_PeW7kkMH5_0;
	wire w_dff_A_eWqVTP6h1_0;
	wire w_dff_A_Pnx97o5o3_0;
	wire w_dff_A_rTCldChL0_0;
	wire w_dff_A_sJGlKoZN8_0;
	wire w_dff_A_wT9ZA0bX7_0;
	wire w_dff_A_8PN1S7Cr2_0;
	wire w_dff_A_uOmmawTv1_0;
	wire w_dff_A_B1BZUJ931_0;
	wire w_dff_A_ftPwKyxt3_1;
	wire w_dff_A_icqAGQ2x4_1;
	wire w_dff_A_T2uWvyeP3_1;
	wire w_dff_A_9IYsCH6a3_1;
	wire w_dff_A_WDKiYE7a3_1;
	wire w_dff_A_cedgfwoZ5_1;
	wire w_dff_A_4bd6Wsb46_1;
	wire w_dff_B_d5cNMmmd5_3;
	wire w_dff_B_kcAU56Im7_3;
	wire w_dff_B_qMjLyACn1_3;
	wire w_dff_B_54y25HS31_3;
	wire w_dff_B_VJKDBgl72_3;
	wire w_dff_B_xxfKP00E7_3;
	wire w_dff_B_EweI4n6z5_3;
	wire w_dff_B_XGQkjbfn8_3;
	wire w_dff_B_yRcC5K3y6_3;
	wire w_dff_B_dZvAHQZL0_3;
	wire w_dff_B_UxWMeUkp0_3;
	wire w_dff_B_zVYBvw3p7_3;
	wire w_dff_B_bs16xm1N2_3;
	wire w_dff_B_750Cn1Mx1_3;
	wire w_dff_B_GJGTG1B15_3;
	wire w_dff_B_kDrnVLV79_3;
	wire w_dff_A_NVfBsJ6J2_0;
	wire w_dff_A_Z6XOJmfD6_0;
	wire w_dff_A_T6Iee2yQ4_0;
	wire w_dff_A_6TPWwDut0_0;
	wire w_dff_A_nDZu8GlS8_0;
	wire w_dff_A_R4IHslOi1_0;
	wire w_dff_A_dMTdSJT36_0;
	wire w_dff_A_T0rZJ28S7_0;
	wire w_dff_A_u1sl0uzd4_0;
	wire w_dff_A_grOjI92V3_0;
	wire w_dff_A_Z0LdavpV1_0;
	wire w_dff_A_9n1cGunY0_0;
	wire w_dff_A_AG6TQukn0_0;
	wire w_dff_A_6g4UUk1S4_0;
	wire w_dff_A_d9VMHloT7_0;
	wire w_dff_A_otwmZ7K66_1;
	wire w_dff_A_XsjyPbYo6_1;
	wire w_dff_A_aYCwG2i71_1;
	wire w_dff_A_n4rZm2Bp4_1;
	wire w_dff_A_eLjLWaAs6_1;
	wire w_dff_A_eeTzjEih8_1;
	wire w_dff_A_SpqyoD0C9_1;
	wire w_dff_A_xzVgzlMI9_1;
	wire w_dff_A_Kc3zzDO38_1;
	wire w_dff_A_uZmpMZ9T5_1;
	wire w_dff_A_2YidaYvC5_1;
	wire w_dff_A_gqVlawb97_1;
	wire w_dff_A_pc9L0pIi1_2;
	wire w_dff_A_eGx7f1Q51_2;
	wire w_dff_A_3DpWNDEr5_2;
	wire w_dff_A_PYxBVZhx8_2;
	wire w_dff_A_p2xDHb3t4_2;
	wire w_dff_A_AnDg3IFC8_2;
	wire w_dff_A_q927HUSt8_2;
	wire w_dff_A_clbAaZkK8_2;
	wire w_dff_A_k2eO1p883_2;
	wire w_dff_A_drC8dM9f7_2;
	wire w_dff_A_znWjcgch0_2;
	wire w_dff_A_UAAT1bQg5_2;
	wire w_dff_A_j2jZPvdg0_2;
	wire w_dff_A_DOKlR9un6_2;
	wire w_dff_A_UYh1kpDt7_2;
	wire w_dff_A_wfDsTIBL0_1;
	wire w_dff_A_USSvfxsm4_1;
	wire w_dff_A_V0WXk8xn0_1;
	wire w_dff_A_ZXve7Bzx4_1;
	wire w_dff_A_7gqzoWAo3_1;
	wire w_dff_A_rRFgyQ5h6_1;
	wire w_dff_A_ldKU0D3X9_1;
	wire w_dff_A_YmuNw9wL0_1;
	wire w_dff_A_gkfyMVve2_1;
	wire w_dff_A_szKKgWPo3_1;
	wire w_dff_A_QVy1HCwZ0_1;
	wire w_dff_A_SkXrW8Wj2_1;
	wire w_dff_A_hFdfcENc6_1;
	wire w_dff_A_UR7pucAm7_1;
	wire w_dff_A_pLDUt66Z5_1;
	wire w_dff_A_V0Gna0CB6_1;
	wire w_dff_A_AiE7RKGB3_2;
	wire w_dff_B_ncci2Lg17_3;
	wire w_dff_A_rf43yoJL4_2;
	wire w_dff_A_DqQ4FdOr5_0;
	wire w_dff_A_t3mlupzd6_0;
	wire w_dff_A_JjbYlYQx7_0;
	wire w_dff_A_rf9kPEQr9_0;
	wire w_dff_A_dDZMe9FQ2_0;
	wire w_dff_A_tDd1w2bm6_0;
	wire w_dff_A_vK3rWXzI0_0;
	wire w_dff_A_lBuhumSC3_2;
	wire w_dff_A_HSJIbGkF4_0;
	wire w_dff_A_VG4lcelf3_0;
	wire w_dff_A_lCnSg9Uv6_0;
	wire w_dff_A_jG2CR8sJ8_0;
	wire w_dff_A_e7giKlnW0_0;
	wire w_dff_A_PEIkaqYm5_0;
	wire w_dff_A_458vZjmV1_0;
	wire w_dff_A_eO18hD5z1_2;
	wire w_dff_A_3kPMnGYT1_0;
	wire w_dff_A_JdYBryj15_0;
	wire w_dff_A_3lUjyb5F3_0;
	wire w_dff_A_wO15XS5a6_0;
	wire w_dff_A_H9S3Zmtk7_0;
	wire w_dff_A_YgWnHk5c8_0;
	wire w_dff_A_JsurAuWB6_0;
	wire w_dff_A_hoBHkjw44_2;
	wire w_dff_A_wdBsn0Ip9_0;
	wire w_dff_A_F9Cz8fkK3_0;
	wire w_dff_A_NM8ne8bv0_0;
	wire w_dff_A_zFFE9N1h1_0;
	wire w_dff_A_4TIpI5nb8_0;
	wire w_dff_A_ftOWdplm3_0;
	wire w_dff_A_nnWLkqy59_0;
	wire w_dff_A_lNq4Cyh81_2;
	wire w_dff_A_8qfaC76O3_0;
	wire w_dff_A_0WwlKeNZ8_0;
	wire w_dff_A_gAiXq8Ze1_0;
	wire w_dff_A_HoAwywnQ6_0;
	wire w_dff_A_yFi0bW4o3_0;
	wire w_dff_A_KuEGRZOL1_0;
	wire w_dff_A_mAnqE5Dy1_0;
	wire w_dff_A_hj6neaL13_2;
	wire w_dff_A_BBVzFjDh6_0;
	wire w_dff_A_fH3JpKnj3_0;
	wire w_dff_A_p7xXiNuJ6_0;
	wire w_dff_A_pLoShYLs1_0;
	wire w_dff_A_KJEoonuq8_0;
	wire w_dff_A_zxFSqyT41_0;
	wire w_dff_A_QtOGY8Mz7_0;
	wire w_dff_A_MQKByHQh7_2;
	wire w_dff_A_3N4nzonT5_0;
	wire w_dff_A_ZOX2T6Mi3_0;
	wire w_dff_A_izmajK9o8_0;
	wire w_dff_A_4CbT9viI2_0;
	wire w_dff_A_6rRrLFjN5_0;
	wire w_dff_A_Oan4keWR6_0;
	wire w_dff_A_QCf0hqno0_0;
	wire w_dff_A_v8v81gOu0_2;
	wire w_dff_A_uVsynPQB4_0;
	wire w_dff_A_pQx3iepF6_0;
	wire w_dff_A_dS6OrFo16_0;
	wire w_dff_A_Gbngxas66_0;
	wire w_dff_A_MDJKZ6ik6_0;
	wire w_dff_A_Kf98beXv8_0;
	wire w_dff_A_VU2Bv5dh1_0;
	wire w_dff_A_6MMl4RMX9_2;
	wire w_dff_A_slnGxkdR8_0;
	wire w_dff_A_9Y4jb4jo2_0;
	wire w_dff_A_PYGZro3Y9_0;
	wire w_dff_A_nGIw7NVE4_0;
	wire w_dff_A_SHB0QNEh5_0;
	wire w_dff_A_vJZ8BV4y7_0;
	wire w_dff_A_7ppUnfnZ6_0;
	wire w_dff_A_I5xO0wr80_2;
	wire w_dff_A_fiHvYHbj9_0;
	wire w_dff_A_E0yHZl4K6_0;
	wire w_dff_A_QgpErsWx5_0;
	wire w_dff_A_WojpYgxi1_0;
	wire w_dff_A_Ka24iUkt3_0;
	wire w_dff_A_NQhAoMm50_0;
	wire w_dff_A_otYwzOBX0_0;
	wire w_dff_A_7zomEpPc3_2;
	wire w_dff_A_qBVdfWZF1_0;
	wire w_dff_A_PYZ2zXnr3_0;
	wire w_dff_A_O9PQebAI8_0;
	wire w_dff_A_PI1MS8eu2_0;
	wire w_dff_A_ar1DRlSm3_0;
	wire w_dff_A_5Yzf6ebd2_0;
	wire w_dff_A_4wG7pdcN0_2;
	wire w_dff_A_53SmPLCM5_0;
	wire w_dff_A_HdiAkpbs7_0;
	wire w_dff_A_TXwxBMh17_0;
	wire w_dff_A_DB8V6ybq5_0;
	wire w_dff_A_p6fKBKuC0_0;
	wire w_dff_A_KyKqygUl2_0;
	wire w_dff_A_5nmiEcia7_0;
	wire w_dff_A_FHZ9zkzZ5_2;
	wire w_dff_A_68mMAGHY6_0;
	wire w_dff_A_ynUaYUQm2_0;
	wire w_dff_A_2SHu7Z7z8_0;
	wire w_dff_A_JDMIB01L9_0;
	wire w_dff_A_wJq8yI2Z8_0;
	wire w_dff_A_H1H5ZwiN7_0;
	wire w_dff_A_SAZMZT7I1_0;
	wire w_dff_A_owRIK1eH7_2;
	wire w_dff_A_kYODZ5Ae6_0;
	wire w_dff_A_UC56cU1K0_0;
	wire w_dff_A_GyP6ThQA8_0;
	wire w_dff_A_p9cqZigD0_0;
	wire w_dff_A_74Ag3JT38_0;
	wire w_dff_A_dvQRztiP1_0;
	wire w_dff_A_KiD3spGf3_0;
	wire w_dff_A_0SkdKhgQ2_2;
	wire w_dff_A_YigTklAD3_0;
	wire w_dff_A_qPs5LhP03_0;
	wire w_dff_A_g3y226p61_0;
	wire w_dff_A_liw3VfIV6_0;
	wire w_dff_A_lO4mnAmy2_0;
	wire w_dff_A_3VkCP3fv2_0;
	wire w_dff_A_svJDJUqM9_0;
	wire w_dff_A_4ZmVwtxX9_2;
	wire w_dff_A_DKLUyJIk1_0;
	wire w_dff_A_e5097vWo3_0;
	wire w_dff_A_krmH0raQ6_0;
	wire w_dff_A_nBDoDcUE8_0;
	wire w_dff_A_bC1GMlB05_0;
	wire w_dff_A_QALXnU1B0_0;
	wire w_dff_A_gGXzisCY3_0;
	wire w_dff_A_FMGvs0En8_2;
	wire w_dff_A_g202tuwu0_2;
	wire w_dff_A_eSfTIwb37_0;
	wire w_dff_A_VvBkGpwi0_2;
	wire w_dff_A_TiRLqdJ76_0;
	wire w_dff_A_IidXqrXl3_2;
	jnot g000(.din(w_G902_3[2]),.dout(n58),.clk(gclk));
	jnot g001(.din(w_G221_0[1]),.dout(n59),.clk(gclk));
	jnot g002(.din(w_G234_1[1]),.dout(n60),.clk(gclk));
	jor g003(.dina(w_G953_2[1]),.dinb(n60),.dout(n61),.clk(gclk));
	jor g004(.dina(n61),.dinb(w_dff_B_MYlh2hkP6_1),.dout(n62),.clk(gclk));
	jnot g005(.din(w_G110_0[2]),.dout(n63),.clk(gclk));
	jxor g006(.dina(w_G119_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jxor g007(.dina(w_dff_B_E2gMzbzZ7_0),.dinb(n62),.dout(n65),.clk(gclk));
	jxor g008(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n66),.clk(gclk));
	jxor g009(.dina(w_n66_0[1]),.dinb(w_G146_0[2]),.dout(n67),.clk(gclk));
	jxor g010(.dina(w_G137_0[2]),.dinb(w_G128_0[2]),.dout(n68),.clk(gclk));
	jxor g011(.dina(w_dff_B_SezSqpel8_0),.dinb(w_n67_0[1]),.dout(n69),.clk(gclk));
	jxor g012(.dina(w_dff_B_fOfk53P32_0),.dinb(n65),.dout(n70),.clk(gclk));
	jand g013(.dina(w_n70_0[1]),.dinb(w_n58_2[2]),.dout(n71),.clk(gclk));
	jand g014(.dina(w_n58_2[1]),.dinb(w_G234_1[0]),.dout(n72),.clk(gclk));
	jnot g015(.din(n72),.dout(n73),.clk(gclk));
	jand g016(.dina(w_n73_0[1]),.dinb(w_G217_0[2]),.dout(n74),.clk(gclk));
	jnot g017(.din(w_n74_0[1]),.dout(n75),.clk(gclk));
	jxor g018(.dina(w_dff_B_gdUnpY1m1_0),.dinb(w_n71_0[1]),.dout(n76),.clk(gclk));
	jxor g019(.dina(w_G143_0[2]),.dinb(w_G128_0[1]),.dout(n77),.clk(gclk));
	jxor g020(.dina(w_n77_0[1]),.dinb(w_G146_0[1]),.dout(n78),.clk(gclk));
	jxor g021(.dina(w_G137_0[1]),.dinb(w_G134_0[2]),.dout(n79),.clk(gclk));
	jxor g022(.dina(n79),.dinb(w_G131_0[2]),.dout(n80),.clk(gclk));
	jxor g023(.dina(n80),.dinb(w_n78_0[1]),.dout(n81),.clk(gclk));
	jnot g024(.din(w_G113_0[2]),.dout(n82),.clk(gclk));
	jxor g025(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g026(.dina(n83),.dinb(n82),.dout(n84),.clk(gclk));
	jnot g027(.din(w_G210_0[2]),.dout(n85),.clk(gclk));
	jor g028(.dina(w_G953_2[0]),.dinb(w_G237_0[2]),.dout(n86),.clk(gclk));
	jor g029(.dina(w_n86_0[1]),.dinb(n85),.dout(n87),.clk(gclk));
	jxor g030(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g031(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g032(.dina(n89),.dinb(w_n81_0[2]),.dout(n90),.clk(gclk));
	jand g033(.dina(w_n90_0[1]),.dinb(w_n58_2[0]),.dout(n91),.clk(gclk));
	jxor g034(.dina(w_n91_0[1]),.dinb(w_G472_0[2]),.dout(n92),.clk(gclk));
	jand g035(.dina(w_n92_1[1]),.dinb(w_n76_1[2]),.dout(n93),.clk(gclk));
	jor g036(.dina(w_G902_3[1]),.dinb(w_G237_0[1]),.dout(n94),.clk(gclk));
	jand g037(.dina(w_n94_0[1]),.dinb(w_G214_0[1]),.dout(n95),.clk(gclk));
	jnot g038(.din(w_n95_1[1]),.dout(n96),.clk(gclk));
	jnot g039(.din(w_G101_0[1]),.dout(n97),.clk(gclk));
	jxor g040(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n98),.clk(gclk));
	jxor g041(.dina(n98),.dinb(n97),.dout(n99),.clk(gclk));
	jxor g042(.dina(w_n99_0[1]),.dinb(w_n84_0[0]),.dout(n100),.clk(gclk));
	jxor g043(.dina(w_G122_1[1]),.dinb(w_G110_0[1]),.dout(n101),.clk(gclk));
	jxor g044(.dina(w_dff_B_tglVqJNZ7_0),.dinb(n100),.dout(n102),.clk(gclk));
	jnot g045(.din(w_G953_1[2]),.dout(n103),.clk(gclk));
	jand g046(.dina(w_n103_3[2]),.dinb(w_G224_0[1]),.dout(n104),.clk(gclk));
	jxor g047(.dina(w_n78_0[0]),.dinb(w_G125_0[1]),.dout(n105),.clk(gclk));
	jxor g048(.dina(n105),.dinb(w_dff_B_OOoXnuC15_1),.dout(n106),.clk(gclk));
	jxor g049(.dina(n106),.dinb(w_n102_0[1]),.dout(n107),.clk(gclk));
	jand g050(.dina(w_n107_0[1]),.dinb(w_n58_1[2]),.dout(n108),.clk(gclk));
	jand g051(.dina(w_n94_0[0]),.dinb(w_G210_0[1]),.dout(n109),.clk(gclk));
	jxor g052(.dina(w_n109_0[1]),.dinb(w_n108_0[1]),.dout(n110),.clk(gclk));
	jand g053(.dina(w_n110_0[1]),.dinb(w_n96_0[2]),.dout(n111),.clk(gclk));
	jand g054(.dina(w_n73_0[0]),.dinb(w_G221_0[0]),.dout(n112),.clk(gclk));
	jnot g055(.din(w_n112_1[1]),.dout(n113),.clk(gclk));
	jand g056(.dina(w_n103_3[1]),.dinb(w_G227_0[1]),.dout(n114),.clk(gclk));
	jxor g057(.dina(w_G140_0[1]),.dinb(w_n63_0[0]),.dout(n115),.clk(gclk));
	jxor g058(.dina(n115),.dinb(n114),.dout(n116),.clk(gclk));
	jxor g059(.dina(n116),.dinb(w_n99_0[0]),.dout(n117),.clk(gclk));
	jxor g060(.dina(n117),.dinb(w_n81_0[1]),.dout(n118),.clk(gclk));
	jand g061(.dina(w_n118_0[1]),.dinb(w_n58_1[1]),.dout(n119),.clk(gclk));
	jxor g062(.dina(w_n119_0[1]),.dinb(w_G469_0[2]),.dout(n120),.clk(gclk));
	jand g063(.dina(w_n120_0[1]),.dinb(w_n113_0[2]),.dout(n121),.clk(gclk));
	jand g064(.dina(w_n121_0[1]),.dinb(w_n111_0[1]),.dout(n122),.clk(gclk));
	jor g065(.dina(w_n103_3[0]),.dinb(w_G898_0[1]),.dout(n123),.clk(gclk));
	jnot g066(.din(n123),.dout(n124),.clk(gclk));
	jand g067(.dina(w_G237_0[0]),.dinb(w_G234_0[2]),.dout(n125),.clk(gclk));
	jnot g068(.din(n125),.dout(n126),.clk(gclk));
	jand g069(.dina(w_n126_0[1]),.dinb(w_G902_3[0]),.dout(n127),.clk(gclk));
	jand g070(.dina(w_n127_0[1]),.dinb(w_n124_0[1]),.dout(n128),.clk(gclk));
	jand g071(.dina(w_n126_0[0]),.dinb(w_G952_0[2]),.dout(n129),.clk(gclk));
	jand g072(.dina(n129),.dinb(w_n103_2[2]),.dout(n130),.clk(gclk));
	jor g073(.dina(w_n130_1[1]),.dinb(n128),.dout(n131),.clk(gclk));
	jnot g074(.din(w_G478_0[2]),.dout(n132),.clk(gclk));
	jxor g075(.dina(w_n77_0[0]),.dinb(w_G134_0[1]),.dout(n133),.clk(gclk));
	jand g076(.dina(w_n103_2[1]),.dinb(w_G234_0[1]),.dout(n134),.clk(gclk));
	jand g077(.dina(n134),.dinb(w_G217_0[1]),.dout(n135),.clk(gclk));
	jxor g078(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n136),.clk(gclk));
	jxor g079(.dina(n136),.dinb(w_G107_0[1]),.dout(n137),.clk(gclk));
	jxor g080(.dina(w_dff_B_0KLhEgVX2_0),.dinb(n135),.dout(n138),.clk(gclk));
	jxor g081(.dina(n138),.dinb(w_dff_B_rGJeMbm67_1),.dout(n139),.clk(gclk));
	jand g082(.dina(w_n139_0[1]),.dinb(w_n58_1[0]),.dout(n140),.clk(gclk));
	jxor g083(.dina(w_n140_0[1]),.dinb(w_dff_B_nKMMM2cI3_1),.dout(n141),.clk(gclk));
	jnot g084(.din(w_G475_0[2]),.dout(n142),.clk(gclk));
	jxor g085(.dina(w_G122_0[2]),.dinb(w_G113_0[1]),.dout(n143),.clk(gclk));
	jxor g086(.dina(n143),.dinb(w_G104_0[1]),.dout(n144),.clk(gclk));
	jnot g087(.din(w_G214_0[0]),.dout(n145),.clk(gclk));
	jor g088(.dina(w_n86_0[0]),.dinb(n145),.dout(n146),.clk(gclk));
	jnot g089(.din(w_G131_0[1]),.dout(n147),.clk(gclk));
	jxor g090(.dina(w_G143_0[1]),.dinb(n147),.dout(n148),.clk(gclk));
	jxor g091(.dina(n148),.dinb(n146),.dout(n149),.clk(gclk));
	jxor g092(.dina(n149),.dinb(w_n67_0[0]),.dout(n150),.clk(gclk));
	jxor g093(.dina(n150),.dinb(w_dff_B_RpTxSUap7_1),.dout(n151),.clk(gclk));
	jand g094(.dina(w_n151_0[2]),.dinb(w_n58_0[2]),.dout(n152),.clk(gclk));
	jxor g095(.dina(w_n152_0[1]),.dinb(w_dff_B_Mxv7YFLo4_1),.dout(n153),.clk(gclk));
	jand g096(.dina(w_n153_1[1]),.dinb(w_n141_1[1]),.dout(n154),.clk(gclk));
	jand g097(.dina(w_n154_1[1]),.dinb(w_n131_1[2]),.dout(n155),.clk(gclk));
	jand g098(.dina(w_n155_0[1]),.dinb(w_n122_1[1]),.dout(n156),.clk(gclk));
	jand g099(.dina(w_n156_0[1]),.dinb(w_n93_1[1]),.dout(n157),.clk(gclk));
	jxor g100(.dina(w_n157_0[1]),.dinb(w_G101_0[0]),.dout(w_dff_A_rf43yoJL4_2),.clk(gclk));
	jnot g101(.din(w_G472_0[1]),.dout(n159),.clk(gclk));
	jxor g102(.dina(w_n91_0[0]),.dinb(w_dff_B_oEXkI1vY7_1),.dout(n160),.clk(gclk));
	jand g103(.dina(w_n160_1[2]),.dinb(w_n76_1[1]),.dout(n161),.clk(gclk));
	jand g104(.dina(w_n161_1[1]),.dinb(w_n122_1[0]),.dout(n162),.clk(gclk));
	jxor g105(.dina(w_n152_0[0]),.dinb(w_G475_0[1]),.dout(n163),.clk(gclk));
	jand g106(.dina(w_n163_1[1]),.dinb(w_n141_1[0]),.dout(n164),.clk(gclk));
	jand g107(.dina(w_n164_0[1]),.dinb(w_n131_1[1]),.dout(n165),.clk(gclk));
	jand g108(.dina(w_n165_0[2]),.dinb(w_n162_0[1]),.dout(n166),.clk(gclk));
	jxor g109(.dina(w_n166_0[1]),.dinb(w_G104_0[0]),.dout(w_dff_A_lBuhumSC3_2),.clk(gclk));
	jxor g110(.dina(w_n140_0[0]),.dinb(w_G478_0[1]),.dout(n168),.clk(gclk));
	jand g111(.dina(w_n153_1[0]),.dinb(w_n168_1[1]),.dout(n169),.clk(gclk));
	jand g112(.dina(w_n169_0[1]),.dinb(w_n131_1[0]),.dout(n170),.clk(gclk));
	jand g113(.dina(w_n170_0[1]),.dinb(w_n162_0[0]),.dout(n171),.clk(gclk));
	jxor g114(.dina(w_n171_0[1]),.dinb(w_G107_0[0]),.dout(w_dff_A_eO18hD5z1_2),.clk(gclk));
	jxor g115(.dina(w_n74_0[0]),.dinb(w_n71_0[0]),.dout(n173),.clk(gclk));
	jand g116(.dina(w_n160_1[1]),.dinb(w_n173_1[1]),.dout(n174),.clk(gclk));
	jand g117(.dina(w_n174_0[1]),.dinb(w_n156_0[0]),.dout(n175),.clk(gclk));
	jxor g118(.dina(w_n175_0[1]),.dinb(w_G110_0[0]),.dout(w_dff_A_hoBHkjw44_2),.clk(gclk));
	jand g119(.dina(w_n92_1[0]),.dinb(w_n173_1[0]),.dout(n177),.clk(gclk));
	jand g120(.dina(w_n177_0[2]),.dinb(w_n122_0[2]),.dout(n178),.clk(gclk));
	jor g121(.dina(w_n103_2[0]),.dinb(w_G900_0[1]),.dout(n179),.clk(gclk));
	jnot g122(.din(n179),.dout(n180),.clk(gclk));
	jand g123(.dina(w_n180_0[1]),.dinb(w_n127_0[0]),.dout(n181),.clk(gclk));
	jor g124(.dina(n181),.dinb(w_n130_1[0]),.dout(n182),.clk(gclk));
	jand g125(.dina(w_n182_1[2]),.dinb(w_n169_0[0]),.dout(n183),.clk(gclk));
	jand g126(.dina(w_n183_0[2]),.dinb(w_n178_0[1]),.dout(n184),.clk(gclk));
	jxor g127(.dina(w_n184_0[1]),.dinb(w_G128_0[0]),.dout(w_dff_A_lNq4Cyh81_2),.clk(gclk));
	jand g128(.dina(w_n163_1[0]),.dinb(w_n168_1[0]),.dout(n186),.clk(gclk));
	jand g129(.dina(w_n186_0[1]),.dinb(w_n93_1[0]),.dout(n187),.clk(gclk));
	jand g130(.dina(n187),.dinb(w_n182_1[1]),.dout(n188),.clk(gclk));
	jand g131(.dina(n188),.dinb(w_n122_0[1]),.dout(n189),.clk(gclk));
	jxor g132(.dina(w_n189_0[1]),.dinb(w_G143_0[0]),.dout(w_dff_A_hj6neaL13_2),.clk(gclk));
	jand g133(.dina(w_n182_1[0]),.dinb(w_n164_0[0]),.dout(n191),.clk(gclk));
	jand g134(.dina(w_n191_0[2]),.dinb(w_n178_0[0]),.dout(n192),.clk(gclk));
	jxor g135(.dina(w_n192_0[2]),.dinb(w_G146_0[0]),.dout(w_dff_A_MQKByHQh7_2),.clk(gclk));
	jnot g136(.din(w_G469_0[1]),.dout(n194),.clk(gclk));
	jxor g137(.dina(w_n119_0[0]),.dinb(w_dff_B_EZajK4Zx4_1),.dout(n195),.clk(gclk));
	jand g138(.dina(w_n195_0[2]),.dinb(w_n113_0[1]),.dout(n196),.clk(gclk));
	jand g139(.dina(n196),.dinb(w_n111_0[0]),.dout(n197),.clk(gclk));
	jand g140(.dina(w_n197_1[1]),.dinb(w_n93_0[2]),.dout(n198),.clk(gclk));
	jand g141(.dina(w_n198_0[1]),.dinb(w_n165_0[1]),.dout(n199),.clk(gclk));
	jxor g142(.dina(w_n199_0[2]),.dinb(w_G113_0[0]),.dout(w_dff_A_v8v81gOu0_2),.clk(gclk));
	jand g143(.dina(w_n198_0[0]),.dinb(w_n170_0[0]),.dout(n201),.clk(gclk));
	jxor g144(.dina(w_n201_0[1]),.dinb(w_G116_0[0]),.dout(w_dff_A_6MMl4RMX9_2),.clk(gclk));
	jand g145(.dina(w_n177_0[1]),.dinb(w_n155_0[0]),.dout(n203),.clk(gclk));
	jand g146(.dina(n203),.dinb(w_n197_1[0]),.dout(n204),.clk(gclk));
	jxor g147(.dina(w_n204_0[1]),.dinb(w_G119_0[0]),.dout(w_dff_A_I5xO0wr80_2),.clk(gclk));
	jand g148(.dina(w_n197_0[2]),.dinb(w_n161_1[0]),.dout(n206),.clk(gclk));
	jand g149(.dina(w_n206_0[1]),.dinb(w_n131_0[2]),.dout(n207),.clk(gclk));
	jand g150(.dina(n207),.dinb(w_n186_0[0]),.dout(n208),.clk(gclk));
	jxor g151(.dina(w_n208_0[1]),.dinb(w_G122_0[1]),.dout(w_dff_A_7zomEpPc3_2),.clk(gclk));
	jand g152(.dina(w_n191_0[1]),.dinb(w_n174_0[0]),.dout(n210),.clk(gclk));
	jand g153(.dina(w_n210_0[1]),.dinb(w_n197_0[1]),.dout(n211),.clk(gclk));
	jxor g154(.dina(w_n211_0[1]),.dinb(w_G125_0[0]),.dout(w_dff_A_4wG7pdcN0_2),.clk(gclk));
	jnot g155(.din(w_n109_0[0]),.dout(n213),.clk(gclk));
	jxor g156(.dina(w_dff_B_9Vd1GOLh7_0),.dinb(w_n108_0[0]),.dout(n214),.clk(gclk));
	jand g157(.dina(w_n214_0[2]),.dinb(w_n96_0[1]),.dout(n215),.clk(gclk));
	jand g158(.dina(n215),.dinb(w_n121_0[0]),.dout(n216),.clk(gclk));
	jand g159(.dina(w_n216_1[1]),.dinb(w_n93_0[1]),.dout(n217),.clk(gclk));
	jand g160(.dina(w_n217_0[1]),.dinb(w_n191_0[0]),.dout(n218),.clk(gclk));
	jxor g161(.dina(w_n218_0[1]),.dinb(w_G131_0[0]),.dout(w_dff_A_FHZ9zkzZ5_2),.clk(gclk));
	jand g162(.dina(w_n217_0[0]),.dinb(w_n183_0[1]),.dout(n220),.clk(gclk));
	jxor g163(.dina(w_n220_0[1]),.dinb(w_G134_0[0]),.dout(w_dff_A_owRIK1eH7_2),.clk(gclk));
	jand g164(.dina(w_n177_0[0]),.dinb(w_n154_1[0]),.dout(n222),.clk(gclk));
	jand g165(.dina(n222),.dinb(w_n182_0[2]),.dout(n223),.clk(gclk));
	jand g166(.dina(n223),.dinb(w_n216_1[0]),.dout(n224),.clk(gclk));
	jxor g167(.dina(w_n224_0[1]),.dinb(w_G137_0[0]),.dout(w_dff_A_0SkdKhgQ2_2),.clk(gclk));
	jand g168(.dina(w_n216_0[2]),.dinb(w_n210_0[0]),.dout(n226),.clk(gclk));
	jxor g169(.dina(w_n226_0[1]),.dinb(w_G140_0[0]),.dout(w_dff_A_4ZmVwtxX9_2),.clk(gclk));
	jor g170(.dina(w_n171_0[0]),.dinb(w_n157_0[0]),.dout(n228),.clk(gclk));
	jor g171(.dina(n228),.dinb(w_n166_0[0]),.dout(n229),.clk(gclk));
	jor g172(.dina(n229),.dinb(w_n208_0[0]),.dout(n230),.clk(gclk));
	jor g173(.dina(w_n204_0[0]),.dinb(w_n201_0[0]),.dout(n231),.clk(gclk));
	jor g174(.dina(n231),.dinb(w_n175_0[0]),.dout(n232),.clk(gclk));
	jor g175(.dina(n232),.dinb(w_n199_0[1]),.dout(n233),.clk(gclk));
	jor g176(.dina(n233),.dinb(n230),.dout(n234),.clk(gclk));
	jor g177(.dina(w_n226_0[0]),.dinb(w_n224_0[0]),.dout(n235),.clk(gclk));
	jor g178(.dina(n235),.dinb(w_n192_0[1]),.dout(n236),.clk(gclk));
	jor g179(.dina(w_n220_0[0]),.dinb(w_n218_0[0]),.dout(n237),.clk(gclk));
	jor g180(.dina(w_n211_0[0]),.dinb(w_n189_0[0]),.dout(n238),.clk(gclk));
	jor g181(.dina(n238),.dinb(w_n184_0[0]),.dout(n239),.clk(gclk));
	jor g182(.dina(n239),.dinb(w_dff_B_8bRbkbHo2_1),.dout(n240),.clk(gclk));
	jor g183(.dina(n240),.dinb(w_dff_B_HfhpR8ps8_1),.dout(n241),.clk(gclk));
	jor g184(.dina(n241),.dinb(n234),.dout(n242),.clk(gclk));
	jand g185(.dina(w_n195_0[1]),.dinb(w_n214_0[1]),.dout(n243),.clk(gclk));
	jxor g186(.dina(w_n112_1[0]),.dinb(w_n95_1[0]),.dout(n244),.clk(gclk));
	jand g187(.dina(w_dff_B_Y7JkvRCC7_0),.dinb(w_n243_0[1]),.dout(n245),.clk(gclk));
	jor g188(.dina(n245),.dinb(w_n216_0[1]),.dout(n246),.clk(gclk));
	jand g189(.dina(n246),.dinb(w_n161_0[2]),.dout(n247),.clk(gclk));
	jand g190(.dina(w_n113_0[0]),.dinb(w_n96_0[0]),.dout(n248),.clk(gclk));
	jand g191(.dina(w_dff_B_rTOt5aZC3_0),.dinb(w_n243_0[0]),.dout(n249),.clk(gclk));
	jxor g192(.dina(w_n160_1[0]),.dinb(w_n76_1[0]),.dout(n250),.clk(gclk));
	jand g193(.dina(w_dff_B_EjutnVrS9_0),.dinb(w_n249_0[1]),.dout(n251),.clk(gclk));
	jor g194(.dina(n251),.dinb(w_n206_0[0]),.dout(n252),.clk(gclk));
	jor g195(.dina(n252),.dinb(n247),.dout(n253),.clk(gclk));
	jand g196(.dina(n253),.dinb(w_n154_0[2]),.dout(n254),.clk(gclk));
	jand g197(.dina(n254),.dinb(w_n130_0[2]),.dout(n255),.clk(gclk));
	jor g198(.dina(w_dff_B_2UGfDtp09_0),.dinb(w_n242_2[2]),.dout(n256),.clk(gclk));
	jand g199(.dina(n256),.dinb(w_G952_0[1]),.dout(n257),.clk(gclk));
	jor g200(.dina(w_n153_0[2]),.dinb(w_n141_0[2]),.dout(n258),.clk(gclk));
	jor g201(.dina(w_n154_0[1]),.dinb(w_n130_0[1]),.dout(n259),.clk(gclk));
	jand g202(.dina(n259),.dinb(w_n258_0[2]),.dout(n260),.clk(gclk));
	jand g203(.dina(n260),.dinb(w_n161_0[1]),.dout(n261),.clk(gclk));
	jand g204(.dina(n261),.dinb(w_n249_0[0]),.dout(n262),.clk(gclk));
	jor g205(.dina(n262),.dinb(w_G953_1[1]),.dout(n263),.clk(gclk));
	jor g206(.dina(w_dff_B_mdhrHRyX3_0),.dinb(n257),.dout(w_dff_A_FMGvs0En8_2),.clk(gclk));
	jor g207(.dina(w_n103_1[2]),.dinb(w_G952_0[0]),.dout(n265),.clk(gclk));
	jand g208(.dina(w_n242_2[1]),.dinb(w_G210_0[0]),.dout(n266),.clk(gclk));
	jand g209(.dina(n266),.dinb(w_G902_2[2]),.dout(n267),.clk(gclk));
	jxor g210(.dina(n267),.dinb(w_n107_0[0]),.dout(n268),.clk(gclk));
	jand g211(.dina(n268),.dinb(w_n265_2[1]),.dout(G51),.clk(gclk));
	jand g212(.dina(w_n242_2[0]),.dinb(w_G469_0[0]),.dout(n270),.clk(gclk));
	jand g213(.dina(n270),.dinb(w_G902_2[1]),.dout(n271),.clk(gclk));
	jxor g214(.dina(n271),.dinb(w_n118_0[0]),.dout(n272),.clk(gclk));
	jand g215(.dina(n272),.dinb(w_n265_2[0]),.dout(G54),.clk(gclk));
	jand g216(.dina(w_G902_2[0]),.dinb(w_G475_0[0]),.dout(n274),.clk(gclk));
	jand g217(.dina(w_n274_0[1]),.dinb(w_n242_1[2]),.dout(n275),.clk(gclk));
	jor g218(.dina(n275),.dinb(w_n151_0[1]),.dout(n276),.clk(gclk));
	jnot g219(.din(w_n151_0[0]),.dout(n277),.clk(gclk));
	jnot g220(.din(w_n131_0[1]),.dout(n278),.clk(gclk));
	jor g221(.dina(w_n92_0[2]),.dinb(w_n173_0[2]),.dout(n279),.clk(gclk));
	jor g222(.dina(w_n214_0[0]),.dinb(w_n95_0[2]),.dout(n280),.clk(gclk));
	jor g223(.dina(w_n120_0[0]),.dinb(w_n112_0[2]),.dout(n281),.clk(gclk));
	jor g224(.dina(n281),.dinb(w_n280_0[1]),.dout(n282),.clk(gclk));
	jor g225(.dina(w_n282_1[1]),.dinb(w_n279_0[1]),.dout(n283),.clk(gclk));
	jor g226(.dina(n283),.dinb(w_n278_0[2]),.dout(n284),.clk(gclk));
	jor g227(.dina(n284),.dinb(w_n258_0[1]),.dout(n285),.clk(gclk));
	jor g228(.dina(w_n195_0[0]),.dinb(w_n112_0[1]),.dout(n286),.clk(gclk));
	jor g229(.dina(w_n286_0[1]),.dinb(w_n280_0[0]),.dout(n287),.clk(gclk));
	jor g230(.dina(w_n279_0[0]),.dinb(w_n287_1[1]),.dout(n288),.clk(gclk));
	jnot g231(.din(w_n165_0[0]),.dout(n289),.clk(gclk));
	jor g232(.dina(n289),.dinb(w_n288_0[1]),.dout(n290),.clk(gclk));
	jor g233(.dina(w_n160_0[2]),.dinb(w_n173_0[1]),.dout(n291),.clk(gclk));
	jor g234(.dina(w_n163_0[2]),.dinb(w_n168_0[2]),.dout(n292),.clk(gclk));
	jor g235(.dina(w_n292_0[1]),.dinb(w_n278_0[1]),.dout(n293),.clk(gclk));
	jor g236(.dina(w_n293_0[1]),.dinb(w_n287_1[0]),.dout(n294),.clk(gclk));
	jor g237(.dina(w_n294_0[1]),.dinb(w_n291_1[1]),.dout(n295),.clk(gclk));
	jor g238(.dina(w_n163_0[1]),.dinb(w_n141_0[1]),.dout(n296),.clk(gclk));
	jor g239(.dina(n296),.dinb(w_n278_0[0]),.dout(n297),.clk(gclk));
	jor g240(.dina(w_n297_0[1]),.dinb(w_n288_0[0]),.dout(n298),.clk(gclk));
	jand g241(.dina(n298),.dinb(n295),.dout(n299),.clk(gclk));
	jand g242(.dina(n299),.dinb(w_dff_B_IBTGc6487_1),.dout(n300),.clk(gclk));
	jand g243(.dina(n300),.dinb(w_dff_B_5rQkiA8U2_1),.dout(n301),.clk(gclk));
	jnot g244(.din(w_n199_0[0]),.dout(n302),.clk(gclk));
	jor g245(.dina(w_n92_0[1]),.dinb(w_n76_0[2]),.dout(n303),.clk(gclk));
	jor g246(.dina(w_n303_0[1]),.dinb(w_n294_0[0]),.dout(n304),.clk(gclk));
	jor g247(.dina(w_n282_1[0]),.dinb(w_n291_1[0]),.dout(n305),.clk(gclk));
	jor g248(.dina(n305),.dinb(w_n297_0[0]),.dout(n306),.clk(gclk));
	jor g249(.dina(w_n160_0[1]),.dinb(w_n76_0[1]),.dout(n307),.clk(gclk));
	jor g250(.dina(w_n307_0[2]),.dinb(w_n293_0[0]),.dout(n308),.clk(gclk));
	jor g251(.dina(n308),.dinb(w_n282_0[2]),.dout(n309),.clk(gclk));
	jand g252(.dina(n309),.dinb(n306),.dout(n310),.clk(gclk));
	jand g253(.dina(n310),.dinb(w_dff_B_XYKnHp0j2_1),.dout(n311),.clk(gclk));
	jand g254(.dina(n311),.dinb(w_dff_B_H0KRGSsn2_1),.dout(n312),.clk(gclk));
	jand g255(.dina(n312),.dinb(n301),.dout(n313),.clk(gclk));
	jnot g256(.din(w_n192_0[0]),.dout(n314),.clk(gclk));
	jor g257(.dina(w_n110_0[0]),.dinb(w_n95_0[1]),.dout(n315),.clk(gclk));
	jor g258(.dina(n315),.dinb(w_n286_0[0]),.dout(n316),.clk(gclk));
	jnot g259(.din(w_n182_0[1]),.dout(n317),.clk(gclk));
	jor g260(.dina(w_n307_0[1]),.dinb(w_n292_0[0]),.dout(n318),.clk(gclk));
	jor g261(.dina(n318),.dinb(w_n317_0[2]),.dout(n319),.clk(gclk));
	jor g262(.dina(n319),.dinb(w_n316_0[2]),.dout(n320),.clk(gclk));
	jor g263(.dina(w_n153_0[1]),.dinb(w_n168_0[1]),.dout(n321),.clk(gclk));
	jor g264(.dina(w_n317_0[1]),.dinb(n321),.dout(n322),.clk(gclk));
	jor g265(.dina(w_n322_0[1]),.dinb(w_n303_0[0]),.dout(n323),.clk(gclk));
	jor g266(.dina(w_n316_0[1]),.dinb(w_n323_0[1]),.dout(n324),.clk(gclk));
	jand g267(.dina(n324),.dinb(n320),.dout(n325),.clk(gclk));
	jand g268(.dina(n325),.dinb(n314),.dout(n326),.clk(gclk));
	jor g269(.dina(w_n316_0[0]),.dinb(w_n291_0[2]),.dout(n327),.clk(gclk));
	jor g270(.dina(w_n327_0[1]),.dinb(w_n322_0[0]),.dout(n328),.clk(gclk));
	jnot g271(.din(w_n183_0[0]),.dout(n329),.clk(gclk));
	jor g272(.dina(w_n327_0[0]),.dinb(w_n329_0[1]),.dout(n330),.clk(gclk));
	jand g273(.dina(n330),.dinb(n328),.dout(n331),.clk(gclk));
	jor g274(.dina(w_n307_0[0]),.dinb(w_n287_0[2]),.dout(n332),.clk(gclk));
	jor g275(.dina(w_n329_0[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jor g276(.dina(w_n258_0[0]),.dinb(w_n291_0[1]),.dout(n334),.clk(gclk));
	jor g277(.dina(n334),.dinb(w_n317_0[0]),.dout(n335),.clk(gclk));
	jor g278(.dina(n335),.dinb(w_n287_0[1]),.dout(n336),.clk(gclk));
	jor g279(.dina(w_n323_0[0]),.dinb(w_n282_0[1]),.dout(n337),.clk(gclk));
	jand g280(.dina(n337),.dinb(n336),.dout(n338),.clk(gclk));
	jand g281(.dina(n338),.dinb(w_dff_B_S6Ympi2H6_1),.dout(n339),.clk(gclk));
	jand g282(.dina(n339),.dinb(w_dff_B_favqS1wC0_1),.dout(n340),.clk(gclk));
	jand g283(.dina(n340),.dinb(w_dff_B_jaVsgVn29_1),.dout(n341),.clk(gclk));
	jand g284(.dina(w_n341_0[1]),.dinb(w_n313_0[1]),.dout(n342),.clk(gclk));
	jnot g285(.din(w_n274_0[0]),.dout(n343),.clk(gclk));
	jor g286(.dina(w_dff_B_xTtMqEP62_0),.dinb(n342),.dout(n344),.clk(gclk));
	jor g287(.dina(n344),.dinb(w_dff_B_Pdmthr8R4_1),.dout(n345),.clk(gclk));
	jand g288(.dina(n345),.dinb(w_n265_1[2]),.dout(n346),.clk(gclk));
	jand g289(.dina(n346),.dinb(w_dff_B_UhkGRgaT1_1),.dout(G60),.clk(gclk));
	jand g290(.dina(w_n242_1[1]),.dinb(w_G478_0[0]),.dout(n348),.clk(gclk));
	jand g291(.dina(n348),.dinb(w_G902_1[2]),.dout(n349),.clk(gclk));
	jxor g292(.dina(n349),.dinb(w_n139_0[0]),.dout(n350),.clk(gclk));
	jand g293(.dina(n350),.dinb(w_n265_1[1]),.dout(G63),.clk(gclk));
	jand g294(.dina(w_n242_1[0]),.dinb(w_G217_0[0]),.dout(n352),.clk(gclk));
	jand g295(.dina(n352),.dinb(w_G902_1[1]),.dout(n353),.clk(gclk));
	jxor g296(.dina(n353),.dinb(w_n70_0[0]),.dout(n354),.clk(gclk));
	jand g297(.dina(n354),.dinb(w_n265_1[0]),.dout(G66),.clk(gclk));
	jor g298(.dina(w_n124_0[0]),.dinb(w_n102_0[0]),.dout(n356),.clk(gclk));
	jor g299(.dina(w_n313_0[0]),.dinb(w_G953_1[0]),.dout(n357),.clk(gclk));
	jand g300(.dina(w_G898_0[0]),.dinb(w_G224_0[0]),.dout(n358),.clk(gclk));
	jor g301(.dina(n358),.dinb(w_n103_1[1]),.dout(n359),.clk(gclk));
	jand g302(.dina(w_dff_B_CT4BKni72_0),.dinb(n357),.dout(n360),.clk(gclk));
	jxor g303(.dina(n360),.dinb(w_dff_B_mm3w6rtw5_1),.dout(w_dff_A_g202tuwu0_2),.clk(gclk));
	jor g304(.dina(w_n341_0[0]),.dinb(w_G953_0[2]),.dout(n362),.clk(gclk));
	jand g305(.dina(w_G900_0[0]),.dinb(w_G227_0[0]),.dout(n363),.clk(gclk));
	jor g306(.dina(n363),.dinb(w_n103_1[0]),.dout(n364),.clk(gclk));
	jand g307(.dina(w_dff_B_XgqYe2sI5_0),.dinb(n362),.dout(n365),.clk(gclk));
	jxor g308(.dina(w_n81_0[0]),.dinb(w_n66_0[0]),.dout(n366),.clk(gclk));
	jor g309(.dina(n366),.dinb(w_n180_0[0]),.dout(n367),.clk(gclk));
	jxor g310(.dina(w_dff_B_pHDAhxtA7_0),.dinb(n365),.dout(w_dff_A_VvBkGpwi0_2),.clk(gclk));
	jand g311(.dina(w_G902_1[0]),.dinb(w_G472_0[0]),.dout(n369),.clk(gclk));
	jand g312(.dina(w_dff_B_iHdfZUwO1_0),.dinb(w_n242_0[2]),.dout(n370),.clk(gclk));
	jxor g313(.dina(n370),.dinb(w_n90_0[0]),.dout(n371),.clk(gclk));
	jand g314(.dina(n371),.dinb(w_n265_0[2]),.dout(w_dff_A_IidXqrXl3_2),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_dff_A_R8YlHE2w3_0),.doutb(w_G101_0[1]),.doutc(w_dff_A_VXWWuc3X5_2),.din(G101));
	jspl3 jspl3_w_G104_0(.douta(w_dff_A_QxyRqpiz9_0),.doutb(w_dff_A_UXNkOvNP1_1),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_dff_A_7X63bgxk9_0),.doutb(w_dff_A_4yWwIPGb3_1),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_dff_A_sEbjAvFW8_0),.doutb(w_G110_0[1]),.doutc(w_G110_0[2]),.din(G110));
	jspl3 jspl3_w_G113_0(.douta(w_dff_A_KDlWnTBC2_0),.doutb(w_G113_0[1]),.doutc(w_G113_0[2]),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_dff_A_rvYggMYV9_0),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_dff_A_I5DHfcvg5_0),.doutb(w_G119_0[1]),.doutc(w_dff_A_0lugVVhC9_2),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_dff_A_uAcqtmzT1_1),.doutc(w_G122_0[2]),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_G122_1[1]),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_dff_A_7Z5JpQnk7_0),.doutb(w_dff_A_L4xYoWA20_1),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_dff_A_jj354q4q8_0),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(G128));
	jspl3 jspl3_w_G131_0(.douta(w_dff_A_UCtd2EQc3_0),.doutb(w_G131_0[1]),.doutc(w_dff_A_kWJYUDkj6_2),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_dff_A_bDdjKQWW9_0),.doutb(w_dff_A_Vr5KbPGm8_1),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_QKqVNlEN5_0),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G140_0(.douta(w_dff_A_n6GAev5Y8_0),.doutb(w_dff_A_6GQaVU096_1),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_dff_A_oEciDPoY5_0),.doutb(w_dff_A_t0QOJokZ5_1),.doutc(w_G143_0[2]),.din(G143));
	jspl3 jspl3_w_G146_0(.douta(w_dff_A_LqyqEvkk1_0),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(w_dff_B_tDf7LaZP8_3));
	jspl3 jspl3_w_G210_0(.douta(w_dff_A_Dvrpoyht9_0),.doutb(w_dff_A_Fnzdoirm6_1),.doutc(w_G210_0[2]),.din(G210));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_dff_A_smhmllAO2_1),.din(G214));
	jspl3 jspl3_w_G217_0(.douta(w_dff_A_MWoF7v4d9_0),.doutb(w_G217_0[1]),.doutc(w_dff_A_u45MO1NO5_2),.din(w_dff_B_n2egPD6k4_3));
	jspl jspl_w_G221_0(.douta(w_dff_A_bfGVxm1p0_0),.doutb(w_G221_0[1]),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_dff_A_wdwqTUD03_1),.din(G224));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_dff_A_PSy1Ef8v9_1),.din(G227));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_dff_A_QulWFVfe7_1),.doutc(w_G234_0[2]),.din(G234));
	jspl jspl_w_G234_1(.douta(w_dff_A_FpyAogCZ2_0),.doutb(w_G234_1[1]),.din(w_G234_0[0]));
	jspl3 jspl3_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.doutc(w_G237_0[2]),.din(G237));
	jspl3 jspl3_w_G469_0(.douta(w_dff_A_Ki5uAwD32_0),.doutb(w_G469_0[1]),.doutc(w_dff_A_Ainhjsqa1_2),.din(G469));
	jspl3 jspl3_w_G472_0(.douta(w_G472_0[0]),.doutb(w_G472_0[1]),.doutc(w_dff_A_ngie6Vjf5_2),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_dff_A_UuWofEKp8_1),.doutc(w_G475_0[2]),.din(G475));
	jspl3 jspl3_w_G478_0(.douta(w_dff_A_B1BZUJ931_0),.doutb(w_dff_A_cedgfwoZ5_1),.doutc(w_G478_0[2]),.din(G478));
	jspl jspl_w_G898_0(.douta(w_G898_0[0]),.doutb(w_dff_A_WgfzuJgN5_1),.din(G898));
	jspl jspl_w_G900_0(.douta(w_G900_0[0]),.doutb(w_dff_A_o5HX76V06_1),.din(G900));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_G902_0[2]),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_dff_A_Xa2aGWVJ7_1),.doutc(w_dff_A_TPWjdESN3_2),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_dff_A_VyTK4dvY7_1),.doutc(w_dff_A_WN7aDri63_2),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_dff_A_KuNoHgdm8_0),.doutb(w_G902_3[1]),.doutc(w_G902_3[2]),.din(w_G902_0[2]));
	jspl3 jspl3_w_G952_0(.douta(w_G952_0[0]),.doutb(w_dff_A_V0Gna0CB6_1),.doutc(w_dff_A_AiE7RKGB3_2),.din(w_dff_B_ncci2Lg17_3));
	jspl3 jspl3_w_G953_0(.douta(w_G953_0[0]),.doutb(w_G953_0[1]),.doutc(w_dff_A_UYh1kpDt7_2),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_dff_A_d9VMHloT7_0),.doutb(w_dff_A_gqVlawb97_1),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl jspl_w_G953_2(.douta(w_G953_2[0]),.doutb(w_dff_A_YMmS6L9s1_1),.din(w_G953_0[1]));
	jspl3 jspl3_w_n58_0(.douta(w_dff_A_iqkRzPY84_0),.doutb(w_n58_0[1]),.doutc(w_dff_A_3N0rDgif6_2),.din(n58));
	jspl3 jspl3_w_n58_1(.douta(w_n58_1[0]),.doutb(w_n58_1[1]),.doutc(w_n58_1[2]),.din(w_n58_0[0]));
	jspl3 jspl3_w_n58_2(.douta(w_dff_A_rQECRfdN9_0),.doutb(w_n58_2[1]),.doutc(w_dff_A_1kggSPbO3_2),.din(w_n58_0[1]));
	jspl jspl_w_n63_0(.douta(w_n63_0[0]),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n66_0(.douta(w_dff_A_YZJPXvwV8_0),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_dff_A_zFmTtjw79_0),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n70_0(.douta(w_dff_A_RtDpuMvy0_0),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n74_0(.douta(w_dff_A_O1ecZPEC7_0),.doutb(w_n74_0[1]),.din(n74));
	jspl3 jspl3_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.doutc(w_n76_0[2]),.din(n76));
	jspl3 jspl3_w_n76_1(.douta(w_n76_1[0]),.doutb(w_n76_1[1]),.doutc(w_n76_1[2]),.din(w_n76_0[0]));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_dff_A_0W73h6m64_1),.doutc(w_dff_A_1jcsAr9G2_2),.din(n81));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_dff_A_DTpVIFKE5_1),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n90_0(.douta(w_dff_A_lDGQmxr08_0),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.din(n91));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n92_1(.douta(w_n92_1[0]),.doutb(w_n92_1[1]),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_dff_A_LhbJ3WDd8_1),.doutc(w_dff_A_OsegNpXQ2_2),.din(n93));
	jspl jspl_w_n93_1(.douta(w_n93_1[0]),.doutb(w_dff_A_gt2VHgWJ4_1),.din(w_n93_0[0]));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n95_0(.douta(w_n95_0[0]),.doutb(w_dff_A_TAIfjDqB5_1),.doutc(w_dff_A_0SNZBjMI2_2),.din(n95));
	jspl jspl_w_n95_1(.douta(w_dff_A_ufFIFDr17_0),.doutb(w_n95_1[1]),.din(w_n95_0[0]));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_dff_A_kiIlB8Vh1_1),.doutc(w_dff_A_H8F0IXdL4_2),.din(w_dff_B_JCHEIWWr5_3));
	jspl jspl_w_n99_0(.douta(w_dff_A_dYQ2sOnO3_0),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n103_1(.douta(w_n103_1[0]),.doutb(w_n103_1[1]),.doutc(w_n103_1[2]),.din(w_n103_0[0]));
	jspl3 jspl3_w_n103_2(.douta(w_n103_2[0]),.doutb(w_n103_2[1]),.doutc(w_dff_A_8Riq3MXW9_2),.din(w_n103_0[1]));
	jspl3 jspl3_w_n103_3(.douta(w_n103_3[0]),.doutb(w_n103_3[1]),.doutc(w_n103_3[2]),.din(w_n103_0[2]));
	jspl jspl_w_n107_0(.douta(w_dff_A_8DSmAR8e6_0),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_dff_A_XXodlFnk5_1),.din(n109));
	jspl jspl_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.din(n110));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_dff_A_szorhQwO6_1),.doutc(w_dff_A_4ZH5GRqy3_2),.din(n112));
	jspl jspl_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_dff_A_pQOq6Uh58_1),.doutc(w_dff_A_glx4b2HU7_2),.din(n113));
	jspl jspl_w_n118_0(.douta(w_dff_A_wqXB6xBt2_0),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_dff_A_BqKbgA812_1),.doutc(w_n122_0[2]),.din(n122));
	jspl jspl_w_n122_1(.douta(w_n122_1[0]),.doutb(w_n122_1[1]),.din(w_n122_0[0]));
	jspl jspl_w_n124_0(.douta(w_dff_A_O9bDVYXm7_0),.doutb(w_n124_0[1]),.din(n124));
	jspl jspl_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.din(n126));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl3 jspl3_w_n130_0(.douta(w_n130_0[0]),.doutb(w_dff_A_yMoIAGfu6_1),.doutc(w_dff_A_EfsTyA2Z4_2),.din(n130));
	jspl jspl_w_n130_1(.douta(w_n130_1[0]),.doutb(w_n130_1[1]),.din(w_n130_0[0]));
	jspl3 jspl3_w_n131_0(.douta(w_dff_A_I8pmQhjl7_0),.doutb(w_n131_0[1]),.doutc(w_dff_A_BGe6APbO8_2),.din(n131));
	jspl3 jspl3_w_n131_1(.douta(w_n131_1[0]),.doutb(w_n131_1[1]),.doutc(w_n131_1[2]),.din(w_n131_0[0]));
	jspl jspl_w_n139_0(.douta(w_dff_A_sOCpEAii1_0),.doutb(w_n139_0[1]),.din(n139));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n141_1(.douta(w_n141_1[0]),.doutb(w_n141_1[1]),.din(w_n141_0[0]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_05lP8yaM7_1),.doutc(w_n151_0[2]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl jspl_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_dff_A_TB3CFVc45_2),.din(n154));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl3 jspl3_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.doutc(w_n160_0[2]),.din(n160));
	jspl3 jspl3_w_n160_1(.douta(w_n160_1[0]),.doutb(w_n160_1[1]),.doutc(w_n160_1[2]),.din(w_n160_0[0]));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_dff_A_4mbwf4eE1_1),.doutc(w_dff_A_Yc2wWo9e0_2),.din(w_dff_B_LUzLjp6Q9_3));
	jspl jspl_w_n161_1(.douta(w_n161_1[0]),.doutb(w_n161_1[1]),.din(w_n161_0[0]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_n163_0[2]),.din(n163));
	jspl jspl_w_n163_1(.douta(w_n163_1[0]),.doutb(w_n163_1[1]),.din(w_n163_0[0]));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_dWLe2s8Q4_1),.doutc(w_dff_A_XBGQncMn4_2),.din(n165));
	jspl jspl_w_n166_0(.douta(w_dff_A_CSeTQGlo6_0),.doutb(w_n166_0[1]),.din(n166));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl jspl_w_n168_1(.douta(w_n168_1[0]),.doutb(w_n168_1[1]),.din(w_n168_0[0]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(w_dff_B_bAL3FZPL7_2));
	jspl jspl_w_n171_0(.douta(w_n171_0[0]),.doutb(w_n171_0[1]),.din(n171));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl jspl_w_n173_1(.douta(w_n173_1[0]),.doutb(w_n173_1[1]),.din(w_n173_0[0]));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_dff_A_H2zQJU8B6_1),.din(w_dff_B_2dksoSKa9_2));
	jspl jspl_w_n175_0(.douta(w_dff_A_Eo3OP6EE2_0),.doutb(w_n175_0[1]),.din(n175));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_dff_A_yuQe9kTT3_1),.doutc(w_dff_A_r82Pybnj4_2),.din(n177));
	jspl jspl_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.din(n178));
	jspl jspl_w_n180_0(.douta(w_dff_A_y3BIuxuQ6_0),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n182_0(.douta(w_dff_A_WL8mdX3K8_0),.doutb(w_n182_0[1]),.doutc(w_dff_A_YoKxsKfO2_2),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_dff_A_QnfWgLoo0_1),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n183_0(.douta(w_n183_0[0]),.doutb(w_dff_A_sdWzoRyN7_1),.doutc(w_dff_A_YL2Miv7Q0_2),.din(n183));
	jspl jspl_w_n184_0(.douta(w_dff_A_nft3XXuY3_0),.doutb(w_n184_0[1]),.din(n184));
	jspl jspl_w_n186_0(.douta(w_dff_A_0S7blAa62_0),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n191_0(.douta(w_dff_A_6H0WDGGA8_0),.doutb(w_n191_0[1]),.doutc(w_dff_A_bCtB2c645_2),.din(n191));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_dff_A_t2ZLaWgT3_1),.doutc(w_n192_0[2]),.din(n192));
	jspl3 jspl3_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.doutc(w_n195_0[2]),.din(n195));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_dff_A_D6wwbt1I7_1),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_dff_A_3UBavrO18_0),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_dff_A_yPIgSjky6_1),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n208_0(.douta(w_dff_A_rQqc1nWU3_0),.doutb(w_n208_0[1]),.din(n208));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.din(n211));
	jspl3 jspl3_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.doutc(w_n214_0[2]),.din(n214));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.doutc(w_dff_A_sehqTj2E5_2),.din(n216));
	jspl jspl_w_n216_1(.douta(w_dff_A_mvYfA7ak6_0),.doutb(w_n216_1[1]),.din(w_n216_0[0]));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl3 jspl3_w_n242_1(.douta(w_n242_1[0]),.doutb(w_n242_1[1]),.doutc(w_n242_1[2]),.din(w_n242_0[0]));
	jspl3 jspl3_w_n242_2(.douta(w_n242_2[0]),.doutb(w_n242_2[1]),.doutc(w_n242_2[2]),.din(w_n242_0[1]));
	jspl jspl_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.din(n243));
	jspl jspl_w_n249_0(.douta(w_dff_A_dSFONKfV8_0),.doutb(w_n249_0[1]),.din(n249));
	jspl3 jspl3_w_n258_0(.douta(w_n258_0[0]),.doutb(w_dff_A_moB27oGJ2_1),.doutc(w_dff_A_MWZ48N6Z3_2),.din(n258));
	jspl3 jspl3_w_n265_0(.douta(w_n265_0[0]),.doutb(w_dff_A_4bd6Wsb46_1),.doutc(w_n265_0[2]),.din(w_dff_B_kDrnVLV79_3));
	jspl3 jspl3_w_n265_1(.douta(w_dff_A_eSyyHdl70_0),.doutb(w_dff_A_ClAuuYEU2_1),.doutc(w_n265_1[2]),.din(w_n265_0[0]));
	jspl jspl_w_n265_2(.douta(w_n265_2[0]),.doutb(w_n265_2[1]),.din(w_n265_0[1]));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_DIdKlfsT9_1),.din(n274));
	jspl3 jspl3_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.doutc(w_dff_A_T9L4824r0_2),.din(w_dff_B_642pIuUB7_3));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(w_dff_B_GBnHB9Zw8_2));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n282_0(.douta(w_n282_0[0]),.doutb(w_dff_A_DEqNbgcH4_1),.doutc(w_dff_A_x6yjkDmP3_2),.din(n282));
	jspl jspl_w_n282_1(.douta(w_n282_1[0]),.doutb(w_n282_1[1]),.din(w_n282_0[0]));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(n286));
	jspl3 jspl3_w_n287_0(.douta(w_n287_0[0]),.doutb(w_dff_A_Ql1RQxrt9_1),.doutc(w_n287_0[2]),.din(n287));
	jspl jspl_w_n287_1(.douta(w_n287_1[0]),.doutb(w_n287_1[1]),.din(w_n287_0[0]));
	jspl jspl_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.din(n288));
	jspl3 jspl3_w_n291_0(.douta(w_dff_A_U0yY5g6B5_0),.doutb(w_n291_0[1]),.doutc(w_dff_A_3bKSKJPS4_2),.din(n291));
	jspl jspl_w_n291_1(.douta(w_n291_1[0]),.doutb(w_dff_A_KyQhiGUQ8_1),.din(w_n291_0[0]));
	jspl jspl_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.din(n292));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n294_0(.douta(w_n294_0[0]),.doutb(w_n294_0[1]),.din(n294));
	jspl jspl_w_n297_0(.douta(w_n297_0[0]),.doutb(w_n297_0[1]),.din(w_dff_B_D7S2f1cO7_2));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_WvrPjgf76_1),.din(w_dff_B_8U3ot9Yd8_2));
	jspl3 jspl3_w_n307_0(.douta(w_dff_A_QwYvSUKV8_0),.doutb(w_n307_0[1]),.doutc(w_dff_A_YwRCZHgK4_2),.din(n307));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n316_0(.douta(w_n316_0[0]),.doutb(w_dff_A_aiYopAbc9_1),.doutc(w_dff_A_4HYK9vc51_2),.din(n316));
	jspl3 jspl3_w_n317_0(.douta(w_dff_A_LnZaJCs82_0),.doutb(w_n317_0[1]),.doutc(w_dff_A_Fxn3f38s5_2),.din(w_dff_B_KSiHxSKO7_3));
	jspl jspl_w_n322_0(.douta(w_dff_A_vRssUqsX6_0),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(n323));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(n327));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n341_0(.douta(w_n341_0[0]),.doutb(w_n341_0[1]),.din(n341));
	jdff dff_B_CdRx2ofj8_0(.din(n263),.dout(w_dff_B_CdRx2ofj8_0),.clk(gclk));
	jdff dff_B_Jofgn1S76_0(.din(w_dff_B_CdRx2ofj8_0),.dout(w_dff_B_Jofgn1S76_0),.clk(gclk));
	jdff dff_B_tSrBdNNg0_0(.din(w_dff_B_Jofgn1S76_0),.dout(w_dff_B_tSrBdNNg0_0),.clk(gclk));
	jdff dff_B_uzJKMgZJ8_0(.din(w_dff_B_tSrBdNNg0_0),.dout(w_dff_B_uzJKMgZJ8_0),.clk(gclk));
	jdff dff_B_mdhrHRyX3_0(.din(w_dff_B_uzJKMgZJ8_0),.dout(w_dff_B_mdhrHRyX3_0),.clk(gclk));
	jdff dff_B_rKkOArAP6_0(.din(n255),.dout(w_dff_B_rKkOArAP6_0),.clk(gclk));
	jdff dff_B_2UGfDtp09_0(.din(w_dff_B_rKkOArAP6_0),.dout(w_dff_B_2UGfDtp09_0),.clk(gclk));
	jdff dff_B_EjutnVrS9_0(.din(n250),.dout(w_dff_B_EjutnVrS9_0),.clk(gclk));
	jdff dff_A_PKCFZb8h0_0(.dout(w_n249_0[0]),.din(w_dff_A_PKCFZb8h0_0),.clk(gclk));
	jdff dff_A_dSFONKfV8_0(.dout(w_dff_A_PKCFZb8h0_0),.din(w_dff_A_dSFONKfV8_0),.clk(gclk));
	jdff dff_B_bWLtcQoM2_0(.din(n248),.dout(w_dff_B_bWLtcQoM2_0),.clk(gclk));
	jdff dff_B_rTOt5aZC3_0(.din(w_dff_B_bWLtcQoM2_0),.dout(w_dff_B_rTOt5aZC3_0),.clk(gclk));
	jdff dff_B_P74BFHHB6_0(.din(n244),.dout(w_dff_B_P74BFHHB6_0),.clk(gclk));
	jdff dff_B_qX0R8aqj3_0(.din(w_dff_B_P74BFHHB6_0),.dout(w_dff_B_qX0R8aqj3_0),.clk(gclk));
	jdff dff_B_Y7JkvRCC7_0(.din(w_dff_B_qX0R8aqj3_0),.dout(w_dff_B_Y7JkvRCC7_0),.clk(gclk));
	jdff dff_B_UhkGRgaT1_1(.din(n276),.dout(w_dff_B_UhkGRgaT1_1),.clk(gclk));
	jdff dff_B_gvI1qoJE5_1(.din(n277),.dout(w_dff_B_gvI1qoJE5_1),.clk(gclk));
	jdff dff_B_Ss4VEQKz8_1(.din(w_dff_B_gvI1qoJE5_1),.dout(w_dff_B_Ss4VEQKz8_1),.clk(gclk));
	jdff dff_B_RoDxmlQO3_1(.din(w_dff_B_Ss4VEQKz8_1),.dout(w_dff_B_RoDxmlQO3_1),.clk(gclk));
	jdff dff_B_noQphQOk8_1(.din(w_dff_B_RoDxmlQO3_1),.dout(w_dff_B_noQphQOk8_1),.clk(gclk));
	jdff dff_B_G6zvj8GB8_1(.din(w_dff_B_noQphQOk8_1),.dout(w_dff_B_G6zvj8GB8_1),.clk(gclk));
	jdff dff_B_33x2tQbN4_1(.din(w_dff_B_G6zvj8GB8_1),.dout(w_dff_B_33x2tQbN4_1),.clk(gclk));
	jdff dff_B_kUGQb4pD9_1(.din(w_dff_B_33x2tQbN4_1),.dout(w_dff_B_kUGQb4pD9_1),.clk(gclk));
	jdff dff_B_SkxkywiX2_1(.din(w_dff_B_kUGQb4pD9_1),.dout(w_dff_B_SkxkywiX2_1),.clk(gclk));
	jdff dff_B_vqkQtcQR0_1(.din(w_dff_B_SkxkywiX2_1),.dout(w_dff_B_vqkQtcQR0_1),.clk(gclk));
	jdff dff_B_GvNAzZn29_1(.din(w_dff_B_vqkQtcQR0_1),.dout(w_dff_B_GvNAzZn29_1),.clk(gclk));
	jdff dff_B_Pdmthr8R4_1(.din(w_dff_B_GvNAzZn29_1),.dout(w_dff_B_Pdmthr8R4_1),.clk(gclk));
	jdff dff_B_E4Ub7aYc9_0(.din(n343),.dout(w_dff_B_E4Ub7aYc9_0),.clk(gclk));
	jdff dff_B_BJZXmpsT4_0(.din(w_dff_B_E4Ub7aYc9_0),.dout(w_dff_B_BJZXmpsT4_0),.clk(gclk));
	jdff dff_B_Rw3IvUap5_0(.din(w_dff_B_BJZXmpsT4_0),.dout(w_dff_B_Rw3IvUap5_0),.clk(gclk));
	jdff dff_B_VQsxdqKi4_0(.din(w_dff_B_Rw3IvUap5_0),.dout(w_dff_B_VQsxdqKi4_0),.clk(gclk));
	jdff dff_B_NAPbsLZ77_0(.din(w_dff_B_VQsxdqKi4_0),.dout(w_dff_B_NAPbsLZ77_0),.clk(gclk));
	jdff dff_B_SNo6lWGV8_0(.din(w_dff_B_NAPbsLZ77_0),.dout(w_dff_B_SNo6lWGV8_0),.clk(gclk));
	jdff dff_B_s02w2U9v6_0(.din(w_dff_B_SNo6lWGV8_0),.dout(w_dff_B_s02w2U9v6_0),.clk(gclk));
	jdff dff_B_lQ3kIVHT5_0(.din(w_dff_B_s02w2U9v6_0),.dout(w_dff_B_lQ3kIVHT5_0),.clk(gclk));
	jdff dff_B_Umxg7UHQ6_0(.din(w_dff_B_lQ3kIVHT5_0),.dout(w_dff_B_Umxg7UHQ6_0),.clk(gclk));
	jdff dff_B_wD9nMmlb6_0(.din(w_dff_B_Umxg7UHQ6_0),.dout(w_dff_B_wD9nMmlb6_0),.clk(gclk));
	jdff dff_B_dMIT6iMI9_0(.din(w_dff_B_wD9nMmlb6_0),.dout(w_dff_B_dMIT6iMI9_0),.clk(gclk));
	jdff dff_B_P7YEjKFB7_0(.din(w_dff_B_dMIT6iMI9_0),.dout(w_dff_B_P7YEjKFB7_0),.clk(gclk));
	jdff dff_B_dEkIWPHf4_0(.din(w_dff_B_P7YEjKFB7_0),.dout(w_dff_B_dEkIWPHf4_0),.clk(gclk));
	jdff dff_B_xTtMqEP62_0(.din(w_dff_B_dEkIWPHf4_0),.dout(w_dff_B_xTtMqEP62_0),.clk(gclk));
	jdff dff_A_01Zlvuku6_1(.dout(w_n274_0[1]),.din(w_dff_A_01Zlvuku6_1),.clk(gclk));
	jdff dff_A_JyQbwjjG5_1(.dout(w_dff_A_01Zlvuku6_1),.din(w_dff_A_JyQbwjjG5_1),.clk(gclk));
	jdff dff_A_RGq2ecjx2_1(.dout(w_dff_A_JyQbwjjG5_1),.din(w_dff_A_RGq2ecjx2_1),.clk(gclk));
	jdff dff_A_BxZUUVZb4_1(.dout(w_dff_A_RGq2ecjx2_1),.din(w_dff_A_BxZUUVZb4_1),.clk(gclk));
	jdff dff_A_BAX7EPEZ4_1(.dout(w_dff_A_BxZUUVZb4_1),.din(w_dff_A_BAX7EPEZ4_1),.clk(gclk));
	jdff dff_A_NiXjGfW73_1(.dout(w_dff_A_BAX7EPEZ4_1),.din(w_dff_A_NiXjGfW73_1),.clk(gclk));
	jdff dff_A_ULNlmOgF4_1(.dout(w_dff_A_NiXjGfW73_1),.din(w_dff_A_ULNlmOgF4_1),.clk(gclk));
	jdff dff_A_IDzbWCqW0_1(.dout(w_dff_A_ULNlmOgF4_1),.din(w_dff_A_IDzbWCqW0_1),.clk(gclk));
	jdff dff_A_Fa6hmuCA7_1(.dout(w_dff_A_IDzbWCqW0_1),.din(w_dff_A_Fa6hmuCA7_1),.clk(gclk));
	jdff dff_A_4FTO6hXT7_1(.dout(w_dff_A_Fa6hmuCA7_1),.din(w_dff_A_4FTO6hXT7_1),.clk(gclk));
	jdff dff_A_2ccFVnGw1_1(.dout(w_dff_A_4FTO6hXT7_1),.din(w_dff_A_2ccFVnGw1_1),.clk(gclk));
	jdff dff_A_9ZosgNHH8_1(.dout(w_dff_A_2ccFVnGw1_1),.din(w_dff_A_9ZosgNHH8_1),.clk(gclk));
	jdff dff_A_W4IyJAAy8_1(.dout(w_dff_A_9ZosgNHH8_1),.din(w_dff_A_W4IyJAAy8_1),.clk(gclk));
	jdff dff_A_46gwKBMl0_1(.dout(w_dff_A_W4IyJAAy8_1),.din(w_dff_A_46gwKBMl0_1),.clk(gclk));
	jdff dff_A_DIdKlfsT9_1(.dout(w_dff_A_46gwKBMl0_1),.din(w_dff_A_DIdKlfsT9_1),.clk(gclk));
	jdff dff_A_Y3wGLXRM6_1(.dout(w_G902_2[1]),.din(w_dff_A_Y3wGLXRM6_1),.clk(gclk));
	jdff dff_A_JgZ3KUDw3_1(.dout(w_dff_A_Y3wGLXRM6_1),.din(w_dff_A_JgZ3KUDw3_1),.clk(gclk));
	jdff dff_A_g9GM441z5_1(.dout(w_dff_A_JgZ3KUDw3_1),.din(w_dff_A_g9GM441z5_1),.clk(gclk));
	jdff dff_A_utWSeLvC1_1(.dout(w_dff_A_g9GM441z5_1),.din(w_dff_A_utWSeLvC1_1),.clk(gclk));
	jdff dff_A_8e7MtCfJ0_1(.dout(w_dff_A_utWSeLvC1_1),.din(w_dff_A_8e7MtCfJ0_1),.clk(gclk));
	jdff dff_A_etSqSXhN7_1(.dout(w_dff_A_8e7MtCfJ0_1),.din(w_dff_A_etSqSXhN7_1),.clk(gclk));
	jdff dff_A_HivJmHxQ4_1(.dout(w_dff_A_etSqSXhN7_1),.din(w_dff_A_HivJmHxQ4_1),.clk(gclk));
	jdff dff_A_scdTvfje6_1(.dout(w_dff_A_HivJmHxQ4_1),.din(w_dff_A_scdTvfje6_1),.clk(gclk));
	jdff dff_A_GGnSifdZ0_1(.dout(w_dff_A_scdTvfje6_1),.din(w_dff_A_GGnSifdZ0_1),.clk(gclk));
	jdff dff_A_iJL4TF6P3_1(.dout(w_dff_A_GGnSifdZ0_1),.din(w_dff_A_iJL4TF6P3_1),.clk(gclk));
	jdff dff_A_6c9bOjaF0_1(.dout(w_dff_A_iJL4TF6P3_1),.din(w_dff_A_6c9bOjaF0_1),.clk(gclk));
	jdff dff_A_6QuDRRlY4_1(.dout(w_dff_A_6c9bOjaF0_1),.din(w_dff_A_6QuDRRlY4_1),.clk(gclk));
	jdff dff_A_LefPmnEp8_1(.dout(w_dff_A_6QuDRRlY4_1),.din(w_dff_A_LefPmnEp8_1),.clk(gclk));
	jdff dff_A_JNikaNm51_1(.dout(w_dff_A_LefPmnEp8_1),.din(w_dff_A_JNikaNm51_1),.clk(gclk));
	jdff dff_A_jg6GCSEe1_1(.dout(w_dff_A_JNikaNm51_1),.din(w_dff_A_jg6GCSEe1_1),.clk(gclk));
	jdff dff_A_Xm3ei6mZ7_1(.dout(w_dff_A_jg6GCSEe1_1),.din(w_dff_A_Xm3ei6mZ7_1),.clk(gclk));
	jdff dff_A_VyTK4dvY7_1(.dout(w_dff_A_Xm3ei6mZ7_1),.din(w_dff_A_VyTK4dvY7_1),.clk(gclk));
	jdff dff_A_97odHxbd8_2(.dout(w_G902_2[2]),.din(w_dff_A_97odHxbd8_2),.clk(gclk));
	jdff dff_A_1geQscUf2_2(.dout(w_dff_A_97odHxbd8_2),.din(w_dff_A_1geQscUf2_2),.clk(gclk));
	jdff dff_A_V2qqzgfI7_2(.dout(w_dff_A_1geQscUf2_2),.din(w_dff_A_V2qqzgfI7_2),.clk(gclk));
	jdff dff_A_IEObQtub7_2(.dout(w_dff_A_V2qqzgfI7_2),.din(w_dff_A_IEObQtub7_2),.clk(gclk));
	jdff dff_A_z0XG4Ye59_2(.dout(w_dff_A_IEObQtub7_2),.din(w_dff_A_z0XG4Ye59_2),.clk(gclk));
	jdff dff_A_M7usmQGk8_2(.dout(w_dff_A_z0XG4Ye59_2),.din(w_dff_A_M7usmQGk8_2),.clk(gclk));
	jdff dff_A_0nY5riSl9_2(.dout(w_dff_A_M7usmQGk8_2),.din(w_dff_A_0nY5riSl9_2),.clk(gclk));
	jdff dff_A_krg8bAKb9_2(.dout(w_dff_A_0nY5riSl9_2),.din(w_dff_A_krg8bAKb9_2),.clk(gclk));
	jdff dff_A_raRC3OMP1_2(.dout(w_dff_A_krg8bAKb9_2),.din(w_dff_A_raRC3OMP1_2),.clk(gclk));
	jdff dff_A_6WVtgcq52_2(.dout(w_dff_A_raRC3OMP1_2),.din(w_dff_A_6WVtgcq52_2),.clk(gclk));
	jdff dff_A_WxVODHg12_2(.dout(w_dff_A_6WVtgcq52_2),.din(w_dff_A_WxVODHg12_2),.clk(gclk));
	jdff dff_A_rkvpdkLv3_2(.dout(w_dff_A_WxVODHg12_2),.din(w_dff_A_rkvpdkLv3_2),.clk(gclk));
	jdff dff_A_DPq1QHOl5_2(.dout(w_dff_A_rkvpdkLv3_2),.din(w_dff_A_DPq1QHOl5_2),.clk(gclk));
	jdff dff_A_HQ7adru01_2(.dout(w_dff_A_DPq1QHOl5_2),.din(w_dff_A_HQ7adru01_2),.clk(gclk));
	jdff dff_A_RXlS4zgb6_2(.dout(w_dff_A_HQ7adru01_2),.din(w_dff_A_RXlS4zgb6_2),.clk(gclk));
	jdff dff_A_PfNa3u4S7_2(.dout(w_dff_A_RXlS4zgb6_2),.din(w_dff_A_PfNa3u4S7_2),.clk(gclk));
	jdff dff_A_WN7aDri63_2(.dout(w_dff_A_PfNa3u4S7_2),.din(w_dff_A_WN7aDri63_2),.clk(gclk));
	jdff dff_A_eSyyHdl70_0(.dout(w_n265_1[0]),.din(w_dff_A_eSyyHdl70_0),.clk(gclk));
	jdff dff_A_ClAuuYEU2_1(.dout(w_n265_1[1]),.din(w_dff_A_ClAuuYEU2_1),.clk(gclk));
	jdff dff_B_KLwBtMBo5_1(.din(n356),.dout(w_dff_B_KLwBtMBo5_1),.clk(gclk));
	jdff dff_B_Pqzg5Onq1_1(.din(w_dff_B_KLwBtMBo5_1),.dout(w_dff_B_Pqzg5Onq1_1),.clk(gclk));
	jdff dff_B_580wu7Pw4_1(.din(w_dff_B_Pqzg5Onq1_1),.dout(w_dff_B_580wu7Pw4_1),.clk(gclk));
	jdff dff_B_8MBa5YkG5_1(.din(w_dff_B_580wu7Pw4_1),.dout(w_dff_B_8MBa5YkG5_1),.clk(gclk));
	jdff dff_B_jCJcTw8x9_1(.din(w_dff_B_8MBa5YkG5_1),.dout(w_dff_B_jCJcTw8x9_1),.clk(gclk));
	jdff dff_B_mNbCnYs29_1(.din(w_dff_B_jCJcTw8x9_1),.dout(w_dff_B_mNbCnYs29_1),.clk(gclk));
	jdff dff_B_Iu3AWsBL9_1(.din(w_dff_B_mNbCnYs29_1),.dout(w_dff_B_Iu3AWsBL9_1),.clk(gclk));
	jdff dff_B_HhoRgETG3_1(.din(w_dff_B_Iu3AWsBL9_1),.dout(w_dff_B_HhoRgETG3_1),.clk(gclk));
	jdff dff_B_ggwC78Ie4_1(.din(w_dff_B_HhoRgETG3_1),.dout(w_dff_B_ggwC78Ie4_1),.clk(gclk));
	jdff dff_B_kddSgT1I0_1(.din(w_dff_B_ggwC78Ie4_1),.dout(w_dff_B_kddSgT1I0_1),.clk(gclk));
	jdff dff_B_32whL4Fq2_1(.din(w_dff_B_kddSgT1I0_1),.dout(w_dff_B_32whL4Fq2_1),.clk(gclk));
	jdff dff_B_mm3w6rtw5_1(.din(w_dff_B_32whL4Fq2_1),.dout(w_dff_B_mm3w6rtw5_1),.clk(gclk));
	jdff dff_B_sZyVdW0g1_0(.din(n359),.dout(w_dff_B_sZyVdW0g1_0),.clk(gclk));
	jdff dff_B_fwm0Thr30_0(.din(w_dff_B_sZyVdW0g1_0),.dout(w_dff_B_fwm0Thr30_0),.clk(gclk));
	jdff dff_B_WKX6vTOm1_0(.din(w_dff_B_fwm0Thr30_0),.dout(w_dff_B_WKX6vTOm1_0),.clk(gclk));
	jdff dff_B_7jWup1Di6_0(.din(w_dff_B_WKX6vTOm1_0),.dout(w_dff_B_7jWup1Di6_0),.clk(gclk));
	jdff dff_B_r5yi4Ilk2_0(.din(w_dff_B_7jWup1Di6_0),.dout(w_dff_B_r5yi4Ilk2_0),.clk(gclk));
	jdff dff_B_7dfcLZX26_0(.din(w_dff_B_r5yi4Ilk2_0),.dout(w_dff_B_7dfcLZX26_0),.clk(gclk));
	jdff dff_B_3vQk8ReK6_0(.din(w_dff_B_7dfcLZX26_0),.dout(w_dff_B_3vQk8ReK6_0),.clk(gclk));
	jdff dff_B_Nf4iurPA5_0(.din(w_dff_B_3vQk8ReK6_0),.dout(w_dff_B_Nf4iurPA5_0),.clk(gclk));
	jdff dff_B_v0JEP4p01_0(.din(w_dff_B_Nf4iurPA5_0),.dout(w_dff_B_v0JEP4p01_0),.clk(gclk));
	jdff dff_B_G059g5QF4_0(.din(w_dff_B_v0JEP4p01_0),.dout(w_dff_B_G059g5QF4_0),.clk(gclk));
	jdff dff_B_OIzh3tr73_0(.din(w_dff_B_G059g5QF4_0),.dout(w_dff_B_OIzh3tr73_0),.clk(gclk));
	jdff dff_B_qMy3jbYl2_0(.din(w_dff_B_OIzh3tr73_0),.dout(w_dff_B_qMy3jbYl2_0),.clk(gclk));
	jdff dff_B_9igCQlhx5_0(.din(w_dff_B_qMy3jbYl2_0),.dout(w_dff_B_9igCQlhx5_0),.clk(gclk));
	jdff dff_B_CT4BKni72_0(.din(w_dff_B_9igCQlhx5_0),.dout(w_dff_B_CT4BKni72_0),.clk(gclk));
	jdff dff_B_H0KRGSsn2_1(.din(n302),.dout(w_dff_B_H0KRGSsn2_1),.clk(gclk));
	jdff dff_B_XYKnHp0j2_1(.din(n304),.dout(w_dff_B_XYKnHp0j2_1),.clk(gclk));
	jdff dff_B_5rQkiA8U2_1(.din(n285),.dout(w_dff_B_5rQkiA8U2_1),.clk(gclk));
	jdff dff_B_IBTGc6487_1(.din(n290),.dout(w_dff_B_IBTGc6487_1),.clk(gclk));
	jdff dff_B_D7S2f1cO7_2(.din(n297),.dout(w_dff_B_D7S2f1cO7_2),.clk(gclk));
	jdff dff_A_KyQhiGUQ8_1(.dout(w_n291_1[1]),.din(w_dff_A_KyQhiGUQ8_1),.clk(gclk));
	jdff dff_B_GBnHB9Zw8_2(.din(n279),.dout(w_dff_B_GBnHB9Zw8_2),.clk(gclk));
	jdff dff_A_E82yDAXB3_2(.dout(w_n278_0[2]),.din(w_dff_A_E82yDAXB3_2),.clk(gclk));
	jdff dff_A_T9L4824r0_2(.dout(w_dff_A_E82yDAXB3_2),.din(w_dff_A_T9L4824r0_2),.clk(gclk));
	jdff dff_B_ZUyHbJGO8_3(.din(n278),.dout(w_dff_B_ZUyHbJGO8_3),.clk(gclk));
	jdff dff_B_642pIuUB7_3(.din(w_dff_B_ZUyHbJGO8_3),.dout(w_dff_B_642pIuUB7_3),.clk(gclk));
	jdff dff_B_bw6JouIo8_0(.din(n367),.dout(w_dff_B_bw6JouIo8_0),.clk(gclk));
	jdff dff_B_nrGvtlF21_0(.din(w_dff_B_bw6JouIo8_0),.dout(w_dff_B_nrGvtlF21_0),.clk(gclk));
	jdff dff_B_dfrEfNZa3_0(.din(w_dff_B_nrGvtlF21_0),.dout(w_dff_B_dfrEfNZa3_0),.clk(gclk));
	jdff dff_B_85COfi2C0_0(.din(w_dff_B_dfrEfNZa3_0),.dout(w_dff_B_85COfi2C0_0),.clk(gclk));
	jdff dff_B_AHPfHRnc0_0(.din(w_dff_B_85COfi2C0_0),.dout(w_dff_B_AHPfHRnc0_0),.clk(gclk));
	jdff dff_B_3V0w02l23_0(.din(w_dff_B_AHPfHRnc0_0),.dout(w_dff_B_3V0w02l23_0),.clk(gclk));
	jdff dff_B_8LlYVvKp9_0(.din(w_dff_B_3V0w02l23_0),.dout(w_dff_B_8LlYVvKp9_0),.clk(gclk));
	jdff dff_B_Rw29LyWx0_0(.din(w_dff_B_8LlYVvKp9_0),.dout(w_dff_B_Rw29LyWx0_0),.clk(gclk));
	jdff dff_B_qr30Hv1l1_0(.din(w_dff_B_Rw29LyWx0_0),.dout(w_dff_B_qr30Hv1l1_0),.clk(gclk));
	jdff dff_B_lRvMcX6T0_0(.din(w_dff_B_qr30Hv1l1_0),.dout(w_dff_B_lRvMcX6T0_0),.clk(gclk));
	jdff dff_B_xlV9W2jf8_0(.din(w_dff_B_lRvMcX6T0_0),.dout(w_dff_B_xlV9W2jf8_0),.clk(gclk));
	jdff dff_B_pHDAhxtA7_0(.din(w_dff_B_xlV9W2jf8_0),.dout(w_dff_B_pHDAhxtA7_0),.clk(gclk));
	jdff dff_B_yr50cWre3_0(.din(n364),.dout(w_dff_B_yr50cWre3_0),.clk(gclk));
	jdff dff_B_aUCGbcsC7_0(.din(w_dff_B_yr50cWre3_0),.dout(w_dff_B_aUCGbcsC7_0),.clk(gclk));
	jdff dff_B_IcUCqYEo6_0(.din(w_dff_B_aUCGbcsC7_0),.dout(w_dff_B_IcUCqYEo6_0),.clk(gclk));
	jdff dff_B_sJs3Z4DR0_0(.din(w_dff_B_IcUCqYEo6_0),.dout(w_dff_B_sJs3Z4DR0_0),.clk(gclk));
	jdff dff_B_RwsggDky2_0(.din(w_dff_B_sJs3Z4DR0_0),.dout(w_dff_B_RwsggDky2_0),.clk(gclk));
	jdff dff_B_n4RqY0dh1_0(.din(w_dff_B_RwsggDky2_0),.dout(w_dff_B_n4RqY0dh1_0),.clk(gclk));
	jdff dff_B_myFuCQOt5_0(.din(w_dff_B_n4RqY0dh1_0),.dout(w_dff_B_myFuCQOt5_0),.clk(gclk));
	jdff dff_B_O9WwE1F88_0(.din(w_dff_B_myFuCQOt5_0),.dout(w_dff_B_O9WwE1F88_0),.clk(gclk));
	jdff dff_B_qlIthqTp6_0(.din(w_dff_B_O9WwE1F88_0),.dout(w_dff_B_qlIthqTp6_0),.clk(gclk));
	jdff dff_B_G6zDwesT8_0(.din(w_dff_B_qlIthqTp6_0),.dout(w_dff_B_G6zDwesT8_0),.clk(gclk));
	jdff dff_B_kPJIySp34_0(.din(w_dff_B_G6zDwesT8_0),.dout(w_dff_B_kPJIySp34_0),.clk(gclk));
	jdff dff_B_MWH7XePi5_0(.din(w_dff_B_kPJIySp34_0),.dout(w_dff_B_MWH7XePi5_0),.clk(gclk));
	jdff dff_B_FJyLm5td2_0(.din(w_dff_B_MWH7XePi5_0),.dout(w_dff_B_FJyLm5td2_0),.clk(gclk));
	jdff dff_B_XgqYe2sI5_0(.din(w_dff_B_FJyLm5td2_0),.dout(w_dff_B_XgqYe2sI5_0),.clk(gclk));
	jdff dff_B_jaVsgVn29_1(.din(n326),.dout(w_dff_B_jaVsgVn29_1),.clk(gclk));
	jdff dff_B_favqS1wC0_1(.din(n331),.dout(w_dff_B_favqS1wC0_1),.clk(gclk));
	jdff dff_B_S6Ympi2H6_1(.din(n333),.dout(w_dff_B_S6Ympi2H6_1),.clk(gclk));
	jdff dff_A_DEqNbgcH4_1(.dout(w_n282_0[1]),.din(w_dff_A_DEqNbgcH4_1),.clk(gclk));
	jdff dff_A_x6yjkDmP3_2(.dout(w_n282_0[2]),.din(w_dff_A_x6yjkDmP3_2),.clk(gclk));
	jdff dff_A_ZODl5Moa2_1(.dout(w_n258_0[1]),.din(w_dff_A_ZODl5Moa2_1),.clk(gclk));
	jdff dff_A_8refZzbe8_1(.dout(w_dff_A_ZODl5Moa2_1),.din(w_dff_A_8refZzbe8_1),.clk(gclk));
	jdff dff_A_moB27oGJ2_1(.dout(w_dff_A_8refZzbe8_1),.din(w_dff_A_moB27oGJ2_1),.clk(gclk));
	jdff dff_A_MWZ48N6Z3_2(.dout(w_n258_0[2]),.din(w_dff_A_MWZ48N6Z3_2),.clk(gclk));
	jdff dff_A_Ql1RQxrt9_1(.dout(w_n287_0[1]),.din(w_dff_A_Ql1RQxrt9_1),.clk(gclk));
	jdff dff_A_U0yY5g6B5_0(.dout(w_n291_0[0]),.din(w_dff_A_U0yY5g6B5_0),.clk(gclk));
	jdff dff_A_3bKSKJPS4_2(.dout(w_n291_0[2]),.din(w_dff_A_3bKSKJPS4_2),.clk(gclk));
	jdff dff_A_vRssUqsX6_0(.dout(w_n322_0[0]),.din(w_dff_A_vRssUqsX6_0),.clk(gclk));
	jdff dff_A_WvrPjgf76_1(.dout(w_n303_0[1]),.din(w_dff_A_WvrPjgf76_1),.clk(gclk));
	jdff dff_B_8U3ot9Yd8_2(.din(n303),.dout(w_dff_B_8U3ot9Yd8_2),.clk(gclk));
	jdff dff_A_QwYvSUKV8_0(.dout(w_n307_0[0]),.din(w_dff_A_QwYvSUKV8_0),.clk(gclk));
	jdff dff_A_YwRCZHgK4_2(.dout(w_n307_0[2]),.din(w_dff_A_YwRCZHgK4_2),.clk(gclk));
	jdff dff_A_LnZaJCs82_0(.dout(w_n317_0[0]),.din(w_dff_A_LnZaJCs82_0),.clk(gclk));
	jdff dff_A_Fxn3f38s5_2(.dout(w_n317_0[2]),.din(w_dff_A_Fxn3f38s5_2),.clk(gclk));
	jdff dff_B_iF8xxByB5_3(.din(n317),.dout(w_dff_B_iF8xxByB5_3),.clk(gclk));
	jdff dff_B_KSiHxSKO7_3(.din(w_dff_B_iF8xxByB5_3),.dout(w_dff_B_KSiHxSKO7_3),.clk(gclk));
	jdff dff_A_aiYopAbc9_1(.dout(w_n316_0[1]),.din(w_dff_A_aiYopAbc9_1),.clk(gclk));
	jdff dff_A_4HYK9vc51_2(.dout(w_n316_0[2]),.din(w_dff_A_4HYK9vc51_2),.clk(gclk));
	jdff dff_B_VMwPWO1d1_0(.din(n369),.dout(w_dff_B_VMwPWO1d1_0),.clk(gclk));
	jdff dff_B_05WJY39F9_0(.din(w_dff_B_VMwPWO1d1_0),.dout(w_dff_B_05WJY39F9_0),.clk(gclk));
	jdff dff_B_F0oEXzHH5_0(.din(w_dff_B_05WJY39F9_0),.dout(w_dff_B_F0oEXzHH5_0),.clk(gclk));
	jdff dff_B_FmogL4Tr6_0(.din(w_dff_B_F0oEXzHH5_0),.dout(w_dff_B_FmogL4Tr6_0),.clk(gclk));
	jdff dff_B_PVEGtvjN1_0(.din(w_dff_B_FmogL4Tr6_0),.dout(w_dff_B_PVEGtvjN1_0),.clk(gclk));
	jdff dff_B_DLzdOQkj4_0(.din(w_dff_B_PVEGtvjN1_0),.dout(w_dff_B_DLzdOQkj4_0),.clk(gclk));
	jdff dff_B_XLT3ylCP2_0(.din(w_dff_B_DLzdOQkj4_0),.dout(w_dff_B_XLT3ylCP2_0),.clk(gclk));
	jdff dff_B_DxleLwwm5_0(.din(w_dff_B_XLT3ylCP2_0),.dout(w_dff_B_DxleLwwm5_0),.clk(gclk));
	jdff dff_B_qnQsVxvs5_0(.din(w_dff_B_DxleLwwm5_0),.dout(w_dff_B_qnQsVxvs5_0),.clk(gclk));
	jdff dff_B_2H44TzEw4_0(.din(w_dff_B_qnQsVxvs5_0),.dout(w_dff_B_2H44TzEw4_0),.clk(gclk));
	jdff dff_B_E2OGXQWx4_0(.din(w_dff_B_2H44TzEw4_0),.dout(w_dff_B_E2OGXQWx4_0),.clk(gclk));
	jdff dff_B_T60XriuG8_0(.din(w_dff_B_E2OGXQWx4_0),.dout(w_dff_B_T60XriuG8_0),.clk(gclk));
	jdff dff_B_dbNB63XD4_0(.din(w_dff_B_T60XriuG8_0),.dout(w_dff_B_dbNB63XD4_0),.clk(gclk));
	jdff dff_B_UcTr2xLm2_0(.din(w_dff_B_dbNB63XD4_0),.dout(w_dff_B_UcTr2xLm2_0),.clk(gclk));
	jdff dff_B_iHdfZUwO1_0(.din(w_dff_B_UcTr2xLm2_0),.dout(w_dff_B_iHdfZUwO1_0),.clk(gclk));
	jdff dff_A_QDdCYJo07_1(.dout(w_G902_1[1]),.din(w_dff_A_QDdCYJo07_1),.clk(gclk));
	jdff dff_A_JRGb2gXD7_1(.dout(w_dff_A_QDdCYJo07_1),.din(w_dff_A_JRGb2gXD7_1),.clk(gclk));
	jdff dff_A_PmhDL7eN5_1(.dout(w_dff_A_JRGb2gXD7_1),.din(w_dff_A_PmhDL7eN5_1),.clk(gclk));
	jdff dff_A_Kr47xTpf5_1(.dout(w_dff_A_PmhDL7eN5_1),.din(w_dff_A_Kr47xTpf5_1),.clk(gclk));
	jdff dff_A_lKPvVncS4_1(.dout(w_dff_A_Kr47xTpf5_1),.din(w_dff_A_lKPvVncS4_1),.clk(gclk));
	jdff dff_A_5q0iiHtL2_1(.dout(w_dff_A_lKPvVncS4_1),.din(w_dff_A_5q0iiHtL2_1),.clk(gclk));
	jdff dff_A_rqkgNDsE1_1(.dout(w_dff_A_5q0iiHtL2_1),.din(w_dff_A_rqkgNDsE1_1),.clk(gclk));
	jdff dff_A_C7DW2jBL0_1(.dout(w_dff_A_rqkgNDsE1_1),.din(w_dff_A_C7DW2jBL0_1),.clk(gclk));
	jdff dff_A_UN8YvMYk7_1(.dout(w_dff_A_C7DW2jBL0_1),.din(w_dff_A_UN8YvMYk7_1),.clk(gclk));
	jdff dff_A_2qnLViUH1_1(.dout(w_dff_A_UN8YvMYk7_1),.din(w_dff_A_2qnLViUH1_1),.clk(gclk));
	jdff dff_A_ZVEVOxHd0_1(.dout(w_dff_A_2qnLViUH1_1),.din(w_dff_A_ZVEVOxHd0_1),.clk(gclk));
	jdff dff_A_fzb2ey0u6_1(.dout(w_dff_A_ZVEVOxHd0_1),.din(w_dff_A_fzb2ey0u6_1),.clk(gclk));
	jdff dff_A_4aRytuxL4_1(.dout(w_dff_A_fzb2ey0u6_1),.din(w_dff_A_4aRytuxL4_1),.clk(gclk));
	jdff dff_A_ayle6BcB5_1(.dout(w_dff_A_4aRytuxL4_1),.din(w_dff_A_ayle6BcB5_1),.clk(gclk));
	jdff dff_A_JKobmPW97_1(.dout(w_dff_A_ayle6BcB5_1),.din(w_dff_A_JKobmPW97_1),.clk(gclk));
	jdff dff_A_b4baawxQ5_1(.dout(w_dff_A_JKobmPW97_1),.din(w_dff_A_b4baawxQ5_1),.clk(gclk));
	jdff dff_A_Xa2aGWVJ7_1(.dout(w_dff_A_b4baawxQ5_1),.din(w_dff_A_Xa2aGWVJ7_1),.clk(gclk));
	jdff dff_A_u7xQmrzd0_2(.dout(w_G902_1[2]),.din(w_dff_A_u7xQmrzd0_2),.clk(gclk));
	jdff dff_A_BipGxom86_2(.dout(w_dff_A_u7xQmrzd0_2),.din(w_dff_A_BipGxom86_2),.clk(gclk));
	jdff dff_A_7MWomFnc0_2(.dout(w_dff_A_BipGxom86_2),.din(w_dff_A_7MWomFnc0_2),.clk(gclk));
	jdff dff_A_aySddW5V9_2(.dout(w_dff_A_7MWomFnc0_2),.din(w_dff_A_aySddW5V9_2),.clk(gclk));
	jdff dff_A_QL6ZRlOf8_2(.dout(w_dff_A_aySddW5V9_2),.din(w_dff_A_QL6ZRlOf8_2),.clk(gclk));
	jdff dff_A_07B2X1Ur5_2(.dout(w_dff_A_QL6ZRlOf8_2),.din(w_dff_A_07B2X1Ur5_2),.clk(gclk));
	jdff dff_A_i60C2Ups4_2(.dout(w_dff_A_07B2X1Ur5_2),.din(w_dff_A_i60C2Ups4_2),.clk(gclk));
	jdff dff_A_Xyp4qGUm3_2(.dout(w_dff_A_i60C2Ups4_2),.din(w_dff_A_Xyp4qGUm3_2),.clk(gclk));
	jdff dff_A_w2vnCVdz4_2(.dout(w_dff_A_Xyp4qGUm3_2),.din(w_dff_A_w2vnCVdz4_2),.clk(gclk));
	jdff dff_A_7Y6mJfUR5_2(.dout(w_dff_A_w2vnCVdz4_2),.din(w_dff_A_7Y6mJfUR5_2),.clk(gclk));
	jdff dff_A_BrrfhQ5v1_2(.dout(w_dff_A_7Y6mJfUR5_2),.din(w_dff_A_BrrfhQ5v1_2),.clk(gclk));
	jdff dff_A_ycwMGVna9_2(.dout(w_dff_A_BrrfhQ5v1_2),.din(w_dff_A_ycwMGVna9_2),.clk(gclk));
	jdff dff_A_eNZWx0B75_2(.dout(w_dff_A_ycwMGVna9_2),.din(w_dff_A_eNZWx0B75_2),.clk(gclk));
	jdff dff_A_jBTPX2LO1_2(.dout(w_dff_A_eNZWx0B75_2),.din(w_dff_A_jBTPX2LO1_2),.clk(gclk));
	jdff dff_A_HFqMOeIh1_2(.dout(w_dff_A_jBTPX2LO1_2),.din(w_dff_A_HFqMOeIh1_2),.clk(gclk));
	jdff dff_A_5z7CCzzn1_2(.dout(w_dff_A_HFqMOeIh1_2),.din(w_dff_A_5z7CCzzn1_2),.clk(gclk));
	jdff dff_A_TPWjdESN3_2(.dout(w_dff_A_5z7CCzzn1_2),.din(w_dff_A_TPWjdESN3_2),.clk(gclk));
	jdff dff_B_HfhpR8ps8_1(.din(n236),.dout(w_dff_B_HfhpR8ps8_1),.clk(gclk));
	jdff dff_B_8bRbkbHo2_1(.din(n237),.dout(w_dff_B_8bRbkbHo2_1),.clk(gclk));
	jdff dff_A_nft3XXuY3_0(.dout(w_n184_0[0]),.din(w_dff_A_nft3XXuY3_0),.clk(gclk));
	jdff dff_A_sdWzoRyN7_1(.dout(w_n183_0[1]),.din(w_dff_A_sdWzoRyN7_1),.clk(gclk));
	jdff dff_A_YL2Miv7Q0_2(.dout(w_n183_0[2]),.din(w_dff_A_YL2Miv7Q0_2),.clk(gclk));
	jdff dff_A_mvYfA7ak6_0(.dout(w_n216_1[0]),.din(w_dff_A_mvYfA7ak6_0),.clk(gclk));
	jdff dff_A_sehqTj2E5_2(.dout(w_n216_0[2]),.din(w_dff_A_sehqTj2E5_2),.clk(gclk));
	jdff dff_B_yc4fuzHt1_0(.din(n213),.dout(w_dff_B_yc4fuzHt1_0),.clk(gclk));
	jdff dff_B_x0dXhVj88_0(.din(w_dff_B_yc4fuzHt1_0),.dout(w_dff_B_x0dXhVj88_0),.clk(gclk));
	jdff dff_B_9Vd1GOLh7_0(.din(w_dff_B_x0dXhVj88_0),.dout(w_dff_B_9Vd1GOLh7_0),.clk(gclk));
	jdff dff_A_t2ZLaWgT3_1(.dout(w_n192_0[1]),.din(w_dff_A_t2ZLaWgT3_1),.clk(gclk));
	jdff dff_A_6H0WDGGA8_0(.dout(w_n191_0[0]),.din(w_dff_A_6H0WDGGA8_0),.clk(gclk));
	jdff dff_A_bCtB2c645_2(.dout(w_n191_0[2]),.din(w_dff_A_bCtB2c645_2),.clk(gclk));
	jdff dff_A_QnfWgLoo0_1(.dout(w_n182_1[1]),.din(w_dff_A_QnfWgLoo0_1),.clk(gclk));
	jdff dff_A_jGjusVUl4_0(.dout(w_n182_0[0]),.din(w_dff_A_jGjusVUl4_0),.clk(gclk));
	jdff dff_A_wGfFCvUd2_0(.dout(w_dff_A_jGjusVUl4_0),.din(w_dff_A_wGfFCvUd2_0),.clk(gclk));
	jdff dff_A_WL8mdX3K8_0(.dout(w_dff_A_wGfFCvUd2_0),.din(w_dff_A_WL8mdX3K8_0),.clk(gclk));
	jdff dff_A_Gf1fOO9v0_2(.dout(w_n182_0[2]),.din(w_dff_A_Gf1fOO9v0_2),.clk(gclk));
	jdff dff_A_4Dnh2owz6_2(.dout(w_dff_A_Gf1fOO9v0_2),.din(w_dff_A_4Dnh2owz6_2),.clk(gclk));
	jdff dff_A_Axm0Vv1I7_2(.dout(w_dff_A_4Dnh2owz6_2),.din(w_dff_A_Axm0Vv1I7_2),.clk(gclk));
	jdff dff_A_YoKxsKfO2_2(.dout(w_dff_A_Axm0Vv1I7_2),.din(w_dff_A_YoKxsKfO2_2),.clk(gclk));
	jdff dff_A_y3BIuxuQ6_0(.dout(w_n180_0[0]),.din(w_dff_A_y3BIuxuQ6_0),.clk(gclk));
	jdff dff_A_o5HX76V06_1(.dout(w_G900_0[1]),.din(w_dff_A_o5HX76V06_1),.clk(gclk));
	jdff dff_A_yuQe9kTT3_1(.dout(w_n177_0[1]),.din(w_dff_A_yuQe9kTT3_1),.clk(gclk));
	jdff dff_A_r82Pybnj4_2(.dout(w_n177_0[2]),.din(w_dff_A_r82Pybnj4_2),.clk(gclk));
	jdff dff_A_Eo3OP6EE2_0(.dout(w_n175_0[0]),.din(w_dff_A_Eo3OP6EE2_0),.clk(gclk));
	jdff dff_A_H2zQJU8B6_1(.dout(w_n174_0[1]),.din(w_dff_A_H2zQJU8B6_1),.clk(gclk));
	jdff dff_B_2dksoSKa9_2(.din(n174),.dout(w_dff_B_2dksoSKa9_2),.clk(gclk));
	jdff dff_A_ljf1Bi7P1_1(.dout(w_n199_0[1]),.din(w_dff_A_ljf1Bi7P1_1),.clk(gclk));
	jdff dff_A_yPIgSjky6_1(.dout(w_dff_A_ljf1Bi7P1_1),.din(w_dff_A_yPIgSjky6_1),.clk(gclk));
	jdff dff_A_3UBavrO18_0(.dout(w_n197_1[0]),.din(w_dff_A_3UBavrO18_0),.clk(gclk));
	jdff dff_B_bAL3FZPL7_2(.din(n170),.dout(w_dff_B_bAL3FZPL7_2),.clk(gclk));
	jdff dff_A_vbbhBETj6_2(.dout(w_n154_0[2]),.din(w_dff_A_vbbhBETj6_2),.clk(gclk));
	jdff dff_A_YQvrdROC5_2(.dout(w_dff_A_vbbhBETj6_2),.din(w_dff_A_YQvrdROC5_2),.clk(gclk));
	jdff dff_A_Rn7lfHCP7_2(.dout(w_dff_A_YQvrdROC5_2),.din(w_dff_A_Rn7lfHCP7_2),.clk(gclk));
	jdff dff_A_TB3CFVc45_2(.dout(w_dff_A_Rn7lfHCP7_2),.din(w_dff_A_TB3CFVc45_2),.clk(gclk));
	jdff dff_B_raM7NCsX4_1(.din(n142),.dout(w_dff_B_raM7NCsX4_1),.clk(gclk));
	jdff dff_B_b594Y2jO9_1(.din(w_dff_B_raM7NCsX4_1),.dout(w_dff_B_b594Y2jO9_1),.clk(gclk));
	jdff dff_B_ztlquN5g3_1(.din(w_dff_B_b594Y2jO9_1),.dout(w_dff_B_ztlquN5g3_1),.clk(gclk));
	jdff dff_B_oA9mZ8LN9_1(.din(w_dff_B_ztlquN5g3_1),.dout(w_dff_B_oA9mZ8LN9_1),.clk(gclk));
	jdff dff_B_Mxv7YFLo4_1(.din(w_dff_B_oA9mZ8LN9_1),.dout(w_dff_B_Mxv7YFLo4_1),.clk(gclk));
	jdff dff_A_bs9puDA28_1(.dout(w_n93_1[1]),.din(w_dff_A_bs9puDA28_1),.clk(gclk));
	jdff dff_A_gt2VHgWJ4_1(.dout(w_dff_A_bs9puDA28_1),.din(w_dff_A_gt2VHgWJ4_1),.clk(gclk));
	jdff dff_A_LhbJ3WDd8_1(.dout(w_n93_0[1]),.din(w_dff_A_LhbJ3WDd8_1),.clk(gclk));
	jdff dff_A_OsegNpXQ2_2(.dout(w_n93_0[2]),.din(w_dff_A_OsegNpXQ2_2),.clk(gclk));
	jdff dff_A_CSeTQGlo6_0(.dout(w_n166_0[0]),.din(w_dff_A_CSeTQGlo6_0),.clk(gclk));
	jdff dff_A_dWLe2s8Q4_1(.dout(w_n165_0[1]),.din(w_dff_A_dWLe2s8Q4_1),.clk(gclk));
	jdff dff_A_XBGQncMn4_2(.dout(w_n165_0[2]),.din(w_dff_A_XBGQncMn4_2),.clk(gclk));
	jdff dff_B_dIolIVmb4_1(.din(n132),.dout(w_dff_B_dIolIVmb4_1),.clk(gclk));
	jdff dff_B_fvnInEzm1_1(.din(w_dff_B_dIolIVmb4_1),.dout(w_dff_B_fvnInEzm1_1),.clk(gclk));
	jdff dff_B_Yg7vPTC64_1(.din(w_dff_B_fvnInEzm1_1),.dout(w_dff_B_Yg7vPTC64_1),.clk(gclk));
	jdff dff_B_dvmuNwsN3_1(.din(w_dff_B_Yg7vPTC64_1),.dout(w_dff_B_dvmuNwsN3_1),.clk(gclk));
	jdff dff_B_nKMMM2cI3_1(.din(w_dff_B_dvmuNwsN3_1),.dout(w_dff_B_nKMMM2cI3_1),.clk(gclk));
	jdff dff_A_BqKbgA812_1(.dout(w_n122_0[1]),.din(w_dff_A_BqKbgA812_1),.clk(gclk));
	jdff dff_A_rQqc1nWU3_0(.dout(w_n208_0[0]),.din(w_dff_A_rQqc1nWU3_0),.clk(gclk));
	jdff dff_A_D6wwbt1I7_1(.dout(w_n197_0[1]),.din(w_dff_A_D6wwbt1I7_1),.clk(gclk));
	jdff dff_B_cYVFmp2Q2_1(.din(n194),.dout(w_dff_B_cYVFmp2Q2_1),.clk(gclk));
	jdff dff_B_AAI2YqKa1_1(.din(w_dff_B_cYVFmp2Q2_1),.dout(w_dff_B_AAI2YqKa1_1),.clk(gclk));
	jdff dff_B_nFzxAVfw5_1(.din(w_dff_B_AAI2YqKa1_1),.dout(w_dff_B_nFzxAVfw5_1),.clk(gclk));
	jdff dff_B_hNv2kRgM7_1(.din(w_dff_B_nFzxAVfw5_1),.dout(w_dff_B_hNv2kRgM7_1),.clk(gclk));
	jdff dff_B_EZajK4Zx4_1(.din(w_dff_B_hNv2kRgM7_1),.dout(w_dff_B_EZajK4Zx4_1),.clk(gclk));
	jdff dff_A_mWbAcvmq0_0(.dout(w_n118_0[0]),.din(w_dff_A_mWbAcvmq0_0),.clk(gclk));
	jdff dff_A_FeUaWPZB4_0(.dout(w_dff_A_mWbAcvmq0_0),.din(w_dff_A_FeUaWPZB4_0),.clk(gclk));
	jdff dff_A_7vFu0o4n8_0(.dout(w_dff_A_FeUaWPZB4_0),.din(w_dff_A_7vFu0o4n8_0),.clk(gclk));
	jdff dff_A_MbAnB5Qd6_0(.dout(w_dff_A_7vFu0o4n8_0),.din(w_dff_A_MbAnB5Qd6_0),.clk(gclk));
	jdff dff_A_MNOQRZPF0_0(.dout(w_dff_A_MbAnB5Qd6_0),.din(w_dff_A_MNOQRZPF0_0),.clk(gclk));
	jdff dff_A_AUxs2JCG2_0(.dout(w_dff_A_MNOQRZPF0_0),.din(w_dff_A_AUxs2JCG2_0),.clk(gclk));
	jdff dff_A_qQ9Fba7L5_0(.dout(w_dff_A_AUxs2JCG2_0),.din(w_dff_A_qQ9Fba7L5_0),.clk(gclk));
	jdff dff_A_knnKQf9j0_0(.dout(w_dff_A_qQ9Fba7L5_0),.din(w_dff_A_knnKQf9j0_0),.clk(gclk));
	jdff dff_A_AAeKoEmm2_0(.dout(w_dff_A_knnKQf9j0_0),.din(w_dff_A_AAeKoEmm2_0),.clk(gclk));
	jdff dff_A_znJYkK2h1_0(.dout(w_dff_A_AAeKoEmm2_0),.din(w_dff_A_znJYkK2h1_0),.clk(gclk));
	jdff dff_A_XtzpvVlA5_0(.dout(w_dff_A_znJYkK2h1_0),.din(w_dff_A_XtzpvVlA5_0),.clk(gclk));
	jdff dff_A_CqFgFXHW0_0(.dout(w_dff_A_XtzpvVlA5_0),.din(w_dff_A_CqFgFXHW0_0),.clk(gclk));
	jdff dff_A_wqXB6xBt2_0(.dout(w_dff_A_CqFgFXHW0_0),.din(w_dff_A_wqXB6xBt2_0),.clk(gclk));
	jdff dff_A_PSy1Ef8v9_1(.dout(w_G227_0[1]),.din(w_dff_A_PSy1Ef8v9_1),.clk(gclk));
	jdff dff_A_fTujv3rS0_0(.dout(w_G469_0[0]),.din(w_dff_A_fTujv3rS0_0),.clk(gclk));
	jdff dff_A_W26QZD3x7_0(.dout(w_dff_A_fTujv3rS0_0),.din(w_dff_A_W26QZD3x7_0),.clk(gclk));
	jdff dff_A_glZCvSbV0_0(.dout(w_dff_A_W26QZD3x7_0),.din(w_dff_A_glZCvSbV0_0),.clk(gclk));
	jdff dff_A_LfdWhR0k2_0(.dout(w_dff_A_glZCvSbV0_0),.din(w_dff_A_LfdWhR0k2_0),.clk(gclk));
	jdff dff_A_BIkT6B4Y6_0(.dout(w_dff_A_LfdWhR0k2_0),.din(w_dff_A_BIkT6B4Y6_0),.clk(gclk));
	jdff dff_A_152QaVWZ4_0(.dout(w_dff_A_BIkT6B4Y6_0),.din(w_dff_A_152QaVWZ4_0),.clk(gclk));
	jdff dff_A_TVAszvr33_0(.dout(w_dff_A_152QaVWZ4_0),.din(w_dff_A_TVAszvr33_0),.clk(gclk));
	jdff dff_A_jQwZCwyL4_0(.dout(w_dff_A_TVAszvr33_0),.din(w_dff_A_jQwZCwyL4_0),.clk(gclk));
	jdff dff_A_RmLCvJR08_0(.dout(w_dff_A_jQwZCwyL4_0),.din(w_dff_A_RmLCvJR08_0),.clk(gclk));
	jdff dff_A_FsXolQU91_0(.dout(w_dff_A_RmLCvJR08_0),.din(w_dff_A_FsXolQU91_0),.clk(gclk));
	jdff dff_A_USbeHMh75_0(.dout(w_dff_A_FsXolQU91_0),.din(w_dff_A_USbeHMh75_0),.clk(gclk));
	jdff dff_A_g0hz9BCR9_0(.dout(w_dff_A_USbeHMh75_0),.din(w_dff_A_g0hz9BCR9_0),.clk(gclk));
	jdff dff_A_jJXHTid63_0(.dout(w_dff_A_g0hz9BCR9_0),.din(w_dff_A_jJXHTid63_0),.clk(gclk));
	jdff dff_A_fts2igdj9_0(.dout(w_dff_A_jJXHTid63_0),.din(w_dff_A_fts2igdj9_0),.clk(gclk));
	jdff dff_A_9afLu5cr4_0(.dout(w_dff_A_fts2igdj9_0),.din(w_dff_A_9afLu5cr4_0),.clk(gclk));
	jdff dff_A_Ki5uAwD32_0(.dout(w_dff_A_9afLu5cr4_0),.din(w_dff_A_Ki5uAwD32_0),.clk(gclk));
	jdff dff_A_qTumxMiU7_2(.dout(w_G469_0[2]),.din(w_dff_A_qTumxMiU7_2),.clk(gclk));
	jdff dff_A_VjfWHbZr1_2(.dout(w_dff_A_qTumxMiU7_2),.din(w_dff_A_VjfWHbZr1_2),.clk(gclk));
	jdff dff_A_4ygaUCMi0_2(.dout(w_dff_A_VjfWHbZr1_2),.din(w_dff_A_4ygaUCMi0_2),.clk(gclk));
	jdff dff_A_OeVzAPap7_2(.dout(w_dff_A_4ygaUCMi0_2),.din(w_dff_A_OeVzAPap7_2),.clk(gclk));
	jdff dff_A_aEk61aJ43_2(.dout(w_dff_A_OeVzAPap7_2),.din(w_dff_A_aEk61aJ43_2),.clk(gclk));
	jdff dff_A_Ainhjsqa1_2(.dout(w_dff_A_aEk61aJ43_2),.din(w_dff_A_Ainhjsqa1_2),.clk(gclk));
	jdff dff_A_Fao2cAqc6_1(.dout(w_n113_0[1]),.din(w_dff_A_Fao2cAqc6_1),.clk(gclk));
	jdff dff_A_pQOq6Uh58_1(.dout(w_dff_A_Fao2cAqc6_1),.din(w_dff_A_pQOq6Uh58_1),.clk(gclk));
	jdff dff_A_37wy3utU9_2(.dout(w_n113_0[2]),.din(w_dff_A_37wy3utU9_2),.clk(gclk));
	jdff dff_A_glx4b2HU7_2(.dout(w_dff_A_37wy3utU9_2),.din(w_dff_A_glx4b2HU7_2),.clk(gclk));
	jdff dff_A_MyexSgyj5_1(.dout(w_n112_0[1]),.din(w_dff_A_MyexSgyj5_1),.clk(gclk));
	jdff dff_A_jsgNo3aG6_1(.dout(w_dff_A_MyexSgyj5_1),.din(w_dff_A_jsgNo3aG6_1),.clk(gclk));
	jdff dff_A_szorhQwO6_1(.dout(w_dff_A_jsgNo3aG6_1),.din(w_dff_A_szorhQwO6_1),.clk(gclk));
	jdff dff_A_Z9JB7D5B1_2(.dout(w_n112_0[2]),.din(w_dff_A_Z9JB7D5B1_2),.clk(gclk));
	jdff dff_A_BMhIXWMj5_2(.dout(w_dff_A_Z9JB7D5B1_2),.din(w_dff_A_BMhIXWMj5_2),.clk(gclk));
	jdff dff_A_4ZH5GRqy3_2(.dout(w_dff_A_BMhIXWMj5_2),.din(w_dff_A_4ZH5GRqy3_2),.clk(gclk));
	jdff dff_A_wxCamwqG0_1(.dout(w_n109_0[1]),.din(w_dff_A_wxCamwqG0_1),.clk(gclk));
	jdff dff_A_vs0lCKW85_1(.dout(w_dff_A_wxCamwqG0_1),.din(w_dff_A_vs0lCKW85_1),.clk(gclk));
	jdff dff_A_PKSGSRMF5_1(.dout(w_dff_A_vs0lCKW85_1),.din(w_dff_A_PKSGSRMF5_1),.clk(gclk));
	jdff dff_A_XXodlFnk5_1(.dout(w_dff_A_PKSGSRMF5_1),.din(w_dff_A_XXodlFnk5_1),.clk(gclk));
	jdff dff_A_Jq81yBNG1_0(.dout(w_n107_0[0]),.din(w_dff_A_Jq81yBNG1_0),.clk(gclk));
	jdff dff_A_mbCLDJc58_0(.dout(w_dff_A_Jq81yBNG1_0),.din(w_dff_A_mbCLDJc58_0),.clk(gclk));
	jdff dff_A_eVJwQ8Rd6_0(.dout(w_dff_A_mbCLDJc58_0),.din(w_dff_A_eVJwQ8Rd6_0),.clk(gclk));
	jdff dff_A_dlUm5GdS9_0(.dout(w_dff_A_eVJwQ8Rd6_0),.din(w_dff_A_dlUm5GdS9_0),.clk(gclk));
	jdff dff_A_5l6aGnp06_0(.dout(w_dff_A_dlUm5GdS9_0),.din(w_dff_A_5l6aGnp06_0),.clk(gclk));
	jdff dff_A_6Znmh7On2_0(.dout(w_dff_A_5l6aGnp06_0),.din(w_dff_A_6Znmh7On2_0),.clk(gclk));
	jdff dff_A_KBIeAkO20_0(.dout(w_dff_A_6Znmh7On2_0),.din(w_dff_A_KBIeAkO20_0),.clk(gclk));
	jdff dff_A_7bhc17KK1_0(.dout(w_dff_A_KBIeAkO20_0),.din(w_dff_A_7bhc17KK1_0),.clk(gclk));
	jdff dff_A_ovrl5xYy2_0(.dout(w_dff_A_7bhc17KK1_0),.din(w_dff_A_ovrl5xYy2_0),.clk(gclk));
	jdff dff_A_MUlJkXFG9_0(.dout(w_dff_A_ovrl5xYy2_0),.din(w_dff_A_MUlJkXFG9_0),.clk(gclk));
	jdff dff_A_koMlqWKZ0_0(.dout(w_dff_A_MUlJkXFG9_0),.din(w_dff_A_koMlqWKZ0_0),.clk(gclk));
	jdff dff_A_ohN5pEQc0_0(.dout(w_dff_A_koMlqWKZ0_0),.din(w_dff_A_ohN5pEQc0_0),.clk(gclk));
	jdff dff_A_8DSmAR8e6_0(.dout(w_dff_A_ohN5pEQc0_0),.din(w_dff_A_8DSmAR8e6_0),.clk(gclk));
	jdff dff_B_OOoXnuC15_1(.din(n104),.dout(w_dff_B_OOoXnuC15_1),.clk(gclk));
	jdff dff_A_wdwqTUD03_1(.dout(w_G224_0[1]),.din(w_dff_A_wdwqTUD03_1),.clk(gclk));
	jdff dff_B_yLgtjOzk6_0(.din(n101),.dout(w_dff_B_yLgtjOzk6_0),.clk(gclk));
	jdff dff_B_tglVqJNZ7_0(.din(w_dff_B_yLgtjOzk6_0),.dout(w_dff_B_tglVqJNZ7_0),.clk(gclk));
	jdff dff_A_dYQ2sOnO3_0(.dout(w_n99_0[0]),.din(w_dff_A_dYQ2sOnO3_0),.clk(gclk));
	jdff dff_A_Jjn2Iy6I8_1(.dout(w_n96_0[1]),.din(w_dff_A_Jjn2Iy6I8_1),.clk(gclk));
	jdff dff_A_kiIlB8Vh1_1(.dout(w_dff_A_Jjn2Iy6I8_1),.din(w_dff_A_kiIlB8Vh1_1),.clk(gclk));
	jdff dff_A_PFqwSlRL6_2(.dout(w_n96_0[2]),.din(w_dff_A_PFqwSlRL6_2),.clk(gclk));
	jdff dff_A_H8F0IXdL4_2(.dout(w_dff_A_PFqwSlRL6_2),.din(w_dff_A_H8F0IXdL4_2),.clk(gclk));
	jdff dff_B_O4s8zUHl7_3(.din(n96),.dout(w_dff_B_O4s8zUHl7_3),.clk(gclk));
	jdff dff_B_JCHEIWWr5_3(.din(w_dff_B_O4s8zUHl7_3),.dout(w_dff_B_JCHEIWWr5_3),.clk(gclk));
	jdff dff_A_5YQM2Dv99_0(.dout(w_n95_1[0]),.din(w_dff_A_5YQM2Dv99_0),.clk(gclk));
	jdff dff_A_ufFIFDr17_0(.dout(w_dff_A_5YQM2Dv99_0),.din(w_dff_A_ufFIFDr17_0),.clk(gclk));
	jdff dff_A_in8rgn4A9_1(.dout(w_n95_0[1]),.din(w_dff_A_in8rgn4A9_1),.clk(gclk));
	jdff dff_A_kvKSfVHq6_1(.dout(w_dff_A_in8rgn4A9_1),.din(w_dff_A_kvKSfVHq6_1),.clk(gclk));
	jdff dff_A_lp5uNfOn0_1(.dout(w_dff_A_kvKSfVHq6_1),.din(w_dff_A_lp5uNfOn0_1),.clk(gclk));
	jdff dff_A_ChyF10g46_1(.dout(w_dff_A_lp5uNfOn0_1),.din(w_dff_A_ChyF10g46_1),.clk(gclk));
	jdff dff_A_TAIfjDqB5_1(.dout(w_dff_A_ChyF10g46_1),.din(w_dff_A_TAIfjDqB5_1),.clk(gclk));
	jdff dff_A_hTI2R2GC7_2(.dout(w_n95_0[2]),.din(w_dff_A_hTI2R2GC7_2),.clk(gclk));
	jdff dff_A_O8CXT4Og7_2(.dout(w_dff_A_hTI2R2GC7_2),.din(w_dff_A_O8CXT4Og7_2),.clk(gclk));
	jdff dff_A_ECJUwDdp2_2(.dout(w_dff_A_O8CXT4Og7_2),.din(w_dff_A_ECJUwDdp2_2),.clk(gclk));
	jdff dff_A_9pp1EhMF8_2(.dout(w_dff_A_ECJUwDdp2_2),.din(w_dff_A_9pp1EhMF8_2),.clk(gclk));
	jdff dff_A_0SNZBjMI2_2(.dout(w_dff_A_9pp1EhMF8_2),.din(w_dff_A_0SNZBjMI2_2),.clk(gclk));
	jdff dff_A_4mbwf4eE1_1(.dout(w_n161_0[1]),.din(w_dff_A_4mbwf4eE1_1),.clk(gclk));
	jdff dff_A_Yc2wWo9e0_2(.dout(w_n161_0[2]),.din(w_dff_A_Yc2wWo9e0_2),.clk(gclk));
	jdff dff_B_LUzLjp6Q9_3(.din(n161),.dout(w_dff_B_LUzLjp6Q9_3),.clk(gclk));
	jdff dff_B_IbDQEo7i1_1(.din(n159),.dout(w_dff_B_IbDQEo7i1_1),.clk(gclk));
	jdff dff_B_hFX4NJtE3_1(.din(w_dff_B_IbDQEo7i1_1),.dout(w_dff_B_hFX4NJtE3_1),.clk(gclk));
	jdff dff_B_YeSQtdKL2_1(.din(w_dff_B_hFX4NJtE3_1),.dout(w_dff_B_YeSQtdKL2_1),.clk(gclk));
	jdff dff_B_373lpKxb8_1(.din(w_dff_B_YeSQtdKL2_1),.dout(w_dff_B_373lpKxb8_1),.clk(gclk));
	jdff dff_B_oEXkI1vY7_1(.din(w_dff_B_373lpKxb8_1),.dout(w_dff_B_oEXkI1vY7_1),.clk(gclk));
	jdff dff_A_IVJjGBzk6_0(.dout(w_n90_0[0]),.din(w_dff_A_IVJjGBzk6_0),.clk(gclk));
	jdff dff_A_XpbkbB1C2_0(.dout(w_dff_A_IVJjGBzk6_0),.din(w_dff_A_XpbkbB1C2_0),.clk(gclk));
	jdff dff_A_fSRLNKkA8_0(.dout(w_dff_A_XpbkbB1C2_0),.din(w_dff_A_fSRLNKkA8_0),.clk(gclk));
	jdff dff_A_HvLa1AXe2_0(.dout(w_dff_A_fSRLNKkA8_0),.din(w_dff_A_HvLa1AXe2_0),.clk(gclk));
	jdff dff_A_uyyNAPEa2_0(.dout(w_dff_A_HvLa1AXe2_0),.din(w_dff_A_uyyNAPEa2_0),.clk(gclk));
	jdff dff_A_3jmxAeI24_0(.dout(w_dff_A_uyyNAPEa2_0),.din(w_dff_A_3jmxAeI24_0),.clk(gclk));
	jdff dff_A_P1ifWpEv2_0(.dout(w_dff_A_3jmxAeI24_0),.din(w_dff_A_P1ifWpEv2_0),.clk(gclk));
	jdff dff_A_Hrd8bJTN3_0(.dout(w_dff_A_P1ifWpEv2_0),.din(w_dff_A_Hrd8bJTN3_0),.clk(gclk));
	jdff dff_A_eS4RkAuC2_0(.dout(w_dff_A_Hrd8bJTN3_0),.din(w_dff_A_eS4RkAuC2_0),.clk(gclk));
	jdff dff_A_cVEwS4jw2_0(.dout(w_dff_A_eS4RkAuC2_0),.din(w_dff_A_cVEwS4jw2_0),.clk(gclk));
	jdff dff_A_bwh7ArJO1_0(.dout(w_dff_A_cVEwS4jw2_0),.din(w_dff_A_bwh7ArJO1_0),.clk(gclk));
	jdff dff_A_lDGQmxr08_0(.dout(w_dff_A_bwh7ArJO1_0),.din(w_dff_A_lDGQmxr08_0),.clk(gclk));
	jdff dff_A_WaaanRHD1_0(.dout(w_G210_0[0]),.din(w_dff_A_WaaanRHD1_0),.clk(gclk));
	jdff dff_A_X4uqIgWo4_0(.dout(w_dff_A_WaaanRHD1_0),.din(w_dff_A_X4uqIgWo4_0),.clk(gclk));
	jdff dff_A_MU7cEkiq8_0(.dout(w_dff_A_X4uqIgWo4_0),.din(w_dff_A_MU7cEkiq8_0),.clk(gclk));
	jdff dff_A_RMZzRwnv4_0(.dout(w_dff_A_MU7cEkiq8_0),.din(w_dff_A_RMZzRwnv4_0),.clk(gclk));
	jdff dff_A_mXfaxYyM3_0(.dout(w_dff_A_RMZzRwnv4_0),.din(w_dff_A_mXfaxYyM3_0),.clk(gclk));
	jdff dff_A_VD3Cy5BD7_0(.dout(w_dff_A_mXfaxYyM3_0),.din(w_dff_A_VD3Cy5BD7_0),.clk(gclk));
	jdff dff_A_AkfgV1Eh4_0(.dout(w_dff_A_VD3Cy5BD7_0),.din(w_dff_A_AkfgV1Eh4_0),.clk(gclk));
	jdff dff_A_Tjz2ZwEm3_0(.dout(w_dff_A_AkfgV1Eh4_0),.din(w_dff_A_Tjz2ZwEm3_0),.clk(gclk));
	jdff dff_A_YCF3mrwO9_0(.dout(w_dff_A_Tjz2ZwEm3_0),.din(w_dff_A_YCF3mrwO9_0),.clk(gclk));
	jdff dff_A_HWNHflyG8_0(.dout(w_dff_A_YCF3mrwO9_0),.din(w_dff_A_HWNHflyG8_0),.clk(gclk));
	jdff dff_A_bDfma8U30_0(.dout(w_dff_A_HWNHflyG8_0),.din(w_dff_A_bDfma8U30_0),.clk(gclk));
	jdff dff_A_Iu1zOiwH6_0(.dout(w_dff_A_bDfma8U30_0),.din(w_dff_A_Iu1zOiwH6_0),.clk(gclk));
	jdff dff_A_TAGELWTD5_0(.dout(w_dff_A_Iu1zOiwH6_0),.din(w_dff_A_TAGELWTD5_0),.clk(gclk));
	jdff dff_A_TfkoPOzq8_0(.dout(w_dff_A_TAGELWTD5_0),.din(w_dff_A_TfkoPOzq8_0),.clk(gclk));
	jdff dff_A_TTg2vcIa2_0(.dout(w_dff_A_TfkoPOzq8_0),.din(w_dff_A_TTg2vcIa2_0),.clk(gclk));
	jdff dff_A_Dvrpoyht9_0(.dout(w_dff_A_TTg2vcIa2_0),.din(w_dff_A_Dvrpoyht9_0),.clk(gclk));
	jdff dff_A_Fnzdoirm6_1(.dout(w_G210_0[1]),.din(w_dff_A_Fnzdoirm6_1),.clk(gclk));
	jdff dff_A_63Xj2V504_0(.dout(w_G101_0[0]),.din(w_dff_A_63Xj2V504_0),.clk(gclk));
	jdff dff_A_7ptXhgKe3_0(.dout(w_dff_A_63Xj2V504_0),.din(w_dff_A_7ptXhgKe3_0),.clk(gclk));
	jdff dff_A_okrlDpS29_0(.dout(w_dff_A_7ptXhgKe3_0),.din(w_dff_A_okrlDpS29_0),.clk(gclk));
	jdff dff_A_I8vmvHrG2_0(.dout(w_dff_A_okrlDpS29_0),.din(w_dff_A_I8vmvHrG2_0),.clk(gclk));
	jdff dff_A_7M5jHN025_0(.dout(w_dff_A_I8vmvHrG2_0),.din(w_dff_A_7M5jHN025_0),.clk(gclk));
	jdff dff_A_7gCRq0WD5_0(.dout(w_dff_A_7M5jHN025_0),.din(w_dff_A_7gCRq0WD5_0),.clk(gclk));
	jdff dff_A_Oo6WF2vO3_0(.dout(w_dff_A_7gCRq0WD5_0),.din(w_dff_A_Oo6WF2vO3_0),.clk(gclk));
	jdff dff_A_vXHwLd4q7_0(.dout(w_dff_A_Oo6WF2vO3_0),.din(w_dff_A_vXHwLd4q7_0),.clk(gclk));
	jdff dff_A_HmwdAIXL9_0(.dout(w_dff_A_vXHwLd4q7_0),.din(w_dff_A_HmwdAIXL9_0),.clk(gclk));
	jdff dff_A_2Se3tiNk8_0(.dout(w_dff_A_HmwdAIXL9_0),.din(w_dff_A_2Se3tiNk8_0),.clk(gclk));
	jdff dff_A_R8YlHE2w3_0(.dout(w_dff_A_2Se3tiNk8_0),.din(w_dff_A_R8YlHE2w3_0),.clk(gclk));
	jdff dff_A_6g28ZD0h5_2(.dout(w_G101_0[2]),.din(w_dff_A_6g28ZD0h5_2),.clk(gclk));
	jdff dff_A_VXWWuc3X5_2(.dout(w_dff_A_6g28ZD0h5_2),.din(w_dff_A_VXWWuc3X5_2),.clk(gclk));
	jdff dff_A_DTpVIFKE5_1(.dout(w_n84_0[1]),.din(w_dff_A_DTpVIFKE5_1),.clk(gclk));
	jdff dff_A_0W73h6m64_1(.dout(w_n81_0[1]),.din(w_dff_A_0W73h6m64_1),.clk(gclk));
	jdff dff_A_1jcsAr9G2_2(.dout(w_n81_0[2]),.din(w_dff_A_1jcsAr9G2_2),.clk(gclk));
	jdff dff_A_hVdLlbEz0_2(.dout(w_G472_0[2]),.din(w_dff_A_hVdLlbEz0_2),.clk(gclk));
	jdff dff_A_hL5gAhwG1_2(.dout(w_dff_A_hVdLlbEz0_2),.din(w_dff_A_hL5gAhwG1_2),.clk(gclk));
	jdff dff_A_XAJyGXLt1_2(.dout(w_dff_A_hL5gAhwG1_2),.din(w_dff_A_XAJyGXLt1_2),.clk(gclk));
	jdff dff_A_4odj30ia1_2(.dout(w_dff_A_XAJyGXLt1_2),.din(w_dff_A_4odj30ia1_2),.clk(gclk));
	jdff dff_A_zpzRYhAj1_2(.dout(w_dff_A_4odj30ia1_2),.din(w_dff_A_zpzRYhAj1_2),.clk(gclk));
	jdff dff_A_ngie6Vjf5_2(.dout(w_dff_A_zpzRYhAj1_2),.din(w_dff_A_ngie6Vjf5_2),.clk(gclk));
	jdff dff_B_gdUnpY1m1_0(.din(n75),.dout(w_dff_B_gdUnpY1m1_0),.clk(gclk));
	jdff dff_A_RwYGsJCT6_0(.dout(w_n74_0[0]),.din(w_dff_A_RwYGsJCT6_0),.clk(gclk));
	jdff dff_A_O1ecZPEC7_0(.dout(w_dff_A_RwYGsJCT6_0),.din(w_dff_A_O1ecZPEC7_0),.clk(gclk));
	jdff dff_A_hgOT9GkU1_0(.dout(w_n70_0[0]),.din(w_dff_A_hgOT9GkU1_0),.clk(gclk));
	jdff dff_A_GXhKf2iZ7_0(.dout(w_dff_A_hgOT9GkU1_0),.din(w_dff_A_GXhKf2iZ7_0),.clk(gclk));
	jdff dff_A_gZQjpllN0_0(.dout(w_dff_A_GXhKf2iZ7_0),.din(w_dff_A_gZQjpllN0_0),.clk(gclk));
	jdff dff_A_TT9wvXy35_0(.dout(w_dff_A_gZQjpllN0_0),.din(w_dff_A_TT9wvXy35_0),.clk(gclk));
	jdff dff_A_yrBFt94H4_0(.dout(w_dff_A_TT9wvXy35_0),.din(w_dff_A_yrBFt94H4_0),.clk(gclk));
	jdff dff_A_lQpPB3ZW5_0(.dout(w_dff_A_yrBFt94H4_0),.din(w_dff_A_lQpPB3ZW5_0),.clk(gclk));
	jdff dff_A_qCeLwvIR4_0(.dout(w_dff_A_lQpPB3ZW5_0),.din(w_dff_A_qCeLwvIR4_0),.clk(gclk));
	jdff dff_A_0rwgrJoI1_0(.dout(w_dff_A_qCeLwvIR4_0),.din(w_dff_A_0rwgrJoI1_0),.clk(gclk));
	jdff dff_A_AXRqwrCx0_0(.dout(w_dff_A_0rwgrJoI1_0),.din(w_dff_A_AXRqwrCx0_0),.clk(gclk));
	jdff dff_A_RSaRzvei8_0(.dout(w_dff_A_AXRqwrCx0_0),.din(w_dff_A_RSaRzvei8_0),.clk(gclk));
	jdff dff_A_QZSIMUtJ3_0(.dout(w_dff_A_RSaRzvei8_0),.din(w_dff_A_QZSIMUtJ3_0),.clk(gclk));
	jdff dff_A_xs6BUOcj4_0(.dout(w_dff_A_QZSIMUtJ3_0),.din(w_dff_A_xs6BUOcj4_0),.clk(gclk));
	jdff dff_A_RtDpuMvy0_0(.dout(w_dff_A_xs6BUOcj4_0),.din(w_dff_A_RtDpuMvy0_0),.clk(gclk));
	jdff dff_B_fOfk53P32_0(.din(n69),.dout(w_dff_B_fOfk53P32_0),.clk(gclk));
	jdff dff_B_SezSqpel8_0(.din(n68),.dout(w_dff_B_SezSqpel8_0),.clk(gclk));
	jdff dff_A_pKZNHe552_0(.dout(w_G137_0[0]),.din(w_dff_A_pKZNHe552_0),.clk(gclk));
	jdff dff_A_3oi60fMZ4_0(.dout(w_dff_A_pKZNHe552_0),.din(w_dff_A_3oi60fMZ4_0),.clk(gclk));
	jdff dff_A_mhuuLXXT6_0(.dout(w_dff_A_3oi60fMZ4_0),.din(w_dff_A_mhuuLXXT6_0),.clk(gclk));
	jdff dff_A_d1KPOBMq1_0(.dout(w_dff_A_mhuuLXXT6_0),.din(w_dff_A_d1KPOBMq1_0),.clk(gclk));
	jdff dff_A_mHAJuHcK2_0(.dout(w_dff_A_d1KPOBMq1_0),.din(w_dff_A_mHAJuHcK2_0),.clk(gclk));
	jdff dff_A_Hpte4vfu5_0(.dout(w_dff_A_mHAJuHcK2_0),.din(w_dff_A_Hpte4vfu5_0),.clk(gclk));
	jdff dff_A_TK4fxhqT6_0(.dout(w_dff_A_Hpte4vfu5_0),.din(w_dff_A_TK4fxhqT6_0),.clk(gclk));
	jdff dff_A_S0XfC0pO6_0(.dout(w_dff_A_TK4fxhqT6_0),.din(w_dff_A_S0XfC0pO6_0),.clk(gclk));
	jdff dff_A_g5sZoqxD7_0(.dout(w_dff_A_S0XfC0pO6_0),.din(w_dff_A_g5sZoqxD7_0),.clk(gclk));
	jdff dff_A_kk5aMkAw7_0(.dout(w_dff_A_g5sZoqxD7_0),.din(w_dff_A_kk5aMkAw7_0),.clk(gclk));
	jdff dff_A_QKqVNlEN5_0(.dout(w_dff_A_kk5aMkAw7_0),.din(w_dff_A_QKqVNlEN5_0),.clk(gclk));
	jdff dff_B_E2gMzbzZ7_0(.din(n64),.dout(w_dff_B_E2gMzbzZ7_0),.clk(gclk));
	jdff dff_A_tNTC83n08_0(.dout(w_G119_0[0]),.din(w_dff_A_tNTC83n08_0),.clk(gclk));
	jdff dff_A_ksZUfEAq9_0(.dout(w_dff_A_tNTC83n08_0),.din(w_dff_A_ksZUfEAq9_0),.clk(gclk));
	jdff dff_A_sJWnaMA38_0(.dout(w_dff_A_ksZUfEAq9_0),.din(w_dff_A_sJWnaMA38_0),.clk(gclk));
	jdff dff_A_j4SrJ4Ch5_0(.dout(w_dff_A_sJWnaMA38_0),.din(w_dff_A_j4SrJ4Ch5_0),.clk(gclk));
	jdff dff_A_btybmDyg1_0(.dout(w_dff_A_j4SrJ4Ch5_0),.din(w_dff_A_btybmDyg1_0),.clk(gclk));
	jdff dff_A_pDflvThv8_0(.dout(w_dff_A_btybmDyg1_0),.din(w_dff_A_pDflvThv8_0),.clk(gclk));
	jdff dff_A_sBiep1zc3_0(.dout(w_dff_A_pDflvThv8_0),.din(w_dff_A_sBiep1zc3_0),.clk(gclk));
	jdff dff_A_OsVdRZSh4_0(.dout(w_dff_A_sBiep1zc3_0),.din(w_dff_A_OsVdRZSh4_0),.clk(gclk));
	jdff dff_A_IfvaPOnB3_0(.dout(w_dff_A_OsVdRZSh4_0),.din(w_dff_A_IfvaPOnB3_0),.clk(gclk));
	jdff dff_A_uAxIQxjG2_0(.dout(w_dff_A_IfvaPOnB3_0),.din(w_dff_A_uAxIQxjG2_0),.clk(gclk));
	jdff dff_A_I5DHfcvg5_0(.dout(w_dff_A_uAxIQxjG2_0),.din(w_dff_A_I5DHfcvg5_0),.clk(gclk));
	jdff dff_A_0lugVVhC9_2(.dout(w_G119_0[2]),.din(w_dff_A_0lugVVhC9_2),.clk(gclk));
	jdff dff_A_5Asyo8uZ5_0(.dout(w_G110_0[0]),.din(w_dff_A_5Asyo8uZ5_0),.clk(gclk));
	jdff dff_A_9eEG8FuC2_0(.dout(w_dff_A_5Asyo8uZ5_0),.din(w_dff_A_9eEG8FuC2_0),.clk(gclk));
	jdff dff_A_OwOH84eF1_0(.dout(w_dff_A_9eEG8FuC2_0),.din(w_dff_A_OwOH84eF1_0),.clk(gclk));
	jdff dff_A_xNDl61YB7_0(.dout(w_dff_A_OwOH84eF1_0),.din(w_dff_A_xNDl61YB7_0),.clk(gclk));
	jdff dff_A_8acG0xR55_0(.dout(w_dff_A_xNDl61YB7_0),.din(w_dff_A_8acG0xR55_0),.clk(gclk));
	jdff dff_A_rRjvU9CP0_0(.dout(w_dff_A_8acG0xR55_0),.din(w_dff_A_rRjvU9CP0_0),.clk(gclk));
	jdff dff_A_FV2sbfqf7_0(.dout(w_dff_A_rRjvU9CP0_0),.din(w_dff_A_FV2sbfqf7_0),.clk(gclk));
	jdff dff_A_WaBbkL3Z2_0(.dout(w_dff_A_FV2sbfqf7_0),.din(w_dff_A_WaBbkL3Z2_0),.clk(gclk));
	jdff dff_A_QQGZNuYD6_0(.dout(w_dff_A_WaBbkL3Z2_0),.din(w_dff_A_QQGZNuYD6_0),.clk(gclk));
	jdff dff_A_JXdWwEvB1_0(.dout(w_dff_A_QQGZNuYD6_0),.din(w_dff_A_JXdWwEvB1_0),.clk(gclk));
	jdff dff_A_sEbjAvFW8_0(.dout(w_dff_A_JXdWwEvB1_0),.din(w_dff_A_sEbjAvFW8_0),.clk(gclk));
	jdff dff_B_MYlh2hkP6_1(.din(n59),.dout(w_dff_B_MYlh2hkP6_1),.clk(gclk));
	jdff dff_A_FpyAogCZ2_0(.dout(w_G234_1[0]),.din(w_dff_A_FpyAogCZ2_0),.clk(gclk));
	jdff dff_A_WuZeBu4y0_0(.dout(w_G221_0[0]),.din(w_dff_A_WuZeBu4y0_0),.clk(gclk));
	jdff dff_A_WxG6asbp1_0(.dout(w_dff_A_WuZeBu4y0_0),.din(w_dff_A_WxG6asbp1_0),.clk(gclk));
	jdff dff_A_bfGVxm1p0_0(.dout(w_dff_A_WxG6asbp1_0),.din(w_dff_A_bfGVxm1p0_0),.clk(gclk));
	jdff dff_A_1X4jttEt0_0(.dout(w_n58_2[0]),.din(w_dff_A_1X4jttEt0_0),.clk(gclk));
	jdff dff_A_ks7Lw3Sr8_0(.dout(w_dff_A_1X4jttEt0_0),.din(w_dff_A_ks7Lw3Sr8_0),.clk(gclk));
	jdff dff_A_PUx7N4Rs1_0(.dout(w_dff_A_ks7Lw3Sr8_0),.din(w_dff_A_PUx7N4Rs1_0),.clk(gclk));
	jdff dff_A_rQECRfdN9_0(.dout(w_dff_A_PUx7N4Rs1_0),.din(w_dff_A_rQECRfdN9_0),.clk(gclk));
	jdff dff_A_JJUYwFe61_2(.dout(w_n58_2[2]),.din(w_dff_A_JJUYwFe61_2),.clk(gclk));
	jdff dff_A_o3ZTjruz8_2(.dout(w_dff_A_JJUYwFe61_2),.din(w_dff_A_o3ZTjruz8_2),.clk(gclk));
	jdff dff_A_RPe0UhA67_2(.dout(w_dff_A_o3ZTjruz8_2),.din(w_dff_A_RPe0UhA67_2),.clk(gclk));
	jdff dff_A_1kggSPbO3_2(.dout(w_dff_A_RPe0UhA67_2),.din(w_dff_A_1kggSPbO3_2),.clk(gclk));
	jdff dff_A_Z90Zwh8F3_0(.dout(w_n131_0[0]),.din(w_dff_A_Z90Zwh8F3_0),.clk(gclk));
	jdff dff_A_n8nmovg17_0(.dout(w_dff_A_Z90Zwh8F3_0),.din(w_dff_A_n8nmovg17_0),.clk(gclk));
	jdff dff_A_I8pmQhjl7_0(.dout(w_dff_A_n8nmovg17_0),.din(w_dff_A_I8pmQhjl7_0),.clk(gclk));
	jdff dff_A_2GMuLE8Z3_2(.dout(w_n131_0[2]),.din(w_dff_A_2GMuLE8Z3_2),.clk(gclk));
	jdff dff_A_lJ5AhLZ90_2(.dout(w_dff_A_2GMuLE8Z3_2),.din(w_dff_A_lJ5AhLZ90_2),.clk(gclk));
	jdff dff_A_J4tJ1UPO0_2(.dout(w_dff_A_lJ5AhLZ90_2),.din(w_dff_A_J4tJ1UPO0_2),.clk(gclk));
	jdff dff_A_hgCRujL88_2(.dout(w_dff_A_J4tJ1UPO0_2),.din(w_dff_A_hgCRujL88_2),.clk(gclk));
	jdff dff_A_BGe6APbO8_2(.dout(w_dff_A_hgCRujL88_2),.din(w_dff_A_BGe6APbO8_2),.clk(gclk));
	jdff dff_A_Uv9nZhjH3_1(.dout(w_n130_0[1]),.din(w_dff_A_Uv9nZhjH3_1),.clk(gclk));
	jdff dff_A_qnLsnTcA7_1(.dout(w_dff_A_Uv9nZhjH3_1),.din(w_dff_A_qnLsnTcA7_1),.clk(gclk));
	jdff dff_A_EGiaBh7U6_1(.dout(w_dff_A_qnLsnTcA7_1),.din(w_dff_A_EGiaBh7U6_1),.clk(gclk));
	jdff dff_A_yMoIAGfu6_1(.dout(w_dff_A_EGiaBh7U6_1),.din(w_dff_A_yMoIAGfu6_1),.clk(gclk));
	jdff dff_A_7XIVxcxE2_2(.dout(w_n130_0[2]),.din(w_dff_A_7XIVxcxE2_2),.clk(gclk));
	jdff dff_A_8o5KYpZZ0_2(.dout(w_dff_A_7XIVxcxE2_2),.din(w_dff_A_8o5KYpZZ0_2),.clk(gclk));
	jdff dff_A_GR1uVg2b9_2(.dout(w_dff_A_8o5KYpZZ0_2),.din(w_dff_A_GR1uVg2b9_2),.clk(gclk));
	jdff dff_A_Bxamrgzn8_2(.dout(w_dff_A_GR1uVg2b9_2),.din(w_dff_A_Bxamrgzn8_2),.clk(gclk));
	jdff dff_A_VWtukREt6_2(.dout(w_dff_A_Bxamrgzn8_2),.din(w_dff_A_VWtukREt6_2),.clk(gclk));
	jdff dff_A_wE6cvfsv4_2(.dout(w_dff_A_VWtukREt6_2),.din(w_dff_A_wE6cvfsv4_2),.clk(gclk));
	jdff dff_A_35AQNABq7_2(.dout(w_dff_A_wE6cvfsv4_2),.din(w_dff_A_35AQNABq7_2),.clk(gclk));
	jdff dff_A_iwleWXhp5_2(.dout(w_dff_A_35AQNABq7_2),.din(w_dff_A_iwleWXhp5_2),.clk(gclk));
	jdff dff_A_EfsTyA2Z4_2(.dout(w_dff_A_iwleWXhp5_2),.din(w_dff_A_EfsTyA2Z4_2),.clk(gclk));
	jdff dff_A_O9bDVYXm7_0(.dout(w_n124_0[0]),.din(w_dff_A_O9bDVYXm7_0),.clk(gclk));
	jdff dff_A_WgfzuJgN5_1(.dout(w_G898_0[1]),.din(w_dff_A_WgfzuJgN5_1),.clk(gclk));
	jdff dff_A_3b2YPRZZ3_0(.dout(w_n186_0[0]),.din(w_dff_A_3b2YPRZZ3_0),.clk(gclk));
	jdff dff_A_cfc6Fpsw1_0(.dout(w_dff_A_3b2YPRZZ3_0),.din(w_dff_A_cfc6Fpsw1_0),.clk(gclk));
	jdff dff_A_0S7blAa62_0(.dout(w_dff_A_cfc6Fpsw1_0),.din(w_dff_A_0S7blAa62_0),.clk(gclk));
	jdff dff_A_KZ7hGh7y2_1(.dout(w_n151_0[1]),.din(w_dff_A_KZ7hGh7y2_1),.clk(gclk));
	jdff dff_A_fwasoT2e1_1(.dout(w_dff_A_KZ7hGh7y2_1),.din(w_dff_A_fwasoT2e1_1),.clk(gclk));
	jdff dff_A_RuHp7h8W7_1(.dout(w_dff_A_fwasoT2e1_1),.din(w_dff_A_RuHp7h8W7_1),.clk(gclk));
	jdff dff_A_xt1G26Iq5_1(.dout(w_dff_A_RuHp7h8W7_1),.din(w_dff_A_xt1G26Iq5_1),.clk(gclk));
	jdff dff_A_ot761LEK5_1(.dout(w_dff_A_xt1G26Iq5_1),.din(w_dff_A_ot761LEK5_1),.clk(gclk));
	jdff dff_A_jucyTyvX1_1(.dout(w_dff_A_ot761LEK5_1),.din(w_dff_A_jucyTyvX1_1),.clk(gclk));
	jdff dff_A_o6nx9h7l6_1(.dout(w_dff_A_jucyTyvX1_1),.din(w_dff_A_o6nx9h7l6_1),.clk(gclk));
	jdff dff_A_0FXadMBX7_1(.dout(w_dff_A_o6nx9h7l6_1),.din(w_dff_A_0FXadMBX7_1),.clk(gclk));
	jdff dff_A_SM2TfiJu9_1(.dout(w_dff_A_0FXadMBX7_1),.din(w_dff_A_SM2TfiJu9_1),.clk(gclk));
	jdff dff_A_fmEMOViY1_1(.dout(w_dff_A_SM2TfiJu9_1),.din(w_dff_A_fmEMOViY1_1),.clk(gclk));
	jdff dff_A_eDYUT59i0_1(.dout(w_dff_A_fmEMOViY1_1),.din(w_dff_A_eDYUT59i0_1),.clk(gclk));
	jdff dff_A_05lP8yaM7_1(.dout(w_dff_A_eDYUT59i0_1),.din(w_dff_A_05lP8yaM7_1),.clk(gclk));
	jdff dff_B_7UJZZigs3_1(.din(n144),.dout(w_dff_B_7UJZZigs3_1),.clk(gclk));
	jdff dff_B_RpTxSUap7_1(.din(w_dff_B_7UJZZigs3_1),.dout(w_dff_B_RpTxSUap7_1),.clk(gclk));
	jdff dff_A_6abGK1HB3_0(.dout(w_G131_0[0]),.din(w_dff_A_6abGK1HB3_0),.clk(gclk));
	jdff dff_A_hoSnWOJF9_0(.dout(w_dff_A_6abGK1HB3_0),.din(w_dff_A_hoSnWOJF9_0),.clk(gclk));
	jdff dff_A_M1pWkXlx1_0(.dout(w_dff_A_hoSnWOJF9_0),.din(w_dff_A_M1pWkXlx1_0),.clk(gclk));
	jdff dff_A_XEpaEkmy8_0(.dout(w_dff_A_M1pWkXlx1_0),.din(w_dff_A_XEpaEkmy8_0),.clk(gclk));
	jdff dff_A_iLf9I2Gs5_0(.dout(w_dff_A_XEpaEkmy8_0),.din(w_dff_A_iLf9I2Gs5_0),.clk(gclk));
	jdff dff_A_9YUT2xh85_0(.dout(w_dff_A_iLf9I2Gs5_0),.din(w_dff_A_9YUT2xh85_0),.clk(gclk));
	jdff dff_A_6ako0U6V3_0(.dout(w_dff_A_9YUT2xh85_0),.din(w_dff_A_6ako0U6V3_0),.clk(gclk));
	jdff dff_A_jXzzJuGt6_0(.dout(w_dff_A_6ako0U6V3_0),.din(w_dff_A_jXzzJuGt6_0),.clk(gclk));
	jdff dff_A_y0Az1ZHM7_0(.dout(w_dff_A_jXzzJuGt6_0),.din(w_dff_A_y0Az1ZHM7_0),.clk(gclk));
	jdff dff_A_IT8zjJY29_0(.dout(w_dff_A_y0Az1ZHM7_0),.din(w_dff_A_IT8zjJY29_0),.clk(gclk));
	jdff dff_A_UCtd2EQc3_0(.dout(w_dff_A_IT8zjJY29_0),.din(w_dff_A_UCtd2EQc3_0),.clk(gclk));
	jdff dff_A_kWJYUDkj6_2(.dout(w_G131_0[2]),.din(w_dff_A_kWJYUDkj6_2),.clk(gclk));
	jdff dff_A_YMmS6L9s1_1(.dout(w_G953_2[1]),.din(w_dff_A_YMmS6L9s1_1),.clk(gclk));
	jdff dff_A_smhmllAO2_1(.dout(w_G214_0[1]),.din(w_dff_A_smhmllAO2_1),.clk(gclk));
	jdff dff_A_zFmTtjw79_0(.dout(w_n67_0[0]),.din(w_dff_A_zFmTtjw79_0),.clk(gclk));
	jdff dff_A_AuvSAvHW6_0(.dout(w_n66_0[0]),.din(w_dff_A_AuvSAvHW6_0),.clk(gclk));
	jdff dff_A_YZJPXvwV8_0(.dout(w_dff_A_AuvSAvHW6_0),.din(w_dff_A_YZJPXvwV8_0),.clk(gclk));
	jdff dff_A_ObWUNuaj5_0(.dout(w_G140_0[0]),.din(w_dff_A_ObWUNuaj5_0),.clk(gclk));
	jdff dff_A_jFmNtVyD2_0(.dout(w_dff_A_ObWUNuaj5_0),.din(w_dff_A_jFmNtVyD2_0),.clk(gclk));
	jdff dff_A_uVJug44B3_0(.dout(w_dff_A_jFmNtVyD2_0),.din(w_dff_A_uVJug44B3_0),.clk(gclk));
	jdff dff_A_O4VLiglz5_0(.dout(w_dff_A_uVJug44B3_0),.din(w_dff_A_O4VLiglz5_0),.clk(gclk));
	jdff dff_A_AkCyC8ka5_0(.dout(w_dff_A_O4VLiglz5_0),.din(w_dff_A_AkCyC8ka5_0),.clk(gclk));
	jdff dff_A_kN6ymnwt2_0(.dout(w_dff_A_AkCyC8ka5_0),.din(w_dff_A_kN6ymnwt2_0),.clk(gclk));
	jdff dff_A_MPRMm5fR2_0(.dout(w_dff_A_kN6ymnwt2_0),.din(w_dff_A_MPRMm5fR2_0),.clk(gclk));
	jdff dff_A_IKjUIpAw9_0(.dout(w_dff_A_MPRMm5fR2_0),.din(w_dff_A_IKjUIpAw9_0),.clk(gclk));
	jdff dff_A_slcVONpW6_0(.dout(w_dff_A_IKjUIpAw9_0),.din(w_dff_A_slcVONpW6_0),.clk(gclk));
	jdff dff_A_o9s3hDUl8_0(.dout(w_dff_A_slcVONpW6_0),.din(w_dff_A_o9s3hDUl8_0),.clk(gclk));
	jdff dff_A_n6GAev5Y8_0(.dout(w_dff_A_o9s3hDUl8_0),.din(w_dff_A_n6GAev5Y8_0),.clk(gclk));
	jdff dff_A_6GQaVU096_1(.dout(w_G140_0[1]),.din(w_dff_A_6GQaVU096_1),.clk(gclk));
	jdff dff_A_iUAE4Xef2_0(.dout(w_G125_0[0]),.din(w_dff_A_iUAE4Xef2_0),.clk(gclk));
	jdff dff_A_gYmzkazS2_0(.dout(w_dff_A_iUAE4Xef2_0),.din(w_dff_A_gYmzkazS2_0),.clk(gclk));
	jdff dff_A_YiaGsrrI9_0(.dout(w_dff_A_gYmzkazS2_0),.din(w_dff_A_YiaGsrrI9_0),.clk(gclk));
	jdff dff_A_qEcDgUcA5_0(.dout(w_dff_A_YiaGsrrI9_0),.din(w_dff_A_qEcDgUcA5_0),.clk(gclk));
	jdff dff_A_pgvuoAmg9_0(.dout(w_dff_A_qEcDgUcA5_0),.din(w_dff_A_pgvuoAmg9_0),.clk(gclk));
	jdff dff_A_sLveICmz3_0(.dout(w_dff_A_pgvuoAmg9_0),.din(w_dff_A_sLveICmz3_0),.clk(gclk));
	jdff dff_A_E3qJyMaQ9_0(.dout(w_dff_A_sLveICmz3_0),.din(w_dff_A_E3qJyMaQ9_0),.clk(gclk));
	jdff dff_A_piWuwKyK9_0(.dout(w_dff_A_E3qJyMaQ9_0),.din(w_dff_A_piWuwKyK9_0),.clk(gclk));
	jdff dff_A_vIvjCqFI3_0(.dout(w_dff_A_piWuwKyK9_0),.din(w_dff_A_vIvjCqFI3_0),.clk(gclk));
	jdff dff_A_x4Y6JPWi6_0(.dout(w_dff_A_vIvjCqFI3_0),.din(w_dff_A_x4Y6JPWi6_0),.clk(gclk));
	jdff dff_A_7Z5JpQnk7_0(.dout(w_dff_A_x4Y6JPWi6_0),.din(w_dff_A_7Z5JpQnk7_0),.clk(gclk));
	jdff dff_A_fOjlT9f56_1(.dout(w_G125_0[1]),.din(w_dff_A_fOjlT9f56_1),.clk(gclk));
	jdff dff_A_L4xYoWA20_1(.dout(w_dff_A_fOjlT9f56_1),.din(w_dff_A_L4xYoWA20_1),.clk(gclk));
	jdff dff_A_JKeSEgmt2_0(.dout(w_G146_0[0]),.din(w_dff_A_JKeSEgmt2_0),.clk(gclk));
	jdff dff_A_0oWuuqk64_0(.dout(w_dff_A_JKeSEgmt2_0),.din(w_dff_A_0oWuuqk64_0),.clk(gclk));
	jdff dff_A_mwKgX20g9_0(.dout(w_dff_A_0oWuuqk64_0),.din(w_dff_A_mwKgX20g9_0),.clk(gclk));
	jdff dff_A_bZol1qMW1_0(.dout(w_dff_A_mwKgX20g9_0),.din(w_dff_A_bZol1qMW1_0),.clk(gclk));
	jdff dff_A_M7Eav1Li4_0(.dout(w_dff_A_bZol1qMW1_0),.din(w_dff_A_M7Eav1Li4_0),.clk(gclk));
	jdff dff_A_Uiorhndm8_0(.dout(w_dff_A_M7Eav1Li4_0),.din(w_dff_A_Uiorhndm8_0),.clk(gclk));
	jdff dff_A_vPPoHPEg1_0(.dout(w_dff_A_Uiorhndm8_0),.din(w_dff_A_vPPoHPEg1_0),.clk(gclk));
	jdff dff_A_C0sjlLTX4_0(.dout(w_dff_A_vPPoHPEg1_0),.din(w_dff_A_C0sjlLTX4_0),.clk(gclk));
	jdff dff_A_MJ64zJmb7_0(.dout(w_dff_A_C0sjlLTX4_0),.din(w_dff_A_MJ64zJmb7_0),.clk(gclk));
	jdff dff_A_LqyqEvkk1_0(.dout(w_dff_A_MJ64zJmb7_0),.din(w_dff_A_LqyqEvkk1_0),.clk(gclk));
	jdff dff_B_tDf7LaZP8_3(.din(G146),.dout(w_dff_B_tDf7LaZP8_3),.clk(gclk));
	jdff dff_A_1ci5hxao0_0(.dout(w_G113_0[0]),.din(w_dff_A_1ci5hxao0_0),.clk(gclk));
	jdff dff_A_17BTM5Yb1_0(.dout(w_dff_A_1ci5hxao0_0),.din(w_dff_A_17BTM5Yb1_0),.clk(gclk));
	jdff dff_A_cuQw0M3q5_0(.dout(w_dff_A_17BTM5Yb1_0),.din(w_dff_A_cuQw0M3q5_0),.clk(gclk));
	jdff dff_A_uoyEAyqJ2_0(.dout(w_dff_A_cuQw0M3q5_0),.din(w_dff_A_uoyEAyqJ2_0),.clk(gclk));
	jdff dff_A_JpVJFe6h4_0(.dout(w_dff_A_uoyEAyqJ2_0),.din(w_dff_A_JpVJFe6h4_0),.clk(gclk));
	jdff dff_A_Ho1MDuCO0_0(.dout(w_dff_A_JpVJFe6h4_0),.din(w_dff_A_Ho1MDuCO0_0),.clk(gclk));
	jdff dff_A_J9OsFp8x5_0(.dout(w_dff_A_Ho1MDuCO0_0),.din(w_dff_A_J9OsFp8x5_0),.clk(gclk));
	jdff dff_A_Fqq7HPkV7_0(.dout(w_dff_A_J9OsFp8x5_0),.din(w_dff_A_Fqq7HPkV7_0),.clk(gclk));
	jdff dff_A_JNmo33VS1_0(.dout(w_dff_A_Fqq7HPkV7_0),.din(w_dff_A_JNmo33VS1_0),.clk(gclk));
	jdff dff_A_VTqvuAUF2_0(.dout(w_dff_A_JNmo33VS1_0),.din(w_dff_A_VTqvuAUF2_0),.clk(gclk));
	jdff dff_A_KDlWnTBC2_0(.dout(w_dff_A_VTqvuAUF2_0),.din(w_dff_A_KDlWnTBC2_0),.clk(gclk));
	jdff dff_A_7cswBw1t9_0(.dout(w_G104_0[0]),.din(w_dff_A_7cswBw1t9_0),.clk(gclk));
	jdff dff_A_d5GERTO76_0(.dout(w_dff_A_7cswBw1t9_0),.din(w_dff_A_d5GERTO76_0),.clk(gclk));
	jdff dff_A_eEk1WIa76_0(.dout(w_dff_A_d5GERTO76_0),.din(w_dff_A_eEk1WIa76_0),.clk(gclk));
	jdff dff_A_7C97W6zW1_0(.dout(w_dff_A_eEk1WIa76_0),.din(w_dff_A_7C97W6zW1_0),.clk(gclk));
	jdff dff_A_DrSQHbmK8_0(.dout(w_dff_A_7C97W6zW1_0),.din(w_dff_A_DrSQHbmK8_0),.clk(gclk));
	jdff dff_A_lErC70C12_0(.dout(w_dff_A_DrSQHbmK8_0),.din(w_dff_A_lErC70C12_0),.clk(gclk));
	jdff dff_A_znjD7QcY3_0(.dout(w_dff_A_lErC70C12_0),.din(w_dff_A_znjD7QcY3_0),.clk(gclk));
	jdff dff_A_3ipr91Wf5_0(.dout(w_dff_A_znjD7QcY3_0),.din(w_dff_A_3ipr91Wf5_0),.clk(gclk));
	jdff dff_A_TzPKrYpL1_0(.dout(w_dff_A_3ipr91Wf5_0),.din(w_dff_A_TzPKrYpL1_0),.clk(gclk));
	jdff dff_A_AXWvgzbM5_0(.dout(w_dff_A_TzPKrYpL1_0),.din(w_dff_A_AXWvgzbM5_0),.clk(gclk));
	jdff dff_A_QxyRqpiz9_0(.dout(w_dff_A_AXWvgzbM5_0),.din(w_dff_A_QxyRqpiz9_0),.clk(gclk));
	jdff dff_A_UXNkOvNP1_1(.dout(w_G104_0[1]),.din(w_dff_A_UXNkOvNP1_1),.clk(gclk));
	jdff dff_A_eRzFMcPL9_1(.dout(w_G475_0[1]),.din(w_dff_A_eRzFMcPL9_1),.clk(gclk));
	jdff dff_A_bfN0Q0R15_1(.dout(w_dff_A_eRzFMcPL9_1),.din(w_dff_A_bfN0Q0R15_1),.clk(gclk));
	jdff dff_A_fCpVzSGy4_1(.dout(w_dff_A_bfN0Q0R15_1),.din(w_dff_A_fCpVzSGy4_1),.clk(gclk));
	jdff dff_A_BdXfqQ4o7_1(.dout(w_dff_A_fCpVzSGy4_1),.din(w_dff_A_BdXfqQ4o7_1),.clk(gclk));
	jdff dff_A_u6rrTcFq6_1(.dout(w_dff_A_BdXfqQ4o7_1),.din(w_dff_A_u6rrTcFq6_1),.clk(gclk));
	jdff dff_A_UuWofEKp8_1(.dout(w_dff_A_u6rrTcFq6_1),.din(w_dff_A_UuWofEKp8_1),.clk(gclk));
	jdff dff_A_yoCtgT8M5_0(.dout(w_n139_0[0]),.din(w_dff_A_yoCtgT8M5_0),.clk(gclk));
	jdff dff_A_WkwsjzLT5_0(.dout(w_dff_A_yoCtgT8M5_0),.din(w_dff_A_WkwsjzLT5_0),.clk(gclk));
	jdff dff_A_kvNusFHk3_0(.dout(w_dff_A_WkwsjzLT5_0),.din(w_dff_A_kvNusFHk3_0),.clk(gclk));
	jdff dff_A_Bi6OkHbp1_0(.dout(w_dff_A_kvNusFHk3_0),.din(w_dff_A_Bi6OkHbp1_0),.clk(gclk));
	jdff dff_A_omCrb17u3_0(.dout(w_dff_A_Bi6OkHbp1_0),.din(w_dff_A_omCrb17u3_0),.clk(gclk));
	jdff dff_A_6ZJLDOnL9_0(.dout(w_dff_A_omCrb17u3_0),.din(w_dff_A_6ZJLDOnL9_0),.clk(gclk));
	jdff dff_A_lQ5MsYHa4_0(.dout(w_dff_A_6ZJLDOnL9_0),.din(w_dff_A_lQ5MsYHa4_0),.clk(gclk));
	jdff dff_A_AoqoFddy4_0(.dout(w_dff_A_lQ5MsYHa4_0),.din(w_dff_A_AoqoFddy4_0),.clk(gclk));
	jdff dff_A_Vramqusf3_0(.dout(w_dff_A_AoqoFddy4_0),.din(w_dff_A_Vramqusf3_0),.clk(gclk));
	jdff dff_A_ExHkzXRH6_0(.dout(w_dff_A_Vramqusf3_0),.din(w_dff_A_ExHkzXRH6_0),.clk(gclk));
	jdff dff_A_tBfZmiO65_0(.dout(w_dff_A_ExHkzXRH6_0),.din(w_dff_A_tBfZmiO65_0),.clk(gclk));
	jdff dff_A_SfD5si6v2_0(.dout(w_dff_A_tBfZmiO65_0),.din(w_dff_A_SfD5si6v2_0),.clk(gclk));
	jdff dff_A_sOCpEAii1_0(.dout(w_dff_A_SfD5si6v2_0),.din(w_dff_A_sOCpEAii1_0),.clk(gclk));
	jdff dff_B_AaC27EVr9_1(.din(n133),.dout(w_dff_B_AaC27EVr9_1),.clk(gclk));
	jdff dff_B_rGJeMbm67_1(.din(w_dff_B_AaC27EVr9_1),.dout(w_dff_B_rGJeMbm67_1),.clk(gclk));
	jdff dff_B_0KLhEgVX2_0(.din(n137),.dout(w_dff_B_0KLhEgVX2_0),.clk(gclk));
	jdff dff_A_FJcUi0DD7_1(.dout(w_G122_0[1]),.din(w_dff_A_FJcUi0DD7_1),.clk(gclk));
	jdff dff_A_zOU00Jo50_1(.dout(w_dff_A_FJcUi0DD7_1),.din(w_dff_A_zOU00Jo50_1),.clk(gclk));
	jdff dff_A_uFRrlYmx5_1(.dout(w_dff_A_zOU00Jo50_1),.din(w_dff_A_uFRrlYmx5_1),.clk(gclk));
	jdff dff_A_HNWrLLCV9_1(.dout(w_dff_A_uFRrlYmx5_1),.din(w_dff_A_HNWrLLCV9_1),.clk(gclk));
	jdff dff_A_8pJLPnNb8_1(.dout(w_dff_A_HNWrLLCV9_1),.din(w_dff_A_8pJLPnNb8_1),.clk(gclk));
	jdff dff_A_lpQKkEot6_1(.dout(w_dff_A_8pJLPnNb8_1),.din(w_dff_A_lpQKkEot6_1),.clk(gclk));
	jdff dff_A_fUfjc2Nt5_1(.dout(w_dff_A_lpQKkEot6_1),.din(w_dff_A_fUfjc2Nt5_1),.clk(gclk));
	jdff dff_A_xzjcm0HP9_1(.dout(w_dff_A_fUfjc2Nt5_1),.din(w_dff_A_xzjcm0HP9_1),.clk(gclk));
	jdff dff_A_pV7U0BwU0_1(.dout(w_dff_A_xzjcm0HP9_1),.din(w_dff_A_pV7U0BwU0_1),.clk(gclk));
	jdff dff_A_1StxXajN7_1(.dout(w_dff_A_pV7U0BwU0_1),.din(w_dff_A_1StxXajN7_1),.clk(gclk));
	jdff dff_A_yJRJj9yl0_1(.dout(w_dff_A_1StxXajN7_1),.din(w_dff_A_yJRJj9yl0_1),.clk(gclk));
	jdff dff_A_uAcqtmzT1_1(.dout(w_dff_A_yJRJj9yl0_1),.din(w_dff_A_uAcqtmzT1_1),.clk(gclk));
	jdff dff_A_CGPkWkbw4_0(.dout(w_G116_0[0]),.din(w_dff_A_CGPkWkbw4_0),.clk(gclk));
	jdff dff_A_rxo7xlto1_0(.dout(w_dff_A_CGPkWkbw4_0),.din(w_dff_A_rxo7xlto1_0),.clk(gclk));
	jdff dff_A_VQGxGIqE0_0(.dout(w_dff_A_rxo7xlto1_0),.din(w_dff_A_VQGxGIqE0_0),.clk(gclk));
	jdff dff_A_AMgOlEnP1_0(.dout(w_dff_A_VQGxGIqE0_0),.din(w_dff_A_AMgOlEnP1_0),.clk(gclk));
	jdff dff_A_9vKkCo9I6_0(.dout(w_dff_A_AMgOlEnP1_0),.din(w_dff_A_9vKkCo9I6_0),.clk(gclk));
	jdff dff_A_gZimZZuF4_0(.dout(w_dff_A_9vKkCo9I6_0),.din(w_dff_A_gZimZZuF4_0),.clk(gclk));
	jdff dff_A_Ze4lYX293_0(.dout(w_dff_A_gZimZZuF4_0),.din(w_dff_A_Ze4lYX293_0),.clk(gclk));
	jdff dff_A_YADflOyV4_0(.dout(w_dff_A_Ze4lYX293_0),.din(w_dff_A_YADflOyV4_0),.clk(gclk));
	jdff dff_A_Jje4ToyZ2_0(.dout(w_dff_A_YADflOyV4_0),.din(w_dff_A_Jje4ToyZ2_0),.clk(gclk));
	jdff dff_A_eyyGZype4_0(.dout(w_dff_A_Jje4ToyZ2_0),.din(w_dff_A_eyyGZype4_0),.clk(gclk));
	jdff dff_A_rvYggMYV9_0(.dout(w_dff_A_eyyGZype4_0),.din(w_dff_A_rvYggMYV9_0),.clk(gclk));
	jdff dff_A_4EsmdIrz9_0(.dout(w_G107_0[0]),.din(w_dff_A_4EsmdIrz9_0),.clk(gclk));
	jdff dff_A_Kuba5AAk3_0(.dout(w_dff_A_4EsmdIrz9_0),.din(w_dff_A_Kuba5AAk3_0),.clk(gclk));
	jdff dff_A_pE3Qa32p8_0(.dout(w_dff_A_Kuba5AAk3_0),.din(w_dff_A_pE3Qa32p8_0),.clk(gclk));
	jdff dff_A_6iiqElcM2_0(.dout(w_dff_A_pE3Qa32p8_0),.din(w_dff_A_6iiqElcM2_0),.clk(gclk));
	jdff dff_A_Af1fojlL4_0(.dout(w_dff_A_6iiqElcM2_0),.din(w_dff_A_Af1fojlL4_0),.clk(gclk));
	jdff dff_A_cl0m71280_0(.dout(w_dff_A_Af1fojlL4_0),.din(w_dff_A_cl0m71280_0),.clk(gclk));
	jdff dff_A_bNj1RzFi8_0(.dout(w_dff_A_cl0m71280_0),.din(w_dff_A_bNj1RzFi8_0),.clk(gclk));
	jdff dff_A_iaoM9yXH4_0(.dout(w_dff_A_bNj1RzFi8_0),.din(w_dff_A_iaoM9yXH4_0),.clk(gclk));
	jdff dff_A_QrVaYf3R7_0(.dout(w_dff_A_iaoM9yXH4_0),.din(w_dff_A_QrVaYf3R7_0),.clk(gclk));
	jdff dff_A_ZaSg8bTT6_0(.dout(w_dff_A_QrVaYf3R7_0),.din(w_dff_A_ZaSg8bTT6_0),.clk(gclk));
	jdff dff_A_7X63bgxk9_0(.dout(w_dff_A_ZaSg8bTT6_0),.din(w_dff_A_7X63bgxk9_0),.clk(gclk));
	jdff dff_A_4yWwIPGb3_1(.dout(w_G107_0[1]),.din(w_dff_A_4yWwIPGb3_1),.clk(gclk));
	jdff dff_A_LCBQVhYw9_2(.dout(w_n103_2[2]),.din(w_dff_A_LCBQVhYw9_2),.clk(gclk));
	jdff dff_A_8Riq3MXW9_2(.dout(w_dff_A_LCBQVhYw9_2),.din(w_dff_A_8Riq3MXW9_2),.clk(gclk));
	jdff dff_A_QulWFVfe7_1(.dout(w_G234_0[1]),.din(w_dff_A_QulWFVfe7_1),.clk(gclk));
	jdff dff_A_LHdbYX1l4_0(.dout(w_G217_0[0]),.din(w_dff_A_LHdbYX1l4_0),.clk(gclk));
	jdff dff_A_fgM0rRkI3_0(.dout(w_dff_A_LHdbYX1l4_0),.din(w_dff_A_fgM0rRkI3_0),.clk(gclk));
	jdff dff_A_9MRPvmYd4_0(.dout(w_dff_A_fgM0rRkI3_0),.din(w_dff_A_9MRPvmYd4_0),.clk(gclk));
	jdff dff_A_thdJSFsO7_0(.dout(w_dff_A_9MRPvmYd4_0),.din(w_dff_A_thdJSFsO7_0),.clk(gclk));
	jdff dff_A_QCy9DNjg5_0(.dout(w_dff_A_thdJSFsO7_0),.din(w_dff_A_QCy9DNjg5_0),.clk(gclk));
	jdff dff_A_xLKU9s3N0_0(.dout(w_dff_A_QCy9DNjg5_0),.din(w_dff_A_xLKU9s3N0_0),.clk(gclk));
	jdff dff_A_gigbAQeI1_0(.dout(w_dff_A_xLKU9s3N0_0),.din(w_dff_A_gigbAQeI1_0),.clk(gclk));
	jdff dff_A_y6u6BAZH1_0(.dout(w_dff_A_gigbAQeI1_0),.din(w_dff_A_y6u6BAZH1_0),.clk(gclk));
	jdff dff_A_xxpNAW7v3_0(.dout(w_dff_A_y6u6BAZH1_0),.din(w_dff_A_xxpNAW7v3_0),.clk(gclk));
	jdff dff_A_O2cWDeTR9_0(.dout(w_dff_A_xxpNAW7v3_0),.din(w_dff_A_O2cWDeTR9_0),.clk(gclk));
	jdff dff_A_qaqcQl2I7_0(.dout(w_dff_A_O2cWDeTR9_0),.din(w_dff_A_qaqcQl2I7_0),.clk(gclk));
	jdff dff_A_Hi1Blwi94_0(.dout(w_dff_A_qaqcQl2I7_0),.din(w_dff_A_Hi1Blwi94_0),.clk(gclk));
	jdff dff_A_95ypSuxk4_0(.dout(w_dff_A_Hi1Blwi94_0),.din(w_dff_A_95ypSuxk4_0),.clk(gclk));
	jdff dff_A_MWoF7v4d9_0(.dout(w_dff_A_95ypSuxk4_0),.din(w_dff_A_MWoF7v4d9_0),.clk(gclk));
	jdff dff_A_u45MO1NO5_2(.dout(w_G217_0[2]),.din(w_dff_A_u45MO1NO5_2),.clk(gclk));
	jdff dff_B_dBsVMmw73_3(.din(G217),.dout(w_dff_B_dBsVMmw73_3),.clk(gclk));
	jdff dff_B_n2egPD6k4_3(.din(w_dff_B_dBsVMmw73_3),.dout(w_dff_B_n2egPD6k4_3),.clk(gclk));
	jdff dff_A_5vbmP3rN7_0(.dout(w_G143_0[0]),.din(w_dff_A_5vbmP3rN7_0),.clk(gclk));
	jdff dff_A_r0TRfFGO6_0(.dout(w_dff_A_5vbmP3rN7_0),.din(w_dff_A_r0TRfFGO6_0),.clk(gclk));
	jdff dff_A_wwTKFn1p7_0(.dout(w_dff_A_r0TRfFGO6_0),.din(w_dff_A_wwTKFn1p7_0),.clk(gclk));
	jdff dff_A_3HY76bT19_0(.dout(w_dff_A_wwTKFn1p7_0),.din(w_dff_A_3HY76bT19_0),.clk(gclk));
	jdff dff_A_43RCmt4a0_0(.dout(w_dff_A_3HY76bT19_0),.din(w_dff_A_43RCmt4a0_0),.clk(gclk));
	jdff dff_A_8BX39smi2_0(.dout(w_dff_A_43RCmt4a0_0),.din(w_dff_A_8BX39smi2_0),.clk(gclk));
	jdff dff_A_z8q9eX0b6_0(.dout(w_dff_A_8BX39smi2_0),.din(w_dff_A_z8q9eX0b6_0),.clk(gclk));
	jdff dff_A_12hBlNlt8_0(.dout(w_dff_A_z8q9eX0b6_0),.din(w_dff_A_12hBlNlt8_0),.clk(gclk));
	jdff dff_A_9CADTxuV0_0(.dout(w_dff_A_12hBlNlt8_0),.din(w_dff_A_9CADTxuV0_0),.clk(gclk));
	jdff dff_A_BhggG4sV1_0(.dout(w_dff_A_9CADTxuV0_0),.din(w_dff_A_BhggG4sV1_0),.clk(gclk));
	jdff dff_A_oEciDPoY5_0(.dout(w_dff_A_BhggG4sV1_0),.din(w_dff_A_oEciDPoY5_0),.clk(gclk));
	jdff dff_A_t0QOJokZ5_1(.dout(w_G143_0[1]),.din(w_dff_A_t0QOJokZ5_1),.clk(gclk));
	jdff dff_A_Wk3nflXf8_0(.dout(w_G128_0[0]),.din(w_dff_A_Wk3nflXf8_0),.clk(gclk));
	jdff dff_A_AcqzBmno9_0(.dout(w_dff_A_Wk3nflXf8_0),.din(w_dff_A_AcqzBmno9_0),.clk(gclk));
	jdff dff_A_ke57k9Ly9_0(.dout(w_dff_A_AcqzBmno9_0),.din(w_dff_A_ke57k9Ly9_0),.clk(gclk));
	jdff dff_A_JzS1N3x26_0(.dout(w_dff_A_ke57k9Ly9_0),.din(w_dff_A_JzS1N3x26_0),.clk(gclk));
	jdff dff_A_ITmY9NBD9_0(.dout(w_dff_A_JzS1N3x26_0),.din(w_dff_A_ITmY9NBD9_0),.clk(gclk));
	jdff dff_A_CoCJX8gk1_0(.dout(w_dff_A_ITmY9NBD9_0),.din(w_dff_A_CoCJX8gk1_0),.clk(gclk));
	jdff dff_A_XuS2VIxY7_0(.dout(w_dff_A_CoCJX8gk1_0),.din(w_dff_A_XuS2VIxY7_0),.clk(gclk));
	jdff dff_A_L2ye1Ak59_0(.dout(w_dff_A_XuS2VIxY7_0),.din(w_dff_A_L2ye1Ak59_0),.clk(gclk));
	jdff dff_A_NEO4XSwV2_0(.dout(w_dff_A_L2ye1Ak59_0),.din(w_dff_A_NEO4XSwV2_0),.clk(gclk));
	jdff dff_A_cKt2JESH7_0(.dout(w_dff_A_NEO4XSwV2_0),.din(w_dff_A_cKt2JESH7_0),.clk(gclk));
	jdff dff_A_jj354q4q8_0(.dout(w_dff_A_cKt2JESH7_0),.din(w_dff_A_jj354q4q8_0),.clk(gclk));
	jdff dff_A_wpf09Gme3_0(.dout(w_G134_0[0]),.din(w_dff_A_wpf09Gme3_0),.clk(gclk));
	jdff dff_A_MxM8sEm29_0(.dout(w_dff_A_wpf09Gme3_0),.din(w_dff_A_MxM8sEm29_0),.clk(gclk));
	jdff dff_A_pEwiFNb82_0(.dout(w_dff_A_MxM8sEm29_0),.din(w_dff_A_pEwiFNb82_0),.clk(gclk));
	jdff dff_A_MV6gKf3u8_0(.dout(w_dff_A_pEwiFNb82_0),.din(w_dff_A_MV6gKf3u8_0),.clk(gclk));
	jdff dff_A_Kp4fMU0B1_0(.dout(w_dff_A_MV6gKf3u8_0),.din(w_dff_A_Kp4fMU0B1_0),.clk(gclk));
	jdff dff_A_oeQf53br4_0(.dout(w_dff_A_Kp4fMU0B1_0),.din(w_dff_A_oeQf53br4_0),.clk(gclk));
	jdff dff_A_O1R10r377_0(.dout(w_dff_A_oeQf53br4_0),.din(w_dff_A_O1R10r377_0),.clk(gclk));
	jdff dff_A_Ux2feFDC8_0(.dout(w_dff_A_O1R10r377_0),.din(w_dff_A_Ux2feFDC8_0),.clk(gclk));
	jdff dff_A_B6l5WYiX2_0(.dout(w_dff_A_Ux2feFDC8_0),.din(w_dff_A_B6l5WYiX2_0),.clk(gclk));
	jdff dff_A_OZdOeCCq2_0(.dout(w_dff_A_B6l5WYiX2_0),.din(w_dff_A_OZdOeCCq2_0),.clk(gclk));
	jdff dff_A_bDdjKQWW9_0(.dout(w_dff_A_OZdOeCCq2_0),.din(w_dff_A_bDdjKQWW9_0),.clk(gclk));
	jdff dff_A_Vr5KbPGm8_1(.dout(w_G134_0[1]),.din(w_dff_A_Vr5KbPGm8_1),.clk(gclk));
	jdff dff_A_JOXvNFby4_0(.dout(w_n58_0[0]),.din(w_dff_A_JOXvNFby4_0),.clk(gclk));
	jdff dff_A_b8WsRpQW0_0(.dout(w_dff_A_JOXvNFby4_0),.din(w_dff_A_b8WsRpQW0_0),.clk(gclk));
	jdff dff_A_WxXg8hHp6_0(.dout(w_dff_A_b8WsRpQW0_0),.din(w_dff_A_WxXg8hHp6_0),.clk(gclk));
	jdff dff_A_iqkRzPY84_0(.dout(w_dff_A_WxXg8hHp6_0),.din(w_dff_A_iqkRzPY84_0),.clk(gclk));
	jdff dff_A_CfEJDDX21_2(.dout(w_n58_0[2]),.din(w_dff_A_CfEJDDX21_2),.clk(gclk));
	jdff dff_A_pErA9So75_2(.dout(w_dff_A_CfEJDDX21_2),.din(w_dff_A_pErA9So75_2),.clk(gclk));
	jdff dff_A_2SsQnHsJ0_2(.dout(w_dff_A_pErA9So75_2),.din(w_dff_A_2SsQnHsJ0_2),.clk(gclk));
	jdff dff_A_3N0rDgif6_2(.dout(w_dff_A_2SsQnHsJ0_2),.din(w_dff_A_3N0rDgif6_2),.clk(gclk));
	jdff dff_A_thEhU3rG8_0(.dout(w_G902_3[0]),.din(w_dff_A_thEhU3rG8_0),.clk(gclk));
	jdff dff_A_KuNoHgdm8_0(.dout(w_dff_A_thEhU3rG8_0),.din(w_dff_A_KuNoHgdm8_0),.clk(gclk));
	jdff dff_A_XO2NXqmB5_0(.dout(w_G478_0[0]),.din(w_dff_A_XO2NXqmB5_0),.clk(gclk));
	jdff dff_A_YLd838JQ1_0(.dout(w_dff_A_XO2NXqmB5_0),.din(w_dff_A_YLd838JQ1_0),.clk(gclk));
	jdff dff_A_Ejkc2pvE5_0(.dout(w_dff_A_YLd838JQ1_0),.din(w_dff_A_Ejkc2pvE5_0),.clk(gclk));
	jdff dff_A_GMhsnH2r1_0(.dout(w_dff_A_Ejkc2pvE5_0),.din(w_dff_A_GMhsnH2r1_0),.clk(gclk));
	jdff dff_A_kBaZRqQp3_0(.dout(w_dff_A_GMhsnH2r1_0),.din(w_dff_A_kBaZRqQp3_0),.clk(gclk));
	jdff dff_A_bq1snYzD8_0(.dout(w_dff_A_kBaZRqQp3_0),.din(w_dff_A_bq1snYzD8_0),.clk(gclk));
	jdff dff_A_UwmH1h3q7_0(.dout(w_dff_A_bq1snYzD8_0),.din(w_dff_A_UwmH1h3q7_0),.clk(gclk));
	jdff dff_A_PeW7kkMH5_0(.dout(w_dff_A_UwmH1h3q7_0),.din(w_dff_A_PeW7kkMH5_0),.clk(gclk));
	jdff dff_A_eWqVTP6h1_0(.dout(w_dff_A_PeW7kkMH5_0),.din(w_dff_A_eWqVTP6h1_0),.clk(gclk));
	jdff dff_A_Pnx97o5o3_0(.dout(w_dff_A_eWqVTP6h1_0),.din(w_dff_A_Pnx97o5o3_0),.clk(gclk));
	jdff dff_A_rTCldChL0_0(.dout(w_dff_A_Pnx97o5o3_0),.din(w_dff_A_rTCldChL0_0),.clk(gclk));
	jdff dff_A_sJGlKoZN8_0(.dout(w_dff_A_rTCldChL0_0),.din(w_dff_A_sJGlKoZN8_0),.clk(gclk));
	jdff dff_A_wT9ZA0bX7_0(.dout(w_dff_A_sJGlKoZN8_0),.din(w_dff_A_wT9ZA0bX7_0),.clk(gclk));
	jdff dff_A_8PN1S7Cr2_0(.dout(w_dff_A_wT9ZA0bX7_0),.din(w_dff_A_8PN1S7Cr2_0),.clk(gclk));
	jdff dff_A_uOmmawTv1_0(.dout(w_dff_A_8PN1S7Cr2_0),.din(w_dff_A_uOmmawTv1_0),.clk(gclk));
	jdff dff_A_B1BZUJ931_0(.dout(w_dff_A_uOmmawTv1_0),.din(w_dff_A_B1BZUJ931_0),.clk(gclk));
	jdff dff_A_ftPwKyxt3_1(.dout(w_G478_0[1]),.din(w_dff_A_ftPwKyxt3_1),.clk(gclk));
	jdff dff_A_icqAGQ2x4_1(.dout(w_dff_A_ftPwKyxt3_1),.din(w_dff_A_icqAGQ2x4_1),.clk(gclk));
	jdff dff_A_T2uWvyeP3_1(.dout(w_dff_A_icqAGQ2x4_1),.din(w_dff_A_T2uWvyeP3_1),.clk(gclk));
	jdff dff_A_9IYsCH6a3_1(.dout(w_dff_A_T2uWvyeP3_1),.din(w_dff_A_9IYsCH6a3_1),.clk(gclk));
	jdff dff_A_WDKiYE7a3_1(.dout(w_dff_A_9IYsCH6a3_1),.din(w_dff_A_WDKiYE7a3_1),.clk(gclk));
	jdff dff_A_cedgfwoZ5_1(.dout(w_dff_A_WDKiYE7a3_1),.din(w_dff_A_cedgfwoZ5_1),.clk(gclk));
	jdff dff_A_4bd6Wsb46_1(.dout(w_n265_0[1]),.din(w_dff_A_4bd6Wsb46_1),.clk(gclk));
	jdff dff_B_d5cNMmmd5_3(.din(n265),.dout(w_dff_B_d5cNMmmd5_3),.clk(gclk));
	jdff dff_B_kcAU56Im7_3(.din(w_dff_B_d5cNMmmd5_3),.dout(w_dff_B_kcAU56Im7_3),.clk(gclk));
	jdff dff_B_qMjLyACn1_3(.din(w_dff_B_kcAU56Im7_3),.dout(w_dff_B_qMjLyACn1_3),.clk(gclk));
	jdff dff_B_54y25HS31_3(.din(w_dff_B_qMjLyACn1_3),.dout(w_dff_B_54y25HS31_3),.clk(gclk));
	jdff dff_B_VJKDBgl72_3(.din(w_dff_B_54y25HS31_3),.dout(w_dff_B_VJKDBgl72_3),.clk(gclk));
	jdff dff_B_xxfKP00E7_3(.din(w_dff_B_VJKDBgl72_3),.dout(w_dff_B_xxfKP00E7_3),.clk(gclk));
	jdff dff_B_EweI4n6z5_3(.din(w_dff_B_xxfKP00E7_3),.dout(w_dff_B_EweI4n6z5_3),.clk(gclk));
	jdff dff_B_XGQkjbfn8_3(.din(w_dff_B_EweI4n6z5_3),.dout(w_dff_B_XGQkjbfn8_3),.clk(gclk));
	jdff dff_B_yRcC5K3y6_3(.din(w_dff_B_XGQkjbfn8_3),.dout(w_dff_B_yRcC5K3y6_3),.clk(gclk));
	jdff dff_B_dZvAHQZL0_3(.din(w_dff_B_yRcC5K3y6_3),.dout(w_dff_B_dZvAHQZL0_3),.clk(gclk));
	jdff dff_B_UxWMeUkp0_3(.din(w_dff_B_dZvAHQZL0_3),.dout(w_dff_B_UxWMeUkp0_3),.clk(gclk));
	jdff dff_B_zVYBvw3p7_3(.din(w_dff_B_UxWMeUkp0_3),.dout(w_dff_B_zVYBvw3p7_3),.clk(gclk));
	jdff dff_B_bs16xm1N2_3(.din(w_dff_B_zVYBvw3p7_3),.dout(w_dff_B_bs16xm1N2_3),.clk(gclk));
	jdff dff_B_750Cn1Mx1_3(.din(w_dff_B_bs16xm1N2_3),.dout(w_dff_B_750Cn1Mx1_3),.clk(gclk));
	jdff dff_B_GJGTG1B15_3(.din(w_dff_B_750Cn1Mx1_3),.dout(w_dff_B_GJGTG1B15_3),.clk(gclk));
	jdff dff_B_kDrnVLV79_3(.din(w_dff_B_GJGTG1B15_3),.dout(w_dff_B_kDrnVLV79_3),.clk(gclk));
	jdff dff_A_NVfBsJ6J2_0(.dout(w_G953_1[0]),.din(w_dff_A_NVfBsJ6J2_0),.clk(gclk));
	jdff dff_A_Z6XOJmfD6_0(.dout(w_dff_A_NVfBsJ6J2_0),.din(w_dff_A_Z6XOJmfD6_0),.clk(gclk));
	jdff dff_A_T6Iee2yQ4_0(.dout(w_dff_A_Z6XOJmfD6_0),.din(w_dff_A_T6Iee2yQ4_0),.clk(gclk));
	jdff dff_A_6TPWwDut0_0(.dout(w_dff_A_T6Iee2yQ4_0),.din(w_dff_A_6TPWwDut0_0),.clk(gclk));
	jdff dff_A_nDZu8GlS8_0(.dout(w_dff_A_6TPWwDut0_0),.din(w_dff_A_nDZu8GlS8_0),.clk(gclk));
	jdff dff_A_R4IHslOi1_0(.dout(w_dff_A_nDZu8GlS8_0),.din(w_dff_A_R4IHslOi1_0),.clk(gclk));
	jdff dff_A_dMTdSJT36_0(.dout(w_dff_A_R4IHslOi1_0),.din(w_dff_A_dMTdSJT36_0),.clk(gclk));
	jdff dff_A_T0rZJ28S7_0(.dout(w_dff_A_dMTdSJT36_0),.din(w_dff_A_T0rZJ28S7_0),.clk(gclk));
	jdff dff_A_u1sl0uzd4_0(.dout(w_dff_A_T0rZJ28S7_0),.din(w_dff_A_u1sl0uzd4_0),.clk(gclk));
	jdff dff_A_grOjI92V3_0(.dout(w_dff_A_u1sl0uzd4_0),.din(w_dff_A_grOjI92V3_0),.clk(gclk));
	jdff dff_A_Z0LdavpV1_0(.dout(w_dff_A_grOjI92V3_0),.din(w_dff_A_Z0LdavpV1_0),.clk(gclk));
	jdff dff_A_9n1cGunY0_0(.dout(w_dff_A_Z0LdavpV1_0),.din(w_dff_A_9n1cGunY0_0),.clk(gclk));
	jdff dff_A_AG6TQukn0_0(.dout(w_dff_A_9n1cGunY0_0),.din(w_dff_A_AG6TQukn0_0),.clk(gclk));
	jdff dff_A_6g4UUk1S4_0(.dout(w_dff_A_AG6TQukn0_0),.din(w_dff_A_6g4UUk1S4_0),.clk(gclk));
	jdff dff_A_d9VMHloT7_0(.dout(w_dff_A_6g4UUk1S4_0),.din(w_dff_A_d9VMHloT7_0),.clk(gclk));
	jdff dff_A_otwmZ7K66_1(.dout(w_G953_1[1]),.din(w_dff_A_otwmZ7K66_1),.clk(gclk));
	jdff dff_A_XsjyPbYo6_1(.dout(w_dff_A_otwmZ7K66_1),.din(w_dff_A_XsjyPbYo6_1),.clk(gclk));
	jdff dff_A_aYCwG2i71_1(.dout(w_dff_A_XsjyPbYo6_1),.din(w_dff_A_aYCwG2i71_1),.clk(gclk));
	jdff dff_A_n4rZm2Bp4_1(.dout(w_dff_A_aYCwG2i71_1),.din(w_dff_A_n4rZm2Bp4_1),.clk(gclk));
	jdff dff_A_eLjLWaAs6_1(.dout(w_dff_A_n4rZm2Bp4_1),.din(w_dff_A_eLjLWaAs6_1),.clk(gclk));
	jdff dff_A_eeTzjEih8_1(.dout(w_dff_A_eLjLWaAs6_1),.din(w_dff_A_eeTzjEih8_1),.clk(gclk));
	jdff dff_A_SpqyoD0C9_1(.dout(w_dff_A_eeTzjEih8_1),.din(w_dff_A_SpqyoD0C9_1),.clk(gclk));
	jdff dff_A_xzVgzlMI9_1(.dout(w_dff_A_SpqyoD0C9_1),.din(w_dff_A_xzVgzlMI9_1),.clk(gclk));
	jdff dff_A_Kc3zzDO38_1(.dout(w_dff_A_xzVgzlMI9_1),.din(w_dff_A_Kc3zzDO38_1),.clk(gclk));
	jdff dff_A_uZmpMZ9T5_1(.dout(w_dff_A_Kc3zzDO38_1),.din(w_dff_A_uZmpMZ9T5_1),.clk(gclk));
	jdff dff_A_2YidaYvC5_1(.dout(w_dff_A_uZmpMZ9T5_1),.din(w_dff_A_2YidaYvC5_1),.clk(gclk));
	jdff dff_A_gqVlawb97_1(.dout(w_dff_A_2YidaYvC5_1),.din(w_dff_A_gqVlawb97_1),.clk(gclk));
	jdff dff_A_pc9L0pIi1_2(.dout(w_G953_0[2]),.din(w_dff_A_pc9L0pIi1_2),.clk(gclk));
	jdff dff_A_eGx7f1Q51_2(.dout(w_dff_A_pc9L0pIi1_2),.din(w_dff_A_eGx7f1Q51_2),.clk(gclk));
	jdff dff_A_3DpWNDEr5_2(.dout(w_dff_A_eGx7f1Q51_2),.din(w_dff_A_3DpWNDEr5_2),.clk(gclk));
	jdff dff_A_PYxBVZhx8_2(.dout(w_dff_A_3DpWNDEr5_2),.din(w_dff_A_PYxBVZhx8_2),.clk(gclk));
	jdff dff_A_p2xDHb3t4_2(.dout(w_dff_A_PYxBVZhx8_2),.din(w_dff_A_p2xDHb3t4_2),.clk(gclk));
	jdff dff_A_AnDg3IFC8_2(.dout(w_dff_A_p2xDHb3t4_2),.din(w_dff_A_AnDg3IFC8_2),.clk(gclk));
	jdff dff_A_q927HUSt8_2(.dout(w_dff_A_AnDg3IFC8_2),.din(w_dff_A_q927HUSt8_2),.clk(gclk));
	jdff dff_A_clbAaZkK8_2(.dout(w_dff_A_q927HUSt8_2),.din(w_dff_A_clbAaZkK8_2),.clk(gclk));
	jdff dff_A_k2eO1p883_2(.dout(w_dff_A_clbAaZkK8_2),.din(w_dff_A_k2eO1p883_2),.clk(gclk));
	jdff dff_A_drC8dM9f7_2(.dout(w_dff_A_k2eO1p883_2),.din(w_dff_A_drC8dM9f7_2),.clk(gclk));
	jdff dff_A_znWjcgch0_2(.dout(w_dff_A_drC8dM9f7_2),.din(w_dff_A_znWjcgch0_2),.clk(gclk));
	jdff dff_A_UAAT1bQg5_2(.dout(w_dff_A_znWjcgch0_2),.din(w_dff_A_UAAT1bQg5_2),.clk(gclk));
	jdff dff_A_j2jZPvdg0_2(.dout(w_dff_A_UAAT1bQg5_2),.din(w_dff_A_j2jZPvdg0_2),.clk(gclk));
	jdff dff_A_DOKlR9un6_2(.dout(w_dff_A_j2jZPvdg0_2),.din(w_dff_A_DOKlR9un6_2),.clk(gclk));
	jdff dff_A_UYh1kpDt7_2(.dout(w_dff_A_DOKlR9un6_2),.din(w_dff_A_UYh1kpDt7_2),.clk(gclk));
	jdff dff_A_wfDsTIBL0_1(.dout(w_G952_0[1]),.din(w_dff_A_wfDsTIBL0_1),.clk(gclk));
	jdff dff_A_USSvfxsm4_1(.dout(w_dff_A_wfDsTIBL0_1),.din(w_dff_A_USSvfxsm4_1),.clk(gclk));
	jdff dff_A_V0WXk8xn0_1(.dout(w_dff_A_USSvfxsm4_1),.din(w_dff_A_V0WXk8xn0_1),.clk(gclk));
	jdff dff_A_ZXve7Bzx4_1(.dout(w_dff_A_V0WXk8xn0_1),.din(w_dff_A_ZXve7Bzx4_1),.clk(gclk));
	jdff dff_A_7gqzoWAo3_1(.dout(w_dff_A_ZXve7Bzx4_1),.din(w_dff_A_7gqzoWAo3_1),.clk(gclk));
	jdff dff_A_rRFgyQ5h6_1(.dout(w_dff_A_7gqzoWAo3_1),.din(w_dff_A_rRFgyQ5h6_1),.clk(gclk));
	jdff dff_A_ldKU0D3X9_1(.dout(w_dff_A_rRFgyQ5h6_1),.din(w_dff_A_ldKU0D3X9_1),.clk(gclk));
	jdff dff_A_YmuNw9wL0_1(.dout(w_dff_A_ldKU0D3X9_1),.din(w_dff_A_YmuNw9wL0_1),.clk(gclk));
	jdff dff_A_gkfyMVve2_1(.dout(w_dff_A_YmuNw9wL0_1),.din(w_dff_A_gkfyMVve2_1),.clk(gclk));
	jdff dff_A_szKKgWPo3_1(.dout(w_dff_A_gkfyMVve2_1),.din(w_dff_A_szKKgWPo3_1),.clk(gclk));
	jdff dff_A_QVy1HCwZ0_1(.dout(w_dff_A_szKKgWPo3_1),.din(w_dff_A_QVy1HCwZ0_1),.clk(gclk));
	jdff dff_A_SkXrW8Wj2_1(.dout(w_dff_A_QVy1HCwZ0_1),.din(w_dff_A_SkXrW8Wj2_1),.clk(gclk));
	jdff dff_A_hFdfcENc6_1(.dout(w_dff_A_SkXrW8Wj2_1),.din(w_dff_A_hFdfcENc6_1),.clk(gclk));
	jdff dff_A_UR7pucAm7_1(.dout(w_dff_A_hFdfcENc6_1),.din(w_dff_A_UR7pucAm7_1),.clk(gclk));
	jdff dff_A_pLDUt66Z5_1(.dout(w_dff_A_UR7pucAm7_1),.din(w_dff_A_pLDUt66Z5_1),.clk(gclk));
	jdff dff_A_V0Gna0CB6_1(.dout(w_dff_A_pLDUt66Z5_1),.din(w_dff_A_V0Gna0CB6_1),.clk(gclk));
	jdff dff_A_AiE7RKGB3_2(.dout(w_G952_0[2]),.din(w_dff_A_AiE7RKGB3_2),.clk(gclk));
	jdff dff_B_ncci2Lg17_3(.din(G952),.dout(w_dff_B_ncci2Lg17_3),.clk(gclk));
	jdff dff_A_rf43yoJL4_2(.dout(w_dff_A_DqQ4FdOr5_0),.din(w_dff_A_rf43yoJL4_2),.clk(gclk));
	jdff dff_A_DqQ4FdOr5_0(.dout(w_dff_A_t3mlupzd6_0),.din(w_dff_A_DqQ4FdOr5_0),.clk(gclk));
	jdff dff_A_t3mlupzd6_0(.dout(w_dff_A_JjbYlYQx7_0),.din(w_dff_A_t3mlupzd6_0),.clk(gclk));
	jdff dff_A_JjbYlYQx7_0(.dout(w_dff_A_rf9kPEQr9_0),.din(w_dff_A_JjbYlYQx7_0),.clk(gclk));
	jdff dff_A_rf9kPEQr9_0(.dout(w_dff_A_dDZMe9FQ2_0),.din(w_dff_A_rf9kPEQr9_0),.clk(gclk));
	jdff dff_A_dDZMe9FQ2_0(.dout(w_dff_A_tDd1w2bm6_0),.din(w_dff_A_dDZMe9FQ2_0),.clk(gclk));
	jdff dff_A_tDd1w2bm6_0(.dout(w_dff_A_vK3rWXzI0_0),.din(w_dff_A_tDd1w2bm6_0),.clk(gclk));
	jdff dff_A_vK3rWXzI0_0(.dout(G3),.din(w_dff_A_vK3rWXzI0_0),.clk(gclk));
	jdff dff_A_lBuhumSC3_2(.dout(w_dff_A_HSJIbGkF4_0),.din(w_dff_A_lBuhumSC3_2),.clk(gclk));
	jdff dff_A_HSJIbGkF4_0(.dout(w_dff_A_VG4lcelf3_0),.din(w_dff_A_HSJIbGkF4_0),.clk(gclk));
	jdff dff_A_VG4lcelf3_0(.dout(w_dff_A_lCnSg9Uv6_0),.din(w_dff_A_VG4lcelf3_0),.clk(gclk));
	jdff dff_A_lCnSg9Uv6_0(.dout(w_dff_A_jG2CR8sJ8_0),.din(w_dff_A_lCnSg9Uv6_0),.clk(gclk));
	jdff dff_A_jG2CR8sJ8_0(.dout(w_dff_A_e7giKlnW0_0),.din(w_dff_A_jG2CR8sJ8_0),.clk(gclk));
	jdff dff_A_e7giKlnW0_0(.dout(w_dff_A_PEIkaqYm5_0),.din(w_dff_A_e7giKlnW0_0),.clk(gclk));
	jdff dff_A_PEIkaqYm5_0(.dout(w_dff_A_458vZjmV1_0),.din(w_dff_A_PEIkaqYm5_0),.clk(gclk));
	jdff dff_A_458vZjmV1_0(.dout(G6),.din(w_dff_A_458vZjmV1_0),.clk(gclk));
	jdff dff_A_eO18hD5z1_2(.dout(w_dff_A_3kPMnGYT1_0),.din(w_dff_A_eO18hD5z1_2),.clk(gclk));
	jdff dff_A_3kPMnGYT1_0(.dout(w_dff_A_JdYBryj15_0),.din(w_dff_A_3kPMnGYT1_0),.clk(gclk));
	jdff dff_A_JdYBryj15_0(.dout(w_dff_A_3lUjyb5F3_0),.din(w_dff_A_JdYBryj15_0),.clk(gclk));
	jdff dff_A_3lUjyb5F3_0(.dout(w_dff_A_wO15XS5a6_0),.din(w_dff_A_3lUjyb5F3_0),.clk(gclk));
	jdff dff_A_wO15XS5a6_0(.dout(w_dff_A_H9S3Zmtk7_0),.din(w_dff_A_wO15XS5a6_0),.clk(gclk));
	jdff dff_A_H9S3Zmtk7_0(.dout(w_dff_A_YgWnHk5c8_0),.din(w_dff_A_H9S3Zmtk7_0),.clk(gclk));
	jdff dff_A_YgWnHk5c8_0(.dout(w_dff_A_JsurAuWB6_0),.din(w_dff_A_YgWnHk5c8_0),.clk(gclk));
	jdff dff_A_JsurAuWB6_0(.dout(G9),.din(w_dff_A_JsurAuWB6_0),.clk(gclk));
	jdff dff_A_hoBHkjw44_2(.dout(w_dff_A_wdBsn0Ip9_0),.din(w_dff_A_hoBHkjw44_2),.clk(gclk));
	jdff dff_A_wdBsn0Ip9_0(.dout(w_dff_A_F9Cz8fkK3_0),.din(w_dff_A_wdBsn0Ip9_0),.clk(gclk));
	jdff dff_A_F9Cz8fkK3_0(.dout(w_dff_A_NM8ne8bv0_0),.din(w_dff_A_F9Cz8fkK3_0),.clk(gclk));
	jdff dff_A_NM8ne8bv0_0(.dout(w_dff_A_zFFE9N1h1_0),.din(w_dff_A_NM8ne8bv0_0),.clk(gclk));
	jdff dff_A_zFFE9N1h1_0(.dout(w_dff_A_4TIpI5nb8_0),.din(w_dff_A_zFFE9N1h1_0),.clk(gclk));
	jdff dff_A_4TIpI5nb8_0(.dout(w_dff_A_ftOWdplm3_0),.din(w_dff_A_4TIpI5nb8_0),.clk(gclk));
	jdff dff_A_ftOWdplm3_0(.dout(w_dff_A_nnWLkqy59_0),.din(w_dff_A_ftOWdplm3_0),.clk(gclk));
	jdff dff_A_nnWLkqy59_0(.dout(G12),.din(w_dff_A_nnWLkqy59_0),.clk(gclk));
	jdff dff_A_lNq4Cyh81_2(.dout(w_dff_A_8qfaC76O3_0),.din(w_dff_A_lNq4Cyh81_2),.clk(gclk));
	jdff dff_A_8qfaC76O3_0(.dout(w_dff_A_0WwlKeNZ8_0),.din(w_dff_A_8qfaC76O3_0),.clk(gclk));
	jdff dff_A_0WwlKeNZ8_0(.dout(w_dff_A_gAiXq8Ze1_0),.din(w_dff_A_0WwlKeNZ8_0),.clk(gclk));
	jdff dff_A_gAiXq8Ze1_0(.dout(w_dff_A_HoAwywnQ6_0),.din(w_dff_A_gAiXq8Ze1_0),.clk(gclk));
	jdff dff_A_HoAwywnQ6_0(.dout(w_dff_A_yFi0bW4o3_0),.din(w_dff_A_HoAwywnQ6_0),.clk(gclk));
	jdff dff_A_yFi0bW4o3_0(.dout(w_dff_A_KuEGRZOL1_0),.din(w_dff_A_yFi0bW4o3_0),.clk(gclk));
	jdff dff_A_KuEGRZOL1_0(.dout(w_dff_A_mAnqE5Dy1_0),.din(w_dff_A_KuEGRZOL1_0),.clk(gclk));
	jdff dff_A_mAnqE5Dy1_0(.dout(G30),.din(w_dff_A_mAnqE5Dy1_0),.clk(gclk));
	jdff dff_A_hj6neaL13_2(.dout(w_dff_A_BBVzFjDh6_0),.din(w_dff_A_hj6neaL13_2),.clk(gclk));
	jdff dff_A_BBVzFjDh6_0(.dout(w_dff_A_fH3JpKnj3_0),.din(w_dff_A_BBVzFjDh6_0),.clk(gclk));
	jdff dff_A_fH3JpKnj3_0(.dout(w_dff_A_p7xXiNuJ6_0),.din(w_dff_A_fH3JpKnj3_0),.clk(gclk));
	jdff dff_A_p7xXiNuJ6_0(.dout(w_dff_A_pLoShYLs1_0),.din(w_dff_A_p7xXiNuJ6_0),.clk(gclk));
	jdff dff_A_pLoShYLs1_0(.dout(w_dff_A_KJEoonuq8_0),.din(w_dff_A_pLoShYLs1_0),.clk(gclk));
	jdff dff_A_KJEoonuq8_0(.dout(w_dff_A_zxFSqyT41_0),.din(w_dff_A_KJEoonuq8_0),.clk(gclk));
	jdff dff_A_zxFSqyT41_0(.dout(w_dff_A_QtOGY8Mz7_0),.din(w_dff_A_zxFSqyT41_0),.clk(gclk));
	jdff dff_A_QtOGY8Mz7_0(.dout(G45),.din(w_dff_A_QtOGY8Mz7_0),.clk(gclk));
	jdff dff_A_MQKByHQh7_2(.dout(w_dff_A_3N4nzonT5_0),.din(w_dff_A_MQKByHQh7_2),.clk(gclk));
	jdff dff_A_3N4nzonT5_0(.dout(w_dff_A_ZOX2T6Mi3_0),.din(w_dff_A_3N4nzonT5_0),.clk(gclk));
	jdff dff_A_ZOX2T6Mi3_0(.dout(w_dff_A_izmajK9o8_0),.din(w_dff_A_ZOX2T6Mi3_0),.clk(gclk));
	jdff dff_A_izmajK9o8_0(.dout(w_dff_A_4CbT9viI2_0),.din(w_dff_A_izmajK9o8_0),.clk(gclk));
	jdff dff_A_4CbT9viI2_0(.dout(w_dff_A_6rRrLFjN5_0),.din(w_dff_A_4CbT9viI2_0),.clk(gclk));
	jdff dff_A_6rRrLFjN5_0(.dout(w_dff_A_Oan4keWR6_0),.din(w_dff_A_6rRrLFjN5_0),.clk(gclk));
	jdff dff_A_Oan4keWR6_0(.dout(w_dff_A_QCf0hqno0_0),.din(w_dff_A_Oan4keWR6_0),.clk(gclk));
	jdff dff_A_QCf0hqno0_0(.dout(G48),.din(w_dff_A_QCf0hqno0_0),.clk(gclk));
	jdff dff_A_v8v81gOu0_2(.dout(w_dff_A_uVsynPQB4_0),.din(w_dff_A_v8v81gOu0_2),.clk(gclk));
	jdff dff_A_uVsynPQB4_0(.dout(w_dff_A_pQx3iepF6_0),.din(w_dff_A_uVsynPQB4_0),.clk(gclk));
	jdff dff_A_pQx3iepF6_0(.dout(w_dff_A_dS6OrFo16_0),.din(w_dff_A_pQx3iepF6_0),.clk(gclk));
	jdff dff_A_dS6OrFo16_0(.dout(w_dff_A_Gbngxas66_0),.din(w_dff_A_dS6OrFo16_0),.clk(gclk));
	jdff dff_A_Gbngxas66_0(.dout(w_dff_A_MDJKZ6ik6_0),.din(w_dff_A_Gbngxas66_0),.clk(gclk));
	jdff dff_A_MDJKZ6ik6_0(.dout(w_dff_A_Kf98beXv8_0),.din(w_dff_A_MDJKZ6ik6_0),.clk(gclk));
	jdff dff_A_Kf98beXv8_0(.dout(w_dff_A_VU2Bv5dh1_0),.din(w_dff_A_Kf98beXv8_0),.clk(gclk));
	jdff dff_A_VU2Bv5dh1_0(.dout(G15),.din(w_dff_A_VU2Bv5dh1_0),.clk(gclk));
	jdff dff_A_6MMl4RMX9_2(.dout(w_dff_A_slnGxkdR8_0),.din(w_dff_A_6MMl4RMX9_2),.clk(gclk));
	jdff dff_A_slnGxkdR8_0(.dout(w_dff_A_9Y4jb4jo2_0),.din(w_dff_A_slnGxkdR8_0),.clk(gclk));
	jdff dff_A_9Y4jb4jo2_0(.dout(w_dff_A_PYGZro3Y9_0),.din(w_dff_A_9Y4jb4jo2_0),.clk(gclk));
	jdff dff_A_PYGZro3Y9_0(.dout(w_dff_A_nGIw7NVE4_0),.din(w_dff_A_PYGZro3Y9_0),.clk(gclk));
	jdff dff_A_nGIw7NVE4_0(.dout(w_dff_A_SHB0QNEh5_0),.din(w_dff_A_nGIw7NVE4_0),.clk(gclk));
	jdff dff_A_SHB0QNEh5_0(.dout(w_dff_A_vJZ8BV4y7_0),.din(w_dff_A_SHB0QNEh5_0),.clk(gclk));
	jdff dff_A_vJZ8BV4y7_0(.dout(w_dff_A_7ppUnfnZ6_0),.din(w_dff_A_vJZ8BV4y7_0),.clk(gclk));
	jdff dff_A_7ppUnfnZ6_0(.dout(G18),.din(w_dff_A_7ppUnfnZ6_0),.clk(gclk));
	jdff dff_A_I5xO0wr80_2(.dout(w_dff_A_fiHvYHbj9_0),.din(w_dff_A_I5xO0wr80_2),.clk(gclk));
	jdff dff_A_fiHvYHbj9_0(.dout(w_dff_A_E0yHZl4K6_0),.din(w_dff_A_fiHvYHbj9_0),.clk(gclk));
	jdff dff_A_E0yHZl4K6_0(.dout(w_dff_A_QgpErsWx5_0),.din(w_dff_A_E0yHZl4K6_0),.clk(gclk));
	jdff dff_A_QgpErsWx5_0(.dout(w_dff_A_WojpYgxi1_0),.din(w_dff_A_QgpErsWx5_0),.clk(gclk));
	jdff dff_A_WojpYgxi1_0(.dout(w_dff_A_Ka24iUkt3_0),.din(w_dff_A_WojpYgxi1_0),.clk(gclk));
	jdff dff_A_Ka24iUkt3_0(.dout(w_dff_A_NQhAoMm50_0),.din(w_dff_A_Ka24iUkt3_0),.clk(gclk));
	jdff dff_A_NQhAoMm50_0(.dout(w_dff_A_otYwzOBX0_0),.din(w_dff_A_NQhAoMm50_0),.clk(gclk));
	jdff dff_A_otYwzOBX0_0(.dout(G21),.din(w_dff_A_otYwzOBX0_0),.clk(gclk));
	jdff dff_A_7zomEpPc3_2(.dout(w_dff_A_qBVdfWZF1_0),.din(w_dff_A_7zomEpPc3_2),.clk(gclk));
	jdff dff_A_qBVdfWZF1_0(.dout(w_dff_A_PYZ2zXnr3_0),.din(w_dff_A_qBVdfWZF1_0),.clk(gclk));
	jdff dff_A_PYZ2zXnr3_0(.dout(w_dff_A_O9PQebAI8_0),.din(w_dff_A_PYZ2zXnr3_0),.clk(gclk));
	jdff dff_A_O9PQebAI8_0(.dout(w_dff_A_PI1MS8eu2_0),.din(w_dff_A_O9PQebAI8_0),.clk(gclk));
	jdff dff_A_PI1MS8eu2_0(.dout(w_dff_A_ar1DRlSm3_0),.din(w_dff_A_PI1MS8eu2_0),.clk(gclk));
	jdff dff_A_ar1DRlSm3_0(.dout(w_dff_A_5Yzf6ebd2_0),.din(w_dff_A_ar1DRlSm3_0),.clk(gclk));
	jdff dff_A_5Yzf6ebd2_0(.dout(G24),.din(w_dff_A_5Yzf6ebd2_0),.clk(gclk));
	jdff dff_A_4wG7pdcN0_2(.dout(w_dff_A_53SmPLCM5_0),.din(w_dff_A_4wG7pdcN0_2),.clk(gclk));
	jdff dff_A_53SmPLCM5_0(.dout(w_dff_A_HdiAkpbs7_0),.din(w_dff_A_53SmPLCM5_0),.clk(gclk));
	jdff dff_A_HdiAkpbs7_0(.dout(w_dff_A_TXwxBMh17_0),.din(w_dff_A_HdiAkpbs7_0),.clk(gclk));
	jdff dff_A_TXwxBMh17_0(.dout(w_dff_A_DB8V6ybq5_0),.din(w_dff_A_TXwxBMh17_0),.clk(gclk));
	jdff dff_A_DB8V6ybq5_0(.dout(w_dff_A_p6fKBKuC0_0),.din(w_dff_A_DB8V6ybq5_0),.clk(gclk));
	jdff dff_A_p6fKBKuC0_0(.dout(w_dff_A_KyKqygUl2_0),.din(w_dff_A_p6fKBKuC0_0),.clk(gclk));
	jdff dff_A_KyKqygUl2_0(.dout(w_dff_A_5nmiEcia7_0),.din(w_dff_A_KyKqygUl2_0),.clk(gclk));
	jdff dff_A_5nmiEcia7_0(.dout(G27),.din(w_dff_A_5nmiEcia7_0),.clk(gclk));
	jdff dff_A_FHZ9zkzZ5_2(.dout(w_dff_A_68mMAGHY6_0),.din(w_dff_A_FHZ9zkzZ5_2),.clk(gclk));
	jdff dff_A_68mMAGHY6_0(.dout(w_dff_A_ynUaYUQm2_0),.din(w_dff_A_68mMAGHY6_0),.clk(gclk));
	jdff dff_A_ynUaYUQm2_0(.dout(w_dff_A_2SHu7Z7z8_0),.din(w_dff_A_ynUaYUQm2_0),.clk(gclk));
	jdff dff_A_2SHu7Z7z8_0(.dout(w_dff_A_JDMIB01L9_0),.din(w_dff_A_2SHu7Z7z8_0),.clk(gclk));
	jdff dff_A_JDMIB01L9_0(.dout(w_dff_A_wJq8yI2Z8_0),.din(w_dff_A_JDMIB01L9_0),.clk(gclk));
	jdff dff_A_wJq8yI2Z8_0(.dout(w_dff_A_H1H5ZwiN7_0),.din(w_dff_A_wJq8yI2Z8_0),.clk(gclk));
	jdff dff_A_H1H5ZwiN7_0(.dout(w_dff_A_SAZMZT7I1_0),.din(w_dff_A_H1H5ZwiN7_0),.clk(gclk));
	jdff dff_A_SAZMZT7I1_0(.dout(G33),.din(w_dff_A_SAZMZT7I1_0),.clk(gclk));
	jdff dff_A_owRIK1eH7_2(.dout(w_dff_A_kYODZ5Ae6_0),.din(w_dff_A_owRIK1eH7_2),.clk(gclk));
	jdff dff_A_kYODZ5Ae6_0(.dout(w_dff_A_UC56cU1K0_0),.din(w_dff_A_kYODZ5Ae6_0),.clk(gclk));
	jdff dff_A_UC56cU1K0_0(.dout(w_dff_A_GyP6ThQA8_0),.din(w_dff_A_UC56cU1K0_0),.clk(gclk));
	jdff dff_A_GyP6ThQA8_0(.dout(w_dff_A_p9cqZigD0_0),.din(w_dff_A_GyP6ThQA8_0),.clk(gclk));
	jdff dff_A_p9cqZigD0_0(.dout(w_dff_A_74Ag3JT38_0),.din(w_dff_A_p9cqZigD0_0),.clk(gclk));
	jdff dff_A_74Ag3JT38_0(.dout(w_dff_A_dvQRztiP1_0),.din(w_dff_A_74Ag3JT38_0),.clk(gclk));
	jdff dff_A_dvQRztiP1_0(.dout(w_dff_A_KiD3spGf3_0),.din(w_dff_A_dvQRztiP1_0),.clk(gclk));
	jdff dff_A_KiD3spGf3_0(.dout(G36),.din(w_dff_A_KiD3spGf3_0),.clk(gclk));
	jdff dff_A_0SkdKhgQ2_2(.dout(w_dff_A_YigTklAD3_0),.din(w_dff_A_0SkdKhgQ2_2),.clk(gclk));
	jdff dff_A_YigTklAD3_0(.dout(w_dff_A_qPs5LhP03_0),.din(w_dff_A_YigTklAD3_0),.clk(gclk));
	jdff dff_A_qPs5LhP03_0(.dout(w_dff_A_g3y226p61_0),.din(w_dff_A_qPs5LhP03_0),.clk(gclk));
	jdff dff_A_g3y226p61_0(.dout(w_dff_A_liw3VfIV6_0),.din(w_dff_A_g3y226p61_0),.clk(gclk));
	jdff dff_A_liw3VfIV6_0(.dout(w_dff_A_lO4mnAmy2_0),.din(w_dff_A_liw3VfIV6_0),.clk(gclk));
	jdff dff_A_lO4mnAmy2_0(.dout(w_dff_A_3VkCP3fv2_0),.din(w_dff_A_lO4mnAmy2_0),.clk(gclk));
	jdff dff_A_3VkCP3fv2_0(.dout(w_dff_A_svJDJUqM9_0),.din(w_dff_A_3VkCP3fv2_0),.clk(gclk));
	jdff dff_A_svJDJUqM9_0(.dout(G39),.din(w_dff_A_svJDJUqM9_0),.clk(gclk));
	jdff dff_A_4ZmVwtxX9_2(.dout(w_dff_A_DKLUyJIk1_0),.din(w_dff_A_4ZmVwtxX9_2),.clk(gclk));
	jdff dff_A_DKLUyJIk1_0(.dout(w_dff_A_e5097vWo3_0),.din(w_dff_A_DKLUyJIk1_0),.clk(gclk));
	jdff dff_A_e5097vWo3_0(.dout(w_dff_A_krmH0raQ6_0),.din(w_dff_A_e5097vWo3_0),.clk(gclk));
	jdff dff_A_krmH0raQ6_0(.dout(w_dff_A_nBDoDcUE8_0),.din(w_dff_A_krmH0raQ6_0),.clk(gclk));
	jdff dff_A_nBDoDcUE8_0(.dout(w_dff_A_bC1GMlB05_0),.din(w_dff_A_nBDoDcUE8_0),.clk(gclk));
	jdff dff_A_bC1GMlB05_0(.dout(w_dff_A_QALXnU1B0_0),.din(w_dff_A_bC1GMlB05_0),.clk(gclk));
	jdff dff_A_QALXnU1B0_0(.dout(w_dff_A_gGXzisCY3_0),.din(w_dff_A_QALXnU1B0_0),.clk(gclk));
	jdff dff_A_gGXzisCY3_0(.dout(G42),.din(w_dff_A_gGXzisCY3_0),.clk(gclk));
	jdff dff_A_FMGvs0En8_2(.dout(G75),.din(w_dff_A_FMGvs0En8_2),.clk(gclk));
	jdff dff_A_g202tuwu0_2(.dout(w_dff_A_eSfTIwb37_0),.din(w_dff_A_g202tuwu0_2),.clk(gclk));
	jdff dff_A_eSfTIwb37_0(.dout(G69),.din(w_dff_A_eSfTIwb37_0),.clk(gclk));
	jdff dff_A_VvBkGpwi0_2(.dout(w_dff_A_TiRLqdJ76_0),.din(w_dff_A_VvBkGpwi0_2),.clk(gclk));
	jdff dff_A_TiRLqdJ76_0(.dout(G72),.din(w_dff_A_TiRLqdJ76_0),.clk(gclk));
	jdff dff_A_IidXqrXl3_2(.dout(G57),.din(w_dff_A_IidXqrXl3_2),.clk(gclk));
endmodule

