/*

c1908:
	jxor: 75
	jspl: 95
	jspl3: 88
	jnot: 40
	jcb: 82
	jdff: 781
	jand: 122

Summary:
	jxor: 75
	jspl: 95
	jspl3: 88
	jnot: 40
	jcb: 82
	jdff: 781
	jand: 122
*/

module c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n170;
	wire n171;
	wire n172;
	wire n174;
	wire n175;
	wire n176;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n193;
	wire n194;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n203;
	wire n205;
	wire n206;
	wire n207;
	wire n209;
	wire n210;
	wire n211;
	wire n213;
	wire n214;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n222;
	wire n224;
	wire n225;
	wire n226;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n275;
	wire n276;
	wire n277;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n353;
	wire n354;
	wire n355;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n374;
	wire n375;
	wire n376;
	wire [2:0] w_G101_0;
	wire [2:0] w_G104_0;
	wire [2:0] w_G107_0;
	wire [2:0] w_G110_0;
	wire [2:0] w_G113_0;
	wire [2:0] w_G116_0;
	wire [2:0] w_G119_0;
	wire [2:0] w_G122_0;
	wire [1:0] w_G122_1;
	wire [2:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [2:0] w_G131_0;
	wire [2:0] w_G134_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G140_0;
	wire [2:0] w_G143_0;
	wire [2:0] w_G146_0;
	wire [2:0] w_G210_0;
	wire [1:0] w_G214_0;
	wire [2:0] w_G217_0;
	wire [1:0] w_G221_0;
	wire [1:0] w_G224_0;
	wire [1:0] w_G227_0;
	wire [2:0] w_G234_0;
	wire [1:0] w_G234_1;
	wire [1:0] w_G237_0;
	wire [1:0] w_G469_0;
	wire [2:0] w_G472_0;
	wire [2:0] w_G475_0;
	wire [1:0] w_G478_0;
	wire [1:0] w_G898_0;
	wire [1:0] w_G900_0;
	wire [2:0] w_G902_0;
	wire [2:0] w_G902_1;
	wire [2:0] w_G902_2;
	wire [2:0] w_G902_3;
	wire [2:0] w_G902_4;
	wire [2:0] w_G952_0;
	wire [2:0] w_G953_0;
	wire [2:0] w_G953_1;
	wire [2:0] w_G953_2;
	wire [1:0] w_G953_3;
	wire [2:0] w_n59_0;
	wire [2:0] w_n59_1;
	wire [1:0] w_n59_2;
	wire [2:0] w_n61_0;
	wire [2:0] w_n61_1;
	wire [2:0] w_n61_2;
	wire [2:0] w_n61_3;
	wire [1:0] w_n65_0;
	wire [1:0] w_n66_0;
	wire [1:0] w_n67_0;
	wire [1:0] w_n71_0;
	wire [1:0] w_n72_0;
	wire [1:0] w_n74_0;
	wire [1:0] w_n75_0;
	wire [2:0] w_n77_0;
	wire [1:0] w_n77_1;
	wire [1:0] w_n78_0;
	wire [1:0] w_n79_0;
	wire [2:0] w_n82_0;
	wire [1:0] w_n84_0;
	wire [2:0] w_n85_0;
	wire [1:0] w_n90_0;
	wire [1:0] w_n91_0;
	wire [2:0] w_n92_0;
	wire [1:0] w_n92_1;
	wire [2:0] w_n93_0;
	wire [1:0] w_n95_0;
	wire [1:0] w_n96_0;
	wire [1:0] w_n98_0;
	wire [2:0] w_n101_0;
	wire [1:0] w_n105_0;
	wire [2:0] w_n108_0;
	wire [2:0] w_n109_0;
	wire [2:0] w_n111_0;
	wire [1:0] w_n119_0;
	wire [2:0] w_n121_0;
	wire [2:0] w_n122_0;
	wire [2:0] w_n123_0;
	wire [1:0] w_n123_1;
	wire [1:0] w_n125_0;
	wire [2:0] w_n128_0;
	wire [1:0] w_n129_0;
	wire [1:0] w_n131_0;
	wire [2:0] w_n134_0;
	wire [2:0] w_n134_1;
	wire [2:0] w_n141_0;
	wire [2:0] w_n143_0;
	wire [2:0] w_n143_1;
	wire [2:0] w_n144_0;
	wire [1:0] w_n144_1;
	wire [2:0] w_n153_0;
	wire [1:0] w_n154_0;
	wire [2:0] w_n155_0;
	wire [2:0] w_n155_1;
	wire [2:0] w_n156_0;
	wire [1:0] w_n156_1;
	wire [1:0] w_n157_0;
	wire [1:0] w_n158_0;
	wire [2:0] w_n159_0;
	wire [2:0] w_n162_0;
	wire [1:0] w_n162_1;
	wire [2:0] w_n163_0;
	wire [1:0] w_n163_1;
	wire [1:0] w_n164_0;
	wire [2:0] w_n165_0;
	wire [1:0] w_n166_0;
	wire [2:0] w_n167_0;
	wire [1:0] w_n168_0;
	wire [1:0] w_n170_0;
	wire [2:0] w_n171_0;
	wire [1:0] w_n172_0;
	wire [2:0] w_n174_0;
	wire [1:0] w_n174_1;
	wire [1:0] w_n175_0;
	wire [1:0] w_n176_0;
	wire [2:0] w_n178_0;
	wire [1:0] w_n179_0;
	wire [1:0] w_n181_0;
	wire [2:0] w_n184_0;
	wire [2:0] w_n184_1;
	wire [2:0] w_n185_0;
	wire [1:0] w_n186_0;
	wire [1:0] w_n188_0;
	wire [1:0] w_n191_0;
	wire [2:0] w_n193_0;
	wire [1:0] w_n194_0;
	wire [1:0] w_n196_0;
	wire [1:0] w_n197_0;
	wire [2:0] w_n198_0;
	wire [2:0] w_n198_1;
	wire [2:0] w_n199_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n201_0;
	wire [1:0] w_n203_0;
	wire [2:0] w_n205_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n211_0;
	wire [1:0] w_n213_0;
	wire [1:0] w_n214_0;
	wire [1:0] w_n216_0;
	wire [2:0] w_n217_0;
	wire [2:0] w_n218_0;
	wire [1:0] w_n218_1;
	wire [1:0] w_n219_0;
	wire [2:0] w_n220_0;
	wire [2:0] w_n222_0;
	wire [1:0] w_n226_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n236_0;
	wire [2:0] w_n244_0;
	wire [2:0] w_n244_1;
	wire [2:0] w_n244_2;
	wire [2:0] w_n247_0;
	wire [1:0] w_n248_0;
	wire [2:0] w_n253_0;
	wire [1:0] w_n253_1;
	wire [1:0] w_n254_0;
	wire [1:0] w_n259_0;
	wire [2:0] w_n269_0;
	wire [2:0] w_n269_1;
	wire [1:0] w_n269_2;
	wire [1:0] w_n279_0;
	wire [2:0] w_n285_0;
	wire [1:0] w_n285_1;
	wire [1:0] w_n286_0;
	wire [1:0] w_n287_0;
	wire [1:0] w_n289_0;
	wire [1:0] w_n296_0;
	wire [1:0] w_n297_0;
	wire [1:0] w_n298_0;
	wire [1:0] w_n300_0;
	wire [1:0] w_n304_0;
	wire [1:0] w_n311_0;
	wire [1:0] w_n313_0;
	wire [2:0] w_n315_0;
	wire [1:0] w_n316_0;
	wire [1:0] w_n321_0;
	wire [1:0] w_n326_0;
	wire [1:0] w_n337_0;
	wire [1:0] w_n338_0;
	wire [1:0] w_n344_0;
	wire w_dff_B_Dk4nmQs10_0;
	wire w_dff_B_OiV1sQ5l7_0;
	wire w_dff_B_YKpfZl1u5_0;
	wire w_dff_B_8Jg4Dzxz2_0;
	wire w_dff_B_ylgErEEf9_0;
	wire w_dff_B_6gIYyRZb2_1;
	wire w_dff_B_MvrFUeGV0_1;
	wire w_dff_B_NjbvnhGJ3_0;
	wire w_dff_B_em63zvdk5_1;
	wire w_dff_B_UY0HwHku7_1;
	wire w_dff_B_U3De3fb42_1;
	wire w_dff_B_kX2MOGrI8_1;
	wire w_dff_B_kXXFVEmg9_1;
	wire w_dff_B_QjdjnfdV3_1;
	wire w_dff_B_T2VrmKJn9_1;
	wire w_dff_B_Itw8uBOB2_1;
	wire w_dff_B_gAJeyiaM8_0;
	wire w_dff_B_PcbmW6ZI7_0;
	wire w_dff_B_UK4GJsiV3_0;
	wire w_dff_B_p8xDgMib8_0;
	wire w_dff_B_rd6nBQVs2_0;
	wire w_dff_B_n697LSWx5_0;
	wire w_dff_B_EB4LNcGZ2_0;
	wire w_dff_B_ts2CxtsM2_0;
	wire w_dff_B_BoWr6wRo6_0;
	wire w_dff_B_BWu6umMX5_0;
	wire w_dff_B_zyjvtZ0X8_0;
	wire w_dff_A_4JaeotOm3_2;
	wire w_dff_A_fvTFRsyf6_1;
	wire w_dff_B_ff8Q1GrI0_1;
	wire w_dff_B_03te53yw1_1;
	wire w_dff_B_GoxgVuQm1_1;
	wire w_dff_B_GxLZSbNy4_1;
	wire w_dff_B_DaoqrbUh7_1;
	wire w_dff_B_Kk1z713U8_1;
	wire w_dff_B_c92ERZF98_1;
	wire w_dff_B_9PlWo8jR6_1;
	wire w_dff_B_Y0mwXCeU4_1;
	wire w_dff_B_XBJ5yhqs2_1;
	wire w_dff_B_gxavRIm69_1;
	wire w_dff_B_c0jutqYs8_1;
	wire w_dff_B_p4MO3Bt46_1;
	wire w_dff_B_WUCWDsxf3_0;
	wire w_dff_B_uSENDypd6_0;
	wire w_dff_B_2RNIIohY6_0;
	wire w_dff_B_cVyJoijz4_0;
	wire w_dff_B_kQZEMinE7_0;
	wire w_dff_B_g2FPmPs22_0;
	wire w_dff_B_ou9mg8HE5_0;
	wire w_dff_B_rG9sL0fK0_0;
	wire w_dff_B_7xA612sE3_0;
	wire w_dff_B_WyNOZNnZ1_0;
	wire w_dff_B_c08gOoFP3_0;
	wire w_dff_B_BtoisHfb7_0;
	wire w_dff_B_zrMQXsVj2_0;
	wire w_dff_B_2xASnDVr2_0;
	wire w_dff_A_EcL0WOZG5_1;
	wire w_dff_A_sEPJfhib7_1;
	wire w_dff_A_rlZF7qFx8_1;
	wire w_dff_A_wxdIY6kZ7_1;
	wire w_dff_A_kUl6HOYn4_1;
	wire w_dff_A_PYfon3DB3_1;
	wire w_dff_A_ibeh9fBD5_1;
	wire w_dff_A_eFB6ihZF5_1;
	wire w_dff_A_UHepSLeq9_1;
	wire w_dff_A_Kfqyqo8a0_1;
	wire w_dff_A_fIkK8fy79_1;
	wire w_dff_B_8fBUTVCq5_1;
	wire w_dff_B_W3BUisI20_1;
	wire w_dff_B_gyGRWXvE0_1;
	wire w_dff_B_dCMRLTmz6_1;
	wire w_dff_B_yKxbtZyX9_1;
	wire w_dff_B_slOzX6yU0_1;
	wire w_dff_B_6KHY34Mi1_1;
	wire w_dff_B_n5iJZUgU0_1;
	wire w_dff_B_wWW4dRvM1_1;
	wire w_dff_B_R9hpgwhr0_1;
	wire w_dff_B_HZMw9LuV2_1;
	wire w_dff_B_ROQ7uGzp9_1;
	wire w_dff_B_PwqUDIoi2_1;
	wire w_dff_B_npYXXQxt5_1;
	wire w_dff_B_OaMo6QT61_1;
	wire w_dff_B_F3DvtgB63_0;
	wire w_dff_B_jnyU4Ckc9_0;
	wire w_dff_B_YlXgNFay8_0;
	wire w_dff_B_qvbMmWX09_0;
	wire w_dff_B_ooPDCouk1_0;
	wire w_dff_B_zvMao9e51_0;
	wire w_dff_B_0aQxesjY8_0;
	wire w_dff_B_agmjxW9b8_0;
	wire w_dff_B_UanMI6PQ5_0;
	wire w_dff_B_0wIwARpR3_0;
	wire w_dff_B_1SozOU5l1_0;
	wire w_dff_B_bhURgl5o7_0;
	wire w_dff_B_JpMHvu8u7_0;
	wire w_dff_B_ZOgbkHDb3_0;
	wire w_dff_A_iWmSOYTH3_1;
	wire w_dff_A_GIDscngr8_1;
	wire w_dff_A_KsALonDl2_1;
	wire w_dff_A_c4dqkhV37_1;
	wire w_dff_A_MBSH6idT0_1;
	wire w_dff_A_UMjil9E39_1;
	wire w_dff_A_tPbWrMP06_1;
	wire w_dff_A_sWuEpO6F0_1;
	wire w_dff_A_ikJaiGE46_1;
	wire w_dff_A_sW092USv9_1;
	wire w_dff_A_7OdfY3Yh9_1;
	wire w_dff_A_fSftLx0k0_1;
	wire w_dff_A_wQFJnKsT9_2;
	wire w_dff_B_12tuOhTj8_0;
	wire w_dff_B_SCNXTHcA9_0;
	wire w_dff_B_34pwF9lI7_0;
	wire w_dff_B_odoxzutY0_0;
	wire w_dff_B_uBEPWvoz9_0;
	wire w_dff_B_e0bCpcWF3_0;
	wire w_dff_B_FzxnJLA86_0;
	wire w_dff_B_R17FHUEx6_0;
	wire w_dff_B_iM9wOI6B4_0;
	wire w_dff_B_FES3Toxd5_0;
	wire w_dff_B_Pcrt2pkk2_0;
	wire w_dff_B_6brJrFNK4_0;
	wire w_dff_B_kOBba82f2_0;
	wire w_dff_B_y0vioXrN2_0;
	wire w_dff_B_Y0kMxlKp3_0;
	wire w_dff_B_MS016RQz8_0;
	wire w_dff_B_lyofbDAS1_0;
	wire w_dff_B_h03GltJP2_0;
	wire w_dff_B_fqBX134S8_0;
	wire w_dff_B_Ad6I2Q6H2_0;
	wire w_dff_B_iIlpi7Af4_0;
	wire w_dff_B_yiyIbJqJ2_0;
	wire w_dff_B_iX483IMn3_0;
	wire w_dff_B_7lY6yjeu8_0;
	wire w_dff_B_0KQt4l9f1_0;
	wire w_dff_B_vMa7JgJg5_0;
	wire w_dff_B_cYj50Ohn8_0;
	wire w_dff_B_GAYwLA6H8_0;
	wire w_dff_A_mOAYSE0e8_1;
	wire w_dff_A_WePsK7ok3_1;
	wire w_dff_B_lDqoR1E15_2;
	wire w_dff_B_hTSCfNiX7_2;
	wire w_dff_B_juXlPDi56_2;
	wire w_dff_B_a5CkEPVo4_0;
	wire w_dff_B_aSJsIa6r1_2;
	wire w_dff_B_Sk0MnWd06_2;
	wire w_dff_A_lCyFUNZz8_1;
	wire w_dff_A_iwoknT9B4_2;
	wire w_dff_B_nz6nYAlU1_0;
	wire w_dff_B_V7dRqMkb6_0;
	wire w_dff_B_TngN26zw1_0;
	wire w_dff_B_xZCUJF3B7_0;
	wire w_dff_B_8sLvhIEi7_0;
	wire w_dff_B_fxz3TBLs6_0;
	wire w_dff_B_nutD5hqc5_0;
	wire w_dff_B_spzrTbcT1_0;
	wire w_dff_B_7wcgNGc58_0;
	wire w_dff_B_qJewMhEt2_0;
	wire w_dff_B_wO5oH2yq7_0;
	wire w_dff_B_I03464Z71_0;
	wire w_dff_B_c9pJwPQJ5_0;
	wire w_dff_B_y2a4YXIC7_0;
	wire w_dff_B_LeQxV6TU7_0;
	wire w_dff_B_eAkV4tXr9_0;
	wire w_dff_B_xErKtZCo4_0;
	wire w_dff_B_fLaqRo0Y6_0;
	wire w_dff_B_iNUBiQYV9_0;
	wire w_dff_B_UVCa8OEN7_0;
	wire w_dff_B_XjSC0c9B5_0;
	wire w_dff_B_WBmJI8q53_0;
	wire w_dff_B_moIPe1Fm6_0;
	wire w_dff_B_pCFVqoTP1_0;
	wire w_dff_B_w1YOFz4z6_0;
	wire w_dff_B_ETtamJp77_0;
	wire w_dff_A_rAEbi5pg6_2;
	wire w_dff_A_mpX9JVRz0_2;
	wire w_dff_A_1JSmv3Xz2_2;
	wire w_dff_A_w1L5U8hZ8_2;
	wire w_dff_A_so2v8p0p3_2;
	wire w_dff_A_jlSTJxON8_2;
	wire w_dff_A_EhNoLLJc3_2;
	wire w_dff_A_tAnzTqMF4_2;
	wire w_dff_A_LBotY2eC5_2;
	wire w_dff_A_whoP7SOZ7_2;
	wire w_dff_A_m6tq2qpa7_2;
	wire w_dff_B_YHUknnpY0_1;
	wire w_dff_B_HOwBZZzy8_1;
	wire w_dff_B_aiRoMdoG5_1;
	wire w_dff_B_ezAnpGU13_1;
	wire w_dff_B_iIqvjNOa3_0;
	wire w_dff_B_pJ5gaPhu0_0;
	wire w_dff_B_n6HfhzeT0_0;
	wire w_dff_B_d4MGz1xW8_1;
	wire w_dff_B_mYZ6SdKZ6_0;
	wire w_dff_A_5eRgs1NA1_0;
	wire w_dff_A_kzyFlC3Z5_0;
	wire w_dff_A_QbYjEiid8_1;
	wire w_dff_B_p6TVTbM01_0;
	wire w_dff_A_xnd6brWN0_1;
	wire w_dff_B_d0hNRf772_3;
	wire w_dff_B_qOkiHl6x6_3;
	wire w_dff_B_BVBFn80e3_3;
	wire w_dff_A_Fk3ksdOx2_0;
	wire w_dff_A_C1rSbdtx0_0;
	wire w_dff_A_E873VoV34_2;
	wire w_dff_A_FweZJOWU1_0;
	wire w_dff_A_seyGBe7W1_0;
	wire w_dff_A_aYCmzNej5_0;
	wire w_dff_A_xqMIXTHk3_0;
	wire w_dff_A_pDYjh9H73_1;
	wire w_dff_A_NrYsuE4t4_1;
	wire w_dff_A_SvPx8n7A4_1;
	wire w_dff_A_PHOxtYAj4_1;
	wire w_dff_B_gpjAV2IP4_0;
	wire w_dff_A_yMeXOukv4_0;
	wire w_dff_A_kiesjfqD5_1;
	wire w_dff_A_lkebg2m49_0;
	wire w_dff_A_saCiEqOW4_0;
	wire w_dff_A_IeajTyD19_2;
	wire w_dff_A_cOP0zIfQ1_2;
	wire w_dff_B_TdvY5iUP8_3;
	wire w_dff_B_vwyHxJUz9_2;
	wire w_dff_A_ALQxHeVA9_1;
	wire w_dff_A_3SgIPXym6_0;
	wire w_dff_A_qdqTPmX23_0;
	wire w_dff_A_8PK2wp6P7_0;
	wire w_dff_A_fu73Tlq03_0;
	wire w_dff_A_lJgjFNBv1_0;
	wire w_dff_A_Kc7QnGub5_2;
	wire w_dff_A_kYqCcBmS4_2;
	wire w_dff_A_VxmxJFC47_2;
	wire w_dff_A_zAzbZurG5_2;
	wire w_dff_A_mkWMQELe8_2;
	wire w_dff_A_JH7mNzYY0_2;
	wire w_dff_A_TkVW8YX26_0;
	wire w_dff_A_6GvLxx1O3_0;
	wire w_dff_B_r8CDHUvp8_1;
	wire w_dff_A_DSmlpsRc5_0;
	wire w_dff_A_CKNJDBMO5_1;
	wire w_dff_B_OTz8mCiT7_3;
	wire w_dff_B_pCvg8te93_3;
	wire w_dff_B_FjK7oy4T4_3;
	wire w_dff_A_FKwiEQCc1_1;
	wire w_dff_B_38toSO1e7_2;
	wire w_dff_B_SuaWyHO09_0;
	wire w_dff_B_POD5FexQ7_2;
	wire w_dff_A_J6r5C7CT5_0;
	wire w_dff_A_3Ik7xgJC2_0;
	wire w_dff_A_zLjQ5DjK5_0;
	wire w_dff_A_COV5c8io0_1;
	wire w_dff_A_R3eqTsLf5_1;
	wire w_dff_A_A5IuR94N6_1;
	wire w_dff_A_Clk3MhQA4_0;
	wire w_dff_A_f7ZbnAm77_2;
	wire w_dff_A_I1kg5hwF5_1;
	wire w_dff_A_TmbHF47T2_2;
	wire w_dff_B_UYS0eS4J9_3;
	wire w_dff_B_WUUlKJsV5_1;
	wire w_dff_B_uklByK084_1;
	wire w_dff_B_YRVpBmOv9_1;
	wire w_dff_B_JZn9NJq96_1;
	wire w_dff_B_5ogbdSgK0_1;
	wire w_dff_B_j1bxsFnM1_1;
	wire w_dff_A_tlUmzFcf7_1;
	wire w_dff_A_WnJsyQ5g5_2;
	wire w_dff_B_XafTWfcB9_1;
	wire w_dff_B_K0R0tMJv5_1;
	wire w_dff_B_FXHEeOVC0_1;
	wire w_dff_B_oYG8wl3J8_1;
	wire w_dff_B_BFqQdm8s5_1;
	wire w_dff_B_CEpUt50U2_1;
	wire w_dff_A_QzJM2grK0_1;
	wire w_dff_A_cTybTbj10_1;
	wire w_dff_A_W3wxZAmc9_1;
	wire w_dff_A_ul88dtbB2_1;
	wire w_dff_A_Vzqp7Vvv8_1;
	wire w_dff_A_8EXInkQS7_1;
	wire w_dff_A_wyUeuZlK6_1;
	wire w_dff_B_WL4qxRGH8_1;
	wire w_dff_B_lk8j5RSt0_1;
	wire w_dff_B_Nga9kcJ61_1;
	wire w_dff_B_8GAf0KfY6_0;
	wire w_dff_B_qVIVlfkD1_0;
	wire w_dff_A_U3yPJwqJ7_1;
	wire w_dff_A_SFvtqPTS6_1;
	wire w_dff_A_0ninUoKv6_1;
	wire w_dff_A_Kd5FgdbA3_1;
	wire w_dff_A_TKaqkm4w4_1;
	wire w_dff_A_fUZ5YBIY0_1;
	wire w_dff_A_tKNjPyhs0_1;
	wire w_dff_B_sFbHan702_3;
	wire w_dff_A_e7HYpYfB3_0;
	wire w_dff_A_r3KvVKkS4_0;
	wire w_dff_A_2BuvrVVT2_1;
	wire w_dff_A_0l7TO2iJ5_1;
	wire w_dff_A_fyMyRoDP8_1;
	wire w_dff_A_P18OMZwK3_1;
	wire w_dff_A_NnGvldnt2_2;
	wire w_dff_A_jA8P3gX08_2;
	wire w_dff_A_58Aotwi94_1;
	wire w_dff_A_fJyzpPt58_1;
	wire w_dff_A_NbZ0Cjgl5_1;
	wire w_dff_A_40Q8aFAP7_1;
	wire w_dff_A_Umaz5U2i0_1;
	wire w_dff_A_KZ1JfUh10_1;
	wire w_dff_A_xpjQbR8o5_1;
	wire w_dff_A_7m5EH2e48_1;
	wire w_dff_A_cvJ4WcHM2_1;
	wire w_dff_B_beFGc0zb8_1;
	wire w_dff_A_M0K3L6hV2_1;
	wire w_dff_A_X7XREVbh4_1;
	wire w_dff_A_axafGabF4_1;
	wire w_dff_A_Tl530lgX9_1;
	wire w_dff_A_FHA5ViFc5_1;
	wire w_dff_A_KBWSiNeo9_0;
	wire w_dff_A_JGGWZiWw8_0;
	wire w_dff_A_tzQcv87I2_0;
	wire w_dff_A_uLz37Kji1_0;
	wire w_dff_A_AccwtbgX6_0;
	wire w_dff_A_u8ECvRTL7_2;
	wire w_dff_A_eylm4DLO2_2;
	wire w_dff_A_jp9X043D2_2;
	wire w_dff_A_I8RaLy6L4_2;
	wire w_dff_A_d3Ly3WpX8_2;
	wire w_dff_A_zQt3MYHd7_0;
	wire w_dff_A_JyL1JZpr0_0;
	wire w_dff_A_zEL2RL1p2_0;
	wire w_dff_A_bDYceyS95_0;
	wire w_dff_A_iVrP5siR5_0;
	wire w_dff_A_XSA9UEDR7_0;
	wire w_dff_A_1YYsurjX7_0;
	wire w_dff_A_KZxb49b16_0;
	wire w_dff_A_UTbR2gQ65_0;
	wire w_dff_A_DkAMU0IW5_0;
	wire w_dff_A_L645vFdR8_0;
	wire w_dff_A_fnjVZbrO0_0;
	wire w_dff_A_HX0s9Wqt5_0;
	wire w_dff_A_C1oU3Xa71_0;
	wire w_dff_B_IUWquhTG7_2;
	wire w_dff_A_Nb8TqsbK3_0;
	wire w_dff_A_Fozfva622_0;
	wire w_dff_A_FlxckdQo0_0;
	wire w_dff_A_yCPGP2PD1_0;
	wire w_dff_A_RuIPQOuh1_0;
	wire w_dff_A_kfeGpP0u2_0;
	wire w_dff_A_TvEj2aQY8_0;
	wire w_dff_A_SvLAo0DM1_0;
	wire w_dff_B_eYBTCMCd2_3;
	wire w_dff_B_dJQNrJGn0_3;
	wire w_dff_A_2NVq1sYn1_1;
	wire w_dff_A_ZtEfrsOh1_1;
	wire w_dff_A_StFfRhm90_1;
	wire w_dff_B_DleYBDfH4_1;
	wire w_dff_B_wKOLTsfF6_1;
	wire w_dff_B_g5j2zA5F0_1;
	wire w_dff_B_VC0glfyq1_1;
	wire w_dff_B_eidb97056_1;
	wire w_dff_A_UGyPXClN7_0;
	wire w_dff_A_N6FXMaXC1_0;
	wire w_dff_A_FRKufGZR2_0;
	wire w_dff_A_lZnqX16A3_0;
	wire w_dff_A_XnJVb39u4_0;
	wire w_dff_A_7svpxIJm4_0;
	wire w_dff_A_8Wr2l8kp8_0;
	wire w_dff_A_inAgN7b92_0;
	wire w_dff_B_fS85srqe2_0;
	wire w_dff_A_P8cvXJkE8_1;
	wire w_dff_A_XaHotoUV6_1;
	wire w_dff_A_pWYZLlQF0_1;
	wire w_dff_A_CDoiX9gV3_1;
	wire w_dff_A_Uz2qX9xz4_1;
	wire w_dff_A_TJQ3WB8z4_1;
	wire w_dff_A_IBug5IEA4_0;
	wire w_dff_A_XbEjRKiI4_0;
	wire w_dff_A_yfToKdmr0_0;
	wire w_dff_A_D9WkKbMJ7_0;
	wire w_dff_A_HcECIPF01_0;
	wire w_dff_A_5cnqSymo7_1;
	wire w_dff_A_NzIIuW7N3_1;
	wire w_dff_A_2JJl2eq21_1;
	wire w_dff_A_4oeNhO5j5_1;
	wire w_dff_A_P6dePn5q4_1;
	wire w_dff_A_U1uDaDXn2_0;
	wire w_dff_A_9I7aLvHq1_0;
	wire w_dff_A_xzHN8wSu2_0;
	wire w_dff_A_tq3evxCx6_1;
	wire w_dff_B_pd0qDGl43_0;
	wire w_dff_B_DKTaPvg74_1;
	wire w_dff_A_U2ppfvjE4_1;
	wire w_dff_A_5ITBupW48_1;
	wire w_dff_A_AJUc31BI1_1;
	wire w_dff_A_7MlgHC1q0_1;
	wire w_dff_A_oBrJVQhk2_1;
	wire w_dff_A_LapVrmbC6_1;
	wire w_dff_A_QykndE3a9_1;
	wire w_dff_A_kHIeJ6Uj7_1;
	wire w_dff_A_YYyDqyYz5_1;
	wire w_dff_A_sBGeQd331_1;
	wire w_dff_A_7w5DLCYU4_1;
	wire w_dff_A_U2HY2R2g0_1;
	wire w_dff_B_1gtld1Sf8_0;
	wire w_dff_A_Ui9PJ5O17_1;
	wire w_dff_A_iohcq6jF2_1;
	wire w_dff_A_s5LjUzUz6_1;
	wire w_dff_A_05OadJCG7_1;
	wire w_dff_A_vD5CDa2t9_1;
	wire w_dff_A_cyhc6bz82_1;
	wire w_dff_A_jXYcU6KF0_1;
	wire w_dff_A_dUMFPHWU8_1;
	wire w_dff_A_WEugoDzi0_1;
	wire w_dff_A_FW6HIXuH1_1;
	wire w_dff_A_lbkTf7lM7_1;
	wire w_dff_A_ttOo4taJ6_1;
	wire w_dff_A_pYAaDC458_1;
	wire w_dff_A_1kv7ps4W5_0;
	wire w_dff_A_bVhzwMjI8_0;
	wire w_dff_A_oySK6syp2_0;
	wire w_dff_A_qACBYdFH4_0;
	wire w_dff_A_7xFuLcjY5_0;
	wire w_dff_A_jlbDLggY5_0;
	wire w_dff_A_BaMYHZHI9_0;
	wire w_dff_A_GsL44PON1_0;
	wire w_dff_A_NtxSgBHr6_0;
	wire w_dff_A_fIKNUMVk9_0;
	wire w_dff_A_mvQDJjhl0_0;
	wire w_dff_A_lFGwgagg5_1;
	wire w_dff_A_QcNN8d9r8_0;
	wire w_dff_A_D8YtNXkA7_0;
	wire w_dff_A_a3NvIrc59_0;
	wire w_dff_A_HNJ7I9yW0_0;
	wire w_dff_A_lkvy8Bwq1_0;
	wire w_dff_A_WDfWyDR46_0;
	wire w_dff_A_bG1umpQW1_0;
	wire w_dff_A_K9TOOPpx4_0;
	wire w_dff_A_IrIcfeQV9_0;
	wire w_dff_A_oTFCBXD72_0;
	wire w_dff_A_ryt0mnN75_0;
	wire w_dff_A_NC3t7dCW0_1;
	wire w_dff_A_WBnHEDFy2_1;
	wire w_dff_A_BSyXgYxY5_1;
	wire w_dff_A_uEvwOPuB5_0;
	wire w_dff_A_pCNrg0vZ5_0;
	wire w_dff_A_Q2jMbFOm1_0;
	wire w_dff_A_3YgReqlg4_1;
	wire w_dff_A_8ddO8xqX1_1;
	wire w_dff_A_ftWgLyG90_1;
	wire w_dff_A_pudfbXUd3_1;
	wire w_dff_A_1rOVvtp43_1;
	wire w_dff_A_npsImUZ42_1;
	wire w_dff_B_VME5RSDq1_2;
	wire w_dff_A_UUgdfLni5_2;
	wire w_dff_A_giDHr2hO0_2;
	wire w_dff_A_2xbg2hI77_0;
	wire w_dff_A_gKwlaWvY7_0;
	wire w_dff_A_6wOHC4WP1_0;
	wire w_dff_A_5FM4vTTV2_0;
	wire w_dff_A_l1t6oyFZ3_0;
	wire w_dff_A_ffJhr80R9_0;
	wire w_dff_A_AkhowQR99_0;
	wire w_dff_A_MXEDLgJw5_0;
	wire w_dff_A_Y0C9aZBy3_0;
	wire w_dff_A_1qEgt9xC6_0;
	wire w_dff_A_AhPFVJ2L0_0;
	wire w_dff_A_gyPgl8wT6_0;
	wire w_dff_A_5RNRl6Vb1_0;
	wire w_dff_A_IeQ2PzdK7_0;
	wire w_dff_A_fYHZdvQU1_0;
	wire w_dff_A_LIZk3YRo9_0;
	wire w_dff_A_3Myj1NgY5_0;
	wire w_dff_A_UoXBNYhe1_0;
	wire w_dff_A_u0r9HC9p1_0;
	wire w_dff_A_t6o6BoYO8_1;
	wire w_dff_A_cSU03OiF5_1;
	wire w_dff_B_5KcbtH9R0_3;
	wire w_dff_A_2RV8VcwV1_0;
	wire w_dff_A_KrZ6EOnd6_2;
	wire w_dff_A_eRzN8rTf6_0;
	wire w_dff_A_AwgT4ywJ4_0;
	wire w_dff_A_IyPAJ7Mx6_0;
	wire w_dff_A_nhBxEeyT8_0;
	wire w_dff_A_fVJcP9a34_0;
	wire w_dff_A_Y9wtmFol1_0;
	wire w_dff_A_cmXUqGba9_0;
	wire w_dff_A_kvPhKXs88_0;
	wire w_dff_A_5YaAlyT65_0;
	wire w_dff_A_OAHrCjFq3_0;
	wire w_dff_A_vhETZMxO6_0;
	wire w_dff_A_v7t7nDrW0_2;
	wire w_dff_A_FtYLZEww0_2;
	wire w_dff_B_y2ks6dKP9_3;
	wire w_dff_A_xxPCt6PZ4_1;
	wire w_dff_A_OwpnqkYD3_1;
	wire w_dff_A_24rS6dwG1_0;
	wire w_dff_A_JuzkRHvL1_0;
	wire w_dff_A_ndAlKMie2_0;
	wire w_dff_A_dRQnyY7x9_0;
	wire w_dff_A_teWS2zCG1_0;
	wire w_dff_A_zf2SE4mo1_0;
	wire w_dff_A_UcxAfrCR0_0;
	wire w_dff_A_f7rNHEMz5_0;
	wire w_dff_A_pluT9Enz8_0;
	wire w_dff_A_OdM7OG2W7_0;
	wire w_dff_A_MS1gN8KP4_0;
	wire w_dff_A_826U4WMO5_0;
	wire w_dff_A_cAGfDvLN2_0;
	wire w_dff_A_e9SMnYKh6_0;
	wire w_dff_A_plsqT4a13_0;
	wire w_dff_A_VyfcBy0g6_0;
	wire w_dff_A_8hrwlRli4_0;
	wire w_dff_A_ITTT5owe8_0;
	wire w_dff_A_u32QCrcr8_0;
	wire w_dff_A_ucaaQgz70_0;
	wire w_dff_A_XQT0xlrj6_0;
	wire w_dff_A_BKpryq4U4_0;
	wire w_dff_A_ZLODwrnj3_2;
	wire w_dff_A_dZrJtdGE4_2;
	wire w_dff_A_FWBvyt5U0_2;
	wire w_dff_A_s4MrnL4K3_0;
	wire w_dff_A_cNSo23I08_0;
	wire w_dff_A_7tprLKZE3_0;
	wire w_dff_A_WrPST0t00_0;
	wire w_dff_A_tw4Tdoqw7_0;
	wire w_dff_A_v1e3CKb47_0;
	wire w_dff_A_wd1xCyMQ7_0;
	wire w_dff_A_c2NcYIJT3_0;
	wire w_dff_A_KQHvbKUM8_0;
	wire w_dff_A_QqfFmQx10_0;
	wire w_dff_A_3HnYfHIg9_0;
	wire w_dff_A_LZJINklu6_1;
	wire w_dff_A_BRpmqw9O3_0;
	wire w_dff_A_VVy7NlmP9_0;
	wire w_dff_A_QEeP222e7_0;
	wire w_dff_A_5WFHONCN6_0;
	wire w_dff_A_BpoZLH6c1_0;
	wire w_dff_A_oT5TMHdb4_0;
	wire w_dff_A_BKSBWluH8_0;
	wire w_dff_A_RRv6MsYz4_0;
	wire w_dff_A_WPsuIQJe9_0;
	wire w_dff_A_GyKhO8CR3_0;
	wire w_dff_A_kBvrLY7q2_0;
	wire w_dff_A_iuCcpqQN4_2;
	wire w_dff_A_1SL49ZY94_0;
	wire w_dff_A_zctUQblE6_0;
	wire w_dff_A_fxNmxl9i1_0;
	wire w_dff_A_dvabvz5G6_0;
	wire w_dff_A_qNzGlO3j2_0;
	wire w_dff_A_qRPjnq8j3_0;
	wire w_dff_A_CfQGplYX8_0;
	wire w_dff_A_V6NZBuYY6_0;
	wire w_dff_A_dSYd7Wko1_0;
	wire w_dff_A_UUIYuLPL5_0;
	wire w_dff_A_obgZl6jG1_0;
	wire w_dff_A_GApTDjgN1_0;
	wire w_dff_A_SNBSiXTw9_0;
	wire w_dff_A_VF7R0M0a8_0;
	wire w_dff_A_ZHudeNIm6_0;
	wire w_dff_A_DtPHaBP40_0;
	wire w_dff_A_xo3NQvQi6_0;
	wire w_dff_A_7ngWHTDD3_0;
	wire w_dff_A_qhxDTkZz0_0;
	wire w_dff_A_kFjFqPnk8_0;
	wire w_dff_A_WsLv4gx42_0;
	wire w_dff_A_QCd9yhUo1_0;
	wire w_dff_A_sXuUSNHX8_0;
	wire w_dff_A_FU9JAAiV3_0;
	wire w_dff_A_m7bR6HhP1_2;
	wire w_dff_A_vALIWXhM6_2;
	wire w_dff_A_cdvz8ir87_2;
	wire w_dff_A_QXjW7J0L2_2;
	wire w_dff_A_OaL2mG203_2;
	wire w_dff_A_rmsSqK9p0_2;
	wire w_dff_A_ICOXnSjx7_2;
	wire w_dff_B_gC6kq2403_3;
	wire w_dff_B_8rLfO2R71_0;
	wire w_dff_B_ahKLhWif8_0;
	wire w_dff_B_YYY2vQAx9_0;
	wire w_dff_A_PxOqAoKK5_0;
	wire w_dff_A_brUGOvlL4_0;
	wire w_dff_A_KhHx9UBa5_0;
	wire w_dff_A_Gxhitpy44_0;
	wire w_dff_A_lIqe7Wt14_0;
	wire w_dff_A_6xYUyHOP2_0;
	wire w_dff_A_z3pJz3030_0;
	wire w_dff_A_s2tO7NjE4_0;
	wire w_dff_A_ycnG1fB95_0;
	wire w_dff_A_HTrla1TD9_0;
	wire w_dff_A_GH1zlFqY8_0;
	wire w_dff_A_oCC99aW00_0;
	wire w_dff_A_Uvr7HL5t3_0;
	wire w_dff_A_p7pPbWTJ5_0;
	wire w_dff_A_xxxnEkvb4_0;
	wire w_dff_A_Gw1p1y5E4_0;
	wire w_dff_A_gdmvXRrI7_2;
	wire w_dff_A_UmtzS4231_0;
	wire w_dff_A_jRr75Cmx9_0;
	wire w_dff_A_DAbspYrE9_0;
	wire w_dff_A_9bilBzyQ2_0;
	wire w_dff_A_wnx3vDL48_0;
	wire w_dff_A_Jk449MZf5_0;
	wire w_dff_A_A92UaAXC8_0;
	wire w_dff_A_SlqB5pf85_0;
	wire w_dff_A_Pnv99A6v3_0;
	wire w_dff_B_Ky51Spd31_1;
	wire w_dff_A_GoMcK60a0_0;
	wire w_dff_A_ju48mgPi5_0;
	wire w_dff_A_5m1Idbjk0_0;
	wire w_dff_A_aYGK7AyO5_0;
	wire w_dff_A_iJsy2A5X6_0;
	wire w_dff_A_p2O1MixS4_0;
	wire w_dff_A_vallSv8x8_0;
	wire w_dff_A_tBEckXBN3_0;
	wire w_dff_A_0KZcFYYb5_0;
	wire w_dff_A_mVMKXJXE7_0;
	wire w_dff_A_HCI87VPS2_0;
	wire w_dff_A_mF7KzgY93_0;
	wire w_dff_A_SJxdXh8r0_2;
	wire w_dff_A_FvvqJ0nI3_0;
	wire w_dff_A_e5vFrYof2_0;
	wire w_dff_A_4FSks8iq8_0;
	wire w_dff_A_xMSghTd98_0;
	wire w_dff_A_N6Pb9mBT2_0;
	wire w_dff_A_e31nRQDY6_0;
	wire w_dff_A_ghKRT1N76_0;
	wire w_dff_A_yTUZHwgc7_0;
	wire w_dff_A_jTfhHgsa5_0;
	wire w_dff_A_vEr9B57F2_0;
	wire w_dff_A_DSi8Rwoj8_0;
	wire w_dff_A_yilBa07N3_0;
	wire w_dff_A_MJ3Mp4tL8_0;
	wire w_dff_A_OeoskeEG5_0;
	wire w_dff_A_Gz4AiwIu0_0;
	wire w_dff_A_llAGGRBC0_0;
	wire w_dff_A_8rGGDLr17_0;
	wire w_dff_A_GTo0dIFo7_0;
	wire w_dff_A_ki44nNqs2_0;
	wire w_dff_A_SVgvjFl49_0;
	wire w_dff_A_Rd0LLEzI0_0;
	wire w_dff_A_gEjCxq0P0_0;
	wire w_dff_A_Uohm0taf4_0;
	wire w_dff_A_kKbp1AZV4_2;
	wire w_dff_A_G3lp0cUe0_2;
	wire w_dff_A_APhnHAiT2_0;
	wire w_dff_B_iPWazfDc1_2;
	wire w_dff_A_RxTxGRxh9_0;
	wire w_dff_A_K3IqHHkr1_0;
	wire w_dff_A_KK7Kz5PD7_0;
	wire w_dff_A_oejqsVYU9_0;
	wire w_dff_A_2cgMUa5v4_0;
	wire w_dff_A_96TMQNo51_0;
	wire w_dff_A_4tSXdq7W5_0;
	wire w_dff_A_djmY2uR50_0;
	wire w_dff_A_hajWMwuI4_0;
	wire w_dff_A_2yLr4S3i8_0;
	wire w_dff_A_ZZH3glHj2_0;
	wire w_dff_A_vxEeDK438_0;
	wire w_dff_A_NKLohOZ70_0;
	wire w_dff_A_IsyiABwm5_0;
	wire w_dff_A_0Lst71Nm1_0;
	wire w_dff_A_t18dTeM72_0;
	wire w_dff_A_kUW22AGN3_0;
	wire w_dff_A_XKEZtip65_0;
	wire w_dff_A_ByBdzqzV6_0;
	wire w_dff_A_6HEV8Rev6_0;
	wire w_dff_A_tU1wH5D77_0;
	wire w_dff_A_V8DD8o0t6_0;
	wire w_dff_A_Xeczaa3W7_0;
	wire w_dff_A_pUzB4IKe8_0;
	wire w_dff_A_AO7eyqxq1_0;
	wire w_dff_A_hAbroMB57_0;
	wire w_dff_A_Pstr7MMN1_1;
	wire w_dff_A_AcWRQco98_1;
	wire w_dff_A_YA06VvK44_0;
	wire w_dff_A_pXsO4R0K4_0;
	wire w_dff_A_eVl1fKW27_0;
	wire w_dff_A_pyNQCoWl4_0;
	wire w_dff_A_P1W2Ql8z9_0;
	wire w_dff_A_e7zaB9HF0_0;
	wire w_dff_A_K4dsJa0A9_0;
	wire w_dff_A_p9bIWyfp6_0;
	wire w_dff_A_62Ctg2Ne2_0;
	wire w_dff_A_GFIt6KrB0_0;
	wire w_dff_B_V41iQZ8u6_3;
	wire w_dff_B_C2m4WaSq7_1;
	wire w_dff_A_ni3v0n9z5_0;
	wire w_dff_A_x4psjkTG0_0;
	wire w_dff_A_dfsJwcK68_0;
	wire w_dff_A_Uh9PD1Lh7_0;
	wire w_dff_A_MflngdFi7_0;
	wire w_dff_A_KDUjAa3E2_0;
	wire w_dff_A_YFxe02qr7_0;
	wire w_dff_A_Aie8JjQ77_0;
	wire w_dff_A_Cr9nVUDA1_0;
	wire w_dff_A_BrWIWytB0_0;
	wire w_dff_A_m8FNkz492_0;
	wire w_dff_A_g5Yaeth48_0;
	wire w_dff_A_iKE1LC3X9_0;
	wire w_dff_A_tREwYbIJ1_0;
	wire w_dff_A_GCmGLdxp6_1;
	wire w_dff_A_6gcsZIfy2_1;
	wire w_dff_A_1z5eNIe28_1;
	wire w_dff_A_1o9DG4HD1_1;
	wire w_dff_A_slIohsjf2_2;
	wire w_dff_A_PSGJPxpB0_2;
	wire w_dff_A_eOiVXpce8_2;
	wire w_dff_A_pltyNh1r3_2;
	wire w_dff_A_SmRkh54p1_2;
	wire w_dff_A_hvpjNHhD4_0;
	wire w_dff_A_FoTLtxJU6_0;
	wire w_dff_A_9gDH7QjS7_0;
	wire w_dff_A_STTiZQIw4_0;
	wire w_dff_A_hC6Riofy9_0;
	wire w_dff_A_EenXafGX8_1;
	wire w_dff_A_DixJRMo74_1;
	wire w_dff_A_UQ5ELU4O9_1;
	wire w_dff_A_OpYzNYPk9_1;
	wire w_dff_A_DX1Jtd824_1;
	wire w_dff_A_F2jV7Pd82_1;
	wire w_dff_A_V6Xc0F5r1_1;
	wire w_dff_A_55eobgb14_1;
	wire w_dff_A_jtykbg1A3_1;
	wire w_dff_A_ImdvI9Mn8_1;
	wire w_dff_A_YN775MRB6_1;
	wire w_dff_A_jYiAAeD65_1;
	wire w_dff_A_hL35ZfMB4_1;
	wire w_dff_A_ZwwODbhB0_1;
	wire w_dff_A_zuPO9N7w4_2;
	wire w_dff_A_730B2bu67_2;
	wire w_dff_A_m7SLLc3W2_2;
	wire w_dff_A_LUYkr2Q20_2;
	wire w_dff_A_NoRgml0h4_2;
	wire w_dff_A_Lf0gwY4J0_2;
	wire w_dff_A_WZFxI3PM5_2;
	wire w_dff_A_jIsy6JS41_2;
	wire w_dff_A_gIGhulHP0_2;
	wire w_dff_A_uvdrltih3_2;
	wire w_dff_A_PSf7OqsH6_2;
	wire w_dff_A_CxHygDJm3_2;
	wire w_dff_A_w6irMycR8_2;
	wire w_dff_A_VyAK8UQF8_2;
	wire w_dff_A_kyALfS8y8_2;
	wire w_dff_A_S93cdf7v1_0;
	wire w_dff_A_T6QzBcsh7_2;
	wire w_dff_B_bSRuW6T07_3;
	wire w_dff_B_QhVnIGew8_3;
	wire w_dff_B_tT049HkM7_3;
	wire w_dff_B_0KDNIxUo6_3;
	wire w_dff_B_vs7CnyFM2_3;
	wire w_dff_B_Wg43Mll57_3;
	wire w_dff_B_vwXDQ3k44_3;
	wire w_dff_B_3rbTZAy59_3;
	wire w_dff_B_3iUJite09_3;
	wire w_dff_B_OKuATHPp5_3;
	wire w_dff_B_D0uIuEKW5_3;
	wire w_dff_B_4jiMGCk33_3;
	wire w_dff_B_xMgHvZ9D3_3;
	wire w_dff_A_PhPMIR101_0;
	wire w_dff_A_PE0GXOYn3_0;
	wire w_dff_A_papfaKOE8_0;
	wire w_dff_A_m0CurfKx7_0;
	wire w_dff_A_wQoLfVjt4_0;
	wire w_dff_A_Jm8wX8NX2_0;
	wire w_dff_A_1eKLivb79_0;
	wire w_dff_A_yekxO9qK3_0;
	wire w_dff_A_QxVqPfhw6_0;
	wire w_dff_A_lZERSlmd7_0;
	wire w_dff_A_zRhpTNeS3_0;
	wire w_dff_A_YmhNpf6I9_0;
	wire w_dff_A_qLXv9ayE6_1;
	wire w_dff_A_NFSuWSaA9_0;
	wire w_dff_A_sm3iMdGl3_1;
	wire w_dff_A_kqCYD7ff0_1;
	wire w_dff_A_LisM0hWW6_1;
	wire w_dff_A_siV0kBdx2_1;
	wire w_dff_A_WCoM8kKN6_1;
	wire w_dff_A_dDm8YGSF9_1;
	wire w_dff_A_IjUh3WNQ5_1;
	wire w_dff_A_jgwiAHf38_1;
	wire w_dff_A_7Izl4Wsj3_1;
	wire w_dff_A_OeAHGV3d7_1;
	wire w_dff_A_EkyAUfKq3_1;
	wire w_dff_A_YKAltODn9_1;
	wire w_dff_A_lX7bwFbg2_1;
	jnot g000(.din(w_G902_4[2]),.dout(n59),.clk(gclk));
	jnot g001(.din(w_G137_0[2]),.dout(n60),.clk(gclk));
	jnot g002(.din(w_G953_3[1]),.dout(n61),.clk(gclk));
	jand g003(.dina(w_G234_1[1]),.dinb(w_G221_0[1]),.dout(n62),.clk(gclk));
	jand g004(.dina(n62),.dinb(w_n61_3[2]),.dout(n63),.clk(gclk));
	jxor g005(.dina(n63),.dinb(w_dff_B_C2m4WaSq7_1),.dout(n64),.clk(gclk));
	jxor g006(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n65),.clk(gclk));
	jxor g007(.dina(w_n65_0[1]),.dinb(w_G146_0[2]),.dout(n66),.clk(gclk));
	jnot g008(.din(w_G110_0[2]),.dout(n67),.clk(gclk));
	jxor g009(.dina(w_G119_0[2]),.dinb(w_n67_0[1]),.dout(n68),.clk(gclk));
	jxor g010(.dina(n68),.dinb(w_G128_0[2]),.dout(n69),.clk(gclk));
	jxor g011(.dina(n69),.dinb(w_n66_0[1]),.dout(n70),.clk(gclk));
	jxor g012(.dina(n70),.dinb(w_dff_B_Ky51Spd31_1),.dout(n71),.clk(gclk));
	jand g013(.dina(w_n71_0[1]),.dinb(w_n59_2[1]),.dout(n72),.clk(gclk));
	jnot g014(.din(w_G234_1[0]),.dout(n73),.clk(gclk));
	jcb g015(.dina(w_G902_4[1]),.dinb(n73),.dout(n74));
	jand g016(.dina(w_n74_0[1]),.dinb(w_G217_0[2]),.dout(n75),.clk(gclk));
	jnot g017(.din(w_n75_0[1]),.dout(n76),.clk(gclk));
	jxor g018(.dina(w_dff_B_YYY2vQAx9_0),.dinb(w_n72_0[1]),.dout(n77),.clk(gclk));
	jxor g019(.dina(w_G143_0[2]),.dinb(w_G128_0[1]),.dout(n78),.clk(gclk));
	jxor g020(.dina(w_n78_0[1]),.dinb(w_G146_0[1]),.dout(n79),.clk(gclk));
	jxor g021(.dina(w_G137_0[1]),.dinb(w_G134_0[2]),.dout(n80),.clk(gclk));
	jxor g022(.dina(n80),.dinb(w_G131_0[2]),.dout(n81),.clk(gclk));
	jxor g023(.dina(n81),.dinb(w_n79_0[1]),.dout(n82),.clk(gclk));
	jxor g024(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g025(.dina(n83),.dinb(w_G113_0[2]),.dout(n84),.clk(gclk));
	jnot g026(.din(w_G237_0[1]),.dout(n85),.clk(gclk));
	jand g027(.dina(w_n61_3[1]),.dinb(w_G210_0[2]),.dout(n86),.clk(gclk));
	jand g028(.dina(n86),.dinb(w_n85_0[2]),.dout(n87),.clk(gclk));
	jxor g029(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g030(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g031(.dina(n89),.dinb(w_n82_0[2]),.dout(n90),.clk(gclk));
	jand g032(.dina(w_n90_0[1]),.dinb(w_n59_2[0]),.dout(n91),.clk(gclk));
	jxor g033(.dina(w_n91_0[1]),.dinb(w_G472_0[2]),.dout(n92),.clk(gclk));
	jand g034(.dina(w_n92_1[1]),.dinb(w_n77_1[1]),.dout(n93),.clk(gclk));
	jand g035(.dina(w_n59_1[2]),.dinb(w_n85_0[1]),.dout(n94),.clk(gclk));
	jnot g036(.din(n94),.dout(n95),.clk(gclk));
	jand g037(.dina(w_n95_0[1]),.dinb(w_G214_0[1]),.dout(n96),.clk(gclk));
	jxor g038(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n97),.clk(gclk));
	jxor g039(.dina(n97),.dinb(w_G101_0[1]),.dout(n98),.clk(gclk));
	jxor g040(.dina(w_n98_0[1]),.dinb(w_n84_0[0]),.dout(n99),.clk(gclk));
	jxor g041(.dina(w_G122_1[1]),.dinb(w_n67_0[0]),.dout(n100),.clk(gclk));
	jxor g042(.dina(w_dff_B_1gtld1Sf8_0),.dinb(n99),.dout(n101),.clk(gclk));
	jand g043(.dina(w_n61_3[0]),.dinb(w_G224_0[1]),.dout(n102),.clk(gclk));
	jxor g044(.dina(w_n79_0[0]),.dinb(w_G125_0[1]),.dout(n103),.clk(gclk));
	jxor g045(.dina(n103),.dinb(w_dff_B_DKTaPvg74_1),.dout(n104),.clk(gclk));
	jxor g046(.dina(n104),.dinb(w_n101_0[2]),.dout(n105),.clk(gclk));
	jcb g047(.dina(w_n105_0[1]),.dinb(w_G902_4[0]),.dout(n106));
	jand g048(.dina(w_n95_0[0]),.dinb(w_G210_0[1]),.dout(n107),.clk(gclk));
	jxor g049(.dina(w_dff_B_pd0qDGl43_0),.dinb(n106),.dout(n108),.clk(gclk));
	jcb g050(.dina(w_n108_0[2]),.dinb(w_n96_0[1]),.dout(n109));
	jnot g051(.din(w_n109_0[2]),.dout(n110),.clk(gclk));
	jand g052(.dina(w_n74_0[0]),.dinb(w_G221_0[0]),.dout(n111),.clk(gclk));
	jnot g053(.din(w_n111_0[2]),.dout(n112),.clk(gclk));
	jnot g054(.din(w_n82_0[1]),.dout(n113),.clk(gclk));
	jnot g055(.din(w_G227_0[1]),.dout(n114),.clk(gclk));
	jcb g056(.dina(w_G953_3[0]),.dinb(n114),.dout(n115));
	jxor g057(.dina(w_G140_0[1]),.dinb(w_G110_0[1]),.dout(n116),.clk(gclk));
	jxor g058(.dina(n116),.dinb(n115),.dout(n117),.clk(gclk));
	jxor g059(.dina(n117),.dinb(w_n98_0[0]),.dout(n118),.clk(gclk));
	jxor g060(.dina(w_dff_B_fS85srqe2_0),.dinb(n113),.dout(n119),.clk(gclk));
	jand g061(.dina(w_n119_0[1]),.dinb(w_n59_1[1]),.dout(n120),.clk(gclk));
	jxor g062(.dina(n120),.dinb(w_G469_0[1]),.dout(n121),.clk(gclk));
	jand g063(.dina(w_n121_0[2]),.dinb(w_dff_B_eidb97056_1),.dout(n122),.clk(gclk));
	jand g064(.dina(w_n122_0[2]),.dinb(w_dff_B_DleYBDfH4_1),.dout(n123),.clk(gclk));
	jnot g065(.din(w_G952_0[2]),.dout(n124),.clk(gclk));
	jand g066(.dina(w_G237_0[0]),.dinb(w_G234_0[2]),.dout(n125),.clk(gclk));
	jcb g067(.dina(w_n125_0[1]),.dinb(n124),.dout(n126));
	jcb g068(.dina(n126),.dinb(w_G953_2[2]),.dout(n127));
	jnot g069(.din(n127),.dout(n128),.clk(gclk));
	jnot g070(.din(w_n125_0[0]),.dout(n129),.clk(gclk));
	jnot g071(.din(w_G898_0[1]),.dout(n130),.clk(gclk));
	jand g072(.dina(w_G953_2[1]),.dinb(n130),.dout(n131),.clk(gclk));
	jand g073(.dina(w_n131_0[1]),.dinb(w_G902_3[2]),.dout(n132),.clk(gclk));
	jand g074(.dina(n132),.dinb(w_n129_0[1]),.dout(n133),.clk(gclk));
	jcb g075(.dina(n133),.dinb(w_n128_0[2]),.dout(n134));
	jand g076(.dina(w_G234_0[1]),.dinb(w_G217_0[1]),.dout(n135),.clk(gclk));
	jand g077(.dina(n135),.dinb(w_n61_2[2]),.dout(n136),.clk(gclk));
	jxor g078(.dina(w_n78_0[0]),.dinb(w_G134_0[1]),.dout(n137),.clk(gclk));
	jxor g079(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n138),.clk(gclk));
	jxor g080(.dina(n138),.dinb(w_G107_0[1]),.dout(n139),.clk(gclk));
	jxor g081(.dina(n139),.dinb(n137),.dout(n140),.clk(gclk));
	jxor g082(.dina(n140),.dinb(w_dff_B_beFGc0zb8_1),.dout(n141),.clk(gclk));
	jand g083(.dina(w_n141_0[2]),.dinb(w_n59_1[0]),.dout(n142),.clk(gclk));
	jxor g084(.dina(n142),.dinb(w_G478_0[1]),.dout(n143),.clk(gclk));
	jnot g085(.din(w_n143_1[2]),.dout(n144),.clk(gclk));
	jnot g086(.din(w_G475_0[2]),.dout(n145),.clk(gclk));
	jxor g087(.dina(w_G122_0[2]),.dinb(w_G113_0[1]),.dout(n146),.clk(gclk));
	jxor g088(.dina(n146),.dinb(w_G104_0[1]),.dout(n147),.clk(gclk));
	jand g089(.dina(w_n61_2[1]),.dinb(w_G214_0[0]),.dout(n148),.clk(gclk));
	jand g090(.dina(n148),.dinb(w_n85_0[0]),.dout(n149),.clk(gclk));
	jxor g091(.dina(w_G143_0[1]),.dinb(w_G131_0[1]),.dout(n150),.clk(gclk));
	jxor g092(.dina(w_dff_B_qVIVlfkD1_0),.dinb(n149),.dout(n151),.clk(gclk));
	jxor g093(.dina(n151),.dinb(w_n66_0[0]),.dout(n152),.clk(gclk));
	jxor g094(.dina(n152),.dinb(w_dff_B_Nga9kcJ61_1),.dout(n153),.clk(gclk));
	jand g095(.dina(w_n153_0[2]),.dinb(w_n59_0[2]),.dout(n154),.clk(gclk));
	jxor g096(.dina(w_n154_0[1]),.dinb(w_dff_B_CEpUt50U2_1),.dout(n155),.clk(gclk));
	jand g097(.dina(w_n155_1[2]),.dinb(w_n144_1[1]),.dout(n156),.clk(gclk));
	jand g098(.dina(w_n156_1[1]),.dinb(w_n134_1[2]),.dout(n157),.clk(gclk));
	jand g099(.dina(w_n157_0[1]),.dinb(w_n123_1[1]),.dout(n158),.clk(gclk));
	jand g100(.dina(w_n158_0[1]),.dinb(w_n93_0[2]),.dout(n159),.clk(gclk));
	jxor g101(.dina(w_n159_0[2]),.dinb(w_G101_0[0]),.dout(G3),.clk(gclk));
	jnot g102(.din(w_G472_0[1]),.dout(n161),.clk(gclk));
	jxor g103(.dina(w_n91_0[0]),.dinb(w_dff_B_j1bxsFnM1_1),.dout(n162),.clk(gclk));
	jand g104(.dina(w_n162_1[1]),.dinb(w_n77_1[0]),.dout(n163),.clk(gclk));
	jand g105(.dina(w_n163_1[1]),.dinb(w_n123_1[0]),.dout(n164),.clk(gclk));
	jxor g106(.dina(w_n154_0[0]),.dinb(w_G475_0[1]),.dout(n165),.clk(gclk));
	jand g107(.dina(w_n165_0[2]),.dinb(w_n144_1[0]),.dout(n166),.clk(gclk));
	jand g108(.dina(w_n166_0[1]),.dinb(w_n134_1[1]),.dout(n167),.clk(gclk));
	jand g109(.dina(w_n167_0[2]),.dinb(w_n164_0[1]),.dout(n168),.clk(gclk));
	jxor g110(.dina(w_n168_0[1]),.dinb(w_G104_0[0]),.dout(G6),.clk(gclk));
	jand g111(.dina(w_n155_1[1]),.dinb(w_n143_1[1]),.dout(n170),.clk(gclk));
	jand g112(.dina(w_n170_0[1]),.dinb(w_n134_1[0]),.dout(n171),.clk(gclk));
	jand g113(.dina(w_n171_0[2]),.dinb(w_n164_0[0]),.dout(n172),.clk(gclk));
	jxor g114(.dina(w_n172_0[1]),.dinb(w_G107_0[0]),.dout(G9),.clk(gclk));
	jxor g115(.dina(w_n75_0[0]),.dinb(w_n72_0[0]),.dout(n174),.clk(gclk));
	jand g116(.dina(w_n162_1[0]),.dinb(w_n174_1[1]),.dout(n175),.clk(gclk));
	jand g117(.dina(w_n175_0[1]),.dinb(w_n158_0[0]),.dout(n176),.clk(gclk));
	jxor g118(.dina(w_n176_0[1]),.dinb(w_G110_0[0]),.dout(G12),.clk(gclk));
	jand g119(.dina(w_n92_1[0]),.dinb(w_n174_1[0]),.dout(n178),.clk(gclk));
	jand g120(.dina(w_n178_0[2]),.dinb(w_n123_0[2]),.dout(n179),.clk(gclk));
	jnot g121(.din(w_G900_0[1]),.dout(n180),.clk(gclk));
	jand g122(.dina(w_G953_2[0]),.dinb(n180),.dout(n181),.clk(gclk));
	jand g123(.dina(w_n181_0[1]),.dinb(w_G902_3[1]),.dout(n182),.clk(gclk));
	jand g124(.dina(n182),.dinb(w_n129_0[0]),.dout(n183),.clk(gclk));
	jcb g125(.dina(n183),.dinb(w_n128_0[1]),.dout(n184));
	jand g126(.dina(w_n184_1[2]),.dinb(w_n170_0[0]),.dout(n185),.clk(gclk));
	jand g127(.dina(w_n185_0[2]),.dinb(w_n179_0[1]),.dout(n186),.clk(gclk));
	jxor g128(.dina(w_n186_0[1]),.dinb(w_G128_0[0]),.dout(G30),.clk(gclk));
	jand g129(.dina(w_n165_0[1]),.dinb(w_n143_1[0]),.dout(n188),.clk(gclk));
	jand g130(.dina(w_n188_0[1]),.dinb(w_n93_0[1]),.dout(n189),.clk(gclk));
	jand g131(.dina(n189),.dinb(w_n184_1[1]),.dout(n190),.clk(gclk));
	jand g132(.dina(n190),.dinb(w_n123_0[1]),.dout(n191),.clk(gclk));
	jxor g133(.dina(w_n191_0[1]),.dinb(w_G143_0[0]),.dout(G45),.clk(gclk));
	jand g134(.dina(w_n184_1[0]),.dinb(w_n166_0[0]),.dout(n193),.clk(gclk));
	jand g135(.dina(w_n193_0[2]),.dinb(w_n179_0[0]),.dout(n194),.clk(gclk));
	jxor g136(.dina(w_n194_0[1]),.dinb(w_G146_0[0]),.dout(G48),.clk(gclk));
	jcb g137(.dina(w_n162_0[2]),.dinb(w_n174_0[2]),.dout(n196));
	jcb g138(.dina(w_n121_0[1]),.dinb(w_n111_0[1]),.dout(n197));
	jcb g139(.dina(w_n197_0[1]),.dinb(w_n109_0[1]),.dout(n198));
	jcb g140(.dina(w_n198_1[2]),.dinb(w_n196_0[1]),.dout(n199));
	jnot g141(.din(w_n199_0[2]),.dout(n200),.clk(gclk));
	jand g142(.dina(w_n200_0[1]),.dinb(w_n167_0[1]),.dout(n201),.clk(gclk));
	jxor g143(.dina(w_n201_0[1]),.dinb(w_G113_0[0]),.dout(G15),.clk(gclk));
	jand g144(.dina(w_n200_0[0]),.dinb(w_n171_0[1]),.dout(n203),.clk(gclk));
	jxor g145(.dina(w_n203_0[1]),.dinb(w_G116_0[0]),.dout(G18),.clk(gclk));
	jnot g146(.din(w_n198_1[1]),.dout(n205),.clk(gclk));
	jand g147(.dina(w_n178_0[1]),.dinb(w_n157_0[0]),.dout(n206),.clk(gclk));
	jand g148(.dina(n206),.dinb(w_n205_0[2]),.dout(n207),.clk(gclk));
	jxor g149(.dina(w_n207_0[1]),.dinb(w_G119_0[0]),.dout(G21),.clk(gclk));
	jand g150(.dina(w_n163_1[0]),.dinb(w_n134_0[2]),.dout(n209),.clk(gclk));
	jand g151(.dina(n209),.dinb(w_n188_0[0]),.dout(n210),.clk(gclk));
	jand g152(.dina(n210),.dinb(w_n205_0[1]),.dout(n211),.clk(gclk));
	jxor g153(.dina(w_n211_0[1]),.dinb(w_G122_0[1]),.dout(G24),.clk(gclk));
	jand g154(.dina(w_n193_0[1]),.dinb(w_n175_0[0]),.dout(n213),.clk(gclk));
	jand g155(.dina(w_n213_0[1]),.dinb(w_n205_0[0]),.dout(n214),.clk(gclk));
	jxor g156(.dina(w_n214_0[1]),.dinb(w_G125_0[0]),.dout(G27),.clk(gclk));
	jnot g157(.din(w_n96_0[0]),.dout(n216),.clk(gclk));
	jand g158(.dina(w_n108_0[1]),.dinb(w_n216_0[1]),.dout(n217),.clk(gclk));
	jand g159(.dina(w_n217_0[2]),.dinb(w_n122_0[1]),.dout(n218),.clk(gclk));
	jand g160(.dina(w_n218_1[1]),.dinb(w_n93_0[0]),.dout(n219),.clk(gclk));
	jand g161(.dina(w_n219_0[1]),.dinb(w_n193_0[0]),.dout(n220),.clk(gclk));
	jxor g162(.dina(w_n220_0[2]),.dinb(w_G131_0[0]),.dout(G33),.clk(gclk));
	jand g163(.dina(w_n219_0[0]),.dinb(w_n185_0[1]),.dout(n222),.clk(gclk));
	jxor g164(.dina(w_n222_0[2]),.dinb(w_G134_0[0]),.dout(G36),.clk(gclk));
	jand g165(.dina(w_n178_0[0]),.dinb(w_n156_1[0]),.dout(n224),.clk(gclk));
	jand g166(.dina(n224),.dinb(w_n184_0[2]),.dout(n225),.clk(gclk));
	jand g167(.dina(n225),.dinb(w_n218_1[0]),.dout(n226),.clk(gclk));
	jxor g168(.dina(w_n226_0[1]),.dinb(w_G137_0[0]),.dout(G39),.clk(gclk));
	jand g169(.dina(w_n218_0[2]),.dinb(w_n213_0[0]),.dout(n228),.clk(gclk));
	jxor g170(.dina(w_n228_0[1]),.dinb(w_G140_0[0]),.dout(G42),.clk(gclk));
	jcb g171(.dina(w_n203_0[0]),.dinb(w_n168_0[0]),.dout(n230));
	jcb g172(.dina(w_dff_B_SuaWyHO09_0),.dinb(w_n159_0[1]),.dout(n231));
	jcb g173(.dina(w_n201_0[0]),.dinb(w_n172_0[0]),.dout(n232));
	jcb g174(.dina(w_n211_0[0]),.dinb(w_n207_0[0]),.dout(n233));
	jcb g175(.dina(n233),.dinb(w_n176_0[0]),.dout(n234));
	jcb g176(.dina(n234),.dinb(w_dff_B_r8CDHUvp8_1),.dout(n235));
	jcb g177(.dina(n235),.dinb(n231),.dout(n236));
	jcb g178(.dina(w_n214_0[0]),.dinb(w_n191_0[0]),.dout(n237));
	jcb g179(.dina(n237),.dinb(w_n194_0[0]),.dout(n238));
	jcb g180(.dina(n238),.dinb(w_n222_0[1]),.dout(n239));
	jcb g181(.dina(w_n228_0[0]),.dinb(w_n226_0[0]),.dout(n240));
	jcb g182(.dina(w_n220_0[1]),.dinb(w_n186_0[0]),.dout(n241));
	jcb g183(.dina(w_dff_B_gpjAV2IP4_0),.dinb(n240),.dout(n242));
	jcb g184(.dina(n242),.dinb(n239),.dout(n243));
	jcb g185(.dina(n243),.dinb(w_n236_0[1]),.dout(n244));
	jxor g186(.dina(w_n121_0[0]),.dinb(w_n111_0[0]),.dout(n245),.clk(gclk));
	jand g187(.dina(n245),.dinb(w_n217_0[1]),.dout(n246),.clk(gclk));
	jcb g188(.dina(w_n92_0[2]),.dinb(w_n174_0[1]),.dout(n247));
	jnot g189(.din(w_n197_0[0]),.dout(n248),.clk(gclk));
	jxor g190(.dina(w_n108_0[0]),.dinb(w_n216_0[0]),.dout(n249),.clk(gclk));
	jand g191(.dina(w_dff_B_NjbvnhGJ3_0),.dinb(w_n248_0[1]),.dout(n250),.clk(gclk));
	jcb g192(.dina(n250),.dinb(w_n247_0[2]),.dout(n251));
	jcb g193(.dina(n251),.dinb(n246),.dout(n252));
	jcb g194(.dina(w_n162_0[1]),.dinb(w_n77_0[2]),.dout(n253));
	jand g195(.dina(w_n217_0[0]),.dinb(w_n248_0[0]),.dout(n254),.clk(gclk));
	jcb g196(.dina(w_n254_0[1]),.dinb(w_n163_0[2]),.dout(n255));
	jand g197(.dina(n255),.dinb(w_n253_1[1]),.dout(n256),.clk(gclk));
	jand g198(.dina(n256),.dinb(w_n156_0[2]),.dout(n257),.clk(gclk));
	jand g199(.dina(n257),.dinb(w_dff_B_MvrFUeGV0_1),.dout(n258),.clk(gclk));
	jand g200(.dina(w_n254_0[0]),.dinb(w_n163_0[1]),.dout(n259),.clk(gclk));
	jxor g201(.dina(w_n155_1[0]),.dinb(w_n144_0[2]),.dout(n260),.clk(gclk));
	jand g202(.dina(w_dff_B_ylgErEEf9_0),.dinb(w_n259_0[1]),.dout(n261),.clk(gclk));
	jcb g203(.dina(w_dff_B_8Jg4Dzxz2_0),.dinb(n258),.dout(n262));
	jand g204(.dina(n262),.dinb(w_n128_0[0]),.dout(n263),.clk(gclk));
	jcb g205(.dina(n263),.dinb(w_n244_2[2]),.dout(n264));
	jand g206(.dina(n264),.dinb(w_G952_0[1]),.dout(n265),.clk(gclk));
	jand g207(.dina(w_n259_0[0]),.dinb(w_n156_0[1]),.dout(n266),.clk(gclk));
	jcb g208(.dina(n266),.dinb(w_G953_1[2]),.dout(n267));
	jcb g209(.dina(w_dff_B_YKpfZl1u5_0),.dinb(n265),.dout(G75));
	jcb g210(.dina(w_n61_2[0]),.dinb(w_G952_0[0]),.dout(n269));
	jnot g211(.din(w_n105_0[0]),.dout(n270),.clk(gclk));
	jand g212(.dina(w_n244_2[1]),.dinb(w_G210_0[0]),.dout(n271),.clk(gclk));
	jand g213(.dina(n271),.dinb(w_G902_3[0]),.dout(n272),.clk(gclk));
	jxor g214(.dina(n272),.dinb(w_dff_B_Itw8uBOB2_1),.dout(n273),.clk(gclk));
	jand g215(.dina(n273),.dinb(w_n269_2[1]),.dout(G51),.clk(gclk));
	jand g216(.dina(w_G902_2[2]),.dinb(w_G469_0[0]),.dout(n275),.clk(gclk));
	jand g217(.dina(w_dff_B_zyjvtZ0X8_0),.dinb(w_n244_2[0]),.dout(n276),.clk(gclk));
	jxor g218(.dina(n276),.dinb(w_n119_0[0]),.dout(n277),.clk(gclk));
	jand g219(.dina(n277),.dinb(w_n269_2[0]),.dout(G54),.clk(gclk));
	jand g220(.dina(w_G902_2[1]),.dinb(w_G475_0[0]),.dout(n279),.clk(gclk));
	jand g221(.dina(w_n279_0[1]),.dinb(w_n244_1[2]),.dout(n280),.clk(gclk));
	jcb g222(.dina(n280),.dinb(w_n153_0[1]),.dout(n281));
	jnot g223(.din(w_n153_0[0]),.dout(n282),.clk(gclk));
	jnot g224(.din(w_n159_0[0]),.dout(n283),.clk(gclk));
	jnot g225(.din(w_n122_0[0]),.dout(n284),.clk(gclk));
	jcb g226(.dina(n284),.dinb(w_n109_0[0]),.dout(n285));
	jcb g227(.dina(w_n247_0[1]),.dinb(w_n285_1[1]),.dout(n286));
	jnot g228(.din(w_n167_0[0]),.dout(n287),.clk(gclk));
	jcb g229(.dina(w_n287_0[1]),.dinb(w_n286_0[1]),.dout(n288));
	jnot g230(.din(w_n171_0[0]),.dout(n289),.clk(gclk));
	jcb g231(.dina(w_n199_0[1]),.dinb(w_n289_0[1]),.dout(n290));
	jand g232(.dina(n290),.dinb(n288),.dout(n291),.clk(gclk));
	jand g233(.dina(w_dff_B_a5CkEPVo4_0),.dinb(n283),.dout(n292),.clk(gclk));
	jcb g234(.dina(w_n289_0[0]),.dinb(w_n286_0[0]),.dout(n293));
	jcb g235(.dina(w_n199_0[0]),.dinb(w_n287_0[0]),.dout(n294));
	jand g236(.dina(n294),.dinb(n293),.dout(n295),.clk(gclk));
	jnot g237(.din(w_n134_0[1]),.dout(n296),.clk(gclk));
	jcb g238(.dina(w_n165_0[0]),.dinb(w_n143_0[2]),.dout(n297));
	jcb g239(.dina(w_n297_0[1]),.dinb(w_n296_0[1]),.dout(n298));
	jcb g240(.dina(w_n298_0[1]),.dinb(w_n285_1[0]),.dout(n299));
	jcb g241(.dina(w_n92_0[1]),.dinb(w_n77_0[1]),.dout(n300));
	jcb g242(.dina(w_n300_0[1]),.dinb(n299),.dout(n301));
	jcb g243(.dina(w_n253_1[0]),.dinb(w_n298_0[0]),.dout(n302));
	jcb g244(.dina(n302),.dinb(w_n198_1[0]),.dout(n303));
	jcb g245(.dina(w_n155_0[2]),.dinb(w_n144_0[1]),.dout(n304));
	jcb g246(.dina(w_n247_0[0]),.dinb(w_n296_0[0]),.dout(n305));
	jcb g247(.dina(n305),.dinb(w_n304_0[1]),.dout(n306));
	jcb g248(.dina(n306),.dinb(w_n198_0[2]),.dout(n307));
	jand g249(.dina(n307),.dinb(n303),.dout(n308),.clk(gclk));
	jand g250(.dina(n308),.dinb(n301),.dout(n309),.clk(gclk));
	jand g251(.dina(w_dff_B_GAYwLA6H8_0),.dinb(n295),.dout(n310),.clk(gclk));
	jand g252(.dina(w_dff_B_vMa7JgJg5_0),.dinb(n292),.dout(n311),.clk(gclk));
	jnot g253(.din(w_n222_0[0]),.dout(n312),.clk(gclk));
	jcb g254(.dina(w_n253_0[2]),.dinb(w_n285_0[2]),.dout(n313));
	jcb g255(.dina(w_n155_0[1]),.dinb(w_n143_0[1]),.dout(n314));
	jnot g256(.din(w_n184_0[1]),.dout(n315),.clk(gclk));
	jcb g257(.dina(w_n315_0[2]),.dinb(n314),.dout(n316));
	jcb g258(.dina(w_n316_0[1]),.dinb(w_n313_0[1]),.dout(n317));
	jcb g259(.dina(w_n304_0[0]),.dinb(w_n196_0[0]),.dout(n318));
	jcb g260(.dina(n318),.dinb(w_n315_0[1]),.dout(n319));
	jcb g261(.dina(w_dff_B_p6TVTbM01_0),.dinb(w_n285_0[1]),.dout(n320));
	jcb g262(.dina(w_n316_0[0]),.dinb(w_n300_0[0]),.dout(n321));
	jcb g263(.dina(w_n321_0[1]),.dinb(w_n198_0[1]),.dout(n322));
	jand g264(.dina(w_dff_B_mYZ6SdKZ6_0),.dinb(n320),.dout(n323),.clk(gclk));
	jand g265(.dina(n323),.dinb(w_dff_B_d4MGz1xW8_1),.dout(n324),.clk(gclk));
	jand g266(.dina(w_dff_B_n6HfhzeT0_0),.dinb(n312),.dout(n325),.clk(gclk));
	jnot g267(.din(w_n218_0[1]),.dout(n326),.clk(gclk));
	jcb g268(.dina(w_n253_0[1]),.dinb(w_n297_0[0]),.dout(n327));
	jcb g269(.dina(n327),.dinb(w_n315_0[0]),.dout(n328));
	jcb g270(.dina(w_dff_B_pJ5gaPhu0_0),.dinb(w_n326_0[1]),.dout(n329));
	jcb g271(.dina(w_n326_0[0]),.dinb(w_n321_0[0]),.dout(n330));
	jand g272(.dina(n330),.dinb(n329),.dout(n331),.clk(gclk));
	jnot g273(.din(w_n185_0[0]),.dout(n332),.clk(gclk));
	jcb g274(.dina(n332),.dinb(w_n313_0[0]),.dout(n333));
	jnot g275(.din(w_n220_0[0]),.dout(n334),.clk(gclk));
	jand g276(.dina(n334),.dinb(w_dff_B_ezAnpGU13_1),.dout(n335),.clk(gclk));
	jand g277(.dina(n335),.dinb(w_dff_B_aiRoMdoG5_1),.dout(n336),.clk(gclk));
	jand g278(.dina(n336),.dinb(w_dff_B_YHUknnpY0_1),.dout(n337),.clk(gclk));
	jand g279(.dina(w_n337_0[1]),.dinb(w_n311_0[1]),.dout(n338),.clk(gclk));
	jnot g280(.din(w_n279_0[0]),.dout(n339),.clk(gclk));
	jcb g281(.dina(w_dff_B_2xASnDVr2_0),.dinb(w_n338_0[1]),.dout(n340));
	jcb g282(.dina(n340),.dinb(w_dff_B_p4MO3Bt46_1),.dout(n341));
	jand g283(.dina(n341),.dinb(w_n269_1[2]),.dout(n342),.clk(gclk));
	jand g284(.dina(n342),.dinb(w_dff_B_GxLZSbNy4_1),.dout(G60),.clk(gclk));
	jand g285(.dina(w_G902_2[0]),.dinb(w_G478_0[0]),.dout(n344),.clk(gclk));
	jand g286(.dina(w_n344_0[1]),.dinb(w_n244_1[1]),.dout(n345),.clk(gclk));
	jcb g287(.dina(n345),.dinb(w_n141_0[1]),.dout(n346));
	jnot g288(.din(w_n141_0[0]),.dout(n347),.clk(gclk));
	jnot g289(.din(w_n344_0[0]),.dout(n348),.clk(gclk));
	jcb g290(.dina(w_dff_B_ZOgbkHDb3_0),.dinb(w_n338_0[0]),.dout(n349));
	jcb g291(.dina(n349),.dinb(w_dff_B_OaMo6QT61_1),.dout(n350));
	jand g292(.dina(n350),.dinb(w_n269_1[1]),.dout(n351),.clk(gclk));
	jand g293(.dina(n351),.dinb(w_dff_B_dCMRLTmz6_1),.dout(G63),.clk(gclk));
	jand g294(.dina(w_n244_1[0]),.dinb(w_G217_0[0]),.dout(n353),.clk(gclk));
	jand g295(.dina(n353),.dinb(w_G902_1[2]),.dout(n354),.clk(gclk));
	jxor g296(.dina(n354),.dinb(w_n71_0[0]),.dout(n355),.clk(gclk));
	jand g297(.dina(n355),.dinb(w_n269_1[0]),.dout(G66),.clk(gclk));
	jcb g298(.dina(w_n311_0[0]),.dinb(w_G953_1[1]),.dout(n357));
	jcb g299(.dina(n357),.dinb(w_n101_0[1]),.dout(n358));
	jand g300(.dina(w_n236_0[0]),.dinb(w_n61_1[2]),.dout(n359),.clk(gclk));
	jnot g301(.din(w_n101_0[0]),.dout(n360),.clk(gclk));
	jcb g302(.dina(w_n131_0[0]),.dinb(n360),.dout(n361));
	jcb g303(.dina(w_dff_B_0KQt4l9f1_0),.dinb(n359),.dout(n362));
	jand g304(.dina(w_dff_B_lyofbDAS1_0),.dinb(n358),.dout(n363),.clk(gclk));
	jand g305(.dina(w_G898_0[0]),.dinb(w_G224_0[0]),.dout(n364),.clk(gclk));
	jcb g306(.dina(n364),.dinb(w_n61_1[1]),.dout(n365));
	jxor g307(.dina(w_dff_B_Y0kMxlKp3_0),.dinb(n363),.dout(G69),.clk(gclk));
	jcb g308(.dina(w_n337_0[0]),.dinb(w_G953_1[0]),.dout(n367));
	jand g309(.dina(w_G900_0[0]),.dinb(w_G227_0[0]),.dout(n368),.clk(gclk));
	jcb g310(.dina(n368),.dinb(w_n61_1[0]),.dout(n369));
	jand g311(.dina(w_dff_B_ETtamJp77_0),.dinb(n367),.dout(n370),.clk(gclk));
	jxor g312(.dina(w_n82_0[0]),.dinb(w_n65_0[0]),.dout(n371),.clk(gclk));
	jcb g313(.dina(n371),.dinb(w_n181_0[0]),.dout(n372));
	jxor g314(.dina(w_dff_B_I03464Z71_0),.dinb(n370),.dout(G72),.clk(gclk));
	jand g315(.dina(w_n244_0[2]),.dinb(w_G472_0[0]),.dout(n374),.clk(gclk));
	jand g316(.dina(n374),.dinb(w_G902_1[1]),.dout(n375),.clk(gclk));
	jxor g317(.dina(n375),.dinb(w_n90_0[0]),.dout(n376),.clk(gclk));
	jand g318(.dina(n376),.dinb(w_n269_0[2]),.dout(G57),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_dff_A_vhETZMxO6_0),.doutb(w_G101_0[1]),.doutc(w_dff_A_FtYLZEww0_2),.din(w_dff_B_y2ks6dKP9_3));
	jspl3 jspl3_w_G104_0(.douta(w_dff_A_ryt0mnN75_0),.doutb(w_dff_A_NC3t7dCW0_1),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_dff_A_mvQDJjhl0_0),.doutb(w_dff_A_lFGwgagg5_1),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_dff_A_yilBa07N3_0),.doutb(w_G110_0[1]),.doutc(w_G110_0[2]),.din(G110));
	jspl3 jspl3_w_G113_0(.douta(w_dff_A_BKpryq4U4_0),.doutb(w_G113_0[1]),.doutc(w_dff_A_ZLODwrnj3_2),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_dff_A_MS1gN8KP4_0),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_dff_A_mF7KzgY93_0),.doutb(w_G119_0[1]),.doutc(w_dff_A_SJxdXh8r0_2),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_dff_A_pYAaDC458_1),.doutc(w_G122_0[2]),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_dff_A_Ui9PJ5O17_1),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_dff_A_hAbroMB57_0),.doutb(w_dff_A_AcWRQco98_1),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_dff_A_Uohm0taf4_0),.doutb(w_G128_0[1]),.doutc(w_dff_A_G3lp0cUe0_2),.din(G128));
	jspl3 jspl3_w_G131_0(.douta(w_dff_A_kBvrLY7q2_0),.doutb(w_G131_0[1]),.doutc(w_dff_A_iuCcpqQN4_2),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_dff_A_3HnYfHIg9_0),.doutb(w_dff_A_LZJINklu6_1),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_iKE1LC3X9_0),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G140_0(.douta(w_dff_A_IsyiABwm5_0),.doutb(w_G140_0[1]),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_dff_A_GApTDjgN1_0),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(G143));
	jspl3 jspl3_w_G146_0(.douta(w_dff_A_GFIt6KrB0_0),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(w_dff_B_V41iQZ8u6_3));
	jspl3 jspl3_w_G210_0(.douta(w_dff_A_u0r9HC9p1_0),.doutb(w_dff_A_cSU03OiF5_1),.doutc(w_G210_0[2]),.din(w_dff_B_5KcbtH9R0_3));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_dff_A_npsImUZ42_1),.din(w_dff_B_VME5RSDq1_2));
	jspl3 jspl3_w_G217_0(.douta(w_dff_A_Gw1p1y5E4_0),.doutb(w_G217_0[1]),.doutc(w_dff_A_gdmvXRrI7_2),.din(G217));
	jspl jspl_w_G221_0(.douta(w_dff_A_ni3v0n9z5_0),.doutb(w_G221_0[1]),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_dff_A_U2ppfvjE4_1),.din(G224));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_G227_0[1]),.din(G227));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_G234_0[2]),.din(G234));
	jspl jspl_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.din(w_G234_0[0]));
	jspl jspl_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.din(G237));
	jspl jspl_w_G469_0(.douta(w_G469_0[0]),.doutb(w_dff_A_TJQ3WB8z4_1),.din(G469));
	jspl3 jspl3_w_G472_0(.douta(w_dff_A_FU9JAAiV3_0),.doutb(w_G472_0[1]),.doutc(w_dff_A_ICOXnSjx7_2),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_dff_A_tKNjPyhs0_1),.doutc(w_G475_0[2]),.din(G475));
	jspl jspl_w_G478_0(.douta(w_G478_0[0]),.doutb(w_dff_A_FHA5ViFc5_1),.din(G478));
	jspl jspl_w_G898_0(.douta(w_G898_0[0]),.doutb(w_G898_0[1]),.din(G898));
	jspl jspl_w_G900_0(.douta(w_G900_0[0]),.doutb(w_G900_0[1]),.din(G900));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_dff_A_kyALfS8y8_2),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_dff_A_ZwwODbhB0_1),.doutc(w_dff_A_w6irMycR8_2),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_G902_2[1]),.doutc(w_G902_2[2]),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_dff_A_C1oU3Xa71_0),.doutb(w_G902_3[1]),.doutc(w_G902_3[2]),.din(w_G902_0[2]));
	jspl3 jspl3_w_G902_4(.douta(w_dff_A_hC6Riofy9_0),.doutb(w_dff_A_EenXafGX8_1),.doutc(w_G902_4[2]),.din(w_G902_1[0]));
	jspl3 jspl3_w_G952_0(.douta(w_dff_A_NFSuWSaA9_0),.doutb(w_dff_A_lX7bwFbg2_1),.doutc(w_G952_0[2]),.din(G952));
	jspl3 jspl3_w_G953_0(.douta(w_dff_A_YmhNpf6I9_0),.doutb(w_dff_A_qLXv9ayE6_1),.doutc(w_G953_0[2]),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_dff_A_xqMIXTHk3_0),.doutb(w_dff_A_PHOxtYAj4_1),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl3 jspl3_w_G953_2(.douta(w_G953_2[0]),.doutb(w_G953_2[1]),.doutc(w_G953_2[2]),.din(w_G953_0[1]));
	jspl jspl_w_G953_3(.douta(w_dff_A_PhPMIR101_0),.doutb(w_G953_3[1]),.din(w_G953_0[2]));
	jspl3 jspl3_w_n59_0(.douta(w_n59_0[0]),.doutb(w_dff_A_1o9DG4HD1_1),.doutc(w_dff_A_SmRkh54p1_2),.din(n59));
	jspl3 jspl3_w_n59_1(.douta(w_dff_A_Q2jMbFOm1_0),.doutb(w_dff_A_pudfbXUd3_1),.doutc(w_n59_1[2]),.din(w_n59_0[0]));
	jspl jspl_w_n59_2(.douta(w_dff_A_tREwYbIJ1_0),.doutb(w_n59_2[1]),.din(w_n59_0[1]));
	jspl3 jspl3_w_n61_0(.douta(w_n61_0[0]),.doutb(w_n61_0[1]),.doutc(w_n61_0[2]),.din(n61));
	jspl3 jspl3_w_n61_1(.douta(w_n61_1[0]),.doutb(w_n61_1[1]),.doutc(w_dff_A_m6tq2qpa7_2),.din(w_n61_0[0]));
	jspl3 jspl3_w_n61_2(.douta(w_n61_2[0]),.doutb(w_n61_2[1]),.doutc(w_n61_2[2]),.din(w_n61_0[1]));
	jspl3 jspl3_w_n61_3(.douta(w_n61_3[0]),.doutb(w_n61_3[1]),.doutc(w_n61_3[2]),.din(w_n61_0[2]));
	jspl jspl_w_n65_0(.douta(w_dff_A_K3IqHHkr1_0),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n66_0(.douta(w_dff_A_APhnHAiT2_0),.doutb(w_n66_0[1]),.din(w_dff_B_iPWazfDc1_2));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n71_0(.douta(w_dff_A_Pnv99A6v3_0),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n72_0(.douta(w_n72_0[0]),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.din(n74));
	jspl jspl_w_n75_0(.douta(w_dff_A_Gxhitpy44_0),.doutb(w_n75_0[1]),.din(n75));
	jspl3 jspl3_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.doutc(w_n77_0[2]),.din(w_dff_B_gC6kq2403_3));
	jspl jspl_w_n77_1(.douta(w_n77_1[0]),.doutb(w_n77_1[1]),.din(w_n77_0[0]));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.din(n79));
	jspl3 jspl3_w_n82_0(.douta(w_n82_0[0]),.doutb(w_n82_0[1]),.doutc(w_dff_A_FWBvyt5U0_2),.din(n82));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_dff_A_OwpnqkYD3_1),.din(n84));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_2RV8VcwV1_0),.doutb(w_n85_0[1]),.doutc(w_dff_A_KrZ6EOnd6_2),.din(n85));
	jspl jspl_w_n90_0(.douta(w_dff_A_MXEDLgJw5_0),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.din(n91));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n92_1(.douta(w_n92_1[0]),.doutb(w_n92_1[1]),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_dff_A_giDHr2hO0_2),.din(n93));
	jspl jspl_w_n95_0(.douta(w_n95_0[0]),.doutb(w_n95_0[1]),.din(n95));
	jspl jspl_w_n96_0(.douta(w_n96_0[0]),.doutb(w_dff_A_BSyXgYxY5_1),.din(n96));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl3 jspl3_w_n101_0(.douta(w_n101_0[0]),.doutb(w_dff_A_U2HY2R2g0_1),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n105_0(.douta(w_n105_0[0]),.doutb(w_n105_0[1]),.din(n105));
	jspl3 jspl3_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.doutc(w_n108_0[2]),.din(n108));
	jspl3 jspl3_w_n109_0(.douta(w_dff_A_xzHN8wSu2_0),.doutb(w_dff_A_tq3evxCx6_1),.doutc(w_n109_0[2]),.din(n109));
	jspl3 jspl3_w_n111_0(.douta(w_dff_A_HcECIPF01_0),.doutb(w_dff_A_P6dePn5q4_1),.doutc(w_n111_0[2]),.din(n111));
	jspl jspl_w_n119_0(.douta(w_dff_A_inAgN7b92_0),.doutb(w_n119_0[1]),.din(n119));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.doutc(w_n122_0[2]),.din(n122));
	jspl3 jspl3_w_n123_0(.douta(w_n123_0[0]),.doutb(w_dff_A_StFfRhm90_1),.doutc(w_n123_0[2]),.din(n123));
	jspl jspl_w_n123_1(.douta(w_n123_1[0]),.doutb(w_dff_A_2NVq1sYn1_1),.din(w_n123_0[0]));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl3 jspl3_w_n128_0(.douta(w_dff_A_SvLAo0DM1_0),.doutb(w_n128_0[1]),.doutc(w_n128_0[2]),.din(w_dff_B_dJQNrJGn0_3));
	jspl jspl_w_n129_0(.douta(w_n129_0[0]),.doutb(w_n129_0[1]),.din(w_dff_B_IUWquhTG7_2));
	jspl jspl_w_n131_0(.douta(w_dff_A_zEL2RL1p2_0),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n134_0(.douta(w_dff_A_AccwtbgX6_0),.doutb(w_n134_0[1]),.doutc(w_dff_A_d3Ly3WpX8_2),.din(n134));
	jspl3 jspl3_w_n134_1(.douta(w_n134_1[0]),.doutb(w_n134_1[1]),.doutc(w_n134_1[2]),.din(w_n134_0[0]));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_dff_A_cvJ4WcHM2_1),.doutc(w_n141_0[2]),.din(n141));
	jspl3 jspl3_w_n143_0(.douta(w_n143_0[0]),.doutb(w_dff_A_P18OMZwK3_1),.doutc(w_dff_A_jA8P3gX08_2),.din(n143));
	jspl3 jspl3_w_n143_1(.douta(w_dff_A_r3KvVKkS4_0),.doutb(w_dff_A_0l7TO2iJ5_1),.doutc(w_n143_1[2]),.din(w_n143_0[0]));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.doutc(w_n144_0[2]),.din(w_dff_B_sFbHan702_3));
	jspl jspl_w_n144_1(.douta(w_n144_1[0]),.doutb(w_n144_1[1]),.din(w_n144_0[0]));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_dff_A_wyUeuZlK6_1),.doutc(w_n153_0[2]),.din(n153));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(n154));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl3 jspl3_w_n155_1(.douta(w_n155_1[0]),.doutb(w_n155_1[1]),.doutc(w_n155_1[2]),.din(w_n155_0[0]));
	jspl3 jspl3_w_n156_0(.douta(w_n156_0[0]),.doutb(w_dff_A_tlUmzFcf7_1),.doutc(w_dff_A_WnJsyQ5g5_2),.din(n156));
	jspl jspl_w_n156_1(.douta(w_n156_1[0]),.doutb(w_n156_1[1]),.din(w_n156_0[0]));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(n158));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl3 jspl3_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.doutc(w_n162_0[2]),.din(n162));
	jspl jspl_w_n162_1(.douta(w_n162_1[0]),.doutb(w_n162_1[1]),.din(w_n162_0[0]));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_n163_0[2]),.din(n163));
	jspl jspl_w_n163_1(.douta(w_n163_1[0]),.doutb(w_n163_1[1]),.din(w_n163_0[0]));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.doutc(w_n165_0[2]),.din(n165));
	jspl jspl_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.din(n166));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.doutc(w_n167_0[2]),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(n170));
	jspl3 jspl3_w_n171_0(.douta(w_n171_0[0]),.doutb(w_n171_0[1]),.doutc(w_n171_0[2]),.din(n171));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl3 jspl3_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.doutc(w_n174_0[2]),.din(w_dff_B_UYS0eS4J9_3));
	jspl jspl_w_n174_1(.douta(w_n174_1[0]),.doutb(w_n174_1[1]),.din(w_n174_0[0]));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_dff_A_FKwiEQCc1_1),.din(w_dff_B_38toSO1e7_2));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl3 jspl3_w_n178_0(.douta(w_n178_0[0]),.doutb(w_dff_A_CKNJDBMO5_1),.doutc(w_n178_0[2]),.din(n178));
	jspl jspl_w_n179_0(.douta(w_n179_0[0]),.doutb(w_n179_0[1]),.din(n179));
	jspl jspl_w_n181_0(.douta(w_dff_A_6GvLxx1O3_0),.doutb(w_n181_0[1]),.din(n181));
	jspl3 jspl3_w_n184_0(.douta(w_dff_A_lJgjFNBv1_0),.doutb(w_n184_0[1]),.doutc(w_dff_A_JH7mNzYY0_2),.din(n184));
	jspl3 jspl3_w_n184_1(.douta(w_n184_1[0]),.doutb(w_dff_A_ALQxHeVA9_1),.doutc(w_n184_1[2]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.doutc(w_n185_0[2]),.din(n185));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n188_0(.douta(w_dff_A_DSmlpsRc5_0),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.din(n191));
	jspl3 jspl3_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.doutc(w_n193_0[2]),.din(n193));
	jspl jspl_w_n194_0(.douta(w_dff_A_yMeXOukv4_0),.doutb(w_n194_0[1]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.din(n196));
	jspl jspl_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.din(n197));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_dff_A_I1kg5hwF5_1),.doutc(w_dff_A_TmbHF47T2_2),.din(n198));
	jspl3 jspl3_w_n198_1(.douta(w_dff_A_Clk3MhQA4_0),.doutb(w_n198_1[1]),.doutc(w_dff_A_f7ZbnAm77_2),.din(w_n198_0[0]));
	jspl3 jspl3_w_n199_0(.douta(w_dff_A_zLjQ5DjK5_0),.doutb(w_dff_A_A5IuR94N6_1),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(w_dff_B_POD5FexQ7_2));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(n203));
	jspl3 jspl3_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.doutc(w_n205_0[2]),.din(w_dff_B_FjK7oy4T4_3));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.din(n211));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl jspl_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.din(n214));
	jspl jspl_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.din(w_dff_B_vwyHxJUz9_2));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(w_dff_B_TdvY5iUP8_3));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_dff_A_cOP0zIfQ1_2),.din(n218));
	jspl jspl_w_n218_1(.douta(w_dff_A_saCiEqOW4_0),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl3 jspl3_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.doutc(w_n220_0[2]),.din(n220));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_dff_A_kiesjfqD5_1),.doutc(w_n222_0[2]),.din(n222));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.din(n236));
	jspl3 jspl3_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.doutc(w_n244_0[2]),.din(n244));
	jspl3 jspl3_w_n244_1(.douta(w_n244_1[0]),.doutb(w_n244_1[1]),.doutc(w_n244_1[2]),.din(w_n244_0[0]));
	jspl3 jspl3_w_n244_2(.douta(w_n244_2[0]),.doutb(w_n244_2[1]),.doutc(w_dff_A_4JaeotOm3_2),.din(w_n244_0[1]));
	jspl3 jspl3_w_n247_0(.douta(w_n247_0[0]),.doutb(w_dff_A_lCyFUNZz8_1),.doutc(w_dff_A_iwoknT9B4_2),.din(n247));
	jspl jspl_w_n248_0(.douta(w_n248_0[0]),.doutb(w_n248_0[1]),.din(n248));
	jspl3 jspl3_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.doutc(w_dff_A_E873VoV34_2),.din(n253));
	jspl jspl_w_n253_1(.douta(w_n253_1[0]),.doutb(w_dff_A_mOAYSE0e8_1),.din(w_n253_0[0]));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl3 jspl3_w_n269_0(.douta(w_dff_A_S93cdf7v1_0),.doutb(w_n269_0[1]),.doutc(w_dff_A_T6QzBcsh7_2),.din(w_dff_B_xMgHvZ9D3_3));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_dff_A_fSftLx0k0_1),.doutc(w_dff_A_wQFJnKsT9_2),.din(w_n269_0[0]));
	jspl jspl_w_n269_2(.douta(w_n269_2[0]),.doutb(w_dff_A_fvTFRsyf6_1),.din(w_n269_0[1]));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_dff_A_fIkK8fy79_1),.din(n279));
	jspl3 jspl3_w_n285_0(.douta(w_n285_0[0]),.doutb(w_n285_0[1]),.doutc(w_n285_0[2]),.din(n285));
	jspl jspl_w_n285_1(.douta(w_n285_1[0]),.doutb(w_n285_1[1]),.din(w_n285_0[0]));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(w_dff_B_Sk0MnWd06_2));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl jspl_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.din(n289));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(w_dff_B_juXlPDi56_2));
	jspl jspl_w_n297_0(.douta(w_n297_0[0]),.doutb(w_n297_0[1]),.din(n297));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_dff_A_WePsK7ok3_1),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_dff_A_QbYjEiid8_1),.din(n300));
	jspl jspl_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.din(n304));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n313_0(.douta(w_dff_A_C1rSbdtx0_0),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.doutc(w_n315_0[2]),.din(w_dff_B_BVBFn80e3_3));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_dff_A_xnd6brWN0_1),.din(n316));
	jspl jspl_w_n321_0(.douta(w_dff_A_kzyFlC3Z5_0),.doutb(w_n321_0[1]),.din(n321));
	jspl jspl_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.din(n326));
	jspl jspl_w_n337_0(.douta(w_n337_0[0]),.doutb(w_n337_0[1]),.din(n337));
	jspl jspl_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.din(n338));
	jspl jspl_w_n344_0(.douta(w_n344_0[0]),.doutb(w_dff_A_7OdfY3Yh9_1),.din(n344));
	jdff dff_B_Dk4nmQs10_0(.din(n267),.dout(w_dff_B_Dk4nmQs10_0),.clk(gclk));
	jdff dff_B_OiV1sQ5l7_0(.din(w_dff_B_Dk4nmQs10_0),.dout(w_dff_B_OiV1sQ5l7_0),.clk(gclk));
	jdff dff_B_YKpfZl1u5_0(.din(w_dff_B_OiV1sQ5l7_0),.dout(w_dff_B_YKpfZl1u5_0),.clk(gclk));
	jdff dff_B_8Jg4Dzxz2_0(.din(n261),.dout(w_dff_B_8Jg4Dzxz2_0),.clk(gclk));
	jdff dff_B_ylgErEEf9_0(.din(n260),.dout(w_dff_B_ylgErEEf9_0),.clk(gclk));
	jdff dff_B_6gIYyRZb2_1(.din(n252),.dout(w_dff_B_6gIYyRZb2_1),.clk(gclk));
	jdff dff_B_MvrFUeGV0_1(.din(w_dff_B_6gIYyRZb2_1),.dout(w_dff_B_MvrFUeGV0_1),.clk(gclk));
	jdff dff_B_NjbvnhGJ3_0(.din(n249),.dout(w_dff_B_NjbvnhGJ3_0),.clk(gclk));
	jdff dff_B_em63zvdk5_1(.din(n270),.dout(w_dff_B_em63zvdk5_1),.clk(gclk));
	jdff dff_B_UY0HwHku7_1(.din(w_dff_B_em63zvdk5_1),.dout(w_dff_B_UY0HwHku7_1),.clk(gclk));
	jdff dff_B_U3De3fb42_1(.din(w_dff_B_UY0HwHku7_1),.dout(w_dff_B_U3De3fb42_1),.clk(gclk));
	jdff dff_B_kX2MOGrI8_1(.din(w_dff_B_U3De3fb42_1),.dout(w_dff_B_kX2MOGrI8_1),.clk(gclk));
	jdff dff_B_kXXFVEmg9_1(.din(w_dff_B_kX2MOGrI8_1),.dout(w_dff_B_kXXFVEmg9_1),.clk(gclk));
	jdff dff_B_QjdjnfdV3_1(.din(w_dff_B_kXXFVEmg9_1),.dout(w_dff_B_QjdjnfdV3_1),.clk(gclk));
	jdff dff_B_T2VrmKJn9_1(.din(w_dff_B_QjdjnfdV3_1),.dout(w_dff_B_T2VrmKJn9_1),.clk(gclk));
	jdff dff_B_Itw8uBOB2_1(.din(w_dff_B_T2VrmKJn9_1),.dout(w_dff_B_Itw8uBOB2_1),.clk(gclk));
	jdff dff_B_gAJeyiaM8_0(.din(n275),.dout(w_dff_B_gAJeyiaM8_0),.clk(gclk));
	jdff dff_B_PcbmW6ZI7_0(.din(w_dff_B_gAJeyiaM8_0),.dout(w_dff_B_PcbmW6ZI7_0),.clk(gclk));
	jdff dff_B_UK4GJsiV3_0(.din(w_dff_B_PcbmW6ZI7_0),.dout(w_dff_B_UK4GJsiV3_0),.clk(gclk));
	jdff dff_B_p8xDgMib8_0(.din(w_dff_B_UK4GJsiV3_0),.dout(w_dff_B_p8xDgMib8_0),.clk(gclk));
	jdff dff_B_rd6nBQVs2_0(.din(w_dff_B_p8xDgMib8_0),.dout(w_dff_B_rd6nBQVs2_0),.clk(gclk));
	jdff dff_B_n697LSWx5_0(.din(w_dff_B_rd6nBQVs2_0),.dout(w_dff_B_n697LSWx5_0),.clk(gclk));
	jdff dff_B_EB4LNcGZ2_0(.din(w_dff_B_n697LSWx5_0),.dout(w_dff_B_EB4LNcGZ2_0),.clk(gclk));
	jdff dff_B_ts2CxtsM2_0(.din(w_dff_B_EB4LNcGZ2_0),.dout(w_dff_B_ts2CxtsM2_0),.clk(gclk));
	jdff dff_B_BoWr6wRo6_0(.din(w_dff_B_ts2CxtsM2_0),.dout(w_dff_B_BoWr6wRo6_0),.clk(gclk));
	jdff dff_B_BWu6umMX5_0(.din(w_dff_B_BoWr6wRo6_0),.dout(w_dff_B_BWu6umMX5_0),.clk(gclk));
	jdff dff_B_zyjvtZ0X8_0(.din(w_dff_B_BWu6umMX5_0),.dout(w_dff_B_zyjvtZ0X8_0),.clk(gclk));
	jdff dff_A_4JaeotOm3_2(.dout(w_n244_2[2]),.din(w_dff_A_4JaeotOm3_2),.clk(gclk));
	jdff dff_A_fvTFRsyf6_1(.dout(w_n269_2[1]),.din(w_dff_A_fvTFRsyf6_1),.clk(gclk));
	jdff dff_B_ff8Q1GrI0_1(.din(n281),.dout(w_dff_B_ff8Q1GrI0_1),.clk(gclk));
	jdff dff_B_03te53yw1_1(.din(w_dff_B_ff8Q1GrI0_1),.dout(w_dff_B_03te53yw1_1),.clk(gclk));
	jdff dff_B_GoxgVuQm1_1(.din(w_dff_B_03te53yw1_1),.dout(w_dff_B_GoxgVuQm1_1),.clk(gclk));
	jdff dff_B_GxLZSbNy4_1(.din(w_dff_B_GoxgVuQm1_1),.dout(w_dff_B_GxLZSbNy4_1),.clk(gclk));
	jdff dff_B_DaoqrbUh7_1(.din(n282),.dout(w_dff_B_DaoqrbUh7_1),.clk(gclk));
	jdff dff_B_Kk1z713U8_1(.din(w_dff_B_DaoqrbUh7_1),.dout(w_dff_B_Kk1z713U8_1),.clk(gclk));
	jdff dff_B_c92ERZF98_1(.din(w_dff_B_Kk1z713U8_1),.dout(w_dff_B_c92ERZF98_1),.clk(gclk));
	jdff dff_B_9PlWo8jR6_1(.din(w_dff_B_c92ERZF98_1),.dout(w_dff_B_9PlWo8jR6_1),.clk(gclk));
	jdff dff_B_Y0mwXCeU4_1(.din(w_dff_B_9PlWo8jR6_1),.dout(w_dff_B_Y0mwXCeU4_1),.clk(gclk));
	jdff dff_B_XBJ5yhqs2_1(.din(w_dff_B_Y0mwXCeU4_1),.dout(w_dff_B_XBJ5yhqs2_1),.clk(gclk));
	jdff dff_B_gxavRIm69_1(.din(w_dff_B_XBJ5yhqs2_1),.dout(w_dff_B_gxavRIm69_1),.clk(gclk));
	jdff dff_B_c0jutqYs8_1(.din(w_dff_B_gxavRIm69_1),.dout(w_dff_B_c0jutqYs8_1),.clk(gclk));
	jdff dff_B_p4MO3Bt46_1(.din(w_dff_B_c0jutqYs8_1),.dout(w_dff_B_p4MO3Bt46_1),.clk(gclk));
	jdff dff_B_WUCWDsxf3_0(.din(n339),.dout(w_dff_B_WUCWDsxf3_0),.clk(gclk));
	jdff dff_B_uSENDypd6_0(.din(w_dff_B_WUCWDsxf3_0),.dout(w_dff_B_uSENDypd6_0),.clk(gclk));
	jdff dff_B_2RNIIohY6_0(.din(w_dff_B_uSENDypd6_0),.dout(w_dff_B_2RNIIohY6_0),.clk(gclk));
	jdff dff_B_cVyJoijz4_0(.din(w_dff_B_2RNIIohY6_0),.dout(w_dff_B_cVyJoijz4_0),.clk(gclk));
	jdff dff_B_kQZEMinE7_0(.din(w_dff_B_cVyJoijz4_0),.dout(w_dff_B_kQZEMinE7_0),.clk(gclk));
	jdff dff_B_g2FPmPs22_0(.din(w_dff_B_kQZEMinE7_0),.dout(w_dff_B_g2FPmPs22_0),.clk(gclk));
	jdff dff_B_ou9mg8HE5_0(.din(w_dff_B_g2FPmPs22_0),.dout(w_dff_B_ou9mg8HE5_0),.clk(gclk));
	jdff dff_B_rG9sL0fK0_0(.din(w_dff_B_ou9mg8HE5_0),.dout(w_dff_B_rG9sL0fK0_0),.clk(gclk));
	jdff dff_B_7xA612sE3_0(.din(w_dff_B_rG9sL0fK0_0),.dout(w_dff_B_7xA612sE3_0),.clk(gclk));
	jdff dff_B_WyNOZNnZ1_0(.din(w_dff_B_7xA612sE3_0),.dout(w_dff_B_WyNOZNnZ1_0),.clk(gclk));
	jdff dff_B_c08gOoFP3_0(.din(w_dff_B_WyNOZNnZ1_0),.dout(w_dff_B_c08gOoFP3_0),.clk(gclk));
	jdff dff_B_BtoisHfb7_0(.din(w_dff_B_c08gOoFP3_0),.dout(w_dff_B_BtoisHfb7_0),.clk(gclk));
	jdff dff_B_zrMQXsVj2_0(.din(w_dff_B_BtoisHfb7_0),.dout(w_dff_B_zrMQXsVj2_0),.clk(gclk));
	jdff dff_B_2xASnDVr2_0(.din(w_dff_B_zrMQXsVj2_0),.dout(w_dff_B_2xASnDVr2_0),.clk(gclk));
	jdff dff_A_EcL0WOZG5_1(.dout(w_n279_0[1]),.din(w_dff_A_EcL0WOZG5_1),.clk(gclk));
	jdff dff_A_sEPJfhib7_1(.dout(w_dff_A_EcL0WOZG5_1),.din(w_dff_A_sEPJfhib7_1),.clk(gclk));
	jdff dff_A_rlZF7qFx8_1(.dout(w_dff_A_sEPJfhib7_1),.din(w_dff_A_rlZF7qFx8_1),.clk(gclk));
	jdff dff_A_wxdIY6kZ7_1(.dout(w_dff_A_rlZF7qFx8_1),.din(w_dff_A_wxdIY6kZ7_1),.clk(gclk));
	jdff dff_A_kUl6HOYn4_1(.dout(w_dff_A_wxdIY6kZ7_1),.din(w_dff_A_kUl6HOYn4_1),.clk(gclk));
	jdff dff_A_PYfon3DB3_1(.dout(w_dff_A_kUl6HOYn4_1),.din(w_dff_A_PYfon3DB3_1),.clk(gclk));
	jdff dff_A_ibeh9fBD5_1(.dout(w_dff_A_PYfon3DB3_1),.din(w_dff_A_ibeh9fBD5_1),.clk(gclk));
	jdff dff_A_eFB6ihZF5_1(.dout(w_dff_A_ibeh9fBD5_1),.din(w_dff_A_eFB6ihZF5_1),.clk(gclk));
	jdff dff_A_UHepSLeq9_1(.dout(w_dff_A_eFB6ihZF5_1),.din(w_dff_A_UHepSLeq9_1),.clk(gclk));
	jdff dff_A_Kfqyqo8a0_1(.dout(w_dff_A_UHepSLeq9_1),.din(w_dff_A_Kfqyqo8a0_1),.clk(gclk));
	jdff dff_A_fIkK8fy79_1(.dout(w_dff_A_Kfqyqo8a0_1),.din(w_dff_A_fIkK8fy79_1),.clk(gclk));
	jdff dff_B_8fBUTVCq5_1(.din(n346),.dout(w_dff_B_8fBUTVCq5_1),.clk(gclk));
	jdff dff_B_W3BUisI20_1(.din(w_dff_B_8fBUTVCq5_1),.dout(w_dff_B_W3BUisI20_1),.clk(gclk));
	jdff dff_B_gyGRWXvE0_1(.din(w_dff_B_W3BUisI20_1),.dout(w_dff_B_gyGRWXvE0_1),.clk(gclk));
	jdff dff_B_dCMRLTmz6_1(.din(w_dff_B_gyGRWXvE0_1),.dout(w_dff_B_dCMRLTmz6_1),.clk(gclk));
	jdff dff_B_yKxbtZyX9_1(.din(n347),.dout(w_dff_B_yKxbtZyX9_1),.clk(gclk));
	jdff dff_B_slOzX6yU0_1(.din(w_dff_B_yKxbtZyX9_1),.dout(w_dff_B_slOzX6yU0_1),.clk(gclk));
	jdff dff_B_6KHY34Mi1_1(.din(w_dff_B_slOzX6yU0_1),.dout(w_dff_B_6KHY34Mi1_1),.clk(gclk));
	jdff dff_B_n5iJZUgU0_1(.din(w_dff_B_6KHY34Mi1_1),.dout(w_dff_B_n5iJZUgU0_1),.clk(gclk));
	jdff dff_B_wWW4dRvM1_1(.din(w_dff_B_n5iJZUgU0_1),.dout(w_dff_B_wWW4dRvM1_1),.clk(gclk));
	jdff dff_B_R9hpgwhr0_1(.din(w_dff_B_wWW4dRvM1_1),.dout(w_dff_B_R9hpgwhr0_1),.clk(gclk));
	jdff dff_B_HZMw9LuV2_1(.din(w_dff_B_R9hpgwhr0_1),.dout(w_dff_B_HZMw9LuV2_1),.clk(gclk));
	jdff dff_B_ROQ7uGzp9_1(.din(w_dff_B_HZMw9LuV2_1),.dout(w_dff_B_ROQ7uGzp9_1),.clk(gclk));
	jdff dff_B_PwqUDIoi2_1(.din(w_dff_B_ROQ7uGzp9_1),.dout(w_dff_B_PwqUDIoi2_1),.clk(gclk));
	jdff dff_B_npYXXQxt5_1(.din(w_dff_B_PwqUDIoi2_1),.dout(w_dff_B_npYXXQxt5_1),.clk(gclk));
	jdff dff_B_OaMo6QT61_1(.din(w_dff_B_npYXXQxt5_1),.dout(w_dff_B_OaMo6QT61_1),.clk(gclk));
	jdff dff_B_F3DvtgB63_0(.din(n348),.dout(w_dff_B_F3DvtgB63_0),.clk(gclk));
	jdff dff_B_jnyU4Ckc9_0(.din(w_dff_B_F3DvtgB63_0),.dout(w_dff_B_jnyU4Ckc9_0),.clk(gclk));
	jdff dff_B_YlXgNFay8_0(.din(w_dff_B_jnyU4Ckc9_0),.dout(w_dff_B_YlXgNFay8_0),.clk(gclk));
	jdff dff_B_qvbMmWX09_0(.din(w_dff_B_YlXgNFay8_0),.dout(w_dff_B_qvbMmWX09_0),.clk(gclk));
	jdff dff_B_ooPDCouk1_0(.din(w_dff_B_qvbMmWX09_0),.dout(w_dff_B_ooPDCouk1_0),.clk(gclk));
	jdff dff_B_zvMao9e51_0(.din(w_dff_B_ooPDCouk1_0),.dout(w_dff_B_zvMao9e51_0),.clk(gclk));
	jdff dff_B_0aQxesjY8_0(.din(w_dff_B_zvMao9e51_0),.dout(w_dff_B_0aQxesjY8_0),.clk(gclk));
	jdff dff_B_agmjxW9b8_0(.din(w_dff_B_0aQxesjY8_0),.dout(w_dff_B_agmjxW9b8_0),.clk(gclk));
	jdff dff_B_UanMI6PQ5_0(.din(w_dff_B_agmjxW9b8_0),.dout(w_dff_B_UanMI6PQ5_0),.clk(gclk));
	jdff dff_B_0wIwARpR3_0(.din(w_dff_B_UanMI6PQ5_0),.dout(w_dff_B_0wIwARpR3_0),.clk(gclk));
	jdff dff_B_1SozOU5l1_0(.din(w_dff_B_0wIwARpR3_0),.dout(w_dff_B_1SozOU5l1_0),.clk(gclk));
	jdff dff_B_bhURgl5o7_0(.din(w_dff_B_1SozOU5l1_0),.dout(w_dff_B_bhURgl5o7_0),.clk(gclk));
	jdff dff_B_JpMHvu8u7_0(.din(w_dff_B_bhURgl5o7_0),.dout(w_dff_B_JpMHvu8u7_0),.clk(gclk));
	jdff dff_B_ZOgbkHDb3_0(.din(w_dff_B_JpMHvu8u7_0),.dout(w_dff_B_ZOgbkHDb3_0),.clk(gclk));
	jdff dff_A_iWmSOYTH3_1(.dout(w_n344_0[1]),.din(w_dff_A_iWmSOYTH3_1),.clk(gclk));
	jdff dff_A_GIDscngr8_1(.dout(w_dff_A_iWmSOYTH3_1),.din(w_dff_A_GIDscngr8_1),.clk(gclk));
	jdff dff_A_KsALonDl2_1(.dout(w_dff_A_GIDscngr8_1),.din(w_dff_A_KsALonDl2_1),.clk(gclk));
	jdff dff_A_c4dqkhV37_1(.dout(w_dff_A_KsALonDl2_1),.din(w_dff_A_c4dqkhV37_1),.clk(gclk));
	jdff dff_A_MBSH6idT0_1(.dout(w_dff_A_c4dqkhV37_1),.din(w_dff_A_MBSH6idT0_1),.clk(gclk));
	jdff dff_A_UMjil9E39_1(.dout(w_dff_A_MBSH6idT0_1),.din(w_dff_A_UMjil9E39_1),.clk(gclk));
	jdff dff_A_tPbWrMP06_1(.dout(w_dff_A_UMjil9E39_1),.din(w_dff_A_tPbWrMP06_1),.clk(gclk));
	jdff dff_A_sWuEpO6F0_1(.dout(w_dff_A_tPbWrMP06_1),.din(w_dff_A_sWuEpO6F0_1),.clk(gclk));
	jdff dff_A_ikJaiGE46_1(.dout(w_dff_A_sWuEpO6F0_1),.din(w_dff_A_ikJaiGE46_1),.clk(gclk));
	jdff dff_A_sW092USv9_1(.dout(w_dff_A_ikJaiGE46_1),.din(w_dff_A_sW092USv9_1),.clk(gclk));
	jdff dff_A_7OdfY3Yh9_1(.dout(w_dff_A_sW092USv9_1),.din(w_dff_A_7OdfY3Yh9_1),.clk(gclk));
	jdff dff_A_fSftLx0k0_1(.dout(w_n269_1[1]),.din(w_dff_A_fSftLx0k0_1),.clk(gclk));
	jdff dff_A_wQFJnKsT9_2(.dout(w_n269_1[2]),.din(w_dff_A_wQFJnKsT9_2),.clk(gclk));
	jdff dff_B_12tuOhTj8_0(.din(n365),.dout(w_dff_B_12tuOhTj8_0),.clk(gclk));
	jdff dff_B_SCNXTHcA9_0(.din(w_dff_B_12tuOhTj8_0),.dout(w_dff_B_SCNXTHcA9_0),.clk(gclk));
	jdff dff_B_34pwF9lI7_0(.din(w_dff_B_SCNXTHcA9_0),.dout(w_dff_B_34pwF9lI7_0),.clk(gclk));
	jdff dff_B_odoxzutY0_0(.din(w_dff_B_34pwF9lI7_0),.dout(w_dff_B_odoxzutY0_0),.clk(gclk));
	jdff dff_B_uBEPWvoz9_0(.din(w_dff_B_odoxzutY0_0),.dout(w_dff_B_uBEPWvoz9_0),.clk(gclk));
	jdff dff_B_e0bCpcWF3_0(.din(w_dff_B_uBEPWvoz9_0),.dout(w_dff_B_e0bCpcWF3_0),.clk(gclk));
	jdff dff_B_FzxnJLA86_0(.din(w_dff_B_e0bCpcWF3_0),.dout(w_dff_B_FzxnJLA86_0),.clk(gclk));
	jdff dff_B_R17FHUEx6_0(.din(w_dff_B_FzxnJLA86_0),.dout(w_dff_B_R17FHUEx6_0),.clk(gclk));
	jdff dff_B_iM9wOI6B4_0(.din(w_dff_B_R17FHUEx6_0),.dout(w_dff_B_iM9wOI6B4_0),.clk(gclk));
	jdff dff_B_FES3Toxd5_0(.din(w_dff_B_iM9wOI6B4_0),.dout(w_dff_B_FES3Toxd5_0),.clk(gclk));
	jdff dff_B_Pcrt2pkk2_0(.din(w_dff_B_FES3Toxd5_0),.dout(w_dff_B_Pcrt2pkk2_0),.clk(gclk));
	jdff dff_B_6brJrFNK4_0(.din(w_dff_B_Pcrt2pkk2_0),.dout(w_dff_B_6brJrFNK4_0),.clk(gclk));
	jdff dff_B_kOBba82f2_0(.din(w_dff_B_6brJrFNK4_0),.dout(w_dff_B_kOBba82f2_0),.clk(gclk));
	jdff dff_B_y0vioXrN2_0(.din(w_dff_B_kOBba82f2_0),.dout(w_dff_B_y0vioXrN2_0),.clk(gclk));
	jdff dff_B_Y0kMxlKp3_0(.din(w_dff_B_y0vioXrN2_0),.dout(w_dff_B_Y0kMxlKp3_0),.clk(gclk));
	jdff dff_B_MS016RQz8_0(.din(n362),.dout(w_dff_B_MS016RQz8_0),.clk(gclk));
	jdff dff_B_lyofbDAS1_0(.din(w_dff_B_MS016RQz8_0),.dout(w_dff_B_lyofbDAS1_0),.clk(gclk));
	jdff dff_B_h03GltJP2_0(.din(n361),.dout(w_dff_B_h03GltJP2_0),.clk(gclk));
	jdff dff_B_fqBX134S8_0(.din(w_dff_B_h03GltJP2_0),.dout(w_dff_B_fqBX134S8_0),.clk(gclk));
	jdff dff_B_Ad6I2Q6H2_0(.din(w_dff_B_fqBX134S8_0),.dout(w_dff_B_Ad6I2Q6H2_0),.clk(gclk));
	jdff dff_B_iIlpi7Af4_0(.din(w_dff_B_Ad6I2Q6H2_0),.dout(w_dff_B_iIlpi7Af4_0),.clk(gclk));
	jdff dff_B_yiyIbJqJ2_0(.din(w_dff_B_iIlpi7Af4_0),.dout(w_dff_B_yiyIbJqJ2_0),.clk(gclk));
	jdff dff_B_iX483IMn3_0(.din(w_dff_B_yiyIbJqJ2_0),.dout(w_dff_B_iX483IMn3_0),.clk(gclk));
	jdff dff_B_7lY6yjeu8_0(.din(w_dff_B_iX483IMn3_0),.dout(w_dff_B_7lY6yjeu8_0),.clk(gclk));
	jdff dff_B_0KQt4l9f1_0(.din(w_dff_B_7lY6yjeu8_0),.dout(w_dff_B_0KQt4l9f1_0),.clk(gclk));
	jdff dff_B_vMa7JgJg5_0(.din(n310),.dout(w_dff_B_vMa7JgJg5_0),.clk(gclk));
	jdff dff_B_cYj50Ohn8_0(.din(n309),.dout(w_dff_B_cYj50Ohn8_0),.clk(gclk));
	jdff dff_B_GAYwLA6H8_0(.din(w_dff_B_cYj50Ohn8_0),.dout(w_dff_B_GAYwLA6H8_0),.clk(gclk));
	jdff dff_A_mOAYSE0e8_1(.dout(w_n253_1[1]),.din(w_dff_A_mOAYSE0e8_1),.clk(gclk));
	jdff dff_A_WePsK7ok3_1(.dout(w_n298_0[1]),.din(w_dff_A_WePsK7ok3_1),.clk(gclk));
	jdff dff_B_lDqoR1E15_2(.din(n296),.dout(w_dff_B_lDqoR1E15_2),.clk(gclk));
	jdff dff_B_hTSCfNiX7_2(.din(w_dff_B_lDqoR1E15_2),.dout(w_dff_B_hTSCfNiX7_2),.clk(gclk));
	jdff dff_B_juXlPDi56_2(.din(w_dff_B_hTSCfNiX7_2),.dout(w_dff_B_juXlPDi56_2),.clk(gclk));
	jdff dff_B_a5CkEPVo4_0(.din(n291),.dout(w_dff_B_a5CkEPVo4_0),.clk(gclk));
	jdff dff_B_aSJsIa6r1_2(.din(n286),.dout(w_dff_B_aSJsIa6r1_2),.clk(gclk));
	jdff dff_B_Sk0MnWd06_2(.din(w_dff_B_aSJsIa6r1_2),.dout(w_dff_B_Sk0MnWd06_2),.clk(gclk));
	jdff dff_A_lCyFUNZz8_1(.dout(w_n247_0[1]),.din(w_dff_A_lCyFUNZz8_1),.clk(gclk));
	jdff dff_A_iwoknT9B4_2(.dout(w_n247_0[2]),.din(w_dff_A_iwoknT9B4_2),.clk(gclk));
	jdff dff_B_nz6nYAlU1_0(.din(n372),.dout(w_dff_B_nz6nYAlU1_0),.clk(gclk));
	jdff dff_B_V7dRqMkb6_0(.din(w_dff_B_nz6nYAlU1_0),.dout(w_dff_B_V7dRqMkb6_0),.clk(gclk));
	jdff dff_B_TngN26zw1_0(.din(w_dff_B_V7dRqMkb6_0),.dout(w_dff_B_TngN26zw1_0),.clk(gclk));
	jdff dff_B_xZCUJF3B7_0(.din(w_dff_B_TngN26zw1_0),.dout(w_dff_B_xZCUJF3B7_0),.clk(gclk));
	jdff dff_B_8sLvhIEi7_0(.din(w_dff_B_xZCUJF3B7_0),.dout(w_dff_B_8sLvhIEi7_0),.clk(gclk));
	jdff dff_B_fxz3TBLs6_0(.din(w_dff_B_8sLvhIEi7_0),.dout(w_dff_B_fxz3TBLs6_0),.clk(gclk));
	jdff dff_B_nutD5hqc5_0(.din(w_dff_B_fxz3TBLs6_0),.dout(w_dff_B_nutD5hqc5_0),.clk(gclk));
	jdff dff_B_spzrTbcT1_0(.din(w_dff_B_nutD5hqc5_0),.dout(w_dff_B_spzrTbcT1_0),.clk(gclk));
	jdff dff_B_7wcgNGc58_0(.din(w_dff_B_spzrTbcT1_0),.dout(w_dff_B_7wcgNGc58_0),.clk(gclk));
	jdff dff_B_qJewMhEt2_0(.din(w_dff_B_7wcgNGc58_0),.dout(w_dff_B_qJewMhEt2_0),.clk(gclk));
	jdff dff_B_wO5oH2yq7_0(.din(w_dff_B_qJewMhEt2_0),.dout(w_dff_B_wO5oH2yq7_0),.clk(gclk));
	jdff dff_B_I03464Z71_0(.din(w_dff_B_wO5oH2yq7_0),.dout(w_dff_B_I03464Z71_0),.clk(gclk));
	jdff dff_B_c9pJwPQJ5_0(.din(n369),.dout(w_dff_B_c9pJwPQJ5_0),.clk(gclk));
	jdff dff_B_y2a4YXIC7_0(.din(w_dff_B_c9pJwPQJ5_0),.dout(w_dff_B_y2a4YXIC7_0),.clk(gclk));
	jdff dff_B_LeQxV6TU7_0(.din(w_dff_B_y2a4YXIC7_0),.dout(w_dff_B_LeQxV6TU7_0),.clk(gclk));
	jdff dff_B_eAkV4tXr9_0(.din(w_dff_B_LeQxV6TU7_0),.dout(w_dff_B_eAkV4tXr9_0),.clk(gclk));
	jdff dff_B_xErKtZCo4_0(.din(w_dff_B_eAkV4tXr9_0),.dout(w_dff_B_xErKtZCo4_0),.clk(gclk));
	jdff dff_B_fLaqRo0Y6_0(.din(w_dff_B_xErKtZCo4_0),.dout(w_dff_B_fLaqRo0Y6_0),.clk(gclk));
	jdff dff_B_iNUBiQYV9_0(.din(w_dff_B_fLaqRo0Y6_0),.dout(w_dff_B_iNUBiQYV9_0),.clk(gclk));
	jdff dff_B_UVCa8OEN7_0(.din(w_dff_B_iNUBiQYV9_0),.dout(w_dff_B_UVCa8OEN7_0),.clk(gclk));
	jdff dff_B_XjSC0c9B5_0(.din(w_dff_B_UVCa8OEN7_0),.dout(w_dff_B_XjSC0c9B5_0),.clk(gclk));
	jdff dff_B_WBmJI8q53_0(.din(w_dff_B_XjSC0c9B5_0),.dout(w_dff_B_WBmJI8q53_0),.clk(gclk));
	jdff dff_B_moIPe1Fm6_0(.din(w_dff_B_WBmJI8q53_0),.dout(w_dff_B_moIPe1Fm6_0),.clk(gclk));
	jdff dff_B_pCFVqoTP1_0(.din(w_dff_B_moIPe1Fm6_0),.dout(w_dff_B_pCFVqoTP1_0),.clk(gclk));
	jdff dff_B_w1YOFz4z6_0(.din(w_dff_B_pCFVqoTP1_0),.dout(w_dff_B_w1YOFz4z6_0),.clk(gclk));
	jdff dff_B_ETtamJp77_0(.din(w_dff_B_w1YOFz4z6_0),.dout(w_dff_B_ETtamJp77_0),.clk(gclk));
	jdff dff_A_rAEbi5pg6_2(.dout(w_n61_1[2]),.din(w_dff_A_rAEbi5pg6_2),.clk(gclk));
	jdff dff_A_mpX9JVRz0_2(.dout(w_dff_A_rAEbi5pg6_2),.din(w_dff_A_mpX9JVRz0_2),.clk(gclk));
	jdff dff_A_1JSmv3Xz2_2(.dout(w_dff_A_mpX9JVRz0_2),.din(w_dff_A_1JSmv3Xz2_2),.clk(gclk));
	jdff dff_A_w1L5U8hZ8_2(.dout(w_dff_A_1JSmv3Xz2_2),.din(w_dff_A_w1L5U8hZ8_2),.clk(gclk));
	jdff dff_A_so2v8p0p3_2(.dout(w_dff_A_w1L5U8hZ8_2),.din(w_dff_A_so2v8p0p3_2),.clk(gclk));
	jdff dff_A_jlSTJxON8_2(.dout(w_dff_A_so2v8p0p3_2),.din(w_dff_A_jlSTJxON8_2),.clk(gclk));
	jdff dff_A_EhNoLLJc3_2(.dout(w_dff_A_jlSTJxON8_2),.din(w_dff_A_EhNoLLJc3_2),.clk(gclk));
	jdff dff_A_tAnzTqMF4_2(.dout(w_dff_A_EhNoLLJc3_2),.din(w_dff_A_tAnzTqMF4_2),.clk(gclk));
	jdff dff_A_LBotY2eC5_2(.dout(w_dff_A_tAnzTqMF4_2),.din(w_dff_A_LBotY2eC5_2),.clk(gclk));
	jdff dff_A_whoP7SOZ7_2(.dout(w_dff_A_LBotY2eC5_2),.din(w_dff_A_whoP7SOZ7_2),.clk(gclk));
	jdff dff_A_m6tq2qpa7_2(.dout(w_dff_A_whoP7SOZ7_2),.din(w_dff_A_m6tq2qpa7_2),.clk(gclk));
	jdff dff_B_YHUknnpY0_1(.din(n325),.dout(w_dff_B_YHUknnpY0_1),.clk(gclk));
	jdff dff_B_HOwBZZzy8_1(.din(n331),.dout(w_dff_B_HOwBZZzy8_1),.clk(gclk));
	jdff dff_B_aiRoMdoG5_1(.din(w_dff_B_HOwBZZzy8_1),.dout(w_dff_B_aiRoMdoG5_1),.clk(gclk));
	jdff dff_B_ezAnpGU13_1(.din(n333),.dout(w_dff_B_ezAnpGU13_1),.clk(gclk));
	jdff dff_B_iIqvjNOa3_0(.din(n328),.dout(w_dff_B_iIqvjNOa3_0),.clk(gclk));
	jdff dff_B_pJ5gaPhu0_0(.din(w_dff_B_iIqvjNOa3_0),.dout(w_dff_B_pJ5gaPhu0_0),.clk(gclk));
	jdff dff_B_n6HfhzeT0_0(.din(n324),.dout(w_dff_B_n6HfhzeT0_0),.clk(gclk));
	jdff dff_B_d4MGz1xW8_1(.din(n317),.dout(w_dff_B_d4MGz1xW8_1),.clk(gclk));
	jdff dff_B_mYZ6SdKZ6_0(.din(n322),.dout(w_dff_B_mYZ6SdKZ6_0),.clk(gclk));
	jdff dff_A_5eRgs1NA1_0(.dout(w_n321_0[0]),.din(w_dff_A_5eRgs1NA1_0),.clk(gclk));
	jdff dff_A_kzyFlC3Z5_0(.dout(w_dff_A_5eRgs1NA1_0),.din(w_dff_A_kzyFlC3Z5_0),.clk(gclk));
	jdff dff_A_QbYjEiid8_1(.dout(w_n300_0[1]),.din(w_dff_A_QbYjEiid8_1),.clk(gclk));
	jdff dff_B_p6TVTbM01_0(.din(n319),.dout(w_dff_B_p6TVTbM01_0),.clk(gclk));
	jdff dff_A_xnd6brWN0_1(.dout(w_n316_0[1]),.din(w_dff_A_xnd6brWN0_1),.clk(gclk));
	jdff dff_B_d0hNRf772_3(.din(n315),.dout(w_dff_B_d0hNRf772_3),.clk(gclk));
	jdff dff_B_qOkiHl6x6_3(.din(w_dff_B_d0hNRf772_3),.dout(w_dff_B_qOkiHl6x6_3),.clk(gclk));
	jdff dff_B_BVBFn80e3_3(.din(w_dff_B_qOkiHl6x6_3),.dout(w_dff_B_BVBFn80e3_3),.clk(gclk));
	jdff dff_A_Fk3ksdOx2_0(.dout(w_n313_0[0]),.din(w_dff_A_Fk3ksdOx2_0),.clk(gclk));
	jdff dff_A_C1rSbdtx0_0(.dout(w_dff_A_Fk3ksdOx2_0),.din(w_dff_A_C1rSbdtx0_0),.clk(gclk));
	jdff dff_A_E873VoV34_2(.dout(w_n253_0[2]),.din(w_dff_A_E873VoV34_2),.clk(gclk));
	jdff dff_A_FweZJOWU1_0(.dout(w_G953_1[0]),.din(w_dff_A_FweZJOWU1_0),.clk(gclk));
	jdff dff_A_seyGBe7W1_0(.dout(w_dff_A_FweZJOWU1_0),.din(w_dff_A_seyGBe7W1_0),.clk(gclk));
	jdff dff_A_aYCmzNej5_0(.dout(w_dff_A_seyGBe7W1_0),.din(w_dff_A_aYCmzNej5_0),.clk(gclk));
	jdff dff_A_xqMIXTHk3_0(.dout(w_dff_A_aYCmzNej5_0),.din(w_dff_A_xqMIXTHk3_0),.clk(gclk));
	jdff dff_A_pDYjh9H73_1(.dout(w_G953_1[1]),.din(w_dff_A_pDYjh9H73_1),.clk(gclk));
	jdff dff_A_NrYsuE4t4_1(.dout(w_dff_A_pDYjh9H73_1),.din(w_dff_A_NrYsuE4t4_1),.clk(gclk));
	jdff dff_A_SvPx8n7A4_1(.dout(w_dff_A_NrYsuE4t4_1),.din(w_dff_A_SvPx8n7A4_1),.clk(gclk));
	jdff dff_A_PHOxtYAj4_1(.dout(w_dff_A_SvPx8n7A4_1),.din(w_dff_A_PHOxtYAj4_1),.clk(gclk));
	jdff dff_B_gpjAV2IP4_0(.din(n241),.dout(w_dff_B_gpjAV2IP4_0),.clk(gclk));
	jdff dff_A_yMeXOukv4_0(.dout(w_n194_0[0]),.din(w_dff_A_yMeXOukv4_0),.clk(gclk));
	jdff dff_A_kiesjfqD5_1(.dout(w_n222_0[1]),.din(w_dff_A_kiesjfqD5_1),.clk(gclk));
	jdff dff_A_lkebg2m49_0(.dout(w_n218_1[0]),.din(w_dff_A_lkebg2m49_0),.clk(gclk));
	jdff dff_A_saCiEqOW4_0(.dout(w_dff_A_lkebg2m49_0),.din(w_dff_A_saCiEqOW4_0),.clk(gclk));
	jdff dff_A_IeajTyD19_2(.dout(w_n218_0[2]),.din(w_dff_A_IeajTyD19_2),.clk(gclk));
	jdff dff_A_cOP0zIfQ1_2(.dout(w_dff_A_IeajTyD19_2),.din(w_dff_A_cOP0zIfQ1_2),.clk(gclk));
	jdff dff_B_TdvY5iUP8_3(.din(n217),.dout(w_dff_B_TdvY5iUP8_3),.clk(gclk));
	jdff dff_B_vwyHxJUz9_2(.din(n216),.dout(w_dff_B_vwyHxJUz9_2),.clk(gclk));
	jdff dff_A_ALQxHeVA9_1(.dout(w_n184_1[1]),.din(w_dff_A_ALQxHeVA9_1),.clk(gclk));
	jdff dff_A_3SgIPXym6_0(.dout(w_n184_0[0]),.din(w_dff_A_3SgIPXym6_0),.clk(gclk));
	jdff dff_A_qdqTPmX23_0(.dout(w_dff_A_3SgIPXym6_0),.din(w_dff_A_qdqTPmX23_0),.clk(gclk));
	jdff dff_A_8PK2wp6P7_0(.dout(w_dff_A_qdqTPmX23_0),.din(w_dff_A_8PK2wp6P7_0),.clk(gclk));
	jdff dff_A_fu73Tlq03_0(.dout(w_dff_A_8PK2wp6P7_0),.din(w_dff_A_fu73Tlq03_0),.clk(gclk));
	jdff dff_A_lJgjFNBv1_0(.dout(w_dff_A_fu73Tlq03_0),.din(w_dff_A_lJgjFNBv1_0),.clk(gclk));
	jdff dff_A_Kc7QnGub5_2(.dout(w_n184_0[2]),.din(w_dff_A_Kc7QnGub5_2),.clk(gclk));
	jdff dff_A_kYqCcBmS4_2(.dout(w_dff_A_Kc7QnGub5_2),.din(w_dff_A_kYqCcBmS4_2),.clk(gclk));
	jdff dff_A_VxmxJFC47_2(.dout(w_dff_A_kYqCcBmS4_2),.din(w_dff_A_VxmxJFC47_2),.clk(gclk));
	jdff dff_A_zAzbZurG5_2(.dout(w_dff_A_VxmxJFC47_2),.din(w_dff_A_zAzbZurG5_2),.clk(gclk));
	jdff dff_A_mkWMQELe8_2(.dout(w_dff_A_zAzbZurG5_2),.din(w_dff_A_mkWMQELe8_2),.clk(gclk));
	jdff dff_A_JH7mNzYY0_2(.dout(w_dff_A_mkWMQELe8_2),.din(w_dff_A_JH7mNzYY0_2),.clk(gclk));
	jdff dff_A_TkVW8YX26_0(.dout(w_n181_0[0]),.din(w_dff_A_TkVW8YX26_0),.clk(gclk));
	jdff dff_A_6GvLxx1O3_0(.dout(w_dff_A_TkVW8YX26_0),.din(w_dff_A_6GvLxx1O3_0),.clk(gclk));
	jdff dff_B_r8CDHUvp8_1(.din(n232),.dout(w_dff_B_r8CDHUvp8_1),.clk(gclk));
	jdff dff_A_DSmlpsRc5_0(.dout(w_n188_0[0]),.din(w_dff_A_DSmlpsRc5_0),.clk(gclk));
	jdff dff_A_CKNJDBMO5_1(.dout(w_n178_0[1]),.din(w_dff_A_CKNJDBMO5_1),.clk(gclk));
	jdff dff_B_OTz8mCiT7_3(.din(n205),.dout(w_dff_B_OTz8mCiT7_3),.clk(gclk));
	jdff dff_B_pCvg8te93_3(.din(w_dff_B_OTz8mCiT7_3),.dout(w_dff_B_pCvg8te93_3),.clk(gclk));
	jdff dff_B_FjK7oy4T4_3(.din(w_dff_B_pCvg8te93_3),.dout(w_dff_B_FjK7oy4T4_3),.clk(gclk));
	jdff dff_A_FKwiEQCc1_1(.dout(w_n175_0[1]),.din(w_dff_A_FKwiEQCc1_1),.clk(gclk));
	jdff dff_B_38toSO1e7_2(.din(n175),.dout(w_dff_B_38toSO1e7_2),.clk(gclk));
	jdff dff_B_SuaWyHO09_0(.din(n230),.dout(w_dff_B_SuaWyHO09_0),.clk(gclk));
	jdff dff_B_POD5FexQ7_2(.din(n200),.dout(w_dff_B_POD5FexQ7_2),.clk(gclk));
	jdff dff_A_J6r5C7CT5_0(.dout(w_n199_0[0]),.din(w_dff_A_J6r5C7CT5_0),.clk(gclk));
	jdff dff_A_3Ik7xgJC2_0(.dout(w_dff_A_J6r5C7CT5_0),.din(w_dff_A_3Ik7xgJC2_0),.clk(gclk));
	jdff dff_A_zLjQ5DjK5_0(.dout(w_dff_A_3Ik7xgJC2_0),.din(w_dff_A_zLjQ5DjK5_0),.clk(gclk));
	jdff dff_A_COV5c8io0_1(.dout(w_n199_0[1]),.din(w_dff_A_COV5c8io0_1),.clk(gclk));
	jdff dff_A_R3eqTsLf5_1(.dout(w_dff_A_COV5c8io0_1),.din(w_dff_A_R3eqTsLf5_1),.clk(gclk));
	jdff dff_A_A5IuR94N6_1(.dout(w_dff_A_R3eqTsLf5_1),.din(w_dff_A_A5IuR94N6_1),.clk(gclk));
	jdff dff_A_Clk3MhQA4_0(.dout(w_n198_1[0]),.din(w_dff_A_Clk3MhQA4_0),.clk(gclk));
	jdff dff_A_f7ZbnAm77_2(.dout(w_n198_1[2]),.din(w_dff_A_f7ZbnAm77_2),.clk(gclk));
	jdff dff_A_I1kg5hwF5_1(.dout(w_n198_0[1]),.din(w_dff_A_I1kg5hwF5_1),.clk(gclk));
	jdff dff_A_TmbHF47T2_2(.dout(w_n198_0[2]),.din(w_dff_A_TmbHF47T2_2),.clk(gclk));
	jdff dff_B_UYS0eS4J9_3(.din(n174),.dout(w_dff_B_UYS0eS4J9_3),.clk(gclk));
	jdff dff_B_WUUlKJsV5_1(.din(n161),.dout(w_dff_B_WUUlKJsV5_1),.clk(gclk));
	jdff dff_B_uklByK084_1(.din(w_dff_B_WUUlKJsV5_1),.dout(w_dff_B_uklByK084_1),.clk(gclk));
	jdff dff_B_YRVpBmOv9_1(.din(w_dff_B_uklByK084_1),.dout(w_dff_B_YRVpBmOv9_1),.clk(gclk));
	jdff dff_B_JZn9NJq96_1(.din(w_dff_B_YRVpBmOv9_1),.dout(w_dff_B_JZn9NJq96_1),.clk(gclk));
	jdff dff_B_5ogbdSgK0_1(.din(w_dff_B_JZn9NJq96_1),.dout(w_dff_B_5ogbdSgK0_1),.clk(gclk));
	jdff dff_B_j1bxsFnM1_1(.din(w_dff_B_5ogbdSgK0_1),.dout(w_dff_B_j1bxsFnM1_1),.clk(gclk));
	jdff dff_A_tlUmzFcf7_1(.dout(w_n156_0[1]),.din(w_dff_A_tlUmzFcf7_1),.clk(gclk));
	jdff dff_A_WnJsyQ5g5_2(.dout(w_n156_0[2]),.din(w_dff_A_WnJsyQ5g5_2),.clk(gclk));
	jdff dff_B_XafTWfcB9_1(.din(n145),.dout(w_dff_B_XafTWfcB9_1),.clk(gclk));
	jdff dff_B_K0R0tMJv5_1(.din(w_dff_B_XafTWfcB9_1),.dout(w_dff_B_K0R0tMJv5_1),.clk(gclk));
	jdff dff_B_FXHEeOVC0_1(.din(w_dff_B_K0R0tMJv5_1),.dout(w_dff_B_FXHEeOVC0_1),.clk(gclk));
	jdff dff_B_oYG8wl3J8_1(.din(w_dff_B_FXHEeOVC0_1),.dout(w_dff_B_oYG8wl3J8_1),.clk(gclk));
	jdff dff_B_BFqQdm8s5_1(.din(w_dff_B_oYG8wl3J8_1),.dout(w_dff_B_BFqQdm8s5_1),.clk(gclk));
	jdff dff_B_CEpUt50U2_1(.din(w_dff_B_BFqQdm8s5_1),.dout(w_dff_B_CEpUt50U2_1),.clk(gclk));
	jdff dff_A_QzJM2grK0_1(.dout(w_n153_0[1]),.din(w_dff_A_QzJM2grK0_1),.clk(gclk));
	jdff dff_A_cTybTbj10_1(.dout(w_dff_A_QzJM2grK0_1),.din(w_dff_A_cTybTbj10_1),.clk(gclk));
	jdff dff_A_W3wxZAmc9_1(.dout(w_dff_A_cTybTbj10_1),.din(w_dff_A_W3wxZAmc9_1),.clk(gclk));
	jdff dff_A_ul88dtbB2_1(.dout(w_dff_A_W3wxZAmc9_1),.din(w_dff_A_ul88dtbB2_1),.clk(gclk));
	jdff dff_A_Vzqp7Vvv8_1(.dout(w_dff_A_ul88dtbB2_1),.din(w_dff_A_Vzqp7Vvv8_1),.clk(gclk));
	jdff dff_A_8EXInkQS7_1(.dout(w_dff_A_Vzqp7Vvv8_1),.din(w_dff_A_8EXInkQS7_1),.clk(gclk));
	jdff dff_A_wyUeuZlK6_1(.dout(w_dff_A_8EXInkQS7_1),.din(w_dff_A_wyUeuZlK6_1),.clk(gclk));
	jdff dff_B_WL4qxRGH8_1(.din(n147),.dout(w_dff_B_WL4qxRGH8_1),.clk(gclk));
	jdff dff_B_lk8j5RSt0_1(.din(w_dff_B_WL4qxRGH8_1),.dout(w_dff_B_lk8j5RSt0_1),.clk(gclk));
	jdff dff_B_Nga9kcJ61_1(.din(w_dff_B_lk8j5RSt0_1),.dout(w_dff_B_Nga9kcJ61_1),.clk(gclk));
	jdff dff_B_8GAf0KfY6_0(.din(n150),.dout(w_dff_B_8GAf0KfY6_0),.clk(gclk));
	jdff dff_B_qVIVlfkD1_0(.din(w_dff_B_8GAf0KfY6_0),.dout(w_dff_B_qVIVlfkD1_0),.clk(gclk));
	jdff dff_A_U3yPJwqJ7_1(.dout(w_G475_0[1]),.din(w_dff_A_U3yPJwqJ7_1),.clk(gclk));
	jdff dff_A_SFvtqPTS6_1(.dout(w_dff_A_U3yPJwqJ7_1),.din(w_dff_A_SFvtqPTS6_1),.clk(gclk));
	jdff dff_A_0ninUoKv6_1(.dout(w_dff_A_SFvtqPTS6_1),.din(w_dff_A_0ninUoKv6_1),.clk(gclk));
	jdff dff_A_Kd5FgdbA3_1(.dout(w_dff_A_0ninUoKv6_1),.din(w_dff_A_Kd5FgdbA3_1),.clk(gclk));
	jdff dff_A_TKaqkm4w4_1(.dout(w_dff_A_Kd5FgdbA3_1),.din(w_dff_A_TKaqkm4w4_1),.clk(gclk));
	jdff dff_A_fUZ5YBIY0_1(.dout(w_dff_A_TKaqkm4w4_1),.din(w_dff_A_fUZ5YBIY0_1),.clk(gclk));
	jdff dff_A_tKNjPyhs0_1(.dout(w_dff_A_fUZ5YBIY0_1),.din(w_dff_A_tKNjPyhs0_1),.clk(gclk));
	jdff dff_B_sFbHan702_3(.din(n144),.dout(w_dff_B_sFbHan702_3),.clk(gclk));
	jdff dff_A_e7HYpYfB3_0(.dout(w_n143_1[0]),.din(w_dff_A_e7HYpYfB3_0),.clk(gclk));
	jdff dff_A_r3KvVKkS4_0(.dout(w_dff_A_e7HYpYfB3_0),.din(w_dff_A_r3KvVKkS4_0),.clk(gclk));
	jdff dff_A_2BuvrVVT2_1(.dout(w_n143_1[1]),.din(w_dff_A_2BuvrVVT2_1),.clk(gclk));
	jdff dff_A_0l7TO2iJ5_1(.dout(w_dff_A_2BuvrVVT2_1),.din(w_dff_A_0l7TO2iJ5_1),.clk(gclk));
	jdff dff_A_fyMyRoDP8_1(.dout(w_n143_0[1]),.din(w_dff_A_fyMyRoDP8_1),.clk(gclk));
	jdff dff_A_P18OMZwK3_1(.dout(w_dff_A_fyMyRoDP8_1),.din(w_dff_A_P18OMZwK3_1),.clk(gclk));
	jdff dff_A_NnGvldnt2_2(.dout(w_n143_0[2]),.din(w_dff_A_NnGvldnt2_2),.clk(gclk));
	jdff dff_A_jA8P3gX08_2(.dout(w_dff_A_NnGvldnt2_2),.din(w_dff_A_jA8P3gX08_2),.clk(gclk));
	jdff dff_A_58Aotwi94_1(.dout(w_n141_0[1]),.din(w_dff_A_58Aotwi94_1),.clk(gclk));
	jdff dff_A_fJyzpPt58_1(.dout(w_dff_A_58Aotwi94_1),.din(w_dff_A_fJyzpPt58_1),.clk(gclk));
	jdff dff_A_NbZ0Cjgl5_1(.dout(w_dff_A_fJyzpPt58_1),.din(w_dff_A_NbZ0Cjgl5_1),.clk(gclk));
	jdff dff_A_40Q8aFAP7_1(.dout(w_dff_A_NbZ0Cjgl5_1),.din(w_dff_A_40Q8aFAP7_1),.clk(gclk));
	jdff dff_A_Umaz5U2i0_1(.dout(w_dff_A_40Q8aFAP7_1),.din(w_dff_A_Umaz5U2i0_1),.clk(gclk));
	jdff dff_A_KZ1JfUh10_1(.dout(w_dff_A_Umaz5U2i0_1),.din(w_dff_A_KZ1JfUh10_1),.clk(gclk));
	jdff dff_A_xpjQbR8o5_1(.dout(w_dff_A_KZ1JfUh10_1),.din(w_dff_A_xpjQbR8o5_1),.clk(gclk));
	jdff dff_A_7m5EH2e48_1(.dout(w_dff_A_xpjQbR8o5_1),.din(w_dff_A_7m5EH2e48_1),.clk(gclk));
	jdff dff_A_cvJ4WcHM2_1(.dout(w_dff_A_7m5EH2e48_1),.din(w_dff_A_cvJ4WcHM2_1),.clk(gclk));
	jdff dff_B_beFGc0zb8_1(.din(n136),.dout(w_dff_B_beFGc0zb8_1),.clk(gclk));
	jdff dff_A_M0K3L6hV2_1(.dout(w_G478_0[1]),.din(w_dff_A_M0K3L6hV2_1),.clk(gclk));
	jdff dff_A_X7XREVbh4_1(.dout(w_dff_A_M0K3L6hV2_1),.din(w_dff_A_X7XREVbh4_1),.clk(gclk));
	jdff dff_A_axafGabF4_1(.dout(w_dff_A_X7XREVbh4_1),.din(w_dff_A_axafGabF4_1),.clk(gclk));
	jdff dff_A_Tl530lgX9_1(.dout(w_dff_A_axafGabF4_1),.din(w_dff_A_Tl530lgX9_1),.clk(gclk));
	jdff dff_A_FHA5ViFc5_1(.dout(w_dff_A_Tl530lgX9_1),.din(w_dff_A_FHA5ViFc5_1),.clk(gclk));
	jdff dff_A_KBWSiNeo9_0(.dout(w_n134_0[0]),.din(w_dff_A_KBWSiNeo9_0),.clk(gclk));
	jdff dff_A_JGGWZiWw8_0(.dout(w_dff_A_KBWSiNeo9_0),.din(w_dff_A_JGGWZiWw8_0),.clk(gclk));
	jdff dff_A_tzQcv87I2_0(.dout(w_dff_A_JGGWZiWw8_0),.din(w_dff_A_tzQcv87I2_0),.clk(gclk));
	jdff dff_A_uLz37Kji1_0(.dout(w_dff_A_tzQcv87I2_0),.din(w_dff_A_uLz37Kji1_0),.clk(gclk));
	jdff dff_A_AccwtbgX6_0(.dout(w_dff_A_uLz37Kji1_0),.din(w_dff_A_AccwtbgX6_0),.clk(gclk));
	jdff dff_A_u8ECvRTL7_2(.dout(w_n134_0[2]),.din(w_dff_A_u8ECvRTL7_2),.clk(gclk));
	jdff dff_A_eylm4DLO2_2(.dout(w_dff_A_u8ECvRTL7_2),.din(w_dff_A_eylm4DLO2_2),.clk(gclk));
	jdff dff_A_jp9X043D2_2(.dout(w_dff_A_eylm4DLO2_2),.din(w_dff_A_jp9X043D2_2),.clk(gclk));
	jdff dff_A_I8RaLy6L4_2(.dout(w_dff_A_jp9X043D2_2),.din(w_dff_A_I8RaLy6L4_2),.clk(gclk));
	jdff dff_A_d3Ly3WpX8_2(.dout(w_dff_A_I8RaLy6L4_2),.din(w_dff_A_d3Ly3WpX8_2),.clk(gclk));
	jdff dff_A_zQt3MYHd7_0(.dout(w_n131_0[0]),.din(w_dff_A_zQt3MYHd7_0),.clk(gclk));
	jdff dff_A_JyL1JZpr0_0(.dout(w_dff_A_zQt3MYHd7_0),.din(w_dff_A_JyL1JZpr0_0),.clk(gclk));
	jdff dff_A_zEL2RL1p2_0(.dout(w_dff_A_JyL1JZpr0_0),.din(w_dff_A_zEL2RL1p2_0),.clk(gclk));
	jdff dff_A_bDYceyS95_0(.dout(w_G902_3[0]),.din(w_dff_A_bDYceyS95_0),.clk(gclk));
	jdff dff_A_iVrP5siR5_0(.dout(w_dff_A_bDYceyS95_0),.din(w_dff_A_iVrP5siR5_0),.clk(gclk));
	jdff dff_A_XSA9UEDR7_0(.dout(w_dff_A_iVrP5siR5_0),.din(w_dff_A_XSA9UEDR7_0),.clk(gclk));
	jdff dff_A_1YYsurjX7_0(.dout(w_dff_A_XSA9UEDR7_0),.din(w_dff_A_1YYsurjX7_0),.clk(gclk));
	jdff dff_A_KZxb49b16_0(.dout(w_dff_A_1YYsurjX7_0),.din(w_dff_A_KZxb49b16_0),.clk(gclk));
	jdff dff_A_UTbR2gQ65_0(.dout(w_dff_A_KZxb49b16_0),.din(w_dff_A_UTbR2gQ65_0),.clk(gclk));
	jdff dff_A_DkAMU0IW5_0(.dout(w_dff_A_UTbR2gQ65_0),.din(w_dff_A_DkAMU0IW5_0),.clk(gclk));
	jdff dff_A_L645vFdR8_0(.dout(w_dff_A_DkAMU0IW5_0),.din(w_dff_A_L645vFdR8_0),.clk(gclk));
	jdff dff_A_fnjVZbrO0_0(.dout(w_dff_A_L645vFdR8_0),.din(w_dff_A_fnjVZbrO0_0),.clk(gclk));
	jdff dff_A_HX0s9Wqt5_0(.dout(w_dff_A_fnjVZbrO0_0),.din(w_dff_A_HX0s9Wqt5_0),.clk(gclk));
	jdff dff_A_C1oU3Xa71_0(.dout(w_dff_A_HX0s9Wqt5_0),.din(w_dff_A_C1oU3Xa71_0),.clk(gclk));
	jdff dff_B_IUWquhTG7_2(.din(n129),.dout(w_dff_B_IUWquhTG7_2),.clk(gclk));
	jdff dff_A_Nb8TqsbK3_0(.dout(w_n128_0[0]),.din(w_dff_A_Nb8TqsbK3_0),.clk(gclk));
	jdff dff_A_Fozfva622_0(.dout(w_dff_A_Nb8TqsbK3_0),.din(w_dff_A_Fozfva622_0),.clk(gclk));
	jdff dff_A_FlxckdQo0_0(.dout(w_dff_A_Fozfva622_0),.din(w_dff_A_FlxckdQo0_0),.clk(gclk));
	jdff dff_A_yCPGP2PD1_0(.dout(w_dff_A_FlxckdQo0_0),.din(w_dff_A_yCPGP2PD1_0),.clk(gclk));
	jdff dff_A_RuIPQOuh1_0(.dout(w_dff_A_yCPGP2PD1_0),.din(w_dff_A_RuIPQOuh1_0),.clk(gclk));
	jdff dff_A_kfeGpP0u2_0(.dout(w_dff_A_RuIPQOuh1_0),.din(w_dff_A_kfeGpP0u2_0),.clk(gclk));
	jdff dff_A_TvEj2aQY8_0(.dout(w_dff_A_kfeGpP0u2_0),.din(w_dff_A_TvEj2aQY8_0),.clk(gclk));
	jdff dff_A_SvLAo0DM1_0(.dout(w_dff_A_TvEj2aQY8_0),.din(w_dff_A_SvLAo0DM1_0),.clk(gclk));
	jdff dff_B_eYBTCMCd2_3(.din(n128),.dout(w_dff_B_eYBTCMCd2_3),.clk(gclk));
	jdff dff_B_dJQNrJGn0_3(.din(w_dff_B_eYBTCMCd2_3),.dout(w_dff_B_dJQNrJGn0_3),.clk(gclk));
	jdff dff_A_2NVq1sYn1_1(.dout(w_n123_1[1]),.din(w_dff_A_2NVq1sYn1_1),.clk(gclk));
	jdff dff_A_ZtEfrsOh1_1(.dout(w_n123_0[1]),.din(w_dff_A_ZtEfrsOh1_1),.clk(gclk));
	jdff dff_A_StFfRhm90_1(.dout(w_dff_A_ZtEfrsOh1_1),.din(w_dff_A_StFfRhm90_1),.clk(gclk));
	jdff dff_B_DleYBDfH4_1(.din(n110),.dout(w_dff_B_DleYBDfH4_1),.clk(gclk));
	jdff dff_B_wKOLTsfF6_1(.din(n112),.dout(w_dff_B_wKOLTsfF6_1),.clk(gclk));
	jdff dff_B_g5j2zA5F0_1(.din(w_dff_B_wKOLTsfF6_1),.dout(w_dff_B_g5j2zA5F0_1),.clk(gclk));
	jdff dff_B_VC0glfyq1_1(.din(w_dff_B_g5j2zA5F0_1),.dout(w_dff_B_VC0glfyq1_1),.clk(gclk));
	jdff dff_B_eidb97056_1(.din(w_dff_B_VC0glfyq1_1),.dout(w_dff_B_eidb97056_1),.clk(gclk));
	jdff dff_A_UGyPXClN7_0(.dout(w_n119_0[0]),.din(w_dff_A_UGyPXClN7_0),.clk(gclk));
	jdff dff_A_N6FXMaXC1_0(.dout(w_dff_A_UGyPXClN7_0),.din(w_dff_A_N6FXMaXC1_0),.clk(gclk));
	jdff dff_A_FRKufGZR2_0(.dout(w_dff_A_N6FXMaXC1_0),.din(w_dff_A_FRKufGZR2_0),.clk(gclk));
	jdff dff_A_lZnqX16A3_0(.dout(w_dff_A_FRKufGZR2_0),.din(w_dff_A_lZnqX16A3_0),.clk(gclk));
	jdff dff_A_XnJVb39u4_0(.dout(w_dff_A_lZnqX16A3_0),.din(w_dff_A_XnJVb39u4_0),.clk(gclk));
	jdff dff_A_7svpxIJm4_0(.dout(w_dff_A_XnJVb39u4_0),.din(w_dff_A_7svpxIJm4_0),.clk(gclk));
	jdff dff_A_8Wr2l8kp8_0(.dout(w_dff_A_7svpxIJm4_0),.din(w_dff_A_8Wr2l8kp8_0),.clk(gclk));
	jdff dff_A_inAgN7b92_0(.dout(w_dff_A_8Wr2l8kp8_0),.din(w_dff_A_inAgN7b92_0),.clk(gclk));
	jdff dff_B_fS85srqe2_0(.din(n118),.dout(w_dff_B_fS85srqe2_0),.clk(gclk));
	jdff dff_A_P8cvXJkE8_1(.dout(w_G469_0[1]),.din(w_dff_A_P8cvXJkE8_1),.clk(gclk));
	jdff dff_A_XaHotoUV6_1(.dout(w_dff_A_P8cvXJkE8_1),.din(w_dff_A_XaHotoUV6_1),.clk(gclk));
	jdff dff_A_pWYZLlQF0_1(.dout(w_dff_A_XaHotoUV6_1),.din(w_dff_A_pWYZLlQF0_1),.clk(gclk));
	jdff dff_A_CDoiX9gV3_1(.dout(w_dff_A_pWYZLlQF0_1),.din(w_dff_A_CDoiX9gV3_1),.clk(gclk));
	jdff dff_A_Uz2qX9xz4_1(.dout(w_dff_A_CDoiX9gV3_1),.din(w_dff_A_Uz2qX9xz4_1),.clk(gclk));
	jdff dff_A_TJQ3WB8z4_1(.dout(w_dff_A_Uz2qX9xz4_1),.din(w_dff_A_TJQ3WB8z4_1),.clk(gclk));
	jdff dff_A_IBug5IEA4_0(.dout(w_n111_0[0]),.din(w_dff_A_IBug5IEA4_0),.clk(gclk));
	jdff dff_A_XbEjRKiI4_0(.dout(w_dff_A_IBug5IEA4_0),.din(w_dff_A_XbEjRKiI4_0),.clk(gclk));
	jdff dff_A_yfToKdmr0_0(.dout(w_dff_A_XbEjRKiI4_0),.din(w_dff_A_yfToKdmr0_0),.clk(gclk));
	jdff dff_A_D9WkKbMJ7_0(.dout(w_dff_A_yfToKdmr0_0),.din(w_dff_A_D9WkKbMJ7_0),.clk(gclk));
	jdff dff_A_HcECIPF01_0(.dout(w_dff_A_D9WkKbMJ7_0),.din(w_dff_A_HcECIPF01_0),.clk(gclk));
	jdff dff_A_5cnqSymo7_1(.dout(w_n111_0[1]),.din(w_dff_A_5cnqSymo7_1),.clk(gclk));
	jdff dff_A_NzIIuW7N3_1(.dout(w_dff_A_5cnqSymo7_1),.din(w_dff_A_NzIIuW7N3_1),.clk(gclk));
	jdff dff_A_2JJl2eq21_1(.dout(w_dff_A_NzIIuW7N3_1),.din(w_dff_A_2JJl2eq21_1),.clk(gclk));
	jdff dff_A_4oeNhO5j5_1(.dout(w_dff_A_2JJl2eq21_1),.din(w_dff_A_4oeNhO5j5_1),.clk(gclk));
	jdff dff_A_P6dePn5q4_1(.dout(w_dff_A_4oeNhO5j5_1),.din(w_dff_A_P6dePn5q4_1),.clk(gclk));
	jdff dff_A_U1uDaDXn2_0(.dout(w_n109_0[0]),.din(w_dff_A_U1uDaDXn2_0),.clk(gclk));
	jdff dff_A_9I7aLvHq1_0(.dout(w_dff_A_U1uDaDXn2_0),.din(w_dff_A_9I7aLvHq1_0),.clk(gclk));
	jdff dff_A_xzHN8wSu2_0(.dout(w_dff_A_9I7aLvHq1_0),.din(w_dff_A_xzHN8wSu2_0),.clk(gclk));
	jdff dff_A_tq3evxCx6_1(.dout(w_n109_0[1]),.din(w_dff_A_tq3evxCx6_1),.clk(gclk));
	jdff dff_B_pd0qDGl43_0(.din(n107),.dout(w_dff_B_pd0qDGl43_0),.clk(gclk));
	jdff dff_B_DKTaPvg74_1(.din(n102),.dout(w_dff_B_DKTaPvg74_1),.clk(gclk));
	jdff dff_A_U2ppfvjE4_1(.dout(w_G224_0[1]),.din(w_dff_A_U2ppfvjE4_1),.clk(gclk));
	jdff dff_A_5ITBupW48_1(.dout(w_n101_0[1]),.din(w_dff_A_5ITBupW48_1),.clk(gclk));
	jdff dff_A_AJUc31BI1_1(.dout(w_dff_A_5ITBupW48_1),.din(w_dff_A_AJUc31BI1_1),.clk(gclk));
	jdff dff_A_7MlgHC1q0_1(.dout(w_dff_A_AJUc31BI1_1),.din(w_dff_A_7MlgHC1q0_1),.clk(gclk));
	jdff dff_A_oBrJVQhk2_1(.dout(w_dff_A_7MlgHC1q0_1),.din(w_dff_A_oBrJVQhk2_1),.clk(gclk));
	jdff dff_A_LapVrmbC6_1(.dout(w_dff_A_oBrJVQhk2_1),.din(w_dff_A_LapVrmbC6_1),.clk(gclk));
	jdff dff_A_QykndE3a9_1(.dout(w_dff_A_LapVrmbC6_1),.din(w_dff_A_QykndE3a9_1),.clk(gclk));
	jdff dff_A_kHIeJ6Uj7_1(.dout(w_dff_A_QykndE3a9_1),.din(w_dff_A_kHIeJ6Uj7_1),.clk(gclk));
	jdff dff_A_YYyDqyYz5_1(.dout(w_dff_A_kHIeJ6Uj7_1),.din(w_dff_A_YYyDqyYz5_1),.clk(gclk));
	jdff dff_A_sBGeQd331_1(.dout(w_dff_A_YYyDqyYz5_1),.din(w_dff_A_sBGeQd331_1),.clk(gclk));
	jdff dff_A_7w5DLCYU4_1(.dout(w_dff_A_sBGeQd331_1),.din(w_dff_A_7w5DLCYU4_1),.clk(gclk));
	jdff dff_A_U2HY2R2g0_1(.dout(w_dff_A_7w5DLCYU4_1),.din(w_dff_A_U2HY2R2g0_1),.clk(gclk));
	jdff dff_B_1gtld1Sf8_0(.din(n100),.dout(w_dff_B_1gtld1Sf8_0),.clk(gclk));
	jdff dff_A_Ui9PJ5O17_1(.dout(w_G122_1[1]),.din(w_dff_A_Ui9PJ5O17_1),.clk(gclk));
	jdff dff_A_iohcq6jF2_1(.dout(w_G122_0[1]),.din(w_dff_A_iohcq6jF2_1),.clk(gclk));
	jdff dff_A_s5LjUzUz6_1(.dout(w_dff_A_iohcq6jF2_1),.din(w_dff_A_s5LjUzUz6_1),.clk(gclk));
	jdff dff_A_05OadJCG7_1(.dout(w_dff_A_s5LjUzUz6_1),.din(w_dff_A_05OadJCG7_1),.clk(gclk));
	jdff dff_A_vD5CDa2t9_1(.dout(w_dff_A_05OadJCG7_1),.din(w_dff_A_vD5CDa2t9_1),.clk(gclk));
	jdff dff_A_cyhc6bz82_1(.dout(w_dff_A_vD5CDa2t9_1),.din(w_dff_A_cyhc6bz82_1),.clk(gclk));
	jdff dff_A_jXYcU6KF0_1(.dout(w_dff_A_cyhc6bz82_1),.din(w_dff_A_jXYcU6KF0_1),.clk(gclk));
	jdff dff_A_dUMFPHWU8_1(.dout(w_dff_A_jXYcU6KF0_1),.din(w_dff_A_dUMFPHWU8_1),.clk(gclk));
	jdff dff_A_WEugoDzi0_1(.dout(w_dff_A_dUMFPHWU8_1),.din(w_dff_A_WEugoDzi0_1),.clk(gclk));
	jdff dff_A_FW6HIXuH1_1(.dout(w_dff_A_WEugoDzi0_1),.din(w_dff_A_FW6HIXuH1_1),.clk(gclk));
	jdff dff_A_lbkTf7lM7_1(.dout(w_dff_A_FW6HIXuH1_1),.din(w_dff_A_lbkTf7lM7_1),.clk(gclk));
	jdff dff_A_ttOo4taJ6_1(.dout(w_dff_A_lbkTf7lM7_1),.din(w_dff_A_ttOo4taJ6_1),.clk(gclk));
	jdff dff_A_pYAaDC458_1(.dout(w_dff_A_ttOo4taJ6_1),.din(w_dff_A_pYAaDC458_1),.clk(gclk));
	jdff dff_A_1kv7ps4W5_0(.dout(w_G107_0[0]),.din(w_dff_A_1kv7ps4W5_0),.clk(gclk));
	jdff dff_A_bVhzwMjI8_0(.dout(w_dff_A_1kv7ps4W5_0),.din(w_dff_A_bVhzwMjI8_0),.clk(gclk));
	jdff dff_A_oySK6syp2_0(.dout(w_dff_A_bVhzwMjI8_0),.din(w_dff_A_oySK6syp2_0),.clk(gclk));
	jdff dff_A_qACBYdFH4_0(.dout(w_dff_A_oySK6syp2_0),.din(w_dff_A_qACBYdFH4_0),.clk(gclk));
	jdff dff_A_7xFuLcjY5_0(.dout(w_dff_A_qACBYdFH4_0),.din(w_dff_A_7xFuLcjY5_0),.clk(gclk));
	jdff dff_A_jlbDLggY5_0(.dout(w_dff_A_7xFuLcjY5_0),.din(w_dff_A_jlbDLggY5_0),.clk(gclk));
	jdff dff_A_BaMYHZHI9_0(.dout(w_dff_A_jlbDLggY5_0),.din(w_dff_A_BaMYHZHI9_0),.clk(gclk));
	jdff dff_A_GsL44PON1_0(.dout(w_dff_A_BaMYHZHI9_0),.din(w_dff_A_GsL44PON1_0),.clk(gclk));
	jdff dff_A_NtxSgBHr6_0(.dout(w_dff_A_GsL44PON1_0),.din(w_dff_A_NtxSgBHr6_0),.clk(gclk));
	jdff dff_A_fIKNUMVk9_0(.dout(w_dff_A_NtxSgBHr6_0),.din(w_dff_A_fIKNUMVk9_0),.clk(gclk));
	jdff dff_A_mvQDJjhl0_0(.dout(w_dff_A_fIKNUMVk9_0),.din(w_dff_A_mvQDJjhl0_0),.clk(gclk));
	jdff dff_A_lFGwgagg5_1(.dout(w_G107_0[1]),.din(w_dff_A_lFGwgagg5_1),.clk(gclk));
	jdff dff_A_QcNN8d9r8_0(.dout(w_G104_0[0]),.din(w_dff_A_QcNN8d9r8_0),.clk(gclk));
	jdff dff_A_D8YtNXkA7_0(.dout(w_dff_A_QcNN8d9r8_0),.din(w_dff_A_D8YtNXkA7_0),.clk(gclk));
	jdff dff_A_a3NvIrc59_0(.dout(w_dff_A_D8YtNXkA7_0),.din(w_dff_A_a3NvIrc59_0),.clk(gclk));
	jdff dff_A_HNJ7I9yW0_0(.dout(w_dff_A_a3NvIrc59_0),.din(w_dff_A_HNJ7I9yW0_0),.clk(gclk));
	jdff dff_A_lkvy8Bwq1_0(.dout(w_dff_A_HNJ7I9yW0_0),.din(w_dff_A_lkvy8Bwq1_0),.clk(gclk));
	jdff dff_A_WDfWyDR46_0(.dout(w_dff_A_lkvy8Bwq1_0),.din(w_dff_A_WDfWyDR46_0),.clk(gclk));
	jdff dff_A_bG1umpQW1_0(.dout(w_dff_A_WDfWyDR46_0),.din(w_dff_A_bG1umpQW1_0),.clk(gclk));
	jdff dff_A_K9TOOPpx4_0(.dout(w_dff_A_bG1umpQW1_0),.din(w_dff_A_K9TOOPpx4_0),.clk(gclk));
	jdff dff_A_IrIcfeQV9_0(.dout(w_dff_A_K9TOOPpx4_0),.din(w_dff_A_IrIcfeQV9_0),.clk(gclk));
	jdff dff_A_oTFCBXD72_0(.dout(w_dff_A_IrIcfeQV9_0),.din(w_dff_A_oTFCBXD72_0),.clk(gclk));
	jdff dff_A_ryt0mnN75_0(.dout(w_dff_A_oTFCBXD72_0),.din(w_dff_A_ryt0mnN75_0),.clk(gclk));
	jdff dff_A_NC3t7dCW0_1(.dout(w_G104_0[1]),.din(w_dff_A_NC3t7dCW0_1),.clk(gclk));
	jdff dff_A_WBnHEDFy2_1(.dout(w_n96_0[1]),.din(w_dff_A_WBnHEDFy2_1),.clk(gclk));
	jdff dff_A_BSyXgYxY5_1(.dout(w_dff_A_WBnHEDFy2_1),.din(w_dff_A_BSyXgYxY5_1),.clk(gclk));
	jdff dff_A_uEvwOPuB5_0(.dout(w_n59_1[0]),.din(w_dff_A_uEvwOPuB5_0),.clk(gclk));
	jdff dff_A_pCNrg0vZ5_0(.dout(w_dff_A_uEvwOPuB5_0),.din(w_dff_A_pCNrg0vZ5_0),.clk(gclk));
	jdff dff_A_Q2jMbFOm1_0(.dout(w_dff_A_pCNrg0vZ5_0),.din(w_dff_A_Q2jMbFOm1_0),.clk(gclk));
	jdff dff_A_3YgReqlg4_1(.dout(w_n59_1[1]),.din(w_dff_A_3YgReqlg4_1),.clk(gclk));
	jdff dff_A_8ddO8xqX1_1(.dout(w_dff_A_3YgReqlg4_1),.din(w_dff_A_8ddO8xqX1_1),.clk(gclk));
	jdff dff_A_ftWgLyG90_1(.dout(w_dff_A_8ddO8xqX1_1),.din(w_dff_A_ftWgLyG90_1),.clk(gclk));
	jdff dff_A_pudfbXUd3_1(.dout(w_dff_A_ftWgLyG90_1),.din(w_dff_A_pudfbXUd3_1),.clk(gclk));
	jdff dff_A_1rOVvtp43_1(.dout(w_G214_0[1]),.din(w_dff_A_1rOVvtp43_1),.clk(gclk));
	jdff dff_A_npsImUZ42_1(.dout(w_dff_A_1rOVvtp43_1),.din(w_dff_A_npsImUZ42_1),.clk(gclk));
	jdff dff_B_VME5RSDq1_2(.din(G214),.dout(w_dff_B_VME5RSDq1_2),.clk(gclk));
	jdff dff_A_UUgdfLni5_2(.dout(w_n93_0[2]),.din(w_dff_A_UUgdfLni5_2),.clk(gclk));
	jdff dff_A_giDHr2hO0_2(.dout(w_dff_A_UUgdfLni5_2),.din(w_dff_A_giDHr2hO0_2),.clk(gclk));
	jdff dff_A_2xbg2hI77_0(.dout(w_n90_0[0]),.din(w_dff_A_2xbg2hI77_0),.clk(gclk));
	jdff dff_A_gKwlaWvY7_0(.dout(w_dff_A_2xbg2hI77_0),.din(w_dff_A_gKwlaWvY7_0),.clk(gclk));
	jdff dff_A_6wOHC4WP1_0(.dout(w_dff_A_gKwlaWvY7_0),.din(w_dff_A_6wOHC4WP1_0),.clk(gclk));
	jdff dff_A_5FM4vTTV2_0(.dout(w_dff_A_6wOHC4WP1_0),.din(w_dff_A_5FM4vTTV2_0),.clk(gclk));
	jdff dff_A_l1t6oyFZ3_0(.dout(w_dff_A_5FM4vTTV2_0),.din(w_dff_A_l1t6oyFZ3_0),.clk(gclk));
	jdff dff_A_ffJhr80R9_0(.dout(w_dff_A_l1t6oyFZ3_0),.din(w_dff_A_ffJhr80R9_0),.clk(gclk));
	jdff dff_A_AkhowQR99_0(.dout(w_dff_A_ffJhr80R9_0),.din(w_dff_A_AkhowQR99_0),.clk(gclk));
	jdff dff_A_MXEDLgJw5_0(.dout(w_dff_A_AkhowQR99_0),.din(w_dff_A_MXEDLgJw5_0),.clk(gclk));
	jdff dff_A_Y0C9aZBy3_0(.dout(w_G210_0[0]),.din(w_dff_A_Y0C9aZBy3_0),.clk(gclk));
	jdff dff_A_1qEgt9xC6_0(.dout(w_dff_A_Y0C9aZBy3_0),.din(w_dff_A_1qEgt9xC6_0),.clk(gclk));
	jdff dff_A_AhPFVJ2L0_0(.dout(w_dff_A_1qEgt9xC6_0),.din(w_dff_A_AhPFVJ2L0_0),.clk(gclk));
	jdff dff_A_gyPgl8wT6_0(.dout(w_dff_A_AhPFVJ2L0_0),.din(w_dff_A_gyPgl8wT6_0),.clk(gclk));
	jdff dff_A_5RNRl6Vb1_0(.dout(w_dff_A_gyPgl8wT6_0),.din(w_dff_A_5RNRl6Vb1_0),.clk(gclk));
	jdff dff_A_IeQ2PzdK7_0(.dout(w_dff_A_5RNRl6Vb1_0),.din(w_dff_A_IeQ2PzdK7_0),.clk(gclk));
	jdff dff_A_fYHZdvQU1_0(.dout(w_dff_A_IeQ2PzdK7_0),.din(w_dff_A_fYHZdvQU1_0),.clk(gclk));
	jdff dff_A_LIZk3YRo9_0(.dout(w_dff_A_fYHZdvQU1_0),.din(w_dff_A_LIZk3YRo9_0),.clk(gclk));
	jdff dff_A_3Myj1NgY5_0(.dout(w_dff_A_LIZk3YRo9_0),.din(w_dff_A_3Myj1NgY5_0),.clk(gclk));
	jdff dff_A_UoXBNYhe1_0(.dout(w_dff_A_3Myj1NgY5_0),.din(w_dff_A_UoXBNYhe1_0),.clk(gclk));
	jdff dff_A_u0r9HC9p1_0(.dout(w_dff_A_UoXBNYhe1_0),.din(w_dff_A_u0r9HC9p1_0),.clk(gclk));
	jdff dff_A_t6o6BoYO8_1(.dout(w_G210_0[1]),.din(w_dff_A_t6o6BoYO8_1),.clk(gclk));
	jdff dff_A_cSU03OiF5_1(.dout(w_dff_A_t6o6BoYO8_1),.din(w_dff_A_cSU03OiF5_1),.clk(gclk));
	jdff dff_B_5KcbtH9R0_3(.din(G210),.dout(w_dff_B_5KcbtH9R0_3),.clk(gclk));
	jdff dff_A_2RV8VcwV1_0(.dout(w_n85_0[0]),.din(w_dff_A_2RV8VcwV1_0),.clk(gclk));
	jdff dff_A_KrZ6EOnd6_2(.dout(w_n85_0[2]),.din(w_dff_A_KrZ6EOnd6_2),.clk(gclk));
	jdff dff_A_eRzN8rTf6_0(.dout(w_G101_0[0]),.din(w_dff_A_eRzN8rTf6_0),.clk(gclk));
	jdff dff_A_AwgT4ywJ4_0(.dout(w_dff_A_eRzN8rTf6_0),.din(w_dff_A_AwgT4ywJ4_0),.clk(gclk));
	jdff dff_A_IyPAJ7Mx6_0(.dout(w_dff_A_AwgT4ywJ4_0),.din(w_dff_A_IyPAJ7Mx6_0),.clk(gclk));
	jdff dff_A_nhBxEeyT8_0(.dout(w_dff_A_IyPAJ7Mx6_0),.din(w_dff_A_nhBxEeyT8_0),.clk(gclk));
	jdff dff_A_fVJcP9a34_0(.dout(w_dff_A_nhBxEeyT8_0),.din(w_dff_A_fVJcP9a34_0),.clk(gclk));
	jdff dff_A_Y9wtmFol1_0(.dout(w_dff_A_fVJcP9a34_0),.din(w_dff_A_Y9wtmFol1_0),.clk(gclk));
	jdff dff_A_cmXUqGba9_0(.dout(w_dff_A_Y9wtmFol1_0),.din(w_dff_A_cmXUqGba9_0),.clk(gclk));
	jdff dff_A_kvPhKXs88_0(.dout(w_dff_A_cmXUqGba9_0),.din(w_dff_A_kvPhKXs88_0),.clk(gclk));
	jdff dff_A_5YaAlyT65_0(.dout(w_dff_A_kvPhKXs88_0),.din(w_dff_A_5YaAlyT65_0),.clk(gclk));
	jdff dff_A_OAHrCjFq3_0(.dout(w_dff_A_5YaAlyT65_0),.din(w_dff_A_OAHrCjFq3_0),.clk(gclk));
	jdff dff_A_vhETZMxO6_0(.dout(w_dff_A_OAHrCjFq3_0),.din(w_dff_A_vhETZMxO6_0),.clk(gclk));
	jdff dff_A_v7t7nDrW0_2(.dout(w_G101_0[2]),.din(w_dff_A_v7t7nDrW0_2),.clk(gclk));
	jdff dff_A_FtYLZEww0_2(.dout(w_dff_A_v7t7nDrW0_2),.din(w_dff_A_FtYLZEww0_2),.clk(gclk));
	jdff dff_B_y2ks6dKP9_3(.din(G101),.dout(w_dff_B_y2ks6dKP9_3),.clk(gclk));
	jdff dff_A_xxPCt6PZ4_1(.dout(w_n84_0[1]),.din(w_dff_A_xxPCt6PZ4_1),.clk(gclk));
	jdff dff_A_OwpnqkYD3_1(.dout(w_dff_A_xxPCt6PZ4_1),.din(w_dff_A_OwpnqkYD3_1),.clk(gclk));
	jdff dff_A_24rS6dwG1_0(.dout(w_G116_0[0]),.din(w_dff_A_24rS6dwG1_0),.clk(gclk));
	jdff dff_A_JuzkRHvL1_0(.dout(w_dff_A_24rS6dwG1_0),.din(w_dff_A_JuzkRHvL1_0),.clk(gclk));
	jdff dff_A_ndAlKMie2_0(.dout(w_dff_A_JuzkRHvL1_0),.din(w_dff_A_ndAlKMie2_0),.clk(gclk));
	jdff dff_A_dRQnyY7x9_0(.dout(w_dff_A_ndAlKMie2_0),.din(w_dff_A_dRQnyY7x9_0),.clk(gclk));
	jdff dff_A_teWS2zCG1_0(.dout(w_dff_A_dRQnyY7x9_0),.din(w_dff_A_teWS2zCG1_0),.clk(gclk));
	jdff dff_A_zf2SE4mo1_0(.dout(w_dff_A_teWS2zCG1_0),.din(w_dff_A_zf2SE4mo1_0),.clk(gclk));
	jdff dff_A_UcxAfrCR0_0(.dout(w_dff_A_zf2SE4mo1_0),.din(w_dff_A_UcxAfrCR0_0),.clk(gclk));
	jdff dff_A_f7rNHEMz5_0(.dout(w_dff_A_UcxAfrCR0_0),.din(w_dff_A_f7rNHEMz5_0),.clk(gclk));
	jdff dff_A_pluT9Enz8_0(.dout(w_dff_A_f7rNHEMz5_0),.din(w_dff_A_pluT9Enz8_0),.clk(gclk));
	jdff dff_A_OdM7OG2W7_0(.dout(w_dff_A_pluT9Enz8_0),.din(w_dff_A_OdM7OG2W7_0),.clk(gclk));
	jdff dff_A_MS1gN8KP4_0(.dout(w_dff_A_OdM7OG2W7_0),.din(w_dff_A_MS1gN8KP4_0),.clk(gclk));
	jdff dff_A_826U4WMO5_0(.dout(w_G113_0[0]),.din(w_dff_A_826U4WMO5_0),.clk(gclk));
	jdff dff_A_cAGfDvLN2_0(.dout(w_dff_A_826U4WMO5_0),.din(w_dff_A_cAGfDvLN2_0),.clk(gclk));
	jdff dff_A_e9SMnYKh6_0(.dout(w_dff_A_cAGfDvLN2_0),.din(w_dff_A_e9SMnYKh6_0),.clk(gclk));
	jdff dff_A_plsqT4a13_0(.dout(w_dff_A_e9SMnYKh6_0),.din(w_dff_A_plsqT4a13_0),.clk(gclk));
	jdff dff_A_VyfcBy0g6_0(.dout(w_dff_A_plsqT4a13_0),.din(w_dff_A_VyfcBy0g6_0),.clk(gclk));
	jdff dff_A_8hrwlRli4_0(.dout(w_dff_A_VyfcBy0g6_0),.din(w_dff_A_8hrwlRli4_0),.clk(gclk));
	jdff dff_A_ITTT5owe8_0(.dout(w_dff_A_8hrwlRli4_0),.din(w_dff_A_ITTT5owe8_0),.clk(gclk));
	jdff dff_A_u32QCrcr8_0(.dout(w_dff_A_ITTT5owe8_0),.din(w_dff_A_u32QCrcr8_0),.clk(gclk));
	jdff dff_A_ucaaQgz70_0(.dout(w_dff_A_u32QCrcr8_0),.din(w_dff_A_ucaaQgz70_0),.clk(gclk));
	jdff dff_A_XQT0xlrj6_0(.dout(w_dff_A_ucaaQgz70_0),.din(w_dff_A_XQT0xlrj6_0),.clk(gclk));
	jdff dff_A_BKpryq4U4_0(.dout(w_dff_A_XQT0xlrj6_0),.din(w_dff_A_BKpryq4U4_0),.clk(gclk));
	jdff dff_A_ZLODwrnj3_2(.dout(w_G113_0[2]),.din(w_dff_A_ZLODwrnj3_2),.clk(gclk));
	jdff dff_A_dZrJtdGE4_2(.dout(w_n82_0[2]),.din(w_dff_A_dZrJtdGE4_2),.clk(gclk));
	jdff dff_A_FWBvyt5U0_2(.dout(w_dff_A_dZrJtdGE4_2),.din(w_dff_A_FWBvyt5U0_2),.clk(gclk));
	jdff dff_A_s4MrnL4K3_0(.dout(w_G134_0[0]),.din(w_dff_A_s4MrnL4K3_0),.clk(gclk));
	jdff dff_A_cNSo23I08_0(.dout(w_dff_A_s4MrnL4K3_0),.din(w_dff_A_cNSo23I08_0),.clk(gclk));
	jdff dff_A_7tprLKZE3_0(.dout(w_dff_A_cNSo23I08_0),.din(w_dff_A_7tprLKZE3_0),.clk(gclk));
	jdff dff_A_WrPST0t00_0(.dout(w_dff_A_7tprLKZE3_0),.din(w_dff_A_WrPST0t00_0),.clk(gclk));
	jdff dff_A_tw4Tdoqw7_0(.dout(w_dff_A_WrPST0t00_0),.din(w_dff_A_tw4Tdoqw7_0),.clk(gclk));
	jdff dff_A_v1e3CKb47_0(.dout(w_dff_A_tw4Tdoqw7_0),.din(w_dff_A_v1e3CKb47_0),.clk(gclk));
	jdff dff_A_wd1xCyMQ7_0(.dout(w_dff_A_v1e3CKb47_0),.din(w_dff_A_wd1xCyMQ7_0),.clk(gclk));
	jdff dff_A_c2NcYIJT3_0(.dout(w_dff_A_wd1xCyMQ7_0),.din(w_dff_A_c2NcYIJT3_0),.clk(gclk));
	jdff dff_A_KQHvbKUM8_0(.dout(w_dff_A_c2NcYIJT3_0),.din(w_dff_A_KQHvbKUM8_0),.clk(gclk));
	jdff dff_A_QqfFmQx10_0(.dout(w_dff_A_KQHvbKUM8_0),.din(w_dff_A_QqfFmQx10_0),.clk(gclk));
	jdff dff_A_3HnYfHIg9_0(.dout(w_dff_A_QqfFmQx10_0),.din(w_dff_A_3HnYfHIg9_0),.clk(gclk));
	jdff dff_A_LZJINklu6_1(.dout(w_G134_0[1]),.din(w_dff_A_LZJINklu6_1),.clk(gclk));
	jdff dff_A_BRpmqw9O3_0(.dout(w_G131_0[0]),.din(w_dff_A_BRpmqw9O3_0),.clk(gclk));
	jdff dff_A_VVy7NlmP9_0(.dout(w_dff_A_BRpmqw9O3_0),.din(w_dff_A_VVy7NlmP9_0),.clk(gclk));
	jdff dff_A_QEeP222e7_0(.dout(w_dff_A_VVy7NlmP9_0),.din(w_dff_A_QEeP222e7_0),.clk(gclk));
	jdff dff_A_5WFHONCN6_0(.dout(w_dff_A_QEeP222e7_0),.din(w_dff_A_5WFHONCN6_0),.clk(gclk));
	jdff dff_A_BpoZLH6c1_0(.dout(w_dff_A_5WFHONCN6_0),.din(w_dff_A_BpoZLH6c1_0),.clk(gclk));
	jdff dff_A_oT5TMHdb4_0(.dout(w_dff_A_BpoZLH6c1_0),.din(w_dff_A_oT5TMHdb4_0),.clk(gclk));
	jdff dff_A_BKSBWluH8_0(.dout(w_dff_A_oT5TMHdb4_0),.din(w_dff_A_BKSBWluH8_0),.clk(gclk));
	jdff dff_A_RRv6MsYz4_0(.dout(w_dff_A_BKSBWluH8_0),.din(w_dff_A_RRv6MsYz4_0),.clk(gclk));
	jdff dff_A_WPsuIQJe9_0(.dout(w_dff_A_RRv6MsYz4_0),.din(w_dff_A_WPsuIQJe9_0),.clk(gclk));
	jdff dff_A_GyKhO8CR3_0(.dout(w_dff_A_WPsuIQJe9_0),.din(w_dff_A_GyKhO8CR3_0),.clk(gclk));
	jdff dff_A_kBvrLY7q2_0(.dout(w_dff_A_GyKhO8CR3_0),.din(w_dff_A_kBvrLY7q2_0),.clk(gclk));
	jdff dff_A_iuCcpqQN4_2(.dout(w_G131_0[2]),.din(w_dff_A_iuCcpqQN4_2),.clk(gclk));
	jdff dff_A_1SL49ZY94_0(.dout(w_G143_0[0]),.din(w_dff_A_1SL49ZY94_0),.clk(gclk));
	jdff dff_A_zctUQblE6_0(.dout(w_dff_A_1SL49ZY94_0),.din(w_dff_A_zctUQblE6_0),.clk(gclk));
	jdff dff_A_fxNmxl9i1_0(.dout(w_dff_A_zctUQblE6_0),.din(w_dff_A_fxNmxl9i1_0),.clk(gclk));
	jdff dff_A_dvabvz5G6_0(.dout(w_dff_A_fxNmxl9i1_0),.din(w_dff_A_dvabvz5G6_0),.clk(gclk));
	jdff dff_A_qNzGlO3j2_0(.dout(w_dff_A_dvabvz5G6_0),.din(w_dff_A_qNzGlO3j2_0),.clk(gclk));
	jdff dff_A_qRPjnq8j3_0(.dout(w_dff_A_qNzGlO3j2_0),.din(w_dff_A_qRPjnq8j3_0),.clk(gclk));
	jdff dff_A_CfQGplYX8_0(.dout(w_dff_A_qRPjnq8j3_0),.din(w_dff_A_CfQGplYX8_0),.clk(gclk));
	jdff dff_A_V6NZBuYY6_0(.dout(w_dff_A_CfQGplYX8_0),.din(w_dff_A_V6NZBuYY6_0),.clk(gclk));
	jdff dff_A_dSYd7Wko1_0(.dout(w_dff_A_V6NZBuYY6_0),.din(w_dff_A_dSYd7Wko1_0),.clk(gclk));
	jdff dff_A_UUIYuLPL5_0(.dout(w_dff_A_dSYd7Wko1_0),.din(w_dff_A_UUIYuLPL5_0),.clk(gclk));
	jdff dff_A_obgZl6jG1_0(.dout(w_dff_A_UUIYuLPL5_0),.din(w_dff_A_obgZl6jG1_0),.clk(gclk));
	jdff dff_A_GApTDjgN1_0(.dout(w_dff_A_obgZl6jG1_0),.din(w_dff_A_GApTDjgN1_0),.clk(gclk));
	jdff dff_A_SNBSiXTw9_0(.dout(w_G472_0[0]),.din(w_dff_A_SNBSiXTw9_0),.clk(gclk));
	jdff dff_A_VF7R0M0a8_0(.dout(w_dff_A_SNBSiXTw9_0),.din(w_dff_A_VF7R0M0a8_0),.clk(gclk));
	jdff dff_A_ZHudeNIm6_0(.dout(w_dff_A_VF7R0M0a8_0),.din(w_dff_A_ZHudeNIm6_0),.clk(gclk));
	jdff dff_A_DtPHaBP40_0(.dout(w_dff_A_ZHudeNIm6_0),.din(w_dff_A_DtPHaBP40_0),.clk(gclk));
	jdff dff_A_xo3NQvQi6_0(.dout(w_dff_A_DtPHaBP40_0),.din(w_dff_A_xo3NQvQi6_0),.clk(gclk));
	jdff dff_A_7ngWHTDD3_0(.dout(w_dff_A_xo3NQvQi6_0),.din(w_dff_A_7ngWHTDD3_0),.clk(gclk));
	jdff dff_A_qhxDTkZz0_0(.dout(w_dff_A_7ngWHTDD3_0),.din(w_dff_A_qhxDTkZz0_0),.clk(gclk));
	jdff dff_A_kFjFqPnk8_0(.dout(w_dff_A_qhxDTkZz0_0),.din(w_dff_A_kFjFqPnk8_0),.clk(gclk));
	jdff dff_A_WsLv4gx42_0(.dout(w_dff_A_kFjFqPnk8_0),.din(w_dff_A_WsLv4gx42_0),.clk(gclk));
	jdff dff_A_QCd9yhUo1_0(.dout(w_dff_A_WsLv4gx42_0),.din(w_dff_A_QCd9yhUo1_0),.clk(gclk));
	jdff dff_A_sXuUSNHX8_0(.dout(w_dff_A_QCd9yhUo1_0),.din(w_dff_A_sXuUSNHX8_0),.clk(gclk));
	jdff dff_A_FU9JAAiV3_0(.dout(w_dff_A_sXuUSNHX8_0),.din(w_dff_A_FU9JAAiV3_0),.clk(gclk));
	jdff dff_A_m7bR6HhP1_2(.dout(w_G472_0[2]),.din(w_dff_A_m7bR6HhP1_2),.clk(gclk));
	jdff dff_A_vALIWXhM6_2(.dout(w_dff_A_m7bR6HhP1_2),.din(w_dff_A_vALIWXhM6_2),.clk(gclk));
	jdff dff_A_cdvz8ir87_2(.dout(w_dff_A_vALIWXhM6_2),.din(w_dff_A_cdvz8ir87_2),.clk(gclk));
	jdff dff_A_QXjW7J0L2_2(.dout(w_dff_A_cdvz8ir87_2),.din(w_dff_A_QXjW7J0L2_2),.clk(gclk));
	jdff dff_A_OaL2mG203_2(.dout(w_dff_A_QXjW7J0L2_2),.din(w_dff_A_OaL2mG203_2),.clk(gclk));
	jdff dff_A_rmsSqK9p0_2(.dout(w_dff_A_OaL2mG203_2),.din(w_dff_A_rmsSqK9p0_2),.clk(gclk));
	jdff dff_A_ICOXnSjx7_2(.dout(w_dff_A_rmsSqK9p0_2),.din(w_dff_A_ICOXnSjx7_2),.clk(gclk));
	jdff dff_B_gC6kq2403_3(.din(n77),.dout(w_dff_B_gC6kq2403_3),.clk(gclk));
	jdff dff_B_8rLfO2R71_0(.din(n76),.dout(w_dff_B_8rLfO2R71_0),.clk(gclk));
	jdff dff_B_ahKLhWif8_0(.din(w_dff_B_8rLfO2R71_0),.dout(w_dff_B_ahKLhWif8_0),.clk(gclk));
	jdff dff_B_YYY2vQAx9_0(.din(w_dff_B_ahKLhWif8_0),.dout(w_dff_B_YYY2vQAx9_0),.clk(gclk));
	jdff dff_A_PxOqAoKK5_0(.dout(w_n75_0[0]),.din(w_dff_A_PxOqAoKK5_0),.clk(gclk));
	jdff dff_A_brUGOvlL4_0(.dout(w_dff_A_PxOqAoKK5_0),.din(w_dff_A_brUGOvlL4_0),.clk(gclk));
	jdff dff_A_KhHx9UBa5_0(.dout(w_dff_A_brUGOvlL4_0),.din(w_dff_A_KhHx9UBa5_0),.clk(gclk));
	jdff dff_A_Gxhitpy44_0(.dout(w_dff_A_KhHx9UBa5_0),.din(w_dff_A_Gxhitpy44_0),.clk(gclk));
	jdff dff_A_lIqe7Wt14_0(.dout(w_G217_0[0]),.din(w_dff_A_lIqe7Wt14_0),.clk(gclk));
	jdff dff_A_6xYUyHOP2_0(.dout(w_dff_A_lIqe7Wt14_0),.din(w_dff_A_6xYUyHOP2_0),.clk(gclk));
	jdff dff_A_z3pJz3030_0(.dout(w_dff_A_6xYUyHOP2_0),.din(w_dff_A_z3pJz3030_0),.clk(gclk));
	jdff dff_A_s2tO7NjE4_0(.dout(w_dff_A_z3pJz3030_0),.din(w_dff_A_s2tO7NjE4_0),.clk(gclk));
	jdff dff_A_ycnG1fB95_0(.dout(w_dff_A_s2tO7NjE4_0),.din(w_dff_A_ycnG1fB95_0),.clk(gclk));
	jdff dff_A_HTrla1TD9_0(.dout(w_dff_A_ycnG1fB95_0),.din(w_dff_A_HTrla1TD9_0),.clk(gclk));
	jdff dff_A_GH1zlFqY8_0(.dout(w_dff_A_HTrla1TD9_0),.din(w_dff_A_GH1zlFqY8_0),.clk(gclk));
	jdff dff_A_oCC99aW00_0(.dout(w_dff_A_GH1zlFqY8_0),.din(w_dff_A_oCC99aW00_0),.clk(gclk));
	jdff dff_A_Uvr7HL5t3_0(.dout(w_dff_A_oCC99aW00_0),.din(w_dff_A_Uvr7HL5t3_0),.clk(gclk));
	jdff dff_A_p7pPbWTJ5_0(.dout(w_dff_A_Uvr7HL5t3_0),.din(w_dff_A_p7pPbWTJ5_0),.clk(gclk));
	jdff dff_A_xxxnEkvb4_0(.dout(w_dff_A_p7pPbWTJ5_0),.din(w_dff_A_xxxnEkvb4_0),.clk(gclk));
	jdff dff_A_Gw1p1y5E4_0(.dout(w_dff_A_xxxnEkvb4_0),.din(w_dff_A_Gw1p1y5E4_0),.clk(gclk));
	jdff dff_A_gdmvXRrI7_2(.dout(w_G217_0[2]),.din(w_dff_A_gdmvXRrI7_2),.clk(gclk));
	jdff dff_A_UmtzS4231_0(.dout(w_n71_0[0]),.din(w_dff_A_UmtzS4231_0),.clk(gclk));
	jdff dff_A_jRr75Cmx9_0(.dout(w_dff_A_UmtzS4231_0),.din(w_dff_A_jRr75Cmx9_0),.clk(gclk));
	jdff dff_A_DAbspYrE9_0(.dout(w_dff_A_jRr75Cmx9_0),.din(w_dff_A_DAbspYrE9_0),.clk(gclk));
	jdff dff_A_9bilBzyQ2_0(.dout(w_dff_A_DAbspYrE9_0),.din(w_dff_A_9bilBzyQ2_0),.clk(gclk));
	jdff dff_A_wnx3vDL48_0(.dout(w_dff_A_9bilBzyQ2_0),.din(w_dff_A_wnx3vDL48_0),.clk(gclk));
	jdff dff_A_Jk449MZf5_0(.dout(w_dff_A_wnx3vDL48_0),.din(w_dff_A_Jk449MZf5_0),.clk(gclk));
	jdff dff_A_A92UaAXC8_0(.dout(w_dff_A_Jk449MZf5_0),.din(w_dff_A_A92UaAXC8_0),.clk(gclk));
	jdff dff_A_SlqB5pf85_0(.dout(w_dff_A_A92UaAXC8_0),.din(w_dff_A_SlqB5pf85_0),.clk(gclk));
	jdff dff_A_Pnv99A6v3_0(.dout(w_dff_A_SlqB5pf85_0),.din(w_dff_A_Pnv99A6v3_0),.clk(gclk));
	jdff dff_B_Ky51Spd31_1(.din(n64),.dout(w_dff_B_Ky51Spd31_1),.clk(gclk));
	jdff dff_A_GoMcK60a0_0(.dout(w_G119_0[0]),.din(w_dff_A_GoMcK60a0_0),.clk(gclk));
	jdff dff_A_ju48mgPi5_0(.dout(w_dff_A_GoMcK60a0_0),.din(w_dff_A_ju48mgPi5_0),.clk(gclk));
	jdff dff_A_5m1Idbjk0_0(.dout(w_dff_A_ju48mgPi5_0),.din(w_dff_A_5m1Idbjk0_0),.clk(gclk));
	jdff dff_A_aYGK7AyO5_0(.dout(w_dff_A_5m1Idbjk0_0),.din(w_dff_A_aYGK7AyO5_0),.clk(gclk));
	jdff dff_A_iJsy2A5X6_0(.dout(w_dff_A_aYGK7AyO5_0),.din(w_dff_A_iJsy2A5X6_0),.clk(gclk));
	jdff dff_A_p2O1MixS4_0(.dout(w_dff_A_iJsy2A5X6_0),.din(w_dff_A_p2O1MixS4_0),.clk(gclk));
	jdff dff_A_vallSv8x8_0(.dout(w_dff_A_p2O1MixS4_0),.din(w_dff_A_vallSv8x8_0),.clk(gclk));
	jdff dff_A_tBEckXBN3_0(.dout(w_dff_A_vallSv8x8_0),.din(w_dff_A_tBEckXBN3_0),.clk(gclk));
	jdff dff_A_0KZcFYYb5_0(.dout(w_dff_A_tBEckXBN3_0),.din(w_dff_A_0KZcFYYb5_0),.clk(gclk));
	jdff dff_A_mVMKXJXE7_0(.dout(w_dff_A_0KZcFYYb5_0),.din(w_dff_A_mVMKXJXE7_0),.clk(gclk));
	jdff dff_A_HCI87VPS2_0(.dout(w_dff_A_mVMKXJXE7_0),.din(w_dff_A_HCI87VPS2_0),.clk(gclk));
	jdff dff_A_mF7KzgY93_0(.dout(w_dff_A_HCI87VPS2_0),.din(w_dff_A_mF7KzgY93_0),.clk(gclk));
	jdff dff_A_SJxdXh8r0_2(.dout(w_G119_0[2]),.din(w_dff_A_SJxdXh8r0_2),.clk(gclk));
	jdff dff_A_FvvqJ0nI3_0(.dout(w_G110_0[0]),.din(w_dff_A_FvvqJ0nI3_0),.clk(gclk));
	jdff dff_A_e5vFrYof2_0(.dout(w_dff_A_FvvqJ0nI3_0),.din(w_dff_A_e5vFrYof2_0),.clk(gclk));
	jdff dff_A_4FSks8iq8_0(.dout(w_dff_A_e5vFrYof2_0),.din(w_dff_A_4FSks8iq8_0),.clk(gclk));
	jdff dff_A_xMSghTd98_0(.dout(w_dff_A_4FSks8iq8_0),.din(w_dff_A_xMSghTd98_0),.clk(gclk));
	jdff dff_A_N6Pb9mBT2_0(.dout(w_dff_A_xMSghTd98_0),.din(w_dff_A_N6Pb9mBT2_0),.clk(gclk));
	jdff dff_A_e31nRQDY6_0(.dout(w_dff_A_N6Pb9mBT2_0),.din(w_dff_A_e31nRQDY6_0),.clk(gclk));
	jdff dff_A_ghKRT1N76_0(.dout(w_dff_A_e31nRQDY6_0),.din(w_dff_A_ghKRT1N76_0),.clk(gclk));
	jdff dff_A_yTUZHwgc7_0(.dout(w_dff_A_ghKRT1N76_0),.din(w_dff_A_yTUZHwgc7_0),.clk(gclk));
	jdff dff_A_jTfhHgsa5_0(.dout(w_dff_A_yTUZHwgc7_0),.din(w_dff_A_jTfhHgsa5_0),.clk(gclk));
	jdff dff_A_vEr9B57F2_0(.dout(w_dff_A_jTfhHgsa5_0),.din(w_dff_A_vEr9B57F2_0),.clk(gclk));
	jdff dff_A_DSi8Rwoj8_0(.dout(w_dff_A_vEr9B57F2_0),.din(w_dff_A_DSi8Rwoj8_0),.clk(gclk));
	jdff dff_A_yilBa07N3_0(.dout(w_dff_A_DSi8Rwoj8_0),.din(w_dff_A_yilBa07N3_0),.clk(gclk));
	jdff dff_A_MJ3Mp4tL8_0(.dout(w_G128_0[0]),.din(w_dff_A_MJ3Mp4tL8_0),.clk(gclk));
	jdff dff_A_OeoskeEG5_0(.dout(w_dff_A_MJ3Mp4tL8_0),.din(w_dff_A_OeoskeEG5_0),.clk(gclk));
	jdff dff_A_Gz4AiwIu0_0(.dout(w_dff_A_OeoskeEG5_0),.din(w_dff_A_Gz4AiwIu0_0),.clk(gclk));
	jdff dff_A_llAGGRBC0_0(.dout(w_dff_A_Gz4AiwIu0_0),.din(w_dff_A_llAGGRBC0_0),.clk(gclk));
	jdff dff_A_8rGGDLr17_0(.dout(w_dff_A_llAGGRBC0_0),.din(w_dff_A_8rGGDLr17_0),.clk(gclk));
	jdff dff_A_GTo0dIFo7_0(.dout(w_dff_A_8rGGDLr17_0),.din(w_dff_A_GTo0dIFo7_0),.clk(gclk));
	jdff dff_A_ki44nNqs2_0(.dout(w_dff_A_GTo0dIFo7_0),.din(w_dff_A_ki44nNqs2_0),.clk(gclk));
	jdff dff_A_SVgvjFl49_0(.dout(w_dff_A_ki44nNqs2_0),.din(w_dff_A_SVgvjFl49_0),.clk(gclk));
	jdff dff_A_Rd0LLEzI0_0(.dout(w_dff_A_SVgvjFl49_0),.din(w_dff_A_Rd0LLEzI0_0),.clk(gclk));
	jdff dff_A_gEjCxq0P0_0(.dout(w_dff_A_Rd0LLEzI0_0),.din(w_dff_A_gEjCxq0P0_0),.clk(gclk));
	jdff dff_A_Uohm0taf4_0(.dout(w_dff_A_gEjCxq0P0_0),.din(w_dff_A_Uohm0taf4_0),.clk(gclk));
	jdff dff_A_kKbp1AZV4_2(.dout(w_G128_0[2]),.din(w_dff_A_kKbp1AZV4_2),.clk(gclk));
	jdff dff_A_G3lp0cUe0_2(.dout(w_dff_A_kKbp1AZV4_2),.din(w_dff_A_G3lp0cUe0_2),.clk(gclk));
	jdff dff_A_APhnHAiT2_0(.dout(w_n66_0[0]),.din(w_dff_A_APhnHAiT2_0),.clk(gclk));
	jdff dff_B_iPWazfDc1_2(.din(n66),.dout(w_dff_B_iPWazfDc1_2),.clk(gclk));
	jdff dff_A_RxTxGRxh9_0(.dout(w_n65_0[0]),.din(w_dff_A_RxTxGRxh9_0),.clk(gclk));
	jdff dff_A_K3IqHHkr1_0(.dout(w_dff_A_RxTxGRxh9_0),.din(w_dff_A_K3IqHHkr1_0),.clk(gclk));
	jdff dff_A_KK7Kz5PD7_0(.dout(w_G140_0[0]),.din(w_dff_A_KK7Kz5PD7_0),.clk(gclk));
	jdff dff_A_oejqsVYU9_0(.dout(w_dff_A_KK7Kz5PD7_0),.din(w_dff_A_oejqsVYU9_0),.clk(gclk));
	jdff dff_A_2cgMUa5v4_0(.dout(w_dff_A_oejqsVYU9_0),.din(w_dff_A_2cgMUa5v4_0),.clk(gclk));
	jdff dff_A_96TMQNo51_0(.dout(w_dff_A_2cgMUa5v4_0),.din(w_dff_A_96TMQNo51_0),.clk(gclk));
	jdff dff_A_4tSXdq7W5_0(.dout(w_dff_A_96TMQNo51_0),.din(w_dff_A_4tSXdq7W5_0),.clk(gclk));
	jdff dff_A_djmY2uR50_0(.dout(w_dff_A_4tSXdq7W5_0),.din(w_dff_A_djmY2uR50_0),.clk(gclk));
	jdff dff_A_hajWMwuI4_0(.dout(w_dff_A_djmY2uR50_0),.din(w_dff_A_hajWMwuI4_0),.clk(gclk));
	jdff dff_A_2yLr4S3i8_0(.dout(w_dff_A_hajWMwuI4_0),.din(w_dff_A_2yLr4S3i8_0),.clk(gclk));
	jdff dff_A_ZZH3glHj2_0(.dout(w_dff_A_2yLr4S3i8_0),.din(w_dff_A_ZZH3glHj2_0),.clk(gclk));
	jdff dff_A_vxEeDK438_0(.dout(w_dff_A_ZZH3glHj2_0),.din(w_dff_A_vxEeDK438_0),.clk(gclk));
	jdff dff_A_NKLohOZ70_0(.dout(w_dff_A_vxEeDK438_0),.din(w_dff_A_NKLohOZ70_0),.clk(gclk));
	jdff dff_A_IsyiABwm5_0(.dout(w_dff_A_NKLohOZ70_0),.din(w_dff_A_IsyiABwm5_0),.clk(gclk));
	jdff dff_A_0Lst71Nm1_0(.dout(w_G125_0[0]),.din(w_dff_A_0Lst71Nm1_0),.clk(gclk));
	jdff dff_A_t18dTeM72_0(.dout(w_dff_A_0Lst71Nm1_0),.din(w_dff_A_t18dTeM72_0),.clk(gclk));
	jdff dff_A_kUW22AGN3_0(.dout(w_dff_A_t18dTeM72_0),.din(w_dff_A_kUW22AGN3_0),.clk(gclk));
	jdff dff_A_XKEZtip65_0(.dout(w_dff_A_kUW22AGN3_0),.din(w_dff_A_XKEZtip65_0),.clk(gclk));
	jdff dff_A_ByBdzqzV6_0(.dout(w_dff_A_XKEZtip65_0),.din(w_dff_A_ByBdzqzV6_0),.clk(gclk));
	jdff dff_A_6HEV8Rev6_0(.dout(w_dff_A_ByBdzqzV6_0),.din(w_dff_A_6HEV8Rev6_0),.clk(gclk));
	jdff dff_A_tU1wH5D77_0(.dout(w_dff_A_6HEV8Rev6_0),.din(w_dff_A_tU1wH5D77_0),.clk(gclk));
	jdff dff_A_V8DD8o0t6_0(.dout(w_dff_A_tU1wH5D77_0),.din(w_dff_A_V8DD8o0t6_0),.clk(gclk));
	jdff dff_A_Xeczaa3W7_0(.dout(w_dff_A_V8DD8o0t6_0),.din(w_dff_A_Xeczaa3W7_0),.clk(gclk));
	jdff dff_A_pUzB4IKe8_0(.dout(w_dff_A_Xeczaa3W7_0),.din(w_dff_A_pUzB4IKe8_0),.clk(gclk));
	jdff dff_A_AO7eyqxq1_0(.dout(w_dff_A_pUzB4IKe8_0),.din(w_dff_A_AO7eyqxq1_0),.clk(gclk));
	jdff dff_A_hAbroMB57_0(.dout(w_dff_A_AO7eyqxq1_0),.din(w_dff_A_hAbroMB57_0),.clk(gclk));
	jdff dff_A_Pstr7MMN1_1(.dout(w_G125_0[1]),.din(w_dff_A_Pstr7MMN1_1),.clk(gclk));
	jdff dff_A_AcWRQco98_1(.dout(w_dff_A_Pstr7MMN1_1),.din(w_dff_A_AcWRQco98_1),.clk(gclk));
	jdff dff_A_YA06VvK44_0(.dout(w_G146_0[0]),.din(w_dff_A_YA06VvK44_0),.clk(gclk));
	jdff dff_A_pXsO4R0K4_0(.dout(w_dff_A_YA06VvK44_0),.din(w_dff_A_pXsO4R0K4_0),.clk(gclk));
	jdff dff_A_eVl1fKW27_0(.dout(w_dff_A_pXsO4R0K4_0),.din(w_dff_A_eVl1fKW27_0),.clk(gclk));
	jdff dff_A_pyNQCoWl4_0(.dout(w_dff_A_eVl1fKW27_0),.din(w_dff_A_pyNQCoWl4_0),.clk(gclk));
	jdff dff_A_P1W2Ql8z9_0(.dout(w_dff_A_pyNQCoWl4_0),.din(w_dff_A_P1W2Ql8z9_0),.clk(gclk));
	jdff dff_A_e7zaB9HF0_0(.dout(w_dff_A_P1W2Ql8z9_0),.din(w_dff_A_e7zaB9HF0_0),.clk(gclk));
	jdff dff_A_K4dsJa0A9_0(.dout(w_dff_A_e7zaB9HF0_0),.din(w_dff_A_K4dsJa0A9_0),.clk(gclk));
	jdff dff_A_p9bIWyfp6_0(.dout(w_dff_A_K4dsJa0A9_0),.din(w_dff_A_p9bIWyfp6_0),.clk(gclk));
	jdff dff_A_62Ctg2Ne2_0(.dout(w_dff_A_p9bIWyfp6_0),.din(w_dff_A_62Ctg2Ne2_0),.clk(gclk));
	jdff dff_A_GFIt6KrB0_0(.dout(w_dff_A_62Ctg2Ne2_0),.din(w_dff_A_GFIt6KrB0_0),.clk(gclk));
	jdff dff_B_V41iQZ8u6_3(.din(G146),.dout(w_dff_B_V41iQZ8u6_3),.clk(gclk));
	jdff dff_B_C2m4WaSq7_1(.din(n60),.dout(w_dff_B_C2m4WaSq7_1),.clk(gclk));
	jdff dff_A_ni3v0n9z5_0(.dout(w_G221_0[0]),.din(w_dff_A_ni3v0n9z5_0),.clk(gclk));
	jdff dff_A_x4psjkTG0_0(.dout(w_G137_0[0]),.din(w_dff_A_x4psjkTG0_0),.clk(gclk));
	jdff dff_A_dfsJwcK68_0(.dout(w_dff_A_x4psjkTG0_0),.din(w_dff_A_dfsJwcK68_0),.clk(gclk));
	jdff dff_A_Uh9PD1Lh7_0(.dout(w_dff_A_dfsJwcK68_0),.din(w_dff_A_Uh9PD1Lh7_0),.clk(gclk));
	jdff dff_A_MflngdFi7_0(.dout(w_dff_A_Uh9PD1Lh7_0),.din(w_dff_A_MflngdFi7_0),.clk(gclk));
	jdff dff_A_KDUjAa3E2_0(.dout(w_dff_A_MflngdFi7_0),.din(w_dff_A_KDUjAa3E2_0),.clk(gclk));
	jdff dff_A_YFxe02qr7_0(.dout(w_dff_A_KDUjAa3E2_0),.din(w_dff_A_YFxe02qr7_0),.clk(gclk));
	jdff dff_A_Aie8JjQ77_0(.dout(w_dff_A_YFxe02qr7_0),.din(w_dff_A_Aie8JjQ77_0),.clk(gclk));
	jdff dff_A_Cr9nVUDA1_0(.dout(w_dff_A_Aie8JjQ77_0),.din(w_dff_A_Cr9nVUDA1_0),.clk(gclk));
	jdff dff_A_BrWIWytB0_0(.dout(w_dff_A_Cr9nVUDA1_0),.din(w_dff_A_BrWIWytB0_0),.clk(gclk));
	jdff dff_A_m8FNkz492_0(.dout(w_dff_A_BrWIWytB0_0),.din(w_dff_A_m8FNkz492_0),.clk(gclk));
	jdff dff_A_g5Yaeth48_0(.dout(w_dff_A_m8FNkz492_0),.din(w_dff_A_g5Yaeth48_0),.clk(gclk));
	jdff dff_A_iKE1LC3X9_0(.dout(w_dff_A_g5Yaeth48_0),.din(w_dff_A_iKE1LC3X9_0),.clk(gclk));
	jdff dff_A_tREwYbIJ1_0(.dout(w_n59_2[0]),.din(w_dff_A_tREwYbIJ1_0),.clk(gclk));
	jdff dff_A_GCmGLdxp6_1(.dout(w_n59_0[1]),.din(w_dff_A_GCmGLdxp6_1),.clk(gclk));
	jdff dff_A_6gcsZIfy2_1(.dout(w_dff_A_GCmGLdxp6_1),.din(w_dff_A_6gcsZIfy2_1),.clk(gclk));
	jdff dff_A_1z5eNIe28_1(.dout(w_dff_A_6gcsZIfy2_1),.din(w_dff_A_1z5eNIe28_1),.clk(gclk));
	jdff dff_A_1o9DG4HD1_1(.dout(w_dff_A_1z5eNIe28_1),.din(w_dff_A_1o9DG4HD1_1),.clk(gclk));
	jdff dff_A_slIohsjf2_2(.dout(w_n59_0[2]),.din(w_dff_A_slIohsjf2_2),.clk(gclk));
	jdff dff_A_PSGJPxpB0_2(.dout(w_dff_A_slIohsjf2_2),.din(w_dff_A_PSGJPxpB0_2),.clk(gclk));
	jdff dff_A_eOiVXpce8_2(.dout(w_dff_A_PSGJPxpB0_2),.din(w_dff_A_eOiVXpce8_2),.clk(gclk));
	jdff dff_A_pltyNh1r3_2(.dout(w_dff_A_eOiVXpce8_2),.din(w_dff_A_pltyNh1r3_2),.clk(gclk));
	jdff dff_A_SmRkh54p1_2(.dout(w_dff_A_pltyNh1r3_2),.din(w_dff_A_SmRkh54p1_2),.clk(gclk));
	jdff dff_A_hvpjNHhD4_0(.dout(w_G902_4[0]),.din(w_dff_A_hvpjNHhD4_0),.clk(gclk));
	jdff dff_A_FoTLtxJU6_0(.dout(w_dff_A_hvpjNHhD4_0),.din(w_dff_A_FoTLtxJU6_0),.clk(gclk));
	jdff dff_A_9gDH7QjS7_0(.dout(w_dff_A_FoTLtxJU6_0),.din(w_dff_A_9gDH7QjS7_0),.clk(gclk));
	jdff dff_A_STTiZQIw4_0(.dout(w_dff_A_9gDH7QjS7_0),.din(w_dff_A_STTiZQIw4_0),.clk(gclk));
	jdff dff_A_hC6Riofy9_0(.dout(w_dff_A_STTiZQIw4_0),.din(w_dff_A_hC6Riofy9_0),.clk(gclk));
	jdff dff_A_EenXafGX8_1(.dout(w_G902_4[1]),.din(w_dff_A_EenXafGX8_1),.clk(gclk));
	jdff dff_A_DixJRMo74_1(.dout(w_G902_1[1]),.din(w_dff_A_DixJRMo74_1),.clk(gclk));
	jdff dff_A_UQ5ELU4O9_1(.dout(w_dff_A_DixJRMo74_1),.din(w_dff_A_UQ5ELU4O9_1),.clk(gclk));
	jdff dff_A_OpYzNYPk9_1(.dout(w_dff_A_UQ5ELU4O9_1),.din(w_dff_A_OpYzNYPk9_1),.clk(gclk));
	jdff dff_A_DX1Jtd824_1(.dout(w_dff_A_OpYzNYPk9_1),.din(w_dff_A_DX1Jtd824_1),.clk(gclk));
	jdff dff_A_F2jV7Pd82_1(.dout(w_dff_A_DX1Jtd824_1),.din(w_dff_A_F2jV7Pd82_1),.clk(gclk));
	jdff dff_A_V6Xc0F5r1_1(.dout(w_dff_A_F2jV7Pd82_1),.din(w_dff_A_V6Xc0F5r1_1),.clk(gclk));
	jdff dff_A_55eobgb14_1(.dout(w_dff_A_V6Xc0F5r1_1),.din(w_dff_A_55eobgb14_1),.clk(gclk));
	jdff dff_A_jtykbg1A3_1(.dout(w_dff_A_55eobgb14_1),.din(w_dff_A_jtykbg1A3_1),.clk(gclk));
	jdff dff_A_ImdvI9Mn8_1(.dout(w_dff_A_jtykbg1A3_1),.din(w_dff_A_ImdvI9Mn8_1),.clk(gclk));
	jdff dff_A_YN775MRB6_1(.dout(w_dff_A_ImdvI9Mn8_1),.din(w_dff_A_YN775MRB6_1),.clk(gclk));
	jdff dff_A_jYiAAeD65_1(.dout(w_dff_A_YN775MRB6_1),.din(w_dff_A_jYiAAeD65_1),.clk(gclk));
	jdff dff_A_hL35ZfMB4_1(.dout(w_dff_A_jYiAAeD65_1),.din(w_dff_A_hL35ZfMB4_1),.clk(gclk));
	jdff dff_A_ZwwODbhB0_1(.dout(w_dff_A_hL35ZfMB4_1),.din(w_dff_A_ZwwODbhB0_1),.clk(gclk));
	jdff dff_A_zuPO9N7w4_2(.dout(w_G902_1[2]),.din(w_dff_A_zuPO9N7w4_2),.clk(gclk));
	jdff dff_A_730B2bu67_2(.dout(w_dff_A_zuPO9N7w4_2),.din(w_dff_A_730B2bu67_2),.clk(gclk));
	jdff dff_A_m7SLLc3W2_2(.dout(w_dff_A_730B2bu67_2),.din(w_dff_A_m7SLLc3W2_2),.clk(gclk));
	jdff dff_A_LUYkr2Q20_2(.dout(w_dff_A_m7SLLc3W2_2),.din(w_dff_A_LUYkr2Q20_2),.clk(gclk));
	jdff dff_A_NoRgml0h4_2(.dout(w_dff_A_LUYkr2Q20_2),.din(w_dff_A_NoRgml0h4_2),.clk(gclk));
	jdff dff_A_Lf0gwY4J0_2(.dout(w_dff_A_NoRgml0h4_2),.din(w_dff_A_Lf0gwY4J0_2),.clk(gclk));
	jdff dff_A_WZFxI3PM5_2(.dout(w_dff_A_Lf0gwY4J0_2),.din(w_dff_A_WZFxI3PM5_2),.clk(gclk));
	jdff dff_A_jIsy6JS41_2(.dout(w_dff_A_WZFxI3PM5_2),.din(w_dff_A_jIsy6JS41_2),.clk(gclk));
	jdff dff_A_gIGhulHP0_2(.dout(w_dff_A_jIsy6JS41_2),.din(w_dff_A_gIGhulHP0_2),.clk(gclk));
	jdff dff_A_uvdrltih3_2(.dout(w_dff_A_gIGhulHP0_2),.din(w_dff_A_uvdrltih3_2),.clk(gclk));
	jdff dff_A_PSf7OqsH6_2(.dout(w_dff_A_uvdrltih3_2),.din(w_dff_A_PSf7OqsH6_2),.clk(gclk));
	jdff dff_A_CxHygDJm3_2(.dout(w_dff_A_PSf7OqsH6_2),.din(w_dff_A_CxHygDJm3_2),.clk(gclk));
	jdff dff_A_w6irMycR8_2(.dout(w_dff_A_CxHygDJm3_2),.din(w_dff_A_w6irMycR8_2),.clk(gclk));
	jdff dff_A_VyAK8UQF8_2(.dout(w_G902_0[2]),.din(w_dff_A_VyAK8UQF8_2),.clk(gclk));
	jdff dff_A_kyALfS8y8_2(.dout(w_dff_A_VyAK8UQF8_2),.din(w_dff_A_kyALfS8y8_2),.clk(gclk));
	jdff dff_A_S93cdf7v1_0(.dout(w_n269_0[0]),.din(w_dff_A_S93cdf7v1_0),.clk(gclk));
	jdff dff_A_T6QzBcsh7_2(.dout(w_n269_0[2]),.din(w_dff_A_T6QzBcsh7_2),.clk(gclk));
	jdff dff_B_bSRuW6T07_3(.din(n269),.dout(w_dff_B_bSRuW6T07_3),.clk(gclk));
	jdff dff_B_QhVnIGew8_3(.din(w_dff_B_bSRuW6T07_3),.dout(w_dff_B_QhVnIGew8_3),.clk(gclk));
	jdff dff_B_tT049HkM7_3(.din(w_dff_B_QhVnIGew8_3),.dout(w_dff_B_tT049HkM7_3),.clk(gclk));
	jdff dff_B_0KDNIxUo6_3(.din(w_dff_B_tT049HkM7_3),.dout(w_dff_B_0KDNIxUo6_3),.clk(gclk));
	jdff dff_B_vs7CnyFM2_3(.din(w_dff_B_0KDNIxUo6_3),.dout(w_dff_B_vs7CnyFM2_3),.clk(gclk));
	jdff dff_B_Wg43Mll57_3(.din(w_dff_B_vs7CnyFM2_3),.dout(w_dff_B_Wg43Mll57_3),.clk(gclk));
	jdff dff_B_vwXDQ3k44_3(.din(w_dff_B_Wg43Mll57_3),.dout(w_dff_B_vwXDQ3k44_3),.clk(gclk));
	jdff dff_B_3rbTZAy59_3(.din(w_dff_B_vwXDQ3k44_3),.dout(w_dff_B_3rbTZAy59_3),.clk(gclk));
	jdff dff_B_3iUJite09_3(.din(w_dff_B_3rbTZAy59_3),.dout(w_dff_B_3iUJite09_3),.clk(gclk));
	jdff dff_B_OKuATHPp5_3(.din(w_dff_B_3iUJite09_3),.dout(w_dff_B_OKuATHPp5_3),.clk(gclk));
	jdff dff_B_D0uIuEKW5_3(.din(w_dff_B_OKuATHPp5_3),.dout(w_dff_B_D0uIuEKW5_3),.clk(gclk));
	jdff dff_B_4jiMGCk33_3(.din(w_dff_B_D0uIuEKW5_3),.dout(w_dff_B_4jiMGCk33_3),.clk(gclk));
	jdff dff_B_xMgHvZ9D3_3(.din(w_dff_B_4jiMGCk33_3),.dout(w_dff_B_xMgHvZ9D3_3),.clk(gclk));
	jdff dff_A_PhPMIR101_0(.dout(w_G953_3[0]),.din(w_dff_A_PhPMIR101_0),.clk(gclk));
	jdff dff_A_PE0GXOYn3_0(.dout(w_G953_0[0]),.din(w_dff_A_PE0GXOYn3_0),.clk(gclk));
	jdff dff_A_papfaKOE8_0(.dout(w_dff_A_PE0GXOYn3_0),.din(w_dff_A_papfaKOE8_0),.clk(gclk));
	jdff dff_A_m0CurfKx7_0(.dout(w_dff_A_papfaKOE8_0),.din(w_dff_A_m0CurfKx7_0),.clk(gclk));
	jdff dff_A_wQoLfVjt4_0(.dout(w_dff_A_m0CurfKx7_0),.din(w_dff_A_wQoLfVjt4_0),.clk(gclk));
	jdff dff_A_Jm8wX8NX2_0(.dout(w_dff_A_wQoLfVjt4_0),.din(w_dff_A_Jm8wX8NX2_0),.clk(gclk));
	jdff dff_A_1eKLivb79_0(.dout(w_dff_A_Jm8wX8NX2_0),.din(w_dff_A_1eKLivb79_0),.clk(gclk));
	jdff dff_A_yekxO9qK3_0(.dout(w_dff_A_1eKLivb79_0),.din(w_dff_A_yekxO9qK3_0),.clk(gclk));
	jdff dff_A_QxVqPfhw6_0(.dout(w_dff_A_yekxO9qK3_0),.din(w_dff_A_QxVqPfhw6_0),.clk(gclk));
	jdff dff_A_lZERSlmd7_0(.dout(w_dff_A_QxVqPfhw6_0),.din(w_dff_A_lZERSlmd7_0),.clk(gclk));
	jdff dff_A_zRhpTNeS3_0(.dout(w_dff_A_lZERSlmd7_0),.din(w_dff_A_zRhpTNeS3_0),.clk(gclk));
	jdff dff_A_YmhNpf6I9_0(.dout(w_dff_A_zRhpTNeS3_0),.din(w_dff_A_YmhNpf6I9_0),.clk(gclk));
	jdff dff_A_qLXv9ayE6_1(.dout(w_G953_0[1]),.din(w_dff_A_qLXv9ayE6_1),.clk(gclk));
	jdff dff_A_NFSuWSaA9_0(.dout(w_G952_0[0]),.din(w_dff_A_NFSuWSaA9_0),.clk(gclk));
	jdff dff_A_sm3iMdGl3_1(.dout(w_G952_0[1]),.din(w_dff_A_sm3iMdGl3_1),.clk(gclk));
	jdff dff_A_kqCYD7ff0_1(.dout(w_dff_A_sm3iMdGl3_1),.din(w_dff_A_kqCYD7ff0_1),.clk(gclk));
	jdff dff_A_LisM0hWW6_1(.dout(w_dff_A_kqCYD7ff0_1),.din(w_dff_A_LisM0hWW6_1),.clk(gclk));
	jdff dff_A_siV0kBdx2_1(.dout(w_dff_A_LisM0hWW6_1),.din(w_dff_A_siV0kBdx2_1),.clk(gclk));
	jdff dff_A_WCoM8kKN6_1(.dout(w_dff_A_siV0kBdx2_1),.din(w_dff_A_WCoM8kKN6_1),.clk(gclk));
	jdff dff_A_dDm8YGSF9_1(.dout(w_dff_A_WCoM8kKN6_1),.din(w_dff_A_dDm8YGSF9_1),.clk(gclk));
	jdff dff_A_IjUh3WNQ5_1(.dout(w_dff_A_dDm8YGSF9_1),.din(w_dff_A_IjUh3WNQ5_1),.clk(gclk));
	jdff dff_A_jgwiAHf38_1(.dout(w_dff_A_IjUh3WNQ5_1),.din(w_dff_A_jgwiAHf38_1),.clk(gclk));
	jdff dff_A_7Izl4Wsj3_1(.dout(w_dff_A_jgwiAHf38_1),.din(w_dff_A_7Izl4Wsj3_1),.clk(gclk));
	jdff dff_A_OeAHGV3d7_1(.dout(w_dff_A_7Izl4Wsj3_1),.din(w_dff_A_OeAHGV3d7_1),.clk(gclk));
	jdff dff_A_EkyAUfKq3_1(.dout(w_dff_A_OeAHGV3d7_1),.din(w_dff_A_EkyAUfKq3_1),.clk(gclk));
	jdff dff_A_YKAltODn9_1(.dout(w_dff_A_EkyAUfKq3_1),.din(w_dff_A_YKAltODn9_1),.clk(gclk));
	jdff dff_A_lX7bwFbg2_1(.dout(w_dff_A_YKAltODn9_1),.din(w_dff_A_lX7bwFbg2_1),.clk(gclk));
endmodule

