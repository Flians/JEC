// Benchmark "c6288" written by ABC on Thu May 07 10:17:59 2020

module c6288 ( 
    G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n86, n87, n88, n89, n90, n91, n92, n93, n94,
    n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n106, n107,
    n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n529, n530, n531, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
    n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
    n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
    n1583, n1584, n1585, n1586, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820;
  jand g0000(.dina(G273gat), .dinb(G1gat), .dout(G545gat));
  jand g0001(.dina(G290gat), .dinb(G18gat), .dout(n65));
  jand g0002(.dina(n65), .dinb(G545gat), .dout(n66));
  jnot g0003(.din(n66), .dout(n67));
  jnot g0004(.din(G18gat), .dout(n68));
  jnot g0005(.din(G273gat), .dout(n69));
  jcb  g0006(.dina(n69), .dinb(n68), .dout(n70));
  jnot g0007(.din(n70), .dout(n71));
  jand g0008(.dina(G290gat), .dinb(G1gat), .dout(n72));
  jcb  g0009(.dina(n72), .dinb(n71), .dout(n73));
  jand g0010(.dina(n73), .dinb(n67), .dout(G1581gat));
  jand g0011(.dina(G307gat), .dinb(G1gat), .dout(n75));
  jnot g0012(.din(n75), .dout(n76));
  jnot g0013(.din(G35gat), .dout(n77));
  jnot g0014(.din(G290gat), .dout(n78));
  jcb  g0015(.dina(n78), .dinb(n77), .dout(n79));
  jcb  g0016(.dina(n79), .dinb(n70), .dout(n80));
  jand g0017(.dina(G273gat), .dinb(G35gat), .dout(n81));
  jcb  g0018(.dina(n81), .dinb(n65), .dout(n82));
  jand g0019(.dina(n82), .dinb(n80), .dout(n83));
  jxor g0020(.dina(n83), .dinb(n67), .dout(n84));
  jxor g0021(.dina(n84), .dinb(n76), .dout(G1901gat));
  jand g0022(.dina(G324gat), .dinb(G1gat), .dout(n86));
  jnot g0023(.din(n86), .dout(n87));
  jcb  g0024(.dina(n83), .dinb(n66), .dout(n88));
  jcb  g0025(.dina(n84), .dinb(n75), .dout(n89));
  jand g0026(.dina(n89), .dinb(n88), .dout(n90));
  jand g0027(.dina(G307gat), .dinb(G18gat), .dout(n91));
  jnot g0028(.din(n91), .dout(n92));
  jnot g0029(.din(n80), .dout(n93));
  jcb  g0030(.dina(n69), .dinb(n77), .dout(n94));
  jnot g0031(.din(G52gat), .dout(n95));
  jcb  g0032(.dina(n78), .dinb(n95), .dout(n96));
  jcb  g0033(.dina(n96), .dinb(n94), .dout(n97));
  jand g0034(.dina(G290gat), .dinb(G35gat), .dout(n98));
  jand g0035(.dina(G273gat), .dinb(G52gat), .dout(n99));
  jcb  g0036(.dina(n99), .dinb(n98), .dout(n100));
  jand g0037(.dina(n100), .dinb(n97), .dout(n101));
  jxor g0038(.dina(n101), .dinb(n93), .dout(n102));
  jxor g0039(.dina(n102), .dinb(n92), .dout(n103));
  jxor g0040(.dina(n103), .dinb(n90), .dout(n104));
  jxor g0041(.dina(n104), .dinb(n87), .dout(G2223gat));
  jand g0042(.dina(G341gat), .dinb(G1gat), .dout(n106));
  jnot g0043(.din(n106), .dout(n107));
  jnot g0044(.din(n103), .dout(n108));
  jcb  g0045(.dina(n108), .dinb(n90), .dout(n109));
  jcb  g0046(.dina(n104), .dinb(n86), .dout(n110));
  jand g0047(.dina(n110), .dinb(n109), .dout(n111));
  jand g0048(.dina(G324gat), .dinb(G18gat), .dout(n112));
  jnot g0049(.din(n112), .dout(n113));
  jcb  g0050(.dina(n101), .dinb(n93), .dout(n114));
  jxor g0051(.dina(n101), .dinb(n80), .dout(n115));
  jcb  g0052(.dina(n115), .dinb(n91), .dout(n116));
  jand g0053(.dina(n116), .dinb(n114), .dout(n117));
  jand g0054(.dina(G307gat), .dinb(G35gat), .dout(n118));
  jnot g0055(.din(n118), .dout(n119));
  jnot g0056(.din(n97), .dout(n120));
  jand g0057(.dina(G290gat), .dinb(G69gat), .dout(n121));
  jand g0058(.dina(n121), .dinb(n99), .dout(n122));
  jnot g0059(.din(n122), .dout(n123));
  jand g0060(.dina(G290gat), .dinb(G52gat), .dout(n124));
  jand g0061(.dina(G273gat), .dinb(G69gat), .dout(n125));
  jcb  g0062(.dina(n125), .dinb(n124), .dout(n126));
  jand g0063(.dina(n126), .dinb(n123), .dout(n127));
  jxor g0064(.dina(n127), .dinb(n120), .dout(n128));
  jxor g0065(.dina(n128), .dinb(n119), .dout(n129));
  jnot g0066(.din(n129), .dout(n130));
  jxor g0067(.dina(n130), .dinb(n117), .dout(n131));
  jxor g0068(.dina(n131), .dinb(n113), .dout(n132));
  jxor g0069(.dina(n132), .dinb(n111), .dout(n133));
  jxor g0070(.dina(n133), .dinb(n107), .dout(G2548gat));
  jand g0071(.dina(G358gat), .dinb(G1gat), .dout(n135));
  jnot g0072(.din(n135), .dout(n136));
  jnot g0073(.din(n132), .dout(n137));
  jcb  g0074(.dina(n137), .dinb(n111), .dout(n138));
  jcb  g0075(.dina(n133), .dinb(n106), .dout(n139));
  jand g0076(.dina(n139), .dinb(n138), .dout(n140));
  jand g0077(.dina(G341gat), .dinb(G18gat), .dout(n141));
  jnot g0078(.din(n141), .dout(n142));
  jcb  g0079(.dina(n130), .dinb(n117), .dout(n143));
  jxor g0080(.dina(n129), .dinb(n117), .dout(n144));
  jcb  g0081(.dina(n144), .dinb(n112), .dout(n145));
  jand g0082(.dina(n145), .dinb(n143), .dout(n146));
  jand g0083(.dina(G324gat), .dinb(G35gat), .dout(n147));
  jnot g0084(.din(n147), .dout(n148));
  jcb  g0085(.dina(n127), .dinb(n120), .dout(n149));
  jnot g0086(.din(n149), .dout(n150));
  jand g0087(.dina(n128), .dinb(n119), .dout(n151));
  jcb  g0088(.dina(n151), .dinb(n150), .dout(n152));
  jand g0089(.dina(G307gat), .dinb(G52gat), .dout(n153));
  jnot g0090(.din(n153), .dout(n154));
  jand g0091(.dina(G290gat), .dinb(G86gat), .dout(n155));
  jand g0092(.dina(n155), .dinb(n125), .dout(n156));
  jnot g0093(.din(n156), .dout(n157));
  jand g0094(.dina(G273gat), .dinb(G86gat), .dout(n158));
  jcb  g0095(.dina(n158), .dinb(n121), .dout(n159));
  jand g0096(.dina(n159), .dinb(n157), .dout(n160));
  jxor g0097(.dina(n160), .dinb(n122), .dout(n161));
  jxor g0098(.dina(n161), .dinb(n154), .dout(n162));
  jxor g0099(.dina(n162), .dinb(n152), .dout(n163));
  jxor g0100(.dina(n163), .dinb(n148), .dout(n164));
  jnot g0101(.din(n164), .dout(n165));
  jxor g0102(.dina(n165), .dinb(n146), .dout(n166));
  jxor g0103(.dina(n166), .dinb(n142), .dout(n167));
  jxor g0104(.dina(n167), .dinb(n140), .dout(n168));
  jxor g0105(.dina(n168), .dinb(n136), .dout(G2877gat));
  jand g0106(.dina(G375gat), .dinb(G1gat), .dout(n170));
  jnot g0107(.din(n170), .dout(n171));
  jnot g0108(.din(n167), .dout(n172));
  jcb  g0109(.dina(n172), .dinb(n140), .dout(n173));
  jcb  g0110(.dina(n168), .dinb(n135), .dout(n174));
  jand g0111(.dina(n174), .dinb(n173), .dout(n175));
  jand g0112(.dina(G358gat), .dinb(G18gat), .dout(n176));
  jnot g0113(.din(n176), .dout(n177));
  jcb  g0114(.dina(n165), .dinb(n146), .dout(n178));
  jxor g0115(.dina(n164), .dinb(n146), .dout(n179));
  jcb  g0116(.dina(n179), .dinb(n141), .dout(n180));
  jand g0117(.dina(n180), .dinb(n178), .dout(n181));
  jand g0118(.dina(G341gat), .dinb(G35gat), .dout(n182));
  jnot g0119(.din(n182), .dout(n183));
  jand g0120(.dina(n162), .dinb(n152), .dout(n184));
  jand g0121(.dina(n163), .dinb(n148), .dout(n185));
  jcb  g0122(.dina(n185), .dinb(n184), .dout(n186));
  jand g0123(.dina(G324gat), .dinb(G52gat), .dout(n187));
  jnot g0124(.din(n187), .dout(n188));
  jnot g0125(.din(n160), .dout(n189));
  jand g0126(.dina(n189), .dinb(n123), .dout(n190));
  jand g0127(.dina(n161), .dinb(n154), .dout(n191));
  jcb  g0128(.dina(n191), .dinb(n190), .dout(n192));
  jand g0129(.dina(G307gat), .dinb(G69gat), .dout(n193));
  jnot g0130(.din(n193), .dout(n194));
  jand g0131(.dina(G290gat), .dinb(G103gat), .dout(n195));
  jand g0132(.dina(n195), .dinb(n158), .dout(n196));
  jnot g0133(.din(n196), .dout(n197));
  jand g0134(.dina(G273gat), .dinb(G103gat), .dout(n198));
  jcb  g0135(.dina(n198), .dinb(n155), .dout(n199));
  jand g0136(.dina(n199), .dinb(n197), .dout(n200));
  jxor g0137(.dina(n200), .dinb(n156), .dout(n201));
  jxor g0138(.dina(n201), .dinb(n194), .dout(n202));
  jxor g0139(.dina(n202), .dinb(n192), .dout(n203));
  jxor g0140(.dina(n203), .dinb(n188), .dout(n204));
  jxor g0141(.dina(n204), .dinb(n186), .dout(n205));
  jxor g0142(.dina(n205), .dinb(n183), .dout(n206));
  jnot g0143(.din(n206), .dout(n207));
  jxor g0144(.dina(n207), .dinb(n181), .dout(n208));
  jxor g0145(.dina(n208), .dinb(n177), .dout(n209));
  jxor g0146(.dina(n209), .dinb(n175), .dout(n210));
  jxor g0147(.dina(n210), .dinb(n171), .dout(G3211gat));
  jand g0148(.dina(G392gat), .dinb(G1gat), .dout(n212));
  jnot g0149(.din(n212), .dout(n213));
  jnot g0150(.din(n209), .dout(n214));
  jcb  g0151(.dina(n214), .dinb(n175), .dout(n215));
  jcb  g0152(.dina(n210), .dinb(n170), .dout(n216));
  jand g0153(.dina(n216), .dinb(n215), .dout(n217));
  jand g0154(.dina(G375gat), .dinb(G18gat), .dout(n218));
  jnot g0155(.din(n218), .dout(n219));
  jcb  g0156(.dina(n207), .dinb(n181), .dout(n220));
  jxor g0157(.dina(n206), .dinb(n181), .dout(n221));
  jcb  g0158(.dina(n221), .dinb(n176), .dout(n222));
  jand g0159(.dina(n222), .dinb(n220), .dout(n223));
  jand g0160(.dina(G358gat), .dinb(G35gat), .dout(n224));
  jnot g0161(.din(n224), .dout(n225));
  jand g0162(.dina(n204), .dinb(n186), .dout(n226));
  jand g0163(.dina(n205), .dinb(n183), .dout(n227));
  jcb  g0164(.dina(n227), .dinb(n226), .dout(n228));
  jand g0165(.dina(G341gat), .dinb(G52gat), .dout(n229));
  jnot g0166(.din(n229), .dout(n230));
  jand g0167(.dina(n202), .dinb(n192), .dout(n231));
  jand g0168(.dina(n203), .dinb(n188), .dout(n232));
  jcb  g0169(.dina(n232), .dinb(n231), .dout(n233));
  jand g0170(.dina(G324gat), .dinb(G69gat), .dout(n234));
  jnot g0171(.din(n234), .dout(n235));
  jnot g0172(.din(n200), .dout(n236));
  jand g0173(.dina(n236), .dinb(n157), .dout(n237));
  jand g0174(.dina(n201), .dinb(n194), .dout(n238));
  jcb  g0175(.dina(n238), .dinb(n237), .dout(n239));
  jand g0176(.dina(G307gat), .dinb(G86gat), .dout(n240));
  jnot g0177(.din(n240), .dout(n241));
  jand g0178(.dina(G290gat), .dinb(G120gat), .dout(n242));
  jand g0179(.dina(n242), .dinb(n198), .dout(n243));
  jnot g0180(.din(n243), .dout(n244));
  jand g0181(.dina(G273gat), .dinb(G120gat), .dout(n245));
  jcb  g0182(.dina(n245), .dinb(n195), .dout(n246));
  jand g0183(.dina(n246), .dinb(n244), .dout(n247));
  jxor g0184(.dina(n247), .dinb(n196), .dout(n248));
  jxor g0185(.dina(n248), .dinb(n241), .dout(n249));
  jxor g0186(.dina(n249), .dinb(n239), .dout(n250));
  jxor g0187(.dina(n250), .dinb(n235), .dout(n251));
  jxor g0188(.dina(n251), .dinb(n233), .dout(n252));
  jxor g0189(.dina(n252), .dinb(n230), .dout(n253));
  jxor g0190(.dina(n253), .dinb(n228), .dout(n254));
  jxor g0191(.dina(n254), .dinb(n225), .dout(n255));
  jnot g0192(.din(n255), .dout(n256));
  jxor g0193(.dina(n256), .dinb(n223), .dout(n257));
  jxor g0194(.dina(n257), .dinb(n219), .dout(n258));
  jxor g0195(.dina(n258), .dinb(n217), .dout(n259));
  jxor g0196(.dina(n259), .dinb(n213), .dout(G3552gat));
  jand g0197(.dina(G409gat), .dinb(G1gat), .dout(n261));
  jnot g0198(.din(n261), .dout(n262));
  jnot g0199(.din(n258), .dout(n263));
  jcb  g0200(.dina(n263), .dinb(n217), .dout(n264));
  jcb  g0201(.dina(n259), .dinb(n212), .dout(n265));
  jand g0202(.dina(n265), .dinb(n264), .dout(n266));
  jand g0203(.dina(G392gat), .dinb(G18gat), .dout(n267));
  jnot g0204(.din(n267), .dout(n268));
  jcb  g0205(.dina(n256), .dinb(n223), .dout(n269));
  jxor g0206(.dina(n255), .dinb(n223), .dout(n270));
  jcb  g0207(.dina(n270), .dinb(n218), .dout(n271));
  jand g0208(.dina(n271), .dinb(n269), .dout(n272));
  jand g0209(.dina(G375gat), .dinb(G35gat), .dout(n273));
  jnot g0210(.din(n273), .dout(n274));
  jand g0211(.dina(n253), .dinb(n228), .dout(n275));
  jand g0212(.dina(n254), .dinb(n225), .dout(n276));
  jcb  g0213(.dina(n276), .dinb(n275), .dout(n277));
  jand g0214(.dina(G358gat), .dinb(G52gat), .dout(n278));
  jnot g0215(.din(n278), .dout(n279));
  jand g0216(.dina(n251), .dinb(n233), .dout(n280));
  jand g0217(.dina(n252), .dinb(n230), .dout(n281));
  jcb  g0218(.dina(n281), .dinb(n280), .dout(n282));
  jand g0219(.dina(G341gat), .dinb(G69gat), .dout(n283));
  jnot g0220(.din(n283), .dout(n284));
  jand g0221(.dina(n249), .dinb(n239), .dout(n285));
  jand g0222(.dina(n250), .dinb(n235), .dout(n286));
  jcb  g0223(.dina(n286), .dinb(n285), .dout(n287));
  jand g0224(.dina(G324gat), .dinb(G86gat), .dout(n288));
  jnot g0225(.din(n288), .dout(n289));
  jcb  g0226(.dina(n247), .dinb(n196), .dout(n290));
  jnot g0227(.din(n290), .dout(n291));
  jand g0228(.dina(n248), .dinb(n241), .dout(n292));
  jcb  g0229(.dina(n292), .dinb(n291), .dout(n293));
  jand g0230(.dina(G307gat), .dinb(G103gat), .dout(n294));
  jnot g0231(.din(n294), .dout(n295));
  jand g0232(.dina(G290gat), .dinb(G137gat), .dout(n296));
  jand g0233(.dina(n296), .dinb(n245), .dout(n297));
  jnot g0234(.din(n297), .dout(n298));
  jand g0235(.dina(G273gat), .dinb(G137gat), .dout(n299));
  jcb  g0236(.dina(n299), .dinb(n242), .dout(n300));
  jand g0237(.dina(n300), .dinb(n298), .dout(n301));
  jxor g0238(.dina(n301), .dinb(n243), .dout(n302));
  jxor g0239(.dina(n302), .dinb(n295), .dout(n303));
  jxor g0240(.dina(n303), .dinb(n293), .dout(n304));
  jxor g0241(.dina(n304), .dinb(n289), .dout(n305));
  jxor g0242(.dina(n305), .dinb(n287), .dout(n306));
  jxor g0243(.dina(n306), .dinb(n284), .dout(n307));
  jxor g0244(.dina(n307), .dinb(n282), .dout(n308));
  jxor g0245(.dina(n308), .dinb(n279), .dout(n309));
  jxor g0246(.dina(n309), .dinb(n277), .dout(n310));
  jxor g0247(.dina(n310), .dinb(n274), .dout(n311));
  jnot g0248(.din(n311), .dout(n312));
  jxor g0249(.dina(n312), .dinb(n272), .dout(n313));
  jxor g0250(.dina(n313), .dinb(n268), .dout(n314));
  jxor g0251(.dina(n314), .dinb(n266), .dout(n315));
  jxor g0252(.dina(n315), .dinb(n262), .dout(G3895gat));
  jand g0253(.dina(G426gat), .dinb(G1gat), .dout(n317));
  jnot g0254(.din(n317), .dout(n318));
  jnot g0255(.din(n314), .dout(n319));
  jcb  g0256(.dina(n319), .dinb(n266), .dout(n320));
  jcb  g0257(.dina(n315), .dinb(n261), .dout(n321));
  jand g0258(.dina(n321), .dinb(n320), .dout(n322));
  jand g0259(.dina(G409gat), .dinb(G18gat), .dout(n323));
  jnot g0260(.din(n323), .dout(n324));
  jcb  g0261(.dina(n312), .dinb(n272), .dout(n325));
  jxor g0262(.dina(n311), .dinb(n272), .dout(n326));
  jcb  g0263(.dina(n326), .dinb(n267), .dout(n327));
  jand g0264(.dina(n327), .dinb(n325), .dout(n328));
  jand g0265(.dina(G392gat), .dinb(G35gat), .dout(n329));
  jnot g0266(.din(n329), .dout(n330));
  jand g0267(.dina(n309), .dinb(n277), .dout(n331));
  jand g0268(.dina(n310), .dinb(n274), .dout(n332));
  jcb  g0269(.dina(n332), .dinb(n331), .dout(n333));
  jand g0270(.dina(G375gat), .dinb(G52gat), .dout(n334));
  jnot g0271(.din(n334), .dout(n335));
  jand g0272(.dina(n307), .dinb(n282), .dout(n336));
  jand g0273(.dina(n308), .dinb(n279), .dout(n337));
  jcb  g0274(.dina(n337), .dinb(n336), .dout(n338));
  jand g0275(.dina(G358gat), .dinb(G69gat), .dout(n339));
  jnot g0276(.din(n339), .dout(n340));
  jand g0277(.dina(n305), .dinb(n287), .dout(n341));
  jand g0278(.dina(n306), .dinb(n284), .dout(n342));
  jcb  g0279(.dina(n342), .dinb(n341), .dout(n343));
  jand g0280(.dina(G341gat), .dinb(G86gat), .dout(n344));
  jnot g0281(.din(n344), .dout(n345));
  jand g0282(.dina(n303), .dinb(n293), .dout(n346));
  jand g0283(.dina(n304), .dinb(n289), .dout(n347));
  jcb  g0284(.dina(n347), .dinb(n346), .dout(n348));
  jand g0285(.dina(G324gat), .dinb(G103gat), .dout(n349));
  jnot g0286(.din(n349), .dout(n350));
  jcb  g0287(.dina(n301), .dinb(n243), .dout(n351));
  jnot g0288(.din(n351), .dout(n352));
  jand g0289(.dina(n302), .dinb(n295), .dout(n353));
  jcb  g0290(.dina(n353), .dinb(n352), .dout(n354));
  jand g0291(.dina(G307gat), .dinb(G120gat), .dout(n355));
  jnot g0292(.din(n355), .dout(n356));
  jand g0293(.dina(G290gat), .dinb(G154gat), .dout(n357));
  jand g0294(.dina(n357), .dinb(n299), .dout(n358));
  jnot g0295(.din(n358), .dout(n359));
  jand g0296(.dina(G273gat), .dinb(G154gat), .dout(n360));
  jcb  g0297(.dina(n360), .dinb(n296), .dout(n361));
  jand g0298(.dina(n361), .dinb(n359), .dout(n362));
  jxor g0299(.dina(n362), .dinb(n297), .dout(n363));
  jxor g0300(.dina(n363), .dinb(n356), .dout(n364));
  jxor g0301(.dina(n364), .dinb(n354), .dout(n365));
  jxor g0302(.dina(n365), .dinb(n350), .dout(n366));
  jxor g0303(.dina(n366), .dinb(n348), .dout(n367));
  jxor g0304(.dina(n367), .dinb(n345), .dout(n368));
  jxor g0305(.dina(n368), .dinb(n343), .dout(n369));
  jxor g0306(.dina(n369), .dinb(n340), .dout(n370));
  jxor g0307(.dina(n370), .dinb(n338), .dout(n371));
  jxor g0308(.dina(n371), .dinb(n335), .dout(n372));
  jxor g0309(.dina(n372), .dinb(n333), .dout(n373));
  jxor g0310(.dina(n373), .dinb(n330), .dout(n374));
  jnot g0311(.din(n374), .dout(n375));
  jxor g0312(.dina(n375), .dinb(n328), .dout(n376));
  jxor g0313(.dina(n376), .dinb(n324), .dout(n377));
  jxor g0314(.dina(n377), .dinb(n322), .dout(n378));
  jxor g0315(.dina(n378), .dinb(n318), .dout(G4241gat));
  jand g0316(.dina(G443gat), .dinb(G1gat), .dout(n380));
  jnot g0317(.din(n380), .dout(n381));
  jnot g0318(.din(n377), .dout(n382));
  jcb  g0319(.dina(n382), .dinb(n322), .dout(n383));
  jcb  g0320(.dina(n378), .dinb(n317), .dout(n384));
  jand g0321(.dina(n384), .dinb(n383), .dout(n385));
  jand g0322(.dina(G426gat), .dinb(G18gat), .dout(n386));
  jnot g0323(.din(n386), .dout(n387));
  jcb  g0324(.dina(n375), .dinb(n328), .dout(n388));
  jxor g0325(.dina(n374), .dinb(n328), .dout(n389));
  jcb  g0326(.dina(n389), .dinb(n323), .dout(n390));
  jand g0327(.dina(n390), .dinb(n388), .dout(n391));
  jand g0328(.dina(G409gat), .dinb(G35gat), .dout(n392));
  jnot g0329(.din(n392), .dout(n393));
  jand g0330(.dina(n372), .dinb(n333), .dout(n394));
  jand g0331(.dina(n373), .dinb(n330), .dout(n395));
  jcb  g0332(.dina(n395), .dinb(n394), .dout(n396));
  jand g0333(.dina(G392gat), .dinb(G52gat), .dout(n397));
  jnot g0334(.din(n397), .dout(n398));
  jand g0335(.dina(n370), .dinb(n338), .dout(n399));
  jand g0336(.dina(n371), .dinb(n335), .dout(n400));
  jcb  g0337(.dina(n400), .dinb(n399), .dout(n401));
  jand g0338(.dina(G375gat), .dinb(G69gat), .dout(n402));
  jnot g0339(.din(n402), .dout(n403));
  jand g0340(.dina(n368), .dinb(n343), .dout(n404));
  jand g0341(.dina(n369), .dinb(n340), .dout(n405));
  jcb  g0342(.dina(n405), .dinb(n404), .dout(n406));
  jand g0343(.dina(G358gat), .dinb(G86gat), .dout(n407));
  jnot g0344(.din(n407), .dout(n408));
  jand g0345(.dina(n366), .dinb(n348), .dout(n409));
  jand g0346(.dina(n367), .dinb(n345), .dout(n410));
  jcb  g0347(.dina(n410), .dinb(n409), .dout(n411));
  jand g0348(.dina(G341gat), .dinb(G103gat), .dout(n412));
  jnot g0349(.din(n412), .dout(n413));
  jand g0350(.dina(n364), .dinb(n354), .dout(n414));
  jand g0351(.dina(n365), .dinb(n350), .dout(n415));
  jcb  g0352(.dina(n415), .dinb(n414), .dout(n416));
  jand g0353(.dina(G324gat), .dinb(G120gat), .dout(n417));
  jnot g0354(.din(n417), .dout(n418));
  jcb  g0355(.dina(n362), .dinb(n297), .dout(n419));
  jand g0356(.dina(n363), .dinb(n356), .dout(n420));
  jnot g0357(.din(n420), .dout(n421));
  jand g0358(.dina(n421), .dinb(n419), .dout(n422));
  jnot g0359(.din(n422), .dout(n423));
  jand g0360(.dina(G307gat), .dinb(G137gat), .dout(n424));
  jnot g0361(.din(n424), .dout(n425));
  jand g0362(.dina(G290gat), .dinb(G171gat), .dout(n426));
  jand g0363(.dina(n426), .dinb(n360), .dout(n427));
  jnot g0364(.din(n427), .dout(n428));
  jand g0365(.dina(G273gat), .dinb(G171gat), .dout(n429));
  jcb  g0366(.dina(n429), .dinb(n357), .dout(n430));
  jand g0367(.dina(n430), .dinb(n428), .dout(n431));
  jxor g0368(.dina(n431), .dinb(n358), .dout(n432));
  jxor g0369(.dina(n432), .dinb(n425), .dout(n433));
  jxor g0370(.dina(n433), .dinb(n423), .dout(n434));
  jxor g0371(.dina(n434), .dinb(n418), .dout(n435));
  jxor g0372(.dina(n435), .dinb(n416), .dout(n436));
  jxor g0373(.dina(n436), .dinb(n413), .dout(n437));
  jxor g0374(.dina(n437), .dinb(n411), .dout(n438));
  jxor g0375(.dina(n438), .dinb(n408), .dout(n439));
  jxor g0376(.dina(n439), .dinb(n406), .dout(n440));
  jxor g0377(.dina(n440), .dinb(n403), .dout(n441));
  jxor g0378(.dina(n441), .dinb(n401), .dout(n442));
  jxor g0379(.dina(n442), .dinb(n398), .dout(n443));
  jxor g0380(.dina(n443), .dinb(n396), .dout(n444));
  jxor g0381(.dina(n444), .dinb(n393), .dout(n445));
  jnot g0382(.din(n445), .dout(n446));
  jxor g0383(.dina(n446), .dinb(n391), .dout(n447));
  jxor g0384(.dina(n447), .dinb(n387), .dout(n448));
  jxor g0385(.dina(n448), .dinb(n385), .dout(n449));
  jxor g0386(.dina(n449), .dinb(n381), .dout(G4591gat));
  jand g0387(.dina(G460gat), .dinb(G1gat), .dout(n451));
  jnot g0388(.din(n451), .dout(n452));
  jnot g0389(.din(n448), .dout(n453));
  jcb  g0390(.dina(n453), .dinb(n385), .dout(n454));
  jcb  g0391(.dina(n449), .dinb(n380), .dout(n455));
  jand g0392(.dina(n455), .dinb(n454), .dout(n456));
  jand g0393(.dina(G443gat), .dinb(G18gat), .dout(n457));
  jnot g0394(.din(n457), .dout(n458));
  jcb  g0395(.dina(n446), .dinb(n391), .dout(n459));
  jxor g0396(.dina(n445), .dinb(n391), .dout(n460));
  jcb  g0397(.dina(n460), .dinb(n386), .dout(n461));
  jand g0398(.dina(n461), .dinb(n459), .dout(n462));
  jand g0399(.dina(G426gat), .dinb(G35gat), .dout(n463));
  jnot g0400(.din(n463), .dout(n464));
  jand g0401(.dina(n443), .dinb(n396), .dout(n465));
  jand g0402(.dina(n444), .dinb(n393), .dout(n466));
  jcb  g0403(.dina(n466), .dinb(n465), .dout(n467));
  jand g0404(.dina(G409gat), .dinb(G52gat), .dout(n468));
  jnot g0405(.din(n468), .dout(n469));
  jand g0406(.dina(n441), .dinb(n401), .dout(n470));
  jand g0407(.dina(n442), .dinb(n398), .dout(n471));
  jcb  g0408(.dina(n471), .dinb(n470), .dout(n472));
  jand g0409(.dina(G392gat), .dinb(G69gat), .dout(n473));
  jnot g0410(.din(n473), .dout(n474));
  jand g0411(.dina(n439), .dinb(n406), .dout(n475));
  jand g0412(.dina(n440), .dinb(n403), .dout(n476));
  jcb  g0413(.dina(n476), .dinb(n475), .dout(n477));
  jand g0414(.dina(G375gat), .dinb(G86gat), .dout(n478));
  jnot g0415(.din(n478), .dout(n479));
  jand g0416(.dina(n437), .dinb(n411), .dout(n480));
  jand g0417(.dina(n438), .dinb(n408), .dout(n481));
  jcb  g0418(.dina(n481), .dinb(n480), .dout(n482));
  jand g0419(.dina(G358gat), .dinb(G103gat), .dout(n483));
  jnot g0420(.din(n483), .dout(n484));
  jand g0421(.dina(n435), .dinb(n416), .dout(n485));
  jand g0422(.dina(n436), .dinb(n413), .dout(n486));
  jcb  g0423(.dina(n486), .dinb(n485), .dout(n487));
  jand g0424(.dina(G341gat), .dinb(G120gat), .dout(n488));
  jnot g0425(.din(n488), .dout(n489));
  jand g0426(.dina(n433), .dinb(n423), .dout(n490));
  jand g0427(.dina(n434), .dinb(n418), .dout(n491));
  jcb  g0428(.dina(n491), .dinb(n490), .dout(n492));
  jand g0429(.dina(G324gat), .dinb(G137gat), .dout(n493));
  jnot g0430(.din(n493), .dout(n494));
  jcb  g0431(.dina(n431), .dinb(n358), .dout(n495));
  jand g0432(.dina(n432), .dinb(n425), .dout(n496));
  jnot g0433(.din(n496), .dout(n497));
  jand g0434(.dina(n497), .dinb(n495), .dout(n498));
  jnot g0435(.din(n498), .dout(n499));
  jand g0436(.dina(G307gat), .dinb(G154gat), .dout(n500));
  jnot g0437(.din(n500), .dout(n501));
  jand g0438(.dina(G290gat), .dinb(G188gat), .dout(n502));
  jand g0439(.dina(n502), .dinb(n429), .dout(n503));
  jnot g0440(.din(n503), .dout(n504));
  jand g0441(.dina(G273gat), .dinb(G188gat), .dout(n505));
  jcb  g0442(.dina(n505), .dinb(n426), .dout(n506));
  jand g0443(.dina(n506), .dinb(n504), .dout(n507));
  jxor g0444(.dina(n507), .dinb(n427), .dout(n508));
  jxor g0445(.dina(n508), .dinb(n501), .dout(n509));
  jxor g0446(.dina(n509), .dinb(n499), .dout(n510));
  jxor g0447(.dina(n510), .dinb(n494), .dout(n511));
  jxor g0448(.dina(n511), .dinb(n492), .dout(n512));
  jxor g0449(.dina(n512), .dinb(n489), .dout(n513));
  jxor g0450(.dina(n513), .dinb(n487), .dout(n514));
  jxor g0451(.dina(n514), .dinb(n484), .dout(n515));
  jxor g0452(.dina(n515), .dinb(n482), .dout(n516));
  jxor g0453(.dina(n516), .dinb(n479), .dout(n517));
  jxor g0454(.dina(n517), .dinb(n477), .dout(n518));
  jxor g0455(.dina(n518), .dinb(n474), .dout(n519));
  jxor g0456(.dina(n519), .dinb(n472), .dout(n520));
  jxor g0457(.dina(n520), .dinb(n469), .dout(n521));
  jxor g0458(.dina(n521), .dinb(n467), .dout(n522));
  jxor g0459(.dina(n522), .dinb(n464), .dout(n523));
  jnot g0460(.din(n523), .dout(n524));
  jxor g0461(.dina(n524), .dinb(n462), .dout(n525));
  jxor g0462(.dina(n525), .dinb(n458), .dout(n526));
  jxor g0463(.dina(n526), .dinb(n456), .dout(n527));
  jxor g0464(.dina(n527), .dinb(n452), .dout(G4946gat));
  jand g0465(.dina(G477gat), .dinb(G1gat), .dout(n529));
  jnot g0466(.din(n529), .dout(n530));
  jnot g0467(.din(n526), .dout(n531));
  jcb  g0468(.dina(n531), .dinb(n456), .dout(n532));
  jcb  g0469(.dina(n527), .dinb(n451), .dout(n533));
  jand g0470(.dina(n533), .dinb(n532), .dout(n534));
  jand g0471(.dina(G460gat), .dinb(G18gat), .dout(n535));
  jnot g0472(.din(n535), .dout(n536));
  jcb  g0473(.dina(n524), .dinb(n462), .dout(n537));
  jxor g0474(.dina(n523), .dinb(n462), .dout(n538));
  jcb  g0475(.dina(n538), .dinb(n457), .dout(n539));
  jand g0476(.dina(n539), .dinb(n537), .dout(n540));
  jand g0477(.dina(G443gat), .dinb(G35gat), .dout(n541));
  jnot g0478(.din(n541), .dout(n542));
  jand g0479(.dina(n521), .dinb(n467), .dout(n543));
  jand g0480(.dina(n522), .dinb(n464), .dout(n544));
  jcb  g0481(.dina(n544), .dinb(n543), .dout(n545));
  jand g0482(.dina(G426gat), .dinb(G52gat), .dout(n546));
  jnot g0483(.din(n546), .dout(n547));
  jand g0484(.dina(n519), .dinb(n472), .dout(n548));
  jand g0485(.dina(n520), .dinb(n469), .dout(n549));
  jcb  g0486(.dina(n549), .dinb(n548), .dout(n550));
  jand g0487(.dina(G409gat), .dinb(G69gat), .dout(n551));
  jnot g0488(.din(n551), .dout(n552));
  jand g0489(.dina(n517), .dinb(n477), .dout(n553));
  jand g0490(.dina(n518), .dinb(n474), .dout(n554));
  jcb  g0491(.dina(n554), .dinb(n553), .dout(n555));
  jand g0492(.dina(G392gat), .dinb(G86gat), .dout(n556));
  jnot g0493(.din(n556), .dout(n557));
  jand g0494(.dina(n515), .dinb(n482), .dout(n558));
  jand g0495(.dina(n516), .dinb(n479), .dout(n559));
  jcb  g0496(.dina(n559), .dinb(n558), .dout(n560));
  jand g0497(.dina(G375gat), .dinb(G103gat), .dout(n561));
  jnot g0498(.din(n561), .dout(n562));
  jand g0499(.dina(n513), .dinb(n487), .dout(n563));
  jand g0500(.dina(n514), .dinb(n484), .dout(n564));
  jcb  g0501(.dina(n564), .dinb(n563), .dout(n565));
  jand g0502(.dina(G358gat), .dinb(G120gat), .dout(n566));
  jnot g0503(.din(n566), .dout(n567));
  jand g0504(.dina(n511), .dinb(n492), .dout(n568));
  jand g0505(.dina(n512), .dinb(n489), .dout(n569));
  jcb  g0506(.dina(n569), .dinb(n568), .dout(n570));
  jand g0507(.dina(G341gat), .dinb(G137gat), .dout(n571));
  jnot g0508(.din(n571), .dout(n572));
  jand g0509(.dina(n509), .dinb(n499), .dout(n573));
  jand g0510(.dina(n510), .dinb(n494), .dout(n574));
  jcb  g0511(.dina(n574), .dinb(n573), .dout(n575));
  jand g0512(.dina(G324gat), .dinb(G154gat), .dout(n576));
  jnot g0513(.din(n576), .dout(n577));
  jcb  g0514(.dina(n507), .dinb(n427), .dout(n578));
  jand g0515(.dina(n508), .dinb(n501), .dout(n579));
  jnot g0516(.din(n579), .dout(n580));
  jand g0517(.dina(n580), .dinb(n578), .dout(n581));
  jnot g0518(.din(n581), .dout(n582));
  jand g0519(.dina(G307gat), .dinb(G171gat), .dout(n583));
  jnot g0520(.din(n583), .dout(n584));
  jand g0521(.dina(G290gat), .dinb(G205gat), .dout(n585));
  jand g0522(.dina(n585), .dinb(n505), .dout(n586));
  jnot g0523(.din(n586), .dout(n587));
  jand g0524(.dina(G273gat), .dinb(G205gat), .dout(n588));
  jcb  g0525(.dina(n588), .dinb(n502), .dout(n589));
  jand g0526(.dina(n589), .dinb(n587), .dout(n590));
  jxor g0527(.dina(n590), .dinb(n503), .dout(n591));
  jxor g0528(.dina(n591), .dinb(n584), .dout(n592));
  jxor g0529(.dina(n592), .dinb(n582), .dout(n593));
  jxor g0530(.dina(n593), .dinb(n577), .dout(n594));
  jxor g0531(.dina(n594), .dinb(n575), .dout(n595));
  jxor g0532(.dina(n595), .dinb(n572), .dout(n596));
  jxor g0533(.dina(n596), .dinb(n570), .dout(n597));
  jxor g0534(.dina(n597), .dinb(n567), .dout(n598));
  jxor g0535(.dina(n598), .dinb(n565), .dout(n599));
  jxor g0536(.dina(n599), .dinb(n562), .dout(n600));
  jxor g0537(.dina(n600), .dinb(n560), .dout(n601));
  jxor g0538(.dina(n601), .dinb(n557), .dout(n602));
  jxor g0539(.dina(n602), .dinb(n555), .dout(n603));
  jxor g0540(.dina(n603), .dinb(n552), .dout(n604));
  jxor g0541(.dina(n604), .dinb(n550), .dout(n605));
  jxor g0542(.dina(n605), .dinb(n547), .dout(n606));
  jxor g0543(.dina(n606), .dinb(n545), .dout(n607));
  jxor g0544(.dina(n607), .dinb(n542), .dout(n608));
  jnot g0545(.din(n608), .dout(n609));
  jxor g0546(.dina(n609), .dinb(n540), .dout(n610));
  jxor g0547(.dina(n610), .dinb(n536), .dout(n611));
  jxor g0548(.dina(n611), .dinb(n534), .dout(n612));
  jxor g0549(.dina(n612), .dinb(n530), .dout(G5308gat));
  jand g0550(.dina(G494gat), .dinb(G1gat), .dout(n614));
  jnot g0551(.din(n614), .dout(n615));
  jnot g0552(.din(n611), .dout(n616));
  jcb  g0553(.dina(n616), .dinb(n534), .dout(n617));
  jcb  g0554(.dina(n612), .dinb(n529), .dout(n618));
  jand g0555(.dina(n618), .dinb(n617), .dout(n619));
  jand g0556(.dina(G477gat), .dinb(G18gat), .dout(n620));
  jnot g0557(.din(n620), .dout(n621));
  jcb  g0558(.dina(n609), .dinb(n540), .dout(n622));
  jxor g0559(.dina(n608), .dinb(n540), .dout(n623));
  jcb  g0560(.dina(n623), .dinb(n535), .dout(n624));
  jand g0561(.dina(n624), .dinb(n622), .dout(n625));
  jand g0562(.dina(G460gat), .dinb(G35gat), .dout(n626));
  jnot g0563(.din(n626), .dout(n627));
  jand g0564(.dina(n606), .dinb(n545), .dout(n628));
  jand g0565(.dina(n607), .dinb(n542), .dout(n629));
  jcb  g0566(.dina(n629), .dinb(n628), .dout(n630));
  jand g0567(.dina(G443gat), .dinb(G52gat), .dout(n631));
  jnot g0568(.din(n631), .dout(n632));
  jand g0569(.dina(n604), .dinb(n550), .dout(n633));
  jand g0570(.dina(n605), .dinb(n547), .dout(n634));
  jcb  g0571(.dina(n634), .dinb(n633), .dout(n635));
  jand g0572(.dina(G426gat), .dinb(G69gat), .dout(n636));
  jnot g0573(.din(n636), .dout(n637));
  jand g0574(.dina(n602), .dinb(n555), .dout(n638));
  jand g0575(.dina(n603), .dinb(n552), .dout(n639));
  jcb  g0576(.dina(n639), .dinb(n638), .dout(n640));
  jand g0577(.dina(G409gat), .dinb(G86gat), .dout(n641));
  jnot g0578(.din(n641), .dout(n642));
  jand g0579(.dina(n600), .dinb(n560), .dout(n643));
  jand g0580(.dina(n601), .dinb(n557), .dout(n644));
  jcb  g0581(.dina(n644), .dinb(n643), .dout(n645));
  jand g0582(.dina(G392gat), .dinb(G103gat), .dout(n646));
  jnot g0583(.din(n646), .dout(n647));
  jand g0584(.dina(n598), .dinb(n565), .dout(n648));
  jand g0585(.dina(n599), .dinb(n562), .dout(n649));
  jcb  g0586(.dina(n649), .dinb(n648), .dout(n650));
  jand g0587(.dina(G375gat), .dinb(G120gat), .dout(n651));
  jnot g0588(.din(n651), .dout(n652));
  jand g0589(.dina(n596), .dinb(n570), .dout(n653));
  jand g0590(.dina(n597), .dinb(n567), .dout(n654));
  jcb  g0591(.dina(n654), .dinb(n653), .dout(n655));
  jand g0592(.dina(G358gat), .dinb(G137gat), .dout(n656));
  jnot g0593(.din(n656), .dout(n657));
  jand g0594(.dina(n594), .dinb(n575), .dout(n658));
  jand g0595(.dina(n595), .dinb(n572), .dout(n659));
  jcb  g0596(.dina(n659), .dinb(n658), .dout(n660));
  jand g0597(.dina(G341gat), .dinb(G154gat), .dout(n661));
  jnot g0598(.din(n661), .dout(n662));
  jand g0599(.dina(n592), .dinb(n582), .dout(n663));
  jand g0600(.dina(n593), .dinb(n577), .dout(n664));
  jcb  g0601(.dina(n664), .dinb(n663), .dout(n665));
  jand g0602(.dina(G324gat), .dinb(G171gat), .dout(n666));
  jnot g0603(.din(n666), .dout(n667));
  jcb  g0604(.dina(n590), .dinb(n503), .dout(n668));
  jand g0605(.dina(n591), .dinb(n584), .dout(n669));
  jnot g0606(.din(n669), .dout(n670));
  jand g0607(.dina(n670), .dinb(n668), .dout(n671));
  jnot g0608(.din(n671), .dout(n672));
  jand g0609(.dina(G307gat), .dinb(G188gat), .dout(n673));
  jnot g0610(.din(n673), .dout(n674));
  jand g0611(.dina(G290gat), .dinb(G222gat), .dout(n675));
  jand g0612(.dina(n675), .dinb(n588), .dout(n676));
  jnot g0613(.din(n676), .dout(n677));
  jand g0614(.dina(G273gat), .dinb(G222gat), .dout(n678));
  jcb  g0615(.dina(n678), .dinb(n585), .dout(n679));
  jand g0616(.dina(n679), .dinb(n677), .dout(n680));
  jxor g0617(.dina(n680), .dinb(n586), .dout(n681));
  jxor g0618(.dina(n681), .dinb(n674), .dout(n682));
  jxor g0619(.dina(n682), .dinb(n672), .dout(n683));
  jxor g0620(.dina(n683), .dinb(n667), .dout(n684));
  jxor g0621(.dina(n684), .dinb(n665), .dout(n685));
  jxor g0622(.dina(n685), .dinb(n662), .dout(n686));
  jxor g0623(.dina(n686), .dinb(n660), .dout(n687));
  jxor g0624(.dina(n687), .dinb(n657), .dout(n688));
  jxor g0625(.dina(n688), .dinb(n655), .dout(n689));
  jxor g0626(.dina(n689), .dinb(n652), .dout(n690));
  jxor g0627(.dina(n690), .dinb(n650), .dout(n691));
  jxor g0628(.dina(n691), .dinb(n647), .dout(n692));
  jxor g0629(.dina(n692), .dinb(n645), .dout(n693));
  jxor g0630(.dina(n693), .dinb(n642), .dout(n694));
  jxor g0631(.dina(n694), .dinb(n640), .dout(n695));
  jxor g0632(.dina(n695), .dinb(n637), .dout(n696));
  jxor g0633(.dina(n696), .dinb(n635), .dout(n697));
  jxor g0634(.dina(n697), .dinb(n632), .dout(n698));
  jxor g0635(.dina(n698), .dinb(n630), .dout(n699));
  jxor g0636(.dina(n699), .dinb(n627), .dout(n700));
  jnot g0637(.din(n700), .dout(n701));
  jxor g0638(.dina(n701), .dinb(n625), .dout(n702));
  jxor g0639(.dina(n702), .dinb(n621), .dout(n703));
  jxor g0640(.dina(n703), .dinb(n619), .dout(n704));
  jxor g0641(.dina(n704), .dinb(n615), .dout(G5672gat));
  jand g0642(.dina(G511gat), .dinb(G1gat), .dout(n706));
  jnot g0643(.din(n706), .dout(n707));
  jnot g0644(.din(n703), .dout(n708));
  jcb  g0645(.dina(n708), .dinb(n619), .dout(n709));
  jcb  g0646(.dina(n704), .dinb(n614), .dout(n710));
  jand g0647(.dina(n710), .dinb(n709), .dout(n711));
  jand g0648(.dina(G494gat), .dinb(G18gat), .dout(n712));
  jnot g0649(.din(n712), .dout(n713));
  jcb  g0650(.dina(n701), .dinb(n625), .dout(n714));
  jxor g0651(.dina(n700), .dinb(n625), .dout(n715));
  jcb  g0652(.dina(n715), .dinb(n620), .dout(n716));
  jand g0653(.dina(n716), .dinb(n714), .dout(n717));
  jand g0654(.dina(G477gat), .dinb(G35gat), .dout(n718));
  jnot g0655(.din(n718), .dout(n719));
  jand g0656(.dina(n698), .dinb(n630), .dout(n720));
  jand g0657(.dina(n699), .dinb(n627), .dout(n721));
  jcb  g0658(.dina(n721), .dinb(n720), .dout(n722));
  jand g0659(.dina(G460gat), .dinb(G52gat), .dout(n723));
  jnot g0660(.din(n723), .dout(n724));
  jand g0661(.dina(n696), .dinb(n635), .dout(n725));
  jand g0662(.dina(n697), .dinb(n632), .dout(n726));
  jcb  g0663(.dina(n726), .dinb(n725), .dout(n727));
  jand g0664(.dina(G443gat), .dinb(G69gat), .dout(n728));
  jnot g0665(.din(n728), .dout(n729));
  jand g0666(.dina(n694), .dinb(n640), .dout(n730));
  jand g0667(.dina(n695), .dinb(n637), .dout(n731));
  jcb  g0668(.dina(n731), .dinb(n730), .dout(n732));
  jand g0669(.dina(G426gat), .dinb(G86gat), .dout(n733));
  jnot g0670(.din(n733), .dout(n734));
  jand g0671(.dina(n692), .dinb(n645), .dout(n735));
  jand g0672(.dina(n693), .dinb(n642), .dout(n736));
  jcb  g0673(.dina(n736), .dinb(n735), .dout(n737));
  jand g0674(.dina(G409gat), .dinb(G103gat), .dout(n738));
  jnot g0675(.din(n738), .dout(n739));
  jand g0676(.dina(n690), .dinb(n650), .dout(n740));
  jand g0677(.dina(n691), .dinb(n647), .dout(n741));
  jcb  g0678(.dina(n741), .dinb(n740), .dout(n742));
  jand g0679(.dina(G392gat), .dinb(G120gat), .dout(n743));
  jnot g0680(.din(n743), .dout(n744));
  jand g0681(.dina(n688), .dinb(n655), .dout(n745));
  jand g0682(.dina(n689), .dinb(n652), .dout(n746));
  jcb  g0683(.dina(n746), .dinb(n745), .dout(n747));
  jand g0684(.dina(G375gat), .dinb(G137gat), .dout(n748));
  jnot g0685(.din(n748), .dout(n749));
  jand g0686(.dina(n686), .dinb(n660), .dout(n750));
  jand g0687(.dina(n687), .dinb(n657), .dout(n751));
  jcb  g0688(.dina(n751), .dinb(n750), .dout(n752));
  jand g0689(.dina(G358gat), .dinb(G154gat), .dout(n753));
  jnot g0690(.din(n753), .dout(n754));
  jand g0691(.dina(n684), .dinb(n665), .dout(n755));
  jand g0692(.dina(n685), .dinb(n662), .dout(n756));
  jcb  g0693(.dina(n756), .dinb(n755), .dout(n757));
  jand g0694(.dina(G341gat), .dinb(G171gat), .dout(n758));
  jnot g0695(.din(n758), .dout(n759));
  jand g0696(.dina(n682), .dinb(n672), .dout(n760));
  jand g0697(.dina(n683), .dinb(n667), .dout(n761));
  jcb  g0698(.dina(n761), .dinb(n760), .dout(n762));
  jand g0699(.dina(G324gat), .dinb(G188gat), .dout(n763));
  jnot g0700(.din(n763), .dout(n764));
  jcb  g0701(.dina(n680), .dinb(n586), .dout(n765));
  jand g0702(.dina(n681), .dinb(n674), .dout(n766));
  jnot g0703(.din(n766), .dout(n767));
  jand g0704(.dina(n767), .dinb(n765), .dout(n768));
  jnot g0705(.din(n768), .dout(n769));
  jand g0706(.dina(G307gat), .dinb(G205gat), .dout(n770));
  jnot g0707(.din(n770), .dout(n771));
  jand g0708(.dina(G290gat), .dinb(G239gat), .dout(n772));
  jand g0709(.dina(n772), .dinb(n678), .dout(n773));
  jnot g0710(.din(n773), .dout(n774));
  jand g0711(.dina(G273gat), .dinb(G239gat), .dout(n775));
  jcb  g0712(.dina(n775), .dinb(n675), .dout(n776));
  jand g0713(.dina(n776), .dinb(n774), .dout(n777));
  jxor g0714(.dina(n777), .dinb(n676), .dout(n778));
  jxor g0715(.dina(n778), .dinb(n771), .dout(n779));
  jxor g0716(.dina(n779), .dinb(n769), .dout(n780));
  jxor g0717(.dina(n780), .dinb(n764), .dout(n781));
  jxor g0718(.dina(n781), .dinb(n762), .dout(n782));
  jxor g0719(.dina(n782), .dinb(n759), .dout(n783));
  jxor g0720(.dina(n783), .dinb(n757), .dout(n784));
  jxor g0721(.dina(n784), .dinb(n754), .dout(n785));
  jxor g0722(.dina(n785), .dinb(n752), .dout(n786));
  jxor g0723(.dina(n786), .dinb(n749), .dout(n787));
  jxor g0724(.dina(n787), .dinb(n747), .dout(n788));
  jxor g0725(.dina(n788), .dinb(n744), .dout(n789));
  jxor g0726(.dina(n789), .dinb(n742), .dout(n790));
  jxor g0727(.dina(n790), .dinb(n739), .dout(n791));
  jxor g0728(.dina(n791), .dinb(n737), .dout(n792));
  jxor g0729(.dina(n792), .dinb(n734), .dout(n793));
  jxor g0730(.dina(n793), .dinb(n732), .dout(n794));
  jxor g0731(.dina(n794), .dinb(n729), .dout(n795));
  jxor g0732(.dina(n795), .dinb(n727), .dout(n796));
  jxor g0733(.dina(n796), .dinb(n724), .dout(n797));
  jxor g0734(.dina(n797), .dinb(n722), .dout(n798));
  jxor g0735(.dina(n798), .dinb(n719), .dout(n799));
  jnot g0736(.din(n799), .dout(n800));
  jxor g0737(.dina(n800), .dinb(n717), .dout(n801));
  jxor g0738(.dina(n801), .dinb(n713), .dout(n802));
  jxor g0739(.dina(n802), .dinb(n711), .dout(n803));
  jxor g0740(.dina(n803), .dinb(n707), .dout(G5971gat));
  jand g0741(.dina(G528gat), .dinb(G1gat), .dout(n805));
  jnot g0742(.din(n805), .dout(n806));
  jnot g0743(.din(n802), .dout(n807));
  jcb  g0744(.dina(n807), .dinb(n711), .dout(n808));
  jcb  g0745(.dina(n803), .dinb(n706), .dout(n809));
  jand g0746(.dina(n809), .dinb(n808), .dout(n810));
  jand g0747(.dina(G511gat), .dinb(G18gat), .dout(n811));
  jcb  g0748(.dina(n800), .dinb(n717), .dout(n812));
  jxor g0749(.dina(n799), .dinb(n717), .dout(n813));
  jcb  g0750(.dina(n813), .dinb(n712), .dout(n814));
  jand g0751(.dina(n814), .dinb(n812), .dout(n815));
  jand g0752(.dina(G494gat), .dinb(G35gat), .dout(n816));
  jnot g0753(.din(n816), .dout(n817));
  jand g0754(.dina(n797), .dinb(n722), .dout(n818));
  jand g0755(.dina(n798), .dinb(n719), .dout(n819));
  jcb  g0756(.dina(n819), .dinb(n818), .dout(n820));
  jand g0757(.dina(G477gat), .dinb(G52gat), .dout(n821));
  jnot g0758(.din(n821), .dout(n822));
  jand g0759(.dina(n795), .dinb(n727), .dout(n823));
  jand g0760(.dina(n796), .dinb(n724), .dout(n824));
  jcb  g0761(.dina(n824), .dinb(n823), .dout(n825));
  jand g0762(.dina(G460gat), .dinb(G69gat), .dout(n826));
  jnot g0763(.din(n826), .dout(n827));
  jand g0764(.dina(n793), .dinb(n732), .dout(n828));
  jand g0765(.dina(n794), .dinb(n729), .dout(n829));
  jcb  g0766(.dina(n829), .dinb(n828), .dout(n830));
  jand g0767(.dina(G443gat), .dinb(G86gat), .dout(n831));
  jnot g0768(.din(n831), .dout(n832));
  jand g0769(.dina(n791), .dinb(n737), .dout(n833));
  jand g0770(.dina(n792), .dinb(n734), .dout(n834));
  jcb  g0771(.dina(n834), .dinb(n833), .dout(n835));
  jand g0772(.dina(G426gat), .dinb(G103gat), .dout(n836));
  jnot g0773(.din(n836), .dout(n837));
  jand g0774(.dina(n789), .dinb(n742), .dout(n838));
  jand g0775(.dina(n790), .dinb(n739), .dout(n839));
  jcb  g0776(.dina(n839), .dinb(n838), .dout(n840));
  jand g0777(.dina(G409gat), .dinb(G120gat), .dout(n841));
  jnot g0778(.din(n841), .dout(n842));
  jand g0779(.dina(n787), .dinb(n747), .dout(n843));
  jand g0780(.dina(n788), .dinb(n744), .dout(n844));
  jcb  g0781(.dina(n844), .dinb(n843), .dout(n845));
  jand g0782(.dina(G392gat), .dinb(G137gat), .dout(n846));
  jnot g0783(.din(n846), .dout(n847));
  jand g0784(.dina(n785), .dinb(n752), .dout(n848));
  jand g0785(.dina(n786), .dinb(n749), .dout(n849));
  jcb  g0786(.dina(n849), .dinb(n848), .dout(n850));
  jand g0787(.dina(G375gat), .dinb(G154gat), .dout(n851));
  jnot g0788(.din(n851), .dout(n852));
  jand g0789(.dina(n783), .dinb(n757), .dout(n853));
  jand g0790(.dina(n784), .dinb(n754), .dout(n854));
  jcb  g0791(.dina(n854), .dinb(n853), .dout(n855));
  jand g0792(.dina(G358gat), .dinb(G171gat), .dout(n856));
  jnot g0793(.din(n856), .dout(n857));
  jand g0794(.dina(n781), .dinb(n762), .dout(n858));
  jand g0795(.dina(n782), .dinb(n759), .dout(n859));
  jcb  g0796(.dina(n859), .dinb(n858), .dout(n860));
  jand g0797(.dina(G341gat), .dinb(G188gat), .dout(n861));
  jnot g0798(.din(n861), .dout(n862));
  jand g0799(.dina(n779), .dinb(n769), .dout(n863));
  jand g0800(.dina(n780), .dinb(n764), .dout(n864));
  jcb  g0801(.dina(n864), .dinb(n863), .dout(n865));
  jand g0802(.dina(G324gat), .dinb(G205gat), .dout(n866));
  jnot g0803(.din(n866), .dout(n867));
  jcb  g0804(.dina(n777), .dinb(n676), .dout(n868));
  jand g0805(.dina(n778), .dinb(n771), .dout(n869));
  jnot g0806(.din(n869), .dout(n870));
  jand g0807(.dina(n870), .dinb(n868), .dout(n871));
  jnot g0808(.din(n871), .dout(n872));
  jand g0809(.dina(G307gat), .dinb(G222gat), .dout(n873));
  jnot g0810(.din(n873), .dout(n874));
  jand g0811(.dina(G273gat), .dinb(G256gat), .dout(n875));
  jxor g0812(.dina(n875), .dinb(n772), .dout(n876));
  jcb  g0813(.dina(n876), .dinb(n773), .dout(n877));
  jcb  g0814(.dina(n875), .dinb(n774), .dout(n878));
  jand g0815(.dina(n878), .dinb(n877), .dout(n879));
  jxor g0816(.dina(n879), .dinb(n874), .dout(n880));
  jxor g0817(.dina(n880), .dinb(n872), .dout(n881));
  jxor g0818(.dina(n881), .dinb(n867), .dout(n882));
  jxor g0819(.dina(n882), .dinb(n865), .dout(n883));
  jxor g0820(.dina(n883), .dinb(n862), .dout(n884));
  jxor g0821(.dina(n884), .dinb(n860), .dout(n885));
  jxor g0822(.dina(n885), .dinb(n857), .dout(n886));
  jxor g0823(.dina(n886), .dinb(n855), .dout(n887));
  jxor g0824(.dina(n887), .dinb(n852), .dout(n888));
  jxor g0825(.dina(n888), .dinb(n850), .dout(n889));
  jxor g0826(.dina(n889), .dinb(n847), .dout(n890));
  jxor g0827(.dina(n890), .dinb(n845), .dout(n891));
  jxor g0828(.dina(n891), .dinb(n842), .dout(n892));
  jxor g0829(.dina(n892), .dinb(n840), .dout(n893));
  jxor g0830(.dina(n893), .dinb(n837), .dout(n894));
  jxor g0831(.dina(n894), .dinb(n835), .dout(n895));
  jxor g0832(.dina(n895), .dinb(n832), .dout(n896));
  jxor g0833(.dina(n896), .dinb(n830), .dout(n897));
  jxor g0834(.dina(n897), .dinb(n827), .dout(n898));
  jxor g0835(.dina(n898), .dinb(n825), .dout(n899));
  jxor g0836(.dina(n899), .dinb(n822), .dout(n900));
  jxor g0837(.dina(n900), .dinb(n820), .dout(n901));
  jxor g0838(.dina(n901), .dinb(n817), .dout(n902));
  jxor g0839(.dina(n902), .dinb(n815), .dout(n903));
  jxor g0840(.dina(n903), .dinb(n811), .dout(n904));
  jxor g0841(.dina(n904), .dinb(n810), .dout(n905));
  jxor g0842(.dina(n905), .dinb(n806), .dout(G6123gat));
  jnot g0843(.din(n904), .dout(n907));
  jcb  g0844(.dina(n907), .dinb(n810), .dout(n908));
  jcb  g0845(.dina(n905), .dinb(n805), .dout(n909));
  jand g0846(.dina(n909), .dinb(n908), .dout(n910));
  jand g0847(.dina(G528gat), .dinb(G18gat), .dout(n911));
  jnot g0848(.din(n902), .dout(n912));
  jcb  g0849(.dina(n912), .dinb(n815), .dout(n913));
  jcb  g0850(.dina(n903), .dinb(n811), .dout(n914));
  jand g0851(.dina(n914), .dinb(n913), .dout(n915));
  jand g0852(.dina(G511gat), .dinb(G35gat), .dout(n916));
  jand g0853(.dina(n900), .dinb(n820), .dout(n917));
  jnot g0854(.din(n917), .dout(n918));
  jnot g0855(.din(n900), .dout(n919));
  jxor g0856(.dina(n919), .dinb(n820), .dout(n920));
  jcb  g0857(.dina(n920), .dinb(n816), .dout(n921));
  jand g0858(.dina(n921), .dinb(n918), .dout(n922));
  jand g0859(.dina(G494gat), .dinb(G52gat), .dout(n923));
  jnot g0860(.din(n923), .dout(n924));
  jand g0861(.dina(n898), .dinb(n825), .dout(n925));
  jand g0862(.dina(n899), .dinb(n822), .dout(n926));
  jcb  g0863(.dina(n926), .dinb(n925), .dout(n927));
  jand g0864(.dina(G477gat), .dinb(G69gat), .dout(n928));
  jnot g0865(.din(n928), .dout(n929));
  jand g0866(.dina(n896), .dinb(n830), .dout(n930));
  jand g0867(.dina(n897), .dinb(n827), .dout(n931));
  jcb  g0868(.dina(n931), .dinb(n930), .dout(n932));
  jand g0869(.dina(G460gat), .dinb(G86gat), .dout(n933));
  jnot g0870(.din(n933), .dout(n934));
  jand g0871(.dina(n894), .dinb(n835), .dout(n935));
  jand g0872(.dina(n895), .dinb(n832), .dout(n936));
  jcb  g0873(.dina(n936), .dinb(n935), .dout(n937));
  jand g0874(.dina(G443gat), .dinb(G103gat), .dout(n938));
  jnot g0875(.din(n938), .dout(n939));
  jand g0876(.dina(n892), .dinb(n840), .dout(n940));
  jand g0877(.dina(n893), .dinb(n837), .dout(n941));
  jcb  g0878(.dina(n941), .dinb(n940), .dout(n942));
  jand g0879(.dina(G426gat), .dinb(G120gat), .dout(n943));
  jnot g0880(.din(n943), .dout(n944));
  jand g0881(.dina(n890), .dinb(n845), .dout(n945));
  jand g0882(.dina(n891), .dinb(n842), .dout(n946));
  jcb  g0883(.dina(n946), .dinb(n945), .dout(n947));
  jand g0884(.dina(G409gat), .dinb(G137gat), .dout(n948));
  jnot g0885(.din(n948), .dout(n949));
  jand g0886(.dina(n888), .dinb(n850), .dout(n950));
  jand g0887(.dina(n889), .dinb(n847), .dout(n951));
  jcb  g0888(.dina(n951), .dinb(n950), .dout(n952));
  jand g0889(.dina(G392gat), .dinb(G154gat), .dout(n953));
  jnot g0890(.din(n953), .dout(n954));
  jand g0891(.dina(n886), .dinb(n855), .dout(n955));
  jand g0892(.dina(n887), .dinb(n852), .dout(n956));
  jcb  g0893(.dina(n956), .dinb(n955), .dout(n957));
  jand g0894(.dina(G375gat), .dinb(G171gat), .dout(n958));
  jnot g0895(.din(n958), .dout(n959));
  jand g0896(.dina(n884), .dinb(n860), .dout(n960));
  jand g0897(.dina(n885), .dinb(n857), .dout(n961));
  jcb  g0898(.dina(n961), .dinb(n960), .dout(n962));
  jand g0899(.dina(G358gat), .dinb(G188gat), .dout(n963));
  jnot g0900(.din(n963), .dout(n964));
  jand g0901(.dina(n882), .dinb(n865), .dout(n965));
  jand g0902(.dina(n883), .dinb(n862), .dout(n966));
  jcb  g0903(.dina(n966), .dinb(n965), .dout(n967));
  jand g0904(.dina(G341gat), .dinb(G205gat), .dout(n968));
  jnot g0905(.din(n968), .dout(n969));
  jand g0906(.dina(n880), .dinb(n872), .dout(n970));
  jand g0907(.dina(n881), .dinb(n867), .dout(n971));
  jcb  g0908(.dina(n971), .dinb(n970), .dout(n972));
  jand g0909(.dina(G324gat), .dinb(G222gat), .dout(n973));
  jnot g0910(.din(n973), .dout(n974));
  jand g0911(.dina(n879), .dinb(n874), .dout(n975));
  jnot g0912(.din(n975), .dout(n976));
  jand g0913(.dina(n976), .dinb(n877), .dout(n977));
  jnot g0914(.din(n977), .dout(n978));
  jnot g0915(.din(n775), .dout(n979));
  jand g0916(.dina(G290gat), .dinb(G256gat), .dout(n980));
  jand g0917(.dina(n980), .dinb(n979), .dout(n981));
  jnot g0918(.din(n981), .dout(n982));
  jand g0919(.dina(G307gat), .dinb(G239gat), .dout(n983));
  jxor g0920(.dina(n983), .dinb(n982), .dout(n984));
  jxor g0921(.dina(n984), .dinb(n978), .dout(n985));
  jxor g0922(.dina(n985), .dinb(n974), .dout(n986));
  jxor g0923(.dina(n986), .dinb(n972), .dout(n987));
  jxor g0924(.dina(n987), .dinb(n969), .dout(n988));
  jxor g0925(.dina(n988), .dinb(n967), .dout(n989));
  jxor g0926(.dina(n989), .dinb(n964), .dout(n990));
  jxor g0927(.dina(n990), .dinb(n962), .dout(n991));
  jxor g0928(.dina(n991), .dinb(n959), .dout(n992));
  jxor g0929(.dina(n992), .dinb(n957), .dout(n993));
  jxor g0930(.dina(n993), .dinb(n954), .dout(n994));
  jxor g0931(.dina(n994), .dinb(n952), .dout(n995));
  jxor g0932(.dina(n995), .dinb(n949), .dout(n996));
  jxor g0933(.dina(n996), .dinb(n947), .dout(n997));
  jxor g0934(.dina(n997), .dinb(n944), .dout(n998));
  jxor g0935(.dina(n998), .dinb(n942), .dout(n999));
  jxor g0936(.dina(n999), .dinb(n939), .dout(n1000));
  jxor g0937(.dina(n1000), .dinb(n937), .dout(n1001));
  jxor g0938(.dina(n1001), .dinb(n934), .dout(n1002));
  jxor g0939(.dina(n1002), .dinb(n932), .dout(n1003));
  jxor g0940(.dina(n1003), .dinb(n929), .dout(n1004));
  jxor g0941(.dina(n1004), .dinb(n927), .dout(n1005));
  jxor g0942(.dina(n1005), .dinb(n924), .dout(n1006));
  jxor g0943(.dina(n1006), .dinb(n922), .dout(n1007));
  jxor g0944(.dina(n1007), .dinb(n916), .dout(n1008));
  jnot g0945(.din(n1008), .dout(n1009));
  jxor g0946(.dina(n1009), .dinb(n915), .dout(n1010));
  jxor g0947(.dina(n1010), .dinb(n911), .dout(n1011));
  jxor g0948(.dina(n1011), .dinb(n910), .dout(G6150gat));
  jand g0949(.dina(n1011), .dinb(n910), .dout(n1013));
  jcb  g0950(.dina(n1009), .dinb(n915), .dout(n1014));
  jxor g0951(.dina(n1008), .dinb(n915), .dout(n1015));
  jcb  g0952(.dina(n1015), .dinb(n911), .dout(n1016));
  jand g0953(.dina(n1016), .dinb(n1014), .dout(n1017));
  jand g0954(.dina(G528gat), .dinb(G35gat), .dout(n1018));
  jnot g0955(.din(n1006), .dout(n1019));
  jcb  g0956(.dina(n1019), .dinb(n922), .dout(n1020));
  jcb  g0957(.dina(n1007), .dinb(n916), .dout(n1021));
  jand g0958(.dina(n1021), .dinb(n1020), .dout(n1022));
  jand g0959(.dina(G511gat), .dinb(G52gat), .dout(n1023));
  jand g0960(.dina(n1004), .dinb(n927), .dout(n1024));
  jand g0961(.dina(n1005), .dinb(n924), .dout(n1025));
  jcb  g0962(.dina(n1025), .dinb(n1024), .dout(n1026));
  jand g0963(.dina(G494gat), .dinb(G69gat), .dout(n1027));
  jnot g0964(.din(n1027), .dout(n1028));
  jand g0965(.dina(n1002), .dinb(n932), .dout(n1029));
  jand g0966(.dina(n1003), .dinb(n929), .dout(n1030));
  jcb  g0967(.dina(n1030), .dinb(n1029), .dout(n1031));
  jand g0968(.dina(G477gat), .dinb(G86gat), .dout(n1032));
  jnot g0969(.din(n1032), .dout(n1033));
  jand g0970(.dina(n1000), .dinb(n937), .dout(n1034));
  jand g0971(.dina(n1001), .dinb(n934), .dout(n1035));
  jcb  g0972(.dina(n1035), .dinb(n1034), .dout(n1036));
  jand g0973(.dina(G460gat), .dinb(G103gat), .dout(n1037));
  jnot g0974(.din(n1037), .dout(n1038));
  jand g0975(.dina(n998), .dinb(n942), .dout(n1039));
  jand g0976(.dina(n999), .dinb(n939), .dout(n1040));
  jcb  g0977(.dina(n1040), .dinb(n1039), .dout(n1041));
  jand g0978(.dina(G443gat), .dinb(G120gat), .dout(n1042));
  jnot g0979(.din(n1042), .dout(n1043));
  jand g0980(.dina(n996), .dinb(n947), .dout(n1044));
  jand g0981(.dina(n997), .dinb(n944), .dout(n1045));
  jcb  g0982(.dina(n1045), .dinb(n1044), .dout(n1046));
  jand g0983(.dina(G426gat), .dinb(G137gat), .dout(n1047));
  jnot g0984(.din(n1047), .dout(n1048));
  jand g0985(.dina(n994), .dinb(n952), .dout(n1049));
  jand g0986(.dina(n995), .dinb(n949), .dout(n1050));
  jcb  g0987(.dina(n1050), .dinb(n1049), .dout(n1051));
  jand g0988(.dina(G409gat), .dinb(G154gat), .dout(n1052));
  jnot g0989(.din(n1052), .dout(n1053));
  jand g0990(.dina(n992), .dinb(n957), .dout(n1054));
  jand g0991(.dina(n993), .dinb(n954), .dout(n1055));
  jcb  g0992(.dina(n1055), .dinb(n1054), .dout(n1056));
  jand g0993(.dina(G392gat), .dinb(G171gat), .dout(n1057));
  jnot g0994(.din(n1057), .dout(n1058));
  jand g0995(.dina(n990), .dinb(n962), .dout(n1059));
  jand g0996(.dina(n991), .dinb(n959), .dout(n1060));
  jcb  g0997(.dina(n1060), .dinb(n1059), .dout(n1061));
  jand g0998(.dina(G375gat), .dinb(G188gat), .dout(n1062));
  jnot g0999(.din(n1062), .dout(n1063));
  jand g1000(.dina(n988), .dinb(n967), .dout(n1064));
  jand g1001(.dina(n989), .dinb(n964), .dout(n1065));
  jcb  g1002(.dina(n1065), .dinb(n1064), .dout(n1066));
  jand g1003(.dina(G358gat), .dinb(G205gat), .dout(n1067));
  jnot g1004(.din(n1067), .dout(n1068));
  jand g1005(.dina(n986), .dinb(n972), .dout(n1069));
  jand g1006(.dina(n987), .dinb(n969), .dout(n1070));
  jcb  g1007(.dina(n1070), .dinb(n1069), .dout(n1071));
  jand g1008(.dina(G341gat), .dinb(G222gat), .dout(n1072));
  jnot g1009(.din(n1072), .dout(n1073));
  jand g1010(.dina(n984), .dinb(n978), .dout(n1074));
  jand g1011(.dina(n985), .dinb(n974), .dout(n1075));
  jcb  g1012(.dina(n1075), .dinb(n1074), .dout(n1076));
  jand g1013(.dina(G324gat), .dinb(G239gat), .dout(n1077));
  jand g1014(.dina(G307gat), .dinb(G256gat), .dout(n1078));
  jcb  g1015(.dina(n983), .dinb(n982), .dout(n1079));
  jand g1016(.dina(n1079), .dinb(n980), .dout(n1080));
  jxor g1017(.dina(n1080), .dinb(n1078), .dout(n1081));
  jnot g1018(.din(n1081), .dout(n1082));
  jxor g1019(.dina(n1082), .dinb(n1077), .dout(n1083));
  jxor g1020(.dina(n1083), .dinb(n1076), .dout(n1084));
  jxor g1021(.dina(n1084), .dinb(n1073), .dout(n1085));
  jxor g1022(.dina(n1085), .dinb(n1071), .dout(n1086));
  jxor g1023(.dina(n1086), .dinb(n1068), .dout(n1087));
  jxor g1024(.dina(n1087), .dinb(n1066), .dout(n1088));
  jxor g1025(.dina(n1088), .dinb(n1063), .dout(n1089));
  jxor g1026(.dina(n1089), .dinb(n1061), .dout(n1090));
  jxor g1027(.dina(n1090), .dinb(n1058), .dout(n1091));
  jxor g1028(.dina(n1091), .dinb(n1056), .dout(n1092));
  jxor g1029(.dina(n1092), .dinb(n1053), .dout(n1093));
  jxor g1030(.dina(n1093), .dinb(n1051), .dout(n1094));
  jxor g1031(.dina(n1094), .dinb(n1048), .dout(n1095));
  jxor g1032(.dina(n1095), .dinb(n1046), .dout(n1096));
  jxor g1033(.dina(n1096), .dinb(n1043), .dout(n1097));
  jxor g1034(.dina(n1097), .dinb(n1041), .dout(n1098));
  jxor g1035(.dina(n1098), .dinb(n1038), .dout(n1099));
  jxor g1036(.dina(n1099), .dinb(n1036), .dout(n1100));
  jxor g1037(.dina(n1100), .dinb(n1033), .dout(n1101));
  jxor g1038(.dina(n1101), .dinb(n1031), .dout(n1102));
  jxor g1039(.dina(n1102), .dinb(n1028), .dout(n1103));
  jxor g1040(.dina(n1103), .dinb(n1026), .dout(n1104));
  jnot g1041(.din(n1104), .dout(n1105));
  jxor g1042(.dina(n1105), .dinb(n1023), .dout(n1106));
  jxor g1043(.dina(n1106), .dinb(n1022), .dout(n1107));
  jxor g1044(.dina(n1107), .dinb(n1018), .dout(n1108));
  jxor g1045(.dina(n1108), .dinb(n1017), .dout(n1109));
  jnot g1046(.din(n1109), .dout(n1110));
  jxor g1047(.dina(n1110), .dinb(n1013), .dout(G6160gat));
  jnot g1048(.din(n1108), .dout(n1112));
  jcb  g1049(.dina(n1112), .dinb(n1017), .dout(n1113));
  jcb  g1050(.dina(n1109), .dinb(n1013), .dout(n1114));
  jand g1051(.dina(n1114), .dinb(n1113), .dout(n1115));
  jnot g1052(.din(n1106), .dout(n1116));
  jcb  g1053(.dina(n1116), .dinb(n1022), .dout(n1117));
  jcb  g1054(.dina(n1107), .dinb(n1018), .dout(n1118));
  jand g1055(.dina(n1118), .dinb(n1117), .dout(n1119));
  jand g1056(.dina(G528gat), .dinb(G52gat), .dout(n1120));
  jand g1057(.dina(n1103), .dinb(n1026), .dout(n1121));
  jnot g1058(.din(n1121), .dout(n1122));
  jcb  g1059(.dina(n1105), .dinb(n1023), .dout(n1123));
  jand g1060(.dina(n1123), .dinb(n1122), .dout(n1124));
  jand g1061(.dina(G511gat), .dinb(G69gat), .dout(n1125));
  jnot g1062(.din(n1125), .dout(n1126));
  jand g1063(.dina(n1101), .dinb(n1031), .dout(n1127));
  jand g1064(.dina(n1102), .dinb(n1028), .dout(n1128));
  jcb  g1065(.dina(n1128), .dinb(n1127), .dout(n1129));
  jand g1066(.dina(G494gat), .dinb(G86gat), .dout(n1130));
  jnot g1067(.din(n1130), .dout(n1131));
  jand g1068(.dina(n1099), .dinb(n1036), .dout(n1132));
  jand g1069(.dina(n1100), .dinb(n1033), .dout(n1133));
  jcb  g1070(.dina(n1133), .dinb(n1132), .dout(n1134));
  jand g1071(.dina(G477gat), .dinb(G103gat), .dout(n1135));
  jnot g1072(.din(n1135), .dout(n1136));
  jand g1073(.dina(n1097), .dinb(n1041), .dout(n1137));
  jand g1074(.dina(n1098), .dinb(n1038), .dout(n1138));
  jcb  g1075(.dina(n1138), .dinb(n1137), .dout(n1139));
  jand g1076(.dina(G460gat), .dinb(G120gat), .dout(n1140));
  jnot g1077(.din(n1140), .dout(n1141));
  jand g1078(.dina(n1095), .dinb(n1046), .dout(n1142));
  jand g1079(.dina(n1096), .dinb(n1043), .dout(n1143));
  jcb  g1080(.dina(n1143), .dinb(n1142), .dout(n1144));
  jand g1081(.dina(G443gat), .dinb(G137gat), .dout(n1145));
  jnot g1082(.din(n1145), .dout(n1146));
  jand g1083(.dina(n1093), .dinb(n1051), .dout(n1147));
  jand g1084(.dina(n1094), .dinb(n1048), .dout(n1148));
  jcb  g1085(.dina(n1148), .dinb(n1147), .dout(n1149));
  jand g1086(.dina(G426gat), .dinb(G154gat), .dout(n1150));
  jnot g1087(.din(n1150), .dout(n1151));
  jand g1088(.dina(n1091), .dinb(n1056), .dout(n1152));
  jand g1089(.dina(n1092), .dinb(n1053), .dout(n1153));
  jcb  g1090(.dina(n1153), .dinb(n1152), .dout(n1154));
  jand g1091(.dina(G409gat), .dinb(G171gat), .dout(n1155));
  jnot g1092(.din(n1155), .dout(n1156));
  jand g1093(.dina(n1089), .dinb(n1061), .dout(n1157));
  jand g1094(.dina(n1090), .dinb(n1058), .dout(n1158));
  jcb  g1095(.dina(n1158), .dinb(n1157), .dout(n1159));
  jand g1096(.dina(G392gat), .dinb(G188gat), .dout(n1160));
  jnot g1097(.din(n1160), .dout(n1161));
  jand g1098(.dina(n1087), .dinb(n1066), .dout(n1162));
  jand g1099(.dina(n1088), .dinb(n1063), .dout(n1163));
  jcb  g1100(.dina(n1163), .dinb(n1162), .dout(n1164));
  jand g1101(.dina(G375gat), .dinb(G205gat), .dout(n1165));
  jnot g1102(.din(n1165), .dout(n1166));
  jand g1103(.dina(n1085), .dinb(n1071), .dout(n1167));
  jand g1104(.dina(n1086), .dinb(n1068), .dout(n1168));
  jcb  g1105(.dina(n1168), .dinb(n1167), .dout(n1169));
  jand g1106(.dina(G358gat), .dinb(G222gat), .dout(n1170));
  jnot g1107(.din(n1170), .dout(n1171));
  jand g1108(.dina(n1083), .dinb(n1076), .dout(n1172));
  jand g1109(.dina(n1084), .dinb(n1073), .dout(n1173));
  jcb  g1110(.dina(n1173), .dinb(n1172), .dout(n1174));
  jand g1111(.dina(G341gat), .dinb(G239gat), .dout(n1175));
  jand g1112(.dina(G324gat), .dinb(G256gat), .dout(n1176));
  jcb  g1113(.dina(n1080), .dinb(n1078), .dout(n1177));
  jcb  g1114(.dina(n1082), .dinb(n1077), .dout(n1178));
  jand g1115(.dina(n1178), .dinb(n1177), .dout(n1179));
  jxor g1116(.dina(n1179), .dinb(n1176), .dout(n1180));
  jnot g1117(.din(n1180), .dout(n1181));
  jxor g1118(.dina(n1181), .dinb(n1175), .dout(n1182));
  jxor g1119(.dina(n1182), .dinb(n1174), .dout(n1183));
  jxor g1120(.dina(n1183), .dinb(n1171), .dout(n1184));
  jxor g1121(.dina(n1184), .dinb(n1169), .dout(n1185));
  jxor g1122(.dina(n1185), .dinb(n1166), .dout(n1186));
  jxor g1123(.dina(n1186), .dinb(n1164), .dout(n1187));
  jxor g1124(.dina(n1187), .dinb(n1161), .dout(n1188));
  jxor g1125(.dina(n1188), .dinb(n1159), .dout(n1189));
  jxor g1126(.dina(n1189), .dinb(n1156), .dout(n1190));
  jxor g1127(.dina(n1190), .dinb(n1154), .dout(n1191));
  jxor g1128(.dina(n1191), .dinb(n1151), .dout(n1192));
  jxor g1129(.dina(n1192), .dinb(n1149), .dout(n1193));
  jxor g1130(.dina(n1193), .dinb(n1146), .dout(n1194));
  jxor g1131(.dina(n1194), .dinb(n1144), .dout(n1195));
  jxor g1132(.dina(n1195), .dinb(n1141), .dout(n1196));
  jxor g1133(.dina(n1196), .dinb(n1139), .dout(n1197));
  jxor g1134(.dina(n1197), .dinb(n1136), .dout(n1198));
  jxor g1135(.dina(n1198), .dinb(n1134), .dout(n1199));
  jxor g1136(.dina(n1199), .dinb(n1131), .dout(n1200));
  jxor g1137(.dina(n1200), .dinb(n1129), .dout(n1201));
  jxor g1138(.dina(n1201), .dinb(n1126), .dout(n1202));
  jnot g1139(.din(n1202), .dout(n1203));
  jxor g1140(.dina(n1203), .dinb(n1124), .dout(n1204));
  jnot g1141(.din(n1204), .dout(n1205));
  jxor g1142(.dina(n1205), .dinb(n1120), .dout(n1206));
  jxor g1143(.dina(n1206), .dinb(n1119), .dout(n1207));
  jnot g1144(.din(n1207), .dout(n1208));
  jxor g1145(.dina(n1208), .dinb(n1115), .dout(G6170gat));
  jnot g1146(.din(n1206), .dout(n1210));
  jcb  g1147(.dina(n1210), .dinb(n1119), .dout(n1211));
  jcb  g1148(.dina(n1207), .dinb(n1115), .dout(n1212));
  jand g1149(.dina(n1212), .dinb(n1211), .dout(n1213));
  jcb  g1150(.dina(n1203), .dinb(n1124), .dout(n1214));
  jcb  g1151(.dina(n1205), .dinb(n1120), .dout(n1215));
  jand g1152(.dina(n1215), .dinb(n1214), .dout(n1216));
  jand g1153(.dina(G528gat), .dinb(G69gat), .dout(n1217));
  jand g1154(.dina(n1200), .dinb(n1129), .dout(n1218));
  jand g1155(.dina(n1201), .dinb(n1126), .dout(n1219));
  jcb  g1156(.dina(n1219), .dinb(n1218), .dout(n1220));
  jand g1157(.dina(G511gat), .dinb(G86gat), .dout(n1221));
  jnot g1158(.din(n1221), .dout(n1222));
  jand g1159(.dina(n1198), .dinb(n1134), .dout(n1223));
  jand g1160(.dina(n1199), .dinb(n1131), .dout(n1224));
  jcb  g1161(.dina(n1224), .dinb(n1223), .dout(n1225));
  jand g1162(.dina(G494gat), .dinb(G103gat), .dout(n1226));
  jnot g1163(.din(n1226), .dout(n1227));
  jand g1164(.dina(n1196), .dinb(n1139), .dout(n1228));
  jand g1165(.dina(n1197), .dinb(n1136), .dout(n1229));
  jcb  g1166(.dina(n1229), .dinb(n1228), .dout(n1230));
  jand g1167(.dina(G477gat), .dinb(G120gat), .dout(n1231));
  jnot g1168(.din(n1231), .dout(n1232));
  jand g1169(.dina(n1194), .dinb(n1144), .dout(n1233));
  jand g1170(.dina(n1195), .dinb(n1141), .dout(n1234));
  jcb  g1171(.dina(n1234), .dinb(n1233), .dout(n1235));
  jand g1172(.dina(G460gat), .dinb(G137gat), .dout(n1236));
  jnot g1173(.din(n1236), .dout(n1237));
  jand g1174(.dina(n1192), .dinb(n1149), .dout(n1238));
  jand g1175(.dina(n1193), .dinb(n1146), .dout(n1239));
  jcb  g1176(.dina(n1239), .dinb(n1238), .dout(n1240));
  jand g1177(.dina(G443gat), .dinb(G154gat), .dout(n1241));
  jnot g1178(.din(n1241), .dout(n1242));
  jand g1179(.dina(n1190), .dinb(n1154), .dout(n1243));
  jand g1180(.dina(n1191), .dinb(n1151), .dout(n1244));
  jcb  g1181(.dina(n1244), .dinb(n1243), .dout(n1245));
  jand g1182(.dina(G426gat), .dinb(G171gat), .dout(n1246));
  jnot g1183(.din(n1246), .dout(n1247));
  jand g1184(.dina(n1188), .dinb(n1159), .dout(n1248));
  jand g1185(.dina(n1189), .dinb(n1156), .dout(n1249));
  jcb  g1186(.dina(n1249), .dinb(n1248), .dout(n1250));
  jand g1187(.dina(G409gat), .dinb(G188gat), .dout(n1251));
  jnot g1188(.din(n1251), .dout(n1252));
  jand g1189(.dina(n1186), .dinb(n1164), .dout(n1253));
  jand g1190(.dina(n1187), .dinb(n1161), .dout(n1254));
  jcb  g1191(.dina(n1254), .dinb(n1253), .dout(n1255));
  jand g1192(.dina(G392gat), .dinb(G205gat), .dout(n1256));
  jnot g1193(.din(n1256), .dout(n1257));
  jand g1194(.dina(n1184), .dinb(n1169), .dout(n1258));
  jand g1195(.dina(n1185), .dinb(n1166), .dout(n1259));
  jcb  g1196(.dina(n1259), .dinb(n1258), .dout(n1260));
  jand g1197(.dina(G375gat), .dinb(G222gat), .dout(n1261));
  jnot g1198(.din(n1261), .dout(n1262));
  jand g1199(.dina(n1182), .dinb(n1174), .dout(n1263));
  jand g1200(.dina(n1183), .dinb(n1171), .dout(n1264));
  jcb  g1201(.dina(n1264), .dinb(n1263), .dout(n1265));
  jand g1202(.dina(G358gat), .dinb(G239gat), .dout(n1266));
  jand g1203(.dina(G341gat), .dinb(G256gat), .dout(n1267));
  jcb  g1204(.dina(n1179), .dinb(n1176), .dout(n1268));
  jcb  g1205(.dina(n1181), .dinb(n1175), .dout(n1269));
  jand g1206(.dina(n1269), .dinb(n1268), .dout(n1270));
  jxor g1207(.dina(n1270), .dinb(n1267), .dout(n1271));
  jnot g1208(.din(n1271), .dout(n1272));
  jxor g1209(.dina(n1272), .dinb(n1266), .dout(n1273));
  jxor g1210(.dina(n1273), .dinb(n1265), .dout(n1274));
  jxor g1211(.dina(n1274), .dinb(n1262), .dout(n1275));
  jxor g1212(.dina(n1275), .dinb(n1260), .dout(n1276));
  jxor g1213(.dina(n1276), .dinb(n1257), .dout(n1277));
  jxor g1214(.dina(n1277), .dinb(n1255), .dout(n1278));
  jxor g1215(.dina(n1278), .dinb(n1252), .dout(n1279));
  jxor g1216(.dina(n1279), .dinb(n1250), .dout(n1280));
  jxor g1217(.dina(n1280), .dinb(n1247), .dout(n1281));
  jxor g1218(.dina(n1281), .dinb(n1245), .dout(n1282));
  jxor g1219(.dina(n1282), .dinb(n1242), .dout(n1283));
  jxor g1220(.dina(n1283), .dinb(n1240), .dout(n1284));
  jxor g1221(.dina(n1284), .dinb(n1237), .dout(n1285));
  jxor g1222(.dina(n1285), .dinb(n1235), .dout(n1286));
  jxor g1223(.dina(n1286), .dinb(n1232), .dout(n1287));
  jxor g1224(.dina(n1287), .dinb(n1230), .dout(n1288));
  jxor g1225(.dina(n1288), .dinb(n1227), .dout(n1289));
  jxor g1226(.dina(n1289), .dinb(n1225), .dout(n1290));
  jxor g1227(.dina(n1290), .dinb(n1222), .dout(n1291));
  jxor g1228(.dina(n1291), .dinb(n1220), .dout(n1292));
  jnot g1229(.din(n1292), .dout(n1293));
  jxor g1230(.dina(n1293), .dinb(n1217), .dout(n1294));
  jxor g1231(.dina(n1294), .dinb(n1216), .dout(n1295));
  jnot g1232(.din(n1295), .dout(n1296));
  jxor g1233(.dina(n1296), .dinb(n1213), .dout(G6180gat));
  jnot g1234(.din(n1294), .dout(n1298));
  jcb  g1235(.dina(n1298), .dinb(n1216), .dout(n1299));
  jcb  g1236(.dina(n1295), .dinb(n1213), .dout(n1300));
  jand g1237(.dina(n1300), .dinb(n1299), .dout(n1301));
  jnot g1238(.din(n1220), .dout(n1302));
  jnot g1239(.din(n1291), .dout(n1303));
  jcb  g1240(.dina(n1303), .dinb(n1302), .dout(n1304));
  jcb  g1241(.dina(n1293), .dinb(n1217), .dout(n1305));
  jand g1242(.dina(n1305), .dinb(n1304), .dout(n1306));
  jand g1243(.dina(G528gat), .dinb(G86gat), .dout(n1307));
  jand g1244(.dina(n1289), .dinb(n1225), .dout(n1308));
  jand g1245(.dina(n1290), .dinb(n1222), .dout(n1309));
  jcb  g1246(.dina(n1309), .dinb(n1308), .dout(n1310));
  jand g1247(.dina(G511gat), .dinb(G103gat), .dout(n1311));
  jnot g1248(.din(n1311), .dout(n1312));
  jand g1249(.dina(n1287), .dinb(n1230), .dout(n1313));
  jand g1250(.dina(n1288), .dinb(n1227), .dout(n1314));
  jcb  g1251(.dina(n1314), .dinb(n1313), .dout(n1315));
  jand g1252(.dina(G494gat), .dinb(G120gat), .dout(n1316));
  jnot g1253(.din(n1316), .dout(n1317));
  jand g1254(.dina(n1285), .dinb(n1235), .dout(n1318));
  jand g1255(.dina(n1286), .dinb(n1232), .dout(n1319));
  jcb  g1256(.dina(n1319), .dinb(n1318), .dout(n1320));
  jand g1257(.dina(G477gat), .dinb(G137gat), .dout(n1321));
  jnot g1258(.din(n1321), .dout(n1322));
  jand g1259(.dina(n1283), .dinb(n1240), .dout(n1323));
  jand g1260(.dina(n1284), .dinb(n1237), .dout(n1324));
  jcb  g1261(.dina(n1324), .dinb(n1323), .dout(n1325));
  jand g1262(.dina(G460gat), .dinb(G154gat), .dout(n1326));
  jnot g1263(.din(n1326), .dout(n1327));
  jand g1264(.dina(n1281), .dinb(n1245), .dout(n1328));
  jand g1265(.dina(n1282), .dinb(n1242), .dout(n1329));
  jcb  g1266(.dina(n1329), .dinb(n1328), .dout(n1330));
  jand g1267(.dina(G443gat), .dinb(G171gat), .dout(n1331));
  jnot g1268(.din(n1331), .dout(n1332));
  jand g1269(.dina(n1279), .dinb(n1250), .dout(n1333));
  jand g1270(.dina(n1280), .dinb(n1247), .dout(n1334));
  jcb  g1271(.dina(n1334), .dinb(n1333), .dout(n1335));
  jand g1272(.dina(G426gat), .dinb(G188gat), .dout(n1336));
  jnot g1273(.din(n1336), .dout(n1337));
  jand g1274(.dina(n1277), .dinb(n1255), .dout(n1338));
  jand g1275(.dina(n1278), .dinb(n1252), .dout(n1339));
  jcb  g1276(.dina(n1339), .dinb(n1338), .dout(n1340));
  jand g1277(.dina(G409gat), .dinb(G205gat), .dout(n1341));
  jnot g1278(.din(n1341), .dout(n1342));
  jand g1279(.dina(n1275), .dinb(n1260), .dout(n1343));
  jand g1280(.dina(n1276), .dinb(n1257), .dout(n1344));
  jcb  g1281(.dina(n1344), .dinb(n1343), .dout(n1345));
  jand g1282(.dina(G392gat), .dinb(G222gat), .dout(n1346));
  jnot g1283(.din(n1346), .dout(n1347));
  jand g1284(.dina(n1273), .dinb(n1265), .dout(n1348));
  jand g1285(.dina(n1274), .dinb(n1262), .dout(n1349));
  jcb  g1286(.dina(n1349), .dinb(n1348), .dout(n1350));
  jand g1287(.dina(G375gat), .dinb(G239gat), .dout(n1351));
  jand g1288(.dina(G358gat), .dinb(G256gat), .dout(n1352));
  jcb  g1289(.dina(n1270), .dinb(n1267), .dout(n1353));
  jcb  g1290(.dina(n1272), .dinb(n1266), .dout(n1354));
  jand g1291(.dina(n1354), .dinb(n1353), .dout(n1355));
  jxor g1292(.dina(n1355), .dinb(n1352), .dout(n1356));
  jnot g1293(.din(n1356), .dout(n1357));
  jxor g1294(.dina(n1357), .dinb(n1351), .dout(n1358));
  jxor g1295(.dina(n1358), .dinb(n1350), .dout(n1359));
  jxor g1296(.dina(n1359), .dinb(n1347), .dout(n1360));
  jxor g1297(.dina(n1360), .dinb(n1345), .dout(n1361));
  jxor g1298(.dina(n1361), .dinb(n1342), .dout(n1362));
  jxor g1299(.dina(n1362), .dinb(n1340), .dout(n1363));
  jxor g1300(.dina(n1363), .dinb(n1337), .dout(n1364));
  jxor g1301(.dina(n1364), .dinb(n1335), .dout(n1365));
  jxor g1302(.dina(n1365), .dinb(n1332), .dout(n1366));
  jxor g1303(.dina(n1366), .dinb(n1330), .dout(n1367));
  jxor g1304(.dina(n1367), .dinb(n1327), .dout(n1368));
  jxor g1305(.dina(n1368), .dinb(n1325), .dout(n1369));
  jxor g1306(.dina(n1369), .dinb(n1322), .dout(n1370));
  jxor g1307(.dina(n1370), .dinb(n1320), .dout(n1371));
  jxor g1308(.dina(n1371), .dinb(n1317), .dout(n1372));
  jxor g1309(.dina(n1372), .dinb(n1315), .dout(n1373));
  jxor g1310(.dina(n1373), .dinb(n1312), .dout(n1374));
  jxor g1311(.dina(n1374), .dinb(n1310), .dout(n1375));
  jnot g1312(.din(n1375), .dout(n1376));
  jxor g1313(.dina(n1376), .dinb(n1307), .dout(n1377));
  jnot g1314(.din(n1377), .dout(n1378));
  jxor g1315(.dina(n1378), .dinb(n1306), .dout(n1379));
  jxor g1316(.dina(n1379), .dinb(n1301), .dout(G6190gat));
  jcb  g1317(.dina(n1378), .dinb(n1306), .dout(n1381));
  jnot g1318(.din(n1379), .dout(n1382));
  jcb  g1319(.dina(n1382), .dinb(n1301), .dout(n1383));
  jand g1320(.dina(n1383), .dinb(n1381), .dout(n1384));
  jnot g1321(.din(n1310), .dout(n1385));
  jnot g1322(.din(n1374), .dout(n1386));
  jcb  g1323(.dina(n1386), .dinb(n1385), .dout(n1387));
  jcb  g1324(.dina(n1376), .dinb(n1307), .dout(n1388));
  jand g1325(.dina(n1388), .dinb(n1387), .dout(n1389));
  jand g1326(.dina(G528gat), .dinb(G103gat), .dout(n1390));
  jand g1327(.dina(n1372), .dinb(n1315), .dout(n1391));
  jand g1328(.dina(n1373), .dinb(n1312), .dout(n1392));
  jcb  g1329(.dina(n1392), .dinb(n1391), .dout(n1393));
  jand g1330(.dina(G511gat), .dinb(G120gat), .dout(n1394));
  jnot g1331(.din(n1394), .dout(n1395));
  jand g1332(.dina(n1370), .dinb(n1320), .dout(n1396));
  jand g1333(.dina(n1371), .dinb(n1317), .dout(n1397));
  jcb  g1334(.dina(n1397), .dinb(n1396), .dout(n1398));
  jand g1335(.dina(G494gat), .dinb(G137gat), .dout(n1399));
  jnot g1336(.din(n1399), .dout(n1400));
  jand g1337(.dina(n1368), .dinb(n1325), .dout(n1401));
  jand g1338(.dina(n1369), .dinb(n1322), .dout(n1402));
  jcb  g1339(.dina(n1402), .dinb(n1401), .dout(n1403));
  jand g1340(.dina(G477gat), .dinb(G154gat), .dout(n1404));
  jnot g1341(.din(n1404), .dout(n1405));
  jand g1342(.dina(n1366), .dinb(n1330), .dout(n1406));
  jand g1343(.dina(n1367), .dinb(n1327), .dout(n1407));
  jcb  g1344(.dina(n1407), .dinb(n1406), .dout(n1408));
  jand g1345(.dina(G460gat), .dinb(G171gat), .dout(n1409));
  jnot g1346(.din(n1409), .dout(n1410));
  jand g1347(.dina(n1364), .dinb(n1335), .dout(n1411));
  jand g1348(.dina(n1365), .dinb(n1332), .dout(n1412));
  jcb  g1349(.dina(n1412), .dinb(n1411), .dout(n1413));
  jand g1350(.dina(G443gat), .dinb(G188gat), .dout(n1414));
  jnot g1351(.din(n1414), .dout(n1415));
  jand g1352(.dina(n1362), .dinb(n1340), .dout(n1416));
  jand g1353(.dina(n1363), .dinb(n1337), .dout(n1417));
  jcb  g1354(.dina(n1417), .dinb(n1416), .dout(n1418));
  jand g1355(.dina(G426gat), .dinb(G205gat), .dout(n1419));
  jnot g1356(.din(n1419), .dout(n1420));
  jand g1357(.dina(n1360), .dinb(n1345), .dout(n1421));
  jand g1358(.dina(n1361), .dinb(n1342), .dout(n1422));
  jcb  g1359(.dina(n1422), .dinb(n1421), .dout(n1423));
  jand g1360(.dina(G409gat), .dinb(G222gat), .dout(n1424));
  jnot g1361(.din(n1424), .dout(n1425));
  jand g1362(.dina(n1358), .dinb(n1350), .dout(n1426));
  jand g1363(.dina(n1359), .dinb(n1347), .dout(n1427));
  jcb  g1364(.dina(n1427), .dinb(n1426), .dout(n1428));
  jand g1365(.dina(G392gat), .dinb(G239gat), .dout(n1429));
  jand g1366(.dina(G375gat), .dinb(G256gat), .dout(n1430));
  jcb  g1367(.dina(n1355), .dinb(n1352), .dout(n1431));
  jcb  g1368(.dina(n1357), .dinb(n1351), .dout(n1432));
  jand g1369(.dina(n1432), .dinb(n1431), .dout(n1433));
  jxor g1370(.dina(n1433), .dinb(n1430), .dout(n1434));
  jnot g1371(.din(n1434), .dout(n1435));
  jxor g1372(.dina(n1435), .dinb(n1429), .dout(n1436));
  jxor g1373(.dina(n1436), .dinb(n1428), .dout(n1437));
  jxor g1374(.dina(n1437), .dinb(n1425), .dout(n1438));
  jxor g1375(.dina(n1438), .dinb(n1423), .dout(n1439));
  jxor g1376(.dina(n1439), .dinb(n1420), .dout(n1440));
  jxor g1377(.dina(n1440), .dinb(n1418), .dout(n1441));
  jxor g1378(.dina(n1441), .dinb(n1415), .dout(n1442));
  jxor g1379(.dina(n1442), .dinb(n1413), .dout(n1443));
  jxor g1380(.dina(n1443), .dinb(n1410), .dout(n1444));
  jxor g1381(.dina(n1444), .dinb(n1408), .dout(n1445));
  jxor g1382(.dina(n1445), .dinb(n1405), .dout(n1446));
  jxor g1383(.dina(n1446), .dinb(n1403), .dout(n1447));
  jxor g1384(.dina(n1447), .dinb(n1400), .dout(n1448));
  jxor g1385(.dina(n1448), .dinb(n1398), .dout(n1449));
  jxor g1386(.dina(n1449), .dinb(n1395), .dout(n1450));
  jxor g1387(.dina(n1450), .dinb(n1393), .dout(n1451));
  jnot g1388(.din(n1451), .dout(n1452));
  jxor g1389(.dina(n1452), .dinb(n1390), .dout(n1453));
  jnot g1390(.din(n1453), .dout(n1454));
  jxor g1391(.dina(n1454), .dinb(n1389), .dout(n1455));
  jxor g1392(.dina(n1455), .dinb(n1384), .dout(G6200gat));
  jcb  g1393(.dina(n1454), .dinb(n1389), .dout(n1457));
  jnot g1394(.din(n1455), .dout(n1458));
  jcb  g1395(.dina(n1458), .dinb(n1384), .dout(n1459));
  jand g1396(.dina(n1459), .dinb(n1457), .dout(n1460));
  jnot g1397(.din(n1393), .dout(n1461));
  jnot g1398(.din(n1450), .dout(n1462));
  jcb  g1399(.dina(n1462), .dinb(n1461), .dout(n1463));
  jcb  g1400(.dina(n1452), .dinb(n1390), .dout(n1464));
  jand g1401(.dina(n1464), .dinb(n1463), .dout(n1465));
  jand g1402(.dina(G528gat), .dinb(G120gat), .dout(n1466));
  jand g1403(.dina(n1448), .dinb(n1398), .dout(n1467));
  jand g1404(.dina(n1449), .dinb(n1395), .dout(n1468));
  jcb  g1405(.dina(n1468), .dinb(n1467), .dout(n1469));
  jand g1406(.dina(G511gat), .dinb(G137gat), .dout(n1470));
  jnot g1407(.din(n1470), .dout(n1471));
  jand g1408(.dina(n1446), .dinb(n1403), .dout(n1472));
  jand g1409(.dina(n1447), .dinb(n1400), .dout(n1473));
  jcb  g1410(.dina(n1473), .dinb(n1472), .dout(n1474));
  jand g1411(.dina(G494gat), .dinb(G154gat), .dout(n1475));
  jnot g1412(.din(n1475), .dout(n1476));
  jand g1413(.dina(n1444), .dinb(n1408), .dout(n1477));
  jand g1414(.dina(n1445), .dinb(n1405), .dout(n1478));
  jcb  g1415(.dina(n1478), .dinb(n1477), .dout(n1479));
  jand g1416(.dina(G477gat), .dinb(G171gat), .dout(n1480));
  jnot g1417(.din(n1480), .dout(n1481));
  jand g1418(.dina(n1442), .dinb(n1413), .dout(n1482));
  jand g1419(.dina(n1443), .dinb(n1410), .dout(n1483));
  jcb  g1420(.dina(n1483), .dinb(n1482), .dout(n1484));
  jand g1421(.dina(G460gat), .dinb(G188gat), .dout(n1485));
  jnot g1422(.din(n1485), .dout(n1486));
  jand g1423(.dina(n1440), .dinb(n1418), .dout(n1487));
  jand g1424(.dina(n1441), .dinb(n1415), .dout(n1488));
  jcb  g1425(.dina(n1488), .dinb(n1487), .dout(n1489));
  jand g1426(.dina(G443gat), .dinb(G205gat), .dout(n1490));
  jnot g1427(.din(n1490), .dout(n1491));
  jand g1428(.dina(n1438), .dinb(n1423), .dout(n1492));
  jand g1429(.dina(n1439), .dinb(n1420), .dout(n1493));
  jcb  g1430(.dina(n1493), .dinb(n1492), .dout(n1494));
  jand g1431(.dina(G426gat), .dinb(G222gat), .dout(n1495));
  jnot g1432(.din(n1495), .dout(n1496));
  jand g1433(.dina(n1436), .dinb(n1428), .dout(n1497));
  jand g1434(.dina(n1437), .dinb(n1425), .dout(n1498));
  jcb  g1435(.dina(n1498), .dinb(n1497), .dout(n1499));
  jand g1436(.dina(G409gat), .dinb(G239gat), .dout(n1500));
  jand g1437(.dina(G392gat), .dinb(G256gat), .dout(n1501));
  jcb  g1438(.dina(n1433), .dinb(n1430), .dout(n1502));
  jcb  g1439(.dina(n1435), .dinb(n1429), .dout(n1503));
  jand g1440(.dina(n1503), .dinb(n1502), .dout(n1504));
  jxor g1441(.dina(n1504), .dinb(n1501), .dout(n1505));
  jnot g1442(.din(n1505), .dout(n1506));
  jxor g1443(.dina(n1506), .dinb(n1500), .dout(n1507));
  jxor g1444(.dina(n1507), .dinb(n1499), .dout(n1508));
  jxor g1445(.dina(n1508), .dinb(n1496), .dout(n1509));
  jxor g1446(.dina(n1509), .dinb(n1494), .dout(n1510));
  jxor g1447(.dina(n1510), .dinb(n1491), .dout(n1511));
  jxor g1448(.dina(n1511), .dinb(n1489), .dout(n1512));
  jxor g1449(.dina(n1512), .dinb(n1486), .dout(n1513));
  jxor g1450(.dina(n1513), .dinb(n1484), .dout(n1514));
  jxor g1451(.dina(n1514), .dinb(n1481), .dout(n1515));
  jxor g1452(.dina(n1515), .dinb(n1479), .dout(n1516));
  jxor g1453(.dina(n1516), .dinb(n1476), .dout(n1517));
  jxor g1454(.dina(n1517), .dinb(n1474), .dout(n1518));
  jxor g1455(.dina(n1518), .dinb(n1471), .dout(n1519));
  jxor g1456(.dina(n1519), .dinb(n1469), .dout(n1520));
  jnot g1457(.din(n1520), .dout(n1521));
  jxor g1458(.dina(n1521), .dinb(n1466), .dout(n1522));
  jnot g1459(.din(n1522), .dout(n1523));
  jxor g1460(.dina(n1523), .dinb(n1465), .dout(n1524));
  jxor g1461(.dina(n1524), .dinb(n1460), .dout(G6210gat));
  jcb  g1462(.dina(n1523), .dinb(n1465), .dout(n1526));
  jnot g1463(.din(n1524), .dout(n1527));
  jcb  g1464(.dina(n1527), .dinb(n1460), .dout(n1528));
  jand g1465(.dina(n1528), .dinb(n1526), .dout(n1529));
  jnot g1466(.din(n1469), .dout(n1530));
  jnot g1467(.din(n1519), .dout(n1531));
  jcb  g1468(.dina(n1531), .dinb(n1530), .dout(n1532));
  jcb  g1469(.dina(n1521), .dinb(n1466), .dout(n1533));
  jand g1470(.dina(n1533), .dinb(n1532), .dout(n1534));
  jand g1471(.dina(G528gat), .dinb(G137gat), .dout(n1535));
  jand g1472(.dina(n1517), .dinb(n1474), .dout(n1536));
  jand g1473(.dina(n1518), .dinb(n1471), .dout(n1537));
  jcb  g1474(.dina(n1537), .dinb(n1536), .dout(n1538));
  jand g1475(.dina(G511gat), .dinb(G154gat), .dout(n1539));
  jnot g1476(.din(n1539), .dout(n1540));
  jand g1477(.dina(n1515), .dinb(n1479), .dout(n1541));
  jand g1478(.dina(n1516), .dinb(n1476), .dout(n1542));
  jcb  g1479(.dina(n1542), .dinb(n1541), .dout(n1543));
  jand g1480(.dina(G494gat), .dinb(G171gat), .dout(n1544));
  jnot g1481(.din(n1544), .dout(n1545));
  jand g1482(.dina(n1513), .dinb(n1484), .dout(n1546));
  jand g1483(.dina(n1514), .dinb(n1481), .dout(n1547));
  jcb  g1484(.dina(n1547), .dinb(n1546), .dout(n1548));
  jand g1485(.dina(G477gat), .dinb(G188gat), .dout(n1549));
  jnot g1486(.din(n1549), .dout(n1550));
  jand g1487(.dina(n1511), .dinb(n1489), .dout(n1551));
  jand g1488(.dina(n1512), .dinb(n1486), .dout(n1552));
  jcb  g1489(.dina(n1552), .dinb(n1551), .dout(n1553));
  jand g1490(.dina(G460gat), .dinb(G205gat), .dout(n1554));
  jnot g1491(.din(n1554), .dout(n1555));
  jand g1492(.dina(n1509), .dinb(n1494), .dout(n1556));
  jand g1493(.dina(n1510), .dinb(n1491), .dout(n1557));
  jcb  g1494(.dina(n1557), .dinb(n1556), .dout(n1558));
  jand g1495(.dina(G443gat), .dinb(G222gat), .dout(n1559));
  jnot g1496(.din(n1559), .dout(n1560));
  jand g1497(.dina(n1507), .dinb(n1499), .dout(n1561));
  jand g1498(.dina(n1508), .dinb(n1496), .dout(n1562));
  jcb  g1499(.dina(n1562), .dinb(n1561), .dout(n1563));
  jand g1500(.dina(G426gat), .dinb(G239gat), .dout(n1564));
  jand g1501(.dina(G409gat), .dinb(G256gat), .dout(n1565));
  jcb  g1502(.dina(n1504), .dinb(n1501), .dout(n1566));
  jcb  g1503(.dina(n1506), .dinb(n1500), .dout(n1567));
  jand g1504(.dina(n1567), .dinb(n1566), .dout(n1568));
  jxor g1505(.dina(n1568), .dinb(n1565), .dout(n1569));
  jnot g1506(.din(n1569), .dout(n1570));
  jxor g1507(.dina(n1570), .dinb(n1564), .dout(n1571));
  jxor g1508(.dina(n1571), .dinb(n1563), .dout(n1572));
  jxor g1509(.dina(n1572), .dinb(n1560), .dout(n1573));
  jxor g1510(.dina(n1573), .dinb(n1558), .dout(n1574));
  jxor g1511(.dina(n1574), .dinb(n1555), .dout(n1575));
  jxor g1512(.dina(n1575), .dinb(n1553), .dout(n1576));
  jxor g1513(.dina(n1576), .dinb(n1550), .dout(n1577));
  jxor g1514(.dina(n1577), .dinb(n1548), .dout(n1578));
  jxor g1515(.dina(n1578), .dinb(n1545), .dout(n1579));
  jxor g1516(.dina(n1579), .dinb(n1543), .dout(n1580));
  jxor g1517(.dina(n1580), .dinb(n1540), .dout(n1581));
  jxor g1518(.dina(n1581), .dinb(n1538), .dout(n1582));
  jnot g1519(.din(n1582), .dout(n1583));
  jxor g1520(.dina(n1583), .dinb(n1535), .dout(n1584));
  jnot g1521(.din(n1584), .dout(n1585));
  jxor g1522(.dina(n1585), .dinb(n1534), .dout(n1586));
  jxor g1523(.dina(n1586), .dinb(n1529), .dout(G6220gat));
  jcb  g1524(.dina(n1585), .dinb(n1534), .dout(n1588));
  jnot g1525(.din(n1586), .dout(n1589));
  jcb  g1526(.dina(n1589), .dinb(n1529), .dout(n1590));
  jand g1527(.dina(n1590), .dinb(n1588), .dout(n1591));
  jnot g1528(.din(n1538), .dout(n1592));
  jnot g1529(.din(n1581), .dout(n1593));
  jcb  g1530(.dina(n1593), .dinb(n1592), .dout(n1594));
  jcb  g1531(.dina(n1583), .dinb(n1535), .dout(n1595));
  jand g1532(.dina(n1595), .dinb(n1594), .dout(n1596));
  jand g1533(.dina(G528gat), .dinb(G154gat), .dout(n1597));
  jand g1534(.dina(n1579), .dinb(n1543), .dout(n1598));
  jand g1535(.dina(n1580), .dinb(n1540), .dout(n1599));
  jcb  g1536(.dina(n1599), .dinb(n1598), .dout(n1600));
  jand g1537(.dina(G511gat), .dinb(G171gat), .dout(n1601));
  jnot g1538(.din(n1601), .dout(n1602));
  jand g1539(.dina(n1577), .dinb(n1548), .dout(n1603));
  jand g1540(.dina(n1578), .dinb(n1545), .dout(n1604));
  jcb  g1541(.dina(n1604), .dinb(n1603), .dout(n1605));
  jand g1542(.dina(G494gat), .dinb(G188gat), .dout(n1606));
  jnot g1543(.din(n1606), .dout(n1607));
  jand g1544(.dina(n1575), .dinb(n1553), .dout(n1608));
  jand g1545(.dina(n1576), .dinb(n1550), .dout(n1609));
  jcb  g1546(.dina(n1609), .dinb(n1608), .dout(n1610));
  jand g1547(.dina(G477gat), .dinb(G205gat), .dout(n1611));
  jnot g1548(.din(n1611), .dout(n1612));
  jand g1549(.dina(n1573), .dinb(n1558), .dout(n1613));
  jand g1550(.dina(n1574), .dinb(n1555), .dout(n1614));
  jcb  g1551(.dina(n1614), .dinb(n1613), .dout(n1615));
  jand g1552(.dina(G460gat), .dinb(G222gat), .dout(n1616));
  jnot g1553(.din(n1616), .dout(n1617));
  jand g1554(.dina(n1571), .dinb(n1563), .dout(n1618));
  jand g1555(.dina(n1572), .dinb(n1560), .dout(n1619));
  jcb  g1556(.dina(n1619), .dinb(n1618), .dout(n1620));
  jand g1557(.dina(G443gat), .dinb(G239gat), .dout(n1621));
  jand g1558(.dina(G426gat), .dinb(G256gat), .dout(n1622));
  jcb  g1559(.dina(n1568), .dinb(n1565), .dout(n1623));
  jcb  g1560(.dina(n1570), .dinb(n1564), .dout(n1624));
  jand g1561(.dina(n1624), .dinb(n1623), .dout(n1625));
  jxor g1562(.dina(n1625), .dinb(n1622), .dout(n1626));
  jnot g1563(.din(n1626), .dout(n1627));
  jxor g1564(.dina(n1627), .dinb(n1621), .dout(n1628));
  jxor g1565(.dina(n1628), .dinb(n1620), .dout(n1629));
  jxor g1566(.dina(n1629), .dinb(n1617), .dout(n1630));
  jxor g1567(.dina(n1630), .dinb(n1615), .dout(n1631));
  jxor g1568(.dina(n1631), .dinb(n1612), .dout(n1632));
  jxor g1569(.dina(n1632), .dinb(n1610), .dout(n1633));
  jxor g1570(.dina(n1633), .dinb(n1607), .dout(n1634));
  jxor g1571(.dina(n1634), .dinb(n1605), .dout(n1635));
  jxor g1572(.dina(n1635), .dinb(n1602), .dout(n1636));
  jxor g1573(.dina(n1636), .dinb(n1600), .dout(n1637));
  jnot g1574(.din(n1637), .dout(n1638));
  jxor g1575(.dina(n1638), .dinb(n1597), .dout(n1639));
  jnot g1576(.din(n1639), .dout(n1640));
  jxor g1577(.dina(n1640), .dinb(n1596), .dout(n1641));
  jxor g1578(.dina(n1641), .dinb(n1591), .dout(G6230gat));
  jcb  g1579(.dina(n1640), .dinb(n1596), .dout(n1643));
  jnot g1580(.din(n1641), .dout(n1644));
  jcb  g1581(.dina(n1644), .dinb(n1591), .dout(n1645));
  jand g1582(.dina(n1645), .dinb(n1643), .dout(n1646));
  jnot g1583(.din(n1600), .dout(n1647));
  jnot g1584(.din(n1636), .dout(n1648));
  jcb  g1585(.dina(n1648), .dinb(n1647), .dout(n1649));
  jcb  g1586(.dina(n1638), .dinb(n1597), .dout(n1650));
  jand g1587(.dina(n1650), .dinb(n1649), .dout(n1651));
  jand g1588(.dina(G528gat), .dinb(G171gat), .dout(n1652));
  jnot g1589(.din(n1652), .dout(n1653));
  jand g1590(.dina(n1634), .dinb(n1605), .dout(n1654));
  jand g1591(.dina(n1635), .dinb(n1602), .dout(n1655));
  jcb  g1592(.dina(n1655), .dinb(n1654), .dout(n1656));
  jand g1593(.dina(G511gat), .dinb(G188gat), .dout(n1657));
  jnot g1594(.din(n1657), .dout(n1658));
  jand g1595(.dina(n1632), .dinb(n1610), .dout(n1659));
  jand g1596(.dina(n1633), .dinb(n1607), .dout(n1660));
  jcb  g1597(.dina(n1660), .dinb(n1659), .dout(n1661));
  jand g1598(.dina(G494gat), .dinb(G205gat), .dout(n1662));
  jnot g1599(.din(n1662), .dout(n1663));
  jand g1600(.dina(n1630), .dinb(n1615), .dout(n1664));
  jand g1601(.dina(n1631), .dinb(n1612), .dout(n1665));
  jcb  g1602(.dina(n1665), .dinb(n1664), .dout(n1666));
  jand g1603(.dina(G477gat), .dinb(G222gat), .dout(n1667));
  jnot g1604(.din(n1667), .dout(n1668));
  jand g1605(.dina(n1628), .dinb(n1620), .dout(n1669));
  jand g1606(.dina(n1629), .dinb(n1617), .dout(n1670));
  jcb  g1607(.dina(n1670), .dinb(n1669), .dout(n1671));
  jand g1608(.dina(G460gat), .dinb(G239gat), .dout(n1672));
  jand g1609(.dina(G443gat), .dinb(G256gat), .dout(n1673));
  jcb  g1610(.dina(n1625), .dinb(n1622), .dout(n1674));
  jcb  g1611(.dina(n1627), .dinb(n1621), .dout(n1675));
  jand g1612(.dina(n1675), .dinb(n1674), .dout(n1676));
  jxor g1613(.dina(n1676), .dinb(n1673), .dout(n1677));
  jnot g1614(.din(n1677), .dout(n1678));
  jxor g1615(.dina(n1678), .dinb(n1672), .dout(n1679));
  jxor g1616(.dina(n1679), .dinb(n1671), .dout(n1680));
  jxor g1617(.dina(n1680), .dinb(n1668), .dout(n1681));
  jxor g1618(.dina(n1681), .dinb(n1666), .dout(n1682));
  jxor g1619(.dina(n1682), .dinb(n1663), .dout(n1683));
  jxor g1620(.dina(n1683), .dinb(n1661), .dout(n1684));
  jxor g1621(.dina(n1684), .dinb(n1658), .dout(n1685));
  jxor g1622(.dina(n1685), .dinb(n1656), .dout(n1686));
  jxor g1623(.dina(n1686), .dinb(n1653), .dout(n1687));
  jnot g1624(.din(n1687), .dout(n1688));
  jxor g1625(.dina(n1688), .dinb(n1651), .dout(n1689));
  jxor g1626(.dina(n1689), .dinb(n1646), .dout(G6240gat));
  jcb  g1627(.dina(n1688), .dinb(n1651), .dout(n1691));
  jnot g1628(.din(n1689), .dout(n1692));
  jcb  g1629(.dina(n1692), .dinb(n1646), .dout(n1693));
  jand g1630(.dina(n1693), .dinb(n1691), .dout(n1694));
  jand g1631(.dina(n1685), .dinb(n1656), .dout(n1695));
  jand g1632(.dina(n1686), .dinb(n1653), .dout(n1696));
  jcb  g1633(.dina(n1696), .dinb(n1695), .dout(n1697));
  jand g1634(.dina(G528gat), .dinb(G188gat), .dout(n1698));
  jnot g1635(.din(n1698), .dout(n1699));
  jand g1636(.dina(n1683), .dinb(n1661), .dout(n1700));
  jand g1637(.dina(n1684), .dinb(n1658), .dout(n1701));
  jcb  g1638(.dina(n1701), .dinb(n1700), .dout(n1702));
  jand g1639(.dina(G511gat), .dinb(G205gat), .dout(n1703));
  jnot g1640(.din(n1703), .dout(n1704));
  jand g1641(.dina(n1681), .dinb(n1666), .dout(n1705));
  jand g1642(.dina(n1682), .dinb(n1663), .dout(n1706));
  jcb  g1643(.dina(n1706), .dinb(n1705), .dout(n1707));
  jand g1644(.dina(G494gat), .dinb(G222gat), .dout(n1708));
  jnot g1645(.din(n1708), .dout(n1709));
  jand g1646(.dina(n1679), .dinb(n1671), .dout(n1710));
  jand g1647(.dina(n1680), .dinb(n1668), .dout(n1711));
  jcb  g1648(.dina(n1711), .dinb(n1710), .dout(n1712));
  jand g1649(.dina(G477gat), .dinb(G239gat), .dout(n1713));
  jand g1650(.dina(G460gat), .dinb(G256gat), .dout(n1714));
  jcb  g1651(.dina(n1676), .dinb(n1673), .dout(n1715));
  jcb  g1652(.dina(n1678), .dinb(n1672), .dout(n1716));
  jand g1653(.dina(n1716), .dinb(n1715), .dout(n1717));
  jxor g1654(.dina(n1717), .dinb(n1714), .dout(n1718));
  jnot g1655(.din(n1718), .dout(n1719));
  jxor g1656(.dina(n1719), .dinb(n1713), .dout(n1720));
  jxor g1657(.dina(n1720), .dinb(n1712), .dout(n1721));
  jxor g1658(.dina(n1721), .dinb(n1709), .dout(n1722));
  jxor g1659(.dina(n1722), .dinb(n1707), .dout(n1723));
  jxor g1660(.dina(n1723), .dinb(n1704), .dout(n1724));
  jxor g1661(.dina(n1724), .dinb(n1702), .dout(n1725));
  jxor g1662(.dina(n1725), .dinb(n1699), .dout(n1726));
  jxor g1663(.dina(n1726), .dinb(n1697), .dout(n1727));
  jxor g1664(.dina(n1727), .dinb(n1694), .dout(G6250gat));
  jnot g1665(.din(n1697), .dout(n1729));
  jnot g1666(.din(n1726), .dout(n1730));
  jcb  g1667(.dina(n1730), .dinb(n1729), .dout(n1731));
  jnot g1668(.din(n1727), .dout(n1732));
  jcb  g1669(.dina(n1732), .dinb(n1694), .dout(n1733));
  jand g1670(.dina(n1733), .dinb(n1731), .dout(n1734));
  jand g1671(.dina(n1724), .dinb(n1702), .dout(n1735));
  jand g1672(.dina(n1725), .dinb(n1699), .dout(n1736));
  jcb  g1673(.dina(n1736), .dinb(n1735), .dout(n1737));
  jand g1674(.dina(G528gat), .dinb(G205gat), .dout(n1738));
  jnot g1675(.din(n1738), .dout(n1739));
  jand g1676(.dina(n1722), .dinb(n1707), .dout(n1740));
  jand g1677(.dina(n1723), .dinb(n1704), .dout(n1741));
  jcb  g1678(.dina(n1741), .dinb(n1740), .dout(n1742));
  jand g1679(.dina(G511gat), .dinb(G222gat), .dout(n1743));
  jnot g1680(.din(n1743), .dout(n1744));
  jand g1681(.dina(n1720), .dinb(n1712), .dout(n1745));
  jand g1682(.dina(n1721), .dinb(n1709), .dout(n1746));
  jcb  g1683(.dina(n1746), .dinb(n1745), .dout(n1747));
  jand g1684(.dina(G494gat), .dinb(G239gat), .dout(n1748));
  jand g1685(.dina(G477gat), .dinb(G256gat), .dout(n1749));
  jcb  g1686(.dina(n1717), .dinb(n1714), .dout(n1750));
  jcb  g1687(.dina(n1719), .dinb(n1713), .dout(n1751));
  jand g1688(.dina(n1751), .dinb(n1750), .dout(n1752));
  jxor g1689(.dina(n1752), .dinb(n1749), .dout(n1753));
  jnot g1690(.din(n1753), .dout(n1754));
  jxor g1691(.dina(n1754), .dinb(n1748), .dout(n1755));
  jxor g1692(.dina(n1755), .dinb(n1747), .dout(n1756));
  jxor g1693(.dina(n1756), .dinb(n1744), .dout(n1757));
  jxor g1694(.dina(n1757), .dinb(n1742), .dout(n1758));
  jxor g1695(.dina(n1758), .dinb(n1739), .dout(n1759));
  jxor g1696(.dina(n1759), .dinb(n1737), .dout(n1760));
  jxor g1697(.dina(n1760), .dinb(n1734), .dout(G6260gat));
  jnot g1698(.din(n1737), .dout(n1762));
  jnot g1699(.din(n1759), .dout(n1763));
  jcb  g1700(.dina(n1763), .dinb(n1762), .dout(n1764));
  jnot g1701(.din(n1760), .dout(n1765));
  jcb  g1702(.dina(n1765), .dinb(n1734), .dout(n1766));
  jand g1703(.dina(n1766), .dinb(n1764), .dout(n1767));
  jand g1704(.dina(n1757), .dinb(n1742), .dout(n1768));
  jand g1705(.dina(n1758), .dinb(n1739), .dout(n1769));
  jcb  g1706(.dina(n1769), .dinb(n1768), .dout(n1770));
  jand g1707(.dina(G528gat), .dinb(G222gat), .dout(n1771));
  jnot g1708(.din(n1771), .dout(n1772));
  jand g1709(.dina(n1755), .dinb(n1747), .dout(n1773));
  jand g1710(.dina(n1756), .dinb(n1744), .dout(n1774));
  jcb  g1711(.dina(n1774), .dinb(n1773), .dout(n1775));
  jand g1712(.dina(G511gat), .dinb(G239gat), .dout(n1776));
  jand g1713(.dina(G494gat), .dinb(G256gat), .dout(n1777));
  jcb  g1714(.dina(n1752), .dinb(n1749), .dout(n1778));
  jcb  g1715(.dina(n1754), .dinb(n1748), .dout(n1779));
  jand g1716(.dina(n1779), .dinb(n1778), .dout(n1780));
  jxor g1717(.dina(n1780), .dinb(n1777), .dout(n1781));
  jnot g1718(.din(n1781), .dout(n1782));
  jxor g1719(.dina(n1782), .dinb(n1776), .dout(n1783));
  jxor g1720(.dina(n1783), .dinb(n1775), .dout(n1784));
  jxor g1721(.dina(n1784), .dinb(n1772), .dout(n1785));
  jxor g1722(.dina(n1785), .dinb(n1770), .dout(n1786));
  jxor g1723(.dina(n1786), .dinb(n1767), .dout(G6270gat));
  jnot g1724(.din(n1770), .dout(n1788));
  jnot g1725(.din(n1785), .dout(n1789));
  jcb  g1726(.dina(n1789), .dinb(n1788), .dout(n1790));
  jnot g1727(.din(n1786), .dout(n1791));
  jcb  g1728(.dina(n1791), .dinb(n1767), .dout(n1792));
  jand g1729(.dina(n1792), .dinb(n1790), .dout(n1793));
  jand g1730(.dina(n1783), .dinb(n1775), .dout(n1794));
  jand g1731(.dina(n1784), .dinb(n1772), .dout(n1795));
  jcb  g1732(.dina(n1795), .dinb(n1794), .dout(n1796));
  jand g1733(.dina(G528gat), .dinb(G239gat), .dout(n1797));
  jand g1734(.dina(G511gat), .dinb(G256gat), .dout(n1798));
  jcb  g1735(.dina(n1780), .dinb(n1777), .dout(n1799));
  jcb  g1736(.dina(n1782), .dinb(n1776), .dout(n1800));
  jand g1737(.dina(n1800), .dinb(n1799), .dout(n1801));
  jxor g1738(.dina(n1801), .dinb(n1798), .dout(n1802));
  jnot g1739(.din(n1802), .dout(n1803));
  jxor g1740(.dina(n1803), .dinb(n1797), .dout(n1804));
  jxor g1741(.dina(n1804), .dinb(n1796), .dout(n1805));
  jxor g1742(.dina(n1805), .dinb(n1793), .dout(G6280gat));
  jand g1743(.dina(G528gat), .dinb(G256gat), .dout(n1807));
  jcb  g1744(.dina(n1801), .dinb(n1798), .dout(n1808));
  jcb  g1745(.dina(n1803), .dinb(n1797), .dout(n1809));
  jand g1746(.dina(n1809), .dinb(n1808), .dout(n1810));
  jcb  g1747(.dina(n1810), .dinb(n1807), .dout(n1811));
  jnot g1748(.din(n1796), .dout(n1812));
  jnot g1749(.din(n1804), .dout(n1813));
  jcb  g1750(.dina(n1813), .dinb(n1812), .dout(n1814));
  jnot g1751(.din(n1805), .dout(n1815));
  jcb  g1752(.dina(n1815), .dinb(n1793), .dout(n1816));
  jand g1753(.dina(n1816), .dinb(n1814), .dout(n1817));
  jxor g1754(.dina(n1810), .dinb(n1807), .dout(n1818));
  jnot g1755(.din(n1818), .dout(n1819));
  jcb  g1756(.dina(n1819), .dinb(n1817), .dout(n1820));
  jand g1757(.dina(n1820), .dinb(n1811), .dout(G6287gat));
  jxor g1758(.dina(n1818), .dinb(n1817), .dout(G6288gat));
endmodule


