// Benchmark "top" written by ABC on Wed May 27 23:37:08 2020

module gf_divisor ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , a16 ,
    a17 , a18 , a19 , a20 , a21 , a22 , a23 , a24 ,
    a25 , a26 , a27 , a28 , a29 , a30 , a31 , a32 ,
    a33 , a34 , a35 , a36 , a37 , a38 , a39 , a40 ,
    a41 , a42 , a43 , a44 , a45 , a46 , a47 , a48 ,
    a49 , a50 , a51 , a52 , a53 , a54 , a55 , a56 ,
    a57 , a58 , a59 , a60 , a61 , a62 , a63 , b0 ,
    b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 , b9 ,
    b10 , b11 , b12 , b13 , b14 , b15 , b16 , b17 ,
    b18 , b19 , b20 , b21 , b22 , b23 , b24 , b25 ,
    b26 , b27 , b28 , b29 , b30 , b31 , b32 , b33 ,
    b34 , b35 , b36 , b37 , b38 , b39 , b40 , b41 ,
    b42 , b43 , b44 , b45 , b46 , b47 , b48 , b49 ,
    b50 , b51 , b52 , b53 , b54 , b55 , b56 , b57 ,
    b58 , b59 , b60 , b61 , b62 , b63 ,
    quotient0 , quotient1 , quotient2 , quotient3 ,
    quotient4 , quotient5 , quotient6 , quotient7 ,
    quotient8 , quotient9 , quotient10 , quotient11 ,
    quotient12 , quotient13 , quotient14 , quotient15 ,
    quotient16 , quotient17 , quotient18 , quotient19 ,
    quotient20 , quotient21 , quotient22 , quotient23 ,
    quotient24 , quotient25 , quotient26 , quotient27 ,
    quotient28 , quotient29 , quotient30 , quotient31 ,
    quotient32 , quotient33 , quotient34 , quotient35 ,
    quotient36 , quotient37 , quotient38 , quotient39 ,
    quotient40 , quotient41 , quotient42 , quotient43 ,
    quotient44 , quotient45 , quotient46 , quotient47 ,
    quotient48 , quotient49 , quotient50 , quotient51 ,
    quotient52 , quotient53 , quotient54 , quotient55 ,
    quotient56 , quotient57 , quotient58 , quotient59 ,
    quotient60 , quotient61 , quotient62 , quotient63 ,
    remainder0 , remainder1 , remainder2 , remainder3 ,
    remainder4 , remainder5 , remainder6 , remainder7 ,
    remainder8 , remainder9 , remainder10 , remainder11 ,
    remainder12 , remainder13 , remainder14 , remainder15 ,
    remainder16 , remainder17 , remainder18 , remainder19 ,
    remainder20 , remainder21 , remainder22 , remainder23 ,
    remainder24 , remainder25 , remainder26 , remainder27 ,
    remainder28 , remainder29 , remainder30 , remainder31 ,
    remainder32 , remainder33 , remainder34 , remainder35 ,
    remainder36 , remainder37 , remainder38 , remainder39 ,
    remainder40 , remainder41 , remainder42 , remainder43 ,
    remainder44 , remainder45 , remainder46 , remainder47 ,
    remainder48 , remainder49 , remainder50 , remainder51 ,
    remainder52 , remainder53 , remainder54 , remainder55 ,
    remainder56 , remainder57 , remainder58 , remainder59 ,
    remainder60 , remainder61 , remainder62 , remainder63   );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    a16 , a17 , a18 , a19 , a20 , a21 , a22 , a23 ,
    a24 , a25 , a26 , a27 , a28 , a29 , a30 , a31 ,
    a32 , a33 , a34 , a35 , a36 , a37 , a38 , a39 ,
    a40 , a41 , a42 , a43 , a44 , a45 , a46 , a47 ,
    a48 , a49 , a50 , a51 , a52 , a53 , a54 , a55 ,
    a56 , a57 , a58 , a59 , a60 , a61 , a62 , a63 ,
    b0 , b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 ,
    b9 , b10 , b11 , b12 , b13 , b14 , b15 , b16 ,
    b17 , b18 , b19 , b20 , b21 , b22 , b23 , b24 ,
    b25 , b26 , b27 , b28 , b29 , b30 , b31 , b32 ,
    b33 , b34 , b35 , b36 , b37 , b38 , b39 , b40 ,
    b41 , b42 , b43 , b44 , b45 , b46 , b47 , b48 ,
    b49 , b50 , b51 , b52 , b53 , b54 , b55 , b56 ,
    b57 , b58 , b59 , b60 , b61 , b62 , b63 ;
  output quotient0 , quotient1 , quotient2 , quotient3 ,
    quotient4 , quotient5 , quotient6 , quotient7 ,
    quotient8 , quotient9 , quotient10 , quotient11 ,
    quotient12 , quotient13 , quotient14 , quotient15 ,
    quotient16 , quotient17 , quotient18 , quotient19 ,
    quotient20 , quotient21 , quotient22 , quotient23 ,
    quotient24 , quotient25 , quotient26 , quotient27 ,
    quotient28 , quotient29 , quotient30 , quotient31 ,
    quotient32 , quotient33 , quotient34 , quotient35 ,
    quotient36 , quotient37 , quotient38 , quotient39 ,
    quotient40 , quotient41 , quotient42 , quotient43 ,
    quotient44 , quotient45 , quotient46 , quotient47 ,
    quotient48 , quotient49 , quotient50 , quotient51 ,
    quotient52 , quotient53 , quotient54 , quotient55 ,
    quotient56 , quotient57 , quotient58 , quotient59 ,
    quotient60 , quotient61 , quotient62 , quotient63 ,
    remainder0 , remainder1 , remainder2 , remainder3 ,
    remainder4 , remainder5 , remainder6 , remainder7 ,
    remainder8 , remainder9 , remainder10 , remainder11 ,
    remainder12 , remainder13 , remainder14 , remainder15 ,
    remainder16 , remainder17 , remainder18 , remainder19 ,
    remainder20 , remainder21 , remainder22 , remainder23 ,
    remainder24 , remainder25 , remainder26 , remainder27 ,
    remainder28 , remainder29 , remainder30 , remainder31 ,
    remainder32 , remainder33 , remainder34 , remainder35 ,
    remainder36 , remainder37 , remainder38 , remainder39 ,
    remainder40 , remainder41 , remainder42 , remainder43 ,
    remainder44 , remainder45 , remainder46 , remainder47 ,
    remainder48 , remainder49 , remainder50 , remainder51 ,
    remainder52 , remainder53 , remainder54 , remainder55 ,
    remainder56 , remainder57 , remainder58 , remainder59 ,
    remainder60 , remainder61 , remainder62 , remainder63 ;
  wire n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n315,
    n316, n317, n318, n319, n320, n324, n325, n326, n327, n328, n329, n331,
    n332, n333, n334, n335, n336, n338, n339, n340, n341, n342, n347, n348,
    n349, n350, n351, n352, n354, n355, n356, n357, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n376, n377, n378, n379, n380, n381, n383, n384, n385, n386, n387, n388,
    n389, n390, n393, n394, n395, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n438, n444, n445, n446, n447, n448, n449,
    n455, n456, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n480, n481, n482, n483, n486, n487,
    n492, n493, n519, n520, n526, n527, n528, n529, n530, n531, n534, n572,
    n573, n574, n579, n580, n583, n589, n590, n591, n610, n648, n649, n650,
    n708, n714, n715, n716, n776, n777, n780, n786, n787, n788, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n914, n915, n916, n951, n952, n998, n999,
    n1002, n1008, n1009, n1010, n1095, n1096, n1104, n1105, n1106, n1207,
    n1208, n1209, n1253, n1254, n1314, n1317, n1323, n1324, n1325, n1429,
    n1430, n1431, n1439, n1440, n1441, n1569, n1570, n1571, n1700, n1706,
    n1707, n1708, n1841, n1842, n1845, n1851, n1852, n1853, n1910, n2001,
    n2002, n2003, n2156, n2162, n2163, n2164, n2315, n2316, n2319, n2325,
    n2326, n2327, n2503, n2504, n2505, n2680, n2681, n2684, n2689, n2690,
    n2691, n2873, n2880, n2881, n2882, n2951, n3076, n3077, n3078, n3157,
    n3158, n3302, n3305, n3310, n3311, n3412, n3469, n3470, n3592, n3593,
    n3600, n3601, n3602, n3678, n3822, n3823, n3824, n3911, n4047, n4053,
    n4054, n4055, n4145, n4277, n4278, n4281, n4287, n4288, n4289, n4540,
    n4541, n4542, n4789, n4795, n4796, n4797, n5042, n5043, n5046, n5052,
    n5053, n5054, n5326, n5327, n5328, n5629, n5630, n5633, n5638, n5639,
    n5777, n6018, n6025, n6026, n6027, n6320, n6321, n6322, n6436, n6437,
    n6653, n6656, n6661, n6662, n6812, n7074, n7075, n7076, n7077, n7084,
    n7085, n7086, n7401, n7402, n7403, n7526, n7527, n7723, n7729, n7730,
    n7731, n8054, n8057, n8063, n8064, n8065, n8446, n8447, n8617, n8923,
    n8924, n8925, n9062, n9273, n9274, n9275, n9424, n9648, n9649, n9650,
    n9795, n9796, n10014, n10015, n10018, n10024, n10025, n10026, n10176,
    n10406, n10407, n10408, n10797, n10798, n10799, n10953, n10954, n11186,
    n11189, n11195, n11196, n11197, n11605, n11606, n11607, n12015, n12016,
    n12017, n12427, n12430, n12436, n12437, n12438, n12863, n12864, n12865,
    n13022, n13025, n13026, n13300, n13301, n13302, n13732, n13735, n13741,
    n13742, n13743, n13910, n13916, n14203, n14204, n14205, n14661, n14662,
    n14663, n15122, n15125, n15131, n15132, n15133, n15612, n15613, n15614,
    n16095, n16096, n16097, n16289, n16585, n16586, n16587, n16769, n17077,
    n17078, n17079, n17269, n17514, n17515, n17523, n17542, n17552, n17559,
    n17570, n17580, n17590, n17591, n17592, n17597, n17602, n17603, n17608,
    n17615, n17625, n17626, n17627, n17632, n17639, n17650, n17660, n17661,
    n17662, n17667, n17672, n17673, n17678, n17683, n17684, n17689, n17696,
    n17707, n17718, n17729, n17740, n17751, n17762, n17772, n17779, n17789,
    n17790, n17801, n17802, n17813, n17814, n17822, n17823, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
    n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
    n17858, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
    n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
    n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
    n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
    n17899, n17900, n17905, n17906, n17907, n17910, n17911, n17912, n17915,
    n17916, n17917, n17920, n17921, n17922, n17928, n17929, n17930, n17931,
    n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17944,
    n17945, n17946, n17949, n17950, n17951, n17957, n17958, n17959, n17960,
    n17961, n17962, n17963, n17968, n17969, n17970, n17973, n17974, n17975,
    n17978, n17979, n17980, n17982, n17983, n17984, n17985, n17986, n17992,
    n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
    n18002, n18003, n18004, n18005, n18006, n18012, n18013, n18014, n18015,
    n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
    n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
    n18037, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
    n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
    n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18066, n18067,
    n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
    n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
    n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
    n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
    n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
    n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
    n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
    n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
    n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
    n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
    n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
    n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
    n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
    n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
    n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
    n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
    n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
    n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
    n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
    n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
    n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
    n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
    n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
    n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
    n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
    n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
    n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
    n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
    n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
    n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
    n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
    n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
    n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
    n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
    n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
    n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
    n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
    n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
    n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
    n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
    n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
    n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
    n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
    n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
    n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
    n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
    n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
    n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
    n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
    n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
    n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
    n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
    n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
    n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
    n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
    n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
    n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
    n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
    n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
    n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
    n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
    n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
    n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
    n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
    n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
    n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
    n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
    n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
    n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
    n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
    n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
    n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
    n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
    n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
    n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
    n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
    n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
    n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
    n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
    n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
    n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
    n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
    n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
    n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
    n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
    n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
    n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
    n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
    n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
    n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
    n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
    n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
    n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
    n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
    n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
    n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
    n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
    n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
    n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
    n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
    n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
    n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
    n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
    n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
    n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
    n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
    n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
    n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
    n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
    n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
    n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
    n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
    n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
    n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
    n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
    n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
    n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
    n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
    n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
    n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
    n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
    n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
    n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
    n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
    n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
    n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
    n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
    n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
    n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
    n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
    n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
    n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
    n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
    n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
    n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
    n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
    n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
    n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
    n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
    n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
    n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
    n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
    n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
    n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
    n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
    n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
    n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
    n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
    n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
    n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
    n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
    n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
    n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
    n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
    n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
    n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
    n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
    n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
    n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
    n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
    n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
    n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
    n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
    n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
    n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
    n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
    n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
    n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
    n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
    n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
    n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
    n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
    n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
    n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
    n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
    n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
    n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
    n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
    n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
    n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
    n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
    n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
    n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
    n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
    n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
    n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
    n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
    n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
    n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
    n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
    n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
    n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
    n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
    n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
    n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
    n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
    n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
    n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
    n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
    n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
    n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
    n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
    n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
    n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
    n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
    n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
    n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
    n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
    n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
    n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
    n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
    n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
    n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
    n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
    n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
    n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
    n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
    n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
    n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
    n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
    n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
    n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
    n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
    n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
    n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
    n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
    n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
    n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
    n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
    n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
    n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
    n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
    n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
    n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
    n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
    n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
    n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
    n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
    n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
    n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
    n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
    n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
    n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
    n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
    n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
    n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
    n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
    n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
    n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
    n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
    n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
    n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
    n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
    n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
    n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
    n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
    n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
    n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
    n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
    n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
    n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
    n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
    n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
    n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
    n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
    n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
    n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
    n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
    n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
    n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
    n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
    n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
    n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
    n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
    n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
    n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
    n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
    n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
    n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
    n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
    n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
    n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
    n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
    n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
    n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
    n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
    n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
    n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
    n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
    n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
    n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
    n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
    n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
    n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
    n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
    n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
    n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
    n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
    n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
    n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
    n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
    n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
    n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
    n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
    n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
    n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
    n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
    n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
    n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
    n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
    n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
    n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
    n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
    n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
    n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
    n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
    n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
    n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
    n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
    n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
    n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
    n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
    n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
    n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
    n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
    n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
    n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
    n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
    n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
    n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
    n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
    n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
    n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
    n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
    n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
    n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
    n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
    n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
    n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
    n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
    n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
    n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
    n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
    n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
    n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
    n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
    n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
    n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
    n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
    n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
    n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
    n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
    n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
    n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
    n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
    n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
    n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
    n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
    n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
    n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
    n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
    n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
    n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
    n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
    n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
    n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
    n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
    n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
    n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
    n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
    n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
    n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
    n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
    n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
    n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054,
    n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
    n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
    n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
    n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
    n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
    n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
    n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
    n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
    n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
    n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
    n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
    n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
    n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
    n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
    n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189,
    n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
    n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
    n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
    n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
    n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
    n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
    n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
    n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261,
    n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
    n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
    n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
    n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
    n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
    n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
    n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
    n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333,
    n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342,
    n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
    n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
    n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
    n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
    n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
    n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396,
    n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405,
    n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414,
    n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
    n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
    n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
    n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
    n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
    n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468,
    n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477,
    n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486,
    n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
    n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,
    n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
    n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
    n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
    n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
    n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549,
    n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558,
    n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
    n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
    n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
    n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
    n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
    n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612,
    n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621,
    n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630,
    n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
    n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,
    n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
    n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
    n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
    n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
    n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702,
    n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
    n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
    n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
    n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
    n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
    n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
    n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765,
    n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774,
    n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
    n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
    n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
    n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
    n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
    n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828,
    n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837,
    n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846,
    n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
    n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
    n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
    n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
    n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
    n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900,
    n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909,
    n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918,
    n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
    n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
    n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
    n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954,
    n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
    n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972,
    n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981,
    n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990,
    n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
    n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
    n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
    n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026,
    n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
    n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044,
    n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053,
    n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062,
    n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
    n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
    n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
    n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098,
    n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
    n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116,
    n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125,
    n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134,
    n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
    n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
    n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
    n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
    n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
    n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188,
    n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197,
    n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206,
    n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
    n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,
    n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
    n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
    n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
    n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260,
    n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269,
    n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278,
    n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
    n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
    n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
    n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
    n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
    n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332,
    n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341,
    n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350,
    n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
    n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
    n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
    n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
    n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
    n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404,
    n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413,
    n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422,
    n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
    n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,
    n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
    n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
    n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
    n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476,
    n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
    n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494,
    n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
    n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,
    n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
    n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
    n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
    n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548,
    n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557,
    n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566,
    n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
    n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,
    n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
    n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602,
    n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
    n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620,
    n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
    n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638,
    n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
    n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656,
    n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
    n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674,
    n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
    n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692,
    n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701,
    n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710,
    n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
    n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728,
    n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
    n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746,
    n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
    n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764,
    n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773,
    n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782,
    n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
    n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800,
    n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
    n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818,
    n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
    n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836,
    n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845,
    n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854,
    n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
    n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872,
    n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
    n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890,
    n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
    n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908,
    n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917,
    n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926,
    n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
    n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,
    n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
    n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
    n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
    n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980,
    n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
    n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998,
    n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
    n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
    n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
    n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034,
    n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
    n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
    n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
    n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070,
    n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
    n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
    n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
    n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
    n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
    n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124,
    n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
    n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
    n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
    n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
    n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
    n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178,
    n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
    n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196,
    n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
    n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
    n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
    n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
    n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
    n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
    n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268,
    n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277,
    n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286,
    n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
    n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
    n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
    n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
    n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
    n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340,
    n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349,
    n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358,
    n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
    n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,
    n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
    n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394,
    n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
    n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412,
    n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421,
    n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430,
    n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
    n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,
    n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
    n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
    n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
    n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484,
    n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493,
    n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502,
    n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
    n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,
    n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
    n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
    n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
    n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556,
    n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565,
    n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574,
    n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
    n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592,
    n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
    n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
    n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
    n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
    n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637,
    n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646,
    n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
    n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664,
    n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
    n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
    n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
    n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700,
    n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709,
    n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718,
    n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
    n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,
    n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
    n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
    n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
    n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772,
    n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781,
    n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790,
    n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799,
    n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808,
    n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
    n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
    n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
    n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
    n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853,
    n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862,
    n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871,
    n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880,
    n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
    n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
    n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
    n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916,
    n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925,
    n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934,
    n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943,
    n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952,
    n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
    n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
    n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
    n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988,
    n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997,
    n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006,
    n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
    n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024,
    n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
    n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
    n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
    n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060,
    n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069,
    n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078,
    n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087,
    n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
    n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
    n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
    n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
    n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132,
    n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141,
    n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150,
    n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
    n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
    n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
    n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
    n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
    n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204,
    n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213,
    n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222,
    n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231,
    n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
    n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
    n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
    n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
    n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276,
    n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285,
    n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294,
    n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303,
    n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
    n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
    n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
    n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
    n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348,
    n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357,
    n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366,
    n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375,
    n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
    n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
    n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
    n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
    n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420,
    n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429,
    n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438,
    n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
    n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
    n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
    n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
    n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
    n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
    n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501,
    n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510,
    n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
    n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
    n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
    n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564,
    n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573,
    n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582,
    n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591,
    n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
    n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
    n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
    n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
    n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636,
    n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654,
    n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663,
    n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
    n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
    n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
    n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
    n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708,
    n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717,
    n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726,
    n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735,
    n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,
    n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
    n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
    n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
    n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780,
    n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789,
    n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798,
    n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807,
    n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,
    n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
    n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
    n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
    n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852,
    n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861,
    n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870,
    n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879,
    n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,
    n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
    n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
    n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
    n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924,
    n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933,
    n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942,
    n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951,
    n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,
    n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
    n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
    n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
    n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996,
    n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014,
    n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,
    n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
    n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
    n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
    n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068,
    n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077,
    n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086,
    n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095,
    n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
    n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
    n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
    n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140,
    n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149,
    n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158,
    n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167,
    n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
    n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
    n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
    n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
    n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212,
    n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221,
    n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230,
    n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239,
    n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,
    n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
    n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
    n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284,
    n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293,
    n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302,
    n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311,
    n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,
    n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
    n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
    n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
    n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356,
    n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365,
    n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374,
    n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383,
    n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
    n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
    n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
    n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
    n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428,
    n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437,
    n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446,
    n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455,
    n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,
    n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
    n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
    n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
    n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500,
    n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518,
    n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
    n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536,
    n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
    n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
    n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572,
    n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590,
    n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,
    n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
    n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644,
    n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653,
    n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662,
    n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
    n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,
    n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
    n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
    n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
    n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
    n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734,
    n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,
    n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
    n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
    n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806,
    n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
    n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
    n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
    n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878,
    n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
    n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
    n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
    n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
    n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932,
    n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941,
    n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950,
    n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
    n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
    n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
    n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
    n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
    n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004,
    n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013,
    n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022,
    n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031,
    n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,
    n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
    n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
    n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
    n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076,
    n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085,
    n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094,
    n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103,
    n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,
    n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
    n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
    n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
    n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
    n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157,
    n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166,
    n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175,
    n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
    n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
    n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
    n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211,
    n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220,
    n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229,
    n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238,
    n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247,
    n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256,
    n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
    n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
    n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283,
    n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292,
    n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301,
    n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310,
    n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319,
    n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328,
    n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
    n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
    n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
    n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364,
    n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373,
    n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382,
    n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391,
    n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400,
    n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
    n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
    n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427,
    n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436,
    n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445,
    n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454,
    n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463,
    n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472,
    n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
    n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490,
    n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499,
    n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508,
    n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517,
    n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526,
    n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535,
    n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544,
    n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
    n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
    n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
    n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580,
    n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589,
    n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598,
    n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607,
    n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616,
    n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
    n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
    n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
    n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652,
    n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661,
    n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670,
    n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679,
    n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688,
    n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
    n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
    n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
    n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724,
    n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733,
    n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742,
    n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751,
    n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760,
    n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
    n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
    n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
    n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796,
    n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805,
    n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814,
    n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823,
    n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832,
    n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
    n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850,
    n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
    n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868,
    n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877,
    n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886,
    n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895,
    n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904,
    n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
    n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922,
    n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
    n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940,
    n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949,
    n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958,
    n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967,
    n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976,
    n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
    n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994,
    n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
    n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012,
    n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021,
    n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030,
    n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039,
    n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048,
    n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
    n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
    n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
    n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
    n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093,
    n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102,
    n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111,
    n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120,
    n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
    n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
    n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
    n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156,
    n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165,
    n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174,
    n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183,
    n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192,
    n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
    n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210,
    n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
    n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228,
    n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237,
    n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246,
    n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255,
    n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264,
    n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
    n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282,
    n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
    n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300,
    n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309,
    n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318,
    n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327,
    n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336,
    n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
    n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354,
    n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
    n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372,
    n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381,
    n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390,
    n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399,
    n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408,
    n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
    n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426,
    n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
    n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444,
    n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453,
    n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462,
    n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471,
    n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480,
    n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
    n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498,
    n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
    n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516,
    n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525,
    n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534,
    n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543,
    n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552,
    n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
    n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570,
    n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
    n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588,
    n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597,
    n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606,
    n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615,
    n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624,
    n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
    n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642,
    n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
    n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660,
    n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669,
    n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678,
    n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687,
    n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696,
    n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
    n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714,
    n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
    n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732,
    n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741,
    n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750,
    n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759,
    n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768,
    n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
    n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786,
    n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
    n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804,
    n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813,
    n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822,
    n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831,
    n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840,
    n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
    n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858,
    n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
    n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876,
    n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885,
    n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894,
    n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903,
    n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912,
    n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
    n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930,
    n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
    n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
    n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966,
    n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984,
    n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
    n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020,
    n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038,
    n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047,
    n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056,
    n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
    n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074,
    n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
    n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092,
    n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110,
    n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
    n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128,
    n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
    n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146,
    n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
    n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164,
    n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173,
    n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182,
    n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191,
    n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200,
    n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
    n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218,
    n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
    n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236,
    n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245,
    n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254,
    n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263,
    n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272,
    n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
    n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290,
    n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299,
    n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308,
    n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317,
    n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326,
    n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335,
    n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344,
    n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
    n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362,
    n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
    n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380,
    n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389,
    n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398,
    n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407,
    n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416,
    n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
    n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434,
    n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443,
    n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452,
    n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461,
    n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470,
    n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479,
    n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488,
    n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
    n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
    n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515,
    n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524,
    n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533,
    n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542,
    n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551,
    n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560,
    n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
    n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578,
    n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
    n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596,
    n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605,
    n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614,
    n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623,
    n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632,
    n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
    n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650,
    n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
    n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668,
    n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677,
    n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686,
    n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695,
    n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704,
    n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
    n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722,
    n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731,
    n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740,
    n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749,
    n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758,
    n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767,
    n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776,
    n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
    n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794,
    n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
    n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812,
    n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821,
    n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830,
    n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839,
    n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848,
    n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
    n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866,
    n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875,
    n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884,
    n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893,
    n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902,
    n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911,
    n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920,
    n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
    n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938,
    n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
    n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956,
    n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965,
    n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974,
    n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983,
    n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992,
    n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
    n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010,
    n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019,
    n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028,
    n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037,
    n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046,
    n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055,
    n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064,
    n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
    n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082,
    n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091,
    n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100,
    n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109,
    n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118,
    n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127,
    n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136,
    n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
    n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154,
    n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163,
    n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172,
    n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181,
    n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190,
    n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199,
    n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208,
    n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
    n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226,
    n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
    n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244,
    n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253,
    n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262,
    n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271,
    n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280,
    n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
    n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298,
    n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
    n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316,
    n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325,
    n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334,
    n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343,
    n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352,
    n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
    n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370,
    n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
    n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388,
    n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397,
    n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406,
    n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415,
    n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424,
    n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
    n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442,
    n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
    n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460,
    n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469,
    n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478,
    n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487,
    n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496,
    n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
    n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514,
    n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523,
    n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532,
    n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541,
    n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550,
    n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559,
    n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568,
    n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
    n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586,
    n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595,
    n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604,
    n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613,
    n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622,
    n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631,
    n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640,
    n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
    n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658,
    n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667,
    n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676,
    n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685,
    n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694,
    n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703,
    n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712,
    n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
    n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730,
    n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739,
    n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748,
    n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757,
    n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766,
    n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775,
    n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784,
    n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
    n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802,
    n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811,
    n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820,
    n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829,
    n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838,
    n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847,
    n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856,
    n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
    n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874,
    n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883,
    n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892,
    n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901,
    n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910,
    n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919,
    n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928,
    n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
    n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946,
    n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955,
    n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964,
    n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973,
    n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982,
    n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991,
    n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000,
    n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
    n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018,
    n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027,
    n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036,
    n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045,
    n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054,
    n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063,
    n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072,
    n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
    n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090,
    n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099,
    n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108,
    n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117,
    n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126,
    n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135,
    n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144,
    n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
    n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162,
    n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171,
    n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180,
    n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189,
    n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198,
    n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207,
    n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216,
    n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
    n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234,
    n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243,
    n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252,
    n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261,
    n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270,
    n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279,
    n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288,
    n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
    n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306,
    n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315,
    n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324,
    n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333,
    n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342,
    n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351,
    n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360,
    n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
    n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378,
    n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387,
    n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396,
    n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405,
    n31406, n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414,
    n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423,
    n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432,
    n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
    n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450,
    n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459,
    n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468,
    n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477,
    n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
    n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495,
    n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504,
    n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
    n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522,
    n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531,
    n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540,
    n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549,
    n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558,
    n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567,
    n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576,
    n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
    n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594,
    n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603,
    n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612,
    n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621,
    n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630,
    n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639,
    n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648,
    n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
    n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666,
    n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675,
    n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684,
    n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693,
    n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702,
    n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711,
    n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720,
    n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
    n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738,
    n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747,
    n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756,
    n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765,
    n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774,
    n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783,
    n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792,
    n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
    n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810,
    n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819,
    n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828,
    n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837,
    n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846,
    n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855,
    n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864,
    n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
    n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882,
    n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891,
    n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900,
    n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909,
    n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918,
    n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927,
    n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936,
    n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
    n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954,
    n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963,
    n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972,
    n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981,
    n31982, n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990,
    n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999,
    n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008,
    n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
    n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026,
    n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035,
    n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044,
    n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053,
    n32054, n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062,
    n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071,
    n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080,
    n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
    n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098,
    n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107,
    n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116,
    n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125,
    n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134,
    n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143,
    n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152,
    n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
    n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170,
    n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179,
    n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188,
    n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197,
    n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206,
    n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215,
    n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224,
    n32225, n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
    n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242,
    n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251,
    n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260,
    n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268, n32269,
    n32270, n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278,
    n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287,
    n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296,
    n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
    n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314,
    n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323,
    n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332,
    n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341,
    n32342, n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350,
    n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359,
    n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368,
    n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
    n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386,
    n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395,
    n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404,
    n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413,
    n32414, n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422,
    n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431,
    n32432, n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440,
    n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
    n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458,
    n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467,
    n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476,
    n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485,
    n32486, n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494,
    n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503,
    n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512,
    n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
    n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530,
    n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539,
    n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548,
    n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557,
    n32558, n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566,
    n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575,
    n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584,
    n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
    n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602,
    n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611,
    n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620,
    n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629,
    n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638,
    n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647,
    n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656,
    n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
    n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674,
    n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683,
    n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692,
    n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701,
    n32702, n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710,
    n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719,
    n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728,
    n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
    n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746,
    n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755,
    n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764,
    n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773,
    n32774, n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782,
    n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791,
    n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800,
    n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
    n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818,
    n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827,
    n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836,
    n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845,
    n32846, n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854,
    n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863,
    n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872,
    n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
    n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890,
    n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899,
    n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908,
    n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916, n32917,
    n32918, n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926,
    n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935,
    n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944,
    n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
    n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962,
    n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971,
    n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980,
    n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32989,
    n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998,
    n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007,
    n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016,
    n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
    n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034,
    n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043,
    n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052,
    n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061,
    n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070,
    n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079,
    n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088,
    n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
    n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106,
    n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115,
    n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124,
    n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133,
    n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142,
    n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151,
    n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160,
    n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
    n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178,
    n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187,
    n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196,
    n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205,
    n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214,
    n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223,
    n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232,
    n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
    n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250,
    n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259,
    n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268,
    n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277,
    n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
    n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295,
    n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304,
    n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
    n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322,
    n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331,
    n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340,
    n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349,
    n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
    n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367,
    n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376,
    n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
    n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394,
    n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403,
    n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412,
    n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421,
    n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430,
    n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439,
    n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448,
    n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
    n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466,
    n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475,
    n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484,
    n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493,
    n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502,
    n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511,
    n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520,
    n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
    n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538,
    n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547,
    n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556,
    n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565,
    n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574,
    n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583,
    n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592,
    n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
    n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610,
    n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619,
    n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628,
    n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637,
    n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646,
    n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655,
    n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664,
    n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
    n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682,
    n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691,
    n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700,
    n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709,
    n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
    n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727,
    n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736,
    n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
    n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754,
    n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763,
    n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772,
    n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781,
    n33782, n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
    n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799,
    n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808,
    n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
    n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826,
    n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
    n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844,
    n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853,
    n33854, n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
    n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871,
    n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880,
    n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
    n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898,
    n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907,
    n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916,
    n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925,
    n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934,
    n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943,
    n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952,
    n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
    n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970,
    n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979,
    n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988,
    n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997,
    n33998, n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006,
    n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015,
    n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024,
    n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
    n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042,
    n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051,
    n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060,
    n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069,
    n34070, n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
    n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087,
    n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096,
    n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
    n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114,
    n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123,
    n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132,
    n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141,
    n34142, n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
    n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159,
    n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168,
    n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
    n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186,
    n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195,
    n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204,
    n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213,
    n34214, n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222,
    n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231,
    n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240,
    n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
    n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258,
    n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267,
    n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276,
    n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285,
    n34286, n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294,
    n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303,
    n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312,
    n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
    n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330,
    n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339,
    n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348,
    n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357,
    n34358, n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366,
    n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375,
    n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384,
    n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
    n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402,
    n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411,
    n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420,
    n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429,
    n34430, n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438,
    n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447,
    n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456,
    n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
    n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474,
    n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483,
    n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492,
    n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501,
    n34502, n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510,
    n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519,
    n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528,
    n34529, n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
    n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546,
    n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555,
    n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564,
    n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573,
    n34574, n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582,
    n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591,
    n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600,
    n34601, n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
    n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618,
    n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627,
    n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636,
    n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644, n34645,
    n34646, n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654,
    n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663,
    n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672,
    n34673, n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
    n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690,
    n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699,
    n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708,
    n34709, n34710, n34711, n34712, n34713, n34714, n34715, n34716, n34717,
    n34718, n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726,
    n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735,
    n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744,
    n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
    n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762,
    n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771,
    n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780,
    n34781, n34782, n34783, n34784, n34785, n34786, n34787, n34788, n34789,
    n34790, n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798,
    n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807,
    n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816,
    n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
    n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834,
    n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843,
    n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852,
    n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860, n34861,
    n34862, n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870,
    n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879,
    n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888,
    n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
    n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906,
    n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915,
    n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924,
    n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932, n34933,
    n34934, n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942,
    n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951,
    n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960,
    n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
    n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978,
    n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987,
    n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996,
    n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004, n35005,
    n35006, n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014,
    n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023,
    n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032,
    n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
    n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050,
    n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059,
    n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068,
    n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076, n35077,
    n35078, n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086,
    n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095,
    n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104,
    n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
    n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122,
    n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131,
    n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140,
    n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148, n35149,
    n35150, n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158,
    n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167,
    n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176,
    n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
    n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194,
    n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203,
    n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212,
    n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220, n35221,
    n35222, n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230,
    n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239,
    n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248,
    n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
    n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266,
    n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275,
    n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284,
    n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292, n35293,
    n35294, n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302,
    n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311,
    n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320,
    n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
    n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338,
    n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347,
    n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356,
    n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364, n35365,
    n35366, n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374,
    n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383,
    n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392,
    n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
    n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410,
    n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419,
    n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428,
    n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436, n35437,
    n35438, n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446,
    n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455,
    n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464,
    n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
    n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482,
    n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491,
    n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500,
    n35501, n35502, n35503, n35504, n35505, n35506, n35507, n35508, n35509,
    n35510, n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518,
    n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527,
    n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536,
    n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
    n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554,
    n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563,
    n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572,
    n35573, n35574, n35575, n35576, n35577, n35578, n35579, n35580, n35581,
    n35582, n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590,
    n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599,
    n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608,
    n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
    n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626,
    n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635,
    n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644,
    n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652, n35653,
    n35654, n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662,
    n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671,
    n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680,
    n35681, n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
    n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698,
    n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707,
    n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716,
    n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724, n35725,
    n35726, n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734,
    n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743,
    n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752,
    n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
    n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770,
    n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779,
    n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788,
    n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796, n35797,
    n35798, n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806,
    n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815,
    n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824,
    n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
    n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842,
    n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851,
    n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860,
    n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868, n35869,
    n35870, n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878,
    n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887,
    n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896,
    n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
    n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914,
    n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923,
    n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932,
    n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941,
    n35942, n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950,
    n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959,
    n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968,
    n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
    n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986,
    n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995,
    n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004,
    n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012, n36013,
    n36014, n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022,
    n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031,
    n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040,
    n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
    n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058,
    n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067,
    n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076,
    n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084, n36085,
    n36086, n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094,
    n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103,
    n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112,
    n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
    n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130,
    n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139,
    n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148,
    n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156, n36157,
    n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166,
    n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175,
    n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184,
    n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
    n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202,
    n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211,
    n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220,
    n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229,
    n36230, n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238,
    n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247,
    n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256,
    n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
    n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274,
    n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283,
    n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291, n36292,
    n36293, n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301,
    n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310,
    n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319,
    n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328,
    n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
    n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346,
    n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355,
    n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364,
    n36365, n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373,
    n36374, n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382,
    n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391,
    n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400,
    n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
    n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418,
    n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427,
    n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436,
    n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445,
    n36446, n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454,
    n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463,
    n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472,
    n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
    n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490,
    n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499,
    n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508,
    n36509, n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517,
    n36518, n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526,
    n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535,
    n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544,
    n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
    n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562,
    n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571,
    n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580,
    n36581, n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589,
    n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598,
    n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607,
    n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616,
    n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
    n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634,
    n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643,
    n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652,
    n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661,
    n36662, n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670,
    n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679,
    n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688,
    n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
    n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706,
    n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715,
    n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724,
    n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733,
    n36734, n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742,
    n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751,
    n36752, n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760,
    n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
    n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778,
    n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787,
    n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796,
    n36797, n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805,
    n36806, n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814,
    n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823,
    n36824, n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832,
    n36833, n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
    n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850,
    n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859,
    n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868,
    n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877,
    n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886,
    n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895,
    n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904,
    n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
    n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922,
    n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931,
    n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940,
    n36941, n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949,
    n36950, n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958,
    n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967,
    n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976,
    n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
    n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994,
    n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003,
    n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012,
    n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021,
    n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030,
    n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039,
    n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048,
    n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
    n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066,
    n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075,
    n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084,
    n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093,
    n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102,
    n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111,
    n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120,
    n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
    n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138,
    n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147,
    n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156,
    n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165,
    n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174,
    n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183,
    n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192,
    n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
    n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210,
    n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219,
    n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228,
    n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237,
    n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246,
    n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255,
    n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264,
    n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
    n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282,
    n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291,
    n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300,
    n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309,
    n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318,
    n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327,
    n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336,
    n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
    n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354,
    n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363,
    n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372,
    n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381,
    n37382, n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390,
    n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399,
    n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408,
    n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
    n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426,
    n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435,
    n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444,
    n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453,
    n37454, n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462,
    n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471,
    n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480,
    n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
    n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498,
    n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507,
    n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516,
    n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525,
    n37526, n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534,
    n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543,
    n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552,
    n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
    n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570,
    n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579,
    n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588,
    n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597,
    n37598, n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606,
    n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615,
    n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624,
    n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
    n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642,
    n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651,
    n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660,
    n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669,
    n37670, n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678,
    n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687,
    n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696,
    n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
    n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714,
    n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723,
    n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732,
    n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741,
    n37742, n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750,
    n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759,
    n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768,
    n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
    n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786,
    n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795,
    n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804,
    n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813,
    n37814, n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822,
    n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831,
    n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840,
    n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
    n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858,
    n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867,
    n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876,
    n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885,
    n37886, n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894,
    n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903,
    n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912,
    n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
    n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930,
    n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939,
    n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948,
    n37949, n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957,
    n37958, n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966,
    n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975,
    n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984,
    n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
    n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002,
    n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011,
    n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020,
    n38021, n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029,
    n38030, n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038,
    n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047,
    n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056,
    n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
    n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074,
    n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083,
    n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092,
    n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101,
    n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110,
    n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119,
    n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128,
    n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
    n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146,
    n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155,
    n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164,
    n38165, n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173,
    n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182,
    n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191,
    n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200,
    n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
    n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218,
    n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227,
    n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236,
    n38237, n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245,
    n38246, n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254,
    n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263,
    n38264, n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272,
    n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
    n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290,
    n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299,
    n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307, n38308,
    n38309, n38310, n38311, n38312, n38313, n38314, n38315, n38316, n38317,
    n38318, n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326,
    n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335,
    n38336, n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344,
    n38345, n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
    n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362,
    n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371,
    n38372, n38373, n38374, n38375, n38376, n38377, n38378, n38379, n38380,
    n38381, n38382, n38383, n38384, n38385, n38386, n38387, n38388, n38389,
    n38390, n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398,
    n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406, n38407,
    n38408, n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416,
    n38417, n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
    n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434,
    n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443,
    n38444, n38445, n38446, n38447, n38448, n38449, n38450, n38451, n38452,
    n38453, n38454, n38455, n38456, n38457, n38458, n38459, n38460, n38461,
    n38462, n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470,
    n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478, n38479,
    n38480, n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488,
    n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
    n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506,
    n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515,
    n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523, n38524,
    n38525, n38526, n38527, n38528, n38529, n38530, n38531, n38532, n38533,
    n38534, n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542,
    n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550, n38551,
    n38552, n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560,
    n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
    n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578,
    n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587,
    n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595, n38596,
    n38597, n38598, n38599, n38600, n38601, n38602, n38603, n38604, n38605,
    n38606, n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614,
    n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622, n38623,
    n38624, n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632,
    n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
    n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650,
    n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659,
    n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667, n38668,
    n38669, n38670, n38671, n38672, n38673, n38674, n38675, n38676, n38677,
    n38678, n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686,
    n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695,
    n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704,
    n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
    n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722,
    n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731,
    n38732, n38733, n38734, n38735, n38736, n38737, n38738, n38739, n38740,
    n38741, n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749,
    n38750, n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758,
    n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767,
    n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776,
    n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
    n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794,
    n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803,
    n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811, n38812,
    n38813, n38814, n38815, n38816, n38817, n38818, n38819, n38820, n38821,
    n38822, n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830,
    n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839,
    n38840, n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848,
    n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
    n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866,
    n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875,
    n38876, n38877, n38878, n38879, n38880, n38881, n38882, n38883, n38884,
    n38885, n38886, n38887, n38888, n38889, n38890, n38891, n38892, n38893,
    n38894, n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902,
    n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911,
    n38912, n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920,
    n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
    n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938,
    n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947,
    n38948, n38949, n38950, n38952, n38953, n38954, n38955, n38956, n38957,
    n38958, n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966,
    n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975,
    n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984,
    n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
    n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002,
    n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011,
    n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019, n39020,
    n39021, n39022, n39023, n39024, n39025, n39026, n39027, n39028, n39029,
    n39030, n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038,
    n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047,
    n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056,
    n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
    n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074,
    n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083,
    n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091, n39092,
    n39093, n39094, n39095, n39096, n39097, n39098, n39099, n39100, n39101,
    n39102, n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110,
    n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119,
    n39120, n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128,
    n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
    n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
    n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155,
    n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163, n39164,
    n39165, n39166, n39167, n39168, n39169, n39170, n39171, n39172, n39173,
    n39174, n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182,
    n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191,
    n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200,
    n39201, n39202, n39203, n39204, n39205, n39207, n39208, n39209, n39210,
    n39212, n39213, n39214, n39216, n39217, n39218, n39220, n39221, n39222,
    n39224, n39225, n39226, n39228, n39229, n39230, n39232, n39233, n39234,
    n39236, n39237, n39238, n39240, n39241, n39242, n39244, n39245, n39246,
    n39248, n39249, n39250, n39252, n39253, n39254, n39256, n39257, n39258,
    n39260, n39261, n39262, n39264, n39265, n39266, n39268, n39269, n39270,
    n39272, n39273, n39274, n39276, n39277, n39278, n39280, n39281, n39282,
    n39284, n39285, n39286, n39288, n39289, n39290, n39292, n39293, n39294,
    n39296, n39297, n39298, n39300, n39301, n39302, n39304, n39305, n39306,
    n39308, n39309, n39310, n39312, n39313, n39314, n39316, n39317, n39318,
    n39320, n39321, n39322, n39324, n39325, n39326, n39328, n39329, n39330,
    n39332, n39333, n39334, n39336, n39337, n39338, n39340, n39341, n39342,
    n39344, n39345, n39346, n39348, n39349, n39350, n39352, n39353, n39354,
    n39356, n39357, n39358, n39360, n39361, n39362, n39364, n39365, n39366,
    n39368, n39369, n39370, n39372, n39373, n39374, n39376, n39377, n39378,
    n39380, n39381, n39382, n39384, n39385, n39386, n39388, n39389, n39390,
    n39392, n39393, n39394, n39396, n39397, n39398, n39400, n39401, n39402,
    n39404, n39405, n39406, n39408, n39409, n39410, n39412, n39413, n39414,
    n39416, n39417, n39418, n39420, n39421, n39422, n39424, n39425, n39426,
    n39428, n39429, n39430, n39432, n39433, n39434, n39436, n39437, n39438,
    n39440, n39441, n39442, n39444, n39445, n39446, n39448, n39449, n39450,
    n39452, n39453;
  jnot g00000(.din(b63 ), .dout(n256));
  jnot g00001(.din(b61 ), .dout(n257));
  jnot g00002(.din(a62 ), .dout(n258));
  jnot g00003(.din(b1 ), .dout(n259));
  jand g00004(.dina(b0 ), .dinb(n258), .dout(n260));
  jnot g00005(.din(n260), .dout(n261));
  jand g00006(.dina(n261), .dinb(n259), .dout(n262));
  jnot g00007(.din(n262), .dout(n263));
  jnot g00008(.din(b3 ), .dout(n264));
  jnot g00009(.din(b7 ), .dout(n265));
  jnot g00010(.din(b18 ), .dout(n266));
  jnot g00011(.din(b19 ), .dout(n267));
  jnot g00012(.din(b23 ), .dout(n268));
  jnot g00013(.din(b25 ), .dout(n269));
  jnot g00014(.din(b26 ), .dout(n270));
  jnot g00015(.din(b27 ), .dout(n271));
  jand g00016(.dina(n271), .dinb(n270), .dout(n272));
  jand g00017(.dina(n272), .dinb(n269), .dout(n273));
  jnot g00018(.din(b24 ), .dout(n274));
  jnot g00019(.din(b31 ), .dout(n275));
  jnot g00020(.din(b35 ), .dout(n276));
  jnot g00021(.din(b39 ), .dout(n277));
  jnot g00022(.din(b40 ), .dout(n278));
  jnot g00023(.din(b41 ), .dout(n279));
  jnot g00024(.din(b42 ), .dout(n280));
  jand g00025(.dina(n280), .dinb(n279), .dout(n281));
  jand g00026(.dina(n281), .dinb(n278), .dout(n282));
  jnot g00027(.din(b43 ), .dout(n283));
  jnot g00028(.din(b47 ), .dout(n284));
  jnot g00029(.din(b48 ), .dout(n285));
  jnot g00030(.din(b49 ), .dout(n286));
  jnot g00031(.din(b50 ), .dout(n287));
  jnot g00032(.din(b51 ), .dout(n288));
  jnot g00033(.din(b52 ), .dout(n289));
  jnot g00034(.din(b53 ), .dout(n290));
  jnot g00035(.din(b54 ), .dout(n291));
  jnot g00036(.din(b55 ), .dout(n292));
  jnot g00037(.din(b56 ), .dout(n293));
  jnot g00038(.din(b57 ), .dout(n294));
  jnot g00039(.din(b58 ), .dout(n295));
  jnot g00040(.din(b59 ), .dout(n296));
  jnot g00041(.din(b60 ), .dout(n297));
  jnot g00042(.din(b62 ), .dout(n298));
  jand g00043(.dina(n256), .dinb(n298), .dout(n299));
  jand g00044(.dina(n299), .dinb(n257), .dout(n300));
  jand g00045(.dina(n300), .dinb(n297), .dout(n301));
  jand g00046(.dina(n301), .dinb(n296), .dout(n302));
  jand g00047(.dina(n302), .dinb(n295), .dout(n303));
  jand g00048(.dina(n303), .dinb(n294), .dout(n304));
  jand g00049(.dina(n304), .dinb(n293), .dout(n305));
  jand g00050(.dina(n305), .dinb(n292), .dout(n306));
  jand g00051(.dina(n306), .dinb(n291), .dout(n307));
  jand g00052(.dina(n307), .dinb(n290), .dout(n308));
  jand g00053(.dina(n308), .dinb(n289), .dout(n309));
  jand g00054(.dina(n309), .dinb(n288), .dout(n310));
  jand g00055(.dina(n310), .dinb(n287), .dout(n311));
  jand g00056(.dina(n311), .dinb(n286), .dout(n312));
  jand g00057(.dina(n312), .dinb(n285), .dout(n313));
  jnot g00058(.din(b44 ), .dout(n315));
  jnot g00059(.din(b45 ), .dout(n316));
  jnot g00060(.din(b46 ), .dout(n317));
  jand g00061(.dina(n317), .dinb(n316), .dout(n318));
  jand g00062(.dina(n318), .dinb(n315), .dout(n319));
  jand g00063(.dina(n319), .dinb(n403), .dout(n320));
  jnot g00064(.din(b36 ), .dout(n324));
  jnot g00065(.din(b37 ), .dout(n325));
  jnot g00066(.din(b38 ), .dout(n326));
  jand g00067(.dina(n326), .dinb(n325), .dout(n327));
  jand g00068(.dina(n327), .dinb(n324), .dout(n328));
  jand g00069(.dina(n328), .dinb(n407), .dout(n329));
  jnot g00070(.din(b32 ), .dout(n331));
  jnot g00071(.din(b33 ), .dout(n332));
  jnot g00072(.din(b34 ), .dout(n333));
  jand g00073(.dina(n333), .dinb(n332), .dout(n334));
  jand g00074(.dina(n334), .dinb(n331), .dout(n335));
  jand g00075(.dina(n335), .dinb(n410), .dout(n336));
  jnot g00076(.din(b28 ), .dout(n338));
  jnot g00077(.din(b29 ), .dout(n339));
  jnot g00078(.din(b30 ), .dout(n340));
  jand g00079(.dina(n340), .dinb(n339), .dout(n341));
  jand g00080(.dina(n341), .dinb(n338), .dout(n342));
  jnot g00081(.din(b20 ), .dout(n347));
  jnot g00082(.din(b21 ), .dout(n348));
  jnot g00083(.din(b22 ), .dout(n349));
  jand g00084(.dina(n349), .dinb(n348), .dout(n350));
  jand g00085(.dina(n350), .dinb(n347), .dout(n351));
  jand g00086(.dina(n351), .dinb(n417), .dout(n352));
  jand g00087(.dina(n1910), .dinb(n266), .dout(n354));
  jnot g00088(.din(b16 ), .dout(n355));
  jnot g00089(.din(b17 ), .dout(n356));
  jand g00090(.dina(n356), .dinb(n355), .dout(n357));
  jnot g00091(.din(b11 ), .dout(n359));
  jnot g00092(.din(b13 ), .dout(n360));
  jnot g00093(.din(b14 ), .dout(n361));
  jand g00094(.dina(n361), .dinb(n360), .dout(n362));
  jnot g00095(.din(b12 ), .dout(n363));
  jnot g00096(.din(b15 ), .dout(n364));
  jand g00097(.dina(n364), .dinb(n363), .dout(n365));
  jand g00098(.dina(n365), .dinb(n362), .dout(n366));
  jnot g00099(.din(b8 ), .dout(n367));
  jnot g00100(.din(b9 ), .dout(n368));
  jnot g00101(.din(b10 ), .dout(n369));
  jand g00102(.dina(n369), .dinb(n368), .dout(n370));
  jand g00103(.dina(n370), .dinb(n367), .dout(n371));
  jand g00104(.dina(n371), .dinb(n366), .dout(n372));
  jand g00105(.dina(n372), .dinb(n359), .dout(n373));
  jand g00106(.dina(n373), .dinb(n1429), .dout(n374));
  jnot g00107(.din(b4 ), .dout(n376));
  jnot g00108(.din(b5 ), .dout(n377));
  jnot g00109(.din(b6 ), .dout(n378));
  jand g00110(.dina(n378), .dinb(n377), .dout(n379));
  jand g00111(.dina(n379), .dinb(n376), .dout(n380));
  jand g00112(.dina(n380), .dinb(n430), .dout(n381));
  jand g00113(.dina(n486), .dinb(b0 ), .dout(n383));
  jnot g00114(.din(a63 ), .dout(n384));
  jand g00115(.dina(b0 ), .dinb(n384), .dout(n385));
  jnot g00116(.din(b2 ), .dout(n386));
  jand g00117(.dina(n386), .dinb(n259), .dout(n387));
  jnot g00118(.din(n387), .dout(n388));
  jor  g00119(.dina(n388), .dinb(n385), .dout(n389));
  jnot g00120(.din(n389), .dout(n390));
  jand g00121(.dina(n260), .dinb(b1 ), .dout(n393));
  jnot g00122(.din(n393), .dout(n394));
  jand g00123(.dina(n394), .dinb(a63 ), .dout(n395));
  jand g00124(.dina(n367), .dinb(n265), .dout(n400));
  jand g00125(.dina(n286), .dinb(n284), .dout(n401));
  jand g00126(.dina(n401), .dinb(n285), .dout(n402));
  jand g00127(.dina(n402), .dinb(n311), .dout(n403));
  jand g00128(.dina(n403), .dinb(n283), .dout(n404));
  jand g00129(.dina(n404), .dinb(n319), .dout(n405));
  jand g00130(.dina(n405), .dinb(n282), .dout(n406));
  jand g00131(.dina(n406), .dinb(n277), .dout(n407));
  jand g00132(.dina(n407), .dinb(n327), .dout(n408));
  jand g00133(.dina(n324), .dinb(n276), .dout(n409));
  jand g00134(.dina(n409), .dinb(n408), .dout(n410));
  jand g00135(.dina(n410), .dinb(n334), .dout(n411));
  jand g00136(.dina(n331), .dinb(n275), .dout(n412));
  jand g00137(.dina(n412), .dinb(n411), .dout(n413));
  jand g00138(.dina(n413), .dinb(n342), .dout(n414));
  jand g00139(.dina(n414), .dinb(n273), .dout(n415));
  jand g00140(.dina(n415), .dinb(n274), .dout(n416));
  jand g00141(.dina(n416), .dinb(n268), .dout(n417));
  jand g00142(.dina(n417), .dinb(n350), .dout(n418));
  jand g00143(.dina(n347), .dinb(n267), .dout(n419));
  jand g00144(.dina(n266), .dinb(n356), .dout(n420));
  jand g00145(.dina(n420), .dinb(n419), .dout(n421));
  jand g00146(.dina(n421), .dinb(n418), .dout(n422));
  jand g00147(.dina(n355), .dinb(n364), .dout(n423));
  jand g00148(.dina(n423), .dinb(n422), .dout(n424));
  jand g00149(.dina(n424), .dinb(n362), .dout(n425));
  jand g00150(.dina(n359), .dinb(n369), .dout(n426));
  jand g00151(.dina(n363), .dinb(n368), .dout(n427));
  jand g00152(.dina(n427), .dinb(n426), .dout(n428));
  jand g00153(.dina(n428), .dinb(n425), .dout(n429));
  jand g00154(.dina(n429), .dinb(n400), .dout(n430));
  jand g00155(.dina(n430), .dinb(n379), .dout(n431));
  jand g00156(.dina(n376), .dinb(b0 ), .dout(n432));
  jand g00157(.dina(n432), .dinb(n431), .dout(n433));
  jand g00158(.dina(n433), .dinb(n264), .dout(n434));
  jand g00159(.dina(n434), .dinb(n386), .dout(n435));
  jand g00160(.dina(n486), .dinb(n386), .dout(n438));
  jnot g00161(.din(a61 ), .dout(n444));
  jand g00162(.dina(b0 ), .dinb(n444), .dout(n445));
  jnot g00163(.din(n445), .dout(n446));
  jand g00164(.dina(n446), .dinb(n259), .dout(n447));
  jand g00165(.dina(n445), .dinb(b1 ), .dout(n448));
  jnot g00166(.din(n448), .dout(n449));
  jand g00167(.dina(n438), .dinb(n263), .dout(n455));
  jand g00168(.dina(n455), .dinb(n394), .dout(n456));
  jnot g00169(.din(n422), .dout(n462));
  jand g00170(.dina(n376), .dinb(n264), .dout(n463));
  jnot g00171(.din(n463), .dout(n464));
  jnot g00172(.din(n362), .dout(n465));
  jnot g00173(.din(n423), .dout(n466));
  jor  g00174(.dina(n466), .dinb(n465), .dout(n467));
  jnot g00175(.din(n379), .dout(n468));
  jnot g00176(.din(n400), .dout(n469));
  jor  g00177(.dina(n469), .dinb(n468), .dout(n470));
  jor  g00178(.dina(n470), .dinb(n448), .dout(n471));
  jnot g00179(.din(n428), .dout(n472));
  jor  g00180(.dina(n447), .dinb(n472), .dout(n473));
  jor  g00181(.dina(n473), .dinb(n471), .dout(n474));
  jor  g00182(.dina(n474), .dinb(n467), .dout(n475));
  jor  g00183(.dina(n475), .dinb(n464), .dout(n476));
  jor  g00184(.dina(n476), .dinb(n462), .dout(n477));
  jnot g00185(.din(a60 ), .dout(n480));
  jand g00186(.dina(b0 ), .dinb(n480), .dout(n481));
  jnot g00187(.din(n481), .dout(n482));
  jand g00188(.dina(n482), .dinb(n259), .dout(n483));
  jand g00189(.dina(n463), .dinb(n431), .dout(n486));
  jand g00190(.dina(n486), .dinb(n445), .dout(n487));
  jand g00191(.dina(n481), .dinb(b1 ), .dout(n492));
  jnot g00192(.din(n492), .dout(n493));
  jand g00193(.dina(n486), .dinb(n18070), .dout(quotient61 ));
  jand g00194(.dina(n18087), .dinb(n381), .dout(quotient60 ));
  jxor g00195(.dina(n481), .dinb(b1 ), .dout(n519));
  jand g00196(.dina(n519), .dinb(n381), .dout(n520));
  jnot g00197(.din(a59 ), .dout(n526));
  jand g00198(.dina(b0 ), .dinb(n526), .dout(n527));
  jnot g00199(.din(n527), .dout(n528));
  jand g00200(.dina(n528), .dinb(n259), .dout(n529));
  jand g00201(.dina(n527), .dinb(b1 ), .dout(n530));
  jnot g00202(.din(n530), .dout(n531));
  jand g00203(.dina(n481), .dinb(n381), .dout(n534));
  jand g00204(.dina(n18177), .dinb(n431), .dout(quotient59 ));
  jnot g00205(.din(n431), .dout(n572));
  jor  g00206(.dina(n529), .dinb(n572), .dout(n573));
  jor  g00207(.dina(n573), .dinb(n530), .dout(n574));
  jand g00208(.dina(n430), .dinb(b0 ), .dout(n579));
  jand g00209(.dina(n579), .dinb(n379), .dout(n580));
  jand g00210(.dina(n527), .dinb(n431), .dout(n583));
  jnot g00211(.din(a58 ), .dout(n589));
  jand g00212(.dina(b0 ), .dinb(n589), .dout(n590));
  jnot g00213(.din(n590), .dout(n591));
  jand g00214(.dina(n430), .dinb(n378), .dout(n610));
  jor  g00215(.dina(n18161), .dinb(n18195), .dout(quotient58 ));
  jnot g00216(.din(a57 ), .dout(n648));
  jand g00217(.dina(b0 ), .dinb(n648), .dout(n649));
  jnot g00218(.din(n649), .dout(n650));
  jand g00219(.dina(n18251), .dinb(n430), .dout(quotient57 ));
  jand g00220(.dina(n649), .dinb(n430), .dout(n708));
  jnot g00221(.din(a56 ), .dout(n714));
  jand g00222(.dina(b0 ), .dinb(n714), .dout(n715));
  jnot g00223(.din(n715), .dout(n716));
  jand g00224(.dina(n18342), .dinb(n374), .dout(quotient56 ));
  jand g00225(.dina(n429), .dinb(b0 ), .dout(n776));
  jand g00226(.dina(n776), .dinb(n367), .dout(n777));
  jand g00227(.dina(n715), .dinb(n374), .dout(n780));
  jnot g00228(.din(a55 ), .dout(n786));
  jand g00229(.dina(b0 ), .dinb(n786), .dout(n787));
  jnot g00230(.din(n787), .dout(n788));
  jnot g00231(.din(n18479), .dout(quotient55 ));
  jnot g00232(.din(n273), .dout(n828));
  jnot g00233(.din(n282), .dout(n829));
  jor  g00234(.dina(b63 ), .dinb(b62 ), .dout(n830));
  jor  g00235(.dina(n830), .dinb(b61 ), .dout(n831));
  jor  g00236(.dina(n831), .dinb(b60 ), .dout(n832));
  jor  g00237(.dina(n832), .dinb(b59 ), .dout(n833));
  jor  g00238(.dina(n833), .dinb(b58 ), .dout(n834));
  jor  g00239(.dina(n834), .dinb(b57 ), .dout(n835));
  jor  g00240(.dina(n835), .dinb(b56 ), .dout(n836));
  jor  g00241(.dina(n836), .dinb(b55 ), .dout(n837));
  jor  g00242(.dina(n837), .dinb(b54 ), .dout(n838));
  jor  g00243(.dina(n838), .dinb(b53 ), .dout(n839));
  jor  g00244(.dina(n839), .dinb(b52 ), .dout(n840));
  jor  g00245(.dina(n840), .dinb(b51 ), .dout(n841));
  jor  g00246(.dina(n841), .dinb(b50 ), .dout(n842));
  jor  g00247(.dina(n842), .dinb(b49 ), .dout(n843));
  jor  g00248(.dina(n843), .dinb(b48 ), .dout(n844));
  jor  g00249(.dina(n844), .dinb(b47 ), .dout(n845));
  jnot g00250(.din(n319), .dout(n846));
  jor  g00251(.dina(n846), .dinb(n845), .dout(n847));
  jor  g00252(.dina(n847), .dinb(b43 ), .dout(n848));
  jor  g00253(.dina(n848), .dinb(n829), .dout(n849));
  jor  g00254(.dina(n849), .dinb(b39 ), .dout(n850));
  jnot g00255(.din(n328), .dout(n851));
  jor  g00256(.dina(n851), .dinb(n850), .dout(n852));
  jor  g00257(.dina(n852), .dinb(b35 ), .dout(n853));
  jnot g00258(.din(n335), .dout(n854));
  jor  g00259(.dina(n854), .dinb(n853), .dout(n855));
  jor  g00260(.dina(n855), .dinb(b31 ), .dout(n856));
  jnot g00261(.din(n342), .dout(n857));
  jor  g00262(.dina(n857), .dinb(n856), .dout(n858));
  jor  g00263(.dina(n858), .dinb(b24 ), .dout(n859));
  jor  g00264(.dina(n859), .dinb(n828), .dout(n860));
  jor  g00265(.dina(n860), .dinb(b23 ), .dout(n861));
  jnot g00266(.din(n351), .dout(n862));
  jor  g00267(.dina(n862), .dinb(n861), .dout(n863));
  jor  g00268(.dina(n863), .dinb(b19 ), .dout(n864));
  jor  g00269(.dina(n864), .dinb(b18 ), .dout(n865));
  jnot g00270(.din(n357), .dout(n866));
  jor  g00271(.dina(n866), .dinb(n865), .dout(n867));
  jnot g00272(.din(n373), .dout(n868));
  jor  g00273(.dina(n868), .dinb(n867), .dout(n869));
  jnot g00274(.din(a54 ), .dout(n914));
  jand g00275(.dina(b0 ), .dinb(n914), .dout(n915));
  jnot g00276(.din(n915), .dout(n916));
  jand g00277(.dina(n18555), .dinb(n998), .dout(quotient54 ));
  jand g00278(.dina(n425), .dinb(n363), .dout(n951));
  jand g00279(.dina(n951), .dinb(n359), .dout(n952));
  jand g00280(.dina(n951), .dinb(n426), .dout(n998));
  jand g00281(.dina(n998), .dinb(b0 ), .dout(n999));
  jand g00282(.dina(n915), .dinb(n998), .dout(n1002));
  jnot g00283(.din(a53 ), .dout(n1008));
  jand g00284(.dina(b0 ), .dinb(n1008), .dout(n1009));
  jnot g00285(.din(n1009), .dout(n1010));
  jand g00286(.dina(n18681), .dinb(n952), .dout(quotient53 ));
  jand g00287(.dina(n951), .dinb(b0 ), .dout(n1095));
  jand g00288(.dina(n1095), .dinb(n359), .dout(n1096));
  jnot g00289(.din(a52 ), .dout(n1104));
  jand g00290(.dina(b0 ), .dinb(n1104), .dout(n1105));
  jnot g00291(.din(n1105), .dout(n1106));
  jnot g00292(.din(n18819), .dout(quotient52 ));
  jnot g00293(.din(a51 ), .dout(n1207));
  jand g00294(.dina(b0 ), .dinb(n1207), .dout(n1208));
  jnot g00295(.din(n1208), .dout(n1209));
  jand g00296(.dina(n18915), .dinb(n425), .dout(quotient51 ));
  jand g00297(.dina(n364), .dinb(n361), .dout(n1253));
  jand g00298(.dina(n1253), .dinb(n1429), .dout(n1254));
  jand g00299(.dina(n425), .dinb(b0 ), .dout(n1314));
  jand g00300(.dina(n1208), .dinb(n425), .dout(n1317));
  jnot g00301(.din(a50 ), .dout(n1323));
  jand g00302(.dina(b0 ), .dinb(n1323), .dout(n1324));
  jnot g00303(.din(n1324), .dout(n1325));
  jand g00304(.dina(n19077), .dinb(n1254), .dout(quotient50 ));
  jand g00305(.dina(n422), .dinb(n355), .dout(n1429));
  jand g00306(.dina(n1429), .dinb(b0 ), .dout(n1430));
  jand g00307(.dina(n1430), .dinb(n1253), .dout(n1431));
  jnot g00308(.din(a49 ), .dout(n1439));
  jand g00309(.dina(b0 ), .dinb(n1439), .dout(n1440));
  jnot g00310(.din(n1440), .dout(n1441));
  jor  g00311(.dina(n19248), .dinb(n19247), .dout(quotient49 ));
  jnot g00312(.din(a48 ), .dout(n1569));
  jand g00313(.dina(b0 ), .dinb(n1569), .dout(n1570));
  jnot g00314(.din(n1570), .dout(n1571));
  jand g00315(.dina(n19373), .dinb(n1429), .dout(quotient48 ));
  jand g00316(.dina(n1570), .dinb(n1429), .dout(n1700));
  jnot g00317(.din(a47 ), .dout(n1706));
  jand g00318(.dina(b0 ), .dinb(n1706), .dout(n1707));
  jnot g00319(.din(n1707), .dout(n1708));
  jand g00320(.dina(n19572), .dinb(n422), .dout(quotient47 ));
  jand g00321(.dina(n1910), .dinb(b0 ), .dout(n1841));
  jand g00322(.dina(n1841), .dinb(n420), .dout(n1842));
  jand g00323(.dina(n1707), .dinb(n422), .dout(n1845));
  jnot g00324(.din(a46 ), .dout(n1851));
  jand g00325(.dina(b0 ), .dinb(n1851), .dout(n1852));
  jnot g00326(.din(n1852), .dout(n1853));
  jor  g00327(.dina(n19782), .dinb(n19583), .dout(quotient46 ));
  jand g00328(.dina(n419), .dinb(n418), .dout(n1910));
  jnot g00329(.din(a45 ), .dout(n2001));
  jand g00330(.dina(b0 ), .dinb(n2001), .dout(n2002));
  jnot g00331(.din(n2002), .dout(n2003));
  jand g00332(.dina(n19929), .dinb(n1910), .dout(quotient45 ));
  jand g00333(.dina(n2002), .dinb(n1910), .dout(n2156));
  jnot g00334(.din(a44 ), .dout(n2162));
  jand g00335(.dina(b0 ), .dinb(n2162), .dout(n2163));
  jnot g00336(.din(n2163), .dout(n2164));
  jand g00337(.dina(n20161), .dinb(n352), .dout(quotient44 ));
  jand g00338(.dina(n351), .dinb(b0 ), .dout(n2315));
  jand g00339(.dina(n2315), .dinb(n417), .dout(n2316));
  jand g00340(.dina(n2163), .dinb(n352), .dout(n2319));
  jnot g00341(.din(a43 ), .dout(n2325));
  jand g00342(.dina(b0 ), .dinb(n2325), .dout(n2326));
  jnot g00343(.din(n2326), .dout(n2327));
  jor  g00344(.dina(n20171), .dinb(n20407), .dout(quotient43 ));
  jnot g00345(.din(a42 ), .dout(n2503));
  jand g00346(.dina(b0 ), .dinb(n2503), .dout(n2504));
  jnot g00347(.din(n2504), .dout(n2505));
  jand g00348(.dina(n20579), .dinb(n2680), .dout(quotient42 ));
  jand g00349(.dina(n417), .dinb(n349), .dout(n2680));
  jand g00350(.dina(n2680), .dinb(b0 ), .dout(n2681));
  jand g00351(.dina(n2504), .dinb(n2680), .dout(n2684));
  jnot g00352(.din(a41 ), .dout(n2689));
  jand g00353(.dina(b0 ), .dinb(n2689), .dout(n2690));
  jnot g00354(.din(n2690), .dout(n2691));
  jnot g00355(.din(n20937), .dout(quotient41 ));
  jand g00356(.dina(n417), .dinb(b0 ), .dout(n2873));
  jnot g00357(.din(a40 ), .dout(n2880));
  jand g00358(.dina(b0 ), .dinb(n2880), .dout(n2881));
  jnot g00359(.din(n2881), .dout(n2882));
  jand g00360(.dina(n20943), .dinb(n417), .dout(n2951));
  jor  g00361(.dina(n2951), .dinb(n21125), .dout(quotient40 ));
  jnot g00362(.din(a39 ), .dout(n3076));
  jand g00363(.dina(b0 ), .dinb(n3076), .dout(n3077));
  jnot g00364(.din(n3077), .dout(n3078));
  jand g00365(.dina(n21323), .dinb(n415), .dout(quotient39 ));
  jand g00366(.dina(n3678), .dinb(n270), .dout(n3157));
  jnot g00367(.din(n3157), .dout(n3158));
  jand g00368(.dina(n415), .dinb(b0 ), .dout(n3302));
  jand g00369(.dina(n3077), .dinb(n415), .dout(n3305));
  jnot g00370(.din(a38 ), .dout(n3310));
  jand g00371(.dina(b0 ), .dinb(n3310), .dout(n3311));
  jnot g00372(.din(n21731), .dout(quotient38 ));
  jnot g00373(.din(n3311), .dout(n3412));
  jand g00374(.dina(n21939), .dinb(n270), .dout(n3469));
  jand g00375(.dina(n3469), .dinb(n3678), .dout(n3470));
  jand g00376(.dina(n414), .dinb(b0 ), .dout(n3592));
  jand g00377(.dina(n3592), .dinb(n272), .dout(n3593));
  jnot g00378(.din(a37 ), .dout(n3600));
  jand g00379(.dina(b0 ), .dinb(n3600), .dout(n3601));
  jnot g00380(.din(n3601), .dout(n3602));
  jand g00381(.dina(n414), .dinb(n271), .dout(n3678));
  jor  g00382(.dina(n21942), .dinb(n3470), .dout(quotient37 ));
  jnot g00383(.din(a36 ), .dout(n3822));
  jand g00384(.dina(b0 ), .dinb(n3822), .dout(n3823));
  jnot g00385(.din(n3823), .dout(n3824));
  jand g00386(.dina(n22167), .dinb(n414), .dout(quotient36 ));
  jand g00387(.dina(n413), .dinb(n341), .dout(n3911));
  jand g00388(.dina(n3823), .dinb(n414), .dout(n4047));
  jnot g00389(.din(a35 ), .dout(n4053));
  jand g00390(.dina(b0 ), .dinb(n4053), .dout(n4054));
  jnot g00391(.din(n4054), .dout(n4055));
  jand g00392(.dina(n22508), .dinb(n3911), .dout(quotient35 ));
  jand g00393(.dina(n413), .dinb(n340), .dout(n4145));
  jand g00394(.dina(n413), .dinb(b0 ), .dout(n4277));
  jand g00395(.dina(n4277), .dinb(n341), .dout(n4278));
  jand g00396(.dina(n4054), .dinb(n3911), .dout(n4281));
  jnot g00397(.din(a34 ), .dout(n4287));
  jand g00398(.dina(b0 ), .dinb(n4287), .dout(n4288));
  jnot g00399(.din(n4288), .dout(n4289));
  jor  g00400(.dina(n22518), .dinb(n22861), .dout(quotient34 ));
  jnot g00401(.din(a33 ), .dout(n4540));
  jand g00402(.dina(b0 ), .dinb(n4540), .dout(n4541));
  jnot g00403(.din(n4541), .dout(n4542));
  jand g00404(.dina(n23104), .dinb(n413), .dout(quotient33 ));
  jand g00405(.dina(n4541), .dinb(n413), .dout(n4789));
  jnot g00406(.din(a32 ), .dout(n4795));
  jand g00407(.dina(b0 ), .dinb(n4795), .dout(n4796));
  jnot g00408(.din(n4796), .dout(n4797));
  jand g00409(.dina(n23482), .dinb(n336), .dout(quotient32 ));
  jand g00410(.dina(n335), .dinb(b0 ), .dout(n5042));
  jand g00411(.dina(n5042), .dinb(n410), .dout(n5043));
  jand g00412(.dina(n4796), .dinb(n336), .dout(n5046));
  jnot g00413(.din(a31 ), .dout(n5052));
  jand g00414(.dina(b0 ), .dinb(n5052), .dout(n5053));
  jnot g00415(.din(n5053), .dout(n5054));
  jor  g00416(.dina(n23492), .dinb(n23871), .dout(quotient31 ));
  jnot g00417(.din(a30 ), .dout(n5326));
  jand g00418(.dina(b0 ), .dinb(n5326), .dout(n5327));
  jnot g00419(.din(n5327), .dout(n5328));
  jand g00420(.dina(n24269), .dinb(n5629), .dout(quotient30 ));
  jand g00421(.dina(n410), .dinb(n333), .dout(n5629));
  jand g00422(.dina(n5629), .dinb(b0 ), .dout(n5630));
  jand g00423(.dina(n5327), .dinb(n5629), .dout(n5633));
  jnot g00424(.din(a29 ), .dout(n5638));
  jand g00425(.dina(b0 ), .dinb(n5638), .dout(n5639));
  jnot g00426(.din(n24820), .dout(quotient29 ));
  jnot g00427(.din(n5639), .dout(n5777));
  jand g00428(.dina(n410), .dinb(b0 ), .dout(n6018));
  jnot g00429(.din(a28 ), .dout(n6025));
  jand g00430(.dina(b0 ), .dinb(n6025), .dout(n6026));
  jnot g00431(.din(n6026), .dout(n6027));
  jor  g00432(.dina(n25105), .dinb(n25106), .dout(quotient28 ));
  jnot g00433(.din(a27 ), .dout(n6320));
  jand g00434(.dina(b0 ), .dinb(n6320), .dout(n6321));
  jnot g00435(.din(n6321), .dout(n6322));
  jand g00436(.dina(n25539), .dinb(n408), .dout(quotient27 ));
  jand g00437(.dina(n407), .dinb(n326), .dout(n6436));
  jnot g00438(.din(n6436), .dout(n6437));
  jand g00439(.dina(n408), .dinb(b0 ), .dout(n6653));
  jand g00440(.dina(n6321), .dinb(n408), .dout(n6656));
  jnot g00441(.din(a26 ), .dout(n6661));
  jand g00442(.dina(b0 ), .dinb(n6661), .dout(n6662));
  jnot g00443(.din(n26138), .dout(quotient26 ));
  jnot g00444(.din(n6662), .dout(n6812));
  jand g00445(.dina(n405), .dinb(b0 ), .dout(n7074));
  jand g00446(.dina(n7074), .dinb(n282), .dout(n7075));
  jand g00447(.dina(n7075), .dinb(n277), .dout(n7076));
  jand g00448(.dina(n7076), .dinb(n326), .dout(n7077));
  jnot g00449(.din(a25 ), .dout(n7084));
  jand g00450(.dina(b0 ), .dinb(n7084), .dout(n7085));
  jnot g00451(.din(n7085), .dout(n7086));
  jor  g00452(.dina(n26446), .dinb(n26445), .dout(quotient25 ));
  jnot g00453(.din(a24 ), .dout(n7401));
  jand g00454(.dina(b0 ), .dinb(n7401), .dout(n7402));
  jnot g00455(.din(n7402), .dout(n7403));
  jand g00456(.dina(n26763), .dinb(n406), .dout(quotient24 ));
  jand g00457(.dina(n405), .dinb(n280), .dout(n7526));
  jand g00458(.dina(n7526), .dinb(n279), .dout(n7527));
  jand g00459(.dina(n7402), .dinb(n406), .dout(n7723));
  jnot g00460(.din(a23 ), .dout(n7729));
  jand g00461(.dina(b0 ), .dinb(n7729), .dout(n7730));
  jnot g00462(.din(n7730), .dout(n7731));
  jand g00463(.dina(n27247), .dinb(n7527), .dout(quotient23 ));
  jand g00464(.dina(n7074), .dinb(n281), .dout(n8054));
  jand g00465(.dina(n7730), .dinb(n7527), .dout(n8057));
  jnot g00466(.din(a22 ), .dout(n8063));
  jand g00467(.dina(b0 ), .dinb(n8063), .dout(n8064));
  jnot g00468(.din(n8064), .dout(n8065));
  jor  g00469(.dina(n27257), .dinb(n27744), .dout(quotient22 ));
  jnot g00470(.din(a21 ), .dout(n8446));
  jand g00471(.dina(b0 ), .dinb(n8446), .dout(n8447));
  jnot g00472(.din(n28419), .dout(quotient21 ));
  jnot g00473(.din(n8447), .dout(n8617));
  jnot g00474(.din(a20 ), .dout(n8923));
  jand g00475(.dina(b0 ), .dinb(n8923), .dout(n8924));
  jnot g00476(.din(n8924), .dout(n8925));
  jor  g00477(.dina(n28768), .dinb(n28426), .dout(quotient20 ));
  jand g00478(.dina(n403), .dinb(n318), .dout(n9062));
  jnot g00479(.din(a19 ), .dout(n9273));
  jand g00480(.dina(b0 ), .dinb(n9273), .dout(n9274));
  jnot g00481(.din(n9274), .dout(n9275));
  jor  g00482(.dina(n29128), .dinb(n29127), .dout(quotient19 ));
  jand g00483(.dina(n403), .dinb(n317), .dout(n9424));
  jnot g00484(.din(a18 ), .dout(n9648));
  jand g00485(.dina(b0 ), .dinb(n9648), .dout(n9649));
  jnot g00486(.din(n9649), .dout(n9650));
  jand g00487(.dina(n29491), .dinb(n9424), .dout(quotient18 ));
  jand g00488(.dina(n29500), .dinb(n317), .dout(n9795));
  jand g00489(.dina(n9795), .dinb(n403), .dout(n9796));
  jand g00490(.dina(n403), .dinb(b0 ), .dout(n10014));
  jand g00491(.dina(n10014), .dinb(n317), .dout(n10015));
  jand g00492(.dina(n9649), .dinb(n9424), .dout(n10018));
  jnot g00493(.din(a17 ), .dout(n10024));
  jand g00494(.dina(b0 ), .dinb(n10024), .dout(n10025));
  jnot g00495(.din(n10025), .dout(n10026));
  jor  g00496(.dina(n30046), .dinb(n9796), .dout(quotient17 ));
  jnot g00497(.din(n9424), .dout(n10176));
  jnot g00498(.din(a16 ), .dout(n10406));
  jand g00499(.dina(b0 ), .dinb(n10406), .dout(n10407));
  jnot g00500(.din(n10407), .dout(n10408));
  jor  g00501(.dina(n30427), .dinb(n30058), .dout(quotient16 ));
  jnot g00502(.din(a15 ), .dout(n10797));
  jand g00503(.dina(b0 ), .dinb(n10797), .dout(n10798));
  jnot g00504(.din(n10798), .dout(n10799));
  jand g00505(.dina(n30816), .dinb(n312), .dout(quotient15 ));
  jand g00506(.dina(n30825), .dinb(n286), .dout(n10953));
  jand g00507(.dina(n10953), .dinb(n311), .dout(n10954));
  jand g00508(.dina(n312), .dinb(b0 ), .dout(n11186));
  jand g00509(.dina(n10798), .dinb(n312), .dout(n11189));
  jnot g00510(.din(a14 ), .dout(n11195));
  jand g00511(.dina(b0 ), .dinb(n11195), .dout(n11196));
  jnot g00512(.din(n11196), .dout(n11197));
  jor  g00513(.dina(n31409), .dinb(n10954), .dout(quotient14 ));
  jnot g00514(.din(a13 ), .dout(n11605));
  jand g00515(.dina(b0 ), .dinb(n11605), .dout(n11606));
  jnot g00516(.din(n11606), .dout(n11607));
  jand g00517(.dina(n31815), .dinb(n310), .dout(quotient13 ));
  jnot g00518(.din(a12 ), .dout(n12015));
  jand g00519(.dina(b0 ), .dinb(n12015), .dout(n12016));
  jnot g00520(.din(n12016), .dout(n12017));
  jand g00521(.dina(n32229), .dinb(n309), .dout(quotient12 ));
  jand g00522(.dina(n309), .dinb(b0 ), .dout(n12427));
  jand g00523(.dina(n12016), .dinb(n309), .dout(n12430));
  jnot g00524(.din(a11 ), .dout(n12436));
  jand g00525(.dina(b0 ), .dinb(n12436), .dout(n12437));
  jnot g00526(.din(n12437), .dout(n12438));
  jand g00527(.dina(n32861), .dinb(n308), .dout(quotient11 ));
  jnot g00528(.din(a10 ), .dout(n12863));
  jand g00529(.dina(b0 ), .dinb(n12863), .dout(n12864));
  jnot g00530(.din(n12864), .dout(n12865));
  jor  g00531(.dina(n33287), .dinb(n32871), .dout(n13022));
  jor  g00532(.dina(n32873), .dinb(n838), .dout(n13025));
  jnot g00533(.din(n13025), .dout(n13026));
  jand g00534(.dina(n13026), .dinb(n13022), .dout(quotient10 ));
  jnot g00535(.din(a9 ), .dout(n13300));
  jand g00536(.dina(b0 ), .dinb(n13300), .dout(n13301));
  jnot g00537(.din(n13301), .dout(n13302));
  jand g00538(.dina(n33725), .dinb(n306), .dout(quotient9 ));
  jand g00539(.dina(n306), .dinb(b0 ), .dout(n13732));
  jand g00540(.dina(n13301), .dinb(n306), .dout(n13735));
  jnot g00541(.din(a8 ), .dout(n13741));
  jand g00542(.dina(b0 ), .dinb(n13741), .dout(n13742));
  jnot g00543(.din(n13742), .dout(n13743));
  jand g00544(.dina(n33735), .dinb(n292), .dout(n13910));
  jand g00545(.dina(n13910), .dinb(n305), .dout(n13916));
  jor  g00546(.dina(n13916), .dinb(n34393), .dout(quotient8 ));
  jnot g00547(.din(a7 ), .dout(n14203));
  jand g00548(.dina(b0 ), .dinb(n14203), .dout(n14204));
  jnot g00549(.din(n14204), .dout(n14205));
  jand g00550(.dina(n34844), .dinb(n304), .dout(quotient7 ));
  jnot g00551(.din(a6 ), .dout(n14661));
  jand g00552(.dina(b0 ), .dinb(n14661), .dout(n14662));
  jnot g00553(.din(n14662), .dout(n14663));
  jand g00554(.dina(n35305), .dinb(n303), .dout(quotient6 ));
  jand g00555(.dina(n303), .dinb(b0 ), .dout(n15122));
  jand g00556(.dina(n14662), .dinb(n303), .dout(n15125));
  jnot g00557(.din(a5 ), .dout(n15131));
  jand g00558(.dina(b0 ), .dinb(n15131), .dout(n15132));
  jnot g00559(.din(n15132), .dout(n15133));
  jor  g00560(.dina(n36008), .dinb(n36009), .dout(quotient5 ));
  jnot g00561(.din(a4 ), .dout(n15612));
  jand g00562(.dina(b0 ), .dinb(n15612), .dout(n15613));
  jnot g00563(.din(n15613), .dout(n15614));
  jand g00564(.dina(n36720), .dinb(n36716), .dout(quotient4 ));
  jnot g00565(.din(a3 ), .dout(n16095));
  jand g00566(.dina(b0 ), .dinb(n16095), .dout(n16096));
  jnot g00567(.din(n16096), .dout(n16097));
  jand g00568(.dina(n37204), .dinb(n37200), .dout(quotient3 ));
  jxor g00569(.dina(n37690), .dinb(n257), .dout(n16289));
  jnot g00570(.din(a2 ), .dout(n16585));
  jand g00571(.dina(b0 ), .dinb(n16585), .dout(n16586));
  jnot g00572(.din(n16586), .dout(n16587));
  jand g00573(.dina(n37938), .dinb(n16289), .dout(n16769));
  jor  g00574(.dina(n37691), .dinb(n16769), .dout(quotient2 ));
  jnot g00575(.din(a1 ), .dout(n17077));
  jand g00576(.dina(b0 ), .dinb(n17077), .dout(n17078));
  jnot g00577(.din(n17078), .dout(n17079));
  jand g00578(.dina(n37935), .dinb(n299), .dout(n17269));
  jxor g00579(.dina(n37935), .dinb(n298), .dout(n17514));
  jand g00580(.dina(n17514), .dinb(n256), .dout(n17515));
  jand g00581(.dina(n17515), .dinb(n38437), .dout(n17523));
  jor  g00582(.dina(n17523), .dinb(n17269), .dout(quotient1 ));
  jor  g00583(.dina(n38460), .dinb(n38465), .dout(n17542));
  jor  g00584(.dina(n38479), .dinb(n294), .dout(n17552));
  jor  g00585(.dina(n38480), .dinb(n38485), .dout(n17559));
  jor  g00586(.dina(n38490), .dinb(n38495), .dout(n17570));
  jor  g00587(.dina(n38509), .dinb(n288), .dout(n17580));
  jor  g00588(.dina(n38519), .dinb(n286), .dout(n17590));
  jor  g00589(.dina(n38514), .dinb(n287), .dout(n17591));
  jand g00590(.dina(n17591), .dinb(n17590), .dout(n17592));
  jor  g00591(.dina(n38529), .dinb(n284), .dout(n17597));
  jor  g00592(.dina(n38524), .dinb(n285), .dout(n17602));
  jand g00593(.dina(n17602), .dinb(n17597), .dout(n17603));
  jor  g00594(.dina(n38539), .dinb(n316), .dout(n17608));
  jor  g00595(.dina(n38540), .dinb(n38545), .dout(n17615));
  jor  g00596(.dina(n38559), .dinb(n279), .dout(n17625));
  jor  g00597(.dina(n38554), .dinb(n280), .dout(n17626));
  jand g00598(.dina(n17626), .dinb(n17625), .dout(n17627));
  jor  g00599(.dina(n38569), .dinb(n277), .dout(n17632));
  jor  g00600(.dina(n38570), .dinb(n38575), .dout(n17639));
  jor  g00601(.dina(n38580), .dinb(n38585), .dout(n17650));
  jor  g00602(.dina(n38599), .dinb(n332), .dout(n17660));
  jor  g00603(.dina(n38594), .dinb(n333), .dout(n17661));
  jand g00604(.dina(n17661), .dinb(n17660), .dout(n17662));
  jor  g00605(.dina(n38609), .dinb(n275), .dout(n17667));
  jor  g00606(.dina(n38604), .dinb(n331), .dout(n17672));
  jand g00607(.dina(n17672), .dinb(n17667), .dout(n17673));
  jor  g00608(.dina(n38619), .dinb(n339), .dout(n17678));
  jor  g00609(.dina(n38614), .dinb(n340), .dout(n17683));
  jand g00610(.dina(n17683), .dinb(n17678), .dout(n17684));
  jor  g00611(.dina(n38629), .dinb(n271), .dout(n17689));
  jor  g00612(.dina(n38630), .dinb(n38635), .dout(n17696));
  jor  g00613(.dina(n38640), .dinb(n38645), .dout(n17707));
  jor  g00614(.dina(n38650), .dinb(n38655), .dout(n17718));
  jor  g00615(.dina(n38660), .dinb(n38665), .dout(n17729));
  jor  g00616(.dina(n38670), .dinb(n38675), .dout(n17740));
  jor  g00617(.dina(n38680), .dinb(n38685), .dout(n17751));
  jor  g00618(.dina(n38690), .dinb(n38695), .dout(n17762));
  jor  g00619(.dina(n38709), .dinb(n359), .dout(n17772));
  jor  g00620(.dina(n38710), .dinb(n38715), .dout(n17779));
  jor  g00621(.dina(n38729), .dinb(n265), .dout(n17789));
  jor  g00622(.dina(n38724), .dinb(n367), .dout(n17790));
  jor  g00623(.dina(n38739), .dinb(n377), .dout(n17801));
  jor  g00624(.dina(n38734), .dinb(n378), .dout(n17802));
  jor  g00625(.dina(n38749), .dinb(n264), .dout(n17813));
  jor  g00626(.dina(n38744), .dinb(n376), .dout(n17814));
  jnot g00627(.din(b0 ), .dout(n17822));
  jor  g00628(.dina(n17822), .dinb(a0 ), .dout(n17823));
  jor  g00629(.dina(n38767), .dinb(n38750), .dout(n17833));
  jand g00630(.dina(n17833), .dinb(n17814), .dout(n17834));
  jand g00631(.dina(n17834), .dinb(n17813), .dout(n17835));
  jor  g00632(.dina(n17835), .dinb(n38740), .dout(n17836));
  jor  g00633(.dina(n17836), .dinb(n38745), .dout(n17837));
  jand g00634(.dina(n17837), .dinb(n17802), .dout(n17838));
  jand g00635(.dina(n17838), .dinb(n17801), .dout(n17839));
  jor  g00636(.dina(n17839), .dinb(n38730), .dout(n17840));
  jor  g00637(.dina(n17840), .dinb(n38735), .dout(n17841));
  jand g00638(.dina(n17841), .dinb(n17790), .dout(n17842));
  jand g00639(.dina(n17842), .dinb(n17789), .dout(n17843));
  jor  g00640(.dina(n38720), .dinb(n17843), .dout(n17849));
  jor  g00641(.dina(n17849), .dinb(n38725), .dout(n17850));
  jor  g00642(.dina(n38719), .dinb(n368), .dout(n17851));
  jor  g00643(.dina(n38714), .dinb(n369), .dout(n17852));
  jand g00644(.dina(n17852), .dinb(n17851), .dout(n17853));
  jand g00645(.dina(n17853), .dinb(n17850), .dout(n17854));
  jor  g00646(.dina(n17854), .dinb(n17779), .dout(n17855));
  jor  g00647(.dina(n38704), .dinb(n363), .dout(n17856));
  jand g00648(.dina(n17856), .dinb(n17855), .dout(n17857));
  jand g00649(.dina(n17857), .dinb(n17772), .dout(n17858));
  jor  g00650(.dina(n38700), .dinb(n17858), .dout(n17864));
  jor  g00651(.dina(n17864), .dinb(n38705), .dout(n17865));
  jor  g00652(.dina(n38699), .dinb(n360), .dout(n17866));
  jor  g00653(.dina(n38694), .dinb(n361), .dout(n17867));
  jand g00654(.dina(n17867), .dinb(n17866), .dout(n17868));
  jand g00655(.dina(n17868), .dinb(n17865), .dout(n17869));
  jor  g00656(.dina(n17869), .dinb(n17762), .dout(n17870));
  jor  g00657(.dina(n38689), .dinb(n364), .dout(n17871));
  jor  g00658(.dina(n38684), .dinb(n355), .dout(n17872));
  jand g00659(.dina(n17872), .dinb(n17871), .dout(n17873));
  jand g00660(.dina(n17873), .dinb(n17870), .dout(n17874));
  jor  g00661(.dina(n17874), .dinb(n17751), .dout(n17875));
  jor  g00662(.dina(n38679), .dinb(n356), .dout(n17876));
  jor  g00663(.dina(n38674), .dinb(n266), .dout(n17877));
  jand g00664(.dina(n17877), .dinb(n17876), .dout(n17878));
  jand g00665(.dina(n17878), .dinb(n17875), .dout(n17879));
  jor  g00666(.dina(n17879), .dinb(n17740), .dout(n17880));
  jor  g00667(.dina(n38669), .dinb(n267), .dout(n17881));
  jor  g00668(.dina(n38664), .dinb(n347), .dout(n17882));
  jand g00669(.dina(n17882), .dinb(n17881), .dout(n17883));
  jand g00670(.dina(n17883), .dinb(n17880), .dout(n17884));
  jor  g00671(.dina(n17884), .dinb(n17729), .dout(n17885));
  jor  g00672(.dina(n38659), .dinb(n348), .dout(n17886));
  jor  g00673(.dina(n38654), .dinb(n349), .dout(n17887));
  jand g00674(.dina(n17887), .dinb(n17886), .dout(n17888));
  jand g00675(.dina(n17888), .dinb(n17885), .dout(n17889));
  jor  g00676(.dina(n17889), .dinb(n17718), .dout(n17890));
  jor  g00677(.dina(n38649), .dinb(n268), .dout(n17891));
  jor  g00678(.dina(n38644), .dinb(n274), .dout(n17892));
  jand g00679(.dina(n17892), .dinb(n17891), .dout(n17893));
  jand g00680(.dina(n17893), .dinb(n17890), .dout(n17894));
  jor  g00681(.dina(n17894), .dinb(n17707), .dout(n17895));
  jor  g00682(.dina(n38639), .dinb(n269), .dout(n17896));
  jor  g00683(.dina(n38634), .dinb(n270), .dout(n17897));
  jand g00684(.dina(n17897), .dinb(n17896), .dout(n17898));
  jand g00685(.dina(n17898), .dinb(n17895), .dout(n17899));
  jor  g00686(.dina(n17899), .dinb(n17696), .dout(n17900));
  jor  g00687(.dina(n38624), .dinb(n338), .dout(n17905));
  jand g00688(.dina(n17905), .dinb(n17900), .dout(n17906));
  jand g00689(.dina(n17906), .dinb(n17689), .dout(n17907));
  jor  g00690(.dina(n38620), .dinb(n38625), .dout(n17910));
  jor  g00691(.dina(n17910), .dinb(n17907), .dout(n17911));
  jand g00692(.dina(n17911), .dinb(n17684), .dout(n17912));
  jor  g00693(.dina(n38610), .dinb(n38615), .dout(n17915));
  jor  g00694(.dina(n17915), .dinb(n17912), .dout(n17916));
  jand g00695(.dina(n17916), .dinb(n17673), .dout(n17917));
  jor  g00696(.dina(n38600), .dinb(n38605), .dout(n17920));
  jor  g00697(.dina(n17920), .dinb(n17917), .dout(n17921));
  jand g00698(.dina(n17921), .dinb(n17662), .dout(n17922));
  jor  g00699(.dina(n38590), .dinb(n17922), .dout(n17928));
  jor  g00700(.dina(n17928), .dinb(n38595), .dout(n17929));
  jor  g00701(.dina(n38589), .dinb(n276), .dout(n17930));
  jor  g00702(.dina(n38584), .dinb(n324), .dout(n17931));
  jand g00703(.dina(n17931), .dinb(n17930), .dout(n17932));
  jand g00704(.dina(n17932), .dinb(n17929), .dout(n17933));
  jor  g00705(.dina(n17933), .dinb(n17650), .dout(n17934));
  jor  g00706(.dina(n38579), .dinb(n325), .dout(n17935));
  jor  g00707(.dina(n38574), .dinb(n326), .dout(n17936));
  jand g00708(.dina(n17936), .dinb(n17935), .dout(n17937));
  jand g00709(.dina(n17937), .dinb(n17934), .dout(n17938));
  jor  g00710(.dina(n17938), .dinb(n17639), .dout(n17939));
  jor  g00711(.dina(n38564), .dinb(n278), .dout(n17944));
  jand g00712(.dina(n17944), .dinb(n17939), .dout(n17945));
  jand g00713(.dina(n17945), .dinb(n17632), .dout(n17946));
  jor  g00714(.dina(n38560), .dinb(n38565), .dout(n17949));
  jor  g00715(.dina(n17949), .dinb(n17946), .dout(n17950));
  jand g00716(.dina(n17950), .dinb(n17627), .dout(n17951));
  jor  g00717(.dina(n38550), .dinb(n17951), .dout(n17957));
  jor  g00718(.dina(n17957), .dinb(n38555), .dout(n17958));
  jor  g00719(.dina(n38549), .dinb(n283), .dout(n17959));
  jor  g00720(.dina(n38544), .dinb(n315), .dout(n17960));
  jand g00721(.dina(n17960), .dinb(n17959), .dout(n17961));
  jand g00722(.dina(n17961), .dinb(n17958), .dout(n17962));
  jor  g00723(.dina(n17962), .dinb(n17615), .dout(n17963));
  jor  g00724(.dina(n38534), .dinb(n317), .dout(n17968));
  jand g00725(.dina(n17968), .dinb(n17963), .dout(n17969));
  jand g00726(.dina(n17969), .dinb(n17608), .dout(n17970));
  jor  g00727(.dina(n38530), .dinb(n38535), .dout(n17973));
  jor  g00728(.dina(n17973), .dinb(n17970), .dout(n17974));
  jand g00729(.dina(n17974), .dinb(n17603), .dout(n17975));
  jor  g00730(.dina(n38520), .dinb(n38525), .dout(n17978));
  jor  g00731(.dina(n17978), .dinb(n17975), .dout(n17979));
  jand g00732(.dina(n17979), .dinb(n17592), .dout(n17980));
  jor  g00733(.dina(n38510), .dinb(n17980), .dout(n17982));
  jor  g00734(.dina(n17982), .dinb(n38515), .dout(n17983));
  jor  g00735(.dina(n38504), .dinb(n289), .dout(n17984));
  jand g00736(.dina(n17984), .dinb(n17983), .dout(n17985));
  jand g00737(.dina(n17985), .dinb(n17580), .dout(n17986));
  jor  g00738(.dina(n38500), .dinb(n17986), .dout(n17992));
  jor  g00739(.dina(n17992), .dinb(n38505), .dout(n17993));
  jor  g00740(.dina(n38499), .dinb(n290), .dout(n17994));
  jor  g00741(.dina(n38494), .dinb(n291), .dout(n17995));
  jand g00742(.dina(n17995), .dinb(n17994), .dout(n17996));
  jand g00743(.dina(n17996), .dinb(n17993), .dout(n17997));
  jor  g00744(.dina(n17997), .dinb(n17570), .dout(n17998));
  jor  g00745(.dina(n38489), .dinb(n292), .dout(n17999));
  jor  g00746(.dina(n38484), .dinb(n293), .dout(n18000));
  jand g00747(.dina(n18000), .dinb(n17999), .dout(n18001));
  jand g00748(.dina(n18001), .dinb(n17998), .dout(n18002));
  jor  g00749(.dina(n18002), .dinb(n17559), .dout(n18003));
  jor  g00750(.dina(n38474), .dinb(n295), .dout(n18004));
  jand g00751(.dina(n18004), .dinb(n18003), .dout(n18005));
  jand g00752(.dina(n18005), .dinb(n17552), .dout(n18006));
  jor  g00753(.dina(n38470), .dinb(n18006), .dout(n18012));
  jor  g00754(.dina(n18012), .dinb(n38475), .dout(n18013));
  jor  g00755(.dina(n38469), .dinb(n296), .dout(n18014));
  jor  g00756(.dina(n38464), .dinb(n297), .dout(n18015));
  jand g00757(.dina(n18015), .dinb(n18014), .dout(n18016));
  jand g00758(.dina(n18016), .dinb(n18013), .dout(n18017));
  jor  g00759(.dina(n18017), .dinb(n17542), .dout(n18018));
  jor  g00760(.dina(n38459), .dinb(n257), .dout(n18019));
  jor  g00761(.dina(n38454), .dinb(n298), .dout(n18020));
  jand g00762(.dina(n18020), .dinb(n18019), .dout(n18021));
  jand g00763(.dina(n18021), .dinb(n18018), .dout(n18022));
  jor  g00764(.dina(n18022), .dinb(n38455), .dout(n18023));
  jand g00765(.dina(n18023), .dinb(n38450), .dout(n18024));
  jor  g00766(.dina(n18024), .dinb(n38448), .dout(quotient0 ));
  jand g00767(.dina(n438), .dinb(n18035), .dout(quotient62 ));
  jand g00768(.dina(n486), .dinb(n390), .dout(quotient63 ));
  jor  g00769(.dina(n869), .dinb(b7 ), .dout(n18028));
  jnot g00770(.din(n380), .dout(n18029));
  jor  g00771(.dina(n18029), .dinb(n18028), .dout(n18030));
  jor  g00772(.dina(n18030), .dinb(b3 ), .dout(n18031));
  jor  g00773(.dina(n18031), .dinb(n17822), .dout(n18032));
  jor  g00774(.dina(n388), .dinb(n18032), .dout(n18033));
  jand g00775(.dina(n18033), .dinb(n395), .dout(n18034));
  jor  g00776(.dina(n18034), .dinb(n262), .dout(n18035));
  jand g00777(.dina(n18035), .dinb(n435), .dout(n18036));
  jor  g00778(.dina(n18036), .dinb(n258), .dout(n18037));
  jnot g00779(.din(n447), .dout(n18041));
  jor  g00780(.dina(n18037), .dinb(n448), .dout(n18042));
  jand g00781(.dina(n18042), .dinb(n18041), .dout(n18043));
  jor  g00782(.dina(n18043), .dinb(b2 ), .dout(n18044));
  jand g00783(.dina(n18033), .dinb(a63 ), .dout(n18045));
  jnot g00784(.din(n18045), .dout(n18046));
  jor  g00785(.dina(n18046), .dinb(n456), .dout(n18047));
  jand g00786(.dina(n18043), .dinb(b2 ), .dout(n18048));
  jor  g00787(.dina(n18048), .dinb(n18047), .dout(n18049));
  jand g00788(.dina(n18049), .dinb(n18044), .dout(n18050));
  jor  g00789(.dina(n18050), .dinb(n477), .dout(n18051));
  jxor g00790(.dina(n18051), .dinb(n18037), .dout(n18052));
  jnot g00791(.din(n18052), .dout(n18053));
  jor  g00792(.dina(n18050), .dinb(n18032), .dout(n18054));
  jand g00793(.dina(n18054), .dinb(a61 ), .dout(n18055));
  jnot g00794(.din(n18044), .dout(n18056));
  jnot g00795(.din(n18047), .dout(n18057));
  jnot g00796(.din(n435), .dout(n18058));
  jnot g00797(.din(n395), .dout(n18059));
  jand g00798(.dina(n387), .dinb(n383), .dout(n18060));
  jor  g00799(.dina(n18060), .dinb(n18059), .dout(n18061));
  jand g00800(.dina(n18061), .dinb(n263), .dout(n18062));
  jor  g00801(.dina(n18062), .dinb(n18058), .dout(n18063));
  jand g00802(.dina(n18063), .dinb(a62 ), .dout(n18064));
  jand g00803(.dina(n18064), .dinb(n449), .dout(n18066));
  jor  g00804(.dina(n18066), .dinb(n447), .dout(n18067));
  jor  g00805(.dina(n18067), .dinb(n386), .dout(n18068));
  jand g00806(.dina(n18068), .dinb(n18057), .dout(n18069));
  jor  g00807(.dina(n18069), .dinb(n18056), .dout(n18070));
  jand g00808(.dina(n18070), .dinb(n487), .dout(n18071));
  jor  g00809(.dina(n18071), .dinb(n18055), .dout(n18072));
  jand g00810(.dina(n18072), .dinb(n493), .dout(n18073));
  jor  g00811(.dina(n18073), .dinb(n483), .dout(n18074));
  jand g00812(.dina(n18074), .dinb(n386), .dout(n18075));
  jor  g00813(.dina(n18074), .dinb(n386), .dout(n18076));
  jand g00814(.dina(n18076), .dinb(n18052), .dout(n18077));
  jor  g00815(.dina(n18077), .dinb(n18075), .dout(n18078));
  jxor g00816(.dina(n18043), .dinb(b2 ), .dout(n18079));
  jand g00817(.dina(n18079), .dinb(n486), .dout(n18080));
  jor  g00818(.dina(n18080), .dinb(n18047), .dout(n18081));
  jand g00819(.dina(n18081), .dinb(b3 ), .dout(n18082));
  jnot g00820(.din(n18082), .dout(n18083));
  jand g00821(.dina(n18083), .dinb(n18078), .dout(n18084));
  jnot g00822(.din(n18081), .dout(n18085));
  jand g00823(.dina(n18085), .dinb(n264), .dout(n18086));
  jor  g00824(.dina(n18086), .dinb(n18084), .dout(n18087));
  jand g00825(.dina(n18087), .dinb(n381), .dout(n18088));
  jxor g00826(.dina(n18074), .dinb(n386), .dout(n18089));
  jand g00827(.dina(n18089), .dinb(n18088), .dout(n18090));
  jxor g00828(.dina(n18090), .dinb(n18053), .dout(n18091));
  jnot g00829(.din(n18091), .dout(n18092));
  jor  g00830(.dina(n18091), .dinb(b3 ), .dout(n18093));
  jand g00831(.dina(n18091), .dinb(b3 ), .dout(n18094));
  jand g00832(.dina(n18087), .dinb(n520), .dout(n18095));
  jxor g00833(.dina(n18095), .dinb(n18072), .dout(n18096));
  jand g00834(.dina(n18096), .dinb(n386), .dout(n18097));
  jnot g00835(.din(n18097), .dout(n18098));
  jnot g00836(.din(n18096), .dout(n18099));
  jand g00837(.dina(n18099), .dinb(b2 ), .dout(n18100));
  jnot g00838(.din(n529), .dout(n18101));
  jand g00839(.dina(n18087), .dinb(n433), .dout(n18102));
  jor  g00840(.dina(n18102), .dinb(n480), .dout(n18103));
  jnot g00841(.din(n534), .dout(n18104));
  jnot g00842(.din(n18075), .dout(n18105));
  jnot g00843(.din(n483), .dout(n18106));
  jand g00844(.dina(n18070), .dinb(n383), .dout(n18107));
  jor  g00845(.dina(n18107), .dinb(n444), .dout(n18108));
  jnot g00846(.din(n487), .dout(n18109));
  jor  g00847(.dina(n18050), .dinb(n18109), .dout(n18110));
  jand g00848(.dina(n18110), .dinb(n18108), .dout(n18111));
  jor  g00849(.dina(n18111), .dinb(n492), .dout(n18112));
  jand g00850(.dina(n18112), .dinb(n18106), .dout(n18113));
  jand g00851(.dina(n18113), .dinb(b2 ), .dout(n18114));
  jor  g00852(.dina(n18114), .dinb(n18053), .dout(n18115));
  jand g00853(.dina(n18115), .dinb(n18105), .dout(n18116));
  jor  g00854(.dina(n18082), .dinb(n18116), .dout(n18117));
  jnot g00855(.din(n18086), .dout(n18118));
  jand g00856(.dina(n18118), .dinb(n18117), .dout(n18119));
  jor  g00857(.dina(n18119), .dinb(n18104), .dout(n18120));
  jand g00858(.dina(n18120), .dinb(n18103), .dout(n18121));
  jor  g00859(.dina(n18121), .dinb(n530), .dout(n18122));
  jand g00860(.dina(n18122), .dinb(n18101), .dout(n18123));
  jor  g00861(.dina(n18123), .dinb(n18100), .dout(n18124));
  jand g00862(.dina(n18124), .dinb(n18098), .dout(n18125));
  jor  g00863(.dina(n18125), .dinb(n18094), .dout(n18126));
  jand g00864(.dina(n18126), .dinb(n18093), .dout(n18127));
  jor  g00865(.dina(n18127), .dinb(b4 ), .dout(n18128));
  jor  g00866(.dina(n18088), .dinb(n18081), .dout(n18129));
  jand g00867(.dina(n18086), .dinb(n18078), .dout(n18130));
  jnot g00868(.din(n18130), .dout(n18131));
  jand g00869(.dina(n18131), .dinb(n18129), .dout(n18132));
  jand g00870(.dina(n18127), .dinb(b4 ), .dout(n18133));
  jor  g00871(.dina(n18133), .dinb(n18132), .dout(n18134));
  jand g00872(.dina(n18134), .dinb(n18128), .dout(n18135));
  jor  g00873(.dina(n18135), .dinb(n572), .dout(n18136));
  jxor g00874(.dina(n18125), .dinb(n264), .dout(n18137));
  jor  g00875(.dina(n18137), .dinb(n18136), .dout(n18138));
  jxor g00876(.dina(n18138), .dinb(n18092), .dout(n18139));
  jnot g00877(.din(n18139), .dout(n18140));
  jnot g00878(.din(n18093), .dout(n18141));
  jnot g00879(.din(n18094), .dout(n18142));
  jnot g00880(.din(n18100), .dout(n18143));
  jnot g00881(.din(n433), .dout(n18144));
  jor  g00882(.dina(n18119), .dinb(n18144), .dout(n18145));
  jand g00883(.dina(n18145), .dinb(a60 ), .dout(n18146));
  jand g00884(.dina(n18087), .dinb(n534), .dout(n18147));
  jor  g00885(.dina(n18147), .dinb(n18146), .dout(n18148));
  jand g00886(.dina(n18148), .dinb(n531), .dout(n18149));
  jor  g00887(.dina(n18149), .dinb(n529), .dout(n18150));
  jand g00888(.dina(n18150), .dinb(n18143), .dout(n18151));
  jor  g00889(.dina(n18151), .dinb(n18097), .dout(n18152));
  jand g00890(.dina(n18152), .dinb(n18142), .dout(n18153));
  jor  g00891(.dina(n18153), .dinb(n18141), .dout(n18154));
  jor  g00892(.dina(n18154), .dinb(n376), .dout(n18155));
  jand g00893(.dina(n18128), .dinb(n431), .dout(n18156));
  jand g00894(.dina(n18156), .dinb(n18155), .dout(n18157));
  jor  g00895(.dina(n18157), .dinb(n18132), .dout(n18158));
  jnot g00896(.din(n18158), .dout(n18159));
  jand g00897(.dina(n18159), .dinb(n377), .dout(n18160));
  jand g00898(.dina(n18160), .dinb(n610), .dout(n18161));
  jand g00899(.dina(n18140), .dinb(n376), .dout(n18162));
  jxor g00900(.dina(n18123), .dinb(n386), .dout(n18163));
  jor  g00901(.dina(n18163), .dinb(n18136), .dout(n18164));
  jxor g00902(.dina(n18164), .dinb(n18099), .dout(n18165));
  jand g00903(.dina(n18165), .dinb(n264), .dout(n18166));
  jor  g00904(.dina(n18135), .dinb(n574), .dout(n18167));
  jxor g00905(.dina(n18167), .dinb(n18148), .dout(n18168));
  jnot g00906(.din(n18168), .dout(n18169));
  jand g00907(.dina(n18169), .dinb(n386), .dout(n18170));
  jnot g00908(.din(n580), .dout(n18171));
  jor  g00909(.dina(n18135), .dinb(n18171), .dout(n18172));
  jand g00910(.dina(n18172), .dinb(a59 ), .dout(n18173));
  jnot g00911(.din(n18128), .dout(n18174));
  jnot g00912(.din(n18132), .dout(n18175));
  jand g00913(.dina(n18155), .dinb(n18175), .dout(n18176));
  jor  g00914(.dina(n18176), .dinb(n18174), .dout(n18177));
  jand g00915(.dina(n18177), .dinb(n583), .dout(n18178));
  jor  g00916(.dina(n18178), .dinb(n18173), .dout(n18179));
  jand g00917(.dina(n18179), .dinb(n259), .dout(n18180));
  jxor g00918(.dina(n18179), .dinb(n259), .dout(n18181));
  jand g00919(.dina(n18181), .dinb(n591), .dout(n18182));
  jor  g00920(.dina(n18182), .dinb(n18180), .dout(n18183));
  jxor g00921(.dina(n18168), .dinb(b2 ), .dout(n18184));
  jand g00922(.dina(n18184), .dinb(n18183), .dout(n18185));
  jor  g00923(.dina(n18185), .dinb(n18170), .dout(n18186));
  jxor g00924(.dina(n18165), .dinb(n264), .dout(n18187));
  jand g00925(.dina(n18187), .dinb(n18186), .dout(n18188));
  jor  g00926(.dina(n18188), .dinb(n18166), .dout(n18189));
  jxor g00927(.dina(n18139), .dinb(b4 ), .dout(n18190));
  jand g00928(.dina(n18190), .dinb(n18189), .dout(n18191));
  jor  g00929(.dina(n18191), .dinb(n18162), .dout(n18192));
  jxor g00930(.dina(n18158), .dinb(b5 ), .dout(n18193));
  jand g00931(.dina(n18193), .dinb(n18192), .dout(n18194));
  jand g00932(.dina(n18194), .dinb(n610), .dout(n18195));
  jor  g00933(.dina(n18195), .dinb(n18161), .dout(n18196));
  jnot g00934(.din(n18196), .dout(n18197));
  jand g00935(.dina(n18197), .dinb(n18140), .dout(n18198));
  jxor g00936(.dina(n18190), .dinb(n18189), .dout(n18199));
  jand g00937(.dina(n18199), .dinb(n18196), .dout(n18200));
  jor  g00938(.dina(n18200), .dinb(n18198), .dout(n18201));
  jxor g00939(.dina(n18193), .dinb(n18192), .dout(n18202));
  jand g00940(.dina(n18202), .dinb(n18161), .dout(n18203));
  jand g00941(.dina(n18197), .dinb(n18159), .dout(n18204));
  jor  g00942(.dina(n18204), .dinb(n18203), .dout(n18205));
  jand g00943(.dina(n18205), .dinb(n378), .dout(n18206));
  jnot g00944(.din(n18205), .dout(n18207));
  jand g00945(.dina(n18207), .dinb(b6 ), .dout(n18208));
  jnot g00946(.din(n18208), .dout(n18209));
  jand g00947(.dina(n18201), .dinb(n377), .dout(n18210));
  jand g00948(.dina(n18197), .dinb(n18165), .dout(n18211));
  jxor g00949(.dina(n18187), .dinb(n18186), .dout(n18212));
  jand g00950(.dina(n18212), .dinb(n18196), .dout(n18213));
  jor  g00951(.dina(n18213), .dinb(n18211), .dout(n18214));
  jand g00952(.dina(n18214), .dinb(n376), .dout(n18215));
  jor  g00953(.dina(n18196), .dinb(n18168), .dout(n18216));
  jxor g00954(.dina(n18184), .dinb(n18183), .dout(n18217));
  jnot g00955(.din(n18217), .dout(n18218));
  jor  g00956(.dina(n18218), .dinb(n18197), .dout(n18219));
  jand g00957(.dina(n18219), .dinb(n18216), .dout(n18220));
  jnot g00958(.din(n18220), .dout(n18221));
  jand g00959(.dina(n18221), .dinb(n264), .dout(n18222));
  jnot g00960(.din(n18179), .dout(n18223));
  jor  g00961(.dina(n18196), .dinb(n18223), .dout(n18224));
  jxor g00962(.dina(n18181), .dinb(n591), .dout(n18225));
  jand g00963(.dina(n18225), .dinb(n18196), .dout(n18226));
  jnot g00964(.din(n18226), .dout(n18227));
  jand g00965(.dina(n18227), .dinb(n18224), .dout(n18228));
  jnot g00966(.din(n18228), .dout(n18229));
  jand g00967(.dina(n18229), .dinb(n386), .dout(n18230));
  jand g00968(.dina(n18196), .dinb(b0 ), .dout(n18231));
  jxor g00969(.dina(n18231), .dinb(a58 ), .dout(n18232));
  jand g00970(.dina(n18232), .dinb(n259), .dout(n18233));
  jxor g00971(.dina(n18231), .dinb(n589), .dout(n18234));
  jxor g00972(.dina(n18234), .dinb(b1 ), .dout(n18235));
  jand g00973(.dina(n18235), .dinb(n650), .dout(n18236));
  jor  g00974(.dina(n18236), .dinb(n18233), .dout(n18237));
  jxor g00975(.dina(n18228), .dinb(b2 ), .dout(n18238));
  jand g00976(.dina(n18238), .dinb(n18237), .dout(n18239));
  jor  g00977(.dina(n18239), .dinb(n18230), .dout(n18240));
  jxor g00978(.dina(n18220), .dinb(b3 ), .dout(n18241));
  jand g00979(.dina(n18241), .dinb(n18240), .dout(n18242));
  jor  g00980(.dina(n18242), .dinb(n18222), .dout(n18243));
  jxor g00981(.dina(n18214), .dinb(n376), .dout(n18244));
  jand g00982(.dina(n18244), .dinb(n18243), .dout(n18245));
  jor  g00983(.dina(n18245), .dinb(n18215), .dout(n18246));
  jxor g00984(.dina(n18201), .dinb(n377), .dout(n18247));
  jand g00985(.dina(n18247), .dinb(n18246), .dout(n18248));
  jor  g00986(.dina(n18248), .dinb(n18210), .dout(n18249));
  jand g00987(.dina(n18249), .dinb(n18209), .dout(n18250));
  jor  g00988(.dina(n18250), .dinb(n18206), .dout(n18251));
  jand g00989(.dina(n18251), .dinb(n430), .dout(n18252));
  jor  g00990(.dina(n18252), .dinb(n18201), .dout(n18253));
  jnot g00991(.din(n18252), .dout(n18254));
  jxor g00992(.dina(n18247), .dinb(n18246), .dout(n18255));
  jor  g00993(.dina(n18255), .dinb(n18254), .dout(n18256));
  jand g00994(.dina(n18256), .dinb(n18253), .dout(n18257));
  jand g00995(.dina(n18254), .dinb(n18205), .dout(n18258));
  jand g00996(.dina(n18249), .dinb(n18206), .dout(n18259));
  jor  g00997(.dina(n18259), .dinb(n18258), .dout(n18260));
  jand g00998(.dina(n18260), .dinb(n265), .dout(n18261));
  jnot g00999(.din(n18260), .dout(n18262));
  jand g01000(.dina(n18262), .dinb(b7 ), .dout(n18263));
  jnot g01001(.din(n18263), .dout(n18264));
  jand g01002(.dina(n18257), .dinb(n378), .dout(n18265));
  jor  g01003(.dina(n18252), .dinb(n18214), .dout(n18266));
  jxor g01004(.dina(n18244), .dinb(n18243), .dout(n18267));
  jor  g01005(.dina(n18267), .dinb(n18254), .dout(n18268));
  jand g01006(.dina(n18268), .dinb(n18266), .dout(n18269));
  jand g01007(.dina(n18269), .dinb(n377), .dout(n18270));
  jand g01008(.dina(n18254), .dinb(n18220), .dout(n18271));
  jnot g01009(.din(n18271), .dout(n18272));
  jxor g01010(.dina(n18241), .dinb(n18240), .dout(n18273));
  jor  g01011(.dina(n18273), .dinb(n18254), .dout(n18274));
  jand g01012(.dina(n18274), .dinb(n18272), .dout(n18275));
  jand g01013(.dina(n18275), .dinb(n376), .dout(n18276));
  jor  g01014(.dina(n18252), .dinb(n18229), .dout(n18277));
  jxor g01015(.dina(n18238), .dinb(n18237), .dout(n18278));
  jor  g01016(.dina(n18278), .dinb(n18254), .dout(n18279));
  jand g01017(.dina(n18279), .dinb(n18277), .dout(n18280));
  jand g01018(.dina(n18280), .dinb(n264), .dout(n18281));
  jxor g01019(.dina(n18235), .dinb(n650), .dout(n18282));
  jand g01020(.dina(n18282), .dinb(n18252), .dout(n18283));
  jnot g01021(.din(n18283), .dout(n18284));
  jor  g01022(.dina(n18252), .dinb(n18234), .dout(n18285));
  jand g01023(.dina(n18285), .dinb(n18284), .dout(n18286));
  jor  g01024(.dina(n18286), .dinb(b2 ), .dout(n18287));
  jnot g01025(.din(n18287), .dout(n18288));
  jnot g01026(.din(n579), .dout(n18289));
  jnot g01027(.din(n18206), .dout(n18290));
  jnot g01028(.din(n18210), .dout(n18291));
  jnot g01029(.din(n18215), .dout(n18292));
  jnot g01030(.din(n18222), .dout(n18293));
  jnot g01031(.din(n18230), .dout(n18294));
  jnot g01032(.din(n18233), .dout(n18295));
  jxor g01033(.dina(n18234), .dinb(n259), .dout(n18296));
  jor  g01034(.dina(n18296), .dinb(n649), .dout(n18297));
  jand g01035(.dina(n18297), .dinb(n18295), .dout(n18298));
  jnot g01036(.din(n18238), .dout(n18299));
  jor  g01037(.dina(n18299), .dinb(n18298), .dout(n18300));
  jand g01038(.dina(n18300), .dinb(n18294), .dout(n18301));
  jnot g01039(.din(n18241), .dout(n18302));
  jor  g01040(.dina(n18302), .dinb(n18301), .dout(n18303));
  jand g01041(.dina(n18303), .dinb(n18293), .dout(n18304));
  jnot g01042(.din(n18244), .dout(n18305));
  jor  g01043(.dina(n18305), .dinb(n18304), .dout(n18306));
  jand g01044(.dina(n18306), .dinb(n18292), .dout(n18307));
  jnot g01045(.din(n18247), .dout(n18308));
  jor  g01046(.dina(n18308), .dinb(n18307), .dout(n18309));
  jand g01047(.dina(n18309), .dinb(n18291), .dout(n18310));
  jor  g01048(.dina(n18310), .dinb(n18208), .dout(n18311));
  jand g01049(.dina(n18311), .dinb(n18290), .dout(n18312));
  jor  g01050(.dina(n18312), .dinb(n18289), .dout(n18313));
  jand g01051(.dina(n18313), .dinb(a57 ), .dout(n18314));
  jnot g01052(.din(n708), .dout(n18315));
  jor  g01053(.dina(n18312), .dinb(n18315), .dout(n18316));
  jnot g01054(.din(n18316), .dout(n18317));
  jor  g01055(.dina(n18317), .dinb(n18314), .dout(n18318));
  jand g01056(.dina(n18318), .dinb(n259), .dout(n18319));
  jand g01057(.dina(n18251), .dinb(n579), .dout(n18320));
  jor  g01058(.dina(n18320), .dinb(n648), .dout(n18321));
  jand g01059(.dina(n18316), .dinb(n18321), .dout(n18322));
  jxor g01060(.dina(n18322), .dinb(b1 ), .dout(n18323));
  jand g01061(.dina(n18323), .dinb(n716), .dout(n18324));
  jor  g01062(.dina(n18324), .dinb(n18319), .dout(n18325));
  jxor g01063(.dina(n18286), .dinb(b2 ), .dout(n18326));
  jand g01064(.dina(n18326), .dinb(n18325), .dout(n18327));
  jor  g01065(.dina(n18327), .dinb(n18288), .dout(n18328));
  jxor g01066(.dina(n18280), .dinb(n264), .dout(n18329));
  jand g01067(.dina(n18329), .dinb(n18328), .dout(n18330));
  jor  g01068(.dina(n18330), .dinb(n18281), .dout(n18331));
  jxor g01069(.dina(n18275), .dinb(n376), .dout(n18332));
  jand g01070(.dina(n18332), .dinb(n18331), .dout(n18333));
  jor  g01071(.dina(n18333), .dinb(n18276), .dout(n18334));
  jxor g01072(.dina(n18269), .dinb(n377), .dout(n18335));
  jand g01073(.dina(n18335), .dinb(n18334), .dout(n18336));
  jor  g01074(.dina(n18336), .dinb(n18270), .dout(n18337));
  jxor g01075(.dina(n18257), .dinb(n378), .dout(n18338));
  jand g01076(.dina(n18338), .dinb(n18337), .dout(n18339));
  jor  g01077(.dina(n18339), .dinb(n18265), .dout(n18340));
  jand g01078(.dina(n18340), .dinb(n18264), .dout(n18341));
  jor  g01079(.dina(n18341), .dinb(n18261), .dout(n18342));
  jand g01080(.dina(n18342), .dinb(n374), .dout(n18343));
  jor  g01081(.dina(n18343), .dinb(n18257), .dout(n18344));
  jnot g01082(.din(n18343), .dout(n18345));
  jxor g01083(.dina(n18338), .dinb(n18337), .dout(n18346));
  jor  g01084(.dina(n18346), .dinb(n18345), .dout(n18347));
  jand g01085(.dina(n18347), .dinb(n18344), .dout(n18348));
  jand g01086(.dina(n18345), .dinb(n18260), .dout(n18349));
  jand g01087(.dina(n18340), .dinb(n18261), .dout(n18350));
  jor  g01088(.dina(n18350), .dinb(n18349), .dout(n18351));
  jand g01089(.dina(n18351), .dinb(n374), .dout(n18352));
  jand g01090(.dina(n18348), .dinb(n265), .dout(n18353));
  jxor g01091(.dina(n18335), .dinb(n18334), .dout(n18354));
  jand g01092(.dina(n18354), .dinb(n18343), .dout(n18355));
  jand g01093(.dina(n18345), .dinb(n18269), .dout(n18356));
  jor  g01094(.dina(n18356), .dinb(n18355), .dout(n18357));
  jand g01095(.dina(n18357), .dinb(n378), .dout(n18358));
  jor  g01096(.dina(n18343), .dinb(n18275), .dout(n18359));
  jxor g01097(.dina(n18332), .dinb(n18331), .dout(n18360));
  jor  g01098(.dina(n18360), .dinb(n18345), .dout(n18361));
  jand g01099(.dina(n18361), .dinb(n18359), .dout(n18362));
  jand g01100(.dina(n18362), .dinb(n377), .dout(n18363));
  jor  g01101(.dina(n18343), .dinb(n18280), .dout(n18364));
  jxor g01102(.dina(n18329), .dinb(n18328), .dout(n18365));
  jor  g01103(.dina(n18365), .dinb(n18345), .dout(n18366));
  jand g01104(.dina(n18366), .dinb(n18364), .dout(n18367));
  jand g01105(.dina(n18367), .dinb(n376), .dout(n18368));
  jxor g01106(.dina(n18326), .dinb(n18325), .dout(n18369));
  jnot g01107(.din(n18369), .dout(n18370));
  jor  g01108(.dina(n18370), .dinb(n18345), .dout(n18371));
  jor  g01109(.dina(n18343), .dinb(n18286), .dout(n18372));
  jand g01110(.dina(n18372), .dinb(n18371), .dout(n18373));
  jnot g01111(.din(n18373), .dout(n18374));
  jand g01112(.dina(n18374), .dinb(n264), .dout(n18375));
  jor  g01113(.dina(n18343), .dinb(n18322), .dout(n18376));
  jxor g01114(.dina(n18323), .dinb(n716), .dout(n18377));
  jand g01115(.dina(n18377), .dinb(n18343), .dout(n18378));
  jnot g01116(.din(n18378), .dout(n18379));
  jand g01117(.dina(n18379), .dinb(n18376), .dout(n18380));
  jnot g01118(.din(n18380), .dout(n18381));
  jand g01119(.dina(n18381), .dinb(n386), .dout(n18382));
  jnot g01120(.din(n777), .dout(n18383));
  jnot g01121(.din(n18261), .dout(n18384));
  jnot g01122(.din(n18265), .dout(n18385));
  jnot g01123(.din(n18270), .dout(n18386));
  jnot g01124(.din(n18276), .dout(n18387));
  jnot g01125(.din(n18281), .dout(n18388));
  jnot g01126(.din(n18319), .dout(n18389));
  jxor g01127(.dina(n18322), .dinb(n259), .dout(n18390));
  jor  g01128(.dina(n18390), .dinb(n715), .dout(n18391));
  jand g01129(.dina(n18391), .dinb(n18389), .dout(n18392));
  jnot g01130(.din(n18326), .dout(n18393));
  jor  g01131(.dina(n18393), .dinb(n18392), .dout(n18394));
  jand g01132(.dina(n18394), .dinb(n18287), .dout(n18395));
  jnot g01133(.din(n18329), .dout(n18396));
  jor  g01134(.dina(n18396), .dinb(n18395), .dout(n18397));
  jand g01135(.dina(n18397), .dinb(n18388), .dout(n18398));
  jnot g01136(.din(n18332), .dout(n18399));
  jor  g01137(.dina(n18399), .dinb(n18398), .dout(n18400));
  jand g01138(.dina(n18400), .dinb(n18387), .dout(n18401));
  jnot g01139(.din(n18335), .dout(n18402));
  jor  g01140(.dina(n18402), .dinb(n18401), .dout(n18403));
  jand g01141(.dina(n18403), .dinb(n18386), .dout(n18404));
  jnot g01142(.din(n18338), .dout(n18405));
  jor  g01143(.dina(n18405), .dinb(n18404), .dout(n18406));
  jand g01144(.dina(n18406), .dinb(n18385), .dout(n18407));
  jor  g01145(.dina(n18407), .dinb(n18263), .dout(n18408));
  jand g01146(.dina(n18408), .dinb(n18384), .dout(n18409));
  jor  g01147(.dina(n18409), .dinb(n18383), .dout(n18410));
  jand g01148(.dina(n18410), .dinb(a56 ), .dout(n18411));
  jnot g01149(.din(n780), .dout(n18412));
  jor  g01150(.dina(n18409), .dinb(n18412), .dout(n18413));
  jnot g01151(.din(n18413), .dout(n18414));
  jor  g01152(.dina(n18414), .dinb(n18411), .dout(n18415));
  jand g01153(.dina(n18415), .dinb(n259), .dout(n18416));
  jand g01154(.dina(n18342), .dinb(n777), .dout(n18417));
  jor  g01155(.dina(n18417), .dinb(n714), .dout(n18418));
  jand g01156(.dina(n18413), .dinb(n18418), .dout(n18419));
  jxor g01157(.dina(n18419), .dinb(b1 ), .dout(n18420));
  jand g01158(.dina(n18420), .dinb(n788), .dout(n18421));
  jor  g01159(.dina(n18421), .dinb(n18416), .dout(n18422));
  jxor g01160(.dina(n18380), .dinb(b2 ), .dout(n18423));
  jand g01161(.dina(n18423), .dinb(n18422), .dout(n18424));
  jor  g01162(.dina(n18424), .dinb(n18382), .dout(n18425));
  jxor g01163(.dina(n18373), .dinb(b3 ), .dout(n18426));
  jand g01164(.dina(n18426), .dinb(n18425), .dout(n18427));
  jor  g01165(.dina(n18427), .dinb(n18375), .dout(n18428));
  jxor g01166(.dina(n18367), .dinb(n376), .dout(n18429));
  jand g01167(.dina(n18429), .dinb(n18428), .dout(n18430));
  jor  g01168(.dina(n18430), .dinb(n18368), .dout(n18431));
  jxor g01169(.dina(n18362), .dinb(n377), .dout(n18432));
  jand g01170(.dina(n18432), .dinb(n18431), .dout(n18433));
  jor  g01171(.dina(n18433), .dinb(n18363), .dout(n18434));
  jxor g01172(.dina(n18357), .dinb(n378), .dout(n18435));
  jand g01173(.dina(n18435), .dinb(n18434), .dout(n18436));
  jor  g01174(.dina(n18436), .dinb(n18358), .dout(n18437));
  jxor g01175(.dina(n18348), .dinb(n265), .dout(n18438));
  jand g01176(.dina(n18438), .dinb(n18437), .dout(n18439));
  jor  g01177(.dina(n18439), .dinb(n18353), .dout(n18440));
  jxor g01178(.dina(n18351), .dinb(b8 ), .dout(n18441));
  jnot g01179(.din(n18441), .dout(n18442));
  jand g01180(.dina(n18442), .dinb(n18440), .dout(n18443));
  jand g01181(.dina(n18443), .dinb(n429), .dout(n18444));
  jor  g01182(.dina(n18444), .dinb(n18352), .dout(n18445));
  jor  g01183(.dina(n18445), .dinb(n18348), .dout(n18446));
  jnot g01184(.din(n18352), .dout(n18447));
  jnot g01185(.din(n429), .dout(n18448));
  jnot g01186(.din(n18353), .dout(n18449));
  jnot g01187(.din(n18358), .dout(n18450));
  jnot g01188(.din(n18363), .dout(n18451));
  jnot g01189(.din(n18368), .dout(n18452));
  jnot g01190(.din(n18375), .dout(n18453));
  jnot g01191(.din(n18382), .dout(n18454));
  jnot g01192(.din(n18416), .dout(n18455));
  jxor g01193(.dina(n18419), .dinb(n259), .dout(n18456));
  jor  g01194(.dina(n18456), .dinb(n787), .dout(n18457));
  jand g01195(.dina(n18457), .dinb(n18455), .dout(n18458));
  jnot g01196(.din(n18423), .dout(n18459));
  jor  g01197(.dina(n18459), .dinb(n18458), .dout(n18460));
  jand g01198(.dina(n18460), .dinb(n18454), .dout(n18461));
  jnot g01199(.din(n18426), .dout(n18462));
  jor  g01200(.dina(n18462), .dinb(n18461), .dout(n18463));
  jand g01201(.dina(n18463), .dinb(n18453), .dout(n18464));
  jnot g01202(.din(n18429), .dout(n18465));
  jor  g01203(.dina(n18465), .dinb(n18464), .dout(n18466));
  jand g01204(.dina(n18466), .dinb(n18452), .dout(n18467));
  jnot g01205(.din(n18432), .dout(n18468));
  jor  g01206(.dina(n18468), .dinb(n18467), .dout(n18469));
  jand g01207(.dina(n18469), .dinb(n18451), .dout(n18470));
  jnot g01208(.din(n18435), .dout(n18471));
  jor  g01209(.dina(n18471), .dinb(n18470), .dout(n18472));
  jand g01210(.dina(n18472), .dinb(n18450), .dout(n18473));
  jnot g01211(.din(n18438), .dout(n18474));
  jor  g01212(.dina(n18474), .dinb(n18473), .dout(n18475));
  jand g01213(.dina(n18475), .dinb(n18449), .dout(n18476));
  jor  g01214(.dina(n18441), .dinb(n18476), .dout(n18477));
  jor  g01215(.dina(n18477), .dinb(n18448), .dout(n18478));
  jand g01216(.dina(n18478), .dinb(n18447), .dout(n18479));
  jxor g01217(.dina(n18438), .dinb(n18437), .dout(n18480));
  jor  g01218(.dina(n18480), .dinb(n18479), .dout(n18481));
  jand g01219(.dina(n18481), .dinb(n18446), .dout(n18482));
  jxor g01220(.dina(n18441), .dinb(n18476), .dout(n18483));
  jor  g01221(.dina(n18483), .dinb(n18479), .dout(n18484));
  jor  g01222(.dina(n18444), .dinb(n18351), .dout(n18485));
  jand g01223(.dina(n18485), .dinb(n18484), .dout(n18486));
  jand g01224(.dina(n18486), .dinb(n368), .dout(n18487));
  jnot g01225(.din(n18486), .dout(n18488));
  jand g01226(.dina(n18488), .dinb(b9 ), .dout(n18489));
  jnot g01227(.din(n18489), .dout(n18490));
  jand g01228(.dina(n18482), .dinb(n367), .dout(n18491));
  jor  g01229(.dina(n18445), .dinb(n18357), .dout(n18492));
  jxor g01230(.dina(n18435), .dinb(n18434), .dout(n18493));
  jor  g01231(.dina(n18493), .dinb(n18479), .dout(n18494));
  jand g01232(.dina(n18494), .dinb(n18492), .dout(n18495));
  jand g01233(.dina(n18495), .dinb(n265), .dout(n18496));
  jor  g01234(.dina(n18445), .dinb(n18362), .dout(n18497));
  jxor g01235(.dina(n18432), .dinb(n18431), .dout(n18498));
  jor  g01236(.dina(n18498), .dinb(n18479), .dout(n18499));
  jand g01237(.dina(n18499), .dinb(n18497), .dout(n18500));
  jand g01238(.dina(n18500), .dinb(n378), .dout(n18501));
  jor  g01239(.dina(n18445), .dinb(n18367), .dout(n18502));
  jxor g01240(.dina(n18429), .dinb(n18428), .dout(n18503));
  jor  g01241(.dina(n18503), .dinb(n18479), .dout(n18504));
  jand g01242(.dina(n18504), .dinb(n18502), .dout(n18505));
  jand g01243(.dina(n18505), .dinb(n377), .dout(n18506));
  jand g01244(.dina(n18479), .dinb(n18373), .dout(n18507));
  jnot g01245(.din(n18507), .dout(n18508));
  jxor g01246(.dina(n18426), .dinb(n18425), .dout(n18509));
  jor  g01247(.dina(n18509), .dinb(n18479), .dout(n18510));
  jand g01248(.dina(n18510), .dinb(n18508), .dout(n18511));
  jand g01249(.dina(n18511), .dinb(n376), .dout(n18512));
  jor  g01250(.dina(n18445), .dinb(n18381), .dout(n18513));
  jxor g01251(.dina(n18423), .dinb(n18422), .dout(n18514));
  jor  g01252(.dina(n18514), .dinb(n18479), .dout(n18515));
  jand g01253(.dina(n18515), .dinb(n18513), .dout(n18516));
  jand g01254(.dina(n18516), .dinb(n264), .dout(n18517));
  jand g01255(.dina(n18456), .dinb(n787), .dout(n18518));
  jor  g01256(.dina(n18479), .dinb(n18421), .dout(n18519));
  jor  g01257(.dina(n18519), .dinb(n18518), .dout(n18520));
  jand g01258(.dina(n18479), .dinb(n18415), .dout(n18521));
  jnot g01259(.din(n18521), .dout(n18522));
  jand g01260(.dina(n18522), .dinb(n18520), .dout(n18523));
  jnot g01261(.din(n18523), .dout(n18524));
  jand g01262(.dina(n18524), .dinb(n386), .dout(n18525));
  jand g01263(.dina(n18445), .dinb(b0 ), .dout(n18526));
  jxor g01264(.dina(n18526), .dinb(a55 ), .dout(n18527));
  jand g01265(.dina(n18527), .dinb(n259), .dout(n18528));
  jxor g01266(.dina(n18526), .dinb(n786), .dout(n18529));
  jxor g01267(.dina(n18529), .dinb(b1 ), .dout(n18530));
  jand g01268(.dina(n18530), .dinb(n916), .dout(n18531));
  jor  g01269(.dina(n18531), .dinb(n18528), .dout(n18532));
  jxor g01270(.dina(n18523), .dinb(b2 ), .dout(n18533));
  jand g01271(.dina(n18533), .dinb(n18532), .dout(n18534));
  jor  g01272(.dina(n18534), .dinb(n18525), .dout(n18535));
  jxor g01273(.dina(n18516), .dinb(n264), .dout(n18536));
  jand g01274(.dina(n18536), .dinb(n18535), .dout(n18537));
  jor  g01275(.dina(n18537), .dinb(n18517), .dout(n18538));
  jxor g01276(.dina(n18511), .dinb(n376), .dout(n18539));
  jand g01277(.dina(n18539), .dinb(n18538), .dout(n18540));
  jor  g01278(.dina(n18540), .dinb(n18512), .dout(n18541));
  jxor g01279(.dina(n18505), .dinb(n377), .dout(n18542));
  jand g01280(.dina(n18542), .dinb(n18541), .dout(n18543));
  jor  g01281(.dina(n18543), .dinb(n18506), .dout(n18544));
  jxor g01282(.dina(n18500), .dinb(n378), .dout(n18545));
  jand g01283(.dina(n18545), .dinb(n18544), .dout(n18546));
  jor  g01284(.dina(n18546), .dinb(n18501), .dout(n18547));
  jxor g01285(.dina(n18495), .dinb(n265), .dout(n18548));
  jand g01286(.dina(n18548), .dinb(n18547), .dout(n18549));
  jor  g01287(.dina(n18549), .dinb(n18496), .dout(n18550));
  jxor g01288(.dina(n18482), .dinb(n367), .dout(n18551));
  jand g01289(.dina(n18551), .dinb(n18550), .dout(n18552));
  jor  g01290(.dina(n18552), .dinb(n18491), .dout(n18553));
  jand g01291(.dina(n18553), .dinb(n18490), .dout(n18554));
  jor  g01292(.dina(n18554), .dinb(n18487), .dout(n18555));
  jand g01293(.dina(n18555), .dinb(n998), .dout(n18556));
  jor  g01294(.dina(n18556), .dinb(n18482), .dout(n18557));
  jnot g01295(.din(n18556), .dout(n18558));
  jxor g01296(.dina(n18551), .dinb(n18550), .dout(n18559));
  jor  g01297(.dina(n18559), .dinb(n18558), .dout(n18560));
  jand g01298(.dina(n18560), .dinb(n18557), .dout(n18561));
  jand g01299(.dina(n18558), .dinb(n18486), .dout(n18562));
  jand g01300(.dina(n18553), .dinb(n18487), .dout(n18563));
  jor  g01301(.dina(n18563), .dinb(n18562), .dout(n18564));
  jand g01302(.dina(n18564), .dinb(n369), .dout(n18565));
  jnot g01303(.din(n18564), .dout(n18566));
  jand g01304(.dina(n18566), .dinb(b10 ), .dout(n18567));
  jnot g01305(.din(n18567), .dout(n18568));
  jand g01306(.dina(n18561), .dinb(n368), .dout(n18569));
  jor  g01307(.dina(n18556), .dinb(n18495), .dout(n18570));
  jxor g01308(.dina(n18548), .dinb(n18547), .dout(n18571));
  jor  g01309(.dina(n18571), .dinb(n18558), .dout(n18572));
  jand g01310(.dina(n18572), .dinb(n18570), .dout(n18573));
  jand g01311(.dina(n18573), .dinb(n367), .dout(n18574));
  jor  g01312(.dina(n18556), .dinb(n18500), .dout(n18575));
  jxor g01313(.dina(n18545), .dinb(n18544), .dout(n18576));
  jor  g01314(.dina(n18576), .dinb(n18558), .dout(n18577));
  jand g01315(.dina(n18577), .dinb(n18575), .dout(n18578));
  jand g01316(.dina(n18578), .dinb(n265), .dout(n18579));
  jor  g01317(.dina(n18556), .dinb(n18505), .dout(n18580));
  jxor g01318(.dina(n18542), .dinb(n18541), .dout(n18581));
  jor  g01319(.dina(n18581), .dinb(n18558), .dout(n18582));
  jand g01320(.dina(n18582), .dinb(n18580), .dout(n18583));
  jand g01321(.dina(n18583), .dinb(n378), .dout(n18584));
  jor  g01322(.dina(n18556), .dinb(n18511), .dout(n18585));
  jxor g01323(.dina(n18539), .dinb(n18538), .dout(n18586));
  jor  g01324(.dina(n18586), .dinb(n18558), .dout(n18587));
  jand g01325(.dina(n18587), .dinb(n18585), .dout(n18588));
  jand g01326(.dina(n18588), .dinb(n377), .dout(n18589));
  jor  g01327(.dina(n18556), .dinb(n18516), .dout(n18590));
  jxor g01328(.dina(n18536), .dinb(n18535), .dout(n18591));
  jor  g01329(.dina(n18591), .dinb(n18558), .dout(n18592));
  jand g01330(.dina(n18592), .dinb(n18590), .dout(n18593));
  jand g01331(.dina(n18593), .dinb(n376), .dout(n18594));
  jor  g01332(.dina(n18556), .dinb(n18524), .dout(n18595));
  jxor g01333(.dina(n18533), .dinb(n18532), .dout(n18596));
  jor  g01334(.dina(n18596), .dinb(n18558), .dout(n18597));
  jand g01335(.dina(n18597), .dinb(n18595), .dout(n18598));
  jand g01336(.dina(n18598), .dinb(n264), .dout(n18599));
  jor  g01337(.dina(n18556), .dinb(n18529), .dout(n18600));
  jxor g01338(.dina(n18530), .dinb(n916), .dout(n18601));
  jand g01339(.dina(n18601), .dinb(n18556), .dout(n18602));
  jnot g01340(.din(n18602), .dout(n18603));
  jand g01341(.dina(n18603), .dinb(n18600), .dout(n18604));
  jor  g01342(.dina(n18604), .dinb(b2 ), .dout(n18605));
  jnot g01343(.din(n18605), .dout(n18606));
  jnot g01344(.din(n999), .dout(n18607));
  jnot g01345(.din(n18487), .dout(n18608));
  jnot g01346(.din(n18491), .dout(n18609));
  jnot g01347(.din(n18496), .dout(n18610));
  jnot g01348(.din(n18501), .dout(n18611));
  jnot g01349(.din(n18506), .dout(n18612));
  jnot g01350(.din(n18512), .dout(n18613));
  jnot g01351(.din(n18517), .dout(n18614));
  jnot g01352(.din(n18525), .dout(n18615));
  jnot g01353(.din(n18528), .dout(n18616));
  jxor g01354(.dina(n18529), .dinb(n259), .dout(n18617));
  jor  g01355(.dina(n18617), .dinb(n915), .dout(n18618));
  jand g01356(.dina(n18618), .dinb(n18616), .dout(n18619));
  jnot g01357(.din(n18533), .dout(n18620));
  jor  g01358(.dina(n18620), .dinb(n18619), .dout(n18621));
  jand g01359(.dina(n18621), .dinb(n18615), .dout(n18622));
  jnot g01360(.din(n18536), .dout(n18623));
  jor  g01361(.dina(n18623), .dinb(n18622), .dout(n18624));
  jand g01362(.dina(n18624), .dinb(n18614), .dout(n18625));
  jnot g01363(.din(n18539), .dout(n18626));
  jor  g01364(.dina(n18626), .dinb(n18625), .dout(n18627));
  jand g01365(.dina(n18627), .dinb(n18613), .dout(n18628));
  jnot g01366(.din(n18542), .dout(n18629));
  jor  g01367(.dina(n18629), .dinb(n18628), .dout(n18630));
  jand g01368(.dina(n18630), .dinb(n18612), .dout(n18631));
  jnot g01369(.din(n18545), .dout(n18632));
  jor  g01370(.dina(n18632), .dinb(n18631), .dout(n18633));
  jand g01371(.dina(n18633), .dinb(n18611), .dout(n18634));
  jnot g01372(.din(n18548), .dout(n18635));
  jor  g01373(.dina(n18635), .dinb(n18634), .dout(n18636));
  jand g01374(.dina(n18636), .dinb(n18610), .dout(n18637));
  jnot g01375(.din(n18551), .dout(n18638));
  jor  g01376(.dina(n18638), .dinb(n18637), .dout(n18639));
  jand g01377(.dina(n18639), .dinb(n18609), .dout(n18640));
  jor  g01378(.dina(n18640), .dinb(n18489), .dout(n18641));
  jand g01379(.dina(n18641), .dinb(n18608), .dout(n18642));
  jor  g01380(.dina(n18642), .dinb(n18607), .dout(n18643));
  jand g01381(.dina(n18643), .dinb(a54 ), .dout(n18644));
  jnot g01382(.din(n1002), .dout(n18645));
  jor  g01383(.dina(n18642), .dinb(n18645), .dout(n18646));
  jnot g01384(.din(n18646), .dout(n18647));
  jor  g01385(.dina(n18647), .dinb(n18644), .dout(n18648));
  jand g01386(.dina(n18648), .dinb(n259), .dout(n18649));
  jand g01387(.dina(n18555), .dinb(n999), .dout(n18650));
  jor  g01388(.dina(n18650), .dinb(n914), .dout(n18651));
  jand g01389(.dina(n18646), .dinb(n18651), .dout(n18652));
  jxor g01390(.dina(n18652), .dinb(b1 ), .dout(n18653));
  jand g01391(.dina(n18653), .dinb(n1010), .dout(n18654));
  jor  g01392(.dina(n18654), .dinb(n18649), .dout(n18655));
  jxor g01393(.dina(n18604), .dinb(b2 ), .dout(n18656));
  jand g01394(.dina(n18656), .dinb(n18655), .dout(n18657));
  jor  g01395(.dina(n18657), .dinb(n18606), .dout(n18658));
  jxor g01396(.dina(n18598), .dinb(n264), .dout(n18659));
  jand g01397(.dina(n18659), .dinb(n18658), .dout(n18660));
  jor  g01398(.dina(n18660), .dinb(n18599), .dout(n18661));
  jxor g01399(.dina(n18593), .dinb(n376), .dout(n18662));
  jand g01400(.dina(n18662), .dinb(n18661), .dout(n18663));
  jor  g01401(.dina(n18663), .dinb(n18594), .dout(n18664));
  jxor g01402(.dina(n18588), .dinb(n377), .dout(n18665));
  jand g01403(.dina(n18665), .dinb(n18664), .dout(n18666));
  jor  g01404(.dina(n18666), .dinb(n18589), .dout(n18667));
  jxor g01405(.dina(n18583), .dinb(n378), .dout(n18668));
  jand g01406(.dina(n18668), .dinb(n18667), .dout(n18669));
  jor  g01407(.dina(n18669), .dinb(n18584), .dout(n18670));
  jxor g01408(.dina(n18578), .dinb(n265), .dout(n18671));
  jand g01409(.dina(n18671), .dinb(n18670), .dout(n18672));
  jor  g01410(.dina(n18672), .dinb(n18579), .dout(n18673));
  jxor g01411(.dina(n18573), .dinb(n367), .dout(n18674));
  jand g01412(.dina(n18674), .dinb(n18673), .dout(n18675));
  jor  g01413(.dina(n18675), .dinb(n18574), .dout(n18676));
  jxor g01414(.dina(n18561), .dinb(n368), .dout(n18677));
  jand g01415(.dina(n18677), .dinb(n18676), .dout(n18678));
  jor  g01416(.dina(n18678), .dinb(n18569), .dout(n18679));
  jand g01417(.dina(n18679), .dinb(n18568), .dout(n18680));
  jor  g01418(.dina(n18680), .dinb(n18565), .dout(n18681));
  jand g01419(.dina(n18681), .dinb(n952), .dout(n18682));
  jor  g01420(.dina(n18682), .dinb(n18561), .dout(n18683));
  jnot g01421(.din(n952), .dout(n18684));
  jnot g01422(.din(n18565), .dout(n18685));
  jnot g01423(.din(n18569), .dout(n18686));
  jnot g01424(.din(n18574), .dout(n18687));
  jnot g01425(.din(n18579), .dout(n18688));
  jnot g01426(.din(n18584), .dout(n18689));
  jnot g01427(.din(n18589), .dout(n18690));
  jnot g01428(.din(n18594), .dout(n18691));
  jnot g01429(.din(n18599), .dout(n18692));
  jor  g01430(.dina(n18652), .dinb(b1 ), .dout(n18693));
  jxor g01431(.dina(n18652), .dinb(n259), .dout(n18694));
  jor  g01432(.dina(n18694), .dinb(n1009), .dout(n18695));
  jand g01433(.dina(n18695), .dinb(n18693), .dout(n18696));
  jxor g01434(.dina(n18604), .dinb(n386), .dout(n18697));
  jor  g01435(.dina(n18697), .dinb(n18696), .dout(n18698));
  jand g01436(.dina(n18698), .dinb(n18605), .dout(n18699));
  jnot g01437(.din(n18659), .dout(n18700));
  jor  g01438(.dina(n18700), .dinb(n18699), .dout(n18701));
  jand g01439(.dina(n18701), .dinb(n18692), .dout(n18702));
  jnot g01440(.din(n18662), .dout(n18703));
  jor  g01441(.dina(n18703), .dinb(n18702), .dout(n18704));
  jand g01442(.dina(n18704), .dinb(n18691), .dout(n18705));
  jnot g01443(.din(n18665), .dout(n18706));
  jor  g01444(.dina(n18706), .dinb(n18705), .dout(n18707));
  jand g01445(.dina(n18707), .dinb(n18690), .dout(n18708));
  jnot g01446(.din(n18668), .dout(n18709));
  jor  g01447(.dina(n18709), .dinb(n18708), .dout(n18710));
  jand g01448(.dina(n18710), .dinb(n18689), .dout(n18711));
  jnot g01449(.din(n18671), .dout(n18712));
  jor  g01450(.dina(n18712), .dinb(n18711), .dout(n18713));
  jand g01451(.dina(n18713), .dinb(n18688), .dout(n18714));
  jnot g01452(.din(n18674), .dout(n18715));
  jor  g01453(.dina(n18715), .dinb(n18714), .dout(n18716));
  jand g01454(.dina(n18716), .dinb(n18687), .dout(n18717));
  jnot g01455(.din(n18677), .dout(n18718));
  jor  g01456(.dina(n18718), .dinb(n18717), .dout(n18719));
  jand g01457(.dina(n18719), .dinb(n18686), .dout(n18720));
  jor  g01458(.dina(n18720), .dinb(n18567), .dout(n18721));
  jand g01459(.dina(n18721), .dinb(n18685), .dout(n18722));
  jor  g01460(.dina(n18722), .dinb(n18684), .dout(n18723));
  jxor g01461(.dina(n18677), .dinb(n18676), .dout(n18724));
  jor  g01462(.dina(n18724), .dinb(n18723), .dout(n18725));
  jand g01463(.dina(n18725), .dinb(n18683), .dout(n18726));
  jand g01464(.dina(n18679), .dinb(n998), .dout(n18727));
  jor  g01465(.dina(n18727), .dinb(n18723), .dout(n18728));
  jand g01466(.dina(n18728), .dinb(n18564), .dout(n18729));
  jand g01467(.dina(n18729), .dinb(n952), .dout(n18730));
  jand g01468(.dina(n18726), .dinb(n369), .dout(n18731));
  jor  g01469(.dina(n18682), .dinb(n18573), .dout(n18732));
  jxor g01470(.dina(n18674), .dinb(n18673), .dout(n18733));
  jor  g01471(.dina(n18733), .dinb(n18723), .dout(n18734));
  jand g01472(.dina(n18734), .dinb(n18732), .dout(n18735));
  jand g01473(.dina(n18735), .dinb(n368), .dout(n18736));
  jor  g01474(.dina(n18682), .dinb(n18578), .dout(n18737));
  jxor g01475(.dina(n18671), .dinb(n18670), .dout(n18738));
  jor  g01476(.dina(n18738), .dinb(n18723), .dout(n18739));
  jand g01477(.dina(n18739), .dinb(n18737), .dout(n18740));
  jand g01478(.dina(n18740), .dinb(n367), .dout(n18741));
  jor  g01479(.dina(n18682), .dinb(n18583), .dout(n18742));
  jxor g01480(.dina(n18668), .dinb(n18667), .dout(n18743));
  jor  g01481(.dina(n18743), .dinb(n18723), .dout(n18744));
  jand g01482(.dina(n18744), .dinb(n18742), .dout(n18745));
  jand g01483(.dina(n18745), .dinb(n265), .dout(n18746));
  jor  g01484(.dina(n18682), .dinb(n18588), .dout(n18747));
  jxor g01485(.dina(n18665), .dinb(n18664), .dout(n18748));
  jor  g01486(.dina(n18748), .dinb(n18723), .dout(n18749));
  jand g01487(.dina(n18749), .dinb(n18747), .dout(n18750));
  jand g01488(.dina(n18750), .dinb(n378), .dout(n18751));
  jor  g01489(.dina(n18682), .dinb(n18593), .dout(n18752));
  jxor g01490(.dina(n18662), .dinb(n18661), .dout(n18753));
  jor  g01491(.dina(n18753), .dinb(n18723), .dout(n18754));
  jand g01492(.dina(n18754), .dinb(n18752), .dout(n18755));
  jand g01493(.dina(n18755), .dinb(n377), .dout(n18756));
  jor  g01494(.dina(n18682), .dinb(n18598), .dout(n18757));
  jxor g01495(.dina(n18659), .dinb(n18658), .dout(n18758));
  jor  g01496(.dina(n18758), .dinb(n18723), .dout(n18759));
  jand g01497(.dina(n18759), .dinb(n18757), .dout(n18760));
  jand g01498(.dina(n18760), .dinb(n376), .dout(n18761));
  jnot g01499(.din(n18604), .dout(n18762));
  jor  g01500(.dina(n18682), .dinb(n18762), .dout(n18763));
  jxor g01501(.dina(n18656), .dinb(n18655), .dout(n18764));
  jor  g01502(.dina(n18764), .dinb(n18723), .dout(n18765));
  jand g01503(.dina(n18765), .dinb(n18763), .dout(n18766));
  jand g01504(.dina(n18766), .dinb(n264), .dout(n18767));
  jand g01505(.dina(n18723), .dinb(n18648), .dout(n18768));
  jxor g01506(.dina(n18653), .dinb(n1010), .dout(n18769));
  jand g01507(.dina(n18769), .dinb(n18682), .dout(n18770));
  jor  g01508(.dina(n18770), .dinb(n18768), .dout(n18771));
  jand g01509(.dina(n18771), .dinb(n386), .dout(n18772));
  jnot g01510(.din(n1096), .dout(n18773));
  jor  g01511(.dina(n18722), .dinb(n18773), .dout(n18774));
  jand g01512(.dina(n18774), .dinb(a53 ), .dout(n18775));
  jand g01513(.dina(n18682), .dinb(n1009), .dout(n18776));
  jor  g01514(.dina(n18776), .dinb(n18775), .dout(n18777));
  jand g01515(.dina(n18777), .dinb(n259), .dout(n18778));
  jand g01516(.dina(n18681), .dinb(n1096), .dout(n18779));
  jor  g01517(.dina(n18779), .dinb(n1008), .dout(n18780));
  jor  g01518(.dina(n18723), .dinb(n1010), .dout(n18781));
  jand g01519(.dina(n18781), .dinb(n18780), .dout(n18782));
  jxor g01520(.dina(n18782), .dinb(b1 ), .dout(n18783));
  jand g01521(.dina(n18783), .dinb(n1106), .dout(n18784));
  jor  g01522(.dina(n18784), .dinb(n18778), .dout(n18785));
  jxor g01523(.dina(n18771), .dinb(n386), .dout(n18786));
  jand g01524(.dina(n18786), .dinb(n18785), .dout(n18787));
  jor  g01525(.dina(n18787), .dinb(n18772), .dout(n18788));
  jxor g01526(.dina(n18766), .dinb(n264), .dout(n18789));
  jand g01527(.dina(n18789), .dinb(n18788), .dout(n18790));
  jor  g01528(.dina(n18790), .dinb(n18767), .dout(n18791));
  jxor g01529(.dina(n18760), .dinb(n376), .dout(n18792));
  jand g01530(.dina(n18792), .dinb(n18791), .dout(n18793));
  jor  g01531(.dina(n18793), .dinb(n18761), .dout(n18794));
  jxor g01532(.dina(n18755), .dinb(n377), .dout(n18795));
  jand g01533(.dina(n18795), .dinb(n18794), .dout(n18796));
  jor  g01534(.dina(n18796), .dinb(n18756), .dout(n18797));
  jxor g01535(.dina(n18750), .dinb(n378), .dout(n18798));
  jand g01536(.dina(n18798), .dinb(n18797), .dout(n18799));
  jor  g01537(.dina(n18799), .dinb(n18751), .dout(n18800));
  jxor g01538(.dina(n18745), .dinb(n265), .dout(n18801));
  jand g01539(.dina(n18801), .dinb(n18800), .dout(n18802));
  jor  g01540(.dina(n18802), .dinb(n18746), .dout(n18803));
  jxor g01541(.dina(n18740), .dinb(n367), .dout(n18804));
  jand g01542(.dina(n18804), .dinb(n18803), .dout(n18805));
  jor  g01543(.dina(n18805), .dinb(n18741), .dout(n18806));
  jxor g01544(.dina(n18735), .dinb(n368), .dout(n18807));
  jand g01545(.dina(n18807), .dinb(n18806), .dout(n18808));
  jor  g01546(.dina(n18808), .dinb(n18736), .dout(n18809));
  jxor g01547(.dina(n18726), .dinb(n369), .dout(n18810));
  jand g01548(.dina(n18810), .dinb(n18809), .dout(n18811));
  jor  g01549(.dina(n18811), .dinb(n18731), .dout(n18812));
  jxor g01550(.dina(n18729), .dinb(b11 ), .dout(n18813));
  jnot g01551(.din(n18813), .dout(n18814));
  jand g01552(.dina(n18814), .dinb(n18812), .dout(n18815));
  jand g01553(.dina(n18815), .dinb(n951), .dout(n18816));
  jor  g01554(.dina(n18816), .dinb(n18730), .dout(n18817));
  jor  g01555(.dina(n18817), .dinb(n18726), .dout(n18818));
  jnot g01556(.din(n18817), .dout(n18819));
  jxor g01557(.dina(n18810), .dinb(n18809), .dout(n18820));
  jor  g01558(.dina(n18820), .dinb(n18819), .dout(n18821));
  jand g01559(.dina(n18821), .dinb(n18818), .dout(n18822));
  jxor g01560(.dina(n18814), .dinb(n18812), .dout(n18823));
  jand g01561(.dina(n18823), .dinb(n18730), .dout(n18824));
  jand g01562(.dina(n18819), .dinb(n18729), .dout(n18825));
  jor  g01563(.dina(n18825), .dinb(n18824), .dout(n18826));
  jand g01564(.dina(n18826), .dinb(n363), .dout(n18827));
  jnot g01565(.din(n18826), .dout(n18828));
  jand g01566(.dina(n18828), .dinb(b12 ), .dout(n18829));
  jnot g01567(.din(n18829), .dout(n18830));
  jand g01568(.dina(n18822), .dinb(n359), .dout(n18831));
  jor  g01569(.dina(n18817), .dinb(n18735), .dout(n18832));
  jxor g01570(.dina(n18807), .dinb(n18806), .dout(n18833));
  jor  g01571(.dina(n18833), .dinb(n18819), .dout(n18834));
  jand g01572(.dina(n18834), .dinb(n18832), .dout(n18835));
  jand g01573(.dina(n18835), .dinb(n369), .dout(n18836));
  jor  g01574(.dina(n18817), .dinb(n18740), .dout(n18837));
  jxor g01575(.dina(n18804), .dinb(n18803), .dout(n18838));
  jor  g01576(.dina(n18838), .dinb(n18819), .dout(n18839));
  jand g01577(.dina(n18839), .dinb(n18837), .dout(n18840));
  jand g01578(.dina(n18840), .dinb(n368), .dout(n18841));
  jor  g01579(.dina(n18817), .dinb(n18745), .dout(n18842));
  jxor g01580(.dina(n18801), .dinb(n18800), .dout(n18843));
  jor  g01581(.dina(n18843), .dinb(n18819), .dout(n18844));
  jand g01582(.dina(n18844), .dinb(n18842), .dout(n18845));
  jand g01583(.dina(n18845), .dinb(n367), .dout(n18846));
  jor  g01584(.dina(n18817), .dinb(n18750), .dout(n18847));
  jxor g01585(.dina(n18798), .dinb(n18797), .dout(n18848));
  jor  g01586(.dina(n18848), .dinb(n18819), .dout(n18849));
  jand g01587(.dina(n18849), .dinb(n18847), .dout(n18850));
  jand g01588(.dina(n18850), .dinb(n265), .dout(n18851));
  jor  g01589(.dina(n18817), .dinb(n18755), .dout(n18852));
  jxor g01590(.dina(n18795), .dinb(n18794), .dout(n18853));
  jor  g01591(.dina(n18853), .dinb(n18819), .dout(n18854));
  jand g01592(.dina(n18854), .dinb(n18852), .dout(n18855));
  jand g01593(.dina(n18855), .dinb(n378), .dout(n18856));
  jor  g01594(.dina(n18817), .dinb(n18760), .dout(n18857));
  jxor g01595(.dina(n18792), .dinb(n18791), .dout(n18858));
  jor  g01596(.dina(n18858), .dinb(n18819), .dout(n18859));
  jand g01597(.dina(n18859), .dinb(n18857), .dout(n18860));
  jand g01598(.dina(n18860), .dinb(n377), .dout(n18861));
  jor  g01599(.dina(n18817), .dinb(n18766), .dout(n18862));
  jxor g01600(.dina(n18789), .dinb(n18788), .dout(n18863));
  jor  g01601(.dina(n18863), .dinb(n18819), .dout(n18864));
  jand g01602(.dina(n18864), .dinb(n18862), .dout(n18865));
  jand g01603(.dina(n18865), .dinb(n376), .dout(n18866));
  jor  g01604(.dina(n18817), .dinb(n18771), .dout(n18867));
  jxor g01605(.dina(n18786), .dinb(n18785), .dout(n18868));
  jor  g01606(.dina(n18868), .dinb(n18819), .dout(n18869));
  jand g01607(.dina(n18869), .dinb(n18867), .dout(n18870));
  jand g01608(.dina(n18870), .dinb(n264), .dout(n18871));
  jor  g01609(.dina(n18817), .dinb(n18777), .dout(n18872));
  jxor g01610(.dina(n18783), .dinb(n1106), .dout(n18873));
  jor  g01611(.dina(n18873), .dinb(n18819), .dout(n18874));
  jand g01612(.dina(n18874), .dinb(n18872), .dout(n18875));
  jand g01613(.dina(n18875), .dinb(n386), .dout(n18876));
  jand g01614(.dina(n18817), .dinb(b0 ), .dout(n18877));
  jxor g01615(.dina(n18877), .dinb(a52 ), .dout(n18878));
  jand g01616(.dina(n18878), .dinb(n259), .dout(n18879));
  jxor g01617(.dina(n18877), .dinb(n1104), .dout(n18880));
  jxor g01618(.dina(n18880), .dinb(b1 ), .dout(n18881));
  jand g01619(.dina(n18881), .dinb(n1209), .dout(n18882));
  jor  g01620(.dina(n18882), .dinb(n18879), .dout(n18883));
  jxor g01621(.dina(n18875), .dinb(n386), .dout(n18884));
  jand g01622(.dina(n18884), .dinb(n18883), .dout(n18885));
  jor  g01623(.dina(n18885), .dinb(n18876), .dout(n18886));
  jxor g01624(.dina(n18870), .dinb(n264), .dout(n18887));
  jand g01625(.dina(n18887), .dinb(n18886), .dout(n18888));
  jor  g01626(.dina(n18888), .dinb(n18871), .dout(n18889));
  jxor g01627(.dina(n18865), .dinb(n376), .dout(n18890));
  jand g01628(.dina(n18890), .dinb(n18889), .dout(n18891));
  jor  g01629(.dina(n18891), .dinb(n18866), .dout(n18892));
  jxor g01630(.dina(n18860), .dinb(n377), .dout(n18893));
  jand g01631(.dina(n18893), .dinb(n18892), .dout(n18894));
  jor  g01632(.dina(n18894), .dinb(n18861), .dout(n18895));
  jxor g01633(.dina(n18855), .dinb(n378), .dout(n18896));
  jand g01634(.dina(n18896), .dinb(n18895), .dout(n18897));
  jor  g01635(.dina(n18897), .dinb(n18856), .dout(n18898));
  jxor g01636(.dina(n18850), .dinb(n265), .dout(n18899));
  jand g01637(.dina(n18899), .dinb(n18898), .dout(n18900));
  jor  g01638(.dina(n18900), .dinb(n18851), .dout(n18901));
  jxor g01639(.dina(n18845), .dinb(n367), .dout(n18902));
  jand g01640(.dina(n18902), .dinb(n18901), .dout(n18903));
  jor  g01641(.dina(n18903), .dinb(n18846), .dout(n18904));
  jxor g01642(.dina(n18840), .dinb(n368), .dout(n18905));
  jand g01643(.dina(n18905), .dinb(n18904), .dout(n18906));
  jor  g01644(.dina(n18906), .dinb(n18841), .dout(n18907));
  jxor g01645(.dina(n18835), .dinb(n369), .dout(n18908));
  jand g01646(.dina(n18908), .dinb(n18907), .dout(n18909));
  jor  g01647(.dina(n18909), .dinb(n18836), .dout(n18910));
  jxor g01648(.dina(n18822), .dinb(n359), .dout(n18911));
  jand g01649(.dina(n18911), .dinb(n18910), .dout(n18912));
  jor  g01650(.dina(n18912), .dinb(n18831), .dout(n18913));
  jand g01651(.dina(n18913), .dinb(n18830), .dout(n18914));
  jor  g01652(.dina(n18914), .dinb(n18827), .dout(n18915));
  jand g01653(.dina(n18915), .dinb(n425), .dout(n18916));
  jor  g01654(.dina(n18916), .dinb(n18822), .dout(n18917));
  jnot g01655(.din(n18916), .dout(n18918));
  jxor g01656(.dina(n18911), .dinb(n18910), .dout(n18919));
  jor  g01657(.dina(n18919), .dinb(n18918), .dout(n18920));
  jand g01658(.dina(n18920), .dinb(n18917), .dout(n18921));
  jand g01659(.dina(n18918), .dinb(n18826), .dout(n18922));
  jand g01660(.dina(n18913), .dinb(n18827), .dout(n18923));
  jor  g01661(.dina(n18923), .dinb(n18922), .dout(n18924));
  jand g01662(.dina(n18924), .dinb(n360), .dout(n18925));
  jnot g01663(.din(n18924), .dout(n18926));
  jand g01664(.dina(n18926), .dinb(b13 ), .dout(n18927));
  jnot g01665(.din(n18927), .dout(n18928));
  jand g01666(.dina(n18921), .dinb(n363), .dout(n18929));
  jor  g01667(.dina(n18916), .dinb(n18835), .dout(n18930));
  jxor g01668(.dina(n18908), .dinb(n18907), .dout(n18931));
  jor  g01669(.dina(n18931), .dinb(n18918), .dout(n18932));
  jand g01670(.dina(n18932), .dinb(n18930), .dout(n18933));
  jand g01671(.dina(n18933), .dinb(n359), .dout(n18934));
  jor  g01672(.dina(n18916), .dinb(n18840), .dout(n18935));
  jxor g01673(.dina(n18905), .dinb(n18904), .dout(n18936));
  jor  g01674(.dina(n18936), .dinb(n18918), .dout(n18937));
  jand g01675(.dina(n18937), .dinb(n18935), .dout(n18938));
  jand g01676(.dina(n18938), .dinb(n369), .dout(n18939));
  jor  g01677(.dina(n18916), .dinb(n18845), .dout(n18940));
  jxor g01678(.dina(n18902), .dinb(n18901), .dout(n18941));
  jor  g01679(.dina(n18941), .dinb(n18918), .dout(n18942));
  jand g01680(.dina(n18942), .dinb(n18940), .dout(n18943));
  jand g01681(.dina(n18943), .dinb(n368), .dout(n18944));
  jor  g01682(.dina(n18916), .dinb(n18850), .dout(n18945));
  jxor g01683(.dina(n18899), .dinb(n18898), .dout(n18946));
  jor  g01684(.dina(n18946), .dinb(n18918), .dout(n18947));
  jand g01685(.dina(n18947), .dinb(n18945), .dout(n18948));
  jand g01686(.dina(n18948), .dinb(n367), .dout(n18949));
  jor  g01687(.dina(n18916), .dinb(n18855), .dout(n18950));
  jxor g01688(.dina(n18896), .dinb(n18895), .dout(n18951));
  jor  g01689(.dina(n18951), .dinb(n18918), .dout(n18952));
  jand g01690(.dina(n18952), .dinb(n18950), .dout(n18953));
  jand g01691(.dina(n18953), .dinb(n265), .dout(n18954));
  jor  g01692(.dina(n18916), .dinb(n18860), .dout(n18955));
  jxor g01693(.dina(n18893), .dinb(n18892), .dout(n18956));
  jor  g01694(.dina(n18956), .dinb(n18918), .dout(n18957));
  jand g01695(.dina(n18957), .dinb(n18955), .dout(n18958));
  jand g01696(.dina(n18958), .dinb(n378), .dout(n18959));
  jor  g01697(.dina(n18916), .dinb(n18865), .dout(n18960));
  jxor g01698(.dina(n18890), .dinb(n18889), .dout(n18961));
  jor  g01699(.dina(n18961), .dinb(n18918), .dout(n18962));
  jand g01700(.dina(n18962), .dinb(n18960), .dout(n18963));
  jand g01701(.dina(n18963), .dinb(n377), .dout(n18964));
  jor  g01702(.dina(n18916), .dinb(n18870), .dout(n18965));
  jxor g01703(.dina(n18887), .dinb(n18886), .dout(n18966));
  jor  g01704(.dina(n18966), .dinb(n18918), .dout(n18967));
  jand g01705(.dina(n18967), .dinb(n18965), .dout(n18968));
  jand g01706(.dina(n18968), .dinb(n376), .dout(n18969));
  jor  g01707(.dina(n18916), .dinb(n18875), .dout(n18970));
  jxor g01708(.dina(n18884), .dinb(n18883), .dout(n18971));
  jor  g01709(.dina(n18971), .dinb(n18918), .dout(n18972));
  jand g01710(.dina(n18972), .dinb(n18970), .dout(n18973));
  jand g01711(.dina(n18973), .dinb(n264), .dout(n18974));
  jor  g01712(.dina(n18916), .dinb(n18880), .dout(n18975));
  jxor g01713(.dina(n18881), .dinb(n1209), .dout(n18976));
  jand g01714(.dina(n18976), .dinb(n18916), .dout(n18977));
  jnot g01715(.din(n18977), .dout(n18978));
  jand g01716(.dina(n18978), .dinb(n18975), .dout(n18979));
  jor  g01717(.dina(n18979), .dinb(b2 ), .dout(n18980));
  jnot g01718(.din(n18980), .dout(n18981));
  jnot g01719(.din(n1314), .dout(n18982));
  jnot g01720(.din(n18827), .dout(n18983));
  jnot g01721(.din(n18831), .dout(n18984));
  jnot g01722(.din(n18836), .dout(n18985));
  jnot g01723(.din(n18841), .dout(n18986));
  jnot g01724(.din(n18846), .dout(n18987));
  jnot g01725(.din(n18851), .dout(n18988));
  jnot g01726(.din(n18856), .dout(n18989));
  jnot g01727(.din(n18861), .dout(n18990));
  jnot g01728(.din(n18866), .dout(n18991));
  jnot g01729(.din(n18871), .dout(n18992));
  jnot g01730(.din(n18876), .dout(n18993));
  jnot g01731(.din(n18879), .dout(n18994));
  jxor g01732(.dina(n18880), .dinb(n259), .dout(n18995));
  jor  g01733(.dina(n18995), .dinb(n1208), .dout(n18996));
  jand g01734(.dina(n18996), .dinb(n18994), .dout(n18997));
  jnot g01735(.din(n18884), .dout(n18998));
  jor  g01736(.dina(n18998), .dinb(n18997), .dout(n18999));
  jand g01737(.dina(n18999), .dinb(n18993), .dout(n19000));
  jnot g01738(.din(n18887), .dout(n19001));
  jor  g01739(.dina(n19001), .dinb(n19000), .dout(n19002));
  jand g01740(.dina(n19002), .dinb(n18992), .dout(n19003));
  jnot g01741(.din(n18890), .dout(n19004));
  jor  g01742(.dina(n19004), .dinb(n19003), .dout(n19005));
  jand g01743(.dina(n19005), .dinb(n18991), .dout(n19006));
  jnot g01744(.din(n18893), .dout(n19007));
  jor  g01745(.dina(n19007), .dinb(n19006), .dout(n19008));
  jand g01746(.dina(n19008), .dinb(n18990), .dout(n19009));
  jnot g01747(.din(n18896), .dout(n19010));
  jor  g01748(.dina(n19010), .dinb(n19009), .dout(n19011));
  jand g01749(.dina(n19011), .dinb(n18989), .dout(n19012));
  jnot g01750(.din(n18899), .dout(n19013));
  jor  g01751(.dina(n19013), .dinb(n19012), .dout(n19014));
  jand g01752(.dina(n19014), .dinb(n18988), .dout(n19015));
  jnot g01753(.din(n18902), .dout(n19016));
  jor  g01754(.dina(n19016), .dinb(n19015), .dout(n19017));
  jand g01755(.dina(n19017), .dinb(n18987), .dout(n19018));
  jnot g01756(.din(n18905), .dout(n19019));
  jor  g01757(.dina(n19019), .dinb(n19018), .dout(n19020));
  jand g01758(.dina(n19020), .dinb(n18986), .dout(n19021));
  jnot g01759(.din(n18908), .dout(n19022));
  jor  g01760(.dina(n19022), .dinb(n19021), .dout(n19023));
  jand g01761(.dina(n19023), .dinb(n18985), .dout(n19024));
  jnot g01762(.din(n18911), .dout(n19025));
  jor  g01763(.dina(n19025), .dinb(n19024), .dout(n19026));
  jand g01764(.dina(n19026), .dinb(n18984), .dout(n19027));
  jor  g01765(.dina(n19027), .dinb(n18829), .dout(n19028));
  jand g01766(.dina(n19028), .dinb(n18983), .dout(n19029));
  jor  g01767(.dina(n19029), .dinb(n18982), .dout(n19030));
  jand g01768(.dina(n19030), .dinb(a51 ), .dout(n19031));
  jnot g01769(.din(n1317), .dout(n19032));
  jor  g01770(.dina(n19029), .dinb(n19032), .dout(n19033));
  jnot g01771(.din(n19033), .dout(n19034));
  jor  g01772(.dina(n19034), .dinb(n19031), .dout(n19035));
  jand g01773(.dina(n19035), .dinb(n259), .dout(n19036));
  jand g01774(.dina(n18915), .dinb(n1314), .dout(n19037));
  jor  g01775(.dina(n19037), .dinb(n1207), .dout(n19038));
  jand g01776(.dina(n19033), .dinb(n19038), .dout(n19039));
  jxor g01777(.dina(n19039), .dinb(b1 ), .dout(n19040));
  jand g01778(.dina(n19040), .dinb(n1325), .dout(n19041));
  jor  g01779(.dina(n19041), .dinb(n19036), .dout(n19042));
  jxor g01780(.dina(n18979), .dinb(b2 ), .dout(n19043));
  jand g01781(.dina(n19043), .dinb(n19042), .dout(n19044));
  jor  g01782(.dina(n19044), .dinb(n18981), .dout(n19045));
  jxor g01783(.dina(n18973), .dinb(n264), .dout(n19046));
  jand g01784(.dina(n19046), .dinb(n19045), .dout(n19047));
  jor  g01785(.dina(n19047), .dinb(n18974), .dout(n19048));
  jxor g01786(.dina(n18968), .dinb(n376), .dout(n19049));
  jand g01787(.dina(n19049), .dinb(n19048), .dout(n19050));
  jor  g01788(.dina(n19050), .dinb(n18969), .dout(n19051));
  jxor g01789(.dina(n18963), .dinb(n377), .dout(n19052));
  jand g01790(.dina(n19052), .dinb(n19051), .dout(n19053));
  jor  g01791(.dina(n19053), .dinb(n18964), .dout(n19054));
  jxor g01792(.dina(n18958), .dinb(n378), .dout(n19055));
  jand g01793(.dina(n19055), .dinb(n19054), .dout(n19056));
  jor  g01794(.dina(n19056), .dinb(n18959), .dout(n19057));
  jxor g01795(.dina(n18953), .dinb(n265), .dout(n19058));
  jand g01796(.dina(n19058), .dinb(n19057), .dout(n19059));
  jor  g01797(.dina(n19059), .dinb(n18954), .dout(n19060));
  jxor g01798(.dina(n18948), .dinb(n367), .dout(n19061));
  jand g01799(.dina(n19061), .dinb(n19060), .dout(n19062));
  jor  g01800(.dina(n19062), .dinb(n18949), .dout(n19063));
  jxor g01801(.dina(n18943), .dinb(n368), .dout(n19064));
  jand g01802(.dina(n19064), .dinb(n19063), .dout(n19065));
  jor  g01803(.dina(n19065), .dinb(n18944), .dout(n19066));
  jxor g01804(.dina(n18938), .dinb(n369), .dout(n19067));
  jand g01805(.dina(n19067), .dinb(n19066), .dout(n19068));
  jor  g01806(.dina(n19068), .dinb(n18939), .dout(n19069));
  jxor g01807(.dina(n18933), .dinb(n359), .dout(n19070));
  jand g01808(.dina(n19070), .dinb(n19069), .dout(n19071));
  jor  g01809(.dina(n19071), .dinb(n18934), .dout(n19072));
  jxor g01810(.dina(n18921), .dinb(n363), .dout(n19073));
  jand g01811(.dina(n19073), .dinb(n19072), .dout(n19074));
  jor  g01812(.dina(n19074), .dinb(n18929), .dout(n19075));
  jand g01813(.dina(n19075), .dinb(n18928), .dout(n19076));
  jor  g01814(.dina(n19076), .dinb(n18925), .dout(n19077));
  jand g01815(.dina(n19077), .dinb(n1254), .dout(n19078));
  jor  g01816(.dina(n19078), .dinb(n18921), .dout(n19079));
  jnot g01817(.din(n1254), .dout(n19080));
  jnot g01818(.din(n18925), .dout(n19081));
  jnot g01819(.din(n18929), .dout(n19082));
  jnot g01820(.din(n18934), .dout(n19083));
  jnot g01821(.din(n18939), .dout(n19084));
  jnot g01822(.din(n18944), .dout(n19085));
  jnot g01823(.din(n18949), .dout(n19086));
  jnot g01824(.din(n18954), .dout(n19087));
  jnot g01825(.din(n18959), .dout(n19088));
  jnot g01826(.din(n18964), .dout(n19089));
  jnot g01827(.din(n18969), .dout(n19090));
  jnot g01828(.din(n18974), .dout(n19091));
  jor  g01829(.dina(n19039), .dinb(b1 ), .dout(n19092));
  jxor g01830(.dina(n19039), .dinb(n259), .dout(n19093));
  jor  g01831(.dina(n19093), .dinb(n1324), .dout(n19094));
  jand g01832(.dina(n19094), .dinb(n19092), .dout(n19095));
  jxor g01833(.dina(n18979), .dinb(n386), .dout(n19096));
  jor  g01834(.dina(n19096), .dinb(n19095), .dout(n19097));
  jand g01835(.dina(n19097), .dinb(n18980), .dout(n19098));
  jnot g01836(.din(n19046), .dout(n19099));
  jor  g01837(.dina(n19099), .dinb(n19098), .dout(n19100));
  jand g01838(.dina(n19100), .dinb(n19091), .dout(n19101));
  jnot g01839(.din(n19049), .dout(n19102));
  jor  g01840(.dina(n19102), .dinb(n19101), .dout(n19103));
  jand g01841(.dina(n19103), .dinb(n19090), .dout(n19104));
  jnot g01842(.din(n19052), .dout(n19105));
  jor  g01843(.dina(n19105), .dinb(n19104), .dout(n19106));
  jand g01844(.dina(n19106), .dinb(n19089), .dout(n19107));
  jnot g01845(.din(n19055), .dout(n19108));
  jor  g01846(.dina(n19108), .dinb(n19107), .dout(n19109));
  jand g01847(.dina(n19109), .dinb(n19088), .dout(n19110));
  jnot g01848(.din(n19058), .dout(n19111));
  jor  g01849(.dina(n19111), .dinb(n19110), .dout(n19112));
  jand g01850(.dina(n19112), .dinb(n19087), .dout(n19113));
  jnot g01851(.din(n19061), .dout(n19114));
  jor  g01852(.dina(n19114), .dinb(n19113), .dout(n19115));
  jand g01853(.dina(n19115), .dinb(n19086), .dout(n19116));
  jnot g01854(.din(n19064), .dout(n19117));
  jor  g01855(.dina(n19117), .dinb(n19116), .dout(n19118));
  jand g01856(.dina(n19118), .dinb(n19085), .dout(n19119));
  jnot g01857(.din(n19067), .dout(n19120));
  jor  g01858(.dina(n19120), .dinb(n19119), .dout(n19121));
  jand g01859(.dina(n19121), .dinb(n19084), .dout(n19122));
  jnot g01860(.din(n19070), .dout(n19123));
  jor  g01861(.dina(n19123), .dinb(n19122), .dout(n19124));
  jand g01862(.dina(n19124), .dinb(n19083), .dout(n19125));
  jnot g01863(.din(n19073), .dout(n19126));
  jor  g01864(.dina(n19126), .dinb(n19125), .dout(n19127));
  jand g01865(.dina(n19127), .dinb(n19082), .dout(n19128));
  jor  g01866(.dina(n19128), .dinb(n18927), .dout(n19129));
  jand g01867(.dina(n19129), .dinb(n19081), .dout(n19130));
  jor  g01868(.dina(n19130), .dinb(n19080), .dout(n19131));
  jxor g01869(.dina(n19073), .dinb(n19072), .dout(n19132));
  jor  g01870(.dina(n19132), .dinb(n19131), .dout(n19133));
  jand g01871(.dina(n19133), .dinb(n19079), .dout(n19134));
  jand g01872(.dina(n19134), .dinb(n360), .dout(n19135));
  jor  g01873(.dina(n19078), .dinb(n18933), .dout(n19136));
  jxor g01874(.dina(n19070), .dinb(n19069), .dout(n19137));
  jor  g01875(.dina(n19137), .dinb(n19131), .dout(n19138));
  jand g01876(.dina(n19138), .dinb(n19136), .dout(n19139));
  jand g01877(.dina(n19139), .dinb(n363), .dout(n19140));
  jor  g01878(.dina(n19078), .dinb(n18938), .dout(n19141));
  jxor g01879(.dina(n19067), .dinb(n19066), .dout(n19142));
  jor  g01880(.dina(n19142), .dinb(n19131), .dout(n19143));
  jand g01881(.dina(n19143), .dinb(n19141), .dout(n19144));
  jand g01882(.dina(n19144), .dinb(n359), .dout(n19145));
  jor  g01883(.dina(n19078), .dinb(n18943), .dout(n19146));
  jxor g01884(.dina(n19064), .dinb(n19063), .dout(n19147));
  jor  g01885(.dina(n19147), .dinb(n19131), .dout(n19148));
  jand g01886(.dina(n19148), .dinb(n19146), .dout(n19149));
  jand g01887(.dina(n19149), .dinb(n369), .dout(n19150));
  jor  g01888(.dina(n19078), .dinb(n18948), .dout(n19151));
  jxor g01889(.dina(n19061), .dinb(n19060), .dout(n19152));
  jor  g01890(.dina(n19152), .dinb(n19131), .dout(n19153));
  jand g01891(.dina(n19153), .dinb(n19151), .dout(n19154));
  jand g01892(.dina(n19154), .dinb(n368), .dout(n19155));
  jor  g01893(.dina(n19078), .dinb(n18953), .dout(n19156));
  jxor g01894(.dina(n19058), .dinb(n19057), .dout(n19157));
  jor  g01895(.dina(n19157), .dinb(n19131), .dout(n19158));
  jand g01896(.dina(n19158), .dinb(n19156), .dout(n19159));
  jand g01897(.dina(n19159), .dinb(n367), .dout(n19160));
  jor  g01898(.dina(n19078), .dinb(n18958), .dout(n19161));
  jxor g01899(.dina(n19055), .dinb(n19054), .dout(n19162));
  jor  g01900(.dina(n19162), .dinb(n19131), .dout(n19163));
  jand g01901(.dina(n19163), .dinb(n19161), .dout(n19164));
  jand g01902(.dina(n19164), .dinb(n265), .dout(n19165));
  jor  g01903(.dina(n19078), .dinb(n18963), .dout(n19166));
  jxor g01904(.dina(n19052), .dinb(n19051), .dout(n19167));
  jor  g01905(.dina(n19167), .dinb(n19131), .dout(n19168));
  jand g01906(.dina(n19168), .dinb(n19166), .dout(n19169));
  jand g01907(.dina(n19169), .dinb(n378), .dout(n19170));
  jor  g01908(.dina(n19078), .dinb(n18968), .dout(n19171));
  jxor g01909(.dina(n19049), .dinb(n19048), .dout(n19172));
  jor  g01910(.dina(n19172), .dinb(n19131), .dout(n19173));
  jand g01911(.dina(n19173), .dinb(n19171), .dout(n19174));
  jand g01912(.dina(n19174), .dinb(n377), .dout(n19175));
  jor  g01913(.dina(n19078), .dinb(n18973), .dout(n19176));
  jxor g01914(.dina(n19046), .dinb(n19045), .dout(n19177));
  jor  g01915(.dina(n19177), .dinb(n19131), .dout(n19178));
  jand g01916(.dina(n19178), .dinb(n19176), .dout(n19179));
  jand g01917(.dina(n19179), .dinb(n376), .dout(n19180));
  jnot g01918(.din(n18979), .dout(n19181));
  jor  g01919(.dina(n19078), .dinb(n19181), .dout(n19182));
  jxor g01920(.dina(n19043), .dinb(n19042), .dout(n19183));
  jor  g01921(.dina(n19183), .dinb(n19131), .dout(n19184));
  jand g01922(.dina(n19184), .dinb(n19182), .dout(n19185));
  jand g01923(.dina(n19185), .dinb(n264), .dout(n19186));
  jand g01924(.dina(n19131), .dinb(n19035), .dout(n19187));
  jxor g01925(.dina(n19040), .dinb(n1325), .dout(n19188));
  jand g01926(.dina(n19188), .dinb(n19078), .dout(n19189));
  jor  g01927(.dina(n19189), .dinb(n19187), .dout(n19190));
  jand g01928(.dina(n19190), .dinb(n386), .dout(n19191));
  jnot g01929(.din(n1431), .dout(n19192));
  jor  g01930(.dina(n19130), .dinb(n19192), .dout(n19193));
  jand g01931(.dina(n19193), .dinb(a50 ), .dout(n19194));
  jand g01932(.dina(n19078), .dinb(n1324), .dout(n19195));
  jor  g01933(.dina(n19195), .dinb(n19194), .dout(n19196));
  jand g01934(.dina(n19196), .dinb(n259), .dout(n19197));
  jand g01935(.dina(n19077), .dinb(n1431), .dout(n19198));
  jor  g01936(.dina(n19198), .dinb(n1323), .dout(n19199));
  jor  g01937(.dina(n19131), .dinb(n1325), .dout(n19200));
  jand g01938(.dina(n19200), .dinb(n19199), .dout(n19201));
  jxor g01939(.dina(n19201), .dinb(b1 ), .dout(n19202));
  jand g01940(.dina(n19202), .dinb(n1441), .dout(n19203));
  jor  g01941(.dina(n19203), .dinb(n19197), .dout(n19204));
  jxor g01942(.dina(n19190), .dinb(n386), .dout(n19205));
  jand g01943(.dina(n19205), .dinb(n19204), .dout(n19206));
  jor  g01944(.dina(n19206), .dinb(n19191), .dout(n19207));
  jxor g01945(.dina(n19185), .dinb(n264), .dout(n19208));
  jand g01946(.dina(n19208), .dinb(n19207), .dout(n19209));
  jor  g01947(.dina(n19209), .dinb(n19186), .dout(n19210));
  jxor g01948(.dina(n19179), .dinb(n376), .dout(n19211));
  jand g01949(.dina(n19211), .dinb(n19210), .dout(n19212));
  jor  g01950(.dina(n19212), .dinb(n19180), .dout(n19213));
  jxor g01951(.dina(n19174), .dinb(n377), .dout(n19214));
  jand g01952(.dina(n19214), .dinb(n19213), .dout(n19215));
  jor  g01953(.dina(n19215), .dinb(n19175), .dout(n19216));
  jxor g01954(.dina(n19169), .dinb(n378), .dout(n19217));
  jand g01955(.dina(n19217), .dinb(n19216), .dout(n19218));
  jor  g01956(.dina(n19218), .dinb(n19170), .dout(n19219));
  jxor g01957(.dina(n19164), .dinb(n265), .dout(n19220));
  jand g01958(.dina(n19220), .dinb(n19219), .dout(n19221));
  jor  g01959(.dina(n19221), .dinb(n19165), .dout(n19222));
  jxor g01960(.dina(n19159), .dinb(n367), .dout(n19223));
  jand g01961(.dina(n19223), .dinb(n19222), .dout(n19224));
  jor  g01962(.dina(n19224), .dinb(n19160), .dout(n19225));
  jxor g01963(.dina(n19154), .dinb(n368), .dout(n19226));
  jand g01964(.dina(n19226), .dinb(n19225), .dout(n19227));
  jor  g01965(.dina(n19227), .dinb(n19155), .dout(n19228));
  jxor g01966(.dina(n19149), .dinb(n369), .dout(n19229));
  jand g01967(.dina(n19229), .dinb(n19228), .dout(n19230));
  jor  g01968(.dina(n19230), .dinb(n19150), .dout(n19231));
  jxor g01969(.dina(n19144), .dinb(n359), .dout(n19232));
  jand g01970(.dina(n19232), .dinb(n19231), .dout(n19233));
  jor  g01971(.dina(n19233), .dinb(n19145), .dout(n19234));
  jxor g01972(.dina(n19139), .dinb(n363), .dout(n19235));
  jand g01973(.dina(n19235), .dinb(n19234), .dout(n19236));
  jor  g01974(.dina(n19236), .dinb(n19140), .dout(n19237));
  jxor g01975(.dina(n19134), .dinb(n360), .dout(n19238));
  jand g01976(.dina(n19238), .dinb(n19237), .dout(n19239));
  jor  g01977(.dina(n19239), .dinb(n19135), .dout(n19240));
  jand g01978(.dina(n19131), .dinb(n18924), .dout(n19241));
  jand g01979(.dina(n19075), .dinb(n18925), .dout(n19242));
  jor  g01980(.dina(n19242), .dinb(n19241), .dout(n19243));
  jxor g01981(.dina(n19243), .dinb(b14 ), .dout(n19244));
  jnot g01982(.din(n19244), .dout(n19245));
  jand g01983(.dina(n19245), .dinb(n19240), .dout(n19246));
  jand g01984(.dina(n19246), .dinb(n424), .dout(n19247));
  jand g01985(.dina(n19243), .dinb(n1254), .dout(n19248));
  jor  g01986(.dina(n19248), .dinb(n19247), .dout(n19249));
  jor  g01987(.dina(n19249), .dinb(n19134), .dout(n19250));
  jnot g01988(.din(n19249), .dout(n19251));
  jxor g01989(.dina(n19238), .dinb(n19237), .dout(n19252));
  jor  g01990(.dina(n19252), .dinb(n19251), .dout(n19253));
  jand g01991(.dina(n19253), .dinb(n19250), .dout(n19254));
  jxor g01992(.dina(n19245), .dinb(n19240), .dout(n19255));
  jor  g01993(.dina(n19255), .dinb(n19251), .dout(n19256));
  jor  g01994(.dina(n19247), .dinb(n19243), .dout(n19257));
  jand g01995(.dina(n19257), .dinb(n19256), .dout(n19258));
  jand g01996(.dina(n19258), .dinb(n364), .dout(n19259));
  jnot g01997(.din(n19258), .dout(n19260));
  jand g01998(.dina(n19260), .dinb(b15 ), .dout(n19261));
  jnot g01999(.din(n19261), .dout(n19262));
  jand g02000(.dina(n19254), .dinb(n361), .dout(n19263));
  jor  g02001(.dina(n19249), .dinb(n19139), .dout(n19264));
  jxor g02002(.dina(n19235), .dinb(n19234), .dout(n19265));
  jor  g02003(.dina(n19265), .dinb(n19251), .dout(n19266));
  jand g02004(.dina(n19266), .dinb(n19264), .dout(n19267));
  jand g02005(.dina(n19267), .dinb(n360), .dout(n19268));
  jor  g02006(.dina(n19249), .dinb(n19144), .dout(n19269));
  jxor g02007(.dina(n19232), .dinb(n19231), .dout(n19270));
  jor  g02008(.dina(n19270), .dinb(n19251), .dout(n19271));
  jand g02009(.dina(n19271), .dinb(n19269), .dout(n19272));
  jand g02010(.dina(n19272), .dinb(n363), .dout(n19273));
  jor  g02011(.dina(n19249), .dinb(n19149), .dout(n19274));
  jxor g02012(.dina(n19229), .dinb(n19228), .dout(n19275));
  jor  g02013(.dina(n19275), .dinb(n19251), .dout(n19276));
  jand g02014(.dina(n19276), .dinb(n19274), .dout(n19277));
  jand g02015(.dina(n19277), .dinb(n359), .dout(n19278));
  jor  g02016(.dina(n19249), .dinb(n19154), .dout(n19279));
  jxor g02017(.dina(n19226), .dinb(n19225), .dout(n19280));
  jor  g02018(.dina(n19280), .dinb(n19251), .dout(n19281));
  jand g02019(.dina(n19281), .dinb(n19279), .dout(n19282));
  jand g02020(.dina(n19282), .dinb(n369), .dout(n19283));
  jor  g02021(.dina(n19249), .dinb(n19159), .dout(n19284));
  jxor g02022(.dina(n19223), .dinb(n19222), .dout(n19285));
  jor  g02023(.dina(n19285), .dinb(n19251), .dout(n19286));
  jand g02024(.dina(n19286), .dinb(n19284), .dout(n19287));
  jand g02025(.dina(n19287), .dinb(n368), .dout(n19288));
  jor  g02026(.dina(n19249), .dinb(n19164), .dout(n19289));
  jxor g02027(.dina(n19220), .dinb(n19219), .dout(n19290));
  jor  g02028(.dina(n19290), .dinb(n19251), .dout(n19291));
  jand g02029(.dina(n19291), .dinb(n19289), .dout(n19292));
  jand g02030(.dina(n19292), .dinb(n367), .dout(n19293));
  jor  g02031(.dina(n19249), .dinb(n19169), .dout(n19294));
  jxor g02032(.dina(n19217), .dinb(n19216), .dout(n19295));
  jor  g02033(.dina(n19295), .dinb(n19251), .dout(n19296));
  jand g02034(.dina(n19296), .dinb(n19294), .dout(n19297));
  jand g02035(.dina(n19297), .dinb(n265), .dout(n19298));
  jor  g02036(.dina(n19249), .dinb(n19174), .dout(n19299));
  jxor g02037(.dina(n19214), .dinb(n19213), .dout(n19300));
  jor  g02038(.dina(n19300), .dinb(n19251), .dout(n19301));
  jand g02039(.dina(n19301), .dinb(n19299), .dout(n19302));
  jand g02040(.dina(n19302), .dinb(n378), .dout(n19303));
  jor  g02041(.dina(n19249), .dinb(n19179), .dout(n19304));
  jxor g02042(.dina(n19211), .dinb(n19210), .dout(n19305));
  jor  g02043(.dina(n19305), .dinb(n19251), .dout(n19306));
  jand g02044(.dina(n19306), .dinb(n19304), .dout(n19307));
  jand g02045(.dina(n19307), .dinb(n377), .dout(n19308));
  jor  g02046(.dina(n19249), .dinb(n19185), .dout(n19309));
  jxor g02047(.dina(n19208), .dinb(n19207), .dout(n19310));
  jor  g02048(.dina(n19310), .dinb(n19251), .dout(n19311));
  jand g02049(.dina(n19311), .dinb(n19309), .dout(n19312));
  jand g02050(.dina(n19312), .dinb(n376), .dout(n19313));
  jor  g02051(.dina(n19249), .dinb(n19190), .dout(n19314));
  jxor g02052(.dina(n19205), .dinb(n19204), .dout(n19315));
  jor  g02053(.dina(n19315), .dinb(n19251), .dout(n19316));
  jand g02054(.dina(n19316), .dinb(n19314), .dout(n19317));
  jand g02055(.dina(n19317), .dinb(n264), .dout(n19318));
  jor  g02056(.dina(n19249), .dinb(n19201), .dout(n19319));
  jxor g02057(.dina(n19202), .dinb(n1441), .dout(n19320));
  jand g02058(.dina(n19320), .dinb(n19249), .dout(n19321));
  jnot g02059(.din(n19321), .dout(n19322));
  jand g02060(.dina(n19322), .dinb(n19319), .dout(n19323));
  jnot g02061(.din(n19323), .dout(n19324));
  jand g02062(.dina(n19324), .dinb(n386), .dout(n19325));
  jand g02063(.dina(n19249), .dinb(b0 ), .dout(n19326));
  jxor g02064(.dina(n19326), .dinb(a49 ), .dout(n19327));
  jand g02065(.dina(n19327), .dinb(n259), .dout(n19328));
  jxor g02066(.dina(n19326), .dinb(n1439), .dout(n19329));
  jxor g02067(.dina(n19329), .dinb(b1 ), .dout(n19330));
  jand g02068(.dina(n19330), .dinb(n1571), .dout(n19331));
  jor  g02069(.dina(n19331), .dinb(n19328), .dout(n19332));
  jxor g02070(.dina(n19323), .dinb(b2 ), .dout(n19333));
  jand g02071(.dina(n19333), .dinb(n19332), .dout(n19334));
  jor  g02072(.dina(n19334), .dinb(n19325), .dout(n19335));
  jxor g02073(.dina(n19317), .dinb(n264), .dout(n19336));
  jand g02074(.dina(n19336), .dinb(n19335), .dout(n19337));
  jor  g02075(.dina(n19337), .dinb(n19318), .dout(n19338));
  jxor g02076(.dina(n19312), .dinb(n376), .dout(n19339));
  jand g02077(.dina(n19339), .dinb(n19338), .dout(n19340));
  jor  g02078(.dina(n19340), .dinb(n19313), .dout(n19341));
  jxor g02079(.dina(n19307), .dinb(n377), .dout(n19342));
  jand g02080(.dina(n19342), .dinb(n19341), .dout(n19343));
  jor  g02081(.dina(n19343), .dinb(n19308), .dout(n19344));
  jxor g02082(.dina(n19302), .dinb(n378), .dout(n19345));
  jand g02083(.dina(n19345), .dinb(n19344), .dout(n19346));
  jor  g02084(.dina(n19346), .dinb(n19303), .dout(n19347));
  jxor g02085(.dina(n19297), .dinb(n265), .dout(n19348));
  jand g02086(.dina(n19348), .dinb(n19347), .dout(n19349));
  jor  g02087(.dina(n19349), .dinb(n19298), .dout(n19350));
  jxor g02088(.dina(n19292), .dinb(n367), .dout(n19351));
  jand g02089(.dina(n19351), .dinb(n19350), .dout(n19352));
  jor  g02090(.dina(n19352), .dinb(n19293), .dout(n19353));
  jxor g02091(.dina(n19287), .dinb(n368), .dout(n19354));
  jand g02092(.dina(n19354), .dinb(n19353), .dout(n19355));
  jor  g02093(.dina(n19355), .dinb(n19288), .dout(n19356));
  jxor g02094(.dina(n19282), .dinb(n369), .dout(n19357));
  jand g02095(.dina(n19357), .dinb(n19356), .dout(n19358));
  jor  g02096(.dina(n19358), .dinb(n19283), .dout(n19359));
  jxor g02097(.dina(n19277), .dinb(n359), .dout(n19360));
  jand g02098(.dina(n19360), .dinb(n19359), .dout(n19361));
  jor  g02099(.dina(n19361), .dinb(n19278), .dout(n19362));
  jxor g02100(.dina(n19272), .dinb(n363), .dout(n19363));
  jand g02101(.dina(n19363), .dinb(n19362), .dout(n19364));
  jor  g02102(.dina(n19364), .dinb(n19273), .dout(n19365));
  jxor g02103(.dina(n19267), .dinb(n360), .dout(n19366));
  jand g02104(.dina(n19366), .dinb(n19365), .dout(n19367));
  jor  g02105(.dina(n19367), .dinb(n19268), .dout(n19368));
  jxor g02106(.dina(n19254), .dinb(n361), .dout(n19369));
  jand g02107(.dina(n19369), .dinb(n19368), .dout(n19370));
  jor  g02108(.dina(n19370), .dinb(n19263), .dout(n19371));
  jand g02109(.dina(n19371), .dinb(n19262), .dout(n19372));
  jor  g02110(.dina(n19372), .dinb(n19259), .dout(n19373));
  jand g02111(.dina(n19373), .dinb(n1429), .dout(n19374));
  jor  g02112(.dina(n19374), .dinb(n19254), .dout(n19375));
  jnot g02113(.din(n19374), .dout(n19376));
  jxor g02114(.dina(n19369), .dinb(n19368), .dout(n19377));
  jor  g02115(.dina(n19377), .dinb(n19376), .dout(n19378));
  jand g02116(.dina(n19378), .dinb(n19375), .dout(n19379));
  jand g02117(.dina(n19371), .dinb(n1429), .dout(n19380));
  jand g02118(.dina(n19380), .dinb(n364), .dout(n19381));
  jor  g02119(.dina(n19381), .dinb(n19376), .dout(n19382));
  jand g02120(.dina(n19382), .dinb(n19258), .dout(n19383));
  jand g02121(.dina(n19383), .dinb(n355), .dout(n19384));
  jnot g02122(.din(n19383), .dout(n19385));
  jand g02123(.dina(n19385), .dinb(b16 ), .dout(n19386));
  jnot g02124(.din(n19386), .dout(n19387));
  jand g02125(.dina(n19379), .dinb(n364), .dout(n19388));
  jor  g02126(.dina(n19374), .dinb(n19267), .dout(n19389));
  jxor g02127(.dina(n19366), .dinb(n19365), .dout(n19390));
  jor  g02128(.dina(n19390), .dinb(n19376), .dout(n19391));
  jand g02129(.dina(n19391), .dinb(n19389), .dout(n19392));
  jand g02130(.dina(n19392), .dinb(n361), .dout(n19393));
  jor  g02131(.dina(n19374), .dinb(n19272), .dout(n19394));
  jxor g02132(.dina(n19363), .dinb(n19362), .dout(n19395));
  jor  g02133(.dina(n19395), .dinb(n19376), .dout(n19396));
  jand g02134(.dina(n19396), .dinb(n19394), .dout(n19397));
  jand g02135(.dina(n19397), .dinb(n360), .dout(n19398));
  jor  g02136(.dina(n19374), .dinb(n19277), .dout(n19399));
  jxor g02137(.dina(n19360), .dinb(n19359), .dout(n19400));
  jor  g02138(.dina(n19400), .dinb(n19376), .dout(n19401));
  jand g02139(.dina(n19401), .dinb(n19399), .dout(n19402));
  jand g02140(.dina(n19402), .dinb(n363), .dout(n19403));
  jor  g02141(.dina(n19374), .dinb(n19282), .dout(n19404));
  jxor g02142(.dina(n19357), .dinb(n19356), .dout(n19405));
  jor  g02143(.dina(n19405), .dinb(n19376), .dout(n19406));
  jand g02144(.dina(n19406), .dinb(n19404), .dout(n19407));
  jand g02145(.dina(n19407), .dinb(n359), .dout(n19408));
  jor  g02146(.dina(n19374), .dinb(n19287), .dout(n19409));
  jxor g02147(.dina(n19354), .dinb(n19353), .dout(n19410));
  jor  g02148(.dina(n19410), .dinb(n19376), .dout(n19411));
  jand g02149(.dina(n19411), .dinb(n19409), .dout(n19412));
  jand g02150(.dina(n19412), .dinb(n369), .dout(n19413));
  jor  g02151(.dina(n19374), .dinb(n19292), .dout(n19414));
  jxor g02152(.dina(n19351), .dinb(n19350), .dout(n19415));
  jor  g02153(.dina(n19415), .dinb(n19376), .dout(n19416));
  jand g02154(.dina(n19416), .dinb(n19414), .dout(n19417));
  jand g02155(.dina(n19417), .dinb(n368), .dout(n19418));
  jor  g02156(.dina(n19374), .dinb(n19297), .dout(n19419));
  jxor g02157(.dina(n19348), .dinb(n19347), .dout(n19420));
  jor  g02158(.dina(n19420), .dinb(n19376), .dout(n19421));
  jand g02159(.dina(n19421), .dinb(n19419), .dout(n19422));
  jand g02160(.dina(n19422), .dinb(n367), .dout(n19423));
  jor  g02161(.dina(n19374), .dinb(n19302), .dout(n19424));
  jxor g02162(.dina(n19345), .dinb(n19344), .dout(n19425));
  jor  g02163(.dina(n19425), .dinb(n19376), .dout(n19426));
  jand g02164(.dina(n19426), .dinb(n19424), .dout(n19427));
  jand g02165(.dina(n19427), .dinb(n265), .dout(n19428));
  jor  g02166(.dina(n19374), .dinb(n19307), .dout(n19429));
  jxor g02167(.dina(n19342), .dinb(n19341), .dout(n19430));
  jor  g02168(.dina(n19430), .dinb(n19376), .dout(n19431));
  jand g02169(.dina(n19431), .dinb(n19429), .dout(n19432));
  jand g02170(.dina(n19432), .dinb(n378), .dout(n19433));
  jor  g02171(.dina(n19374), .dinb(n19312), .dout(n19434));
  jxor g02172(.dina(n19339), .dinb(n19338), .dout(n19435));
  jor  g02173(.dina(n19435), .dinb(n19376), .dout(n19436));
  jand g02174(.dina(n19436), .dinb(n19434), .dout(n19437));
  jand g02175(.dina(n19437), .dinb(n377), .dout(n19438));
  jor  g02176(.dina(n19374), .dinb(n19317), .dout(n19439));
  jxor g02177(.dina(n19336), .dinb(n19335), .dout(n19440));
  jor  g02178(.dina(n19440), .dinb(n19376), .dout(n19441));
  jand g02179(.dina(n19441), .dinb(n19439), .dout(n19442));
  jand g02180(.dina(n19442), .dinb(n376), .dout(n19443));
  jor  g02181(.dina(n19374), .dinb(n19324), .dout(n19444));
  jxor g02182(.dina(n19333), .dinb(n19332), .dout(n19445));
  jor  g02183(.dina(n19445), .dinb(n19376), .dout(n19446));
  jand g02184(.dina(n19446), .dinb(n19444), .dout(n19447));
  jand g02185(.dina(n19447), .dinb(n264), .dout(n19448));
  jor  g02186(.dina(n19374), .dinb(n19329), .dout(n19449));
  jxor g02187(.dina(n19330), .dinb(n1571), .dout(n19450));
  jand g02188(.dina(n19450), .dinb(n19374), .dout(n19451));
  jnot g02189(.din(n19451), .dout(n19452));
  jand g02190(.dina(n19452), .dinb(n19449), .dout(n19453));
  jnot g02191(.din(n19453), .dout(n19454));
  jand g02192(.dina(n19454), .dinb(n386), .dout(n19455));
  jnot g02193(.din(n1430), .dout(n19456));
  jnot g02194(.din(n19259), .dout(n19457));
  jnot g02195(.din(n19263), .dout(n19458));
  jnot g02196(.din(n19268), .dout(n19459));
  jnot g02197(.din(n19273), .dout(n19460));
  jnot g02198(.din(n19278), .dout(n19461));
  jnot g02199(.din(n19283), .dout(n19462));
  jnot g02200(.din(n19288), .dout(n19463));
  jnot g02201(.din(n19293), .dout(n19464));
  jnot g02202(.din(n19298), .dout(n19465));
  jnot g02203(.din(n19303), .dout(n19466));
  jnot g02204(.din(n19308), .dout(n19467));
  jnot g02205(.din(n19313), .dout(n19468));
  jnot g02206(.din(n19318), .dout(n19469));
  jnot g02207(.din(n19325), .dout(n19470));
  jnot g02208(.din(n19328), .dout(n19471));
  jxor g02209(.dina(n19329), .dinb(n259), .dout(n19472));
  jor  g02210(.dina(n19472), .dinb(n1570), .dout(n19473));
  jand g02211(.dina(n19473), .dinb(n19471), .dout(n19474));
  jnot g02212(.din(n19333), .dout(n19475));
  jor  g02213(.dina(n19475), .dinb(n19474), .dout(n19476));
  jand g02214(.dina(n19476), .dinb(n19470), .dout(n19477));
  jnot g02215(.din(n19336), .dout(n19478));
  jor  g02216(.dina(n19478), .dinb(n19477), .dout(n19479));
  jand g02217(.dina(n19479), .dinb(n19469), .dout(n19480));
  jnot g02218(.din(n19339), .dout(n19481));
  jor  g02219(.dina(n19481), .dinb(n19480), .dout(n19482));
  jand g02220(.dina(n19482), .dinb(n19468), .dout(n19483));
  jnot g02221(.din(n19342), .dout(n19484));
  jor  g02222(.dina(n19484), .dinb(n19483), .dout(n19485));
  jand g02223(.dina(n19485), .dinb(n19467), .dout(n19486));
  jnot g02224(.din(n19345), .dout(n19487));
  jor  g02225(.dina(n19487), .dinb(n19486), .dout(n19488));
  jand g02226(.dina(n19488), .dinb(n19466), .dout(n19489));
  jnot g02227(.din(n19348), .dout(n19490));
  jor  g02228(.dina(n19490), .dinb(n19489), .dout(n19491));
  jand g02229(.dina(n19491), .dinb(n19465), .dout(n19492));
  jnot g02230(.din(n19351), .dout(n19493));
  jor  g02231(.dina(n19493), .dinb(n19492), .dout(n19494));
  jand g02232(.dina(n19494), .dinb(n19464), .dout(n19495));
  jnot g02233(.din(n19354), .dout(n19496));
  jor  g02234(.dina(n19496), .dinb(n19495), .dout(n19497));
  jand g02235(.dina(n19497), .dinb(n19463), .dout(n19498));
  jnot g02236(.din(n19357), .dout(n19499));
  jor  g02237(.dina(n19499), .dinb(n19498), .dout(n19500));
  jand g02238(.dina(n19500), .dinb(n19462), .dout(n19501));
  jnot g02239(.din(n19360), .dout(n19502));
  jor  g02240(.dina(n19502), .dinb(n19501), .dout(n19503));
  jand g02241(.dina(n19503), .dinb(n19461), .dout(n19504));
  jnot g02242(.din(n19363), .dout(n19505));
  jor  g02243(.dina(n19505), .dinb(n19504), .dout(n19506));
  jand g02244(.dina(n19506), .dinb(n19460), .dout(n19507));
  jnot g02245(.din(n19366), .dout(n19508));
  jor  g02246(.dina(n19508), .dinb(n19507), .dout(n19509));
  jand g02247(.dina(n19509), .dinb(n19459), .dout(n19510));
  jnot g02248(.din(n19369), .dout(n19511));
  jor  g02249(.dina(n19511), .dinb(n19510), .dout(n19512));
  jand g02250(.dina(n19512), .dinb(n19458), .dout(n19513));
  jor  g02251(.dina(n19513), .dinb(n19261), .dout(n19514));
  jand g02252(.dina(n19514), .dinb(n19457), .dout(n19515));
  jor  g02253(.dina(n19515), .dinb(n19456), .dout(n19516));
  jand g02254(.dina(n19516), .dinb(a48 ), .dout(n19517));
  jnot g02255(.din(n1700), .dout(n19518));
  jor  g02256(.dina(n19515), .dinb(n19518), .dout(n19519));
  jnot g02257(.din(n19519), .dout(n19520));
  jor  g02258(.dina(n19520), .dinb(n19517), .dout(n19521));
  jand g02259(.dina(n19521), .dinb(n259), .dout(n19522));
  jand g02260(.dina(n19373), .dinb(n1430), .dout(n19523));
  jor  g02261(.dina(n19523), .dinb(n1569), .dout(n19524));
  jand g02262(.dina(n19519), .dinb(n19524), .dout(n19525));
  jxor g02263(.dina(n19525), .dinb(b1 ), .dout(n19526));
  jand g02264(.dina(n19526), .dinb(n1708), .dout(n19527));
  jor  g02265(.dina(n19527), .dinb(n19522), .dout(n19528));
  jxor g02266(.dina(n19453), .dinb(b2 ), .dout(n19529));
  jand g02267(.dina(n19529), .dinb(n19528), .dout(n19530));
  jor  g02268(.dina(n19530), .dinb(n19455), .dout(n19531));
  jxor g02269(.dina(n19447), .dinb(n264), .dout(n19532));
  jand g02270(.dina(n19532), .dinb(n19531), .dout(n19533));
  jor  g02271(.dina(n19533), .dinb(n19448), .dout(n19534));
  jxor g02272(.dina(n19442), .dinb(n376), .dout(n19535));
  jand g02273(.dina(n19535), .dinb(n19534), .dout(n19536));
  jor  g02274(.dina(n19536), .dinb(n19443), .dout(n19537));
  jxor g02275(.dina(n19437), .dinb(n377), .dout(n19538));
  jand g02276(.dina(n19538), .dinb(n19537), .dout(n19539));
  jor  g02277(.dina(n19539), .dinb(n19438), .dout(n19540));
  jxor g02278(.dina(n19432), .dinb(n378), .dout(n19541));
  jand g02279(.dina(n19541), .dinb(n19540), .dout(n19542));
  jor  g02280(.dina(n19542), .dinb(n19433), .dout(n19543));
  jxor g02281(.dina(n19427), .dinb(n265), .dout(n19544));
  jand g02282(.dina(n19544), .dinb(n19543), .dout(n19545));
  jor  g02283(.dina(n19545), .dinb(n19428), .dout(n19546));
  jxor g02284(.dina(n19422), .dinb(n367), .dout(n19547));
  jand g02285(.dina(n19547), .dinb(n19546), .dout(n19548));
  jor  g02286(.dina(n19548), .dinb(n19423), .dout(n19549));
  jxor g02287(.dina(n19417), .dinb(n368), .dout(n19550));
  jand g02288(.dina(n19550), .dinb(n19549), .dout(n19551));
  jor  g02289(.dina(n19551), .dinb(n19418), .dout(n19552));
  jxor g02290(.dina(n19412), .dinb(n369), .dout(n19553));
  jand g02291(.dina(n19553), .dinb(n19552), .dout(n19554));
  jor  g02292(.dina(n19554), .dinb(n19413), .dout(n19555));
  jxor g02293(.dina(n19407), .dinb(n359), .dout(n19556));
  jand g02294(.dina(n19556), .dinb(n19555), .dout(n19557));
  jor  g02295(.dina(n19557), .dinb(n19408), .dout(n19558));
  jxor g02296(.dina(n19402), .dinb(n363), .dout(n19559));
  jand g02297(.dina(n19559), .dinb(n19558), .dout(n19560));
  jor  g02298(.dina(n19560), .dinb(n19403), .dout(n19561));
  jxor g02299(.dina(n19397), .dinb(n360), .dout(n19562));
  jand g02300(.dina(n19562), .dinb(n19561), .dout(n19563));
  jor  g02301(.dina(n19563), .dinb(n19398), .dout(n19564));
  jxor g02302(.dina(n19392), .dinb(n361), .dout(n19565));
  jand g02303(.dina(n19565), .dinb(n19564), .dout(n19566));
  jor  g02304(.dina(n19566), .dinb(n19393), .dout(n19567));
  jxor g02305(.dina(n19379), .dinb(n364), .dout(n19568));
  jand g02306(.dina(n19568), .dinb(n19567), .dout(n19569));
  jor  g02307(.dina(n19569), .dinb(n19388), .dout(n19570));
  jand g02308(.dina(n19570), .dinb(n19387), .dout(n19571));
  jor  g02309(.dina(n19571), .dinb(n19384), .dout(n19572));
  jand g02310(.dina(n19572), .dinb(n422), .dout(n19573));
  jor  g02311(.dina(n19573), .dinb(n19379), .dout(n19574));
  jnot g02312(.din(n19573), .dout(n19575));
  jxor g02313(.dina(n19568), .dinb(n19567), .dout(n19576));
  jor  g02314(.dina(n19576), .dinb(n19575), .dout(n19577));
  jand g02315(.dina(n19577), .dinb(n19574), .dout(n19578));
  jand g02316(.dina(n19575), .dinb(n19383), .dout(n19579));
  jand g02317(.dina(n19570), .dinb(n19384), .dout(n19580));
  jand g02318(.dina(n19580), .dinb(n422), .dout(n19581));
  jor  g02319(.dina(n19581), .dinb(n19579), .dout(n19582));
  jand g02320(.dina(n19582), .dinb(n422), .dout(n19583));
  jand g02321(.dina(n19578), .dinb(n355), .dout(n19584));
  jor  g02322(.dina(n19573), .dinb(n19392), .dout(n19585));
  jxor g02323(.dina(n19565), .dinb(n19564), .dout(n19586));
  jor  g02324(.dina(n19586), .dinb(n19575), .dout(n19587));
  jand g02325(.dina(n19587), .dinb(n19585), .dout(n19588));
  jand g02326(.dina(n19588), .dinb(n364), .dout(n19589));
  jor  g02327(.dina(n19573), .dinb(n19397), .dout(n19590));
  jxor g02328(.dina(n19562), .dinb(n19561), .dout(n19591));
  jor  g02329(.dina(n19591), .dinb(n19575), .dout(n19592));
  jand g02330(.dina(n19592), .dinb(n19590), .dout(n19593));
  jand g02331(.dina(n19593), .dinb(n361), .dout(n19594));
  jor  g02332(.dina(n19573), .dinb(n19402), .dout(n19595));
  jxor g02333(.dina(n19559), .dinb(n19558), .dout(n19596));
  jor  g02334(.dina(n19596), .dinb(n19575), .dout(n19597));
  jand g02335(.dina(n19597), .dinb(n19595), .dout(n19598));
  jand g02336(.dina(n19598), .dinb(n360), .dout(n19599));
  jor  g02337(.dina(n19573), .dinb(n19407), .dout(n19600));
  jxor g02338(.dina(n19556), .dinb(n19555), .dout(n19601));
  jor  g02339(.dina(n19601), .dinb(n19575), .dout(n19602));
  jand g02340(.dina(n19602), .dinb(n19600), .dout(n19603));
  jand g02341(.dina(n19603), .dinb(n363), .dout(n19604));
  jor  g02342(.dina(n19573), .dinb(n19412), .dout(n19605));
  jxor g02343(.dina(n19553), .dinb(n19552), .dout(n19606));
  jor  g02344(.dina(n19606), .dinb(n19575), .dout(n19607));
  jand g02345(.dina(n19607), .dinb(n19605), .dout(n19608));
  jand g02346(.dina(n19608), .dinb(n359), .dout(n19609));
  jor  g02347(.dina(n19573), .dinb(n19417), .dout(n19610));
  jxor g02348(.dina(n19550), .dinb(n19549), .dout(n19611));
  jor  g02349(.dina(n19611), .dinb(n19575), .dout(n19612));
  jand g02350(.dina(n19612), .dinb(n19610), .dout(n19613));
  jand g02351(.dina(n19613), .dinb(n369), .dout(n19614));
  jor  g02352(.dina(n19573), .dinb(n19422), .dout(n19615));
  jxor g02353(.dina(n19547), .dinb(n19546), .dout(n19616));
  jor  g02354(.dina(n19616), .dinb(n19575), .dout(n19617));
  jand g02355(.dina(n19617), .dinb(n19615), .dout(n19618));
  jand g02356(.dina(n19618), .dinb(n368), .dout(n19619));
  jor  g02357(.dina(n19573), .dinb(n19427), .dout(n19620));
  jxor g02358(.dina(n19544), .dinb(n19543), .dout(n19621));
  jor  g02359(.dina(n19621), .dinb(n19575), .dout(n19622));
  jand g02360(.dina(n19622), .dinb(n19620), .dout(n19623));
  jand g02361(.dina(n19623), .dinb(n367), .dout(n19624));
  jor  g02362(.dina(n19573), .dinb(n19432), .dout(n19625));
  jxor g02363(.dina(n19541), .dinb(n19540), .dout(n19626));
  jor  g02364(.dina(n19626), .dinb(n19575), .dout(n19627));
  jand g02365(.dina(n19627), .dinb(n19625), .dout(n19628));
  jand g02366(.dina(n19628), .dinb(n265), .dout(n19629));
  jor  g02367(.dina(n19573), .dinb(n19437), .dout(n19630));
  jxor g02368(.dina(n19538), .dinb(n19537), .dout(n19631));
  jor  g02369(.dina(n19631), .dinb(n19575), .dout(n19632));
  jand g02370(.dina(n19632), .dinb(n19630), .dout(n19633));
  jand g02371(.dina(n19633), .dinb(n378), .dout(n19634));
  jor  g02372(.dina(n19573), .dinb(n19442), .dout(n19635));
  jxor g02373(.dina(n19535), .dinb(n19534), .dout(n19636));
  jor  g02374(.dina(n19636), .dinb(n19575), .dout(n19637));
  jand g02375(.dina(n19637), .dinb(n19635), .dout(n19638));
  jand g02376(.dina(n19638), .dinb(n377), .dout(n19639));
  jor  g02377(.dina(n19573), .dinb(n19447), .dout(n19640));
  jxor g02378(.dina(n19532), .dinb(n19531), .dout(n19641));
  jor  g02379(.dina(n19641), .dinb(n19575), .dout(n19642));
  jand g02380(.dina(n19642), .dinb(n19640), .dout(n19643));
  jand g02381(.dina(n19643), .dinb(n376), .dout(n19644));
  jor  g02382(.dina(n19573), .dinb(n19454), .dout(n19645));
  jxor g02383(.dina(n19529), .dinb(n19528), .dout(n19646));
  jor  g02384(.dina(n19646), .dinb(n19575), .dout(n19647));
  jand g02385(.dina(n19647), .dinb(n19645), .dout(n19648));
  jand g02386(.dina(n19648), .dinb(n264), .dout(n19649));
  jor  g02387(.dina(n19573), .dinb(n19525), .dout(n19650));
  jxor g02388(.dina(n19526), .dinb(n1708), .dout(n19651));
  jand g02389(.dina(n19651), .dinb(n19573), .dout(n19652));
  jnot g02390(.din(n19652), .dout(n19653));
  jand g02391(.dina(n19653), .dinb(n19650), .dout(n19654));
  jnot g02392(.din(n19654), .dout(n19655));
  jand g02393(.dina(n19655), .dinb(n386), .dout(n19656));
  jnot g02394(.din(n1842), .dout(n19657));
  jnot g02395(.din(n19384), .dout(n19658));
  jnot g02396(.din(n19388), .dout(n19659));
  jnot g02397(.din(n19393), .dout(n19660));
  jnot g02398(.din(n19398), .dout(n19661));
  jnot g02399(.din(n19403), .dout(n19662));
  jnot g02400(.din(n19408), .dout(n19663));
  jnot g02401(.din(n19413), .dout(n19664));
  jnot g02402(.din(n19418), .dout(n19665));
  jnot g02403(.din(n19423), .dout(n19666));
  jnot g02404(.din(n19428), .dout(n19667));
  jnot g02405(.din(n19433), .dout(n19668));
  jnot g02406(.din(n19438), .dout(n19669));
  jnot g02407(.din(n19443), .dout(n19670));
  jnot g02408(.din(n19448), .dout(n19671));
  jnot g02409(.din(n19455), .dout(n19672));
  jnot g02410(.din(n19522), .dout(n19673));
  jxor g02411(.dina(n19525), .dinb(n259), .dout(n19674));
  jor  g02412(.dina(n19674), .dinb(n1707), .dout(n19675));
  jand g02413(.dina(n19675), .dinb(n19673), .dout(n19676));
  jnot g02414(.din(n19529), .dout(n19677));
  jor  g02415(.dina(n19677), .dinb(n19676), .dout(n19678));
  jand g02416(.dina(n19678), .dinb(n19672), .dout(n19679));
  jnot g02417(.din(n19532), .dout(n19680));
  jor  g02418(.dina(n19680), .dinb(n19679), .dout(n19681));
  jand g02419(.dina(n19681), .dinb(n19671), .dout(n19682));
  jnot g02420(.din(n19535), .dout(n19683));
  jor  g02421(.dina(n19683), .dinb(n19682), .dout(n19684));
  jand g02422(.dina(n19684), .dinb(n19670), .dout(n19685));
  jnot g02423(.din(n19538), .dout(n19686));
  jor  g02424(.dina(n19686), .dinb(n19685), .dout(n19687));
  jand g02425(.dina(n19687), .dinb(n19669), .dout(n19688));
  jnot g02426(.din(n19541), .dout(n19689));
  jor  g02427(.dina(n19689), .dinb(n19688), .dout(n19690));
  jand g02428(.dina(n19690), .dinb(n19668), .dout(n19691));
  jnot g02429(.din(n19544), .dout(n19692));
  jor  g02430(.dina(n19692), .dinb(n19691), .dout(n19693));
  jand g02431(.dina(n19693), .dinb(n19667), .dout(n19694));
  jnot g02432(.din(n19547), .dout(n19695));
  jor  g02433(.dina(n19695), .dinb(n19694), .dout(n19696));
  jand g02434(.dina(n19696), .dinb(n19666), .dout(n19697));
  jnot g02435(.din(n19550), .dout(n19698));
  jor  g02436(.dina(n19698), .dinb(n19697), .dout(n19699));
  jand g02437(.dina(n19699), .dinb(n19665), .dout(n19700));
  jnot g02438(.din(n19553), .dout(n19701));
  jor  g02439(.dina(n19701), .dinb(n19700), .dout(n19702));
  jand g02440(.dina(n19702), .dinb(n19664), .dout(n19703));
  jnot g02441(.din(n19556), .dout(n19704));
  jor  g02442(.dina(n19704), .dinb(n19703), .dout(n19705));
  jand g02443(.dina(n19705), .dinb(n19663), .dout(n19706));
  jnot g02444(.din(n19559), .dout(n19707));
  jor  g02445(.dina(n19707), .dinb(n19706), .dout(n19708));
  jand g02446(.dina(n19708), .dinb(n19662), .dout(n19709));
  jnot g02447(.din(n19562), .dout(n19710));
  jor  g02448(.dina(n19710), .dinb(n19709), .dout(n19711));
  jand g02449(.dina(n19711), .dinb(n19661), .dout(n19712));
  jnot g02450(.din(n19565), .dout(n19713));
  jor  g02451(.dina(n19713), .dinb(n19712), .dout(n19714));
  jand g02452(.dina(n19714), .dinb(n19660), .dout(n19715));
  jnot g02453(.din(n19568), .dout(n19716));
  jor  g02454(.dina(n19716), .dinb(n19715), .dout(n19717));
  jand g02455(.dina(n19717), .dinb(n19659), .dout(n19718));
  jor  g02456(.dina(n19718), .dinb(n19386), .dout(n19719));
  jand g02457(.dina(n19719), .dinb(n19658), .dout(n19720));
  jor  g02458(.dina(n19720), .dinb(n19657), .dout(n19721));
  jand g02459(.dina(n19721), .dinb(a47 ), .dout(n19722));
  jnot g02460(.din(n1845), .dout(n19723));
  jor  g02461(.dina(n19720), .dinb(n19723), .dout(n19724));
  jnot g02462(.din(n19724), .dout(n19725));
  jor  g02463(.dina(n19725), .dinb(n19722), .dout(n19726));
  jand g02464(.dina(n19726), .dinb(n259), .dout(n19727));
  jand g02465(.dina(n19572), .dinb(n1842), .dout(n19728));
  jor  g02466(.dina(n19728), .dinb(n1706), .dout(n19729));
  jand g02467(.dina(n19724), .dinb(n19729), .dout(n19730));
  jxor g02468(.dina(n19730), .dinb(b1 ), .dout(n19731));
  jand g02469(.dina(n19731), .dinb(n1853), .dout(n19732));
  jor  g02470(.dina(n19732), .dinb(n19727), .dout(n19733));
  jxor g02471(.dina(n19654), .dinb(b2 ), .dout(n19734));
  jand g02472(.dina(n19734), .dinb(n19733), .dout(n19735));
  jor  g02473(.dina(n19735), .dinb(n19656), .dout(n19736));
  jxor g02474(.dina(n19648), .dinb(n264), .dout(n19737));
  jand g02475(.dina(n19737), .dinb(n19736), .dout(n19738));
  jor  g02476(.dina(n19738), .dinb(n19649), .dout(n19739));
  jxor g02477(.dina(n19643), .dinb(n376), .dout(n19740));
  jand g02478(.dina(n19740), .dinb(n19739), .dout(n19741));
  jor  g02479(.dina(n19741), .dinb(n19644), .dout(n19742));
  jxor g02480(.dina(n19638), .dinb(n377), .dout(n19743));
  jand g02481(.dina(n19743), .dinb(n19742), .dout(n19744));
  jor  g02482(.dina(n19744), .dinb(n19639), .dout(n19745));
  jxor g02483(.dina(n19633), .dinb(n378), .dout(n19746));
  jand g02484(.dina(n19746), .dinb(n19745), .dout(n19747));
  jor  g02485(.dina(n19747), .dinb(n19634), .dout(n19748));
  jxor g02486(.dina(n19628), .dinb(n265), .dout(n19749));
  jand g02487(.dina(n19749), .dinb(n19748), .dout(n19750));
  jor  g02488(.dina(n19750), .dinb(n19629), .dout(n19751));
  jxor g02489(.dina(n19623), .dinb(n367), .dout(n19752));
  jand g02490(.dina(n19752), .dinb(n19751), .dout(n19753));
  jor  g02491(.dina(n19753), .dinb(n19624), .dout(n19754));
  jxor g02492(.dina(n19618), .dinb(n368), .dout(n19755));
  jand g02493(.dina(n19755), .dinb(n19754), .dout(n19756));
  jor  g02494(.dina(n19756), .dinb(n19619), .dout(n19757));
  jxor g02495(.dina(n19613), .dinb(n369), .dout(n19758));
  jand g02496(.dina(n19758), .dinb(n19757), .dout(n19759));
  jor  g02497(.dina(n19759), .dinb(n19614), .dout(n19760));
  jxor g02498(.dina(n19608), .dinb(n359), .dout(n19761));
  jand g02499(.dina(n19761), .dinb(n19760), .dout(n19762));
  jor  g02500(.dina(n19762), .dinb(n19609), .dout(n19763));
  jxor g02501(.dina(n19603), .dinb(n363), .dout(n19764));
  jand g02502(.dina(n19764), .dinb(n19763), .dout(n19765));
  jor  g02503(.dina(n19765), .dinb(n19604), .dout(n19766));
  jxor g02504(.dina(n19598), .dinb(n360), .dout(n19767));
  jand g02505(.dina(n19767), .dinb(n19766), .dout(n19768));
  jor  g02506(.dina(n19768), .dinb(n19599), .dout(n19769));
  jxor g02507(.dina(n19593), .dinb(n361), .dout(n19770));
  jand g02508(.dina(n19770), .dinb(n19769), .dout(n19771));
  jor  g02509(.dina(n19771), .dinb(n19594), .dout(n19772));
  jxor g02510(.dina(n19588), .dinb(n364), .dout(n19773));
  jand g02511(.dina(n19773), .dinb(n19772), .dout(n19774));
  jor  g02512(.dina(n19774), .dinb(n19589), .dout(n19775));
  jxor g02513(.dina(n19578), .dinb(n355), .dout(n19776));
  jand g02514(.dina(n19776), .dinb(n19775), .dout(n19777));
  jor  g02515(.dina(n19777), .dinb(n19584), .dout(n19778));
  jxor g02516(.dina(n19582), .dinb(b17 ), .dout(n19779));
  jnot g02517(.din(n19779), .dout(n19780));
  jand g02518(.dina(n19780), .dinb(n19778), .dout(n19781));
  jand g02519(.dina(n19781), .dinb(n354), .dout(n19782));
  jor  g02520(.dina(n19782), .dinb(n19583), .dout(n19783));
  jor  g02521(.dina(n19783), .dinb(n19578), .dout(n19784));
  jnot g02522(.din(n19783), .dout(n19785));
  jxor g02523(.dina(n19776), .dinb(n19775), .dout(n19786));
  jor  g02524(.dina(n19786), .dinb(n19785), .dout(n19787));
  jand g02525(.dina(n19787), .dinb(n19784), .dout(n19788));
  jxor g02526(.dina(n19780), .dinb(n19778), .dout(n19789));
  jor  g02527(.dina(n19789), .dinb(n19785), .dout(n19790));
  jor  g02528(.dina(n19782), .dinb(n19582), .dout(n19791));
  jand g02529(.dina(n19791), .dinb(n19790), .dout(n19792));
  jand g02530(.dina(n19792), .dinb(n266), .dout(n19793));
  jnot g02531(.din(n19792), .dout(n19794));
  jand g02532(.dina(n19794), .dinb(b18 ), .dout(n19795));
  jnot g02533(.din(n19795), .dout(n19796));
  jand g02534(.dina(n19788), .dinb(n356), .dout(n19797));
  jor  g02535(.dina(n19783), .dinb(n19588), .dout(n19798));
  jxor g02536(.dina(n19773), .dinb(n19772), .dout(n19799));
  jor  g02537(.dina(n19799), .dinb(n19785), .dout(n19800));
  jand g02538(.dina(n19800), .dinb(n19798), .dout(n19801));
  jand g02539(.dina(n19801), .dinb(n355), .dout(n19802));
  jor  g02540(.dina(n19783), .dinb(n19593), .dout(n19803));
  jxor g02541(.dina(n19770), .dinb(n19769), .dout(n19804));
  jor  g02542(.dina(n19804), .dinb(n19785), .dout(n19805));
  jand g02543(.dina(n19805), .dinb(n19803), .dout(n19806));
  jand g02544(.dina(n19806), .dinb(n364), .dout(n19807));
  jor  g02545(.dina(n19783), .dinb(n19598), .dout(n19808));
  jxor g02546(.dina(n19767), .dinb(n19766), .dout(n19809));
  jor  g02547(.dina(n19809), .dinb(n19785), .dout(n19810));
  jand g02548(.dina(n19810), .dinb(n19808), .dout(n19811));
  jand g02549(.dina(n19811), .dinb(n361), .dout(n19812));
  jor  g02550(.dina(n19783), .dinb(n19603), .dout(n19813));
  jxor g02551(.dina(n19764), .dinb(n19763), .dout(n19814));
  jor  g02552(.dina(n19814), .dinb(n19785), .dout(n19815));
  jand g02553(.dina(n19815), .dinb(n19813), .dout(n19816));
  jand g02554(.dina(n19816), .dinb(n360), .dout(n19817));
  jor  g02555(.dina(n19783), .dinb(n19608), .dout(n19818));
  jxor g02556(.dina(n19761), .dinb(n19760), .dout(n19819));
  jor  g02557(.dina(n19819), .dinb(n19785), .dout(n19820));
  jand g02558(.dina(n19820), .dinb(n19818), .dout(n19821));
  jand g02559(.dina(n19821), .dinb(n363), .dout(n19822));
  jor  g02560(.dina(n19783), .dinb(n19613), .dout(n19823));
  jxor g02561(.dina(n19758), .dinb(n19757), .dout(n19824));
  jor  g02562(.dina(n19824), .dinb(n19785), .dout(n19825));
  jand g02563(.dina(n19825), .dinb(n19823), .dout(n19826));
  jand g02564(.dina(n19826), .dinb(n359), .dout(n19827));
  jor  g02565(.dina(n19783), .dinb(n19618), .dout(n19828));
  jxor g02566(.dina(n19755), .dinb(n19754), .dout(n19829));
  jor  g02567(.dina(n19829), .dinb(n19785), .dout(n19830));
  jand g02568(.dina(n19830), .dinb(n19828), .dout(n19831));
  jand g02569(.dina(n19831), .dinb(n369), .dout(n19832));
  jor  g02570(.dina(n19783), .dinb(n19623), .dout(n19833));
  jxor g02571(.dina(n19752), .dinb(n19751), .dout(n19834));
  jor  g02572(.dina(n19834), .dinb(n19785), .dout(n19835));
  jand g02573(.dina(n19835), .dinb(n19833), .dout(n19836));
  jand g02574(.dina(n19836), .dinb(n368), .dout(n19837));
  jor  g02575(.dina(n19783), .dinb(n19628), .dout(n19838));
  jxor g02576(.dina(n19749), .dinb(n19748), .dout(n19839));
  jor  g02577(.dina(n19839), .dinb(n19785), .dout(n19840));
  jand g02578(.dina(n19840), .dinb(n19838), .dout(n19841));
  jand g02579(.dina(n19841), .dinb(n367), .dout(n19842));
  jor  g02580(.dina(n19783), .dinb(n19633), .dout(n19843));
  jxor g02581(.dina(n19746), .dinb(n19745), .dout(n19844));
  jor  g02582(.dina(n19844), .dinb(n19785), .dout(n19845));
  jand g02583(.dina(n19845), .dinb(n19843), .dout(n19846));
  jand g02584(.dina(n19846), .dinb(n265), .dout(n19847));
  jor  g02585(.dina(n19783), .dinb(n19638), .dout(n19848));
  jxor g02586(.dina(n19743), .dinb(n19742), .dout(n19849));
  jor  g02587(.dina(n19849), .dinb(n19785), .dout(n19850));
  jand g02588(.dina(n19850), .dinb(n19848), .dout(n19851));
  jand g02589(.dina(n19851), .dinb(n378), .dout(n19852));
  jor  g02590(.dina(n19783), .dinb(n19643), .dout(n19853));
  jxor g02591(.dina(n19740), .dinb(n19739), .dout(n19854));
  jor  g02592(.dina(n19854), .dinb(n19785), .dout(n19855));
  jand g02593(.dina(n19855), .dinb(n19853), .dout(n19856));
  jand g02594(.dina(n19856), .dinb(n377), .dout(n19857));
  jor  g02595(.dina(n19783), .dinb(n19648), .dout(n19858));
  jxor g02596(.dina(n19737), .dinb(n19736), .dout(n19859));
  jor  g02597(.dina(n19859), .dinb(n19785), .dout(n19860));
  jand g02598(.dina(n19860), .dinb(n19858), .dout(n19861));
  jand g02599(.dina(n19861), .dinb(n376), .dout(n19862));
  jor  g02600(.dina(n19783), .dinb(n19655), .dout(n19863));
  jxor g02601(.dina(n19734), .dinb(n19733), .dout(n19864));
  jor  g02602(.dina(n19864), .dinb(n19785), .dout(n19865));
  jand g02603(.dina(n19865), .dinb(n19863), .dout(n19866));
  jand g02604(.dina(n19866), .dinb(n264), .dout(n19867));
  jor  g02605(.dina(n19783), .dinb(n19726), .dout(n19868));
  jxor g02606(.dina(n19731), .dinb(n1853), .dout(n19869));
  jor  g02607(.dina(n19869), .dinb(n19785), .dout(n19870));
  jand g02608(.dina(n19870), .dinb(n19868), .dout(n19871));
  jand g02609(.dina(n19871), .dinb(n386), .dout(n19872));
  jand g02610(.dina(n19783), .dinb(b0 ), .dout(n19873));
  jxor g02611(.dina(n19873), .dinb(a46 ), .dout(n19874));
  jand g02612(.dina(n19874), .dinb(n259), .dout(n19875));
  jxor g02613(.dina(n19873), .dinb(n1851), .dout(n19876));
  jxor g02614(.dina(n19876), .dinb(b1 ), .dout(n19877));
  jand g02615(.dina(n19877), .dinb(n2003), .dout(n19878));
  jor  g02616(.dina(n19878), .dinb(n19875), .dout(n19879));
  jxor g02617(.dina(n19871), .dinb(n386), .dout(n19880));
  jand g02618(.dina(n19880), .dinb(n19879), .dout(n19881));
  jor  g02619(.dina(n19881), .dinb(n19872), .dout(n19882));
  jxor g02620(.dina(n19866), .dinb(n264), .dout(n19883));
  jand g02621(.dina(n19883), .dinb(n19882), .dout(n19884));
  jor  g02622(.dina(n19884), .dinb(n19867), .dout(n19885));
  jxor g02623(.dina(n19861), .dinb(n376), .dout(n19886));
  jand g02624(.dina(n19886), .dinb(n19885), .dout(n19887));
  jor  g02625(.dina(n19887), .dinb(n19862), .dout(n19888));
  jxor g02626(.dina(n19856), .dinb(n377), .dout(n19889));
  jand g02627(.dina(n19889), .dinb(n19888), .dout(n19890));
  jor  g02628(.dina(n19890), .dinb(n19857), .dout(n19891));
  jxor g02629(.dina(n19851), .dinb(n378), .dout(n19892));
  jand g02630(.dina(n19892), .dinb(n19891), .dout(n19893));
  jor  g02631(.dina(n19893), .dinb(n19852), .dout(n19894));
  jxor g02632(.dina(n19846), .dinb(n265), .dout(n19895));
  jand g02633(.dina(n19895), .dinb(n19894), .dout(n19896));
  jor  g02634(.dina(n19896), .dinb(n19847), .dout(n19897));
  jxor g02635(.dina(n19841), .dinb(n367), .dout(n19898));
  jand g02636(.dina(n19898), .dinb(n19897), .dout(n19899));
  jor  g02637(.dina(n19899), .dinb(n19842), .dout(n19900));
  jxor g02638(.dina(n19836), .dinb(n368), .dout(n19901));
  jand g02639(.dina(n19901), .dinb(n19900), .dout(n19902));
  jor  g02640(.dina(n19902), .dinb(n19837), .dout(n19903));
  jxor g02641(.dina(n19831), .dinb(n369), .dout(n19904));
  jand g02642(.dina(n19904), .dinb(n19903), .dout(n19905));
  jor  g02643(.dina(n19905), .dinb(n19832), .dout(n19906));
  jxor g02644(.dina(n19826), .dinb(n359), .dout(n19907));
  jand g02645(.dina(n19907), .dinb(n19906), .dout(n19908));
  jor  g02646(.dina(n19908), .dinb(n19827), .dout(n19909));
  jxor g02647(.dina(n19821), .dinb(n363), .dout(n19910));
  jand g02648(.dina(n19910), .dinb(n19909), .dout(n19911));
  jor  g02649(.dina(n19911), .dinb(n19822), .dout(n19912));
  jxor g02650(.dina(n19816), .dinb(n360), .dout(n19913));
  jand g02651(.dina(n19913), .dinb(n19912), .dout(n19914));
  jor  g02652(.dina(n19914), .dinb(n19817), .dout(n19915));
  jxor g02653(.dina(n19811), .dinb(n361), .dout(n19916));
  jand g02654(.dina(n19916), .dinb(n19915), .dout(n19917));
  jor  g02655(.dina(n19917), .dinb(n19812), .dout(n19918));
  jxor g02656(.dina(n19806), .dinb(n364), .dout(n19919));
  jand g02657(.dina(n19919), .dinb(n19918), .dout(n19920));
  jor  g02658(.dina(n19920), .dinb(n19807), .dout(n19921));
  jxor g02659(.dina(n19801), .dinb(n355), .dout(n19922));
  jand g02660(.dina(n19922), .dinb(n19921), .dout(n19923));
  jor  g02661(.dina(n19923), .dinb(n19802), .dout(n19924));
  jxor g02662(.dina(n19788), .dinb(n356), .dout(n19925));
  jand g02663(.dina(n19925), .dinb(n19924), .dout(n19926));
  jor  g02664(.dina(n19926), .dinb(n19797), .dout(n19927));
  jand g02665(.dina(n19927), .dinb(n19796), .dout(n19928));
  jor  g02666(.dina(n19928), .dinb(n19793), .dout(n19929));
  jand g02667(.dina(n19929), .dinb(n1910), .dout(n19930));
  jor  g02668(.dina(n19930), .dinb(n19788), .dout(n19931));
  jnot g02669(.din(n19930), .dout(n19932));
  jxor g02670(.dina(n19925), .dinb(n19924), .dout(n19933));
  jor  g02671(.dina(n19933), .dinb(n19932), .dout(n19934));
  jand g02672(.dina(n19934), .dinb(n19931), .dout(n19935));
  jand g02673(.dina(n19932), .dinb(n19792), .dout(n19936));
  jand g02674(.dina(n19927), .dinb(n19793), .dout(n19937));
  jor  g02675(.dina(n19937), .dinb(n19936), .dout(n19938));
  jand g02676(.dina(n19938), .dinb(n267), .dout(n19939));
  jnot g02677(.din(n19938), .dout(n19940));
  jand g02678(.dina(n19940), .dinb(b19 ), .dout(n19941));
  jnot g02679(.din(n19941), .dout(n19942));
  jand g02680(.dina(n19935), .dinb(n266), .dout(n19943));
  jor  g02681(.dina(n19930), .dinb(n19801), .dout(n19944));
  jxor g02682(.dina(n19922), .dinb(n19921), .dout(n19945));
  jor  g02683(.dina(n19945), .dinb(n19932), .dout(n19946));
  jand g02684(.dina(n19946), .dinb(n19944), .dout(n19947));
  jand g02685(.dina(n19947), .dinb(n356), .dout(n19948));
  jor  g02686(.dina(n19930), .dinb(n19806), .dout(n19949));
  jxor g02687(.dina(n19919), .dinb(n19918), .dout(n19950));
  jor  g02688(.dina(n19950), .dinb(n19932), .dout(n19951));
  jand g02689(.dina(n19951), .dinb(n19949), .dout(n19952));
  jand g02690(.dina(n19952), .dinb(n355), .dout(n19953));
  jor  g02691(.dina(n19930), .dinb(n19811), .dout(n19954));
  jxor g02692(.dina(n19916), .dinb(n19915), .dout(n19955));
  jor  g02693(.dina(n19955), .dinb(n19932), .dout(n19956));
  jand g02694(.dina(n19956), .dinb(n19954), .dout(n19957));
  jand g02695(.dina(n19957), .dinb(n364), .dout(n19958));
  jor  g02696(.dina(n19930), .dinb(n19816), .dout(n19959));
  jxor g02697(.dina(n19913), .dinb(n19912), .dout(n19960));
  jor  g02698(.dina(n19960), .dinb(n19932), .dout(n19961));
  jand g02699(.dina(n19961), .dinb(n19959), .dout(n19962));
  jand g02700(.dina(n19962), .dinb(n361), .dout(n19963));
  jor  g02701(.dina(n19930), .dinb(n19821), .dout(n19964));
  jxor g02702(.dina(n19910), .dinb(n19909), .dout(n19965));
  jor  g02703(.dina(n19965), .dinb(n19932), .dout(n19966));
  jand g02704(.dina(n19966), .dinb(n19964), .dout(n19967));
  jand g02705(.dina(n19967), .dinb(n360), .dout(n19968));
  jor  g02706(.dina(n19930), .dinb(n19826), .dout(n19969));
  jxor g02707(.dina(n19907), .dinb(n19906), .dout(n19970));
  jor  g02708(.dina(n19970), .dinb(n19932), .dout(n19971));
  jand g02709(.dina(n19971), .dinb(n19969), .dout(n19972));
  jand g02710(.dina(n19972), .dinb(n363), .dout(n19973));
  jor  g02711(.dina(n19930), .dinb(n19831), .dout(n19974));
  jxor g02712(.dina(n19904), .dinb(n19903), .dout(n19975));
  jor  g02713(.dina(n19975), .dinb(n19932), .dout(n19976));
  jand g02714(.dina(n19976), .dinb(n19974), .dout(n19977));
  jand g02715(.dina(n19977), .dinb(n359), .dout(n19978));
  jor  g02716(.dina(n19930), .dinb(n19836), .dout(n19979));
  jxor g02717(.dina(n19901), .dinb(n19900), .dout(n19980));
  jor  g02718(.dina(n19980), .dinb(n19932), .dout(n19981));
  jand g02719(.dina(n19981), .dinb(n19979), .dout(n19982));
  jand g02720(.dina(n19982), .dinb(n369), .dout(n19983));
  jor  g02721(.dina(n19930), .dinb(n19841), .dout(n19984));
  jxor g02722(.dina(n19898), .dinb(n19897), .dout(n19985));
  jor  g02723(.dina(n19985), .dinb(n19932), .dout(n19986));
  jand g02724(.dina(n19986), .dinb(n19984), .dout(n19987));
  jand g02725(.dina(n19987), .dinb(n368), .dout(n19988));
  jor  g02726(.dina(n19930), .dinb(n19846), .dout(n19989));
  jxor g02727(.dina(n19895), .dinb(n19894), .dout(n19990));
  jor  g02728(.dina(n19990), .dinb(n19932), .dout(n19991));
  jand g02729(.dina(n19991), .dinb(n19989), .dout(n19992));
  jand g02730(.dina(n19992), .dinb(n367), .dout(n19993));
  jor  g02731(.dina(n19930), .dinb(n19851), .dout(n19994));
  jxor g02732(.dina(n19892), .dinb(n19891), .dout(n19995));
  jor  g02733(.dina(n19995), .dinb(n19932), .dout(n19996));
  jand g02734(.dina(n19996), .dinb(n19994), .dout(n19997));
  jand g02735(.dina(n19997), .dinb(n265), .dout(n19998));
  jor  g02736(.dina(n19930), .dinb(n19856), .dout(n19999));
  jxor g02737(.dina(n19889), .dinb(n19888), .dout(n20000));
  jor  g02738(.dina(n20000), .dinb(n19932), .dout(n20001));
  jand g02739(.dina(n20001), .dinb(n19999), .dout(n20002));
  jand g02740(.dina(n20002), .dinb(n378), .dout(n20003));
  jor  g02741(.dina(n19930), .dinb(n19861), .dout(n20004));
  jxor g02742(.dina(n19886), .dinb(n19885), .dout(n20005));
  jor  g02743(.dina(n20005), .dinb(n19932), .dout(n20006));
  jand g02744(.dina(n20006), .dinb(n20004), .dout(n20007));
  jand g02745(.dina(n20007), .dinb(n377), .dout(n20008));
  jor  g02746(.dina(n19930), .dinb(n19866), .dout(n20009));
  jxor g02747(.dina(n19883), .dinb(n19882), .dout(n20010));
  jor  g02748(.dina(n20010), .dinb(n19932), .dout(n20011));
  jand g02749(.dina(n20011), .dinb(n20009), .dout(n20012));
  jand g02750(.dina(n20012), .dinb(n376), .dout(n20013));
  jor  g02751(.dina(n19930), .dinb(n19871), .dout(n20014));
  jxor g02752(.dina(n19880), .dinb(n19879), .dout(n20015));
  jor  g02753(.dina(n20015), .dinb(n19932), .dout(n20016));
  jand g02754(.dina(n20016), .dinb(n20014), .dout(n20017));
  jand g02755(.dina(n20017), .dinb(n264), .dout(n20018));
  jor  g02756(.dina(n19930), .dinb(n19874), .dout(n20019));
  jxor g02757(.dina(n19877), .dinb(n2003), .dout(n20020));
  jor  g02758(.dina(n20020), .dinb(n19932), .dout(n20021));
  jand g02759(.dina(n20021), .dinb(n20019), .dout(n20022));
  jand g02760(.dina(n20022), .dinb(n386), .dout(n20023));
  jnot g02761(.din(n1841), .dout(n20024));
  jnot g02762(.din(n19793), .dout(n20025));
  jnot g02763(.din(n19797), .dout(n20026));
  jnot g02764(.din(n19802), .dout(n20027));
  jnot g02765(.din(n19807), .dout(n20028));
  jnot g02766(.din(n19812), .dout(n20029));
  jnot g02767(.din(n19817), .dout(n20030));
  jnot g02768(.din(n19822), .dout(n20031));
  jnot g02769(.din(n19827), .dout(n20032));
  jnot g02770(.din(n19832), .dout(n20033));
  jnot g02771(.din(n19837), .dout(n20034));
  jnot g02772(.din(n19842), .dout(n20035));
  jnot g02773(.din(n19847), .dout(n20036));
  jnot g02774(.din(n19852), .dout(n20037));
  jnot g02775(.din(n19857), .dout(n20038));
  jnot g02776(.din(n19862), .dout(n20039));
  jnot g02777(.din(n19867), .dout(n20040));
  jnot g02778(.din(n19872), .dout(n20041));
  jnot g02779(.din(n19875), .dout(n20042));
  jxor g02780(.dina(n19876), .dinb(n259), .dout(n20043));
  jor  g02781(.dina(n20043), .dinb(n2002), .dout(n20044));
  jand g02782(.dina(n20044), .dinb(n20042), .dout(n20045));
  jnot g02783(.din(n19880), .dout(n20046));
  jor  g02784(.dina(n20046), .dinb(n20045), .dout(n20047));
  jand g02785(.dina(n20047), .dinb(n20041), .dout(n20048));
  jnot g02786(.din(n19883), .dout(n20049));
  jor  g02787(.dina(n20049), .dinb(n20048), .dout(n20050));
  jand g02788(.dina(n20050), .dinb(n20040), .dout(n20051));
  jnot g02789(.din(n19886), .dout(n20052));
  jor  g02790(.dina(n20052), .dinb(n20051), .dout(n20053));
  jand g02791(.dina(n20053), .dinb(n20039), .dout(n20054));
  jnot g02792(.din(n19889), .dout(n20055));
  jor  g02793(.dina(n20055), .dinb(n20054), .dout(n20056));
  jand g02794(.dina(n20056), .dinb(n20038), .dout(n20057));
  jnot g02795(.din(n19892), .dout(n20058));
  jor  g02796(.dina(n20058), .dinb(n20057), .dout(n20059));
  jand g02797(.dina(n20059), .dinb(n20037), .dout(n20060));
  jnot g02798(.din(n19895), .dout(n20061));
  jor  g02799(.dina(n20061), .dinb(n20060), .dout(n20062));
  jand g02800(.dina(n20062), .dinb(n20036), .dout(n20063));
  jnot g02801(.din(n19898), .dout(n20064));
  jor  g02802(.dina(n20064), .dinb(n20063), .dout(n20065));
  jand g02803(.dina(n20065), .dinb(n20035), .dout(n20066));
  jnot g02804(.din(n19901), .dout(n20067));
  jor  g02805(.dina(n20067), .dinb(n20066), .dout(n20068));
  jand g02806(.dina(n20068), .dinb(n20034), .dout(n20069));
  jnot g02807(.din(n19904), .dout(n20070));
  jor  g02808(.dina(n20070), .dinb(n20069), .dout(n20071));
  jand g02809(.dina(n20071), .dinb(n20033), .dout(n20072));
  jnot g02810(.din(n19907), .dout(n20073));
  jor  g02811(.dina(n20073), .dinb(n20072), .dout(n20074));
  jand g02812(.dina(n20074), .dinb(n20032), .dout(n20075));
  jnot g02813(.din(n19910), .dout(n20076));
  jor  g02814(.dina(n20076), .dinb(n20075), .dout(n20077));
  jand g02815(.dina(n20077), .dinb(n20031), .dout(n20078));
  jnot g02816(.din(n19913), .dout(n20079));
  jor  g02817(.dina(n20079), .dinb(n20078), .dout(n20080));
  jand g02818(.dina(n20080), .dinb(n20030), .dout(n20081));
  jnot g02819(.din(n19916), .dout(n20082));
  jor  g02820(.dina(n20082), .dinb(n20081), .dout(n20083));
  jand g02821(.dina(n20083), .dinb(n20029), .dout(n20084));
  jnot g02822(.din(n19919), .dout(n20085));
  jor  g02823(.dina(n20085), .dinb(n20084), .dout(n20086));
  jand g02824(.dina(n20086), .dinb(n20028), .dout(n20087));
  jnot g02825(.din(n19922), .dout(n20088));
  jor  g02826(.dina(n20088), .dinb(n20087), .dout(n20089));
  jand g02827(.dina(n20089), .dinb(n20027), .dout(n20090));
  jnot g02828(.din(n19925), .dout(n20091));
  jor  g02829(.dina(n20091), .dinb(n20090), .dout(n20092));
  jand g02830(.dina(n20092), .dinb(n20026), .dout(n20093));
  jor  g02831(.dina(n20093), .dinb(n19795), .dout(n20094));
  jand g02832(.dina(n20094), .dinb(n20025), .dout(n20095));
  jor  g02833(.dina(n20095), .dinb(n20024), .dout(n20096));
  jand g02834(.dina(n20096), .dinb(a45 ), .dout(n20097));
  jnot g02835(.din(n2156), .dout(n20098));
  jor  g02836(.dina(n20095), .dinb(n20098), .dout(n20099));
  jnot g02837(.din(n20099), .dout(n20100));
  jor  g02838(.dina(n20100), .dinb(n20097), .dout(n20101));
  jand g02839(.dina(n20101), .dinb(n259), .dout(n20102));
  jand g02840(.dina(n19929), .dinb(n1841), .dout(n20103));
  jor  g02841(.dina(n20103), .dinb(n2001), .dout(n20104));
  jand g02842(.dina(n20099), .dinb(n20104), .dout(n20105));
  jxor g02843(.dina(n20105), .dinb(b1 ), .dout(n20106));
  jand g02844(.dina(n20106), .dinb(n2164), .dout(n20107));
  jor  g02845(.dina(n20107), .dinb(n20102), .dout(n20108));
  jxor g02846(.dina(n20022), .dinb(n386), .dout(n20109));
  jand g02847(.dina(n20109), .dinb(n20108), .dout(n20110));
  jor  g02848(.dina(n20110), .dinb(n20023), .dout(n20111));
  jxor g02849(.dina(n20017), .dinb(n264), .dout(n20112));
  jand g02850(.dina(n20112), .dinb(n20111), .dout(n20113));
  jor  g02851(.dina(n20113), .dinb(n20018), .dout(n20114));
  jxor g02852(.dina(n20012), .dinb(n376), .dout(n20115));
  jand g02853(.dina(n20115), .dinb(n20114), .dout(n20116));
  jor  g02854(.dina(n20116), .dinb(n20013), .dout(n20117));
  jxor g02855(.dina(n20007), .dinb(n377), .dout(n20118));
  jand g02856(.dina(n20118), .dinb(n20117), .dout(n20119));
  jor  g02857(.dina(n20119), .dinb(n20008), .dout(n20120));
  jxor g02858(.dina(n20002), .dinb(n378), .dout(n20121));
  jand g02859(.dina(n20121), .dinb(n20120), .dout(n20122));
  jor  g02860(.dina(n20122), .dinb(n20003), .dout(n20123));
  jxor g02861(.dina(n19997), .dinb(n265), .dout(n20124));
  jand g02862(.dina(n20124), .dinb(n20123), .dout(n20125));
  jor  g02863(.dina(n20125), .dinb(n19998), .dout(n20126));
  jxor g02864(.dina(n19992), .dinb(n367), .dout(n20127));
  jand g02865(.dina(n20127), .dinb(n20126), .dout(n20128));
  jor  g02866(.dina(n20128), .dinb(n19993), .dout(n20129));
  jxor g02867(.dina(n19987), .dinb(n368), .dout(n20130));
  jand g02868(.dina(n20130), .dinb(n20129), .dout(n20131));
  jor  g02869(.dina(n20131), .dinb(n19988), .dout(n20132));
  jxor g02870(.dina(n19982), .dinb(n369), .dout(n20133));
  jand g02871(.dina(n20133), .dinb(n20132), .dout(n20134));
  jor  g02872(.dina(n20134), .dinb(n19983), .dout(n20135));
  jxor g02873(.dina(n19977), .dinb(n359), .dout(n20136));
  jand g02874(.dina(n20136), .dinb(n20135), .dout(n20137));
  jor  g02875(.dina(n20137), .dinb(n19978), .dout(n20138));
  jxor g02876(.dina(n19972), .dinb(n363), .dout(n20139));
  jand g02877(.dina(n20139), .dinb(n20138), .dout(n20140));
  jor  g02878(.dina(n20140), .dinb(n19973), .dout(n20141));
  jxor g02879(.dina(n19967), .dinb(n360), .dout(n20142));
  jand g02880(.dina(n20142), .dinb(n20141), .dout(n20143));
  jor  g02881(.dina(n20143), .dinb(n19968), .dout(n20144));
  jxor g02882(.dina(n19962), .dinb(n361), .dout(n20145));
  jand g02883(.dina(n20145), .dinb(n20144), .dout(n20146));
  jor  g02884(.dina(n20146), .dinb(n19963), .dout(n20147));
  jxor g02885(.dina(n19957), .dinb(n364), .dout(n20148));
  jand g02886(.dina(n20148), .dinb(n20147), .dout(n20149));
  jor  g02887(.dina(n20149), .dinb(n19958), .dout(n20150));
  jxor g02888(.dina(n19952), .dinb(n355), .dout(n20151));
  jand g02889(.dina(n20151), .dinb(n20150), .dout(n20152));
  jor  g02890(.dina(n20152), .dinb(n19953), .dout(n20153));
  jxor g02891(.dina(n19947), .dinb(n356), .dout(n20154));
  jand g02892(.dina(n20154), .dinb(n20153), .dout(n20155));
  jor  g02893(.dina(n20155), .dinb(n19948), .dout(n20156));
  jxor g02894(.dina(n19935), .dinb(n266), .dout(n20157));
  jand g02895(.dina(n20157), .dinb(n20156), .dout(n20158));
  jor  g02896(.dina(n20158), .dinb(n19943), .dout(n20159));
  jand g02897(.dina(n20159), .dinb(n19942), .dout(n20160));
  jor  g02898(.dina(n20160), .dinb(n19939), .dout(n20161));
  jand g02899(.dina(n20161), .dinb(n352), .dout(n20162));
  jor  g02900(.dina(n20162), .dinb(n19935), .dout(n20163));
  jnot g02901(.din(n20162), .dout(n20164));
  jxor g02902(.dina(n20157), .dinb(n20156), .dout(n20165));
  jor  g02903(.dina(n20165), .dinb(n20164), .dout(n20166));
  jand g02904(.dina(n20166), .dinb(n20163), .dout(n20167));
  jand g02905(.dina(n20164), .dinb(n19938), .dout(n20168));
  jand g02906(.dina(n20159), .dinb(n19939), .dout(n20169));
  jor  g02907(.dina(n20169), .dinb(n20168), .dout(n20170));
  jand g02908(.dina(n20170), .dinb(n352), .dout(n20171));
  jand g02909(.dina(n20167), .dinb(n267), .dout(n20172));
  jor  g02910(.dina(n20162), .dinb(n19947), .dout(n20173));
  jxor g02911(.dina(n20154), .dinb(n20153), .dout(n20174));
  jor  g02912(.dina(n20174), .dinb(n20164), .dout(n20175));
  jand g02913(.dina(n20175), .dinb(n20173), .dout(n20176));
  jand g02914(.dina(n20176), .dinb(n266), .dout(n20177));
  jor  g02915(.dina(n20162), .dinb(n19952), .dout(n20178));
  jxor g02916(.dina(n20151), .dinb(n20150), .dout(n20179));
  jor  g02917(.dina(n20179), .dinb(n20164), .dout(n20180));
  jand g02918(.dina(n20180), .dinb(n20178), .dout(n20181));
  jand g02919(.dina(n20181), .dinb(n356), .dout(n20182));
  jor  g02920(.dina(n20162), .dinb(n19957), .dout(n20183));
  jxor g02921(.dina(n20148), .dinb(n20147), .dout(n20184));
  jor  g02922(.dina(n20184), .dinb(n20164), .dout(n20185));
  jand g02923(.dina(n20185), .dinb(n20183), .dout(n20186));
  jand g02924(.dina(n20186), .dinb(n355), .dout(n20187));
  jor  g02925(.dina(n20162), .dinb(n19962), .dout(n20188));
  jxor g02926(.dina(n20145), .dinb(n20144), .dout(n20189));
  jor  g02927(.dina(n20189), .dinb(n20164), .dout(n20190));
  jand g02928(.dina(n20190), .dinb(n20188), .dout(n20191));
  jand g02929(.dina(n20191), .dinb(n364), .dout(n20192));
  jor  g02930(.dina(n20162), .dinb(n19967), .dout(n20193));
  jxor g02931(.dina(n20142), .dinb(n20141), .dout(n20194));
  jor  g02932(.dina(n20194), .dinb(n20164), .dout(n20195));
  jand g02933(.dina(n20195), .dinb(n20193), .dout(n20196));
  jand g02934(.dina(n20196), .dinb(n361), .dout(n20197));
  jor  g02935(.dina(n20162), .dinb(n19972), .dout(n20198));
  jxor g02936(.dina(n20139), .dinb(n20138), .dout(n20199));
  jor  g02937(.dina(n20199), .dinb(n20164), .dout(n20200));
  jand g02938(.dina(n20200), .dinb(n20198), .dout(n20201));
  jand g02939(.dina(n20201), .dinb(n360), .dout(n20202));
  jor  g02940(.dina(n20162), .dinb(n19977), .dout(n20203));
  jxor g02941(.dina(n20136), .dinb(n20135), .dout(n20204));
  jor  g02942(.dina(n20204), .dinb(n20164), .dout(n20205));
  jand g02943(.dina(n20205), .dinb(n20203), .dout(n20206));
  jand g02944(.dina(n20206), .dinb(n363), .dout(n20207));
  jor  g02945(.dina(n20162), .dinb(n19982), .dout(n20208));
  jxor g02946(.dina(n20133), .dinb(n20132), .dout(n20209));
  jor  g02947(.dina(n20209), .dinb(n20164), .dout(n20210));
  jand g02948(.dina(n20210), .dinb(n20208), .dout(n20211));
  jand g02949(.dina(n20211), .dinb(n359), .dout(n20212));
  jor  g02950(.dina(n20162), .dinb(n19987), .dout(n20213));
  jxor g02951(.dina(n20130), .dinb(n20129), .dout(n20214));
  jor  g02952(.dina(n20214), .dinb(n20164), .dout(n20215));
  jand g02953(.dina(n20215), .dinb(n20213), .dout(n20216));
  jand g02954(.dina(n20216), .dinb(n369), .dout(n20217));
  jor  g02955(.dina(n20162), .dinb(n19992), .dout(n20218));
  jxor g02956(.dina(n20127), .dinb(n20126), .dout(n20219));
  jor  g02957(.dina(n20219), .dinb(n20164), .dout(n20220));
  jand g02958(.dina(n20220), .dinb(n20218), .dout(n20221));
  jand g02959(.dina(n20221), .dinb(n368), .dout(n20222));
  jor  g02960(.dina(n20162), .dinb(n19997), .dout(n20223));
  jxor g02961(.dina(n20124), .dinb(n20123), .dout(n20224));
  jor  g02962(.dina(n20224), .dinb(n20164), .dout(n20225));
  jand g02963(.dina(n20225), .dinb(n20223), .dout(n20226));
  jand g02964(.dina(n20226), .dinb(n367), .dout(n20227));
  jor  g02965(.dina(n20162), .dinb(n20002), .dout(n20228));
  jxor g02966(.dina(n20121), .dinb(n20120), .dout(n20229));
  jor  g02967(.dina(n20229), .dinb(n20164), .dout(n20230));
  jand g02968(.dina(n20230), .dinb(n20228), .dout(n20231));
  jand g02969(.dina(n20231), .dinb(n265), .dout(n20232));
  jor  g02970(.dina(n20162), .dinb(n20007), .dout(n20233));
  jxor g02971(.dina(n20118), .dinb(n20117), .dout(n20234));
  jor  g02972(.dina(n20234), .dinb(n20164), .dout(n20235));
  jand g02973(.dina(n20235), .dinb(n20233), .dout(n20236));
  jand g02974(.dina(n20236), .dinb(n378), .dout(n20237));
  jor  g02975(.dina(n20162), .dinb(n20012), .dout(n20238));
  jxor g02976(.dina(n20115), .dinb(n20114), .dout(n20239));
  jor  g02977(.dina(n20239), .dinb(n20164), .dout(n20240));
  jand g02978(.dina(n20240), .dinb(n20238), .dout(n20241));
  jand g02979(.dina(n20241), .dinb(n377), .dout(n20242));
  jor  g02980(.dina(n20162), .dinb(n20017), .dout(n20243));
  jxor g02981(.dina(n20112), .dinb(n20111), .dout(n20244));
  jor  g02982(.dina(n20244), .dinb(n20164), .dout(n20245));
  jand g02983(.dina(n20245), .dinb(n20243), .dout(n20246));
  jand g02984(.dina(n20246), .dinb(n376), .dout(n20247));
  jor  g02985(.dina(n20162), .dinb(n20022), .dout(n20248));
  jxor g02986(.dina(n20109), .dinb(n20108), .dout(n20249));
  jor  g02987(.dina(n20249), .dinb(n20164), .dout(n20250));
  jand g02988(.dina(n20250), .dinb(n20248), .dout(n20251));
  jand g02989(.dina(n20251), .dinb(n264), .dout(n20252));
  jor  g02990(.dina(n20162), .dinb(n20105), .dout(n20253));
  jxor g02991(.dina(n20106), .dinb(n2164), .dout(n20254));
  jand g02992(.dina(n20254), .dinb(n20162), .dout(n20255));
  jnot g02993(.din(n20255), .dout(n20256));
  jand g02994(.dina(n20256), .dinb(n20253), .dout(n20257));
  jnot g02995(.din(n20257), .dout(n20258));
  jand g02996(.dina(n20258), .dinb(n386), .dout(n20259));
  jnot g02997(.din(n2316), .dout(n20260));
  jnot g02998(.din(n19939), .dout(n20261));
  jnot g02999(.din(n19943), .dout(n20262));
  jnot g03000(.din(n19948), .dout(n20263));
  jnot g03001(.din(n19953), .dout(n20264));
  jnot g03002(.din(n19958), .dout(n20265));
  jnot g03003(.din(n19963), .dout(n20266));
  jnot g03004(.din(n19968), .dout(n20267));
  jnot g03005(.din(n19973), .dout(n20268));
  jnot g03006(.din(n19978), .dout(n20269));
  jnot g03007(.din(n19983), .dout(n20270));
  jnot g03008(.din(n19988), .dout(n20271));
  jnot g03009(.din(n19993), .dout(n20272));
  jnot g03010(.din(n19998), .dout(n20273));
  jnot g03011(.din(n20003), .dout(n20274));
  jnot g03012(.din(n20008), .dout(n20275));
  jnot g03013(.din(n20013), .dout(n20276));
  jnot g03014(.din(n20018), .dout(n20277));
  jnot g03015(.din(n20023), .dout(n20278));
  jnot g03016(.din(n20102), .dout(n20279));
  jxor g03017(.dina(n20105), .dinb(n259), .dout(n20280));
  jor  g03018(.dina(n20280), .dinb(n2163), .dout(n20281));
  jand g03019(.dina(n20281), .dinb(n20279), .dout(n20282));
  jnot g03020(.din(n20109), .dout(n20283));
  jor  g03021(.dina(n20283), .dinb(n20282), .dout(n20284));
  jand g03022(.dina(n20284), .dinb(n20278), .dout(n20285));
  jnot g03023(.din(n20112), .dout(n20286));
  jor  g03024(.dina(n20286), .dinb(n20285), .dout(n20287));
  jand g03025(.dina(n20287), .dinb(n20277), .dout(n20288));
  jnot g03026(.din(n20115), .dout(n20289));
  jor  g03027(.dina(n20289), .dinb(n20288), .dout(n20290));
  jand g03028(.dina(n20290), .dinb(n20276), .dout(n20291));
  jnot g03029(.din(n20118), .dout(n20292));
  jor  g03030(.dina(n20292), .dinb(n20291), .dout(n20293));
  jand g03031(.dina(n20293), .dinb(n20275), .dout(n20294));
  jnot g03032(.din(n20121), .dout(n20295));
  jor  g03033(.dina(n20295), .dinb(n20294), .dout(n20296));
  jand g03034(.dina(n20296), .dinb(n20274), .dout(n20297));
  jnot g03035(.din(n20124), .dout(n20298));
  jor  g03036(.dina(n20298), .dinb(n20297), .dout(n20299));
  jand g03037(.dina(n20299), .dinb(n20273), .dout(n20300));
  jnot g03038(.din(n20127), .dout(n20301));
  jor  g03039(.dina(n20301), .dinb(n20300), .dout(n20302));
  jand g03040(.dina(n20302), .dinb(n20272), .dout(n20303));
  jnot g03041(.din(n20130), .dout(n20304));
  jor  g03042(.dina(n20304), .dinb(n20303), .dout(n20305));
  jand g03043(.dina(n20305), .dinb(n20271), .dout(n20306));
  jnot g03044(.din(n20133), .dout(n20307));
  jor  g03045(.dina(n20307), .dinb(n20306), .dout(n20308));
  jand g03046(.dina(n20308), .dinb(n20270), .dout(n20309));
  jnot g03047(.din(n20136), .dout(n20310));
  jor  g03048(.dina(n20310), .dinb(n20309), .dout(n20311));
  jand g03049(.dina(n20311), .dinb(n20269), .dout(n20312));
  jnot g03050(.din(n20139), .dout(n20313));
  jor  g03051(.dina(n20313), .dinb(n20312), .dout(n20314));
  jand g03052(.dina(n20314), .dinb(n20268), .dout(n20315));
  jnot g03053(.din(n20142), .dout(n20316));
  jor  g03054(.dina(n20316), .dinb(n20315), .dout(n20317));
  jand g03055(.dina(n20317), .dinb(n20267), .dout(n20318));
  jnot g03056(.din(n20145), .dout(n20319));
  jor  g03057(.dina(n20319), .dinb(n20318), .dout(n20320));
  jand g03058(.dina(n20320), .dinb(n20266), .dout(n20321));
  jnot g03059(.din(n20148), .dout(n20322));
  jor  g03060(.dina(n20322), .dinb(n20321), .dout(n20323));
  jand g03061(.dina(n20323), .dinb(n20265), .dout(n20324));
  jnot g03062(.din(n20151), .dout(n20325));
  jor  g03063(.dina(n20325), .dinb(n20324), .dout(n20326));
  jand g03064(.dina(n20326), .dinb(n20264), .dout(n20327));
  jnot g03065(.din(n20154), .dout(n20328));
  jor  g03066(.dina(n20328), .dinb(n20327), .dout(n20329));
  jand g03067(.dina(n20329), .dinb(n20263), .dout(n20330));
  jnot g03068(.din(n20157), .dout(n20331));
  jor  g03069(.dina(n20331), .dinb(n20330), .dout(n20332));
  jand g03070(.dina(n20332), .dinb(n20262), .dout(n20333));
  jor  g03071(.dina(n20333), .dinb(n19941), .dout(n20334));
  jand g03072(.dina(n20334), .dinb(n20261), .dout(n20335));
  jor  g03073(.dina(n20335), .dinb(n20260), .dout(n20336));
  jand g03074(.dina(n20336), .dinb(a44 ), .dout(n20337));
  jnot g03075(.din(n2319), .dout(n20338));
  jor  g03076(.dina(n20335), .dinb(n20338), .dout(n20339));
  jnot g03077(.din(n20339), .dout(n20340));
  jor  g03078(.dina(n20340), .dinb(n20337), .dout(n20341));
  jand g03079(.dina(n20341), .dinb(n259), .dout(n20342));
  jand g03080(.dina(n20161), .dinb(n2316), .dout(n20343));
  jor  g03081(.dina(n20343), .dinb(n2162), .dout(n20344));
  jand g03082(.dina(n20339), .dinb(n20344), .dout(n20345));
  jxor g03083(.dina(n20345), .dinb(b1 ), .dout(n20346));
  jand g03084(.dina(n20346), .dinb(n2327), .dout(n20347));
  jor  g03085(.dina(n20347), .dinb(n20342), .dout(n20348));
  jxor g03086(.dina(n20257), .dinb(b2 ), .dout(n20349));
  jand g03087(.dina(n20349), .dinb(n20348), .dout(n20350));
  jor  g03088(.dina(n20350), .dinb(n20259), .dout(n20351));
  jxor g03089(.dina(n20251), .dinb(n264), .dout(n20352));
  jand g03090(.dina(n20352), .dinb(n20351), .dout(n20353));
  jor  g03091(.dina(n20353), .dinb(n20252), .dout(n20354));
  jxor g03092(.dina(n20246), .dinb(n376), .dout(n20355));
  jand g03093(.dina(n20355), .dinb(n20354), .dout(n20356));
  jor  g03094(.dina(n20356), .dinb(n20247), .dout(n20357));
  jxor g03095(.dina(n20241), .dinb(n377), .dout(n20358));
  jand g03096(.dina(n20358), .dinb(n20357), .dout(n20359));
  jor  g03097(.dina(n20359), .dinb(n20242), .dout(n20360));
  jxor g03098(.dina(n20236), .dinb(n378), .dout(n20361));
  jand g03099(.dina(n20361), .dinb(n20360), .dout(n20362));
  jor  g03100(.dina(n20362), .dinb(n20237), .dout(n20363));
  jxor g03101(.dina(n20231), .dinb(n265), .dout(n20364));
  jand g03102(.dina(n20364), .dinb(n20363), .dout(n20365));
  jor  g03103(.dina(n20365), .dinb(n20232), .dout(n20366));
  jxor g03104(.dina(n20226), .dinb(n367), .dout(n20367));
  jand g03105(.dina(n20367), .dinb(n20366), .dout(n20368));
  jor  g03106(.dina(n20368), .dinb(n20227), .dout(n20369));
  jxor g03107(.dina(n20221), .dinb(n368), .dout(n20370));
  jand g03108(.dina(n20370), .dinb(n20369), .dout(n20371));
  jor  g03109(.dina(n20371), .dinb(n20222), .dout(n20372));
  jxor g03110(.dina(n20216), .dinb(n369), .dout(n20373));
  jand g03111(.dina(n20373), .dinb(n20372), .dout(n20374));
  jor  g03112(.dina(n20374), .dinb(n20217), .dout(n20375));
  jxor g03113(.dina(n20211), .dinb(n359), .dout(n20376));
  jand g03114(.dina(n20376), .dinb(n20375), .dout(n20377));
  jor  g03115(.dina(n20377), .dinb(n20212), .dout(n20378));
  jxor g03116(.dina(n20206), .dinb(n363), .dout(n20379));
  jand g03117(.dina(n20379), .dinb(n20378), .dout(n20380));
  jor  g03118(.dina(n20380), .dinb(n20207), .dout(n20381));
  jxor g03119(.dina(n20201), .dinb(n360), .dout(n20382));
  jand g03120(.dina(n20382), .dinb(n20381), .dout(n20383));
  jor  g03121(.dina(n20383), .dinb(n20202), .dout(n20384));
  jxor g03122(.dina(n20196), .dinb(n361), .dout(n20385));
  jand g03123(.dina(n20385), .dinb(n20384), .dout(n20386));
  jor  g03124(.dina(n20386), .dinb(n20197), .dout(n20387));
  jxor g03125(.dina(n20191), .dinb(n364), .dout(n20388));
  jand g03126(.dina(n20388), .dinb(n20387), .dout(n20389));
  jor  g03127(.dina(n20389), .dinb(n20192), .dout(n20390));
  jxor g03128(.dina(n20186), .dinb(n355), .dout(n20391));
  jand g03129(.dina(n20391), .dinb(n20390), .dout(n20392));
  jor  g03130(.dina(n20392), .dinb(n20187), .dout(n20393));
  jxor g03131(.dina(n20181), .dinb(n356), .dout(n20394));
  jand g03132(.dina(n20394), .dinb(n20393), .dout(n20395));
  jor  g03133(.dina(n20395), .dinb(n20182), .dout(n20396));
  jxor g03134(.dina(n20176), .dinb(n266), .dout(n20397));
  jand g03135(.dina(n20397), .dinb(n20396), .dout(n20398));
  jor  g03136(.dina(n20398), .dinb(n20177), .dout(n20399));
  jxor g03137(.dina(n20167), .dinb(n267), .dout(n20400));
  jand g03138(.dina(n20400), .dinb(n20399), .dout(n20401));
  jor  g03139(.dina(n20401), .dinb(n20172), .dout(n20402));
  jnot g03140(.din(n418), .dout(n20403));
  jxor g03141(.dina(n20170), .dinb(b20 ), .dout(n20404));
  jor  g03142(.dina(n20404), .dinb(n20403), .dout(n20405));
  jnot g03143(.din(n20405), .dout(n20406));
  jand g03144(.dina(n20406), .dinb(n20402), .dout(n20407));
  jor  g03145(.dina(n20407), .dinb(n20171), .dout(n20408));
  jor  g03146(.dina(n20408), .dinb(n20167), .dout(n20409));
  jnot g03147(.din(n20408), .dout(n20410));
  jxor g03148(.dina(n20400), .dinb(n20399), .dout(n20411));
  jor  g03149(.dina(n20411), .dinb(n20410), .dout(n20412));
  jand g03150(.dina(n20412), .dinb(n20409), .dout(n20413));
  jand g03151(.dina(n20410), .dinb(n20170), .dout(n20414));
  jnot g03152(.din(n20404), .dout(n20415));
  jxor g03153(.dina(n20415), .dinb(n20402), .dout(n20416));
  jand g03154(.dina(n20416), .dinb(n20171), .dout(n20417));
  jor  g03155(.dina(n20417), .dinb(n20414), .dout(n20418));
  jand g03156(.dina(n20418), .dinb(n348), .dout(n20419));
  jnot g03157(.din(n20418), .dout(n20420));
  jand g03158(.dina(n20420), .dinb(b21 ), .dout(n20421));
  jnot g03159(.din(n20421), .dout(n20422));
  jand g03160(.dina(n20413), .dinb(n347), .dout(n20423));
  jor  g03161(.dina(n20408), .dinb(n20176), .dout(n20424));
  jxor g03162(.dina(n20397), .dinb(n20396), .dout(n20425));
  jor  g03163(.dina(n20425), .dinb(n20410), .dout(n20426));
  jand g03164(.dina(n20426), .dinb(n20424), .dout(n20427));
  jand g03165(.dina(n20427), .dinb(n267), .dout(n20428));
  jor  g03166(.dina(n20408), .dinb(n20181), .dout(n20429));
  jxor g03167(.dina(n20394), .dinb(n20393), .dout(n20430));
  jor  g03168(.dina(n20430), .dinb(n20410), .dout(n20431));
  jand g03169(.dina(n20431), .dinb(n20429), .dout(n20432));
  jand g03170(.dina(n20432), .dinb(n266), .dout(n20433));
  jor  g03171(.dina(n20408), .dinb(n20186), .dout(n20434));
  jxor g03172(.dina(n20391), .dinb(n20390), .dout(n20435));
  jor  g03173(.dina(n20435), .dinb(n20410), .dout(n20436));
  jand g03174(.dina(n20436), .dinb(n20434), .dout(n20437));
  jand g03175(.dina(n20437), .dinb(n356), .dout(n20438));
  jor  g03176(.dina(n20408), .dinb(n20191), .dout(n20439));
  jxor g03177(.dina(n20388), .dinb(n20387), .dout(n20440));
  jor  g03178(.dina(n20440), .dinb(n20410), .dout(n20441));
  jand g03179(.dina(n20441), .dinb(n20439), .dout(n20442));
  jand g03180(.dina(n20442), .dinb(n355), .dout(n20443));
  jor  g03181(.dina(n20408), .dinb(n20196), .dout(n20444));
  jxor g03182(.dina(n20385), .dinb(n20384), .dout(n20445));
  jor  g03183(.dina(n20445), .dinb(n20410), .dout(n20446));
  jand g03184(.dina(n20446), .dinb(n20444), .dout(n20447));
  jand g03185(.dina(n20447), .dinb(n364), .dout(n20448));
  jor  g03186(.dina(n20408), .dinb(n20201), .dout(n20449));
  jxor g03187(.dina(n20382), .dinb(n20381), .dout(n20450));
  jor  g03188(.dina(n20450), .dinb(n20410), .dout(n20451));
  jand g03189(.dina(n20451), .dinb(n20449), .dout(n20452));
  jand g03190(.dina(n20452), .dinb(n361), .dout(n20453));
  jor  g03191(.dina(n20408), .dinb(n20206), .dout(n20454));
  jxor g03192(.dina(n20379), .dinb(n20378), .dout(n20455));
  jor  g03193(.dina(n20455), .dinb(n20410), .dout(n20456));
  jand g03194(.dina(n20456), .dinb(n20454), .dout(n20457));
  jand g03195(.dina(n20457), .dinb(n360), .dout(n20458));
  jor  g03196(.dina(n20408), .dinb(n20211), .dout(n20459));
  jxor g03197(.dina(n20376), .dinb(n20375), .dout(n20460));
  jor  g03198(.dina(n20460), .dinb(n20410), .dout(n20461));
  jand g03199(.dina(n20461), .dinb(n20459), .dout(n20462));
  jand g03200(.dina(n20462), .dinb(n363), .dout(n20463));
  jor  g03201(.dina(n20408), .dinb(n20216), .dout(n20464));
  jxor g03202(.dina(n20373), .dinb(n20372), .dout(n20465));
  jor  g03203(.dina(n20465), .dinb(n20410), .dout(n20466));
  jand g03204(.dina(n20466), .dinb(n20464), .dout(n20467));
  jand g03205(.dina(n20467), .dinb(n359), .dout(n20468));
  jor  g03206(.dina(n20408), .dinb(n20221), .dout(n20469));
  jxor g03207(.dina(n20370), .dinb(n20369), .dout(n20470));
  jor  g03208(.dina(n20470), .dinb(n20410), .dout(n20471));
  jand g03209(.dina(n20471), .dinb(n20469), .dout(n20472));
  jand g03210(.dina(n20472), .dinb(n369), .dout(n20473));
  jor  g03211(.dina(n20408), .dinb(n20226), .dout(n20474));
  jxor g03212(.dina(n20367), .dinb(n20366), .dout(n20475));
  jor  g03213(.dina(n20475), .dinb(n20410), .dout(n20476));
  jand g03214(.dina(n20476), .dinb(n20474), .dout(n20477));
  jand g03215(.dina(n20477), .dinb(n368), .dout(n20478));
  jor  g03216(.dina(n20408), .dinb(n20231), .dout(n20479));
  jxor g03217(.dina(n20364), .dinb(n20363), .dout(n20480));
  jor  g03218(.dina(n20480), .dinb(n20410), .dout(n20481));
  jand g03219(.dina(n20481), .dinb(n20479), .dout(n20482));
  jand g03220(.dina(n20482), .dinb(n367), .dout(n20483));
  jor  g03221(.dina(n20408), .dinb(n20236), .dout(n20484));
  jxor g03222(.dina(n20361), .dinb(n20360), .dout(n20485));
  jor  g03223(.dina(n20485), .dinb(n20410), .dout(n20486));
  jand g03224(.dina(n20486), .dinb(n20484), .dout(n20487));
  jand g03225(.dina(n20487), .dinb(n265), .dout(n20488));
  jor  g03226(.dina(n20408), .dinb(n20241), .dout(n20489));
  jxor g03227(.dina(n20358), .dinb(n20357), .dout(n20490));
  jor  g03228(.dina(n20490), .dinb(n20410), .dout(n20491));
  jand g03229(.dina(n20491), .dinb(n20489), .dout(n20492));
  jand g03230(.dina(n20492), .dinb(n378), .dout(n20493));
  jor  g03231(.dina(n20408), .dinb(n20246), .dout(n20494));
  jxor g03232(.dina(n20355), .dinb(n20354), .dout(n20495));
  jor  g03233(.dina(n20495), .dinb(n20410), .dout(n20496));
  jand g03234(.dina(n20496), .dinb(n20494), .dout(n20497));
  jand g03235(.dina(n20497), .dinb(n377), .dout(n20498));
  jor  g03236(.dina(n20408), .dinb(n20251), .dout(n20499));
  jxor g03237(.dina(n20352), .dinb(n20351), .dout(n20500));
  jor  g03238(.dina(n20500), .dinb(n20410), .dout(n20501));
  jand g03239(.dina(n20501), .dinb(n20499), .dout(n20502));
  jand g03240(.dina(n20502), .dinb(n376), .dout(n20503));
  jor  g03241(.dina(n20408), .dinb(n20258), .dout(n20504));
  jxor g03242(.dina(n20349), .dinb(n20348), .dout(n20505));
  jor  g03243(.dina(n20505), .dinb(n20410), .dout(n20506));
  jand g03244(.dina(n20506), .dinb(n20504), .dout(n20507));
  jand g03245(.dina(n20507), .dinb(n264), .dout(n20508));
  jor  g03246(.dina(n20408), .dinb(n20341), .dout(n20509));
  jxor g03247(.dina(n20346), .dinb(n2327), .dout(n20510));
  jor  g03248(.dina(n20510), .dinb(n20410), .dout(n20511));
  jand g03249(.dina(n20511), .dinb(n20509), .dout(n20512));
  jand g03250(.dina(n20512), .dinb(n386), .dout(n20513));
  jand g03251(.dina(n20408), .dinb(b0 ), .dout(n20514));
  jxor g03252(.dina(n20514), .dinb(a43 ), .dout(n20515));
  jand g03253(.dina(n20515), .dinb(n259), .dout(n20516));
  jxor g03254(.dina(n20514), .dinb(n2325), .dout(n20517));
  jxor g03255(.dina(n20517), .dinb(b1 ), .dout(n20518));
  jand g03256(.dina(n20518), .dinb(n2505), .dout(n20519));
  jor  g03257(.dina(n20519), .dinb(n20516), .dout(n20520));
  jxor g03258(.dina(n20512), .dinb(n386), .dout(n20521));
  jand g03259(.dina(n20521), .dinb(n20520), .dout(n20522));
  jor  g03260(.dina(n20522), .dinb(n20513), .dout(n20523));
  jxor g03261(.dina(n20507), .dinb(n264), .dout(n20524));
  jand g03262(.dina(n20524), .dinb(n20523), .dout(n20525));
  jor  g03263(.dina(n20525), .dinb(n20508), .dout(n20526));
  jxor g03264(.dina(n20502), .dinb(n376), .dout(n20527));
  jand g03265(.dina(n20527), .dinb(n20526), .dout(n20528));
  jor  g03266(.dina(n20528), .dinb(n20503), .dout(n20529));
  jxor g03267(.dina(n20497), .dinb(n377), .dout(n20530));
  jand g03268(.dina(n20530), .dinb(n20529), .dout(n20531));
  jor  g03269(.dina(n20531), .dinb(n20498), .dout(n20532));
  jxor g03270(.dina(n20492), .dinb(n378), .dout(n20533));
  jand g03271(.dina(n20533), .dinb(n20532), .dout(n20534));
  jor  g03272(.dina(n20534), .dinb(n20493), .dout(n20535));
  jxor g03273(.dina(n20487), .dinb(n265), .dout(n20536));
  jand g03274(.dina(n20536), .dinb(n20535), .dout(n20537));
  jor  g03275(.dina(n20537), .dinb(n20488), .dout(n20538));
  jxor g03276(.dina(n20482), .dinb(n367), .dout(n20539));
  jand g03277(.dina(n20539), .dinb(n20538), .dout(n20540));
  jor  g03278(.dina(n20540), .dinb(n20483), .dout(n20541));
  jxor g03279(.dina(n20477), .dinb(n368), .dout(n20542));
  jand g03280(.dina(n20542), .dinb(n20541), .dout(n20543));
  jor  g03281(.dina(n20543), .dinb(n20478), .dout(n20544));
  jxor g03282(.dina(n20472), .dinb(n369), .dout(n20545));
  jand g03283(.dina(n20545), .dinb(n20544), .dout(n20546));
  jor  g03284(.dina(n20546), .dinb(n20473), .dout(n20547));
  jxor g03285(.dina(n20467), .dinb(n359), .dout(n20548));
  jand g03286(.dina(n20548), .dinb(n20547), .dout(n20549));
  jor  g03287(.dina(n20549), .dinb(n20468), .dout(n20550));
  jxor g03288(.dina(n20462), .dinb(n363), .dout(n20551));
  jand g03289(.dina(n20551), .dinb(n20550), .dout(n20552));
  jor  g03290(.dina(n20552), .dinb(n20463), .dout(n20553));
  jxor g03291(.dina(n20457), .dinb(n360), .dout(n20554));
  jand g03292(.dina(n20554), .dinb(n20553), .dout(n20555));
  jor  g03293(.dina(n20555), .dinb(n20458), .dout(n20556));
  jxor g03294(.dina(n20452), .dinb(n361), .dout(n20557));
  jand g03295(.dina(n20557), .dinb(n20556), .dout(n20558));
  jor  g03296(.dina(n20558), .dinb(n20453), .dout(n20559));
  jxor g03297(.dina(n20447), .dinb(n364), .dout(n20560));
  jand g03298(.dina(n20560), .dinb(n20559), .dout(n20561));
  jor  g03299(.dina(n20561), .dinb(n20448), .dout(n20562));
  jxor g03300(.dina(n20442), .dinb(n355), .dout(n20563));
  jand g03301(.dina(n20563), .dinb(n20562), .dout(n20564));
  jor  g03302(.dina(n20564), .dinb(n20443), .dout(n20565));
  jxor g03303(.dina(n20437), .dinb(n356), .dout(n20566));
  jand g03304(.dina(n20566), .dinb(n20565), .dout(n20567));
  jor  g03305(.dina(n20567), .dinb(n20438), .dout(n20568));
  jxor g03306(.dina(n20432), .dinb(n266), .dout(n20569));
  jand g03307(.dina(n20569), .dinb(n20568), .dout(n20570));
  jor  g03308(.dina(n20570), .dinb(n20433), .dout(n20571));
  jxor g03309(.dina(n20427), .dinb(n267), .dout(n20572));
  jand g03310(.dina(n20572), .dinb(n20571), .dout(n20573));
  jor  g03311(.dina(n20573), .dinb(n20428), .dout(n20574));
  jxor g03312(.dina(n20413), .dinb(n347), .dout(n20575));
  jand g03313(.dina(n20575), .dinb(n20574), .dout(n20576));
  jor  g03314(.dina(n20576), .dinb(n20423), .dout(n20577));
  jand g03315(.dina(n20577), .dinb(n20422), .dout(n20578));
  jor  g03316(.dina(n20578), .dinb(n20419), .dout(n20579));
  jand g03317(.dina(n20579), .dinb(n2680), .dout(n20580));
  jor  g03318(.dina(n20580), .dinb(n20413), .dout(n20581));
  jnot g03319(.din(n20580), .dout(n20582));
  jxor g03320(.dina(n20575), .dinb(n20574), .dout(n20583));
  jor  g03321(.dina(n20583), .dinb(n20582), .dout(n20584));
  jand g03322(.dina(n20584), .dinb(n20581), .dout(n20585));
  jand g03323(.dina(n20582), .dinb(n20418), .dout(n20586));
  jand g03324(.dina(n20577), .dinb(n20419), .dout(n20587));
  jor  g03325(.dina(n20587), .dinb(n20586), .dout(n20588));
  jand g03326(.dina(n20588), .dinb(n349), .dout(n20589));
  jnot g03327(.din(n20588), .dout(n20590));
  jand g03328(.dina(n20590), .dinb(b22 ), .dout(n20591));
  jnot g03329(.din(n20591), .dout(n20592));
  jand g03330(.dina(n20585), .dinb(n348), .dout(n20593));
  jor  g03331(.dina(n20580), .dinb(n20427), .dout(n20594));
  jxor g03332(.dina(n20572), .dinb(n20571), .dout(n20595));
  jor  g03333(.dina(n20595), .dinb(n20582), .dout(n20596));
  jand g03334(.dina(n20596), .dinb(n20594), .dout(n20597));
  jand g03335(.dina(n20597), .dinb(n347), .dout(n20598));
  jor  g03336(.dina(n20580), .dinb(n20432), .dout(n20599));
  jxor g03337(.dina(n20569), .dinb(n20568), .dout(n20600));
  jor  g03338(.dina(n20600), .dinb(n20582), .dout(n20601));
  jand g03339(.dina(n20601), .dinb(n20599), .dout(n20602));
  jand g03340(.dina(n20602), .dinb(n267), .dout(n20603));
  jor  g03341(.dina(n20580), .dinb(n20437), .dout(n20604));
  jxor g03342(.dina(n20566), .dinb(n20565), .dout(n20605));
  jor  g03343(.dina(n20605), .dinb(n20582), .dout(n20606));
  jand g03344(.dina(n20606), .dinb(n20604), .dout(n20607));
  jand g03345(.dina(n20607), .dinb(n266), .dout(n20608));
  jor  g03346(.dina(n20580), .dinb(n20442), .dout(n20609));
  jxor g03347(.dina(n20563), .dinb(n20562), .dout(n20610));
  jor  g03348(.dina(n20610), .dinb(n20582), .dout(n20611));
  jand g03349(.dina(n20611), .dinb(n20609), .dout(n20612));
  jand g03350(.dina(n20612), .dinb(n356), .dout(n20613));
  jor  g03351(.dina(n20580), .dinb(n20447), .dout(n20614));
  jxor g03352(.dina(n20560), .dinb(n20559), .dout(n20615));
  jor  g03353(.dina(n20615), .dinb(n20582), .dout(n20616));
  jand g03354(.dina(n20616), .dinb(n20614), .dout(n20617));
  jand g03355(.dina(n20617), .dinb(n355), .dout(n20618));
  jor  g03356(.dina(n20580), .dinb(n20452), .dout(n20619));
  jxor g03357(.dina(n20557), .dinb(n20556), .dout(n20620));
  jor  g03358(.dina(n20620), .dinb(n20582), .dout(n20621));
  jand g03359(.dina(n20621), .dinb(n20619), .dout(n20622));
  jand g03360(.dina(n20622), .dinb(n364), .dout(n20623));
  jor  g03361(.dina(n20580), .dinb(n20457), .dout(n20624));
  jxor g03362(.dina(n20554), .dinb(n20553), .dout(n20625));
  jor  g03363(.dina(n20625), .dinb(n20582), .dout(n20626));
  jand g03364(.dina(n20626), .dinb(n20624), .dout(n20627));
  jand g03365(.dina(n20627), .dinb(n361), .dout(n20628));
  jor  g03366(.dina(n20580), .dinb(n20462), .dout(n20629));
  jxor g03367(.dina(n20551), .dinb(n20550), .dout(n20630));
  jor  g03368(.dina(n20630), .dinb(n20582), .dout(n20631));
  jand g03369(.dina(n20631), .dinb(n20629), .dout(n20632));
  jand g03370(.dina(n20632), .dinb(n360), .dout(n20633));
  jor  g03371(.dina(n20580), .dinb(n20467), .dout(n20634));
  jxor g03372(.dina(n20548), .dinb(n20547), .dout(n20635));
  jor  g03373(.dina(n20635), .dinb(n20582), .dout(n20636));
  jand g03374(.dina(n20636), .dinb(n20634), .dout(n20637));
  jand g03375(.dina(n20637), .dinb(n363), .dout(n20638));
  jor  g03376(.dina(n20580), .dinb(n20472), .dout(n20639));
  jxor g03377(.dina(n20545), .dinb(n20544), .dout(n20640));
  jor  g03378(.dina(n20640), .dinb(n20582), .dout(n20641));
  jand g03379(.dina(n20641), .dinb(n20639), .dout(n20642));
  jand g03380(.dina(n20642), .dinb(n359), .dout(n20643));
  jor  g03381(.dina(n20580), .dinb(n20477), .dout(n20644));
  jxor g03382(.dina(n20542), .dinb(n20541), .dout(n20645));
  jor  g03383(.dina(n20645), .dinb(n20582), .dout(n20646));
  jand g03384(.dina(n20646), .dinb(n20644), .dout(n20647));
  jand g03385(.dina(n20647), .dinb(n369), .dout(n20648));
  jor  g03386(.dina(n20580), .dinb(n20482), .dout(n20649));
  jxor g03387(.dina(n20539), .dinb(n20538), .dout(n20650));
  jor  g03388(.dina(n20650), .dinb(n20582), .dout(n20651));
  jand g03389(.dina(n20651), .dinb(n20649), .dout(n20652));
  jand g03390(.dina(n20652), .dinb(n368), .dout(n20653));
  jor  g03391(.dina(n20580), .dinb(n20487), .dout(n20654));
  jxor g03392(.dina(n20536), .dinb(n20535), .dout(n20655));
  jor  g03393(.dina(n20655), .dinb(n20582), .dout(n20656));
  jand g03394(.dina(n20656), .dinb(n20654), .dout(n20657));
  jand g03395(.dina(n20657), .dinb(n367), .dout(n20658));
  jor  g03396(.dina(n20580), .dinb(n20492), .dout(n20659));
  jxor g03397(.dina(n20533), .dinb(n20532), .dout(n20660));
  jor  g03398(.dina(n20660), .dinb(n20582), .dout(n20661));
  jand g03399(.dina(n20661), .dinb(n20659), .dout(n20662));
  jand g03400(.dina(n20662), .dinb(n265), .dout(n20663));
  jor  g03401(.dina(n20580), .dinb(n20497), .dout(n20664));
  jxor g03402(.dina(n20530), .dinb(n20529), .dout(n20665));
  jor  g03403(.dina(n20665), .dinb(n20582), .dout(n20666));
  jand g03404(.dina(n20666), .dinb(n20664), .dout(n20667));
  jand g03405(.dina(n20667), .dinb(n378), .dout(n20668));
  jor  g03406(.dina(n20580), .dinb(n20502), .dout(n20669));
  jxor g03407(.dina(n20527), .dinb(n20526), .dout(n20670));
  jor  g03408(.dina(n20670), .dinb(n20582), .dout(n20671));
  jand g03409(.dina(n20671), .dinb(n20669), .dout(n20672));
  jand g03410(.dina(n20672), .dinb(n377), .dout(n20673));
  jor  g03411(.dina(n20580), .dinb(n20507), .dout(n20674));
  jxor g03412(.dina(n20524), .dinb(n20523), .dout(n20675));
  jor  g03413(.dina(n20675), .dinb(n20582), .dout(n20676));
  jand g03414(.dina(n20676), .dinb(n20674), .dout(n20677));
  jand g03415(.dina(n20677), .dinb(n376), .dout(n20678));
  jor  g03416(.dina(n20580), .dinb(n20512), .dout(n20679));
  jxor g03417(.dina(n20521), .dinb(n20520), .dout(n20680));
  jor  g03418(.dina(n20680), .dinb(n20582), .dout(n20681));
  jand g03419(.dina(n20681), .dinb(n20679), .dout(n20682));
  jand g03420(.dina(n20682), .dinb(n264), .dout(n20683));
  jor  g03421(.dina(n20580), .dinb(n20515), .dout(n20684));
  jxor g03422(.dina(n20518), .dinb(n2505), .dout(n20685));
  jor  g03423(.dina(n20685), .dinb(n20582), .dout(n20686));
  jand g03424(.dina(n20686), .dinb(n20684), .dout(n20687));
  jand g03425(.dina(n20687), .dinb(n386), .dout(n20688));
  jnot g03426(.din(n2681), .dout(n20689));
  jnot g03427(.din(n20419), .dout(n20690));
  jnot g03428(.din(n20423), .dout(n20691));
  jnot g03429(.din(n20428), .dout(n20692));
  jnot g03430(.din(n20433), .dout(n20693));
  jnot g03431(.din(n20438), .dout(n20694));
  jnot g03432(.din(n20443), .dout(n20695));
  jnot g03433(.din(n20448), .dout(n20696));
  jnot g03434(.din(n20453), .dout(n20697));
  jnot g03435(.din(n20458), .dout(n20698));
  jnot g03436(.din(n20463), .dout(n20699));
  jnot g03437(.din(n20468), .dout(n20700));
  jnot g03438(.din(n20473), .dout(n20701));
  jnot g03439(.din(n20478), .dout(n20702));
  jnot g03440(.din(n20483), .dout(n20703));
  jnot g03441(.din(n20488), .dout(n20704));
  jnot g03442(.din(n20493), .dout(n20705));
  jnot g03443(.din(n20498), .dout(n20706));
  jnot g03444(.din(n20503), .dout(n20707));
  jnot g03445(.din(n20508), .dout(n20708));
  jnot g03446(.din(n20513), .dout(n20709));
  jnot g03447(.din(n20516), .dout(n20710));
  jxor g03448(.dina(n20517), .dinb(n259), .dout(n20711));
  jor  g03449(.dina(n20711), .dinb(n2504), .dout(n20712));
  jand g03450(.dina(n20712), .dinb(n20710), .dout(n20713));
  jnot g03451(.din(n20521), .dout(n20714));
  jor  g03452(.dina(n20714), .dinb(n20713), .dout(n20715));
  jand g03453(.dina(n20715), .dinb(n20709), .dout(n20716));
  jnot g03454(.din(n20524), .dout(n20717));
  jor  g03455(.dina(n20717), .dinb(n20716), .dout(n20718));
  jand g03456(.dina(n20718), .dinb(n20708), .dout(n20719));
  jnot g03457(.din(n20527), .dout(n20720));
  jor  g03458(.dina(n20720), .dinb(n20719), .dout(n20721));
  jand g03459(.dina(n20721), .dinb(n20707), .dout(n20722));
  jnot g03460(.din(n20530), .dout(n20723));
  jor  g03461(.dina(n20723), .dinb(n20722), .dout(n20724));
  jand g03462(.dina(n20724), .dinb(n20706), .dout(n20725));
  jnot g03463(.din(n20533), .dout(n20726));
  jor  g03464(.dina(n20726), .dinb(n20725), .dout(n20727));
  jand g03465(.dina(n20727), .dinb(n20705), .dout(n20728));
  jnot g03466(.din(n20536), .dout(n20729));
  jor  g03467(.dina(n20729), .dinb(n20728), .dout(n20730));
  jand g03468(.dina(n20730), .dinb(n20704), .dout(n20731));
  jnot g03469(.din(n20539), .dout(n20732));
  jor  g03470(.dina(n20732), .dinb(n20731), .dout(n20733));
  jand g03471(.dina(n20733), .dinb(n20703), .dout(n20734));
  jnot g03472(.din(n20542), .dout(n20735));
  jor  g03473(.dina(n20735), .dinb(n20734), .dout(n20736));
  jand g03474(.dina(n20736), .dinb(n20702), .dout(n20737));
  jnot g03475(.din(n20545), .dout(n20738));
  jor  g03476(.dina(n20738), .dinb(n20737), .dout(n20739));
  jand g03477(.dina(n20739), .dinb(n20701), .dout(n20740));
  jnot g03478(.din(n20548), .dout(n20741));
  jor  g03479(.dina(n20741), .dinb(n20740), .dout(n20742));
  jand g03480(.dina(n20742), .dinb(n20700), .dout(n20743));
  jnot g03481(.din(n20551), .dout(n20744));
  jor  g03482(.dina(n20744), .dinb(n20743), .dout(n20745));
  jand g03483(.dina(n20745), .dinb(n20699), .dout(n20746));
  jnot g03484(.din(n20554), .dout(n20747));
  jor  g03485(.dina(n20747), .dinb(n20746), .dout(n20748));
  jand g03486(.dina(n20748), .dinb(n20698), .dout(n20749));
  jnot g03487(.din(n20557), .dout(n20750));
  jor  g03488(.dina(n20750), .dinb(n20749), .dout(n20751));
  jand g03489(.dina(n20751), .dinb(n20697), .dout(n20752));
  jnot g03490(.din(n20560), .dout(n20753));
  jor  g03491(.dina(n20753), .dinb(n20752), .dout(n20754));
  jand g03492(.dina(n20754), .dinb(n20696), .dout(n20755));
  jnot g03493(.din(n20563), .dout(n20756));
  jor  g03494(.dina(n20756), .dinb(n20755), .dout(n20757));
  jand g03495(.dina(n20757), .dinb(n20695), .dout(n20758));
  jnot g03496(.din(n20566), .dout(n20759));
  jor  g03497(.dina(n20759), .dinb(n20758), .dout(n20760));
  jand g03498(.dina(n20760), .dinb(n20694), .dout(n20761));
  jnot g03499(.din(n20569), .dout(n20762));
  jor  g03500(.dina(n20762), .dinb(n20761), .dout(n20763));
  jand g03501(.dina(n20763), .dinb(n20693), .dout(n20764));
  jnot g03502(.din(n20572), .dout(n20765));
  jor  g03503(.dina(n20765), .dinb(n20764), .dout(n20766));
  jand g03504(.dina(n20766), .dinb(n20692), .dout(n20767));
  jnot g03505(.din(n20575), .dout(n20768));
  jor  g03506(.dina(n20768), .dinb(n20767), .dout(n20769));
  jand g03507(.dina(n20769), .dinb(n20691), .dout(n20770));
  jor  g03508(.dina(n20770), .dinb(n20421), .dout(n20771));
  jand g03509(.dina(n20771), .dinb(n20690), .dout(n20772));
  jor  g03510(.dina(n20772), .dinb(n20689), .dout(n20773));
  jand g03511(.dina(n20773), .dinb(a42 ), .dout(n20774));
  jnot g03512(.din(n2684), .dout(n20775));
  jor  g03513(.dina(n20772), .dinb(n20775), .dout(n20776));
  jnot g03514(.din(n20776), .dout(n20777));
  jor  g03515(.dina(n20777), .dinb(n20774), .dout(n20778));
  jand g03516(.dina(n20778), .dinb(n259), .dout(n20779));
  jand g03517(.dina(n20579), .dinb(n2681), .dout(n20780));
  jor  g03518(.dina(n20780), .dinb(n2503), .dout(n20781));
  jand g03519(.dina(n20776), .dinb(n20781), .dout(n20782));
  jxor g03520(.dina(n20782), .dinb(b1 ), .dout(n20783));
  jand g03521(.dina(n20783), .dinb(n2691), .dout(n20784));
  jor  g03522(.dina(n20784), .dinb(n20779), .dout(n20785));
  jxor g03523(.dina(n20687), .dinb(n386), .dout(n20786));
  jand g03524(.dina(n20786), .dinb(n20785), .dout(n20787));
  jor  g03525(.dina(n20787), .dinb(n20688), .dout(n20788));
  jxor g03526(.dina(n20682), .dinb(n264), .dout(n20789));
  jand g03527(.dina(n20789), .dinb(n20788), .dout(n20790));
  jor  g03528(.dina(n20790), .dinb(n20683), .dout(n20791));
  jxor g03529(.dina(n20677), .dinb(n376), .dout(n20792));
  jand g03530(.dina(n20792), .dinb(n20791), .dout(n20793));
  jor  g03531(.dina(n20793), .dinb(n20678), .dout(n20794));
  jxor g03532(.dina(n20672), .dinb(n377), .dout(n20795));
  jand g03533(.dina(n20795), .dinb(n20794), .dout(n20796));
  jor  g03534(.dina(n20796), .dinb(n20673), .dout(n20797));
  jxor g03535(.dina(n20667), .dinb(n378), .dout(n20798));
  jand g03536(.dina(n20798), .dinb(n20797), .dout(n20799));
  jor  g03537(.dina(n20799), .dinb(n20668), .dout(n20800));
  jxor g03538(.dina(n20662), .dinb(n265), .dout(n20801));
  jand g03539(.dina(n20801), .dinb(n20800), .dout(n20802));
  jor  g03540(.dina(n20802), .dinb(n20663), .dout(n20803));
  jxor g03541(.dina(n20657), .dinb(n367), .dout(n20804));
  jand g03542(.dina(n20804), .dinb(n20803), .dout(n20805));
  jor  g03543(.dina(n20805), .dinb(n20658), .dout(n20806));
  jxor g03544(.dina(n20652), .dinb(n368), .dout(n20807));
  jand g03545(.dina(n20807), .dinb(n20806), .dout(n20808));
  jor  g03546(.dina(n20808), .dinb(n20653), .dout(n20809));
  jxor g03547(.dina(n20647), .dinb(n369), .dout(n20810));
  jand g03548(.dina(n20810), .dinb(n20809), .dout(n20811));
  jor  g03549(.dina(n20811), .dinb(n20648), .dout(n20812));
  jxor g03550(.dina(n20642), .dinb(n359), .dout(n20813));
  jand g03551(.dina(n20813), .dinb(n20812), .dout(n20814));
  jor  g03552(.dina(n20814), .dinb(n20643), .dout(n20815));
  jxor g03553(.dina(n20637), .dinb(n363), .dout(n20816));
  jand g03554(.dina(n20816), .dinb(n20815), .dout(n20817));
  jor  g03555(.dina(n20817), .dinb(n20638), .dout(n20818));
  jxor g03556(.dina(n20632), .dinb(n360), .dout(n20819));
  jand g03557(.dina(n20819), .dinb(n20818), .dout(n20820));
  jor  g03558(.dina(n20820), .dinb(n20633), .dout(n20821));
  jxor g03559(.dina(n20627), .dinb(n361), .dout(n20822));
  jand g03560(.dina(n20822), .dinb(n20821), .dout(n20823));
  jor  g03561(.dina(n20823), .dinb(n20628), .dout(n20824));
  jxor g03562(.dina(n20622), .dinb(n364), .dout(n20825));
  jand g03563(.dina(n20825), .dinb(n20824), .dout(n20826));
  jor  g03564(.dina(n20826), .dinb(n20623), .dout(n20827));
  jxor g03565(.dina(n20617), .dinb(n355), .dout(n20828));
  jand g03566(.dina(n20828), .dinb(n20827), .dout(n20829));
  jor  g03567(.dina(n20829), .dinb(n20618), .dout(n20830));
  jxor g03568(.dina(n20612), .dinb(n356), .dout(n20831));
  jand g03569(.dina(n20831), .dinb(n20830), .dout(n20832));
  jor  g03570(.dina(n20832), .dinb(n20613), .dout(n20833));
  jxor g03571(.dina(n20607), .dinb(n266), .dout(n20834));
  jand g03572(.dina(n20834), .dinb(n20833), .dout(n20835));
  jor  g03573(.dina(n20835), .dinb(n20608), .dout(n20836));
  jxor g03574(.dina(n20602), .dinb(n267), .dout(n20837));
  jand g03575(.dina(n20837), .dinb(n20836), .dout(n20838));
  jor  g03576(.dina(n20838), .dinb(n20603), .dout(n20839));
  jxor g03577(.dina(n20597), .dinb(n347), .dout(n20840));
  jand g03578(.dina(n20840), .dinb(n20839), .dout(n20841));
  jor  g03579(.dina(n20841), .dinb(n20598), .dout(n20842));
  jxor g03580(.dina(n20585), .dinb(n348), .dout(n20843));
  jand g03581(.dina(n20843), .dinb(n20842), .dout(n20844));
  jor  g03582(.dina(n20844), .dinb(n20593), .dout(n20845));
  jand g03583(.dina(n20845), .dinb(n20592), .dout(n20846));
  jor  g03584(.dina(n20846), .dinb(n20589), .dout(n20847));
  jand g03585(.dina(n20847), .dinb(n417), .dout(n20848));
  jor  g03586(.dina(n20848), .dinb(n20585), .dout(n20849));
  jnot g03587(.din(n20589), .dout(n20850));
  jnot g03588(.din(n20593), .dout(n20851));
  jnot g03589(.din(n20598), .dout(n20852));
  jnot g03590(.din(n20603), .dout(n20853));
  jnot g03591(.din(n20608), .dout(n20854));
  jnot g03592(.din(n20613), .dout(n20855));
  jnot g03593(.din(n20618), .dout(n20856));
  jnot g03594(.din(n20623), .dout(n20857));
  jnot g03595(.din(n20628), .dout(n20858));
  jnot g03596(.din(n20633), .dout(n20859));
  jnot g03597(.din(n20638), .dout(n20860));
  jnot g03598(.din(n20643), .dout(n20861));
  jnot g03599(.din(n20648), .dout(n20862));
  jnot g03600(.din(n20653), .dout(n20863));
  jnot g03601(.din(n20658), .dout(n20864));
  jnot g03602(.din(n20663), .dout(n20865));
  jnot g03603(.din(n20668), .dout(n20866));
  jnot g03604(.din(n20673), .dout(n20867));
  jnot g03605(.din(n20678), .dout(n20868));
  jnot g03606(.din(n20683), .dout(n20869));
  jnot g03607(.din(n20688), .dout(n20870));
  jor  g03608(.dina(n20782), .dinb(b1 ), .dout(n20871));
  jxor g03609(.dina(n20782), .dinb(n259), .dout(n20872));
  jor  g03610(.dina(n20872), .dinb(n2690), .dout(n20873));
  jand g03611(.dina(n20873), .dinb(n20871), .dout(n20874));
  jxor g03612(.dina(n20687), .dinb(b2 ), .dout(n20875));
  jor  g03613(.dina(n20875), .dinb(n20874), .dout(n20876));
  jand g03614(.dina(n20876), .dinb(n20870), .dout(n20877));
  jnot g03615(.din(n20789), .dout(n20878));
  jor  g03616(.dina(n20878), .dinb(n20877), .dout(n20879));
  jand g03617(.dina(n20879), .dinb(n20869), .dout(n20880));
  jnot g03618(.din(n20792), .dout(n20881));
  jor  g03619(.dina(n20881), .dinb(n20880), .dout(n20882));
  jand g03620(.dina(n20882), .dinb(n20868), .dout(n20883));
  jnot g03621(.din(n20795), .dout(n20884));
  jor  g03622(.dina(n20884), .dinb(n20883), .dout(n20885));
  jand g03623(.dina(n20885), .dinb(n20867), .dout(n20886));
  jnot g03624(.din(n20798), .dout(n20887));
  jor  g03625(.dina(n20887), .dinb(n20886), .dout(n20888));
  jand g03626(.dina(n20888), .dinb(n20866), .dout(n20889));
  jnot g03627(.din(n20801), .dout(n20890));
  jor  g03628(.dina(n20890), .dinb(n20889), .dout(n20891));
  jand g03629(.dina(n20891), .dinb(n20865), .dout(n20892));
  jnot g03630(.din(n20804), .dout(n20893));
  jor  g03631(.dina(n20893), .dinb(n20892), .dout(n20894));
  jand g03632(.dina(n20894), .dinb(n20864), .dout(n20895));
  jnot g03633(.din(n20807), .dout(n20896));
  jor  g03634(.dina(n20896), .dinb(n20895), .dout(n20897));
  jand g03635(.dina(n20897), .dinb(n20863), .dout(n20898));
  jnot g03636(.din(n20810), .dout(n20899));
  jor  g03637(.dina(n20899), .dinb(n20898), .dout(n20900));
  jand g03638(.dina(n20900), .dinb(n20862), .dout(n20901));
  jnot g03639(.din(n20813), .dout(n20902));
  jor  g03640(.dina(n20902), .dinb(n20901), .dout(n20903));
  jand g03641(.dina(n20903), .dinb(n20861), .dout(n20904));
  jnot g03642(.din(n20816), .dout(n20905));
  jor  g03643(.dina(n20905), .dinb(n20904), .dout(n20906));
  jand g03644(.dina(n20906), .dinb(n20860), .dout(n20907));
  jnot g03645(.din(n20819), .dout(n20908));
  jor  g03646(.dina(n20908), .dinb(n20907), .dout(n20909));
  jand g03647(.dina(n20909), .dinb(n20859), .dout(n20910));
  jnot g03648(.din(n20822), .dout(n20911));
  jor  g03649(.dina(n20911), .dinb(n20910), .dout(n20912));
  jand g03650(.dina(n20912), .dinb(n20858), .dout(n20913));
  jnot g03651(.din(n20825), .dout(n20914));
  jor  g03652(.dina(n20914), .dinb(n20913), .dout(n20915));
  jand g03653(.dina(n20915), .dinb(n20857), .dout(n20916));
  jnot g03654(.din(n20828), .dout(n20917));
  jor  g03655(.dina(n20917), .dinb(n20916), .dout(n20918));
  jand g03656(.dina(n20918), .dinb(n20856), .dout(n20919));
  jnot g03657(.din(n20831), .dout(n20920));
  jor  g03658(.dina(n20920), .dinb(n20919), .dout(n20921));
  jand g03659(.dina(n20921), .dinb(n20855), .dout(n20922));
  jnot g03660(.din(n20834), .dout(n20923));
  jor  g03661(.dina(n20923), .dinb(n20922), .dout(n20924));
  jand g03662(.dina(n20924), .dinb(n20854), .dout(n20925));
  jnot g03663(.din(n20837), .dout(n20926));
  jor  g03664(.dina(n20926), .dinb(n20925), .dout(n20927));
  jand g03665(.dina(n20927), .dinb(n20853), .dout(n20928));
  jnot g03666(.din(n20840), .dout(n20929));
  jor  g03667(.dina(n20929), .dinb(n20928), .dout(n20930));
  jand g03668(.dina(n20930), .dinb(n20852), .dout(n20931));
  jnot g03669(.din(n20843), .dout(n20932));
  jor  g03670(.dina(n20932), .dinb(n20931), .dout(n20933));
  jand g03671(.dina(n20933), .dinb(n20851), .dout(n20934));
  jor  g03672(.dina(n20934), .dinb(n20591), .dout(n20935));
  jand g03673(.dina(n20935), .dinb(n20850), .dout(n20936));
  jor  g03674(.dina(n20936), .dinb(n861), .dout(n20937));
  jxor g03675(.dina(n20843), .dinb(n20842), .dout(n20938));
  jor  g03676(.dina(n20938), .dinb(n20937), .dout(n20939));
  jand g03677(.dina(n20939), .dinb(n20849), .dout(n20940));
  jand g03678(.dina(n20937), .dinb(n20588), .dout(n20941));
  jand g03679(.dina(n20845), .dinb(n20589), .dout(n20942));
  jor  g03680(.dina(n20942), .dinb(n20941), .dout(n20943));
  jand g03681(.dina(n20943), .dinb(n268), .dout(n20944));
  jand g03682(.dina(n20944), .dinb(n416), .dout(n20945));
  jand g03683(.dina(n20940), .dinb(n349), .dout(n20946));
  jor  g03684(.dina(n20848), .dinb(n20597), .dout(n20947));
  jxor g03685(.dina(n20840), .dinb(n20839), .dout(n20948));
  jor  g03686(.dina(n20948), .dinb(n20937), .dout(n20949));
  jand g03687(.dina(n20949), .dinb(n20947), .dout(n20950));
  jand g03688(.dina(n20950), .dinb(n348), .dout(n20951));
  jor  g03689(.dina(n20848), .dinb(n20602), .dout(n20952));
  jxor g03690(.dina(n20837), .dinb(n20836), .dout(n20953));
  jor  g03691(.dina(n20953), .dinb(n20937), .dout(n20954));
  jand g03692(.dina(n20954), .dinb(n20952), .dout(n20955));
  jand g03693(.dina(n20955), .dinb(n347), .dout(n20956));
  jor  g03694(.dina(n20848), .dinb(n20607), .dout(n20957));
  jxor g03695(.dina(n20834), .dinb(n20833), .dout(n20958));
  jor  g03696(.dina(n20958), .dinb(n20937), .dout(n20959));
  jand g03697(.dina(n20959), .dinb(n20957), .dout(n20960));
  jand g03698(.dina(n20960), .dinb(n267), .dout(n20961));
  jor  g03699(.dina(n20848), .dinb(n20612), .dout(n20962));
  jxor g03700(.dina(n20831), .dinb(n20830), .dout(n20963));
  jor  g03701(.dina(n20963), .dinb(n20937), .dout(n20964));
  jand g03702(.dina(n20964), .dinb(n20962), .dout(n20965));
  jand g03703(.dina(n20965), .dinb(n266), .dout(n20966));
  jor  g03704(.dina(n20848), .dinb(n20617), .dout(n20967));
  jxor g03705(.dina(n20828), .dinb(n20827), .dout(n20968));
  jor  g03706(.dina(n20968), .dinb(n20937), .dout(n20969));
  jand g03707(.dina(n20969), .dinb(n20967), .dout(n20970));
  jand g03708(.dina(n20970), .dinb(n356), .dout(n20971));
  jor  g03709(.dina(n20848), .dinb(n20622), .dout(n20972));
  jxor g03710(.dina(n20825), .dinb(n20824), .dout(n20973));
  jor  g03711(.dina(n20973), .dinb(n20937), .dout(n20974));
  jand g03712(.dina(n20974), .dinb(n20972), .dout(n20975));
  jand g03713(.dina(n20975), .dinb(n355), .dout(n20976));
  jor  g03714(.dina(n20848), .dinb(n20627), .dout(n20977));
  jxor g03715(.dina(n20822), .dinb(n20821), .dout(n20978));
  jor  g03716(.dina(n20978), .dinb(n20937), .dout(n20979));
  jand g03717(.dina(n20979), .dinb(n20977), .dout(n20980));
  jand g03718(.dina(n20980), .dinb(n364), .dout(n20981));
  jor  g03719(.dina(n20848), .dinb(n20632), .dout(n20982));
  jxor g03720(.dina(n20819), .dinb(n20818), .dout(n20983));
  jor  g03721(.dina(n20983), .dinb(n20937), .dout(n20984));
  jand g03722(.dina(n20984), .dinb(n20982), .dout(n20985));
  jand g03723(.dina(n20985), .dinb(n361), .dout(n20986));
  jor  g03724(.dina(n20848), .dinb(n20637), .dout(n20987));
  jxor g03725(.dina(n20816), .dinb(n20815), .dout(n20988));
  jor  g03726(.dina(n20988), .dinb(n20937), .dout(n20989));
  jand g03727(.dina(n20989), .dinb(n20987), .dout(n20990));
  jand g03728(.dina(n20990), .dinb(n360), .dout(n20991));
  jor  g03729(.dina(n20848), .dinb(n20642), .dout(n20992));
  jxor g03730(.dina(n20813), .dinb(n20812), .dout(n20993));
  jor  g03731(.dina(n20993), .dinb(n20937), .dout(n20994));
  jand g03732(.dina(n20994), .dinb(n20992), .dout(n20995));
  jand g03733(.dina(n20995), .dinb(n363), .dout(n20996));
  jor  g03734(.dina(n20848), .dinb(n20647), .dout(n20997));
  jxor g03735(.dina(n20810), .dinb(n20809), .dout(n20998));
  jor  g03736(.dina(n20998), .dinb(n20937), .dout(n20999));
  jand g03737(.dina(n20999), .dinb(n20997), .dout(n21000));
  jand g03738(.dina(n21000), .dinb(n359), .dout(n21001));
  jor  g03739(.dina(n20848), .dinb(n20652), .dout(n21002));
  jxor g03740(.dina(n20807), .dinb(n20806), .dout(n21003));
  jor  g03741(.dina(n21003), .dinb(n20937), .dout(n21004));
  jand g03742(.dina(n21004), .dinb(n21002), .dout(n21005));
  jand g03743(.dina(n21005), .dinb(n369), .dout(n21006));
  jor  g03744(.dina(n20848), .dinb(n20657), .dout(n21007));
  jxor g03745(.dina(n20804), .dinb(n20803), .dout(n21008));
  jor  g03746(.dina(n21008), .dinb(n20937), .dout(n21009));
  jand g03747(.dina(n21009), .dinb(n21007), .dout(n21010));
  jand g03748(.dina(n21010), .dinb(n368), .dout(n21011));
  jor  g03749(.dina(n20848), .dinb(n20662), .dout(n21012));
  jxor g03750(.dina(n20801), .dinb(n20800), .dout(n21013));
  jor  g03751(.dina(n21013), .dinb(n20937), .dout(n21014));
  jand g03752(.dina(n21014), .dinb(n21012), .dout(n21015));
  jand g03753(.dina(n21015), .dinb(n367), .dout(n21016));
  jor  g03754(.dina(n20848), .dinb(n20667), .dout(n21017));
  jxor g03755(.dina(n20798), .dinb(n20797), .dout(n21018));
  jor  g03756(.dina(n21018), .dinb(n20937), .dout(n21019));
  jand g03757(.dina(n21019), .dinb(n21017), .dout(n21020));
  jand g03758(.dina(n21020), .dinb(n265), .dout(n21021));
  jor  g03759(.dina(n20848), .dinb(n20672), .dout(n21022));
  jxor g03760(.dina(n20795), .dinb(n20794), .dout(n21023));
  jor  g03761(.dina(n21023), .dinb(n20937), .dout(n21024));
  jand g03762(.dina(n21024), .dinb(n21022), .dout(n21025));
  jand g03763(.dina(n21025), .dinb(n378), .dout(n21026));
  jor  g03764(.dina(n20848), .dinb(n20677), .dout(n21027));
  jxor g03765(.dina(n20792), .dinb(n20791), .dout(n21028));
  jor  g03766(.dina(n21028), .dinb(n20937), .dout(n21029));
  jand g03767(.dina(n21029), .dinb(n21027), .dout(n21030));
  jand g03768(.dina(n21030), .dinb(n377), .dout(n21031));
  jor  g03769(.dina(n20848), .dinb(n20682), .dout(n21032));
  jxor g03770(.dina(n20789), .dinb(n20788), .dout(n21033));
  jor  g03771(.dina(n21033), .dinb(n20937), .dout(n21034));
  jand g03772(.dina(n21034), .dinb(n21032), .dout(n21035));
  jand g03773(.dina(n21035), .dinb(n376), .dout(n21036));
  jor  g03774(.dina(n20848), .dinb(n20687), .dout(n21037));
  jxor g03775(.dina(n20786), .dinb(n20785), .dout(n21038));
  jor  g03776(.dina(n21038), .dinb(n20937), .dout(n21039));
  jand g03777(.dina(n21039), .dinb(n21037), .dout(n21040));
  jand g03778(.dina(n21040), .dinb(n264), .dout(n21041));
  jand g03779(.dina(n20937), .dinb(n20778), .dout(n21042));
  jxor g03780(.dina(n20783), .dinb(n2691), .dout(n21043));
  jand g03781(.dina(n21043), .dinb(n20848), .dout(n21044));
  jor  g03782(.dina(n21044), .dinb(n21042), .dout(n21045));
  jand g03783(.dina(n21045), .dinb(n386), .dout(n21046));
  jnot g03784(.din(n2873), .dout(n21047));
  jor  g03785(.dina(n20936), .dinb(n21047), .dout(n21048));
  jand g03786(.dina(n21048), .dinb(a41 ), .dout(n21049));
  jand g03787(.dina(n20848), .dinb(n2690), .dout(n21050));
  jor  g03788(.dina(n21050), .dinb(n21049), .dout(n21051));
  jand g03789(.dina(n21051), .dinb(n259), .dout(n21052));
  jand g03790(.dina(n20847), .dinb(n2873), .dout(n21053));
  jor  g03791(.dina(n21053), .dinb(n2689), .dout(n21054));
  jor  g03792(.dina(n20937), .dinb(n2691), .dout(n21055));
  jand g03793(.dina(n21055), .dinb(n21054), .dout(n21056));
  jxor g03794(.dina(n21056), .dinb(b1 ), .dout(n21057));
  jand g03795(.dina(n21057), .dinb(n2882), .dout(n21058));
  jor  g03796(.dina(n21058), .dinb(n21052), .dout(n21059));
  jxor g03797(.dina(n21045), .dinb(n386), .dout(n21060));
  jand g03798(.dina(n21060), .dinb(n21059), .dout(n21061));
  jor  g03799(.dina(n21061), .dinb(n21046), .dout(n21062));
  jxor g03800(.dina(n21040), .dinb(n264), .dout(n21063));
  jand g03801(.dina(n21063), .dinb(n21062), .dout(n21064));
  jor  g03802(.dina(n21064), .dinb(n21041), .dout(n21065));
  jxor g03803(.dina(n21035), .dinb(n376), .dout(n21066));
  jand g03804(.dina(n21066), .dinb(n21065), .dout(n21067));
  jor  g03805(.dina(n21067), .dinb(n21036), .dout(n21068));
  jxor g03806(.dina(n21030), .dinb(n377), .dout(n21069));
  jand g03807(.dina(n21069), .dinb(n21068), .dout(n21070));
  jor  g03808(.dina(n21070), .dinb(n21031), .dout(n21071));
  jxor g03809(.dina(n21025), .dinb(n378), .dout(n21072));
  jand g03810(.dina(n21072), .dinb(n21071), .dout(n21073));
  jor  g03811(.dina(n21073), .dinb(n21026), .dout(n21074));
  jxor g03812(.dina(n21020), .dinb(n265), .dout(n21075));
  jand g03813(.dina(n21075), .dinb(n21074), .dout(n21076));
  jor  g03814(.dina(n21076), .dinb(n21021), .dout(n21077));
  jxor g03815(.dina(n21015), .dinb(n367), .dout(n21078));
  jand g03816(.dina(n21078), .dinb(n21077), .dout(n21079));
  jor  g03817(.dina(n21079), .dinb(n21016), .dout(n21080));
  jxor g03818(.dina(n21010), .dinb(n368), .dout(n21081));
  jand g03819(.dina(n21081), .dinb(n21080), .dout(n21082));
  jor  g03820(.dina(n21082), .dinb(n21011), .dout(n21083));
  jxor g03821(.dina(n21005), .dinb(n369), .dout(n21084));
  jand g03822(.dina(n21084), .dinb(n21083), .dout(n21085));
  jor  g03823(.dina(n21085), .dinb(n21006), .dout(n21086));
  jxor g03824(.dina(n21000), .dinb(n359), .dout(n21087));
  jand g03825(.dina(n21087), .dinb(n21086), .dout(n21088));
  jor  g03826(.dina(n21088), .dinb(n21001), .dout(n21089));
  jxor g03827(.dina(n20995), .dinb(n363), .dout(n21090));
  jand g03828(.dina(n21090), .dinb(n21089), .dout(n21091));
  jor  g03829(.dina(n21091), .dinb(n20996), .dout(n21092));
  jxor g03830(.dina(n20990), .dinb(n360), .dout(n21093));
  jand g03831(.dina(n21093), .dinb(n21092), .dout(n21094));
  jor  g03832(.dina(n21094), .dinb(n20991), .dout(n21095));
  jxor g03833(.dina(n20985), .dinb(n361), .dout(n21096));
  jand g03834(.dina(n21096), .dinb(n21095), .dout(n21097));
  jor  g03835(.dina(n21097), .dinb(n20986), .dout(n21098));
  jxor g03836(.dina(n20980), .dinb(n364), .dout(n21099));
  jand g03837(.dina(n21099), .dinb(n21098), .dout(n21100));
  jor  g03838(.dina(n21100), .dinb(n20981), .dout(n21101));
  jxor g03839(.dina(n20975), .dinb(n355), .dout(n21102));
  jand g03840(.dina(n21102), .dinb(n21101), .dout(n21103));
  jor  g03841(.dina(n21103), .dinb(n20976), .dout(n21104));
  jxor g03842(.dina(n20970), .dinb(n356), .dout(n21105));
  jand g03843(.dina(n21105), .dinb(n21104), .dout(n21106));
  jor  g03844(.dina(n21106), .dinb(n20971), .dout(n21107));
  jxor g03845(.dina(n20965), .dinb(n266), .dout(n21108));
  jand g03846(.dina(n21108), .dinb(n21107), .dout(n21109));
  jor  g03847(.dina(n21109), .dinb(n20966), .dout(n21110));
  jxor g03848(.dina(n20960), .dinb(n267), .dout(n21111));
  jand g03849(.dina(n21111), .dinb(n21110), .dout(n21112));
  jor  g03850(.dina(n21112), .dinb(n20961), .dout(n21113));
  jxor g03851(.dina(n20955), .dinb(n347), .dout(n21114));
  jand g03852(.dina(n21114), .dinb(n21113), .dout(n21115));
  jor  g03853(.dina(n21115), .dinb(n20956), .dout(n21116));
  jxor g03854(.dina(n20950), .dinb(n348), .dout(n21117));
  jand g03855(.dina(n21117), .dinb(n21116), .dout(n21118));
  jor  g03856(.dina(n21118), .dinb(n20951), .dout(n21119));
  jxor g03857(.dina(n20940), .dinb(n349), .dout(n21120));
  jand g03858(.dina(n21120), .dinb(n21119), .dout(n21121));
  jor  g03859(.dina(n21121), .dinb(n20946), .dout(n21122));
  jxor g03860(.dina(n20943), .dinb(n268), .dout(n21123));
  jand g03861(.dina(n21123), .dinb(n416), .dout(n21124));
  jand g03862(.dina(n21124), .dinb(n21122), .dout(n21125));
  jor  g03863(.dina(n21125), .dinb(n20945), .dout(n21126));
  jor  g03864(.dina(n21126), .dinb(n20940), .dout(n21127));
  jnot g03865(.din(n21126), .dout(n21128));
  jxor g03866(.dina(n21120), .dinb(n21119), .dout(n21129));
  jor  g03867(.dina(n21129), .dinb(n21128), .dout(n21130));
  jand g03868(.dina(n21130), .dinb(n21127), .dout(n21131));
  jand g03869(.dina(n21128), .dinb(n20943), .dout(n21132));
  jxor g03870(.dina(n21123), .dinb(n21122), .dout(n21133));
  jand g03871(.dina(n21133), .dinb(n20945), .dout(n21134));
  jor  g03872(.dina(n21134), .dinb(n21132), .dout(n21135));
  jand g03873(.dina(n21135), .dinb(n274), .dout(n21136));
  jnot g03874(.din(n21135), .dout(n21137));
  jand g03875(.dina(n21137), .dinb(b24 ), .dout(n21138));
  jnot g03876(.din(n21138), .dout(n21139));
  jand g03877(.dina(n21131), .dinb(n268), .dout(n21140));
  jor  g03878(.dina(n21126), .dinb(n20950), .dout(n21141));
  jxor g03879(.dina(n21117), .dinb(n21116), .dout(n21142));
  jor  g03880(.dina(n21142), .dinb(n21128), .dout(n21143));
  jand g03881(.dina(n21143), .dinb(n21141), .dout(n21144));
  jand g03882(.dina(n21144), .dinb(n349), .dout(n21145));
  jor  g03883(.dina(n21126), .dinb(n20955), .dout(n21146));
  jxor g03884(.dina(n21114), .dinb(n21113), .dout(n21147));
  jor  g03885(.dina(n21147), .dinb(n21128), .dout(n21148));
  jand g03886(.dina(n21148), .dinb(n21146), .dout(n21149));
  jand g03887(.dina(n21149), .dinb(n348), .dout(n21150));
  jor  g03888(.dina(n21126), .dinb(n20960), .dout(n21151));
  jxor g03889(.dina(n21111), .dinb(n21110), .dout(n21152));
  jor  g03890(.dina(n21152), .dinb(n21128), .dout(n21153));
  jand g03891(.dina(n21153), .dinb(n21151), .dout(n21154));
  jand g03892(.dina(n21154), .dinb(n347), .dout(n21155));
  jor  g03893(.dina(n21126), .dinb(n20965), .dout(n21156));
  jxor g03894(.dina(n21108), .dinb(n21107), .dout(n21157));
  jor  g03895(.dina(n21157), .dinb(n21128), .dout(n21158));
  jand g03896(.dina(n21158), .dinb(n21156), .dout(n21159));
  jand g03897(.dina(n21159), .dinb(n267), .dout(n21160));
  jor  g03898(.dina(n21126), .dinb(n20970), .dout(n21161));
  jxor g03899(.dina(n21105), .dinb(n21104), .dout(n21162));
  jor  g03900(.dina(n21162), .dinb(n21128), .dout(n21163));
  jand g03901(.dina(n21163), .dinb(n21161), .dout(n21164));
  jand g03902(.dina(n21164), .dinb(n266), .dout(n21165));
  jor  g03903(.dina(n21126), .dinb(n20975), .dout(n21166));
  jxor g03904(.dina(n21102), .dinb(n21101), .dout(n21167));
  jor  g03905(.dina(n21167), .dinb(n21128), .dout(n21168));
  jand g03906(.dina(n21168), .dinb(n21166), .dout(n21169));
  jand g03907(.dina(n21169), .dinb(n356), .dout(n21170));
  jor  g03908(.dina(n21126), .dinb(n20980), .dout(n21171));
  jxor g03909(.dina(n21099), .dinb(n21098), .dout(n21172));
  jor  g03910(.dina(n21172), .dinb(n21128), .dout(n21173));
  jand g03911(.dina(n21173), .dinb(n21171), .dout(n21174));
  jand g03912(.dina(n21174), .dinb(n355), .dout(n21175));
  jor  g03913(.dina(n21126), .dinb(n20985), .dout(n21176));
  jxor g03914(.dina(n21096), .dinb(n21095), .dout(n21177));
  jor  g03915(.dina(n21177), .dinb(n21128), .dout(n21178));
  jand g03916(.dina(n21178), .dinb(n21176), .dout(n21179));
  jand g03917(.dina(n21179), .dinb(n364), .dout(n21180));
  jor  g03918(.dina(n21126), .dinb(n20990), .dout(n21181));
  jxor g03919(.dina(n21093), .dinb(n21092), .dout(n21182));
  jor  g03920(.dina(n21182), .dinb(n21128), .dout(n21183));
  jand g03921(.dina(n21183), .dinb(n21181), .dout(n21184));
  jand g03922(.dina(n21184), .dinb(n361), .dout(n21185));
  jor  g03923(.dina(n21126), .dinb(n20995), .dout(n21186));
  jxor g03924(.dina(n21090), .dinb(n21089), .dout(n21187));
  jor  g03925(.dina(n21187), .dinb(n21128), .dout(n21188));
  jand g03926(.dina(n21188), .dinb(n21186), .dout(n21189));
  jand g03927(.dina(n21189), .dinb(n360), .dout(n21190));
  jor  g03928(.dina(n21126), .dinb(n21000), .dout(n21191));
  jxor g03929(.dina(n21087), .dinb(n21086), .dout(n21192));
  jor  g03930(.dina(n21192), .dinb(n21128), .dout(n21193));
  jand g03931(.dina(n21193), .dinb(n21191), .dout(n21194));
  jand g03932(.dina(n21194), .dinb(n363), .dout(n21195));
  jor  g03933(.dina(n21126), .dinb(n21005), .dout(n21196));
  jxor g03934(.dina(n21084), .dinb(n21083), .dout(n21197));
  jor  g03935(.dina(n21197), .dinb(n21128), .dout(n21198));
  jand g03936(.dina(n21198), .dinb(n21196), .dout(n21199));
  jand g03937(.dina(n21199), .dinb(n359), .dout(n21200));
  jor  g03938(.dina(n21126), .dinb(n21010), .dout(n21201));
  jxor g03939(.dina(n21081), .dinb(n21080), .dout(n21202));
  jor  g03940(.dina(n21202), .dinb(n21128), .dout(n21203));
  jand g03941(.dina(n21203), .dinb(n21201), .dout(n21204));
  jand g03942(.dina(n21204), .dinb(n369), .dout(n21205));
  jor  g03943(.dina(n21126), .dinb(n21015), .dout(n21206));
  jxor g03944(.dina(n21078), .dinb(n21077), .dout(n21207));
  jor  g03945(.dina(n21207), .dinb(n21128), .dout(n21208));
  jand g03946(.dina(n21208), .dinb(n21206), .dout(n21209));
  jand g03947(.dina(n21209), .dinb(n368), .dout(n21210));
  jor  g03948(.dina(n21126), .dinb(n21020), .dout(n21211));
  jxor g03949(.dina(n21075), .dinb(n21074), .dout(n21212));
  jor  g03950(.dina(n21212), .dinb(n21128), .dout(n21213));
  jand g03951(.dina(n21213), .dinb(n21211), .dout(n21214));
  jand g03952(.dina(n21214), .dinb(n367), .dout(n21215));
  jor  g03953(.dina(n21126), .dinb(n21025), .dout(n21216));
  jxor g03954(.dina(n21072), .dinb(n21071), .dout(n21217));
  jor  g03955(.dina(n21217), .dinb(n21128), .dout(n21218));
  jand g03956(.dina(n21218), .dinb(n21216), .dout(n21219));
  jand g03957(.dina(n21219), .dinb(n265), .dout(n21220));
  jor  g03958(.dina(n21126), .dinb(n21030), .dout(n21221));
  jxor g03959(.dina(n21069), .dinb(n21068), .dout(n21222));
  jor  g03960(.dina(n21222), .dinb(n21128), .dout(n21223));
  jand g03961(.dina(n21223), .dinb(n21221), .dout(n21224));
  jand g03962(.dina(n21224), .dinb(n378), .dout(n21225));
  jor  g03963(.dina(n21126), .dinb(n21035), .dout(n21226));
  jxor g03964(.dina(n21066), .dinb(n21065), .dout(n21227));
  jor  g03965(.dina(n21227), .dinb(n21128), .dout(n21228));
  jand g03966(.dina(n21228), .dinb(n21226), .dout(n21229));
  jand g03967(.dina(n21229), .dinb(n377), .dout(n21230));
  jor  g03968(.dina(n21126), .dinb(n21040), .dout(n21231));
  jxor g03969(.dina(n21063), .dinb(n21062), .dout(n21232));
  jor  g03970(.dina(n21232), .dinb(n21128), .dout(n21233));
  jand g03971(.dina(n21233), .dinb(n21231), .dout(n21234));
  jand g03972(.dina(n21234), .dinb(n376), .dout(n21235));
  jxor g03973(.dina(n21060), .dinb(n21059), .dout(n21236));
  jnot g03974(.din(n21236), .dout(n21237));
  jor  g03975(.dina(n21237), .dinb(n21128), .dout(n21238));
  jnot g03976(.din(n21045), .dout(n21239));
  jor  g03977(.dina(n21126), .dinb(n21239), .dout(n21240));
  jand g03978(.dina(n21240), .dinb(n21238), .dout(n21241));
  jnot g03979(.din(n21241), .dout(n21242));
  jand g03980(.dina(n21242), .dinb(n264), .dout(n21243));
  jor  g03981(.dina(n21126), .dinb(n21051), .dout(n21244));
  jxor g03982(.dina(n21057), .dinb(n2882), .dout(n21245));
  jor  g03983(.dina(n21245), .dinb(n21128), .dout(n21246));
  jand g03984(.dina(n21246), .dinb(n21244), .dout(n21247));
  jand g03985(.dina(n21247), .dinb(n386), .dout(n21248));
  jand g03986(.dina(n21126), .dinb(b0 ), .dout(n21249));
  jxor g03987(.dina(n21249), .dinb(a40 ), .dout(n21250));
  jand g03988(.dina(n21250), .dinb(n259), .dout(n21251));
  jxor g03989(.dina(n21249), .dinb(n2880), .dout(n21252));
  jxor g03990(.dina(n21252), .dinb(b1 ), .dout(n21253));
  jand g03991(.dina(n21253), .dinb(n3078), .dout(n21254));
  jor  g03992(.dina(n21254), .dinb(n21251), .dout(n21255));
  jxor g03993(.dina(n21247), .dinb(n386), .dout(n21256));
  jand g03994(.dina(n21256), .dinb(n21255), .dout(n21257));
  jor  g03995(.dina(n21257), .dinb(n21248), .dout(n21258));
  jxor g03996(.dina(n21241), .dinb(b3 ), .dout(n21259));
  jand g03997(.dina(n21259), .dinb(n21258), .dout(n21260));
  jor  g03998(.dina(n21260), .dinb(n21243), .dout(n21261));
  jxor g03999(.dina(n21234), .dinb(n376), .dout(n21262));
  jand g04000(.dina(n21262), .dinb(n21261), .dout(n21263));
  jor  g04001(.dina(n21263), .dinb(n21235), .dout(n21264));
  jxor g04002(.dina(n21229), .dinb(n377), .dout(n21265));
  jand g04003(.dina(n21265), .dinb(n21264), .dout(n21266));
  jor  g04004(.dina(n21266), .dinb(n21230), .dout(n21267));
  jxor g04005(.dina(n21224), .dinb(n378), .dout(n21268));
  jand g04006(.dina(n21268), .dinb(n21267), .dout(n21269));
  jor  g04007(.dina(n21269), .dinb(n21225), .dout(n21270));
  jxor g04008(.dina(n21219), .dinb(n265), .dout(n21271));
  jand g04009(.dina(n21271), .dinb(n21270), .dout(n21272));
  jor  g04010(.dina(n21272), .dinb(n21220), .dout(n21273));
  jxor g04011(.dina(n21214), .dinb(n367), .dout(n21274));
  jand g04012(.dina(n21274), .dinb(n21273), .dout(n21275));
  jor  g04013(.dina(n21275), .dinb(n21215), .dout(n21276));
  jxor g04014(.dina(n21209), .dinb(n368), .dout(n21277));
  jand g04015(.dina(n21277), .dinb(n21276), .dout(n21278));
  jor  g04016(.dina(n21278), .dinb(n21210), .dout(n21279));
  jxor g04017(.dina(n21204), .dinb(n369), .dout(n21280));
  jand g04018(.dina(n21280), .dinb(n21279), .dout(n21281));
  jor  g04019(.dina(n21281), .dinb(n21205), .dout(n21282));
  jxor g04020(.dina(n21199), .dinb(n359), .dout(n21283));
  jand g04021(.dina(n21283), .dinb(n21282), .dout(n21284));
  jor  g04022(.dina(n21284), .dinb(n21200), .dout(n21285));
  jxor g04023(.dina(n21194), .dinb(n363), .dout(n21286));
  jand g04024(.dina(n21286), .dinb(n21285), .dout(n21287));
  jor  g04025(.dina(n21287), .dinb(n21195), .dout(n21288));
  jxor g04026(.dina(n21189), .dinb(n360), .dout(n21289));
  jand g04027(.dina(n21289), .dinb(n21288), .dout(n21290));
  jor  g04028(.dina(n21290), .dinb(n21190), .dout(n21291));
  jxor g04029(.dina(n21184), .dinb(n361), .dout(n21292));
  jand g04030(.dina(n21292), .dinb(n21291), .dout(n21293));
  jor  g04031(.dina(n21293), .dinb(n21185), .dout(n21294));
  jxor g04032(.dina(n21179), .dinb(n364), .dout(n21295));
  jand g04033(.dina(n21295), .dinb(n21294), .dout(n21296));
  jor  g04034(.dina(n21296), .dinb(n21180), .dout(n21297));
  jxor g04035(.dina(n21174), .dinb(n355), .dout(n21298));
  jand g04036(.dina(n21298), .dinb(n21297), .dout(n21299));
  jor  g04037(.dina(n21299), .dinb(n21175), .dout(n21300));
  jxor g04038(.dina(n21169), .dinb(n356), .dout(n21301));
  jand g04039(.dina(n21301), .dinb(n21300), .dout(n21302));
  jor  g04040(.dina(n21302), .dinb(n21170), .dout(n21303));
  jxor g04041(.dina(n21164), .dinb(n266), .dout(n21304));
  jand g04042(.dina(n21304), .dinb(n21303), .dout(n21305));
  jor  g04043(.dina(n21305), .dinb(n21165), .dout(n21306));
  jxor g04044(.dina(n21159), .dinb(n267), .dout(n21307));
  jand g04045(.dina(n21307), .dinb(n21306), .dout(n21308));
  jor  g04046(.dina(n21308), .dinb(n21160), .dout(n21309));
  jxor g04047(.dina(n21154), .dinb(n347), .dout(n21310));
  jand g04048(.dina(n21310), .dinb(n21309), .dout(n21311));
  jor  g04049(.dina(n21311), .dinb(n21155), .dout(n21312));
  jxor g04050(.dina(n21149), .dinb(n348), .dout(n21313));
  jand g04051(.dina(n21313), .dinb(n21312), .dout(n21314));
  jor  g04052(.dina(n21314), .dinb(n21150), .dout(n21315));
  jxor g04053(.dina(n21144), .dinb(n349), .dout(n21316));
  jand g04054(.dina(n21316), .dinb(n21315), .dout(n21317));
  jor  g04055(.dina(n21317), .dinb(n21145), .dout(n21318));
  jxor g04056(.dina(n21131), .dinb(n268), .dout(n21319));
  jand g04057(.dina(n21319), .dinb(n21318), .dout(n21320));
  jor  g04058(.dina(n21320), .dinb(n21140), .dout(n21321));
  jand g04059(.dina(n21321), .dinb(n21139), .dout(n21322));
  jor  g04060(.dina(n21322), .dinb(n21136), .dout(n21323));
  jand g04061(.dina(n21323), .dinb(n415), .dout(n21324));
  jor  g04062(.dina(n21324), .dinb(n21131), .dout(n21325));
  jnot g04063(.din(n21324), .dout(n21326));
  jxor g04064(.dina(n21319), .dinb(n21318), .dout(n21327));
  jor  g04065(.dina(n21327), .dinb(n21326), .dout(n21328));
  jand g04066(.dina(n21328), .dinb(n21325), .dout(n21329));
  jand g04067(.dina(n21326), .dinb(n21135), .dout(n21330));
  jand g04068(.dina(n21321), .dinb(n21136), .dout(n21331));
  jor  g04069(.dina(n21331), .dinb(n21330), .dout(n21332));
  jand g04070(.dina(n21332), .dinb(n269), .dout(n21333));
  jnot g04071(.din(n21332), .dout(n21334));
  jand g04072(.dina(n21334), .dinb(b25 ), .dout(n21335));
  jnot g04073(.din(n21335), .dout(n21336));
  jand g04074(.dina(n21329), .dinb(n274), .dout(n21337));
  jor  g04075(.dina(n21324), .dinb(n21144), .dout(n21338));
  jxor g04076(.dina(n21316), .dinb(n21315), .dout(n21339));
  jor  g04077(.dina(n21339), .dinb(n21326), .dout(n21340));
  jand g04078(.dina(n21340), .dinb(n21338), .dout(n21341));
  jand g04079(.dina(n21341), .dinb(n268), .dout(n21342));
  jor  g04080(.dina(n21324), .dinb(n21149), .dout(n21343));
  jxor g04081(.dina(n21313), .dinb(n21312), .dout(n21344));
  jor  g04082(.dina(n21344), .dinb(n21326), .dout(n21345));
  jand g04083(.dina(n21345), .dinb(n21343), .dout(n21346));
  jand g04084(.dina(n21346), .dinb(n349), .dout(n21347));
  jor  g04085(.dina(n21324), .dinb(n21154), .dout(n21348));
  jxor g04086(.dina(n21310), .dinb(n21309), .dout(n21349));
  jor  g04087(.dina(n21349), .dinb(n21326), .dout(n21350));
  jand g04088(.dina(n21350), .dinb(n21348), .dout(n21351));
  jand g04089(.dina(n21351), .dinb(n348), .dout(n21352));
  jor  g04090(.dina(n21324), .dinb(n21159), .dout(n21353));
  jxor g04091(.dina(n21307), .dinb(n21306), .dout(n21354));
  jor  g04092(.dina(n21354), .dinb(n21326), .dout(n21355));
  jand g04093(.dina(n21355), .dinb(n21353), .dout(n21356));
  jand g04094(.dina(n21356), .dinb(n347), .dout(n21357));
  jor  g04095(.dina(n21324), .dinb(n21164), .dout(n21358));
  jxor g04096(.dina(n21304), .dinb(n21303), .dout(n21359));
  jor  g04097(.dina(n21359), .dinb(n21326), .dout(n21360));
  jand g04098(.dina(n21360), .dinb(n21358), .dout(n21361));
  jand g04099(.dina(n21361), .dinb(n267), .dout(n21362));
  jor  g04100(.dina(n21324), .dinb(n21169), .dout(n21363));
  jxor g04101(.dina(n21301), .dinb(n21300), .dout(n21364));
  jor  g04102(.dina(n21364), .dinb(n21326), .dout(n21365));
  jand g04103(.dina(n21365), .dinb(n21363), .dout(n21366));
  jand g04104(.dina(n21366), .dinb(n266), .dout(n21367));
  jor  g04105(.dina(n21324), .dinb(n21174), .dout(n21368));
  jxor g04106(.dina(n21298), .dinb(n21297), .dout(n21369));
  jor  g04107(.dina(n21369), .dinb(n21326), .dout(n21370));
  jand g04108(.dina(n21370), .dinb(n21368), .dout(n21371));
  jand g04109(.dina(n21371), .dinb(n356), .dout(n21372));
  jor  g04110(.dina(n21324), .dinb(n21179), .dout(n21373));
  jxor g04111(.dina(n21295), .dinb(n21294), .dout(n21374));
  jor  g04112(.dina(n21374), .dinb(n21326), .dout(n21375));
  jand g04113(.dina(n21375), .dinb(n21373), .dout(n21376));
  jand g04114(.dina(n21376), .dinb(n355), .dout(n21377));
  jor  g04115(.dina(n21324), .dinb(n21184), .dout(n21378));
  jxor g04116(.dina(n21292), .dinb(n21291), .dout(n21379));
  jor  g04117(.dina(n21379), .dinb(n21326), .dout(n21380));
  jand g04118(.dina(n21380), .dinb(n21378), .dout(n21381));
  jand g04119(.dina(n21381), .dinb(n364), .dout(n21382));
  jor  g04120(.dina(n21324), .dinb(n21189), .dout(n21383));
  jxor g04121(.dina(n21289), .dinb(n21288), .dout(n21384));
  jor  g04122(.dina(n21384), .dinb(n21326), .dout(n21385));
  jand g04123(.dina(n21385), .dinb(n21383), .dout(n21386));
  jand g04124(.dina(n21386), .dinb(n361), .dout(n21387));
  jor  g04125(.dina(n21324), .dinb(n21194), .dout(n21388));
  jxor g04126(.dina(n21286), .dinb(n21285), .dout(n21389));
  jor  g04127(.dina(n21389), .dinb(n21326), .dout(n21390));
  jand g04128(.dina(n21390), .dinb(n21388), .dout(n21391));
  jand g04129(.dina(n21391), .dinb(n360), .dout(n21392));
  jor  g04130(.dina(n21324), .dinb(n21199), .dout(n21393));
  jxor g04131(.dina(n21283), .dinb(n21282), .dout(n21394));
  jor  g04132(.dina(n21394), .dinb(n21326), .dout(n21395));
  jand g04133(.dina(n21395), .dinb(n21393), .dout(n21396));
  jand g04134(.dina(n21396), .dinb(n363), .dout(n21397));
  jor  g04135(.dina(n21324), .dinb(n21204), .dout(n21398));
  jxor g04136(.dina(n21280), .dinb(n21279), .dout(n21399));
  jor  g04137(.dina(n21399), .dinb(n21326), .dout(n21400));
  jand g04138(.dina(n21400), .dinb(n21398), .dout(n21401));
  jand g04139(.dina(n21401), .dinb(n359), .dout(n21402));
  jor  g04140(.dina(n21324), .dinb(n21209), .dout(n21403));
  jxor g04141(.dina(n21277), .dinb(n21276), .dout(n21404));
  jor  g04142(.dina(n21404), .dinb(n21326), .dout(n21405));
  jand g04143(.dina(n21405), .dinb(n21403), .dout(n21406));
  jand g04144(.dina(n21406), .dinb(n369), .dout(n21407));
  jor  g04145(.dina(n21324), .dinb(n21214), .dout(n21408));
  jxor g04146(.dina(n21274), .dinb(n21273), .dout(n21409));
  jor  g04147(.dina(n21409), .dinb(n21326), .dout(n21410));
  jand g04148(.dina(n21410), .dinb(n21408), .dout(n21411));
  jand g04149(.dina(n21411), .dinb(n368), .dout(n21412));
  jor  g04150(.dina(n21324), .dinb(n21219), .dout(n21413));
  jxor g04151(.dina(n21271), .dinb(n21270), .dout(n21414));
  jor  g04152(.dina(n21414), .dinb(n21326), .dout(n21415));
  jand g04153(.dina(n21415), .dinb(n21413), .dout(n21416));
  jand g04154(.dina(n21416), .dinb(n367), .dout(n21417));
  jor  g04155(.dina(n21324), .dinb(n21224), .dout(n21418));
  jxor g04156(.dina(n21268), .dinb(n21267), .dout(n21419));
  jor  g04157(.dina(n21419), .dinb(n21326), .dout(n21420));
  jand g04158(.dina(n21420), .dinb(n21418), .dout(n21421));
  jand g04159(.dina(n21421), .dinb(n265), .dout(n21422));
  jor  g04160(.dina(n21324), .dinb(n21229), .dout(n21423));
  jxor g04161(.dina(n21265), .dinb(n21264), .dout(n21424));
  jor  g04162(.dina(n21424), .dinb(n21326), .dout(n21425));
  jand g04163(.dina(n21425), .dinb(n21423), .dout(n21426));
  jand g04164(.dina(n21426), .dinb(n378), .dout(n21427));
  jor  g04165(.dina(n21324), .dinb(n21234), .dout(n21428));
  jxor g04166(.dina(n21262), .dinb(n21261), .dout(n21429));
  jor  g04167(.dina(n21429), .dinb(n21326), .dout(n21430));
  jand g04168(.dina(n21430), .dinb(n21428), .dout(n21431));
  jand g04169(.dina(n21431), .dinb(n377), .dout(n21432));
  jand g04170(.dina(n21326), .dinb(n21241), .dout(n21433));
  jnot g04171(.din(n21433), .dout(n21434));
  jxor g04172(.dina(n21259), .dinb(n21258), .dout(n21435));
  jor  g04173(.dina(n21435), .dinb(n21326), .dout(n21436));
  jand g04174(.dina(n21436), .dinb(n21434), .dout(n21437));
  jand g04175(.dina(n21437), .dinb(n376), .dout(n21438));
  jor  g04176(.dina(n21324), .dinb(n21247), .dout(n21439));
  jxor g04177(.dina(n21256), .dinb(n21255), .dout(n21440));
  jor  g04178(.dina(n21440), .dinb(n21326), .dout(n21441));
  jand g04179(.dina(n21441), .dinb(n21439), .dout(n21442));
  jand g04180(.dina(n21442), .dinb(n264), .dout(n21443));
  jor  g04181(.dina(n21324), .dinb(n21252), .dout(n21444));
  jxor g04182(.dina(n21253), .dinb(n3078), .dout(n21445));
  jand g04183(.dina(n21445), .dinb(n21324), .dout(n21446));
  jnot g04184(.din(n21446), .dout(n21447));
  jand g04185(.dina(n21447), .dinb(n21444), .dout(n21448));
  jor  g04186(.dina(n21448), .dinb(b2 ), .dout(n21449));
  jnot g04187(.din(n21449), .dout(n21450));
  jnot g04188(.din(n3302), .dout(n21451));
  jnot g04189(.din(n21136), .dout(n21452));
  jnot g04190(.din(n21140), .dout(n21453));
  jnot g04191(.din(n21145), .dout(n21454));
  jnot g04192(.din(n21150), .dout(n21455));
  jnot g04193(.din(n21155), .dout(n21456));
  jnot g04194(.din(n21160), .dout(n21457));
  jnot g04195(.din(n21165), .dout(n21458));
  jnot g04196(.din(n21170), .dout(n21459));
  jnot g04197(.din(n21175), .dout(n21460));
  jnot g04198(.din(n21180), .dout(n21461));
  jnot g04199(.din(n21185), .dout(n21462));
  jnot g04200(.din(n21190), .dout(n21463));
  jnot g04201(.din(n21195), .dout(n21464));
  jnot g04202(.din(n21200), .dout(n21465));
  jnot g04203(.din(n21205), .dout(n21466));
  jnot g04204(.din(n21210), .dout(n21467));
  jnot g04205(.din(n21215), .dout(n21468));
  jnot g04206(.din(n21220), .dout(n21469));
  jnot g04207(.din(n21225), .dout(n21470));
  jnot g04208(.din(n21230), .dout(n21471));
  jnot g04209(.din(n21235), .dout(n21472));
  jnot g04210(.din(n21243), .dout(n21473));
  jnot g04211(.din(n21248), .dout(n21474));
  jnot g04212(.din(n21251), .dout(n21475));
  jxor g04213(.dina(n21252), .dinb(n259), .dout(n21476));
  jor  g04214(.dina(n21476), .dinb(n3077), .dout(n21477));
  jand g04215(.dina(n21477), .dinb(n21475), .dout(n21478));
  jnot g04216(.din(n21256), .dout(n21479));
  jor  g04217(.dina(n21479), .dinb(n21478), .dout(n21480));
  jand g04218(.dina(n21480), .dinb(n21474), .dout(n21481));
  jnot g04219(.din(n21259), .dout(n21482));
  jor  g04220(.dina(n21482), .dinb(n21481), .dout(n21483));
  jand g04221(.dina(n21483), .dinb(n21473), .dout(n21484));
  jnot g04222(.din(n21262), .dout(n21485));
  jor  g04223(.dina(n21485), .dinb(n21484), .dout(n21486));
  jand g04224(.dina(n21486), .dinb(n21472), .dout(n21487));
  jnot g04225(.din(n21265), .dout(n21488));
  jor  g04226(.dina(n21488), .dinb(n21487), .dout(n21489));
  jand g04227(.dina(n21489), .dinb(n21471), .dout(n21490));
  jnot g04228(.din(n21268), .dout(n21491));
  jor  g04229(.dina(n21491), .dinb(n21490), .dout(n21492));
  jand g04230(.dina(n21492), .dinb(n21470), .dout(n21493));
  jnot g04231(.din(n21271), .dout(n21494));
  jor  g04232(.dina(n21494), .dinb(n21493), .dout(n21495));
  jand g04233(.dina(n21495), .dinb(n21469), .dout(n21496));
  jnot g04234(.din(n21274), .dout(n21497));
  jor  g04235(.dina(n21497), .dinb(n21496), .dout(n21498));
  jand g04236(.dina(n21498), .dinb(n21468), .dout(n21499));
  jnot g04237(.din(n21277), .dout(n21500));
  jor  g04238(.dina(n21500), .dinb(n21499), .dout(n21501));
  jand g04239(.dina(n21501), .dinb(n21467), .dout(n21502));
  jnot g04240(.din(n21280), .dout(n21503));
  jor  g04241(.dina(n21503), .dinb(n21502), .dout(n21504));
  jand g04242(.dina(n21504), .dinb(n21466), .dout(n21505));
  jnot g04243(.din(n21283), .dout(n21506));
  jor  g04244(.dina(n21506), .dinb(n21505), .dout(n21507));
  jand g04245(.dina(n21507), .dinb(n21465), .dout(n21508));
  jnot g04246(.din(n21286), .dout(n21509));
  jor  g04247(.dina(n21509), .dinb(n21508), .dout(n21510));
  jand g04248(.dina(n21510), .dinb(n21464), .dout(n21511));
  jnot g04249(.din(n21289), .dout(n21512));
  jor  g04250(.dina(n21512), .dinb(n21511), .dout(n21513));
  jand g04251(.dina(n21513), .dinb(n21463), .dout(n21514));
  jnot g04252(.din(n21292), .dout(n21515));
  jor  g04253(.dina(n21515), .dinb(n21514), .dout(n21516));
  jand g04254(.dina(n21516), .dinb(n21462), .dout(n21517));
  jnot g04255(.din(n21295), .dout(n21518));
  jor  g04256(.dina(n21518), .dinb(n21517), .dout(n21519));
  jand g04257(.dina(n21519), .dinb(n21461), .dout(n21520));
  jnot g04258(.din(n21298), .dout(n21521));
  jor  g04259(.dina(n21521), .dinb(n21520), .dout(n21522));
  jand g04260(.dina(n21522), .dinb(n21460), .dout(n21523));
  jnot g04261(.din(n21301), .dout(n21524));
  jor  g04262(.dina(n21524), .dinb(n21523), .dout(n21525));
  jand g04263(.dina(n21525), .dinb(n21459), .dout(n21526));
  jnot g04264(.din(n21304), .dout(n21527));
  jor  g04265(.dina(n21527), .dinb(n21526), .dout(n21528));
  jand g04266(.dina(n21528), .dinb(n21458), .dout(n21529));
  jnot g04267(.din(n21307), .dout(n21530));
  jor  g04268(.dina(n21530), .dinb(n21529), .dout(n21531));
  jand g04269(.dina(n21531), .dinb(n21457), .dout(n21532));
  jnot g04270(.din(n21310), .dout(n21533));
  jor  g04271(.dina(n21533), .dinb(n21532), .dout(n21534));
  jand g04272(.dina(n21534), .dinb(n21456), .dout(n21535));
  jnot g04273(.din(n21313), .dout(n21536));
  jor  g04274(.dina(n21536), .dinb(n21535), .dout(n21537));
  jand g04275(.dina(n21537), .dinb(n21455), .dout(n21538));
  jnot g04276(.din(n21316), .dout(n21539));
  jor  g04277(.dina(n21539), .dinb(n21538), .dout(n21540));
  jand g04278(.dina(n21540), .dinb(n21454), .dout(n21541));
  jnot g04279(.din(n21319), .dout(n21542));
  jor  g04280(.dina(n21542), .dinb(n21541), .dout(n21543));
  jand g04281(.dina(n21543), .dinb(n21453), .dout(n21544));
  jor  g04282(.dina(n21544), .dinb(n21138), .dout(n21545));
  jand g04283(.dina(n21545), .dinb(n21452), .dout(n21546));
  jor  g04284(.dina(n21546), .dinb(n21451), .dout(n21547));
  jand g04285(.dina(n21547), .dinb(a39 ), .dout(n21548));
  jnot g04286(.din(n3305), .dout(n21549));
  jor  g04287(.dina(n21546), .dinb(n21549), .dout(n21550));
  jnot g04288(.din(n21550), .dout(n21551));
  jor  g04289(.dina(n21551), .dinb(n21548), .dout(n21552));
  jand g04290(.dina(n21552), .dinb(n259), .dout(n21553));
  jand g04291(.dina(n21323), .dinb(n3302), .dout(n21554));
  jor  g04292(.dina(n21554), .dinb(n3076), .dout(n21555));
  jand g04293(.dina(n21550), .dinb(n21555), .dout(n21556));
  jxor g04294(.dina(n21556), .dinb(b1 ), .dout(n21557));
  jand g04295(.dina(n21557), .dinb(n3412), .dout(n21558));
  jor  g04296(.dina(n21558), .dinb(n21553), .dout(n21559));
  jxor g04297(.dina(n21448), .dinb(b2 ), .dout(n21560));
  jand g04298(.dina(n21560), .dinb(n21559), .dout(n21561));
  jor  g04299(.dina(n21561), .dinb(n21450), .dout(n21562));
  jxor g04300(.dina(n21442), .dinb(n264), .dout(n21563));
  jand g04301(.dina(n21563), .dinb(n21562), .dout(n21564));
  jor  g04302(.dina(n21564), .dinb(n21443), .dout(n21565));
  jxor g04303(.dina(n21437), .dinb(n376), .dout(n21566));
  jand g04304(.dina(n21566), .dinb(n21565), .dout(n21567));
  jor  g04305(.dina(n21567), .dinb(n21438), .dout(n21568));
  jxor g04306(.dina(n21431), .dinb(n377), .dout(n21569));
  jand g04307(.dina(n21569), .dinb(n21568), .dout(n21570));
  jor  g04308(.dina(n21570), .dinb(n21432), .dout(n21571));
  jxor g04309(.dina(n21426), .dinb(n378), .dout(n21572));
  jand g04310(.dina(n21572), .dinb(n21571), .dout(n21573));
  jor  g04311(.dina(n21573), .dinb(n21427), .dout(n21574));
  jxor g04312(.dina(n21421), .dinb(n265), .dout(n21575));
  jand g04313(.dina(n21575), .dinb(n21574), .dout(n21576));
  jor  g04314(.dina(n21576), .dinb(n21422), .dout(n21577));
  jxor g04315(.dina(n21416), .dinb(n367), .dout(n21578));
  jand g04316(.dina(n21578), .dinb(n21577), .dout(n21579));
  jor  g04317(.dina(n21579), .dinb(n21417), .dout(n21580));
  jxor g04318(.dina(n21411), .dinb(n368), .dout(n21581));
  jand g04319(.dina(n21581), .dinb(n21580), .dout(n21582));
  jor  g04320(.dina(n21582), .dinb(n21412), .dout(n21583));
  jxor g04321(.dina(n21406), .dinb(n369), .dout(n21584));
  jand g04322(.dina(n21584), .dinb(n21583), .dout(n21585));
  jor  g04323(.dina(n21585), .dinb(n21407), .dout(n21586));
  jxor g04324(.dina(n21401), .dinb(n359), .dout(n21587));
  jand g04325(.dina(n21587), .dinb(n21586), .dout(n21588));
  jor  g04326(.dina(n21588), .dinb(n21402), .dout(n21589));
  jxor g04327(.dina(n21396), .dinb(n363), .dout(n21590));
  jand g04328(.dina(n21590), .dinb(n21589), .dout(n21591));
  jor  g04329(.dina(n21591), .dinb(n21397), .dout(n21592));
  jxor g04330(.dina(n21391), .dinb(n360), .dout(n21593));
  jand g04331(.dina(n21593), .dinb(n21592), .dout(n21594));
  jor  g04332(.dina(n21594), .dinb(n21392), .dout(n21595));
  jxor g04333(.dina(n21386), .dinb(n361), .dout(n21596));
  jand g04334(.dina(n21596), .dinb(n21595), .dout(n21597));
  jor  g04335(.dina(n21597), .dinb(n21387), .dout(n21598));
  jxor g04336(.dina(n21381), .dinb(n364), .dout(n21599));
  jand g04337(.dina(n21599), .dinb(n21598), .dout(n21600));
  jor  g04338(.dina(n21600), .dinb(n21382), .dout(n21601));
  jxor g04339(.dina(n21376), .dinb(n355), .dout(n21602));
  jand g04340(.dina(n21602), .dinb(n21601), .dout(n21603));
  jor  g04341(.dina(n21603), .dinb(n21377), .dout(n21604));
  jxor g04342(.dina(n21371), .dinb(n356), .dout(n21605));
  jand g04343(.dina(n21605), .dinb(n21604), .dout(n21606));
  jor  g04344(.dina(n21606), .dinb(n21372), .dout(n21607));
  jxor g04345(.dina(n21366), .dinb(n266), .dout(n21608));
  jand g04346(.dina(n21608), .dinb(n21607), .dout(n21609));
  jor  g04347(.dina(n21609), .dinb(n21367), .dout(n21610));
  jxor g04348(.dina(n21361), .dinb(n267), .dout(n21611));
  jand g04349(.dina(n21611), .dinb(n21610), .dout(n21612));
  jor  g04350(.dina(n21612), .dinb(n21362), .dout(n21613));
  jxor g04351(.dina(n21356), .dinb(n347), .dout(n21614));
  jand g04352(.dina(n21614), .dinb(n21613), .dout(n21615));
  jor  g04353(.dina(n21615), .dinb(n21357), .dout(n21616));
  jxor g04354(.dina(n21351), .dinb(n348), .dout(n21617));
  jand g04355(.dina(n21617), .dinb(n21616), .dout(n21618));
  jor  g04356(.dina(n21618), .dinb(n21352), .dout(n21619));
  jxor g04357(.dina(n21346), .dinb(n349), .dout(n21620));
  jand g04358(.dina(n21620), .dinb(n21619), .dout(n21621));
  jor  g04359(.dina(n21621), .dinb(n21347), .dout(n21622));
  jxor g04360(.dina(n21341), .dinb(n268), .dout(n21623));
  jand g04361(.dina(n21623), .dinb(n21622), .dout(n21624));
  jor  g04362(.dina(n21624), .dinb(n21342), .dout(n21625));
  jxor g04363(.dina(n21329), .dinb(n274), .dout(n21626));
  jand g04364(.dina(n21626), .dinb(n21625), .dout(n21627));
  jor  g04365(.dina(n21627), .dinb(n21337), .dout(n21628));
  jand g04366(.dina(n21628), .dinb(n21336), .dout(n21629));
  jor  g04367(.dina(n21629), .dinb(n21333), .dout(n21630));
  jand g04368(.dina(n21630), .dinb(n3157), .dout(n21631));
  jor  g04369(.dina(n21631), .dinb(n21329), .dout(n21632));
  jnot g04370(.din(n21333), .dout(n21633));
  jnot g04371(.din(n21337), .dout(n21634));
  jnot g04372(.din(n21342), .dout(n21635));
  jnot g04373(.din(n21347), .dout(n21636));
  jnot g04374(.din(n21352), .dout(n21637));
  jnot g04375(.din(n21357), .dout(n21638));
  jnot g04376(.din(n21362), .dout(n21639));
  jnot g04377(.din(n21367), .dout(n21640));
  jnot g04378(.din(n21372), .dout(n21641));
  jnot g04379(.din(n21377), .dout(n21642));
  jnot g04380(.din(n21382), .dout(n21643));
  jnot g04381(.din(n21387), .dout(n21644));
  jnot g04382(.din(n21392), .dout(n21645));
  jnot g04383(.din(n21397), .dout(n21646));
  jnot g04384(.din(n21402), .dout(n21647));
  jnot g04385(.din(n21407), .dout(n21648));
  jnot g04386(.din(n21412), .dout(n21649));
  jnot g04387(.din(n21417), .dout(n21650));
  jnot g04388(.din(n21422), .dout(n21651));
  jnot g04389(.din(n21427), .dout(n21652));
  jnot g04390(.din(n21432), .dout(n21653));
  jnot g04391(.din(n21438), .dout(n21654));
  jnot g04392(.din(n21443), .dout(n21655));
  jor  g04393(.dina(n21556), .dinb(b1 ), .dout(n21656));
  jxor g04394(.dina(n21556), .dinb(n259), .dout(n21657));
  jor  g04395(.dina(n21657), .dinb(n3311), .dout(n21658));
  jand g04396(.dina(n21658), .dinb(n21656), .dout(n21659));
  jxor g04397(.dina(n21448), .dinb(n386), .dout(n21660));
  jor  g04398(.dina(n21660), .dinb(n21659), .dout(n21661));
  jand g04399(.dina(n21661), .dinb(n21449), .dout(n21662));
  jnot g04400(.din(n21563), .dout(n21663));
  jor  g04401(.dina(n21663), .dinb(n21662), .dout(n21664));
  jand g04402(.dina(n21664), .dinb(n21655), .dout(n21665));
  jnot g04403(.din(n21566), .dout(n21666));
  jor  g04404(.dina(n21666), .dinb(n21665), .dout(n21667));
  jand g04405(.dina(n21667), .dinb(n21654), .dout(n21668));
  jnot g04406(.din(n21569), .dout(n21669));
  jor  g04407(.dina(n21669), .dinb(n21668), .dout(n21670));
  jand g04408(.dina(n21670), .dinb(n21653), .dout(n21671));
  jnot g04409(.din(n21572), .dout(n21672));
  jor  g04410(.dina(n21672), .dinb(n21671), .dout(n21673));
  jand g04411(.dina(n21673), .dinb(n21652), .dout(n21674));
  jnot g04412(.din(n21575), .dout(n21675));
  jor  g04413(.dina(n21675), .dinb(n21674), .dout(n21676));
  jand g04414(.dina(n21676), .dinb(n21651), .dout(n21677));
  jnot g04415(.din(n21578), .dout(n21678));
  jor  g04416(.dina(n21678), .dinb(n21677), .dout(n21679));
  jand g04417(.dina(n21679), .dinb(n21650), .dout(n21680));
  jnot g04418(.din(n21581), .dout(n21681));
  jor  g04419(.dina(n21681), .dinb(n21680), .dout(n21682));
  jand g04420(.dina(n21682), .dinb(n21649), .dout(n21683));
  jnot g04421(.din(n21584), .dout(n21684));
  jor  g04422(.dina(n21684), .dinb(n21683), .dout(n21685));
  jand g04423(.dina(n21685), .dinb(n21648), .dout(n21686));
  jnot g04424(.din(n21587), .dout(n21687));
  jor  g04425(.dina(n21687), .dinb(n21686), .dout(n21688));
  jand g04426(.dina(n21688), .dinb(n21647), .dout(n21689));
  jnot g04427(.din(n21590), .dout(n21690));
  jor  g04428(.dina(n21690), .dinb(n21689), .dout(n21691));
  jand g04429(.dina(n21691), .dinb(n21646), .dout(n21692));
  jnot g04430(.din(n21593), .dout(n21693));
  jor  g04431(.dina(n21693), .dinb(n21692), .dout(n21694));
  jand g04432(.dina(n21694), .dinb(n21645), .dout(n21695));
  jnot g04433(.din(n21596), .dout(n21696));
  jor  g04434(.dina(n21696), .dinb(n21695), .dout(n21697));
  jand g04435(.dina(n21697), .dinb(n21644), .dout(n21698));
  jnot g04436(.din(n21599), .dout(n21699));
  jor  g04437(.dina(n21699), .dinb(n21698), .dout(n21700));
  jand g04438(.dina(n21700), .dinb(n21643), .dout(n21701));
  jnot g04439(.din(n21602), .dout(n21702));
  jor  g04440(.dina(n21702), .dinb(n21701), .dout(n21703));
  jand g04441(.dina(n21703), .dinb(n21642), .dout(n21704));
  jnot g04442(.din(n21605), .dout(n21705));
  jor  g04443(.dina(n21705), .dinb(n21704), .dout(n21706));
  jand g04444(.dina(n21706), .dinb(n21641), .dout(n21707));
  jnot g04445(.din(n21608), .dout(n21708));
  jor  g04446(.dina(n21708), .dinb(n21707), .dout(n21709));
  jand g04447(.dina(n21709), .dinb(n21640), .dout(n21710));
  jnot g04448(.din(n21611), .dout(n21711));
  jor  g04449(.dina(n21711), .dinb(n21710), .dout(n21712));
  jand g04450(.dina(n21712), .dinb(n21639), .dout(n21713));
  jnot g04451(.din(n21614), .dout(n21714));
  jor  g04452(.dina(n21714), .dinb(n21713), .dout(n21715));
  jand g04453(.dina(n21715), .dinb(n21638), .dout(n21716));
  jnot g04454(.din(n21617), .dout(n21717));
  jor  g04455(.dina(n21717), .dinb(n21716), .dout(n21718));
  jand g04456(.dina(n21718), .dinb(n21637), .dout(n21719));
  jnot g04457(.din(n21620), .dout(n21720));
  jor  g04458(.dina(n21720), .dinb(n21719), .dout(n21721));
  jand g04459(.dina(n21721), .dinb(n21636), .dout(n21722));
  jnot g04460(.din(n21623), .dout(n21723));
  jor  g04461(.dina(n21723), .dinb(n21722), .dout(n21724));
  jand g04462(.dina(n21724), .dinb(n21635), .dout(n21725));
  jnot g04463(.din(n21626), .dout(n21726));
  jor  g04464(.dina(n21726), .dinb(n21725), .dout(n21727));
  jand g04465(.dina(n21727), .dinb(n21634), .dout(n21728));
  jor  g04466(.dina(n21728), .dinb(n21335), .dout(n21729));
  jand g04467(.dina(n21729), .dinb(n21633), .dout(n21730));
  jor  g04468(.dina(n21730), .dinb(n3158), .dout(n21731));
  jxor g04469(.dina(n21626), .dinb(n21625), .dout(n21732));
  jor  g04470(.dina(n21732), .dinb(n21731), .dout(n21733));
  jand g04471(.dina(n21733), .dinb(n21632), .dout(n21734));
  jand g04472(.dina(n21734), .dinb(n269), .dout(n21735));
  jor  g04473(.dina(n21631), .dinb(n21341), .dout(n21736));
  jxor g04474(.dina(n21623), .dinb(n21622), .dout(n21737));
  jor  g04475(.dina(n21737), .dinb(n21731), .dout(n21738));
  jand g04476(.dina(n21738), .dinb(n21736), .dout(n21739));
  jand g04477(.dina(n21739), .dinb(n274), .dout(n21740));
  jor  g04478(.dina(n21631), .dinb(n21346), .dout(n21741));
  jxor g04479(.dina(n21620), .dinb(n21619), .dout(n21742));
  jor  g04480(.dina(n21742), .dinb(n21731), .dout(n21743));
  jand g04481(.dina(n21743), .dinb(n21741), .dout(n21744));
  jand g04482(.dina(n21744), .dinb(n268), .dout(n21745));
  jor  g04483(.dina(n21631), .dinb(n21351), .dout(n21746));
  jxor g04484(.dina(n21617), .dinb(n21616), .dout(n21747));
  jor  g04485(.dina(n21747), .dinb(n21731), .dout(n21748));
  jand g04486(.dina(n21748), .dinb(n21746), .dout(n21749));
  jand g04487(.dina(n21749), .dinb(n349), .dout(n21750));
  jor  g04488(.dina(n21631), .dinb(n21356), .dout(n21751));
  jxor g04489(.dina(n21614), .dinb(n21613), .dout(n21752));
  jor  g04490(.dina(n21752), .dinb(n21731), .dout(n21753));
  jand g04491(.dina(n21753), .dinb(n21751), .dout(n21754));
  jand g04492(.dina(n21754), .dinb(n348), .dout(n21755));
  jor  g04493(.dina(n21631), .dinb(n21361), .dout(n21756));
  jxor g04494(.dina(n21611), .dinb(n21610), .dout(n21757));
  jor  g04495(.dina(n21757), .dinb(n21731), .dout(n21758));
  jand g04496(.dina(n21758), .dinb(n21756), .dout(n21759));
  jand g04497(.dina(n21759), .dinb(n347), .dout(n21760));
  jor  g04498(.dina(n21631), .dinb(n21366), .dout(n21761));
  jxor g04499(.dina(n21608), .dinb(n21607), .dout(n21762));
  jor  g04500(.dina(n21762), .dinb(n21731), .dout(n21763));
  jand g04501(.dina(n21763), .dinb(n21761), .dout(n21764));
  jand g04502(.dina(n21764), .dinb(n267), .dout(n21765));
  jor  g04503(.dina(n21631), .dinb(n21371), .dout(n21766));
  jxor g04504(.dina(n21605), .dinb(n21604), .dout(n21767));
  jor  g04505(.dina(n21767), .dinb(n21731), .dout(n21768));
  jand g04506(.dina(n21768), .dinb(n21766), .dout(n21769));
  jand g04507(.dina(n21769), .dinb(n266), .dout(n21770));
  jor  g04508(.dina(n21631), .dinb(n21376), .dout(n21771));
  jxor g04509(.dina(n21602), .dinb(n21601), .dout(n21772));
  jor  g04510(.dina(n21772), .dinb(n21731), .dout(n21773));
  jand g04511(.dina(n21773), .dinb(n21771), .dout(n21774));
  jand g04512(.dina(n21774), .dinb(n356), .dout(n21775));
  jor  g04513(.dina(n21631), .dinb(n21381), .dout(n21776));
  jxor g04514(.dina(n21599), .dinb(n21598), .dout(n21777));
  jor  g04515(.dina(n21777), .dinb(n21731), .dout(n21778));
  jand g04516(.dina(n21778), .dinb(n21776), .dout(n21779));
  jand g04517(.dina(n21779), .dinb(n355), .dout(n21780));
  jor  g04518(.dina(n21631), .dinb(n21386), .dout(n21781));
  jxor g04519(.dina(n21596), .dinb(n21595), .dout(n21782));
  jor  g04520(.dina(n21782), .dinb(n21731), .dout(n21783));
  jand g04521(.dina(n21783), .dinb(n21781), .dout(n21784));
  jand g04522(.dina(n21784), .dinb(n364), .dout(n21785));
  jor  g04523(.dina(n21631), .dinb(n21391), .dout(n21786));
  jxor g04524(.dina(n21593), .dinb(n21592), .dout(n21787));
  jor  g04525(.dina(n21787), .dinb(n21731), .dout(n21788));
  jand g04526(.dina(n21788), .dinb(n21786), .dout(n21789));
  jand g04527(.dina(n21789), .dinb(n361), .dout(n21790));
  jor  g04528(.dina(n21631), .dinb(n21396), .dout(n21791));
  jxor g04529(.dina(n21590), .dinb(n21589), .dout(n21792));
  jor  g04530(.dina(n21792), .dinb(n21731), .dout(n21793));
  jand g04531(.dina(n21793), .dinb(n21791), .dout(n21794));
  jand g04532(.dina(n21794), .dinb(n360), .dout(n21795));
  jor  g04533(.dina(n21631), .dinb(n21401), .dout(n21796));
  jxor g04534(.dina(n21587), .dinb(n21586), .dout(n21797));
  jor  g04535(.dina(n21797), .dinb(n21731), .dout(n21798));
  jand g04536(.dina(n21798), .dinb(n21796), .dout(n21799));
  jand g04537(.dina(n21799), .dinb(n363), .dout(n21800));
  jor  g04538(.dina(n21631), .dinb(n21406), .dout(n21801));
  jxor g04539(.dina(n21584), .dinb(n21583), .dout(n21802));
  jor  g04540(.dina(n21802), .dinb(n21731), .dout(n21803));
  jand g04541(.dina(n21803), .dinb(n21801), .dout(n21804));
  jand g04542(.dina(n21804), .dinb(n359), .dout(n21805));
  jor  g04543(.dina(n21631), .dinb(n21411), .dout(n21806));
  jxor g04544(.dina(n21581), .dinb(n21580), .dout(n21807));
  jor  g04545(.dina(n21807), .dinb(n21731), .dout(n21808));
  jand g04546(.dina(n21808), .dinb(n21806), .dout(n21809));
  jand g04547(.dina(n21809), .dinb(n369), .dout(n21810));
  jor  g04548(.dina(n21631), .dinb(n21416), .dout(n21811));
  jxor g04549(.dina(n21578), .dinb(n21577), .dout(n21812));
  jor  g04550(.dina(n21812), .dinb(n21731), .dout(n21813));
  jand g04551(.dina(n21813), .dinb(n21811), .dout(n21814));
  jand g04552(.dina(n21814), .dinb(n368), .dout(n21815));
  jor  g04553(.dina(n21631), .dinb(n21421), .dout(n21816));
  jxor g04554(.dina(n21575), .dinb(n21574), .dout(n21817));
  jor  g04555(.dina(n21817), .dinb(n21731), .dout(n21818));
  jand g04556(.dina(n21818), .dinb(n21816), .dout(n21819));
  jand g04557(.dina(n21819), .dinb(n367), .dout(n21820));
  jor  g04558(.dina(n21631), .dinb(n21426), .dout(n21821));
  jxor g04559(.dina(n21572), .dinb(n21571), .dout(n21822));
  jor  g04560(.dina(n21822), .dinb(n21731), .dout(n21823));
  jand g04561(.dina(n21823), .dinb(n21821), .dout(n21824));
  jand g04562(.dina(n21824), .dinb(n265), .dout(n21825));
  jor  g04563(.dina(n21631), .dinb(n21431), .dout(n21826));
  jxor g04564(.dina(n21569), .dinb(n21568), .dout(n21827));
  jor  g04565(.dina(n21827), .dinb(n21731), .dout(n21828));
  jand g04566(.dina(n21828), .dinb(n21826), .dout(n21829));
  jand g04567(.dina(n21829), .dinb(n378), .dout(n21830));
  jor  g04568(.dina(n21631), .dinb(n21437), .dout(n21831));
  jxor g04569(.dina(n21566), .dinb(n21565), .dout(n21832));
  jor  g04570(.dina(n21832), .dinb(n21731), .dout(n21833));
  jand g04571(.dina(n21833), .dinb(n21831), .dout(n21834));
  jand g04572(.dina(n21834), .dinb(n377), .dout(n21835));
  jor  g04573(.dina(n21631), .dinb(n21442), .dout(n21836));
  jxor g04574(.dina(n21563), .dinb(n21562), .dout(n21837));
  jor  g04575(.dina(n21837), .dinb(n21731), .dout(n21838));
  jand g04576(.dina(n21838), .dinb(n21836), .dout(n21839));
  jand g04577(.dina(n21839), .dinb(n376), .dout(n21840));
  jnot g04578(.din(n21448), .dout(n21841));
  jor  g04579(.dina(n21631), .dinb(n21841), .dout(n21842));
  jxor g04580(.dina(n21560), .dinb(n21559), .dout(n21843));
  jor  g04581(.dina(n21843), .dinb(n21731), .dout(n21844));
  jand g04582(.dina(n21844), .dinb(n21842), .dout(n21845));
  jand g04583(.dina(n21845), .dinb(n264), .dout(n21846));
  jand g04584(.dina(n21731), .dinb(n21552), .dout(n21847));
  jxor g04585(.dina(n21557), .dinb(n3412), .dout(n21848));
  jand g04586(.dina(n21848), .dinb(n21631), .dout(n21849));
  jor  g04587(.dina(n21849), .dinb(n21847), .dout(n21850));
  jand g04588(.dina(n21850), .dinb(n386), .dout(n21851));
  jnot g04589(.din(n3593), .dout(n21852));
  jor  g04590(.dina(n21730), .dinb(n21852), .dout(n21853));
  jand g04591(.dina(n21853), .dinb(a38 ), .dout(n21854));
  jand g04592(.dina(n21631), .dinb(n3311), .dout(n21855));
  jor  g04593(.dina(n21855), .dinb(n21854), .dout(n21856));
  jand g04594(.dina(n21856), .dinb(n259), .dout(n21857));
  jand g04595(.dina(n21630), .dinb(n3593), .dout(n21858));
  jor  g04596(.dina(n21858), .dinb(n3310), .dout(n21859));
  jor  g04597(.dina(n21731), .dinb(n3412), .dout(n21860));
  jand g04598(.dina(n21860), .dinb(n21859), .dout(n21861));
  jxor g04599(.dina(n21861), .dinb(b1 ), .dout(n21862));
  jand g04600(.dina(n21862), .dinb(n3602), .dout(n21863));
  jor  g04601(.dina(n21863), .dinb(n21857), .dout(n21864));
  jxor g04602(.dina(n21850), .dinb(n386), .dout(n21865));
  jand g04603(.dina(n21865), .dinb(n21864), .dout(n21866));
  jor  g04604(.dina(n21866), .dinb(n21851), .dout(n21867));
  jxor g04605(.dina(n21845), .dinb(n264), .dout(n21868));
  jand g04606(.dina(n21868), .dinb(n21867), .dout(n21869));
  jor  g04607(.dina(n21869), .dinb(n21846), .dout(n21870));
  jxor g04608(.dina(n21839), .dinb(n376), .dout(n21871));
  jand g04609(.dina(n21871), .dinb(n21870), .dout(n21872));
  jor  g04610(.dina(n21872), .dinb(n21840), .dout(n21873));
  jxor g04611(.dina(n21834), .dinb(n377), .dout(n21874));
  jand g04612(.dina(n21874), .dinb(n21873), .dout(n21875));
  jor  g04613(.dina(n21875), .dinb(n21835), .dout(n21876));
  jxor g04614(.dina(n21829), .dinb(n378), .dout(n21877));
  jand g04615(.dina(n21877), .dinb(n21876), .dout(n21878));
  jor  g04616(.dina(n21878), .dinb(n21830), .dout(n21879));
  jxor g04617(.dina(n21824), .dinb(n265), .dout(n21880));
  jand g04618(.dina(n21880), .dinb(n21879), .dout(n21881));
  jor  g04619(.dina(n21881), .dinb(n21825), .dout(n21882));
  jxor g04620(.dina(n21819), .dinb(n367), .dout(n21883));
  jand g04621(.dina(n21883), .dinb(n21882), .dout(n21884));
  jor  g04622(.dina(n21884), .dinb(n21820), .dout(n21885));
  jxor g04623(.dina(n21814), .dinb(n368), .dout(n21886));
  jand g04624(.dina(n21886), .dinb(n21885), .dout(n21887));
  jor  g04625(.dina(n21887), .dinb(n21815), .dout(n21888));
  jxor g04626(.dina(n21809), .dinb(n369), .dout(n21889));
  jand g04627(.dina(n21889), .dinb(n21888), .dout(n21890));
  jor  g04628(.dina(n21890), .dinb(n21810), .dout(n21891));
  jxor g04629(.dina(n21804), .dinb(n359), .dout(n21892));
  jand g04630(.dina(n21892), .dinb(n21891), .dout(n21893));
  jor  g04631(.dina(n21893), .dinb(n21805), .dout(n21894));
  jxor g04632(.dina(n21799), .dinb(n363), .dout(n21895));
  jand g04633(.dina(n21895), .dinb(n21894), .dout(n21896));
  jor  g04634(.dina(n21896), .dinb(n21800), .dout(n21897));
  jxor g04635(.dina(n21794), .dinb(n360), .dout(n21898));
  jand g04636(.dina(n21898), .dinb(n21897), .dout(n21899));
  jor  g04637(.dina(n21899), .dinb(n21795), .dout(n21900));
  jxor g04638(.dina(n21789), .dinb(n361), .dout(n21901));
  jand g04639(.dina(n21901), .dinb(n21900), .dout(n21902));
  jor  g04640(.dina(n21902), .dinb(n21790), .dout(n21903));
  jxor g04641(.dina(n21784), .dinb(n364), .dout(n21904));
  jand g04642(.dina(n21904), .dinb(n21903), .dout(n21905));
  jor  g04643(.dina(n21905), .dinb(n21785), .dout(n21906));
  jxor g04644(.dina(n21779), .dinb(n355), .dout(n21907));
  jand g04645(.dina(n21907), .dinb(n21906), .dout(n21908));
  jor  g04646(.dina(n21908), .dinb(n21780), .dout(n21909));
  jxor g04647(.dina(n21774), .dinb(n356), .dout(n21910));
  jand g04648(.dina(n21910), .dinb(n21909), .dout(n21911));
  jor  g04649(.dina(n21911), .dinb(n21775), .dout(n21912));
  jxor g04650(.dina(n21769), .dinb(n266), .dout(n21913));
  jand g04651(.dina(n21913), .dinb(n21912), .dout(n21914));
  jor  g04652(.dina(n21914), .dinb(n21770), .dout(n21915));
  jxor g04653(.dina(n21764), .dinb(n267), .dout(n21916));
  jand g04654(.dina(n21916), .dinb(n21915), .dout(n21917));
  jor  g04655(.dina(n21917), .dinb(n21765), .dout(n21918));
  jxor g04656(.dina(n21759), .dinb(n347), .dout(n21919));
  jand g04657(.dina(n21919), .dinb(n21918), .dout(n21920));
  jor  g04658(.dina(n21920), .dinb(n21760), .dout(n21921));
  jxor g04659(.dina(n21754), .dinb(n348), .dout(n21922));
  jand g04660(.dina(n21922), .dinb(n21921), .dout(n21923));
  jor  g04661(.dina(n21923), .dinb(n21755), .dout(n21924));
  jxor g04662(.dina(n21749), .dinb(n349), .dout(n21925));
  jand g04663(.dina(n21925), .dinb(n21924), .dout(n21926));
  jor  g04664(.dina(n21926), .dinb(n21750), .dout(n21927));
  jxor g04665(.dina(n21744), .dinb(n268), .dout(n21928));
  jand g04666(.dina(n21928), .dinb(n21927), .dout(n21929));
  jor  g04667(.dina(n21929), .dinb(n21745), .dout(n21930));
  jxor g04668(.dina(n21739), .dinb(n274), .dout(n21931));
  jand g04669(.dina(n21931), .dinb(n21930), .dout(n21932));
  jor  g04670(.dina(n21932), .dinb(n21740), .dout(n21933));
  jxor g04671(.dina(n21734), .dinb(n269), .dout(n21934));
  jand g04672(.dina(n21934), .dinb(n21933), .dout(n21935));
  jor  g04673(.dina(n21935), .dinb(n21735), .dout(n21936));
  jand g04674(.dina(n21628), .dinb(n415), .dout(n21937));
  jor  g04675(.dina(n21937), .dinb(n21731), .dout(n21938));
  jand g04676(.dina(n21938), .dinb(n21332), .dout(n21939));
  jxor g04677(.dina(n21939), .dinb(n270), .dout(n21940));
  jand g04678(.dina(n21940), .dinb(n21936), .dout(n21941));
  jand g04679(.dina(n21941), .dinb(n3678), .dout(n21942));
  jand g04680(.dina(n21939), .dinb(n3157), .dout(n21943));
  jor  g04681(.dina(n21943), .dinb(n21942), .dout(n21944));
  jor  g04682(.dina(n21944), .dinb(n21734), .dout(n21945));
  jnot g04683(.din(n21944), .dout(n21946));
  jxor g04684(.dina(n21934), .dinb(n21933), .dout(n21947));
  jor  g04685(.dina(n21947), .dinb(n21946), .dout(n21948));
  jand g04686(.dina(n21948), .dinb(n21945), .dout(n21949));
  jxor g04687(.dina(n21940), .dinb(n21936), .dout(n21950));
  jor  g04688(.dina(n21950), .dinb(n21946), .dout(n21951));
  jor  g04689(.dina(n21942), .dinb(n21939), .dout(n21952));
  jand g04690(.dina(n21952), .dinb(n21951), .dout(n21953));
  jand g04691(.dina(n21953), .dinb(n271), .dout(n21954));
  jnot g04692(.din(n21953), .dout(n21955));
  jand g04693(.dina(n21955), .dinb(b27 ), .dout(n21956));
  jnot g04694(.din(n21956), .dout(n21957));
  jand g04695(.dina(n21949), .dinb(n270), .dout(n21958));
  jor  g04696(.dina(n21944), .dinb(n21739), .dout(n21959));
  jxor g04697(.dina(n21931), .dinb(n21930), .dout(n21960));
  jor  g04698(.dina(n21960), .dinb(n21946), .dout(n21961));
  jand g04699(.dina(n21961), .dinb(n21959), .dout(n21962));
  jand g04700(.dina(n21962), .dinb(n269), .dout(n21963));
  jor  g04701(.dina(n21944), .dinb(n21744), .dout(n21964));
  jxor g04702(.dina(n21928), .dinb(n21927), .dout(n21965));
  jor  g04703(.dina(n21965), .dinb(n21946), .dout(n21966));
  jand g04704(.dina(n21966), .dinb(n21964), .dout(n21967));
  jand g04705(.dina(n21967), .dinb(n274), .dout(n21968));
  jor  g04706(.dina(n21944), .dinb(n21749), .dout(n21969));
  jxor g04707(.dina(n21925), .dinb(n21924), .dout(n21970));
  jor  g04708(.dina(n21970), .dinb(n21946), .dout(n21971));
  jand g04709(.dina(n21971), .dinb(n21969), .dout(n21972));
  jand g04710(.dina(n21972), .dinb(n268), .dout(n21973));
  jor  g04711(.dina(n21944), .dinb(n21754), .dout(n21974));
  jxor g04712(.dina(n21922), .dinb(n21921), .dout(n21975));
  jor  g04713(.dina(n21975), .dinb(n21946), .dout(n21976));
  jand g04714(.dina(n21976), .dinb(n21974), .dout(n21977));
  jand g04715(.dina(n21977), .dinb(n349), .dout(n21978));
  jor  g04716(.dina(n21944), .dinb(n21759), .dout(n21979));
  jxor g04717(.dina(n21919), .dinb(n21918), .dout(n21980));
  jor  g04718(.dina(n21980), .dinb(n21946), .dout(n21981));
  jand g04719(.dina(n21981), .dinb(n21979), .dout(n21982));
  jand g04720(.dina(n21982), .dinb(n348), .dout(n21983));
  jor  g04721(.dina(n21944), .dinb(n21764), .dout(n21984));
  jxor g04722(.dina(n21916), .dinb(n21915), .dout(n21985));
  jor  g04723(.dina(n21985), .dinb(n21946), .dout(n21986));
  jand g04724(.dina(n21986), .dinb(n21984), .dout(n21987));
  jand g04725(.dina(n21987), .dinb(n347), .dout(n21988));
  jor  g04726(.dina(n21944), .dinb(n21769), .dout(n21989));
  jxor g04727(.dina(n21913), .dinb(n21912), .dout(n21990));
  jor  g04728(.dina(n21990), .dinb(n21946), .dout(n21991));
  jand g04729(.dina(n21991), .dinb(n21989), .dout(n21992));
  jand g04730(.dina(n21992), .dinb(n267), .dout(n21993));
  jor  g04731(.dina(n21944), .dinb(n21774), .dout(n21994));
  jxor g04732(.dina(n21910), .dinb(n21909), .dout(n21995));
  jor  g04733(.dina(n21995), .dinb(n21946), .dout(n21996));
  jand g04734(.dina(n21996), .dinb(n21994), .dout(n21997));
  jand g04735(.dina(n21997), .dinb(n266), .dout(n21998));
  jor  g04736(.dina(n21944), .dinb(n21779), .dout(n21999));
  jxor g04737(.dina(n21907), .dinb(n21906), .dout(n22000));
  jor  g04738(.dina(n22000), .dinb(n21946), .dout(n22001));
  jand g04739(.dina(n22001), .dinb(n21999), .dout(n22002));
  jand g04740(.dina(n22002), .dinb(n356), .dout(n22003));
  jor  g04741(.dina(n21944), .dinb(n21784), .dout(n22004));
  jxor g04742(.dina(n21904), .dinb(n21903), .dout(n22005));
  jor  g04743(.dina(n22005), .dinb(n21946), .dout(n22006));
  jand g04744(.dina(n22006), .dinb(n22004), .dout(n22007));
  jand g04745(.dina(n22007), .dinb(n355), .dout(n22008));
  jor  g04746(.dina(n21944), .dinb(n21789), .dout(n22009));
  jxor g04747(.dina(n21901), .dinb(n21900), .dout(n22010));
  jor  g04748(.dina(n22010), .dinb(n21946), .dout(n22011));
  jand g04749(.dina(n22011), .dinb(n22009), .dout(n22012));
  jand g04750(.dina(n22012), .dinb(n364), .dout(n22013));
  jor  g04751(.dina(n21944), .dinb(n21794), .dout(n22014));
  jxor g04752(.dina(n21898), .dinb(n21897), .dout(n22015));
  jor  g04753(.dina(n22015), .dinb(n21946), .dout(n22016));
  jand g04754(.dina(n22016), .dinb(n22014), .dout(n22017));
  jand g04755(.dina(n22017), .dinb(n361), .dout(n22018));
  jor  g04756(.dina(n21944), .dinb(n21799), .dout(n22019));
  jxor g04757(.dina(n21895), .dinb(n21894), .dout(n22020));
  jor  g04758(.dina(n22020), .dinb(n21946), .dout(n22021));
  jand g04759(.dina(n22021), .dinb(n22019), .dout(n22022));
  jand g04760(.dina(n22022), .dinb(n360), .dout(n22023));
  jor  g04761(.dina(n21944), .dinb(n21804), .dout(n22024));
  jxor g04762(.dina(n21892), .dinb(n21891), .dout(n22025));
  jor  g04763(.dina(n22025), .dinb(n21946), .dout(n22026));
  jand g04764(.dina(n22026), .dinb(n22024), .dout(n22027));
  jand g04765(.dina(n22027), .dinb(n363), .dout(n22028));
  jor  g04766(.dina(n21944), .dinb(n21809), .dout(n22029));
  jxor g04767(.dina(n21889), .dinb(n21888), .dout(n22030));
  jor  g04768(.dina(n22030), .dinb(n21946), .dout(n22031));
  jand g04769(.dina(n22031), .dinb(n22029), .dout(n22032));
  jand g04770(.dina(n22032), .dinb(n359), .dout(n22033));
  jor  g04771(.dina(n21944), .dinb(n21814), .dout(n22034));
  jxor g04772(.dina(n21886), .dinb(n21885), .dout(n22035));
  jor  g04773(.dina(n22035), .dinb(n21946), .dout(n22036));
  jand g04774(.dina(n22036), .dinb(n22034), .dout(n22037));
  jand g04775(.dina(n22037), .dinb(n369), .dout(n22038));
  jor  g04776(.dina(n21944), .dinb(n21819), .dout(n22039));
  jxor g04777(.dina(n21883), .dinb(n21882), .dout(n22040));
  jor  g04778(.dina(n22040), .dinb(n21946), .dout(n22041));
  jand g04779(.dina(n22041), .dinb(n22039), .dout(n22042));
  jand g04780(.dina(n22042), .dinb(n368), .dout(n22043));
  jor  g04781(.dina(n21944), .dinb(n21824), .dout(n22044));
  jxor g04782(.dina(n21880), .dinb(n21879), .dout(n22045));
  jor  g04783(.dina(n22045), .dinb(n21946), .dout(n22046));
  jand g04784(.dina(n22046), .dinb(n22044), .dout(n22047));
  jand g04785(.dina(n22047), .dinb(n367), .dout(n22048));
  jor  g04786(.dina(n21944), .dinb(n21829), .dout(n22049));
  jxor g04787(.dina(n21877), .dinb(n21876), .dout(n22050));
  jor  g04788(.dina(n22050), .dinb(n21946), .dout(n22051));
  jand g04789(.dina(n22051), .dinb(n22049), .dout(n22052));
  jand g04790(.dina(n22052), .dinb(n265), .dout(n22053));
  jor  g04791(.dina(n21944), .dinb(n21834), .dout(n22054));
  jxor g04792(.dina(n21874), .dinb(n21873), .dout(n22055));
  jor  g04793(.dina(n22055), .dinb(n21946), .dout(n22056));
  jand g04794(.dina(n22056), .dinb(n22054), .dout(n22057));
  jand g04795(.dina(n22057), .dinb(n378), .dout(n22058));
  jor  g04796(.dina(n21944), .dinb(n21839), .dout(n22059));
  jxor g04797(.dina(n21871), .dinb(n21870), .dout(n22060));
  jor  g04798(.dina(n22060), .dinb(n21946), .dout(n22061));
  jand g04799(.dina(n22061), .dinb(n22059), .dout(n22062));
  jand g04800(.dina(n22062), .dinb(n377), .dout(n22063));
  jor  g04801(.dina(n21944), .dinb(n21845), .dout(n22064));
  jxor g04802(.dina(n21868), .dinb(n21867), .dout(n22065));
  jor  g04803(.dina(n22065), .dinb(n21946), .dout(n22066));
  jand g04804(.dina(n22066), .dinb(n22064), .dout(n22067));
  jand g04805(.dina(n22067), .dinb(n376), .dout(n22068));
  jxor g04806(.dina(n21865), .dinb(n21864), .dout(n22069));
  jnot g04807(.din(n22069), .dout(n22070));
  jor  g04808(.dina(n22070), .dinb(n21946), .dout(n22071));
  jnot g04809(.din(n21850), .dout(n22072));
  jor  g04810(.dina(n21944), .dinb(n22072), .dout(n22073));
  jand g04811(.dina(n22073), .dinb(n22071), .dout(n22074));
  jnot g04812(.din(n22074), .dout(n22075));
  jand g04813(.dina(n22075), .dinb(n264), .dout(n22076));
  jor  g04814(.dina(n21944), .dinb(n21861), .dout(n22077));
  jxor g04815(.dina(n21862), .dinb(n3602), .dout(n22078));
  jand g04816(.dina(n22078), .dinb(n21944), .dout(n22079));
  jnot g04817(.din(n22079), .dout(n22080));
  jand g04818(.dina(n22080), .dinb(n22077), .dout(n22081));
  jnot g04819(.din(n22081), .dout(n22082));
  jand g04820(.dina(n22082), .dinb(n386), .dout(n22083));
  jand g04821(.dina(n21944), .dinb(b0 ), .dout(n22084));
  jxor g04822(.dina(n22084), .dinb(a37 ), .dout(n22085));
  jand g04823(.dina(n22085), .dinb(n259), .dout(n22086));
  jxor g04824(.dina(n22084), .dinb(n3600), .dout(n22087));
  jxor g04825(.dina(n22087), .dinb(b1 ), .dout(n22088));
  jand g04826(.dina(n22088), .dinb(n3824), .dout(n22089));
  jor  g04827(.dina(n22089), .dinb(n22086), .dout(n22090));
  jxor g04828(.dina(n22081), .dinb(b2 ), .dout(n22091));
  jand g04829(.dina(n22091), .dinb(n22090), .dout(n22092));
  jor  g04830(.dina(n22092), .dinb(n22083), .dout(n22093));
  jxor g04831(.dina(n22074), .dinb(b3 ), .dout(n22094));
  jand g04832(.dina(n22094), .dinb(n22093), .dout(n22095));
  jor  g04833(.dina(n22095), .dinb(n22076), .dout(n22096));
  jxor g04834(.dina(n22067), .dinb(n376), .dout(n22097));
  jand g04835(.dina(n22097), .dinb(n22096), .dout(n22098));
  jor  g04836(.dina(n22098), .dinb(n22068), .dout(n22099));
  jxor g04837(.dina(n22062), .dinb(n377), .dout(n22100));
  jand g04838(.dina(n22100), .dinb(n22099), .dout(n22101));
  jor  g04839(.dina(n22101), .dinb(n22063), .dout(n22102));
  jxor g04840(.dina(n22057), .dinb(n378), .dout(n22103));
  jand g04841(.dina(n22103), .dinb(n22102), .dout(n22104));
  jor  g04842(.dina(n22104), .dinb(n22058), .dout(n22105));
  jxor g04843(.dina(n22052), .dinb(n265), .dout(n22106));
  jand g04844(.dina(n22106), .dinb(n22105), .dout(n22107));
  jor  g04845(.dina(n22107), .dinb(n22053), .dout(n22108));
  jxor g04846(.dina(n22047), .dinb(n367), .dout(n22109));
  jand g04847(.dina(n22109), .dinb(n22108), .dout(n22110));
  jor  g04848(.dina(n22110), .dinb(n22048), .dout(n22111));
  jxor g04849(.dina(n22042), .dinb(n368), .dout(n22112));
  jand g04850(.dina(n22112), .dinb(n22111), .dout(n22113));
  jor  g04851(.dina(n22113), .dinb(n22043), .dout(n22114));
  jxor g04852(.dina(n22037), .dinb(n369), .dout(n22115));
  jand g04853(.dina(n22115), .dinb(n22114), .dout(n22116));
  jor  g04854(.dina(n22116), .dinb(n22038), .dout(n22117));
  jxor g04855(.dina(n22032), .dinb(n359), .dout(n22118));
  jand g04856(.dina(n22118), .dinb(n22117), .dout(n22119));
  jor  g04857(.dina(n22119), .dinb(n22033), .dout(n22120));
  jxor g04858(.dina(n22027), .dinb(n363), .dout(n22121));
  jand g04859(.dina(n22121), .dinb(n22120), .dout(n22122));
  jor  g04860(.dina(n22122), .dinb(n22028), .dout(n22123));
  jxor g04861(.dina(n22022), .dinb(n360), .dout(n22124));
  jand g04862(.dina(n22124), .dinb(n22123), .dout(n22125));
  jor  g04863(.dina(n22125), .dinb(n22023), .dout(n22126));
  jxor g04864(.dina(n22017), .dinb(n361), .dout(n22127));
  jand g04865(.dina(n22127), .dinb(n22126), .dout(n22128));
  jor  g04866(.dina(n22128), .dinb(n22018), .dout(n22129));
  jxor g04867(.dina(n22012), .dinb(n364), .dout(n22130));
  jand g04868(.dina(n22130), .dinb(n22129), .dout(n22131));
  jor  g04869(.dina(n22131), .dinb(n22013), .dout(n22132));
  jxor g04870(.dina(n22007), .dinb(n355), .dout(n22133));
  jand g04871(.dina(n22133), .dinb(n22132), .dout(n22134));
  jor  g04872(.dina(n22134), .dinb(n22008), .dout(n22135));
  jxor g04873(.dina(n22002), .dinb(n356), .dout(n22136));
  jand g04874(.dina(n22136), .dinb(n22135), .dout(n22137));
  jor  g04875(.dina(n22137), .dinb(n22003), .dout(n22138));
  jxor g04876(.dina(n21997), .dinb(n266), .dout(n22139));
  jand g04877(.dina(n22139), .dinb(n22138), .dout(n22140));
  jor  g04878(.dina(n22140), .dinb(n21998), .dout(n22141));
  jxor g04879(.dina(n21992), .dinb(n267), .dout(n22142));
  jand g04880(.dina(n22142), .dinb(n22141), .dout(n22143));
  jor  g04881(.dina(n22143), .dinb(n21993), .dout(n22144));
  jxor g04882(.dina(n21987), .dinb(n347), .dout(n22145));
  jand g04883(.dina(n22145), .dinb(n22144), .dout(n22146));
  jor  g04884(.dina(n22146), .dinb(n21988), .dout(n22147));
  jxor g04885(.dina(n21982), .dinb(n348), .dout(n22148));
  jand g04886(.dina(n22148), .dinb(n22147), .dout(n22149));
  jor  g04887(.dina(n22149), .dinb(n21983), .dout(n22150));
  jxor g04888(.dina(n21977), .dinb(n349), .dout(n22151));
  jand g04889(.dina(n22151), .dinb(n22150), .dout(n22152));
  jor  g04890(.dina(n22152), .dinb(n21978), .dout(n22153));
  jxor g04891(.dina(n21972), .dinb(n268), .dout(n22154));
  jand g04892(.dina(n22154), .dinb(n22153), .dout(n22155));
  jor  g04893(.dina(n22155), .dinb(n21973), .dout(n22156));
  jxor g04894(.dina(n21967), .dinb(n274), .dout(n22157));
  jand g04895(.dina(n22157), .dinb(n22156), .dout(n22158));
  jor  g04896(.dina(n22158), .dinb(n21968), .dout(n22159));
  jxor g04897(.dina(n21962), .dinb(n269), .dout(n22160));
  jand g04898(.dina(n22160), .dinb(n22159), .dout(n22161));
  jor  g04899(.dina(n22161), .dinb(n21963), .dout(n22162));
  jxor g04900(.dina(n21949), .dinb(n270), .dout(n22163));
  jand g04901(.dina(n22163), .dinb(n22162), .dout(n22164));
  jor  g04902(.dina(n22164), .dinb(n21958), .dout(n22165));
  jand g04903(.dina(n22165), .dinb(n21957), .dout(n22166));
  jor  g04904(.dina(n22166), .dinb(n21954), .dout(n22167));
  jand g04905(.dina(n22167), .dinb(n414), .dout(n22168));
  jor  g04906(.dina(n22168), .dinb(n21949), .dout(n22169));
  jnot g04907(.din(n22168), .dout(n22170));
  jxor g04908(.dina(n22163), .dinb(n22162), .dout(n22171));
  jor  g04909(.dina(n22171), .dinb(n22170), .dout(n22172));
  jand g04910(.dina(n22172), .dinb(n22169), .dout(n22173));
  jand g04911(.dina(n22170), .dinb(n21953), .dout(n22174));
  jand g04912(.dina(n22165), .dinb(n21954), .dout(n22175));
  jor  g04913(.dina(n22175), .dinb(n22174), .dout(n22176));
  jand g04914(.dina(n22176), .dinb(n338), .dout(n22177));
  jnot g04915(.din(n22176), .dout(n22178));
  jand g04916(.dina(n22178), .dinb(b28 ), .dout(n22179));
  jnot g04917(.din(n22179), .dout(n22180));
  jand g04918(.dina(n22173), .dinb(n271), .dout(n22181));
  jor  g04919(.dina(n22168), .dinb(n21962), .dout(n22182));
  jxor g04920(.dina(n22160), .dinb(n22159), .dout(n22183));
  jor  g04921(.dina(n22183), .dinb(n22170), .dout(n22184));
  jand g04922(.dina(n22184), .dinb(n22182), .dout(n22185));
  jand g04923(.dina(n22185), .dinb(n270), .dout(n22186));
  jor  g04924(.dina(n22168), .dinb(n21967), .dout(n22187));
  jxor g04925(.dina(n22157), .dinb(n22156), .dout(n22188));
  jor  g04926(.dina(n22188), .dinb(n22170), .dout(n22189));
  jand g04927(.dina(n22189), .dinb(n22187), .dout(n22190));
  jand g04928(.dina(n22190), .dinb(n269), .dout(n22191));
  jor  g04929(.dina(n22168), .dinb(n21972), .dout(n22192));
  jxor g04930(.dina(n22154), .dinb(n22153), .dout(n22193));
  jor  g04931(.dina(n22193), .dinb(n22170), .dout(n22194));
  jand g04932(.dina(n22194), .dinb(n22192), .dout(n22195));
  jand g04933(.dina(n22195), .dinb(n274), .dout(n22196));
  jor  g04934(.dina(n22168), .dinb(n21977), .dout(n22197));
  jxor g04935(.dina(n22151), .dinb(n22150), .dout(n22198));
  jor  g04936(.dina(n22198), .dinb(n22170), .dout(n22199));
  jand g04937(.dina(n22199), .dinb(n22197), .dout(n22200));
  jand g04938(.dina(n22200), .dinb(n268), .dout(n22201));
  jor  g04939(.dina(n22168), .dinb(n21982), .dout(n22202));
  jxor g04940(.dina(n22148), .dinb(n22147), .dout(n22203));
  jor  g04941(.dina(n22203), .dinb(n22170), .dout(n22204));
  jand g04942(.dina(n22204), .dinb(n22202), .dout(n22205));
  jand g04943(.dina(n22205), .dinb(n349), .dout(n22206));
  jor  g04944(.dina(n22168), .dinb(n21987), .dout(n22207));
  jxor g04945(.dina(n22145), .dinb(n22144), .dout(n22208));
  jor  g04946(.dina(n22208), .dinb(n22170), .dout(n22209));
  jand g04947(.dina(n22209), .dinb(n22207), .dout(n22210));
  jand g04948(.dina(n22210), .dinb(n348), .dout(n22211));
  jor  g04949(.dina(n22168), .dinb(n21992), .dout(n22212));
  jxor g04950(.dina(n22142), .dinb(n22141), .dout(n22213));
  jor  g04951(.dina(n22213), .dinb(n22170), .dout(n22214));
  jand g04952(.dina(n22214), .dinb(n22212), .dout(n22215));
  jand g04953(.dina(n22215), .dinb(n347), .dout(n22216));
  jor  g04954(.dina(n22168), .dinb(n21997), .dout(n22217));
  jxor g04955(.dina(n22139), .dinb(n22138), .dout(n22218));
  jor  g04956(.dina(n22218), .dinb(n22170), .dout(n22219));
  jand g04957(.dina(n22219), .dinb(n22217), .dout(n22220));
  jand g04958(.dina(n22220), .dinb(n267), .dout(n22221));
  jor  g04959(.dina(n22168), .dinb(n22002), .dout(n22222));
  jxor g04960(.dina(n22136), .dinb(n22135), .dout(n22223));
  jor  g04961(.dina(n22223), .dinb(n22170), .dout(n22224));
  jand g04962(.dina(n22224), .dinb(n22222), .dout(n22225));
  jand g04963(.dina(n22225), .dinb(n266), .dout(n22226));
  jor  g04964(.dina(n22168), .dinb(n22007), .dout(n22227));
  jxor g04965(.dina(n22133), .dinb(n22132), .dout(n22228));
  jor  g04966(.dina(n22228), .dinb(n22170), .dout(n22229));
  jand g04967(.dina(n22229), .dinb(n22227), .dout(n22230));
  jand g04968(.dina(n22230), .dinb(n356), .dout(n22231));
  jor  g04969(.dina(n22168), .dinb(n22012), .dout(n22232));
  jxor g04970(.dina(n22130), .dinb(n22129), .dout(n22233));
  jor  g04971(.dina(n22233), .dinb(n22170), .dout(n22234));
  jand g04972(.dina(n22234), .dinb(n22232), .dout(n22235));
  jand g04973(.dina(n22235), .dinb(n355), .dout(n22236));
  jor  g04974(.dina(n22168), .dinb(n22017), .dout(n22237));
  jxor g04975(.dina(n22127), .dinb(n22126), .dout(n22238));
  jor  g04976(.dina(n22238), .dinb(n22170), .dout(n22239));
  jand g04977(.dina(n22239), .dinb(n22237), .dout(n22240));
  jand g04978(.dina(n22240), .dinb(n364), .dout(n22241));
  jor  g04979(.dina(n22168), .dinb(n22022), .dout(n22242));
  jxor g04980(.dina(n22124), .dinb(n22123), .dout(n22243));
  jor  g04981(.dina(n22243), .dinb(n22170), .dout(n22244));
  jand g04982(.dina(n22244), .dinb(n22242), .dout(n22245));
  jand g04983(.dina(n22245), .dinb(n361), .dout(n22246));
  jor  g04984(.dina(n22168), .dinb(n22027), .dout(n22247));
  jxor g04985(.dina(n22121), .dinb(n22120), .dout(n22248));
  jor  g04986(.dina(n22248), .dinb(n22170), .dout(n22249));
  jand g04987(.dina(n22249), .dinb(n22247), .dout(n22250));
  jand g04988(.dina(n22250), .dinb(n360), .dout(n22251));
  jor  g04989(.dina(n22168), .dinb(n22032), .dout(n22252));
  jxor g04990(.dina(n22118), .dinb(n22117), .dout(n22253));
  jor  g04991(.dina(n22253), .dinb(n22170), .dout(n22254));
  jand g04992(.dina(n22254), .dinb(n22252), .dout(n22255));
  jand g04993(.dina(n22255), .dinb(n363), .dout(n22256));
  jor  g04994(.dina(n22168), .dinb(n22037), .dout(n22257));
  jxor g04995(.dina(n22115), .dinb(n22114), .dout(n22258));
  jor  g04996(.dina(n22258), .dinb(n22170), .dout(n22259));
  jand g04997(.dina(n22259), .dinb(n22257), .dout(n22260));
  jand g04998(.dina(n22260), .dinb(n359), .dout(n22261));
  jor  g04999(.dina(n22168), .dinb(n22042), .dout(n22262));
  jxor g05000(.dina(n22112), .dinb(n22111), .dout(n22263));
  jor  g05001(.dina(n22263), .dinb(n22170), .dout(n22264));
  jand g05002(.dina(n22264), .dinb(n22262), .dout(n22265));
  jand g05003(.dina(n22265), .dinb(n369), .dout(n22266));
  jor  g05004(.dina(n22168), .dinb(n22047), .dout(n22267));
  jxor g05005(.dina(n22109), .dinb(n22108), .dout(n22268));
  jor  g05006(.dina(n22268), .dinb(n22170), .dout(n22269));
  jand g05007(.dina(n22269), .dinb(n22267), .dout(n22270));
  jand g05008(.dina(n22270), .dinb(n368), .dout(n22271));
  jor  g05009(.dina(n22168), .dinb(n22052), .dout(n22272));
  jxor g05010(.dina(n22106), .dinb(n22105), .dout(n22273));
  jor  g05011(.dina(n22273), .dinb(n22170), .dout(n22274));
  jand g05012(.dina(n22274), .dinb(n22272), .dout(n22275));
  jand g05013(.dina(n22275), .dinb(n367), .dout(n22276));
  jor  g05014(.dina(n22168), .dinb(n22057), .dout(n22277));
  jxor g05015(.dina(n22103), .dinb(n22102), .dout(n22278));
  jor  g05016(.dina(n22278), .dinb(n22170), .dout(n22279));
  jand g05017(.dina(n22279), .dinb(n22277), .dout(n22280));
  jand g05018(.dina(n22280), .dinb(n265), .dout(n22281));
  jor  g05019(.dina(n22168), .dinb(n22062), .dout(n22282));
  jxor g05020(.dina(n22100), .dinb(n22099), .dout(n22283));
  jor  g05021(.dina(n22283), .dinb(n22170), .dout(n22284));
  jand g05022(.dina(n22284), .dinb(n22282), .dout(n22285));
  jand g05023(.dina(n22285), .dinb(n378), .dout(n22286));
  jor  g05024(.dina(n22168), .dinb(n22067), .dout(n22287));
  jxor g05025(.dina(n22097), .dinb(n22096), .dout(n22288));
  jor  g05026(.dina(n22288), .dinb(n22170), .dout(n22289));
  jand g05027(.dina(n22289), .dinb(n22287), .dout(n22290));
  jand g05028(.dina(n22290), .dinb(n377), .dout(n22291));
  jand g05029(.dina(n22170), .dinb(n22074), .dout(n22292));
  jnot g05030(.din(n22292), .dout(n22293));
  jxor g05031(.dina(n22094), .dinb(n22093), .dout(n22294));
  jor  g05032(.dina(n22294), .dinb(n22170), .dout(n22295));
  jand g05033(.dina(n22295), .dinb(n22293), .dout(n22296));
  jand g05034(.dina(n22296), .dinb(n376), .dout(n22297));
  jor  g05035(.dina(n22168), .dinb(n22082), .dout(n22298));
  jxor g05036(.dina(n22091), .dinb(n22090), .dout(n22299));
  jor  g05037(.dina(n22299), .dinb(n22170), .dout(n22300));
  jand g05038(.dina(n22300), .dinb(n22298), .dout(n22301));
  jand g05039(.dina(n22301), .dinb(n264), .dout(n22302));
  jor  g05040(.dina(n22168), .dinb(n22085), .dout(n22303));
  jxor g05041(.dina(n22088), .dinb(n3824), .dout(n22304));
  jor  g05042(.dina(n22304), .dinb(n22170), .dout(n22305));
  jand g05043(.dina(n22305), .dinb(n22303), .dout(n22306));
  jand g05044(.dina(n22306), .dinb(n386), .dout(n22307));
  jnot g05045(.din(n3592), .dout(n22308));
  jnot g05046(.din(n21954), .dout(n22309));
  jnot g05047(.din(n21958), .dout(n22310));
  jnot g05048(.din(n21963), .dout(n22311));
  jnot g05049(.din(n21968), .dout(n22312));
  jnot g05050(.din(n21973), .dout(n22313));
  jnot g05051(.din(n21978), .dout(n22314));
  jnot g05052(.din(n21983), .dout(n22315));
  jnot g05053(.din(n21988), .dout(n22316));
  jnot g05054(.din(n21993), .dout(n22317));
  jnot g05055(.din(n21998), .dout(n22318));
  jnot g05056(.din(n22003), .dout(n22319));
  jnot g05057(.din(n22008), .dout(n22320));
  jnot g05058(.din(n22013), .dout(n22321));
  jnot g05059(.din(n22018), .dout(n22322));
  jnot g05060(.din(n22023), .dout(n22323));
  jnot g05061(.din(n22028), .dout(n22324));
  jnot g05062(.din(n22033), .dout(n22325));
  jnot g05063(.din(n22038), .dout(n22326));
  jnot g05064(.din(n22043), .dout(n22327));
  jnot g05065(.din(n22048), .dout(n22328));
  jnot g05066(.din(n22053), .dout(n22329));
  jnot g05067(.din(n22058), .dout(n22330));
  jnot g05068(.din(n22063), .dout(n22331));
  jnot g05069(.din(n22068), .dout(n22332));
  jnot g05070(.din(n22076), .dout(n22333));
  jnot g05071(.din(n22083), .dout(n22334));
  jnot g05072(.din(n22086), .dout(n22335));
  jxor g05073(.dina(n22087), .dinb(n259), .dout(n22336));
  jor  g05074(.dina(n22336), .dinb(n3823), .dout(n22337));
  jand g05075(.dina(n22337), .dinb(n22335), .dout(n22338));
  jnot g05076(.din(n22091), .dout(n22339));
  jor  g05077(.dina(n22339), .dinb(n22338), .dout(n22340));
  jand g05078(.dina(n22340), .dinb(n22334), .dout(n22341));
  jnot g05079(.din(n22094), .dout(n22342));
  jor  g05080(.dina(n22342), .dinb(n22341), .dout(n22343));
  jand g05081(.dina(n22343), .dinb(n22333), .dout(n22344));
  jnot g05082(.din(n22097), .dout(n22345));
  jor  g05083(.dina(n22345), .dinb(n22344), .dout(n22346));
  jand g05084(.dina(n22346), .dinb(n22332), .dout(n22347));
  jnot g05085(.din(n22100), .dout(n22348));
  jor  g05086(.dina(n22348), .dinb(n22347), .dout(n22349));
  jand g05087(.dina(n22349), .dinb(n22331), .dout(n22350));
  jnot g05088(.din(n22103), .dout(n22351));
  jor  g05089(.dina(n22351), .dinb(n22350), .dout(n22352));
  jand g05090(.dina(n22352), .dinb(n22330), .dout(n22353));
  jnot g05091(.din(n22106), .dout(n22354));
  jor  g05092(.dina(n22354), .dinb(n22353), .dout(n22355));
  jand g05093(.dina(n22355), .dinb(n22329), .dout(n22356));
  jnot g05094(.din(n22109), .dout(n22357));
  jor  g05095(.dina(n22357), .dinb(n22356), .dout(n22358));
  jand g05096(.dina(n22358), .dinb(n22328), .dout(n22359));
  jnot g05097(.din(n22112), .dout(n22360));
  jor  g05098(.dina(n22360), .dinb(n22359), .dout(n22361));
  jand g05099(.dina(n22361), .dinb(n22327), .dout(n22362));
  jnot g05100(.din(n22115), .dout(n22363));
  jor  g05101(.dina(n22363), .dinb(n22362), .dout(n22364));
  jand g05102(.dina(n22364), .dinb(n22326), .dout(n22365));
  jnot g05103(.din(n22118), .dout(n22366));
  jor  g05104(.dina(n22366), .dinb(n22365), .dout(n22367));
  jand g05105(.dina(n22367), .dinb(n22325), .dout(n22368));
  jnot g05106(.din(n22121), .dout(n22369));
  jor  g05107(.dina(n22369), .dinb(n22368), .dout(n22370));
  jand g05108(.dina(n22370), .dinb(n22324), .dout(n22371));
  jnot g05109(.din(n22124), .dout(n22372));
  jor  g05110(.dina(n22372), .dinb(n22371), .dout(n22373));
  jand g05111(.dina(n22373), .dinb(n22323), .dout(n22374));
  jnot g05112(.din(n22127), .dout(n22375));
  jor  g05113(.dina(n22375), .dinb(n22374), .dout(n22376));
  jand g05114(.dina(n22376), .dinb(n22322), .dout(n22377));
  jnot g05115(.din(n22130), .dout(n22378));
  jor  g05116(.dina(n22378), .dinb(n22377), .dout(n22379));
  jand g05117(.dina(n22379), .dinb(n22321), .dout(n22380));
  jnot g05118(.din(n22133), .dout(n22381));
  jor  g05119(.dina(n22381), .dinb(n22380), .dout(n22382));
  jand g05120(.dina(n22382), .dinb(n22320), .dout(n22383));
  jnot g05121(.din(n22136), .dout(n22384));
  jor  g05122(.dina(n22384), .dinb(n22383), .dout(n22385));
  jand g05123(.dina(n22385), .dinb(n22319), .dout(n22386));
  jnot g05124(.din(n22139), .dout(n22387));
  jor  g05125(.dina(n22387), .dinb(n22386), .dout(n22388));
  jand g05126(.dina(n22388), .dinb(n22318), .dout(n22389));
  jnot g05127(.din(n22142), .dout(n22390));
  jor  g05128(.dina(n22390), .dinb(n22389), .dout(n22391));
  jand g05129(.dina(n22391), .dinb(n22317), .dout(n22392));
  jnot g05130(.din(n22145), .dout(n22393));
  jor  g05131(.dina(n22393), .dinb(n22392), .dout(n22394));
  jand g05132(.dina(n22394), .dinb(n22316), .dout(n22395));
  jnot g05133(.din(n22148), .dout(n22396));
  jor  g05134(.dina(n22396), .dinb(n22395), .dout(n22397));
  jand g05135(.dina(n22397), .dinb(n22315), .dout(n22398));
  jnot g05136(.din(n22151), .dout(n22399));
  jor  g05137(.dina(n22399), .dinb(n22398), .dout(n22400));
  jand g05138(.dina(n22400), .dinb(n22314), .dout(n22401));
  jnot g05139(.din(n22154), .dout(n22402));
  jor  g05140(.dina(n22402), .dinb(n22401), .dout(n22403));
  jand g05141(.dina(n22403), .dinb(n22313), .dout(n22404));
  jnot g05142(.din(n22157), .dout(n22405));
  jor  g05143(.dina(n22405), .dinb(n22404), .dout(n22406));
  jand g05144(.dina(n22406), .dinb(n22312), .dout(n22407));
  jnot g05145(.din(n22160), .dout(n22408));
  jor  g05146(.dina(n22408), .dinb(n22407), .dout(n22409));
  jand g05147(.dina(n22409), .dinb(n22311), .dout(n22410));
  jnot g05148(.din(n22163), .dout(n22411));
  jor  g05149(.dina(n22411), .dinb(n22410), .dout(n22412));
  jand g05150(.dina(n22412), .dinb(n22310), .dout(n22413));
  jor  g05151(.dina(n22413), .dinb(n21956), .dout(n22414));
  jand g05152(.dina(n22414), .dinb(n22309), .dout(n22415));
  jor  g05153(.dina(n22415), .dinb(n22308), .dout(n22416));
  jand g05154(.dina(n22416), .dinb(a36 ), .dout(n22417));
  jnot g05155(.din(n4047), .dout(n22418));
  jor  g05156(.dina(n22415), .dinb(n22418), .dout(n22419));
  jnot g05157(.din(n22419), .dout(n22420));
  jor  g05158(.dina(n22420), .dinb(n22417), .dout(n22421));
  jand g05159(.dina(n22421), .dinb(n259), .dout(n22422));
  jand g05160(.dina(n22167), .dinb(n3592), .dout(n22423));
  jor  g05161(.dina(n22423), .dinb(n3822), .dout(n22424));
  jand g05162(.dina(n22419), .dinb(n22424), .dout(n22425));
  jxor g05163(.dina(n22425), .dinb(b1 ), .dout(n22426));
  jand g05164(.dina(n22426), .dinb(n4055), .dout(n22427));
  jor  g05165(.dina(n22427), .dinb(n22422), .dout(n22428));
  jxor g05166(.dina(n22306), .dinb(n386), .dout(n22429));
  jand g05167(.dina(n22429), .dinb(n22428), .dout(n22430));
  jor  g05168(.dina(n22430), .dinb(n22307), .dout(n22431));
  jxor g05169(.dina(n22301), .dinb(n264), .dout(n22432));
  jand g05170(.dina(n22432), .dinb(n22431), .dout(n22433));
  jor  g05171(.dina(n22433), .dinb(n22302), .dout(n22434));
  jxor g05172(.dina(n22296), .dinb(n376), .dout(n22435));
  jand g05173(.dina(n22435), .dinb(n22434), .dout(n22436));
  jor  g05174(.dina(n22436), .dinb(n22297), .dout(n22437));
  jxor g05175(.dina(n22290), .dinb(n377), .dout(n22438));
  jand g05176(.dina(n22438), .dinb(n22437), .dout(n22439));
  jor  g05177(.dina(n22439), .dinb(n22291), .dout(n22440));
  jxor g05178(.dina(n22285), .dinb(n378), .dout(n22441));
  jand g05179(.dina(n22441), .dinb(n22440), .dout(n22442));
  jor  g05180(.dina(n22442), .dinb(n22286), .dout(n22443));
  jxor g05181(.dina(n22280), .dinb(n265), .dout(n22444));
  jand g05182(.dina(n22444), .dinb(n22443), .dout(n22445));
  jor  g05183(.dina(n22445), .dinb(n22281), .dout(n22446));
  jxor g05184(.dina(n22275), .dinb(n367), .dout(n22447));
  jand g05185(.dina(n22447), .dinb(n22446), .dout(n22448));
  jor  g05186(.dina(n22448), .dinb(n22276), .dout(n22449));
  jxor g05187(.dina(n22270), .dinb(n368), .dout(n22450));
  jand g05188(.dina(n22450), .dinb(n22449), .dout(n22451));
  jor  g05189(.dina(n22451), .dinb(n22271), .dout(n22452));
  jxor g05190(.dina(n22265), .dinb(n369), .dout(n22453));
  jand g05191(.dina(n22453), .dinb(n22452), .dout(n22454));
  jor  g05192(.dina(n22454), .dinb(n22266), .dout(n22455));
  jxor g05193(.dina(n22260), .dinb(n359), .dout(n22456));
  jand g05194(.dina(n22456), .dinb(n22455), .dout(n22457));
  jor  g05195(.dina(n22457), .dinb(n22261), .dout(n22458));
  jxor g05196(.dina(n22255), .dinb(n363), .dout(n22459));
  jand g05197(.dina(n22459), .dinb(n22458), .dout(n22460));
  jor  g05198(.dina(n22460), .dinb(n22256), .dout(n22461));
  jxor g05199(.dina(n22250), .dinb(n360), .dout(n22462));
  jand g05200(.dina(n22462), .dinb(n22461), .dout(n22463));
  jor  g05201(.dina(n22463), .dinb(n22251), .dout(n22464));
  jxor g05202(.dina(n22245), .dinb(n361), .dout(n22465));
  jand g05203(.dina(n22465), .dinb(n22464), .dout(n22466));
  jor  g05204(.dina(n22466), .dinb(n22246), .dout(n22467));
  jxor g05205(.dina(n22240), .dinb(n364), .dout(n22468));
  jand g05206(.dina(n22468), .dinb(n22467), .dout(n22469));
  jor  g05207(.dina(n22469), .dinb(n22241), .dout(n22470));
  jxor g05208(.dina(n22235), .dinb(n355), .dout(n22471));
  jand g05209(.dina(n22471), .dinb(n22470), .dout(n22472));
  jor  g05210(.dina(n22472), .dinb(n22236), .dout(n22473));
  jxor g05211(.dina(n22230), .dinb(n356), .dout(n22474));
  jand g05212(.dina(n22474), .dinb(n22473), .dout(n22475));
  jor  g05213(.dina(n22475), .dinb(n22231), .dout(n22476));
  jxor g05214(.dina(n22225), .dinb(n266), .dout(n22477));
  jand g05215(.dina(n22477), .dinb(n22476), .dout(n22478));
  jor  g05216(.dina(n22478), .dinb(n22226), .dout(n22479));
  jxor g05217(.dina(n22220), .dinb(n267), .dout(n22480));
  jand g05218(.dina(n22480), .dinb(n22479), .dout(n22481));
  jor  g05219(.dina(n22481), .dinb(n22221), .dout(n22482));
  jxor g05220(.dina(n22215), .dinb(n347), .dout(n22483));
  jand g05221(.dina(n22483), .dinb(n22482), .dout(n22484));
  jor  g05222(.dina(n22484), .dinb(n22216), .dout(n22485));
  jxor g05223(.dina(n22210), .dinb(n348), .dout(n22486));
  jand g05224(.dina(n22486), .dinb(n22485), .dout(n22487));
  jor  g05225(.dina(n22487), .dinb(n22211), .dout(n22488));
  jxor g05226(.dina(n22205), .dinb(n349), .dout(n22489));
  jand g05227(.dina(n22489), .dinb(n22488), .dout(n22490));
  jor  g05228(.dina(n22490), .dinb(n22206), .dout(n22491));
  jxor g05229(.dina(n22200), .dinb(n268), .dout(n22492));
  jand g05230(.dina(n22492), .dinb(n22491), .dout(n22493));
  jor  g05231(.dina(n22493), .dinb(n22201), .dout(n22494));
  jxor g05232(.dina(n22195), .dinb(n274), .dout(n22495));
  jand g05233(.dina(n22495), .dinb(n22494), .dout(n22496));
  jor  g05234(.dina(n22496), .dinb(n22196), .dout(n22497));
  jxor g05235(.dina(n22190), .dinb(n269), .dout(n22498));
  jand g05236(.dina(n22498), .dinb(n22497), .dout(n22499));
  jor  g05237(.dina(n22499), .dinb(n22191), .dout(n22500));
  jxor g05238(.dina(n22185), .dinb(n270), .dout(n22501));
  jand g05239(.dina(n22501), .dinb(n22500), .dout(n22502));
  jor  g05240(.dina(n22502), .dinb(n22186), .dout(n22503));
  jxor g05241(.dina(n22173), .dinb(n271), .dout(n22504));
  jand g05242(.dina(n22504), .dinb(n22503), .dout(n22505));
  jor  g05243(.dina(n22505), .dinb(n22181), .dout(n22506));
  jand g05244(.dina(n22506), .dinb(n22180), .dout(n22507));
  jor  g05245(.dina(n22507), .dinb(n22177), .dout(n22508));
  jand g05246(.dina(n22508), .dinb(n3911), .dout(n22509));
  jor  g05247(.dina(n22509), .dinb(n22173), .dout(n22510));
  jnot g05248(.din(n22509), .dout(n22511));
  jxor g05249(.dina(n22504), .dinb(n22503), .dout(n22512));
  jor  g05250(.dina(n22512), .dinb(n22511), .dout(n22513));
  jand g05251(.dina(n22513), .dinb(n22510), .dout(n22514));
  jand g05252(.dina(n22506), .dinb(n414), .dout(n22515));
  jor  g05253(.dina(n22515), .dinb(n22511), .dout(n22516));
  jand g05254(.dina(n22516), .dinb(n22176), .dout(n22517));
  jand g05255(.dina(n22517), .dinb(n3911), .dout(n22518));
  jand g05256(.dina(n22514), .dinb(n338), .dout(n22519));
  jor  g05257(.dina(n22509), .dinb(n22185), .dout(n22520));
  jxor g05258(.dina(n22501), .dinb(n22500), .dout(n22521));
  jor  g05259(.dina(n22521), .dinb(n22511), .dout(n22522));
  jand g05260(.dina(n22522), .dinb(n22520), .dout(n22523));
  jand g05261(.dina(n22523), .dinb(n271), .dout(n22524));
  jor  g05262(.dina(n22509), .dinb(n22190), .dout(n22525));
  jxor g05263(.dina(n22498), .dinb(n22497), .dout(n22526));
  jor  g05264(.dina(n22526), .dinb(n22511), .dout(n22527));
  jand g05265(.dina(n22527), .dinb(n22525), .dout(n22528));
  jand g05266(.dina(n22528), .dinb(n270), .dout(n22529));
  jor  g05267(.dina(n22509), .dinb(n22195), .dout(n22530));
  jxor g05268(.dina(n22495), .dinb(n22494), .dout(n22531));
  jor  g05269(.dina(n22531), .dinb(n22511), .dout(n22532));
  jand g05270(.dina(n22532), .dinb(n22530), .dout(n22533));
  jand g05271(.dina(n22533), .dinb(n269), .dout(n22534));
  jor  g05272(.dina(n22509), .dinb(n22200), .dout(n22535));
  jxor g05273(.dina(n22492), .dinb(n22491), .dout(n22536));
  jor  g05274(.dina(n22536), .dinb(n22511), .dout(n22537));
  jand g05275(.dina(n22537), .dinb(n22535), .dout(n22538));
  jand g05276(.dina(n22538), .dinb(n274), .dout(n22539));
  jor  g05277(.dina(n22509), .dinb(n22205), .dout(n22540));
  jxor g05278(.dina(n22489), .dinb(n22488), .dout(n22541));
  jor  g05279(.dina(n22541), .dinb(n22511), .dout(n22542));
  jand g05280(.dina(n22542), .dinb(n22540), .dout(n22543));
  jand g05281(.dina(n22543), .dinb(n268), .dout(n22544));
  jor  g05282(.dina(n22509), .dinb(n22210), .dout(n22545));
  jxor g05283(.dina(n22486), .dinb(n22485), .dout(n22546));
  jor  g05284(.dina(n22546), .dinb(n22511), .dout(n22547));
  jand g05285(.dina(n22547), .dinb(n22545), .dout(n22548));
  jand g05286(.dina(n22548), .dinb(n349), .dout(n22549));
  jor  g05287(.dina(n22509), .dinb(n22215), .dout(n22550));
  jxor g05288(.dina(n22483), .dinb(n22482), .dout(n22551));
  jor  g05289(.dina(n22551), .dinb(n22511), .dout(n22552));
  jand g05290(.dina(n22552), .dinb(n22550), .dout(n22553));
  jand g05291(.dina(n22553), .dinb(n348), .dout(n22554));
  jor  g05292(.dina(n22509), .dinb(n22220), .dout(n22555));
  jxor g05293(.dina(n22480), .dinb(n22479), .dout(n22556));
  jor  g05294(.dina(n22556), .dinb(n22511), .dout(n22557));
  jand g05295(.dina(n22557), .dinb(n22555), .dout(n22558));
  jand g05296(.dina(n22558), .dinb(n347), .dout(n22559));
  jor  g05297(.dina(n22509), .dinb(n22225), .dout(n22560));
  jxor g05298(.dina(n22477), .dinb(n22476), .dout(n22561));
  jor  g05299(.dina(n22561), .dinb(n22511), .dout(n22562));
  jand g05300(.dina(n22562), .dinb(n22560), .dout(n22563));
  jand g05301(.dina(n22563), .dinb(n267), .dout(n22564));
  jor  g05302(.dina(n22509), .dinb(n22230), .dout(n22565));
  jxor g05303(.dina(n22474), .dinb(n22473), .dout(n22566));
  jor  g05304(.dina(n22566), .dinb(n22511), .dout(n22567));
  jand g05305(.dina(n22567), .dinb(n22565), .dout(n22568));
  jand g05306(.dina(n22568), .dinb(n266), .dout(n22569));
  jor  g05307(.dina(n22509), .dinb(n22235), .dout(n22570));
  jxor g05308(.dina(n22471), .dinb(n22470), .dout(n22571));
  jor  g05309(.dina(n22571), .dinb(n22511), .dout(n22572));
  jand g05310(.dina(n22572), .dinb(n22570), .dout(n22573));
  jand g05311(.dina(n22573), .dinb(n356), .dout(n22574));
  jor  g05312(.dina(n22509), .dinb(n22240), .dout(n22575));
  jxor g05313(.dina(n22468), .dinb(n22467), .dout(n22576));
  jor  g05314(.dina(n22576), .dinb(n22511), .dout(n22577));
  jand g05315(.dina(n22577), .dinb(n22575), .dout(n22578));
  jand g05316(.dina(n22578), .dinb(n355), .dout(n22579));
  jor  g05317(.dina(n22509), .dinb(n22245), .dout(n22580));
  jxor g05318(.dina(n22465), .dinb(n22464), .dout(n22581));
  jor  g05319(.dina(n22581), .dinb(n22511), .dout(n22582));
  jand g05320(.dina(n22582), .dinb(n22580), .dout(n22583));
  jand g05321(.dina(n22583), .dinb(n364), .dout(n22584));
  jor  g05322(.dina(n22509), .dinb(n22250), .dout(n22585));
  jxor g05323(.dina(n22462), .dinb(n22461), .dout(n22586));
  jor  g05324(.dina(n22586), .dinb(n22511), .dout(n22587));
  jand g05325(.dina(n22587), .dinb(n22585), .dout(n22588));
  jand g05326(.dina(n22588), .dinb(n361), .dout(n22589));
  jor  g05327(.dina(n22509), .dinb(n22255), .dout(n22590));
  jxor g05328(.dina(n22459), .dinb(n22458), .dout(n22591));
  jor  g05329(.dina(n22591), .dinb(n22511), .dout(n22592));
  jand g05330(.dina(n22592), .dinb(n22590), .dout(n22593));
  jand g05331(.dina(n22593), .dinb(n360), .dout(n22594));
  jor  g05332(.dina(n22509), .dinb(n22260), .dout(n22595));
  jxor g05333(.dina(n22456), .dinb(n22455), .dout(n22596));
  jor  g05334(.dina(n22596), .dinb(n22511), .dout(n22597));
  jand g05335(.dina(n22597), .dinb(n22595), .dout(n22598));
  jand g05336(.dina(n22598), .dinb(n363), .dout(n22599));
  jor  g05337(.dina(n22509), .dinb(n22265), .dout(n22600));
  jxor g05338(.dina(n22453), .dinb(n22452), .dout(n22601));
  jor  g05339(.dina(n22601), .dinb(n22511), .dout(n22602));
  jand g05340(.dina(n22602), .dinb(n22600), .dout(n22603));
  jand g05341(.dina(n22603), .dinb(n359), .dout(n22604));
  jor  g05342(.dina(n22509), .dinb(n22270), .dout(n22605));
  jxor g05343(.dina(n22450), .dinb(n22449), .dout(n22606));
  jor  g05344(.dina(n22606), .dinb(n22511), .dout(n22607));
  jand g05345(.dina(n22607), .dinb(n22605), .dout(n22608));
  jand g05346(.dina(n22608), .dinb(n369), .dout(n22609));
  jor  g05347(.dina(n22509), .dinb(n22275), .dout(n22610));
  jxor g05348(.dina(n22447), .dinb(n22446), .dout(n22611));
  jor  g05349(.dina(n22611), .dinb(n22511), .dout(n22612));
  jand g05350(.dina(n22612), .dinb(n22610), .dout(n22613));
  jand g05351(.dina(n22613), .dinb(n368), .dout(n22614));
  jor  g05352(.dina(n22509), .dinb(n22280), .dout(n22615));
  jxor g05353(.dina(n22444), .dinb(n22443), .dout(n22616));
  jor  g05354(.dina(n22616), .dinb(n22511), .dout(n22617));
  jand g05355(.dina(n22617), .dinb(n22615), .dout(n22618));
  jand g05356(.dina(n22618), .dinb(n367), .dout(n22619));
  jor  g05357(.dina(n22509), .dinb(n22285), .dout(n22620));
  jxor g05358(.dina(n22441), .dinb(n22440), .dout(n22621));
  jor  g05359(.dina(n22621), .dinb(n22511), .dout(n22622));
  jand g05360(.dina(n22622), .dinb(n22620), .dout(n22623));
  jand g05361(.dina(n22623), .dinb(n265), .dout(n22624));
  jor  g05362(.dina(n22509), .dinb(n22290), .dout(n22625));
  jxor g05363(.dina(n22438), .dinb(n22437), .dout(n22626));
  jor  g05364(.dina(n22626), .dinb(n22511), .dout(n22627));
  jand g05365(.dina(n22627), .dinb(n22625), .dout(n22628));
  jand g05366(.dina(n22628), .dinb(n378), .dout(n22629));
  jor  g05367(.dina(n22509), .dinb(n22296), .dout(n22630));
  jxor g05368(.dina(n22435), .dinb(n22434), .dout(n22631));
  jor  g05369(.dina(n22631), .dinb(n22511), .dout(n22632));
  jand g05370(.dina(n22632), .dinb(n22630), .dout(n22633));
  jand g05371(.dina(n22633), .dinb(n377), .dout(n22634));
  jor  g05372(.dina(n22509), .dinb(n22301), .dout(n22635));
  jxor g05373(.dina(n22432), .dinb(n22431), .dout(n22636));
  jor  g05374(.dina(n22636), .dinb(n22511), .dout(n22637));
  jand g05375(.dina(n22637), .dinb(n22635), .dout(n22638));
  jand g05376(.dina(n22638), .dinb(n376), .dout(n22639));
  jor  g05377(.dina(n22509), .dinb(n22306), .dout(n22640));
  jxor g05378(.dina(n22429), .dinb(n22428), .dout(n22641));
  jor  g05379(.dina(n22641), .dinb(n22511), .dout(n22642));
  jand g05380(.dina(n22642), .dinb(n22640), .dout(n22643));
  jand g05381(.dina(n22643), .dinb(n264), .dout(n22644));
  jor  g05382(.dina(n22509), .dinb(n22425), .dout(n22645));
  jxor g05383(.dina(n22426), .dinb(n4055), .dout(n22646));
  jand g05384(.dina(n22646), .dinb(n22509), .dout(n22647));
  jnot g05385(.din(n22647), .dout(n22648));
  jand g05386(.dina(n22648), .dinb(n22645), .dout(n22649));
  jnot g05387(.din(n22649), .dout(n22650));
  jand g05388(.dina(n22650), .dinb(n386), .dout(n22651));
  jnot g05389(.din(n4278), .dout(n22652));
  jnot g05390(.din(n22177), .dout(n22653));
  jnot g05391(.din(n22181), .dout(n22654));
  jnot g05392(.din(n22186), .dout(n22655));
  jnot g05393(.din(n22191), .dout(n22656));
  jnot g05394(.din(n22196), .dout(n22657));
  jnot g05395(.din(n22201), .dout(n22658));
  jnot g05396(.din(n22206), .dout(n22659));
  jnot g05397(.din(n22211), .dout(n22660));
  jnot g05398(.din(n22216), .dout(n22661));
  jnot g05399(.din(n22221), .dout(n22662));
  jnot g05400(.din(n22226), .dout(n22663));
  jnot g05401(.din(n22231), .dout(n22664));
  jnot g05402(.din(n22236), .dout(n22665));
  jnot g05403(.din(n22241), .dout(n22666));
  jnot g05404(.din(n22246), .dout(n22667));
  jnot g05405(.din(n22251), .dout(n22668));
  jnot g05406(.din(n22256), .dout(n22669));
  jnot g05407(.din(n22261), .dout(n22670));
  jnot g05408(.din(n22266), .dout(n22671));
  jnot g05409(.din(n22271), .dout(n22672));
  jnot g05410(.din(n22276), .dout(n22673));
  jnot g05411(.din(n22281), .dout(n22674));
  jnot g05412(.din(n22286), .dout(n22675));
  jnot g05413(.din(n22291), .dout(n22676));
  jnot g05414(.din(n22297), .dout(n22677));
  jnot g05415(.din(n22302), .dout(n22678));
  jnot g05416(.din(n22307), .dout(n22679));
  jnot g05417(.din(n22422), .dout(n22680));
  jxor g05418(.dina(n22425), .dinb(n259), .dout(n22681));
  jor  g05419(.dina(n22681), .dinb(n4054), .dout(n22682));
  jand g05420(.dina(n22682), .dinb(n22680), .dout(n22683));
  jnot g05421(.din(n22429), .dout(n22684));
  jor  g05422(.dina(n22684), .dinb(n22683), .dout(n22685));
  jand g05423(.dina(n22685), .dinb(n22679), .dout(n22686));
  jnot g05424(.din(n22432), .dout(n22687));
  jor  g05425(.dina(n22687), .dinb(n22686), .dout(n22688));
  jand g05426(.dina(n22688), .dinb(n22678), .dout(n22689));
  jnot g05427(.din(n22435), .dout(n22690));
  jor  g05428(.dina(n22690), .dinb(n22689), .dout(n22691));
  jand g05429(.dina(n22691), .dinb(n22677), .dout(n22692));
  jnot g05430(.din(n22438), .dout(n22693));
  jor  g05431(.dina(n22693), .dinb(n22692), .dout(n22694));
  jand g05432(.dina(n22694), .dinb(n22676), .dout(n22695));
  jnot g05433(.din(n22441), .dout(n22696));
  jor  g05434(.dina(n22696), .dinb(n22695), .dout(n22697));
  jand g05435(.dina(n22697), .dinb(n22675), .dout(n22698));
  jnot g05436(.din(n22444), .dout(n22699));
  jor  g05437(.dina(n22699), .dinb(n22698), .dout(n22700));
  jand g05438(.dina(n22700), .dinb(n22674), .dout(n22701));
  jnot g05439(.din(n22447), .dout(n22702));
  jor  g05440(.dina(n22702), .dinb(n22701), .dout(n22703));
  jand g05441(.dina(n22703), .dinb(n22673), .dout(n22704));
  jnot g05442(.din(n22450), .dout(n22705));
  jor  g05443(.dina(n22705), .dinb(n22704), .dout(n22706));
  jand g05444(.dina(n22706), .dinb(n22672), .dout(n22707));
  jnot g05445(.din(n22453), .dout(n22708));
  jor  g05446(.dina(n22708), .dinb(n22707), .dout(n22709));
  jand g05447(.dina(n22709), .dinb(n22671), .dout(n22710));
  jnot g05448(.din(n22456), .dout(n22711));
  jor  g05449(.dina(n22711), .dinb(n22710), .dout(n22712));
  jand g05450(.dina(n22712), .dinb(n22670), .dout(n22713));
  jnot g05451(.din(n22459), .dout(n22714));
  jor  g05452(.dina(n22714), .dinb(n22713), .dout(n22715));
  jand g05453(.dina(n22715), .dinb(n22669), .dout(n22716));
  jnot g05454(.din(n22462), .dout(n22717));
  jor  g05455(.dina(n22717), .dinb(n22716), .dout(n22718));
  jand g05456(.dina(n22718), .dinb(n22668), .dout(n22719));
  jnot g05457(.din(n22465), .dout(n22720));
  jor  g05458(.dina(n22720), .dinb(n22719), .dout(n22721));
  jand g05459(.dina(n22721), .dinb(n22667), .dout(n22722));
  jnot g05460(.din(n22468), .dout(n22723));
  jor  g05461(.dina(n22723), .dinb(n22722), .dout(n22724));
  jand g05462(.dina(n22724), .dinb(n22666), .dout(n22725));
  jnot g05463(.din(n22471), .dout(n22726));
  jor  g05464(.dina(n22726), .dinb(n22725), .dout(n22727));
  jand g05465(.dina(n22727), .dinb(n22665), .dout(n22728));
  jnot g05466(.din(n22474), .dout(n22729));
  jor  g05467(.dina(n22729), .dinb(n22728), .dout(n22730));
  jand g05468(.dina(n22730), .dinb(n22664), .dout(n22731));
  jnot g05469(.din(n22477), .dout(n22732));
  jor  g05470(.dina(n22732), .dinb(n22731), .dout(n22733));
  jand g05471(.dina(n22733), .dinb(n22663), .dout(n22734));
  jnot g05472(.din(n22480), .dout(n22735));
  jor  g05473(.dina(n22735), .dinb(n22734), .dout(n22736));
  jand g05474(.dina(n22736), .dinb(n22662), .dout(n22737));
  jnot g05475(.din(n22483), .dout(n22738));
  jor  g05476(.dina(n22738), .dinb(n22737), .dout(n22739));
  jand g05477(.dina(n22739), .dinb(n22661), .dout(n22740));
  jnot g05478(.din(n22486), .dout(n22741));
  jor  g05479(.dina(n22741), .dinb(n22740), .dout(n22742));
  jand g05480(.dina(n22742), .dinb(n22660), .dout(n22743));
  jnot g05481(.din(n22489), .dout(n22744));
  jor  g05482(.dina(n22744), .dinb(n22743), .dout(n22745));
  jand g05483(.dina(n22745), .dinb(n22659), .dout(n22746));
  jnot g05484(.din(n22492), .dout(n22747));
  jor  g05485(.dina(n22747), .dinb(n22746), .dout(n22748));
  jand g05486(.dina(n22748), .dinb(n22658), .dout(n22749));
  jnot g05487(.din(n22495), .dout(n22750));
  jor  g05488(.dina(n22750), .dinb(n22749), .dout(n22751));
  jand g05489(.dina(n22751), .dinb(n22657), .dout(n22752));
  jnot g05490(.din(n22498), .dout(n22753));
  jor  g05491(.dina(n22753), .dinb(n22752), .dout(n22754));
  jand g05492(.dina(n22754), .dinb(n22656), .dout(n22755));
  jnot g05493(.din(n22501), .dout(n22756));
  jor  g05494(.dina(n22756), .dinb(n22755), .dout(n22757));
  jand g05495(.dina(n22757), .dinb(n22655), .dout(n22758));
  jnot g05496(.din(n22504), .dout(n22759));
  jor  g05497(.dina(n22759), .dinb(n22758), .dout(n22760));
  jand g05498(.dina(n22760), .dinb(n22654), .dout(n22761));
  jor  g05499(.dina(n22761), .dinb(n22179), .dout(n22762));
  jand g05500(.dina(n22762), .dinb(n22653), .dout(n22763));
  jor  g05501(.dina(n22763), .dinb(n22652), .dout(n22764));
  jand g05502(.dina(n22764), .dinb(a35 ), .dout(n22765));
  jnot g05503(.din(n4281), .dout(n22766));
  jor  g05504(.dina(n22763), .dinb(n22766), .dout(n22767));
  jnot g05505(.din(n22767), .dout(n22768));
  jor  g05506(.dina(n22768), .dinb(n22765), .dout(n22769));
  jand g05507(.dina(n22769), .dinb(n259), .dout(n22770));
  jand g05508(.dina(n22508), .dinb(n4278), .dout(n22771));
  jor  g05509(.dina(n22771), .dinb(n4053), .dout(n22772));
  jand g05510(.dina(n22767), .dinb(n22772), .dout(n22773));
  jxor g05511(.dina(n22773), .dinb(b1 ), .dout(n22774));
  jand g05512(.dina(n22774), .dinb(n4289), .dout(n22775));
  jor  g05513(.dina(n22775), .dinb(n22770), .dout(n22776));
  jxor g05514(.dina(n22649), .dinb(b2 ), .dout(n22777));
  jand g05515(.dina(n22777), .dinb(n22776), .dout(n22778));
  jor  g05516(.dina(n22778), .dinb(n22651), .dout(n22779));
  jxor g05517(.dina(n22643), .dinb(n264), .dout(n22780));
  jand g05518(.dina(n22780), .dinb(n22779), .dout(n22781));
  jor  g05519(.dina(n22781), .dinb(n22644), .dout(n22782));
  jxor g05520(.dina(n22638), .dinb(n376), .dout(n22783));
  jand g05521(.dina(n22783), .dinb(n22782), .dout(n22784));
  jor  g05522(.dina(n22784), .dinb(n22639), .dout(n22785));
  jxor g05523(.dina(n22633), .dinb(n377), .dout(n22786));
  jand g05524(.dina(n22786), .dinb(n22785), .dout(n22787));
  jor  g05525(.dina(n22787), .dinb(n22634), .dout(n22788));
  jxor g05526(.dina(n22628), .dinb(n378), .dout(n22789));
  jand g05527(.dina(n22789), .dinb(n22788), .dout(n22790));
  jor  g05528(.dina(n22790), .dinb(n22629), .dout(n22791));
  jxor g05529(.dina(n22623), .dinb(n265), .dout(n22792));
  jand g05530(.dina(n22792), .dinb(n22791), .dout(n22793));
  jor  g05531(.dina(n22793), .dinb(n22624), .dout(n22794));
  jxor g05532(.dina(n22618), .dinb(n367), .dout(n22795));
  jand g05533(.dina(n22795), .dinb(n22794), .dout(n22796));
  jor  g05534(.dina(n22796), .dinb(n22619), .dout(n22797));
  jxor g05535(.dina(n22613), .dinb(n368), .dout(n22798));
  jand g05536(.dina(n22798), .dinb(n22797), .dout(n22799));
  jor  g05537(.dina(n22799), .dinb(n22614), .dout(n22800));
  jxor g05538(.dina(n22608), .dinb(n369), .dout(n22801));
  jand g05539(.dina(n22801), .dinb(n22800), .dout(n22802));
  jor  g05540(.dina(n22802), .dinb(n22609), .dout(n22803));
  jxor g05541(.dina(n22603), .dinb(n359), .dout(n22804));
  jand g05542(.dina(n22804), .dinb(n22803), .dout(n22805));
  jor  g05543(.dina(n22805), .dinb(n22604), .dout(n22806));
  jxor g05544(.dina(n22598), .dinb(n363), .dout(n22807));
  jand g05545(.dina(n22807), .dinb(n22806), .dout(n22808));
  jor  g05546(.dina(n22808), .dinb(n22599), .dout(n22809));
  jxor g05547(.dina(n22593), .dinb(n360), .dout(n22810));
  jand g05548(.dina(n22810), .dinb(n22809), .dout(n22811));
  jor  g05549(.dina(n22811), .dinb(n22594), .dout(n22812));
  jxor g05550(.dina(n22588), .dinb(n361), .dout(n22813));
  jand g05551(.dina(n22813), .dinb(n22812), .dout(n22814));
  jor  g05552(.dina(n22814), .dinb(n22589), .dout(n22815));
  jxor g05553(.dina(n22583), .dinb(n364), .dout(n22816));
  jand g05554(.dina(n22816), .dinb(n22815), .dout(n22817));
  jor  g05555(.dina(n22817), .dinb(n22584), .dout(n22818));
  jxor g05556(.dina(n22578), .dinb(n355), .dout(n22819));
  jand g05557(.dina(n22819), .dinb(n22818), .dout(n22820));
  jor  g05558(.dina(n22820), .dinb(n22579), .dout(n22821));
  jxor g05559(.dina(n22573), .dinb(n356), .dout(n22822));
  jand g05560(.dina(n22822), .dinb(n22821), .dout(n22823));
  jor  g05561(.dina(n22823), .dinb(n22574), .dout(n22824));
  jxor g05562(.dina(n22568), .dinb(n266), .dout(n22825));
  jand g05563(.dina(n22825), .dinb(n22824), .dout(n22826));
  jor  g05564(.dina(n22826), .dinb(n22569), .dout(n22827));
  jxor g05565(.dina(n22563), .dinb(n267), .dout(n22828));
  jand g05566(.dina(n22828), .dinb(n22827), .dout(n22829));
  jor  g05567(.dina(n22829), .dinb(n22564), .dout(n22830));
  jxor g05568(.dina(n22558), .dinb(n347), .dout(n22831));
  jand g05569(.dina(n22831), .dinb(n22830), .dout(n22832));
  jor  g05570(.dina(n22832), .dinb(n22559), .dout(n22833));
  jxor g05571(.dina(n22553), .dinb(n348), .dout(n22834));
  jand g05572(.dina(n22834), .dinb(n22833), .dout(n22835));
  jor  g05573(.dina(n22835), .dinb(n22554), .dout(n22836));
  jxor g05574(.dina(n22548), .dinb(n349), .dout(n22837));
  jand g05575(.dina(n22837), .dinb(n22836), .dout(n22838));
  jor  g05576(.dina(n22838), .dinb(n22549), .dout(n22839));
  jxor g05577(.dina(n22543), .dinb(n268), .dout(n22840));
  jand g05578(.dina(n22840), .dinb(n22839), .dout(n22841));
  jor  g05579(.dina(n22841), .dinb(n22544), .dout(n22842));
  jxor g05580(.dina(n22538), .dinb(n274), .dout(n22843));
  jand g05581(.dina(n22843), .dinb(n22842), .dout(n22844));
  jor  g05582(.dina(n22844), .dinb(n22539), .dout(n22845));
  jxor g05583(.dina(n22533), .dinb(n269), .dout(n22846));
  jand g05584(.dina(n22846), .dinb(n22845), .dout(n22847));
  jor  g05585(.dina(n22847), .dinb(n22534), .dout(n22848));
  jxor g05586(.dina(n22528), .dinb(n270), .dout(n22849));
  jand g05587(.dina(n22849), .dinb(n22848), .dout(n22850));
  jor  g05588(.dina(n22850), .dinb(n22529), .dout(n22851));
  jxor g05589(.dina(n22523), .dinb(n271), .dout(n22852));
  jand g05590(.dina(n22852), .dinb(n22851), .dout(n22853));
  jor  g05591(.dina(n22853), .dinb(n22524), .dout(n22854));
  jxor g05592(.dina(n22514), .dinb(n338), .dout(n22855));
  jand g05593(.dina(n22855), .dinb(n22854), .dout(n22856));
  jor  g05594(.dina(n22856), .dinb(n22519), .dout(n22857));
  jxor g05595(.dina(n22517), .dinb(b29 ), .dout(n22858));
  jnot g05596(.din(n22858), .dout(n22859));
  jand g05597(.dina(n22859), .dinb(n22857), .dout(n22860));
  jand g05598(.dina(n22860), .dinb(n4145), .dout(n22861));
  jor  g05599(.dina(n22861), .dinb(n22518), .dout(n22862));
  jor  g05600(.dina(n22862), .dinb(n22514), .dout(n22863));
  jnot g05601(.din(n22862), .dout(n22864));
  jxor g05602(.dina(n22855), .dinb(n22854), .dout(n22865));
  jor  g05603(.dina(n22865), .dinb(n22864), .dout(n22866));
  jand g05604(.dina(n22866), .dinb(n22863), .dout(n22867));
  jxor g05605(.dina(n22859), .dinb(n22857), .dout(n22868));
  jand g05606(.dina(n22868), .dinb(n22518), .dout(n22869));
  jand g05607(.dina(n22864), .dinb(n22517), .dout(n22870));
  jor  g05608(.dina(n22870), .dinb(n22869), .dout(n22871));
  jand g05609(.dina(n22871), .dinb(n340), .dout(n22872));
  jnot g05610(.din(n22871), .dout(n22873));
  jand g05611(.dina(n22873), .dinb(b30 ), .dout(n22874));
  jnot g05612(.din(n22874), .dout(n22875));
  jand g05613(.dina(n22867), .dinb(n339), .dout(n22876));
  jor  g05614(.dina(n22862), .dinb(n22523), .dout(n22877));
  jxor g05615(.dina(n22852), .dinb(n22851), .dout(n22878));
  jor  g05616(.dina(n22878), .dinb(n22864), .dout(n22879));
  jand g05617(.dina(n22879), .dinb(n22877), .dout(n22880));
  jand g05618(.dina(n22880), .dinb(n338), .dout(n22881));
  jor  g05619(.dina(n22862), .dinb(n22528), .dout(n22882));
  jxor g05620(.dina(n22849), .dinb(n22848), .dout(n22883));
  jor  g05621(.dina(n22883), .dinb(n22864), .dout(n22884));
  jand g05622(.dina(n22884), .dinb(n22882), .dout(n22885));
  jand g05623(.dina(n22885), .dinb(n271), .dout(n22886));
  jor  g05624(.dina(n22862), .dinb(n22533), .dout(n22887));
  jxor g05625(.dina(n22846), .dinb(n22845), .dout(n22888));
  jor  g05626(.dina(n22888), .dinb(n22864), .dout(n22889));
  jand g05627(.dina(n22889), .dinb(n22887), .dout(n22890));
  jand g05628(.dina(n22890), .dinb(n270), .dout(n22891));
  jor  g05629(.dina(n22862), .dinb(n22538), .dout(n22892));
  jxor g05630(.dina(n22843), .dinb(n22842), .dout(n22893));
  jor  g05631(.dina(n22893), .dinb(n22864), .dout(n22894));
  jand g05632(.dina(n22894), .dinb(n22892), .dout(n22895));
  jand g05633(.dina(n22895), .dinb(n269), .dout(n22896));
  jor  g05634(.dina(n22862), .dinb(n22543), .dout(n22897));
  jxor g05635(.dina(n22840), .dinb(n22839), .dout(n22898));
  jor  g05636(.dina(n22898), .dinb(n22864), .dout(n22899));
  jand g05637(.dina(n22899), .dinb(n22897), .dout(n22900));
  jand g05638(.dina(n22900), .dinb(n274), .dout(n22901));
  jor  g05639(.dina(n22862), .dinb(n22548), .dout(n22902));
  jxor g05640(.dina(n22837), .dinb(n22836), .dout(n22903));
  jor  g05641(.dina(n22903), .dinb(n22864), .dout(n22904));
  jand g05642(.dina(n22904), .dinb(n22902), .dout(n22905));
  jand g05643(.dina(n22905), .dinb(n268), .dout(n22906));
  jor  g05644(.dina(n22862), .dinb(n22553), .dout(n22907));
  jxor g05645(.dina(n22834), .dinb(n22833), .dout(n22908));
  jor  g05646(.dina(n22908), .dinb(n22864), .dout(n22909));
  jand g05647(.dina(n22909), .dinb(n22907), .dout(n22910));
  jand g05648(.dina(n22910), .dinb(n349), .dout(n22911));
  jor  g05649(.dina(n22862), .dinb(n22558), .dout(n22912));
  jxor g05650(.dina(n22831), .dinb(n22830), .dout(n22913));
  jor  g05651(.dina(n22913), .dinb(n22864), .dout(n22914));
  jand g05652(.dina(n22914), .dinb(n22912), .dout(n22915));
  jand g05653(.dina(n22915), .dinb(n348), .dout(n22916));
  jor  g05654(.dina(n22862), .dinb(n22563), .dout(n22917));
  jxor g05655(.dina(n22828), .dinb(n22827), .dout(n22918));
  jor  g05656(.dina(n22918), .dinb(n22864), .dout(n22919));
  jand g05657(.dina(n22919), .dinb(n22917), .dout(n22920));
  jand g05658(.dina(n22920), .dinb(n347), .dout(n22921));
  jor  g05659(.dina(n22862), .dinb(n22568), .dout(n22922));
  jxor g05660(.dina(n22825), .dinb(n22824), .dout(n22923));
  jor  g05661(.dina(n22923), .dinb(n22864), .dout(n22924));
  jand g05662(.dina(n22924), .dinb(n22922), .dout(n22925));
  jand g05663(.dina(n22925), .dinb(n267), .dout(n22926));
  jor  g05664(.dina(n22862), .dinb(n22573), .dout(n22927));
  jxor g05665(.dina(n22822), .dinb(n22821), .dout(n22928));
  jor  g05666(.dina(n22928), .dinb(n22864), .dout(n22929));
  jand g05667(.dina(n22929), .dinb(n22927), .dout(n22930));
  jand g05668(.dina(n22930), .dinb(n266), .dout(n22931));
  jor  g05669(.dina(n22862), .dinb(n22578), .dout(n22932));
  jxor g05670(.dina(n22819), .dinb(n22818), .dout(n22933));
  jor  g05671(.dina(n22933), .dinb(n22864), .dout(n22934));
  jand g05672(.dina(n22934), .dinb(n22932), .dout(n22935));
  jand g05673(.dina(n22935), .dinb(n356), .dout(n22936));
  jor  g05674(.dina(n22862), .dinb(n22583), .dout(n22937));
  jxor g05675(.dina(n22816), .dinb(n22815), .dout(n22938));
  jor  g05676(.dina(n22938), .dinb(n22864), .dout(n22939));
  jand g05677(.dina(n22939), .dinb(n22937), .dout(n22940));
  jand g05678(.dina(n22940), .dinb(n355), .dout(n22941));
  jor  g05679(.dina(n22862), .dinb(n22588), .dout(n22942));
  jxor g05680(.dina(n22813), .dinb(n22812), .dout(n22943));
  jor  g05681(.dina(n22943), .dinb(n22864), .dout(n22944));
  jand g05682(.dina(n22944), .dinb(n22942), .dout(n22945));
  jand g05683(.dina(n22945), .dinb(n364), .dout(n22946));
  jor  g05684(.dina(n22862), .dinb(n22593), .dout(n22947));
  jxor g05685(.dina(n22810), .dinb(n22809), .dout(n22948));
  jor  g05686(.dina(n22948), .dinb(n22864), .dout(n22949));
  jand g05687(.dina(n22949), .dinb(n22947), .dout(n22950));
  jand g05688(.dina(n22950), .dinb(n361), .dout(n22951));
  jor  g05689(.dina(n22862), .dinb(n22598), .dout(n22952));
  jxor g05690(.dina(n22807), .dinb(n22806), .dout(n22953));
  jor  g05691(.dina(n22953), .dinb(n22864), .dout(n22954));
  jand g05692(.dina(n22954), .dinb(n22952), .dout(n22955));
  jand g05693(.dina(n22955), .dinb(n360), .dout(n22956));
  jor  g05694(.dina(n22862), .dinb(n22603), .dout(n22957));
  jxor g05695(.dina(n22804), .dinb(n22803), .dout(n22958));
  jor  g05696(.dina(n22958), .dinb(n22864), .dout(n22959));
  jand g05697(.dina(n22959), .dinb(n22957), .dout(n22960));
  jand g05698(.dina(n22960), .dinb(n363), .dout(n22961));
  jor  g05699(.dina(n22862), .dinb(n22608), .dout(n22962));
  jxor g05700(.dina(n22801), .dinb(n22800), .dout(n22963));
  jor  g05701(.dina(n22963), .dinb(n22864), .dout(n22964));
  jand g05702(.dina(n22964), .dinb(n22962), .dout(n22965));
  jand g05703(.dina(n22965), .dinb(n359), .dout(n22966));
  jor  g05704(.dina(n22862), .dinb(n22613), .dout(n22967));
  jxor g05705(.dina(n22798), .dinb(n22797), .dout(n22968));
  jor  g05706(.dina(n22968), .dinb(n22864), .dout(n22969));
  jand g05707(.dina(n22969), .dinb(n22967), .dout(n22970));
  jand g05708(.dina(n22970), .dinb(n369), .dout(n22971));
  jor  g05709(.dina(n22862), .dinb(n22618), .dout(n22972));
  jxor g05710(.dina(n22795), .dinb(n22794), .dout(n22973));
  jor  g05711(.dina(n22973), .dinb(n22864), .dout(n22974));
  jand g05712(.dina(n22974), .dinb(n22972), .dout(n22975));
  jand g05713(.dina(n22975), .dinb(n368), .dout(n22976));
  jor  g05714(.dina(n22862), .dinb(n22623), .dout(n22977));
  jxor g05715(.dina(n22792), .dinb(n22791), .dout(n22978));
  jor  g05716(.dina(n22978), .dinb(n22864), .dout(n22979));
  jand g05717(.dina(n22979), .dinb(n22977), .dout(n22980));
  jand g05718(.dina(n22980), .dinb(n367), .dout(n22981));
  jor  g05719(.dina(n22862), .dinb(n22628), .dout(n22982));
  jxor g05720(.dina(n22789), .dinb(n22788), .dout(n22983));
  jor  g05721(.dina(n22983), .dinb(n22864), .dout(n22984));
  jand g05722(.dina(n22984), .dinb(n22982), .dout(n22985));
  jand g05723(.dina(n22985), .dinb(n265), .dout(n22986));
  jor  g05724(.dina(n22862), .dinb(n22633), .dout(n22987));
  jxor g05725(.dina(n22786), .dinb(n22785), .dout(n22988));
  jor  g05726(.dina(n22988), .dinb(n22864), .dout(n22989));
  jand g05727(.dina(n22989), .dinb(n22987), .dout(n22990));
  jand g05728(.dina(n22990), .dinb(n378), .dout(n22991));
  jor  g05729(.dina(n22862), .dinb(n22638), .dout(n22992));
  jxor g05730(.dina(n22783), .dinb(n22782), .dout(n22993));
  jor  g05731(.dina(n22993), .dinb(n22864), .dout(n22994));
  jand g05732(.dina(n22994), .dinb(n22992), .dout(n22995));
  jand g05733(.dina(n22995), .dinb(n377), .dout(n22996));
  jor  g05734(.dina(n22862), .dinb(n22643), .dout(n22997));
  jxor g05735(.dina(n22780), .dinb(n22779), .dout(n22998));
  jor  g05736(.dina(n22998), .dinb(n22864), .dout(n22999));
  jand g05737(.dina(n22999), .dinb(n22997), .dout(n23000));
  jand g05738(.dina(n23000), .dinb(n376), .dout(n23001));
  jor  g05739(.dina(n22862), .dinb(n22650), .dout(n23002));
  jxor g05740(.dina(n22777), .dinb(n22776), .dout(n23003));
  jor  g05741(.dina(n23003), .dinb(n22864), .dout(n23004));
  jand g05742(.dina(n23004), .dinb(n23002), .dout(n23005));
  jand g05743(.dina(n23005), .dinb(n264), .dout(n23006));
  jor  g05744(.dina(n22862), .dinb(n22769), .dout(n23007));
  jxor g05745(.dina(n22774), .dinb(n4289), .dout(n23008));
  jor  g05746(.dina(n23008), .dinb(n22864), .dout(n23009));
  jand g05747(.dina(n23009), .dinb(n23007), .dout(n23010));
  jand g05748(.dina(n23010), .dinb(n386), .dout(n23011));
  jand g05749(.dina(n22862), .dinb(b0 ), .dout(n23012));
  jxor g05750(.dina(n23012), .dinb(a34 ), .dout(n23013));
  jand g05751(.dina(n23013), .dinb(n259), .dout(n23014));
  jxor g05752(.dina(n23012), .dinb(n4287), .dout(n23015));
  jxor g05753(.dina(n23015), .dinb(b1 ), .dout(n23016));
  jand g05754(.dina(n23016), .dinb(n4542), .dout(n23017));
  jor  g05755(.dina(n23017), .dinb(n23014), .dout(n23018));
  jxor g05756(.dina(n23010), .dinb(n386), .dout(n23019));
  jand g05757(.dina(n23019), .dinb(n23018), .dout(n23020));
  jor  g05758(.dina(n23020), .dinb(n23011), .dout(n23021));
  jxor g05759(.dina(n23005), .dinb(n264), .dout(n23022));
  jand g05760(.dina(n23022), .dinb(n23021), .dout(n23023));
  jor  g05761(.dina(n23023), .dinb(n23006), .dout(n23024));
  jxor g05762(.dina(n23000), .dinb(n376), .dout(n23025));
  jand g05763(.dina(n23025), .dinb(n23024), .dout(n23026));
  jor  g05764(.dina(n23026), .dinb(n23001), .dout(n23027));
  jxor g05765(.dina(n22995), .dinb(n377), .dout(n23028));
  jand g05766(.dina(n23028), .dinb(n23027), .dout(n23029));
  jor  g05767(.dina(n23029), .dinb(n22996), .dout(n23030));
  jxor g05768(.dina(n22990), .dinb(n378), .dout(n23031));
  jand g05769(.dina(n23031), .dinb(n23030), .dout(n23032));
  jor  g05770(.dina(n23032), .dinb(n22991), .dout(n23033));
  jxor g05771(.dina(n22985), .dinb(n265), .dout(n23034));
  jand g05772(.dina(n23034), .dinb(n23033), .dout(n23035));
  jor  g05773(.dina(n23035), .dinb(n22986), .dout(n23036));
  jxor g05774(.dina(n22980), .dinb(n367), .dout(n23037));
  jand g05775(.dina(n23037), .dinb(n23036), .dout(n23038));
  jor  g05776(.dina(n23038), .dinb(n22981), .dout(n23039));
  jxor g05777(.dina(n22975), .dinb(n368), .dout(n23040));
  jand g05778(.dina(n23040), .dinb(n23039), .dout(n23041));
  jor  g05779(.dina(n23041), .dinb(n22976), .dout(n23042));
  jxor g05780(.dina(n22970), .dinb(n369), .dout(n23043));
  jand g05781(.dina(n23043), .dinb(n23042), .dout(n23044));
  jor  g05782(.dina(n23044), .dinb(n22971), .dout(n23045));
  jxor g05783(.dina(n22965), .dinb(n359), .dout(n23046));
  jand g05784(.dina(n23046), .dinb(n23045), .dout(n23047));
  jor  g05785(.dina(n23047), .dinb(n22966), .dout(n23048));
  jxor g05786(.dina(n22960), .dinb(n363), .dout(n23049));
  jand g05787(.dina(n23049), .dinb(n23048), .dout(n23050));
  jor  g05788(.dina(n23050), .dinb(n22961), .dout(n23051));
  jxor g05789(.dina(n22955), .dinb(n360), .dout(n23052));
  jand g05790(.dina(n23052), .dinb(n23051), .dout(n23053));
  jor  g05791(.dina(n23053), .dinb(n22956), .dout(n23054));
  jxor g05792(.dina(n22950), .dinb(n361), .dout(n23055));
  jand g05793(.dina(n23055), .dinb(n23054), .dout(n23056));
  jor  g05794(.dina(n23056), .dinb(n22951), .dout(n23057));
  jxor g05795(.dina(n22945), .dinb(n364), .dout(n23058));
  jand g05796(.dina(n23058), .dinb(n23057), .dout(n23059));
  jor  g05797(.dina(n23059), .dinb(n22946), .dout(n23060));
  jxor g05798(.dina(n22940), .dinb(n355), .dout(n23061));
  jand g05799(.dina(n23061), .dinb(n23060), .dout(n23062));
  jor  g05800(.dina(n23062), .dinb(n22941), .dout(n23063));
  jxor g05801(.dina(n22935), .dinb(n356), .dout(n23064));
  jand g05802(.dina(n23064), .dinb(n23063), .dout(n23065));
  jor  g05803(.dina(n23065), .dinb(n22936), .dout(n23066));
  jxor g05804(.dina(n22930), .dinb(n266), .dout(n23067));
  jand g05805(.dina(n23067), .dinb(n23066), .dout(n23068));
  jor  g05806(.dina(n23068), .dinb(n22931), .dout(n23069));
  jxor g05807(.dina(n22925), .dinb(n267), .dout(n23070));
  jand g05808(.dina(n23070), .dinb(n23069), .dout(n23071));
  jor  g05809(.dina(n23071), .dinb(n22926), .dout(n23072));
  jxor g05810(.dina(n22920), .dinb(n347), .dout(n23073));
  jand g05811(.dina(n23073), .dinb(n23072), .dout(n23074));
  jor  g05812(.dina(n23074), .dinb(n22921), .dout(n23075));
  jxor g05813(.dina(n22915), .dinb(n348), .dout(n23076));
  jand g05814(.dina(n23076), .dinb(n23075), .dout(n23077));
  jor  g05815(.dina(n23077), .dinb(n22916), .dout(n23078));
  jxor g05816(.dina(n22910), .dinb(n349), .dout(n23079));
  jand g05817(.dina(n23079), .dinb(n23078), .dout(n23080));
  jor  g05818(.dina(n23080), .dinb(n22911), .dout(n23081));
  jxor g05819(.dina(n22905), .dinb(n268), .dout(n23082));
  jand g05820(.dina(n23082), .dinb(n23081), .dout(n23083));
  jor  g05821(.dina(n23083), .dinb(n22906), .dout(n23084));
  jxor g05822(.dina(n22900), .dinb(n274), .dout(n23085));
  jand g05823(.dina(n23085), .dinb(n23084), .dout(n23086));
  jor  g05824(.dina(n23086), .dinb(n22901), .dout(n23087));
  jxor g05825(.dina(n22895), .dinb(n269), .dout(n23088));
  jand g05826(.dina(n23088), .dinb(n23087), .dout(n23089));
  jor  g05827(.dina(n23089), .dinb(n22896), .dout(n23090));
  jxor g05828(.dina(n22890), .dinb(n270), .dout(n23091));
  jand g05829(.dina(n23091), .dinb(n23090), .dout(n23092));
  jor  g05830(.dina(n23092), .dinb(n22891), .dout(n23093));
  jxor g05831(.dina(n22885), .dinb(n271), .dout(n23094));
  jand g05832(.dina(n23094), .dinb(n23093), .dout(n23095));
  jor  g05833(.dina(n23095), .dinb(n22886), .dout(n23096));
  jxor g05834(.dina(n22880), .dinb(n338), .dout(n23097));
  jand g05835(.dina(n23097), .dinb(n23096), .dout(n23098));
  jor  g05836(.dina(n23098), .dinb(n22881), .dout(n23099));
  jxor g05837(.dina(n22867), .dinb(n339), .dout(n23100));
  jand g05838(.dina(n23100), .dinb(n23099), .dout(n23101));
  jor  g05839(.dina(n23101), .dinb(n22876), .dout(n23102));
  jand g05840(.dina(n23102), .dinb(n22875), .dout(n23103));
  jor  g05841(.dina(n23103), .dinb(n22872), .dout(n23104));
  jand g05842(.dina(n23104), .dinb(n413), .dout(n23105));
  jor  g05843(.dina(n23105), .dinb(n22867), .dout(n23106));
  jnot g05844(.din(n23105), .dout(n23107));
  jxor g05845(.dina(n23100), .dinb(n23099), .dout(n23108));
  jor  g05846(.dina(n23108), .dinb(n23107), .dout(n23109));
  jand g05847(.dina(n23109), .dinb(n23106), .dout(n23110));
  jand g05848(.dina(n23107), .dinb(n22871), .dout(n23111));
  jand g05849(.dina(n23102), .dinb(n22872), .dout(n23112));
  jor  g05850(.dina(n23112), .dinb(n23111), .dout(n23113));
  jand g05851(.dina(n23113), .dinb(n275), .dout(n23114));
  jnot g05852(.din(n23113), .dout(n23115));
  jand g05853(.dina(n23115), .dinb(b31 ), .dout(n23116));
  jnot g05854(.din(n23116), .dout(n23117));
  jand g05855(.dina(n23110), .dinb(n340), .dout(n23118));
  jor  g05856(.dina(n23105), .dinb(n22880), .dout(n23119));
  jxor g05857(.dina(n23097), .dinb(n23096), .dout(n23120));
  jor  g05858(.dina(n23120), .dinb(n23107), .dout(n23121));
  jand g05859(.dina(n23121), .dinb(n23119), .dout(n23122));
  jand g05860(.dina(n23122), .dinb(n339), .dout(n23123));
  jor  g05861(.dina(n23105), .dinb(n22885), .dout(n23124));
  jxor g05862(.dina(n23094), .dinb(n23093), .dout(n23125));
  jor  g05863(.dina(n23125), .dinb(n23107), .dout(n23126));
  jand g05864(.dina(n23126), .dinb(n23124), .dout(n23127));
  jand g05865(.dina(n23127), .dinb(n338), .dout(n23128));
  jor  g05866(.dina(n23105), .dinb(n22890), .dout(n23129));
  jxor g05867(.dina(n23091), .dinb(n23090), .dout(n23130));
  jor  g05868(.dina(n23130), .dinb(n23107), .dout(n23131));
  jand g05869(.dina(n23131), .dinb(n23129), .dout(n23132));
  jand g05870(.dina(n23132), .dinb(n271), .dout(n23133));
  jor  g05871(.dina(n23105), .dinb(n22895), .dout(n23134));
  jxor g05872(.dina(n23088), .dinb(n23087), .dout(n23135));
  jor  g05873(.dina(n23135), .dinb(n23107), .dout(n23136));
  jand g05874(.dina(n23136), .dinb(n23134), .dout(n23137));
  jand g05875(.dina(n23137), .dinb(n270), .dout(n23138));
  jor  g05876(.dina(n23105), .dinb(n22900), .dout(n23139));
  jxor g05877(.dina(n23085), .dinb(n23084), .dout(n23140));
  jor  g05878(.dina(n23140), .dinb(n23107), .dout(n23141));
  jand g05879(.dina(n23141), .dinb(n23139), .dout(n23142));
  jand g05880(.dina(n23142), .dinb(n269), .dout(n23143));
  jor  g05881(.dina(n23105), .dinb(n22905), .dout(n23144));
  jxor g05882(.dina(n23082), .dinb(n23081), .dout(n23145));
  jor  g05883(.dina(n23145), .dinb(n23107), .dout(n23146));
  jand g05884(.dina(n23146), .dinb(n23144), .dout(n23147));
  jand g05885(.dina(n23147), .dinb(n274), .dout(n23148));
  jor  g05886(.dina(n23105), .dinb(n22910), .dout(n23149));
  jxor g05887(.dina(n23079), .dinb(n23078), .dout(n23150));
  jor  g05888(.dina(n23150), .dinb(n23107), .dout(n23151));
  jand g05889(.dina(n23151), .dinb(n23149), .dout(n23152));
  jand g05890(.dina(n23152), .dinb(n268), .dout(n23153));
  jor  g05891(.dina(n23105), .dinb(n22915), .dout(n23154));
  jxor g05892(.dina(n23076), .dinb(n23075), .dout(n23155));
  jor  g05893(.dina(n23155), .dinb(n23107), .dout(n23156));
  jand g05894(.dina(n23156), .dinb(n23154), .dout(n23157));
  jand g05895(.dina(n23157), .dinb(n349), .dout(n23158));
  jor  g05896(.dina(n23105), .dinb(n22920), .dout(n23159));
  jxor g05897(.dina(n23073), .dinb(n23072), .dout(n23160));
  jor  g05898(.dina(n23160), .dinb(n23107), .dout(n23161));
  jand g05899(.dina(n23161), .dinb(n23159), .dout(n23162));
  jand g05900(.dina(n23162), .dinb(n348), .dout(n23163));
  jor  g05901(.dina(n23105), .dinb(n22925), .dout(n23164));
  jxor g05902(.dina(n23070), .dinb(n23069), .dout(n23165));
  jor  g05903(.dina(n23165), .dinb(n23107), .dout(n23166));
  jand g05904(.dina(n23166), .dinb(n23164), .dout(n23167));
  jand g05905(.dina(n23167), .dinb(n347), .dout(n23168));
  jor  g05906(.dina(n23105), .dinb(n22930), .dout(n23169));
  jxor g05907(.dina(n23067), .dinb(n23066), .dout(n23170));
  jor  g05908(.dina(n23170), .dinb(n23107), .dout(n23171));
  jand g05909(.dina(n23171), .dinb(n23169), .dout(n23172));
  jand g05910(.dina(n23172), .dinb(n267), .dout(n23173));
  jor  g05911(.dina(n23105), .dinb(n22935), .dout(n23174));
  jxor g05912(.dina(n23064), .dinb(n23063), .dout(n23175));
  jor  g05913(.dina(n23175), .dinb(n23107), .dout(n23176));
  jand g05914(.dina(n23176), .dinb(n23174), .dout(n23177));
  jand g05915(.dina(n23177), .dinb(n266), .dout(n23178));
  jor  g05916(.dina(n23105), .dinb(n22940), .dout(n23179));
  jxor g05917(.dina(n23061), .dinb(n23060), .dout(n23180));
  jor  g05918(.dina(n23180), .dinb(n23107), .dout(n23181));
  jand g05919(.dina(n23181), .dinb(n23179), .dout(n23182));
  jand g05920(.dina(n23182), .dinb(n356), .dout(n23183));
  jor  g05921(.dina(n23105), .dinb(n22945), .dout(n23184));
  jxor g05922(.dina(n23058), .dinb(n23057), .dout(n23185));
  jor  g05923(.dina(n23185), .dinb(n23107), .dout(n23186));
  jand g05924(.dina(n23186), .dinb(n23184), .dout(n23187));
  jand g05925(.dina(n23187), .dinb(n355), .dout(n23188));
  jor  g05926(.dina(n23105), .dinb(n22950), .dout(n23189));
  jxor g05927(.dina(n23055), .dinb(n23054), .dout(n23190));
  jor  g05928(.dina(n23190), .dinb(n23107), .dout(n23191));
  jand g05929(.dina(n23191), .dinb(n23189), .dout(n23192));
  jand g05930(.dina(n23192), .dinb(n364), .dout(n23193));
  jor  g05931(.dina(n23105), .dinb(n22955), .dout(n23194));
  jxor g05932(.dina(n23052), .dinb(n23051), .dout(n23195));
  jor  g05933(.dina(n23195), .dinb(n23107), .dout(n23196));
  jand g05934(.dina(n23196), .dinb(n23194), .dout(n23197));
  jand g05935(.dina(n23197), .dinb(n361), .dout(n23198));
  jor  g05936(.dina(n23105), .dinb(n22960), .dout(n23199));
  jxor g05937(.dina(n23049), .dinb(n23048), .dout(n23200));
  jor  g05938(.dina(n23200), .dinb(n23107), .dout(n23201));
  jand g05939(.dina(n23201), .dinb(n23199), .dout(n23202));
  jand g05940(.dina(n23202), .dinb(n360), .dout(n23203));
  jor  g05941(.dina(n23105), .dinb(n22965), .dout(n23204));
  jxor g05942(.dina(n23046), .dinb(n23045), .dout(n23205));
  jor  g05943(.dina(n23205), .dinb(n23107), .dout(n23206));
  jand g05944(.dina(n23206), .dinb(n23204), .dout(n23207));
  jand g05945(.dina(n23207), .dinb(n363), .dout(n23208));
  jor  g05946(.dina(n23105), .dinb(n22970), .dout(n23209));
  jxor g05947(.dina(n23043), .dinb(n23042), .dout(n23210));
  jor  g05948(.dina(n23210), .dinb(n23107), .dout(n23211));
  jand g05949(.dina(n23211), .dinb(n23209), .dout(n23212));
  jand g05950(.dina(n23212), .dinb(n359), .dout(n23213));
  jor  g05951(.dina(n23105), .dinb(n22975), .dout(n23214));
  jxor g05952(.dina(n23040), .dinb(n23039), .dout(n23215));
  jor  g05953(.dina(n23215), .dinb(n23107), .dout(n23216));
  jand g05954(.dina(n23216), .dinb(n23214), .dout(n23217));
  jand g05955(.dina(n23217), .dinb(n369), .dout(n23218));
  jor  g05956(.dina(n23105), .dinb(n22980), .dout(n23219));
  jxor g05957(.dina(n23037), .dinb(n23036), .dout(n23220));
  jor  g05958(.dina(n23220), .dinb(n23107), .dout(n23221));
  jand g05959(.dina(n23221), .dinb(n23219), .dout(n23222));
  jand g05960(.dina(n23222), .dinb(n368), .dout(n23223));
  jor  g05961(.dina(n23105), .dinb(n22985), .dout(n23224));
  jxor g05962(.dina(n23034), .dinb(n23033), .dout(n23225));
  jor  g05963(.dina(n23225), .dinb(n23107), .dout(n23226));
  jand g05964(.dina(n23226), .dinb(n23224), .dout(n23227));
  jand g05965(.dina(n23227), .dinb(n367), .dout(n23228));
  jor  g05966(.dina(n23105), .dinb(n22990), .dout(n23229));
  jxor g05967(.dina(n23031), .dinb(n23030), .dout(n23230));
  jor  g05968(.dina(n23230), .dinb(n23107), .dout(n23231));
  jand g05969(.dina(n23231), .dinb(n23229), .dout(n23232));
  jand g05970(.dina(n23232), .dinb(n265), .dout(n23233));
  jor  g05971(.dina(n23105), .dinb(n22995), .dout(n23234));
  jxor g05972(.dina(n23028), .dinb(n23027), .dout(n23235));
  jor  g05973(.dina(n23235), .dinb(n23107), .dout(n23236));
  jand g05974(.dina(n23236), .dinb(n23234), .dout(n23237));
  jand g05975(.dina(n23237), .dinb(n378), .dout(n23238));
  jor  g05976(.dina(n23105), .dinb(n23000), .dout(n23239));
  jxor g05977(.dina(n23025), .dinb(n23024), .dout(n23240));
  jor  g05978(.dina(n23240), .dinb(n23107), .dout(n23241));
  jand g05979(.dina(n23241), .dinb(n23239), .dout(n23242));
  jand g05980(.dina(n23242), .dinb(n377), .dout(n23243));
  jor  g05981(.dina(n23105), .dinb(n23005), .dout(n23244));
  jxor g05982(.dina(n23022), .dinb(n23021), .dout(n23245));
  jor  g05983(.dina(n23245), .dinb(n23107), .dout(n23246));
  jand g05984(.dina(n23246), .dinb(n23244), .dout(n23247));
  jand g05985(.dina(n23247), .dinb(n376), .dout(n23248));
  jor  g05986(.dina(n23105), .dinb(n23010), .dout(n23249));
  jxor g05987(.dina(n23019), .dinb(n23018), .dout(n23250));
  jor  g05988(.dina(n23250), .dinb(n23107), .dout(n23251));
  jand g05989(.dina(n23251), .dinb(n23249), .dout(n23252));
  jand g05990(.dina(n23252), .dinb(n264), .dout(n23253));
  jor  g05991(.dina(n23105), .dinb(n23015), .dout(n23254));
  jxor g05992(.dina(n23016), .dinb(n4542), .dout(n23255));
  jand g05993(.dina(n23255), .dinb(n23105), .dout(n23256));
  jnot g05994(.din(n23256), .dout(n23257));
  jand g05995(.dina(n23257), .dinb(n23254), .dout(n23258));
  jnot g05996(.din(n23258), .dout(n23259));
  jand g05997(.dina(n23259), .dinb(n386), .dout(n23260));
  jnot g05998(.din(n4277), .dout(n23261));
  jnot g05999(.din(n22872), .dout(n23262));
  jnot g06000(.din(n22876), .dout(n23263));
  jnot g06001(.din(n22881), .dout(n23264));
  jnot g06002(.din(n22886), .dout(n23265));
  jnot g06003(.din(n22891), .dout(n23266));
  jnot g06004(.din(n22896), .dout(n23267));
  jnot g06005(.din(n22901), .dout(n23268));
  jnot g06006(.din(n22906), .dout(n23269));
  jnot g06007(.din(n22911), .dout(n23270));
  jnot g06008(.din(n22916), .dout(n23271));
  jnot g06009(.din(n22921), .dout(n23272));
  jnot g06010(.din(n22926), .dout(n23273));
  jnot g06011(.din(n22931), .dout(n23274));
  jnot g06012(.din(n22936), .dout(n23275));
  jnot g06013(.din(n22941), .dout(n23276));
  jnot g06014(.din(n22946), .dout(n23277));
  jnot g06015(.din(n22951), .dout(n23278));
  jnot g06016(.din(n22956), .dout(n23279));
  jnot g06017(.din(n22961), .dout(n23280));
  jnot g06018(.din(n22966), .dout(n23281));
  jnot g06019(.din(n22971), .dout(n23282));
  jnot g06020(.din(n22976), .dout(n23283));
  jnot g06021(.din(n22981), .dout(n23284));
  jnot g06022(.din(n22986), .dout(n23285));
  jnot g06023(.din(n22991), .dout(n23286));
  jnot g06024(.din(n22996), .dout(n23287));
  jnot g06025(.din(n23001), .dout(n23288));
  jnot g06026(.din(n23006), .dout(n23289));
  jnot g06027(.din(n23011), .dout(n23290));
  jnot g06028(.din(n23014), .dout(n23291));
  jxor g06029(.dina(n23015), .dinb(n259), .dout(n23292));
  jor  g06030(.dina(n23292), .dinb(n4541), .dout(n23293));
  jand g06031(.dina(n23293), .dinb(n23291), .dout(n23294));
  jnot g06032(.din(n23019), .dout(n23295));
  jor  g06033(.dina(n23295), .dinb(n23294), .dout(n23296));
  jand g06034(.dina(n23296), .dinb(n23290), .dout(n23297));
  jnot g06035(.din(n23022), .dout(n23298));
  jor  g06036(.dina(n23298), .dinb(n23297), .dout(n23299));
  jand g06037(.dina(n23299), .dinb(n23289), .dout(n23300));
  jnot g06038(.din(n23025), .dout(n23301));
  jor  g06039(.dina(n23301), .dinb(n23300), .dout(n23302));
  jand g06040(.dina(n23302), .dinb(n23288), .dout(n23303));
  jnot g06041(.din(n23028), .dout(n23304));
  jor  g06042(.dina(n23304), .dinb(n23303), .dout(n23305));
  jand g06043(.dina(n23305), .dinb(n23287), .dout(n23306));
  jnot g06044(.din(n23031), .dout(n23307));
  jor  g06045(.dina(n23307), .dinb(n23306), .dout(n23308));
  jand g06046(.dina(n23308), .dinb(n23286), .dout(n23309));
  jnot g06047(.din(n23034), .dout(n23310));
  jor  g06048(.dina(n23310), .dinb(n23309), .dout(n23311));
  jand g06049(.dina(n23311), .dinb(n23285), .dout(n23312));
  jnot g06050(.din(n23037), .dout(n23313));
  jor  g06051(.dina(n23313), .dinb(n23312), .dout(n23314));
  jand g06052(.dina(n23314), .dinb(n23284), .dout(n23315));
  jnot g06053(.din(n23040), .dout(n23316));
  jor  g06054(.dina(n23316), .dinb(n23315), .dout(n23317));
  jand g06055(.dina(n23317), .dinb(n23283), .dout(n23318));
  jnot g06056(.din(n23043), .dout(n23319));
  jor  g06057(.dina(n23319), .dinb(n23318), .dout(n23320));
  jand g06058(.dina(n23320), .dinb(n23282), .dout(n23321));
  jnot g06059(.din(n23046), .dout(n23322));
  jor  g06060(.dina(n23322), .dinb(n23321), .dout(n23323));
  jand g06061(.dina(n23323), .dinb(n23281), .dout(n23324));
  jnot g06062(.din(n23049), .dout(n23325));
  jor  g06063(.dina(n23325), .dinb(n23324), .dout(n23326));
  jand g06064(.dina(n23326), .dinb(n23280), .dout(n23327));
  jnot g06065(.din(n23052), .dout(n23328));
  jor  g06066(.dina(n23328), .dinb(n23327), .dout(n23329));
  jand g06067(.dina(n23329), .dinb(n23279), .dout(n23330));
  jnot g06068(.din(n23055), .dout(n23331));
  jor  g06069(.dina(n23331), .dinb(n23330), .dout(n23332));
  jand g06070(.dina(n23332), .dinb(n23278), .dout(n23333));
  jnot g06071(.din(n23058), .dout(n23334));
  jor  g06072(.dina(n23334), .dinb(n23333), .dout(n23335));
  jand g06073(.dina(n23335), .dinb(n23277), .dout(n23336));
  jnot g06074(.din(n23061), .dout(n23337));
  jor  g06075(.dina(n23337), .dinb(n23336), .dout(n23338));
  jand g06076(.dina(n23338), .dinb(n23276), .dout(n23339));
  jnot g06077(.din(n23064), .dout(n23340));
  jor  g06078(.dina(n23340), .dinb(n23339), .dout(n23341));
  jand g06079(.dina(n23341), .dinb(n23275), .dout(n23342));
  jnot g06080(.din(n23067), .dout(n23343));
  jor  g06081(.dina(n23343), .dinb(n23342), .dout(n23344));
  jand g06082(.dina(n23344), .dinb(n23274), .dout(n23345));
  jnot g06083(.din(n23070), .dout(n23346));
  jor  g06084(.dina(n23346), .dinb(n23345), .dout(n23347));
  jand g06085(.dina(n23347), .dinb(n23273), .dout(n23348));
  jnot g06086(.din(n23073), .dout(n23349));
  jor  g06087(.dina(n23349), .dinb(n23348), .dout(n23350));
  jand g06088(.dina(n23350), .dinb(n23272), .dout(n23351));
  jnot g06089(.din(n23076), .dout(n23352));
  jor  g06090(.dina(n23352), .dinb(n23351), .dout(n23353));
  jand g06091(.dina(n23353), .dinb(n23271), .dout(n23354));
  jnot g06092(.din(n23079), .dout(n23355));
  jor  g06093(.dina(n23355), .dinb(n23354), .dout(n23356));
  jand g06094(.dina(n23356), .dinb(n23270), .dout(n23357));
  jnot g06095(.din(n23082), .dout(n23358));
  jor  g06096(.dina(n23358), .dinb(n23357), .dout(n23359));
  jand g06097(.dina(n23359), .dinb(n23269), .dout(n23360));
  jnot g06098(.din(n23085), .dout(n23361));
  jor  g06099(.dina(n23361), .dinb(n23360), .dout(n23362));
  jand g06100(.dina(n23362), .dinb(n23268), .dout(n23363));
  jnot g06101(.din(n23088), .dout(n23364));
  jor  g06102(.dina(n23364), .dinb(n23363), .dout(n23365));
  jand g06103(.dina(n23365), .dinb(n23267), .dout(n23366));
  jnot g06104(.din(n23091), .dout(n23367));
  jor  g06105(.dina(n23367), .dinb(n23366), .dout(n23368));
  jand g06106(.dina(n23368), .dinb(n23266), .dout(n23369));
  jnot g06107(.din(n23094), .dout(n23370));
  jor  g06108(.dina(n23370), .dinb(n23369), .dout(n23371));
  jand g06109(.dina(n23371), .dinb(n23265), .dout(n23372));
  jnot g06110(.din(n23097), .dout(n23373));
  jor  g06111(.dina(n23373), .dinb(n23372), .dout(n23374));
  jand g06112(.dina(n23374), .dinb(n23264), .dout(n23375));
  jnot g06113(.din(n23100), .dout(n23376));
  jor  g06114(.dina(n23376), .dinb(n23375), .dout(n23377));
  jand g06115(.dina(n23377), .dinb(n23263), .dout(n23378));
  jor  g06116(.dina(n23378), .dinb(n22874), .dout(n23379));
  jand g06117(.dina(n23379), .dinb(n23262), .dout(n23380));
  jor  g06118(.dina(n23380), .dinb(n23261), .dout(n23381));
  jand g06119(.dina(n23381), .dinb(a33 ), .dout(n23382));
  jnot g06120(.din(n4789), .dout(n23383));
  jor  g06121(.dina(n23380), .dinb(n23383), .dout(n23384));
  jnot g06122(.din(n23384), .dout(n23385));
  jor  g06123(.dina(n23385), .dinb(n23382), .dout(n23386));
  jand g06124(.dina(n23386), .dinb(n259), .dout(n23387));
  jand g06125(.dina(n23104), .dinb(n4277), .dout(n23388));
  jor  g06126(.dina(n23388), .dinb(n4540), .dout(n23389));
  jand g06127(.dina(n23384), .dinb(n23389), .dout(n23390));
  jxor g06128(.dina(n23390), .dinb(b1 ), .dout(n23391));
  jand g06129(.dina(n23391), .dinb(n4797), .dout(n23392));
  jor  g06130(.dina(n23392), .dinb(n23387), .dout(n23393));
  jxor g06131(.dina(n23258), .dinb(b2 ), .dout(n23394));
  jand g06132(.dina(n23394), .dinb(n23393), .dout(n23395));
  jor  g06133(.dina(n23395), .dinb(n23260), .dout(n23396));
  jxor g06134(.dina(n23252), .dinb(n264), .dout(n23397));
  jand g06135(.dina(n23397), .dinb(n23396), .dout(n23398));
  jor  g06136(.dina(n23398), .dinb(n23253), .dout(n23399));
  jxor g06137(.dina(n23247), .dinb(n376), .dout(n23400));
  jand g06138(.dina(n23400), .dinb(n23399), .dout(n23401));
  jor  g06139(.dina(n23401), .dinb(n23248), .dout(n23402));
  jxor g06140(.dina(n23242), .dinb(n377), .dout(n23403));
  jand g06141(.dina(n23403), .dinb(n23402), .dout(n23404));
  jor  g06142(.dina(n23404), .dinb(n23243), .dout(n23405));
  jxor g06143(.dina(n23237), .dinb(n378), .dout(n23406));
  jand g06144(.dina(n23406), .dinb(n23405), .dout(n23407));
  jor  g06145(.dina(n23407), .dinb(n23238), .dout(n23408));
  jxor g06146(.dina(n23232), .dinb(n265), .dout(n23409));
  jand g06147(.dina(n23409), .dinb(n23408), .dout(n23410));
  jor  g06148(.dina(n23410), .dinb(n23233), .dout(n23411));
  jxor g06149(.dina(n23227), .dinb(n367), .dout(n23412));
  jand g06150(.dina(n23412), .dinb(n23411), .dout(n23413));
  jor  g06151(.dina(n23413), .dinb(n23228), .dout(n23414));
  jxor g06152(.dina(n23222), .dinb(n368), .dout(n23415));
  jand g06153(.dina(n23415), .dinb(n23414), .dout(n23416));
  jor  g06154(.dina(n23416), .dinb(n23223), .dout(n23417));
  jxor g06155(.dina(n23217), .dinb(n369), .dout(n23418));
  jand g06156(.dina(n23418), .dinb(n23417), .dout(n23419));
  jor  g06157(.dina(n23419), .dinb(n23218), .dout(n23420));
  jxor g06158(.dina(n23212), .dinb(n359), .dout(n23421));
  jand g06159(.dina(n23421), .dinb(n23420), .dout(n23422));
  jor  g06160(.dina(n23422), .dinb(n23213), .dout(n23423));
  jxor g06161(.dina(n23207), .dinb(n363), .dout(n23424));
  jand g06162(.dina(n23424), .dinb(n23423), .dout(n23425));
  jor  g06163(.dina(n23425), .dinb(n23208), .dout(n23426));
  jxor g06164(.dina(n23202), .dinb(n360), .dout(n23427));
  jand g06165(.dina(n23427), .dinb(n23426), .dout(n23428));
  jor  g06166(.dina(n23428), .dinb(n23203), .dout(n23429));
  jxor g06167(.dina(n23197), .dinb(n361), .dout(n23430));
  jand g06168(.dina(n23430), .dinb(n23429), .dout(n23431));
  jor  g06169(.dina(n23431), .dinb(n23198), .dout(n23432));
  jxor g06170(.dina(n23192), .dinb(n364), .dout(n23433));
  jand g06171(.dina(n23433), .dinb(n23432), .dout(n23434));
  jor  g06172(.dina(n23434), .dinb(n23193), .dout(n23435));
  jxor g06173(.dina(n23187), .dinb(n355), .dout(n23436));
  jand g06174(.dina(n23436), .dinb(n23435), .dout(n23437));
  jor  g06175(.dina(n23437), .dinb(n23188), .dout(n23438));
  jxor g06176(.dina(n23182), .dinb(n356), .dout(n23439));
  jand g06177(.dina(n23439), .dinb(n23438), .dout(n23440));
  jor  g06178(.dina(n23440), .dinb(n23183), .dout(n23441));
  jxor g06179(.dina(n23177), .dinb(n266), .dout(n23442));
  jand g06180(.dina(n23442), .dinb(n23441), .dout(n23443));
  jor  g06181(.dina(n23443), .dinb(n23178), .dout(n23444));
  jxor g06182(.dina(n23172), .dinb(n267), .dout(n23445));
  jand g06183(.dina(n23445), .dinb(n23444), .dout(n23446));
  jor  g06184(.dina(n23446), .dinb(n23173), .dout(n23447));
  jxor g06185(.dina(n23167), .dinb(n347), .dout(n23448));
  jand g06186(.dina(n23448), .dinb(n23447), .dout(n23449));
  jor  g06187(.dina(n23449), .dinb(n23168), .dout(n23450));
  jxor g06188(.dina(n23162), .dinb(n348), .dout(n23451));
  jand g06189(.dina(n23451), .dinb(n23450), .dout(n23452));
  jor  g06190(.dina(n23452), .dinb(n23163), .dout(n23453));
  jxor g06191(.dina(n23157), .dinb(n349), .dout(n23454));
  jand g06192(.dina(n23454), .dinb(n23453), .dout(n23455));
  jor  g06193(.dina(n23455), .dinb(n23158), .dout(n23456));
  jxor g06194(.dina(n23152), .dinb(n268), .dout(n23457));
  jand g06195(.dina(n23457), .dinb(n23456), .dout(n23458));
  jor  g06196(.dina(n23458), .dinb(n23153), .dout(n23459));
  jxor g06197(.dina(n23147), .dinb(n274), .dout(n23460));
  jand g06198(.dina(n23460), .dinb(n23459), .dout(n23461));
  jor  g06199(.dina(n23461), .dinb(n23148), .dout(n23462));
  jxor g06200(.dina(n23142), .dinb(n269), .dout(n23463));
  jand g06201(.dina(n23463), .dinb(n23462), .dout(n23464));
  jor  g06202(.dina(n23464), .dinb(n23143), .dout(n23465));
  jxor g06203(.dina(n23137), .dinb(n270), .dout(n23466));
  jand g06204(.dina(n23466), .dinb(n23465), .dout(n23467));
  jor  g06205(.dina(n23467), .dinb(n23138), .dout(n23468));
  jxor g06206(.dina(n23132), .dinb(n271), .dout(n23469));
  jand g06207(.dina(n23469), .dinb(n23468), .dout(n23470));
  jor  g06208(.dina(n23470), .dinb(n23133), .dout(n23471));
  jxor g06209(.dina(n23127), .dinb(n338), .dout(n23472));
  jand g06210(.dina(n23472), .dinb(n23471), .dout(n23473));
  jor  g06211(.dina(n23473), .dinb(n23128), .dout(n23474));
  jxor g06212(.dina(n23122), .dinb(n339), .dout(n23475));
  jand g06213(.dina(n23475), .dinb(n23474), .dout(n23476));
  jor  g06214(.dina(n23476), .dinb(n23123), .dout(n23477));
  jxor g06215(.dina(n23110), .dinb(n340), .dout(n23478));
  jand g06216(.dina(n23478), .dinb(n23477), .dout(n23479));
  jor  g06217(.dina(n23479), .dinb(n23118), .dout(n23480));
  jand g06218(.dina(n23480), .dinb(n23117), .dout(n23481));
  jor  g06219(.dina(n23481), .dinb(n23114), .dout(n23482));
  jand g06220(.dina(n23482), .dinb(n336), .dout(n23483));
  jor  g06221(.dina(n23483), .dinb(n23110), .dout(n23484));
  jnot g06222(.din(n23483), .dout(n23485));
  jxor g06223(.dina(n23478), .dinb(n23477), .dout(n23486));
  jor  g06224(.dina(n23486), .dinb(n23485), .dout(n23487));
  jand g06225(.dina(n23487), .dinb(n23484), .dout(n23488));
  jand g06226(.dina(n23485), .dinb(n23113), .dout(n23489));
  jand g06227(.dina(n23480), .dinb(n23114), .dout(n23490));
  jor  g06228(.dina(n23490), .dinb(n23489), .dout(n23491));
  jand g06229(.dina(n23491), .dinb(n336), .dout(n23492));
  jand g06230(.dina(n23488), .dinb(n275), .dout(n23493));
  jor  g06231(.dina(n23483), .dinb(n23122), .dout(n23494));
  jxor g06232(.dina(n23475), .dinb(n23474), .dout(n23495));
  jor  g06233(.dina(n23495), .dinb(n23485), .dout(n23496));
  jand g06234(.dina(n23496), .dinb(n23494), .dout(n23497));
  jand g06235(.dina(n23497), .dinb(n340), .dout(n23498));
  jor  g06236(.dina(n23483), .dinb(n23127), .dout(n23499));
  jxor g06237(.dina(n23472), .dinb(n23471), .dout(n23500));
  jor  g06238(.dina(n23500), .dinb(n23485), .dout(n23501));
  jand g06239(.dina(n23501), .dinb(n23499), .dout(n23502));
  jand g06240(.dina(n23502), .dinb(n339), .dout(n23503));
  jor  g06241(.dina(n23483), .dinb(n23132), .dout(n23504));
  jxor g06242(.dina(n23469), .dinb(n23468), .dout(n23505));
  jor  g06243(.dina(n23505), .dinb(n23485), .dout(n23506));
  jand g06244(.dina(n23506), .dinb(n23504), .dout(n23507));
  jand g06245(.dina(n23507), .dinb(n338), .dout(n23508));
  jor  g06246(.dina(n23483), .dinb(n23137), .dout(n23509));
  jxor g06247(.dina(n23466), .dinb(n23465), .dout(n23510));
  jor  g06248(.dina(n23510), .dinb(n23485), .dout(n23511));
  jand g06249(.dina(n23511), .dinb(n23509), .dout(n23512));
  jand g06250(.dina(n23512), .dinb(n271), .dout(n23513));
  jor  g06251(.dina(n23483), .dinb(n23142), .dout(n23514));
  jxor g06252(.dina(n23463), .dinb(n23462), .dout(n23515));
  jor  g06253(.dina(n23515), .dinb(n23485), .dout(n23516));
  jand g06254(.dina(n23516), .dinb(n23514), .dout(n23517));
  jand g06255(.dina(n23517), .dinb(n270), .dout(n23518));
  jor  g06256(.dina(n23483), .dinb(n23147), .dout(n23519));
  jxor g06257(.dina(n23460), .dinb(n23459), .dout(n23520));
  jor  g06258(.dina(n23520), .dinb(n23485), .dout(n23521));
  jand g06259(.dina(n23521), .dinb(n23519), .dout(n23522));
  jand g06260(.dina(n23522), .dinb(n269), .dout(n23523));
  jor  g06261(.dina(n23483), .dinb(n23152), .dout(n23524));
  jxor g06262(.dina(n23457), .dinb(n23456), .dout(n23525));
  jor  g06263(.dina(n23525), .dinb(n23485), .dout(n23526));
  jand g06264(.dina(n23526), .dinb(n23524), .dout(n23527));
  jand g06265(.dina(n23527), .dinb(n274), .dout(n23528));
  jor  g06266(.dina(n23483), .dinb(n23157), .dout(n23529));
  jxor g06267(.dina(n23454), .dinb(n23453), .dout(n23530));
  jor  g06268(.dina(n23530), .dinb(n23485), .dout(n23531));
  jand g06269(.dina(n23531), .dinb(n23529), .dout(n23532));
  jand g06270(.dina(n23532), .dinb(n268), .dout(n23533));
  jor  g06271(.dina(n23483), .dinb(n23162), .dout(n23534));
  jxor g06272(.dina(n23451), .dinb(n23450), .dout(n23535));
  jor  g06273(.dina(n23535), .dinb(n23485), .dout(n23536));
  jand g06274(.dina(n23536), .dinb(n23534), .dout(n23537));
  jand g06275(.dina(n23537), .dinb(n349), .dout(n23538));
  jor  g06276(.dina(n23483), .dinb(n23167), .dout(n23539));
  jxor g06277(.dina(n23448), .dinb(n23447), .dout(n23540));
  jor  g06278(.dina(n23540), .dinb(n23485), .dout(n23541));
  jand g06279(.dina(n23541), .dinb(n23539), .dout(n23542));
  jand g06280(.dina(n23542), .dinb(n348), .dout(n23543));
  jor  g06281(.dina(n23483), .dinb(n23172), .dout(n23544));
  jxor g06282(.dina(n23445), .dinb(n23444), .dout(n23545));
  jor  g06283(.dina(n23545), .dinb(n23485), .dout(n23546));
  jand g06284(.dina(n23546), .dinb(n23544), .dout(n23547));
  jand g06285(.dina(n23547), .dinb(n347), .dout(n23548));
  jor  g06286(.dina(n23483), .dinb(n23177), .dout(n23549));
  jxor g06287(.dina(n23442), .dinb(n23441), .dout(n23550));
  jor  g06288(.dina(n23550), .dinb(n23485), .dout(n23551));
  jand g06289(.dina(n23551), .dinb(n23549), .dout(n23552));
  jand g06290(.dina(n23552), .dinb(n267), .dout(n23553));
  jor  g06291(.dina(n23483), .dinb(n23182), .dout(n23554));
  jxor g06292(.dina(n23439), .dinb(n23438), .dout(n23555));
  jor  g06293(.dina(n23555), .dinb(n23485), .dout(n23556));
  jand g06294(.dina(n23556), .dinb(n23554), .dout(n23557));
  jand g06295(.dina(n23557), .dinb(n266), .dout(n23558));
  jor  g06296(.dina(n23483), .dinb(n23187), .dout(n23559));
  jxor g06297(.dina(n23436), .dinb(n23435), .dout(n23560));
  jor  g06298(.dina(n23560), .dinb(n23485), .dout(n23561));
  jand g06299(.dina(n23561), .dinb(n23559), .dout(n23562));
  jand g06300(.dina(n23562), .dinb(n356), .dout(n23563));
  jor  g06301(.dina(n23483), .dinb(n23192), .dout(n23564));
  jxor g06302(.dina(n23433), .dinb(n23432), .dout(n23565));
  jor  g06303(.dina(n23565), .dinb(n23485), .dout(n23566));
  jand g06304(.dina(n23566), .dinb(n23564), .dout(n23567));
  jand g06305(.dina(n23567), .dinb(n355), .dout(n23568));
  jor  g06306(.dina(n23483), .dinb(n23197), .dout(n23569));
  jxor g06307(.dina(n23430), .dinb(n23429), .dout(n23570));
  jor  g06308(.dina(n23570), .dinb(n23485), .dout(n23571));
  jand g06309(.dina(n23571), .dinb(n23569), .dout(n23572));
  jand g06310(.dina(n23572), .dinb(n364), .dout(n23573));
  jor  g06311(.dina(n23483), .dinb(n23202), .dout(n23574));
  jxor g06312(.dina(n23427), .dinb(n23426), .dout(n23575));
  jor  g06313(.dina(n23575), .dinb(n23485), .dout(n23576));
  jand g06314(.dina(n23576), .dinb(n23574), .dout(n23577));
  jand g06315(.dina(n23577), .dinb(n361), .dout(n23578));
  jor  g06316(.dina(n23483), .dinb(n23207), .dout(n23579));
  jxor g06317(.dina(n23424), .dinb(n23423), .dout(n23580));
  jor  g06318(.dina(n23580), .dinb(n23485), .dout(n23581));
  jand g06319(.dina(n23581), .dinb(n23579), .dout(n23582));
  jand g06320(.dina(n23582), .dinb(n360), .dout(n23583));
  jor  g06321(.dina(n23483), .dinb(n23212), .dout(n23584));
  jxor g06322(.dina(n23421), .dinb(n23420), .dout(n23585));
  jor  g06323(.dina(n23585), .dinb(n23485), .dout(n23586));
  jand g06324(.dina(n23586), .dinb(n23584), .dout(n23587));
  jand g06325(.dina(n23587), .dinb(n363), .dout(n23588));
  jor  g06326(.dina(n23483), .dinb(n23217), .dout(n23589));
  jxor g06327(.dina(n23418), .dinb(n23417), .dout(n23590));
  jor  g06328(.dina(n23590), .dinb(n23485), .dout(n23591));
  jand g06329(.dina(n23591), .dinb(n23589), .dout(n23592));
  jand g06330(.dina(n23592), .dinb(n359), .dout(n23593));
  jor  g06331(.dina(n23483), .dinb(n23222), .dout(n23594));
  jxor g06332(.dina(n23415), .dinb(n23414), .dout(n23595));
  jor  g06333(.dina(n23595), .dinb(n23485), .dout(n23596));
  jand g06334(.dina(n23596), .dinb(n23594), .dout(n23597));
  jand g06335(.dina(n23597), .dinb(n369), .dout(n23598));
  jor  g06336(.dina(n23483), .dinb(n23227), .dout(n23599));
  jxor g06337(.dina(n23412), .dinb(n23411), .dout(n23600));
  jor  g06338(.dina(n23600), .dinb(n23485), .dout(n23601));
  jand g06339(.dina(n23601), .dinb(n23599), .dout(n23602));
  jand g06340(.dina(n23602), .dinb(n368), .dout(n23603));
  jor  g06341(.dina(n23483), .dinb(n23232), .dout(n23604));
  jxor g06342(.dina(n23409), .dinb(n23408), .dout(n23605));
  jor  g06343(.dina(n23605), .dinb(n23485), .dout(n23606));
  jand g06344(.dina(n23606), .dinb(n23604), .dout(n23607));
  jand g06345(.dina(n23607), .dinb(n367), .dout(n23608));
  jor  g06346(.dina(n23483), .dinb(n23237), .dout(n23609));
  jxor g06347(.dina(n23406), .dinb(n23405), .dout(n23610));
  jor  g06348(.dina(n23610), .dinb(n23485), .dout(n23611));
  jand g06349(.dina(n23611), .dinb(n23609), .dout(n23612));
  jand g06350(.dina(n23612), .dinb(n265), .dout(n23613));
  jor  g06351(.dina(n23483), .dinb(n23242), .dout(n23614));
  jxor g06352(.dina(n23403), .dinb(n23402), .dout(n23615));
  jor  g06353(.dina(n23615), .dinb(n23485), .dout(n23616));
  jand g06354(.dina(n23616), .dinb(n23614), .dout(n23617));
  jand g06355(.dina(n23617), .dinb(n378), .dout(n23618));
  jor  g06356(.dina(n23483), .dinb(n23247), .dout(n23619));
  jxor g06357(.dina(n23400), .dinb(n23399), .dout(n23620));
  jor  g06358(.dina(n23620), .dinb(n23485), .dout(n23621));
  jand g06359(.dina(n23621), .dinb(n23619), .dout(n23622));
  jand g06360(.dina(n23622), .dinb(n377), .dout(n23623));
  jor  g06361(.dina(n23483), .dinb(n23252), .dout(n23624));
  jxor g06362(.dina(n23397), .dinb(n23396), .dout(n23625));
  jor  g06363(.dina(n23625), .dinb(n23485), .dout(n23626));
  jand g06364(.dina(n23626), .dinb(n23624), .dout(n23627));
  jand g06365(.dina(n23627), .dinb(n376), .dout(n23628));
  jor  g06366(.dina(n23483), .dinb(n23259), .dout(n23629));
  jxor g06367(.dina(n23394), .dinb(n23393), .dout(n23630));
  jor  g06368(.dina(n23630), .dinb(n23485), .dout(n23631));
  jand g06369(.dina(n23631), .dinb(n23629), .dout(n23632));
  jand g06370(.dina(n23632), .dinb(n264), .dout(n23633));
  jor  g06371(.dina(n23483), .dinb(n23390), .dout(n23634));
  jxor g06372(.dina(n23391), .dinb(n4797), .dout(n23635));
  jand g06373(.dina(n23635), .dinb(n23483), .dout(n23636));
  jnot g06374(.din(n23636), .dout(n23637));
  jand g06375(.dina(n23637), .dinb(n23634), .dout(n23638));
  jnot g06376(.din(n23638), .dout(n23639));
  jand g06377(.dina(n23639), .dinb(n386), .dout(n23640));
  jnot g06378(.din(n5043), .dout(n23641));
  jnot g06379(.din(n23114), .dout(n23642));
  jnot g06380(.din(n23118), .dout(n23643));
  jnot g06381(.din(n23123), .dout(n23644));
  jnot g06382(.din(n23128), .dout(n23645));
  jnot g06383(.din(n23133), .dout(n23646));
  jnot g06384(.din(n23138), .dout(n23647));
  jnot g06385(.din(n23143), .dout(n23648));
  jnot g06386(.din(n23148), .dout(n23649));
  jnot g06387(.din(n23153), .dout(n23650));
  jnot g06388(.din(n23158), .dout(n23651));
  jnot g06389(.din(n23163), .dout(n23652));
  jnot g06390(.din(n23168), .dout(n23653));
  jnot g06391(.din(n23173), .dout(n23654));
  jnot g06392(.din(n23178), .dout(n23655));
  jnot g06393(.din(n23183), .dout(n23656));
  jnot g06394(.din(n23188), .dout(n23657));
  jnot g06395(.din(n23193), .dout(n23658));
  jnot g06396(.din(n23198), .dout(n23659));
  jnot g06397(.din(n23203), .dout(n23660));
  jnot g06398(.din(n23208), .dout(n23661));
  jnot g06399(.din(n23213), .dout(n23662));
  jnot g06400(.din(n23218), .dout(n23663));
  jnot g06401(.din(n23223), .dout(n23664));
  jnot g06402(.din(n23228), .dout(n23665));
  jnot g06403(.din(n23233), .dout(n23666));
  jnot g06404(.din(n23238), .dout(n23667));
  jnot g06405(.din(n23243), .dout(n23668));
  jnot g06406(.din(n23248), .dout(n23669));
  jnot g06407(.din(n23253), .dout(n23670));
  jnot g06408(.din(n23260), .dout(n23671));
  jnot g06409(.din(n23387), .dout(n23672));
  jxor g06410(.dina(n23390), .dinb(n259), .dout(n23673));
  jor  g06411(.dina(n23673), .dinb(n4796), .dout(n23674));
  jand g06412(.dina(n23674), .dinb(n23672), .dout(n23675));
  jnot g06413(.din(n23394), .dout(n23676));
  jor  g06414(.dina(n23676), .dinb(n23675), .dout(n23677));
  jand g06415(.dina(n23677), .dinb(n23671), .dout(n23678));
  jnot g06416(.din(n23397), .dout(n23679));
  jor  g06417(.dina(n23679), .dinb(n23678), .dout(n23680));
  jand g06418(.dina(n23680), .dinb(n23670), .dout(n23681));
  jnot g06419(.din(n23400), .dout(n23682));
  jor  g06420(.dina(n23682), .dinb(n23681), .dout(n23683));
  jand g06421(.dina(n23683), .dinb(n23669), .dout(n23684));
  jnot g06422(.din(n23403), .dout(n23685));
  jor  g06423(.dina(n23685), .dinb(n23684), .dout(n23686));
  jand g06424(.dina(n23686), .dinb(n23668), .dout(n23687));
  jnot g06425(.din(n23406), .dout(n23688));
  jor  g06426(.dina(n23688), .dinb(n23687), .dout(n23689));
  jand g06427(.dina(n23689), .dinb(n23667), .dout(n23690));
  jnot g06428(.din(n23409), .dout(n23691));
  jor  g06429(.dina(n23691), .dinb(n23690), .dout(n23692));
  jand g06430(.dina(n23692), .dinb(n23666), .dout(n23693));
  jnot g06431(.din(n23412), .dout(n23694));
  jor  g06432(.dina(n23694), .dinb(n23693), .dout(n23695));
  jand g06433(.dina(n23695), .dinb(n23665), .dout(n23696));
  jnot g06434(.din(n23415), .dout(n23697));
  jor  g06435(.dina(n23697), .dinb(n23696), .dout(n23698));
  jand g06436(.dina(n23698), .dinb(n23664), .dout(n23699));
  jnot g06437(.din(n23418), .dout(n23700));
  jor  g06438(.dina(n23700), .dinb(n23699), .dout(n23701));
  jand g06439(.dina(n23701), .dinb(n23663), .dout(n23702));
  jnot g06440(.din(n23421), .dout(n23703));
  jor  g06441(.dina(n23703), .dinb(n23702), .dout(n23704));
  jand g06442(.dina(n23704), .dinb(n23662), .dout(n23705));
  jnot g06443(.din(n23424), .dout(n23706));
  jor  g06444(.dina(n23706), .dinb(n23705), .dout(n23707));
  jand g06445(.dina(n23707), .dinb(n23661), .dout(n23708));
  jnot g06446(.din(n23427), .dout(n23709));
  jor  g06447(.dina(n23709), .dinb(n23708), .dout(n23710));
  jand g06448(.dina(n23710), .dinb(n23660), .dout(n23711));
  jnot g06449(.din(n23430), .dout(n23712));
  jor  g06450(.dina(n23712), .dinb(n23711), .dout(n23713));
  jand g06451(.dina(n23713), .dinb(n23659), .dout(n23714));
  jnot g06452(.din(n23433), .dout(n23715));
  jor  g06453(.dina(n23715), .dinb(n23714), .dout(n23716));
  jand g06454(.dina(n23716), .dinb(n23658), .dout(n23717));
  jnot g06455(.din(n23436), .dout(n23718));
  jor  g06456(.dina(n23718), .dinb(n23717), .dout(n23719));
  jand g06457(.dina(n23719), .dinb(n23657), .dout(n23720));
  jnot g06458(.din(n23439), .dout(n23721));
  jor  g06459(.dina(n23721), .dinb(n23720), .dout(n23722));
  jand g06460(.dina(n23722), .dinb(n23656), .dout(n23723));
  jnot g06461(.din(n23442), .dout(n23724));
  jor  g06462(.dina(n23724), .dinb(n23723), .dout(n23725));
  jand g06463(.dina(n23725), .dinb(n23655), .dout(n23726));
  jnot g06464(.din(n23445), .dout(n23727));
  jor  g06465(.dina(n23727), .dinb(n23726), .dout(n23728));
  jand g06466(.dina(n23728), .dinb(n23654), .dout(n23729));
  jnot g06467(.din(n23448), .dout(n23730));
  jor  g06468(.dina(n23730), .dinb(n23729), .dout(n23731));
  jand g06469(.dina(n23731), .dinb(n23653), .dout(n23732));
  jnot g06470(.din(n23451), .dout(n23733));
  jor  g06471(.dina(n23733), .dinb(n23732), .dout(n23734));
  jand g06472(.dina(n23734), .dinb(n23652), .dout(n23735));
  jnot g06473(.din(n23454), .dout(n23736));
  jor  g06474(.dina(n23736), .dinb(n23735), .dout(n23737));
  jand g06475(.dina(n23737), .dinb(n23651), .dout(n23738));
  jnot g06476(.din(n23457), .dout(n23739));
  jor  g06477(.dina(n23739), .dinb(n23738), .dout(n23740));
  jand g06478(.dina(n23740), .dinb(n23650), .dout(n23741));
  jnot g06479(.din(n23460), .dout(n23742));
  jor  g06480(.dina(n23742), .dinb(n23741), .dout(n23743));
  jand g06481(.dina(n23743), .dinb(n23649), .dout(n23744));
  jnot g06482(.din(n23463), .dout(n23745));
  jor  g06483(.dina(n23745), .dinb(n23744), .dout(n23746));
  jand g06484(.dina(n23746), .dinb(n23648), .dout(n23747));
  jnot g06485(.din(n23466), .dout(n23748));
  jor  g06486(.dina(n23748), .dinb(n23747), .dout(n23749));
  jand g06487(.dina(n23749), .dinb(n23647), .dout(n23750));
  jnot g06488(.din(n23469), .dout(n23751));
  jor  g06489(.dina(n23751), .dinb(n23750), .dout(n23752));
  jand g06490(.dina(n23752), .dinb(n23646), .dout(n23753));
  jnot g06491(.din(n23472), .dout(n23754));
  jor  g06492(.dina(n23754), .dinb(n23753), .dout(n23755));
  jand g06493(.dina(n23755), .dinb(n23645), .dout(n23756));
  jnot g06494(.din(n23475), .dout(n23757));
  jor  g06495(.dina(n23757), .dinb(n23756), .dout(n23758));
  jand g06496(.dina(n23758), .dinb(n23644), .dout(n23759));
  jnot g06497(.din(n23478), .dout(n23760));
  jor  g06498(.dina(n23760), .dinb(n23759), .dout(n23761));
  jand g06499(.dina(n23761), .dinb(n23643), .dout(n23762));
  jor  g06500(.dina(n23762), .dinb(n23116), .dout(n23763));
  jand g06501(.dina(n23763), .dinb(n23642), .dout(n23764));
  jor  g06502(.dina(n23764), .dinb(n23641), .dout(n23765));
  jand g06503(.dina(n23765), .dinb(a32 ), .dout(n23766));
  jnot g06504(.din(n5046), .dout(n23767));
  jor  g06505(.dina(n23764), .dinb(n23767), .dout(n23768));
  jnot g06506(.din(n23768), .dout(n23769));
  jor  g06507(.dina(n23769), .dinb(n23766), .dout(n23770));
  jand g06508(.dina(n23770), .dinb(n259), .dout(n23771));
  jand g06509(.dina(n23482), .dinb(n5043), .dout(n23772));
  jor  g06510(.dina(n23772), .dinb(n4795), .dout(n23773));
  jand g06511(.dina(n23768), .dinb(n23773), .dout(n23774));
  jxor g06512(.dina(n23774), .dinb(b1 ), .dout(n23775));
  jand g06513(.dina(n23775), .dinb(n5054), .dout(n23776));
  jor  g06514(.dina(n23776), .dinb(n23771), .dout(n23777));
  jxor g06515(.dina(n23638), .dinb(b2 ), .dout(n23778));
  jand g06516(.dina(n23778), .dinb(n23777), .dout(n23779));
  jor  g06517(.dina(n23779), .dinb(n23640), .dout(n23780));
  jxor g06518(.dina(n23632), .dinb(n264), .dout(n23781));
  jand g06519(.dina(n23781), .dinb(n23780), .dout(n23782));
  jor  g06520(.dina(n23782), .dinb(n23633), .dout(n23783));
  jxor g06521(.dina(n23627), .dinb(n376), .dout(n23784));
  jand g06522(.dina(n23784), .dinb(n23783), .dout(n23785));
  jor  g06523(.dina(n23785), .dinb(n23628), .dout(n23786));
  jxor g06524(.dina(n23622), .dinb(n377), .dout(n23787));
  jand g06525(.dina(n23787), .dinb(n23786), .dout(n23788));
  jor  g06526(.dina(n23788), .dinb(n23623), .dout(n23789));
  jxor g06527(.dina(n23617), .dinb(n378), .dout(n23790));
  jand g06528(.dina(n23790), .dinb(n23789), .dout(n23791));
  jor  g06529(.dina(n23791), .dinb(n23618), .dout(n23792));
  jxor g06530(.dina(n23612), .dinb(n265), .dout(n23793));
  jand g06531(.dina(n23793), .dinb(n23792), .dout(n23794));
  jor  g06532(.dina(n23794), .dinb(n23613), .dout(n23795));
  jxor g06533(.dina(n23607), .dinb(n367), .dout(n23796));
  jand g06534(.dina(n23796), .dinb(n23795), .dout(n23797));
  jor  g06535(.dina(n23797), .dinb(n23608), .dout(n23798));
  jxor g06536(.dina(n23602), .dinb(n368), .dout(n23799));
  jand g06537(.dina(n23799), .dinb(n23798), .dout(n23800));
  jor  g06538(.dina(n23800), .dinb(n23603), .dout(n23801));
  jxor g06539(.dina(n23597), .dinb(n369), .dout(n23802));
  jand g06540(.dina(n23802), .dinb(n23801), .dout(n23803));
  jor  g06541(.dina(n23803), .dinb(n23598), .dout(n23804));
  jxor g06542(.dina(n23592), .dinb(n359), .dout(n23805));
  jand g06543(.dina(n23805), .dinb(n23804), .dout(n23806));
  jor  g06544(.dina(n23806), .dinb(n23593), .dout(n23807));
  jxor g06545(.dina(n23587), .dinb(n363), .dout(n23808));
  jand g06546(.dina(n23808), .dinb(n23807), .dout(n23809));
  jor  g06547(.dina(n23809), .dinb(n23588), .dout(n23810));
  jxor g06548(.dina(n23582), .dinb(n360), .dout(n23811));
  jand g06549(.dina(n23811), .dinb(n23810), .dout(n23812));
  jor  g06550(.dina(n23812), .dinb(n23583), .dout(n23813));
  jxor g06551(.dina(n23577), .dinb(n361), .dout(n23814));
  jand g06552(.dina(n23814), .dinb(n23813), .dout(n23815));
  jor  g06553(.dina(n23815), .dinb(n23578), .dout(n23816));
  jxor g06554(.dina(n23572), .dinb(n364), .dout(n23817));
  jand g06555(.dina(n23817), .dinb(n23816), .dout(n23818));
  jor  g06556(.dina(n23818), .dinb(n23573), .dout(n23819));
  jxor g06557(.dina(n23567), .dinb(n355), .dout(n23820));
  jand g06558(.dina(n23820), .dinb(n23819), .dout(n23821));
  jor  g06559(.dina(n23821), .dinb(n23568), .dout(n23822));
  jxor g06560(.dina(n23562), .dinb(n356), .dout(n23823));
  jand g06561(.dina(n23823), .dinb(n23822), .dout(n23824));
  jor  g06562(.dina(n23824), .dinb(n23563), .dout(n23825));
  jxor g06563(.dina(n23557), .dinb(n266), .dout(n23826));
  jand g06564(.dina(n23826), .dinb(n23825), .dout(n23827));
  jor  g06565(.dina(n23827), .dinb(n23558), .dout(n23828));
  jxor g06566(.dina(n23552), .dinb(n267), .dout(n23829));
  jand g06567(.dina(n23829), .dinb(n23828), .dout(n23830));
  jor  g06568(.dina(n23830), .dinb(n23553), .dout(n23831));
  jxor g06569(.dina(n23547), .dinb(n347), .dout(n23832));
  jand g06570(.dina(n23832), .dinb(n23831), .dout(n23833));
  jor  g06571(.dina(n23833), .dinb(n23548), .dout(n23834));
  jxor g06572(.dina(n23542), .dinb(n348), .dout(n23835));
  jand g06573(.dina(n23835), .dinb(n23834), .dout(n23836));
  jor  g06574(.dina(n23836), .dinb(n23543), .dout(n23837));
  jxor g06575(.dina(n23537), .dinb(n349), .dout(n23838));
  jand g06576(.dina(n23838), .dinb(n23837), .dout(n23839));
  jor  g06577(.dina(n23839), .dinb(n23538), .dout(n23840));
  jxor g06578(.dina(n23532), .dinb(n268), .dout(n23841));
  jand g06579(.dina(n23841), .dinb(n23840), .dout(n23842));
  jor  g06580(.dina(n23842), .dinb(n23533), .dout(n23843));
  jxor g06581(.dina(n23527), .dinb(n274), .dout(n23844));
  jand g06582(.dina(n23844), .dinb(n23843), .dout(n23845));
  jor  g06583(.dina(n23845), .dinb(n23528), .dout(n23846));
  jxor g06584(.dina(n23522), .dinb(n269), .dout(n23847));
  jand g06585(.dina(n23847), .dinb(n23846), .dout(n23848));
  jor  g06586(.dina(n23848), .dinb(n23523), .dout(n23849));
  jxor g06587(.dina(n23517), .dinb(n270), .dout(n23850));
  jand g06588(.dina(n23850), .dinb(n23849), .dout(n23851));
  jor  g06589(.dina(n23851), .dinb(n23518), .dout(n23852));
  jxor g06590(.dina(n23512), .dinb(n271), .dout(n23853));
  jand g06591(.dina(n23853), .dinb(n23852), .dout(n23854));
  jor  g06592(.dina(n23854), .dinb(n23513), .dout(n23855));
  jxor g06593(.dina(n23507), .dinb(n338), .dout(n23856));
  jand g06594(.dina(n23856), .dinb(n23855), .dout(n23857));
  jor  g06595(.dina(n23857), .dinb(n23508), .dout(n23858));
  jxor g06596(.dina(n23502), .dinb(n339), .dout(n23859));
  jand g06597(.dina(n23859), .dinb(n23858), .dout(n23860));
  jor  g06598(.dina(n23860), .dinb(n23503), .dout(n23861));
  jxor g06599(.dina(n23497), .dinb(n340), .dout(n23862));
  jand g06600(.dina(n23862), .dinb(n23861), .dout(n23863));
  jor  g06601(.dina(n23863), .dinb(n23498), .dout(n23864));
  jxor g06602(.dina(n23488), .dinb(n275), .dout(n23865));
  jand g06603(.dina(n23865), .dinb(n23864), .dout(n23866));
  jor  g06604(.dina(n23866), .dinb(n23493), .dout(n23867));
  jxor g06605(.dina(n23491), .dinb(b32 ), .dout(n23868));
  jnot g06606(.din(n23868), .dout(n23869));
  jand g06607(.dina(n23869), .dinb(n23867), .dout(n23870));
  jand g06608(.dina(n23870), .dinb(n411), .dout(n23871));
  jor  g06609(.dina(n23871), .dinb(n23492), .dout(n23872));
  jor  g06610(.dina(n23872), .dinb(n23488), .dout(n23873));
  jnot g06611(.din(n23492), .dout(n23874));
  jnot g06612(.din(n411), .dout(n23875));
  jnot g06613(.din(n23493), .dout(n23876));
  jnot g06614(.din(n23498), .dout(n23877));
  jnot g06615(.din(n23503), .dout(n23878));
  jnot g06616(.din(n23508), .dout(n23879));
  jnot g06617(.din(n23513), .dout(n23880));
  jnot g06618(.din(n23518), .dout(n23881));
  jnot g06619(.din(n23523), .dout(n23882));
  jnot g06620(.din(n23528), .dout(n23883));
  jnot g06621(.din(n23533), .dout(n23884));
  jnot g06622(.din(n23538), .dout(n23885));
  jnot g06623(.din(n23543), .dout(n23886));
  jnot g06624(.din(n23548), .dout(n23887));
  jnot g06625(.din(n23553), .dout(n23888));
  jnot g06626(.din(n23558), .dout(n23889));
  jnot g06627(.din(n23563), .dout(n23890));
  jnot g06628(.din(n23568), .dout(n23891));
  jnot g06629(.din(n23573), .dout(n23892));
  jnot g06630(.din(n23578), .dout(n23893));
  jnot g06631(.din(n23583), .dout(n23894));
  jnot g06632(.din(n23588), .dout(n23895));
  jnot g06633(.din(n23593), .dout(n23896));
  jnot g06634(.din(n23598), .dout(n23897));
  jnot g06635(.din(n23603), .dout(n23898));
  jnot g06636(.din(n23608), .dout(n23899));
  jnot g06637(.din(n23613), .dout(n23900));
  jnot g06638(.din(n23618), .dout(n23901));
  jnot g06639(.din(n23623), .dout(n23902));
  jnot g06640(.din(n23628), .dout(n23903));
  jnot g06641(.din(n23633), .dout(n23904));
  jnot g06642(.din(n23640), .dout(n23905));
  jnot g06643(.din(n23771), .dout(n23906));
  jxor g06644(.dina(n23774), .dinb(n259), .dout(n23907));
  jor  g06645(.dina(n23907), .dinb(n5053), .dout(n23908));
  jand g06646(.dina(n23908), .dinb(n23906), .dout(n23909));
  jnot g06647(.din(n23778), .dout(n23910));
  jor  g06648(.dina(n23910), .dinb(n23909), .dout(n23911));
  jand g06649(.dina(n23911), .dinb(n23905), .dout(n23912));
  jnot g06650(.din(n23781), .dout(n23913));
  jor  g06651(.dina(n23913), .dinb(n23912), .dout(n23914));
  jand g06652(.dina(n23914), .dinb(n23904), .dout(n23915));
  jnot g06653(.din(n23784), .dout(n23916));
  jor  g06654(.dina(n23916), .dinb(n23915), .dout(n23917));
  jand g06655(.dina(n23917), .dinb(n23903), .dout(n23918));
  jnot g06656(.din(n23787), .dout(n23919));
  jor  g06657(.dina(n23919), .dinb(n23918), .dout(n23920));
  jand g06658(.dina(n23920), .dinb(n23902), .dout(n23921));
  jnot g06659(.din(n23790), .dout(n23922));
  jor  g06660(.dina(n23922), .dinb(n23921), .dout(n23923));
  jand g06661(.dina(n23923), .dinb(n23901), .dout(n23924));
  jnot g06662(.din(n23793), .dout(n23925));
  jor  g06663(.dina(n23925), .dinb(n23924), .dout(n23926));
  jand g06664(.dina(n23926), .dinb(n23900), .dout(n23927));
  jnot g06665(.din(n23796), .dout(n23928));
  jor  g06666(.dina(n23928), .dinb(n23927), .dout(n23929));
  jand g06667(.dina(n23929), .dinb(n23899), .dout(n23930));
  jnot g06668(.din(n23799), .dout(n23931));
  jor  g06669(.dina(n23931), .dinb(n23930), .dout(n23932));
  jand g06670(.dina(n23932), .dinb(n23898), .dout(n23933));
  jnot g06671(.din(n23802), .dout(n23934));
  jor  g06672(.dina(n23934), .dinb(n23933), .dout(n23935));
  jand g06673(.dina(n23935), .dinb(n23897), .dout(n23936));
  jnot g06674(.din(n23805), .dout(n23937));
  jor  g06675(.dina(n23937), .dinb(n23936), .dout(n23938));
  jand g06676(.dina(n23938), .dinb(n23896), .dout(n23939));
  jnot g06677(.din(n23808), .dout(n23940));
  jor  g06678(.dina(n23940), .dinb(n23939), .dout(n23941));
  jand g06679(.dina(n23941), .dinb(n23895), .dout(n23942));
  jnot g06680(.din(n23811), .dout(n23943));
  jor  g06681(.dina(n23943), .dinb(n23942), .dout(n23944));
  jand g06682(.dina(n23944), .dinb(n23894), .dout(n23945));
  jnot g06683(.din(n23814), .dout(n23946));
  jor  g06684(.dina(n23946), .dinb(n23945), .dout(n23947));
  jand g06685(.dina(n23947), .dinb(n23893), .dout(n23948));
  jnot g06686(.din(n23817), .dout(n23949));
  jor  g06687(.dina(n23949), .dinb(n23948), .dout(n23950));
  jand g06688(.dina(n23950), .dinb(n23892), .dout(n23951));
  jnot g06689(.din(n23820), .dout(n23952));
  jor  g06690(.dina(n23952), .dinb(n23951), .dout(n23953));
  jand g06691(.dina(n23953), .dinb(n23891), .dout(n23954));
  jnot g06692(.din(n23823), .dout(n23955));
  jor  g06693(.dina(n23955), .dinb(n23954), .dout(n23956));
  jand g06694(.dina(n23956), .dinb(n23890), .dout(n23957));
  jnot g06695(.din(n23826), .dout(n23958));
  jor  g06696(.dina(n23958), .dinb(n23957), .dout(n23959));
  jand g06697(.dina(n23959), .dinb(n23889), .dout(n23960));
  jnot g06698(.din(n23829), .dout(n23961));
  jor  g06699(.dina(n23961), .dinb(n23960), .dout(n23962));
  jand g06700(.dina(n23962), .dinb(n23888), .dout(n23963));
  jnot g06701(.din(n23832), .dout(n23964));
  jor  g06702(.dina(n23964), .dinb(n23963), .dout(n23965));
  jand g06703(.dina(n23965), .dinb(n23887), .dout(n23966));
  jnot g06704(.din(n23835), .dout(n23967));
  jor  g06705(.dina(n23967), .dinb(n23966), .dout(n23968));
  jand g06706(.dina(n23968), .dinb(n23886), .dout(n23969));
  jnot g06707(.din(n23838), .dout(n23970));
  jor  g06708(.dina(n23970), .dinb(n23969), .dout(n23971));
  jand g06709(.dina(n23971), .dinb(n23885), .dout(n23972));
  jnot g06710(.din(n23841), .dout(n23973));
  jor  g06711(.dina(n23973), .dinb(n23972), .dout(n23974));
  jand g06712(.dina(n23974), .dinb(n23884), .dout(n23975));
  jnot g06713(.din(n23844), .dout(n23976));
  jor  g06714(.dina(n23976), .dinb(n23975), .dout(n23977));
  jand g06715(.dina(n23977), .dinb(n23883), .dout(n23978));
  jnot g06716(.din(n23847), .dout(n23979));
  jor  g06717(.dina(n23979), .dinb(n23978), .dout(n23980));
  jand g06718(.dina(n23980), .dinb(n23882), .dout(n23981));
  jnot g06719(.din(n23850), .dout(n23982));
  jor  g06720(.dina(n23982), .dinb(n23981), .dout(n23983));
  jand g06721(.dina(n23983), .dinb(n23881), .dout(n23984));
  jnot g06722(.din(n23853), .dout(n23985));
  jor  g06723(.dina(n23985), .dinb(n23984), .dout(n23986));
  jand g06724(.dina(n23986), .dinb(n23880), .dout(n23987));
  jnot g06725(.din(n23856), .dout(n23988));
  jor  g06726(.dina(n23988), .dinb(n23987), .dout(n23989));
  jand g06727(.dina(n23989), .dinb(n23879), .dout(n23990));
  jnot g06728(.din(n23859), .dout(n23991));
  jor  g06729(.dina(n23991), .dinb(n23990), .dout(n23992));
  jand g06730(.dina(n23992), .dinb(n23878), .dout(n23993));
  jnot g06731(.din(n23862), .dout(n23994));
  jor  g06732(.dina(n23994), .dinb(n23993), .dout(n23995));
  jand g06733(.dina(n23995), .dinb(n23877), .dout(n23996));
  jnot g06734(.din(n23865), .dout(n23997));
  jor  g06735(.dina(n23997), .dinb(n23996), .dout(n23998));
  jand g06736(.dina(n23998), .dinb(n23876), .dout(n23999));
  jor  g06737(.dina(n23868), .dinb(n23999), .dout(n24000));
  jor  g06738(.dina(n24000), .dinb(n23875), .dout(n24001));
  jand g06739(.dina(n24001), .dinb(n23874), .dout(n24002));
  jxor g06740(.dina(n23865), .dinb(n23864), .dout(n24003));
  jor  g06741(.dina(n24003), .dinb(n24002), .dout(n24004));
  jand g06742(.dina(n24004), .dinb(n23873), .dout(n24005));
  jxor g06743(.dina(n23868), .dinb(n23999), .dout(n24006));
  jor  g06744(.dina(n24006), .dinb(n24002), .dout(n24007));
  jor  g06745(.dina(n23871), .dinb(n23491), .dout(n24008));
  jand g06746(.dina(n24008), .dinb(n24007), .dout(n24009));
  jand g06747(.dina(n24009), .dinb(n332), .dout(n24010));
  jnot g06748(.din(n24009), .dout(n24011));
  jand g06749(.dina(n24011), .dinb(b33 ), .dout(n24012));
  jnot g06750(.din(n24012), .dout(n24013));
  jand g06751(.dina(n24005), .dinb(n331), .dout(n24014));
  jor  g06752(.dina(n23872), .dinb(n23497), .dout(n24015));
  jxor g06753(.dina(n23862), .dinb(n23861), .dout(n24016));
  jor  g06754(.dina(n24016), .dinb(n24002), .dout(n24017));
  jand g06755(.dina(n24017), .dinb(n24015), .dout(n24018));
  jand g06756(.dina(n24018), .dinb(n275), .dout(n24019));
  jor  g06757(.dina(n23872), .dinb(n23502), .dout(n24020));
  jxor g06758(.dina(n23859), .dinb(n23858), .dout(n24021));
  jor  g06759(.dina(n24021), .dinb(n24002), .dout(n24022));
  jand g06760(.dina(n24022), .dinb(n24020), .dout(n24023));
  jand g06761(.dina(n24023), .dinb(n340), .dout(n24024));
  jor  g06762(.dina(n23872), .dinb(n23507), .dout(n24025));
  jxor g06763(.dina(n23856), .dinb(n23855), .dout(n24026));
  jor  g06764(.dina(n24026), .dinb(n24002), .dout(n24027));
  jand g06765(.dina(n24027), .dinb(n24025), .dout(n24028));
  jand g06766(.dina(n24028), .dinb(n339), .dout(n24029));
  jor  g06767(.dina(n23872), .dinb(n23512), .dout(n24030));
  jxor g06768(.dina(n23853), .dinb(n23852), .dout(n24031));
  jor  g06769(.dina(n24031), .dinb(n24002), .dout(n24032));
  jand g06770(.dina(n24032), .dinb(n24030), .dout(n24033));
  jand g06771(.dina(n24033), .dinb(n338), .dout(n24034));
  jor  g06772(.dina(n23872), .dinb(n23517), .dout(n24035));
  jxor g06773(.dina(n23850), .dinb(n23849), .dout(n24036));
  jor  g06774(.dina(n24036), .dinb(n24002), .dout(n24037));
  jand g06775(.dina(n24037), .dinb(n24035), .dout(n24038));
  jand g06776(.dina(n24038), .dinb(n271), .dout(n24039));
  jor  g06777(.dina(n23872), .dinb(n23522), .dout(n24040));
  jxor g06778(.dina(n23847), .dinb(n23846), .dout(n24041));
  jor  g06779(.dina(n24041), .dinb(n24002), .dout(n24042));
  jand g06780(.dina(n24042), .dinb(n24040), .dout(n24043));
  jand g06781(.dina(n24043), .dinb(n270), .dout(n24044));
  jor  g06782(.dina(n23872), .dinb(n23527), .dout(n24045));
  jxor g06783(.dina(n23844), .dinb(n23843), .dout(n24046));
  jor  g06784(.dina(n24046), .dinb(n24002), .dout(n24047));
  jand g06785(.dina(n24047), .dinb(n24045), .dout(n24048));
  jand g06786(.dina(n24048), .dinb(n269), .dout(n24049));
  jor  g06787(.dina(n23872), .dinb(n23532), .dout(n24050));
  jxor g06788(.dina(n23841), .dinb(n23840), .dout(n24051));
  jor  g06789(.dina(n24051), .dinb(n24002), .dout(n24052));
  jand g06790(.dina(n24052), .dinb(n24050), .dout(n24053));
  jand g06791(.dina(n24053), .dinb(n274), .dout(n24054));
  jor  g06792(.dina(n23872), .dinb(n23537), .dout(n24055));
  jxor g06793(.dina(n23838), .dinb(n23837), .dout(n24056));
  jor  g06794(.dina(n24056), .dinb(n24002), .dout(n24057));
  jand g06795(.dina(n24057), .dinb(n24055), .dout(n24058));
  jand g06796(.dina(n24058), .dinb(n268), .dout(n24059));
  jor  g06797(.dina(n23872), .dinb(n23542), .dout(n24060));
  jxor g06798(.dina(n23835), .dinb(n23834), .dout(n24061));
  jor  g06799(.dina(n24061), .dinb(n24002), .dout(n24062));
  jand g06800(.dina(n24062), .dinb(n24060), .dout(n24063));
  jand g06801(.dina(n24063), .dinb(n349), .dout(n24064));
  jor  g06802(.dina(n23872), .dinb(n23547), .dout(n24065));
  jxor g06803(.dina(n23832), .dinb(n23831), .dout(n24066));
  jor  g06804(.dina(n24066), .dinb(n24002), .dout(n24067));
  jand g06805(.dina(n24067), .dinb(n24065), .dout(n24068));
  jand g06806(.dina(n24068), .dinb(n348), .dout(n24069));
  jor  g06807(.dina(n23872), .dinb(n23552), .dout(n24070));
  jxor g06808(.dina(n23829), .dinb(n23828), .dout(n24071));
  jor  g06809(.dina(n24071), .dinb(n24002), .dout(n24072));
  jand g06810(.dina(n24072), .dinb(n24070), .dout(n24073));
  jand g06811(.dina(n24073), .dinb(n347), .dout(n24074));
  jor  g06812(.dina(n23872), .dinb(n23557), .dout(n24075));
  jxor g06813(.dina(n23826), .dinb(n23825), .dout(n24076));
  jor  g06814(.dina(n24076), .dinb(n24002), .dout(n24077));
  jand g06815(.dina(n24077), .dinb(n24075), .dout(n24078));
  jand g06816(.dina(n24078), .dinb(n267), .dout(n24079));
  jor  g06817(.dina(n23872), .dinb(n23562), .dout(n24080));
  jxor g06818(.dina(n23823), .dinb(n23822), .dout(n24081));
  jor  g06819(.dina(n24081), .dinb(n24002), .dout(n24082));
  jand g06820(.dina(n24082), .dinb(n24080), .dout(n24083));
  jand g06821(.dina(n24083), .dinb(n266), .dout(n24084));
  jor  g06822(.dina(n23872), .dinb(n23567), .dout(n24085));
  jxor g06823(.dina(n23820), .dinb(n23819), .dout(n24086));
  jor  g06824(.dina(n24086), .dinb(n24002), .dout(n24087));
  jand g06825(.dina(n24087), .dinb(n24085), .dout(n24088));
  jand g06826(.dina(n24088), .dinb(n356), .dout(n24089));
  jor  g06827(.dina(n23872), .dinb(n23572), .dout(n24090));
  jxor g06828(.dina(n23817), .dinb(n23816), .dout(n24091));
  jor  g06829(.dina(n24091), .dinb(n24002), .dout(n24092));
  jand g06830(.dina(n24092), .dinb(n24090), .dout(n24093));
  jand g06831(.dina(n24093), .dinb(n355), .dout(n24094));
  jor  g06832(.dina(n23872), .dinb(n23577), .dout(n24095));
  jxor g06833(.dina(n23814), .dinb(n23813), .dout(n24096));
  jor  g06834(.dina(n24096), .dinb(n24002), .dout(n24097));
  jand g06835(.dina(n24097), .dinb(n24095), .dout(n24098));
  jand g06836(.dina(n24098), .dinb(n364), .dout(n24099));
  jor  g06837(.dina(n23872), .dinb(n23582), .dout(n24100));
  jxor g06838(.dina(n23811), .dinb(n23810), .dout(n24101));
  jor  g06839(.dina(n24101), .dinb(n24002), .dout(n24102));
  jand g06840(.dina(n24102), .dinb(n24100), .dout(n24103));
  jand g06841(.dina(n24103), .dinb(n361), .dout(n24104));
  jor  g06842(.dina(n23872), .dinb(n23587), .dout(n24105));
  jxor g06843(.dina(n23808), .dinb(n23807), .dout(n24106));
  jor  g06844(.dina(n24106), .dinb(n24002), .dout(n24107));
  jand g06845(.dina(n24107), .dinb(n24105), .dout(n24108));
  jand g06846(.dina(n24108), .dinb(n360), .dout(n24109));
  jor  g06847(.dina(n23872), .dinb(n23592), .dout(n24110));
  jxor g06848(.dina(n23805), .dinb(n23804), .dout(n24111));
  jor  g06849(.dina(n24111), .dinb(n24002), .dout(n24112));
  jand g06850(.dina(n24112), .dinb(n24110), .dout(n24113));
  jand g06851(.dina(n24113), .dinb(n363), .dout(n24114));
  jor  g06852(.dina(n23872), .dinb(n23597), .dout(n24115));
  jxor g06853(.dina(n23802), .dinb(n23801), .dout(n24116));
  jor  g06854(.dina(n24116), .dinb(n24002), .dout(n24117));
  jand g06855(.dina(n24117), .dinb(n24115), .dout(n24118));
  jand g06856(.dina(n24118), .dinb(n359), .dout(n24119));
  jor  g06857(.dina(n23872), .dinb(n23602), .dout(n24120));
  jxor g06858(.dina(n23799), .dinb(n23798), .dout(n24121));
  jor  g06859(.dina(n24121), .dinb(n24002), .dout(n24122));
  jand g06860(.dina(n24122), .dinb(n24120), .dout(n24123));
  jand g06861(.dina(n24123), .dinb(n369), .dout(n24124));
  jor  g06862(.dina(n23872), .dinb(n23607), .dout(n24125));
  jxor g06863(.dina(n23796), .dinb(n23795), .dout(n24126));
  jor  g06864(.dina(n24126), .dinb(n24002), .dout(n24127));
  jand g06865(.dina(n24127), .dinb(n24125), .dout(n24128));
  jand g06866(.dina(n24128), .dinb(n368), .dout(n24129));
  jor  g06867(.dina(n23872), .dinb(n23612), .dout(n24130));
  jxor g06868(.dina(n23793), .dinb(n23792), .dout(n24131));
  jor  g06869(.dina(n24131), .dinb(n24002), .dout(n24132));
  jand g06870(.dina(n24132), .dinb(n24130), .dout(n24133));
  jand g06871(.dina(n24133), .dinb(n367), .dout(n24134));
  jor  g06872(.dina(n23872), .dinb(n23617), .dout(n24135));
  jxor g06873(.dina(n23790), .dinb(n23789), .dout(n24136));
  jor  g06874(.dina(n24136), .dinb(n24002), .dout(n24137));
  jand g06875(.dina(n24137), .dinb(n24135), .dout(n24138));
  jand g06876(.dina(n24138), .dinb(n265), .dout(n24139));
  jor  g06877(.dina(n23872), .dinb(n23622), .dout(n24140));
  jxor g06878(.dina(n23787), .dinb(n23786), .dout(n24141));
  jor  g06879(.dina(n24141), .dinb(n24002), .dout(n24142));
  jand g06880(.dina(n24142), .dinb(n24140), .dout(n24143));
  jand g06881(.dina(n24143), .dinb(n378), .dout(n24144));
  jor  g06882(.dina(n23872), .dinb(n23627), .dout(n24145));
  jxor g06883(.dina(n23784), .dinb(n23783), .dout(n24146));
  jor  g06884(.dina(n24146), .dinb(n24002), .dout(n24147));
  jand g06885(.dina(n24147), .dinb(n24145), .dout(n24148));
  jand g06886(.dina(n24148), .dinb(n377), .dout(n24149));
  jor  g06887(.dina(n23872), .dinb(n23632), .dout(n24150));
  jxor g06888(.dina(n23781), .dinb(n23780), .dout(n24151));
  jor  g06889(.dina(n24151), .dinb(n24002), .dout(n24152));
  jand g06890(.dina(n24152), .dinb(n24150), .dout(n24153));
  jand g06891(.dina(n24153), .dinb(n376), .dout(n24154));
  jor  g06892(.dina(n23872), .dinb(n23639), .dout(n24155));
  jxor g06893(.dina(n23778), .dinb(n23777), .dout(n24156));
  jor  g06894(.dina(n24156), .dinb(n24002), .dout(n24157));
  jand g06895(.dina(n24157), .dinb(n24155), .dout(n24158));
  jand g06896(.dina(n24158), .dinb(n264), .dout(n24159));
  jand g06897(.dina(n23907), .dinb(n5053), .dout(n24160));
  jor  g06898(.dina(n24002), .dinb(n23776), .dout(n24161));
  jor  g06899(.dina(n24161), .dinb(n24160), .dout(n24162));
  jand g06900(.dina(n24002), .dinb(n23770), .dout(n24163));
  jnot g06901(.din(n24163), .dout(n24164));
  jand g06902(.dina(n24164), .dinb(n24162), .dout(n24165));
  jnot g06903(.din(n24165), .dout(n24166));
  jand g06904(.dina(n24166), .dinb(n386), .dout(n24167));
  jand g06905(.dina(n23872), .dinb(b0 ), .dout(n24168));
  jxor g06906(.dina(n24168), .dinb(a31 ), .dout(n24169));
  jand g06907(.dina(n24169), .dinb(n259), .dout(n24170));
  jxor g06908(.dina(n24168), .dinb(n5052), .dout(n24171));
  jxor g06909(.dina(n24171), .dinb(b1 ), .dout(n24172));
  jand g06910(.dina(n24172), .dinb(n5328), .dout(n24173));
  jor  g06911(.dina(n24173), .dinb(n24170), .dout(n24174));
  jxor g06912(.dina(n24165), .dinb(b2 ), .dout(n24175));
  jand g06913(.dina(n24175), .dinb(n24174), .dout(n24176));
  jor  g06914(.dina(n24176), .dinb(n24167), .dout(n24177));
  jxor g06915(.dina(n24158), .dinb(n264), .dout(n24178));
  jand g06916(.dina(n24178), .dinb(n24177), .dout(n24179));
  jor  g06917(.dina(n24179), .dinb(n24159), .dout(n24180));
  jxor g06918(.dina(n24153), .dinb(n376), .dout(n24181));
  jand g06919(.dina(n24181), .dinb(n24180), .dout(n24182));
  jor  g06920(.dina(n24182), .dinb(n24154), .dout(n24183));
  jxor g06921(.dina(n24148), .dinb(n377), .dout(n24184));
  jand g06922(.dina(n24184), .dinb(n24183), .dout(n24185));
  jor  g06923(.dina(n24185), .dinb(n24149), .dout(n24186));
  jxor g06924(.dina(n24143), .dinb(n378), .dout(n24187));
  jand g06925(.dina(n24187), .dinb(n24186), .dout(n24188));
  jor  g06926(.dina(n24188), .dinb(n24144), .dout(n24189));
  jxor g06927(.dina(n24138), .dinb(n265), .dout(n24190));
  jand g06928(.dina(n24190), .dinb(n24189), .dout(n24191));
  jor  g06929(.dina(n24191), .dinb(n24139), .dout(n24192));
  jxor g06930(.dina(n24133), .dinb(n367), .dout(n24193));
  jand g06931(.dina(n24193), .dinb(n24192), .dout(n24194));
  jor  g06932(.dina(n24194), .dinb(n24134), .dout(n24195));
  jxor g06933(.dina(n24128), .dinb(n368), .dout(n24196));
  jand g06934(.dina(n24196), .dinb(n24195), .dout(n24197));
  jor  g06935(.dina(n24197), .dinb(n24129), .dout(n24198));
  jxor g06936(.dina(n24123), .dinb(n369), .dout(n24199));
  jand g06937(.dina(n24199), .dinb(n24198), .dout(n24200));
  jor  g06938(.dina(n24200), .dinb(n24124), .dout(n24201));
  jxor g06939(.dina(n24118), .dinb(n359), .dout(n24202));
  jand g06940(.dina(n24202), .dinb(n24201), .dout(n24203));
  jor  g06941(.dina(n24203), .dinb(n24119), .dout(n24204));
  jxor g06942(.dina(n24113), .dinb(n363), .dout(n24205));
  jand g06943(.dina(n24205), .dinb(n24204), .dout(n24206));
  jor  g06944(.dina(n24206), .dinb(n24114), .dout(n24207));
  jxor g06945(.dina(n24108), .dinb(n360), .dout(n24208));
  jand g06946(.dina(n24208), .dinb(n24207), .dout(n24209));
  jor  g06947(.dina(n24209), .dinb(n24109), .dout(n24210));
  jxor g06948(.dina(n24103), .dinb(n361), .dout(n24211));
  jand g06949(.dina(n24211), .dinb(n24210), .dout(n24212));
  jor  g06950(.dina(n24212), .dinb(n24104), .dout(n24213));
  jxor g06951(.dina(n24098), .dinb(n364), .dout(n24214));
  jand g06952(.dina(n24214), .dinb(n24213), .dout(n24215));
  jor  g06953(.dina(n24215), .dinb(n24099), .dout(n24216));
  jxor g06954(.dina(n24093), .dinb(n355), .dout(n24217));
  jand g06955(.dina(n24217), .dinb(n24216), .dout(n24218));
  jor  g06956(.dina(n24218), .dinb(n24094), .dout(n24219));
  jxor g06957(.dina(n24088), .dinb(n356), .dout(n24220));
  jand g06958(.dina(n24220), .dinb(n24219), .dout(n24221));
  jor  g06959(.dina(n24221), .dinb(n24089), .dout(n24222));
  jxor g06960(.dina(n24083), .dinb(n266), .dout(n24223));
  jand g06961(.dina(n24223), .dinb(n24222), .dout(n24224));
  jor  g06962(.dina(n24224), .dinb(n24084), .dout(n24225));
  jxor g06963(.dina(n24078), .dinb(n267), .dout(n24226));
  jand g06964(.dina(n24226), .dinb(n24225), .dout(n24227));
  jor  g06965(.dina(n24227), .dinb(n24079), .dout(n24228));
  jxor g06966(.dina(n24073), .dinb(n347), .dout(n24229));
  jand g06967(.dina(n24229), .dinb(n24228), .dout(n24230));
  jor  g06968(.dina(n24230), .dinb(n24074), .dout(n24231));
  jxor g06969(.dina(n24068), .dinb(n348), .dout(n24232));
  jand g06970(.dina(n24232), .dinb(n24231), .dout(n24233));
  jor  g06971(.dina(n24233), .dinb(n24069), .dout(n24234));
  jxor g06972(.dina(n24063), .dinb(n349), .dout(n24235));
  jand g06973(.dina(n24235), .dinb(n24234), .dout(n24236));
  jor  g06974(.dina(n24236), .dinb(n24064), .dout(n24237));
  jxor g06975(.dina(n24058), .dinb(n268), .dout(n24238));
  jand g06976(.dina(n24238), .dinb(n24237), .dout(n24239));
  jor  g06977(.dina(n24239), .dinb(n24059), .dout(n24240));
  jxor g06978(.dina(n24053), .dinb(n274), .dout(n24241));
  jand g06979(.dina(n24241), .dinb(n24240), .dout(n24242));
  jor  g06980(.dina(n24242), .dinb(n24054), .dout(n24243));
  jxor g06981(.dina(n24048), .dinb(n269), .dout(n24244));
  jand g06982(.dina(n24244), .dinb(n24243), .dout(n24245));
  jor  g06983(.dina(n24245), .dinb(n24049), .dout(n24246));
  jxor g06984(.dina(n24043), .dinb(n270), .dout(n24247));
  jand g06985(.dina(n24247), .dinb(n24246), .dout(n24248));
  jor  g06986(.dina(n24248), .dinb(n24044), .dout(n24249));
  jxor g06987(.dina(n24038), .dinb(n271), .dout(n24250));
  jand g06988(.dina(n24250), .dinb(n24249), .dout(n24251));
  jor  g06989(.dina(n24251), .dinb(n24039), .dout(n24252));
  jxor g06990(.dina(n24033), .dinb(n338), .dout(n24253));
  jand g06991(.dina(n24253), .dinb(n24252), .dout(n24254));
  jor  g06992(.dina(n24254), .dinb(n24034), .dout(n24255));
  jxor g06993(.dina(n24028), .dinb(n339), .dout(n24256));
  jand g06994(.dina(n24256), .dinb(n24255), .dout(n24257));
  jor  g06995(.dina(n24257), .dinb(n24029), .dout(n24258));
  jxor g06996(.dina(n24023), .dinb(n340), .dout(n24259));
  jand g06997(.dina(n24259), .dinb(n24258), .dout(n24260));
  jor  g06998(.dina(n24260), .dinb(n24024), .dout(n24261));
  jxor g06999(.dina(n24018), .dinb(n275), .dout(n24262));
  jand g07000(.dina(n24262), .dinb(n24261), .dout(n24263));
  jor  g07001(.dina(n24263), .dinb(n24019), .dout(n24264));
  jxor g07002(.dina(n24005), .dinb(n331), .dout(n24265));
  jand g07003(.dina(n24265), .dinb(n24264), .dout(n24266));
  jor  g07004(.dina(n24266), .dinb(n24014), .dout(n24267));
  jand g07005(.dina(n24267), .dinb(n24013), .dout(n24268));
  jor  g07006(.dina(n24268), .dinb(n24010), .dout(n24269));
  jand g07007(.dina(n24269), .dinb(n5629), .dout(n24270));
  jor  g07008(.dina(n24270), .dinb(n24005), .dout(n24271));
  jnot g07009(.din(n24270), .dout(n24272));
  jxor g07010(.dina(n24265), .dinb(n24264), .dout(n24273));
  jor  g07011(.dina(n24273), .dinb(n24272), .dout(n24274));
  jand g07012(.dina(n24274), .dinb(n24271), .dout(n24275));
  jand g07013(.dina(n24011), .dinb(b34 ), .dout(n24276));
  jnot g07014(.din(n24276), .dout(n24277));
  jand g07015(.dina(n24267), .dinb(n5629), .dout(n24278));
  jand g07016(.dina(n24278), .dinb(n332), .dout(n24279));
  jor  g07017(.dina(n24279), .dinb(n24272), .dout(n24280));
  jand g07018(.dina(n24280), .dinb(n24009), .dout(n24281));
  jand g07019(.dina(n24281), .dinb(n333), .dout(n24282));
  jand g07020(.dina(n24275), .dinb(n332), .dout(n24283));
  jor  g07021(.dina(n24270), .dinb(n24018), .dout(n24284));
  jxor g07022(.dina(n24262), .dinb(n24261), .dout(n24285));
  jor  g07023(.dina(n24285), .dinb(n24272), .dout(n24286));
  jand g07024(.dina(n24286), .dinb(n24284), .dout(n24287));
  jand g07025(.dina(n24287), .dinb(n331), .dout(n24288));
  jor  g07026(.dina(n24270), .dinb(n24023), .dout(n24289));
  jxor g07027(.dina(n24259), .dinb(n24258), .dout(n24290));
  jor  g07028(.dina(n24290), .dinb(n24272), .dout(n24291));
  jand g07029(.dina(n24291), .dinb(n24289), .dout(n24292));
  jand g07030(.dina(n24292), .dinb(n275), .dout(n24293));
  jor  g07031(.dina(n24270), .dinb(n24028), .dout(n24294));
  jxor g07032(.dina(n24256), .dinb(n24255), .dout(n24295));
  jor  g07033(.dina(n24295), .dinb(n24272), .dout(n24296));
  jand g07034(.dina(n24296), .dinb(n24294), .dout(n24297));
  jand g07035(.dina(n24297), .dinb(n340), .dout(n24298));
  jor  g07036(.dina(n24270), .dinb(n24033), .dout(n24299));
  jxor g07037(.dina(n24253), .dinb(n24252), .dout(n24300));
  jor  g07038(.dina(n24300), .dinb(n24272), .dout(n24301));
  jand g07039(.dina(n24301), .dinb(n24299), .dout(n24302));
  jand g07040(.dina(n24302), .dinb(n339), .dout(n24303));
  jor  g07041(.dina(n24270), .dinb(n24038), .dout(n24304));
  jxor g07042(.dina(n24250), .dinb(n24249), .dout(n24305));
  jor  g07043(.dina(n24305), .dinb(n24272), .dout(n24306));
  jand g07044(.dina(n24306), .dinb(n24304), .dout(n24307));
  jand g07045(.dina(n24307), .dinb(n338), .dout(n24308));
  jor  g07046(.dina(n24270), .dinb(n24043), .dout(n24309));
  jxor g07047(.dina(n24247), .dinb(n24246), .dout(n24310));
  jor  g07048(.dina(n24310), .dinb(n24272), .dout(n24311));
  jand g07049(.dina(n24311), .dinb(n24309), .dout(n24312));
  jand g07050(.dina(n24312), .dinb(n271), .dout(n24313));
  jor  g07051(.dina(n24270), .dinb(n24048), .dout(n24314));
  jxor g07052(.dina(n24244), .dinb(n24243), .dout(n24315));
  jor  g07053(.dina(n24315), .dinb(n24272), .dout(n24316));
  jand g07054(.dina(n24316), .dinb(n24314), .dout(n24317));
  jand g07055(.dina(n24317), .dinb(n270), .dout(n24318));
  jor  g07056(.dina(n24270), .dinb(n24053), .dout(n24319));
  jxor g07057(.dina(n24241), .dinb(n24240), .dout(n24320));
  jor  g07058(.dina(n24320), .dinb(n24272), .dout(n24321));
  jand g07059(.dina(n24321), .dinb(n24319), .dout(n24322));
  jand g07060(.dina(n24322), .dinb(n269), .dout(n24323));
  jor  g07061(.dina(n24270), .dinb(n24058), .dout(n24324));
  jxor g07062(.dina(n24238), .dinb(n24237), .dout(n24325));
  jor  g07063(.dina(n24325), .dinb(n24272), .dout(n24326));
  jand g07064(.dina(n24326), .dinb(n24324), .dout(n24327));
  jand g07065(.dina(n24327), .dinb(n274), .dout(n24328));
  jor  g07066(.dina(n24270), .dinb(n24063), .dout(n24329));
  jxor g07067(.dina(n24235), .dinb(n24234), .dout(n24330));
  jor  g07068(.dina(n24330), .dinb(n24272), .dout(n24331));
  jand g07069(.dina(n24331), .dinb(n24329), .dout(n24332));
  jand g07070(.dina(n24332), .dinb(n268), .dout(n24333));
  jor  g07071(.dina(n24270), .dinb(n24068), .dout(n24334));
  jxor g07072(.dina(n24232), .dinb(n24231), .dout(n24335));
  jor  g07073(.dina(n24335), .dinb(n24272), .dout(n24336));
  jand g07074(.dina(n24336), .dinb(n24334), .dout(n24337));
  jand g07075(.dina(n24337), .dinb(n349), .dout(n24338));
  jor  g07076(.dina(n24270), .dinb(n24073), .dout(n24339));
  jxor g07077(.dina(n24229), .dinb(n24228), .dout(n24340));
  jor  g07078(.dina(n24340), .dinb(n24272), .dout(n24341));
  jand g07079(.dina(n24341), .dinb(n24339), .dout(n24342));
  jand g07080(.dina(n24342), .dinb(n348), .dout(n24343));
  jor  g07081(.dina(n24270), .dinb(n24078), .dout(n24344));
  jxor g07082(.dina(n24226), .dinb(n24225), .dout(n24345));
  jor  g07083(.dina(n24345), .dinb(n24272), .dout(n24346));
  jand g07084(.dina(n24346), .dinb(n24344), .dout(n24347));
  jand g07085(.dina(n24347), .dinb(n347), .dout(n24348));
  jor  g07086(.dina(n24270), .dinb(n24083), .dout(n24349));
  jxor g07087(.dina(n24223), .dinb(n24222), .dout(n24350));
  jor  g07088(.dina(n24350), .dinb(n24272), .dout(n24351));
  jand g07089(.dina(n24351), .dinb(n24349), .dout(n24352));
  jand g07090(.dina(n24352), .dinb(n267), .dout(n24353));
  jor  g07091(.dina(n24270), .dinb(n24088), .dout(n24354));
  jxor g07092(.dina(n24220), .dinb(n24219), .dout(n24355));
  jor  g07093(.dina(n24355), .dinb(n24272), .dout(n24356));
  jand g07094(.dina(n24356), .dinb(n24354), .dout(n24357));
  jand g07095(.dina(n24357), .dinb(n266), .dout(n24358));
  jor  g07096(.dina(n24270), .dinb(n24093), .dout(n24359));
  jxor g07097(.dina(n24217), .dinb(n24216), .dout(n24360));
  jor  g07098(.dina(n24360), .dinb(n24272), .dout(n24361));
  jand g07099(.dina(n24361), .dinb(n24359), .dout(n24362));
  jand g07100(.dina(n24362), .dinb(n356), .dout(n24363));
  jor  g07101(.dina(n24270), .dinb(n24098), .dout(n24364));
  jxor g07102(.dina(n24214), .dinb(n24213), .dout(n24365));
  jor  g07103(.dina(n24365), .dinb(n24272), .dout(n24366));
  jand g07104(.dina(n24366), .dinb(n24364), .dout(n24367));
  jand g07105(.dina(n24367), .dinb(n355), .dout(n24368));
  jor  g07106(.dina(n24270), .dinb(n24103), .dout(n24369));
  jxor g07107(.dina(n24211), .dinb(n24210), .dout(n24370));
  jor  g07108(.dina(n24370), .dinb(n24272), .dout(n24371));
  jand g07109(.dina(n24371), .dinb(n24369), .dout(n24372));
  jand g07110(.dina(n24372), .dinb(n364), .dout(n24373));
  jor  g07111(.dina(n24270), .dinb(n24108), .dout(n24374));
  jxor g07112(.dina(n24208), .dinb(n24207), .dout(n24375));
  jor  g07113(.dina(n24375), .dinb(n24272), .dout(n24376));
  jand g07114(.dina(n24376), .dinb(n24374), .dout(n24377));
  jand g07115(.dina(n24377), .dinb(n361), .dout(n24378));
  jor  g07116(.dina(n24270), .dinb(n24113), .dout(n24379));
  jxor g07117(.dina(n24205), .dinb(n24204), .dout(n24380));
  jor  g07118(.dina(n24380), .dinb(n24272), .dout(n24381));
  jand g07119(.dina(n24381), .dinb(n24379), .dout(n24382));
  jand g07120(.dina(n24382), .dinb(n360), .dout(n24383));
  jor  g07121(.dina(n24270), .dinb(n24118), .dout(n24384));
  jxor g07122(.dina(n24202), .dinb(n24201), .dout(n24385));
  jor  g07123(.dina(n24385), .dinb(n24272), .dout(n24386));
  jand g07124(.dina(n24386), .dinb(n24384), .dout(n24387));
  jand g07125(.dina(n24387), .dinb(n363), .dout(n24388));
  jor  g07126(.dina(n24270), .dinb(n24123), .dout(n24389));
  jxor g07127(.dina(n24199), .dinb(n24198), .dout(n24390));
  jor  g07128(.dina(n24390), .dinb(n24272), .dout(n24391));
  jand g07129(.dina(n24391), .dinb(n24389), .dout(n24392));
  jand g07130(.dina(n24392), .dinb(n359), .dout(n24393));
  jor  g07131(.dina(n24270), .dinb(n24128), .dout(n24394));
  jxor g07132(.dina(n24196), .dinb(n24195), .dout(n24395));
  jor  g07133(.dina(n24395), .dinb(n24272), .dout(n24396));
  jand g07134(.dina(n24396), .dinb(n24394), .dout(n24397));
  jand g07135(.dina(n24397), .dinb(n369), .dout(n24398));
  jor  g07136(.dina(n24270), .dinb(n24133), .dout(n24399));
  jxor g07137(.dina(n24193), .dinb(n24192), .dout(n24400));
  jor  g07138(.dina(n24400), .dinb(n24272), .dout(n24401));
  jand g07139(.dina(n24401), .dinb(n24399), .dout(n24402));
  jand g07140(.dina(n24402), .dinb(n368), .dout(n24403));
  jor  g07141(.dina(n24270), .dinb(n24138), .dout(n24404));
  jxor g07142(.dina(n24190), .dinb(n24189), .dout(n24405));
  jor  g07143(.dina(n24405), .dinb(n24272), .dout(n24406));
  jand g07144(.dina(n24406), .dinb(n24404), .dout(n24407));
  jand g07145(.dina(n24407), .dinb(n367), .dout(n24408));
  jor  g07146(.dina(n24270), .dinb(n24143), .dout(n24409));
  jxor g07147(.dina(n24187), .dinb(n24186), .dout(n24410));
  jor  g07148(.dina(n24410), .dinb(n24272), .dout(n24411));
  jand g07149(.dina(n24411), .dinb(n24409), .dout(n24412));
  jand g07150(.dina(n24412), .dinb(n265), .dout(n24413));
  jor  g07151(.dina(n24270), .dinb(n24148), .dout(n24414));
  jxor g07152(.dina(n24184), .dinb(n24183), .dout(n24415));
  jor  g07153(.dina(n24415), .dinb(n24272), .dout(n24416));
  jand g07154(.dina(n24416), .dinb(n24414), .dout(n24417));
  jand g07155(.dina(n24417), .dinb(n378), .dout(n24418));
  jor  g07156(.dina(n24270), .dinb(n24153), .dout(n24419));
  jxor g07157(.dina(n24181), .dinb(n24180), .dout(n24420));
  jor  g07158(.dina(n24420), .dinb(n24272), .dout(n24421));
  jand g07159(.dina(n24421), .dinb(n24419), .dout(n24422));
  jand g07160(.dina(n24422), .dinb(n377), .dout(n24423));
  jor  g07161(.dina(n24270), .dinb(n24158), .dout(n24424));
  jxor g07162(.dina(n24178), .dinb(n24177), .dout(n24425));
  jor  g07163(.dina(n24425), .dinb(n24272), .dout(n24426));
  jand g07164(.dina(n24426), .dinb(n24424), .dout(n24427));
  jand g07165(.dina(n24427), .dinb(n376), .dout(n24428));
  jor  g07166(.dina(n24270), .dinb(n24166), .dout(n24429));
  jxor g07167(.dina(n24175), .dinb(n24174), .dout(n24430));
  jor  g07168(.dina(n24430), .dinb(n24272), .dout(n24431));
  jand g07169(.dina(n24431), .dinb(n24429), .dout(n24432));
  jand g07170(.dina(n24432), .dinb(n264), .dout(n24433));
  jor  g07171(.dina(n24270), .dinb(n24171), .dout(n24434));
  jxor g07172(.dina(n24172), .dinb(n5328), .dout(n24435));
  jand g07173(.dina(n24435), .dinb(n24270), .dout(n24436));
  jnot g07174(.din(n24436), .dout(n24437));
  jand g07175(.dina(n24437), .dinb(n24434), .dout(n24438));
  jor  g07176(.dina(n24438), .dinb(b2 ), .dout(n24439));
  jnot g07177(.din(n24439), .dout(n24440));
  jnot g07178(.din(n5630), .dout(n24441));
  jnot g07179(.din(n24010), .dout(n24442));
  jnot g07180(.din(n24014), .dout(n24443));
  jnot g07181(.din(n24019), .dout(n24444));
  jnot g07182(.din(n24024), .dout(n24445));
  jnot g07183(.din(n24029), .dout(n24446));
  jnot g07184(.din(n24034), .dout(n24447));
  jnot g07185(.din(n24039), .dout(n24448));
  jnot g07186(.din(n24044), .dout(n24449));
  jnot g07187(.din(n24049), .dout(n24450));
  jnot g07188(.din(n24054), .dout(n24451));
  jnot g07189(.din(n24059), .dout(n24452));
  jnot g07190(.din(n24064), .dout(n24453));
  jnot g07191(.din(n24069), .dout(n24454));
  jnot g07192(.din(n24074), .dout(n24455));
  jnot g07193(.din(n24079), .dout(n24456));
  jnot g07194(.din(n24084), .dout(n24457));
  jnot g07195(.din(n24089), .dout(n24458));
  jnot g07196(.din(n24094), .dout(n24459));
  jnot g07197(.din(n24099), .dout(n24460));
  jnot g07198(.din(n24104), .dout(n24461));
  jnot g07199(.din(n24109), .dout(n24462));
  jnot g07200(.din(n24114), .dout(n24463));
  jnot g07201(.din(n24119), .dout(n24464));
  jnot g07202(.din(n24124), .dout(n24465));
  jnot g07203(.din(n24129), .dout(n24466));
  jnot g07204(.din(n24134), .dout(n24467));
  jnot g07205(.din(n24139), .dout(n24468));
  jnot g07206(.din(n24144), .dout(n24469));
  jnot g07207(.din(n24149), .dout(n24470));
  jnot g07208(.din(n24154), .dout(n24471));
  jnot g07209(.din(n24159), .dout(n24472));
  jnot g07210(.din(n24167), .dout(n24473));
  jnot g07211(.din(n24170), .dout(n24474));
  jxor g07212(.dina(n24171), .dinb(n259), .dout(n24475));
  jor  g07213(.dina(n24475), .dinb(n5327), .dout(n24476));
  jand g07214(.dina(n24476), .dinb(n24474), .dout(n24477));
  jnot g07215(.din(n24175), .dout(n24478));
  jor  g07216(.dina(n24478), .dinb(n24477), .dout(n24479));
  jand g07217(.dina(n24479), .dinb(n24473), .dout(n24480));
  jnot g07218(.din(n24178), .dout(n24481));
  jor  g07219(.dina(n24481), .dinb(n24480), .dout(n24482));
  jand g07220(.dina(n24482), .dinb(n24472), .dout(n24483));
  jnot g07221(.din(n24181), .dout(n24484));
  jor  g07222(.dina(n24484), .dinb(n24483), .dout(n24485));
  jand g07223(.dina(n24485), .dinb(n24471), .dout(n24486));
  jnot g07224(.din(n24184), .dout(n24487));
  jor  g07225(.dina(n24487), .dinb(n24486), .dout(n24488));
  jand g07226(.dina(n24488), .dinb(n24470), .dout(n24489));
  jnot g07227(.din(n24187), .dout(n24490));
  jor  g07228(.dina(n24490), .dinb(n24489), .dout(n24491));
  jand g07229(.dina(n24491), .dinb(n24469), .dout(n24492));
  jnot g07230(.din(n24190), .dout(n24493));
  jor  g07231(.dina(n24493), .dinb(n24492), .dout(n24494));
  jand g07232(.dina(n24494), .dinb(n24468), .dout(n24495));
  jnot g07233(.din(n24193), .dout(n24496));
  jor  g07234(.dina(n24496), .dinb(n24495), .dout(n24497));
  jand g07235(.dina(n24497), .dinb(n24467), .dout(n24498));
  jnot g07236(.din(n24196), .dout(n24499));
  jor  g07237(.dina(n24499), .dinb(n24498), .dout(n24500));
  jand g07238(.dina(n24500), .dinb(n24466), .dout(n24501));
  jnot g07239(.din(n24199), .dout(n24502));
  jor  g07240(.dina(n24502), .dinb(n24501), .dout(n24503));
  jand g07241(.dina(n24503), .dinb(n24465), .dout(n24504));
  jnot g07242(.din(n24202), .dout(n24505));
  jor  g07243(.dina(n24505), .dinb(n24504), .dout(n24506));
  jand g07244(.dina(n24506), .dinb(n24464), .dout(n24507));
  jnot g07245(.din(n24205), .dout(n24508));
  jor  g07246(.dina(n24508), .dinb(n24507), .dout(n24509));
  jand g07247(.dina(n24509), .dinb(n24463), .dout(n24510));
  jnot g07248(.din(n24208), .dout(n24511));
  jor  g07249(.dina(n24511), .dinb(n24510), .dout(n24512));
  jand g07250(.dina(n24512), .dinb(n24462), .dout(n24513));
  jnot g07251(.din(n24211), .dout(n24514));
  jor  g07252(.dina(n24514), .dinb(n24513), .dout(n24515));
  jand g07253(.dina(n24515), .dinb(n24461), .dout(n24516));
  jnot g07254(.din(n24214), .dout(n24517));
  jor  g07255(.dina(n24517), .dinb(n24516), .dout(n24518));
  jand g07256(.dina(n24518), .dinb(n24460), .dout(n24519));
  jnot g07257(.din(n24217), .dout(n24520));
  jor  g07258(.dina(n24520), .dinb(n24519), .dout(n24521));
  jand g07259(.dina(n24521), .dinb(n24459), .dout(n24522));
  jnot g07260(.din(n24220), .dout(n24523));
  jor  g07261(.dina(n24523), .dinb(n24522), .dout(n24524));
  jand g07262(.dina(n24524), .dinb(n24458), .dout(n24525));
  jnot g07263(.din(n24223), .dout(n24526));
  jor  g07264(.dina(n24526), .dinb(n24525), .dout(n24527));
  jand g07265(.dina(n24527), .dinb(n24457), .dout(n24528));
  jnot g07266(.din(n24226), .dout(n24529));
  jor  g07267(.dina(n24529), .dinb(n24528), .dout(n24530));
  jand g07268(.dina(n24530), .dinb(n24456), .dout(n24531));
  jnot g07269(.din(n24229), .dout(n24532));
  jor  g07270(.dina(n24532), .dinb(n24531), .dout(n24533));
  jand g07271(.dina(n24533), .dinb(n24455), .dout(n24534));
  jnot g07272(.din(n24232), .dout(n24535));
  jor  g07273(.dina(n24535), .dinb(n24534), .dout(n24536));
  jand g07274(.dina(n24536), .dinb(n24454), .dout(n24537));
  jnot g07275(.din(n24235), .dout(n24538));
  jor  g07276(.dina(n24538), .dinb(n24537), .dout(n24539));
  jand g07277(.dina(n24539), .dinb(n24453), .dout(n24540));
  jnot g07278(.din(n24238), .dout(n24541));
  jor  g07279(.dina(n24541), .dinb(n24540), .dout(n24542));
  jand g07280(.dina(n24542), .dinb(n24452), .dout(n24543));
  jnot g07281(.din(n24241), .dout(n24544));
  jor  g07282(.dina(n24544), .dinb(n24543), .dout(n24545));
  jand g07283(.dina(n24545), .dinb(n24451), .dout(n24546));
  jnot g07284(.din(n24244), .dout(n24547));
  jor  g07285(.dina(n24547), .dinb(n24546), .dout(n24548));
  jand g07286(.dina(n24548), .dinb(n24450), .dout(n24549));
  jnot g07287(.din(n24247), .dout(n24550));
  jor  g07288(.dina(n24550), .dinb(n24549), .dout(n24551));
  jand g07289(.dina(n24551), .dinb(n24449), .dout(n24552));
  jnot g07290(.din(n24250), .dout(n24553));
  jor  g07291(.dina(n24553), .dinb(n24552), .dout(n24554));
  jand g07292(.dina(n24554), .dinb(n24448), .dout(n24555));
  jnot g07293(.din(n24253), .dout(n24556));
  jor  g07294(.dina(n24556), .dinb(n24555), .dout(n24557));
  jand g07295(.dina(n24557), .dinb(n24447), .dout(n24558));
  jnot g07296(.din(n24256), .dout(n24559));
  jor  g07297(.dina(n24559), .dinb(n24558), .dout(n24560));
  jand g07298(.dina(n24560), .dinb(n24446), .dout(n24561));
  jnot g07299(.din(n24259), .dout(n24562));
  jor  g07300(.dina(n24562), .dinb(n24561), .dout(n24563));
  jand g07301(.dina(n24563), .dinb(n24445), .dout(n24564));
  jnot g07302(.din(n24262), .dout(n24565));
  jor  g07303(.dina(n24565), .dinb(n24564), .dout(n24566));
  jand g07304(.dina(n24566), .dinb(n24444), .dout(n24567));
  jnot g07305(.din(n24265), .dout(n24568));
  jor  g07306(.dina(n24568), .dinb(n24567), .dout(n24569));
  jand g07307(.dina(n24569), .dinb(n24443), .dout(n24570));
  jor  g07308(.dina(n24570), .dinb(n24012), .dout(n24571));
  jand g07309(.dina(n24571), .dinb(n24442), .dout(n24572));
  jor  g07310(.dina(n24572), .dinb(n24441), .dout(n24573));
  jand g07311(.dina(n24573), .dinb(a30 ), .dout(n24574));
  jnot g07312(.din(n5633), .dout(n24575));
  jor  g07313(.dina(n24572), .dinb(n24575), .dout(n24576));
  jnot g07314(.din(n24576), .dout(n24577));
  jor  g07315(.dina(n24577), .dinb(n24574), .dout(n24578));
  jand g07316(.dina(n24578), .dinb(n259), .dout(n24579));
  jand g07317(.dina(n24269), .dinb(n5630), .dout(n24580));
  jor  g07318(.dina(n24580), .dinb(n5326), .dout(n24581));
  jand g07319(.dina(n24576), .dinb(n24581), .dout(n24582));
  jxor g07320(.dina(n24582), .dinb(b1 ), .dout(n24583));
  jand g07321(.dina(n24583), .dinb(n5777), .dout(n24584));
  jor  g07322(.dina(n24584), .dinb(n24579), .dout(n24585));
  jxor g07323(.dina(n24438), .dinb(b2 ), .dout(n24586));
  jand g07324(.dina(n24586), .dinb(n24585), .dout(n24587));
  jor  g07325(.dina(n24587), .dinb(n24440), .dout(n24588));
  jxor g07326(.dina(n24432), .dinb(n264), .dout(n24589));
  jand g07327(.dina(n24589), .dinb(n24588), .dout(n24590));
  jor  g07328(.dina(n24590), .dinb(n24433), .dout(n24591));
  jxor g07329(.dina(n24427), .dinb(n376), .dout(n24592));
  jand g07330(.dina(n24592), .dinb(n24591), .dout(n24593));
  jor  g07331(.dina(n24593), .dinb(n24428), .dout(n24594));
  jxor g07332(.dina(n24422), .dinb(n377), .dout(n24595));
  jand g07333(.dina(n24595), .dinb(n24594), .dout(n24596));
  jor  g07334(.dina(n24596), .dinb(n24423), .dout(n24597));
  jxor g07335(.dina(n24417), .dinb(n378), .dout(n24598));
  jand g07336(.dina(n24598), .dinb(n24597), .dout(n24599));
  jor  g07337(.dina(n24599), .dinb(n24418), .dout(n24600));
  jxor g07338(.dina(n24412), .dinb(n265), .dout(n24601));
  jand g07339(.dina(n24601), .dinb(n24600), .dout(n24602));
  jor  g07340(.dina(n24602), .dinb(n24413), .dout(n24603));
  jxor g07341(.dina(n24407), .dinb(n367), .dout(n24604));
  jand g07342(.dina(n24604), .dinb(n24603), .dout(n24605));
  jor  g07343(.dina(n24605), .dinb(n24408), .dout(n24606));
  jxor g07344(.dina(n24402), .dinb(n368), .dout(n24607));
  jand g07345(.dina(n24607), .dinb(n24606), .dout(n24608));
  jor  g07346(.dina(n24608), .dinb(n24403), .dout(n24609));
  jxor g07347(.dina(n24397), .dinb(n369), .dout(n24610));
  jand g07348(.dina(n24610), .dinb(n24609), .dout(n24611));
  jor  g07349(.dina(n24611), .dinb(n24398), .dout(n24612));
  jxor g07350(.dina(n24392), .dinb(n359), .dout(n24613));
  jand g07351(.dina(n24613), .dinb(n24612), .dout(n24614));
  jor  g07352(.dina(n24614), .dinb(n24393), .dout(n24615));
  jxor g07353(.dina(n24387), .dinb(n363), .dout(n24616));
  jand g07354(.dina(n24616), .dinb(n24615), .dout(n24617));
  jor  g07355(.dina(n24617), .dinb(n24388), .dout(n24618));
  jxor g07356(.dina(n24382), .dinb(n360), .dout(n24619));
  jand g07357(.dina(n24619), .dinb(n24618), .dout(n24620));
  jor  g07358(.dina(n24620), .dinb(n24383), .dout(n24621));
  jxor g07359(.dina(n24377), .dinb(n361), .dout(n24622));
  jand g07360(.dina(n24622), .dinb(n24621), .dout(n24623));
  jor  g07361(.dina(n24623), .dinb(n24378), .dout(n24624));
  jxor g07362(.dina(n24372), .dinb(n364), .dout(n24625));
  jand g07363(.dina(n24625), .dinb(n24624), .dout(n24626));
  jor  g07364(.dina(n24626), .dinb(n24373), .dout(n24627));
  jxor g07365(.dina(n24367), .dinb(n355), .dout(n24628));
  jand g07366(.dina(n24628), .dinb(n24627), .dout(n24629));
  jor  g07367(.dina(n24629), .dinb(n24368), .dout(n24630));
  jxor g07368(.dina(n24362), .dinb(n356), .dout(n24631));
  jand g07369(.dina(n24631), .dinb(n24630), .dout(n24632));
  jor  g07370(.dina(n24632), .dinb(n24363), .dout(n24633));
  jxor g07371(.dina(n24357), .dinb(n266), .dout(n24634));
  jand g07372(.dina(n24634), .dinb(n24633), .dout(n24635));
  jor  g07373(.dina(n24635), .dinb(n24358), .dout(n24636));
  jxor g07374(.dina(n24352), .dinb(n267), .dout(n24637));
  jand g07375(.dina(n24637), .dinb(n24636), .dout(n24638));
  jor  g07376(.dina(n24638), .dinb(n24353), .dout(n24639));
  jxor g07377(.dina(n24347), .dinb(n347), .dout(n24640));
  jand g07378(.dina(n24640), .dinb(n24639), .dout(n24641));
  jor  g07379(.dina(n24641), .dinb(n24348), .dout(n24642));
  jxor g07380(.dina(n24342), .dinb(n348), .dout(n24643));
  jand g07381(.dina(n24643), .dinb(n24642), .dout(n24644));
  jor  g07382(.dina(n24644), .dinb(n24343), .dout(n24645));
  jxor g07383(.dina(n24337), .dinb(n349), .dout(n24646));
  jand g07384(.dina(n24646), .dinb(n24645), .dout(n24647));
  jor  g07385(.dina(n24647), .dinb(n24338), .dout(n24648));
  jxor g07386(.dina(n24332), .dinb(n268), .dout(n24649));
  jand g07387(.dina(n24649), .dinb(n24648), .dout(n24650));
  jor  g07388(.dina(n24650), .dinb(n24333), .dout(n24651));
  jxor g07389(.dina(n24327), .dinb(n274), .dout(n24652));
  jand g07390(.dina(n24652), .dinb(n24651), .dout(n24653));
  jor  g07391(.dina(n24653), .dinb(n24328), .dout(n24654));
  jxor g07392(.dina(n24322), .dinb(n269), .dout(n24655));
  jand g07393(.dina(n24655), .dinb(n24654), .dout(n24656));
  jor  g07394(.dina(n24656), .dinb(n24323), .dout(n24657));
  jxor g07395(.dina(n24317), .dinb(n270), .dout(n24658));
  jand g07396(.dina(n24658), .dinb(n24657), .dout(n24659));
  jor  g07397(.dina(n24659), .dinb(n24318), .dout(n24660));
  jxor g07398(.dina(n24312), .dinb(n271), .dout(n24661));
  jand g07399(.dina(n24661), .dinb(n24660), .dout(n24662));
  jor  g07400(.dina(n24662), .dinb(n24313), .dout(n24663));
  jxor g07401(.dina(n24307), .dinb(n338), .dout(n24664));
  jand g07402(.dina(n24664), .dinb(n24663), .dout(n24665));
  jor  g07403(.dina(n24665), .dinb(n24308), .dout(n24666));
  jxor g07404(.dina(n24302), .dinb(n339), .dout(n24667));
  jand g07405(.dina(n24667), .dinb(n24666), .dout(n24668));
  jor  g07406(.dina(n24668), .dinb(n24303), .dout(n24669));
  jxor g07407(.dina(n24297), .dinb(n340), .dout(n24670));
  jand g07408(.dina(n24670), .dinb(n24669), .dout(n24671));
  jor  g07409(.dina(n24671), .dinb(n24298), .dout(n24672));
  jxor g07410(.dina(n24292), .dinb(n275), .dout(n24673));
  jand g07411(.dina(n24673), .dinb(n24672), .dout(n24674));
  jor  g07412(.dina(n24674), .dinb(n24293), .dout(n24675));
  jxor g07413(.dina(n24287), .dinb(n331), .dout(n24676));
  jand g07414(.dina(n24676), .dinb(n24675), .dout(n24677));
  jor  g07415(.dina(n24677), .dinb(n24288), .dout(n24678));
  jxor g07416(.dina(n24275), .dinb(n332), .dout(n24679));
  jand g07417(.dina(n24679), .dinb(n24678), .dout(n24680));
  jor  g07418(.dina(n24680), .dinb(n24283), .dout(n24681));
  jor  g07419(.dina(n24681), .dinb(n24282), .dout(n24682));
  jand g07420(.dina(n24682), .dinb(n24277), .dout(n24683));
  jand g07421(.dina(n24683), .dinb(n410), .dout(n24684));
  jor  g07422(.dina(n24684), .dinb(n24275), .dout(n24685));
  jnot g07423(.din(n24282), .dout(n24686));
  jnot g07424(.din(n24283), .dout(n24687));
  jnot g07425(.din(n24288), .dout(n24688));
  jnot g07426(.din(n24293), .dout(n24689));
  jnot g07427(.din(n24298), .dout(n24690));
  jnot g07428(.din(n24303), .dout(n24691));
  jnot g07429(.din(n24308), .dout(n24692));
  jnot g07430(.din(n24313), .dout(n24693));
  jnot g07431(.din(n24318), .dout(n24694));
  jnot g07432(.din(n24323), .dout(n24695));
  jnot g07433(.din(n24328), .dout(n24696));
  jnot g07434(.din(n24333), .dout(n24697));
  jnot g07435(.din(n24338), .dout(n24698));
  jnot g07436(.din(n24343), .dout(n24699));
  jnot g07437(.din(n24348), .dout(n24700));
  jnot g07438(.din(n24353), .dout(n24701));
  jnot g07439(.din(n24358), .dout(n24702));
  jnot g07440(.din(n24363), .dout(n24703));
  jnot g07441(.din(n24368), .dout(n24704));
  jnot g07442(.din(n24373), .dout(n24705));
  jnot g07443(.din(n24378), .dout(n24706));
  jnot g07444(.din(n24383), .dout(n24707));
  jnot g07445(.din(n24388), .dout(n24708));
  jnot g07446(.din(n24393), .dout(n24709));
  jnot g07447(.din(n24398), .dout(n24710));
  jnot g07448(.din(n24403), .dout(n24711));
  jnot g07449(.din(n24408), .dout(n24712));
  jnot g07450(.din(n24413), .dout(n24713));
  jnot g07451(.din(n24418), .dout(n24714));
  jnot g07452(.din(n24423), .dout(n24715));
  jnot g07453(.din(n24428), .dout(n24716));
  jnot g07454(.din(n24433), .dout(n24717));
  jor  g07455(.dina(n24582), .dinb(b1 ), .dout(n24718));
  jxor g07456(.dina(n24582), .dinb(n259), .dout(n24719));
  jor  g07457(.dina(n24719), .dinb(n5639), .dout(n24720));
  jand g07458(.dina(n24720), .dinb(n24718), .dout(n24721));
  jxor g07459(.dina(n24438), .dinb(n386), .dout(n24722));
  jor  g07460(.dina(n24722), .dinb(n24721), .dout(n24723));
  jand g07461(.dina(n24723), .dinb(n24439), .dout(n24724));
  jnot g07462(.din(n24589), .dout(n24725));
  jor  g07463(.dina(n24725), .dinb(n24724), .dout(n24726));
  jand g07464(.dina(n24726), .dinb(n24717), .dout(n24727));
  jnot g07465(.din(n24592), .dout(n24728));
  jor  g07466(.dina(n24728), .dinb(n24727), .dout(n24729));
  jand g07467(.dina(n24729), .dinb(n24716), .dout(n24730));
  jnot g07468(.din(n24595), .dout(n24731));
  jor  g07469(.dina(n24731), .dinb(n24730), .dout(n24732));
  jand g07470(.dina(n24732), .dinb(n24715), .dout(n24733));
  jnot g07471(.din(n24598), .dout(n24734));
  jor  g07472(.dina(n24734), .dinb(n24733), .dout(n24735));
  jand g07473(.dina(n24735), .dinb(n24714), .dout(n24736));
  jnot g07474(.din(n24601), .dout(n24737));
  jor  g07475(.dina(n24737), .dinb(n24736), .dout(n24738));
  jand g07476(.dina(n24738), .dinb(n24713), .dout(n24739));
  jnot g07477(.din(n24604), .dout(n24740));
  jor  g07478(.dina(n24740), .dinb(n24739), .dout(n24741));
  jand g07479(.dina(n24741), .dinb(n24712), .dout(n24742));
  jnot g07480(.din(n24607), .dout(n24743));
  jor  g07481(.dina(n24743), .dinb(n24742), .dout(n24744));
  jand g07482(.dina(n24744), .dinb(n24711), .dout(n24745));
  jnot g07483(.din(n24610), .dout(n24746));
  jor  g07484(.dina(n24746), .dinb(n24745), .dout(n24747));
  jand g07485(.dina(n24747), .dinb(n24710), .dout(n24748));
  jnot g07486(.din(n24613), .dout(n24749));
  jor  g07487(.dina(n24749), .dinb(n24748), .dout(n24750));
  jand g07488(.dina(n24750), .dinb(n24709), .dout(n24751));
  jnot g07489(.din(n24616), .dout(n24752));
  jor  g07490(.dina(n24752), .dinb(n24751), .dout(n24753));
  jand g07491(.dina(n24753), .dinb(n24708), .dout(n24754));
  jnot g07492(.din(n24619), .dout(n24755));
  jor  g07493(.dina(n24755), .dinb(n24754), .dout(n24756));
  jand g07494(.dina(n24756), .dinb(n24707), .dout(n24757));
  jnot g07495(.din(n24622), .dout(n24758));
  jor  g07496(.dina(n24758), .dinb(n24757), .dout(n24759));
  jand g07497(.dina(n24759), .dinb(n24706), .dout(n24760));
  jnot g07498(.din(n24625), .dout(n24761));
  jor  g07499(.dina(n24761), .dinb(n24760), .dout(n24762));
  jand g07500(.dina(n24762), .dinb(n24705), .dout(n24763));
  jnot g07501(.din(n24628), .dout(n24764));
  jor  g07502(.dina(n24764), .dinb(n24763), .dout(n24765));
  jand g07503(.dina(n24765), .dinb(n24704), .dout(n24766));
  jnot g07504(.din(n24631), .dout(n24767));
  jor  g07505(.dina(n24767), .dinb(n24766), .dout(n24768));
  jand g07506(.dina(n24768), .dinb(n24703), .dout(n24769));
  jnot g07507(.din(n24634), .dout(n24770));
  jor  g07508(.dina(n24770), .dinb(n24769), .dout(n24771));
  jand g07509(.dina(n24771), .dinb(n24702), .dout(n24772));
  jnot g07510(.din(n24637), .dout(n24773));
  jor  g07511(.dina(n24773), .dinb(n24772), .dout(n24774));
  jand g07512(.dina(n24774), .dinb(n24701), .dout(n24775));
  jnot g07513(.din(n24640), .dout(n24776));
  jor  g07514(.dina(n24776), .dinb(n24775), .dout(n24777));
  jand g07515(.dina(n24777), .dinb(n24700), .dout(n24778));
  jnot g07516(.din(n24643), .dout(n24779));
  jor  g07517(.dina(n24779), .dinb(n24778), .dout(n24780));
  jand g07518(.dina(n24780), .dinb(n24699), .dout(n24781));
  jnot g07519(.din(n24646), .dout(n24782));
  jor  g07520(.dina(n24782), .dinb(n24781), .dout(n24783));
  jand g07521(.dina(n24783), .dinb(n24698), .dout(n24784));
  jnot g07522(.din(n24649), .dout(n24785));
  jor  g07523(.dina(n24785), .dinb(n24784), .dout(n24786));
  jand g07524(.dina(n24786), .dinb(n24697), .dout(n24787));
  jnot g07525(.din(n24652), .dout(n24788));
  jor  g07526(.dina(n24788), .dinb(n24787), .dout(n24789));
  jand g07527(.dina(n24789), .dinb(n24696), .dout(n24790));
  jnot g07528(.din(n24655), .dout(n24791));
  jor  g07529(.dina(n24791), .dinb(n24790), .dout(n24792));
  jand g07530(.dina(n24792), .dinb(n24695), .dout(n24793));
  jnot g07531(.din(n24658), .dout(n24794));
  jor  g07532(.dina(n24794), .dinb(n24793), .dout(n24795));
  jand g07533(.dina(n24795), .dinb(n24694), .dout(n24796));
  jnot g07534(.din(n24661), .dout(n24797));
  jor  g07535(.dina(n24797), .dinb(n24796), .dout(n24798));
  jand g07536(.dina(n24798), .dinb(n24693), .dout(n24799));
  jnot g07537(.din(n24664), .dout(n24800));
  jor  g07538(.dina(n24800), .dinb(n24799), .dout(n24801));
  jand g07539(.dina(n24801), .dinb(n24692), .dout(n24802));
  jnot g07540(.din(n24667), .dout(n24803));
  jor  g07541(.dina(n24803), .dinb(n24802), .dout(n24804));
  jand g07542(.dina(n24804), .dinb(n24691), .dout(n24805));
  jnot g07543(.din(n24670), .dout(n24806));
  jor  g07544(.dina(n24806), .dinb(n24805), .dout(n24807));
  jand g07545(.dina(n24807), .dinb(n24690), .dout(n24808));
  jnot g07546(.din(n24673), .dout(n24809));
  jor  g07547(.dina(n24809), .dinb(n24808), .dout(n24810));
  jand g07548(.dina(n24810), .dinb(n24689), .dout(n24811));
  jnot g07549(.din(n24676), .dout(n24812));
  jor  g07550(.dina(n24812), .dinb(n24811), .dout(n24813));
  jand g07551(.dina(n24813), .dinb(n24688), .dout(n24814));
  jnot g07552(.din(n24679), .dout(n24815));
  jor  g07553(.dina(n24815), .dinb(n24814), .dout(n24816));
  jand g07554(.dina(n24816), .dinb(n24687), .dout(n24817));
  jand g07555(.dina(n24817), .dinb(n24686), .dout(n24818));
  jor  g07556(.dina(n24818), .dinb(n24276), .dout(n24819));
  jor  g07557(.dina(n24819), .dinb(n853), .dout(n24820));
  jxor g07558(.dina(n24679), .dinb(n24678), .dout(n24821));
  jor  g07559(.dina(n24821), .dinb(n24820), .dout(n24822));
  jand g07560(.dina(n24822), .dinb(n24685), .dout(n24823));
  jand g07561(.dina(n24823), .dinb(n333), .dout(n24824));
  jor  g07562(.dina(n24684), .dinb(n24287), .dout(n24825));
  jxor g07563(.dina(n24676), .dinb(n24675), .dout(n24826));
  jor  g07564(.dina(n24826), .dinb(n24820), .dout(n24827));
  jand g07565(.dina(n24827), .dinb(n24825), .dout(n24828));
  jand g07566(.dina(n24828), .dinb(n332), .dout(n24829));
  jor  g07567(.dina(n24684), .dinb(n24292), .dout(n24830));
  jxor g07568(.dina(n24673), .dinb(n24672), .dout(n24831));
  jor  g07569(.dina(n24831), .dinb(n24820), .dout(n24832));
  jand g07570(.dina(n24832), .dinb(n24830), .dout(n24833));
  jand g07571(.dina(n24833), .dinb(n331), .dout(n24834));
  jor  g07572(.dina(n24684), .dinb(n24297), .dout(n24835));
  jxor g07573(.dina(n24670), .dinb(n24669), .dout(n24836));
  jor  g07574(.dina(n24836), .dinb(n24820), .dout(n24837));
  jand g07575(.dina(n24837), .dinb(n24835), .dout(n24838));
  jand g07576(.dina(n24838), .dinb(n275), .dout(n24839));
  jor  g07577(.dina(n24684), .dinb(n24302), .dout(n24840));
  jxor g07578(.dina(n24667), .dinb(n24666), .dout(n24841));
  jor  g07579(.dina(n24841), .dinb(n24820), .dout(n24842));
  jand g07580(.dina(n24842), .dinb(n24840), .dout(n24843));
  jand g07581(.dina(n24843), .dinb(n340), .dout(n24844));
  jor  g07582(.dina(n24684), .dinb(n24307), .dout(n24845));
  jxor g07583(.dina(n24664), .dinb(n24663), .dout(n24846));
  jor  g07584(.dina(n24846), .dinb(n24820), .dout(n24847));
  jand g07585(.dina(n24847), .dinb(n24845), .dout(n24848));
  jand g07586(.dina(n24848), .dinb(n339), .dout(n24849));
  jor  g07587(.dina(n24684), .dinb(n24312), .dout(n24850));
  jxor g07588(.dina(n24661), .dinb(n24660), .dout(n24851));
  jor  g07589(.dina(n24851), .dinb(n24820), .dout(n24852));
  jand g07590(.dina(n24852), .dinb(n24850), .dout(n24853));
  jand g07591(.dina(n24853), .dinb(n338), .dout(n24854));
  jor  g07592(.dina(n24684), .dinb(n24317), .dout(n24855));
  jxor g07593(.dina(n24658), .dinb(n24657), .dout(n24856));
  jor  g07594(.dina(n24856), .dinb(n24820), .dout(n24857));
  jand g07595(.dina(n24857), .dinb(n24855), .dout(n24858));
  jand g07596(.dina(n24858), .dinb(n271), .dout(n24859));
  jor  g07597(.dina(n24684), .dinb(n24322), .dout(n24860));
  jxor g07598(.dina(n24655), .dinb(n24654), .dout(n24861));
  jor  g07599(.dina(n24861), .dinb(n24820), .dout(n24862));
  jand g07600(.dina(n24862), .dinb(n24860), .dout(n24863));
  jand g07601(.dina(n24863), .dinb(n270), .dout(n24864));
  jor  g07602(.dina(n24684), .dinb(n24327), .dout(n24865));
  jxor g07603(.dina(n24652), .dinb(n24651), .dout(n24866));
  jor  g07604(.dina(n24866), .dinb(n24820), .dout(n24867));
  jand g07605(.dina(n24867), .dinb(n24865), .dout(n24868));
  jand g07606(.dina(n24868), .dinb(n269), .dout(n24869));
  jor  g07607(.dina(n24684), .dinb(n24332), .dout(n24870));
  jxor g07608(.dina(n24649), .dinb(n24648), .dout(n24871));
  jor  g07609(.dina(n24871), .dinb(n24820), .dout(n24872));
  jand g07610(.dina(n24872), .dinb(n24870), .dout(n24873));
  jand g07611(.dina(n24873), .dinb(n274), .dout(n24874));
  jor  g07612(.dina(n24684), .dinb(n24337), .dout(n24875));
  jxor g07613(.dina(n24646), .dinb(n24645), .dout(n24876));
  jor  g07614(.dina(n24876), .dinb(n24820), .dout(n24877));
  jand g07615(.dina(n24877), .dinb(n24875), .dout(n24878));
  jand g07616(.dina(n24878), .dinb(n268), .dout(n24879));
  jor  g07617(.dina(n24684), .dinb(n24342), .dout(n24880));
  jxor g07618(.dina(n24643), .dinb(n24642), .dout(n24881));
  jor  g07619(.dina(n24881), .dinb(n24820), .dout(n24882));
  jand g07620(.dina(n24882), .dinb(n24880), .dout(n24883));
  jand g07621(.dina(n24883), .dinb(n349), .dout(n24884));
  jor  g07622(.dina(n24684), .dinb(n24347), .dout(n24885));
  jxor g07623(.dina(n24640), .dinb(n24639), .dout(n24886));
  jor  g07624(.dina(n24886), .dinb(n24820), .dout(n24887));
  jand g07625(.dina(n24887), .dinb(n24885), .dout(n24888));
  jand g07626(.dina(n24888), .dinb(n348), .dout(n24889));
  jor  g07627(.dina(n24684), .dinb(n24352), .dout(n24890));
  jxor g07628(.dina(n24637), .dinb(n24636), .dout(n24891));
  jor  g07629(.dina(n24891), .dinb(n24820), .dout(n24892));
  jand g07630(.dina(n24892), .dinb(n24890), .dout(n24893));
  jand g07631(.dina(n24893), .dinb(n347), .dout(n24894));
  jor  g07632(.dina(n24684), .dinb(n24357), .dout(n24895));
  jxor g07633(.dina(n24634), .dinb(n24633), .dout(n24896));
  jor  g07634(.dina(n24896), .dinb(n24820), .dout(n24897));
  jand g07635(.dina(n24897), .dinb(n24895), .dout(n24898));
  jand g07636(.dina(n24898), .dinb(n267), .dout(n24899));
  jor  g07637(.dina(n24684), .dinb(n24362), .dout(n24900));
  jxor g07638(.dina(n24631), .dinb(n24630), .dout(n24901));
  jor  g07639(.dina(n24901), .dinb(n24820), .dout(n24902));
  jand g07640(.dina(n24902), .dinb(n24900), .dout(n24903));
  jand g07641(.dina(n24903), .dinb(n266), .dout(n24904));
  jor  g07642(.dina(n24684), .dinb(n24367), .dout(n24905));
  jxor g07643(.dina(n24628), .dinb(n24627), .dout(n24906));
  jor  g07644(.dina(n24906), .dinb(n24820), .dout(n24907));
  jand g07645(.dina(n24907), .dinb(n24905), .dout(n24908));
  jand g07646(.dina(n24908), .dinb(n356), .dout(n24909));
  jor  g07647(.dina(n24684), .dinb(n24372), .dout(n24910));
  jxor g07648(.dina(n24625), .dinb(n24624), .dout(n24911));
  jor  g07649(.dina(n24911), .dinb(n24820), .dout(n24912));
  jand g07650(.dina(n24912), .dinb(n24910), .dout(n24913));
  jand g07651(.dina(n24913), .dinb(n355), .dout(n24914));
  jor  g07652(.dina(n24684), .dinb(n24377), .dout(n24915));
  jxor g07653(.dina(n24622), .dinb(n24621), .dout(n24916));
  jor  g07654(.dina(n24916), .dinb(n24820), .dout(n24917));
  jand g07655(.dina(n24917), .dinb(n24915), .dout(n24918));
  jand g07656(.dina(n24918), .dinb(n364), .dout(n24919));
  jor  g07657(.dina(n24684), .dinb(n24382), .dout(n24920));
  jxor g07658(.dina(n24619), .dinb(n24618), .dout(n24921));
  jor  g07659(.dina(n24921), .dinb(n24820), .dout(n24922));
  jand g07660(.dina(n24922), .dinb(n24920), .dout(n24923));
  jand g07661(.dina(n24923), .dinb(n361), .dout(n24924));
  jor  g07662(.dina(n24684), .dinb(n24387), .dout(n24925));
  jxor g07663(.dina(n24616), .dinb(n24615), .dout(n24926));
  jor  g07664(.dina(n24926), .dinb(n24820), .dout(n24927));
  jand g07665(.dina(n24927), .dinb(n24925), .dout(n24928));
  jand g07666(.dina(n24928), .dinb(n360), .dout(n24929));
  jor  g07667(.dina(n24684), .dinb(n24392), .dout(n24930));
  jxor g07668(.dina(n24613), .dinb(n24612), .dout(n24931));
  jor  g07669(.dina(n24931), .dinb(n24820), .dout(n24932));
  jand g07670(.dina(n24932), .dinb(n24930), .dout(n24933));
  jand g07671(.dina(n24933), .dinb(n363), .dout(n24934));
  jor  g07672(.dina(n24684), .dinb(n24397), .dout(n24935));
  jxor g07673(.dina(n24610), .dinb(n24609), .dout(n24936));
  jor  g07674(.dina(n24936), .dinb(n24820), .dout(n24937));
  jand g07675(.dina(n24937), .dinb(n24935), .dout(n24938));
  jand g07676(.dina(n24938), .dinb(n359), .dout(n24939));
  jor  g07677(.dina(n24684), .dinb(n24402), .dout(n24940));
  jxor g07678(.dina(n24607), .dinb(n24606), .dout(n24941));
  jor  g07679(.dina(n24941), .dinb(n24820), .dout(n24942));
  jand g07680(.dina(n24942), .dinb(n24940), .dout(n24943));
  jand g07681(.dina(n24943), .dinb(n369), .dout(n24944));
  jor  g07682(.dina(n24684), .dinb(n24407), .dout(n24945));
  jxor g07683(.dina(n24604), .dinb(n24603), .dout(n24946));
  jor  g07684(.dina(n24946), .dinb(n24820), .dout(n24947));
  jand g07685(.dina(n24947), .dinb(n24945), .dout(n24948));
  jand g07686(.dina(n24948), .dinb(n368), .dout(n24949));
  jor  g07687(.dina(n24684), .dinb(n24412), .dout(n24950));
  jxor g07688(.dina(n24601), .dinb(n24600), .dout(n24951));
  jor  g07689(.dina(n24951), .dinb(n24820), .dout(n24952));
  jand g07690(.dina(n24952), .dinb(n24950), .dout(n24953));
  jand g07691(.dina(n24953), .dinb(n367), .dout(n24954));
  jor  g07692(.dina(n24684), .dinb(n24417), .dout(n24955));
  jxor g07693(.dina(n24598), .dinb(n24597), .dout(n24956));
  jor  g07694(.dina(n24956), .dinb(n24820), .dout(n24957));
  jand g07695(.dina(n24957), .dinb(n24955), .dout(n24958));
  jand g07696(.dina(n24958), .dinb(n265), .dout(n24959));
  jor  g07697(.dina(n24684), .dinb(n24422), .dout(n24960));
  jxor g07698(.dina(n24595), .dinb(n24594), .dout(n24961));
  jor  g07699(.dina(n24961), .dinb(n24820), .dout(n24962));
  jand g07700(.dina(n24962), .dinb(n24960), .dout(n24963));
  jand g07701(.dina(n24963), .dinb(n378), .dout(n24964));
  jor  g07702(.dina(n24684), .dinb(n24427), .dout(n24965));
  jxor g07703(.dina(n24592), .dinb(n24591), .dout(n24966));
  jor  g07704(.dina(n24966), .dinb(n24820), .dout(n24967));
  jand g07705(.dina(n24967), .dinb(n24965), .dout(n24968));
  jand g07706(.dina(n24968), .dinb(n377), .dout(n24969));
  jor  g07707(.dina(n24684), .dinb(n24432), .dout(n24970));
  jxor g07708(.dina(n24589), .dinb(n24588), .dout(n24971));
  jor  g07709(.dina(n24971), .dinb(n24820), .dout(n24972));
  jand g07710(.dina(n24972), .dinb(n24970), .dout(n24973));
  jand g07711(.dina(n24973), .dinb(n376), .dout(n24974));
  jnot g07712(.din(n24438), .dout(n24975));
  jor  g07713(.dina(n24684), .dinb(n24975), .dout(n24976));
  jxor g07714(.dina(n24586), .dinb(n24585), .dout(n24977));
  jor  g07715(.dina(n24977), .dinb(n24820), .dout(n24978));
  jand g07716(.dina(n24978), .dinb(n24976), .dout(n24979));
  jand g07717(.dina(n24979), .dinb(n264), .dout(n24980));
  jand g07718(.dina(n24820), .dinb(n24578), .dout(n24981));
  jxor g07719(.dina(n24583), .dinb(n5777), .dout(n24982));
  jand g07720(.dina(n24982), .dinb(n24684), .dout(n24983));
  jor  g07721(.dina(n24983), .dinb(n24981), .dout(n24984));
  jand g07722(.dina(n24984), .dinb(n386), .dout(n24985));
  jnot g07723(.din(n6018), .dout(n24986));
  jor  g07724(.dina(n24819), .dinb(n24986), .dout(n24987));
  jand g07725(.dina(n24987), .dinb(a29 ), .dout(n24988));
  jand g07726(.dina(n24684), .dinb(n5639), .dout(n24989));
  jor  g07727(.dina(n24989), .dinb(n24988), .dout(n24990));
  jand g07728(.dina(n24990), .dinb(n259), .dout(n24991));
  jand g07729(.dina(n24683), .dinb(n6018), .dout(n24992));
  jor  g07730(.dina(n24992), .dinb(n5638), .dout(n24993));
  jor  g07731(.dina(n24820), .dinb(n5777), .dout(n24994));
  jand g07732(.dina(n24994), .dinb(n24993), .dout(n24995));
  jxor g07733(.dina(n24995), .dinb(b1 ), .dout(n24996));
  jand g07734(.dina(n24996), .dinb(n6027), .dout(n24997));
  jor  g07735(.dina(n24997), .dinb(n24991), .dout(n24998));
  jxor g07736(.dina(n24984), .dinb(n386), .dout(n24999));
  jand g07737(.dina(n24999), .dinb(n24998), .dout(n25000));
  jor  g07738(.dina(n25000), .dinb(n24985), .dout(n25001));
  jxor g07739(.dina(n24979), .dinb(n264), .dout(n25002));
  jand g07740(.dina(n25002), .dinb(n25001), .dout(n25003));
  jor  g07741(.dina(n25003), .dinb(n24980), .dout(n25004));
  jxor g07742(.dina(n24973), .dinb(n376), .dout(n25005));
  jand g07743(.dina(n25005), .dinb(n25004), .dout(n25006));
  jor  g07744(.dina(n25006), .dinb(n24974), .dout(n25007));
  jxor g07745(.dina(n24968), .dinb(n377), .dout(n25008));
  jand g07746(.dina(n25008), .dinb(n25007), .dout(n25009));
  jor  g07747(.dina(n25009), .dinb(n24969), .dout(n25010));
  jxor g07748(.dina(n24963), .dinb(n378), .dout(n25011));
  jand g07749(.dina(n25011), .dinb(n25010), .dout(n25012));
  jor  g07750(.dina(n25012), .dinb(n24964), .dout(n25013));
  jxor g07751(.dina(n24958), .dinb(n265), .dout(n25014));
  jand g07752(.dina(n25014), .dinb(n25013), .dout(n25015));
  jor  g07753(.dina(n25015), .dinb(n24959), .dout(n25016));
  jxor g07754(.dina(n24953), .dinb(n367), .dout(n25017));
  jand g07755(.dina(n25017), .dinb(n25016), .dout(n25018));
  jor  g07756(.dina(n25018), .dinb(n24954), .dout(n25019));
  jxor g07757(.dina(n24948), .dinb(n368), .dout(n25020));
  jand g07758(.dina(n25020), .dinb(n25019), .dout(n25021));
  jor  g07759(.dina(n25021), .dinb(n24949), .dout(n25022));
  jxor g07760(.dina(n24943), .dinb(n369), .dout(n25023));
  jand g07761(.dina(n25023), .dinb(n25022), .dout(n25024));
  jor  g07762(.dina(n25024), .dinb(n24944), .dout(n25025));
  jxor g07763(.dina(n24938), .dinb(n359), .dout(n25026));
  jand g07764(.dina(n25026), .dinb(n25025), .dout(n25027));
  jor  g07765(.dina(n25027), .dinb(n24939), .dout(n25028));
  jxor g07766(.dina(n24933), .dinb(n363), .dout(n25029));
  jand g07767(.dina(n25029), .dinb(n25028), .dout(n25030));
  jor  g07768(.dina(n25030), .dinb(n24934), .dout(n25031));
  jxor g07769(.dina(n24928), .dinb(n360), .dout(n25032));
  jand g07770(.dina(n25032), .dinb(n25031), .dout(n25033));
  jor  g07771(.dina(n25033), .dinb(n24929), .dout(n25034));
  jxor g07772(.dina(n24923), .dinb(n361), .dout(n25035));
  jand g07773(.dina(n25035), .dinb(n25034), .dout(n25036));
  jor  g07774(.dina(n25036), .dinb(n24924), .dout(n25037));
  jxor g07775(.dina(n24918), .dinb(n364), .dout(n25038));
  jand g07776(.dina(n25038), .dinb(n25037), .dout(n25039));
  jor  g07777(.dina(n25039), .dinb(n24919), .dout(n25040));
  jxor g07778(.dina(n24913), .dinb(n355), .dout(n25041));
  jand g07779(.dina(n25041), .dinb(n25040), .dout(n25042));
  jor  g07780(.dina(n25042), .dinb(n24914), .dout(n25043));
  jxor g07781(.dina(n24908), .dinb(n356), .dout(n25044));
  jand g07782(.dina(n25044), .dinb(n25043), .dout(n25045));
  jor  g07783(.dina(n25045), .dinb(n24909), .dout(n25046));
  jxor g07784(.dina(n24903), .dinb(n266), .dout(n25047));
  jand g07785(.dina(n25047), .dinb(n25046), .dout(n25048));
  jor  g07786(.dina(n25048), .dinb(n24904), .dout(n25049));
  jxor g07787(.dina(n24898), .dinb(n267), .dout(n25050));
  jand g07788(.dina(n25050), .dinb(n25049), .dout(n25051));
  jor  g07789(.dina(n25051), .dinb(n24899), .dout(n25052));
  jxor g07790(.dina(n24893), .dinb(n347), .dout(n25053));
  jand g07791(.dina(n25053), .dinb(n25052), .dout(n25054));
  jor  g07792(.dina(n25054), .dinb(n24894), .dout(n25055));
  jxor g07793(.dina(n24888), .dinb(n348), .dout(n25056));
  jand g07794(.dina(n25056), .dinb(n25055), .dout(n25057));
  jor  g07795(.dina(n25057), .dinb(n24889), .dout(n25058));
  jxor g07796(.dina(n24883), .dinb(n349), .dout(n25059));
  jand g07797(.dina(n25059), .dinb(n25058), .dout(n25060));
  jor  g07798(.dina(n25060), .dinb(n24884), .dout(n25061));
  jxor g07799(.dina(n24878), .dinb(n268), .dout(n25062));
  jand g07800(.dina(n25062), .dinb(n25061), .dout(n25063));
  jor  g07801(.dina(n25063), .dinb(n24879), .dout(n25064));
  jxor g07802(.dina(n24873), .dinb(n274), .dout(n25065));
  jand g07803(.dina(n25065), .dinb(n25064), .dout(n25066));
  jor  g07804(.dina(n25066), .dinb(n24874), .dout(n25067));
  jxor g07805(.dina(n24868), .dinb(n269), .dout(n25068));
  jand g07806(.dina(n25068), .dinb(n25067), .dout(n25069));
  jor  g07807(.dina(n25069), .dinb(n24869), .dout(n25070));
  jxor g07808(.dina(n24863), .dinb(n270), .dout(n25071));
  jand g07809(.dina(n25071), .dinb(n25070), .dout(n25072));
  jor  g07810(.dina(n25072), .dinb(n24864), .dout(n25073));
  jxor g07811(.dina(n24858), .dinb(n271), .dout(n25074));
  jand g07812(.dina(n25074), .dinb(n25073), .dout(n25075));
  jor  g07813(.dina(n25075), .dinb(n24859), .dout(n25076));
  jxor g07814(.dina(n24853), .dinb(n338), .dout(n25077));
  jand g07815(.dina(n25077), .dinb(n25076), .dout(n25078));
  jor  g07816(.dina(n25078), .dinb(n24854), .dout(n25079));
  jxor g07817(.dina(n24848), .dinb(n339), .dout(n25080));
  jand g07818(.dina(n25080), .dinb(n25079), .dout(n25081));
  jor  g07819(.dina(n25081), .dinb(n24849), .dout(n25082));
  jxor g07820(.dina(n24843), .dinb(n340), .dout(n25083));
  jand g07821(.dina(n25083), .dinb(n25082), .dout(n25084));
  jor  g07822(.dina(n25084), .dinb(n24844), .dout(n25085));
  jxor g07823(.dina(n24838), .dinb(n275), .dout(n25086));
  jand g07824(.dina(n25086), .dinb(n25085), .dout(n25087));
  jor  g07825(.dina(n25087), .dinb(n24839), .dout(n25088));
  jxor g07826(.dina(n24833), .dinb(n331), .dout(n25089));
  jand g07827(.dina(n25089), .dinb(n25088), .dout(n25090));
  jor  g07828(.dina(n25090), .dinb(n24834), .dout(n25091));
  jxor g07829(.dina(n24828), .dinb(n332), .dout(n25092));
  jand g07830(.dina(n25092), .dinb(n25091), .dout(n25093));
  jor  g07831(.dina(n25093), .dinb(n24829), .dout(n25094));
  jxor g07832(.dina(n24823), .dinb(n333), .dout(n25095));
  jand g07833(.dina(n25095), .dinb(n25094), .dout(n25096));
  jor  g07834(.dina(n25096), .dinb(n24824), .dout(n25097));
  jand g07835(.dina(n24820), .dinb(n24281), .dout(n25098));
  jand g07836(.dina(n24681), .dinb(n24282), .dout(n25099));
  jand g07837(.dina(n25099), .dinb(n410), .dout(n25100));
  jor  g07838(.dina(n25100), .dinb(n25098), .dout(n25101));
  jxor g07839(.dina(n25101), .dinb(b35 ), .dout(n25102));
  jnot g07840(.din(n25102), .dout(n25103));
  jand g07841(.dina(n25103), .dinb(n25097), .dout(n25104));
  jand g07842(.dina(n25104), .dinb(n329), .dout(n25105));
  jand g07843(.dina(n25101), .dinb(n410), .dout(n25106));
  jor  g07844(.dina(n25106), .dinb(n25105), .dout(n25107));
  jor  g07845(.dina(n25107), .dinb(n24823), .dout(n25108));
  jnot g07846(.din(n24824), .dout(n25109));
  jnot g07847(.din(n24829), .dout(n25110));
  jnot g07848(.din(n24834), .dout(n25111));
  jnot g07849(.din(n24839), .dout(n25112));
  jnot g07850(.din(n24844), .dout(n25113));
  jnot g07851(.din(n24849), .dout(n25114));
  jnot g07852(.din(n24854), .dout(n25115));
  jnot g07853(.din(n24859), .dout(n25116));
  jnot g07854(.din(n24864), .dout(n25117));
  jnot g07855(.din(n24869), .dout(n25118));
  jnot g07856(.din(n24874), .dout(n25119));
  jnot g07857(.din(n24879), .dout(n25120));
  jnot g07858(.din(n24884), .dout(n25121));
  jnot g07859(.din(n24889), .dout(n25122));
  jnot g07860(.din(n24894), .dout(n25123));
  jnot g07861(.din(n24899), .dout(n25124));
  jnot g07862(.din(n24904), .dout(n25125));
  jnot g07863(.din(n24909), .dout(n25126));
  jnot g07864(.din(n24914), .dout(n25127));
  jnot g07865(.din(n24919), .dout(n25128));
  jnot g07866(.din(n24924), .dout(n25129));
  jnot g07867(.din(n24929), .dout(n25130));
  jnot g07868(.din(n24934), .dout(n25131));
  jnot g07869(.din(n24939), .dout(n25132));
  jnot g07870(.din(n24944), .dout(n25133));
  jnot g07871(.din(n24949), .dout(n25134));
  jnot g07872(.din(n24954), .dout(n25135));
  jnot g07873(.din(n24959), .dout(n25136));
  jnot g07874(.din(n24964), .dout(n25137));
  jnot g07875(.din(n24969), .dout(n25138));
  jnot g07876(.din(n24974), .dout(n25139));
  jnot g07877(.din(n24980), .dout(n25140));
  jnot g07878(.din(n24985), .dout(n25141));
  jnot g07879(.din(n24991), .dout(n25142));
  jxor g07880(.dina(n24995), .dinb(n259), .dout(n25143));
  jor  g07881(.dina(n25143), .dinb(n6026), .dout(n25144));
  jand g07882(.dina(n25144), .dinb(n25142), .dout(n25145));
  jnot g07883(.din(n24999), .dout(n25146));
  jor  g07884(.dina(n25146), .dinb(n25145), .dout(n25147));
  jand g07885(.dina(n25147), .dinb(n25141), .dout(n25148));
  jnot g07886(.din(n25002), .dout(n25149));
  jor  g07887(.dina(n25149), .dinb(n25148), .dout(n25150));
  jand g07888(.dina(n25150), .dinb(n25140), .dout(n25151));
  jnot g07889(.din(n25005), .dout(n25152));
  jor  g07890(.dina(n25152), .dinb(n25151), .dout(n25153));
  jand g07891(.dina(n25153), .dinb(n25139), .dout(n25154));
  jnot g07892(.din(n25008), .dout(n25155));
  jor  g07893(.dina(n25155), .dinb(n25154), .dout(n25156));
  jand g07894(.dina(n25156), .dinb(n25138), .dout(n25157));
  jnot g07895(.din(n25011), .dout(n25158));
  jor  g07896(.dina(n25158), .dinb(n25157), .dout(n25159));
  jand g07897(.dina(n25159), .dinb(n25137), .dout(n25160));
  jnot g07898(.din(n25014), .dout(n25161));
  jor  g07899(.dina(n25161), .dinb(n25160), .dout(n25162));
  jand g07900(.dina(n25162), .dinb(n25136), .dout(n25163));
  jnot g07901(.din(n25017), .dout(n25164));
  jor  g07902(.dina(n25164), .dinb(n25163), .dout(n25165));
  jand g07903(.dina(n25165), .dinb(n25135), .dout(n25166));
  jnot g07904(.din(n25020), .dout(n25167));
  jor  g07905(.dina(n25167), .dinb(n25166), .dout(n25168));
  jand g07906(.dina(n25168), .dinb(n25134), .dout(n25169));
  jnot g07907(.din(n25023), .dout(n25170));
  jor  g07908(.dina(n25170), .dinb(n25169), .dout(n25171));
  jand g07909(.dina(n25171), .dinb(n25133), .dout(n25172));
  jnot g07910(.din(n25026), .dout(n25173));
  jor  g07911(.dina(n25173), .dinb(n25172), .dout(n25174));
  jand g07912(.dina(n25174), .dinb(n25132), .dout(n25175));
  jnot g07913(.din(n25029), .dout(n25176));
  jor  g07914(.dina(n25176), .dinb(n25175), .dout(n25177));
  jand g07915(.dina(n25177), .dinb(n25131), .dout(n25178));
  jnot g07916(.din(n25032), .dout(n25179));
  jor  g07917(.dina(n25179), .dinb(n25178), .dout(n25180));
  jand g07918(.dina(n25180), .dinb(n25130), .dout(n25181));
  jnot g07919(.din(n25035), .dout(n25182));
  jor  g07920(.dina(n25182), .dinb(n25181), .dout(n25183));
  jand g07921(.dina(n25183), .dinb(n25129), .dout(n25184));
  jnot g07922(.din(n25038), .dout(n25185));
  jor  g07923(.dina(n25185), .dinb(n25184), .dout(n25186));
  jand g07924(.dina(n25186), .dinb(n25128), .dout(n25187));
  jnot g07925(.din(n25041), .dout(n25188));
  jor  g07926(.dina(n25188), .dinb(n25187), .dout(n25189));
  jand g07927(.dina(n25189), .dinb(n25127), .dout(n25190));
  jnot g07928(.din(n25044), .dout(n25191));
  jor  g07929(.dina(n25191), .dinb(n25190), .dout(n25192));
  jand g07930(.dina(n25192), .dinb(n25126), .dout(n25193));
  jnot g07931(.din(n25047), .dout(n25194));
  jor  g07932(.dina(n25194), .dinb(n25193), .dout(n25195));
  jand g07933(.dina(n25195), .dinb(n25125), .dout(n25196));
  jnot g07934(.din(n25050), .dout(n25197));
  jor  g07935(.dina(n25197), .dinb(n25196), .dout(n25198));
  jand g07936(.dina(n25198), .dinb(n25124), .dout(n25199));
  jnot g07937(.din(n25053), .dout(n25200));
  jor  g07938(.dina(n25200), .dinb(n25199), .dout(n25201));
  jand g07939(.dina(n25201), .dinb(n25123), .dout(n25202));
  jnot g07940(.din(n25056), .dout(n25203));
  jor  g07941(.dina(n25203), .dinb(n25202), .dout(n25204));
  jand g07942(.dina(n25204), .dinb(n25122), .dout(n25205));
  jnot g07943(.din(n25059), .dout(n25206));
  jor  g07944(.dina(n25206), .dinb(n25205), .dout(n25207));
  jand g07945(.dina(n25207), .dinb(n25121), .dout(n25208));
  jnot g07946(.din(n25062), .dout(n25209));
  jor  g07947(.dina(n25209), .dinb(n25208), .dout(n25210));
  jand g07948(.dina(n25210), .dinb(n25120), .dout(n25211));
  jnot g07949(.din(n25065), .dout(n25212));
  jor  g07950(.dina(n25212), .dinb(n25211), .dout(n25213));
  jand g07951(.dina(n25213), .dinb(n25119), .dout(n25214));
  jnot g07952(.din(n25068), .dout(n25215));
  jor  g07953(.dina(n25215), .dinb(n25214), .dout(n25216));
  jand g07954(.dina(n25216), .dinb(n25118), .dout(n25217));
  jnot g07955(.din(n25071), .dout(n25218));
  jor  g07956(.dina(n25218), .dinb(n25217), .dout(n25219));
  jand g07957(.dina(n25219), .dinb(n25117), .dout(n25220));
  jnot g07958(.din(n25074), .dout(n25221));
  jor  g07959(.dina(n25221), .dinb(n25220), .dout(n25222));
  jand g07960(.dina(n25222), .dinb(n25116), .dout(n25223));
  jnot g07961(.din(n25077), .dout(n25224));
  jor  g07962(.dina(n25224), .dinb(n25223), .dout(n25225));
  jand g07963(.dina(n25225), .dinb(n25115), .dout(n25226));
  jnot g07964(.din(n25080), .dout(n25227));
  jor  g07965(.dina(n25227), .dinb(n25226), .dout(n25228));
  jand g07966(.dina(n25228), .dinb(n25114), .dout(n25229));
  jnot g07967(.din(n25083), .dout(n25230));
  jor  g07968(.dina(n25230), .dinb(n25229), .dout(n25231));
  jand g07969(.dina(n25231), .dinb(n25113), .dout(n25232));
  jnot g07970(.din(n25086), .dout(n25233));
  jor  g07971(.dina(n25233), .dinb(n25232), .dout(n25234));
  jand g07972(.dina(n25234), .dinb(n25112), .dout(n25235));
  jnot g07973(.din(n25089), .dout(n25236));
  jor  g07974(.dina(n25236), .dinb(n25235), .dout(n25237));
  jand g07975(.dina(n25237), .dinb(n25111), .dout(n25238));
  jnot g07976(.din(n25092), .dout(n25239));
  jor  g07977(.dina(n25239), .dinb(n25238), .dout(n25240));
  jand g07978(.dina(n25240), .dinb(n25110), .dout(n25241));
  jnot g07979(.din(n25095), .dout(n25242));
  jor  g07980(.dina(n25242), .dinb(n25241), .dout(n25243));
  jand g07981(.dina(n25243), .dinb(n25109), .dout(n25244));
  jor  g07982(.dina(n25102), .dinb(n25244), .dout(n25245));
  jor  g07983(.dina(n25245), .dinb(n852), .dout(n25246));
  jnot g07984(.din(n25106), .dout(n25247));
  jand g07985(.dina(n25247), .dinb(n25246), .dout(n25248));
  jxor g07986(.dina(n25095), .dinb(n25094), .dout(n25249));
  jor  g07987(.dina(n25249), .dinb(n25248), .dout(n25250));
  jand g07988(.dina(n25250), .dinb(n25108), .dout(n25251));
  jxor g07989(.dina(n25102), .dinb(n25244), .dout(n25252));
  jor  g07990(.dina(n25252), .dinb(n25248), .dout(n25253));
  jor  g07991(.dina(n25105), .dinb(n25101), .dout(n25254));
  jand g07992(.dina(n25254), .dinb(n25253), .dout(n25255));
  jand g07993(.dina(n25255), .dinb(n324), .dout(n25256));
  jnot g07994(.din(n25255), .dout(n25257));
  jand g07995(.dina(n25257), .dinb(b36 ), .dout(n25258));
  jnot g07996(.din(n25258), .dout(n25259));
  jand g07997(.dina(n25251), .dinb(n276), .dout(n25260));
  jor  g07998(.dina(n25107), .dinb(n24828), .dout(n25261));
  jxor g07999(.dina(n25092), .dinb(n25091), .dout(n25262));
  jor  g08000(.dina(n25262), .dinb(n25248), .dout(n25263));
  jand g08001(.dina(n25263), .dinb(n25261), .dout(n25264));
  jand g08002(.dina(n25264), .dinb(n333), .dout(n25265));
  jor  g08003(.dina(n25107), .dinb(n24833), .dout(n25266));
  jxor g08004(.dina(n25089), .dinb(n25088), .dout(n25267));
  jor  g08005(.dina(n25267), .dinb(n25248), .dout(n25268));
  jand g08006(.dina(n25268), .dinb(n25266), .dout(n25269));
  jand g08007(.dina(n25269), .dinb(n332), .dout(n25270));
  jor  g08008(.dina(n25107), .dinb(n24838), .dout(n25271));
  jxor g08009(.dina(n25086), .dinb(n25085), .dout(n25272));
  jor  g08010(.dina(n25272), .dinb(n25248), .dout(n25273));
  jand g08011(.dina(n25273), .dinb(n25271), .dout(n25274));
  jand g08012(.dina(n25274), .dinb(n331), .dout(n25275));
  jor  g08013(.dina(n25107), .dinb(n24843), .dout(n25276));
  jxor g08014(.dina(n25083), .dinb(n25082), .dout(n25277));
  jor  g08015(.dina(n25277), .dinb(n25248), .dout(n25278));
  jand g08016(.dina(n25278), .dinb(n25276), .dout(n25279));
  jand g08017(.dina(n25279), .dinb(n275), .dout(n25280));
  jor  g08018(.dina(n25107), .dinb(n24848), .dout(n25281));
  jxor g08019(.dina(n25080), .dinb(n25079), .dout(n25282));
  jor  g08020(.dina(n25282), .dinb(n25248), .dout(n25283));
  jand g08021(.dina(n25283), .dinb(n25281), .dout(n25284));
  jand g08022(.dina(n25284), .dinb(n340), .dout(n25285));
  jor  g08023(.dina(n25107), .dinb(n24853), .dout(n25286));
  jxor g08024(.dina(n25077), .dinb(n25076), .dout(n25287));
  jor  g08025(.dina(n25287), .dinb(n25248), .dout(n25288));
  jand g08026(.dina(n25288), .dinb(n25286), .dout(n25289));
  jand g08027(.dina(n25289), .dinb(n339), .dout(n25290));
  jor  g08028(.dina(n25107), .dinb(n24858), .dout(n25291));
  jxor g08029(.dina(n25074), .dinb(n25073), .dout(n25292));
  jor  g08030(.dina(n25292), .dinb(n25248), .dout(n25293));
  jand g08031(.dina(n25293), .dinb(n25291), .dout(n25294));
  jand g08032(.dina(n25294), .dinb(n338), .dout(n25295));
  jor  g08033(.dina(n25107), .dinb(n24863), .dout(n25296));
  jxor g08034(.dina(n25071), .dinb(n25070), .dout(n25297));
  jor  g08035(.dina(n25297), .dinb(n25248), .dout(n25298));
  jand g08036(.dina(n25298), .dinb(n25296), .dout(n25299));
  jand g08037(.dina(n25299), .dinb(n271), .dout(n25300));
  jor  g08038(.dina(n25107), .dinb(n24868), .dout(n25301));
  jxor g08039(.dina(n25068), .dinb(n25067), .dout(n25302));
  jor  g08040(.dina(n25302), .dinb(n25248), .dout(n25303));
  jand g08041(.dina(n25303), .dinb(n25301), .dout(n25304));
  jand g08042(.dina(n25304), .dinb(n270), .dout(n25305));
  jor  g08043(.dina(n25107), .dinb(n24873), .dout(n25306));
  jxor g08044(.dina(n25065), .dinb(n25064), .dout(n25307));
  jor  g08045(.dina(n25307), .dinb(n25248), .dout(n25308));
  jand g08046(.dina(n25308), .dinb(n25306), .dout(n25309));
  jand g08047(.dina(n25309), .dinb(n269), .dout(n25310));
  jor  g08048(.dina(n25107), .dinb(n24878), .dout(n25311));
  jxor g08049(.dina(n25062), .dinb(n25061), .dout(n25312));
  jor  g08050(.dina(n25312), .dinb(n25248), .dout(n25313));
  jand g08051(.dina(n25313), .dinb(n25311), .dout(n25314));
  jand g08052(.dina(n25314), .dinb(n274), .dout(n25315));
  jor  g08053(.dina(n25107), .dinb(n24883), .dout(n25316));
  jxor g08054(.dina(n25059), .dinb(n25058), .dout(n25317));
  jor  g08055(.dina(n25317), .dinb(n25248), .dout(n25318));
  jand g08056(.dina(n25318), .dinb(n25316), .dout(n25319));
  jand g08057(.dina(n25319), .dinb(n268), .dout(n25320));
  jor  g08058(.dina(n25107), .dinb(n24888), .dout(n25321));
  jxor g08059(.dina(n25056), .dinb(n25055), .dout(n25322));
  jor  g08060(.dina(n25322), .dinb(n25248), .dout(n25323));
  jand g08061(.dina(n25323), .dinb(n25321), .dout(n25324));
  jand g08062(.dina(n25324), .dinb(n349), .dout(n25325));
  jor  g08063(.dina(n25107), .dinb(n24893), .dout(n25326));
  jxor g08064(.dina(n25053), .dinb(n25052), .dout(n25327));
  jor  g08065(.dina(n25327), .dinb(n25248), .dout(n25328));
  jand g08066(.dina(n25328), .dinb(n25326), .dout(n25329));
  jand g08067(.dina(n25329), .dinb(n348), .dout(n25330));
  jor  g08068(.dina(n25107), .dinb(n24898), .dout(n25331));
  jxor g08069(.dina(n25050), .dinb(n25049), .dout(n25332));
  jor  g08070(.dina(n25332), .dinb(n25248), .dout(n25333));
  jand g08071(.dina(n25333), .dinb(n25331), .dout(n25334));
  jand g08072(.dina(n25334), .dinb(n347), .dout(n25335));
  jor  g08073(.dina(n25107), .dinb(n24903), .dout(n25336));
  jxor g08074(.dina(n25047), .dinb(n25046), .dout(n25337));
  jor  g08075(.dina(n25337), .dinb(n25248), .dout(n25338));
  jand g08076(.dina(n25338), .dinb(n25336), .dout(n25339));
  jand g08077(.dina(n25339), .dinb(n267), .dout(n25340));
  jor  g08078(.dina(n25107), .dinb(n24908), .dout(n25341));
  jxor g08079(.dina(n25044), .dinb(n25043), .dout(n25342));
  jor  g08080(.dina(n25342), .dinb(n25248), .dout(n25343));
  jand g08081(.dina(n25343), .dinb(n25341), .dout(n25344));
  jand g08082(.dina(n25344), .dinb(n266), .dout(n25345));
  jor  g08083(.dina(n25107), .dinb(n24913), .dout(n25346));
  jxor g08084(.dina(n25041), .dinb(n25040), .dout(n25347));
  jor  g08085(.dina(n25347), .dinb(n25248), .dout(n25348));
  jand g08086(.dina(n25348), .dinb(n25346), .dout(n25349));
  jand g08087(.dina(n25349), .dinb(n356), .dout(n25350));
  jor  g08088(.dina(n25107), .dinb(n24918), .dout(n25351));
  jxor g08089(.dina(n25038), .dinb(n25037), .dout(n25352));
  jor  g08090(.dina(n25352), .dinb(n25248), .dout(n25353));
  jand g08091(.dina(n25353), .dinb(n25351), .dout(n25354));
  jand g08092(.dina(n25354), .dinb(n355), .dout(n25355));
  jor  g08093(.dina(n25107), .dinb(n24923), .dout(n25356));
  jxor g08094(.dina(n25035), .dinb(n25034), .dout(n25357));
  jor  g08095(.dina(n25357), .dinb(n25248), .dout(n25358));
  jand g08096(.dina(n25358), .dinb(n25356), .dout(n25359));
  jand g08097(.dina(n25359), .dinb(n364), .dout(n25360));
  jor  g08098(.dina(n25107), .dinb(n24928), .dout(n25361));
  jxor g08099(.dina(n25032), .dinb(n25031), .dout(n25362));
  jor  g08100(.dina(n25362), .dinb(n25248), .dout(n25363));
  jand g08101(.dina(n25363), .dinb(n25361), .dout(n25364));
  jand g08102(.dina(n25364), .dinb(n361), .dout(n25365));
  jor  g08103(.dina(n25107), .dinb(n24933), .dout(n25366));
  jxor g08104(.dina(n25029), .dinb(n25028), .dout(n25367));
  jor  g08105(.dina(n25367), .dinb(n25248), .dout(n25368));
  jand g08106(.dina(n25368), .dinb(n25366), .dout(n25369));
  jand g08107(.dina(n25369), .dinb(n360), .dout(n25370));
  jor  g08108(.dina(n25107), .dinb(n24938), .dout(n25371));
  jxor g08109(.dina(n25026), .dinb(n25025), .dout(n25372));
  jor  g08110(.dina(n25372), .dinb(n25248), .dout(n25373));
  jand g08111(.dina(n25373), .dinb(n25371), .dout(n25374));
  jand g08112(.dina(n25374), .dinb(n363), .dout(n25375));
  jor  g08113(.dina(n25107), .dinb(n24943), .dout(n25376));
  jxor g08114(.dina(n25023), .dinb(n25022), .dout(n25377));
  jor  g08115(.dina(n25377), .dinb(n25248), .dout(n25378));
  jand g08116(.dina(n25378), .dinb(n25376), .dout(n25379));
  jand g08117(.dina(n25379), .dinb(n359), .dout(n25380));
  jor  g08118(.dina(n25107), .dinb(n24948), .dout(n25381));
  jxor g08119(.dina(n25020), .dinb(n25019), .dout(n25382));
  jor  g08120(.dina(n25382), .dinb(n25248), .dout(n25383));
  jand g08121(.dina(n25383), .dinb(n25381), .dout(n25384));
  jand g08122(.dina(n25384), .dinb(n369), .dout(n25385));
  jor  g08123(.dina(n25107), .dinb(n24953), .dout(n25386));
  jxor g08124(.dina(n25017), .dinb(n25016), .dout(n25387));
  jor  g08125(.dina(n25387), .dinb(n25248), .dout(n25388));
  jand g08126(.dina(n25388), .dinb(n25386), .dout(n25389));
  jand g08127(.dina(n25389), .dinb(n368), .dout(n25390));
  jor  g08128(.dina(n25107), .dinb(n24958), .dout(n25391));
  jxor g08129(.dina(n25014), .dinb(n25013), .dout(n25392));
  jor  g08130(.dina(n25392), .dinb(n25248), .dout(n25393));
  jand g08131(.dina(n25393), .dinb(n25391), .dout(n25394));
  jand g08132(.dina(n25394), .dinb(n367), .dout(n25395));
  jor  g08133(.dina(n25107), .dinb(n24963), .dout(n25396));
  jxor g08134(.dina(n25011), .dinb(n25010), .dout(n25397));
  jor  g08135(.dina(n25397), .dinb(n25248), .dout(n25398));
  jand g08136(.dina(n25398), .dinb(n25396), .dout(n25399));
  jand g08137(.dina(n25399), .dinb(n265), .dout(n25400));
  jor  g08138(.dina(n25107), .dinb(n24968), .dout(n25401));
  jxor g08139(.dina(n25008), .dinb(n25007), .dout(n25402));
  jor  g08140(.dina(n25402), .dinb(n25248), .dout(n25403));
  jand g08141(.dina(n25403), .dinb(n25401), .dout(n25404));
  jand g08142(.dina(n25404), .dinb(n378), .dout(n25405));
  jor  g08143(.dina(n25107), .dinb(n24973), .dout(n25406));
  jxor g08144(.dina(n25005), .dinb(n25004), .dout(n25407));
  jor  g08145(.dina(n25407), .dinb(n25248), .dout(n25408));
  jand g08146(.dina(n25408), .dinb(n25406), .dout(n25409));
  jand g08147(.dina(n25409), .dinb(n377), .dout(n25410));
  jor  g08148(.dina(n25107), .dinb(n24979), .dout(n25411));
  jxor g08149(.dina(n25002), .dinb(n25001), .dout(n25412));
  jor  g08150(.dina(n25412), .dinb(n25248), .dout(n25413));
  jand g08151(.dina(n25413), .dinb(n25411), .dout(n25414));
  jand g08152(.dina(n25414), .dinb(n376), .dout(n25415));
  jor  g08153(.dina(n25107), .dinb(n24984), .dout(n25416));
  jxor g08154(.dina(n24999), .dinb(n24998), .dout(n25417));
  jor  g08155(.dina(n25417), .dinb(n25248), .dout(n25418));
  jand g08156(.dina(n25418), .dinb(n25416), .dout(n25419));
  jand g08157(.dina(n25419), .dinb(n264), .dout(n25420));
  jand g08158(.dina(n25143), .dinb(n6026), .dout(n25421));
  jor  g08159(.dina(n25248), .dinb(n24997), .dout(n25422));
  jor  g08160(.dina(n25422), .dinb(n25421), .dout(n25423));
  jand g08161(.dina(n25248), .dinb(n24990), .dout(n25424));
  jnot g08162(.din(n25424), .dout(n25425));
  jand g08163(.dina(n25425), .dinb(n25423), .dout(n25426));
  jnot g08164(.din(n25426), .dout(n25427));
  jand g08165(.dina(n25427), .dinb(n386), .dout(n25428));
  jand g08166(.dina(n25107), .dinb(b0 ), .dout(n25429));
  jxor g08167(.dina(n25429), .dinb(a28 ), .dout(n25430));
  jand g08168(.dina(n25430), .dinb(n259), .dout(n25431));
  jxor g08169(.dina(n25429), .dinb(n6025), .dout(n25432));
  jxor g08170(.dina(n25432), .dinb(b1 ), .dout(n25433));
  jand g08171(.dina(n25433), .dinb(n6322), .dout(n25434));
  jor  g08172(.dina(n25434), .dinb(n25431), .dout(n25435));
  jxor g08173(.dina(n25426), .dinb(b2 ), .dout(n25436));
  jand g08174(.dina(n25436), .dinb(n25435), .dout(n25437));
  jor  g08175(.dina(n25437), .dinb(n25428), .dout(n25438));
  jxor g08176(.dina(n25419), .dinb(n264), .dout(n25439));
  jand g08177(.dina(n25439), .dinb(n25438), .dout(n25440));
  jor  g08178(.dina(n25440), .dinb(n25420), .dout(n25441));
  jxor g08179(.dina(n25414), .dinb(n376), .dout(n25442));
  jand g08180(.dina(n25442), .dinb(n25441), .dout(n25443));
  jor  g08181(.dina(n25443), .dinb(n25415), .dout(n25444));
  jxor g08182(.dina(n25409), .dinb(n377), .dout(n25445));
  jand g08183(.dina(n25445), .dinb(n25444), .dout(n25446));
  jor  g08184(.dina(n25446), .dinb(n25410), .dout(n25447));
  jxor g08185(.dina(n25404), .dinb(n378), .dout(n25448));
  jand g08186(.dina(n25448), .dinb(n25447), .dout(n25449));
  jor  g08187(.dina(n25449), .dinb(n25405), .dout(n25450));
  jxor g08188(.dina(n25399), .dinb(n265), .dout(n25451));
  jand g08189(.dina(n25451), .dinb(n25450), .dout(n25452));
  jor  g08190(.dina(n25452), .dinb(n25400), .dout(n25453));
  jxor g08191(.dina(n25394), .dinb(n367), .dout(n25454));
  jand g08192(.dina(n25454), .dinb(n25453), .dout(n25455));
  jor  g08193(.dina(n25455), .dinb(n25395), .dout(n25456));
  jxor g08194(.dina(n25389), .dinb(n368), .dout(n25457));
  jand g08195(.dina(n25457), .dinb(n25456), .dout(n25458));
  jor  g08196(.dina(n25458), .dinb(n25390), .dout(n25459));
  jxor g08197(.dina(n25384), .dinb(n369), .dout(n25460));
  jand g08198(.dina(n25460), .dinb(n25459), .dout(n25461));
  jor  g08199(.dina(n25461), .dinb(n25385), .dout(n25462));
  jxor g08200(.dina(n25379), .dinb(n359), .dout(n25463));
  jand g08201(.dina(n25463), .dinb(n25462), .dout(n25464));
  jor  g08202(.dina(n25464), .dinb(n25380), .dout(n25465));
  jxor g08203(.dina(n25374), .dinb(n363), .dout(n25466));
  jand g08204(.dina(n25466), .dinb(n25465), .dout(n25467));
  jor  g08205(.dina(n25467), .dinb(n25375), .dout(n25468));
  jxor g08206(.dina(n25369), .dinb(n360), .dout(n25469));
  jand g08207(.dina(n25469), .dinb(n25468), .dout(n25470));
  jor  g08208(.dina(n25470), .dinb(n25370), .dout(n25471));
  jxor g08209(.dina(n25364), .dinb(n361), .dout(n25472));
  jand g08210(.dina(n25472), .dinb(n25471), .dout(n25473));
  jor  g08211(.dina(n25473), .dinb(n25365), .dout(n25474));
  jxor g08212(.dina(n25359), .dinb(n364), .dout(n25475));
  jand g08213(.dina(n25475), .dinb(n25474), .dout(n25476));
  jor  g08214(.dina(n25476), .dinb(n25360), .dout(n25477));
  jxor g08215(.dina(n25354), .dinb(n355), .dout(n25478));
  jand g08216(.dina(n25478), .dinb(n25477), .dout(n25479));
  jor  g08217(.dina(n25479), .dinb(n25355), .dout(n25480));
  jxor g08218(.dina(n25349), .dinb(n356), .dout(n25481));
  jand g08219(.dina(n25481), .dinb(n25480), .dout(n25482));
  jor  g08220(.dina(n25482), .dinb(n25350), .dout(n25483));
  jxor g08221(.dina(n25344), .dinb(n266), .dout(n25484));
  jand g08222(.dina(n25484), .dinb(n25483), .dout(n25485));
  jor  g08223(.dina(n25485), .dinb(n25345), .dout(n25486));
  jxor g08224(.dina(n25339), .dinb(n267), .dout(n25487));
  jand g08225(.dina(n25487), .dinb(n25486), .dout(n25488));
  jor  g08226(.dina(n25488), .dinb(n25340), .dout(n25489));
  jxor g08227(.dina(n25334), .dinb(n347), .dout(n25490));
  jand g08228(.dina(n25490), .dinb(n25489), .dout(n25491));
  jor  g08229(.dina(n25491), .dinb(n25335), .dout(n25492));
  jxor g08230(.dina(n25329), .dinb(n348), .dout(n25493));
  jand g08231(.dina(n25493), .dinb(n25492), .dout(n25494));
  jor  g08232(.dina(n25494), .dinb(n25330), .dout(n25495));
  jxor g08233(.dina(n25324), .dinb(n349), .dout(n25496));
  jand g08234(.dina(n25496), .dinb(n25495), .dout(n25497));
  jor  g08235(.dina(n25497), .dinb(n25325), .dout(n25498));
  jxor g08236(.dina(n25319), .dinb(n268), .dout(n25499));
  jand g08237(.dina(n25499), .dinb(n25498), .dout(n25500));
  jor  g08238(.dina(n25500), .dinb(n25320), .dout(n25501));
  jxor g08239(.dina(n25314), .dinb(n274), .dout(n25502));
  jand g08240(.dina(n25502), .dinb(n25501), .dout(n25503));
  jor  g08241(.dina(n25503), .dinb(n25315), .dout(n25504));
  jxor g08242(.dina(n25309), .dinb(n269), .dout(n25505));
  jand g08243(.dina(n25505), .dinb(n25504), .dout(n25506));
  jor  g08244(.dina(n25506), .dinb(n25310), .dout(n25507));
  jxor g08245(.dina(n25304), .dinb(n270), .dout(n25508));
  jand g08246(.dina(n25508), .dinb(n25507), .dout(n25509));
  jor  g08247(.dina(n25509), .dinb(n25305), .dout(n25510));
  jxor g08248(.dina(n25299), .dinb(n271), .dout(n25511));
  jand g08249(.dina(n25511), .dinb(n25510), .dout(n25512));
  jor  g08250(.dina(n25512), .dinb(n25300), .dout(n25513));
  jxor g08251(.dina(n25294), .dinb(n338), .dout(n25514));
  jand g08252(.dina(n25514), .dinb(n25513), .dout(n25515));
  jor  g08253(.dina(n25515), .dinb(n25295), .dout(n25516));
  jxor g08254(.dina(n25289), .dinb(n339), .dout(n25517));
  jand g08255(.dina(n25517), .dinb(n25516), .dout(n25518));
  jor  g08256(.dina(n25518), .dinb(n25290), .dout(n25519));
  jxor g08257(.dina(n25284), .dinb(n340), .dout(n25520));
  jand g08258(.dina(n25520), .dinb(n25519), .dout(n25521));
  jor  g08259(.dina(n25521), .dinb(n25285), .dout(n25522));
  jxor g08260(.dina(n25279), .dinb(n275), .dout(n25523));
  jand g08261(.dina(n25523), .dinb(n25522), .dout(n25524));
  jor  g08262(.dina(n25524), .dinb(n25280), .dout(n25525));
  jxor g08263(.dina(n25274), .dinb(n331), .dout(n25526));
  jand g08264(.dina(n25526), .dinb(n25525), .dout(n25527));
  jor  g08265(.dina(n25527), .dinb(n25275), .dout(n25528));
  jxor g08266(.dina(n25269), .dinb(n332), .dout(n25529));
  jand g08267(.dina(n25529), .dinb(n25528), .dout(n25530));
  jor  g08268(.dina(n25530), .dinb(n25270), .dout(n25531));
  jxor g08269(.dina(n25264), .dinb(n333), .dout(n25532));
  jand g08270(.dina(n25532), .dinb(n25531), .dout(n25533));
  jor  g08271(.dina(n25533), .dinb(n25265), .dout(n25534));
  jxor g08272(.dina(n25251), .dinb(n276), .dout(n25535));
  jand g08273(.dina(n25535), .dinb(n25534), .dout(n25536));
  jor  g08274(.dina(n25536), .dinb(n25260), .dout(n25537));
  jand g08275(.dina(n25537), .dinb(n25259), .dout(n25538));
  jor  g08276(.dina(n25538), .dinb(n25256), .dout(n25539));
  jand g08277(.dina(n25539), .dinb(n408), .dout(n25540));
  jor  g08278(.dina(n25540), .dinb(n25251), .dout(n25541));
  jnot g08279(.din(n25540), .dout(n25542));
  jxor g08280(.dina(n25535), .dinb(n25534), .dout(n25543));
  jor  g08281(.dina(n25543), .dinb(n25542), .dout(n25544));
  jand g08282(.dina(n25544), .dinb(n25541), .dout(n25545));
  jand g08283(.dina(n25537), .dinb(n408), .dout(n25546));
  jand g08284(.dina(n25546), .dinb(n324), .dout(n25547));
  jor  g08285(.dina(n25547), .dinb(n25542), .dout(n25548));
  jand g08286(.dina(n25548), .dinb(n25255), .dout(n25549));
  jand g08287(.dina(n25549), .dinb(n325), .dout(n25550));
  jnot g08288(.din(n25549), .dout(n25551));
  jand g08289(.dina(n25551), .dinb(b37 ), .dout(n25552));
  jnot g08290(.din(n25552), .dout(n25553));
  jand g08291(.dina(n25545), .dinb(n324), .dout(n25554));
  jor  g08292(.dina(n25540), .dinb(n25264), .dout(n25555));
  jxor g08293(.dina(n25532), .dinb(n25531), .dout(n25556));
  jor  g08294(.dina(n25556), .dinb(n25542), .dout(n25557));
  jand g08295(.dina(n25557), .dinb(n25555), .dout(n25558));
  jand g08296(.dina(n25558), .dinb(n276), .dout(n25559));
  jor  g08297(.dina(n25540), .dinb(n25269), .dout(n25560));
  jxor g08298(.dina(n25529), .dinb(n25528), .dout(n25561));
  jor  g08299(.dina(n25561), .dinb(n25542), .dout(n25562));
  jand g08300(.dina(n25562), .dinb(n25560), .dout(n25563));
  jand g08301(.dina(n25563), .dinb(n333), .dout(n25564));
  jor  g08302(.dina(n25540), .dinb(n25274), .dout(n25565));
  jxor g08303(.dina(n25526), .dinb(n25525), .dout(n25566));
  jor  g08304(.dina(n25566), .dinb(n25542), .dout(n25567));
  jand g08305(.dina(n25567), .dinb(n25565), .dout(n25568));
  jand g08306(.dina(n25568), .dinb(n332), .dout(n25569));
  jor  g08307(.dina(n25540), .dinb(n25279), .dout(n25570));
  jxor g08308(.dina(n25523), .dinb(n25522), .dout(n25571));
  jor  g08309(.dina(n25571), .dinb(n25542), .dout(n25572));
  jand g08310(.dina(n25572), .dinb(n25570), .dout(n25573));
  jand g08311(.dina(n25573), .dinb(n331), .dout(n25574));
  jor  g08312(.dina(n25540), .dinb(n25284), .dout(n25575));
  jxor g08313(.dina(n25520), .dinb(n25519), .dout(n25576));
  jor  g08314(.dina(n25576), .dinb(n25542), .dout(n25577));
  jand g08315(.dina(n25577), .dinb(n25575), .dout(n25578));
  jand g08316(.dina(n25578), .dinb(n275), .dout(n25579));
  jor  g08317(.dina(n25540), .dinb(n25289), .dout(n25580));
  jxor g08318(.dina(n25517), .dinb(n25516), .dout(n25581));
  jor  g08319(.dina(n25581), .dinb(n25542), .dout(n25582));
  jand g08320(.dina(n25582), .dinb(n25580), .dout(n25583));
  jand g08321(.dina(n25583), .dinb(n340), .dout(n25584));
  jor  g08322(.dina(n25540), .dinb(n25294), .dout(n25585));
  jxor g08323(.dina(n25514), .dinb(n25513), .dout(n25586));
  jor  g08324(.dina(n25586), .dinb(n25542), .dout(n25587));
  jand g08325(.dina(n25587), .dinb(n25585), .dout(n25588));
  jand g08326(.dina(n25588), .dinb(n339), .dout(n25589));
  jor  g08327(.dina(n25540), .dinb(n25299), .dout(n25590));
  jxor g08328(.dina(n25511), .dinb(n25510), .dout(n25591));
  jor  g08329(.dina(n25591), .dinb(n25542), .dout(n25592));
  jand g08330(.dina(n25592), .dinb(n25590), .dout(n25593));
  jand g08331(.dina(n25593), .dinb(n338), .dout(n25594));
  jor  g08332(.dina(n25540), .dinb(n25304), .dout(n25595));
  jxor g08333(.dina(n25508), .dinb(n25507), .dout(n25596));
  jor  g08334(.dina(n25596), .dinb(n25542), .dout(n25597));
  jand g08335(.dina(n25597), .dinb(n25595), .dout(n25598));
  jand g08336(.dina(n25598), .dinb(n271), .dout(n25599));
  jor  g08337(.dina(n25540), .dinb(n25309), .dout(n25600));
  jxor g08338(.dina(n25505), .dinb(n25504), .dout(n25601));
  jor  g08339(.dina(n25601), .dinb(n25542), .dout(n25602));
  jand g08340(.dina(n25602), .dinb(n25600), .dout(n25603));
  jand g08341(.dina(n25603), .dinb(n270), .dout(n25604));
  jor  g08342(.dina(n25540), .dinb(n25314), .dout(n25605));
  jxor g08343(.dina(n25502), .dinb(n25501), .dout(n25606));
  jor  g08344(.dina(n25606), .dinb(n25542), .dout(n25607));
  jand g08345(.dina(n25607), .dinb(n25605), .dout(n25608));
  jand g08346(.dina(n25608), .dinb(n269), .dout(n25609));
  jor  g08347(.dina(n25540), .dinb(n25319), .dout(n25610));
  jxor g08348(.dina(n25499), .dinb(n25498), .dout(n25611));
  jor  g08349(.dina(n25611), .dinb(n25542), .dout(n25612));
  jand g08350(.dina(n25612), .dinb(n25610), .dout(n25613));
  jand g08351(.dina(n25613), .dinb(n274), .dout(n25614));
  jor  g08352(.dina(n25540), .dinb(n25324), .dout(n25615));
  jxor g08353(.dina(n25496), .dinb(n25495), .dout(n25616));
  jor  g08354(.dina(n25616), .dinb(n25542), .dout(n25617));
  jand g08355(.dina(n25617), .dinb(n25615), .dout(n25618));
  jand g08356(.dina(n25618), .dinb(n268), .dout(n25619));
  jor  g08357(.dina(n25540), .dinb(n25329), .dout(n25620));
  jxor g08358(.dina(n25493), .dinb(n25492), .dout(n25621));
  jor  g08359(.dina(n25621), .dinb(n25542), .dout(n25622));
  jand g08360(.dina(n25622), .dinb(n25620), .dout(n25623));
  jand g08361(.dina(n25623), .dinb(n349), .dout(n25624));
  jor  g08362(.dina(n25540), .dinb(n25334), .dout(n25625));
  jxor g08363(.dina(n25490), .dinb(n25489), .dout(n25626));
  jor  g08364(.dina(n25626), .dinb(n25542), .dout(n25627));
  jand g08365(.dina(n25627), .dinb(n25625), .dout(n25628));
  jand g08366(.dina(n25628), .dinb(n348), .dout(n25629));
  jor  g08367(.dina(n25540), .dinb(n25339), .dout(n25630));
  jxor g08368(.dina(n25487), .dinb(n25486), .dout(n25631));
  jor  g08369(.dina(n25631), .dinb(n25542), .dout(n25632));
  jand g08370(.dina(n25632), .dinb(n25630), .dout(n25633));
  jand g08371(.dina(n25633), .dinb(n347), .dout(n25634));
  jor  g08372(.dina(n25540), .dinb(n25344), .dout(n25635));
  jxor g08373(.dina(n25484), .dinb(n25483), .dout(n25636));
  jor  g08374(.dina(n25636), .dinb(n25542), .dout(n25637));
  jand g08375(.dina(n25637), .dinb(n25635), .dout(n25638));
  jand g08376(.dina(n25638), .dinb(n267), .dout(n25639));
  jor  g08377(.dina(n25540), .dinb(n25349), .dout(n25640));
  jxor g08378(.dina(n25481), .dinb(n25480), .dout(n25641));
  jor  g08379(.dina(n25641), .dinb(n25542), .dout(n25642));
  jand g08380(.dina(n25642), .dinb(n25640), .dout(n25643));
  jand g08381(.dina(n25643), .dinb(n266), .dout(n25644));
  jor  g08382(.dina(n25540), .dinb(n25354), .dout(n25645));
  jxor g08383(.dina(n25478), .dinb(n25477), .dout(n25646));
  jor  g08384(.dina(n25646), .dinb(n25542), .dout(n25647));
  jand g08385(.dina(n25647), .dinb(n25645), .dout(n25648));
  jand g08386(.dina(n25648), .dinb(n356), .dout(n25649));
  jor  g08387(.dina(n25540), .dinb(n25359), .dout(n25650));
  jxor g08388(.dina(n25475), .dinb(n25474), .dout(n25651));
  jor  g08389(.dina(n25651), .dinb(n25542), .dout(n25652));
  jand g08390(.dina(n25652), .dinb(n25650), .dout(n25653));
  jand g08391(.dina(n25653), .dinb(n355), .dout(n25654));
  jor  g08392(.dina(n25540), .dinb(n25364), .dout(n25655));
  jxor g08393(.dina(n25472), .dinb(n25471), .dout(n25656));
  jor  g08394(.dina(n25656), .dinb(n25542), .dout(n25657));
  jand g08395(.dina(n25657), .dinb(n25655), .dout(n25658));
  jand g08396(.dina(n25658), .dinb(n364), .dout(n25659));
  jor  g08397(.dina(n25540), .dinb(n25369), .dout(n25660));
  jxor g08398(.dina(n25469), .dinb(n25468), .dout(n25661));
  jor  g08399(.dina(n25661), .dinb(n25542), .dout(n25662));
  jand g08400(.dina(n25662), .dinb(n25660), .dout(n25663));
  jand g08401(.dina(n25663), .dinb(n361), .dout(n25664));
  jor  g08402(.dina(n25540), .dinb(n25374), .dout(n25665));
  jxor g08403(.dina(n25466), .dinb(n25465), .dout(n25666));
  jor  g08404(.dina(n25666), .dinb(n25542), .dout(n25667));
  jand g08405(.dina(n25667), .dinb(n25665), .dout(n25668));
  jand g08406(.dina(n25668), .dinb(n360), .dout(n25669));
  jor  g08407(.dina(n25540), .dinb(n25379), .dout(n25670));
  jxor g08408(.dina(n25463), .dinb(n25462), .dout(n25671));
  jor  g08409(.dina(n25671), .dinb(n25542), .dout(n25672));
  jand g08410(.dina(n25672), .dinb(n25670), .dout(n25673));
  jand g08411(.dina(n25673), .dinb(n363), .dout(n25674));
  jor  g08412(.dina(n25540), .dinb(n25384), .dout(n25675));
  jxor g08413(.dina(n25460), .dinb(n25459), .dout(n25676));
  jor  g08414(.dina(n25676), .dinb(n25542), .dout(n25677));
  jand g08415(.dina(n25677), .dinb(n25675), .dout(n25678));
  jand g08416(.dina(n25678), .dinb(n359), .dout(n25679));
  jor  g08417(.dina(n25540), .dinb(n25389), .dout(n25680));
  jxor g08418(.dina(n25457), .dinb(n25456), .dout(n25681));
  jor  g08419(.dina(n25681), .dinb(n25542), .dout(n25682));
  jand g08420(.dina(n25682), .dinb(n25680), .dout(n25683));
  jand g08421(.dina(n25683), .dinb(n369), .dout(n25684));
  jor  g08422(.dina(n25540), .dinb(n25394), .dout(n25685));
  jxor g08423(.dina(n25454), .dinb(n25453), .dout(n25686));
  jor  g08424(.dina(n25686), .dinb(n25542), .dout(n25687));
  jand g08425(.dina(n25687), .dinb(n25685), .dout(n25688));
  jand g08426(.dina(n25688), .dinb(n368), .dout(n25689));
  jor  g08427(.dina(n25540), .dinb(n25399), .dout(n25690));
  jxor g08428(.dina(n25451), .dinb(n25450), .dout(n25691));
  jor  g08429(.dina(n25691), .dinb(n25542), .dout(n25692));
  jand g08430(.dina(n25692), .dinb(n25690), .dout(n25693));
  jand g08431(.dina(n25693), .dinb(n367), .dout(n25694));
  jor  g08432(.dina(n25540), .dinb(n25404), .dout(n25695));
  jxor g08433(.dina(n25448), .dinb(n25447), .dout(n25696));
  jor  g08434(.dina(n25696), .dinb(n25542), .dout(n25697));
  jand g08435(.dina(n25697), .dinb(n25695), .dout(n25698));
  jand g08436(.dina(n25698), .dinb(n265), .dout(n25699));
  jor  g08437(.dina(n25540), .dinb(n25409), .dout(n25700));
  jxor g08438(.dina(n25445), .dinb(n25444), .dout(n25701));
  jor  g08439(.dina(n25701), .dinb(n25542), .dout(n25702));
  jand g08440(.dina(n25702), .dinb(n25700), .dout(n25703));
  jand g08441(.dina(n25703), .dinb(n378), .dout(n25704));
  jor  g08442(.dina(n25540), .dinb(n25414), .dout(n25705));
  jxor g08443(.dina(n25442), .dinb(n25441), .dout(n25706));
  jor  g08444(.dina(n25706), .dinb(n25542), .dout(n25707));
  jand g08445(.dina(n25707), .dinb(n25705), .dout(n25708));
  jand g08446(.dina(n25708), .dinb(n377), .dout(n25709));
  jor  g08447(.dina(n25540), .dinb(n25419), .dout(n25710));
  jxor g08448(.dina(n25439), .dinb(n25438), .dout(n25711));
  jor  g08449(.dina(n25711), .dinb(n25542), .dout(n25712));
  jand g08450(.dina(n25712), .dinb(n25710), .dout(n25713));
  jand g08451(.dina(n25713), .dinb(n376), .dout(n25714));
  jor  g08452(.dina(n25540), .dinb(n25427), .dout(n25715));
  jxor g08453(.dina(n25436), .dinb(n25435), .dout(n25716));
  jor  g08454(.dina(n25716), .dinb(n25542), .dout(n25717));
  jand g08455(.dina(n25717), .dinb(n25715), .dout(n25718));
  jand g08456(.dina(n25718), .dinb(n264), .dout(n25719));
  jor  g08457(.dina(n25540), .dinb(n25430), .dout(n25720));
  jxor g08458(.dina(n25433), .dinb(n6322), .dout(n25721));
  jor  g08459(.dina(n25721), .dinb(n25542), .dout(n25722));
  jand g08460(.dina(n25722), .dinb(n25720), .dout(n25723));
  jand g08461(.dina(n25723), .dinb(n386), .dout(n25724));
  jnot g08462(.din(n6653), .dout(n25725));
  jnot g08463(.din(n25256), .dout(n25726));
  jnot g08464(.din(n25260), .dout(n25727));
  jnot g08465(.din(n25265), .dout(n25728));
  jnot g08466(.din(n25270), .dout(n25729));
  jnot g08467(.din(n25275), .dout(n25730));
  jnot g08468(.din(n25280), .dout(n25731));
  jnot g08469(.din(n25285), .dout(n25732));
  jnot g08470(.din(n25290), .dout(n25733));
  jnot g08471(.din(n25295), .dout(n25734));
  jnot g08472(.din(n25300), .dout(n25735));
  jnot g08473(.din(n25305), .dout(n25736));
  jnot g08474(.din(n25310), .dout(n25737));
  jnot g08475(.din(n25315), .dout(n25738));
  jnot g08476(.din(n25320), .dout(n25739));
  jnot g08477(.din(n25325), .dout(n25740));
  jnot g08478(.din(n25330), .dout(n25741));
  jnot g08479(.din(n25335), .dout(n25742));
  jnot g08480(.din(n25340), .dout(n25743));
  jnot g08481(.din(n25345), .dout(n25744));
  jnot g08482(.din(n25350), .dout(n25745));
  jnot g08483(.din(n25355), .dout(n25746));
  jnot g08484(.din(n25360), .dout(n25747));
  jnot g08485(.din(n25365), .dout(n25748));
  jnot g08486(.din(n25370), .dout(n25749));
  jnot g08487(.din(n25375), .dout(n25750));
  jnot g08488(.din(n25380), .dout(n25751));
  jnot g08489(.din(n25385), .dout(n25752));
  jnot g08490(.din(n25390), .dout(n25753));
  jnot g08491(.din(n25395), .dout(n25754));
  jnot g08492(.din(n25400), .dout(n25755));
  jnot g08493(.din(n25405), .dout(n25756));
  jnot g08494(.din(n25410), .dout(n25757));
  jnot g08495(.din(n25415), .dout(n25758));
  jnot g08496(.din(n25420), .dout(n25759));
  jnot g08497(.din(n25428), .dout(n25760));
  jnot g08498(.din(n25431), .dout(n25761));
  jxor g08499(.dina(n25432), .dinb(n259), .dout(n25762));
  jor  g08500(.dina(n25762), .dinb(n6321), .dout(n25763));
  jand g08501(.dina(n25763), .dinb(n25761), .dout(n25764));
  jnot g08502(.din(n25436), .dout(n25765));
  jor  g08503(.dina(n25765), .dinb(n25764), .dout(n25766));
  jand g08504(.dina(n25766), .dinb(n25760), .dout(n25767));
  jnot g08505(.din(n25439), .dout(n25768));
  jor  g08506(.dina(n25768), .dinb(n25767), .dout(n25769));
  jand g08507(.dina(n25769), .dinb(n25759), .dout(n25770));
  jnot g08508(.din(n25442), .dout(n25771));
  jor  g08509(.dina(n25771), .dinb(n25770), .dout(n25772));
  jand g08510(.dina(n25772), .dinb(n25758), .dout(n25773));
  jnot g08511(.din(n25445), .dout(n25774));
  jor  g08512(.dina(n25774), .dinb(n25773), .dout(n25775));
  jand g08513(.dina(n25775), .dinb(n25757), .dout(n25776));
  jnot g08514(.din(n25448), .dout(n25777));
  jor  g08515(.dina(n25777), .dinb(n25776), .dout(n25778));
  jand g08516(.dina(n25778), .dinb(n25756), .dout(n25779));
  jnot g08517(.din(n25451), .dout(n25780));
  jor  g08518(.dina(n25780), .dinb(n25779), .dout(n25781));
  jand g08519(.dina(n25781), .dinb(n25755), .dout(n25782));
  jnot g08520(.din(n25454), .dout(n25783));
  jor  g08521(.dina(n25783), .dinb(n25782), .dout(n25784));
  jand g08522(.dina(n25784), .dinb(n25754), .dout(n25785));
  jnot g08523(.din(n25457), .dout(n25786));
  jor  g08524(.dina(n25786), .dinb(n25785), .dout(n25787));
  jand g08525(.dina(n25787), .dinb(n25753), .dout(n25788));
  jnot g08526(.din(n25460), .dout(n25789));
  jor  g08527(.dina(n25789), .dinb(n25788), .dout(n25790));
  jand g08528(.dina(n25790), .dinb(n25752), .dout(n25791));
  jnot g08529(.din(n25463), .dout(n25792));
  jor  g08530(.dina(n25792), .dinb(n25791), .dout(n25793));
  jand g08531(.dina(n25793), .dinb(n25751), .dout(n25794));
  jnot g08532(.din(n25466), .dout(n25795));
  jor  g08533(.dina(n25795), .dinb(n25794), .dout(n25796));
  jand g08534(.dina(n25796), .dinb(n25750), .dout(n25797));
  jnot g08535(.din(n25469), .dout(n25798));
  jor  g08536(.dina(n25798), .dinb(n25797), .dout(n25799));
  jand g08537(.dina(n25799), .dinb(n25749), .dout(n25800));
  jnot g08538(.din(n25472), .dout(n25801));
  jor  g08539(.dina(n25801), .dinb(n25800), .dout(n25802));
  jand g08540(.dina(n25802), .dinb(n25748), .dout(n25803));
  jnot g08541(.din(n25475), .dout(n25804));
  jor  g08542(.dina(n25804), .dinb(n25803), .dout(n25805));
  jand g08543(.dina(n25805), .dinb(n25747), .dout(n25806));
  jnot g08544(.din(n25478), .dout(n25807));
  jor  g08545(.dina(n25807), .dinb(n25806), .dout(n25808));
  jand g08546(.dina(n25808), .dinb(n25746), .dout(n25809));
  jnot g08547(.din(n25481), .dout(n25810));
  jor  g08548(.dina(n25810), .dinb(n25809), .dout(n25811));
  jand g08549(.dina(n25811), .dinb(n25745), .dout(n25812));
  jnot g08550(.din(n25484), .dout(n25813));
  jor  g08551(.dina(n25813), .dinb(n25812), .dout(n25814));
  jand g08552(.dina(n25814), .dinb(n25744), .dout(n25815));
  jnot g08553(.din(n25487), .dout(n25816));
  jor  g08554(.dina(n25816), .dinb(n25815), .dout(n25817));
  jand g08555(.dina(n25817), .dinb(n25743), .dout(n25818));
  jnot g08556(.din(n25490), .dout(n25819));
  jor  g08557(.dina(n25819), .dinb(n25818), .dout(n25820));
  jand g08558(.dina(n25820), .dinb(n25742), .dout(n25821));
  jnot g08559(.din(n25493), .dout(n25822));
  jor  g08560(.dina(n25822), .dinb(n25821), .dout(n25823));
  jand g08561(.dina(n25823), .dinb(n25741), .dout(n25824));
  jnot g08562(.din(n25496), .dout(n25825));
  jor  g08563(.dina(n25825), .dinb(n25824), .dout(n25826));
  jand g08564(.dina(n25826), .dinb(n25740), .dout(n25827));
  jnot g08565(.din(n25499), .dout(n25828));
  jor  g08566(.dina(n25828), .dinb(n25827), .dout(n25829));
  jand g08567(.dina(n25829), .dinb(n25739), .dout(n25830));
  jnot g08568(.din(n25502), .dout(n25831));
  jor  g08569(.dina(n25831), .dinb(n25830), .dout(n25832));
  jand g08570(.dina(n25832), .dinb(n25738), .dout(n25833));
  jnot g08571(.din(n25505), .dout(n25834));
  jor  g08572(.dina(n25834), .dinb(n25833), .dout(n25835));
  jand g08573(.dina(n25835), .dinb(n25737), .dout(n25836));
  jnot g08574(.din(n25508), .dout(n25837));
  jor  g08575(.dina(n25837), .dinb(n25836), .dout(n25838));
  jand g08576(.dina(n25838), .dinb(n25736), .dout(n25839));
  jnot g08577(.din(n25511), .dout(n25840));
  jor  g08578(.dina(n25840), .dinb(n25839), .dout(n25841));
  jand g08579(.dina(n25841), .dinb(n25735), .dout(n25842));
  jnot g08580(.din(n25514), .dout(n25843));
  jor  g08581(.dina(n25843), .dinb(n25842), .dout(n25844));
  jand g08582(.dina(n25844), .dinb(n25734), .dout(n25845));
  jnot g08583(.din(n25517), .dout(n25846));
  jor  g08584(.dina(n25846), .dinb(n25845), .dout(n25847));
  jand g08585(.dina(n25847), .dinb(n25733), .dout(n25848));
  jnot g08586(.din(n25520), .dout(n25849));
  jor  g08587(.dina(n25849), .dinb(n25848), .dout(n25850));
  jand g08588(.dina(n25850), .dinb(n25732), .dout(n25851));
  jnot g08589(.din(n25523), .dout(n25852));
  jor  g08590(.dina(n25852), .dinb(n25851), .dout(n25853));
  jand g08591(.dina(n25853), .dinb(n25731), .dout(n25854));
  jnot g08592(.din(n25526), .dout(n25855));
  jor  g08593(.dina(n25855), .dinb(n25854), .dout(n25856));
  jand g08594(.dina(n25856), .dinb(n25730), .dout(n25857));
  jnot g08595(.din(n25529), .dout(n25858));
  jor  g08596(.dina(n25858), .dinb(n25857), .dout(n25859));
  jand g08597(.dina(n25859), .dinb(n25729), .dout(n25860));
  jnot g08598(.din(n25532), .dout(n25861));
  jor  g08599(.dina(n25861), .dinb(n25860), .dout(n25862));
  jand g08600(.dina(n25862), .dinb(n25728), .dout(n25863));
  jnot g08601(.din(n25535), .dout(n25864));
  jor  g08602(.dina(n25864), .dinb(n25863), .dout(n25865));
  jand g08603(.dina(n25865), .dinb(n25727), .dout(n25866));
  jor  g08604(.dina(n25866), .dinb(n25258), .dout(n25867));
  jand g08605(.dina(n25867), .dinb(n25726), .dout(n25868));
  jor  g08606(.dina(n25868), .dinb(n25725), .dout(n25869));
  jand g08607(.dina(n25869), .dinb(a27 ), .dout(n25870));
  jnot g08608(.din(n6656), .dout(n25871));
  jor  g08609(.dina(n25868), .dinb(n25871), .dout(n25872));
  jnot g08610(.din(n25872), .dout(n25873));
  jor  g08611(.dina(n25873), .dinb(n25870), .dout(n25874));
  jand g08612(.dina(n25874), .dinb(n259), .dout(n25875));
  jand g08613(.dina(n25539), .dinb(n6653), .dout(n25876));
  jor  g08614(.dina(n25876), .dinb(n6320), .dout(n25877));
  jand g08615(.dina(n25872), .dinb(n25877), .dout(n25878));
  jxor g08616(.dina(n25878), .dinb(b1 ), .dout(n25879));
  jand g08617(.dina(n25879), .dinb(n6812), .dout(n25880));
  jor  g08618(.dina(n25880), .dinb(n25875), .dout(n25881));
  jxor g08619(.dina(n25723), .dinb(n386), .dout(n25882));
  jand g08620(.dina(n25882), .dinb(n25881), .dout(n25883));
  jor  g08621(.dina(n25883), .dinb(n25724), .dout(n25884));
  jxor g08622(.dina(n25718), .dinb(n264), .dout(n25885));
  jand g08623(.dina(n25885), .dinb(n25884), .dout(n25886));
  jor  g08624(.dina(n25886), .dinb(n25719), .dout(n25887));
  jxor g08625(.dina(n25713), .dinb(n376), .dout(n25888));
  jand g08626(.dina(n25888), .dinb(n25887), .dout(n25889));
  jor  g08627(.dina(n25889), .dinb(n25714), .dout(n25890));
  jxor g08628(.dina(n25708), .dinb(n377), .dout(n25891));
  jand g08629(.dina(n25891), .dinb(n25890), .dout(n25892));
  jor  g08630(.dina(n25892), .dinb(n25709), .dout(n25893));
  jxor g08631(.dina(n25703), .dinb(n378), .dout(n25894));
  jand g08632(.dina(n25894), .dinb(n25893), .dout(n25895));
  jor  g08633(.dina(n25895), .dinb(n25704), .dout(n25896));
  jxor g08634(.dina(n25698), .dinb(n265), .dout(n25897));
  jand g08635(.dina(n25897), .dinb(n25896), .dout(n25898));
  jor  g08636(.dina(n25898), .dinb(n25699), .dout(n25899));
  jxor g08637(.dina(n25693), .dinb(n367), .dout(n25900));
  jand g08638(.dina(n25900), .dinb(n25899), .dout(n25901));
  jor  g08639(.dina(n25901), .dinb(n25694), .dout(n25902));
  jxor g08640(.dina(n25688), .dinb(n368), .dout(n25903));
  jand g08641(.dina(n25903), .dinb(n25902), .dout(n25904));
  jor  g08642(.dina(n25904), .dinb(n25689), .dout(n25905));
  jxor g08643(.dina(n25683), .dinb(n369), .dout(n25906));
  jand g08644(.dina(n25906), .dinb(n25905), .dout(n25907));
  jor  g08645(.dina(n25907), .dinb(n25684), .dout(n25908));
  jxor g08646(.dina(n25678), .dinb(n359), .dout(n25909));
  jand g08647(.dina(n25909), .dinb(n25908), .dout(n25910));
  jor  g08648(.dina(n25910), .dinb(n25679), .dout(n25911));
  jxor g08649(.dina(n25673), .dinb(n363), .dout(n25912));
  jand g08650(.dina(n25912), .dinb(n25911), .dout(n25913));
  jor  g08651(.dina(n25913), .dinb(n25674), .dout(n25914));
  jxor g08652(.dina(n25668), .dinb(n360), .dout(n25915));
  jand g08653(.dina(n25915), .dinb(n25914), .dout(n25916));
  jor  g08654(.dina(n25916), .dinb(n25669), .dout(n25917));
  jxor g08655(.dina(n25663), .dinb(n361), .dout(n25918));
  jand g08656(.dina(n25918), .dinb(n25917), .dout(n25919));
  jor  g08657(.dina(n25919), .dinb(n25664), .dout(n25920));
  jxor g08658(.dina(n25658), .dinb(n364), .dout(n25921));
  jand g08659(.dina(n25921), .dinb(n25920), .dout(n25922));
  jor  g08660(.dina(n25922), .dinb(n25659), .dout(n25923));
  jxor g08661(.dina(n25653), .dinb(n355), .dout(n25924));
  jand g08662(.dina(n25924), .dinb(n25923), .dout(n25925));
  jor  g08663(.dina(n25925), .dinb(n25654), .dout(n25926));
  jxor g08664(.dina(n25648), .dinb(n356), .dout(n25927));
  jand g08665(.dina(n25927), .dinb(n25926), .dout(n25928));
  jor  g08666(.dina(n25928), .dinb(n25649), .dout(n25929));
  jxor g08667(.dina(n25643), .dinb(n266), .dout(n25930));
  jand g08668(.dina(n25930), .dinb(n25929), .dout(n25931));
  jor  g08669(.dina(n25931), .dinb(n25644), .dout(n25932));
  jxor g08670(.dina(n25638), .dinb(n267), .dout(n25933));
  jand g08671(.dina(n25933), .dinb(n25932), .dout(n25934));
  jor  g08672(.dina(n25934), .dinb(n25639), .dout(n25935));
  jxor g08673(.dina(n25633), .dinb(n347), .dout(n25936));
  jand g08674(.dina(n25936), .dinb(n25935), .dout(n25937));
  jor  g08675(.dina(n25937), .dinb(n25634), .dout(n25938));
  jxor g08676(.dina(n25628), .dinb(n348), .dout(n25939));
  jand g08677(.dina(n25939), .dinb(n25938), .dout(n25940));
  jor  g08678(.dina(n25940), .dinb(n25629), .dout(n25941));
  jxor g08679(.dina(n25623), .dinb(n349), .dout(n25942));
  jand g08680(.dina(n25942), .dinb(n25941), .dout(n25943));
  jor  g08681(.dina(n25943), .dinb(n25624), .dout(n25944));
  jxor g08682(.dina(n25618), .dinb(n268), .dout(n25945));
  jand g08683(.dina(n25945), .dinb(n25944), .dout(n25946));
  jor  g08684(.dina(n25946), .dinb(n25619), .dout(n25947));
  jxor g08685(.dina(n25613), .dinb(n274), .dout(n25948));
  jand g08686(.dina(n25948), .dinb(n25947), .dout(n25949));
  jor  g08687(.dina(n25949), .dinb(n25614), .dout(n25950));
  jxor g08688(.dina(n25608), .dinb(n269), .dout(n25951));
  jand g08689(.dina(n25951), .dinb(n25950), .dout(n25952));
  jor  g08690(.dina(n25952), .dinb(n25609), .dout(n25953));
  jxor g08691(.dina(n25603), .dinb(n270), .dout(n25954));
  jand g08692(.dina(n25954), .dinb(n25953), .dout(n25955));
  jor  g08693(.dina(n25955), .dinb(n25604), .dout(n25956));
  jxor g08694(.dina(n25598), .dinb(n271), .dout(n25957));
  jand g08695(.dina(n25957), .dinb(n25956), .dout(n25958));
  jor  g08696(.dina(n25958), .dinb(n25599), .dout(n25959));
  jxor g08697(.dina(n25593), .dinb(n338), .dout(n25960));
  jand g08698(.dina(n25960), .dinb(n25959), .dout(n25961));
  jor  g08699(.dina(n25961), .dinb(n25594), .dout(n25962));
  jxor g08700(.dina(n25588), .dinb(n339), .dout(n25963));
  jand g08701(.dina(n25963), .dinb(n25962), .dout(n25964));
  jor  g08702(.dina(n25964), .dinb(n25589), .dout(n25965));
  jxor g08703(.dina(n25583), .dinb(n340), .dout(n25966));
  jand g08704(.dina(n25966), .dinb(n25965), .dout(n25967));
  jor  g08705(.dina(n25967), .dinb(n25584), .dout(n25968));
  jxor g08706(.dina(n25578), .dinb(n275), .dout(n25969));
  jand g08707(.dina(n25969), .dinb(n25968), .dout(n25970));
  jor  g08708(.dina(n25970), .dinb(n25579), .dout(n25971));
  jxor g08709(.dina(n25573), .dinb(n331), .dout(n25972));
  jand g08710(.dina(n25972), .dinb(n25971), .dout(n25973));
  jor  g08711(.dina(n25973), .dinb(n25574), .dout(n25974));
  jxor g08712(.dina(n25568), .dinb(n332), .dout(n25975));
  jand g08713(.dina(n25975), .dinb(n25974), .dout(n25976));
  jor  g08714(.dina(n25976), .dinb(n25569), .dout(n25977));
  jxor g08715(.dina(n25563), .dinb(n333), .dout(n25978));
  jand g08716(.dina(n25978), .dinb(n25977), .dout(n25979));
  jor  g08717(.dina(n25979), .dinb(n25564), .dout(n25980));
  jxor g08718(.dina(n25558), .dinb(n276), .dout(n25981));
  jand g08719(.dina(n25981), .dinb(n25980), .dout(n25982));
  jor  g08720(.dina(n25982), .dinb(n25559), .dout(n25983));
  jxor g08721(.dina(n25545), .dinb(n324), .dout(n25984));
  jand g08722(.dina(n25984), .dinb(n25983), .dout(n25985));
  jor  g08723(.dina(n25985), .dinb(n25554), .dout(n25986));
  jand g08724(.dina(n25986), .dinb(n25553), .dout(n25987));
  jor  g08725(.dina(n25987), .dinb(n25550), .dout(n25988));
  jand g08726(.dina(n25988), .dinb(n6436), .dout(n25989));
  jor  g08727(.dina(n25989), .dinb(n25545), .dout(n25990));
  jnot g08728(.din(n25550), .dout(n25991));
  jnot g08729(.din(n25554), .dout(n25992));
  jnot g08730(.din(n25559), .dout(n25993));
  jnot g08731(.din(n25564), .dout(n25994));
  jnot g08732(.din(n25569), .dout(n25995));
  jnot g08733(.din(n25574), .dout(n25996));
  jnot g08734(.din(n25579), .dout(n25997));
  jnot g08735(.din(n25584), .dout(n25998));
  jnot g08736(.din(n25589), .dout(n25999));
  jnot g08737(.din(n25594), .dout(n26000));
  jnot g08738(.din(n25599), .dout(n26001));
  jnot g08739(.din(n25604), .dout(n26002));
  jnot g08740(.din(n25609), .dout(n26003));
  jnot g08741(.din(n25614), .dout(n26004));
  jnot g08742(.din(n25619), .dout(n26005));
  jnot g08743(.din(n25624), .dout(n26006));
  jnot g08744(.din(n25629), .dout(n26007));
  jnot g08745(.din(n25634), .dout(n26008));
  jnot g08746(.din(n25639), .dout(n26009));
  jnot g08747(.din(n25644), .dout(n26010));
  jnot g08748(.din(n25649), .dout(n26011));
  jnot g08749(.din(n25654), .dout(n26012));
  jnot g08750(.din(n25659), .dout(n26013));
  jnot g08751(.din(n25664), .dout(n26014));
  jnot g08752(.din(n25669), .dout(n26015));
  jnot g08753(.din(n25674), .dout(n26016));
  jnot g08754(.din(n25679), .dout(n26017));
  jnot g08755(.din(n25684), .dout(n26018));
  jnot g08756(.din(n25689), .dout(n26019));
  jnot g08757(.din(n25694), .dout(n26020));
  jnot g08758(.din(n25699), .dout(n26021));
  jnot g08759(.din(n25704), .dout(n26022));
  jnot g08760(.din(n25709), .dout(n26023));
  jnot g08761(.din(n25714), .dout(n26024));
  jnot g08762(.din(n25719), .dout(n26025));
  jnot g08763(.din(n25724), .dout(n26026));
  jor  g08764(.dina(n25878), .dinb(b1 ), .dout(n26027));
  jxor g08765(.dina(n25878), .dinb(n259), .dout(n26028));
  jor  g08766(.dina(n26028), .dinb(n6662), .dout(n26029));
  jand g08767(.dina(n26029), .dinb(n26027), .dout(n26030));
  jxor g08768(.dina(n25723), .dinb(b2 ), .dout(n26031));
  jor  g08769(.dina(n26031), .dinb(n26030), .dout(n26032));
  jand g08770(.dina(n26032), .dinb(n26026), .dout(n26033));
  jnot g08771(.din(n25885), .dout(n26034));
  jor  g08772(.dina(n26034), .dinb(n26033), .dout(n26035));
  jand g08773(.dina(n26035), .dinb(n26025), .dout(n26036));
  jnot g08774(.din(n25888), .dout(n26037));
  jor  g08775(.dina(n26037), .dinb(n26036), .dout(n26038));
  jand g08776(.dina(n26038), .dinb(n26024), .dout(n26039));
  jnot g08777(.din(n25891), .dout(n26040));
  jor  g08778(.dina(n26040), .dinb(n26039), .dout(n26041));
  jand g08779(.dina(n26041), .dinb(n26023), .dout(n26042));
  jnot g08780(.din(n25894), .dout(n26043));
  jor  g08781(.dina(n26043), .dinb(n26042), .dout(n26044));
  jand g08782(.dina(n26044), .dinb(n26022), .dout(n26045));
  jnot g08783(.din(n25897), .dout(n26046));
  jor  g08784(.dina(n26046), .dinb(n26045), .dout(n26047));
  jand g08785(.dina(n26047), .dinb(n26021), .dout(n26048));
  jnot g08786(.din(n25900), .dout(n26049));
  jor  g08787(.dina(n26049), .dinb(n26048), .dout(n26050));
  jand g08788(.dina(n26050), .dinb(n26020), .dout(n26051));
  jnot g08789(.din(n25903), .dout(n26052));
  jor  g08790(.dina(n26052), .dinb(n26051), .dout(n26053));
  jand g08791(.dina(n26053), .dinb(n26019), .dout(n26054));
  jnot g08792(.din(n25906), .dout(n26055));
  jor  g08793(.dina(n26055), .dinb(n26054), .dout(n26056));
  jand g08794(.dina(n26056), .dinb(n26018), .dout(n26057));
  jnot g08795(.din(n25909), .dout(n26058));
  jor  g08796(.dina(n26058), .dinb(n26057), .dout(n26059));
  jand g08797(.dina(n26059), .dinb(n26017), .dout(n26060));
  jnot g08798(.din(n25912), .dout(n26061));
  jor  g08799(.dina(n26061), .dinb(n26060), .dout(n26062));
  jand g08800(.dina(n26062), .dinb(n26016), .dout(n26063));
  jnot g08801(.din(n25915), .dout(n26064));
  jor  g08802(.dina(n26064), .dinb(n26063), .dout(n26065));
  jand g08803(.dina(n26065), .dinb(n26015), .dout(n26066));
  jnot g08804(.din(n25918), .dout(n26067));
  jor  g08805(.dina(n26067), .dinb(n26066), .dout(n26068));
  jand g08806(.dina(n26068), .dinb(n26014), .dout(n26069));
  jnot g08807(.din(n25921), .dout(n26070));
  jor  g08808(.dina(n26070), .dinb(n26069), .dout(n26071));
  jand g08809(.dina(n26071), .dinb(n26013), .dout(n26072));
  jnot g08810(.din(n25924), .dout(n26073));
  jor  g08811(.dina(n26073), .dinb(n26072), .dout(n26074));
  jand g08812(.dina(n26074), .dinb(n26012), .dout(n26075));
  jnot g08813(.din(n25927), .dout(n26076));
  jor  g08814(.dina(n26076), .dinb(n26075), .dout(n26077));
  jand g08815(.dina(n26077), .dinb(n26011), .dout(n26078));
  jnot g08816(.din(n25930), .dout(n26079));
  jor  g08817(.dina(n26079), .dinb(n26078), .dout(n26080));
  jand g08818(.dina(n26080), .dinb(n26010), .dout(n26081));
  jnot g08819(.din(n25933), .dout(n26082));
  jor  g08820(.dina(n26082), .dinb(n26081), .dout(n26083));
  jand g08821(.dina(n26083), .dinb(n26009), .dout(n26084));
  jnot g08822(.din(n25936), .dout(n26085));
  jor  g08823(.dina(n26085), .dinb(n26084), .dout(n26086));
  jand g08824(.dina(n26086), .dinb(n26008), .dout(n26087));
  jnot g08825(.din(n25939), .dout(n26088));
  jor  g08826(.dina(n26088), .dinb(n26087), .dout(n26089));
  jand g08827(.dina(n26089), .dinb(n26007), .dout(n26090));
  jnot g08828(.din(n25942), .dout(n26091));
  jor  g08829(.dina(n26091), .dinb(n26090), .dout(n26092));
  jand g08830(.dina(n26092), .dinb(n26006), .dout(n26093));
  jnot g08831(.din(n25945), .dout(n26094));
  jor  g08832(.dina(n26094), .dinb(n26093), .dout(n26095));
  jand g08833(.dina(n26095), .dinb(n26005), .dout(n26096));
  jnot g08834(.din(n25948), .dout(n26097));
  jor  g08835(.dina(n26097), .dinb(n26096), .dout(n26098));
  jand g08836(.dina(n26098), .dinb(n26004), .dout(n26099));
  jnot g08837(.din(n25951), .dout(n26100));
  jor  g08838(.dina(n26100), .dinb(n26099), .dout(n26101));
  jand g08839(.dina(n26101), .dinb(n26003), .dout(n26102));
  jnot g08840(.din(n25954), .dout(n26103));
  jor  g08841(.dina(n26103), .dinb(n26102), .dout(n26104));
  jand g08842(.dina(n26104), .dinb(n26002), .dout(n26105));
  jnot g08843(.din(n25957), .dout(n26106));
  jor  g08844(.dina(n26106), .dinb(n26105), .dout(n26107));
  jand g08845(.dina(n26107), .dinb(n26001), .dout(n26108));
  jnot g08846(.din(n25960), .dout(n26109));
  jor  g08847(.dina(n26109), .dinb(n26108), .dout(n26110));
  jand g08848(.dina(n26110), .dinb(n26000), .dout(n26111));
  jnot g08849(.din(n25963), .dout(n26112));
  jor  g08850(.dina(n26112), .dinb(n26111), .dout(n26113));
  jand g08851(.dina(n26113), .dinb(n25999), .dout(n26114));
  jnot g08852(.din(n25966), .dout(n26115));
  jor  g08853(.dina(n26115), .dinb(n26114), .dout(n26116));
  jand g08854(.dina(n26116), .dinb(n25998), .dout(n26117));
  jnot g08855(.din(n25969), .dout(n26118));
  jor  g08856(.dina(n26118), .dinb(n26117), .dout(n26119));
  jand g08857(.dina(n26119), .dinb(n25997), .dout(n26120));
  jnot g08858(.din(n25972), .dout(n26121));
  jor  g08859(.dina(n26121), .dinb(n26120), .dout(n26122));
  jand g08860(.dina(n26122), .dinb(n25996), .dout(n26123));
  jnot g08861(.din(n25975), .dout(n26124));
  jor  g08862(.dina(n26124), .dinb(n26123), .dout(n26125));
  jand g08863(.dina(n26125), .dinb(n25995), .dout(n26126));
  jnot g08864(.din(n25978), .dout(n26127));
  jor  g08865(.dina(n26127), .dinb(n26126), .dout(n26128));
  jand g08866(.dina(n26128), .dinb(n25994), .dout(n26129));
  jnot g08867(.din(n25981), .dout(n26130));
  jor  g08868(.dina(n26130), .dinb(n26129), .dout(n26131));
  jand g08869(.dina(n26131), .dinb(n25993), .dout(n26132));
  jnot g08870(.din(n25984), .dout(n26133));
  jor  g08871(.dina(n26133), .dinb(n26132), .dout(n26134));
  jand g08872(.dina(n26134), .dinb(n25992), .dout(n26135));
  jor  g08873(.dina(n26135), .dinb(n25552), .dout(n26136));
  jand g08874(.dina(n26136), .dinb(n25991), .dout(n26137));
  jor  g08875(.dina(n26137), .dinb(n6437), .dout(n26138));
  jxor g08876(.dina(n25984), .dinb(n25983), .dout(n26139));
  jor  g08877(.dina(n26139), .dinb(n26138), .dout(n26140));
  jand g08878(.dina(n26140), .dinb(n25990), .dout(n26141));
  jand g08879(.dina(n26141), .dinb(n325), .dout(n26142));
  jor  g08880(.dina(n25989), .dinb(n25558), .dout(n26143));
  jxor g08881(.dina(n25981), .dinb(n25980), .dout(n26144));
  jor  g08882(.dina(n26144), .dinb(n26138), .dout(n26145));
  jand g08883(.dina(n26145), .dinb(n26143), .dout(n26146));
  jand g08884(.dina(n26146), .dinb(n324), .dout(n26147));
  jor  g08885(.dina(n25989), .dinb(n25563), .dout(n26148));
  jxor g08886(.dina(n25978), .dinb(n25977), .dout(n26149));
  jor  g08887(.dina(n26149), .dinb(n26138), .dout(n26150));
  jand g08888(.dina(n26150), .dinb(n26148), .dout(n26151));
  jand g08889(.dina(n26151), .dinb(n276), .dout(n26152));
  jor  g08890(.dina(n25989), .dinb(n25568), .dout(n26153));
  jxor g08891(.dina(n25975), .dinb(n25974), .dout(n26154));
  jor  g08892(.dina(n26154), .dinb(n26138), .dout(n26155));
  jand g08893(.dina(n26155), .dinb(n26153), .dout(n26156));
  jand g08894(.dina(n26156), .dinb(n333), .dout(n26157));
  jor  g08895(.dina(n25989), .dinb(n25573), .dout(n26158));
  jxor g08896(.dina(n25972), .dinb(n25971), .dout(n26159));
  jor  g08897(.dina(n26159), .dinb(n26138), .dout(n26160));
  jand g08898(.dina(n26160), .dinb(n26158), .dout(n26161));
  jand g08899(.dina(n26161), .dinb(n332), .dout(n26162));
  jor  g08900(.dina(n25989), .dinb(n25578), .dout(n26163));
  jxor g08901(.dina(n25969), .dinb(n25968), .dout(n26164));
  jor  g08902(.dina(n26164), .dinb(n26138), .dout(n26165));
  jand g08903(.dina(n26165), .dinb(n26163), .dout(n26166));
  jand g08904(.dina(n26166), .dinb(n331), .dout(n26167));
  jor  g08905(.dina(n25989), .dinb(n25583), .dout(n26168));
  jxor g08906(.dina(n25966), .dinb(n25965), .dout(n26169));
  jor  g08907(.dina(n26169), .dinb(n26138), .dout(n26170));
  jand g08908(.dina(n26170), .dinb(n26168), .dout(n26171));
  jand g08909(.dina(n26171), .dinb(n275), .dout(n26172));
  jor  g08910(.dina(n25989), .dinb(n25588), .dout(n26173));
  jxor g08911(.dina(n25963), .dinb(n25962), .dout(n26174));
  jor  g08912(.dina(n26174), .dinb(n26138), .dout(n26175));
  jand g08913(.dina(n26175), .dinb(n26173), .dout(n26176));
  jand g08914(.dina(n26176), .dinb(n340), .dout(n26177));
  jor  g08915(.dina(n25989), .dinb(n25593), .dout(n26178));
  jxor g08916(.dina(n25960), .dinb(n25959), .dout(n26179));
  jor  g08917(.dina(n26179), .dinb(n26138), .dout(n26180));
  jand g08918(.dina(n26180), .dinb(n26178), .dout(n26181));
  jand g08919(.dina(n26181), .dinb(n339), .dout(n26182));
  jor  g08920(.dina(n25989), .dinb(n25598), .dout(n26183));
  jxor g08921(.dina(n25957), .dinb(n25956), .dout(n26184));
  jor  g08922(.dina(n26184), .dinb(n26138), .dout(n26185));
  jand g08923(.dina(n26185), .dinb(n26183), .dout(n26186));
  jand g08924(.dina(n26186), .dinb(n338), .dout(n26187));
  jor  g08925(.dina(n25989), .dinb(n25603), .dout(n26188));
  jxor g08926(.dina(n25954), .dinb(n25953), .dout(n26189));
  jor  g08927(.dina(n26189), .dinb(n26138), .dout(n26190));
  jand g08928(.dina(n26190), .dinb(n26188), .dout(n26191));
  jand g08929(.dina(n26191), .dinb(n271), .dout(n26192));
  jor  g08930(.dina(n25989), .dinb(n25608), .dout(n26193));
  jxor g08931(.dina(n25951), .dinb(n25950), .dout(n26194));
  jor  g08932(.dina(n26194), .dinb(n26138), .dout(n26195));
  jand g08933(.dina(n26195), .dinb(n26193), .dout(n26196));
  jand g08934(.dina(n26196), .dinb(n270), .dout(n26197));
  jor  g08935(.dina(n25989), .dinb(n25613), .dout(n26198));
  jxor g08936(.dina(n25948), .dinb(n25947), .dout(n26199));
  jor  g08937(.dina(n26199), .dinb(n26138), .dout(n26200));
  jand g08938(.dina(n26200), .dinb(n26198), .dout(n26201));
  jand g08939(.dina(n26201), .dinb(n269), .dout(n26202));
  jor  g08940(.dina(n25989), .dinb(n25618), .dout(n26203));
  jxor g08941(.dina(n25945), .dinb(n25944), .dout(n26204));
  jor  g08942(.dina(n26204), .dinb(n26138), .dout(n26205));
  jand g08943(.dina(n26205), .dinb(n26203), .dout(n26206));
  jand g08944(.dina(n26206), .dinb(n274), .dout(n26207));
  jor  g08945(.dina(n25989), .dinb(n25623), .dout(n26208));
  jxor g08946(.dina(n25942), .dinb(n25941), .dout(n26209));
  jor  g08947(.dina(n26209), .dinb(n26138), .dout(n26210));
  jand g08948(.dina(n26210), .dinb(n26208), .dout(n26211));
  jand g08949(.dina(n26211), .dinb(n268), .dout(n26212));
  jor  g08950(.dina(n25989), .dinb(n25628), .dout(n26213));
  jxor g08951(.dina(n25939), .dinb(n25938), .dout(n26214));
  jor  g08952(.dina(n26214), .dinb(n26138), .dout(n26215));
  jand g08953(.dina(n26215), .dinb(n26213), .dout(n26216));
  jand g08954(.dina(n26216), .dinb(n349), .dout(n26217));
  jor  g08955(.dina(n25989), .dinb(n25633), .dout(n26218));
  jxor g08956(.dina(n25936), .dinb(n25935), .dout(n26219));
  jor  g08957(.dina(n26219), .dinb(n26138), .dout(n26220));
  jand g08958(.dina(n26220), .dinb(n26218), .dout(n26221));
  jand g08959(.dina(n26221), .dinb(n348), .dout(n26222));
  jor  g08960(.dina(n25989), .dinb(n25638), .dout(n26223));
  jxor g08961(.dina(n25933), .dinb(n25932), .dout(n26224));
  jor  g08962(.dina(n26224), .dinb(n26138), .dout(n26225));
  jand g08963(.dina(n26225), .dinb(n26223), .dout(n26226));
  jand g08964(.dina(n26226), .dinb(n347), .dout(n26227));
  jor  g08965(.dina(n25989), .dinb(n25643), .dout(n26228));
  jxor g08966(.dina(n25930), .dinb(n25929), .dout(n26229));
  jor  g08967(.dina(n26229), .dinb(n26138), .dout(n26230));
  jand g08968(.dina(n26230), .dinb(n26228), .dout(n26231));
  jand g08969(.dina(n26231), .dinb(n267), .dout(n26232));
  jor  g08970(.dina(n25989), .dinb(n25648), .dout(n26233));
  jxor g08971(.dina(n25927), .dinb(n25926), .dout(n26234));
  jor  g08972(.dina(n26234), .dinb(n26138), .dout(n26235));
  jand g08973(.dina(n26235), .dinb(n26233), .dout(n26236));
  jand g08974(.dina(n26236), .dinb(n266), .dout(n26237));
  jor  g08975(.dina(n25989), .dinb(n25653), .dout(n26238));
  jxor g08976(.dina(n25924), .dinb(n25923), .dout(n26239));
  jor  g08977(.dina(n26239), .dinb(n26138), .dout(n26240));
  jand g08978(.dina(n26240), .dinb(n26238), .dout(n26241));
  jand g08979(.dina(n26241), .dinb(n356), .dout(n26242));
  jor  g08980(.dina(n25989), .dinb(n25658), .dout(n26243));
  jxor g08981(.dina(n25921), .dinb(n25920), .dout(n26244));
  jor  g08982(.dina(n26244), .dinb(n26138), .dout(n26245));
  jand g08983(.dina(n26245), .dinb(n26243), .dout(n26246));
  jand g08984(.dina(n26246), .dinb(n355), .dout(n26247));
  jor  g08985(.dina(n25989), .dinb(n25663), .dout(n26248));
  jxor g08986(.dina(n25918), .dinb(n25917), .dout(n26249));
  jor  g08987(.dina(n26249), .dinb(n26138), .dout(n26250));
  jand g08988(.dina(n26250), .dinb(n26248), .dout(n26251));
  jand g08989(.dina(n26251), .dinb(n364), .dout(n26252));
  jor  g08990(.dina(n25989), .dinb(n25668), .dout(n26253));
  jxor g08991(.dina(n25915), .dinb(n25914), .dout(n26254));
  jor  g08992(.dina(n26254), .dinb(n26138), .dout(n26255));
  jand g08993(.dina(n26255), .dinb(n26253), .dout(n26256));
  jand g08994(.dina(n26256), .dinb(n361), .dout(n26257));
  jor  g08995(.dina(n25989), .dinb(n25673), .dout(n26258));
  jxor g08996(.dina(n25912), .dinb(n25911), .dout(n26259));
  jor  g08997(.dina(n26259), .dinb(n26138), .dout(n26260));
  jand g08998(.dina(n26260), .dinb(n26258), .dout(n26261));
  jand g08999(.dina(n26261), .dinb(n360), .dout(n26262));
  jor  g09000(.dina(n25989), .dinb(n25678), .dout(n26263));
  jxor g09001(.dina(n25909), .dinb(n25908), .dout(n26264));
  jor  g09002(.dina(n26264), .dinb(n26138), .dout(n26265));
  jand g09003(.dina(n26265), .dinb(n26263), .dout(n26266));
  jand g09004(.dina(n26266), .dinb(n363), .dout(n26267));
  jor  g09005(.dina(n25989), .dinb(n25683), .dout(n26268));
  jxor g09006(.dina(n25906), .dinb(n25905), .dout(n26269));
  jor  g09007(.dina(n26269), .dinb(n26138), .dout(n26270));
  jand g09008(.dina(n26270), .dinb(n26268), .dout(n26271));
  jand g09009(.dina(n26271), .dinb(n359), .dout(n26272));
  jor  g09010(.dina(n25989), .dinb(n25688), .dout(n26273));
  jxor g09011(.dina(n25903), .dinb(n25902), .dout(n26274));
  jor  g09012(.dina(n26274), .dinb(n26138), .dout(n26275));
  jand g09013(.dina(n26275), .dinb(n26273), .dout(n26276));
  jand g09014(.dina(n26276), .dinb(n369), .dout(n26277));
  jor  g09015(.dina(n25989), .dinb(n25693), .dout(n26278));
  jxor g09016(.dina(n25900), .dinb(n25899), .dout(n26279));
  jor  g09017(.dina(n26279), .dinb(n26138), .dout(n26280));
  jand g09018(.dina(n26280), .dinb(n26278), .dout(n26281));
  jand g09019(.dina(n26281), .dinb(n368), .dout(n26282));
  jor  g09020(.dina(n25989), .dinb(n25698), .dout(n26283));
  jxor g09021(.dina(n25897), .dinb(n25896), .dout(n26284));
  jor  g09022(.dina(n26284), .dinb(n26138), .dout(n26285));
  jand g09023(.dina(n26285), .dinb(n26283), .dout(n26286));
  jand g09024(.dina(n26286), .dinb(n367), .dout(n26287));
  jor  g09025(.dina(n25989), .dinb(n25703), .dout(n26288));
  jxor g09026(.dina(n25894), .dinb(n25893), .dout(n26289));
  jor  g09027(.dina(n26289), .dinb(n26138), .dout(n26290));
  jand g09028(.dina(n26290), .dinb(n26288), .dout(n26291));
  jand g09029(.dina(n26291), .dinb(n265), .dout(n26292));
  jor  g09030(.dina(n25989), .dinb(n25708), .dout(n26293));
  jxor g09031(.dina(n25891), .dinb(n25890), .dout(n26294));
  jor  g09032(.dina(n26294), .dinb(n26138), .dout(n26295));
  jand g09033(.dina(n26295), .dinb(n26293), .dout(n26296));
  jand g09034(.dina(n26296), .dinb(n378), .dout(n26297));
  jor  g09035(.dina(n25989), .dinb(n25713), .dout(n26298));
  jxor g09036(.dina(n25888), .dinb(n25887), .dout(n26299));
  jor  g09037(.dina(n26299), .dinb(n26138), .dout(n26300));
  jand g09038(.dina(n26300), .dinb(n26298), .dout(n26301));
  jand g09039(.dina(n26301), .dinb(n377), .dout(n26302));
  jor  g09040(.dina(n25989), .dinb(n25718), .dout(n26303));
  jxor g09041(.dina(n25885), .dinb(n25884), .dout(n26304));
  jor  g09042(.dina(n26304), .dinb(n26138), .dout(n26305));
  jand g09043(.dina(n26305), .dinb(n26303), .dout(n26306));
  jand g09044(.dina(n26306), .dinb(n376), .dout(n26307));
  jor  g09045(.dina(n25989), .dinb(n25723), .dout(n26308));
  jxor g09046(.dina(n25882), .dinb(n25881), .dout(n26309));
  jor  g09047(.dina(n26309), .dinb(n26138), .dout(n26310));
  jand g09048(.dina(n26310), .dinb(n26308), .dout(n26311));
  jand g09049(.dina(n26311), .dinb(n264), .dout(n26312));
  jand g09050(.dina(n26138), .dinb(n25874), .dout(n26313));
  jxor g09051(.dina(n25879), .dinb(n6812), .dout(n26314));
  jand g09052(.dina(n26314), .dinb(n25989), .dout(n26315));
  jor  g09053(.dina(n26315), .dinb(n26313), .dout(n26316));
  jand g09054(.dina(n26316), .dinb(n386), .dout(n26317));
  jnot g09055(.din(n7077), .dout(n26318));
  jor  g09056(.dina(n26137), .dinb(n26318), .dout(n26319));
  jand g09057(.dina(n26319), .dinb(a26 ), .dout(n26320));
  jand g09058(.dina(n25989), .dinb(n6662), .dout(n26321));
  jor  g09059(.dina(n26321), .dinb(n26320), .dout(n26322));
  jand g09060(.dina(n26322), .dinb(n259), .dout(n26323));
  jand g09061(.dina(n25988), .dinb(n7077), .dout(n26324));
  jor  g09062(.dina(n26324), .dinb(n6661), .dout(n26325));
  jor  g09063(.dina(n26138), .dinb(n6812), .dout(n26326));
  jand g09064(.dina(n26326), .dinb(n26325), .dout(n26327));
  jxor g09065(.dina(n26327), .dinb(b1 ), .dout(n26328));
  jand g09066(.dina(n26328), .dinb(n7086), .dout(n26329));
  jor  g09067(.dina(n26329), .dinb(n26323), .dout(n26330));
  jxor g09068(.dina(n26316), .dinb(n386), .dout(n26331));
  jand g09069(.dina(n26331), .dinb(n26330), .dout(n26332));
  jor  g09070(.dina(n26332), .dinb(n26317), .dout(n26333));
  jxor g09071(.dina(n26311), .dinb(n264), .dout(n26334));
  jand g09072(.dina(n26334), .dinb(n26333), .dout(n26335));
  jor  g09073(.dina(n26335), .dinb(n26312), .dout(n26336));
  jxor g09074(.dina(n26306), .dinb(n376), .dout(n26337));
  jand g09075(.dina(n26337), .dinb(n26336), .dout(n26338));
  jor  g09076(.dina(n26338), .dinb(n26307), .dout(n26339));
  jxor g09077(.dina(n26301), .dinb(n377), .dout(n26340));
  jand g09078(.dina(n26340), .dinb(n26339), .dout(n26341));
  jor  g09079(.dina(n26341), .dinb(n26302), .dout(n26342));
  jxor g09080(.dina(n26296), .dinb(n378), .dout(n26343));
  jand g09081(.dina(n26343), .dinb(n26342), .dout(n26344));
  jor  g09082(.dina(n26344), .dinb(n26297), .dout(n26345));
  jxor g09083(.dina(n26291), .dinb(n265), .dout(n26346));
  jand g09084(.dina(n26346), .dinb(n26345), .dout(n26347));
  jor  g09085(.dina(n26347), .dinb(n26292), .dout(n26348));
  jxor g09086(.dina(n26286), .dinb(n367), .dout(n26349));
  jand g09087(.dina(n26349), .dinb(n26348), .dout(n26350));
  jor  g09088(.dina(n26350), .dinb(n26287), .dout(n26351));
  jxor g09089(.dina(n26281), .dinb(n368), .dout(n26352));
  jand g09090(.dina(n26352), .dinb(n26351), .dout(n26353));
  jor  g09091(.dina(n26353), .dinb(n26282), .dout(n26354));
  jxor g09092(.dina(n26276), .dinb(n369), .dout(n26355));
  jand g09093(.dina(n26355), .dinb(n26354), .dout(n26356));
  jor  g09094(.dina(n26356), .dinb(n26277), .dout(n26357));
  jxor g09095(.dina(n26271), .dinb(n359), .dout(n26358));
  jand g09096(.dina(n26358), .dinb(n26357), .dout(n26359));
  jor  g09097(.dina(n26359), .dinb(n26272), .dout(n26360));
  jxor g09098(.dina(n26266), .dinb(n363), .dout(n26361));
  jand g09099(.dina(n26361), .dinb(n26360), .dout(n26362));
  jor  g09100(.dina(n26362), .dinb(n26267), .dout(n26363));
  jxor g09101(.dina(n26261), .dinb(n360), .dout(n26364));
  jand g09102(.dina(n26364), .dinb(n26363), .dout(n26365));
  jor  g09103(.dina(n26365), .dinb(n26262), .dout(n26366));
  jxor g09104(.dina(n26256), .dinb(n361), .dout(n26367));
  jand g09105(.dina(n26367), .dinb(n26366), .dout(n26368));
  jor  g09106(.dina(n26368), .dinb(n26257), .dout(n26369));
  jxor g09107(.dina(n26251), .dinb(n364), .dout(n26370));
  jand g09108(.dina(n26370), .dinb(n26369), .dout(n26371));
  jor  g09109(.dina(n26371), .dinb(n26252), .dout(n26372));
  jxor g09110(.dina(n26246), .dinb(n355), .dout(n26373));
  jand g09111(.dina(n26373), .dinb(n26372), .dout(n26374));
  jor  g09112(.dina(n26374), .dinb(n26247), .dout(n26375));
  jxor g09113(.dina(n26241), .dinb(n356), .dout(n26376));
  jand g09114(.dina(n26376), .dinb(n26375), .dout(n26377));
  jor  g09115(.dina(n26377), .dinb(n26242), .dout(n26378));
  jxor g09116(.dina(n26236), .dinb(n266), .dout(n26379));
  jand g09117(.dina(n26379), .dinb(n26378), .dout(n26380));
  jor  g09118(.dina(n26380), .dinb(n26237), .dout(n26381));
  jxor g09119(.dina(n26231), .dinb(n267), .dout(n26382));
  jand g09120(.dina(n26382), .dinb(n26381), .dout(n26383));
  jor  g09121(.dina(n26383), .dinb(n26232), .dout(n26384));
  jxor g09122(.dina(n26226), .dinb(n347), .dout(n26385));
  jand g09123(.dina(n26385), .dinb(n26384), .dout(n26386));
  jor  g09124(.dina(n26386), .dinb(n26227), .dout(n26387));
  jxor g09125(.dina(n26221), .dinb(n348), .dout(n26388));
  jand g09126(.dina(n26388), .dinb(n26387), .dout(n26389));
  jor  g09127(.dina(n26389), .dinb(n26222), .dout(n26390));
  jxor g09128(.dina(n26216), .dinb(n349), .dout(n26391));
  jand g09129(.dina(n26391), .dinb(n26390), .dout(n26392));
  jor  g09130(.dina(n26392), .dinb(n26217), .dout(n26393));
  jxor g09131(.dina(n26211), .dinb(n268), .dout(n26394));
  jand g09132(.dina(n26394), .dinb(n26393), .dout(n26395));
  jor  g09133(.dina(n26395), .dinb(n26212), .dout(n26396));
  jxor g09134(.dina(n26206), .dinb(n274), .dout(n26397));
  jand g09135(.dina(n26397), .dinb(n26396), .dout(n26398));
  jor  g09136(.dina(n26398), .dinb(n26207), .dout(n26399));
  jxor g09137(.dina(n26201), .dinb(n269), .dout(n26400));
  jand g09138(.dina(n26400), .dinb(n26399), .dout(n26401));
  jor  g09139(.dina(n26401), .dinb(n26202), .dout(n26402));
  jxor g09140(.dina(n26196), .dinb(n270), .dout(n26403));
  jand g09141(.dina(n26403), .dinb(n26402), .dout(n26404));
  jor  g09142(.dina(n26404), .dinb(n26197), .dout(n26405));
  jxor g09143(.dina(n26191), .dinb(n271), .dout(n26406));
  jand g09144(.dina(n26406), .dinb(n26405), .dout(n26407));
  jor  g09145(.dina(n26407), .dinb(n26192), .dout(n26408));
  jxor g09146(.dina(n26186), .dinb(n338), .dout(n26409));
  jand g09147(.dina(n26409), .dinb(n26408), .dout(n26410));
  jor  g09148(.dina(n26410), .dinb(n26187), .dout(n26411));
  jxor g09149(.dina(n26181), .dinb(n339), .dout(n26412));
  jand g09150(.dina(n26412), .dinb(n26411), .dout(n26413));
  jor  g09151(.dina(n26413), .dinb(n26182), .dout(n26414));
  jxor g09152(.dina(n26176), .dinb(n340), .dout(n26415));
  jand g09153(.dina(n26415), .dinb(n26414), .dout(n26416));
  jor  g09154(.dina(n26416), .dinb(n26177), .dout(n26417));
  jxor g09155(.dina(n26171), .dinb(n275), .dout(n26418));
  jand g09156(.dina(n26418), .dinb(n26417), .dout(n26419));
  jor  g09157(.dina(n26419), .dinb(n26172), .dout(n26420));
  jxor g09158(.dina(n26166), .dinb(n331), .dout(n26421));
  jand g09159(.dina(n26421), .dinb(n26420), .dout(n26422));
  jor  g09160(.dina(n26422), .dinb(n26167), .dout(n26423));
  jxor g09161(.dina(n26161), .dinb(n332), .dout(n26424));
  jand g09162(.dina(n26424), .dinb(n26423), .dout(n26425));
  jor  g09163(.dina(n26425), .dinb(n26162), .dout(n26426));
  jxor g09164(.dina(n26156), .dinb(n333), .dout(n26427));
  jand g09165(.dina(n26427), .dinb(n26426), .dout(n26428));
  jor  g09166(.dina(n26428), .dinb(n26157), .dout(n26429));
  jxor g09167(.dina(n26151), .dinb(n276), .dout(n26430));
  jand g09168(.dina(n26430), .dinb(n26429), .dout(n26431));
  jor  g09169(.dina(n26431), .dinb(n26152), .dout(n26432));
  jxor g09170(.dina(n26146), .dinb(n324), .dout(n26433));
  jand g09171(.dina(n26433), .dinb(n26432), .dout(n26434));
  jor  g09172(.dina(n26434), .dinb(n26147), .dout(n26435));
  jxor g09173(.dina(n26141), .dinb(n325), .dout(n26436));
  jand g09174(.dina(n26436), .dinb(n26435), .dout(n26437));
  jor  g09175(.dina(n26437), .dinb(n26142), .dout(n26438));
  jand g09176(.dina(n25986), .dinb(n408), .dout(n26439));
  jor  g09177(.dina(n26439), .dinb(n26138), .dout(n26440));
  jand g09178(.dina(n26440), .dinb(n25549), .dout(n26441));
  jxor g09179(.dina(n26441), .dinb(b38 ), .dout(n26442));
  jnot g09180(.din(n26442), .dout(n26443));
  jand g09181(.dina(n26443), .dinb(n26438), .dout(n26444));
  jand g09182(.dina(n26444), .dinb(n407), .dout(n26445));
  jand g09183(.dina(n26441), .dinb(n6436), .dout(n26446));
  jor  g09184(.dina(n26446), .dinb(n26445), .dout(n26447));
  jor  g09185(.dina(n26447), .dinb(n26141), .dout(n26448));
  jnot g09186(.din(n26447), .dout(n26449));
  jxor g09187(.dina(n26436), .dinb(n26435), .dout(n26450));
  jor  g09188(.dina(n26450), .dinb(n26449), .dout(n26451));
  jand g09189(.dina(n26451), .dinb(n26448), .dout(n26452));
  jand g09190(.dina(n26449), .dinb(n26441), .dout(n26453));
  jxor g09191(.dina(n26443), .dinb(n26438), .dout(n26454));
  jand g09192(.dina(n26454), .dinb(n26447), .dout(n26455));
  jor  g09193(.dina(n26455), .dinb(n26453), .dout(n26456));
  jand g09194(.dina(n26456), .dinb(n277), .dout(n26457));
  jnot g09195(.din(n26456), .dout(n26458));
  jand g09196(.dina(n26458), .dinb(b39 ), .dout(n26459));
  jnot g09197(.din(n26459), .dout(n26460));
  jand g09198(.dina(n26452), .dinb(n326), .dout(n26461));
  jor  g09199(.dina(n26447), .dinb(n26146), .dout(n26462));
  jxor g09200(.dina(n26433), .dinb(n26432), .dout(n26463));
  jor  g09201(.dina(n26463), .dinb(n26449), .dout(n26464));
  jand g09202(.dina(n26464), .dinb(n26462), .dout(n26465));
  jand g09203(.dina(n26465), .dinb(n325), .dout(n26466));
  jor  g09204(.dina(n26447), .dinb(n26151), .dout(n26467));
  jxor g09205(.dina(n26430), .dinb(n26429), .dout(n26468));
  jor  g09206(.dina(n26468), .dinb(n26449), .dout(n26469));
  jand g09207(.dina(n26469), .dinb(n26467), .dout(n26470));
  jand g09208(.dina(n26470), .dinb(n324), .dout(n26471));
  jor  g09209(.dina(n26447), .dinb(n26156), .dout(n26472));
  jxor g09210(.dina(n26427), .dinb(n26426), .dout(n26473));
  jor  g09211(.dina(n26473), .dinb(n26449), .dout(n26474));
  jand g09212(.dina(n26474), .dinb(n26472), .dout(n26475));
  jand g09213(.dina(n26475), .dinb(n276), .dout(n26476));
  jor  g09214(.dina(n26447), .dinb(n26161), .dout(n26477));
  jxor g09215(.dina(n26424), .dinb(n26423), .dout(n26478));
  jor  g09216(.dina(n26478), .dinb(n26449), .dout(n26479));
  jand g09217(.dina(n26479), .dinb(n26477), .dout(n26480));
  jand g09218(.dina(n26480), .dinb(n333), .dout(n26481));
  jor  g09219(.dina(n26447), .dinb(n26166), .dout(n26482));
  jxor g09220(.dina(n26421), .dinb(n26420), .dout(n26483));
  jor  g09221(.dina(n26483), .dinb(n26449), .dout(n26484));
  jand g09222(.dina(n26484), .dinb(n26482), .dout(n26485));
  jand g09223(.dina(n26485), .dinb(n332), .dout(n26486));
  jor  g09224(.dina(n26447), .dinb(n26171), .dout(n26487));
  jxor g09225(.dina(n26418), .dinb(n26417), .dout(n26488));
  jor  g09226(.dina(n26488), .dinb(n26449), .dout(n26489));
  jand g09227(.dina(n26489), .dinb(n26487), .dout(n26490));
  jand g09228(.dina(n26490), .dinb(n331), .dout(n26491));
  jor  g09229(.dina(n26447), .dinb(n26176), .dout(n26492));
  jxor g09230(.dina(n26415), .dinb(n26414), .dout(n26493));
  jor  g09231(.dina(n26493), .dinb(n26449), .dout(n26494));
  jand g09232(.dina(n26494), .dinb(n26492), .dout(n26495));
  jand g09233(.dina(n26495), .dinb(n275), .dout(n26496));
  jor  g09234(.dina(n26447), .dinb(n26181), .dout(n26497));
  jxor g09235(.dina(n26412), .dinb(n26411), .dout(n26498));
  jor  g09236(.dina(n26498), .dinb(n26449), .dout(n26499));
  jand g09237(.dina(n26499), .dinb(n26497), .dout(n26500));
  jand g09238(.dina(n26500), .dinb(n340), .dout(n26501));
  jor  g09239(.dina(n26447), .dinb(n26186), .dout(n26502));
  jxor g09240(.dina(n26409), .dinb(n26408), .dout(n26503));
  jor  g09241(.dina(n26503), .dinb(n26449), .dout(n26504));
  jand g09242(.dina(n26504), .dinb(n26502), .dout(n26505));
  jand g09243(.dina(n26505), .dinb(n339), .dout(n26506));
  jor  g09244(.dina(n26447), .dinb(n26191), .dout(n26507));
  jxor g09245(.dina(n26406), .dinb(n26405), .dout(n26508));
  jor  g09246(.dina(n26508), .dinb(n26449), .dout(n26509));
  jand g09247(.dina(n26509), .dinb(n26507), .dout(n26510));
  jand g09248(.dina(n26510), .dinb(n338), .dout(n26511));
  jor  g09249(.dina(n26447), .dinb(n26196), .dout(n26512));
  jxor g09250(.dina(n26403), .dinb(n26402), .dout(n26513));
  jor  g09251(.dina(n26513), .dinb(n26449), .dout(n26514));
  jand g09252(.dina(n26514), .dinb(n26512), .dout(n26515));
  jand g09253(.dina(n26515), .dinb(n271), .dout(n26516));
  jor  g09254(.dina(n26447), .dinb(n26201), .dout(n26517));
  jxor g09255(.dina(n26400), .dinb(n26399), .dout(n26518));
  jor  g09256(.dina(n26518), .dinb(n26449), .dout(n26519));
  jand g09257(.dina(n26519), .dinb(n26517), .dout(n26520));
  jand g09258(.dina(n26520), .dinb(n270), .dout(n26521));
  jor  g09259(.dina(n26447), .dinb(n26206), .dout(n26522));
  jxor g09260(.dina(n26397), .dinb(n26396), .dout(n26523));
  jor  g09261(.dina(n26523), .dinb(n26449), .dout(n26524));
  jand g09262(.dina(n26524), .dinb(n26522), .dout(n26525));
  jand g09263(.dina(n26525), .dinb(n269), .dout(n26526));
  jor  g09264(.dina(n26447), .dinb(n26211), .dout(n26527));
  jxor g09265(.dina(n26394), .dinb(n26393), .dout(n26528));
  jor  g09266(.dina(n26528), .dinb(n26449), .dout(n26529));
  jand g09267(.dina(n26529), .dinb(n26527), .dout(n26530));
  jand g09268(.dina(n26530), .dinb(n274), .dout(n26531));
  jor  g09269(.dina(n26447), .dinb(n26216), .dout(n26532));
  jxor g09270(.dina(n26391), .dinb(n26390), .dout(n26533));
  jor  g09271(.dina(n26533), .dinb(n26449), .dout(n26534));
  jand g09272(.dina(n26534), .dinb(n26532), .dout(n26535));
  jand g09273(.dina(n26535), .dinb(n268), .dout(n26536));
  jor  g09274(.dina(n26447), .dinb(n26221), .dout(n26537));
  jxor g09275(.dina(n26388), .dinb(n26387), .dout(n26538));
  jor  g09276(.dina(n26538), .dinb(n26449), .dout(n26539));
  jand g09277(.dina(n26539), .dinb(n26537), .dout(n26540));
  jand g09278(.dina(n26540), .dinb(n349), .dout(n26541));
  jor  g09279(.dina(n26447), .dinb(n26226), .dout(n26542));
  jxor g09280(.dina(n26385), .dinb(n26384), .dout(n26543));
  jor  g09281(.dina(n26543), .dinb(n26449), .dout(n26544));
  jand g09282(.dina(n26544), .dinb(n26542), .dout(n26545));
  jand g09283(.dina(n26545), .dinb(n348), .dout(n26546));
  jor  g09284(.dina(n26447), .dinb(n26231), .dout(n26547));
  jxor g09285(.dina(n26382), .dinb(n26381), .dout(n26548));
  jor  g09286(.dina(n26548), .dinb(n26449), .dout(n26549));
  jand g09287(.dina(n26549), .dinb(n26547), .dout(n26550));
  jand g09288(.dina(n26550), .dinb(n347), .dout(n26551));
  jor  g09289(.dina(n26447), .dinb(n26236), .dout(n26552));
  jxor g09290(.dina(n26379), .dinb(n26378), .dout(n26553));
  jor  g09291(.dina(n26553), .dinb(n26449), .dout(n26554));
  jand g09292(.dina(n26554), .dinb(n26552), .dout(n26555));
  jand g09293(.dina(n26555), .dinb(n267), .dout(n26556));
  jor  g09294(.dina(n26447), .dinb(n26241), .dout(n26557));
  jxor g09295(.dina(n26376), .dinb(n26375), .dout(n26558));
  jor  g09296(.dina(n26558), .dinb(n26449), .dout(n26559));
  jand g09297(.dina(n26559), .dinb(n26557), .dout(n26560));
  jand g09298(.dina(n26560), .dinb(n266), .dout(n26561));
  jor  g09299(.dina(n26447), .dinb(n26246), .dout(n26562));
  jxor g09300(.dina(n26373), .dinb(n26372), .dout(n26563));
  jor  g09301(.dina(n26563), .dinb(n26449), .dout(n26564));
  jand g09302(.dina(n26564), .dinb(n26562), .dout(n26565));
  jand g09303(.dina(n26565), .dinb(n356), .dout(n26566));
  jor  g09304(.dina(n26447), .dinb(n26251), .dout(n26567));
  jxor g09305(.dina(n26370), .dinb(n26369), .dout(n26568));
  jor  g09306(.dina(n26568), .dinb(n26449), .dout(n26569));
  jand g09307(.dina(n26569), .dinb(n26567), .dout(n26570));
  jand g09308(.dina(n26570), .dinb(n355), .dout(n26571));
  jor  g09309(.dina(n26447), .dinb(n26256), .dout(n26572));
  jxor g09310(.dina(n26367), .dinb(n26366), .dout(n26573));
  jor  g09311(.dina(n26573), .dinb(n26449), .dout(n26574));
  jand g09312(.dina(n26574), .dinb(n26572), .dout(n26575));
  jand g09313(.dina(n26575), .dinb(n364), .dout(n26576));
  jor  g09314(.dina(n26447), .dinb(n26261), .dout(n26577));
  jxor g09315(.dina(n26364), .dinb(n26363), .dout(n26578));
  jor  g09316(.dina(n26578), .dinb(n26449), .dout(n26579));
  jand g09317(.dina(n26579), .dinb(n26577), .dout(n26580));
  jand g09318(.dina(n26580), .dinb(n361), .dout(n26581));
  jor  g09319(.dina(n26447), .dinb(n26266), .dout(n26582));
  jxor g09320(.dina(n26361), .dinb(n26360), .dout(n26583));
  jor  g09321(.dina(n26583), .dinb(n26449), .dout(n26584));
  jand g09322(.dina(n26584), .dinb(n26582), .dout(n26585));
  jand g09323(.dina(n26585), .dinb(n360), .dout(n26586));
  jor  g09324(.dina(n26447), .dinb(n26271), .dout(n26587));
  jxor g09325(.dina(n26358), .dinb(n26357), .dout(n26588));
  jor  g09326(.dina(n26588), .dinb(n26449), .dout(n26589));
  jand g09327(.dina(n26589), .dinb(n26587), .dout(n26590));
  jand g09328(.dina(n26590), .dinb(n363), .dout(n26591));
  jor  g09329(.dina(n26447), .dinb(n26276), .dout(n26592));
  jxor g09330(.dina(n26355), .dinb(n26354), .dout(n26593));
  jor  g09331(.dina(n26593), .dinb(n26449), .dout(n26594));
  jand g09332(.dina(n26594), .dinb(n26592), .dout(n26595));
  jand g09333(.dina(n26595), .dinb(n359), .dout(n26596));
  jor  g09334(.dina(n26447), .dinb(n26281), .dout(n26597));
  jxor g09335(.dina(n26352), .dinb(n26351), .dout(n26598));
  jor  g09336(.dina(n26598), .dinb(n26449), .dout(n26599));
  jand g09337(.dina(n26599), .dinb(n26597), .dout(n26600));
  jand g09338(.dina(n26600), .dinb(n369), .dout(n26601));
  jor  g09339(.dina(n26447), .dinb(n26286), .dout(n26602));
  jxor g09340(.dina(n26349), .dinb(n26348), .dout(n26603));
  jor  g09341(.dina(n26603), .dinb(n26449), .dout(n26604));
  jand g09342(.dina(n26604), .dinb(n26602), .dout(n26605));
  jand g09343(.dina(n26605), .dinb(n368), .dout(n26606));
  jor  g09344(.dina(n26447), .dinb(n26291), .dout(n26607));
  jxor g09345(.dina(n26346), .dinb(n26345), .dout(n26608));
  jor  g09346(.dina(n26608), .dinb(n26449), .dout(n26609));
  jand g09347(.dina(n26609), .dinb(n26607), .dout(n26610));
  jand g09348(.dina(n26610), .dinb(n367), .dout(n26611));
  jor  g09349(.dina(n26447), .dinb(n26296), .dout(n26612));
  jxor g09350(.dina(n26343), .dinb(n26342), .dout(n26613));
  jor  g09351(.dina(n26613), .dinb(n26449), .dout(n26614));
  jand g09352(.dina(n26614), .dinb(n26612), .dout(n26615));
  jand g09353(.dina(n26615), .dinb(n265), .dout(n26616));
  jor  g09354(.dina(n26447), .dinb(n26301), .dout(n26617));
  jxor g09355(.dina(n26340), .dinb(n26339), .dout(n26618));
  jor  g09356(.dina(n26618), .dinb(n26449), .dout(n26619));
  jand g09357(.dina(n26619), .dinb(n26617), .dout(n26620));
  jand g09358(.dina(n26620), .dinb(n378), .dout(n26621));
  jor  g09359(.dina(n26447), .dinb(n26306), .dout(n26622));
  jxor g09360(.dina(n26337), .dinb(n26336), .dout(n26623));
  jor  g09361(.dina(n26623), .dinb(n26449), .dout(n26624));
  jand g09362(.dina(n26624), .dinb(n26622), .dout(n26625));
  jand g09363(.dina(n26625), .dinb(n377), .dout(n26626));
  jor  g09364(.dina(n26447), .dinb(n26311), .dout(n26627));
  jxor g09365(.dina(n26334), .dinb(n26333), .dout(n26628));
  jor  g09366(.dina(n26628), .dinb(n26449), .dout(n26629));
  jand g09367(.dina(n26629), .dinb(n26627), .dout(n26630));
  jand g09368(.dina(n26630), .dinb(n376), .dout(n26631));
  jor  g09369(.dina(n26447), .dinb(n26316), .dout(n26632));
  jxor g09370(.dina(n26331), .dinb(n26330), .dout(n26633));
  jor  g09371(.dina(n26633), .dinb(n26449), .dout(n26634));
  jand g09372(.dina(n26634), .dinb(n26632), .dout(n26635));
  jand g09373(.dina(n26635), .dinb(n264), .dout(n26636));
  jor  g09374(.dina(n26447), .dinb(n26327), .dout(n26637));
  jxor g09375(.dina(n26328), .dinb(n7086), .dout(n26638));
  jand g09376(.dina(n26638), .dinb(n26447), .dout(n26639));
  jnot g09377(.din(n26639), .dout(n26640));
  jand g09378(.dina(n26640), .dinb(n26637), .dout(n26641));
  jnot g09379(.din(n26641), .dout(n26642));
  jand g09380(.dina(n26642), .dinb(n386), .dout(n26643));
  jand g09381(.dina(n26447), .dinb(b0 ), .dout(n26644));
  jxor g09382(.dina(n26644), .dinb(a25 ), .dout(n26645));
  jand g09383(.dina(n26645), .dinb(n259), .dout(n26646));
  jxor g09384(.dina(n26644), .dinb(n7084), .dout(n26647));
  jxor g09385(.dina(n26647), .dinb(b1 ), .dout(n26648));
  jand g09386(.dina(n26648), .dinb(n7403), .dout(n26649));
  jor  g09387(.dina(n26649), .dinb(n26646), .dout(n26650));
  jxor g09388(.dina(n26641), .dinb(b2 ), .dout(n26651));
  jand g09389(.dina(n26651), .dinb(n26650), .dout(n26652));
  jor  g09390(.dina(n26652), .dinb(n26643), .dout(n26653));
  jxor g09391(.dina(n26635), .dinb(n264), .dout(n26654));
  jand g09392(.dina(n26654), .dinb(n26653), .dout(n26655));
  jor  g09393(.dina(n26655), .dinb(n26636), .dout(n26656));
  jxor g09394(.dina(n26630), .dinb(n376), .dout(n26657));
  jand g09395(.dina(n26657), .dinb(n26656), .dout(n26658));
  jor  g09396(.dina(n26658), .dinb(n26631), .dout(n26659));
  jxor g09397(.dina(n26625), .dinb(n377), .dout(n26660));
  jand g09398(.dina(n26660), .dinb(n26659), .dout(n26661));
  jor  g09399(.dina(n26661), .dinb(n26626), .dout(n26662));
  jxor g09400(.dina(n26620), .dinb(n378), .dout(n26663));
  jand g09401(.dina(n26663), .dinb(n26662), .dout(n26664));
  jor  g09402(.dina(n26664), .dinb(n26621), .dout(n26665));
  jxor g09403(.dina(n26615), .dinb(n265), .dout(n26666));
  jand g09404(.dina(n26666), .dinb(n26665), .dout(n26667));
  jor  g09405(.dina(n26667), .dinb(n26616), .dout(n26668));
  jxor g09406(.dina(n26610), .dinb(n367), .dout(n26669));
  jand g09407(.dina(n26669), .dinb(n26668), .dout(n26670));
  jor  g09408(.dina(n26670), .dinb(n26611), .dout(n26671));
  jxor g09409(.dina(n26605), .dinb(n368), .dout(n26672));
  jand g09410(.dina(n26672), .dinb(n26671), .dout(n26673));
  jor  g09411(.dina(n26673), .dinb(n26606), .dout(n26674));
  jxor g09412(.dina(n26600), .dinb(n369), .dout(n26675));
  jand g09413(.dina(n26675), .dinb(n26674), .dout(n26676));
  jor  g09414(.dina(n26676), .dinb(n26601), .dout(n26677));
  jxor g09415(.dina(n26595), .dinb(n359), .dout(n26678));
  jand g09416(.dina(n26678), .dinb(n26677), .dout(n26679));
  jor  g09417(.dina(n26679), .dinb(n26596), .dout(n26680));
  jxor g09418(.dina(n26590), .dinb(n363), .dout(n26681));
  jand g09419(.dina(n26681), .dinb(n26680), .dout(n26682));
  jor  g09420(.dina(n26682), .dinb(n26591), .dout(n26683));
  jxor g09421(.dina(n26585), .dinb(n360), .dout(n26684));
  jand g09422(.dina(n26684), .dinb(n26683), .dout(n26685));
  jor  g09423(.dina(n26685), .dinb(n26586), .dout(n26686));
  jxor g09424(.dina(n26580), .dinb(n361), .dout(n26687));
  jand g09425(.dina(n26687), .dinb(n26686), .dout(n26688));
  jor  g09426(.dina(n26688), .dinb(n26581), .dout(n26689));
  jxor g09427(.dina(n26575), .dinb(n364), .dout(n26690));
  jand g09428(.dina(n26690), .dinb(n26689), .dout(n26691));
  jor  g09429(.dina(n26691), .dinb(n26576), .dout(n26692));
  jxor g09430(.dina(n26570), .dinb(n355), .dout(n26693));
  jand g09431(.dina(n26693), .dinb(n26692), .dout(n26694));
  jor  g09432(.dina(n26694), .dinb(n26571), .dout(n26695));
  jxor g09433(.dina(n26565), .dinb(n356), .dout(n26696));
  jand g09434(.dina(n26696), .dinb(n26695), .dout(n26697));
  jor  g09435(.dina(n26697), .dinb(n26566), .dout(n26698));
  jxor g09436(.dina(n26560), .dinb(n266), .dout(n26699));
  jand g09437(.dina(n26699), .dinb(n26698), .dout(n26700));
  jor  g09438(.dina(n26700), .dinb(n26561), .dout(n26701));
  jxor g09439(.dina(n26555), .dinb(n267), .dout(n26702));
  jand g09440(.dina(n26702), .dinb(n26701), .dout(n26703));
  jor  g09441(.dina(n26703), .dinb(n26556), .dout(n26704));
  jxor g09442(.dina(n26550), .dinb(n347), .dout(n26705));
  jand g09443(.dina(n26705), .dinb(n26704), .dout(n26706));
  jor  g09444(.dina(n26706), .dinb(n26551), .dout(n26707));
  jxor g09445(.dina(n26545), .dinb(n348), .dout(n26708));
  jand g09446(.dina(n26708), .dinb(n26707), .dout(n26709));
  jor  g09447(.dina(n26709), .dinb(n26546), .dout(n26710));
  jxor g09448(.dina(n26540), .dinb(n349), .dout(n26711));
  jand g09449(.dina(n26711), .dinb(n26710), .dout(n26712));
  jor  g09450(.dina(n26712), .dinb(n26541), .dout(n26713));
  jxor g09451(.dina(n26535), .dinb(n268), .dout(n26714));
  jand g09452(.dina(n26714), .dinb(n26713), .dout(n26715));
  jor  g09453(.dina(n26715), .dinb(n26536), .dout(n26716));
  jxor g09454(.dina(n26530), .dinb(n274), .dout(n26717));
  jand g09455(.dina(n26717), .dinb(n26716), .dout(n26718));
  jor  g09456(.dina(n26718), .dinb(n26531), .dout(n26719));
  jxor g09457(.dina(n26525), .dinb(n269), .dout(n26720));
  jand g09458(.dina(n26720), .dinb(n26719), .dout(n26721));
  jor  g09459(.dina(n26721), .dinb(n26526), .dout(n26722));
  jxor g09460(.dina(n26520), .dinb(n270), .dout(n26723));
  jand g09461(.dina(n26723), .dinb(n26722), .dout(n26724));
  jor  g09462(.dina(n26724), .dinb(n26521), .dout(n26725));
  jxor g09463(.dina(n26515), .dinb(n271), .dout(n26726));
  jand g09464(.dina(n26726), .dinb(n26725), .dout(n26727));
  jor  g09465(.dina(n26727), .dinb(n26516), .dout(n26728));
  jxor g09466(.dina(n26510), .dinb(n338), .dout(n26729));
  jand g09467(.dina(n26729), .dinb(n26728), .dout(n26730));
  jor  g09468(.dina(n26730), .dinb(n26511), .dout(n26731));
  jxor g09469(.dina(n26505), .dinb(n339), .dout(n26732));
  jand g09470(.dina(n26732), .dinb(n26731), .dout(n26733));
  jor  g09471(.dina(n26733), .dinb(n26506), .dout(n26734));
  jxor g09472(.dina(n26500), .dinb(n340), .dout(n26735));
  jand g09473(.dina(n26735), .dinb(n26734), .dout(n26736));
  jor  g09474(.dina(n26736), .dinb(n26501), .dout(n26737));
  jxor g09475(.dina(n26495), .dinb(n275), .dout(n26738));
  jand g09476(.dina(n26738), .dinb(n26737), .dout(n26739));
  jor  g09477(.dina(n26739), .dinb(n26496), .dout(n26740));
  jxor g09478(.dina(n26490), .dinb(n331), .dout(n26741));
  jand g09479(.dina(n26741), .dinb(n26740), .dout(n26742));
  jor  g09480(.dina(n26742), .dinb(n26491), .dout(n26743));
  jxor g09481(.dina(n26485), .dinb(n332), .dout(n26744));
  jand g09482(.dina(n26744), .dinb(n26743), .dout(n26745));
  jor  g09483(.dina(n26745), .dinb(n26486), .dout(n26746));
  jxor g09484(.dina(n26480), .dinb(n333), .dout(n26747));
  jand g09485(.dina(n26747), .dinb(n26746), .dout(n26748));
  jor  g09486(.dina(n26748), .dinb(n26481), .dout(n26749));
  jxor g09487(.dina(n26475), .dinb(n276), .dout(n26750));
  jand g09488(.dina(n26750), .dinb(n26749), .dout(n26751));
  jor  g09489(.dina(n26751), .dinb(n26476), .dout(n26752));
  jxor g09490(.dina(n26470), .dinb(n324), .dout(n26753));
  jand g09491(.dina(n26753), .dinb(n26752), .dout(n26754));
  jor  g09492(.dina(n26754), .dinb(n26471), .dout(n26755));
  jxor g09493(.dina(n26465), .dinb(n325), .dout(n26756));
  jand g09494(.dina(n26756), .dinb(n26755), .dout(n26757));
  jor  g09495(.dina(n26757), .dinb(n26466), .dout(n26758));
  jxor g09496(.dina(n26452), .dinb(n326), .dout(n26759));
  jand g09497(.dina(n26759), .dinb(n26758), .dout(n26760));
  jor  g09498(.dina(n26760), .dinb(n26461), .dout(n26761));
  jand g09499(.dina(n26761), .dinb(n26460), .dout(n26762));
  jor  g09500(.dina(n26762), .dinb(n26457), .dout(n26763));
  jand g09501(.dina(n26763), .dinb(n406), .dout(n26764));
  jor  g09502(.dina(n26764), .dinb(n26452), .dout(n26765));
  jnot g09503(.din(n26764), .dout(n26766));
  jxor g09504(.dina(n26759), .dinb(n26758), .dout(n26767));
  jor  g09505(.dina(n26767), .dinb(n26766), .dout(n26768));
  jand g09506(.dina(n26768), .dinb(n26765), .dout(n26769));
  jand g09507(.dina(n26766), .dinb(n26456), .dout(n26770));
  jand g09508(.dina(n26761), .dinb(n26457), .dout(n26771));
  jor  g09509(.dina(n26771), .dinb(n26770), .dout(n26772));
  jand g09510(.dina(n26772), .dinb(n278), .dout(n26773));
  jnot g09511(.din(n26772), .dout(n26774));
  jand g09512(.dina(n26774), .dinb(b40 ), .dout(n26775));
  jnot g09513(.din(n26775), .dout(n26776));
  jand g09514(.dina(n26769), .dinb(n277), .dout(n26777));
  jor  g09515(.dina(n26764), .dinb(n26465), .dout(n26778));
  jxor g09516(.dina(n26756), .dinb(n26755), .dout(n26779));
  jor  g09517(.dina(n26779), .dinb(n26766), .dout(n26780));
  jand g09518(.dina(n26780), .dinb(n26778), .dout(n26781));
  jand g09519(.dina(n26781), .dinb(n326), .dout(n26782));
  jor  g09520(.dina(n26764), .dinb(n26470), .dout(n26783));
  jxor g09521(.dina(n26753), .dinb(n26752), .dout(n26784));
  jor  g09522(.dina(n26784), .dinb(n26766), .dout(n26785));
  jand g09523(.dina(n26785), .dinb(n26783), .dout(n26786));
  jand g09524(.dina(n26786), .dinb(n325), .dout(n26787));
  jor  g09525(.dina(n26764), .dinb(n26475), .dout(n26788));
  jxor g09526(.dina(n26750), .dinb(n26749), .dout(n26789));
  jor  g09527(.dina(n26789), .dinb(n26766), .dout(n26790));
  jand g09528(.dina(n26790), .dinb(n26788), .dout(n26791));
  jand g09529(.dina(n26791), .dinb(n324), .dout(n26792));
  jor  g09530(.dina(n26764), .dinb(n26480), .dout(n26793));
  jxor g09531(.dina(n26747), .dinb(n26746), .dout(n26794));
  jor  g09532(.dina(n26794), .dinb(n26766), .dout(n26795));
  jand g09533(.dina(n26795), .dinb(n26793), .dout(n26796));
  jand g09534(.dina(n26796), .dinb(n276), .dout(n26797));
  jor  g09535(.dina(n26764), .dinb(n26485), .dout(n26798));
  jxor g09536(.dina(n26744), .dinb(n26743), .dout(n26799));
  jor  g09537(.dina(n26799), .dinb(n26766), .dout(n26800));
  jand g09538(.dina(n26800), .dinb(n26798), .dout(n26801));
  jand g09539(.dina(n26801), .dinb(n333), .dout(n26802));
  jor  g09540(.dina(n26764), .dinb(n26490), .dout(n26803));
  jxor g09541(.dina(n26741), .dinb(n26740), .dout(n26804));
  jor  g09542(.dina(n26804), .dinb(n26766), .dout(n26805));
  jand g09543(.dina(n26805), .dinb(n26803), .dout(n26806));
  jand g09544(.dina(n26806), .dinb(n332), .dout(n26807));
  jor  g09545(.dina(n26764), .dinb(n26495), .dout(n26808));
  jxor g09546(.dina(n26738), .dinb(n26737), .dout(n26809));
  jor  g09547(.dina(n26809), .dinb(n26766), .dout(n26810));
  jand g09548(.dina(n26810), .dinb(n26808), .dout(n26811));
  jand g09549(.dina(n26811), .dinb(n331), .dout(n26812));
  jor  g09550(.dina(n26764), .dinb(n26500), .dout(n26813));
  jxor g09551(.dina(n26735), .dinb(n26734), .dout(n26814));
  jor  g09552(.dina(n26814), .dinb(n26766), .dout(n26815));
  jand g09553(.dina(n26815), .dinb(n26813), .dout(n26816));
  jand g09554(.dina(n26816), .dinb(n275), .dout(n26817));
  jor  g09555(.dina(n26764), .dinb(n26505), .dout(n26818));
  jxor g09556(.dina(n26732), .dinb(n26731), .dout(n26819));
  jor  g09557(.dina(n26819), .dinb(n26766), .dout(n26820));
  jand g09558(.dina(n26820), .dinb(n26818), .dout(n26821));
  jand g09559(.dina(n26821), .dinb(n340), .dout(n26822));
  jor  g09560(.dina(n26764), .dinb(n26510), .dout(n26823));
  jxor g09561(.dina(n26729), .dinb(n26728), .dout(n26824));
  jor  g09562(.dina(n26824), .dinb(n26766), .dout(n26825));
  jand g09563(.dina(n26825), .dinb(n26823), .dout(n26826));
  jand g09564(.dina(n26826), .dinb(n339), .dout(n26827));
  jor  g09565(.dina(n26764), .dinb(n26515), .dout(n26828));
  jxor g09566(.dina(n26726), .dinb(n26725), .dout(n26829));
  jor  g09567(.dina(n26829), .dinb(n26766), .dout(n26830));
  jand g09568(.dina(n26830), .dinb(n26828), .dout(n26831));
  jand g09569(.dina(n26831), .dinb(n338), .dout(n26832));
  jor  g09570(.dina(n26764), .dinb(n26520), .dout(n26833));
  jxor g09571(.dina(n26723), .dinb(n26722), .dout(n26834));
  jor  g09572(.dina(n26834), .dinb(n26766), .dout(n26835));
  jand g09573(.dina(n26835), .dinb(n26833), .dout(n26836));
  jand g09574(.dina(n26836), .dinb(n271), .dout(n26837));
  jor  g09575(.dina(n26764), .dinb(n26525), .dout(n26838));
  jxor g09576(.dina(n26720), .dinb(n26719), .dout(n26839));
  jor  g09577(.dina(n26839), .dinb(n26766), .dout(n26840));
  jand g09578(.dina(n26840), .dinb(n26838), .dout(n26841));
  jand g09579(.dina(n26841), .dinb(n270), .dout(n26842));
  jor  g09580(.dina(n26764), .dinb(n26530), .dout(n26843));
  jxor g09581(.dina(n26717), .dinb(n26716), .dout(n26844));
  jor  g09582(.dina(n26844), .dinb(n26766), .dout(n26845));
  jand g09583(.dina(n26845), .dinb(n26843), .dout(n26846));
  jand g09584(.dina(n26846), .dinb(n269), .dout(n26847));
  jor  g09585(.dina(n26764), .dinb(n26535), .dout(n26848));
  jxor g09586(.dina(n26714), .dinb(n26713), .dout(n26849));
  jor  g09587(.dina(n26849), .dinb(n26766), .dout(n26850));
  jand g09588(.dina(n26850), .dinb(n26848), .dout(n26851));
  jand g09589(.dina(n26851), .dinb(n274), .dout(n26852));
  jor  g09590(.dina(n26764), .dinb(n26540), .dout(n26853));
  jxor g09591(.dina(n26711), .dinb(n26710), .dout(n26854));
  jor  g09592(.dina(n26854), .dinb(n26766), .dout(n26855));
  jand g09593(.dina(n26855), .dinb(n26853), .dout(n26856));
  jand g09594(.dina(n26856), .dinb(n268), .dout(n26857));
  jor  g09595(.dina(n26764), .dinb(n26545), .dout(n26858));
  jxor g09596(.dina(n26708), .dinb(n26707), .dout(n26859));
  jor  g09597(.dina(n26859), .dinb(n26766), .dout(n26860));
  jand g09598(.dina(n26860), .dinb(n26858), .dout(n26861));
  jand g09599(.dina(n26861), .dinb(n349), .dout(n26862));
  jor  g09600(.dina(n26764), .dinb(n26550), .dout(n26863));
  jxor g09601(.dina(n26705), .dinb(n26704), .dout(n26864));
  jor  g09602(.dina(n26864), .dinb(n26766), .dout(n26865));
  jand g09603(.dina(n26865), .dinb(n26863), .dout(n26866));
  jand g09604(.dina(n26866), .dinb(n348), .dout(n26867));
  jor  g09605(.dina(n26764), .dinb(n26555), .dout(n26868));
  jxor g09606(.dina(n26702), .dinb(n26701), .dout(n26869));
  jor  g09607(.dina(n26869), .dinb(n26766), .dout(n26870));
  jand g09608(.dina(n26870), .dinb(n26868), .dout(n26871));
  jand g09609(.dina(n26871), .dinb(n347), .dout(n26872));
  jor  g09610(.dina(n26764), .dinb(n26560), .dout(n26873));
  jxor g09611(.dina(n26699), .dinb(n26698), .dout(n26874));
  jor  g09612(.dina(n26874), .dinb(n26766), .dout(n26875));
  jand g09613(.dina(n26875), .dinb(n26873), .dout(n26876));
  jand g09614(.dina(n26876), .dinb(n267), .dout(n26877));
  jor  g09615(.dina(n26764), .dinb(n26565), .dout(n26878));
  jxor g09616(.dina(n26696), .dinb(n26695), .dout(n26879));
  jor  g09617(.dina(n26879), .dinb(n26766), .dout(n26880));
  jand g09618(.dina(n26880), .dinb(n26878), .dout(n26881));
  jand g09619(.dina(n26881), .dinb(n266), .dout(n26882));
  jor  g09620(.dina(n26764), .dinb(n26570), .dout(n26883));
  jxor g09621(.dina(n26693), .dinb(n26692), .dout(n26884));
  jor  g09622(.dina(n26884), .dinb(n26766), .dout(n26885));
  jand g09623(.dina(n26885), .dinb(n26883), .dout(n26886));
  jand g09624(.dina(n26886), .dinb(n356), .dout(n26887));
  jor  g09625(.dina(n26764), .dinb(n26575), .dout(n26888));
  jxor g09626(.dina(n26690), .dinb(n26689), .dout(n26889));
  jor  g09627(.dina(n26889), .dinb(n26766), .dout(n26890));
  jand g09628(.dina(n26890), .dinb(n26888), .dout(n26891));
  jand g09629(.dina(n26891), .dinb(n355), .dout(n26892));
  jor  g09630(.dina(n26764), .dinb(n26580), .dout(n26893));
  jxor g09631(.dina(n26687), .dinb(n26686), .dout(n26894));
  jor  g09632(.dina(n26894), .dinb(n26766), .dout(n26895));
  jand g09633(.dina(n26895), .dinb(n26893), .dout(n26896));
  jand g09634(.dina(n26896), .dinb(n364), .dout(n26897));
  jor  g09635(.dina(n26764), .dinb(n26585), .dout(n26898));
  jxor g09636(.dina(n26684), .dinb(n26683), .dout(n26899));
  jor  g09637(.dina(n26899), .dinb(n26766), .dout(n26900));
  jand g09638(.dina(n26900), .dinb(n26898), .dout(n26901));
  jand g09639(.dina(n26901), .dinb(n361), .dout(n26902));
  jor  g09640(.dina(n26764), .dinb(n26590), .dout(n26903));
  jxor g09641(.dina(n26681), .dinb(n26680), .dout(n26904));
  jor  g09642(.dina(n26904), .dinb(n26766), .dout(n26905));
  jand g09643(.dina(n26905), .dinb(n26903), .dout(n26906));
  jand g09644(.dina(n26906), .dinb(n360), .dout(n26907));
  jor  g09645(.dina(n26764), .dinb(n26595), .dout(n26908));
  jxor g09646(.dina(n26678), .dinb(n26677), .dout(n26909));
  jor  g09647(.dina(n26909), .dinb(n26766), .dout(n26910));
  jand g09648(.dina(n26910), .dinb(n26908), .dout(n26911));
  jand g09649(.dina(n26911), .dinb(n363), .dout(n26912));
  jor  g09650(.dina(n26764), .dinb(n26600), .dout(n26913));
  jxor g09651(.dina(n26675), .dinb(n26674), .dout(n26914));
  jor  g09652(.dina(n26914), .dinb(n26766), .dout(n26915));
  jand g09653(.dina(n26915), .dinb(n26913), .dout(n26916));
  jand g09654(.dina(n26916), .dinb(n359), .dout(n26917));
  jor  g09655(.dina(n26764), .dinb(n26605), .dout(n26918));
  jxor g09656(.dina(n26672), .dinb(n26671), .dout(n26919));
  jor  g09657(.dina(n26919), .dinb(n26766), .dout(n26920));
  jand g09658(.dina(n26920), .dinb(n26918), .dout(n26921));
  jand g09659(.dina(n26921), .dinb(n369), .dout(n26922));
  jor  g09660(.dina(n26764), .dinb(n26610), .dout(n26923));
  jxor g09661(.dina(n26669), .dinb(n26668), .dout(n26924));
  jor  g09662(.dina(n26924), .dinb(n26766), .dout(n26925));
  jand g09663(.dina(n26925), .dinb(n26923), .dout(n26926));
  jand g09664(.dina(n26926), .dinb(n368), .dout(n26927));
  jor  g09665(.dina(n26764), .dinb(n26615), .dout(n26928));
  jxor g09666(.dina(n26666), .dinb(n26665), .dout(n26929));
  jor  g09667(.dina(n26929), .dinb(n26766), .dout(n26930));
  jand g09668(.dina(n26930), .dinb(n26928), .dout(n26931));
  jand g09669(.dina(n26931), .dinb(n367), .dout(n26932));
  jor  g09670(.dina(n26764), .dinb(n26620), .dout(n26933));
  jxor g09671(.dina(n26663), .dinb(n26662), .dout(n26934));
  jor  g09672(.dina(n26934), .dinb(n26766), .dout(n26935));
  jand g09673(.dina(n26935), .dinb(n26933), .dout(n26936));
  jand g09674(.dina(n26936), .dinb(n265), .dout(n26937));
  jor  g09675(.dina(n26764), .dinb(n26625), .dout(n26938));
  jxor g09676(.dina(n26660), .dinb(n26659), .dout(n26939));
  jor  g09677(.dina(n26939), .dinb(n26766), .dout(n26940));
  jand g09678(.dina(n26940), .dinb(n26938), .dout(n26941));
  jand g09679(.dina(n26941), .dinb(n378), .dout(n26942));
  jor  g09680(.dina(n26764), .dinb(n26630), .dout(n26943));
  jxor g09681(.dina(n26657), .dinb(n26656), .dout(n26944));
  jor  g09682(.dina(n26944), .dinb(n26766), .dout(n26945));
  jand g09683(.dina(n26945), .dinb(n26943), .dout(n26946));
  jand g09684(.dina(n26946), .dinb(n377), .dout(n26947));
  jor  g09685(.dina(n26764), .dinb(n26635), .dout(n26948));
  jxor g09686(.dina(n26654), .dinb(n26653), .dout(n26949));
  jor  g09687(.dina(n26949), .dinb(n26766), .dout(n26950));
  jand g09688(.dina(n26950), .dinb(n26948), .dout(n26951));
  jand g09689(.dina(n26951), .dinb(n376), .dout(n26952));
  jor  g09690(.dina(n26764), .dinb(n26642), .dout(n26953));
  jxor g09691(.dina(n26651), .dinb(n26650), .dout(n26954));
  jor  g09692(.dina(n26954), .dinb(n26766), .dout(n26955));
  jand g09693(.dina(n26955), .dinb(n26953), .dout(n26956));
  jand g09694(.dina(n26956), .dinb(n264), .dout(n26957));
  jor  g09695(.dina(n26764), .dinb(n26645), .dout(n26958));
  jxor g09696(.dina(n26648), .dinb(n7403), .dout(n26959));
  jor  g09697(.dina(n26959), .dinb(n26766), .dout(n26960));
  jand g09698(.dina(n26960), .dinb(n26958), .dout(n26961));
  jand g09699(.dina(n26961), .dinb(n386), .dout(n26962));
  jnot g09700(.din(n7075), .dout(n26963));
  jnot g09701(.din(n26457), .dout(n26964));
  jnot g09702(.din(n26461), .dout(n26965));
  jnot g09703(.din(n26466), .dout(n26966));
  jnot g09704(.din(n26471), .dout(n26967));
  jnot g09705(.din(n26476), .dout(n26968));
  jnot g09706(.din(n26481), .dout(n26969));
  jnot g09707(.din(n26486), .dout(n26970));
  jnot g09708(.din(n26491), .dout(n26971));
  jnot g09709(.din(n26496), .dout(n26972));
  jnot g09710(.din(n26501), .dout(n26973));
  jnot g09711(.din(n26506), .dout(n26974));
  jnot g09712(.din(n26511), .dout(n26975));
  jnot g09713(.din(n26516), .dout(n26976));
  jnot g09714(.din(n26521), .dout(n26977));
  jnot g09715(.din(n26526), .dout(n26978));
  jnot g09716(.din(n26531), .dout(n26979));
  jnot g09717(.din(n26536), .dout(n26980));
  jnot g09718(.din(n26541), .dout(n26981));
  jnot g09719(.din(n26546), .dout(n26982));
  jnot g09720(.din(n26551), .dout(n26983));
  jnot g09721(.din(n26556), .dout(n26984));
  jnot g09722(.din(n26561), .dout(n26985));
  jnot g09723(.din(n26566), .dout(n26986));
  jnot g09724(.din(n26571), .dout(n26987));
  jnot g09725(.din(n26576), .dout(n26988));
  jnot g09726(.din(n26581), .dout(n26989));
  jnot g09727(.din(n26586), .dout(n26990));
  jnot g09728(.din(n26591), .dout(n26991));
  jnot g09729(.din(n26596), .dout(n26992));
  jnot g09730(.din(n26601), .dout(n26993));
  jnot g09731(.din(n26606), .dout(n26994));
  jnot g09732(.din(n26611), .dout(n26995));
  jnot g09733(.din(n26616), .dout(n26996));
  jnot g09734(.din(n26621), .dout(n26997));
  jnot g09735(.din(n26626), .dout(n26998));
  jnot g09736(.din(n26631), .dout(n26999));
  jnot g09737(.din(n26636), .dout(n27000));
  jnot g09738(.din(n26643), .dout(n27001));
  jnot g09739(.din(n26646), .dout(n27002));
  jxor g09740(.dina(n26647), .dinb(n259), .dout(n27003));
  jor  g09741(.dina(n27003), .dinb(n7402), .dout(n27004));
  jand g09742(.dina(n27004), .dinb(n27002), .dout(n27005));
  jnot g09743(.din(n26651), .dout(n27006));
  jor  g09744(.dina(n27006), .dinb(n27005), .dout(n27007));
  jand g09745(.dina(n27007), .dinb(n27001), .dout(n27008));
  jnot g09746(.din(n26654), .dout(n27009));
  jor  g09747(.dina(n27009), .dinb(n27008), .dout(n27010));
  jand g09748(.dina(n27010), .dinb(n27000), .dout(n27011));
  jnot g09749(.din(n26657), .dout(n27012));
  jor  g09750(.dina(n27012), .dinb(n27011), .dout(n27013));
  jand g09751(.dina(n27013), .dinb(n26999), .dout(n27014));
  jnot g09752(.din(n26660), .dout(n27015));
  jor  g09753(.dina(n27015), .dinb(n27014), .dout(n27016));
  jand g09754(.dina(n27016), .dinb(n26998), .dout(n27017));
  jnot g09755(.din(n26663), .dout(n27018));
  jor  g09756(.dina(n27018), .dinb(n27017), .dout(n27019));
  jand g09757(.dina(n27019), .dinb(n26997), .dout(n27020));
  jnot g09758(.din(n26666), .dout(n27021));
  jor  g09759(.dina(n27021), .dinb(n27020), .dout(n27022));
  jand g09760(.dina(n27022), .dinb(n26996), .dout(n27023));
  jnot g09761(.din(n26669), .dout(n27024));
  jor  g09762(.dina(n27024), .dinb(n27023), .dout(n27025));
  jand g09763(.dina(n27025), .dinb(n26995), .dout(n27026));
  jnot g09764(.din(n26672), .dout(n27027));
  jor  g09765(.dina(n27027), .dinb(n27026), .dout(n27028));
  jand g09766(.dina(n27028), .dinb(n26994), .dout(n27029));
  jnot g09767(.din(n26675), .dout(n27030));
  jor  g09768(.dina(n27030), .dinb(n27029), .dout(n27031));
  jand g09769(.dina(n27031), .dinb(n26993), .dout(n27032));
  jnot g09770(.din(n26678), .dout(n27033));
  jor  g09771(.dina(n27033), .dinb(n27032), .dout(n27034));
  jand g09772(.dina(n27034), .dinb(n26992), .dout(n27035));
  jnot g09773(.din(n26681), .dout(n27036));
  jor  g09774(.dina(n27036), .dinb(n27035), .dout(n27037));
  jand g09775(.dina(n27037), .dinb(n26991), .dout(n27038));
  jnot g09776(.din(n26684), .dout(n27039));
  jor  g09777(.dina(n27039), .dinb(n27038), .dout(n27040));
  jand g09778(.dina(n27040), .dinb(n26990), .dout(n27041));
  jnot g09779(.din(n26687), .dout(n27042));
  jor  g09780(.dina(n27042), .dinb(n27041), .dout(n27043));
  jand g09781(.dina(n27043), .dinb(n26989), .dout(n27044));
  jnot g09782(.din(n26690), .dout(n27045));
  jor  g09783(.dina(n27045), .dinb(n27044), .dout(n27046));
  jand g09784(.dina(n27046), .dinb(n26988), .dout(n27047));
  jnot g09785(.din(n26693), .dout(n27048));
  jor  g09786(.dina(n27048), .dinb(n27047), .dout(n27049));
  jand g09787(.dina(n27049), .dinb(n26987), .dout(n27050));
  jnot g09788(.din(n26696), .dout(n27051));
  jor  g09789(.dina(n27051), .dinb(n27050), .dout(n27052));
  jand g09790(.dina(n27052), .dinb(n26986), .dout(n27053));
  jnot g09791(.din(n26699), .dout(n27054));
  jor  g09792(.dina(n27054), .dinb(n27053), .dout(n27055));
  jand g09793(.dina(n27055), .dinb(n26985), .dout(n27056));
  jnot g09794(.din(n26702), .dout(n27057));
  jor  g09795(.dina(n27057), .dinb(n27056), .dout(n27058));
  jand g09796(.dina(n27058), .dinb(n26984), .dout(n27059));
  jnot g09797(.din(n26705), .dout(n27060));
  jor  g09798(.dina(n27060), .dinb(n27059), .dout(n27061));
  jand g09799(.dina(n27061), .dinb(n26983), .dout(n27062));
  jnot g09800(.din(n26708), .dout(n27063));
  jor  g09801(.dina(n27063), .dinb(n27062), .dout(n27064));
  jand g09802(.dina(n27064), .dinb(n26982), .dout(n27065));
  jnot g09803(.din(n26711), .dout(n27066));
  jor  g09804(.dina(n27066), .dinb(n27065), .dout(n27067));
  jand g09805(.dina(n27067), .dinb(n26981), .dout(n27068));
  jnot g09806(.din(n26714), .dout(n27069));
  jor  g09807(.dina(n27069), .dinb(n27068), .dout(n27070));
  jand g09808(.dina(n27070), .dinb(n26980), .dout(n27071));
  jnot g09809(.din(n26717), .dout(n27072));
  jor  g09810(.dina(n27072), .dinb(n27071), .dout(n27073));
  jand g09811(.dina(n27073), .dinb(n26979), .dout(n27074));
  jnot g09812(.din(n26720), .dout(n27075));
  jor  g09813(.dina(n27075), .dinb(n27074), .dout(n27076));
  jand g09814(.dina(n27076), .dinb(n26978), .dout(n27077));
  jnot g09815(.din(n26723), .dout(n27078));
  jor  g09816(.dina(n27078), .dinb(n27077), .dout(n27079));
  jand g09817(.dina(n27079), .dinb(n26977), .dout(n27080));
  jnot g09818(.din(n26726), .dout(n27081));
  jor  g09819(.dina(n27081), .dinb(n27080), .dout(n27082));
  jand g09820(.dina(n27082), .dinb(n26976), .dout(n27083));
  jnot g09821(.din(n26729), .dout(n27084));
  jor  g09822(.dina(n27084), .dinb(n27083), .dout(n27085));
  jand g09823(.dina(n27085), .dinb(n26975), .dout(n27086));
  jnot g09824(.din(n26732), .dout(n27087));
  jor  g09825(.dina(n27087), .dinb(n27086), .dout(n27088));
  jand g09826(.dina(n27088), .dinb(n26974), .dout(n27089));
  jnot g09827(.din(n26735), .dout(n27090));
  jor  g09828(.dina(n27090), .dinb(n27089), .dout(n27091));
  jand g09829(.dina(n27091), .dinb(n26973), .dout(n27092));
  jnot g09830(.din(n26738), .dout(n27093));
  jor  g09831(.dina(n27093), .dinb(n27092), .dout(n27094));
  jand g09832(.dina(n27094), .dinb(n26972), .dout(n27095));
  jnot g09833(.din(n26741), .dout(n27096));
  jor  g09834(.dina(n27096), .dinb(n27095), .dout(n27097));
  jand g09835(.dina(n27097), .dinb(n26971), .dout(n27098));
  jnot g09836(.din(n26744), .dout(n27099));
  jor  g09837(.dina(n27099), .dinb(n27098), .dout(n27100));
  jand g09838(.dina(n27100), .dinb(n26970), .dout(n27101));
  jnot g09839(.din(n26747), .dout(n27102));
  jor  g09840(.dina(n27102), .dinb(n27101), .dout(n27103));
  jand g09841(.dina(n27103), .dinb(n26969), .dout(n27104));
  jnot g09842(.din(n26750), .dout(n27105));
  jor  g09843(.dina(n27105), .dinb(n27104), .dout(n27106));
  jand g09844(.dina(n27106), .dinb(n26968), .dout(n27107));
  jnot g09845(.din(n26753), .dout(n27108));
  jor  g09846(.dina(n27108), .dinb(n27107), .dout(n27109));
  jand g09847(.dina(n27109), .dinb(n26967), .dout(n27110));
  jnot g09848(.din(n26756), .dout(n27111));
  jor  g09849(.dina(n27111), .dinb(n27110), .dout(n27112));
  jand g09850(.dina(n27112), .dinb(n26966), .dout(n27113));
  jnot g09851(.din(n26759), .dout(n27114));
  jor  g09852(.dina(n27114), .dinb(n27113), .dout(n27115));
  jand g09853(.dina(n27115), .dinb(n26965), .dout(n27116));
  jor  g09854(.dina(n27116), .dinb(n26459), .dout(n27117));
  jand g09855(.dina(n27117), .dinb(n26964), .dout(n27118));
  jor  g09856(.dina(n27118), .dinb(n26963), .dout(n27119));
  jand g09857(.dina(n27119), .dinb(a24 ), .dout(n27120));
  jnot g09858(.din(n7723), .dout(n27121));
  jor  g09859(.dina(n27118), .dinb(n27121), .dout(n27122));
  jnot g09860(.din(n27122), .dout(n27123));
  jor  g09861(.dina(n27123), .dinb(n27120), .dout(n27124));
  jand g09862(.dina(n27124), .dinb(n259), .dout(n27125));
  jand g09863(.dina(n26763), .dinb(n7075), .dout(n27126));
  jor  g09864(.dina(n27126), .dinb(n7401), .dout(n27127));
  jand g09865(.dina(n27122), .dinb(n27127), .dout(n27128));
  jxor g09866(.dina(n27128), .dinb(b1 ), .dout(n27129));
  jand g09867(.dina(n27129), .dinb(n7731), .dout(n27130));
  jor  g09868(.dina(n27130), .dinb(n27125), .dout(n27131));
  jxor g09869(.dina(n26961), .dinb(n386), .dout(n27132));
  jand g09870(.dina(n27132), .dinb(n27131), .dout(n27133));
  jor  g09871(.dina(n27133), .dinb(n26962), .dout(n27134));
  jxor g09872(.dina(n26956), .dinb(n264), .dout(n27135));
  jand g09873(.dina(n27135), .dinb(n27134), .dout(n27136));
  jor  g09874(.dina(n27136), .dinb(n26957), .dout(n27137));
  jxor g09875(.dina(n26951), .dinb(n376), .dout(n27138));
  jand g09876(.dina(n27138), .dinb(n27137), .dout(n27139));
  jor  g09877(.dina(n27139), .dinb(n26952), .dout(n27140));
  jxor g09878(.dina(n26946), .dinb(n377), .dout(n27141));
  jand g09879(.dina(n27141), .dinb(n27140), .dout(n27142));
  jor  g09880(.dina(n27142), .dinb(n26947), .dout(n27143));
  jxor g09881(.dina(n26941), .dinb(n378), .dout(n27144));
  jand g09882(.dina(n27144), .dinb(n27143), .dout(n27145));
  jor  g09883(.dina(n27145), .dinb(n26942), .dout(n27146));
  jxor g09884(.dina(n26936), .dinb(n265), .dout(n27147));
  jand g09885(.dina(n27147), .dinb(n27146), .dout(n27148));
  jor  g09886(.dina(n27148), .dinb(n26937), .dout(n27149));
  jxor g09887(.dina(n26931), .dinb(n367), .dout(n27150));
  jand g09888(.dina(n27150), .dinb(n27149), .dout(n27151));
  jor  g09889(.dina(n27151), .dinb(n26932), .dout(n27152));
  jxor g09890(.dina(n26926), .dinb(n368), .dout(n27153));
  jand g09891(.dina(n27153), .dinb(n27152), .dout(n27154));
  jor  g09892(.dina(n27154), .dinb(n26927), .dout(n27155));
  jxor g09893(.dina(n26921), .dinb(n369), .dout(n27156));
  jand g09894(.dina(n27156), .dinb(n27155), .dout(n27157));
  jor  g09895(.dina(n27157), .dinb(n26922), .dout(n27158));
  jxor g09896(.dina(n26916), .dinb(n359), .dout(n27159));
  jand g09897(.dina(n27159), .dinb(n27158), .dout(n27160));
  jor  g09898(.dina(n27160), .dinb(n26917), .dout(n27161));
  jxor g09899(.dina(n26911), .dinb(n363), .dout(n27162));
  jand g09900(.dina(n27162), .dinb(n27161), .dout(n27163));
  jor  g09901(.dina(n27163), .dinb(n26912), .dout(n27164));
  jxor g09902(.dina(n26906), .dinb(n360), .dout(n27165));
  jand g09903(.dina(n27165), .dinb(n27164), .dout(n27166));
  jor  g09904(.dina(n27166), .dinb(n26907), .dout(n27167));
  jxor g09905(.dina(n26901), .dinb(n361), .dout(n27168));
  jand g09906(.dina(n27168), .dinb(n27167), .dout(n27169));
  jor  g09907(.dina(n27169), .dinb(n26902), .dout(n27170));
  jxor g09908(.dina(n26896), .dinb(n364), .dout(n27171));
  jand g09909(.dina(n27171), .dinb(n27170), .dout(n27172));
  jor  g09910(.dina(n27172), .dinb(n26897), .dout(n27173));
  jxor g09911(.dina(n26891), .dinb(n355), .dout(n27174));
  jand g09912(.dina(n27174), .dinb(n27173), .dout(n27175));
  jor  g09913(.dina(n27175), .dinb(n26892), .dout(n27176));
  jxor g09914(.dina(n26886), .dinb(n356), .dout(n27177));
  jand g09915(.dina(n27177), .dinb(n27176), .dout(n27178));
  jor  g09916(.dina(n27178), .dinb(n26887), .dout(n27179));
  jxor g09917(.dina(n26881), .dinb(n266), .dout(n27180));
  jand g09918(.dina(n27180), .dinb(n27179), .dout(n27181));
  jor  g09919(.dina(n27181), .dinb(n26882), .dout(n27182));
  jxor g09920(.dina(n26876), .dinb(n267), .dout(n27183));
  jand g09921(.dina(n27183), .dinb(n27182), .dout(n27184));
  jor  g09922(.dina(n27184), .dinb(n26877), .dout(n27185));
  jxor g09923(.dina(n26871), .dinb(n347), .dout(n27186));
  jand g09924(.dina(n27186), .dinb(n27185), .dout(n27187));
  jor  g09925(.dina(n27187), .dinb(n26872), .dout(n27188));
  jxor g09926(.dina(n26866), .dinb(n348), .dout(n27189));
  jand g09927(.dina(n27189), .dinb(n27188), .dout(n27190));
  jor  g09928(.dina(n27190), .dinb(n26867), .dout(n27191));
  jxor g09929(.dina(n26861), .dinb(n349), .dout(n27192));
  jand g09930(.dina(n27192), .dinb(n27191), .dout(n27193));
  jor  g09931(.dina(n27193), .dinb(n26862), .dout(n27194));
  jxor g09932(.dina(n26856), .dinb(n268), .dout(n27195));
  jand g09933(.dina(n27195), .dinb(n27194), .dout(n27196));
  jor  g09934(.dina(n27196), .dinb(n26857), .dout(n27197));
  jxor g09935(.dina(n26851), .dinb(n274), .dout(n27198));
  jand g09936(.dina(n27198), .dinb(n27197), .dout(n27199));
  jor  g09937(.dina(n27199), .dinb(n26852), .dout(n27200));
  jxor g09938(.dina(n26846), .dinb(n269), .dout(n27201));
  jand g09939(.dina(n27201), .dinb(n27200), .dout(n27202));
  jor  g09940(.dina(n27202), .dinb(n26847), .dout(n27203));
  jxor g09941(.dina(n26841), .dinb(n270), .dout(n27204));
  jand g09942(.dina(n27204), .dinb(n27203), .dout(n27205));
  jor  g09943(.dina(n27205), .dinb(n26842), .dout(n27206));
  jxor g09944(.dina(n26836), .dinb(n271), .dout(n27207));
  jand g09945(.dina(n27207), .dinb(n27206), .dout(n27208));
  jor  g09946(.dina(n27208), .dinb(n26837), .dout(n27209));
  jxor g09947(.dina(n26831), .dinb(n338), .dout(n27210));
  jand g09948(.dina(n27210), .dinb(n27209), .dout(n27211));
  jor  g09949(.dina(n27211), .dinb(n26832), .dout(n27212));
  jxor g09950(.dina(n26826), .dinb(n339), .dout(n27213));
  jand g09951(.dina(n27213), .dinb(n27212), .dout(n27214));
  jor  g09952(.dina(n27214), .dinb(n26827), .dout(n27215));
  jxor g09953(.dina(n26821), .dinb(n340), .dout(n27216));
  jand g09954(.dina(n27216), .dinb(n27215), .dout(n27217));
  jor  g09955(.dina(n27217), .dinb(n26822), .dout(n27218));
  jxor g09956(.dina(n26816), .dinb(n275), .dout(n27219));
  jand g09957(.dina(n27219), .dinb(n27218), .dout(n27220));
  jor  g09958(.dina(n27220), .dinb(n26817), .dout(n27221));
  jxor g09959(.dina(n26811), .dinb(n331), .dout(n27222));
  jand g09960(.dina(n27222), .dinb(n27221), .dout(n27223));
  jor  g09961(.dina(n27223), .dinb(n26812), .dout(n27224));
  jxor g09962(.dina(n26806), .dinb(n332), .dout(n27225));
  jand g09963(.dina(n27225), .dinb(n27224), .dout(n27226));
  jor  g09964(.dina(n27226), .dinb(n26807), .dout(n27227));
  jxor g09965(.dina(n26801), .dinb(n333), .dout(n27228));
  jand g09966(.dina(n27228), .dinb(n27227), .dout(n27229));
  jor  g09967(.dina(n27229), .dinb(n26802), .dout(n27230));
  jxor g09968(.dina(n26796), .dinb(n276), .dout(n27231));
  jand g09969(.dina(n27231), .dinb(n27230), .dout(n27232));
  jor  g09970(.dina(n27232), .dinb(n26797), .dout(n27233));
  jxor g09971(.dina(n26791), .dinb(n324), .dout(n27234));
  jand g09972(.dina(n27234), .dinb(n27233), .dout(n27235));
  jor  g09973(.dina(n27235), .dinb(n26792), .dout(n27236));
  jxor g09974(.dina(n26786), .dinb(n325), .dout(n27237));
  jand g09975(.dina(n27237), .dinb(n27236), .dout(n27238));
  jor  g09976(.dina(n27238), .dinb(n26787), .dout(n27239));
  jxor g09977(.dina(n26781), .dinb(n326), .dout(n27240));
  jand g09978(.dina(n27240), .dinb(n27239), .dout(n27241));
  jor  g09979(.dina(n27241), .dinb(n26782), .dout(n27242));
  jxor g09980(.dina(n26769), .dinb(n277), .dout(n27243));
  jand g09981(.dina(n27243), .dinb(n27242), .dout(n27244));
  jor  g09982(.dina(n27244), .dinb(n26777), .dout(n27245));
  jand g09983(.dina(n27245), .dinb(n26776), .dout(n27246));
  jor  g09984(.dina(n27246), .dinb(n26773), .dout(n27247));
  jand g09985(.dina(n27247), .dinb(n7527), .dout(n27248));
  jor  g09986(.dina(n27248), .dinb(n26769), .dout(n27249));
  jnot g09987(.din(n27248), .dout(n27250));
  jxor g09988(.dina(n27243), .dinb(n27242), .dout(n27251));
  jor  g09989(.dina(n27251), .dinb(n27250), .dout(n27252));
  jand g09990(.dina(n27252), .dinb(n27249), .dout(n27253));
  jand g09991(.dina(n27245), .dinb(n406), .dout(n27254));
  jor  g09992(.dina(n27254), .dinb(n27250), .dout(n27255));
  jand g09993(.dina(n27255), .dinb(n26772), .dout(n27256));
  jand g09994(.dina(n27256), .dinb(n7527), .dout(n27257));
  jand g09995(.dina(n27253), .dinb(n278), .dout(n27258));
  jor  g09996(.dina(n27248), .dinb(n26781), .dout(n27259));
  jxor g09997(.dina(n27240), .dinb(n27239), .dout(n27260));
  jor  g09998(.dina(n27260), .dinb(n27250), .dout(n27261));
  jand g09999(.dina(n27261), .dinb(n27259), .dout(n27262));
  jand g10000(.dina(n27262), .dinb(n277), .dout(n27263));
  jor  g10001(.dina(n27248), .dinb(n26786), .dout(n27264));
  jxor g10002(.dina(n27237), .dinb(n27236), .dout(n27265));
  jor  g10003(.dina(n27265), .dinb(n27250), .dout(n27266));
  jand g10004(.dina(n27266), .dinb(n27264), .dout(n27267));
  jand g10005(.dina(n27267), .dinb(n326), .dout(n27268));
  jor  g10006(.dina(n27248), .dinb(n26791), .dout(n27269));
  jxor g10007(.dina(n27234), .dinb(n27233), .dout(n27270));
  jor  g10008(.dina(n27270), .dinb(n27250), .dout(n27271));
  jand g10009(.dina(n27271), .dinb(n27269), .dout(n27272));
  jand g10010(.dina(n27272), .dinb(n325), .dout(n27273));
  jor  g10011(.dina(n27248), .dinb(n26796), .dout(n27274));
  jxor g10012(.dina(n27231), .dinb(n27230), .dout(n27275));
  jor  g10013(.dina(n27275), .dinb(n27250), .dout(n27276));
  jand g10014(.dina(n27276), .dinb(n27274), .dout(n27277));
  jand g10015(.dina(n27277), .dinb(n324), .dout(n27278));
  jor  g10016(.dina(n27248), .dinb(n26801), .dout(n27279));
  jxor g10017(.dina(n27228), .dinb(n27227), .dout(n27280));
  jor  g10018(.dina(n27280), .dinb(n27250), .dout(n27281));
  jand g10019(.dina(n27281), .dinb(n27279), .dout(n27282));
  jand g10020(.dina(n27282), .dinb(n276), .dout(n27283));
  jor  g10021(.dina(n27248), .dinb(n26806), .dout(n27284));
  jxor g10022(.dina(n27225), .dinb(n27224), .dout(n27285));
  jor  g10023(.dina(n27285), .dinb(n27250), .dout(n27286));
  jand g10024(.dina(n27286), .dinb(n27284), .dout(n27287));
  jand g10025(.dina(n27287), .dinb(n333), .dout(n27288));
  jor  g10026(.dina(n27248), .dinb(n26811), .dout(n27289));
  jxor g10027(.dina(n27222), .dinb(n27221), .dout(n27290));
  jor  g10028(.dina(n27290), .dinb(n27250), .dout(n27291));
  jand g10029(.dina(n27291), .dinb(n27289), .dout(n27292));
  jand g10030(.dina(n27292), .dinb(n332), .dout(n27293));
  jor  g10031(.dina(n27248), .dinb(n26816), .dout(n27294));
  jxor g10032(.dina(n27219), .dinb(n27218), .dout(n27295));
  jor  g10033(.dina(n27295), .dinb(n27250), .dout(n27296));
  jand g10034(.dina(n27296), .dinb(n27294), .dout(n27297));
  jand g10035(.dina(n27297), .dinb(n331), .dout(n27298));
  jor  g10036(.dina(n27248), .dinb(n26821), .dout(n27299));
  jxor g10037(.dina(n27216), .dinb(n27215), .dout(n27300));
  jor  g10038(.dina(n27300), .dinb(n27250), .dout(n27301));
  jand g10039(.dina(n27301), .dinb(n27299), .dout(n27302));
  jand g10040(.dina(n27302), .dinb(n275), .dout(n27303));
  jor  g10041(.dina(n27248), .dinb(n26826), .dout(n27304));
  jxor g10042(.dina(n27213), .dinb(n27212), .dout(n27305));
  jor  g10043(.dina(n27305), .dinb(n27250), .dout(n27306));
  jand g10044(.dina(n27306), .dinb(n27304), .dout(n27307));
  jand g10045(.dina(n27307), .dinb(n340), .dout(n27308));
  jor  g10046(.dina(n27248), .dinb(n26831), .dout(n27309));
  jxor g10047(.dina(n27210), .dinb(n27209), .dout(n27310));
  jor  g10048(.dina(n27310), .dinb(n27250), .dout(n27311));
  jand g10049(.dina(n27311), .dinb(n27309), .dout(n27312));
  jand g10050(.dina(n27312), .dinb(n339), .dout(n27313));
  jor  g10051(.dina(n27248), .dinb(n26836), .dout(n27314));
  jxor g10052(.dina(n27207), .dinb(n27206), .dout(n27315));
  jor  g10053(.dina(n27315), .dinb(n27250), .dout(n27316));
  jand g10054(.dina(n27316), .dinb(n27314), .dout(n27317));
  jand g10055(.dina(n27317), .dinb(n338), .dout(n27318));
  jor  g10056(.dina(n27248), .dinb(n26841), .dout(n27319));
  jxor g10057(.dina(n27204), .dinb(n27203), .dout(n27320));
  jor  g10058(.dina(n27320), .dinb(n27250), .dout(n27321));
  jand g10059(.dina(n27321), .dinb(n27319), .dout(n27322));
  jand g10060(.dina(n27322), .dinb(n271), .dout(n27323));
  jor  g10061(.dina(n27248), .dinb(n26846), .dout(n27324));
  jxor g10062(.dina(n27201), .dinb(n27200), .dout(n27325));
  jor  g10063(.dina(n27325), .dinb(n27250), .dout(n27326));
  jand g10064(.dina(n27326), .dinb(n27324), .dout(n27327));
  jand g10065(.dina(n27327), .dinb(n270), .dout(n27328));
  jor  g10066(.dina(n27248), .dinb(n26851), .dout(n27329));
  jxor g10067(.dina(n27198), .dinb(n27197), .dout(n27330));
  jor  g10068(.dina(n27330), .dinb(n27250), .dout(n27331));
  jand g10069(.dina(n27331), .dinb(n27329), .dout(n27332));
  jand g10070(.dina(n27332), .dinb(n269), .dout(n27333));
  jor  g10071(.dina(n27248), .dinb(n26856), .dout(n27334));
  jxor g10072(.dina(n27195), .dinb(n27194), .dout(n27335));
  jor  g10073(.dina(n27335), .dinb(n27250), .dout(n27336));
  jand g10074(.dina(n27336), .dinb(n27334), .dout(n27337));
  jand g10075(.dina(n27337), .dinb(n274), .dout(n27338));
  jor  g10076(.dina(n27248), .dinb(n26861), .dout(n27339));
  jxor g10077(.dina(n27192), .dinb(n27191), .dout(n27340));
  jor  g10078(.dina(n27340), .dinb(n27250), .dout(n27341));
  jand g10079(.dina(n27341), .dinb(n27339), .dout(n27342));
  jand g10080(.dina(n27342), .dinb(n268), .dout(n27343));
  jor  g10081(.dina(n27248), .dinb(n26866), .dout(n27344));
  jxor g10082(.dina(n27189), .dinb(n27188), .dout(n27345));
  jor  g10083(.dina(n27345), .dinb(n27250), .dout(n27346));
  jand g10084(.dina(n27346), .dinb(n27344), .dout(n27347));
  jand g10085(.dina(n27347), .dinb(n349), .dout(n27348));
  jor  g10086(.dina(n27248), .dinb(n26871), .dout(n27349));
  jxor g10087(.dina(n27186), .dinb(n27185), .dout(n27350));
  jor  g10088(.dina(n27350), .dinb(n27250), .dout(n27351));
  jand g10089(.dina(n27351), .dinb(n27349), .dout(n27352));
  jand g10090(.dina(n27352), .dinb(n348), .dout(n27353));
  jor  g10091(.dina(n27248), .dinb(n26876), .dout(n27354));
  jxor g10092(.dina(n27183), .dinb(n27182), .dout(n27355));
  jor  g10093(.dina(n27355), .dinb(n27250), .dout(n27356));
  jand g10094(.dina(n27356), .dinb(n27354), .dout(n27357));
  jand g10095(.dina(n27357), .dinb(n347), .dout(n27358));
  jor  g10096(.dina(n27248), .dinb(n26881), .dout(n27359));
  jxor g10097(.dina(n27180), .dinb(n27179), .dout(n27360));
  jor  g10098(.dina(n27360), .dinb(n27250), .dout(n27361));
  jand g10099(.dina(n27361), .dinb(n27359), .dout(n27362));
  jand g10100(.dina(n27362), .dinb(n267), .dout(n27363));
  jor  g10101(.dina(n27248), .dinb(n26886), .dout(n27364));
  jxor g10102(.dina(n27177), .dinb(n27176), .dout(n27365));
  jor  g10103(.dina(n27365), .dinb(n27250), .dout(n27366));
  jand g10104(.dina(n27366), .dinb(n27364), .dout(n27367));
  jand g10105(.dina(n27367), .dinb(n266), .dout(n27368));
  jor  g10106(.dina(n27248), .dinb(n26891), .dout(n27369));
  jxor g10107(.dina(n27174), .dinb(n27173), .dout(n27370));
  jor  g10108(.dina(n27370), .dinb(n27250), .dout(n27371));
  jand g10109(.dina(n27371), .dinb(n27369), .dout(n27372));
  jand g10110(.dina(n27372), .dinb(n356), .dout(n27373));
  jor  g10111(.dina(n27248), .dinb(n26896), .dout(n27374));
  jxor g10112(.dina(n27171), .dinb(n27170), .dout(n27375));
  jor  g10113(.dina(n27375), .dinb(n27250), .dout(n27376));
  jand g10114(.dina(n27376), .dinb(n27374), .dout(n27377));
  jand g10115(.dina(n27377), .dinb(n355), .dout(n27378));
  jor  g10116(.dina(n27248), .dinb(n26901), .dout(n27379));
  jxor g10117(.dina(n27168), .dinb(n27167), .dout(n27380));
  jor  g10118(.dina(n27380), .dinb(n27250), .dout(n27381));
  jand g10119(.dina(n27381), .dinb(n27379), .dout(n27382));
  jand g10120(.dina(n27382), .dinb(n364), .dout(n27383));
  jor  g10121(.dina(n27248), .dinb(n26906), .dout(n27384));
  jxor g10122(.dina(n27165), .dinb(n27164), .dout(n27385));
  jor  g10123(.dina(n27385), .dinb(n27250), .dout(n27386));
  jand g10124(.dina(n27386), .dinb(n27384), .dout(n27387));
  jand g10125(.dina(n27387), .dinb(n361), .dout(n27388));
  jor  g10126(.dina(n27248), .dinb(n26911), .dout(n27389));
  jxor g10127(.dina(n27162), .dinb(n27161), .dout(n27390));
  jor  g10128(.dina(n27390), .dinb(n27250), .dout(n27391));
  jand g10129(.dina(n27391), .dinb(n27389), .dout(n27392));
  jand g10130(.dina(n27392), .dinb(n360), .dout(n27393));
  jor  g10131(.dina(n27248), .dinb(n26916), .dout(n27394));
  jxor g10132(.dina(n27159), .dinb(n27158), .dout(n27395));
  jor  g10133(.dina(n27395), .dinb(n27250), .dout(n27396));
  jand g10134(.dina(n27396), .dinb(n27394), .dout(n27397));
  jand g10135(.dina(n27397), .dinb(n363), .dout(n27398));
  jor  g10136(.dina(n27248), .dinb(n26921), .dout(n27399));
  jxor g10137(.dina(n27156), .dinb(n27155), .dout(n27400));
  jor  g10138(.dina(n27400), .dinb(n27250), .dout(n27401));
  jand g10139(.dina(n27401), .dinb(n27399), .dout(n27402));
  jand g10140(.dina(n27402), .dinb(n359), .dout(n27403));
  jor  g10141(.dina(n27248), .dinb(n26926), .dout(n27404));
  jxor g10142(.dina(n27153), .dinb(n27152), .dout(n27405));
  jor  g10143(.dina(n27405), .dinb(n27250), .dout(n27406));
  jand g10144(.dina(n27406), .dinb(n27404), .dout(n27407));
  jand g10145(.dina(n27407), .dinb(n369), .dout(n27408));
  jor  g10146(.dina(n27248), .dinb(n26931), .dout(n27409));
  jxor g10147(.dina(n27150), .dinb(n27149), .dout(n27410));
  jor  g10148(.dina(n27410), .dinb(n27250), .dout(n27411));
  jand g10149(.dina(n27411), .dinb(n27409), .dout(n27412));
  jand g10150(.dina(n27412), .dinb(n368), .dout(n27413));
  jor  g10151(.dina(n27248), .dinb(n26936), .dout(n27414));
  jxor g10152(.dina(n27147), .dinb(n27146), .dout(n27415));
  jor  g10153(.dina(n27415), .dinb(n27250), .dout(n27416));
  jand g10154(.dina(n27416), .dinb(n27414), .dout(n27417));
  jand g10155(.dina(n27417), .dinb(n367), .dout(n27418));
  jor  g10156(.dina(n27248), .dinb(n26941), .dout(n27419));
  jxor g10157(.dina(n27144), .dinb(n27143), .dout(n27420));
  jor  g10158(.dina(n27420), .dinb(n27250), .dout(n27421));
  jand g10159(.dina(n27421), .dinb(n27419), .dout(n27422));
  jand g10160(.dina(n27422), .dinb(n265), .dout(n27423));
  jor  g10161(.dina(n27248), .dinb(n26946), .dout(n27424));
  jxor g10162(.dina(n27141), .dinb(n27140), .dout(n27425));
  jor  g10163(.dina(n27425), .dinb(n27250), .dout(n27426));
  jand g10164(.dina(n27426), .dinb(n27424), .dout(n27427));
  jand g10165(.dina(n27427), .dinb(n378), .dout(n27428));
  jor  g10166(.dina(n27248), .dinb(n26951), .dout(n27429));
  jxor g10167(.dina(n27138), .dinb(n27137), .dout(n27430));
  jor  g10168(.dina(n27430), .dinb(n27250), .dout(n27431));
  jand g10169(.dina(n27431), .dinb(n27429), .dout(n27432));
  jand g10170(.dina(n27432), .dinb(n377), .dout(n27433));
  jor  g10171(.dina(n27248), .dinb(n26956), .dout(n27434));
  jxor g10172(.dina(n27135), .dinb(n27134), .dout(n27435));
  jor  g10173(.dina(n27435), .dinb(n27250), .dout(n27436));
  jand g10174(.dina(n27436), .dinb(n27434), .dout(n27437));
  jand g10175(.dina(n27437), .dinb(n376), .dout(n27438));
  jor  g10176(.dina(n27248), .dinb(n26961), .dout(n27439));
  jxor g10177(.dina(n27132), .dinb(n27131), .dout(n27440));
  jor  g10178(.dina(n27440), .dinb(n27250), .dout(n27441));
  jand g10179(.dina(n27441), .dinb(n27439), .dout(n27442));
  jand g10180(.dina(n27442), .dinb(n264), .dout(n27443));
  jor  g10181(.dina(n27248), .dinb(n27128), .dout(n27444));
  jxor g10182(.dina(n27129), .dinb(n7731), .dout(n27445));
  jand g10183(.dina(n27445), .dinb(n27248), .dout(n27446));
  jnot g10184(.din(n27446), .dout(n27447));
  jand g10185(.dina(n27447), .dinb(n27444), .dout(n27448));
  jnot g10186(.din(n27448), .dout(n27449));
  jand g10187(.dina(n27449), .dinb(n386), .dout(n27450));
  jnot g10188(.din(n8054), .dout(n27451));
  jnot g10189(.din(n26773), .dout(n27452));
  jnot g10190(.din(n26777), .dout(n27453));
  jnot g10191(.din(n26782), .dout(n27454));
  jnot g10192(.din(n26787), .dout(n27455));
  jnot g10193(.din(n26792), .dout(n27456));
  jnot g10194(.din(n26797), .dout(n27457));
  jnot g10195(.din(n26802), .dout(n27458));
  jnot g10196(.din(n26807), .dout(n27459));
  jnot g10197(.din(n26812), .dout(n27460));
  jnot g10198(.din(n26817), .dout(n27461));
  jnot g10199(.din(n26822), .dout(n27462));
  jnot g10200(.din(n26827), .dout(n27463));
  jnot g10201(.din(n26832), .dout(n27464));
  jnot g10202(.din(n26837), .dout(n27465));
  jnot g10203(.din(n26842), .dout(n27466));
  jnot g10204(.din(n26847), .dout(n27467));
  jnot g10205(.din(n26852), .dout(n27468));
  jnot g10206(.din(n26857), .dout(n27469));
  jnot g10207(.din(n26862), .dout(n27470));
  jnot g10208(.din(n26867), .dout(n27471));
  jnot g10209(.din(n26872), .dout(n27472));
  jnot g10210(.din(n26877), .dout(n27473));
  jnot g10211(.din(n26882), .dout(n27474));
  jnot g10212(.din(n26887), .dout(n27475));
  jnot g10213(.din(n26892), .dout(n27476));
  jnot g10214(.din(n26897), .dout(n27477));
  jnot g10215(.din(n26902), .dout(n27478));
  jnot g10216(.din(n26907), .dout(n27479));
  jnot g10217(.din(n26912), .dout(n27480));
  jnot g10218(.din(n26917), .dout(n27481));
  jnot g10219(.din(n26922), .dout(n27482));
  jnot g10220(.din(n26927), .dout(n27483));
  jnot g10221(.din(n26932), .dout(n27484));
  jnot g10222(.din(n26937), .dout(n27485));
  jnot g10223(.din(n26942), .dout(n27486));
  jnot g10224(.din(n26947), .dout(n27487));
  jnot g10225(.din(n26952), .dout(n27488));
  jnot g10226(.din(n26957), .dout(n27489));
  jnot g10227(.din(n26962), .dout(n27490));
  jnot g10228(.din(n27125), .dout(n27491));
  jxor g10229(.dina(n27128), .dinb(n259), .dout(n27492));
  jor  g10230(.dina(n27492), .dinb(n7730), .dout(n27493));
  jand g10231(.dina(n27493), .dinb(n27491), .dout(n27494));
  jnot g10232(.din(n27132), .dout(n27495));
  jor  g10233(.dina(n27495), .dinb(n27494), .dout(n27496));
  jand g10234(.dina(n27496), .dinb(n27490), .dout(n27497));
  jnot g10235(.din(n27135), .dout(n27498));
  jor  g10236(.dina(n27498), .dinb(n27497), .dout(n27499));
  jand g10237(.dina(n27499), .dinb(n27489), .dout(n27500));
  jnot g10238(.din(n27138), .dout(n27501));
  jor  g10239(.dina(n27501), .dinb(n27500), .dout(n27502));
  jand g10240(.dina(n27502), .dinb(n27488), .dout(n27503));
  jnot g10241(.din(n27141), .dout(n27504));
  jor  g10242(.dina(n27504), .dinb(n27503), .dout(n27505));
  jand g10243(.dina(n27505), .dinb(n27487), .dout(n27506));
  jnot g10244(.din(n27144), .dout(n27507));
  jor  g10245(.dina(n27507), .dinb(n27506), .dout(n27508));
  jand g10246(.dina(n27508), .dinb(n27486), .dout(n27509));
  jnot g10247(.din(n27147), .dout(n27510));
  jor  g10248(.dina(n27510), .dinb(n27509), .dout(n27511));
  jand g10249(.dina(n27511), .dinb(n27485), .dout(n27512));
  jnot g10250(.din(n27150), .dout(n27513));
  jor  g10251(.dina(n27513), .dinb(n27512), .dout(n27514));
  jand g10252(.dina(n27514), .dinb(n27484), .dout(n27515));
  jnot g10253(.din(n27153), .dout(n27516));
  jor  g10254(.dina(n27516), .dinb(n27515), .dout(n27517));
  jand g10255(.dina(n27517), .dinb(n27483), .dout(n27518));
  jnot g10256(.din(n27156), .dout(n27519));
  jor  g10257(.dina(n27519), .dinb(n27518), .dout(n27520));
  jand g10258(.dina(n27520), .dinb(n27482), .dout(n27521));
  jnot g10259(.din(n27159), .dout(n27522));
  jor  g10260(.dina(n27522), .dinb(n27521), .dout(n27523));
  jand g10261(.dina(n27523), .dinb(n27481), .dout(n27524));
  jnot g10262(.din(n27162), .dout(n27525));
  jor  g10263(.dina(n27525), .dinb(n27524), .dout(n27526));
  jand g10264(.dina(n27526), .dinb(n27480), .dout(n27527));
  jnot g10265(.din(n27165), .dout(n27528));
  jor  g10266(.dina(n27528), .dinb(n27527), .dout(n27529));
  jand g10267(.dina(n27529), .dinb(n27479), .dout(n27530));
  jnot g10268(.din(n27168), .dout(n27531));
  jor  g10269(.dina(n27531), .dinb(n27530), .dout(n27532));
  jand g10270(.dina(n27532), .dinb(n27478), .dout(n27533));
  jnot g10271(.din(n27171), .dout(n27534));
  jor  g10272(.dina(n27534), .dinb(n27533), .dout(n27535));
  jand g10273(.dina(n27535), .dinb(n27477), .dout(n27536));
  jnot g10274(.din(n27174), .dout(n27537));
  jor  g10275(.dina(n27537), .dinb(n27536), .dout(n27538));
  jand g10276(.dina(n27538), .dinb(n27476), .dout(n27539));
  jnot g10277(.din(n27177), .dout(n27540));
  jor  g10278(.dina(n27540), .dinb(n27539), .dout(n27541));
  jand g10279(.dina(n27541), .dinb(n27475), .dout(n27542));
  jnot g10280(.din(n27180), .dout(n27543));
  jor  g10281(.dina(n27543), .dinb(n27542), .dout(n27544));
  jand g10282(.dina(n27544), .dinb(n27474), .dout(n27545));
  jnot g10283(.din(n27183), .dout(n27546));
  jor  g10284(.dina(n27546), .dinb(n27545), .dout(n27547));
  jand g10285(.dina(n27547), .dinb(n27473), .dout(n27548));
  jnot g10286(.din(n27186), .dout(n27549));
  jor  g10287(.dina(n27549), .dinb(n27548), .dout(n27550));
  jand g10288(.dina(n27550), .dinb(n27472), .dout(n27551));
  jnot g10289(.din(n27189), .dout(n27552));
  jor  g10290(.dina(n27552), .dinb(n27551), .dout(n27553));
  jand g10291(.dina(n27553), .dinb(n27471), .dout(n27554));
  jnot g10292(.din(n27192), .dout(n27555));
  jor  g10293(.dina(n27555), .dinb(n27554), .dout(n27556));
  jand g10294(.dina(n27556), .dinb(n27470), .dout(n27557));
  jnot g10295(.din(n27195), .dout(n27558));
  jor  g10296(.dina(n27558), .dinb(n27557), .dout(n27559));
  jand g10297(.dina(n27559), .dinb(n27469), .dout(n27560));
  jnot g10298(.din(n27198), .dout(n27561));
  jor  g10299(.dina(n27561), .dinb(n27560), .dout(n27562));
  jand g10300(.dina(n27562), .dinb(n27468), .dout(n27563));
  jnot g10301(.din(n27201), .dout(n27564));
  jor  g10302(.dina(n27564), .dinb(n27563), .dout(n27565));
  jand g10303(.dina(n27565), .dinb(n27467), .dout(n27566));
  jnot g10304(.din(n27204), .dout(n27567));
  jor  g10305(.dina(n27567), .dinb(n27566), .dout(n27568));
  jand g10306(.dina(n27568), .dinb(n27466), .dout(n27569));
  jnot g10307(.din(n27207), .dout(n27570));
  jor  g10308(.dina(n27570), .dinb(n27569), .dout(n27571));
  jand g10309(.dina(n27571), .dinb(n27465), .dout(n27572));
  jnot g10310(.din(n27210), .dout(n27573));
  jor  g10311(.dina(n27573), .dinb(n27572), .dout(n27574));
  jand g10312(.dina(n27574), .dinb(n27464), .dout(n27575));
  jnot g10313(.din(n27213), .dout(n27576));
  jor  g10314(.dina(n27576), .dinb(n27575), .dout(n27577));
  jand g10315(.dina(n27577), .dinb(n27463), .dout(n27578));
  jnot g10316(.din(n27216), .dout(n27579));
  jor  g10317(.dina(n27579), .dinb(n27578), .dout(n27580));
  jand g10318(.dina(n27580), .dinb(n27462), .dout(n27581));
  jnot g10319(.din(n27219), .dout(n27582));
  jor  g10320(.dina(n27582), .dinb(n27581), .dout(n27583));
  jand g10321(.dina(n27583), .dinb(n27461), .dout(n27584));
  jnot g10322(.din(n27222), .dout(n27585));
  jor  g10323(.dina(n27585), .dinb(n27584), .dout(n27586));
  jand g10324(.dina(n27586), .dinb(n27460), .dout(n27587));
  jnot g10325(.din(n27225), .dout(n27588));
  jor  g10326(.dina(n27588), .dinb(n27587), .dout(n27589));
  jand g10327(.dina(n27589), .dinb(n27459), .dout(n27590));
  jnot g10328(.din(n27228), .dout(n27591));
  jor  g10329(.dina(n27591), .dinb(n27590), .dout(n27592));
  jand g10330(.dina(n27592), .dinb(n27458), .dout(n27593));
  jnot g10331(.din(n27231), .dout(n27594));
  jor  g10332(.dina(n27594), .dinb(n27593), .dout(n27595));
  jand g10333(.dina(n27595), .dinb(n27457), .dout(n27596));
  jnot g10334(.din(n27234), .dout(n27597));
  jor  g10335(.dina(n27597), .dinb(n27596), .dout(n27598));
  jand g10336(.dina(n27598), .dinb(n27456), .dout(n27599));
  jnot g10337(.din(n27237), .dout(n27600));
  jor  g10338(.dina(n27600), .dinb(n27599), .dout(n27601));
  jand g10339(.dina(n27601), .dinb(n27455), .dout(n27602));
  jnot g10340(.din(n27240), .dout(n27603));
  jor  g10341(.dina(n27603), .dinb(n27602), .dout(n27604));
  jand g10342(.dina(n27604), .dinb(n27454), .dout(n27605));
  jnot g10343(.din(n27243), .dout(n27606));
  jor  g10344(.dina(n27606), .dinb(n27605), .dout(n27607));
  jand g10345(.dina(n27607), .dinb(n27453), .dout(n27608));
  jor  g10346(.dina(n27608), .dinb(n26775), .dout(n27609));
  jand g10347(.dina(n27609), .dinb(n27452), .dout(n27610));
  jor  g10348(.dina(n27610), .dinb(n27451), .dout(n27611));
  jand g10349(.dina(n27611), .dinb(a23 ), .dout(n27612));
  jnot g10350(.din(n8057), .dout(n27613));
  jor  g10351(.dina(n27610), .dinb(n27613), .dout(n27614));
  jnot g10352(.din(n27614), .dout(n27615));
  jor  g10353(.dina(n27615), .dinb(n27612), .dout(n27616));
  jand g10354(.dina(n27616), .dinb(n259), .dout(n27617));
  jand g10355(.dina(n27247), .dinb(n8054), .dout(n27618));
  jor  g10356(.dina(n27618), .dinb(n7729), .dout(n27619));
  jand g10357(.dina(n27614), .dinb(n27619), .dout(n27620));
  jxor g10358(.dina(n27620), .dinb(b1 ), .dout(n27621));
  jand g10359(.dina(n27621), .dinb(n8065), .dout(n27622));
  jor  g10360(.dina(n27622), .dinb(n27617), .dout(n27623));
  jxor g10361(.dina(n27448), .dinb(b2 ), .dout(n27624));
  jand g10362(.dina(n27624), .dinb(n27623), .dout(n27625));
  jor  g10363(.dina(n27625), .dinb(n27450), .dout(n27626));
  jxor g10364(.dina(n27442), .dinb(n264), .dout(n27627));
  jand g10365(.dina(n27627), .dinb(n27626), .dout(n27628));
  jor  g10366(.dina(n27628), .dinb(n27443), .dout(n27629));
  jxor g10367(.dina(n27437), .dinb(n376), .dout(n27630));
  jand g10368(.dina(n27630), .dinb(n27629), .dout(n27631));
  jor  g10369(.dina(n27631), .dinb(n27438), .dout(n27632));
  jxor g10370(.dina(n27432), .dinb(n377), .dout(n27633));
  jand g10371(.dina(n27633), .dinb(n27632), .dout(n27634));
  jor  g10372(.dina(n27634), .dinb(n27433), .dout(n27635));
  jxor g10373(.dina(n27427), .dinb(n378), .dout(n27636));
  jand g10374(.dina(n27636), .dinb(n27635), .dout(n27637));
  jor  g10375(.dina(n27637), .dinb(n27428), .dout(n27638));
  jxor g10376(.dina(n27422), .dinb(n265), .dout(n27639));
  jand g10377(.dina(n27639), .dinb(n27638), .dout(n27640));
  jor  g10378(.dina(n27640), .dinb(n27423), .dout(n27641));
  jxor g10379(.dina(n27417), .dinb(n367), .dout(n27642));
  jand g10380(.dina(n27642), .dinb(n27641), .dout(n27643));
  jor  g10381(.dina(n27643), .dinb(n27418), .dout(n27644));
  jxor g10382(.dina(n27412), .dinb(n368), .dout(n27645));
  jand g10383(.dina(n27645), .dinb(n27644), .dout(n27646));
  jor  g10384(.dina(n27646), .dinb(n27413), .dout(n27647));
  jxor g10385(.dina(n27407), .dinb(n369), .dout(n27648));
  jand g10386(.dina(n27648), .dinb(n27647), .dout(n27649));
  jor  g10387(.dina(n27649), .dinb(n27408), .dout(n27650));
  jxor g10388(.dina(n27402), .dinb(n359), .dout(n27651));
  jand g10389(.dina(n27651), .dinb(n27650), .dout(n27652));
  jor  g10390(.dina(n27652), .dinb(n27403), .dout(n27653));
  jxor g10391(.dina(n27397), .dinb(n363), .dout(n27654));
  jand g10392(.dina(n27654), .dinb(n27653), .dout(n27655));
  jor  g10393(.dina(n27655), .dinb(n27398), .dout(n27656));
  jxor g10394(.dina(n27392), .dinb(n360), .dout(n27657));
  jand g10395(.dina(n27657), .dinb(n27656), .dout(n27658));
  jor  g10396(.dina(n27658), .dinb(n27393), .dout(n27659));
  jxor g10397(.dina(n27387), .dinb(n361), .dout(n27660));
  jand g10398(.dina(n27660), .dinb(n27659), .dout(n27661));
  jor  g10399(.dina(n27661), .dinb(n27388), .dout(n27662));
  jxor g10400(.dina(n27382), .dinb(n364), .dout(n27663));
  jand g10401(.dina(n27663), .dinb(n27662), .dout(n27664));
  jor  g10402(.dina(n27664), .dinb(n27383), .dout(n27665));
  jxor g10403(.dina(n27377), .dinb(n355), .dout(n27666));
  jand g10404(.dina(n27666), .dinb(n27665), .dout(n27667));
  jor  g10405(.dina(n27667), .dinb(n27378), .dout(n27668));
  jxor g10406(.dina(n27372), .dinb(n356), .dout(n27669));
  jand g10407(.dina(n27669), .dinb(n27668), .dout(n27670));
  jor  g10408(.dina(n27670), .dinb(n27373), .dout(n27671));
  jxor g10409(.dina(n27367), .dinb(n266), .dout(n27672));
  jand g10410(.dina(n27672), .dinb(n27671), .dout(n27673));
  jor  g10411(.dina(n27673), .dinb(n27368), .dout(n27674));
  jxor g10412(.dina(n27362), .dinb(n267), .dout(n27675));
  jand g10413(.dina(n27675), .dinb(n27674), .dout(n27676));
  jor  g10414(.dina(n27676), .dinb(n27363), .dout(n27677));
  jxor g10415(.dina(n27357), .dinb(n347), .dout(n27678));
  jand g10416(.dina(n27678), .dinb(n27677), .dout(n27679));
  jor  g10417(.dina(n27679), .dinb(n27358), .dout(n27680));
  jxor g10418(.dina(n27352), .dinb(n348), .dout(n27681));
  jand g10419(.dina(n27681), .dinb(n27680), .dout(n27682));
  jor  g10420(.dina(n27682), .dinb(n27353), .dout(n27683));
  jxor g10421(.dina(n27347), .dinb(n349), .dout(n27684));
  jand g10422(.dina(n27684), .dinb(n27683), .dout(n27685));
  jor  g10423(.dina(n27685), .dinb(n27348), .dout(n27686));
  jxor g10424(.dina(n27342), .dinb(n268), .dout(n27687));
  jand g10425(.dina(n27687), .dinb(n27686), .dout(n27688));
  jor  g10426(.dina(n27688), .dinb(n27343), .dout(n27689));
  jxor g10427(.dina(n27337), .dinb(n274), .dout(n27690));
  jand g10428(.dina(n27690), .dinb(n27689), .dout(n27691));
  jor  g10429(.dina(n27691), .dinb(n27338), .dout(n27692));
  jxor g10430(.dina(n27332), .dinb(n269), .dout(n27693));
  jand g10431(.dina(n27693), .dinb(n27692), .dout(n27694));
  jor  g10432(.dina(n27694), .dinb(n27333), .dout(n27695));
  jxor g10433(.dina(n27327), .dinb(n270), .dout(n27696));
  jand g10434(.dina(n27696), .dinb(n27695), .dout(n27697));
  jor  g10435(.dina(n27697), .dinb(n27328), .dout(n27698));
  jxor g10436(.dina(n27322), .dinb(n271), .dout(n27699));
  jand g10437(.dina(n27699), .dinb(n27698), .dout(n27700));
  jor  g10438(.dina(n27700), .dinb(n27323), .dout(n27701));
  jxor g10439(.dina(n27317), .dinb(n338), .dout(n27702));
  jand g10440(.dina(n27702), .dinb(n27701), .dout(n27703));
  jor  g10441(.dina(n27703), .dinb(n27318), .dout(n27704));
  jxor g10442(.dina(n27312), .dinb(n339), .dout(n27705));
  jand g10443(.dina(n27705), .dinb(n27704), .dout(n27706));
  jor  g10444(.dina(n27706), .dinb(n27313), .dout(n27707));
  jxor g10445(.dina(n27307), .dinb(n340), .dout(n27708));
  jand g10446(.dina(n27708), .dinb(n27707), .dout(n27709));
  jor  g10447(.dina(n27709), .dinb(n27308), .dout(n27710));
  jxor g10448(.dina(n27302), .dinb(n275), .dout(n27711));
  jand g10449(.dina(n27711), .dinb(n27710), .dout(n27712));
  jor  g10450(.dina(n27712), .dinb(n27303), .dout(n27713));
  jxor g10451(.dina(n27297), .dinb(n331), .dout(n27714));
  jand g10452(.dina(n27714), .dinb(n27713), .dout(n27715));
  jor  g10453(.dina(n27715), .dinb(n27298), .dout(n27716));
  jxor g10454(.dina(n27292), .dinb(n332), .dout(n27717));
  jand g10455(.dina(n27717), .dinb(n27716), .dout(n27718));
  jor  g10456(.dina(n27718), .dinb(n27293), .dout(n27719));
  jxor g10457(.dina(n27287), .dinb(n333), .dout(n27720));
  jand g10458(.dina(n27720), .dinb(n27719), .dout(n27721));
  jor  g10459(.dina(n27721), .dinb(n27288), .dout(n27722));
  jxor g10460(.dina(n27282), .dinb(n276), .dout(n27723));
  jand g10461(.dina(n27723), .dinb(n27722), .dout(n27724));
  jor  g10462(.dina(n27724), .dinb(n27283), .dout(n27725));
  jxor g10463(.dina(n27277), .dinb(n324), .dout(n27726));
  jand g10464(.dina(n27726), .dinb(n27725), .dout(n27727));
  jor  g10465(.dina(n27727), .dinb(n27278), .dout(n27728));
  jxor g10466(.dina(n27272), .dinb(n325), .dout(n27729));
  jand g10467(.dina(n27729), .dinb(n27728), .dout(n27730));
  jor  g10468(.dina(n27730), .dinb(n27273), .dout(n27731));
  jxor g10469(.dina(n27267), .dinb(n326), .dout(n27732));
  jand g10470(.dina(n27732), .dinb(n27731), .dout(n27733));
  jor  g10471(.dina(n27733), .dinb(n27268), .dout(n27734));
  jxor g10472(.dina(n27262), .dinb(n277), .dout(n27735));
  jand g10473(.dina(n27735), .dinb(n27734), .dout(n27736));
  jor  g10474(.dina(n27736), .dinb(n27263), .dout(n27737));
  jxor g10475(.dina(n27253), .dinb(n278), .dout(n27738));
  jand g10476(.dina(n27738), .dinb(n27737), .dout(n27739));
  jor  g10477(.dina(n27739), .dinb(n27258), .dout(n27740));
  jxor g10478(.dina(n27256), .dinb(b41 ), .dout(n27741));
  jnot g10479(.din(n27741), .dout(n27742));
  jand g10480(.dina(n27742), .dinb(n27740), .dout(n27743));
  jand g10481(.dina(n27743), .dinb(n7526), .dout(n27744));
  jor  g10482(.dina(n27744), .dinb(n27257), .dout(n27745));
  jor  g10483(.dina(n27745), .dinb(n27253), .dout(n27746));
  jnot g10484(.din(n27257), .dout(n27747));
  jnot g10485(.din(n7526), .dout(n27748));
  jnot g10486(.din(n27258), .dout(n27749));
  jnot g10487(.din(n27263), .dout(n27750));
  jnot g10488(.din(n27268), .dout(n27751));
  jnot g10489(.din(n27273), .dout(n27752));
  jnot g10490(.din(n27278), .dout(n27753));
  jnot g10491(.din(n27283), .dout(n27754));
  jnot g10492(.din(n27288), .dout(n27755));
  jnot g10493(.din(n27293), .dout(n27756));
  jnot g10494(.din(n27298), .dout(n27757));
  jnot g10495(.din(n27303), .dout(n27758));
  jnot g10496(.din(n27308), .dout(n27759));
  jnot g10497(.din(n27313), .dout(n27760));
  jnot g10498(.din(n27318), .dout(n27761));
  jnot g10499(.din(n27323), .dout(n27762));
  jnot g10500(.din(n27328), .dout(n27763));
  jnot g10501(.din(n27333), .dout(n27764));
  jnot g10502(.din(n27338), .dout(n27765));
  jnot g10503(.din(n27343), .dout(n27766));
  jnot g10504(.din(n27348), .dout(n27767));
  jnot g10505(.din(n27353), .dout(n27768));
  jnot g10506(.din(n27358), .dout(n27769));
  jnot g10507(.din(n27363), .dout(n27770));
  jnot g10508(.din(n27368), .dout(n27771));
  jnot g10509(.din(n27373), .dout(n27772));
  jnot g10510(.din(n27378), .dout(n27773));
  jnot g10511(.din(n27383), .dout(n27774));
  jnot g10512(.din(n27388), .dout(n27775));
  jnot g10513(.din(n27393), .dout(n27776));
  jnot g10514(.din(n27398), .dout(n27777));
  jnot g10515(.din(n27403), .dout(n27778));
  jnot g10516(.din(n27408), .dout(n27779));
  jnot g10517(.din(n27413), .dout(n27780));
  jnot g10518(.din(n27418), .dout(n27781));
  jnot g10519(.din(n27423), .dout(n27782));
  jnot g10520(.din(n27428), .dout(n27783));
  jnot g10521(.din(n27433), .dout(n27784));
  jnot g10522(.din(n27438), .dout(n27785));
  jnot g10523(.din(n27443), .dout(n27786));
  jnot g10524(.din(n27450), .dout(n27787));
  jnot g10525(.din(n27617), .dout(n27788));
  jxor g10526(.dina(n27620), .dinb(n259), .dout(n27789));
  jor  g10527(.dina(n27789), .dinb(n8064), .dout(n27790));
  jand g10528(.dina(n27790), .dinb(n27788), .dout(n27791));
  jnot g10529(.din(n27624), .dout(n27792));
  jor  g10530(.dina(n27792), .dinb(n27791), .dout(n27793));
  jand g10531(.dina(n27793), .dinb(n27787), .dout(n27794));
  jnot g10532(.din(n27627), .dout(n27795));
  jor  g10533(.dina(n27795), .dinb(n27794), .dout(n27796));
  jand g10534(.dina(n27796), .dinb(n27786), .dout(n27797));
  jnot g10535(.din(n27630), .dout(n27798));
  jor  g10536(.dina(n27798), .dinb(n27797), .dout(n27799));
  jand g10537(.dina(n27799), .dinb(n27785), .dout(n27800));
  jnot g10538(.din(n27633), .dout(n27801));
  jor  g10539(.dina(n27801), .dinb(n27800), .dout(n27802));
  jand g10540(.dina(n27802), .dinb(n27784), .dout(n27803));
  jnot g10541(.din(n27636), .dout(n27804));
  jor  g10542(.dina(n27804), .dinb(n27803), .dout(n27805));
  jand g10543(.dina(n27805), .dinb(n27783), .dout(n27806));
  jnot g10544(.din(n27639), .dout(n27807));
  jor  g10545(.dina(n27807), .dinb(n27806), .dout(n27808));
  jand g10546(.dina(n27808), .dinb(n27782), .dout(n27809));
  jnot g10547(.din(n27642), .dout(n27810));
  jor  g10548(.dina(n27810), .dinb(n27809), .dout(n27811));
  jand g10549(.dina(n27811), .dinb(n27781), .dout(n27812));
  jnot g10550(.din(n27645), .dout(n27813));
  jor  g10551(.dina(n27813), .dinb(n27812), .dout(n27814));
  jand g10552(.dina(n27814), .dinb(n27780), .dout(n27815));
  jnot g10553(.din(n27648), .dout(n27816));
  jor  g10554(.dina(n27816), .dinb(n27815), .dout(n27817));
  jand g10555(.dina(n27817), .dinb(n27779), .dout(n27818));
  jnot g10556(.din(n27651), .dout(n27819));
  jor  g10557(.dina(n27819), .dinb(n27818), .dout(n27820));
  jand g10558(.dina(n27820), .dinb(n27778), .dout(n27821));
  jnot g10559(.din(n27654), .dout(n27822));
  jor  g10560(.dina(n27822), .dinb(n27821), .dout(n27823));
  jand g10561(.dina(n27823), .dinb(n27777), .dout(n27824));
  jnot g10562(.din(n27657), .dout(n27825));
  jor  g10563(.dina(n27825), .dinb(n27824), .dout(n27826));
  jand g10564(.dina(n27826), .dinb(n27776), .dout(n27827));
  jnot g10565(.din(n27660), .dout(n27828));
  jor  g10566(.dina(n27828), .dinb(n27827), .dout(n27829));
  jand g10567(.dina(n27829), .dinb(n27775), .dout(n27830));
  jnot g10568(.din(n27663), .dout(n27831));
  jor  g10569(.dina(n27831), .dinb(n27830), .dout(n27832));
  jand g10570(.dina(n27832), .dinb(n27774), .dout(n27833));
  jnot g10571(.din(n27666), .dout(n27834));
  jor  g10572(.dina(n27834), .dinb(n27833), .dout(n27835));
  jand g10573(.dina(n27835), .dinb(n27773), .dout(n27836));
  jnot g10574(.din(n27669), .dout(n27837));
  jor  g10575(.dina(n27837), .dinb(n27836), .dout(n27838));
  jand g10576(.dina(n27838), .dinb(n27772), .dout(n27839));
  jnot g10577(.din(n27672), .dout(n27840));
  jor  g10578(.dina(n27840), .dinb(n27839), .dout(n27841));
  jand g10579(.dina(n27841), .dinb(n27771), .dout(n27842));
  jnot g10580(.din(n27675), .dout(n27843));
  jor  g10581(.dina(n27843), .dinb(n27842), .dout(n27844));
  jand g10582(.dina(n27844), .dinb(n27770), .dout(n27845));
  jnot g10583(.din(n27678), .dout(n27846));
  jor  g10584(.dina(n27846), .dinb(n27845), .dout(n27847));
  jand g10585(.dina(n27847), .dinb(n27769), .dout(n27848));
  jnot g10586(.din(n27681), .dout(n27849));
  jor  g10587(.dina(n27849), .dinb(n27848), .dout(n27850));
  jand g10588(.dina(n27850), .dinb(n27768), .dout(n27851));
  jnot g10589(.din(n27684), .dout(n27852));
  jor  g10590(.dina(n27852), .dinb(n27851), .dout(n27853));
  jand g10591(.dina(n27853), .dinb(n27767), .dout(n27854));
  jnot g10592(.din(n27687), .dout(n27855));
  jor  g10593(.dina(n27855), .dinb(n27854), .dout(n27856));
  jand g10594(.dina(n27856), .dinb(n27766), .dout(n27857));
  jnot g10595(.din(n27690), .dout(n27858));
  jor  g10596(.dina(n27858), .dinb(n27857), .dout(n27859));
  jand g10597(.dina(n27859), .dinb(n27765), .dout(n27860));
  jnot g10598(.din(n27693), .dout(n27861));
  jor  g10599(.dina(n27861), .dinb(n27860), .dout(n27862));
  jand g10600(.dina(n27862), .dinb(n27764), .dout(n27863));
  jnot g10601(.din(n27696), .dout(n27864));
  jor  g10602(.dina(n27864), .dinb(n27863), .dout(n27865));
  jand g10603(.dina(n27865), .dinb(n27763), .dout(n27866));
  jnot g10604(.din(n27699), .dout(n27867));
  jor  g10605(.dina(n27867), .dinb(n27866), .dout(n27868));
  jand g10606(.dina(n27868), .dinb(n27762), .dout(n27869));
  jnot g10607(.din(n27702), .dout(n27870));
  jor  g10608(.dina(n27870), .dinb(n27869), .dout(n27871));
  jand g10609(.dina(n27871), .dinb(n27761), .dout(n27872));
  jnot g10610(.din(n27705), .dout(n27873));
  jor  g10611(.dina(n27873), .dinb(n27872), .dout(n27874));
  jand g10612(.dina(n27874), .dinb(n27760), .dout(n27875));
  jnot g10613(.din(n27708), .dout(n27876));
  jor  g10614(.dina(n27876), .dinb(n27875), .dout(n27877));
  jand g10615(.dina(n27877), .dinb(n27759), .dout(n27878));
  jnot g10616(.din(n27711), .dout(n27879));
  jor  g10617(.dina(n27879), .dinb(n27878), .dout(n27880));
  jand g10618(.dina(n27880), .dinb(n27758), .dout(n27881));
  jnot g10619(.din(n27714), .dout(n27882));
  jor  g10620(.dina(n27882), .dinb(n27881), .dout(n27883));
  jand g10621(.dina(n27883), .dinb(n27757), .dout(n27884));
  jnot g10622(.din(n27717), .dout(n27885));
  jor  g10623(.dina(n27885), .dinb(n27884), .dout(n27886));
  jand g10624(.dina(n27886), .dinb(n27756), .dout(n27887));
  jnot g10625(.din(n27720), .dout(n27888));
  jor  g10626(.dina(n27888), .dinb(n27887), .dout(n27889));
  jand g10627(.dina(n27889), .dinb(n27755), .dout(n27890));
  jnot g10628(.din(n27723), .dout(n27891));
  jor  g10629(.dina(n27891), .dinb(n27890), .dout(n27892));
  jand g10630(.dina(n27892), .dinb(n27754), .dout(n27893));
  jnot g10631(.din(n27726), .dout(n27894));
  jor  g10632(.dina(n27894), .dinb(n27893), .dout(n27895));
  jand g10633(.dina(n27895), .dinb(n27753), .dout(n27896));
  jnot g10634(.din(n27729), .dout(n27897));
  jor  g10635(.dina(n27897), .dinb(n27896), .dout(n27898));
  jand g10636(.dina(n27898), .dinb(n27752), .dout(n27899));
  jnot g10637(.din(n27732), .dout(n27900));
  jor  g10638(.dina(n27900), .dinb(n27899), .dout(n27901));
  jand g10639(.dina(n27901), .dinb(n27751), .dout(n27902));
  jnot g10640(.din(n27735), .dout(n27903));
  jor  g10641(.dina(n27903), .dinb(n27902), .dout(n27904));
  jand g10642(.dina(n27904), .dinb(n27750), .dout(n27905));
  jnot g10643(.din(n27738), .dout(n27906));
  jor  g10644(.dina(n27906), .dinb(n27905), .dout(n27907));
  jand g10645(.dina(n27907), .dinb(n27749), .dout(n27908));
  jor  g10646(.dina(n27741), .dinb(n27908), .dout(n27909));
  jor  g10647(.dina(n27909), .dinb(n27748), .dout(n27910));
  jand g10648(.dina(n27910), .dinb(n27747), .dout(n27911));
  jxor g10649(.dina(n27738), .dinb(n27737), .dout(n27912));
  jor  g10650(.dina(n27912), .dinb(n27911), .dout(n27913));
  jand g10651(.dina(n27913), .dinb(n27746), .dout(n27914));
  jxor g10652(.dina(n27741), .dinb(n27908), .dout(n27915));
  jand g10653(.dina(n27915), .dinb(n27257), .dout(n27916));
  jand g10654(.dina(n27911), .dinb(n27256), .dout(n27917));
  jor  g10655(.dina(n27917), .dinb(n27916), .dout(n27918));
  jand g10656(.dina(n27918), .dinb(n280), .dout(n27919));
  jnot g10657(.din(n27918), .dout(n27920));
  jand g10658(.dina(n27920), .dinb(b42 ), .dout(n27921));
  jnot g10659(.din(n27921), .dout(n27922));
  jand g10660(.dina(n27914), .dinb(n279), .dout(n27923));
  jor  g10661(.dina(n27745), .dinb(n27262), .dout(n27924));
  jxor g10662(.dina(n27735), .dinb(n27734), .dout(n27925));
  jor  g10663(.dina(n27925), .dinb(n27911), .dout(n27926));
  jand g10664(.dina(n27926), .dinb(n27924), .dout(n27927));
  jand g10665(.dina(n27927), .dinb(n278), .dout(n27928));
  jor  g10666(.dina(n27745), .dinb(n27267), .dout(n27929));
  jxor g10667(.dina(n27732), .dinb(n27731), .dout(n27930));
  jor  g10668(.dina(n27930), .dinb(n27911), .dout(n27931));
  jand g10669(.dina(n27931), .dinb(n27929), .dout(n27932));
  jand g10670(.dina(n27932), .dinb(n277), .dout(n27933));
  jor  g10671(.dina(n27745), .dinb(n27272), .dout(n27934));
  jxor g10672(.dina(n27729), .dinb(n27728), .dout(n27935));
  jor  g10673(.dina(n27935), .dinb(n27911), .dout(n27936));
  jand g10674(.dina(n27936), .dinb(n27934), .dout(n27937));
  jand g10675(.dina(n27937), .dinb(n326), .dout(n27938));
  jor  g10676(.dina(n27745), .dinb(n27277), .dout(n27939));
  jxor g10677(.dina(n27726), .dinb(n27725), .dout(n27940));
  jor  g10678(.dina(n27940), .dinb(n27911), .dout(n27941));
  jand g10679(.dina(n27941), .dinb(n27939), .dout(n27942));
  jand g10680(.dina(n27942), .dinb(n325), .dout(n27943));
  jor  g10681(.dina(n27745), .dinb(n27282), .dout(n27944));
  jxor g10682(.dina(n27723), .dinb(n27722), .dout(n27945));
  jor  g10683(.dina(n27945), .dinb(n27911), .dout(n27946));
  jand g10684(.dina(n27946), .dinb(n27944), .dout(n27947));
  jand g10685(.dina(n27947), .dinb(n324), .dout(n27948));
  jor  g10686(.dina(n27745), .dinb(n27287), .dout(n27949));
  jxor g10687(.dina(n27720), .dinb(n27719), .dout(n27950));
  jor  g10688(.dina(n27950), .dinb(n27911), .dout(n27951));
  jand g10689(.dina(n27951), .dinb(n27949), .dout(n27952));
  jand g10690(.dina(n27952), .dinb(n276), .dout(n27953));
  jor  g10691(.dina(n27745), .dinb(n27292), .dout(n27954));
  jxor g10692(.dina(n27717), .dinb(n27716), .dout(n27955));
  jor  g10693(.dina(n27955), .dinb(n27911), .dout(n27956));
  jand g10694(.dina(n27956), .dinb(n27954), .dout(n27957));
  jand g10695(.dina(n27957), .dinb(n333), .dout(n27958));
  jor  g10696(.dina(n27745), .dinb(n27297), .dout(n27959));
  jxor g10697(.dina(n27714), .dinb(n27713), .dout(n27960));
  jor  g10698(.dina(n27960), .dinb(n27911), .dout(n27961));
  jand g10699(.dina(n27961), .dinb(n27959), .dout(n27962));
  jand g10700(.dina(n27962), .dinb(n332), .dout(n27963));
  jor  g10701(.dina(n27745), .dinb(n27302), .dout(n27964));
  jxor g10702(.dina(n27711), .dinb(n27710), .dout(n27965));
  jor  g10703(.dina(n27965), .dinb(n27911), .dout(n27966));
  jand g10704(.dina(n27966), .dinb(n27964), .dout(n27967));
  jand g10705(.dina(n27967), .dinb(n331), .dout(n27968));
  jor  g10706(.dina(n27745), .dinb(n27307), .dout(n27969));
  jxor g10707(.dina(n27708), .dinb(n27707), .dout(n27970));
  jor  g10708(.dina(n27970), .dinb(n27911), .dout(n27971));
  jand g10709(.dina(n27971), .dinb(n27969), .dout(n27972));
  jand g10710(.dina(n27972), .dinb(n275), .dout(n27973));
  jor  g10711(.dina(n27745), .dinb(n27312), .dout(n27974));
  jxor g10712(.dina(n27705), .dinb(n27704), .dout(n27975));
  jor  g10713(.dina(n27975), .dinb(n27911), .dout(n27976));
  jand g10714(.dina(n27976), .dinb(n27974), .dout(n27977));
  jand g10715(.dina(n27977), .dinb(n340), .dout(n27978));
  jor  g10716(.dina(n27745), .dinb(n27317), .dout(n27979));
  jxor g10717(.dina(n27702), .dinb(n27701), .dout(n27980));
  jor  g10718(.dina(n27980), .dinb(n27911), .dout(n27981));
  jand g10719(.dina(n27981), .dinb(n27979), .dout(n27982));
  jand g10720(.dina(n27982), .dinb(n339), .dout(n27983));
  jor  g10721(.dina(n27745), .dinb(n27322), .dout(n27984));
  jxor g10722(.dina(n27699), .dinb(n27698), .dout(n27985));
  jor  g10723(.dina(n27985), .dinb(n27911), .dout(n27986));
  jand g10724(.dina(n27986), .dinb(n27984), .dout(n27987));
  jand g10725(.dina(n27987), .dinb(n338), .dout(n27988));
  jor  g10726(.dina(n27745), .dinb(n27327), .dout(n27989));
  jxor g10727(.dina(n27696), .dinb(n27695), .dout(n27990));
  jor  g10728(.dina(n27990), .dinb(n27911), .dout(n27991));
  jand g10729(.dina(n27991), .dinb(n27989), .dout(n27992));
  jand g10730(.dina(n27992), .dinb(n271), .dout(n27993));
  jor  g10731(.dina(n27745), .dinb(n27332), .dout(n27994));
  jxor g10732(.dina(n27693), .dinb(n27692), .dout(n27995));
  jor  g10733(.dina(n27995), .dinb(n27911), .dout(n27996));
  jand g10734(.dina(n27996), .dinb(n27994), .dout(n27997));
  jand g10735(.dina(n27997), .dinb(n270), .dout(n27998));
  jor  g10736(.dina(n27745), .dinb(n27337), .dout(n27999));
  jxor g10737(.dina(n27690), .dinb(n27689), .dout(n28000));
  jor  g10738(.dina(n28000), .dinb(n27911), .dout(n28001));
  jand g10739(.dina(n28001), .dinb(n27999), .dout(n28002));
  jand g10740(.dina(n28002), .dinb(n269), .dout(n28003));
  jor  g10741(.dina(n27745), .dinb(n27342), .dout(n28004));
  jxor g10742(.dina(n27687), .dinb(n27686), .dout(n28005));
  jor  g10743(.dina(n28005), .dinb(n27911), .dout(n28006));
  jand g10744(.dina(n28006), .dinb(n28004), .dout(n28007));
  jand g10745(.dina(n28007), .dinb(n274), .dout(n28008));
  jor  g10746(.dina(n27745), .dinb(n27347), .dout(n28009));
  jxor g10747(.dina(n27684), .dinb(n27683), .dout(n28010));
  jor  g10748(.dina(n28010), .dinb(n27911), .dout(n28011));
  jand g10749(.dina(n28011), .dinb(n28009), .dout(n28012));
  jand g10750(.dina(n28012), .dinb(n268), .dout(n28013));
  jor  g10751(.dina(n27745), .dinb(n27352), .dout(n28014));
  jxor g10752(.dina(n27681), .dinb(n27680), .dout(n28015));
  jor  g10753(.dina(n28015), .dinb(n27911), .dout(n28016));
  jand g10754(.dina(n28016), .dinb(n28014), .dout(n28017));
  jand g10755(.dina(n28017), .dinb(n349), .dout(n28018));
  jor  g10756(.dina(n27745), .dinb(n27357), .dout(n28019));
  jxor g10757(.dina(n27678), .dinb(n27677), .dout(n28020));
  jor  g10758(.dina(n28020), .dinb(n27911), .dout(n28021));
  jand g10759(.dina(n28021), .dinb(n28019), .dout(n28022));
  jand g10760(.dina(n28022), .dinb(n348), .dout(n28023));
  jor  g10761(.dina(n27745), .dinb(n27362), .dout(n28024));
  jxor g10762(.dina(n27675), .dinb(n27674), .dout(n28025));
  jor  g10763(.dina(n28025), .dinb(n27911), .dout(n28026));
  jand g10764(.dina(n28026), .dinb(n28024), .dout(n28027));
  jand g10765(.dina(n28027), .dinb(n347), .dout(n28028));
  jor  g10766(.dina(n27745), .dinb(n27367), .dout(n28029));
  jxor g10767(.dina(n27672), .dinb(n27671), .dout(n28030));
  jor  g10768(.dina(n28030), .dinb(n27911), .dout(n28031));
  jand g10769(.dina(n28031), .dinb(n28029), .dout(n28032));
  jand g10770(.dina(n28032), .dinb(n267), .dout(n28033));
  jor  g10771(.dina(n27745), .dinb(n27372), .dout(n28034));
  jxor g10772(.dina(n27669), .dinb(n27668), .dout(n28035));
  jor  g10773(.dina(n28035), .dinb(n27911), .dout(n28036));
  jand g10774(.dina(n28036), .dinb(n28034), .dout(n28037));
  jand g10775(.dina(n28037), .dinb(n266), .dout(n28038));
  jor  g10776(.dina(n27745), .dinb(n27377), .dout(n28039));
  jxor g10777(.dina(n27666), .dinb(n27665), .dout(n28040));
  jor  g10778(.dina(n28040), .dinb(n27911), .dout(n28041));
  jand g10779(.dina(n28041), .dinb(n28039), .dout(n28042));
  jand g10780(.dina(n28042), .dinb(n356), .dout(n28043));
  jor  g10781(.dina(n27745), .dinb(n27382), .dout(n28044));
  jxor g10782(.dina(n27663), .dinb(n27662), .dout(n28045));
  jor  g10783(.dina(n28045), .dinb(n27911), .dout(n28046));
  jand g10784(.dina(n28046), .dinb(n28044), .dout(n28047));
  jand g10785(.dina(n28047), .dinb(n355), .dout(n28048));
  jor  g10786(.dina(n27745), .dinb(n27387), .dout(n28049));
  jxor g10787(.dina(n27660), .dinb(n27659), .dout(n28050));
  jor  g10788(.dina(n28050), .dinb(n27911), .dout(n28051));
  jand g10789(.dina(n28051), .dinb(n28049), .dout(n28052));
  jand g10790(.dina(n28052), .dinb(n364), .dout(n28053));
  jor  g10791(.dina(n27745), .dinb(n27392), .dout(n28054));
  jxor g10792(.dina(n27657), .dinb(n27656), .dout(n28055));
  jor  g10793(.dina(n28055), .dinb(n27911), .dout(n28056));
  jand g10794(.dina(n28056), .dinb(n28054), .dout(n28057));
  jand g10795(.dina(n28057), .dinb(n361), .dout(n28058));
  jor  g10796(.dina(n27745), .dinb(n27397), .dout(n28059));
  jxor g10797(.dina(n27654), .dinb(n27653), .dout(n28060));
  jor  g10798(.dina(n28060), .dinb(n27911), .dout(n28061));
  jand g10799(.dina(n28061), .dinb(n28059), .dout(n28062));
  jand g10800(.dina(n28062), .dinb(n360), .dout(n28063));
  jor  g10801(.dina(n27745), .dinb(n27402), .dout(n28064));
  jxor g10802(.dina(n27651), .dinb(n27650), .dout(n28065));
  jor  g10803(.dina(n28065), .dinb(n27911), .dout(n28066));
  jand g10804(.dina(n28066), .dinb(n28064), .dout(n28067));
  jand g10805(.dina(n28067), .dinb(n363), .dout(n28068));
  jor  g10806(.dina(n27745), .dinb(n27407), .dout(n28069));
  jxor g10807(.dina(n27648), .dinb(n27647), .dout(n28070));
  jor  g10808(.dina(n28070), .dinb(n27911), .dout(n28071));
  jand g10809(.dina(n28071), .dinb(n28069), .dout(n28072));
  jand g10810(.dina(n28072), .dinb(n359), .dout(n28073));
  jor  g10811(.dina(n27745), .dinb(n27412), .dout(n28074));
  jxor g10812(.dina(n27645), .dinb(n27644), .dout(n28075));
  jor  g10813(.dina(n28075), .dinb(n27911), .dout(n28076));
  jand g10814(.dina(n28076), .dinb(n28074), .dout(n28077));
  jand g10815(.dina(n28077), .dinb(n369), .dout(n28078));
  jor  g10816(.dina(n27745), .dinb(n27417), .dout(n28079));
  jxor g10817(.dina(n27642), .dinb(n27641), .dout(n28080));
  jor  g10818(.dina(n28080), .dinb(n27911), .dout(n28081));
  jand g10819(.dina(n28081), .dinb(n28079), .dout(n28082));
  jand g10820(.dina(n28082), .dinb(n368), .dout(n28083));
  jor  g10821(.dina(n27745), .dinb(n27422), .dout(n28084));
  jxor g10822(.dina(n27639), .dinb(n27638), .dout(n28085));
  jor  g10823(.dina(n28085), .dinb(n27911), .dout(n28086));
  jand g10824(.dina(n28086), .dinb(n28084), .dout(n28087));
  jand g10825(.dina(n28087), .dinb(n367), .dout(n28088));
  jor  g10826(.dina(n27745), .dinb(n27427), .dout(n28089));
  jxor g10827(.dina(n27636), .dinb(n27635), .dout(n28090));
  jor  g10828(.dina(n28090), .dinb(n27911), .dout(n28091));
  jand g10829(.dina(n28091), .dinb(n28089), .dout(n28092));
  jand g10830(.dina(n28092), .dinb(n265), .dout(n28093));
  jor  g10831(.dina(n27745), .dinb(n27432), .dout(n28094));
  jxor g10832(.dina(n27633), .dinb(n27632), .dout(n28095));
  jor  g10833(.dina(n28095), .dinb(n27911), .dout(n28096));
  jand g10834(.dina(n28096), .dinb(n28094), .dout(n28097));
  jand g10835(.dina(n28097), .dinb(n378), .dout(n28098));
  jor  g10836(.dina(n27745), .dinb(n27437), .dout(n28099));
  jxor g10837(.dina(n27630), .dinb(n27629), .dout(n28100));
  jor  g10838(.dina(n28100), .dinb(n27911), .dout(n28101));
  jand g10839(.dina(n28101), .dinb(n28099), .dout(n28102));
  jand g10840(.dina(n28102), .dinb(n377), .dout(n28103));
  jor  g10841(.dina(n27745), .dinb(n27442), .dout(n28104));
  jxor g10842(.dina(n27627), .dinb(n27626), .dout(n28105));
  jor  g10843(.dina(n28105), .dinb(n27911), .dout(n28106));
  jand g10844(.dina(n28106), .dinb(n28104), .dout(n28107));
  jand g10845(.dina(n28107), .dinb(n376), .dout(n28108));
  jor  g10846(.dina(n27745), .dinb(n27449), .dout(n28109));
  jxor g10847(.dina(n27624), .dinb(n27623), .dout(n28110));
  jor  g10848(.dina(n28110), .dinb(n27911), .dout(n28111));
  jand g10849(.dina(n28111), .dinb(n28109), .dout(n28112));
  jand g10850(.dina(n28112), .dinb(n264), .dout(n28113));
  jand g10851(.dina(n27789), .dinb(n8064), .dout(n28114));
  jor  g10852(.dina(n27911), .dinb(n27622), .dout(n28115));
  jor  g10853(.dina(n28115), .dinb(n28114), .dout(n28116));
  jand g10854(.dina(n27911), .dinb(n27616), .dout(n28117));
  jnot g10855(.din(n28117), .dout(n28118));
  jand g10856(.dina(n28118), .dinb(n28116), .dout(n28119));
  jor  g10857(.dina(n28119), .dinb(b2 ), .dout(n28120));
  jnot g10858(.din(n28120), .dout(n28121));
  jand g10859(.dina(n27745), .dinb(b0 ), .dout(n28122));
  jxor g10860(.dina(n28122), .dinb(a22 ), .dout(n28123));
  jand g10861(.dina(n28123), .dinb(n259), .dout(n28124));
  jxor g10862(.dina(n28122), .dinb(n8063), .dout(n28125));
  jxor g10863(.dina(n28125), .dinb(b1 ), .dout(n28126));
  jand g10864(.dina(n28126), .dinb(n8617), .dout(n28127));
  jor  g10865(.dina(n28127), .dinb(n28124), .dout(n28128));
  jxor g10866(.dina(n28119), .dinb(b2 ), .dout(n28129));
  jand g10867(.dina(n28129), .dinb(n28128), .dout(n28130));
  jor  g10868(.dina(n28130), .dinb(n28121), .dout(n28131));
  jxor g10869(.dina(n28112), .dinb(n264), .dout(n28132));
  jand g10870(.dina(n28132), .dinb(n28131), .dout(n28133));
  jor  g10871(.dina(n28133), .dinb(n28113), .dout(n28134));
  jxor g10872(.dina(n28107), .dinb(n376), .dout(n28135));
  jand g10873(.dina(n28135), .dinb(n28134), .dout(n28136));
  jor  g10874(.dina(n28136), .dinb(n28108), .dout(n28137));
  jxor g10875(.dina(n28102), .dinb(n377), .dout(n28138));
  jand g10876(.dina(n28138), .dinb(n28137), .dout(n28139));
  jor  g10877(.dina(n28139), .dinb(n28103), .dout(n28140));
  jxor g10878(.dina(n28097), .dinb(n378), .dout(n28141));
  jand g10879(.dina(n28141), .dinb(n28140), .dout(n28142));
  jor  g10880(.dina(n28142), .dinb(n28098), .dout(n28143));
  jxor g10881(.dina(n28092), .dinb(n265), .dout(n28144));
  jand g10882(.dina(n28144), .dinb(n28143), .dout(n28145));
  jor  g10883(.dina(n28145), .dinb(n28093), .dout(n28146));
  jxor g10884(.dina(n28087), .dinb(n367), .dout(n28147));
  jand g10885(.dina(n28147), .dinb(n28146), .dout(n28148));
  jor  g10886(.dina(n28148), .dinb(n28088), .dout(n28149));
  jxor g10887(.dina(n28082), .dinb(n368), .dout(n28150));
  jand g10888(.dina(n28150), .dinb(n28149), .dout(n28151));
  jor  g10889(.dina(n28151), .dinb(n28083), .dout(n28152));
  jxor g10890(.dina(n28077), .dinb(n369), .dout(n28153));
  jand g10891(.dina(n28153), .dinb(n28152), .dout(n28154));
  jor  g10892(.dina(n28154), .dinb(n28078), .dout(n28155));
  jxor g10893(.dina(n28072), .dinb(n359), .dout(n28156));
  jand g10894(.dina(n28156), .dinb(n28155), .dout(n28157));
  jor  g10895(.dina(n28157), .dinb(n28073), .dout(n28158));
  jxor g10896(.dina(n28067), .dinb(n363), .dout(n28159));
  jand g10897(.dina(n28159), .dinb(n28158), .dout(n28160));
  jor  g10898(.dina(n28160), .dinb(n28068), .dout(n28161));
  jxor g10899(.dina(n28062), .dinb(n360), .dout(n28162));
  jand g10900(.dina(n28162), .dinb(n28161), .dout(n28163));
  jor  g10901(.dina(n28163), .dinb(n28063), .dout(n28164));
  jxor g10902(.dina(n28057), .dinb(n361), .dout(n28165));
  jand g10903(.dina(n28165), .dinb(n28164), .dout(n28166));
  jor  g10904(.dina(n28166), .dinb(n28058), .dout(n28167));
  jxor g10905(.dina(n28052), .dinb(n364), .dout(n28168));
  jand g10906(.dina(n28168), .dinb(n28167), .dout(n28169));
  jor  g10907(.dina(n28169), .dinb(n28053), .dout(n28170));
  jxor g10908(.dina(n28047), .dinb(n355), .dout(n28171));
  jand g10909(.dina(n28171), .dinb(n28170), .dout(n28172));
  jor  g10910(.dina(n28172), .dinb(n28048), .dout(n28173));
  jxor g10911(.dina(n28042), .dinb(n356), .dout(n28174));
  jand g10912(.dina(n28174), .dinb(n28173), .dout(n28175));
  jor  g10913(.dina(n28175), .dinb(n28043), .dout(n28176));
  jxor g10914(.dina(n28037), .dinb(n266), .dout(n28177));
  jand g10915(.dina(n28177), .dinb(n28176), .dout(n28178));
  jor  g10916(.dina(n28178), .dinb(n28038), .dout(n28179));
  jxor g10917(.dina(n28032), .dinb(n267), .dout(n28180));
  jand g10918(.dina(n28180), .dinb(n28179), .dout(n28181));
  jor  g10919(.dina(n28181), .dinb(n28033), .dout(n28182));
  jxor g10920(.dina(n28027), .dinb(n347), .dout(n28183));
  jand g10921(.dina(n28183), .dinb(n28182), .dout(n28184));
  jor  g10922(.dina(n28184), .dinb(n28028), .dout(n28185));
  jxor g10923(.dina(n28022), .dinb(n348), .dout(n28186));
  jand g10924(.dina(n28186), .dinb(n28185), .dout(n28187));
  jor  g10925(.dina(n28187), .dinb(n28023), .dout(n28188));
  jxor g10926(.dina(n28017), .dinb(n349), .dout(n28189));
  jand g10927(.dina(n28189), .dinb(n28188), .dout(n28190));
  jor  g10928(.dina(n28190), .dinb(n28018), .dout(n28191));
  jxor g10929(.dina(n28012), .dinb(n268), .dout(n28192));
  jand g10930(.dina(n28192), .dinb(n28191), .dout(n28193));
  jor  g10931(.dina(n28193), .dinb(n28013), .dout(n28194));
  jxor g10932(.dina(n28007), .dinb(n274), .dout(n28195));
  jand g10933(.dina(n28195), .dinb(n28194), .dout(n28196));
  jor  g10934(.dina(n28196), .dinb(n28008), .dout(n28197));
  jxor g10935(.dina(n28002), .dinb(n269), .dout(n28198));
  jand g10936(.dina(n28198), .dinb(n28197), .dout(n28199));
  jor  g10937(.dina(n28199), .dinb(n28003), .dout(n28200));
  jxor g10938(.dina(n27997), .dinb(n270), .dout(n28201));
  jand g10939(.dina(n28201), .dinb(n28200), .dout(n28202));
  jor  g10940(.dina(n28202), .dinb(n27998), .dout(n28203));
  jxor g10941(.dina(n27992), .dinb(n271), .dout(n28204));
  jand g10942(.dina(n28204), .dinb(n28203), .dout(n28205));
  jor  g10943(.dina(n28205), .dinb(n27993), .dout(n28206));
  jxor g10944(.dina(n27987), .dinb(n338), .dout(n28207));
  jand g10945(.dina(n28207), .dinb(n28206), .dout(n28208));
  jor  g10946(.dina(n28208), .dinb(n27988), .dout(n28209));
  jxor g10947(.dina(n27982), .dinb(n339), .dout(n28210));
  jand g10948(.dina(n28210), .dinb(n28209), .dout(n28211));
  jor  g10949(.dina(n28211), .dinb(n27983), .dout(n28212));
  jxor g10950(.dina(n27977), .dinb(n340), .dout(n28213));
  jand g10951(.dina(n28213), .dinb(n28212), .dout(n28214));
  jor  g10952(.dina(n28214), .dinb(n27978), .dout(n28215));
  jxor g10953(.dina(n27972), .dinb(n275), .dout(n28216));
  jand g10954(.dina(n28216), .dinb(n28215), .dout(n28217));
  jor  g10955(.dina(n28217), .dinb(n27973), .dout(n28218));
  jxor g10956(.dina(n27967), .dinb(n331), .dout(n28219));
  jand g10957(.dina(n28219), .dinb(n28218), .dout(n28220));
  jor  g10958(.dina(n28220), .dinb(n27968), .dout(n28221));
  jxor g10959(.dina(n27962), .dinb(n332), .dout(n28222));
  jand g10960(.dina(n28222), .dinb(n28221), .dout(n28223));
  jor  g10961(.dina(n28223), .dinb(n27963), .dout(n28224));
  jxor g10962(.dina(n27957), .dinb(n333), .dout(n28225));
  jand g10963(.dina(n28225), .dinb(n28224), .dout(n28226));
  jor  g10964(.dina(n28226), .dinb(n27958), .dout(n28227));
  jxor g10965(.dina(n27952), .dinb(n276), .dout(n28228));
  jand g10966(.dina(n28228), .dinb(n28227), .dout(n28229));
  jor  g10967(.dina(n28229), .dinb(n27953), .dout(n28230));
  jxor g10968(.dina(n27947), .dinb(n324), .dout(n28231));
  jand g10969(.dina(n28231), .dinb(n28230), .dout(n28232));
  jor  g10970(.dina(n28232), .dinb(n27948), .dout(n28233));
  jxor g10971(.dina(n27942), .dinb(n325), .dout(n28234));
  jand g10972(.dina(n28234), .dinb(n28233), .dout(n28235));
  jor  g10973(.dina(n28235), .dinb(n27943), .dout(n28236));
  jxor g10974(.dina(n27937), .dinb(n326), .dout(n28237));
  jand g10975(.dina(n28237), .dinb(n28236), .dout(n28238));
  jor  g10976(.dina(n28238), .dinb(n27938), .dout(n28239));
  jxor g10977(.dina(n27932), .dinb(n277), .dout(n28240));
  jand g10978(.dina(n28240), .dinb(n28239), .dout(n28241));
  jor  g10979(.dina(n28241), .dinb(n27933), .dout(n28242));
  jxor g10980(.dina(n27927), .dinb(n278), .dout(n28243));
  jand g10981(.dina(n28243), .dinb(n28242), .dout(n28244));
  jor  g10982(.dina(n28244), .dinb(n27928), .dout(n28245));
  jxor g10983(.dina(n27914), .dinb(n279), .dout(n28246));
  jand g10984(.dina(n28246), .dinb(n28245), .dout(n28247));
  jor  g10985(.dina(n28247), .dinb(n27923), .dout(n28248));
  jand g10986(.dina(n28248), .dinb(n27922), .dout(n28249));
  jor  g10987(.dina(n28249), .dinb(n27919), .dout(n28250));
  jand g10988(.dina(n28250), .dinb(n405), .dout(n28251));
  jor  g10989(.dina(n28251), .dinb(n27914), .dout(n28252));
  jnot g10990(.din(n27919), .dout(n28253));
  jnot g10991(.din(n27923), .dout(n28254));
  jnot g10992(.din(n27928), .dout(n28255));
  jnot g10993(.din(n27933), .dout(n28256));
  jnot g10994(.din(n27938), .dout(n28257));
  jnot g10995(.din(n27943), .dout(n28258));
  jnot g10996(.din(n27948), .dout(n28259));
  jnot g10997(.din(n27953), .dout(n28260));
  jnot g10998(.din(n27958), .dout(n28261));
  jnot g10999(.din(n27963), .dout(n28262));
  jnot g11000(.din(n27968), .dout(n28263));
  jnot g11001(.din(n27973), .dout(n28264));
  jnot g11002(.din(n27978), .dout(n28265));
  jnot g11003(.din(n27983), .dout(n28266));
  jnot g11004(.din(n27988), .dout(n28267));
  jnot g11005(.din(n27993), .dout(n28268));
  jnot g11006(.din(n27998), .dout(n28269));
  jnot g11007(.din(n28003), .dout(n28270));
  jnot g11008(.din(n28008), .dout(n28271));
  jnot g11009(.din(n28013), .dout(n28272));
  jnot g11010(.din(n28018), .dout(n28273));
  jnot g11011(.din(n28023), .dout(n28274));
  jnot g11012(.din(n28028), .dout(n28275));
  jnot g11013(.din(n28033), .dout(n28276));
  jnot g11014(.din(n28038), .dout(n28277));
  jnot g11015(.din(n28043), .dout(n28278));
  jnot g11016(.din(n28048), .dout(n28279));
  jnot g11017(.din(n28053), .dout(n28280));
  jnot g11018(.din(n28058), .dout(n28281));
  jnot g11019(.din(n28063), .dout(n28282));
  jnot g11020(.din(n28068), .dout(n28283));
  jnot g11021(.din(n28073), .dout(n28284));
  jnot g11022(.din(n28078), .dout(n28285));
  jnot g11023(.din(n28083), .dout(n28286));
  jnot g11024(.din(n28088), .dout(n28287));
  jnot g11025(.din(n28093), .dout(n28288));
  jnot g11026(.din(n28098), .dout(n28289));
  jnot g11027(.din(n28103), .dout(n28290));
  jnot g11028(.din(n28108), .dout(n28291));
  jnot g11029(.din(n28113), .dout(n28292));
  jor  g11030(.dina(n28125), .dinb(b1 ), .dout(n28293));
  jxor g11031(.dina(n28125), .dinb(n259), .dout(n28294));
  jor  g11032(.dina(n28294), .dinb(n8447), .dout(n28295));
  jand g11033(.dina(n28295), .dinb(n28293), .dout(n28296));
  jxor g11034(.dina(n28119), .dinb(n386), .dout(n28297));
  jor  g11035(.dina(n28297), .dinb(n28296), .dout(n28298));
  jand g11036(.dina(n28298), .dinb(n28120), .dout(n28299));
  jnot g11037(.din(n28132), .dout(n28300));
  jor  g11038(.dina(n28300), .dinb(n28299), .dout(n28301));
  jand g11039(.dina(n28301), .dinb(n28292), .dout(n28302));
  jnot g11040(.din(n28135), .dout(n28303));
  jor  g11041(.dina(n28303), .dinb(n28302), .dout(n28304));
  jand g11042(.dina(n28304), .dinb(n28291), .dout(n28305));
  jnot g11043(.din(n28138), .dout(n28306));
  jor  g11044(.dina(n28306), .dinb(n28305), .dout(n28307));
  jand g11045(.dina(n28307), .dinb(n28290), .dout(n28308));
  jnot g11046(.din(n28141), .dout(n28309));
  jor  g11047(.dina(n28309), .dinb(n28308), .dout(n28310));
  jand g11048(.dina(n28310), .dinb(n28289), .dout(n28311));
  jnot g11049(.din(n28144), .dout(n28312));
  jor  g11050(.dina(n28312), .dinb(n28311), .dout(n28313));
  jand g11051(.dina(n28313), .dinb(n28288), .dout(n28314));
  jnot g11052(.din(n28147), .dout(n28315));
  jor  g11053(.dina(n28315), .dinb(n28314), .dout(n28316));
  jand g11054(.dina(n28316), .dinb(n28287), .dout(n28317));
  jnot g11055(.din(n28150), .dout(n28318));
  jor  g11056(.dina(n28318), .dinb(n28317), .dout(n28319));
  jand g11057(.dina(n28319), .dinb(n28286), .dout(n28320));
  jnot g11058(.din(n28153), .dout(n28321));
  jor  g11059(.dina(n28321), .dinb(n28320), .dout(n28322));
  jand g11060(.dina(n28322), .dinb(n28285), .dout(n28323));
  jnot g11061(.din(n28156), .dout(n28324));
  jor  g11062(.dina(n28324), .dinb(n28323), .dout(n28325));
  jand g11063(.dina(n28325), .dinb(n28284), .dout(n28326));
  jnot g11064(.din(n28159), .dout(n28327));
  jor  g11065(.dina(n28327), .dinb(n28326), .dout(n28328));
  jand g11066(.dina(n28328), .dinb(n28283), .dout(n28329));
  jnot g11067(.din(n28162), .dout(n28330));
  jor  g11068(.dina(n28330), .dinb(n28329), .dout(n28331));
  jand g11069(.dina(n28331), .dinb(n28282), .dout(n28332));
  jnot g11070(.din(n28165), .dout(n28333));
  jor  g11071(.dina(n28333), .dinb(n28332), .dout(n28334));
  jand g11072(.dina(n28334), .dinb(n28281), .dout(n28335));
  jnot g11073(.din(n28168), .dout(n28336));
  jor  g11074(.dina(n28336), .dinb(n28335), .dout(n28337));
  jand g11075(.dina(n28337), .dinb(n28280), .dout(n28338));
  jnot g11076(.din(n28171), .dout(n28339));
  jor  g11077(.dina(n28339), .dinb(n28338), .dout(n28340));
  jand g11078(.dina(n28340), .dinb(n28279), .dout(n28341));
  jnot g11079(.din(n28174), .dout(n28342));
  jor  g11080(.dina(n28342), .dinb(n28341), .dout(n28343));
  jand g11081(.dina(n28343), .dinb(n28278), .dout(n28344));
  jnot g11082(.din(n28177), .dout(n28345));
  jor  g11083(.dina(n28345), .dinb(n28344), .dout(n28346));
  jand g11084(.dina(n28346), .dinb(n28277), .dout(n28347));
  jnot g11085(.din(n28180), .dout(n28348));
  jor  g11086(.dina(n28348), .dinb(n28347), .dout(n28349));
  jand g11087(.dina(n28349), .dinb(n28276), .dout(n28350));
  jnot g11088(.din(n28183), .dout(n28351));
  jor  g11089(.dina(n28351), .dinb(n28350), .dout(n28352));
  jand g11090(.dina(n28352), .dinb(n28275), .dout(n28353));
  jnot g11091(.din(n28186), .dout(n28354));
  jor  g11092(.dina(n28354), .dinb(n28353), .dout(n28355));
  jand g11093(.dina(n28355), .dinb(n28274), .dout(n28356));
  jnot g11094(.din(n28189), .dout(n28357));
  jor  g11095(.dina(n28357), .dinb(n28356), .dout(n28358));
  jand g11096(.dina(n28358), .dinb(n28273), .dout(n28359));
  jnot g11097(.din(n28192), .dout(n28360));
  jor  g11098(.dina(n28360), .dinb(n28359), .dout(n28361));
  jand g11099(.dina(n28361), .dinb(n28272), .dout(n28362));
  jnot g11100(.din(n28195), .dout(n28363));
  jor  g11101(.dina(n28363), .dinb(n28362), .dout(n28364));
  jand g11102(.dina(n28364), .dinb(n28271), .dout(n28365));
  jnot g11103(.din(n28198), .dout(n28366));
  jor  g11104(.dina(n28366), .dinb(n28365), .dout(n28367));
  jand g11105(.dina(n28367), .dinb(n28270), .dout(n28368));
  jnot g11106(.din(n28201), .dout(n28369));
  jor  g11107(.dina(n28369), .dinb(n28368), .dout(n28370));
  jand g11108(.dina(n28370), .dinb(n28269), .dout(n28371));
  jnot g11109(.din(n28204), .dout(n28372));
  jor  g11110(.dina(n28372), .dinb(n28371), .dout(n28373));
  jand g11111(.dina(n28373), .dinb(n28268), .dout(n28374));
  jnot g11112(.din(n28207), .dout(n28375));
  jor  g11113(.dina(n28375), .dinb(n28374), .dout(n28376));
  jand g11114(.dina(n28376), .dinb(n28267), .dout(n28377));
  jnot g11115(.din(n28210), .dout(n28378));
  jor  g11116(.dina(n28378), .dinb(n28377), .dout(n28379));
  jand g11117(.dina(n28379), .dinb(n28266), .dout(n28380));
  jnot g11118(.din(n28213), .dout(n28381));
  jor  g11119(.dina(n28381), .dinb(n28380), .dout(n28382));
  jand g11120(.dina(n28382), .dinb(n28265), .dout(n28383));
  jnot g11121(.din(n28216), .dout(n28384));
  jor  g11122(.dina(n28384), .dinb(n28383), .dout(n28385));
  jand g11123(.dina(n28385), .dinb(n28264), .dout(n28386));
  jnot g11124(.din(n28219), .dout(n28387));
  jor  g11125(.dina(n28387), .dinb(n28386), .dout(n28388));
  jand g11126(.dina(n28388), .dinb(n28263), .dout(n28389));
  jnot g11127(.din(n28222), .dout(n28390));
  jor  g11128(.dina(n28390), .dinb(n28389), .dout(n28391));
  jand g11129(.dina(n28391), .dinb(n28262), .dout(n28392));
  jnot g11130(.din(n28225), .dout(n28393));
  jor  g11131(.dina(n28393), .dinb(n28392), .dout(n28394));
  jand g11132(.dina(n28394), .dinb(n28261), .dout(n28395));
  jnot g11133(.din(n28228), .dout(n28396));
  jor  g11134(.dina(n28396), .dinb(n28395), .dout(n28397));
  jand g11135(.dina(n28397), .dinb(n28260), .dout(n28398));
  jnot g11136(.din(n28231), .dout(n28399));
  jor  g11137(.dina(n28399), .dinb(n28398), .dout(n28400));
  jand g11138(.dina(n28400), .dinb(n28259), .dout(n28401));
  jnot g11139(.din(n28234), .dout(n28402));
  jor  g11140(.dina(n28402), .dinb(n28401), .dout(n28403));
  jand g11141(.dina(n28403), .dinb(n28258), .dout(n28404));
  jnot g11142(.din(n28237), .dout(n28405));
  jor  g11143(.dina(n28405), .dinb(n28404), .dout(n28406));
  jand g11144(.dina(n28406), .dinb(n28257), .dout(n28407));
  jnot g11145(.din(n28240), .dout(n28408));
  jor  g11146(.dina(n28408), .dinb(n28407), .dout(n28409));
  jand g11147(.dina(n28409), .dinb(n28256), .dout(n28410));
  jnot g11148(.din(n28243), .dout(n28411));
  jor  g11149(.dina(n28411), .dinb(n28410), .dout(n28412));
  jand g11150(.dina(n28412), .dinb(n28255), .dout(n28413));
  jnot g11151(.din(n28246), .dout(n28414));
  jor  g11152(.dina(n28414), .dinb(n28413), .dout(n28415));
  jand g11153(.dina(n28415), .dinb(n28254), .dout(n28416));
  jor  g11154(.dina(n28416), .dinb(n27921), .dout(n28417));
  jand g11155(.dina(n28417), .dinb(n28253), .dout(n28418));
  jor  g11156(.dina(n28418), .dinb(n848), .dout(n28419));
  jxor g11157(.dina(n28246), .dinb(n28245), .dout(n28420));
  jor  g11158(.dina(n28420), .dinb(n28419), .dout(n28421));
  jand g11159(.dina(n28421), .dinb(n28252), .dout(n28422));
  jand g11160(.dina(n28419), .dinb(n27918), .dout(n28423));
  jand g11161(.dina(n28248), .dinb(n27919), .dout(n28424));
  jor  g11162(.dina(n28424), .dinb(n28423), .dout(n28425));
  jand g11163(.dina(n28425), .dinb(n405), .dout(n28426));
  jand g11164(.dina(n28422), .dinb(n280), .dout(n28427));
  jor  g11165(.dina(n28251), .dinb(n27927), .dout(n28428));
  jxor g11166(.dina(n28243), .dinb(n28242), .dout(n28429));
  jor  g11167(.dina(n28429), .dinb(n28419), .dout(n28430));
  jand g11168(.dina(n28430), .dinb(n28428), .dout(n28431));
  jand g11169(.dina(n28431), .dinb(n279), .dout(n28432));
  jor  g11170(.dina(n28251), .dinb(n27932), .dout(n28433));
  jxor g11171(.dina(n28240), .dinb(n28239), .dout(n28434));
  jor  g11172(.dina(n28434), .dinb(n28419), .dout(n28435));
  jand g11173(.dina(n28435), .dinb(n28433), .dout(n28436));
  jand g11174(.dina(n28436), .dinb(n278), .dout(n28437));
  jor  g11175(.dina(n28251), .dinb(n27937), .dout(n28438));
  jxor g11176(.dina(n28237), .dinb(n28236), .dout(n28439));
  jor  g11177(.dina(n28439), .dinb(n28419), .dout(n28440));
  jand g11178(.dina(n28440), .dinb(n28438), .dout(n28441));
  jand g11179(.dina(n28441), .dinb(n277), .dout(n28442));
  jor  g11180(.dina(n28251), .dinb(n27942), .dout(n28443));
  jxor g11181(.dina(n28234), .dinb(n28233), .dout(n28444));
  jor  g11182(.dina(n28444), .dinb(n28419), .dout(n28445));
  jand g11183(.dina(n28445), .dinb(n28443), .dout(n28446));
  jand g11184(.dina(n28446), .dinb(n326), .dout(n28447));
  jor  g11185(.dina(n28251), .dinb(n27947), .dout(n28448));
  jxor g11186(.dina(n28231), .dinb(n28230), .dout(n28449));
  jor  g11187(.dina(n28449), .dinb(n28419), .dout(n28450));
  jand g11188(.dina(n28450), .dinb(n28448), .dout(n28451));
  jand g11189(.dina(n28451), .dinb(n325), .dout(n28452));
  jor  g11190(.dina(n28251), .dinb(n27952), .dout(n28453));
  jxor g11191(.dina(n28228), .dinb(n28227), .dout(n28454));
  jor  g11192(.dina(n28454), .dinb(n28419), .dout(n28455));
  jand g11193(.dina(n28455), .dinb(n28453), .dout(n28456));
  jand g11194(.dina(n28456), .dinb(n324), .dout(n28457));
  jor  g11195(.dina(n28251), .dinb(n27957), .dout(n28458));
  jxor g11196(.dina(n28225), .dinb(n28224), .dout(n28459));
  jor  g11197(.dina(n28459), .dinb(n28419), .dout(n28460));
  jand g11198(.dina(n28460), .dinb(n28458), .dout(n28461));
  jand g11199(.dina(n28461), .dinb(n276), .dout(n28462));
  jor  g11200(.dina(n28251), .dinb(n27962), .dout(n28463));
  jxor g11201(.dina(n28222), .dinb(n28221), .dout(n28464));
  jor  g11202(.dina(n28464), .dinb(n28419), .dout(n28465));
  jand g11203(.dina(n28465), .dinb(n28463), .dout(n28466));
  jand g11204(.dina(n28466), .dinb(n333), .dout(n28467));
  jor  g11205(.dina(n28251), .dinb(n27967), .dout(n28468));
  jxor g11206(.dina(n28219), .dinb(n28218), .dout(n28469));
  jor  g11207(.dina(n28469), .dinb(n28419), .dout(n28470));
  jand g11208(.dina(n28470), .dinb(n28468), .dout(n28471));
  jand g11209(.dina(n28471), .dinb(n332), .dout(n28472));
  jor  g11210(.dina(n28251), .dinb(n27972), .dout(n28473));
  jxor g11211(.dina(n28216), .dinb(n28215), .dout(n28474));
  jor  g11212(.dina(n28474), .dinb(n28419), .dout(n28475));
  jand g11213(.dina(n28475), .dinb(n28473), .dout(n28476));
  jand g11214(.dina(n28476), .dinb(n331), .dout(n28477));
  jor  g11215(.dina(n28251), .dinb(n27977), .dout(n28478));
  jxor g11216(.dina(n28213), .dinb(n28212), .dout(n28479));
  jor  g11217(.dina(n28479), .dinb(n28419), .dout(n28480));
  jand g11218(.dina(n28480), .dinb(n28478), .dout(n28481));
  jand g11219(.dina(n28481), .dinb(n275), .dout(n28482));
  jor  g11220(.dina(n28251), .dinb(n27982), .dout(n28483));
  jxor g11221(.dina(n28210), .dinb(n28209), .dout(n28484));
  jor  g11222(.dina(n28484), .dinb(n28419), .dout(n28485));
  jand g11223(.dina(n28485), .dinb(n28483), .dout(n28486));
  jand g11224(.dina(n28486), .dinb(n340), .dout(n28487));
  jor  g11225(.dina(n28251), .dinb(n27987), .dout(n28488));
  jxor g11226(.dina(n28207), .dinb(n28206), .dout(n28489));
  jor  g11227(.dina(n28489), .dinb(n28419), .dout(n28490));
  jand g11228(.dina(n28490), .dinb(n28488), .dout(n28491));
  jand g11229(.dina(n28491), .dinb(n339), .dout(n28492));
  jor  g11230(.dina(n28251), .dinb(n27992), .dout(n28493));
  jxor g11231(.dina(n28204), .dinb(n28203), .dout(n28494));
  jor  g11232(.dina(n28494), .dinb(n28419), .dout(n28495));
  jand g11233(.dina(n28495), .dinb(n28493), .dout(n28496));
  jand g11234(.dina(n28496), .dinb(n338), .dout(n28497));
  jor  g11235(.dina(n28251), .dinb(n27997), .dout(n28498));
  jxor g11236(.dina(n28201), .dinb(n28200), .dout(n28499));
  jor  g11237(.dina(n28499), .dinb(n28419), .dout(n28500));
  jand g11238(.dina(n28500), .dinb(n28498), .dout(n28501));
  jand g11239(.dina(n28501), .dinb(n271), .dout(n28502));
  jor  g11240(.dina(n28251), .dinb(n28002), .dout(n28503));
  jxor g11241(.dina(n28198), .dinb(n28197), .dout(n28504));
  jor  g11242(.dina(n28504), .dinb(n28419), .dout(n28505));
  jand g11243(.dina(n28505), .dinb(n28503), .dout(n28506));
  jand g11244(.dina(n28506), .dinb(n270), .dout(n28507));
  jor  g11245(.dina(n28251), .dinb(n28007), .dout(n28508));
  jxor g11246(.dina(n28195), .dinb(n28194), .dout(n28509));
  jor  g11247(.dina(n28509), .dinb(n28419), .dout(n28510));
  jand g11248(.dina(n28510), .dinb(n28508), .dout(n28511));
  jand g11249(.dina(n28511), .dinb(n269), .dout(n28512));
  jor  g11250(.dina(n28251), .dinb(n28012), .dout(n28513));
  jxor g11251(.dina(n28192), .dinb(n28191), .dout(n28514));
  jor  g11252(.dina(n28514), .dinb(n28419), .dout(n28515));
  jand g11253(.dina(n28515), .dinb(n28513), .dout(n28516));
  jand g11254(.dina(n28516), .dinb(n274), .dout(n28517));
  jor  g11255(.dina(n28251), .dinb(n28017), .dout(n28518));
  jxor g11256(.dina(n28189), .dinb(n28188), .dout(n28519));
  jor  g11257(.dina(n28519), .dinb(n28419), .dout(n28520));
  jand g11258(.dina(n28520), .dinb(n28518), .dout(n28521));
  jand g11259(.dina(n28521), .dinb(n268), .dout(n28522));
  jor  g11260(.dina(n28251), .dinb(n28022), .dout(n28523));
  jxor g11261(.dina(n28186), .dinb(n28185), .dout(n28524));
  jor  g11262(.dina(n28524), .dinb(n28419), .dout(n28525));
  jand g11263(.dina(n28525), .dinb(n28523), .dout(n28526));
  jand g11264(.dina(n28526), .dinb(n349), .dout(n28527));
  jor  g11265(.dina(n28251), .dinb(n28027), .dout(n28528));
  jxor g11266(.dina(n28183), .dinb(n28182), .dout(n28529));
  jor  g11267(.dina(n28529), .dinb(n28419), .dout(n28530));
  jand g11268(.dina(n28530), .dinb(n28528), .dout(n28531));
  jand g11269(.dina(n28531), .dinb(n348), .dout(n28532));
  jor  g11270(.dina(n28251), .dinb(n28032), .dout(n28533));
  jxor g11271(.dina(n28180), .dinb(n28179), .dout(n28534));
  jor  g11272(.dina(n28534), .dinb(n28419), .dout(n28535));
  jand g11273(.dina(n28535), .dinb(n28533), .dout(n28536));
  jand g11274(.dina(n28536), .dinb(n347), .dout(n28537));
  jor  g11275(.dina(n28251), .dinb(n28037), .dout(n28538));
  jxor g11276(.dina(n28177), .dinb(n28176), .dout(n28539));
  jor  g11277(.dina(n28539), .dinb(n28419), .dout(n28540));
  jand g11278(.dina(n28540), .dinb(n28538), .dout(n28541));
  jand g11279(.dina(n28541), .dinb(n267), .dout(n28542));
  jor  g11280(.dina(n28251), .dinb(n28042), .dout(n28543));
  jxor g11281(.dina(n28174), .dinb(n28173), .dout(n28544));
  jor  g11282(.dina(n28544), .dinb(n28419), .dout(n28545));
  jand g11283(.dina(n28545), .dinb(n28543), .dout(n28546));
  jand g11284(.dina(n28546), .dinb(n266), .dout(n28547));
  jor  g11285(.dina(n28251), .dinb(n28047), .dout(n28548));
  jxor g11286(.dina(n28171), .dinb(n28170), .dout(n28549));
  jor  g11287(.dina(n28549), .dinb(n28419), .dout(n28550));
  jand g11288(.dina(n28550), .dinb(n28548), .dout(n28551));
  jand g11289(.dina(n28551), .dinb(n356), .dout(n28552));
  jor  g11290(.dina(n28251), .dinb(n28052), .dout(n28553));
  jxor g11291(.dina(n28168), .dinb(n28167), .dout(n28554));
  jor  g11292(.dina(n28554), .dinb(n28419), .dout(n28555));
  jand g11293(.dina(n28555), .dinb(n28553), .dout(n28556));
  jand g11294(.dina(n28556), .dinb(n355), .dout(n28557));
  jor  g11295(.dina(n28251), .dinb(n28057), .dout(n28558));
  jxor g11296(.dina(n28165), .dinb(n28164), .dout(n28559));
  jor  g11297(.dina(n28559), .dinb(n28419), .dout(n28560));
  jand g11298(.dina(n28560), .dinb(n28558), .dout(n28561));
  jand g11299(.dina(n28561), .dinb(n364), .dout(n28562));
  jor  g11300(.dina(n28251), .dinb(n28062), .dout(n28563));
  jxor g11301(.dina(n28162), .dinb(n28161), .dout(n28564));
  jor  g11302(.dina(n28564), .dinb(n28419), .dout(n28565));
  jand g11303(.dina(n28565), .dinb(n28563), .dout(n28566));
  jand g11304(.dina(n28566), .dinb(n361), .dout(n28567));
  jor  g11305(.dina(n28251), .dinb(n28067), .dout(n28568));
  jxor g11306(.dina(n28159), .dinb(n28158), .dout(n28569));
  jor  g11307(.dina(n28569), .dinb(n28419), .dout(n28570));
  jand g11308(.dina(n28570), .dinb(n28568), .dout(n28571));
  jand g11309(.dina(n28571), .dinb(n360), .dout(n28572));
  jor  g11310(.dina(n28251), .dinb(n28072), .dout(n28573));
  jxor g11311(.dina(n28156), .dinb(n28155), .dout(n28574));
  jor  g11312(.dina(n28574), .dinb(n28419), .dout(n28575));
  jand g11313(.dina(n28575), .dinb(n28573), .dout(n28576));
  jand g11314(.dina(n28576), .dinb(n363), .dout(n28577));
  jor  g11315(.dina(n28251), .dinb(n28077), .dout(n28578));
  jxor g11316(.dina(n28153), .dinb(n28152), .dout(n28579));
  jor  g11317(.dina(n28579), .dinb(n28419), .dout(n28580));
  jand g11318(.dina(n28580), .dinb(n28578), .dout(n28581));
  jand g11319(.dina(n28581), .dinb(n359), .dout(n28582));
  jor  g11320(.dina(n28251), .dinb(n28082), .dout(n28583));
  jxor g11321(.dina(n28150), .dinb(n28149), .dout(n28584));
  jor  g11322(.dina(n28584), .dinb(n28419), .dout(n28585));
  jand g11323(.dina(n28585), .dinb(n28583), .dout(n28586));
  jand g11324(.dina(n28586), .dinb(n369), .dout(n28587));
  jor  g11325(.dina(n28251), .dinb(n28087), .dout(n28588));
  jxor g11326(.dina(n28147), .dinb(n28146), .dout(n28589));
  jor  g11327(.dina(n28589), .dinb(n28419), .dout(n28590));
  jand g11328(.dina(n28590), .dinb(n28588), .dout(n28591));
  jand g11329(.dina(n28591), .dinb(n368), .dout(n28592));
  jor  g11330(.dina(n28251), .dinb(n28092), .dout(n28593));
  jxor g11331(.dina(n28144), .dinb(n28143), .dout(n28594));
  jor  g11332(.dina(n28594), .dinb(n28419), .dout(n28595));
  jand g11333(.dina(n28595), .dinb(n28593), .dout(n28596));
  jand g11334(.dina(n28596), .dinb(n367), .dout(n28597));
  jor  g11335(.dina(n28251), .dinb(n28097), .dout(n28598));
  jxor g11336(.dina(n28141), .dinb(n28140), .dout(n28599));
  jor  g11337(.dina(n28599), .dinb(n28419), .dout(n28600));
  jand g11338(.dina(n28600), .dinb(n28598), .dout(n28601));
  jand g11339(.dina(n28601), .dinb(n265), .dout(n28602));
  jor  g11340(.dina(n28251), .dinb(n28102), .dout(n28603));
  jxor g11341(.dina(n28138), .dinb(n28137), .dout(n28604));
  jor  g11342(.dina(n28604), .dinb(n28419), .dout(n28605));
  jand g11343(.dina(n28605), .dinb(n28603), .dout(n28606));
  jand g11344(.dina(n28606), .dinb(n378), .dout(n28607));
  jor  g11345(.dina(n28251), .dinb(n28107), .dout(n28608));
  jxor g11346(.dina(n28135), .dinb(n28134), .dout(n28609));
  jor  g11347(.dina(n28609), .dinb(n28419), .dout(n28610));
  jand g11348(.dina(n28610), .dinb(n28608), .dout(n28611));
  jand g11349(.dina(n28611), .dinb(n377), .dout(n28612));
  jor  g11350(.dina(n28251), .dinb(n28112), .dout(n28613));
  jxor g11351(.dina(n28132), .dinb(n28131), .dout(n28614));
  jor  g11352(.dina(n28614), .dinb(n28419), .dout(n28615));
  jand g11353(.dina(n28615), .dinb(n28613), .dout(n28616));
  jand g11354(.dina(n28616), .dinb(n376), .dout(n28617));
  jnot g11355(.din(n28119), .dout(n28618));
  jor  g11356(.dina(n28251), .dinb(n28618), .dout(n28619));
  jxor g11357(.dina(n28129), .dinb(n28128), .dout(n28620));
  jor  g11358(.dina(n28620), .dinb(n28419), .dout(n28621));
  jand g11359(.dina(n28621), .dinb(n28619), .dout(n28622));
  jand g11360(.dina(n28622), .dinb(n264), .dout(n28623));
  jand g11361(.dina(n28419), .dinb(n28123), .dout(n28624));
  jxor g11362(.dina(n28126), .dinb(n8617), .dout(n28625));
  jand g11363(.dina(n28625), .dinb(n28251), .dout(n28626));
  jor  g11364(.dina(n28626), .dinb(n28624), .dout(n28627));
  jand g11365(.dina(n28627), .dinb(n386), .dout(n28628));
  jnot g11366(.din(n7074), .dout(n28629));
  jor  g11367(.dina(n28418), .dinb(n28629), .dout(n28630));
  jand g11368(.dina(n28630), .dinb(a21 ), .dout(n28631));
  jand g11369(.dina(n28251), .dinb(n8447), .dout(n28632));
  jor  g11370(.dina(n28632), .dinb(n28631), .dout(n28633));
  jand g11371(.dina(n28633), .dinb(n259), .dout(n28634));
  jand g11372(.dina(n28250), .dinb(n7074), .dout(n28635));
  jor  g11373(.dina(n28635), .dinb(n8446), .dout(n28636));
  jor  g11374(.dina(n28419), .dinb(n8617), .dout(n28637));
  jand g11375(.dina(n28637), .dinb(n28636), .dout(n28638));
  jxor g11376(.dina(n28638), .dinb(b1 ), .dout(n28639));
  jand g11377(.dina(n28639), .dinb(n8925), .dout(n28640));
  jor  g11378(.dina(n28640), .dinb(n28634), .dout(n28641));
  jxor g11379(.dina(n28627), .dinb(n386), .dout(n28642));
  jand g11380(.dina(n28642), .dinb(n28641), .dout(n28643));
  jor  g11381(.dina(n28643), .dinb(n28628), .dout(n28644));
  jxor g11382(.dina(n28622), .dinb(n264), .dout(n28645));
  jand g11383(.dina(n28645), .dinb(n28644), .dout(n28646));
  jor  g11384(.dina(n28646), .dinb(n28623), .dout(n28647));
  jxor g11385(.dina(n28616), .dinb(n376), .dout(n28648));
  jand g11386(.dina(n28648), .dinb(n28647), .dout(n28649));
  jor  g11387(.dina(n28649), .dinb(n28617), .dout(n28650));
  jxor g11388(.dina(n28611), .dinb(n377), .dout(n28651));
  jand g11389(.dina(n28651), .dinb(n28650), .dout(n28652));
  jor  g11390(.dina(n28652), .dinb(n28612), .dout(n28653));
  jxor g11391(.dina(n28606), .dinb(n378), .dout(n28654));
  jand g11392(.dina(n28654), .dinb(n28653), .dout(n28655));
  jor  g11393(.dina(n28655), .dinb(n28607), .dout(n28656));
  jxor g11394(.dina(n28601), .dinb(n265), .dout(n28657));
  jand g11395(.dina(n28657), .dinb(n28656), .dout(n28658));
  jor  g11396(.dina(n28658), .dinb(n28602), .dout(n28659));
  jxor g11397(.dina(n28596), .dinb(n367), .dout(n28660));
  jand g11398(.dina(n28660), .dinb(n28659), .dout(n28661));
  jor  g11399(.dina(n28661), .dinb(n28597), .dout(n28662));
  jxor g11400(.dina(n28591), .dinb(n368), .dout(n28663));
  jand g11401(.dina(n28663), .dinb(n28662), .dout(n28664));
  jor  g11402(.dina(n28664), .dinb(n28592), .dout(n28665));
  jxor g11403(.dina(n28586), .dinb(n369), .dout(n28666));
  jand g11404(.dina(n28666), .dinb(n28665), .dout(n28667));
  jor  g11405(.dina(n28667), .dinb(n28587), .dout(n28668));
  jxor g11406(.dina(n28581), .dinb(n359), .dout(n28669));
  jand g11407(.dina(n28669), .dinb(n28668), .dout(n28670));
  jor  g11408(.dina(n28670), .dinb(n28582), .dout(n28671));
  jxor g11409(.dina(n28576), .dinb(n363), .dout(n28672));
  jand g11410(.dina(n28672), .dinb(n28671), .dout(n28673));
  jor  g11411(.dina(n28673), .dinb(n28577), .dout(n28674));
  jxor g11412(.dina(n28571), .dinb(n360), .dout(n28675));
  jand g11413(.dina(n28675), .dinb(n28674), .dout(n28676));
  jor  g11414(.dina(n28676), .dinb(n28572), .dout(n28677));
  jxor g11415(.dina(n28566), .dinb(n361), .dout(n28678));
  jand g11416(.dina(n28678), .dinb(n28677), .dout(n28679));
  jor  g11417(.dina(n28679), .dinb(n28567), .dout(n28680));
  jxor g11418(.dina(n28561), .dinb(n364), .dout(n28681));
  jand g11419(.dina(n28681), .dinb(n28680), .dout(n28682));
  jor  g11420(.dina(n28682), .dinb(n28562), .dout(n28683));
  jxor g11421(.dina(n28556), .dinb(n355), .dout(n28684));
  jand g11422(.dina(n28684), .dinb(n28683), .dout(n28685));
  jor  g11423(.dina(n28685), .dinb(n28557), .dout(n28686));
  jxor g11424(.dina(n28551), .dinb(n356), .dout(n28687));
  jand g11425(.dina(n28687), .dinb(n28686), .dout(n28688));
  jor  g11426(.dina(n28688), .dinb(n28552), .dout(n28689));
  jxor g11427(.dina(n28546), .dinb(n266), .dout(n28690));
  jand g11428(.dina(n28690), .dinb(n28689), .dout(n28691));
  jor  g11429(.dina(n28691), .dinb(n28547), .dout(n28692));
  jxor g11430(.dina(n28541), .dinb(n267), .dout(n28693));
  jand g11431(.dina(n28693), .dinb(n28692), .dout(n28694));
  jor  g11432(.dina(n28694), .dinb(n28542), .dout(n28695));
  jxor g11433(.dina(n28536), .dinb(n347), .dout(n28696));
  jand g11434(.dina(n28696), .dinb(n28695), .dout(n28697));
  jor  g11435(.dina(n28697), .dinb(n28537), .dout(n28698));
  jxor g11436(.dina(n28531), .dinb(n348), .dout(n28699));
  jand g11437(.dina(n28699), .dinb(n28698), .dout(n28700));
  jor  g11438(.dina(n28700), .dinb(n28532), .dout(n28701));
  jxor g11439(.dina(n28526), .dinb(n349), .dout(n28702));
  jand g11440(.dina(n28702), .dinb(n28701), .dout(n28703));
  jor  g11441(.dina(n28703), .dinb(n28527), .dout(n28704));
  jxor g11442(.dina(n28521), .dinb(n268), .dout(n28705));
  jand g11443(.dina(n28705), .dinb(n28704), .dout(n28706));
  jor  g11444(.dina(n28706), .dinb(n28522), .dout(n28707));
  jxor g11445(.dina(n28516), .dinb(n274), .dout(n28708));
  jand g11446(.dina(n28708), .dinb(n28707), .dout(n28709));
  jor  g11447(.dina(n28709), .dinb(n28517), .dout(n28710));
  jxor g11448(.dina(n28511), .dinb(n269), .dout(n28711));
  jand g11449(.dina(n28711), .dinb(n28710), .dout(n28712));
  jor  g11450(.dina(n28712), .dinb(n28512), .dout(n28713));
  jxor g11451(.dina(n28506), .dinb(n270), .dout(n28714));
  jand g11452(.dina(n28714), .dinb(n28713), .dout(n28715));
  jor  g11453(.dina(n28715), .dinb(n28507), .dout(n28716));
  jxor g11454(.dina(n28501), .dinb(n271), .dout(n28717));
  jand g11455(.dina(n28717), .dinb(n28716), .dout(n28718));
  jor  g11456(.dina(n28718), .dinb(n28502), .dout(n28719));
  jxor g11457(.dina(n28496), .dinb(n338), .dout(n28720));
  jand g11458(.dina(n28720), .dinb(n28719), .dout(n28721));
  jor  g11459(.dina(n28721), .dinb(n28497), .dout(n28722));
  jxor g11460(.dina(n28491), .dinb(n339), .dout(n28723));
  jand g11461(.dina(n28723), .dinb(n28722), .dout(n28724));
  jor  g11462(.dina(n28724), .dinb(n28492), .dout(n28725));
  jxor g11463(.dina(n28486), .dinb(n340), .dout(n28726));
  jand g11464(.dina(n28726), .dinb(n28725), .dout(n28727));
  jor  g11465(.dina(n28727), .dinb(n28487), .dout(n28728));
  jxor g11466(.dina(n28481), .dinb(n275), .dout(n28729));
  jand g11467(.dina(n28729), .dinb(n28728), .dout(n28730));
  jor  g11468(.dina(n28730), .dinb(n28482), .dout(n28731));
  jxor g11469(.dina(n28476), .dinb(n331), .dout(n28732));
  jand g11470(.dina(n28732), .dinb(n28731), .dout(n28733));
  jor  g11471(.dina(n28733), .dinb(n28477), .dout(n28734));
  jxor g11472(.dina(n28471), .dinb(n332), .dout(n28735));
  jand g11473(.dina(n28735), .dinb(n28734), .dout(n28736));
  jor  g11474(.dina(n28736), .dinb(n28472), .dout(n28737));
  jxor g11475(.dina(n28466), .dinb(n333), .dout(n28738));
  jand g11476(.dina(n28738), .dinb(n28737), .dout(n28739));
  jor  g11477(.dina(n28739), .dinb(n28467), .dout(n28740));
  jxor g11478(.dina(n28461), .dinb(n276), .dout(n28741));
  jand g11479(.dina(n28741), .dinb(n28740), .dout(n28742));
  jor  g11480(.dina(n28742), .dinb(n28462), .dout(n28743));
  jxor g11481(.dina(n28456), .dinb(n324), .dout(n28744));
  jand g11482(.dina(n28744), .dinb(n28743), .dout(n28745));
  jor  g11483(.dina(n28745), .dinb(n28457), .dout(n28746));
  jxor g11484(.dina(n28451), .dinb(n325), .dout(n28747));
  jand g11485(.dina(n28747), .dinb(n28746), .dout(n28748));
  jor  g11486(.dina(n28748), .dinb(n28452), .dout(n28749));
  jxor g11487(.dina(n28446), .dinb(n326), .dout(n28750));
  jand g11488(.dina(n28750), .dinb(n28749), .dout(n28751));
  jor  g11489(.dina(n28751), .dinb(n28447), .dout(n28752));
  jxor g11490(.dina(n28441), .dinb(n277), .dout(n28753));
  jand g11491(.dina(n28753), .dinb(n28752), .dout(n28754));
  jor  g11492(.dina(n28754), .dinb(n28442), .dout(n28755));
  jxor g11493(.dina(n28436), .dinb(n278), .dout(n28756));
  jand g11494(.dina(n28756), .dinb(n28755), .dout(n28757));
  jor  g11495(.dina(n28757), .dinb(n28437), .dout(n28758));
  jxor g11496(.dina(n28431), .dinb(n279), .dout(n28759));
  jand g11497(.dina(n28759), .dinb(n28758), .dout(n28760));
  jor  g11498(.dina(n28760), .dinb(n28432), .dout(n28761));
  jxor g11499(.dina(n28422), .dinb(n280), .dout(n28762));
  jand g11500(.dina(n28762), .dinb(n28761), .dout(n28763));
  jor  g11501(.dina(n28763), .dinb(n28427), .dout(n28764));
  jxor g11502(.dina(n28425), .dinb(b43 ), .dout(n28765));
  jnot g11503(.din(n28765), .dout(n28766));
  jand g11504(.dina(n28766), .dinb(n28764), .dout(n28767));
  jand g11505(.dina(n28767), .dinb(n320), .dout(n28768));
  jor  g11506(.dina(n28768), .dinb(n28426), .dout(n28769));
  jor  g11507(.dina(n28769), .dinb(n28422), .dout(n28770));
  jnot g11508(.din(n28769), .dout(n28771));
  jxor g11509(.dina(n28762), .dinb(n28761), .dout(n28772));
  jor  g11510(.dina(n28772), .dinb(n28771), .dout(n28773));
  jand g11511(.dina(n28773), .dinb(n28770), .dout(n28774));
  jand g11512(.dina(n28774), .dinb(n283), .dout(n28775));
  jor  g11513(.dina(n28769), .dinb(n28431), .dout(n28776));
  jxor g11514(.dina(n28759), .dinb(n28758), .dout(n28777));
  jor  g11515(.dina(n28777), .dinb(n28771), .dout(n28778));
  jand g11516(.dina(n28778), .dinb(n28776), .dout(n28779));
  jand g11517(.dina(n28779), .dinb(n280), .dout(n28780));
  jor  g11518(.dina(n28769), .dinb(n28436), .dout(n28781));
  jxor g11519(.dina(n28756), .dinb(n28755), .dout(n28782));
  jor  g11520(.dina(n28782), .dinb(n28771), .dout(n28783));
  jand g11521(.dina(n28783), .dinb(n28781), .dout(n28784));
  jand g11522(.dina(n28784), .dinb(n279), .dout(n28785));
  jor  g11523(.dina(n28769), .dinb(n28441), .dout(n28786));
  jxor g11524(.dina(n28753), .dinb(n28752), .dout(n28787));
  jor  g11525(.dina(n28787), .dinb(n28771), .dout(n28788));
  jand g11526(.dina(n28788), .dinb(n28786), .dout(n28789));
  jand g11527(.dina(n28789), .dinb(n278), .dout(n28790));
  jor  g11528(.dina(n28769), .dinb(n28446), .dout(n28791));
  jxor g11529(.dina(n28750), .dinb(n28749), .dout(n28792));
  jor  g11530(.dina(n28792), .dinb(n28771), .dout(n28793));
  jand g11531(.dina(n28793), .dinb(n28791), .dout(n28794));
  jand g11532(.dina(n28794), .dinb(n277), .dout(n28795));
  jor  g11533(.dina(n28769), .dinb(n28451), .dout(n28796));
  jxor g11534(.dina(n28747), .dinb(n28746), .dout(n28797));
  jor  g11535(.dina(n28797), .dinb(n28771), .dout(n28798));
  jand g11536(.dina(n28798), .dinb(n28796), .dout(n28799));
  jand g11537(.dina(n28799), .dinb(n326), .dout(n28800));
  jor  g11538(.dina(n28769), .dinb(n28456), .dout(n28801));
  jxor g11539(.dina(n28744), .dinb(n28743), .dout(n28802));
  jor  g11540(.dina(n28802), .dinb(n28771), .dout(n28803));
  jand g11541(.dina(n28803), .dinb(n28801), .dout(n28804));
  jand g11542(.dina(n28804), .dinb(n325), .dout(n28805));
  jor  g11543(.dina(n28769), .dinb(n28461), .dout(n28806));
  jxor g11544(.dina(n28741), .dinb(n28740), .dout(n28807));
  jor  g11545(.dina(n28807), .dinb(n28771), .dout(n28808));
  jand g11546(.dina(n28808), .dinb(n28806), .dout(n28809));
  jand g11547(.dina(n28809), .dinb(n324), .dout(n28810));
  jor  g11548(.dina(n28769), .dinb(n28466), .dout(n28811));
  jxor g11549(.dina(n28738), .dinb(n28737), .dout(n28812));
  jor  g11550(.dina(n28812), .dinb(n28771), .dout(n28813));
  jand g11551(.dina(n28813), .dinb(n28811), .dout(n28814));
  jand g11552(.dina(n28814), .dinb(n276), .dout(n28815));
  jor  g11553(.dina(n28769), .dinb(n28471), .dout(n28816));
  jxor g11554(.dina(n28735), .dinb(n28734), .dout(n28817));
  jor  g11555(.dina(n28817), .dinb(n28771), .dout(n28818));
  jand g11556(.dina(n28818), .dinb(n28816), .dout(n28819));
  jand g11557(.dina(n28819), .dinb(n333), .dout(n28820));
  jor  g11558(.dina(n28769), .dinb(n28476), .dout(n28821));
  jxor g11559(.dina(n28732), .dinb(n28731), .dout(n28822));
  jor  g11560(.dina(n28822), .dinb(n28771), .dout(n28823));
  jand g11561(.dina(n28823), .dinb(n28821), .dout(n28824));
  jand g11562(.dina(n28824), .dinb(n332), .dout(n28825));
  jor  g11563(.dina(n28769), .dinb(n28481), .dout(n28826));
  jxor g11564(.dina(n28729), .dinb(n28728), .dout(n28827));
  jor  g11565(.dina(n28827), .dinb(n28771), .dout(n28828));
  jand g11566(.dina(n28828), .dinb(n28826), .dout(n28829));
  jand g11567(.dina(n28829), .dinb(n331), .dout(n28830));
  jor  g11568(.dina(n28769), .dinb(n28486), .dout(n28831));
  jxor g11569(.dina(n28726), .dinb(n28725), .dout(n28832));
  jor  g11570(.dina(n28832), .dinb(n28771), .dout(n28833));
  jand g11571(.dina(n28833), .dinb(n28831), .dout(n28834));
  jand g11572(.dina(n28834), .dinb(n275), .dout(n28835));
  jor  g11573(.dina(n28769), .dinb(n28491), .dout(n28836));
  jxor g11574(.dina(n28723), .dinb(n28722), .dout(n28837));
  jor  g11575(.dina(n28837), .dinb(n28771), .dout(n28838));
  jand g11576(.dina(n28838), .dinb(n28836), .dout(n28839));
  jand g11577(.dina(n28839), .dinb(n340), .dout(n28840));
  jor  g11578(.dina(n28769), .dinb(n28496), .dout(n28841));
  jxor g11579(.dina(n28720), .dinb(n28719), .dout(n28842));
  jor  g11580(.dina(n28842), .dinb(n28771), .dout(n28843));
  jand g11581(.dina(n28843), .dinb(n28841), .dout(n28844));
  jand g11582(.dina(n28844), .dinb(n339), .dout(n28845));
  jor  g11583(.dina(n28769), .dinb(n28501), .dout(n28846));
  jxor g11584(.dina(n28717), .dinb(n28716), .dout(n28847));
  jor  g11585(.dina(n28847), .dinb(n28771), .dout(n28848));
  jand g11586(.dina(n28848), .dinb(n28846), .dout(n28849));
  jand g11587(.dina(n28849), .dinb(n338), .dout(n28850));
  jor  g11588(.dina(n28769), .dinb(n28506), .dout(n28851));
  jxor g11589(.dina(n28714), .dinb(n28713), .dout(n28852));
  jor  g11590(.dina(n28852), .dinb(n28771), .dout(n28853));
  jand g11591(.dina(n28853), .dinb(n28851), .dout(n28854));
  jand g11592(.dina(n28854), .dinb(n271), .dout(n28855));
  jor  g11593(.dina(n28769), .dinb(n28511), .dout(n28856));
  jxor g11594(.dina(n28711), .dinb(n28710), .dout(n28857));
  jor  g11595(.dina(n28857), .dinb(n28771), .dout(n28858));
  jand g11596(.dina(n28858), .dinb(n28856), .dout(n28859));
  jand g11597(.dina(n28859), .dinb(n270), .dout(n28860));
  jor  g11598(.dina(n28769), .dinb(n28516), .dout(n28861));
  jxor g11599(.dina(n28708), .dinb(n28707), .dout(n28862));
  jor  g11600(.dina(n28862), .dinb(n28771), .dout(n28863));
  jand g11601(.dina(n28863), .dinb(n28861), .dout(n28864));
  jand g11602(.dina(n28864), .dinb(n269), .dout(n28865));
  jor  g11603(.dina(n28769), .dinb(n28521), .dout(n28866));
  jxor g11604(.dina(n28705), .dinb(n28704), .dout(n28867));
  jor  g11605(.dina(n28867), .dinb(n28771), .dout(n28868));
  jand g11606(.dina(n28868), .dinb(n28866), .dout(n28869));
  jand g11607(.dina(n28869), .dinb(n274), .dout(n28870));
  jor  g11608(.dina(n28769), .dinb(n28526), .dout(n28871));
  jxor g11609(.dina(n28702), .dinb(n28701), .dout(n28872));
  jor  g11610(.dina(n28872), .dinb(n28771), .dout(n28873));
  jand g11611(.dina(n28873), .dinb(n28871), .dout(n28874));
  jand g11612(.dina(n28874), .dinb(n268), .dout(n28875));
  jor  g11613(.dina(n28769), .dinb(n28531), .dout(n28876));
  jxor g11614(.dina(n28699), .dinb(n28698), .dout(n28877));
  jor  g11615(.dina(n28877), .dinb(n28771), .dout(n28878));
  jand g11616(.dina(n28878), .dinb(n28876), .dout(n28879));
  jand g11617(.dina(n28879), .dinb(n349), .dout(n28880));
  jor  g11618(.dina(n28769), .dinb(n28536), .dout(n28881));
  jxor g11619(.dina(n28696), .dinb(n28695), .dout(n28882));
  jor  g11620(.dina(n28882), .dinb(n28771), .dout(n28883));
  jand g11621(.dina(n28883), .dinb(n28881), .dout(n28884));
  jand g11622(.dina(n28884), .dinb(n348), .dout(n28885));
  jor  g11623(.dina(n28769), .dinb(n28541), .dout(n28886));
  jxor g11624(.dina(n28693), .dinb(n28692), .dout(n28887));
  jor  g11625(.dina(n28887), .dinb(n28771), .dout(n28888));
  jand g11626(.dina(n28888), .dinb(n28886), .dout(n28889));
  jand g11627(.dina(n28889), .dinb(n347), .dout(n28890));
  jor  g11628(.dina(n28769), .dinb(n28546), .dout(n28891));
  jxor g11629(.dina(n28690), .dinb(n28689), .dout(n28892));
  jor  g11630(.dina(n28892), .dinb(n28771), .dout(n28893));
  jand g11631(.dina(n28893), .dinb(n28891), .dout(n28894));
  jand g11632(.dina(n28894), .dinb(n267), .dout(n28895));
  jor  g11633(.dina(n28769), .dinb(n28551), .dout(n28896));
  jxor g11634(.dina(n28687), .dinb(n28686), .dout(n28897));
  jor  g11635(.dina(n28897), .dinb(n28771), .dout(n28898));
  jand g11636(.dina(n28898), .dinb(n28896), .dout(n28899));
  jand g11637(.dina(n28899), .dinb(n266), .dout(n28900));
  jor  g11638(.dina(n28769), .dinb(n28556), .dout(n28901));
  jxor g11639(.dina(n28684), .dinb(n28683), .dout(n28902));
  jor  g11640(.dina(n28902), .dinb(n28771), .dout(n28903));
  jand g11641(.dina(n28903), .dinb(n28901), .dout(n28904));
  jand g11642(.dina(n28904), .dinb(n356), .dout(n28905));
  jor  g11643(.dina(n28769), .dinb(n28561), .dout(n28906));
  jxor g11644(.dina(n28681), .dinb(n28680), .dout(n28907));
  jor  g11645(.dina(n28907), .dinb(n28771), .dout(n28908));
  jand g11646(.dina(n28908), .dinb(n28906), .dout(n28909));
  jand g11647(.dina(n28909), .dinb(n355), .dout(n28910));
  jor  g11648(.dina(n28769), .dinb(n28566), .dout(n28911));
  jxor g11649(.dina(n28678), .dinb(n28677), .dout(n28912));
  jor  g11650(.dina(n28912), .dinb(n28771), .dout(n28913));
  jand g11651(.dina(n28913), .dinb(n28911), .dout(n28914));
  jand g11652(.dina(n28914), .dinb(n364), .dout(n28915));
  jor  g11653(.dina(n28769), .dinb(n28571), .dout(n28916));
  jxor g11654(.dina(n28675), .dinb(n28674), .dout(n28917));
  jor  g11655(.dina(n28917), .dinb(n28771), .dout(n28918));
  jand g11656(.dina(n28918), .dinb(n28916), .dout(n28919));
  jand g11657(.dina(n28919), .dinb(n361), .dout(n28920));
  jor  g11658(.dina(n28769), .dinb(n28576), .dout(n28921));
  jxor g11659(.dina(n28672), .dinb(n28671), .dout(n28922));
  jor  g11660(.dina(n28922), .dinb(n28771), .dout(n28923));
  jand g11661(.dina(n28923), .dinb(n28921), .dout(n28924));
  jand g11662(.dina(n28924), .dinb(n360), .dout(n28925));
  jor  g11663(.dina(n28769), .dinb(n28581), .dout(n28926));
  jxor g11664(.dina(n28669), .dinb(n28668), .dout(n28927));
  jor  g11665(.dina(n28927), .dinb(n28771), .dout(n28928));
  jand g11666(.dina(n28928), .dinb(n28926), .dout(n28929));
  jand g11667(.dina(n28929), .dinb(n363), .dout(n28930));
  jor  g11668(.dina(n28769), .dinb(n28586), .dout(n28931));
  jxor g11669(.dina(n28666), .dinb(n28665), .dout(n28932));
  jor  g11670(.dina(n28932), .dinb(n28771), .dout(n28933));
  jand g11671(.dina(n28933), .dinb(n28931), .dout(n28934));
  jand g11672(.dina(n28934), .dinb(n359), .dout(n28935));
  jor  g11673(.dina(n28769), .dinb(n28591), .dout(n28936));
  jxor g11674(.dina(n28663), .dinb(n28662), .dout(n28937));
  jor  g11675(.dina(n28937), .dinb(n28771), .dout(n28938));
  jand g11676(.dina(n28938), .dinb(n28936), .dout(n28939));
  jand g11677(.dina(n28939), .dinb(n369), .dout(n28940));
  jor  g11678(.dina(n28769), .dinb(n28596), .dout(n28941));
  jxor g11679(.dina(n28660), .dinb(n28659), .dout(n28942));
  jor  g11680(.dina(n28942), .dinb(n28771), .dout(n28943));
  jand g11681(.dina(n28943), .dinb(n28941), .dout(n28944));
  jand g11682(.dina(n28944), .dinb(n368), .dout(n28945));
  jor  g11683(.dina(n28769), .dinb(n28601), .dout(n28946));
  jxor g11684(.dina(n28657), .dinb(n28656), .dout(n28947));
  jor  g11685(.dina(n28947), .dinb(n28771), .dout(n28948));
  jand g11686(.dina(n28948), .dinb(n28946), .dout(n28949));
  jand g11687(.dina(n28949), .dinb(n367), .dout(n28950));
  jor  g11688(.dina(n28769), .dinb(n28606), .dout(n28951));
  jxor g11689(.dina(n28654), .dinb(n28653), .dout(n28952));
  jor  g11690(.dina(n28952), .dinb(n28771), .dout(n28953));
  jand g11691(.dina(n28953), .dinb(n28951), .dout(n28954));
  jand g11692(.dina(n28954), .dinb(n265), .dout(n28955));
  jor  g11693(.dina(n28769), .dinb(n28611), .dout(n28956));
  jxor g11694(.dina(n28651), .dinb(n28650), .dout(n28957));
  jor  g11695(.dina(n28957), .dinb(n28771), .dout(n28958));
  jand g11696(.dina(n28958), .dinb(n28956), .dout(n28959));
  jand g11697(.dina(n28959), .dinb(n378), .dout(n28960));
  jor  g11698(.dina(n28769), .dinb(n28616), .dout(n28961));
  jxor g11699(.dina(n28648), .dinb(n28647), .dout(n28962));
  jor  g11700(.dina(n28962), .dinb(n28771), .dout(n28963));
  jand g11701(.dina(n28963), .dinb(n28961), .dout(n28964));
  jand g11702(.dina(n28964), .dinb(n377), .dout(n28965));
  jor  g11703(.dina(n28769), .dinb(n28622), .dout(n28966));
  jxor g11704(.dina(n28645), .dinb(n28644), .dout(n28967));
  jor  g11705(.dina(n28967), .dinb(n28771), .dout(n28968));
  jand g11706(.dina(n28968), .dinb(n28966), .dout(n28969));
  jand g11707(.dina(n28969), .dinb(n376), .dout(n28970));
  jor  g11708(.dina(n28769), .dinb(n28627), .dout(n28971));
  jxor g11709(.dina(n28642), .dinb(n28641), .dout(n28972));
  jor  g11710(.dina(n28972), .dinb(n28771), .dout(n28973));
  jand g11711(.dina(n28973), .dinb(n28971), .dout(n28974));
  jand g11712(.dina(n28974), .dinb(n264), .dout(n28975));
  jor  g11713(.dina(n28769), .dinb(n28633), .dout(n28976));
  jxor g11714(.dina(n28639), .dinb(n8925), .dout(n28977));
  jor  g11715(.dina(n28977), .dinb(n28771), .dout(n28978));
  jand g11716(.dina(n28978), .dinb(n28976), .dout(n28979));
  jand g11717(.dina(n28979), .dinb(n386), .dout(n28980));
  jand g11718(.dina(n28769), .dinb(b0 ), .dout(n28981));
  jxor g11719(.dina(n28981), .dinb(a20 ), .dout(n28982));
  jand g11720(.dina(n28982), .dinb(n259), .dout(n28983));
  jxor g11721(.dina(n28981), .dinb(n8923), .dout(n28984));
  jxor g11722(.dina(n28984), .dinb(b1 ), .dout(n28985));
  jand g11723(.dina(n28985), .dinb(n9275), .dout(n28986));
  jor  g11724(.dina(n28986), .dinb(n28983), .dout(n28987));
  jxor g11725(.dina(n28979), .dinb(n386), .dout(n28988));
  jand g11726(.dina(n28988), .dinb(n28987), .dout(n28989));
  jor  g11727(.dina(n28989), .dinb(n28980), .dout(n28990));
  jxor g11728(.dina(n28974), .dinb(n264), .dout(n28991));
  jand g11729(.dina(n28991), .dinb(n28990), .dout(n28992));
  jor  g11730(.dina(n28992), .dinb(n28975), .dout(n28993));
  jxor g11731(.dina(n28969), .dinb(n376), .dout(n28994));
  jand g11732(.dina(n28994), .dinb(n28993), .dout(n28995));
  jor  g11733(.dina(n28995), .dinb(n28970), .dout(n28996));
  jxor g11734(.dina(n28964), .dinb(n377), .dout(n28997));
  jand g11735(.dina(n28997), .dinb(n28996), .dout(n28998));
  jor  g11736(.dina(n28998), .dinb(n28965), .dout(n28999));
  jxor g11737(.dina(n28959), .dinb(n378), .dout(n29000));
  jand g11738(.dina(n29000), .dinb(n28999), .dout(n29001));
  jor  g11739(.dina(n29001), .dinb(n28960), .dout(n29002));
  jxor g11740(.dina(n28954), .dinb(n265), .dout(n29003));
  jand g11741(.dina(n29003), .dinb(n29002), .dout(n29004));
  jor  g11742(.dina(n29004), .dinb(n28955), .dout(n29005));
  jxor g11743(.dina(n28949), .dinb(n367), .dout(n29006));
  jand g11744(.dina(n29006), .dinb(n29005), .dout(n29007));
  jor  g11745(.dina(n29007), .dinb(n28950), .dout(n29008));
  jxor g11746(.dina(n28944), .dinb(n368), .dout(n29009));
  jand g11747(.dina(n29009), .dinb(n29008), .dout(n29010));
  jor  g11748(.dina(n29010), .dinb(n28945), .dout(n29011));
  jxor g11749(.dina(n28939), .dinb(n369), .dout(n29012));
  jand g11750(.dina(n29012), .dinb(n29011), .dout(n29013));
  jor  g11751(.dina(n29013), .dinb(n28940), .dout(n29014));
  jxor g11752(.dina(n28934), .dinb(n359), .dout(n29015));
  jand g11753(.dina(n29015), .dinb(n29014), .dout(n29016));
  jor  g11754(.dina(n29016), .dinb(n28935), .dout(n29017));
  jxor g11755(.dina(n28929), .dinb(n363), .dout(n29018));
  jand g11756(.dina(n29018), .dinb(n29017), .dout(n29019));
  jor  g11757(.dina(n29019), .dinb(n28930), .dout(n29020));
  jxor g11758(.dina(n28924), .dinb(n360), .dout(n29021));
  jand g11759(.dina(n29021), .dinb(n29020), .dout(n29022));
  jor  g11760(.dina(n29022), .dinb(n28925), .dout(n29023));
  jxor g11761(.dina(n28919), .dinb(n361), .dout(n29024));
  jand g11762(.dina(n29024), .dinb(n29023), .dout(n29025));
  jor  g11763(.dina(n29025), .dinb(n28920), .dout(n29026));
  jxor g11764(.dina(n28914), .dinb(n364), .dout(n29027));
  jand g11765(.dina(n29027), .dinb(n29026), .dout(n29028));
  jor  g11766(.dina(n29028), .dinb(n28915), .dout(n29029));
  jxor g11767(.dina(n28909), .dinb(n355), .dout(n29030));
  jand g11768(.dina(n29030), .dinb(n29029), .dout(n29031));
  jor  g11769(.dina(n29031), .dinb(n28910), .dout(n29032));
  jxor g11770(.dina(n28904), .dinb(n356), .dout(n29033));
  jand g11771(.dina(n29033), .dinb(n29032), .dout(n29034));
  jor  g11772(.dina(n29034), .dinb(n28905), .dout(n29035));
  jxor g11773(.dina(n28899), .dinb(n266), .dout(n29036));
  jand g11774(.dina(n29036), .dinb(n29035), .dout(n29037));
  jor  g11775(.dina(n29037), .dinb(n28900), .dout(n29038));
  jxor g11776(.dina(n28894), .dinb(n267), .dout(n29039));
  jand g11777(.dina(n29039), .dinb(n29038), .dout(n29040));
  jor  g11778(.dina(n29040), .dinb(n28895), .dout(n29041));
  jxor g11779(.dina(n28889), .dinb(n347), .dout(n29042));
  jand g11780(.dina(n29042), .dinb(n29041), .dout(n29043));
  jor  g11781(.dina(n29043), .dinb(n28890), .dout(n29044));
  jxor g11782(.dina(n28884), .dinb(n348), .dout(n29045));
  jand g11783(.dina(n29045), .dinb(n29044), .dout(n29046));
  jor  g11784(.dina(n29046), .dinb(n28885), .dout(n29047));
  jxor g11785(.dina(n28879), .dinb(n349), .dout(n29048));
  jand g11786(.dina(n29048), .dinb(n29047), .dout(n29049));
  jor  g11787(.dina(n29049), .dinb(n28880), .dout(n29050));
  jxor g11788(.dina(n28874), .dinb(n268), .dout(n29051));
  jand g11789(.dina(n29051), .dinb(n29050), .dout(n29052));
  jor  g11790(.dina(n29052), .dinb(n28875), .dout(n29053));
  jxor g11791(.dina(n28869), .dinb(n274), .dout(n29054));
  jand g11792(.dina(n29054), .dinb(n29053), .dout(n29055));
  jor  g11793(.dina(n29055), .dinb(n28870), .dout(n29056));
  jxor g11794(.dina(n28864), .dinb(n269), .dout(n29057));
  jand g11795(.dina(n29057), .dinb(n29056), .dout(n29058));
  jor  g11796(.dina(n29058), .dinb(n28865), .dout(n29059));
  jxor g11797(.dina(n28859), .dinb(n270), .dout(n29060));
  jand g11798(.dina(n29060), .dinb(n29059), .dout(n29061));
  jor  g11799(.dina(n29061), .dinb(n28860), .dout(n29062));
  jxor g11800(.dina(n28854), .dinb(n271), .dout(n29063));
  jand g11801(.dina(n29063), .dinb(n29062), .dout(n29064));
  jor  g11802(.dina(n29064), .dinb(n28855), .dout(n29065));
  jxor g11803(.dina(n28849), .dinb(n338), .dout(n29066));
  jand g11804(.dina(n29066), .dinb(n29065), .dout(n29067));
  jor  g11805(.dina(n29067), .dinb(n28850), .dout(n29068));
  jxor g11806(.dina(n28844), .dinb(n339), .dout(n29069));
  jand g11807(.dina(n29069), .dinb(n29068), .dout(n29070));
  jor  g11808(.dina(n29070), .dinb(n28845), .dout(n29071));
  jxor g11809(.dina(n28839), .dinb(n340), .dout(n29072));
  jand g11810(.dina(n29072), .dinb(n29071), .dout(n29073));
  jor  g11811(.dina(n29073), .dinb(n28840), .dout(n29074));
  jxor g11812(.dina(n28834), .dinb(n275), .dout(n29075));
  jand g11813(.dina(n29075), .dinb(n29074), .dout(n29076));
  jor  g11814(.dina(n29076), .dinb(n28835), .dout(n29077));
  jxor g11815(.dina(n28829), .dinb(n331), .dout(n29078));
  jand g11816(.dina(n29078), .dinb(n29077), .dout(n29079));
  jor  g11817(.dina(n29079), .dinb(n28830), .dout(n29080));
  jxor g11818(.dina(n28824), .dinb(n332), .dout(n29081));
  jand g11819(.dina(n29081), .dinb(n29080), .dout(n29082));
  jor  g11820(.dina(n29082), .dinb(n28825), .dout(n29083));
  jxor g11821(.dina(n28819), .dinb(n333), .dout(n29084));
  jand g11822(.dina(n29084), .dinb(n29083), .dout(n29085));
  jor  g11823(.dina(n29085), .dinb(n28820), .dout(n29086));
  jxor g11824(.dina(n28814), .dinb(n276), .dout(n29087));
  jand g11825(.dina(n29087), .dinb(n29086), .dout(n29088));
  jor  g11826(.dina(n29088), .dinb(n28815), .dout(n29089));
  jxor g11827(.dina(n28809), .dinb(n324), .dout(n29090));
  jand g11828(.dina(n29090), .dinb(n29089), .dout(n29091));
  jor  g11829(.dina(n29091), .dinb(n28810), .dout(n29092));
  jxor g11830(.dina(n28804), .dinb(n325), .dout(n29093));
  jand g11831(.dina(n29093), .dinb(n29092), .dout(n29094));
  jor  g11832(.dina(n29094), .dinb(n28805), .dout(n29095));
  jxor g11833(.dina(n28799), .dinb(n326), .dout(n29096));
  jand g11834(.dina(n29096), .dinb(n29095), .dout(n29097));
  jor  g11835(.dina(n29097), .dinb(n28800), .dout(n29098));
  jxor g11836(.dina(n28794), .dinb(n277), .dout(n29099));
  jand g11837(.dina(n29099), .dinb(n29098), .dout(n29100));
  jor  g11838(.dina(n29100), .dinb(n28795), .dout(n29101));
  jxor g11839(.dina(n28789), .dinb(n278), .dout(n29102));
  jand g11840(.dina(n29102), .dinb(n29101), .dout(n29103));
  jor  g11841(.dina(n29103), .dinb(n28790), .dout(n29104));
  jxor g11842(.dina(n28784), .dinb(n279), .dout(n29105));
  jand g11843(.dina(n29105), .dinb(n29104), .dout(n29106));
  jor  g11844(.dina(n29106), .dinb(n28785), .dout(n29107));
  jxor g11845(.dina(n28779), .dinb(n280), .dout(n29108));
  jand g11846(.dina(n29108), .dinb(n29107), .dout(n29109));
  jor  g11847(.dina(n29109), .dinb(n28780), .dout(n29110));
  jxor g11848(.dina(n28774), .dinb(n283), .dout(n29111));
  jand g11849(.dina(n29111), .dinb(n29110), .dout(n29112));
  jor  g11850(.dina(n29112), .dinb(n28775), .dout(n29113));
  jnot g11851(.din(n28764), .dout(n29114));
  jand g11852(.dina(n29114), .dinb(n283), .dout(n29115));
  jnot g11853(.din(n29115), .dout(n29116));
  jnot g11854(.din(n28767), .dout(n29117));
  jand g11855(.dina(n29117), .dinb(n28426), .dout(n29118));
  jand g11856(.dina(n29118), .dinb(n29116), .dout(n29119));
  jnot g11857(.din(n28768), .dout(n29120));
  jand g11858(.dina(n27918), .dinb(n848), .dout(n29121));
  jand g11859(.dina(n29121), .dinb(n29120), .dout(n29122));
  jor  g11860(.dina(n29122), .dinb(n29119), .dout(n29123));
  jxor g11861(.dina(n29123), .dinb(b44 ), .dout(n29124));
  jnot g11862(.din(n29124), .dout(n29125));
  jand g11863(.dina(n29125), .dinb(n29113), .dout(n29126));
  jand g11864(.dina(n29126), .dinb(n9062), .dout(n29127));
  jand g11865(.dina(n29123), .dinb(n320), .dout(n29128));
  jor  g11866(.dina(n29128), .dinb(n29127), .dout(n29129));
  jor  g11867(.dina(n29129), .dinb(n28774), .dout(n29130));
  jnot g11868(.din(n29129), .dout(n29131));
  jxor g11869(.dina(n29111), .dinb(n29110), .dout(n29132));
  jor  g11870(.dina(n29132), .dinb(n29131), .dout(n29133));
  jand g11871(.dina(n29133), .dinb(n29130), .dout(n29134));
  jxor g11872(.dina(n29125), .dinb(n29113), .dout(n29135));
  jor  g11873(.dina(n29135), .dinb(n29131), .dout(n29136));
  jor  g11874(.dina(n29127), .dinb(n29123), .dout(n29137));
  jand g11875(.dina(n29137), .dinb(n29136), .dout(n29138));
  jand g11876(.dina(n29138), .dinb(n316), .dout(n29139));
  jnot g11877(.din(n29138), .dout(n29140));
  jand g11878(.dina(n29140), .dinb(b45 ), .dout(n29141));
  jnot g11879(.din(n29141), .dout(n29142));
  jand g11880(.dina(n29134), .dinb(n315), .dout(n29143));
  jor  g11881(.dina(n29129), .dinb(n28779), .dout(n29144));
  jxor g11882(.dina(n29108), .dinb(n29107), .dout(n29145));
  jor  g11883(.dina(n29145), .dinb(n29131), .dout(n29146));
  jand g11884(.dina(n29146), .dinb(n29144), .dout(n29147));
  jand g11885(.dina(n29147), .dinb(n283), .dout(n29148));
  jor  g11886(.dina(n29129), .dinb(n28784), .dout(n29149));
  jxor g11887(.dina(n29105), .dinb(n29104), .dout(n29150));
  jor  g11888(.dina(n29150), .dinb(n29131), .dout(n29151));
  jand g11889(.dina(n29151), .dinb(n29149), .dout(n29152));
  jand g11890(.dina(n29152), .dinb(n280), .dout(n29153));
  jor  g11891(.dina(n29129), .dinb(n28789), .dout(n29154));
  jxor g11892(.dina(n29102), .dinb(n29101), .dout(n29155));
  jor  g11893(.dina(n29155), .dinb(n29131), .dout(n29156));
  jand g11894(.dina(n29156), .dinb(n29154), .dout(n29157));
  jand g11895(.dina(n29157), .dinb(n279), .dout(n29158));
  jor  g11896(.dina(n29129), .dinb(n28794), .dout(n29159));
  jxor g11897(.dina(n29099), .dinb(n29098), .dout(n29160));
  jor  g11898(.dina(n29160), .dinb(n29131), .dout(n29161));
  jand g11899(.dina(n29161), .dinb(n29159), .dout(n29162));
  jand g11900(.dina(n29162), .dinb(n278), .dout(n29163));
  jor  g11901(.dina(n29129), .dinb(n28799), .dout(n29164));
  jxor g11902(.dina(n29096), .dinb(n29095), .dout(n29165));
  jor  g11903(.dina(n29165), .dinb(n29131), .dout(n29166));
  jand g11904(.dina(n29166), .dinb(n29164), .dout(n29167));
  jand g11905(.dina(n29167), .dinb(n277), .dout(n29168));
  jor  g11906(.dina(n29129), .dinb(n28804), .dout(n29169));
  jxor g11907(.dina(n29093), .dinb(n29092), .dout(n29170));
  jor  g11908(.dina(n29170), .dinb(n29131), .dout(n29171));
  jand g11909(.dina(n29171), .dinb(n29169), .dout(n29172));
  jand g11910(.dina(n29172), .dinb(n326), .dout(n29173));
  jor  g11911(.dina(n29129), .dinb(n28809), .dout(n29174));
  jxor g11912(.dina(n29090), .dinb(n29089), .dout(n29175));
  jor  g11913(.dina(n29175), .dinb(n29131), .dout(n29176));
  jand g11914(.dina(n29176), .dinb(n29174), .dout(n29177));
  jand g11915(.dina(n29177), .dinb(n325), .dout(n29178));
  jor  g11916(.dina(n29129), .dinb(n28814), .dout(n29179));
  jxor g11917(.dina(n29087), .dinb(n29086), .dout(n29180));
  jor  g11918(.dina(n29180), .dinb(n29131), .dout(n29181));
  jand g11919(.dina(n29181), .dinb(n29179), .dout(n29182));
  jand g11920(.dina(n29182), .dinb(n324), .dout(n29183));
  jor  g11921(.dina(n29129), .dinb(n28819), .dout(n29184));
  jxor g11922(.dina(n29084), .dinb(n29083), .dout(n29185));
  jor  g11923(.dina(n29185), .dinb(n29131), .dout(n29186));
  jand g11924(.dina(n29186), .dinb(n29184), .dout(n29187));
  jand g11925(.dina(n29187), .dinb(n276), .dout(n29188));
  jor  g11926(.dina(n29129), .dinb(n28824), .dout(n29189));
  jxor g11927(.dina(n29081), .dinb(n29080), .dout(n29190));
  jor  g11928(.dina(n29190), .dinb(n29131), .dout(n29191));
  jand g11929(.dina(n29191), .dinb(n29189), .dout(n29192));
  jand g11930(.dina(n29192), .dinb(n333), .dout(n29193));
  jor  g11931(.dina(n29129), .dinb(n28829), .dout(n29194));
  jxor g11932(.dina(n29078), .dinb(n29077), .dout(n29195));
  jor  g11933(.dina(n29195), .dinb(n29131), .dout(n29196));
  jand g11934(.dina(n29196), .dinb(n29194), .dout(n29197));
  jand g11935(.dina(n29197), .dinb(n332), .dout(n29198));
  jor  g11936(.dina(n29129), .dinb(n28834), .dout(n29199));
  jxor g11937(.dina(n29075), .dinb(n29074), .dout(n29200));
  jor  g11938(.dina(n29200), .dinb(n29131), .dout(n29201));
  jand g11939(.dina(n29201), .dinb(n29199), .dout(n29202));
  jand g11940(.dina(n29202), .dinb(n331), .dout(n29203));
  jor  g11941(.dina(n29129), .dinb(n28839), .dout(n29204));
  jxor g11942(.dina(n29072), .dinb(n29071), .dout(n29205));
  jor  g11943(.dina(n29205), .dinb(n29131), .dout(n29206));
  jand g11944(.dina(n29206), .dinb(n29204), .dout(n29207));
  jand g11945(.dina(n29207), .dinb(n275), .dout(n29208));
  jor  g11946(.dina(n29129), .dinb(n28844), .dout(n29209));
  jxor g11947(.dina(n29069), .dinb(n29068), .dout(n29210));
  jor  g11948(.dina(n29210), .dinb(n29131), .dout(n29211));
  jand g11949(.dina(n29211), .dinb(n29209), .dout(n29212));
  jand g11950(.dina(n29212), .dinb(n340), .dout(n29213));
  jor  g11951(.dina(n29129), .dinb(n28849), .dout(n29214));
  jxor g11952(.dina(n29066), .dinb(n29065), .dout(n29215));
  jor  g11953(.dina(n29215), .dinb(n29131), .dout(n29216));
  jand g11954(.dina(n29216), .dinb(n29214), .dout(n29217));
  jand g11955(.dina(n29217), .dinb(n339), .dout(n29218));
  jor  g11956(.dina(n29129), .dinb(n28854), .dout(n29219));
  jxor g11957(.dina(n29063), .dinb(n29062), .dout(n29220));
  jor  g11958(.dina(n29220), .dinb(n29131), .dout(n29221));
  jand g11959(.dina(n29221), .dinb(n29219), .dout(n29222));
  jand g11960(.dina(n29222), .dinb(n338), .dout(n29223));
  jor  g11961(.dina(n29129), .dinb(n28859), .dout(n29224));
  jxor g11962(.dina(n29060), .dinb(n29059), .dout(n29225));
  jor  g11963(.dina(n29225), .dinb(n29131), .dout(n29226));
  jand g11964(.dina(n29226), .dinb(n29224), .dout(n29227));
  jand g11965(.dina(n29227), .dinb(n271), .dout(n29228));
  jor  g11966(.dina(n29129), .dinb(n28864), .dout(n29229));
  jxor g11967(.dina(n29057), .dinb(n29056), .dout(n29230));
  jor  g11968(.dina(n29230), .dinb(n29131), .dout(n29231));
  jand g11969(.dina(n29231), .dinb(n29229), .dout(n29232));
  jand g11970(.dina(n29232), .dinb(n270), .dout(n29233));
  jor  g11971(.dina(n29129), .dinb(n28869), .dout(n29234));
  jxor g11972(.dina(n29054), .dinb(n29053), .dout(n29235));
  jor  g11973(.dina(n29235), .dinb(n29131), .dout(n29236));
  jand g11974(.dina(n29236), .dinb(n29234), .dout(n29237));
  jand g11975(.dina(n29237), .dinb(n269), .dout(n29238));
  jor  g11976(.dina(n29129), .dinb(n28874), .dout(n29239));
  jxor g11977(.dina(n29051), .dinb(n29050), .dout(n29240));
  jor  g11978(.dina(n29240), .dinb(n29131), .dout(n29241));
  jand g11979(.dina(n29241), .dinb(n29239), .dout(n29242));
  jand g11980(.dina(n29242), .dinb(n274), .dout(n29243));
  jor  g11981(.dina(n29129), .dinb(n28879), .dout(n29244));
  jxor g11982(.dina(n29048), .dinb(n29047), .dout(n29245));
  jor  g11983(.dina(n29245), .dinb(n29131), .dout(n29246));
  jand g11984(.dina(n29246), .dinb(n29244), .dout(n29247));
  jand g11985(.dina(n29247), .dinb(n268), .dout(n29248));
  jor  g11986(.dina(n29129), .dinb(n28884), .dout(n29249));
  jxor g11987(.dina(n29045), .dinb(n29044), .dout(n29250));
  jor  g11988(.dina(n29250), .dinb(n29131), .dout(n29251));
  jand g11989(.dina(n29251), .dinb(n29249), .dout(n29252));
  jand g11990(.dina(n29252), .dinb(n349), .dout(n29253));
  jor  g11991(.dina(n29129), .dinb(n28889), .dout(n29254));
  jxor g11992(.dina(n29042), .dinb(n29041), .dout(n29255));
  jor  g11993(.dina(n29255), .dinb(n29131), .dout(n29256));
  jand g11994(.dina(n29256), .dinb(n29254), .dout(n29257));
  jand g11995(.dina(n29257), .dinb(n348), .dout(n29258));
  jor  g11996(.dina(n29129), .dinb(n28894), .dout(n29259));
  jxor g11997(.dina(n29039), .dinb(n29038), .dout(n29260));
  jor  g11998(.dina(n29260), .dinb(n29131), .dout(n29261));
  jand g11999(.dina(n29261), .dinb(n29259), .dout(n29262));
  jand g12000(.dina(n29262), .dinb(n347), .dout(n29263));
  jor  g12001(.dina(n29129), .dinb(n28899), .dout(n29264));
  jxor g12002(.dina(n29036), .dinb(n29035), .dout(n29265));
  jor  g12003(.dina(n29265), .dinb(n29131), .dout(n29266));
  jand g12004(.dina(n29266), .dinb(n29264), .dout(n29267));
  jand g12005(.dina(n29267), .dinb(n267), .dout(n29268));
  jor  g12006(.dina(n29129), .dinb(n28904), .dout(n29269));
  jxor g12007(.dina(n29033), .dinb(n29032), .dout(n29270));
  jor  g12008(.dina(n29270), .dinb(n29131), .dout(n29271));
  jand g12009(.dina(n29271), .dinb(n29269), .dout(n29272));
  jand g12010(.dina(n29272), .dinb(n266), .dout(n29273));
  jor  g12011(.dina(n29129), .dinb(n28909), .dout(n29274));
  jxor g12012(.dina(n29030), .dinb(n29029), .dout(n29275));
  jor  g12013(.dina(n29275), .dinb(n29131), .dout(n29276));
  jand g12014(.dina(n29276), .dinb(n29274), .dout(n29277));
  jand g12015(.dina(n29277), .dinb(n356), .dout(n29278));
  jor  g12016(.dina(n29129), .dinb(n28914), .dout(n29279));
  jxor g12017(.dina(n29027), .dinb(n29026), .dout(n29280));
  jor  g12018(.dina(n29280), .dinb(n29131), .dout(n29281));
  jand g12019(.dina(n29281), .dinb(n29279), .dout(n29282));
  jand g12020(.dina(n29282), .dinb(n355), .dout(n29283));
  jor  g12021(.dina(n29129), .dinb(n28919), .dout(n29284));
  jxor g12022(.dina(n29024), .dinb(n29023), .dout(n29285));
  jor  g12023(.dina(n29285), .dinb(n29131), .dout(n29286));
  jand g12024(.dina(n29286), .dinb(n29284), .dout(n29287));
  jand g12025(.dina(n29287), .dinb(n364), .dout(n29288));
  jor  g12026(.dina(n29129), .dinb(n28924), .dout(n29289));
  jxor g12027(.dina(n29021), .dinb(n29020), .dout(n29290));
  jor  g12028(.dina(n29290), .dinb(n29131), .dout(n29291));
  jand g12029(.dina(n29291), .dinb(n29289), .dout(n29292));
  jand g12030(.dina(n29292), .dinb(n361), .dout(n29293));
  jor  g12031(.dina(n29129), .dinb(n28929), .dout(n29294));
  jxor g12032(.dina(n29018), .dinb(n29017), .dout(n29295));
  jor  g12033(.dina(n29295), .dinb(n29131), .dout(n29296));
  jand g12034(.dina(n29296), .dinb(n29294), .dout(n29297));
  jand g12035(.dina(n29297), .dinb(n360), .dout(n29298));
  jor  g12036(.dina(n29129), .dinb(n28934), .dout(n29299));
  jxor g12037(.dina(n29015), .dinb(n29014), .dout(n29300));
  jor  g12038(.dina(n29300), .dinb(n29131), .dout(n29301));
  jand g12039(.dina(n29301), .dinb(n29299), .dout(n29302));
  jand g12040(.dina(n29302), .dinb(n363), .dout(n29303));
  jor  g12041(.dina(n29129), .dinb(n28939), .dout(n29304));
  jxor g12042(.dina(n29012), .dinb(n29011), .dout(n29305));
  jor  g12043(.dina(n29305), .dinb(n29131), .dout(n29306));
  jand g12044(.dina(n29306), .dinb(n29304), .dout(n29307));
  jand g12045(.dina(n29307), .dinb(n359), .dout(n29308));
  jor  g12046(.dina(n29129), .dinb(n28944), .dout(n29309));
  jxor g12047(.dina(n29009), .dinb(n29008), .dout(n29310));
  jor  g12048(.dina(n29310), .dinb(n29131), .dout(n29311));
  jand g12049(.dina(n29311), .dinb(n29309), .dout(n29312));
  jand g12050(.dina(n29312), .dinb(n369), .dout(n29313));
  jor  g12051(.dina(n29129), .dinb(n28949), .dout(n29314));
  jxor g12052(.dina(n29006), .dinb(n29005), .dout(n29315));
  jor  g12053(.dina(n29315), .dinb(n29131), .dout(n29316));
  jand g12054(.dina(n29316), .dinb(n29314), .dout(n29317));
  jand g12055(.dina(n29317), .dinb(n368), .dout(n29318));
  jor  g12056(.dina(n29129), .dinb(n28954), .dout(n29319));
  jxor g12057(.dina(n29003), .dinb(n29002), .dout(n29320));
  jor  g12058(.dina(n29320), .dinb(n29131), .dout(n29321));
  jand g12059(.dina(n29321), .dinb(n29319), .dout(n29322));
  jand g12060(.dina(n29322), .dinb(n367), .dout(n29323));
  jor  g12061(.dina(n29129), .dinb(n28959), .dout(n29324));
  jxor g12062(.dina(n29000), .dinb(n28999), .dout(n29325));
  jor  g12063(.dina(n29325), .dinb(n29131), .dout(n29326));
  jand g12064(.dina(n29326), .dinb(n29324), .dout(n29327));
  jand g12065(.dina(n29327), .dinb(n265), .dout(n29328));
  jor  g12066(.dina(n29129), .dinb(n28964), .dout(n29329));
  jxor g12067(.dina(n28997), .dinb(n28996), .dout(n29330));
  jor  g12068(.dina(n29330), .dinb(n29131), .dout(n29331));
  jand g12069(.dina(n29331), .dinb(n29329), .dout(n29332));
  jand g12070(.dina(n29332), .dinb(n378), .dout(n29333));
  jor  g12071(.dina(n29129), .dinb(n28969), .dout(n29334));
  jxor g12072(.dina(n28994), .dinb(n28993), .dout(n29335));
  jor  g12073(.dina(n29335), .dinb(n29131), .dout(n29336));
  jand g12074(.dina(n29336), .dinb(n29334), .dout(n29337));
  jand g12075(.dina(n29337), .dinb(n377), .dout(n29338));
  jor  g12076(.dina(n29129), .dinb(n28974), .dout(n29339));
  jxor g12077(.dina(n28991), .dinb(n28990), .dout(n29340));
  jor  g12078(.dina(n29340), .dinb(n29131), .dout(n29341));
  jand g12079(.dina(n29341), .dinb(n29339), .dout(n29342));
  jand g12080(.dina(n29342), .dinb(n376), .dout(n29343));
  jor  g12081(.dina(n29129), .dinb(n28979), .dout(n29344));
  jxor g12082(.dina(n28988), .dinb(n28987), .dout(n29345));
  jor  g12083(.dina(n29345), .dinb(n29131), .dout(n29346));
  jand g12084(.dina(n29346), .dinb(n29344), .dout(n29347));
  jand g12085(.dina(n29347), .dinb(n264), .dout(n29348));
  jor  g12086(.dina(n29129), .dinb(n28982), .dout(n29349));
  jxor g12087(.dina(n28985), .dinb(n9275), .dout(n29350));
  jor  g12088(.dina(n29350), .dinb(n29131), .dout(n29351));
  jand g12089(.dina(n29351), .dinb(n29349), .dout(n29352));
  jand g12090(.dina(n29352), .dinb(n386), .dout(n29353));
  jand g12091(.dina(n29129), .dinb(b0 ), .dout(n29354));
  jxor g12092(.dina(n29354), .dinb(a19 ), .dout(n29355));
  jand g12093(.dina(n29355), .dinb(n259), .dout(n29356));
  jxor g12094(.dina(n29354), .dinb(n9273), .dout(n29357));
  jxor g12095(.dina(n29357), .dinb(b1 ), .dout(n29358));
  jand g12096(.dina(n29358), .dinb(n9650), .dout(n29359));
  jor  g12097(.dina(n29359), .dinb(n29356), .dout(n29360));
  jxor g12098(.dina(n29352), .dinb(n386), .dout(n29361));
  jand g12099(.dina(n29361), .dinb(n29360), .dout(n29362));
  jor  g12100(.dina(n29362), .dinb(n29353), .dout(n29363));
  jxor g12101(.dina(n29347), .dinb(n264), .dout(n29364));
  jand g12102(.dina(n29364), .dinb(n29363), .dout(n29365));
  jor  g12103(.dina(n29365), .dinb(n29348), .dout(n29366));
  jxor g12104(.dina(n29342), .dinb(n376), .dout(n29367));
  jand g12105(.dina(n29367), .dinb(n29366), .dout(n29368));
  jor  g12106(.dina(n29368), .dinb(n29343), .dout(n29369));
  jxor g12107(.dina(n29337), .dinb(n377), .dout(n29370));
  jand g12108(.dina(n29370), .dinb(n29369), .dout(n29371));
  jor  g12109(.dina(n29371), .dinb(n29338), .dout(n29372));
  jxor g12110(.dina(n29332), .dinb(n378), .dout(n29373));
  jand g12111(.dina(n29373), .dinb(n29372), .dout(n29374));
  jor  g12112(.dina(n29374), .dinb(n29333), .dout(n29375));
  jxor g12113(.dina(n29327), .dinb(n265), .dout(n29376));
  jand g12114(.dina(n29376), .dinb(n29375), .dout(n29377));
  jor  g12115(.dina(n29377), .dinb(n29328), .dout(n29378));
  jxor g12116(.dina(n29322), .dinb(n367), .dout(n29379));
  jand g12117(.dina(n29379), .dinb(n29378), .dout(n29380));
  jor  g12118(.dina(n29380), .dinb(n29323), .dout(n29381));
  jxor g12119(.dina(n29317), .dinb(n368), .dout(n29382));
  jand g12120(.dina(n29382), .dinb(n29381), .dout(n29383));
  jor  g12121(.dina(n29383), .dinb(n29318), .dout(n29384));
  jxor g12122(.dina(n29312), .dinb(n369), .dout(n29385));
  jand g12123(.dina(n29385), .dinb(n29384), .dout(n29386));
  jor  g12124(.dina(n29386), .dinb(n29313), .dout(n29387));
  jxor g12125(.dina(n29307), .dinb(n359), .dout(n29388));
  jand g12126(.dina(n29388), .dinb(n29387), .dout(n29389));
  jor  g12127(.dina(n29389), .dinb(n29308), .dout(n29390));
  jxor g12128(.dina(n29302), .dinb(n363), .dout(n29391));
  jand g12129(.dina(n29391), .dinb(n29390), .dout(n29392));
  jor  g12130(.dina(n29392), .dinb(n29303), .dout(n29393));
  jxor g12131(.dina(n29297), .dinb(n360), .dout(n29394));
  jand g12132(.dina(n29394), .dinb(n29393), .dout(n29395));
  jor  g12133(.dina(n29395), .dinb(n29298), .dout(n29396));
  jxor g12134(.dina(n29292), .dinb(n361), .dout(n29397));
  jand g12135(.dina(n29397), .dinb(n29396), .dout(n29398));
  jor  g12136(.dina(n29398), .dinb(n29293), .dout(n29399));
  jxor g12137(.dina(n29287), .dinb(n364), .dout(n29400));
  jand g12138(.dina(n29400), .dinb(n29399), .dout(n29401));
  jor  g12139(.dina(n29401), .dinb(n29288), .dout(n29402));
  jxor g12140(.dina(n29282), .dinb(n355), .dout(n29403));
  jand g12141(.dina(n29403), .dinb(n29402), .dout(n29404));
  jor  g12142(.dina(n29404), .dinb(n29283), .dout(n29405));
  jxor g12143(.dina(n29277), .dinb(n356), .dout(n29406));
  jand g12144(.dina(n29406), .dinb(n29405), .dout(n29407));
  jor  g12145(.dina(n29407), .dinb(n29278), .dout(n29408));
  jxor g12146(.dina(n29272), .dinb(n266), .dout(n29409));
  jand g12147(.dina(n29409), .dinb(n29408), .dout(n29410));
  jor  g12148(.dina(n29410), .dinb(n29273), .dout(n29411));
  jxor g12149(.dina(n29267), .dinb(n267), .dout(n29412));
  jand g12150(.dina(n29412), .dinb(n29411), .dout(n29413));
  jor  g12151(.dina(n29413), .dinb(n29268), .dout(n29414));
  jxor g12152(.dina(n29262), .dinb(n347), .dout(n29415));
  jand g12153(.dina(n29415), .dinb(n29414), .dout(n29416));
  jor  g12154(.dina(n29416), .dinb(n29263), .dout(n29417));
  jxor g12155(.dina(n29257), .dinb(n348), .dout(n29418));
  jand g12156(.dina(n29418), .dinb(n29417), .dout(n29419));
  jor  g12157(.dina(n29419), .dinb(n29258), .dout(n29420));
  jxor g12158(.dina(n29252), .dinb(n349), .dout(n29421));
  jand g12159(.dina(n29421), .dinb(n29420), .dout(n29422));
  jor  g12160(.dina(n29422), .dinb(n29253), .dout(n29423));
  jxor g12161(.dina(n29247), .dinb(n268), .dout(n29424));
  jand g12162(.dina(n29424), .dinb(n29423), .dout(n29425));
  jor  g12163(.dina(n29425), .dinb(n29248), .dout(n29426));
  jxor g12164(.dina(n29242), .dinb(n274), .dout(n29427));
  jand g12165(.dina(n29427), .dinb(n29426), .dout(n29428));
  jor  g12166(.dina(n29428), .dinb(n29243), .dout(n29429));
  jxor g12167(.dina(n29237), .dinb(n269), .dout(n29430));
  jand g12168(.dina(n29430), .dinb(n29429), .dout(n29431));
  jor  g12169(.dina(n29431), .dinb(n29238), .dout(n29432));
  jxor g12170(.dina(n29232), .dinb(n270), .dout(n29433));
  jand g12171(.dina(n29433), .dinb(n29432), .dout(n29434));
  jor  g12172(.dina(n29434), .dinb(n29233), .dout(n29435));
  jxor g12173(.dina(n29227), .dinb(n271), .dout(n29436));
  jand g12174(.dina(n29436), .dinb(n29435), .dout(n29437));
  jor  g12175(.dina(n29437), .dinb(n29228), .dout(n29438));
  jxor g12176(.dina(n29222), .dinb(n338), .dout(n29439));
  jand g12177(.dina(n29439), .dinb(n29438), .dout(n29440));
  jor  g12178(.dina(n29440), .dinb(n29223), .dout(n29441));
  jxor g12179(.dina(n29217), .dinb(n339), .dout(n29442));
  jand g12180(.dina(n29442), .dinb(n29441), .dout(n29443));
  jor  g12181(.dina(n29443), .dinb(n29218), .dout(n29444));
  jxor g12182(.dina(n29212), .dinb(n340), .dout(n29445));
  jand g12183(.dina(n29445), .dinb(n29444), .dout(n29446));
  jor  g12184(.dina(n29446), .dinb(n29213), .dout(n29447));
  jxor g12185(.dina(n29207), .dinb(n275), .dout(n29448));
  jand g12186(.dina(n29448), .dinb(n29447), .dout(n29449));
  jor  g12187(.dina(n29449), .dinb(n29208), .dout(n29450));
  jxor g12188(.dina(n29202), .dinb(n331), .dout(n29451));
  jand g12189(.dina(n29451), .dinb(n29450), .dout(n29452));
  jor  g12190(.dina(n29452), .dinb(n29203), .dout(n29453));
  jxor g12191(.dina(n29197), .dinb(n332), .dout(n29454));
  jand g12192(.dina(n29454), .dinb(n29453), .dout(n29455));
  jor  g12193(.dina(n29455), .dinb(n29198), .dout(n29456));
  jxor g12194(.dina(n29192), .dinb(n333), .dout(n29457));
  jand g12195(.dina(n29457), .dinb(n29456), .dout(n29458));
  jor  g12196(.dina(n29458), .dinb(n29193), .dout(n29459));
  jxor g12197(.dina(n29187), .dinb(n276), .dout(n29460));
  jand g12198(.dina(n29460), .dinb(n29459), .dout(n29461));
  jor  g12199(.dina(n29461), .dinb(n29188), .dout(n29462));
  jxor g12200(.dina(n29182), .dinb(n324), .dout(n29463));
  jand g12201(.dina(n29463), .dinb(n29462), .dout(n29464));
  jor  g12202(.dina(n29464), .dinb(n29183), .dout(n29465));
  jxor g12203(.dina(n29177), .dinb(n325), .dout(n29466));
  jand g12204(.dina(n29466), .dinb(n29465), .dout(n29467));
  jor  g12205(.dina(n29467), .dinb(n29178), .dout(n29468));
  jxor g12206(.dina(n29172), .dinb(n326), .dout(n29469));
  jand g12207(.dina(n29469), .dinb(n29468), .dout(n29470));
  jor  g12208(.dina(n29470), .dinb(n29173), .dout(n29471));
  jxor g12209(.dina(n29167), .dinb(n277), .dout(n29472));
  jand g12210(.dina(n29472), .dinb(n29471), .dout(n29473));
  jor  g12211(.dina(n29473), .dinb(n29168), .dout(n29474));
  jxor g12212(.dina(n29162), .dinb(n278), .dout(n29475));
  jand g12213(.dina(n29475), .dinb(n29474), .dout(n29476));
  jor  g12214(.dina(n29476), .dinb(n29163), .dout(n29477));
  jxor g12215(.dina(n29157), .dinb(n279), .dout(n29478));
  jand g12216(.dina(n29478), .dinb(n29477), .dout(n29479));
  jor  g12217(.dina(n29479), .dinb(n29158), .dout(n29480));
  jxor g12218(.dina(n29152), .dinb(n280), .dout(n29481));
  jand g12219(.dina(n29481), .dinb(n29480), .dout(n29482));
  jor  g12220(.dina(n29482), .dinb(n29153), .dout(n29483));
  jxor g12221(.dina(n29147), .dinb(n283), .dout(n29484));
  jand g12222(.dina(n29484), .dinb(n29483), .dout(n29485));
  jor  g12223(.dina(n29485), .dinb(n29148), .dout(n29486));
  jxor g12224(.dina(n29134), .dinb(n315), .dout(n29487));
  jand g12225(.dina(n29487), .dinb(n29486), .dout(n29488));
  jor  g12226(.dina(n29488), .dinb(n29143), .dout(n29489));
  jand g12227(.dina(n29489), .dinb(n29142), .dout(n29490));
  jor  g12228(.dina(n29490), .dinb(n29139), .dout(n29491));
  jand g12229(.dina(n29491), .dinb(n9424), .dout(n29492));
  jor  g12230(.dina(n29492), .dinb(n29134), .dout(n29493));
  jnot g12231(.din(n29492), .dout(n29494));
  jxor g12232(.dina(n29487), .dinb(n29486), .dout(n29495));
  jor  g12233(.dina(n29495), .dinb(n29494), .dout(n29496));
  jand g12234(.dina(n29496), .dinb(n29493), .dout(n29497));
  jand g12235(.dina(n29494), .dinb(n29138), .dout(n29498));
  jand g12236(.dina(n29489), .dinb(n29139), .dout(n29499));
  jor  g12237(.dina(n29499), .dinb(n29498), .dout(n29500));
  jand g12238(.dina(n29500), .dinb(n9424), .dout(n29501));
  jand g12239(.dina(n29497), .dinb(n316), .dout(n29502));
  jor  g12240(.dina(n29492), .dinb(n29147), .dout(n29503));
  jxor g12241(.dina(n29484), .dinb(n29483), .dout(n29504));
  jor  g12242(.dina(n29504), .dinb(n29494), .dout(n29505));
  jand g12243(.dina(n29505), .dinb(n29503), .dout(n29506));
  jand g12244(.dina(n29506), .dinb(n315), .dout(n29507));
  jor  g12245(.dina(n29492), .dinb(n29152), .dout(n29508));
  jxor g12246(.dina(n29481), .dinb(n29480), .dout(n29509));
  jor  g12247(.dina(n29509), .dinb(n29494), .dout(n29510));
  jand g12248(.dina(n29510), .dinb(n29508), .dout(n29511));
  jand g12249(.dina(n29511), .dinb(n283), .dout(n29512));
  jor  g12250(.dina(n29492), .dinb(n29157), .dout(n29513));
  jxor g12251(.dina(n29478), .dinb(n29477), .dout(n29514));
  jor  g12252(.dina(n29514), .dinb(n29494), .dout(n29515));
  jand g12253(.dina(n29515), .dinb(n29513), .dout(n29516));
  jand g12254(.dina(n29516), .dinb(n280), .dout(n29517));
  jor  g12255(.dina(n29492), .dinb(n29162), .dout(n29518));
  jxor g12256(.dina(n29475), .dinb(n29474), .dout(n29519));
  jor  g12257(.dina(n29519), .dinb(n29494), .dout(n29520));
  jand g12258(.dina(n29520), .dinb(n29518), .dout(n29521));
  jand g12259(.dina(n29521), .dinb(n279), .dout(n29522));
  jor  g12260(.dina(n29492), .dinb(n29167), .dout(n29523));
  jxor g12261(.dina(n29472), .dinb(n29471), .dout(n29524));
  jor  g12262(.dina(n29524), .dinb(n29494), .dout(n29525));
  jand g12263(.dina(n29525), .dinb(n29523), .dout(n29526));
  jand g12264(.dina(n29526), .dinb(n278), .dout(n29527));
  jor  g12265(.dina(n29492), .dinb(n29172), .dout(n29528));
  jxor g12266(.dina(n29469), .dinb(n29468), .dout(n29529));
  jor  g12267(.dina(n29529), .dinb(n29494), .dout(n29530));
  jand g12268(.dina(n29530), .dinb(n29528), .dout(n29531));
  jand g12269(.dina(n29531), .dinb(n277), .dout(n29532));
  jor  g12270(.dina(n29492), .dinb(n29177), .dout(n29533));
  jxor g12271(.dina(n29466), .dinb(n29465), .dout(n29534));
  jor  g12272(.dina(n29534), .dinb(n29494), .dout(n29535));
  jand g12273(.dina(n29535), .dinb(n29533), .dout(n29536));
  jand g12274(.dina(n29536), .dinb(n326), .dout(n29537));
  jor  g12275(.dina(n29492), .dinb(n29182), .dout(n29538));
  jxor g12276(.dina(n29463), .dinb(n29462), .dout(n29539));
  jor  g12277(.dina(n29539), .dinb(n29494), .dout(n29540));
  jand g12278(.dina(n29540), .dinb(n29538), .dout(n29541));
  jand g12279(.dina(n29541), .dinb(n325), .dout(n29542));
  jor  g12280(.dina(n29492), .dinb(n29187), .dout(n29543));
  jxor g12281(.dina(n29460), .dinb(n29459), .dout(n29544));
  jor  g12282(.dina(n29544), .dinb(n29494), .dout(n29545));
  jand g12283(.dina(n29545), .dinb(n29543), .dout(n29546));
  jand g12284(.dina(n29546), .dinb(n324), .dout(n29547));
  jor  g12285(.dina(n29492), .dinb(n29192), .dout(n29548));
  jxor g12286(.dina(n29457), .dinb(n29456), .dout(n29549));
  jor  g12287(.dina(n29549), .dinb(n29494), .dout(n29550));
  jand g12288(.dina(n29550), .dinb(n29548), .dout(n29551));
  jand g12289(.dina(n29551), .dinb(n276), .dout(n29552));
  jor  g12290(.dina(n29492), .dinb(n29197), .dout(n29553));
  jxor g12291(.dina(n29454), .dinb(n29453), .dout(n29554));
  jor  g12292(.dina(n29554), .dinb(n29494), .dout(n29555));
  jand g12293(.dina(n29555), .dinb(n29553), .dout(n29556));
  jand g12294(.dina(n29556), .dinb(n333), .dout(n29557));
  jor  g12295(.dina(n29492), .dinb(n29202), .dout(n29558));
  jxor g12296(.dina(n29451), .dinb(n29450), .dout(n29559));
  jor  g12297(.dina(n29559), .dinb(n29494), .dout(n29560));
  jand g12298(.dina(n29560), .dinb(n29558), .dout(n29561));
  jand g12299(.dina(n29561), .dinb(n332), .dout(n29562));
  jor  g12300(.dina(n29492), .dinb(n29207), .dout(n29563));
  jxor g12301(.dina(n29448), .dinb(n29447), .dout(n29564));
  jor  g12302(.dina(n29564), .dinb(n29494), .dout(n29565));
  jand g12303(.dina(n29565), .dinb(n29563), .dout(n29566));
  jand g12304(.dina(n29566), .dinb(n331), .dout(n29567));
  jor  g12305(.dina(n29492), .dinb(n29212), .dout(n29568));
  jxor g12306(.dina(n29445), .dinb(n29444), .dout(n29569));
  jor  g12307(.dina(n29569), .dinb(n29494), .dout(n29570));
  jand g12308(.dina(n29570), .dinb(n29568), .dout(n29571));
  jand g12309(.dina(n29571), .dinb(n275), .dout(n29572));
  jor  g12310(.dina(n29492), .dinb(n29217), .dout(n29573));
  jxor g12311(.dina(n29442), .dinb(n29441), .dout(n29574));
  jor  g12312(.dina(n29574), .dinb(n29494), .dout(n29575));
  jand g12313(.dina(n29575), .dinb(n29573), .dout(n29576));
  jand g12314(.dina(n29576), .dinb(n340), .dout(n29577));
  jor  g12315(.dina(n29492), .dinb(n29222), .dout(n29578));
  jxor g12316(.dina(n29439), .dinb(n29438), .dout(n29579));
  jor  g12317(.dina(n29579), .dinb(n29494), .dout(n29580));
  jand g12318(.dina(n29580), .dinb(n29578), .dout(n29581));
  jand g12319(.dina(n29581), .dinb(n339), .dout(n29582));
  jor  g12320(.dina(n29492), .dinb(n29227), .dout(n29583));
  jxor g12321(.dina(n29436), .dinb(n29435), .dout(n29584));
  jor  g12322(.dina(n29584), .dinb(n29494), .dout(n29585));
  jand g12323(.dina(n29585), .dinb(n29583), .dout(n29586));
  jand g12324(.dina(n29586), .dinb(n338), .dout(n29587));
  jor  g12325(.dina(n29492), .dinb(n29232), .dout(n29588));
  jxor g12326(.dina(n29433), .dinb(n29432), .dout(n29589));
  jor  g12327(.dina(n29589), .dinb(n29494), .dout(n29590));
  jand g12328(.dina(n29590), .dinb(n29588), .dout(n29591));
  jand g12329(.dina(n29591), .dinb(n271), .dout(n29592));
  jor  g12330(.dina(n29492), .dinb(n29237), .dout(n29593));
  jxor g12331(.dina(n29430), .dinb(n29429), .dout(n29594));
  jor  g12332(.dina(n29594), .dinb(n29494), .dout(n29595));
  jand g12333(.dina(n29595), .dinb(n29593), .dout(n29596));
  jand g12334(.dina(n29596), .dinb(n270), .dout(n29597));
  jor  g12335(.dina(n29492), .dinb(n29242), .dout(n29598));
  jxor g12336(.dina(n29427), .dinb(n29426), .dout(n29599));
  jor  g12337(.dina(n29599), .dinb(n29494), .dout(n29600));
  jand g12338(.dina(n29600), .dinb(n29598), .dout(n29601));
  jand g12339(.dina(n29601), .dinb(n269), .dout(n29602));
  jor  g12340(.dina(n29492), .dinb(n29247), .dout(n29603));
  jxor g12341(.dina(n29424), .dinb(n29423), .dout(n29604));
  jor  g12342(.dina(n29604), .dinb(n29494), .dout(n29605));
  jand g12343(.dina(n29605), .dinb(n29603), .dout(n29606));
  jand g12344(.dina(n29606), .dinb(n274), .dout(n29607));
  jor  g12345(.dina(n29492), .dinb(n29252), .dout(n29608));
  jxor g12346(.dina(n29421), .dinb(n29420), .dout(n29609));
  jor  g12347(.dina(n29609), .dinb(n29494), .dout(n29610));
  jand g12348(.dina(n29610), .dinb(n29608), .dout(n29611));
  jand g12349(.dina(n29611), .dinb(n268), .dout(n29612));
  jor  g12350(.dina(n29492), .dinb(n29257), .dout(n29613));
  jxor g12351(.dina(n29418), .dinb(n29417), .dout(n29614));
  jor  g12352(.dina(n29614), .dinb(n29494), .dout(n29615));
  jand g12353(.dina(n29615), .dinb(n29613), .dout(n29616));
  jand g12354(.dina(n29616), .dinb(n349), .dout(n29617));
  jor  g12355(.dina(n29492), .dinb(n29262), .dout(n29618));
  jxor g12356(.dina(n29415), .dinb(n29414), .dout(n29619));
  jor  g12357(.dina(n29619), .dinb(n29494), .dout(n29620));
  jand g12358(.dina(n29620), .dinb(n29618), .dout(n29621));
  jand g12359(.dina(n29621), .dinb(n348), .dout(n29622));
  jor  g12360(.dina(n29492), .dinb(n29267), .dout(n29623));
  jxor g12361(.dina(n29412), .dinb(n29411), .dout(n29624));
  jor  g12362(.dina(n29624), .dinb(n29494), .dout(n29625));
  jand g12363(.dina(n29625), .dinb(n29623), .dout(n29626));
  jand g12364(.dina(n29626), .dinb(n347), .dout(n29627));
  jor  g12365(.dina(n29492), .dinb(n29272), .dout(n29628));
  jxor g12366(.dina(n29409), .dinb(n29408), .dout(n29629));
  jor  g12367(.dina(n29629), .dinb(n29494), .dout(n29630));
  jand g12368(.dina(n29630), .dinb(n29628), .dout(n29631));
  jand g12369(.dina(n29631), .dinb(n267), .dout(n29632));
  jor  g12370(.dina(n29492), .dinb(n29277), .dout(n29633));
  jxor g12371(.dina(n29406), .dinb(n29405), .dout(n29634));
  jor  g12372(.dina(n29634), .dinb(n29494), .dout(n29635));
  jand g12373(.dina(n29635), .dinb(n29633), .dout(n29636));
  jand g12374(.dina(n29636), .dinb(n266), .dout(n29637));
  jor  g12375(.dina(n29492), .dinb(n29282), .dout(n29638));
  jxor g12376(.dina(n29403), .dinb(n29402), .dout(n29639));
  jor  g12377(.dina(n29639), .dinb(n29494), .dout(n29640));
  jand g12378(.dina(n29640), .dinb(n29638), .dout(n29641));
  jand g12379(.dina(n29641), .dinb(n356), .dout(n29642));
  jor  g12380(.dina(n29492), .dinb(n29287), .dout(n29643));
  jxor g12381(.dina(n29400), .dinb(n29399), .dout(n29644));
  jor  g12382(.dina(n29644), .dinb(n29494), .dout(n29645));
  jand g12383(.dina(n29645), .dinb(n29643), .dout(n29646));
  jand g12384(.dina(n29646), .dinb(n355), .dout(n29647));
  jor  g12385(.dina(n29492), .dinb(n29292), .dout(n29648));
  jxor g12386(.dina(n29397), .dinb(n29396), .dout(n29649));
  jor  g12387(.dina(n29649), .dinb(n29494), .dout(n29650));
  jand g12388(.dina(n29650), .dinb(n29648), .dout(n29651));
  jand g12389(.dina(n29651), .dinb(n364), .dout(n29652));
  jor  g12390(.dina(n29492), .dinb(n29297), .dout(n29653));
  jxor g12391(.dina(n29394), .dinb(n29393), .dout(n29654));
  jor  g12392(.dina(n29654), .dinb(n29494), .dout(n29655));
  jand g12393(.dina(n29655), .dinb(n29653), .dout(n29656));
  jand g12394(.dina(n29656), .dinb(n361), .dout(n29657));
  jor  g12395(.dina(n29492), .dinb(n29302), .dout(n29658));
  jxor g12396(.dina(n29391), .dinb(n29390), .dout(n29659));
  jor  g12397(.dina(n29659), .dinb(n29494), .dout(n29660));
  jand g12398(.dina(n29660), .dinb(n29658), .dout(n29661));
  jand g12399(.dina(n29661), .dinb(n360), .dout(n29662));
  jor  g12400(.dina(n29492), .dinb(n29307), .dout(n29663));
  jxor g12401(.dina(n29388), .dinb(n29387), .dout(n29664));
  jor  g12402(.dina(n29664), .dinb(n29494), .dout(n29665));
  jand g12403(.dina(n29665), .dinb(n29663), .dout(n29666));
  jand g12404(.dina(n29666), .dinb(n363), .dout(n29667));
  jor  g12405(.dina(n29492), .dinb(n29312), .dout(n29668));
  jxor g12406(.dina(n29385), .dinb(n29384), .dout(n29669));
  jor  g12407(.dina(n29669), .dinb(n29494), .dout(n29670));
  jand g12408(.dina(n29670), .dinb(n29668), .dout(n29671));
  jand g12409(.dina(n29671), .dinb(n359), .dout(n29672));
  jor  g12410(.dina(n29492), .dinb(n29317), .dout(n29673));
  jxor g12411(.dina(n29382), .dinb(n29381), .dout(n29674));
  jor  g12412(.dina(n29674), .dinb(n29494), .dout(n29675));
  jand g12413(.dina(n29675), .dinb(n29673), .dout(n29676));
  jand g12414(.dina(n29676), .dinb(n369), .dout(n29677));
  jor  g12415(.dina(n29492), .dinb(n29322), .dout(n29678));
  jxor g12416(.dina(n29379), .dinb(n29378), .dout(n29679));
  jor  g12417(.dina(n29679), .dinb(n29494), .dout(n29680));
  jand g12418(.dina(n29680), .dinb(n29678), .dout(n29681));
  jand g12419(.dina(n29681), .dinb(n368), .dout(n29682));
  jor  g12420(.dina(n29492), .dinb(n29327), .dout(n29683));
  jxor g12421(.dina(n29376), .dinb(n29375), .dout(n29684));
  jor  g12422(.dina(n29684), .dinb(n29494), .dout(n29685));
  jand g12423(.dina(n29685), .dinb(n29683), .dout(n29686));
  jand g12424(.dina(n29686), .dinb(n367), .dout(n29687));
  jor  g12425(.dina(n29492), .dinb(n29332), .dout(n29688));
  jxor g12426(.dina(n29373), .dinb(n29372), .dout(n29689));
  jor  g12427(.dina(n29689), .dinb(n29494), .dout(n29690));
  jand g12428(.dina(n29690), .dinb(n29688), .dout(n29691));
  jand g12429(.dina(n29691), .dinb(n265), .dout(n29692));
  jor  g12430(.dina(n29492), .dinb(n29337), .dout(n29693));
  jxor g12431(.dina(n29370), .dinb(n29369), .dout(n29694));
  jor  g12432(.dina(n29694), .dinb(n29494), .dout(n29695));
  jand g12433(.dina(n29695), .dinb(n29693), .dout(n29696));
  jand g12434(.dina(n29696), .dinb(n378), .dout(n29697));
  jor  g12435(.dina(n29492), .dinb(n29342), .dout(n29698));
  jxor g12436(.dina(n29367), .dinb(n29366), .dout(n29699));
  jor  g12437(.dina(n29699), .dinb(n29494), .dout(n29700));
  jand g12438(.dina(n29700), .dinb(n29698), .dout(n29701));
  jand g12439(.dina(n29701), .dinb(n377), .dout(n29702));
  jor  g12440(.dina(n29492), .dinb(n29347), .dout(n29703));
  jxor g12441(.dina(n29364), .dinb(n29363), .dout(n29704));
  jor  g12442(.dina(n29704), .dinb(n29494), .dout(n29705));
  jand g12443(.dina(n29705), .dinb(n29703), .dout(n29706));
  jand g12444(.dina(n29706), .dinb(n376), .dout(n29707));
  jor  g12445(.dina(n29492), .dinb(n29352), .dout(n29708));
  jxor g12446(.dina(n29361), .dinb(n29360), .dout(n29709));
  jor  g12447(.dina(n29709), .dinb(n29494), .dout(n29710));
  jand g12448(.dina(n29710), .dinb(n29708), .dout(n29711));
  jand g12449(.dina(n29711), .dinb(n264), .dout(n29712));
  jor  g12450(.dina(n29492), .dinb(n29355), .dout(n29713));
  jxor g12451(.dina(n29358), .dinb(n9650), .dout(n29714));
  jor  g12452(.dina(n29714), .dinb(n29494), .dout(n29715));
  jand g12453(.dina(n29715), .dinb(n29713), .dout(n29716));
  jand g12454(.dina(n29716), .dinb(n386), .dout(n29717));
  jnot g12455(.din(n10015), .dout(n29718));
  jnot g12456(.din(n29139), .dout(n29719));
  jnot g12457(.din(n29143), .dout(n29720));
  jnot g12458(.din(n29148), .dout(n29721));
  jnot g12459(.din(n29153), .dout(n29722));
  jnot g12460(.din(n29158), .dout(n29723));
  jnot g12461(.din(n29163), .dout(n29724));
  jnot g12462(.din(n29168), .dout(n29725));
  jnot g12463(.din(n29173), .dout(n29726));
  jnot g12464(.din(n29178), .dout(n29727));
  jnot g12465(.din(n29183), .dout(n29728));
  jnot g12466(.din(n29188), .dout(n29729));
  jnot g12467(.din(n29193), .dout(n29730));
  jnot g12468(.din(n29198), .dout(n29731));
  jnot g12469(.din(n29203), .dout(n29732));
  jnot g12470(.din(n29208), .dout(n29733));
  jnot g12471(.din(n29213), .dout(n29734));
  jnot g12472(.din(n29218), .dout(n29735));
  jnot g12473(.din(n29223), .dout(n29736));
  jnot g12474(.din(n29228), .dout(n29737));
  jnot g12475(.din(n29233), .dout(n29738));
  jnot g12476(.din(n29238), .dout(n29739));
  jnot g12477(.din(n29243), .dout(n29740));
  jnot g12478(.din(n29248), .dout(n29741));
  jnot g12479(.din(n29253), .dout(n29742));
  jnot g12480(.din(n29258), .dout(n29743));
  jnot g12481(.din(n29263), .dout(n29744));
  jnot g12482(.din(n29268), .dout(n29745));
  jnot g12483(.din(n29273), .dout(n29746));
  jnot g12484(.din(n29278), .dout(n29747));
  jnot g12485(.din(n29283), .dout(n29748));
  jnot g12486(.din(n29288), .dout(n29749));
  jnot g12487(.din(n29293), .dout(n29750));
  jnot g12488(.din(n29298), .dout(n29751));
  jnot g12489(.din(n29303), .dout(n29752));
  jnot g12490(.din(n29308), .dout(n29753));
  jnot g12491(.din(n29313), .dout(n29754));
  jnot g12492(.din(n29318), .dout(n29755));
  jnot g12493(.din(n29323), .dout(n29756));
  jnot g12494(.din(n29328), .dout(n29757));
  jnot g12495(.din(n29333), .dout(n29758));
  jnot g12496(.din(n29338), .dout(n29759));
  jnot g12497(.din(n29343), .dout(n29760));
  jnot g12498(.din(n29348), .dout(n29761));
  jnot g12499(.din(n29353), .dout(n29762));
  jnot g12500(.din(n29356), .dout(n29763));
  jxor g12501(.dina(n29357), .dinb(n259), .dout(n29764));
  jor  g12502(.dina(n29764), .dinb(n9649), .dout(n29765));
  jand g12503(.dina(n29765), .dinb(n29763), .dout(n29766));
  jnot g12504(.din(n29361), .dout(n29767));
  jor  g12505(.dina(n29767), .dinb(n29766), .dout(n29768));
  jand g12506(.dina(n29768), .dinb(n29762), .dout(n29769));
  jnot g12507(.din(n29364), .dout(n29770));
  jor  g12508(.dina(n29770), .dinb(n29769), .dout(n29771));
  jand g12509(.dina(n29771), .dinb(n29761), .dout(n29772));
  jnot g12510(.din(n29367), .dout(n29773));
  jor  g12511(.dina(n29773), .dinb(n29772), .dout(n29774));
  jand g12512(.dina(n29774), .dinb(n29760), .dout(n29775));
  jnot g12513(.din(n29370), .dout(n29776));
  jor  g12514(.dina(n29776), .dinb(n29775), .dout(n29777));
  jand g12515(.dina(n29777), .dinb(n29759), .dout(n29778));
  jnot g12516(.din(n29373), .dout(n29779));
  jor  g12517(.dina(n29779), .dinb(n29778), .dout(n29780));
  jand g12518(.dina(n29780), .dinb(n29758), .dout(n29781));
  jnot g12519(.din(n29376), .dout(n29782));
  jor  g12520(.dina(n29782), .dinb(n29781), .dout(n29783));
  jand g12521(.dina(n29783), .dinb(n29757), .dout(n29784));
  jnot g12522(.din(n29379), .dout(n29785));
  jor  g12523(.dina(n29785), .dinb(n29784), .dout(n29786));
  jand g12524(.dina(n29786), .dinb(n29756), .dout(n29787));
  jnot g12525(.din(n29382), .dout(n29788));
  jor  g12526(.dina(n29788), .dinb(n29787), .dout(n29789));
  jand g12527(.dina(n29789), .dinb(n29755), .dout(n29790));
  jnot g12528(.din(n29385), .dout(n29791));
  jor  g12529(.dina(n29791), .dinb(n29790), .dout(n29792));
  jand g12530(.dina(n29792), .dinb(n29754), .dout(n29793));
  jnot g12531(.din(n29388), .dout(n29794));
  jor  g12532(.dina(n29794), .dinb(n29793), .dout(n29795));
  jand g12533(.dina(n29795), .dinb(n29753), .dout(n29796));
  jnot g12534(.din(n29391), .dout(n29797));
  jor  g12535(.dina(n29797), .dinb(n29796), .dout(n29798));
  jand g12536(.dina(n29798), .dinb(n29752), .dout(n29799));
  jnot g12537(.din(n29394), .dout(n29800));
  jor  g12538(.dina(n29800), .dinb(n29799), .dout(n29801));
  jand g12539(.dina(n29801), .dinb(n29751), .dout(n29802));
  jnot g12540(.din(n29397), .dout(n29803));
  jor  g12541(.dina(n29803), .dinb(n29802), .dout(n29804));
  jand g12542(.dina(n29804), .dinb(n29750), .dout(n29805));
  jnot g12543(.din(n29400), .dout(n29806));
  jor  g12544(.dina(n29806), .dinb(n29805), .dout(n29807));
  jand g12545(.dina(n29807), .dinb(n29749), .dout(n29808));
  jnot g12546(.din(n29403), .dout(n29809));
  jor  g12547(.dina(n29809), .dinb(n29808), .dout(n29810));
  jand g12548(.dina(n29810), .dinb(n29748), .dout(n29811));
  jnot g12549(.din(n29406), .dout(n29812));
  jor  g12550(.dina(n29812), .dinb(n29811), .dout(n29813));
  jand g12551(.dina(n29813), .dinb(n29747), .dout(n29814));
  jnot g12552(.din(n29409), .dout(n29815));
  jor  g12553(.dina(n29815), .dinb(n29814), .dout(n29816));
  jand g12554(.dina(n29816), .dinb(n29746), .dout(n29817));
  jnot g12555(.din(n29412), .dout(n29818));
  jor  g12556(.dina(n29818), .dinb(n29817), .dout(n29819));
  jand g12557(.dina(n29819), .dinb(n29745), .dout(n29820));
  jnot g12558(.din(n29415), .dout(n29821));
  jor  g12559(.dina(n29821), .dinb(n29820), .dout(n29822));
  jand g12560(.dina(n29822), .dinb(n29744), .dout(n29823));
  jnot g12561(.din(n29418), .dout(n29824));
  jor  g12562(.dina(n29824), .dinb(n29823), .dout(n29825));
  jand g12563(.dina(n29825), .dinb(n29743), .dout(n29826));
  jnot g12564(.din(n29421), .dout(n29827));
  jor  g12565(.dina(n29827), .dinb(n29826), .dout(n29828));
  jand g12566(.dina(n29828), .dinb(n29742), .dout(n29829));
  jnot g12567(.din(n29424), .dout(n29830));
  jor  g12568(.dina(n29830), .dinb(n29829), .dout(n29831));
  jand g12569(.dina(n29831), .dinb(n29741), .dout(n29832));
  jnot g12570(.din(n29427), .dout(n29833));
  jor  g12571(.dina(n29833), .dinb(n29832), .dout(n29834));
  jand g12572(.dina(n29834), .dinb(n29740), .dout(n29835));
  jnot g12573(.din(n29430), .dout(n29836));
  jor  g12574(.dina(n29836), .dinb(n29835), .dout(n29837));
  jand g12575(.dina(n29837), .dinb(n29739), .dout(n29838));
  jnot g12576(.din(n29433), .dout(n29839));
  jor  g12577(.dina(n29839), .dinb(n29838), .dout(n29840));
  jand g12578(.dina(n29840), .dinb(n29738), .dout(n29841));
  jnot g12579(.din(n29436), .dout(n29842));
  jor  g12580(.dina(n29842), .dinb(n29841), .dout(n29843));
  jand g12581(.dina(n29843), .dinb(n29737), .dout(n29844));
  jnot g12582(.din(n29439), .dout(n29845));
  jor  g12583(.dina(n29845), .dinb(n29844), .dout(n29846));
  jand g12584(.dina(n29846), .dinb(n29736), .dout(n29847));
  jnot g12585(.din(n29442), .dout(n29848));
  jor  g12586(.dina(n29848), .dinb(n29847), .dout(n29849));
  jand g12587(.dina(n29849), .dinb(n29735), .dout(n29850));
  jnot g12588(.din(n29445), .dout(n29851));
  jor  g12589(.dina(n29851), .dinb(n29850), .dout(n29852));
  jand g12590(.dina(n29852), .dinb(n29734), .dout(n29853));
  jnot g12591(.din(n29448), .dout(n29854));
  jor  g12592(.dina(n29854), .dinb(n29853), .dout(n29855));
  jand g12593(.dina(n29855), .dinb(n29733), .dout(n29856));
  jnot g12594(.din(n29451), .dout(n29857));
  jor  g12595(.dina(n29857), .dinb(n29856), .dout(n29858));
  jand g12596(.dina(n29858), .dinb(n29732), .dout(n29859));
  jnot g12597(.din(n29454), .dout(n29860));
  jor  g12598(.dina(n29860), .dinb(n29859), .dout(n29861));
  jand g12599(.dina(n29861), .dinb(n29731), .dout(n29862));
  jnot g12600(.din(n29457), .dout(n29863));
  jor  g12601(.dina(n29863), .dinb(n29862), .dout(n29864));
  jand g12602(.dina(n29864), .dinb(n29730), .dout(n29865));
  jnot g12603(.din(n29460), .dout(n29866));
  jor  g12604(.dina(n29866), .dinb(n29865), .dout(n29867));
  jand g12605(.dina(n29867), .dinb(n29729), .dout(n29868));
  jnot g12606(.din(n29463), .dout(n29869));
  jor  g12607(.dina(n29869), .dinb(n29868), .dout(n29870));
  jand g12608(.dina(n29870), .dinb(n29728), .dout(n29871));
  jnot g12609(.din(n29466), .dout(n29872));
  jor  g12610(.dina(n29872), .dinb(n29871), .dout(n29873));
  jand g12611(.dina(n29873), .dinb(n29727), .dout(n29874));
  jnot g12612(.din(n29469), .dout(n29875));
  jor  g12613(.dina(n29875), .dinb(n29874), .dout(n29876));
  jand g12614(.dina(n29876), .dinb(n29726), .dout(n29877));
  jnot g12615(.din(n29472), .dout(n29878));
  jor  g12616(.dina(n29878), .dinb(n29877), .dout(n29879));
  jand g12617(.dina(n29879), .dinb(n29725), .dout(n29880));
  jnot g12618(.din(n29475), .dout(n29881));
  jor  g12619(.dina(n29881), .dinb(n29880), .dout(n29882));
  jand g12620(.dina(n29882), .dinb(n29724), .dout(n29883));
  jnot g12621(.din(n29478), .dout(n29884));
  jor  g12622(.dina(n29884), .dinb(n29883), .dout(n29885));
  jand g12623(.dina(n29885), .dinb(n29723), .dout(n29886));
  jnot g12624(.din(n29481), .dout(n29887));
  jor  g12625(.dina(n29887), .dinb(n29886), .dout(n29888));
  jand g12626(.dina(n29888), .dinb(n29722), .dout(n29889));
  jnot g12627(.din(n29484), .dout(n29890));
  jor  g12628(.dina(n29890), .dinb(n29889), .dout(n29891));
  jand g12629(.dina(n29891), .dinb(n29721), .dout(n29892));
  jnot g12630(.din(n29487), .dout(n29893));
  jor  g12631(.dina(n29893), .dinb(n29892), .dout(n29894));
  jand g12632(.dina(n29894), .dinb(n29720), .dout(n29895));
  jor  g12633(.dina(n29895), .dinb(n29141), .dout(n29896));
  jand g12634(.dina(n29896), .dinb(n29719), .dout(n29897));
  jor  g12635(.dina(n29897), .dinb(n29718), .dout(n29898));
  jand g12636(.dina(n29898), .dinb(a18 ), .dout(n29899));
  jnot g12637(.din(n10018), .dout(n29900));
  jor  g12638(.dina(n29897), .dinb(n29900), .dout(n29901));
  jnot g12639(.din(n29901), .dout(n29902));
  jor  g12640(.dina(n29902), .dinb(n29899), .dout(n29903));
  jand g12641(.dina(n29903), .dinb(n259), .dout(n29904));
  jand g12642(.dina(n29491), .dinb(n10015), .dout(n29905));
  jor  g12643(.dina(n29905), .dinb(n9648), .dout(n29906));
  jand g12644(.dina(n29901), .dinb(n29906), .dout(n29907));
  jxor g12645(.dina(n29907), .dinb(b1 ), .dout(n29908));
  jand g12646(.dina(n29908), .dinb(n10026), .dout(n29909));
  jor  g12647(.dina(n29909), .dinb(n29904), .dout(n29910));
  jxor g12648(.dina(n29716), .dinb(n386), .dout(n29911));
  jand g12649(.dina(n29911), .dinb(n29910), .dout(n29912));
  jor  g12650(.dina(n29912), .dinb(n29717), .dout(n29913));
  jxor g12651(.dina(n29711), .dinb(n264), .dout(n29914));
  jand g12652(.dina(n29914), .dinb(n29913), .dout(n29915));
  jor  g12653(.dina(n29915), .dinb(n29712), .dout(n29916));
  jxor g12654(.dina(n29706), .dinb(n376), .dout(n29917));
  jand g12655(.dina(n29917), .dinb(n29916), .dout(n29918));
  jor  g12656(.dina(n29918), .dinb(n29707), .dout(n29919));
  jxor g12657(.dina(n29701), .dinb(n377), .dout(n29920));
  jand g12658(.dina(n29920), .dinb(n29919), .dout(n29921));
  jor  g12659(.dina(n29921), .dinb(n29702), .dout(n29922));
  jxor g12660(.dina(n29696), .dinb(n378), .dout(n29923));
  jand g12661(.dina(n29923), .dinb(n29922), .dout(n29924));
  jor  g12662(.dina(n29924), .dinb(n29697), .dout(n29925));
  jxor g12663(.dina(n29691), .dinb(n265), .dout(n29926));
  jand g12664(.dina(n29926), .dinb(n29925), .dout(n29927));
  jor  g12665(.dina(n29927), .dinb(n29692), .dout(n29928));
  jxor g12666(.dina(n29686), .dinb(n367), .dout(n29929));
  jand g12667(.dina(n29929), .dinb(n29928), .dout(n29930));
  jor  g12668(.dina(n29930), .dinb(n29687), .dout(n29931));
  jxor g12669(.dina(n29681), .dinb(n368), .dout(n29932));
  jand g12670(.dina(n29932), .dinb(n29931), .dout(n29933));
  jor  g12671(.dina(n29933), .dinb(n29682), .dout(n29934));
  jxor g12672(.dina(n29676), .dinb(n369), .dout(n29935));
  jand g12673(.dina(n29935), .dinb(n29934), .dout(n29936));
  jor  g12674(.dina(n29936), .dinb(n29677), .dout(n29937));
  jxor g12675(.dina(n29671), .dinb(n359), .dout(n29938));
  jand g12676(.dina(n29938), .dinb(n29937), .dout(n29939));
  jor  g12677(.dina(n29939), .dinb(n29672), .dout(n29940));
  jxor g12678(.dina(n29666), .dinb(n363), .dout(n29941));
  jand g12679(.dina(n29941), .dinb(n29940), .dout(n29942));
  jor  g12680(.dina(n29942), .dinb(n29667), .dout(n29943));
  jxor g12681(.dina(n29661), .dinb(n360), .dout(n29944));
  jand g12682(.dina(n29944), .dinb(n29943), .dout(n29945));
  jor  g12683(.dina(n29945), .dinb(n29662), .dout(n29946));
  jxor g12684(.dina(n29656), .dinb(n361), .dout(n29947));
  jand g12685(.dina(n29947), .dinb(n29946), .dout(n29948));
  jor  g12686(.dina(n29948), .dinb(n29657), .dout(n29949));
  jxor g12687(.dina(n29651), .dinb(n364), .dout(n29950));
  jand g12688(.dina(n29950), .dinb(n29949), .dout(n29951));
  jor  g12689(.dina(n29951), .dinb(n29652), .dout(n29952));
  jxor g12690(.dina(n29646), .dinb(n355), .dout(n29953));
  jand g12691(.dina(n29953), .dinb(n29952), .dout(n29954));
  jor  g12692(.dina(n29954), .dinb(n29647), .dout(n29955));
  jxor g12693(.dina(n29641), .dinb(n356), .dout(n29956));
  jand g12694(.dina(n29956), .dinb(n29955), .dout(n29957));
  jor  g12695(.dina(n29957), .dinb(n29642), .dout(n29958));
  jxor g12696(.dina(n29636), .dinb(n266), .dout(n29959));
  jand g12697(.dina(n29959), .dinb(n29958), .dout(n29960));
  jor  g12698(.dina(n29960), .dinb(n29637), .dout(n29961));
  jxor g12699(.dina(n29631), .dinb(n267), .dout(n29962));
  jand g12700(.dina(n29962), .dinb(n29961), .dout(n29963));
  jor  g12701(.dina(n29963), .dinb(n29632), .dout(n29964));
  jxor g12702(.dina(n29626), .dinb(n347), .dout(n29965));
  jand g12703(.dina(n29965), .dinb(n29964), .dout(n29966));
  jor  g12704(.dina(n29966), .dinb(n29627), .dout(n29967));
  jxor g12705(.dina(n29621), .dinb(n348), .dout(n29968));
  jand g12706(.dina(n29968), .dinb(n29967), .dout(n29969));
  jor  g12707(.dina(n29969), .dinb(n29622), .dout(n29970));
  jxor g12708(.dina(n29616), .dinb(n349), .dout(n29971));
  jand g12709(.dina(n29971), .dinb(n29970), .dout(n29972));
  jor  g12710(.dina(n29972), .dinb(n29617), .dout(n29973));
  jxor g12711(.dina(n29611), .dinb(n268), .dout(n29974));
  jand g12712(.dina(n29974), .dinb(n29973), .dout(n29975));
  jor  g12713(.dina(n29975), .dinb(n29612), .dout(n29976));
  jxor g12714(.dina(n29606), .dinb(n274), .dout(n29977));
  jand g12715(.dina(n29977), .dinb(n29976), .dout(n29978));
  jor  g12716(.dina(n29978), .dinb(n29607), .dout(n29979));
  jxor g12717(.dina(n29601), .dinb(n269), .dout(n29980));
  jand g12718(.dina(n29980), .dinb(n29979), .dout(n29981));
  jor  g12719(.dina(n29981), .dinb(n29602), .dout(n29982));
  jxor g12720(.dina(n29596), .dinb(n270), .dout(n29983));
  jand g12721(.dina(n29983), .dinb(n29982), .dout(n29984));
  jor  g12722(.dina(n29984), .dinb(n29597), .dout(n29985));
  jxor g12723(.dina(n29591), .dinb(n271), .dout(n29986));
  jand g12724(.dina(n29986), .dinb(n29985), .dout(n29987));
  jor  g12725(.dina(n29987), .dinb(n29592), .dout(n29988));
  jxor g12726(.dina(n29586), .dinb(n338), .dout(n29989));
  jand g12727(.dina(n29989), .dinb(n29988), .dout(n29990));
  jor  g12728(.dina(n29990), .dinb(n29587), .dout(n29991));
  jxor g12729(.dina(n29581), .dinb(n339), .dout(n29992));
  jand g12730(.dina(n29992), .dinb(n29991), .dout(n29993));
  jor  g12731(.dina(n29993), .dinb(n29582), .dout(n29994));
  jxor g12732(.dina(n29576), .dinb(n340), .dout(n29995));
  jand g12733(.dina(n29995), .dinb(n29994), .dout(n29996));
  jor  g12734(.dina(n29996), .dinb(n29577), .dout(n29997));
  jxor g12735(.dina(n29571), .dinb(n275), .dout(n29998));
  jand g12736(.dina(n29998), .dinb(n29997), .dout(n29999));
  jor  g12737(.dina(n29999), .dinb(n29572), .dout(n30000));
  jxor g12738(.dina(n29566), .dinb(n331), .dout(n30001));
  jand g12739(.dina(n30001), .dinb(n30000), .dout(n30002));
  jor  g12740(.dina(n30002), .dinb(n29567), .dout(n30003));
  jxor g12741(.dina(n29561), .dinb(n332), .dout(n30004));
  jand g12742(.dina(n30004), .dinb(n30003), .dout(n30005));
  jor  g12743(.dina(n30005), .dinb(n29562), .dout(n30006));
  jxor g12744(.dina(n29556), .dinb(n333), .dout(n30007));
  jand g12745(.dina(n30007), .dinb(n30006), .dout(n30008));
  jor  g12746(.dina(n30008), .dinb(n29557), .dout(n30009));
  jxor g12747(.dina(n29551), .dinb(n276), .dout(n30010));
  jand g12748(.dina(n30010), .dinb(n30009), .dout(n30011));
  jor  g12749(.dina(n30011), .dinb(n29552), .dout(n30012));
  jxor g12750(.dina(n29546), .dinb(n324), .dout(n30013));
  jand g12751(.dina(n30013), .dinb(n30012), .dout(n30014));
  jor  g12752(.dina(n30014), .dinb(n29547), .dout(n30015));
  jxor g12753(.dina(n29541), .dinb(n325), .dout(n30016));
  jand g12754(.dina(n30016), .dinb(n30015), .dout(n30017));
  jor  g12755(.dina(n30017), .dinb(n29542), .dout(n30018));
  jxor g12756(.dina(n29536), .dinb(n326), .dout(n30019));
  jand g12757(.dina(n30019), .dinb(n30018), .dout(n30020));
  jor  g12758(.dina(n30020), .dinb(n29537), .dout(n30021));
  jxor g12759(.dina(n29531), .dinb(n277), .dout(n30022));
  jand g12760(.dina(n30022), .dinb(n30021), .dout(n30023));
  jor  g12761(.dina(n30023), .dinb(n29532), .dout(n30024));
  jxor g12762(.dina(n29526), .dinb(n278), .dout(n30025));
  jand g12763(.dina(n30025), .dinb(n30024), .dout(n30026));
  jor  g12764(.dina(n30026), .dinb(n29527), .dout(n30027));
  jxor g12765(.dina(n29521), .dinb(n279), .dout(n30028));
  jand g12766(.dina(n30028), .dinb(n30027), .dout(n30029));
  jor  g12767(.dina(n30029), .dinb(n29522), .dout(n30030));
  jxor g12768(.dina(n29516), .dinb(n280), .dout(n30031));
  jand g12769(.dina(n30031), .dinb(n30030), .dout(n30032));
  jor  g12770(.dina(n30032), .dinb(n29517), .dout(n30033));
  jxor g12771(.dina(n29511), .dinb(n283), .dout(n30034));
  jand g12772(.dina(n30034), .dinb(n30033), .dout(n30035));
  jor  g12773(.dina(n30035), .dinb(n29512), .dout(n30036));
  jxor g12774(.dina(n29506), .dinb(n315), .dout(n30037));
  jand g12775(.dina(n30037), .dinb(n30036), .dout(n30038));
  jor  g12776(.dina(n30038), .dinb(n29507), .dout(n30039));
  jxor g12777(.dina(n29497), .dinb(n316), .dout(n30040));
  jand g12778(.dina(n30040), .dinb(n30039), .dout(n30041));
  jor  g12779(.dina(n30041), .dinb(n29502), .dout(n30042));
  jxor g12780(.dina(n29500), .dinb(b46 ), .dout(n30043));
  jnot g12781(.din(n30043), .dout(n30044));
  jand g12782(.dina(n30044), .dinb(n30042), .dout(n30045));
  jand g12783(.dina(n30045), .dinb(n403), .dout(n30046));
  jor  g12784(.dina(n30046), .dinb(n29501), .dout(n30047));
  jor  g12785(.dina(n30047), .dinb(n29497), .dout(n30048));
  jnot g12786(.din(n30047), .dout(n30049));
  jxor g12787(.dina(n30040), .dinb(n30039), .dout(n30050));
  jor  g12788(.dina(n30050), .dinb(n30049), .dout(n30051));
  jand g12789(.dina(n30051), .dinb(n30048), .dout(n30052));
  jand g12790(.dina(n30042), .dinb(n29501), .dout(n30053));
  jnot g12791(.din(n30046), .dout(n30054));
  jand g12792(.dina(n29138), .dinb(n10176), .dout(n30055));
  jand g12793(.dina(n30055), .dinb(n30054), .dout(n30056));
  jor  g12794(.dina(n30056), .dinb(n30053), .dout(n30057));
  jand g12795(.dina(n30057), .dinb(n403), .dout(n30058));
  jand g12796(.dina(n30052), .dinb(n317), .dout(n30059));
  jor  g12797(.dina(n30047), .dinb(n29506), .dout(n30060));
  jxor g12798(.dina(n30037), .dinb(n30036), .dout(n30061));
  jor  g12799(.dina(n30061), .dinb(n30049), .dout(n30062));
  jand g12800(.dina(n30062), .dinb(n30060), .dout(n30063));
  jand g12801(.dina(n30063), .dinb(n316), .dout(n30064));
  jor  g12802(.dina(n30047), .dinb(n29511), .dout(n30065));
  jxor g12803(.dina(n30034), .dinb(n30033), .dout(n30066));
  jor  g12804(.dina(n30066), .dinb(n30049), .dout(n30067));
  jand g12805(.dina(n30067), .dinb(n30065), .dout(n30068));
  jand g12806(.dina(n30068), .dinb(n315), .dout(n30069));
  jor  g12807(.dina(n30047), .dinb(n29516), .dout(n30070));
  jxor g12808(.dina(n30031), .dinb(n30030), .dout(n30071));
  jor  g12809(.dina(n30071), .dinb(n30049), .dout(n30072));
  jand g12810(.dina(n30072), .dinb(n30070), .dout(n30073));
  jand g12811(.dina(n30073), .dinb(n283), .dout(n30074));
  jor  g12812(.dina(n30047), .dinb(n29521), .dout(n30075));
  jxor g12813(.dina(n30028), .dinb(n30027), .dout(n30076));
  jor  g12814(.dina(n30076), .dinb(n30049), .dout(n30077));
  jand g12815(.dina(n30077), .dinb(n30075), .dout(n30078));
  jand g12816(.dina(n30078), .dinb(n280), .dout(n30079));
  jor  g12817(.dina(n30047), .dinb(n29526), .dout(n30080));
  jxor g12818(.dina(n30025), .dinb(n30024), .dout(n30081));
  jor  g12819(.dina(n30081), .dinb(n30049), .dout(n30082));
  jand g12820(.dina(n30082), .dinb(n30080), .dout(n30083));
  jand g12821(.dina(n30083), .dinb(n279), .dout(n30084));
  jor  g12822(.dina(n30047), .dinb(n29531), .dout(n30085));
  jxor g12823(.dina(n30022), .dinb(n30021), .dout(n30086));
  jor  g12824(.dina(n30086), .dinb(n30049), .dout(n30087));
  jand g12825(.dina(n30087), .dinb(n30085), .dout(n30088));
  jand g12826(.dina(n30088), .dinb(n278), .dout(n30089));
  jor  g12827(.dina(n30047), .dinb(n29536), .dout(n30090));
  jxor g12828(.dina(n30019), .dinb(n30018), .dout(n30091));
  jor  g12829(.dina(n30091), .dinb(n30049), .dout(n30092));
  jand g12830(.dina(n30092), .dinb(n30090), .dout(n30093));
  jand g12831(.dina(n30093), .dinb(n277), .dout(n30094));
  jor  g12832(.dina(n30047), .dinb(n29541), .dout(n30095));
  jxor g12833(.dina(n30016), .dinb(n30015), .dout(n30096));
  jor  g12834(.dina(n30096), .dinb(n30049), .dout(n30097));
  jand g12835(.dina(n30097), .dinb(n30095), .dout(n30098));
  jand g12836(.dina(n30098), .dinb(n326), .dout(n30099));
  jor  g12837(.dina(n30047), .dinb(n29546), .dout(n30100));
  jxor g12838(.dina(n30013), .dinb(n30012), .dout(n30101));
  jor  g12839(.dina(n30101), .dinb(n30049), .dout(n30102));
  jand g12840(.dina(n30102), .dinb(n30100), .dout(n30103));
  jand g12841(.dina(n30103), .dinb(n325), .dout(n30104));
  jor  g12842(.dina(n30047), .dinb(n29551), .dout(n30105));
  jxor g12843(.dina(n30010), .dinb(n30009), .dout(n30106));
  jor  g12844(.dina(n30106), .dinb(n30049), .dout(n30107));
  jand g12845(.dina(n30107), .dinb(n30105), .dout(n30108));
  jand g12846(.dina(n30108), .dinb(n324), .dout(n30109));
  jor  g12847(.dina(n30047), .dinb(n29556), .dout(n30110));
  jxor g12848(.dina(n30007), .dinb(n30006), .dout(n30111));
  jor  g12849(.dina(n30111), .dinb(n30049), .dout(n30112));
  jand g12850(.dina(n30112), .dinb(n30110), .dout(n30113));
  jand g12851(.dina(n30113), .dinb(n276), .dout(n30114));
  jor  g12852(.dina(n30047), .dinb(n29561), .dout(n30115));
  jxor g12853(.dina(n30004), .dinb(n30003), .dout(n30116));
  jor  g12854(.dina(n30116), .dinb(n30049), .dout(n30117));
  jand g12855(.dina(n30117), .dinb(n30115), .dout(n30118));
  jand g12856(.dina(n30118), .dinb(n333), .dout(n30119));
  jor  g12857(.dina(n30047), .dinb(n29566), .dout(n30120));
  jxor g12858(.dina(n30001), .dinb(n30000), .dout(n30121));
  jor  g12859(.dina(n30121), .dinb(n30049), .dout(n30122));
  jand g12860(.dina(n30122), .dinb(n30120), .dout(n30123));
  jand g12861(.dina(n30123), .dinb(n332), .dout(n30124));
  jor  g12862(.dina(n30047), .dinb(n29571), .dout(n30125));
  jxor g12863(.dina(n29998), .dinb(n29997), .dout(n30126));
  jor  g12864(.dina(n30126), .dinb(n30049), .dout(n30127));
  jand g12865(.dina(n30127), .dinb(n30125), .dout(n30128));
  jand g12866(.dina(n30128), .dinb(n331), .dout(n30129));
  jor  g12867(.dina(n30047), .dinb(n29576), .dout(n30130));
  jxor g12868(.dina(n29995), .dinb(n29994), .dout(n30131));
  jor  g12869(.dina(n30131), .dinb(n30049), .dout(n30132));
  jand g12870(.dina(n30132), .dinb(n30130), .dout(n30133));
  jand g12871(.dina(n30133), .dinb(n275), .dout(n30134));
  jor  g12872(.dina(n30047), .dinb(n29581), .dout(n30135));
  jxor g12873(.dina(n29992), .dinb(n29991), .dout(n30136));
  jor  g12874(.dina(n30136), .dinb(n30049), .dout(n30137));
  jand g12875(.dina(n30137), .dinb(n30135), .dout(n30138));
  jand g12876(.dina(n30138), .dinb(n340), .dout(n30139));
  jor  g12877(.dina(n30047), .dinb(n29586), .dout(n30140));
  jxor g12878(.dina(n29989), .dinb(n29988), .dout(n30141));
  jor  g12879(.dina(n30141), .dinb(n30049), .dout(n30142));
  jand g12880(.dina(n30142), .dinb(n30140), .dout(n30143));
  jand g12881(.dina(n30143), .dinb(n339), .dout(n30144));
  jor  g12882(.dina(n30047), .dinb(n29591), .dout(n30145));
  jxor g12883(.dina(n29986), .dinb(n29985), .dout(n30146));
  jor  g12884(.dina(n30146), .dinb(n30049), .dout(n30147));
  jand g12885(.dina(n30147), .dinb(n30145), .dout(n30148));
  jand g12886(.dina(n30148), .dinb(n338), .dout(n30149));
  jor  g12887(.dina(n30047), .dinb(n29596), .dout(n30150));
  jxor g12888(.dina(n29983), .dinb(n29982), .dout(n30151));
  jor  g12889(.dina(n30151), .dinb(n30049), .dout(n30152));
  jand g12890(.dina(n30152), .dinb(n30150), .dout(n30153));
  jand g12891(.dina(n30153), .dinb(n271), .dout(n30154));
  jor  g12892(.dina(n30047), .dinb(n29601), .dout(n30155));
  jxor g12893(.dina(n29980), .dinb(n29979), .dout(n30156));
  jor  g12894(.dina(n30156), .dinb(n30049), .dout(n30157));
  jand g12895(.dina(n30157), .dinb(n30155), .dout(n30158));
  jand g12896(.dina(n30158), .dinb(n270), .dout(n30159));
  jor  g12897(.dina(n30047), .dinb(n29606), .dout(n30160));
  jxor g12898(.dina(n29977), .dinb(n29976), .dout(n30161));
  jor  g12899(.dina(n30161), .dinb(n30049), .dout(n30162));
  jand g12900(.dina(n30162), .dinb(n30160), .dout(n30163));
  jand g12901(.dina(n30163), .dinb(n269), .dout(n30164));
  jor  g12902(.dina(n30047), .dinb(n29611), .dout(n30165));
  jxor g12903(.dina(n29974), .dinb(n29973), .dout(n30166));
  jor  g12904(.dina(n30166), .dinb(n30049), .dout(n30167));
  jand g12905(.dina(n30167), .dinb(n30165), .dout(n30168));
  jand g12906(.dina(n30168), .dinb(n274), .dout(n30169));
  jor  g12907(.dina(n30047), .dinb(n29616), .dout(n30170));
  jxor g12908(.dina(n29971), .dinb(n29970), .dout(n30171));
  jor  g12909(.dina(n30171), .dinb(n30049), .dout(n30172));
  jand g12910(.dina(n30172), .dinb(n30170), .dout(n30173));
  jand g12911(.dina(n30173), .dinb(n268), .dout(n30174));
  jor  g12912(.dina(n30047), .dinb(n29621), .dout(n30175));
  jxor g12913(.dina(n29968), .dinb(n29967), .dout(n30176));
  jor  g12914(.dina(n30176), .dinb(n30049), .dout(n30177));
  jand g12915(.dina(n30177), .dinb(n30175), .dout(n30178));
  jand g12916(.dina(n30178), .dinb(n349), .dout(n30179));
  jor  g12917(.dina(n30047), .dinb(n29626), .dout(n30180));
  jxor g12918(.dina(n29965), .dinb(n29964), .dout(n30181));
  jor  g12919(.dina(n30181), .dinb(n30049), .dout(n30182));
  jand g12920(.dina(n30182), .dinb(n30180), .dout(n30183));
  jand g12921(.dina(n30183), .dinb(n348), .dout(n30184));
  jor  g12922(.dina(n30047), .dinb(n29631), .dout(n30185));
  jxor g12923(.dina(n29962), .dinb(n29961), .dout(n30186));
  jor  g12924(.dina(n30186), .dinb(n30049), .dout(n30187));
  jand g12925(.dina(n30187), .dinb(n30185), .dout(n30188));
  jand g12926(.dina(n30188), .dinb(n347), .dout(n30189));
  jor  g12927(.dina(n30047), .dinb(n29636), .dout(n30190));
  jxor g12928(.dina(n29959), .dinb(n29958), .dout(n30191));
  jor  g12929(.dina(n30191), .dinb(n30049), .dout(n30192));
  jand g12930(.dina(n30192), .dinb(n30190), .dout(n30193));
  jand g12931(.dina(n30193), .dinb(n267), .dout(n30194));
  jor  g12932(.dina(n30047), .dinb(n29641), .dout(n30195));
  jxor g12933(.dina(n29956), .dinb(n29955), .dout(n30196));
  jor  g12934(.dina(n30196), .dinb(n30049), .dout(n30197));
  jand g12935(.dina(n30197), .dinb(n30195), .dout(n30198));
  jand g12936(.dina(n30198), .dinb(n266), .dout(n30199));
  jor  g12937(.dina(n30047), .dinb(n29646), .dout(n30200));
  jxor g12938(.dina(n29953), .dinb(n29952), .dout(n30201));
  jor  g12939(.dina(n30201), .dinb(n30049), .dout(n30202));
  jand g12940(.dina(n30202), .dinb(n30200), .dout(n30203));
  jand g12941(.dina(n30203), .dinb(n356), .dout(n30204));
  jor  g12942(.dina(n30047), .dinb(n29651), .dout(n30205));
  jxor g12943(.dina(n29950), .dinb(n29949), .dout(n30206));
  jor  g12944(.dina(n30206), .dinb(n30049), .dout(n30207));
  jand g12945(.dina(n30207), .dinb(n30205), .dout(n30208));
  jand g12946(.dina(n30208), .dinb(n355), .dout(n30209));
  jor  g12947(.dina(n30047), .dinb(n29656), .dout(n30210));
  jxor g12948(.dina(n29947), .dinb(n29946), .dout(n30211));
  jor  g12949(.dina(n30211), .dinb(n30049), .dout(n30212));
  jand g12950(.dina(n30212), .dinb(n30210), .dout(n30213));
  jand g12951(.dina(n30213), .dinb(n364), .dout(n30214));
  jor  g12952(.dina(n30047), .dinb(n29661), .dout(n30215));
  jxor g12953(.dina(n29944), .dinb(n29943), .dout(n30216));
  jor  g12954(.dina(n30216), .dinb(n30049), .dout(n30217));
  jand g12955(.dina(n30217), .dinb(n30215), .dout(n30218));
  jand g12956(.dina(n30218), .dinb(n361), .dout(n30219));
  jor  g12957(.dina(n30047), .dinb(n29666), .dout(n30220));
  jxor g12958(.dina(n29941), .dinb(n29940), .dout(n30221));
  jor  g12959(.dina(n30221), .dinb(n30049), .dout(n30222));
  jand g12960(.dina(n30222), .dinb(n30220), .dout(n30223));
  jand g12961(.dina(n30223), .dinb(n360), .dout(n30224));
  jor  g12962(.dina(n30047), .dinb(n29671), .dout(n30225));
  jxor g12963(.dina(n29938), .dinb(n29937), .dout(n30226));
  jor  g12964(.dina(n30226), .dinb(n30049), .dout(n30227));
  jand g12965(.dina(n30227), .dinb(n30225), .dout(n30228));
  jand g12966(.dina(n30228), .dinb(n363), .dout(n30229));
  jor  g12967(.dina(n30047), .dinb(n29676), .dout(n30230));
  jxor g12968(.dina(n29935), .dinb(n29934), .dout(n30231));
  jor  g12969(.dina(n30231), .dinb(n30049), .dout(n30232));
  jand g12970(.dina(n30232), .dinb(n30230), .dout(n30233));
  jand g12971(.dina(n30233), .dinb(n359), .dout(n30234));
  jor  g12972(.dina(n30047), .dinb(n29681), .dout(n30235));
  jxor g12973(.dina(n29932), .dinb(n29931), .dout(n30236));
  jor  g12974(.dina(n30236), .dinb(n30049), .dout(n30237));
  jand g12975(.dina(n30237), .dinb(n30235), .dout(n30238));
  jand g12976(.dina(n30238), .dinb(n369), .dout(n30239));
  jor  g12977(.dina(n30047), .dinb(n29686), .dout(n30240));
  jxor g12978(.dina(n29929), .dinb(n29928), .dout(n30241));
  jor  g12979(.dina(n30241), .dinb(n30049), .dout(n30242));
  jand g12980(.dina(n30242), .dinb(n30240), .dout(n30243));
  jand g12981(.dina(n30243), .dinb(n368), .dout(n30244));
  jor  g12982(.dina(n30047), .dinb(n29691), .dout(n30245));
  jxor g12983(.dina(n29926), .dinb(n29925), .dout(n30246));
  jor  g12984(.dina(n30246), .dinb(n30049), .dout(n30247));
  jand g12985(.dina(n30247), .dinb(n30245), .dout(n30248));
  jand g12986(.dina(n30248), .dinb(n367), .dout(n30249));
  jor  g12987(.dina(n30047), .dinb(n29696), .dout(n30250));
  jxor g12988(.dina(n29923), .dinb(n29922), .dout(n30251));
  jor  g12989(.dina(n30251), .dinb(n30049), .dout(n30252));
  jand g12990(.dina(n30252), .dinb(n30250), .dout(n30253));
  jand g12991(.dina(n30253), .dinb(n265), .dout(n30254));
  jor  g12992(.dina(n30047), .dinb(n29701), .dout(n30255));
  jxor g12993(.dina(n29920), .dinb(n29919), .dout(n30256));
  jor  g12994(.dina(n30256), .dinb(n30049), .dout(n30257));
  jand g12995(.dina(n30257), .dinb(n30255), .dout(n30258));
  jand g12996(.dina(n30258), .dinb(n378), .dout(n30259));
  jor  g12997(.dina(n30047), .dinb(n29706), .dout(n30260));
  jxor g12998(.dina(n29917), .dinb(n29916), .dout(n30261));
  jor  g12999(.dina(n30261), .dinb(n30049), .dout(n30262));
  jand g13000(.dina(n30262), .dinb(n30260), .dout(n30263));
  jand g13001(.dina(n30263), .dinb(n377), .dout(n30264));
  jor  g13002(.dina(n30047), .dinb(n29711), .dout(n30265));
  jxor g13003(.dina(n29914), .dinb(n29913), .dout(n30266));
  jor  g13004(.dina(n30266), .dinb(n30049), .dout(n30267));
  jand g13005(.dina(n30267), .dinb(n30265), .dout(n30268));
  jand g13006(.dina(n30268), .dinb(n376), .dout(n30269));
  jor  g13007(.dina(n30047), .dinb(n29716), .dout(n30270));
  jxor g13008(.dina(n29911), .dinb(n29910), .dout(n30271));
  jor  g13009(.dina(n30271), .dinb(n30049), .dout(n30272));
  jand g13010(.dina(n30272), .dinb(n30270), .dout(n30273));
  jand g13011(.dina(n30273), .dinb(n264), .dout(n30274));
  jor  g13012(.dina(n30047), .dinb(n29907), .dout(n30275));
  jxor g13013(.dina(n29908), .dinb(n10026), .dout(n30276));
  jand g13014(.dina(n30276), .dinb(n30047), .dout(n30277));
  jnot g13015(.din(n30277), .dout(n30278));
  jand g13016(.dina(n30278), .dinb(n30275), .dout(n30279));
  jnot g13017(.din(n30279), .dout(n30280));
  jand g13018(.dina(n30280), .dinb(n386), .dout(n30281));
  jand g13019(.dina(n30047), .dinb(b0 ), .dout(n30282));
  jxor g13020(.dina(n30282), .dinb(a17 ), .dout(n30283));
  jand g13021(.dina(n30283), .dinb(n259), .dout(n30284));
  jxor g13022(.dina(n30282), .dinb(n10024), .dout(n30285));
  jxor g13023(.dina(n30285), .dinb(b1 ), .dout(n30286));
  jand g13024(.dina(n30286), .dinb(n10408), .dout(n30287));
  jor  g13025(.dina(n30287), .dinb(n30284), .dout(n30288));
  jxor g13026(.dina(n30279), .dinb(b2 ), .dout(n30289));
  jand g13027(.dina(n30289), .dinb(n30288), .dout(n30290));
  jor  g13028(.dina(n30290), .dinb(n30281), .dout(n30291));
  jxor g13029(.dina(n30273), .dinb(n264), .dout(n30292));
  jand g13030(.dina(n30292), .dinb(n30291), .dout(n30293));
  jor  g13031(.dina(n30293), .dinb(n30274), .dout(n30294));
  jxor g13032(.dina(n30268), .dinb(n376), .dout(n30295));
  jand g13033(.dina(n30295), .dinb(n30294), .dout(n30296));
  jor  g13034(.dina(n30296), .dinb(n30269), .dout(n30297));
  jxor g13035(.dina(n30263), .dinb(n377), .dout(n30298));
  jand g13036(.dina(n30298), .dinb(n30297), .dout(n30299));
  jor  g13037(.dina(n30299), .dinb(n30264), .dout(n30300));
  jxor g13038(.dina(n30258), .dinb(n378), .dout(n30301));
  jand g13039(.dina(n30301), .dinb(n30300), .dout(n30302));
  jor  g13040(.dina(n30302), .dinb(n30259), .dout(n30303));
  jxor g13041(.dina(n30253), .dinb(n265), .dout(n30304));
  jand g13042(.dina(n30304), .dinb(n30303), .dout(n30305));
  jor  g13043(.dina(n30305), .dinb(n30254), .dout(n30306));
  jxor g13044(.dina(n30248), .dinb(n367), .dout(n30307));
  jand g13045(.dina(n30307), .dinb(n30306), .dout(n30308));
  jor  g13046(.dina(n30308), .dinb(n30249), .dout(n30309));
  jxor g13047(.dina(n30243), .dinb(n368), .dout(n30310));
  jand g13048(.dina(n30310), .dinb(n30309), .dout(n30311));
  jor  g13049(.dina(n30311), .dinb(n30244), .dout(n30312));
  jxor g13050(.dina(n30238), .dinb(n369), .dout(n30313));
  jand g13051(.dina(n30313), .dinb(n30312), .dout(n30314));
  jor  g13052(.dina(n30314), .dinb(n30239), .dout(n30315));
  jxor g13053(.dina(n30233), .dinb(n359), .dout(n30316));
  jand g13054(.dina(n30316), .dinb(n30315), .dout(n30317));
  jor  g13055(.dina(n30317), .dinb(n30234), .dout(n30318));
  jxor g13056(.dina(n30228), .dinb(n363), .dout(n30319));
  jand g13057(.dina(n30319), .dinb(n30318), .dout(n30320));
  jor  g13058(.dina(n30320), .dinb(n30229), .dout(n30321));
  jxor g13059(.dina(n30223), .dinb(n360), .dout(n30322));
  jand g13060(.dina(n30322), .dinb(n30321), .dout(n30323));
  jor  g13061(.dina(n30323), .dinb(n30224), .dout(n30324));
  jxor g13062(.dina(n30218), .dinb(n361), .dout(n30325));
  jand g13063(.dina(n30325), .dinb(n30324), .dout(n30326));
  jor  g13064(.dina(n30326), .dinb(n30219), .dout(n30327));
  jxor g13065(.dina(n30213), .dinb(n364), .dout(n30328));
  jand g13066(.dina(n30328), .dinb(n30327), .dout(n30329));
  jor  g13067(.dina(n30329), .dinb(n30214), .dout(n30330));
  jxor g13068(.dina(n30208), .dinb(n355), .dout(n30331));
  jand g13069(.dina(n30331), .dinb(n30330), .dout(n30332));
  jor  g13070(.dina(n30332), .dinb(n30209), .dout(n30333));
  jxor g13071(.dina(n30203), .dinb(n356), .dout(n30334));
  jand g13072(.dina(n30334), .dinb(n30333), .dout(n30335));
  jor  g13073(.dina(n30335), .dinb(n30204), .dout(n30336));
  jxor g13074(.dina(n30198), .dinb(n266), .dout(n30337));
  jand g13075(.dina(n30337), .dinb(n30336), .dout(n30338));
  jor  g13076(.dina(n30338), .dinb(n30199), .dout(n30339));
  jxor g13077(.dina(n30193), .dinb(n267), .dout(n30340));
  jand g13078(.dina(n30340), .dinb(n30339), .dout(n30341));
  jor  g13079(.dina(n30341), .dinb(n30194), .dout(n30342));
  jxor g13080(.dina(n30188), .dinb(n347), .dout(n30343));
  jand g13081(.dina(n30343), .dinb(n30342), .dout(n30344));
  jor  g13082(.dina(n30344), .dinb(n30189), .dout(n30345));
  jxor g13083(.dina(n30183), .dinb(n348), .dout(n30346));
  jand g13084(.dina(n30346), .dinb(n30345), .dout(n30347));
  jor  g13085(.dina(n30347), .dinb(n30184), .dout(n30348));
  jxor g13086(.dina(n30178), .dinb(n349), .dout(n30349));
  jand g13087(.dina(n30349), .dinb(n30348), .dout(n30350));
  jor  g13088(.dina(n30350), .dinb(n30179), .dout(n30351));
  jxor g13089(.dina(n30173), .dinb(n268), .dout(n30352));
  jand g13090(.dina(n30352), .dinb(n30351), .dout(n30353));
  jor  g13091(.dina(n30353), .dinb(n30174), .dout(n30354));
  jxor g13092(.dina(n30168), .dinb(n274), .dout(n30355));
  jand g13093(.dina(n30355), .dinb(n30354), .dout(n30356));
  jor  g13094(.dina(n30356), .dinb(n30169), .dout(n30357));
  jxor g13095(.dina(n30163), .dinb(n269), .dout(n30358));
  jand g13096(.dina(n30358), .dinb(n30357), .dout(n30359));
  jor  g13097(.dina(n30359), .dinb(n30164), .dout(n30360));
  jxor g13098(.dina(n30158), .dinb(n270), .dout(n30361));
  jand g13099(.dina(n30361), .dinb(n30360), .dout(n30362));
  jor  g13100(.dina(n30362), .dinb(n30159), .dout(n30363));
  jxor g13101(.dina(n30153), .dinb(n271), .dout(n30364));
  jand g13102(.dina(n30364), .dinb(n30363), .dout(n30365));
  jor  g13103(.dina(n30365), .dinb(n30154), .dout(n30366));
  jxor g13104(.dina(n30148), .dinb(n338), .dout(n30367));
  jand g13105(.dina(n30367), .dinb(n30366), .dout(n30368));
  jor  g13106(.dina(n30368), .dinb(n30149), .dout(n30369));
  jxor g13107(.dina(n30143), .dinb(n339), .dout(n30370));
  jand g13108(.dina(n30370), .dinb(n30369), .dout(n30371));
  jor  g13109(.dina(n30371), .dinb(n30144), .dout(n30372));
  jxor g13110(.dina(n30138), .dinb(n340), .dout(n30373));
  jand g13111(.dina(n30373), .dinb(n30372), .dout(n30374));
  jor  g13112(.dina(n30374), .dinb(n30139), .dout(n30375));
  jxor g13113(.dina(n30133), .dinb(n275), .dout(n30376));
  jand g13114(.dina(n30376), .dinb(n30375), .dout(n30377));
  jor  g13115(.dina(n30377), .dinb(n30134), .dout(n30378));
  jxor g13116(.dina(n30128), .dinb(n331), .dout(n30379));
  jand g13117(.dina(n30379), .dinb(n30378), .dout(n30380));
  jor  g13118(.dina(n30380), .dinb(n30129), .dout(n30381));
  jxor g13119(.dina(n30123), .dinb(n332), .dout(n30382));
  jand g13120(.dina(n30382), .dinb(n30381), .dout(n30383));
  jor  g13121(.dina(n30383), .dinb(n30124), .dout(n30384));
  jxor g13122(.dina(n30118), .dinb(n333), .dout(n30385));
  jand g13123(.dina(n30385), .dinb(n30384), .dout(n30386));
  jor  g13124(.dina(n30386), .dinb(n30119), .dout(n30387));
  jxor g13125(.dina(n30113), .dinb(n276), .dout(n30388));
  jand g13126(.dina(n30388), .dinb(n30387), .dout(n30389));
  jor  g13127(.dina(n30389), .dinb(n30114), .dout(n30390));
  jxor g13128(.dina(n30108), .dinb(n324), .dout(n30391));
  jand g13129(.dina(n30391), .dinb(n30390), .dout(n30392));
  jor  g13130(.dina(n30392), .dinb(n30109), .dout(n30393));
  jxor g13131(.dina(n30103), .dinb(n325), .dout(n30394));
  jand g13132(.dina(n30394), .dinb(n30393), .dout(n30395));
  jor  g13133(.dina(n30395), .dinb(n30104), .dout(n30396));
  jxor g13134(.dina(n30098), .dinb(n326), .dout(n30397));
  jand g13135(.dina(n30397), .dinb(n30396), .dout(n30398));
  jor  g13136(.dina(n30398), .dinb(n30099), .dout(n30399));
  jxor g13137(.dina(n30093), .dinb(n277), .dout(n30400));
  jand g13138(.dina(n30400), .dinb(n30399), .dout(n30401));
  jor  g13139(.dina(n30401), .dinb(n30094), .dout(n30402));
  jxor g13140(.dina(n30088), .dinb(n278), .dout(n30403));
  jand g13141(.dina(n30403), .dinb(n30402), .dout(n30404));
  jor  g13142(.dina(n30404), .dinb(n30089), .dout(n30405));
  jxor g13143(.dina(n30083), .dinb(n279), .dout(n30406));
  jand g13144(.dina(n30406), .dinb(n30405), .dout(n30407));
  jor  g13145(.dina(n30407), .dinb(n30084), .dout(n30408));
  jxor g13146(.dina(n30078), .dinb(n280), .dout(n30409));
  jand g13147(.dina(n30409), .dinb(n30408), .dout(n30410));
  jor  g13148(.dina(n30410), .dinb(n30079), .dout(n30411));
  jxor g13149(.dina(n30073), .dinb(n283), .dout(n30412));
  jand g13150(.dina(n30412), .dinb(n30411), .dout(n30413));
  jor  g13151(.dina(n30413), .dinb(n30074), .dout(n30414));
  jxor g13152(.dina(n30068), .dinb(n315), .dout(n30415));
  jand g13153(.dina(n30415), .dinb(n30414), .dout(n30416));
  jor  g13154(.dina(n30416), .dinb(n30069), .dout(n30417));
  jxor g13155(.dina(n30063), .dinb(n316), .dout(n30418));
  jand g13156(.dina(n30418), .dinb(n30417), .dout(n30419));
  jor  g13157(.dina(n30419), .dinb(n30064), .dout(n30420));
  jxor g13158(.dina(n30052), .dinb(n317), .dout(n30421));
  jand g13159(.dina(n30421), .dinb(n30420), .dout(n30422));
  jor  g13160(.dina(n30422), .dinb(n30059), .dout(n30423));
  jxor g13161(.dina(n30057), .dinb(b47 ), .dout(n30424));
  jnot g13162(.din(n30424), .dout(n30425));
  jand g13163(.dina(n30425), .dinb(n30423), .dout(n30426));
  jand g13164(.dina(n30426), .dinb(n313), .dout(n30427));
  jor  g13165(.dina(n30427), .dinb(n30058), .dout(n30428));
  jor  g13166(.dina(n30428), .dinb(n30052), .dout(n30429));
  jnot g13167(.din(n30428), .dout(n30430));
  jxor g13168(.dina(n30421), .dinb(n30420), .dout(n30431));
  jor  g13169(.dina(n30431), .dinb(n30430), .dout(n30432));
  jand g13170(.dina(n30432), .dinb(n30429), .dout(n30433));
  jxor g13171(.dina(n30425), .dinb(n30423), .dout(n30434));
  jor  g13172(.dina(n30434), .dinb(n30430), .dout(n30435));
  jor  g13173(.dina(n30427), .dinb(n30057), .dout(n30436));
  jand g13174(.dina(n30436), .dinb(n30435), .dout(n30437));
  jand g13175(.dina(n30437), .dinb(n285), .dout(n30438));
  jnot g13176(.din(n30437), .dout(n30439));
  jand g13177(.dina(n30439), .dinb(b48 ), .dout(n30440));
  jnot g13178(.din(n30440), .dout(n30441));
  jand g13179(.dina(n30433), .dinb(n284), .dout(n30442));
  jor  g13180(.dina(n30428), .dinb(n30063), .dout(n30443));
  jxor g13181(.dina(n30418), .dinb(n30417), .dout(n30444));
  jor  g13182(.dina(n30444), .dinb(n30430), .dout(n30445));
  jand g13183(.dina(n30445), .dinb(n30443), .dout(n30446));
  jand g13184(.dina(n30446), .dinb(n317), .dout(n30447));
  jor  g13185(.dina(n30428), .dinb(n30068), .dout(n30448));
  jxor g13186(.dina(n30415), .dinb(n30414), .dout(n30449));
  jor  g13187(.dina(n30449), .dinb(n30430), .dout(n30450));
  jand g13188(.dina(n30450), .dinb(n30448), .dout(n30451));
  jand g13189(.dina(n30451), .dinb(n316), .dout(n30452));
  jor  g13190(.dina(n30428), .dinb(n30073), .dout(n30453));
  jxor g13191(.dina(n30412), .dinb(n30411), .dout(n30454));
  jor  g13192(.dina(n30454), .dinb(n30430), .dout(n30455));
  jand g13193(.dina(n30455), .dinb(n30453), .dout(n30456));
  jand g13194(.dina(n30456), .dinb(n315), .dout(n30457));
  jor  g13195(.dina(n30428), .dinb(n30078), .dout(n30458));
  jxor g13196(.dina(n30409), .dinb(n30408), .dout(n30459));
  jor  g13197(.dina(n30459), .dinb(n30430), .dout(n30460));
  jand g13198(.dina(n30460), .dinb(n30458), .dout(n30461));
  jand g13199(.dina(n30461), .dinb(n283), .dout(n30462));
  jor  g13200(.dina(n30428), .dinb(n30083), .dout(n30463));
  jxor g13201(.dina(n30406), .dinb(n30405), .dout(n30464));
  jor  g13202(.dina(n30464), .dinb(n30430), .dout(n30465));
  jand g13203(.dina(n30465), .dinb(n30463), .dout(n30466));
  jand g13204(.dina(n30466), .dinb(n280), .dout(n30467));
  jor  g13205(.dina(n30428), .dinb(n30088), .dout(n30468));
  jxor g13206(.dina(n30403), .dinb(n30402), .dout(n30469));
  jor  g13207(.dina(n30469), .dinb(n30430), .dout(n30470));
  jand g13208(.dina(n30470), .dinb(n30468), .dout(n30471));
  jand g13209(.dina(n30471), .dinb(n279), .dout(n30472));
  jor  g13210(.dina(n30428), .dinb(n30093), .dout(n30473));
  jxor g13211(.dina(n30400), .dinb(n30399), .dout(n30474));
  jor  g13212(.dina(n30474), .dinb(n30430), .dout(n30475));
  jand g13213(.dina(n30475), .dinb(n30473), .dout(n30476));
  jand g13214(.dina(n30476), .dinb(n278), .dout(n30477));
  jor  g13215(.dina(n30428), .dinb(n30098), .dout(n30478));
  jxor g13216(.dina(n30397), .dinb(n30396), .dout(n30479));
  jor  g13217(.dina(n30479), .dinb(n30430), .dout(n30480));
  jand g13218(.dina(n30480), .dinb(n30478), .dout(n30481));
  jand g13219(.dina(n30481), .dinb(n277), .dout(n30482));
  jor  g13220(.dina(n30428), .dinb(n30103), .dout(n30483));
  jxor g13221(.dina(n30394), .dinb(n30393), .dout(n30484));
  jor  g13222(.dina(n30484), .dinb(n30430), .dout(n30485));
  jand g13223(.dina(n30485), .dinb(n30483), .dout(n30486));
  jand g13224(.dina(n30486), .dinb(n326), .dout(n30487));
  jor  g13225(.dina(n30428), .dinb(n30108), .dout(n30488));
  jxor g13226(.dina(n30391), .dinb(n30390), .dout(n30489));
  jor  g13227(.dina(n30489), .dinb(n30430), .dout(n30490));
  jand g13228(.dina(n30490), .dinb(n30488), .dout(n30491));
  jand g13229(.dina(n30491), .dinb(n325), .dout(n30492));
  jor  g13230(.dina(n30428), .dinb(n30113), .dout(n30493));
  jxor g13231(.dina(n30388), .dinb(n30387), .dout(n30494));
  jor  g13232(.dina(n30494), .dinb(n30430), .dout(n30495));
  jand g13233(.dina(n30495), .dinb(n30493), .dout(n30496));
  jand g13234(.dina(n30496), .dinb(n324), .dout(n30497));
  jor  g13235(.dina(n30428), .dinb(n30118), .dout(n30498));
  jxor g13236(.dina(n30385), .dinb(n30384), .dout(n30499));
  jor  g13237(.dina(n30499), .dinb(n30430), .dout(n30500));
  jand g13238(.dina(n30500), .dinb(n30498), .dout(n30501));
  jand g13239(.dina(n30501), .dinb(n276), .dout(n30502));
  jor  g13240(.dina(n30428), .dinb(n30123), .dout(n30503));
  jxor g13241(.dina(n30382), .dinb(n30381), .dout(n30504));
  jor  g13242(.dina(n30504), .dinb(n30430), .dout(n30505));
  jand g13243(.dina(n30505), .dinb(n30503), .dout(n30506));
  jand g13244(.dina(n30506), .dinb(n333), .dout(n30507));
  jor  g13245(.dina(n30428), .dinb(n30128), .dout(n30508));
  jxor g13246(.dina(n30379), .dinb(n30378), .dout(n30509));
  jor  g13247(.dina(n30509), .dinb(n30430), .dout(n30510));
  jand g13248(.dina(n30510), .dinb(n30508), .dout(n30511));
  jand g13249(.dina(n30511), .dinb(n332), .dout(n30512));
  jor  g13250(.dina(n30428), .dinb(n30133), .dout(n30513));
  jxor g13251(.dina(n30376), .dinb(n30375), .dout(n30514));
  jor  g13252(.dina(n30514), .dinb(n30430), .dout(n30515));
  jand g13253(.dina(n30515), .dinb(n30513), .dout(n30516));
  jand g13254(.dina(n30516), .dinb(n331), .dout(n30517));
  jor  g13255(.dina(n30428), .dinb(n30138), .dout(n30518));
  jxor g13256(.dina(n30373), .dinb(n30372), .dout(n30519));
  jor  g13257(.dina(n30519), .dinb(n30430), .dout(n30520));
  jand g13258(.dina(n30520), .dinb(n30518), .dout(n30521));
  jand g13259(.dina(n30521), .dinb(n275), .dout(n30522));
  jor  g13260(.dina(n30428), .dinb(n30143), .dout(n30523));
  jxor g13261(.dina(n30370), .dinb(n30369), .dout(n30524));
  jor  g13262(.dina(n30524), .dinb(n30430), .dout(n30525));
  jand g13263(.dina(n30525), .dinb(n30523), .dout(n30526));
  jand g13264(.dina(n30526), .dinb(n340), .dout(n30527));
  jor  g13265(.dina(n30428), .dinb(n30148), .dout(n30528));
  jxor g13266(.dina(n30367), .dinb(n30366), .dout(n30529));
  jor  g13267(.dina(n30529), .dinb(n30430), .dout(n30530));
  jand g13268(.dina(n30530), .dinb(n30528), .dout(n30531));
  jand g13269(.dina(n30531), .dinb(n339), .dout(n30532));
  jor  g13270(.dina(n30428), .dinb(n30153), .dout(n30533));
  jxor g13271(.dina(n30364), .dinb(n30363), .dout(n30534));
  jor  g13272(.dina(n30534), .dinb(n30430), .dout(n30535));
  jand g13273(.dina(n30535), .dinb(n30533), .dout(n30536));
  jand g13274(.dina(n30536), .dinb(n338), .dout(n30537));
  jor  g13275(.dina(n30428), .dinb(n30158), .dout(n30538));
  jxor g13276(.dina(n30361), .dinb(n30360), .dout(n30539));
  jor  g13277(.dina(n30539), .dinb(n30430), .dout(n30540));
  jand g13278(.dina(n30540), .dinb(n30538), .dout(n30541));
  jand g13279(.dina(n30541), .dinb(n271), .dout(n30542));
  jor  g13280(.dina(n30428), .dinb(n30163), .dout(n30543));
  jxor g13281(.dina(n30358), .dinb(n30357), .dout(n30544));
  jor  g13282(.dina(n30544), .dinb(n30430), .dout(n30545));
  jand g13283(.dina(n30545), .dinb(n30543), .dout(n30546));
  jand g13284(.dina(n30546), .dinb(n270), .dout(n30547));
  jor  g13285(.dina(n30428), .dinb(n30168), .dout(n30548));
  jxor g13286(.dina(n30355), .dinb(n30354), .dout(n30549));
  jor  g13287(.dina(n30549), .dinb(n30430), .dout(n30550));
  jand g13288(.dina(n30550), .dinb(n30548), .dout(n30551));
  jand g13289(.dina(n30551), .dinb(n269), .dout(n30552));
  jor  g13290(.dina(n30428), .dinb(n30173), .dout(n30553));
  jxor g13291(.dina(n30352), .dinb(n30351), .dout(n30554));
  jor  g13292(.dina(n30554), .dinb(n30430), .dout(n30555));
  jand g13293(.dina(n30555), .dinb(n30553), .dout(n30556));
  jand g13294(.dina(n30556), .dinb(n274), .dout(n30557));
  jor  g13295(.dina(n30428), .dinb(n30178), .dout(n30558));
  jxor g13296(.dina(n30349), .dinb(n30348), .dout(n30559));
  jor  g13297(.dina(n30559), .dinb(n30430), .dout(n30560));
  jand g13298(.dina(n30560), .dinb(n30558), .dout(n30561));
  jand g13299(.dina(n30561), .dinb(n268), .dout(n30562));
  jor  g13300(.dina(n30428), .dinb(n30183), .dout(n30563));
  jxor g13301(.dina(n30346), .dinb(n30345), .dout(n30564));
  jor  g13302(.dina(n30564), .dinb(n30430), .dout(n30565));
  jand g13303(.dina(n30565), .dinb(n30563), .dout(n30566));
  jand g13304(.dina(n30566), .dinb(n349), .dout(n30567));
  jor  g13305(.dina(n30428), .dinb(n30188), .dout(n30568));
  jxor g13306(.dina(n30343), .dinb(n30342), .dout(n30569));
  jor  g13307(.dina(n30569), .dinb(n30430), .dout(n30570));
  jand g13308(.dina(n30570), .dinb(n30568), .dout(n30571));
  jand g13309(.dina(n30571), .dinb(n348), .dout(n30572));
  jor  g13310(.dina(n30428), .dinb(n30193), .dout(n30573));
  jxor g13311(.dina(n30340), .dinb(n30339), .dout(n30574));
  jor  g13312(.dina(n30574), .dinb(n30430), .dout(n30575));
  jand g13313(.dina(n30575), .dinb(n30573), .dout(n30576));
  jand g13314(.dina(n30576), .dinb(n347), .dout(n30577));
  jor  g13315(.dina(n30428), .dinb(n30198), .dout(n30578));
  jxor g13316(.dina(n30337), .dinb(n30336), .dout(n30579));
  jor  g13317(.dina(n30579), .dinb(n30430), .dout(n30580));
  jand g13318(.dina(n30580), .dinb(n30578), .dout(n30581));
  jand g13319(.dina(n30581), .dinb(n267), .dout(n30582));
  jor  g13320(.dina(n30428), .dinb(n30203), .dout(n30583));
  jxor g13321(.dina(n30334), .dinb(n30333), .dout(n30584));
  jor  g13322(.dina(n30584), .dinb(n30430), .dout(n30585));
  jand g13323(.dina(n30585), .dinb(n30583), .dout(n30586));
  jand g13324(.dina(n30586), .dinb(n266), .dout(n30587));
  jor  g13325(.dina(n30428), .dinb(n30208), .dout(n30588));
  jxor g13326(.dina(n30331), .dinb(n30330), .dout(n30589));
  jor  g13327(.dina(n30589), .dinb(n30430), .dout(n30590));
  jand g13328(.dina(n30590), .dinb(n30588), .dout(n30591));
  jand g13329(.dina(n30591), .dinb(n356), .dout(n30592));
  jor  g13330(.dina(n30428), .dinb(n30213), .dout(n30593));
  jxor g13331(.dina(n30328), .dinb(n30327), .dout(n30594));
  jor  g13332(.dina(n30594), .dinb(n30430), .dout(n30595));
  jand g13333(.dina(n30595), .dinb(n30593), .dout(n30596));
  jand g13334(.dina(n30596), .dinb(n355), .dout(n30597));
  jor  g13335(.dina(n30428), .dinb(n30218), .dout(n30598));
  jxor g13336(.dina(n30325), .dinb(n30324), .dout(n30599));
  jor  g13337(.dina(n30599), .dinb(n30430), .dout(n30600));
  jand g13338(.dina(n30600), .dinb(n30598), .dout(n30601));
  jand g13339(.dina(n30601), .dinb(n364), .dout(n30602));
  jor  g13340(.dina(n30428), .dinb(n30223), .dout(n30603));
  jxor g13341(.dina(n30322), .dinb(n30321), .dout(n30604));
  jor  g13342(.dina(n30604), .dinb(n30430), .dout(n30605));
  jand g13343(.dina(n30605), .dinb(n30603), .dout(n30606));
  jand g13344(.dina(n30606), .dinb(n361), .dout(n30607));
  jor  g13345(.dina(n30428), .dinb(n30228), .dout(n30608));
  jxor g13346(.dina(n30319), .dinb(n30318), .dout(n30609));
  jor  g13347(.dina(n30609), .dinb(n30430), .dout(n30610));
  jand g13348(.dina(n30610), .dinb(n30608), .dout(n30611));
  jand g13349(.dina(n30611), .dinb(n360), .dout(n30612));
  jor  g13350(.dina(n30428), .dinb(n30233), .dout(n30613));
  jxor g13351(.dina(n30316), .dinb(n30315), .dout(n30614));
  jor  g13352(.dina(n30614), .dinb(n30430), .dout(n30615));
  jand g13353(.dina(n30615), .dinb(n30613), .dout(n30616));
  jand g13354(.dina(n30616), .dinb(n363), .dout(n30617));
  jor  g13355(.dina(n30428), .dinb(n30238), .dout(n30618));
  jxor g13356(.dina(n30313), .dinb(n30312), .dout(n30619));
  jor  g13357(.dina(n30619), .dinb(n30430), .dout(n30620));
  jand g13358(.dina(n30620), .dinb(n30618), .dout(n30621));
  jand g13359(.dina(n30621), .dinb(n359), .dout(n30622));
  jor  g13360(.dina(n30428), .dinb(n30243), .dout(n30623));
  jxor g13361(.dina(n30310), .dinb(n30309), .dout(n30624));
  jor  g13362(.dina(n30624), .dinb(n30430), .dout(n30625));
  jand g13363(.dina(n30625), .dinb(n30623), .dout(n30626));
  jand g13364(.dina(n30626), .dinb(n369), .dout(n30627));
  jor  g13365(.dina(n30428), .dinb(n30248), .dout(n30628));
  jxor g13366(.dina(n30307), .dinb(n30306), .dout(n30629));
  jor  g13367(.dina(n30629), .dinb(n30430), .dout(n30630));
  jand g13368(.dina(n30630), .dinb(n30628), .dout(n30631));
  jand g13369(.dina(n30631), .dinb(n368), .dout(n30632));
  jor  g13370(.dina(n30428), .dinb(n30253), .dout(n30633));
  jxor g13371(.dina(n30304), .dinb(n30303), .dout(n30634));
  jor  g13372(.dina(n30634), .dinb(n30430), .dout(n30635));
  jand g13373(.dina(n30635), .dinb(n30633), .dout(n30636));
  jand g13374(.dina(n30636), .dinb(n367), .dout(n30637));
  jor  g13375(.dina(n30428), .dinb(n30258), .dout(n30638));
  jxor g13376(.dina(n30301), .dinb(n30300), .dout(n30639));
  jor  g13377(.dina(n30639), .dinb(n30430), .dout(n30640));
  jand g13378(.dina(n30640), .dinb(n30638), .dout(n30641));
  jand g13379(.dina(n30641), .dinb(n265), .dout(n30642));
  jor  g13380(.dina(n30428), .dinb(n30263), .dout(n30643));
  jxor g13381(.dina(n30298), .dinb(n30297), .dout(n30644));
  jor  g13382(.dina(n30644), .dinb(n30430), .dout(n30645));
  jand g13383(.dina(n30645), .dinb(n30643), .dout(n30646));
  jand g13384(.dina(n30646), .dinb(n378), .dout(n30647));
  jor  g13385(.dina(n30428), .dinb(n30268), .dout(n30648));
  jxor g13386(.dina(n30295), .dinb(n30294), .dout(n30649));
  jor  g13387(.dina(n30649), .dinb(n30430), .dout(n30650));
  jand g13388(.dina(n30650), .dinb(n30648), .dout(n30651));
  jand g13389(.dina(n30651), .dinb(n377), .dout(n30652));
  jor  g13390(.dina(n30428), .dinb(n30273), .dout(n30653));
  jxor g13391(.dina(n30292), .dinb(n30291), .dout(n30654));
  jor  g13392(.dina(n30654), .dinb(n30430), .dout(n30655));
  jand g13393(.dina(n30655), .dinb(n30653), .dout(n30656));
  jand g13394(.dina(n30656), .dinb(n376), .dout(n30657));
  jor  g13395(.dina(n30428), .dinb(n30280), .dout(n30658));
  jxor g13396(.dina(n30289), .dinb(n30288), .dout(n30659));
  jor  g13397(.dina(n30659), .dinb(n30430), .dout(n30660));
  jand g13398(.dina(n30660), .dinb(n30658), .dout(n30661));
  jand g13399(.dina(n30661), .dinb(n264), .dout(n30662));
  jxor g13400(.dina(n30286), .dinb(n10408), .dout(n30663));
  jand g13401(.dina(n30663), .dinb(n30428), .dout(n30664));
  jnot g13402(.din(n30664), .dout(n30665));
  jor  g13403(.dina(n30428), .dinb(n30285), .dout(n30666));
  jand g13404(.dina(n30666), .dinb(n30665), .dout(n30667));
  jnot g13405(.din(n30667), .dout(n30668));
  jand g13406(.dina(n30668), .dinb(n386), .dout(n30669));
  jand g13407(.dina(n30428), .dinb(b0 ), .dout(n30670));
  jxor g13408(.dina(n30670), .dinb(a16 ), .dout(n30671));
  jand g13409(.dina(n30671), .dinb(n259), .dout(n30672));
  jxor g13410(.dina(n30670), .dinb(n10406), .dout(n30673));
  jxor g13411(.dina(n30673), .dinb(b1 ), .dout(n30674));
  jand g13412(.dina(n30674), .dinb(n10799), .dout(n30675));
  jor  g13413(.dina(n30675), .dinb(n30672), .dout(n30676));
  jxor g13414(.dina(n30667), .dinb(b2 ), .dout(n30677));
  jand g13415(.dina(n30677), .dinb(n30676), .dout(n30678));
  jor  g13416(.dina(n30678), .dinb(n30669), .dout(n30679));
  jxor g13417(.dina(n30661), .dinb(n264), .dout(n30680));
  jand g13418(.dina(n30680), .dinb(n30679), .dout(n30681));
  jor  g13419(.dina(n30681), .dinb(n30662), .dout(n30682));
  jxor g13420(.dina(n30656), .dinb(n376), .dout(n30683));
  jand g13421(.dina(n30683), .dinb(n30682), .dout(n30684));
  jor  g13422(.dina(n30684), .dinb(n30657), .dout(n30685));
  jxor g13423(.dina(n30651), .dinb(n377), .dout(n30686));
  jand g13424(.dina(n30686), .dinb(n30685), .dout(n30687));
  jor  g13425(.dina(n30687), .dinb(n30652), .dout(n30688));
  jxor g13426(.dina(n30646), .dinb(n378), .dout(n30689));
  jand g13427(.dina(n30689), .dinb(n30688), .dout(n30690));
  jor  g13428(.dina(n30690), .dinb(n30647), .dout(n30691));
  jxor g13429(.dina(n30641), .dinb(n265), .dout(n30692));
  jand g13430(.dina(n30692), .dinb(n30691), .dout(n30693));
  jor  g13431(.dina(n30693), .dinb(n30642), .dout(n30694));
  jxor g13432(.dina(n30636), .dinb(n367), .dout(n30695));
  jand g13433(.dina(n30695), .dinb(n30694), .dout(n30696));
  jor  g13434(.dina(n30696), .dinb(n30637), .dout(n30697));
  jxor g13435(.dina(n30631), .dinb(n368), .dout(n30698));
  jand g13436(.dina(n30698), .dinb(n30697), .dout(n30699));
  jor  g13437(.dina(n30699), .dinb(n30632), .dout(n30700));
  jxor g13438(.dina(n30626), .dinb(n369), .dout(n30701));
  jand g13439(.dina(n30701), .dinb(n30700), .dout(n30702));
  jor  g13440(.dina(n30702), .dinb(n30627), .dout(n30703));
  jxor g13441(.dina(n30621), .dinb(n359), .dout(n30704));
  jand g13442(.dina(n30704), .dinb(n30703), .dout(n30705));
  jor  g13443(.dina(n30705), .dinb(n30622), .dout(n30706));
  jxor g13444(.dina(n30616), .dinb(n363), .dout(n30707));
  jand g13445(.dina(n30707), .dinb(n30706), .dout(n30708));
  jor  g13446(.dina(n30708), .dinb(n30617), .dout(n30709));
  jxor g13447(.dina(n30611), .dinb(n360), .dout(n30710));
  jand g13448(.dina(n30710), .dinb(n30709), .dout(n30711));
  jor  g13449(.dina(n30711), .dinb(n30612), .dout(n30712));
  jxor g13450(.dina(n30606), .dinb(n361), .dout(n30713));
  jand g13451(.dina(n30713), .dinb(n30712), .dout(n30714));
  jor  g13452(.dina(n30714), .dinb(n30607), .dout(n30715));
  jxor g13453(.dina(n30601), .dinb(n364), .dout(n30716));
  jand g13454(.dina(n30716), .dinb(n30715), .dout(n30717));
  jor  g13455(.dina(n30717), .dinb(n30602), .dout(n30718));
  jxor g13456(.dina(n30596), .dinb(n355), .dout(n30719));
  jand g13457(.dina(n30719), .dinb(n30718), .dout(n30720));
  jor  g13458(.dina(n30720), .dinb(n30597), .dout(n30721));
  jxor g13459(.dina(n30591), .dinb(n356), .dout(n30722));
  jand g13460(.dina(n30722), .dinb(n30721), .dout(n30723));
  jor  g13461(.dina(n30723), .dinb(n30592), .dout(n30724));
  jxor g13462(.dina(n30586), .dinb(n266), .dout(n30725));
  jand g13463(.dina(n30725), .dinb(n30724), .dout(n30726));
  jor  g13464(.dina(n30726), .dinb(n30587), .dout(n30727));
  jxor g13465(.dina(n30581), .dinb(n267), .dout(n30728));
  jand g13466(.dina(n30728), .dinb(n30727), .dout(n30729));
  jor  g13467(.dina(n30729), .dinb(n30582), .dout(n30730));
  jxor g13468(.dina(n30576), .dinb(n347), .dout(n30731));
  jand g13469(.dina(n30731), .dinb(n30730), .dout(n30732));
  jor  g13470(.dina(n30732), .dinb(n30577), .dout(n30733));
  jxor g13471(.dina(n30571), .dinb(n348), .dout(n30734));
  jand g13472(.dina(n30734), .dinb(n30733), .dout(n30735));
  jor  g13473(.dina(n30735), .dinb(n30572), .dout(n30736));
  jxor g13474(.dina(n30566), .dinb(n349), .dout(n30737));
  jand g13475(.dina(n30737), .dinb(n30736), .dout(n30738));
  jor  g13476(.dina(n30738), .dinb(n30567), .dout(n30739));
  jxor g13477(.dina(n30561), .dinb(n268), .dout(n30740));
  jand g13478(.dina(n30740), .dinb(n30739), .dout(n30741));
  jor  g13479(.dina(n30741), .dinb(n30562), .dout(n30742));
  jxor g13480(.dina(n30556), .dinb(n274), .dout(n30743));
  jand g13481(.dina(n30743), .dinb(n30742), .dout(n30744));
  jor  g13482(.dina(n30744), .dinb(n30557), .dout(n30745));
  jxor g13483(.dina(n30551), .dinb(n269), .dout(n30746));
  jand g13484(.dina(n30746), .dinb(n30745), .dout(n30747));
  jor  g13485(.dina(n30747), .dinb(n30552), .dout(n30748));
  jxor g13486(.dina(n30546), .dinb(n270), .dout(n30749));
  jand g13487(.dina(n30749), .dinb(n30748), .dout(n30750));
  jor  g13488(.dina(n30750), .dinb(n30547), .dout(n30751));
  jxor g13489(.dina(n30541), .dinb(n271), .dout(n30752));
  jand g13490(.dina(n30752), .dinb(n30751), .dout(n30753));
  jor  g13491(.dina(n30753), .dinb(n30542), .dout(n30754));
  jxor g13492(.dina(n30536), .dinb(n338), .dout(n30755));
  jand g13493(.dina(n30755), .dinb(n30754), .dout(n30756));
  jor  g13494(.dina(n30756), .dinb(n30537), .dout(n30757));
  jxor g13495(.dina(n30531), .dinb(n339), .dout(n30758));
  jand g13496(.dina(n30758), .dinb(n30757), .dout(n30759));
  jor  g13497(.dina(n30759), .dinb(n30532), .dout(n30760));
  jxor g13498(.dina(n30526), .dinb(n340), .dout(n30761));
  jand g13499(.dina(n30761), .dinb(n30760), .dout(n30762));
  jor  g13500(.dina(n30762), .dinb(n30527), .dout(n30763));
  jxor g13501(.dina(n30521), .dinb(n275), .dout(n30764));
  jand g13502(.dina(n30764), .dinb(n30763), .dout(n30765));
  jor  g13503(.dina(n30765), .dinb(n30522), .dout(n30766));
  jxor g13504(.dina(n30516), .dinb(n331), .dout(n30767));
  jand g13505(.dina(n30767), .dinb(n30766), .dout(n30768));
  jor  g13506(.dina(n30768), .dinb(n30517), .dout(n30769));
  jxor g13507(.dina(n30511), .dinb(n332), .dout(n30770));
  jand g13508(.dina(n30770), .dinb(n30769), .dout(n30771));
  jor  g13509(.dina(n30771), .dinb(n30512), .dout(n30772));
  jxor g13510(.dina(n30506), .dinb(n333), .dout(n30773));
  jand g13511(.dina(n30773), .dinb(n30772), .dout(n30774));
  jor  g13512(.dina(n30774), .dinb(n30507), .dout(n30775));
  jxor g13513(.dina(n30501), .dinb(n276), .dout(n30776));
  jand g13514(.dina(n30776), .dinb(n30775), .dout(n30777));
  jor  g13515(.dina(n30777), .dinb(n30502), .dout(n30778));
  jxor g13516(.dina(n30496), .dinb(n324), .dout(n30779));
  jand g13517(.dina(n30779), .dinb(n30778), .dout(n30780));
  jor  g13518(.dina(n30780), .dinb(n30497), .dout(n30781));
  jxor g13519(.dina(n30491), .dinb(n325), .dout(n30782));
  jand g13520(.dina(n30782), .dinb(n30781), .dout(n30783));
  jor  g13521(.dina(n30783), .dinb(n30492), .dout(n30784));
  jxor g13522(.dina(n30486), .dinb(n326), .dout(n30785));
  jand g13523(.dina(n30785), .dinb(n30784), .dout(n30786));
  jor  g13524(.dina(n30786), .dinb(n30487), .dout(n30787));
  jxor g13525(.dina(n30481), .dinb(n277), .dout(n30788));
  jand g13526(.dina(n30788), .dinb(n30787), .dout(n30789));
  jor  g13527(.dina(n30789), .dinb(n30482), .dout(n30790));
  jxor g13528(.dina(n30476), .dinb(n278), .dout(n30791));
  jand g13529(.dina(n30791), .dinb(n30790), .dout(n30792));
  jor  g13530(.dina(n30792), .dinb(n30477), .dout(n30793));
  jxor g13531(.dina(n30471), .dinb(n279), .dout(n30794));
  jand g13532(.dina(n30794), .dinb(n30793), .dout(n30795));
  jor  g13533(.dina(n30795), .dinb(n30472), .dout(n30796));
  jxor g13534(.dina(n30466), .dinb(n280), .dout(n30797));
  jand g13535(.dina(n30797), .dinb(n30796), .dout(n30798));
  jor  g13536(.dina(n30798), .dinb(n30467), .dout(n30799));
  jxor g13537(.dina(n30461), .dinb(n283), .dout(n30800));
  jand g13538(.dina(n30800), .dinb(n30799), .dout(n30801));
  jor  g13539(.dina(n30801), .dinb(n30462), .dout(n30802));
  jxor g13540(.dina(n30456), .dinb(n315), .dout(n30803));
  jand g13541(.dina(n30803), .dinb(n30802), .dout(n30804));
  jor  g13542(.dina(n30804), .dinb(n30457), .dout(n30805));
  jxor g13543(.dina(n30451), .dinb(n316), .dout(n30806));
  jand g13544(.dina(n30806), .dinb(n30805), .dout(n30807));
  jor  g13545(.dina(n30807), .dinb(n30452), .dout(n30808));
  jxor g13546(.dina(n30446), .dinb(n317), .dout(n30809));
  jand g13547(.dina(n30809), .dinb(n30808), .dout(n30810));
  jor  g13548(.dina(n30810), .dinb(n30447), .dout(n30811));
  jxor g13549(.dina(n30433), .dinb(n284), .dout(n30812));
  jand g13550(.dina(n30812), .dinb(n30811), .dout(n30813));
  jor  g13551(.dina(n30813), .dinb(n30442), .dout(n30814));
  jand g13552(.dina(n30814), .dinb(n30441), .dout(n30815));
  jor  g13553(.dina(n30815), .dinb(n30438), .dout(n30816));
  jand g13554(.dina(n30816), .dinb(n312), .dout(n30817));
  jor  g13555(.dina(n30817), .dinb(n30433), .dout(n30818));
  jnot g13556(.din(n30817), .dout(n30819));
  jxor g13557(.dina(n30812), .dinb(n30811), .dout(n30820));
  jor  g13558(.dina(n30820), .dinb(n30819), .dout(n30821));
  jand g13559(.dina(n30821), .dinb(n30818), .dout(n30822));
  jand g13560(.dina(n30819), .dinb(n30437), .dout(n30823));
  jand g13561(.dina(n30814), .dinb(n30438), .dout(n30824));
  jor  g13562(.dina(n30824), .dinb(n30823), .dout(n30825));
  jand g13563(.dina(n30825), .dinb(n312), .dout(n30826));
  jand g13564(.dina(n30822), .dinb(n285), .dout(n30827));
  jor  g13565(.dina(n30817), .dinb(n30446), .dout(n30828));
  jxor g13566(.dina(n30809), .dinb(n30808), .dout(n30829));
  jor  g13567(.dina(n30829), .dinb(n30819), .dout(n30830));
  jand g13568(.dina(n30830), .dinb(n30828), .dout(n30831));
  jand g13569(.dina(n30831), .dinb(n284), .dout(n30832));
  jor  g13570(.dina(n30817), .dinb(n30451), .dout(n30833));
  jxor g13571(.dina(n30806), .dinb(n30805), .dout(n30834));
  jor  g13572(.dina(n30834), .dinb(n30819), .dout(n30835));
  jand g13573(.dina(n30835), .dinb(n30833), .dout(n30836));
  jand g13574(.dina(n30836), .dinb(n317), .dout(n30837));
  jor  g13575(.dina(n30817), .dinb(n30456), .dout(n30838));
  jxor g13576(.dina(n30803), .dinb(n30802), .dout(n30839));
  jor  g13577(.dina(n30839), .dinb(n30819), .dout(n30840));
  jand g13578(.dina(n30840), .dinb(n30838), .dout(n30841));
  jand g13579(.dina(n30841), .dinb(n316), .dout(n30842));
  jor  g13580(.dina(n30817), .dinb(n30461), .dout(n30843));
  jxor g13581(.dina(n30800), .dinb(n30799), .dout(n30844));
  jor  g13582(.dina(n30844), .dinb(n30819), .dout(n30845));
  jand g13583(.dina(n30845), .dinb(n30843), .dout(n30846));
  jand g13584(.dina(n30846), .dinb(n315), .dout(n30847));
  jor  g13585(.dina(n30817), .dinb(n30466), .dout(n30848));
  jxor g13586(.dina(n30797), .dinb(n30796), .dout(n30849));
  jor  g13587(.dina(n30849), .dinb(n30819), .dout(n30850));
  jand g13588(.dina(n30850), .dinb(n30848), .dout(n30851));
  jand g13589(.dina(n30851), .dinb(n283), .dout(n30852));
  jor  g13590(.dina(n30817), .dinb(n30471), .dout(n30853));
  jxor g13591(.dina(n30794), .dinb(n30793), .dout(n30854));
  jor  g13592(.dina(n30854), .dinb(n30819), .dout(n30855));
  jand g13593(.dina(n30855), .dinb(n30853), .dout(n30856));
  jand g13594(.dina(n30856), .dinb(n280), .dout(n30857));
  jor  g13595(.dina(n30817), .dinb(n30476), .dout(n30858));
  jxor g13596(.dina(n30791), .dinb(n30790), .dout(n30859));
  jor  g13597(.dina(n30859), .dinb(n30819), .dout(n30860));
  jand g13598(.dina(n30860), .dinb(n30858), .dout(n30861));
  jand g13599(.dina(n30861), .dinb(n279), .dout(n30862));
  jor  g13600(.dina(n30817), .dinb(n30481), .dout(n30863));
  jxor g13601(.dina(n30788), .dinb(n30787), .dout(n30864));
  jor  g13602(.dina(n30864), .dinb(n30819), .dout(n30865));
  jand g13603(.dina(n30865), .dinb(n30863), .dout(n30866));
  jand g13604(.dina(n30866), .dinb(n278), .dout(n30867));
  jor  g13605(.dina(n30817), .dinb(n30486), .dout(n30868));
  jxor g13606(.dina(n30785), .dinb(n30784), .dout(n30869));
  jor  g13607(.dina(n30869), .dinb(n30819), .dout(n30870));
  jand g13608(.dina(n30870), .dinb(n30868), .dout(n30871));
  jand g13609(.dina(n30871), .dinb(n277), .dout(n30872));
  jor  g13610(.dina(n30817), .dinb(n30491), .dout(n30873));
  jxor g13611(.dina(n30782), .dinb(n30781), .dout(n30874));
  jor  g13612(.dina(n30874), .dinb(n30819), .dout(n30875));
  jand g13613(.dina(n30875), .dinb(n30873), .dout(n30876));
  jand g13614(.dina(n30876), .dinb(n326), .dout(n30877));
  jor  g13615(.dina(n30817), .dinb(n30496), .dout(n30878));
  jxor g13616(.dina(n30779), .dinb(n30778), .dout(n30879));
  jor  g13617(.dina(n30879), .dinb(n30819), .dout(n30880));
  jand g13618(.dina(n30880), .dinb(n30878), .dout(n30881));
  jand g13619(.dina(n30881), .dinb(n325), .dout(n30882));
  jor  g13620(.dina(n30817), .dinb(n30501), .dout(n30883));
  jxor g13621(.dina(n30776), .dinb(n30775), .dout(n30884));
  jor  g13622(.dina(n30884), .dinb(n30819), .dout(n30885));
  jand g13623(.dina(n30885), .dinb(n30883), .dout(n30886));
  jand g13624(.dina(n30886), .dinb(n324), .dout(n30887));
  jor  g13625(.dina(n30817), .dinb(n30506), .dout(n30888));
  jxor g13626(.dina(n30773), .dinb(n30772), .dout(n30889));
  jor  g13627(.dina(n30889), .dinb(n30819), .dout(n30890));
  jand g13628(.dina(n30890), .dinb(n30888), .dout(n30891));
  jand g13629(.dina(n30891), .dinb(n276), .dout(n30892));
  jor  g13630(.dina(n30817), .dinb(n30511), .dout(n30893));
  jxor g13631(.dina(n30770), .dinb(n30769), .dout(n30894));
  jor  g13632(.dina(n30894), .dinb(n30819), .dout(n30895));
  jand g13633(.dina(n30895), .dinb(n30893), .dout(n30896));
  jand g13634(.dina(n30896), .dinb(n333), .dout(n30897));
  jor  g13635(.dina(n30817), .dinb(n30516), .dout(n30898));
  jxor g13636(.dina(n30767), .dinb(n30766), .dout(n30899));
  jor  g13637(.dina(n30899), .dinb(n30819), .dout(n30900));
  jand g13638(.dina(n30900), .dinb(n30898), .dout(n30901));
  jand g13639(.dina(n30901), .dinb(n332), .dout(n30902));
  jor  g13640(.dina(n30817), .dinb(n30521), .dout(n30903));
  jxor g13641(.dina(n30764), .dinb(n30763), .dout(n30904));
  jor  g13642(.dina(n30904), .dinb(n30819), .dout(n30905));
  jand g13643(.dina(n30905), .dinb(n30903), .dout(n30906));
  jand g13644(.dina(n30906), .dinb(n331), .dout(n30907));
  jor  g13645(.dina(n30817), .dinb(n30526), .dout(n30908));
  jxor g13646(.dina(n30761), .dinb(n30760), .dout(n30909));
  jor  g13647(.dina(n30909), .dinb(n30819), .dout(n30910));
  jand g13648(.dina(n30910), .dinb(n30908), .dout(n30911));
  jand g13649(.dina(n30911), .dinb(n275), .dout(n30912));
  jor  g13650(.dina(n30817), .dinb(n30531), .dout(n30913));
  jxor g13651(.dina(n30758), .dinb(n30757), .dout(n30914));
  jor  g13652(.dina(n30914), .dinb(n30819), .dout(n30915));
  jand g13653(.dina(n30915), .dinb(n30913), .dout(n30916));
  jand g13654(.dina(n30916), .dinb(n340), .dout(n30917));
  jor  g13655(.dina(n30817), .dinb(n30536), .dout(n30918));
  jxor g13656(.dina(n30755), .dinb(n30754), .dout(n30919));
  jor  g13657(.dina(n30919), .dinb(n30819), .dout(n30920));
  jand g13658(.dina(n30920), .dinb(n30918), .dout(n30921));
  jand g13659(.dina(n30921), .dinb(n339), .dout(n30922));
  jor  g13660(.dina(n30817), .dinb(n30541), .dout(n30923));
  jxor g13661(.dina(n30752), .dinb(n30751), .dout(n30924));
  jor  g13662(.dina(n30924), .dinb(n30819), .dout(n30925));
  jand g13663(.dina(n30925), .dinb(n30923), .dout(n30926));
  jand g13664(.dina(n30926), .dinb(n338), .dout(n30927));
  jor  g13665(.dina(n30817), .dinb(n30546), .dout(n30928));
  jxor g13666(.dina(n30749), .dinb(n30748), .dout(n30929));
  jor  g13667(.dina(n30929), .dinb(n30819), .dout(n30930));
  jand g13668(.dina(n30930), .dinb(n30928), .dout(n30931));
  jand g13669(.dina(n30931), .dinb(n271), .dout(n30932));
  jor  g13670(.dina(n30817), .dinb(n30551), .dout(n30933));
  jxor g13671(.dina(n30746), .dinb(n30745), .dout(n30934));
  jor  g13672(.dina(n30934), .dinb(n30819), .dout(n30935));
  jand g13673(.dina(n30935), .dinb(n30933), .dout(n30936));
  jand g13674(.dina(n30936), .dinb(n270), .dout(n30937));
  jor  g13675(.dina(n30817), .dinb(n30556), .dout(n30938));
  jxor g13676(.dina(n30743), .dinb(n30742), .dout(n30939));
  jor  g13677(.dina(n30939), .dinb(n30819), .dout(n30940));
  jand g13678(.dina(n30940), .dinb(n30938), .dout(n30941));
  jand g13679(.dina(n30941), .dinb(n269), .dout(n30942));
  jor  g13680(.dina(n30817), .dinb(n30561), .dout(n30943));
  jxor g13681(.dina(n30740), .dinb(n30739), .dout(n30944));
  jor  g13682(.dina(n30944), .dinb(n30819), .dout(n30945));
  jand g13683(.dina(n30945), .dinb(n30943), .dout(n30946));
  jand g13684(.dina(n30946), .dinb(n274), .dout(n30947));
  jor  g13685(.dina(n30817), .dinb(n30566), .dout(n30948));
  jxor g13686(.dina(n30737), .dinb(n30736), .dout(n30949));
  jor  g13687(.dina(n30949), .dinb(n30819), .dout(n30950));
  jand g13688(.dina(n30950), .dinb(n30948), .dout(n30951));
  jand g13689(.dina(n30951), .dinb(n268), .dout(n30952));
  jor  g13690(.dina(n30817), .dinb(n30571), .dout(n30953));
  jxor g13691(.dina(n30734), .dinb(n30733), .dout(n30954));
  jor  g13692(.dina(n30954), .dinb(n30819), .dout(n30955));
  jand g13693(.dina(n30955), .dinb(n30953), .dout(n30956));
  jand g13694(.dina(n30956), .dinb(n349), .dout(n30957));
  jor  g13695(.dina(n30817), .dinb(n30576), .dout(n30958));
  jxor g13696(.dina(n30731), .dinb(n30730), .dout(n30959));
  jor  g13697(.dina(n30959), .dinb(n30819), .dout(n30960));
  jand g13698(.dina(n30960), .dinb(n30958), .dout(n30961));
  jand g13699(.dina(n30961), .dinb(n348), .dout(n30962));
  jor  g13700(.dina(n30817), .dinb(n30581), .dout(n30963));
  jxor g13701(.dina(n30728), .dinb(n30727), .dout(n30964));
  jor  g13702(.dina(n30964), .dinb(n30819), .dout(n30965));
  jand g13703(.dina(n30965), .dinb(n30963), .dout(n30966));
  jand g13704(.dina(n30966), .dinb(n347), .dout(n30967));
  jor  g13705(.dina(n30817), .dinb(n30586), .dout(n30968));
  jxor g13706(.dina(n30725), .dinb(n30724), .dout(n30969));
  jor  g13707(.dina(n30969), .dinb(n30819), .dout(n30970));
  jand g13708(.dina(n30970), .dinb(n30968), .dout(n30971));
  jand g13709(.dina(n30971), .dinb(n267), .dout(n30972));
  jor  g13710(.dina(n30817), .dinb(n30591), .dout(n30973));
  jxor g13711(.dina(n30722), .dinb(n30721), .dout(n30974));
  jor  g13712(.dina(n30974), .dinb(n30819), .dout(n30975));
  jand g13713(.dina(n30975), .dinb(n30973), .dout(n30976));
  jand g13714(.dina(n30976), .dinb(n266), .dout(n30977));
  jor  g13715(.dina(n30817), .dinb(n30596), .dout(n30978));
  jxor g13716(.dina(n30719), .dinb(n30718), .dout(n30979));
  jor  g13717(.dina(n30979), .dinb(n30819), .dout(n30980));
  jand g13718(.dina(n30980), .dinb(n30978), .dout(n30981));
  jand g13719(.dina(n30981), .dinb(n356), .dout(n30982));
  jor  g13720(.dina(n30817), .dinb(n30601), .dout(n30983));
  jxor g13721(.dina(n30716), .dinb(n30715), .dout(n30984));
  jor  g13722(.dina(n30984), .dinb(n30819), .dout(n30985));
  jand g13723(.dina(n30985), .dinb(n30983), .dout(n30986));
  jand g13724(.dina(n30986), .dinb(n355), .dout(n30987));
  jor  g13725(.dina(n30817), .dinb(n30606), .dout(n30988));
  jxor g13726(.dina(n30713), .dinb(n30712), .dout(n30989));
  jor  g13727(.dina(n30989), .dinb(n30819), .dout(n30990));
  jand g13728(.dina(n30990), .dinb(n30988), .dout(n30991));
  jand g13729(.dina(n30991), .dinb(n364), .dout(n30992));
  jor  g13730(.dina(n30817), .dinb(n30611), .dout(n30993));
  jxor g13731(.dina(n30710), .dinb(n30709), .dout(n30994));
  jor  g13732(.dina(n30994), .dinb(n30819), .dout(n30995));
  jand g13733(.dina(n30995), .dinb(n30993), .dout(n30996));
  jand g13734(.dina(n30996), .dinb(n361), .dout(n30997));
  jor  g13735(.dina(n30817), .dinb(n30616), .dout(n30998));
  jxor g13736(.dina(n30707), .dinb(n30706), .dout(n30999));
  jor  g13737(.dina(n30999), .dinb(n30819), .dout(n31000));
  jand g13738(.dina(n31000), .dinb(n30998), .dout(n31001));
  jand g13739(.dina(n31001), .dinb(n360), .dout(n31002));
  jor  g13740(.dina(n30817), .dinb(n30621), .dout(n31003));
  jxor g13741(.dina(n30704), .dinb(n30703), .dout(n31004));
  jor  g13742(.dina(n31004), .dinb(n30819), .dout(n31005));
  jand g13743(.dina(n31005), .dinb(n31003), .dout(n31006));
  jand g13744(.dina(n31006), .dinb(n363), .dout(n31007));
  jor  g13745(.dina(n30817), .dinb(n30626), .dout(n31008));
  jxor g13746(.dina(n30701), .dinb(n30700), .dout(n31009));
  jor  g13747(.dina(n31009), .dinb(n30819), .dout(n31010));
  jand g13748(.dina(n31010), .dinb(n31008), .dout(n31011));
  jand g13749(.dina(n31011), .dinb(n359), .dout(n31012));
  jor  g13750(.dina(n30817), .dinb(n30631), .dout(n31013));
  jxor g13751(.dina(n30698), .dinb(n30697), .dout(n31014));
  jor  g13752(.dina(n31014), .dinb(n30819), .dout(n31015));
  jand g13753(.dina(n31015), .dinb(n31013), .dout(n31016));
  jand g13754(.dina(n31016), .dinb(n369), .dout(n31017));
  jor  g13755(.dina(n30817), .dinb(n30636), .dout(n31018));
  jxor g13756(.dina(n30695), .dinb(n30694), .dout(n31019));
  jor  g13757(.dina(n31019), .dinb(n30819), .dout(n31020));
  jand g13758(.dina(n31020), .dinb(n31018), .dout(n31021));
  jand g13759(.dina(n31021), .dinb(n368), .dout(n31022));
  jor  g13760(.dina(n30817), .dinb(n30641), .dout(n31023));
  jxor g13761(.dina(n30692), .dinb(n30691), .dout(n31024));
  jor  g13762(.dina(n31024), .dinb(n30819), .dout(n31025));
  jand g13763(.dina(n31025), .dinb(n31023), .dout(n31026));
  jand g13764(.dina(n31026), .dinb(n367), .dout(n31027));
  jor  g13765(.dina(n30817), .dinb(n30646), .dout(n31028));
  jxor g13766(.dina(n30689), .dinb(n30688), .dout(n31029));
  jor  g13767(.dina(n31029), .dinb(n30819), .dout(n31030));
  jand g13768(.dina(n31030), .dinb(n31028), .dout(n31031));
  jand g13769(.dina(n31031), .dinb(n265), .dout(n31032));
  jor  g13770(.dina(n30817), .dinb(n30651), .dout(n31033));
  jxor g13771(.dina(n30686), .dinb(n30685), .dout(n31034));
  jor  g13772(.dina(n31034), .dinb(n30819), .dout(n31035));
  jand g13773(.dina(n31035), .dinb(n31033), .dout(n31036));
  jand g13774(.dina(n31036), .dinb(n378), .dout(n31037));
  jor  g13775(.dina(n30817), .dinb(n30656), .dout(n31038));
  jxor g13776(.dina(n30683), .dinb(n30682), .dout(n31039));
  jor  g13777(.dina(n31039), .dinb(n30819), .dout(n31040));
  jand g13778(.dina(n31040), .dinb(n31038), .dout(n31041));
  jand g13779(.dina(n31041), .dinb(n377), .dout(n31042));
  jor  g13780(.dina(n30817), .dinb(n30661), .dout(n31043));
  jxor g13781(.dina(n30680), .dinb(n30679), .dout(n31044));
  jor  g13782(.dina(n31044), .dinb(n30819), .dout(n31045));
  jand g13783(.dina(n31045), .dinb(n31043), .dout(n31046));
  jand g13784(.dina(n31046), .dinb(n376), .dout(n31047));
  jor  g13785(.dina(n30817), .dinb(n30668), .dout(n31048));
  jxor g13786(.dina(n30677), .dinb(n30676), .dout(n31049));
  jor  g13787(.dina(n31049), .dinb(n30819), .dout(n31050));
  jand g13788(.dina(n31050), .dinb(n31048), .dout(n31051));
  jand g13789(.dina(n31051), .dinb(n264), .dout(n31052));
  jor  g13790(.dina(n30817), .dinb(n30673), .dout(n31053));
  jxor g13791(.dina(n30674), .dinb(n10799), .dout(n31054));
  jand g13792(.dina(n31054), .dinb(n30817), .dout(n31055));
  jnot g13793(.din(n31055), .dout(n31056));
  jand g13794(.dina(n31056), .dinb(n31053), .dout(n31057));
  jnot g13795(.din(n31057), .dout(n31058));
  jand g13796(.dina(n31058), .dinb(n386), .dout(n31059));
  jnot g13797(.din(n11186), .dout(n31060));
  jnot g13798(.din(n30438), .dout(n31061));
  jnot g13799(.din(n30442), .dout(n31062));
  jnot g13800(.din(n30447), .dout(n31063));
  jnot g13801(.din(n30452), .dout(n31064));
  jnot g13802(.din(n30457), .dout(n31065));
  jnot g13803(.din(n30462), .dout(n31066));
  jnot g13804(.din(n30467), .dout(n31067));
  jnot g13805(.din(n30472), .dout(n31068));
  jnot g13806(.din(n30477), .dout(n31069));
  jnot g13807(.din(n30482), .dout(n31070));
  jnot g13808(.din(n30487), .dout(n31071));
  jnot g13809(.din(n30492), .dout(n31072));
  jnot g13810(.din(n30497), .dout(n31073));
  jnot g13811(.din(n30502), .dout(n31074));
  jnot g13812(.din(n30507), .dout(n31075));
  jnot g13813(.din(n30512), .dout(n31076));
  jnot g13814(.din(n30517), .dout(n31077));
  jnot g13815(.din(n30522), .dout(n31078));
  jnot g13816(.din(n30527), .dout(n31079));
  jnot g13817(.din(n30532), .dout(n31080));
  jnot g13818(.din(n30537), .dout(n31081));
  jnot g13819(.din(n30542), .dout(n31082));
  jnot g13820(.din(n30547), .dout(n31083));
  jnot g13821(.din(n30552), .dout(n31084));
  jnot g13822(.din(n30557), .dout(n31085));
  jnot g13823(.din(n30562), .dout(n31086));
  jnot g13824(.din(n30567), .dout(n31087));
  jnot g13825(.din(n30572), .dout(n31088));
  jnot g13826(.din(n30577), .dout(n31089));
  jnot g13827(.din(n30582), .dout(n31090));
  jnot g13828(.din(n30587), .dout(n31091));
  jnot g13829(.din(n30592), .dout(n31092));
  jnot g13830(.din(n30597), .dout(n31093));
  jnot g13831(.din(n30602), .dout(n31094));
  jnot g13832(.din(n30607), .dout(n31095));
  jnot g13833(.din(n30612), .dout(n31096));
  jnot g13834(.din(n30617), .dout(n31097));
  jnot g13835(.din(n30622), .dout(n31098));
  jnot g13836(.din(n30627), .dout(n31099));
  jnot g13837(.din(n30632), .dout(n31100));
  jnot g13838(.din(n30637), .dout(n31101));
  jnot g13839(.din(n30642), .dout(n31102));
  jnot g13840(.din(n30647), .dout(n31103));
  jnot g13841(.din(n30652), .dout(n31104));
  jnot g13842(.din(n30657), .dout(n31105));
  jnot g13843(.din(n30662), .dout(n31106));
  jnot g13844(.din(n30669), .dout(n31107));
  jnot g13845(.din(n30672), .dout(n31108));
  jxor g13846(.dina(n30673), .dinb(n259), .dout(n31109));
  jor  g13847(.dina(n31109), .dinb(n10798), .dout(n31110));
  jand g13848(.dina(n31110), .dinb(n31108), .dout(n31111));
  jnot g13849(.din(n30677), .dout(n31112));
  jor  g13850(.dina(n31112), .dinb(n31111), .dout(n31113));
  jand g13851(.dina(n31113), .dinb(n31107), .dout(n31114));
  jnot g13852(.din(n30680), .dout(n31115));
  jor  g13853(.dina(n31115), .dinb(n31114), .dout(n31116));
  jand g13854(.dina(n31116), .dinb(n31106), .dout(n31117));
  jnot g13855(.din(n30683), .dout(n31118));
  jor  g13856(.dina(n31118), .dinb(n31117), .dout(n31119));
  jand g13857(.dina(n31119), .dinb(n31105), .dout(n31120));
  jnot g13858(.din(n30686), .dout(n31121));
  jor  g13859(.dina(n31121), .dinb(n31120), .dout(n31122));
  jand g13860(.dina(n31122), .dinb(n31104), .dout(n31123));
  jnot g13861(.din(n30689), .dout(n31124));
  jor  g13862(.dina(n31124), .dinb(n31123), .dout(n31125));
  jand g13863(.dina(n31125), .dinb(n31103), .dout(n31126));
  jnot g13864(.din(n30692), .dout(n31127));
  jor  g13865(.dina(n31127), .dinb(n31126), .dout(n31128));
  jand g13866(.dina(n31128), .dinb(n31102), .dout(n31129));
  jnot g13867(.din(n30695), .dout(n31130));
  jor  g13868(.dina(n31130), .dinb(n31129), .dout(n31131));
  jand g13869(.dina(n31131), .dinb(n31101), .dout(n31132));
  jnot g13870(.din(n30698), .dout(n31133));
  jor  g13871(.dina(n31133), .dinb(n31132), .dout(n31134));
  jand g13872(.dina(n31134), .dinb(n31100), .dout(n31135));
  jnot g13873(.din(n30701), .dout(n31136));
  jor  g13874(.dina(n31136), .dinb(n31135), .dout(n31137));
  jand g13875(.dina(n31137), .dinb(n31099), .dout(n31138));
  jnot g13876(.din(n30704), .dout(n31139));
  jor  g13877(.dina(n31139), .dinb(n31138), .dout(n31140));
  jand g13878(.dina(n31140), .dinb(n31098), .dout(n31141));
  jnot g13879(.din(n30707), .dout(n31142));
  jor  g13880(.dina(n31142), .dinb(n31141), .dout(n31143));
  jand g13881(.dina(n31143), .dinb(n31097), .dout(n31144));
  jnot g13882(.din(n30710), .dout(n31145));
  jor  g13883(.dina(n31145), .dinb(n31144), .dout(n31146));
  jand g13884(.dina(n31146), .dinb(n31096), .dout(n31147));
  jnot g13885(.din(n30713), .dout(n31148));
  jor  g13886(.dina(n31148), .dinb(n31147), .dout(n31149));
  jand g13887(.dina(n31149), .dinb(n31095), .dout(n31150));
  jnot g13888(.din(n30716), .dout(n31151));
  jor  g13889(.dina(n31151), .dinb(n31150), .dout(n31152));
  jand g13890(.dina(n31152), .dinb(n31094), .dout(n31153));
  jnot g13891(.din(n30719), .dout(n31154));
  jor  g13892(.dina(n31154), .dinb(n31153), .dout(n31155));
  jand g13893(.dina(n31155), .dinb(n31093), .dout(n31156));
  jnot g13894(.din(n30722), .dout(n31157));
  jor  g13895(.dina(n31157), .dinb(n31156), .dout(n31158));
  jand g13896(.dina(n31158), .dinb(n31092), .dout(n31159));
  jnot g13897(.din(n30725), .dout(n31160));
  jor  g13898(.dina(n31160), .dinb(n31159), .dout(n31161));
  jand g13899(.dina(n31161), .dinb(n31091), .dout(n31162));
  jnot g13900(.din(n30728), .dout(n31163));
  jor  g13901(.dina(n31163), .dinb(n31162), .dout(n31164));
  jand g13902(.dina(n31164), .dinb(n31090), .dout(n31165));
  jnot g13903(.din(n30731), .dout(n31166));
  jor  g13904(.dina(n31166), .dinb(n31165), .dout(n31167));
  jand g13905(.dina(n31167), .dinb(n31089), .dout(n31168));
  jnot g13906(.din(n30734), .dout(n31169));
  jor  g13907(.dina(n31169), .dinb(n31168), .dout(n31170));
  jand g13908(.dina(n31170), .dinb(n31088), .dout(n31171));
  jnot g13909(.din(n30737), .dout(n31172));
  jor  g13910(.dina(n31172), .dinb(n31171), .dout(n31173));
  jand g13911(.dina(n31173), .dinb(n31087), .dout(n31174));
  jnot g13912(.din(n30740), .dout(n31175));
  jor  g13913(.dina(n31175), .dinb(n31174), .dout(n31176));
  jand g13914(.dina(n31176), .dinb(n31086), .dout(n31177));
  jnot g13915(.din(n30743), .dout(n31178));
  jor  g13916(.dina(n31178), .dinb(n31177), .dout(n31179));
  jand g13917(.dina(n31179), .dinb(n31085), .dout(n31180));
  jnot g13918(.din(n30746), .dout(n31181));
  jor  g13919(.dina(n31181), .dinb(n31180), .dout(n31182));
  jand g13920(.dina(n31182), .dinb(n31084), .dout(n31183));
  jnot g13921(.din(n30749), .dout(n31184));
  jor  g13922(.dina(n31184), .dinb(n31183), .dout(n31185));
  jand g13923(.dina(n31185), .dinb(n31083), .dout(n31186));
  jnot g13924(.din(n30752), .dout(n31187));
  jor  g13925(.dina(n31187), .dinb(n31186), .dout(n31188));
  jand g13926(.dina(n31188), .dinb(n31082), .dout(n31189));
  jnot g13927(.din(n30755), .dout(n31190));
  jor  g13928(.dina(n31190), .dinb(n31189), .dout(n31191));
  jand g13929(.dina(n31191), .dinb(n31081), .dout(n31192));
  jnot g13930(.din(n30758), .dout(n31193));
  jor  g13931(.dina(n31193), .dinb(n31192), .dout(n31194));
  jand g13932(.dina(n31194), .dinb(n31080), .dout(n31195));
  jnot g13933(.din(n30761), .dout(n31196));
  jor  g13934(.dina(n31196), .dinb(n31195), .dout(n31197));
  jand g13935(.dina(n31197), .dinb(n31079), .dout(n31198));
  jnot g13936(.din(n30764), .dout(n31199));
  jor  g13937(.dina(n31199), .dinb(n31198), .dout(n31200));
  jand g13938(.dina(n31200), .dinb(n31078), .dout(n31201));
  jnot g13939(.din(n30767), .dout(n31202));
  jor  g13940(.dina(n31202), .dinb(n31201), .dout(n31203));
  jand g13941(.dina(n31203), .dinb(n31077), .dout(n31204));
  jnot g13942(.din(n30770), .dout(n31205));
  jor  g13943(.dina(n31205), .dinb(n31204), .dout(n31206));
  jand g13944(.dina(n31206), .dinb(n31076), .dout(n31207));
  jnot g13945(.din(n30773), .dout(n31208));
  jor  g13946(.dina(n31208), .dinb(n31207), .dout(n31209));
  jand g13947(.dina(n31209), .dinb(n31075), .dout(n31210));
  jnot g13948(.din(n30776), .dout(n31211));
  jor  g13949(.dina(n31211), .dinb(n31210), .dout(n31212));
  jand g13950(.dina(n31212), .dinb(n31074), .dout(n31213));
  jnot g13951(.din(n30779), .dout(n31214));
  jor  g13952(.dina(n31214), .dinb(n31213), .dout(n31215));
  jand g13953(.dina(n31215), .dinb(n31073), .dout(n31216));
  jnot g13954(.din(n30782), .dout(n31217));
  jor  g13955(.dina(n31217), .dinb(n31216), .dout(n31218));
  jand g13956(.dina(n31218), .dinb(n31072), .dout(n31219));
  jnot g13957(.din(n30785), .dout(n31220));
  jor  g13958(.dina(n31220), .dinb(n31219), .dout(n31221));
  jand g13959(.dina(n31221), .dinb(n31071), .dout(n31222));
  jnot g13960(.din(n30788), .dout(n31223));
  jor  g13961(.dina(n31223), .dinb(n31222), .dout(n31224));
  jand g13962(.dina(n31224), .dinb(n31070), .dout(n31225));
  jnot g13963(.din(n30791), .dout(n31226));
  jor  g13964(.dina(n31226), .dinb(n31225), .dout(n31227));
  jand g13965(.dina(n31227), .dinb(n31069), .dout(n31228));
  jnot g13966(.din(n30794), .dout(n31229));
  jor  g13967(.dina(n31229), .dinb(n31228), .dout(n31230));
  jand g13968(.dina(n31230), .dinb(n31068), .dout(n31231));
  jnot g13969(.din(n30797), .dout(n31232));
  jor  g13970(.dina(n31232), .dinb(n31231), .dout(n31233));
  jand g13971(.dina(n31233), .dinb(n31067), .dout(n31234));
  jnot g13972(.din(n30800), .dout(n31235));
  jor  g13973(.dina(n31235), .dinb(n31234), .dout(n31236));
  jand g13974(.dina(n31236), .dinb(n31066), .dout(n31237));
  jnot g13975(.din(n30803), .dout(n31238));
  jor  g13976(.dina(n31238), .dinb(n31237), .dout(n31239));
  jand g13977(.dina(n31239), .dinb(n31065), .dout(n31240));
  jnot g13978(.din(n30806), .dout(n31241));
  jor  g13979(.dina(n31241), .dinb(n31240), .dout(n31242));
  jand g13980(.dina(n31242), .dinb(n31064), .dout(n31243));
  jnot g13981(.din(n30809), .dout(n31244));
  jor  g13982(.dina(n31244), .dinb(n31243), .dout(n31245));
  jand g13983(.dina(n31245), .dinb(n31063), .dout(n31246));
  jnot g13984(.din(n30812), .dout(n31247));
  jor  g13985(.dina(n31247), .dinb(n31246), .dout(n31248));
  jand g13986(.dina(n31248), .dinb(n31062), .dout(n31249));
  jor  g13987(.dina(n31249), .dinb(n30440), .dout(n31250));
  jand g13988(.dina(n31250), .dinb(n31061), .dout(n31251));
  jor  g13989(.dina(n31251), .dinb(n31060), .dout(n31252));
  jand g13990(.dina(n31252), .dinb(a15 ), .dout(n31253));
  jnot g13991(.din(n11189), .dout(n31254));
  jor  g13992(.dina(n31251), .dinb(n31254), .dout(n31255));
  jnot g13993(.din(n31255), .dout(n31256));
  jor  g13994(.dina(n31256), .dinb(n31253), .dout(n31257));
  jand g13995(.dina(n31257), .dinb(n259), .dout(n31258));
  jand g13996(.dina(n30816), .dinb(n11186), .dout(n31259));
  jor  g13997(.dina(n31259), .dinb(n10797), .dout(n31260));
  jand g13998(.dina(n31255), .dinb(n31260), .dout(n31261));
  jxor g13999(.dina(n31261), .dinb(b1 ), .dout(n31262));
  jand g14000(.dina(n31262), .dinb(n11197), .dout(n31263));
  jor  g14001(.dina(n31263), .dinb(n31258), .dout(n31264));
  jxor g14002(.dina(n31057), .dinb(b2 ), .dout(n31265));
  jand g14003(.dina(n31265), .dinb(n31264), .dout(n31266));
  jor  g14004(.dina(n31266), .dinb(n31059), .dout(n31267));
  jxor g14005(.dina(n31051), .dinb(n264), .dout(n31268));
  jand g14006(.dina(n31268), .dinb(n31267), .dout(n31269));
  jor  g14007(.dina(n31269), .dinb(n31052), .dout(n31270));
  jxor g14008(.dina(n31046), .dinb(n376), .dout(n31271));
  jand g14009(.dina(n31271), .dinb(n31270), .dout(n31272));
  jor  g14010(.dina(n31272), .dinb(n31047), .dout(n31273));
  jxor g14011(.dina(n31041), .dinb(n377), .dout(n31274));
  jand g14012(.dina(n31274), .dinb(n31273), .dout(n31275));
  jor  g14013(.dina(n31275), .dinb(n31042), .dout(n31276));
  jxor g14014(.dina(n31036), .dinb(n378), .dout(n31277));
  jand g14015(.dina(n31277), .dinb(n31276), .dout(n31278));
  jor  g14016(.dina(n31278), .dinb(n31037), .dout(n31279));
  jxor g14017(.dina(n31031), .dinb(n265), .dout(n31280));
  jand g14018(.dina(n31280), .dinb(n31279), .dout(n31281));
  jor  g14019(.dina(n31281), .dinb(n31032), .dout(n31282));
  jxor g14020(.dina(n31026), .dinb(n367), .dout(n31283));
  jand g14021(.dina(n31283), .dinb(n31282), .dout(n31284));
  jor  g14022(.dina(n31284), .dinb(n31027), .dout(n31285));
  jxor g14023(.dina(n31021), .dinb(n368), .dout(n31286));
  jand g14024(.dina(n31286), .dinb(n31285), .dout(n31287));
  jor  g14025(.dina(n31287), .dinb(n31022), .dout(n31288));
  jxor g14026(.dina(n31016), .dinb(n369), .dout(n31289));
  jand g14027(.dina(n31289), .dinb(n31288), .dout(n31290));
  jor  g14028(.dina(n31290), .dinb(n31017), .dout(n31291));
  jxor g14029(.dina(n31011), .dinb(n359), .dout(n31292));
  jand g14030(.dina(n31292), .dinb(n31291), .dout(n31293));
  jor  g14031(.dina(n31293), .dinb(n31012), .dout(n31294));
  jxor g14032(.dina(n31006), .dinb(n363), .dout(n31295));
  jand g14033(.dina(n31295), .dinb(n31294), .dout(n31296));
  jor  g14034(.dina(n31296), .dinb(n31007), .dout(n31297));
  jxor g14035(.dina(n31001), .dinb(n360), .dout(n31298));
  jand g14036(.dina(n31298), .dinb(n31297), .dout(n31299));
  jor  g14037(.dina(n31299), .dinb(n31002), .dout(n31300));
  jxor g14038(.dina(n30996), .dinb(n361), .dout(n31301));
  jand g14039(.dina(n31301), .dinb(n31300), .dout(n31302));
  jor  g14040(.dina(n31302), .dinb(n30997), .dout(n31303));
  jxor g14041(.dina(n30991), .dinb(n364), .dout(n31304));
  jand g14042(.dina(n31304), .dinb(n31303), .dout(n31305));
  jor  g14043(.dina(n31305), .dinb(n30992), .dout(n31306));
  jxor g14044(.dina(n30986), .dinb(n355), .dout(n31307));
  jand g14045(.dina(n31307), .dinb(n31306), .dout(n31308));
  jor  g14046(.dina(n31308), .dinb(n30987), .dout(n31309));
  jxor g14047(.dina(n30981), .dinb(n356), .dout(n31310));
  jand g14048(.dina(n31310), .dinb(n31309), .dout(n31311));
  jor  g14049(.dina(n31311), .dinb(n30982), .dout(n31312));
  jxor g14050(.dina(n30976), .dinb(n266), .dout(n31313));
  jand g14051(.dina(n31313), .dinb(n31312), .dout(n31314));
  jor  g14052(.dina(n31314), .dinb(n30977), .dout(n31315));
  jxor g14053(.dina(n30971), .dinb(n267), .dout(n31316));
  jand g14054(.dina(n31316), .dinb(n31315), .dout(n31317));
  jor  g14055(.dina(n31317), .dinb(n30972), .dout(n31318));
  jxor g14056(.dina(n30966), .dinb(n347), .dout(n31319));
  jand g14057(.dina(n31319), .dinb(n31318), .dout(n31320));
  jor  g14058(.dina(n31320), .dinb(n30967), .dout(n31321));
  jxor g14059(.dina(n30961), .dinb(n348), .dout(n31322));
  jand g14060(.dina(n31322), .dinb(n31321), .dout(n31323));
  jor  g14061(.dina(n31323), .dinb(n30962), .dout(n31324));
  jxor g14062(.dina(n30956), .dinb(n349), .dout(n31325));
  jand g14063(.dina(n31325), .dinb(n31324), .dout(n31326));
  jor  g14064(.dina(n31326), .dinb(n30957), .dout(n31327));
  jxor g14065(.dina(n30951), .dinb(n268), .dout(n31328));
  jand g14066(.dina(n31328), .dinb(n31327), .dout(n31329));
  jor  g14067(.dina(n31329), .dinb(n30952), .dout(n31330));
  jxor g14068(.dina(n30946), .dinb(n274), .dout(n31331));
  jand g14069(.dina(n31331), .dinb(n31330), .dout(n31332));
  jor  g14070(.dina(n31332), .dinb(n30947), .dout(n31333));
  jxor g14071(.dina(n30941), .dinb(n269), .dout(n31334));
  jand g14072(.dina(n31334), .dinb(n31333), .dout(n31335));
  jor  g14073(.dina(n31335), .dinb(n30942), .dout(n31336));
  jxor g14074(.dina(n30936), .dinb(n270), .dout(n31337));
  jand g14075(.dina(n31337), .dinb(n31336), .dout(n31338));
  jor  g14076(.dina(n31338), .dinb(n30937), .dout(n31339));
  jxor g14077(.dina(n30931), .dinb(n271), .dout(n31340));
  jand g14078(.dina(n31340), .dinb(n31339), .dout(n31341));
  jor  g14079(.dina(n31341), .dinb(n30932), .dout(n31342));
  jxor g14080(.dina(n30926), .dinb(n338), .dout(n31343));
  jand g14081(.dina(n31343), .dinb(n31342), .dout(n31344));
  jor  g14082(.dina(n31344), .dinb(n30927), .dout(n31345));
  jxor g14083(.dina(n30921), .dinb(n339), .dout(n31346));
  jand g14084(.dina(n31346), .dinb(n31345), .dout(n31347));
  jor  g14085(.dina(n31347), .dinb(n30922), .dout(n31348));
  jxor g14086(.dina(n30916), .dinb(n340), .dout(n31349));
  jand g14087(.dina(n31349), .dinb(n31348), .dout(n31350));
  jor  g14088(.dina(n31350), .dinb(n30917), .dout(n31351));
  jxor g14089(.dina(n30911), .dinb(n275), .dout(n31352));
  jand g14090(.dina(n31352), .dinb(n31351), .dout(n31353));
  jor  g14091(.dina(n31353), .dinb(n30912), .dout(n31354));
  jxor g14092(.dina(n30906), .dinb(n331), .dout(n31355));
  jand g14093(.dina(n31355), .dinb(n31354), .dout(n31356));
  jor  g14094(.dina(n31356), .dinb(n30907), .dout(n31357));
  jxor g14095(.dina(n30901), .dinb(n332), .dout(n31358));
  jand g14096(.dina(n31358), .dinb(n31357), .dout(n31359));
  jor  g14097(.dina(n31359), .dinb(n30902), .dout(n31360));
  jxor g14098(.dina(n30896), .dinb(n333), .dout(n31361));
  jand g14099(.dina(n31361), .dinb(n31360), .dout(n31362));
  jor  g14100(.dina(n31362), .dinb(n30897), .dout(n31363));
  jxor g14101(.dina(n30891), .dinb(n276), .dout(n31364));
  jand g14102(.dina(n31364), .dinb(n31363), .dout(n31365));
  jor  g14103(.dina(n31365), .dinb(n30892), .dout(n31366));
  jxor g14104(.dina(n30886), .dinb(n324), .dout(n31367));
  jand g14105(.dina(n31367), .dinb(n31366), .dout(n31368));
  jor  g14106(.dina(n31368), .dinb(n30887), .dout(n31369));
  jxor g14107(.dina(n30881), .dinb(n325), .dout(n31370));
  jand g14108(.dina(n31370), .dinb(n31369), .dout(n31371));
  jor  g14109(.dina(n31371), .dinb(n30882), .dout(n31372));
  jxor g14110(.dina(n30876), .dinb(n326), .dout(n31373));
  jand g14111(.dina(n31373), .dinb(n31372), .dout(n31374));
  jor  g14112(.dina(n31374), .dinb(n30877), .dout(n31375));
  jxor g14113(.dina(n30871), .dinb(n277), .dout(n31376));
  jand g14114(.dina(n31376), .dinb(n31375), .dout(n31377));
  jor  g14115(.dina(n31377), .dinb(n30872), .dout(n31378));
  jxor g14116(.dina(n30866), .dinb(n278), .dout(n31379));
  jand g14117(.dina(n31379), .dinb(n31378), .dout(n31380));
  jor  g14118(.dina(n31380), .dinb(n30867), .dout(n31381));
  jxor g14119(.dina(n30861), .dinb(n279), .dout(n31382));
  jand g14120(.dina(n31382), .dinb(n31381), .dout(n31383));
  jor  g14121(.dina(n31383), .dinb(n30862), .dout(n31384));
  jxor g14122(.dina(n30856), .dinb(n280), .dout(n31385));
  jand g14123(.dina(n31385), .dinb(n31384), .dout(n31386));
  jor  g14124(.dina(n31386), .dinb(n30857), .dout(n31387));
  jxor g14125(.dina(n30851), .dinb(n283), .dout(n31388));
  jand g14126(.dina(n31388), .dinb(n31387), .dout(n31389));
  jor  g14127(.dina(n31389), .dinb(n30852), .dout(n31390));
  jxor g14128(.dina(n30846), .dinb(n315), .dout(n31391));
  jand g14129(.dina(n31391), .dinb(n31390), .dout(n31392));
  jor  g14130(.dina(n31392), .dinb(n30847), .dout(n31393));
  jxor g14131(.dina(n30841), .dinb(n316), .dout(n31394));
  jand g14132(.dina(n31394), .dinb(n31393), .dout(n31395));
  jor  g14133(.dina(n31395), .dinb(n30842), .dout(n31396));
  jxor g14134(.dina(n30836), .dinb(n317), .dout(n31397));
  jand g14135(.dina(n31397), .dinb(n31396), .dout(n31398));
  jor  g14136(.dina(n31398), .dinb(n30837), .dout(n31399));
  jxor g14137(.dina(n30831), .dinb(n284), .dout(n31400));
  jand g14138(.dina(n31400), .dinb(n31399), .dout(n31401));
  jor  g14139(.dina(n31401), .dinb(n30832), .dout(n31402));
  jxor g14140(.dina(n30822), .dinb(n285), .dout(n31403));
  jand g14141(.dina(n31403), .dinb(n31402), .dout(n31404));
  jor  g14142(.dina(n31404), .dinb(n30827), .dout(n31405));
  jxor g14143(.dina(n30825), .dinb(b49 ), .dout(n31406));
  jnot g14144(.din(n31406), .dout(n31407));
  jand g14145(.dina(n31407), .dinb(n31405), .dout(n31408));
  jand g14146(.dina(n31408), .dinb(n311), .dout(n31409));
  jor  g14147(.dina(n31409), .dinb(n30826), .dout(n31410));
  jor  g14148(.dina(n31410), .dinb(n30822), .dout(n31411));
  jnot g14149(.din(n31410), .dout(n31412));
  jxor g14150(.dina(n31403), .dinb(n31402), .dout(n31413));
  jor  g14151(.dina(n31413), .dinb(n31412), .dout(n31414));
  jand g14152(.dina(n31414), .dinb(n31411), .dout(n31415));
  jand g14153(.dina(n31405), .dinb(n30826), .dout(n31416));
  jnot g14154(.din(n31409), .dout(n31417));
  jand g14155(.dina(n31417), .dinb(n30437), .dout(n31418));
  jand g14156(.dina(n31418), .dinb(n843), .dout(n31419));
  jor  g14157(.dina(n31419), .dinb(n31416), .dout(n31420));
  jand g14158(.dina(n31420), .dinb(n287), .dout(n31421));
  jnot g14159(.din(n31420), .dout(n31422));
  jand g14160(.dina(n31422), .dinb(b50 ), .dout(n31423));
  jnot g14161(.din(n31423), .dout(n31424));
  jand g14162(.dina(n31415), .dinb(n286), .dout(n31425));
  jor  g14163(.dina(n31410), .dinb(n30831), .dout(n31426));
  jxor g14164(.dina(n31400), .dinb(n31399), .dout(n31427));
  jor  g14165(.dina(n31427), .dinb(n31412), .dout(n31428));
  jand g14166(.dina(n31428), .dinb(n31426), .dout(n31429));
  jand g14167(.dina(n31429), .dinb(n285), .dout(n31430));
  jor  g14168(.dina(n31410), .dinb(n30836), .dout(n31431));
  jxor g14169(.dina(n31397), .dinb(n31396), .dout(n31432));
  jor  g14170(.dina(n31432), .dinb(n31412), .dout(n31433));
  jand g14171(.dina(n31433), .dinb(n31431), .dout(n31434));
  jand g14172(.dina(n31434), .dinb(n284), .dout(n31435));
  jor  g14173(.dina(n31410), .dinb(n30841), .dout(n31436));
  jxor g14174(.dina(n31394), .dinb(n31393), .dout(n31437));
  jor  g14175(.dina(n31437), .dinb(n31412), .dout(n31438));
  jand g14176(.dina(n31438), .dinb(n31436), .dout(n31439));
  jand g14177(.dina(n31439), .dinb(n317), .dout(n31440));
  jor  g14178(.dina(n31410), .dinb(n30846), .dout(n31441));
  jxor g14179(.dina(n31391), .dinb(n31390), .dout(n31442));
  jor  g14180(.dina(n31442), .dinb(n31412), .dout(n31443));
  jand g14181(.dina(n31443), .dinb(n31441), .dout(n31444));
  jand g14182(.dina(n31444), .dinb(n316), .dout(n31445));
  jor  g14183(.dina(n31410), .dinb(n30851), .dout(n31446));
  jxor g14184(.dina(n31388), .dinb(n31387), .dout(n31447));
  jor  g14185(.dina(n31447), .dinb(n31412), .dout(n31448));
  jand g14186(.dina(n31448), .dinb(n31446), .dout(n31449));
  jand g14187(.dina(n31449), .dinb(n315), .dout(n31450));
  jor  g14188(.dina(n31410), .dinb(n30856), .dout(n31451));
  jxor g14189(.dina(n31385), .dinb(n31384), .dout(n31452));
  jor  g14190(.dina(n31452), .dinb(n31412), .dout(n31453));
  jand g14191(.dina(n31453), .dinb(n31451), .dout(n31454));
  jand g14192(.dina(n31454), .dinb(n283), .dout(n31455));
  jor  g14193(.dina(n31410), .dinb(n30861), .dout(n31456));
  jxor g14194(.dina(n31382), .dinb(n31381), .dout(n31457));
  jor  g14195(.dina(n31457), .dinb(n31412), .dout(n31458));
  jand g14196(.dina(n31458), .dinb(n31456), .dout(n31459));
  jand g14197(.dina(n31459), .dinb(n280), .dout(n31460));
  jor  g14198(.dina(n31410), .dinb(n30866), .dout(n31461));
  jxor g14199(.dina(n31379), .dinb(n31378), .dout(n31462));
  jor  g14200(.dina(n31462), .dinb(n31412), .dout(n31463));
  jand g14201(.dina(n31463), .dinb(n31461), .dout(n31464));
  jand g14202(.dina(n31464), .dinb(n279), .dout(n31465));
  jor  g14203(.dina(n31410), .dinb(n30871), .dout(n31466));
  jxor g14204(.dina(n31376), .dinb(n31375), .dout(n31467));
  jor  g14205(.dina(n31467), .dinb(n31412), .dout(n31468));
  jand g14206(.dina(n31468), .dinb(n31466), .dout(n31469));
  jand g14207(.dina(n31469), .dinb(n278), .dout(n31470));
  jor  g14208(.dina(n31410), .dinb(n30876), .dout(n31471));
  jxor g14209(.dina(n31373), .dinb(n31372), .dout(n31472));
  jor  g14210(.dina(n31472), .dinb(n31412), .dout(n31473));
  jand g14211(.dina(n31473), .dinb(n31471), .dout(n31474));
  jand g14212(.dina(n31474), .dinb(n277), .dout(n31475));
  jor  g14213(.dina(n31410), .dinb(n30881), .dout(n31476));
  jxor g14214(.dina(n31370), .dinb(n31369), .dout(n31477));
  jor  g14215(.dina(n31477), .dinb(n31412), .dout(n31478));
  jand g14216(.dina(n31478), .dinb(n31476), .dout(n31479));
  jand g14217(.dina(n31479), .dinb(n326), .dout(n31480));
  jor  g14218(.dina(n31410), .dinb(n30886), .dout(n31481));
  jxor g14219(.dina(n31367), .dinb(n31366), .dout(n31482));
  jor  g14220(.dina(n31482), .dinb(n31412), .dout(n31483));
  jand g14221(.dina(n31483), .dinb(n31481), .dout(n31484));
  jand g14222(.dina(n31484), .dinb(n325), .dout(n31485));
  jor  g14223(.dina(n31410), .dinb(n30891), .dout(n31486));
  jxor g14224(.dina(n31364), .dinb(n31363), .dout(n31487));
  jor  g14225(.dina(n31487), .dinb(n31412), .dout(n31488));
  jand g14226(.dina(n31488), .dinb(n31486), .dout(n31489));
  jand g14227(.dina(n31489), .dinb(n324), .dout(n31490));
  jor  g14228(.dina(n31410), .dinb(n30896), .dout(n31491));
  jxor g14229(.dina(n31361), .dinb(n31360), .dout(n31492));
  jor  g14230(.dina(n31492), .dinb(n31412), .dout(n31493));
  jand g14231(.dina(n31493), .dinb(n31491), .dout(n31494));
  jand g14232(.dina(n31494), .dinb(n276), .dout(n31495));
  jor  g14233(.dina(n31410), .dinb(n30901), .dout(n31496));
  jxor g14234(.dina(n31358), .dinb(n31357), .dout(n31497));
  jor  g14235(.dina(n31497), .dinb(n31412), .dout(n31498));
  jand g14236(.dina(n31498), .dinb(n31496), .dout(n31499));
  jand g14237(.dina(n31499), .dinb(n333), .dout(n31500));
  jor  g14238(.dina(n31410), .dinb(n30906), .dout(n31501));
  jxor g14239(.dina(n31355), .dinb(n31354), .dout(n31502));
  jor  g14240(.dina(n31502), .dinb(n31412), .dout(n31503));
  jand g14241(.dina(n31503), .dinb(n31501), .dout(n31504));
  jand g14242(.dina(n31504), .dinb(n332), .dout(n31505));
  jor  g14243(.dina(n31410), .dinb(n30911), .dout(n31506));
  jxor g14244(.dina(n31352), .dinb(n31351), .dout(n31507));
  jor  g14245(.dina(n31507), .dinb(n31412), .dout(n31508));
  jand g14246(.dina(n31508), .dinb(n31506), .dout(n31509));
  jand g14247(.dina(n31509), .dinb(n331), .dout(n31510));
  jor  g14248(.dina(n31410), .dinb(n30916), .dout(n31511));
  jxor g14249(.dina(n31349), .dinb(n31348), .dout(n31512));
  jor  g14250(.dina(n31512), .dinb(n31412), .dout(n31513));
  jand g14251(.dina(n31513), .dinb(n31511), .dout(n31514));
  jand g14252(.dina(n31514), .dinb(n275), .dout(n31515));
  jor  g14253(.dina(n31410), .dinb(n30921), .dout(n31516));
  jxor g14254(.dina(n31346), .dinb(n31345), .dout(n31517));
  jor  g14255(.dina(n31517), .dinb(n31412), .dout(n31518));
  jand g14256(.dina(n31518), .dinb(n31516), .dout(n31519));
  jand g14257(.dina(n31519), .dinb(n340), .dout(n31520));
  jor  g14258(.dina(n31410), .dinb(n30926), .dout(n31521));
  jxor g14259(.dina(n31343), .dinb(n31342), .dout(n31522));
  jor  g14260(.dina(n31522), .dinb(n31412), .dout(n31523));
  jand g14261(.dina(n31523), .dinb(n31521), .dout(n31524));
  jand g14262(.dina(n31524), .dinb(n339), .dout(n31525));
  jor  g14263(.dina(n31410), .dinb(n30931), .dout(n31526));
  jxor g14264(.dina(n31340), .dinb(n31339), .dout(n31527));
  jor  g14265(.dina(n31527), .dinb(n31412), .dout(n31528));
  jand g14266(.dina(n31528), .dinb(n31526), .dout(n31529));
  jand g14267(.dina(n31529), .dinb(n338), .dout(n31530));
  jor  g14268(.dina(n31410), .dinb(n30936), .dout(n31531));
  jxor g14269(.dina(n31337), .dinb(n31336), .dout(n31532));
  jor  g14270(.dina(n31532), .dinb(n31412), .dout(n31533));
  jand g14271(.dina(n31533), .dinb(n31531), .dout(n31534));
  jand g14272(.dina(n31534), .dinb(n271), .dout(n31535));
  jor  g14273(.dina(n31410), .dinb(n30941), .dout(n31536));
  jxor g14274(.dina(n31334), .dinb(n31333), .dout(n31537));
  jor  g14275(.dina(n31537), .dinb(n31412), .dout(n31538));
  jand g14276(.dina(n31538), .dinb(n31536), .dout(n31539));
  jand g14277(.dina(n31539), .dinb(n270), .dout(n31540));
  jor  g14278(.dina(n31410), .dinb(n30946), .dout(n31541));
  jxor g14279(.dina(n31331), .dinb(n31330), .dout(n31542));
  jor  g14280(.dina(n31542), .dinb(n31412), .dout(n31543));
  jand g14281(.dina(n31543), .dinb(n31541), .dout(n31544));
  jand g14282(.dina(n31544), .dinb(n269), .dout(n31545));
  jor  g14283(.dina(n31410), .dinb(n30951), .dout(n31546));
  jxor g14284(.dina(n31328), .dinb(n31327), .dout(n31547));
  jor  g14285(.dina(n31547), .dinb(n31412), .dout(n31548));
  jand g14286(.dina(n31548), .dinb(n31546), .dout(n31549));
  jand g14287(.dina(n31549), .dinb(n274), .dout(n31550));
  jor  g14288(.dina(n31410), .dinb(n30956), .dout(n31551));
  jxor g14289(.dina(n31325), .dinb(n31324), .dout(n31552));
  jor  g14290(.dina(n31552), .dinb(n31412), .dout(n31553));
  jand g14291(.dina(n31553), .dinb(n31551), .dout(n31554));
  jand g14292(.dina(n31554), .dinb(n268), .dout(n31555));
  jor  g14293(.dina(n31410), .dinb(n30961), .dout(n31556));
  jxor g14294(.dina(n31322), .dinb(n31321), .dout(n31557));
  jor  g14295(.dina(n31557), .dinb(n31412), .dout(n31558));
  jand g14296(.dina(n31558), .dinb(n31556), .dout(n31559));
  jand g14297(.dina(n31559), .dinb(n349), .dout(n31560));
  jor  g14298(.dina(n31410), .dinb(n30966), .dout(n31561));
  jxor g14299(.dina(n31319), .dinb(n31318), .dout(n31562));
  jor  g14300(.dina(n31562), .dinb(n31412), .dout(n31563));
  jand g14301(.dina(n31563), .dinb(n31561), .dout(n31564));
  jand g14302(.dina(n31564), .dinb(n348), .dout(n31565));
  jor  g14303(.dina(n31410), .dinb(n30971), .dout(n31566));
  jxor g14304(.dina(n31316), .dinb(n31315), .dout(n31567));
  jor  g14305(.dina(n31567), .dinb(n31412), .dout(n31568));
  jand g14306(.dina(n31568), .dinb(n31566), .dout(n31569));
  jand g14307(.dina(n31569), .dinb(n347), .dout(n31570));
  jor  g14308(.dina(n31410), .dinb(n30976), .dout(n31571));
  jxor g14309(.dina(n31313), .dinb(n31312), .dout(n31572));
  jor  g14310(.dina(n31572), .dinb(n31412), .dout(n31573));
  jand g14311(.dina(n31573), .dinb(n31571), .dout(n31574));
  jand g14312(.dina(n31574), .dinb(n267), .dout(n31575));
  jor  g14313(.dina(n31410), .dinb(n30981), .dout(n31576));
  jxor g14314(.dina(n31310), .dinb(n31309), .dout(n31577));
  jor  g14315(.dina(n31577), .dinb(n31412), .dout(n31578));
  jand g14316(.dina(n31578), .dinb(n31576), .dout(n31579));
  jand g14317(.dina(n31579), .dinb(n266), .dout(n31580));
  jor  g14318(.dina(n31410), .dinb(n30986), .dout(n31581));
  jxor g14319(.dina(n31307), .dinb(n31306), .dout(n31582));
  jor  g14320(.dina(n31582), .dinb(n31412), .dout(n31583));
  jand g14321(.dina(n31583), .dinb(n31581), .dout(n31584));
  jand g14322(.dina(n31584), .dinb(n356), .dout(n31585));
  jor  g14323(.dina(n31410), .dinb(n30991), .dout(n31586));
  jxor g14324(.dina(n31304), .dinb(n31303), .dout(n31587));
  jor  g14325(.dina(n31587), .dinb(n31412), .dout(n31588));
  jand g14326(.dina(n31588), .dinb(n31586), .dout(n31589));
  jand g14327(.dina(n31589), .dinb(n355), .dout(n31590));
  jor  g14328(.dina(n31410), .dinb(n30996), .dout(n31591));
  jxor g14329(.dina(n31301), .dinb(n31300), .dout(n31592));
  jor  g14330(.dina(n31592), .dinb(n31412), .dout(n31593));
  jand g14331(.dina(n31593), .dinb(n31591), .dout(n31594));
  jand g14332(.dina(n31594), .dinb(n364), .dout(n31595));
  jor  g14333(.dina(n31410), .dinb(n31001), .dout(n31596));
  jxor g14334(.dina(n31298), .dinb(n31297), .dout(n31597));
  jor  g14335(.dina(n31597), .dinb(n31412), .dout(n31598));
  jand g14336(.dina(n31598), .dinb(n31596), .dout(n31599));
  jand g14337(.dina(n31599), .dinb(n361), .dout(n31600));
  jor  g14338(.dina(n31410), .dinb(n31006), .dout(n31601));
  jxor g14339(.dina(n31295), .dinb(n31294), .dout(n31602));
  jor  g14340(.dina(n31602), .dinb(n31412), .dout(n31603));
  jand g14341(.dina(n31603), .dinb(n31601), .dout(n31604));
  jand g14342(.dina(n31604), .dinb(n360), .dout(n31605));
  jor  g14343(.dina(n31410), .dinb(n31011), .dout(n31606));
  jxor g14344(.dina(n31292), .dinb(n31291), .dout(n31607));
  jor  g14345(.dina(n31607), .dinb(n31412), .dout(n31608));
  jand g14346(.dina(n31608), .dinb(n31606), .dout(n31609));
  jand g14347(.dina(n31609), .dinb(n363), .dout(n31610));
  jor  g14348(.dina(n31410), .dinb(n31016), .dout(n31611));
  jxor g14349(.dina(n31289), .dinb(n31288), .dout(n31612));
  jor  g14350(.dina(n31612), .dinb(n31412), .dout(n31613));
  jand g14351(.dina(n31613), .dinb(n31611), .dout(n31614));
  jand g14352(.dina(n31614), .dinb(n359), .dout(n31615));
  jor  g14353(.dina(n31410), .dinb(n31021), .dout(n31616));
  jxor g14354(.dina(n31286), .dinb(n31285), .dout(n31617));
  jor  g14355(.dina(n31617), .dinb(n31412), .dout(n31618));
  jand g14356(.dina(n31618), .dinb(n31616), .dout(n31619));
  jand g14357(.dina(n31619), .dinb(n369), .dout(n31620));
  jor  g14358(.dina(n31410), .dinb(n31026), .dout(n31621));
  jxor g14359(.dina(n31283), .dinb(n31282), .dout(n31622));
  jor  g14360(.dina(n31622), .dinb(n31412), .dout(n31623));
  jand g14361(.dina(n31623), .dinb(n31621), .dout(n31624));
  jand g14362(.dina(n31624), .dinb(n368), .dout(n31625));
  jor  g14363(.dina(n31410), .dinb(n31031), .dout(n31626));
  jxor g14364(.dina(n31280), .dinb(n31279), .dout(n31627));
  jor  g14365(.dina(n31627), .dinb(n31412), .dout(n31628));
  jand g14366(.dina(n31628), .dinb(n31626), .dout(n31629));
  jand g14367(.dina(n31629), .dinb(n367), .dout(n31630));
  jor  g14368(.dina(n31410), .dinb(n31036), .dout(n31631));
  jxor g14369(.dina(n31277), .dinb(n31276), .dout(n31632));
  jor  g14370(.dina(n31632), .dinb(n31412), .dout(n31633));
  jand g14371(.dina(n31633), .dinb(n31631), .dout(n31634));
  jand g14372(.dina(n31634), .dinb(n265), .dout(n31635));
  jor  g14373(.dina(n31410), .dinb(n31041), .dout(n31636));
  jxor g14374(.dina(n31274), .dinb(n31273), .dout(n31637));
  jor  g14375(.dina(n31637), .dinb(n31412), .dout(n31638));
  jand g14376(.dina(n31638), .dinb(n31636), .dout(n31639));
  jand g14377(.dina(n31639), .dinb(n378), .dout(n31640));
  jor  g14378(.dina(n31410), .dinb(n31046), .dout(n31641));
  jxor g14379(.dina(n31271), .dinb(n31270), .dout(n31642));
  jor  g14380(.dina(n31642), .dinb(n31412), .dout(n31643));
  jand g14381(.dina(n31643), .dinb(n31641), .dout(n31644));
  jand g14382(.dina(n31644), .dinb(n377), .dout(n31645));
  jor  g14383(.dina(n31410), .dinb(n31051), .dout(n31646));
  jxor g14384(.dina(n31268), .dinb(n31267), .dout(n31647));
  jor  g14385(.dina(n31647), .dinb(n31412), .dout(n31648));
  jand g14386(.dina(n31648), .dinb(n31646), .dout(n31649));
  jand g14387(.dina(n31649), .dinb(n376), .dout(n31650));
  jor  g14388(.dina(n31410), .dinb(n31058), .dout(n31651));
  jxor g14389(.dina(n31265), .dinb(n31264), .dout(n31652));
  jor  g14390(.dina(n31652), .dinb(n31412), .dout(n31653));
  jand g14391(.dina(n31653), .dinb(n31651), .dout(n31654));
  jand g14392(.dina(n31654), .dinb(n264), .dout(n31655));
  jor  g14393(.dina(n31410), .dinb(n31261), .dout(n31656));
  jxor g14394(.dina(n31262), .dinb(n11197), .dout(n31657));
  jand g14395(.dina(n31657), .dinb(n31410), .dout(n31658));
  jnot g14396(.din(n31658), .dout(n31659));
  jand g14397(.dina(n31659), .dinb(n31656), .dout(n31660));
  jnot g14398(.din(n31660), .dout(n31661));
  jand g14399(.dina(n31661), .dinb(n386), .dout(n31662));
  jand g14400(.dina(n31410), .dinb(b0 ), .dout(n31663));
  jxor g14401(.dina(n31663), .dinb(a14 ), .dout(n31664));
  jand g14402(.dina(n31664), .dinb(n259), .dout(n31665));
  jxor g14403(.dina(n31663), .dinb(n11195), .dout(n31666));
  jxor g14404(.dina(n31666), .dinb(b1 ), .dout(n31667));
  jand g14405(.dina(n31667), .dinb(n11607), .dout(n31668));
  jor  g14406(.dina(n31668), .dinb(n31665), .dout(n31669));
  jxor g14407(.dina(n31660), .dinb(b2 ), .dout(n31670));
  jand g14408(.dina(n31670), .dinb(n31669), .dout(n31671));
  jor  g14409(.dina(n31671), .dinb(n31662), .dout(n31672));
  jxor g14410(.dina(n31654), .dinb(n264), .dout(n31673));
  jand g14411(.dina(n31673), .dinb(n31672), .dout(n31674));
  jor  g14412(.dina(n31674), .dinb(n31655), .dout(n31675));
  jxor g14413(.dina(n31649), .dinb(n376), .dout(n31676));
  jand g14414(.dina(n31676), .dinb(n31675), .dout(n31677));
  jor  g14415(.dina(n31677), .dinb(n31650), .dout(n31678));
  jxor g14416(.dina(n31644), .dinb(n377), .dout(n31679));
  jand g14417(.dina(n31679), .dinb(n31678), .dout(n31680));
  jor  g14418(.dina(n31680), .dinb(n31645), .dout(n31681));
  jxor g14419(.dina(n31639), .dinb(n378), .dout(n31682));
  jand g14420(.dina(n31682), .dinb(n31681), .dout(n31683));
  jor  g14421(.dina(n31683), .dinb(n31640), .dout(n31684));
  jxor g14422(.dina(n31634), .dinb(n265), .dout(n31685));
  jand g14423(.dina(n31685), .dinb(n31684), .dout(n31686));
  jor  g14424(.dina(n31686), .dinb(n31635), .dout(n31687));
  jxor g14425(.dina(n31629), .dinb(n367), .dout(n31688));
  jand g14426(.dina(n31688), .dinb(n31687), .dout(n31689));
  jor  g14427(.dina(n31689), .dinb(n31630), .dout(n31690));
  jxor g14428(.dina(n31624), .dinb(n368), .dout(n31691));
  jand g14429(.dina(n31691), .dinb(n31690), .dout(n31692));
  jor  g14430(.dina(n31692), .dinb(n31625), .dout(n31693));
  jxor g14431(.dina(n31619), .dinb(n369), .dout(n31694));
  jand g14432(.dina(n31694), .dinb(n31693), .dout(n31695));
  jor  g14433(.dina(n31695), .dinb(n31620), .dout(n31696));
  jxor g14434(.dina(n31614), .dinb(n359), .dout(n31697));
  jand g14435(.dina(n31697), .dinb(n31696), .dout(n31698));
  jor  g14436(.dina(n31698), .dinb(n31615), .dout(n31699));
  jxor g14437(.dina(n31609), .dinb(n363), .dout(n31700));
  jand g14438(.dina(n31700), .dinb(n31699), .dout(n31701));
  jor  g14439(.dina(n31701), .dinb(n31610), .dout(n31702));
  jxor g14440(.dina(n31604), .dinb(n360), .dout(n31703));
  jand g14441(.dina(n31703), .dinb(n31702), .dout(n31704));
  jor  g14442(.dina(n31704), .dinb(n31605), .dout(n31705));
  jxor g14443(.dina(n31599), .dinb(n361), .dout(n31706));
  jand g14444(.dina(n31706), .dinb(n31705), .dout(n31707));
  jor  g14445(.dina(n31707), .dinb(n31600), .dout(n31708));
  jxor g14446(.dina(n31594), .dinb(n364), .dout(n31709));
  jand g14447(.dina(n31709), .dinb(n31708), .dout(n31710));
  jor  g14448(.dina(n31710), .dinb(n31595), .dout(n31711));
  jxor g14449(.dina(n31589), .dinb(n355), .dout(n31712));
  jand g14450(.dina(n31712), .dinb(n31711), .dout(n31713));
  jor  g14451(.dina(n31713), .dinb(n31590), .dout(n31714));
  jxor g14452(.dina(n31584), .dinb(n356), .dout(n31715));
  jand g14453(.dina(n31715), .dinb(n31714), .dout(n31716));
  jor  g14454(.dina(n31716), .dinb(n31585), .dout(n31717));
  jxor g14455(.dina(n31579), .dinb(n266), .dout(n31718));
  jand g14456(.dina(n31718), .dinb(n31717), .dout(n31719));
  jor  g14457(.dina(n31719), .dinb(n31580), .dout(n31720));
  jxor g14458(.dina(n31574), .dinb(n267), .dout(n31721));
  jand g14459(.dina(n31721), .dinb(n31720), .dout(n31722));
  jor  g14460(.dina(n31722), .dinb(n31575), .dout(n31723));
  jxor g14461(.dina(n31569), .dinb(n347), .dout(n31724));
  jand g14462(.dina(n31724), .dinb(n31723), .dout(n31725));
  jor  g14463(.dina(n31725), .dinb(n31570), .dout(n31726));
  jxor g14464(.dina(n31564), .dinb(n348), .dout(n31727));
  jand g14465(.dina(n31727), .dinb(n31726), .dout(n31728));
  jor  g14466(.dina(n31728), .dinb(n31565), .dout(n31729));
  jxor g14467(.dina(n31559), .dinb(n349), .dout(n31730));
  jand g14468(.dina(n31730), .dinb(n31729), .dout(n31731));
  jor  g14469(.dina(n31731), .dinb(n31560), .dout(n31732));
  jxor g14470(.dina(n31554), .dinb(n268), .dout(n31733));
  jand g14471(.dina(n31733), .dinb(n31732), .dout(n31734));
  jor  g14472(.dina(n31734), .dinb(n31555), .dout(n31735));
  jxor g14473(.dina(n31549), .dinb(n274), .dout(n31736));
  jand g14474(.dina(n31736), .dinb(n31735), .dout(n31737));
  jor  g14475(.dina(n31737), .dinb(n31550), .dout(n31738));
  jxor g14476(.dina(n31544), .dinb(n269), .dout(n31739));
  jand g14477(.dina(n31739), .dinb(n31738), .dout(n31740));
  jor  g14478(.dina(n31740), .dinb(n31545), .dout(n31741));
  jxor g14479(.dina(n31539), .dinb(n270), .dout(n31742));
  jand g14480(.dina(n31742), .dinb(n31741), .dout(n31743));
  jor  g14481(.dina(n31743), .dinb(n31540), .dout(n31744));
  jxor g14482(.dina(n31534), .dinb(n271), .dout(n31745));
  jand g14483(.dina(n31745), .dinb(n31744), .dout(n31746));
  jor  g14484(.dina(n31746), .dinb(n31535), .dout(n31747));
  jxor g14485(.dina(n31529), .dinb(n338), .dout(n31748));
  jand g14486(.dina(n31748), .dinb(n31747), .dout(n31749));
  jor  g14487(.dina(n31749), .dinb(n31530), .dout(n31750));
  jxor g14488(.dina(n31524), .dinb(n339), .dout(n31751));
  jand g14489(.dina(n31751), .dinb(n31750), .dout(n31752));
  jor  g14490(.dina(n31752), .dinb(n31525), .dout(n31753));
  jxor g14491(.dina(n31519), .dinb(n340), .dout(n31754));
  jand g14492(.dina(n31754), .dinb(n31753), .dout(n31755));
  jor  g14493(.dina(n31755), .dinb(n31520), .dout(n31756));
  jxor g14494(.dina(n31514), .dinb(n275), .dout(n31757));
  jand g14495(.dina(n31757), .dinb(n31756), .dout(n31758));
  jor  g14496(.dina(n31758), .dinb(n31515), .dout(n31759));
  jxor g14497(.dina(n31509), .dinb(n331), .dout(n31760));
  jand g14498(.dina(n31760), .dinb(n31759), .dout(n31761));
  jor  g14499(.dina(n31761), .dinb(n31510), .dout(n31762));
  jxor g14500(.dina(n31504), .dinb(n332), .dout(n31763));
  jand g14501(.dina(n31763), .dinb(n31762), .dout(n31764));
  jor  g14502(.dina(n31764), .dinb(n31505), .dout(n31765));
  jxor g14503(.dina(n31499), .dinb(n333), .dout(n31766));
  jand g14504(.dina(n31766), .dinb(n31765), .dout(n31767));
  jor  g14505(.dina(n31767), .dinb(n31500), .dout(n31768));
  jxor g14506(.dina(n31494), .dinb(n276), .dout(n31769));
  jand g14507(.dina(n31769), .dinb(n31768), .dout(n31770));
  jor  g14508(.dina(n31770), .dinb(n31495), .dout(n31771));
  jxor g14509(.dina(n31489), .dinb(n324), .dout(n31772));
  jand g14510(.dina(n31772), .dinb(n31771), .dout(n31773));
  jor  g14511(.dina(n31773), .dinb(n31490), .dout(n31774));
  jxor g14512(.dina(n31484), .dinb(n325), .dout(n31775));
  jand g14513(.dina(n31775), .dinb(n31774), .dout(n31776));
  jor  g14514(.dina(n31776), .dinb(n31485), .dout(n31777));
  jxor g14515(.dina(n31479), .dinb(n326), .dout(n31778));
  jand g14516(.dina(n31778), .dinb(n31777), .dout(n31779));
  jor  g14517(.dina(n31779), .dinb(n31480), .dout(n31780));
  jxor g14518(.dina(n31474), .dinb(n277), .dout(n31781));
  jand g14519(.dina(n31781), .dinb(n31780), .dout(n31782));
  jor  g14520(.dina(n31782), .dinb(n31475), .dout(n31783));
  jxor g14521(.dina(n31469), .dinb(n278), .dout(n31784));
  jand g14522(.dina(n31784), .dinb(n31783), .dout(n31785));
  jor  g14523(.dina(n31785), .dinb(n31470), .dout(n31786));
  jxor g14524(.dina(n31464), .dinb(n279), .dout(n31787));
  jand g14525(.dina(n31787), .dinb(n31786), .dout(n31788));
  jor  g14526(.dina(n31788), .dinb(n31465), .dout(n31789));
  jxor g14527(.dina(n31459), .dinb(n280), .dout(n31790));
  jand g14528(.dina(n31790), .dinb(n31789), .dout(n31791));
  jor  g14529(.dina(n31791), .dinb(n31460), .dout(n31792));
  jxor g14530(.dina(n31454), .dinb(n283), .dout(n31793));
  jand g14531(.dina(n31793), .dinb(n31792), .dout(n31794));
  jor  g14532(.dina(n31794), .dinb(n31455), .dout(n31795));
  jxor g14533(.dina(n31449), .dinb(n315), .dout(n31796));
  jand g14534(.dina(n31796), .dinb(n31795), .dout(n31797));
  jor  g14535(.dina(n31797), .dinb(n31450), .dout(n31798));
  jxor g14536(.dina(n31444), .dinb(n316), .dout(n31799));
  jand g14537(.dina(n31799), .dinb(n31798), .dout(n31800));
  jor  g14538(.dina(n31800), .dinb(n31445), .dout(n31801));
  jxor g14539(.dina(n31439), .dinb(n317), .dout(n31802));
  jand g14540(.dina(n31802), .dinb(n31801), .dout(n31803));
  jor  g14541(.dina(n31803), .dinb(n31440), .dout(n31804));
  jxor g14542(.dina(n31434), .dinb(n284), .dout(n31805));
  jand g14543(.dina(n31805), .dinb(n31804), .dout(n31806));
  jor  g14544(.dina(n31806), .dinb(n31435), .dout(n31807));
  jxor g14545(.dina(n31429), .dinb(n285), .dout(n31808));
  jand g14546(.dina(n31808), .dinb(n31807), .dout(n31809));
  jor  g14547(.dina(n31809), .dinb(n31430), .dout(n31810));
  jxor g14548(.dina(n31415), .dinb(n286), .dout(n31811));
  jand g14549(.dina(n31811), .dinb(n31810), .dout(n31812));
  jor  g14550(.dina(n31812), .dinb(n31425), .dout(n31813));
  jand g14551(.dina(n31813), .dinb(n31424), .dout(n31814));
  jor  g14552(.dina(n31814), .dinb(n31421), .dout(n31815));
  jand g14553(.dina(n31815), .dinb(n310), .dout(n31816));
  jnot g14554(.din(n31816), .dout(n31817));
  jand g14555(.dina(n31817), .dinb(n31415), .dout(n31818));
  jxor g14556(.dina(n31811), .dinb(n31810), .dout(n31819));
  jand g14557(.dina(n31819), .dinb(n31816), .dout(n31820));
  jor  g14558(.dina(n31820), .dinb(n31818), .dout(n31821));
  jand g14559(.dina(n31817), .dinb(n31420), .dout(n31822));
  jand g14560(.dina(n31813), .dinb(n31421), .dout(n31823));
  jor  g14561(.dina(n31823), .dinb(n31822), .dout(n31824));
  jand g14562(.dina(n31824), .dinb(n288), .dout(n31825));
  jnot g14563(.din(n31824), .dout(n31826));
  jand g14564(.dina(n31826), .dinb(b51 ), .dout(n31827));
  jnot g14565(.din(n31827), .dout(n31828));
  jand g14566(.dina(n31821), .dinb(n287), .dout(n31829));
  jand g14567(.dina(n31817), .dinb(n31429), .dout(n31830));
  jxor g14568(.dina(n31808), .dinb(n31807), .dout(n31831));
  jand g14569(.dina(n31831), .dinb(n31816), .dout(n31832));
  jor  g14570(.dina(n31832), .dinb(n31830), .dout(n31833));
  jand g14571(.dina(n31833), .dinb(n286), .dout(n31834));
  jand g14572(.dina(n31817), .dinb(n31434), .dout(n31835));
  jxor g14573(.dina(n31805), .dinb(n31804), .dout(n31836));
  jand g14574(.dina(n31836), .dinb(n31816), .dout(n31837));
  jor  g14575(.dina(n31837), .dinb(n31835), .dout(n31838));
  jand g14576(.dina(n31838), .dinb(n285), .dout(n31839));
  jand g14577(.dina(n31817), .dinb(n31439), .dout(n31840));
  jxor g14578(.dina(n31802), .dinb(n31801), .dout(n31841));
  jand g14579(.dina(n31841), .dinb(n31816), .dout(n31842));
  jor  g14580(.dina(n31842), .dinb(n31840), .dout(n31843));
  jand g14581(.dina(n31843), .dinb(n284), .dout(n31844));
  jand g14582(.dina(n31817), .dinb(n31444), .dout(n31845));
  jxor g14583(.dina(n31799), .dinb(n31798), .dout(n31846));
  jand g14584(.dina(n31846), .dinb(n31816), .dout(n31847));
  jor  g14585(.dina(n31847), .dinb(n31845), .dout(n31848));
  jand g14586(.dina(n31848), .dinb(n317), .dout(n31849));
  jand g14587(.dina(n31817), .dinb(n31449), .dout(n31850));
  jxor g14588(.dina(n31796), .dinb(n31795), .dout(n31851));
  jand g14589(.dina(n31851), .dinb(n31816), .dout(n31852));
  jor  g14590(.dina(n31852), .dinb(n31850), .dout(n31853));
  jand g14591(.dina(n31853), .dinb(n316), .dout(n31854));
  jor  g14592(.dina(n31816), .dinb(n31454), .dout(n31855));
  jxor g14593(.dina(n31793), .dinb(n31792), .dout(n31856));
  jor  g14594(.dina(n31856), .dinb(n31817), .dout(n31857));
  jand g14595(.dina(n31857), .dinb(n31855), .dout(n31858));
  jand g14596(.dina(n31858), .dinb(n315), .dout(n31859));
  jand g14597(.dina(n31817), .dinb(n31459), .dout(n31860));
  jxor g14598(.dina(n31790), .dinb(n31789), .dout(n31861));
  jand g14599(.dina(n31861), .dinb(n31816), .dout(n31862));
  jor  g14600(.dina(n31862), .dinb(n31860), .dout(n31863));
  jand g14601(.dina(n31863), .dinb(n283), .dout(n31864));
  jand g14602(.dina(n31817), .dinb(n31464), .dout(n31865));
  jxor g14603(.dina(n31787), .dinb(n31786), .dout(n31866));
  jand g14604(.dina(n31866), .dinb(n31816), .dout(n31867));
  jor  g14605(.dina(n31867), .dinb(n31865), .dout(n31868));
  jand g14606(.dina(n31868), .dinb(n280), .dout(n31869));
  jand g14607(.dina(n31817), .dinb(n31469), .dout(n31870));
  jxor g14608(.dina(n31784), .dinb(n31783), .dout(n31871));
  jand g14609(.dina(n31871), .dinb(n31816), .dout(n31872));
  jor  g14610(.dina(n31872), .dinb(n31870), .dout(n31873));
  jand g14611(.dina(n31873), .dinb(n279), .dout(n31874));
  jor  g14612(.dina(n31816), .dinb(n31474), .dout(n31875));
  jxor g14613(.dina(n31781), .dinb(n31780), .dout(n31876));
  jor  g14614(.dina(n31876), .dinb(n31817), .dout(n31877));
  jand g14615(.dina(n31877), .dinb(n31875), .dout(n31878));
  jand g14616(.dina(n31878), .dinb(n278), .dout(n31879));
  jor  g14617(.dina(n31816), .dinb(n31479), .dout(n31880));
  jxor g14618(.dina(n31778), .dinb(n31777), .dout(n31881));
  jor  g14619(.dina(n31881), .dinb(n31817), .dout(n31882));
  jand g14620(.dina(n31882), .dinb(n31880), .dout(n31883));
  jand g14621(.dina(n31883), .dinb(n277), .dout(n31884));
  jand g14622(.dina(n31817), .dinb(n31484), .dout(n31885));
  jxor g14623(.dina(n31775), .dinb(n31774), .dout(n31886));
  jand g14624(.dina(n31886), .dinb(n31816), .dout(n31887));
  jor  g14625(.dina(n31887), .dinb(n31885), .dout(n31888));
  jand g14626(.dina(n31888), .dinb(n326), .dout(n31889));
  jor  g14627(.dina(n31816), .dinb(n31489), .dout(n31890));
  jxor g14628(.dina(n31772), .dinb(n31771), .dout(n31891));
  jor  g14629(.dina(n31891), .dinb(n31817), .dout(n31892));
  jand g14630(.dina(n31892), .dinb(n31890), .dout(n31893));
  jand g14631(.dina(n31893), .dinb(n325), .dout(n31894));
  jand g14632(.dina(n31817), .dinb(n31494), .dout(n31895));
  jxor g14633(.dina(n31769), .dinb(n31768), .dout(n31896));
  jand g14634(.dina(n31896), .dinb(n31816), .dout(n31897));
  jor  g14635(.dina(n31897), .dinb(n31895), .dout(n31898));
  jand g14636(.dina(n31898), .dinb(n324), .dout(n31899));
  jand g14637(.dina(n31817), .dinb(n31499), .dout(n31900));
  jxor g14638(.dina(n31766), .dinb(n31765), .dout(n31901));
  jand g14639(.dina(n31901), .dinb(n31816), .dout(n31902));
  jor  g14640(.dina(n31902), .dinb(n31900), .dout(n31903));
  jand g14641(.dina(n31903), .dinb(n276), .dout(n31904));
  jand g14642(.dina(n31817), .dinb(n31504), .dout(n31905));
  jxor g14643(.dina(n31763), .dinb(n31762), .dout(n31906));
  jand g14644(.dina(n31906), .dinb(n31816), .dout(n31907));
  jor  g14645(.dina(n31907), .dinb(n31905), .dout(n31908));
  jand g14646(.dina(n31908), .dinb(n333), .dout(n31909));
  jand g14647(.dina(n31817), .dinb(n31509), .dout(n31910));
  jxor g14648(.dina(n31760), .dinb(n31759), .dout(n31911));
  jand g14649(.dina(n31911), .dinb(n31816), .dout(n31912));
  jor  g14650(.dina(n31912), .dinb(n31910), .dout(n31913));
  jand g14651(.dina(n31913), .dinb(n332), .dout(n31914));
  jand g14652(.dina(n31817), .dinb(n31514), .dout(n31915));
  jxor g14653(.dina(n31757), .dinb(n31756), .dout(n31916));
  jand g14654(.dina(n31916), .dinb(n31816), .dout(n31917));
  jor  g14655(.dina(n31917), .dinb(n31915), .dout(n31918));
  jand g14656(.dina(n31918), .dinb(n331), .dout(n31919));
  jor  g14657(.dina(n31816), .dinb(n31519), .dout(n31920));
  jxor g14658(.dina(n31754), .dinb(n31753), .dout(n31921));
  jor  g14659(.dina(n31921), .dinb(n31817), .dout(n31922));
  jand g14660(.dina(n31922), .dinb(n31920), .dout(n31923));
  jand g14661(.dina(n31923), .dinb(n275), .dout(n31924));
  jand g14662(.dina(n31817), .dinb(n31524), .dout(n31925));
  jxor g14663(.dina(n31751), .dinb(n31750), .dout(n31926));
  jand g14664(.dina(n31926), .dinb(n31816), .dout(n31927));
  jor  g14665(.dina(n31927), .dinb(n31925), .dout(n31928));
  jand g14666(.dina(n31928), .dinb(n340), .dout(n31929));
  jor  g14667(.dina(n31816), .dinb(n31529), .dout(n31930));
  jxor g14668(.dina(n31748), .dinb(n31747), .dout(n31931));
  jor  g14669(.dina(n31931), .dinb(n31817), .dout(n31932));
  jand g14670(.dina(n31932), .dinb(n31930), .dout(n31933));
  jand g14671(.dina(n31933), .dinb(n339), .dout(n31934));
  jor  g14672(.dina(n31816), .dinb(n31534), .dout(n31935));
  jxor g14673(.dina(n31745), .dinb(n31744), .dout(n31936));
  jor  g14674(.dina(n31936), .dinb(n31817), .dout(n31937));
  jand g14675(.dina(n31937), .dinb(n31935), .dout(n31938));
  jand g14676(.dina(n31938), .dinb(n338), .dout(n31939));
  jand g14677(.dina(n31817), .dinb(n31539), .dout(n31940));
  jxor g14678(.dina(n31742), .dinb(n31741), .dout(n31941));
  jand g14679(.dina(n31941), .dinb(n31816), .dout(n31942));
  jor  g14680(.dina(n31942), .dinb(n31940), .dout(n31943));
  jand g14681(.dina(n31943), .dinb(n271), .dout(n31944));
  jand g14682(.dina(n31817), .dinb(n31544), .dout(n31945));
  jxor g14683(.dina(n31739), .dinb(n31738), .dout(n31946));
  jand g14684(.dina(n31946), .dinb(n31816), .dout(n31947));
  jor  g14685(.dina(n31947), .dinb(n31945), .dout(n31948));
  jand g14686(.dina(n31948), .dinb(n270), .dout(n31949));
  jand g14687(.dina(n31817), .dinb(n31549), .dout(n31950));
  jxor g14688(.dina(n31736), .dinb(n31735), .dout(n31951));
  jand g14689(.dina(n31951), .dinb(n31816), .dout(n31952));
  jor  g14690(.dina(n31952), .dinb(n31950), .dout(n31953));
  jand g14691(.dina(n31953), .dinb(n269), .dout(n31954));
  jor  g14692(.dina(n31816), .dinb(n31554), .dout(n31955));
  jxor g14693(.dina(n31733), .dinb(n31732), .dout(n31956));
  jor  g14694(.dina(n31956), .dinb(n31817), .dout(n31957));
  jand g14695(.dina(n31957), .dinb(n31955), .dout(n31958));
  jand g14696(.dina(n31958), .dinb(n274), .dout(n31959));
  jor  g14697(.dina(n31816), .dinb(n31559), .dout(n31960));
  jxor g14698(.dina(n31730), .dinb(n31729), .dout(n31961));
  jor  g14699(.dina(n31961), .dinb(n31817), .dout(n31962));
  jand g14700(.dina(n31962), .dinb(n31960), .dout(n31963));
  jand g14701(.dina(n31963), .dinb(n268), .dout(n31964));
  jand g14702(.dina(n31817), .dinb(n31564), .dout(n31965));
  jxor g14703(.dina(n31727), .dinb(n31726), .dout(n31966));
  jand g14704(.dina(n31966), .dinb(n31816), .dout(n31967));
  jor  g14705(.dina(n31967), .dinb(n31965), .dout(n31968));
  jand g14706(.dina(n31968), .dinb(n349), .dout(n31969));
  jor  g14707(.dina(n31816), .dinb(n31569), .dout(n31970));
  jxor g14708(.dina(n31724), .dinb(n31723), .dout(n31971));
  jor  g14709(.dina(n31971), .dinb(n31817), .dout(n31972));
  jand g14710(.dina(n31972), .dinb(n31970), .dout(n31973));
  jand g14711(.dina(n31973), .dinb(n348), .dout(n31974));
  jor  g14712(.dina(n31816), .dinb(n31574), .dout(n31975));
  jxor g14713(.dina(n31721), .dinb(n31720), .dout(n31976));
  jor  g14714(.dina(n31976), .dinb(n31817), .dout(n31977));
  jand g14715(.dina(n31977), .dinb(n31975), .dout(n31978));
  jand g14716(.dina(n31978), .dinb(n347), .dout(n31979));
  jor  g14717(.dina(n31816), .dinb(n31579), .dout(n31980));
  jxor g14718(.dina(n31718), .dinb(n31717), .dout(n31981));
  jor  g14719(.dina(n31981), .dinb(n31817), .dout(n31982));
  jand g14720(.dina(n31982), .dinb(n31980), .dout(n31983));
  jand g14721(.dina(n31983), .dinb(n267), .dout(n31984));
  jand g14722(.dina(n31817), .dinb(n31584), .dout(n31985));
  jxor g14723(.dina(n31715), .dinb(n31714), .dout(n31986));
  jand g14724(.dina(n31986), .dinb(n31816), .dout(n31987));
  jor  g14725(.dina(n31987), .dinb(n31985), .dout(n31988));
  jand g14726(.dina(n31988), .dinb(n266), .dout(n31989));
  jand g14727(.dina(n31817), .dinb(n31589), .dout(n31990));
  jxor g14728(.dina(n31712), .dinb(n31711), .dout(n31991));
  jand g14729(.dina(n31991), .dinb(n31816), .dout(n31992));
  jor  g14730(.dina(n31992), .dinb(n31990), .dout(n31993));
  jand g14731(.dina(n31993), .dinb(n356), .dout(n31994));
  jand g14732(.dina(n31817), .dinb(n31594), .dout(n31995));
  jxor g14733(.dina(n31709), .dinb(n31708), .dout(n31996));
  jand g14734(.dina(n31996), .dinb(n31816), .dout(n31997));
  jor  g14735(.dina(n31997), .dinb(n31995), .dout(n31998));
  jand g14736(.dina(n31998), .dinb(n355), .dout(n31999));
  jand g14737(.dina(n31817), .dinb(n31599), .dout(n32000));
  jxor g14738(.dina(n31706), .dinb(n31705), .dout(n32001));
  jand g14739(.dina(n32001), .dinb(n31816), .dout(n32002));
  jor  g14740(.dina(n32002), .dinb(n32000), .dout(n32003));
  jand g14741(.dina(n32003), .dinb(n364), .dout(n32004));
  jand g14742(.dina(n31817), .dinb(n31604), .dout(n32005));
  jxor g14743(.dina(n31703), .dinb(n31702), .dout(n32006));
  jand g14744(.dina(n32006), .dinb(n31816), .dout(n32007));
  jor  g14745(.dina(n32007), .dinb(n32005), .dout(n32008));
  jand g14746(.dina(n32008), .dinb(n361), .dout(n32009));
  jand g14747(.dina(n31817), .dinb(n31609), .dout(n32010));
  jxor g14748(.dina(n31700), .dinb(n31699), .dout(n32011));
  jand g14749(.dina(n32011), .dinb(n31816), .dout(n32012));
  jor  g14750(.dina(n32012), .dinb(n32010), .dout(n32013));
  jand g14751(.dina(n32013), .dinb(n360), .dout(n32014));
  jor  g14752(.dina(n31816), .dinb(n31614), .dout(n32015));
  jxor g14753(.dina(n31697), .dinb(n31696), .dout(n32016));
  jor  g14754(.dina(n32016), .dinb(n31817), .dout(n32017));
  jand g14755(.dina(n32017), .dinb(n32015), .dout(n32018));
  jand g14756(.dina(n32018), .dinb(n363), .dout(n32019));
  jand g14757(.dina(n31817), .dinb(n31619), .dout(n32020));
  jxor g14758(.dina(n31694), .dinb(n31693), .dout(n32021));
  jand g14759(.dina(n32021), .dinb(n31816), .dout(n32022));
  jor  g14760(.dina(n32022), .dinb(n32020), .dout(n32023));
  jand g14761(.dina(n32023), .dinb(n359), .dout(n32024));
  jand g14762(.dina(n31817), .dinb(n31624), .dout(n32025));
  jxor g14763(.dina(n31691), .dinb(n31690), .dout(n32026));
  jand g14764(.dina(n32026), .dinb(n31816), .dout(n32027));
  jor  g14765(.dina(n32027), .dinb(n32025), .dout(n32028));
  jand g14766(.dina(n32028), .dinb(n369), .dout(n32029));
  jand g14767(.dina(n31817), .dinb(n31629), .dout(n32030));
  jxor g14768(.dina(n31688), .dinb(n31687), .dout(n32031));
  jand g14769(.dina(n32031), .dinb(n31816), .dout(n32032));
  jor  g14770(.dina(n32032), .dinb(n32030), .dout(n32033));
  jand g14771(.dina(n32033), .dinb(n368), .dout(n32034));
  jor  g14772(.dina(n31816), .dinb(n31634), .dout(n32035));
  jxor g14773(.dina(n31685), .dinb(n31684), .dout(n32036));
  jor  g14774(.dina(n32036), .dinb(n31817), .dout(n32037));
  jand g14775(.dina(n32037), .dinb(n32035), .dout(n32038));
  jand g14776(.dina(n32038), .dinb(n367), .dout(n32039));
  jor  g14777(.dina(n31816), .dinb(n31639), .dout(n32040));
  jxor g14778(.dina(n31682), .dinb(n31681), .dout(n32041));
  jor  g14779(.dina(n32041), .dinb(n31817), .dout(n32042));
  jand g14780(.dina(n32042), .dinb(n32040), .dout(n32043));
  jand g14781(.dina(n32043), .dinb(n265), .dout(n32044));
  jand g14782(.dina(n31817), .dinb(n31644), .dout(n32045));
  jxor g14783(.dina(n31679), .dinb(n31678), .dout(n32046));
  jand g14784(.dina(n32046), .dinb(n31816), .dout(n32047));
  jor  g14785(.dina(n32047), .dinb(n32045), .dout(n32048));
  jand g14786(.dina(n32048), .dinb(n378), .dout(n32049));
  jor  g14787(.dina(n31816), .dinb(n31649), .dout(n32050));
  jxor g14788(.dina(n31676), .dinb(n31675), .dout(n32051));
  jor  g14789(.dina(n32051), .dinb(n31817), .dout(n32052));
  jand g14790(.dina(n32052), .dinb(n32050), .dout(n32053));
  jand g14791(.dina(n32053), .dinb(n377), .dout(n32054));
  jand g14792(.dina(n31817), .dinb(n31654), .dout(n32055));
  jxor g14793(.dina(n31673), .dinb(n31672), .dout(n32056));
  jand g14794(.dina(n32056), .dinb(n31816), .dout(n32057));
  jor  g14795(.dina(n32057), .dinb(n32055), .dout(n32058));
  jand g14796(.dina(n32058), .dinb(n376), .dout(n32059));
  jor  g14797(.dina(n31816), .dinb(n31660), .dout(n32060));
  jxor g14798(.dina(n31670), .dinb(n31669), .dout(n32061));
  jnot g14799(.din(n32061), .dout(n32062));
  jor  g14800(.dina(n32062), .dinb(n31817), .dout(n32063));
  jand g14801(.dina(n32063), .dinb(n32060), .dout(n32064));
  jnot g14802(.din(n32064), .dout(n32065));
  jand g14803(.dina(n32065), .dinb(n264), .dout(n32066));
  jxor g14804(.dina(n31667), .dinb(n11607), .dout(n32067));
  jand g14805(.dina(n32067), .dinb(n31816), .dout(n32068));
  jnot g14806(.din(n32068), .dout(n32069));
  jor  g14807(.dina(n31816), .dinb(n31666), .dout(n32070));
  jand g14808(.dina(n32070), .dinb(n32069), .dout(n32071));
  jnot g14809(.din(n32071), .dout(n32072));
  jand g14810(.dina(n32072), .dinb(n386), .dout(n32073));
  jand g14811(.dina(n31816), .dinb(b0 ), .dout(n32074));
  jxor g14812(.dina(n32074), .dinb(a13 ), .dout(n32075));
  jand g14813(.dina(n32075), .dinb(n259), .dout(n32076));
  jxor g14814(.dina(n32074), .dinb(n11605), .dout(n32077));
  jxor g14815(.dina(n32077), .dinb(b1 ), .dout(n32078));
  jand g14816(.dina(n32078), .dinb(n12017), .dout(n32079));
  jor  g14817(.dina(n32079), .dinb(n32076), .dout(n32080));
  jxor g14818(.dina(n32071), .dinb(b2 ), .dout(n32081));
  jand g14819(.dina(n32081), .dinb(n32080), .dout(n32082));
  jor  g14820(.dina(n32082), .dinb(n32073), .dout(n32083));
  jxor g14821(.dina(n32064), .dinb(b3 ), .dout(n32084));
  jand g14822(.dina(n32084), .dinb(n32083), .dout(n32085));
  jor  g14823(.dina(n32085), .dinb(n32066), .dout(n32086));
  jxor g14824(.dina(n32058), .dinb(n376), .dout(n32087));
  jand g14825(.dina(n32087), .dinb(n32086), .dout(n32088));
  jor  g14826(.dina(n32088), .dinb(n32059), .dout(n32089));
  jxor g14827(.dina(n32053), .dinb(n377), .dout(n32090));
  jand g14828(.dina(n32090), .dinb(n32089), .dout(n32091));
  jor  g14829(.dina(n32091), .dinb(n32054), .dout(n32092));
  jxor g14830(.dina(n32048), .dinb(n378), .dout(n32093));
  jand g14831(.dina(n32093), .dinb(n32092), .dout(n32094));
  jor  g14832(.dina(n32094), .dinb(n32049), .dout(n32095));
  jxor g14833(.dina(n32043), .dinb(n265), .dout(n32096));
  jand g14834(.dina(n32096), .dinb(n32095), .dout(n32097));
  jor  g14835(.dina(n32097), .dinb(n32044), .dout(n32098));
  jxor g14836(.dina(n32038), .dinb(n367), .dout(n32099));
  jand g14837(.dina(n32099), .dinb(n32098), .dout(n32100));
  jor  g14838(.dina(n32100), .dinb(n32039), .dout(n32101));
  jxor g14839(.dina(n32033), .dinb(n368), .dout(n32102));
  jand g14840(.dina(n32102), .dinb(n32101), .dout(n32103));
  jor  g14841(.dina(n32103), .dinb(n32034), .dout(n32104));
  jxor g14842(.dina(n32028), .dinb(n369), .dout(n32105));
  jand g14843(.dina(n32105), .dinb(n32104), .dout(n32106));
  jor  g14844(.dina(n32106), .dinb(n32029), .dout(n32107));
  jxor g14845(.dina(n32023), .dinb(n359), .dout(n32108));
  jand g14846(.dina(n32108), .dinb(n32107), .dout(n32109));
  jor  g14847(.dina(n32109), .dinb(n32024), .dout(n32110));
  jxor g14848(.dina(n32018), .dinb(n363), .dout(n32111));
  jand g14849(.dina(n32111), .dinb(n32110), .dout(n32112));
  jor  g14850(.dina(n32112), .dinb(n32019), .dout(n32113));
  jxor g14851(.dina(n32013), .dinb(n360), .dout(n32114));
  jand g14852(.dina(n32114), .dinb(n32113), .dout(n32115));
  jor  g14853(.dina(n32115), .dinb(n32014), .dout(n32116));
  jxor g14854(.dina(n32008), .dinb(n361), .dout(n32117));
  jand g14855(.dina(n32117), .dinb(n32116), .dout(n32118));
  jor  g14856(.dina(n32118), .dinb(n32009), .dout(n32119));
  jxor g14857(.dina(n32003), .dinb(n364), .dout(n32120));
  jand g14858(.dina(n32120), .dinb(n32119), .dout(n32121));
  jor  g14859(.dina(n32121), .dinb(n32004), .dout(n32122));
  jxor g14860(.dina(n31998), .dinb(n355), .dout(n32123));
  jand g14861(.dina(n32123), .dinb(n32122), .dout(n32124));
  jor  g14862(.dina(n32124), .dinb(n31999), .dout(n32125));
  jxor g14863(.dina(n31993), .dinb(n356), .dout(n32126));
  jand g14864(.dina(n32126), .dinb(n32125), .dout(n32127));
  jor  g14865(.dina(n32127), .dinb(n31994), .dout(n32128));
  jxor g14866(.dina(n31988), .dinb(n266), .dout(n32129));
  jand g14867(.dina(n32129), .dinb(n32128), .dout(n32130));
  jor  g14868(.dina(n32130), .dinb(n31989), .dout(n32131));
  jxor g14869(.dina(n31983), .dinb(n267), .dout(n32132));
  jand g14870(.dina(n32132), .dinb(n32131), .dout(n32133));
  jor  g14871(.dina(n32133), .dinb(n31984), .dout(n32134));
  jxor g14872(.dina(n31978), .dinb(n347), .dout(n32135));
  jand g14873(.dina(n32135), .dinb(n32134), .dout(n32136));
  jor  g14874(.dina(n32136), .dinb(n31979), .dout(n32137));
  jxor g14875(.dina(n31973), .dinb(n348), .dout(n32138));
  jand g14876(.dina(n32138), .dinb(n32137), .dout(n32139));
  jor  g14877(.dina(n32139), .dinb(n31974), .dout(n32140));
  jxor g14878(.dina(n31968), .dinb(n349), .dout(n32141));
  jand g14879(.dina(n32141), .dinb(n32140), .dout(n32142));
  jor  g14880(.dina(n32142), .dinb(n31969), .dout(n32143));
  jxor g14881(.dina(n31963), .dinb(n268), .dout(n32144));
  jand g14882(.dina(n32144), .dinb(n32143), .dout(n32145));
  jor  g14883(.dina(n32145), .dinb(n31964), .dout(n32146));
  jxor g14884(.dina(n31958), .dinb(n274), .dout(n32147));
  jand g14885(.dina(n32147), .dinb(n32146), .dout(n32148));
  jor  g14886(.dina(n32148), .dinb(n31959), .dout(n32149));
  jxor g14887(.dina(n31953), .dinb(n269), .dout(n32150));
  jand g14888(.dina(n32150), .dinb(n32149), .dout(n32151));
  jor  g14889(.dina(n32151), .dinb(n31954), .dout(n32152));
  jxor g14890(.dina(n31948), .dinb(n270), .dout(n32153));
  jand g14891(.dina(n32153), .dinb(n32152), .dout(n32154));
  jor  g14892(.dina(n32154), .dinb(n31949), .dout(n32155));
  jxor g14893(.dina(n31943), .dinb(n271), .dout(n32156));
  jand g14894(.dina(n32156), .dinb(n32155), .dout(n32157));
  jor  g14895(.dina(n32157), .dinb(n31944), .dout(n32158));
  jxor g14896(.dina(n31938), .dinb(n338), .dout(n32159));
  jand g14897(.dina(n32159), .dinb(n32158), .dout(n32160));
  jor  g14898(.dina(n32160), .dinb(n31939), .dout(n32161));
  jxor g14899(.dina(n31933), .dinb(n339), .dout(n32162));
  jand g14900(.dina(n32162), .dinb(n32161), .dout(n32163));
  jor  g14901(.dina(n32163), .dinb(n31934), .dout(n32164));
  jxor g14902(.dina(n31928), .dinb(n340), .dout(n32165));
  jand g14903(.dina(n32165), .dinb(n32164), .dout(n32166));
  jor  g14904(.dina(n32166), .dinb(n31929), .dout(n32167));
  jxor g14905(.dina(n31923), .dinb(n275), .dout(n32168));
  jand g14906(.dina(n32168), .dinb(n32167), .dout(n32169));
  jor  g14907(.dina(n32169), .dinb(n31924), .dout(n32170));
  jxor g14908(.dina(n31918), .dinb(n331), .dout(n32171));
  jand g14909(.dina(n32171), .dinb(n32170), .dout(n32172));
  jor  g14910(.dina(n32172), .dinb(n31919), .dout(n32173));
  jxor g14911(.dina(n31913), .dinb(n332), .dout(n32174));
  jand g14912(.dina(n32174), .dinb(n32173), .dout(n32175));
  jor  g14913(.dina(n32175), .dinb(n31914), .dout(n32176));
  jxor g14914(.dina(n31908), .dinb(n333), .dout(n32177));
  jand g14915(.dina(n32177), .dinb(n32176), .dout(n32178));
  jor  g14916(.dina(n32178), .dinb(n31909), .dout(n32179));
  jxor g14917(.dina(n31903), .dinb(n276), .dout(n32180));
  jand g14918(.dina(n32180), .dinb(n32179), .dout(n32181));
  jor  g14919(.dina(n32181), .dinb(n31904), .dout(n32182));
  jxor g14920(.dina(n31898), .dinb(n324), .dout(n32183));
  jand g14921(.dina(n32183), .dinb(n32182), .dout(n32184));
  jor  g14922(.dina(n32184), .dinb(n31899), .dout(n32185));
  jxor g14923(.dina(n31893), .dinb(n325), .dout(n32186));
  jand g14924(.dina(n32186), .dinb(n32185), .dout(n32187));
  jor  g14925(.dina(n32187), .dinb(n31894), .dout(n32188));
  jxor g14926(.dina(n31888), .dinb(n326), .dout(n32189));
  jand g14927(.dina(n32189), .dinb(n32188), .dout(n32190));
  jor  g14928(.dina(n32190), .dinb(n31889), .dout(n32191));
  jxor g14929(.dina(n31883), .dinb(n277), .dout(n32192));
  jand g14930(.dina(n32192), .dinb(n32191), .dout(n32193));
  jor  g14931(.dina(n32193), .dinb(n31884), .dout(n32194));
  jxor g14932(.dina(n31878), .dinb(n278), .dout(n32195));
  jand g14933(.dina(n32195), .dinb(n32194), .dout(n32196));
  jor  g14934(.dina(n32196), .dinb(n31879), .dout(n32197));
  jxor g14935(.dina(n31873), .dinb(n279), .dout(n32198));
  jand g14936(.dina(n32198), .dinb(n32197), .dout(n32199));
  jor  g14937(.dina(n32199), .dinb(n31874), .dout(n32200));
  jxor g14938(.dina(n31868), .dinb(n280), .dout(n32201));
  jand g14939(.dina(n32201), .dinb(n32200), .dout(n32202));
  jor  g14940(.dina(n32202), .dinb(n31869), .dout(n32203));
  jxor g14941(.dina(n31863), .dinb(n283), .dout(n32204));
  jand g14942(.dina(n32204), .dinb(n32203), .dout(n32205));
  jor  g14943(.dina(n32205), .dinb(n31864), .dout(n32206));
  jxor g14944(.dina(n31858), .dinb(n315), .dout(n32207));
  jand g14945(.dina(n32207), .dinb(n32206), .dout(n32208));
  jor  g14946(.dina(n32208), .dinb(n31859), .dout(n32209));
  jxor g14947(.dina(n31853), .dinb(n316), .dout(n32210));
  jand g14948(.dina(n32210), .dinb(n32209), .dout(n32211));
  jor  g14949(.dina(n32211), .dinb(n31854), .dout(n32212));
  jxor g14950(.dina(n31848), .dinb(n317), .dout(n32213));
  jand g14951(.dina(n32213), .dinb(n32212), .dout(n32214));
  jor  g14952(.dina(n32214), .dinb(n31849), .dout(n32215));
  jxor g14953(.dina(n31843), .dinb(n284), .dout(n32216));
  jand g14954(.dina(n32216), .dinb(n32215), .dout(n32217));
  jor  g14955(.dina(n32217), .dinb(n31844), .dout(n32218));
  jxor g14956(.dina(n31838), .dinb(n285), .dout(n32219));
  jand g14957(.dina(n32219), .dinb(n32218), .dout(n32220));
  jor  g14958(.dina(n32220), .dinb(n31839), .dout(n32221));
  jxor g14959(.dina(n31833), .dinb(n286), .dout(n32222));
  jand g14960(.dina(n32222), .dinb(n32221), .dout(n32223));
  jor  g14961(.dina(n32223), .dinb(n31834), .dout(n32224));
  jxor g14962(.dina(n31821), .dinb(n287), .dout(n32225));
  jand g14963(.dina(n32225), .dinb(n32224), .dout(n32226));
  jor  g14964(.dina(n32226), .dinb(n31829), .dout(n32227));
  jand g14965(.dina(n32227), .dinb(n31828), .dout(n32228));
  jor  g14966(.dina(n32228), .dinb(n31825), .dout(n32229));
  jand g14967(.dina(n32229), .dinb(n309), .dout(n32230));
  jor  g14968(.dina(n32230), .dinb(n31821), .dout(n32231));
  jnot g14969(.din(n32230), .dout(n32232));
  jxor g14970(.dina(n32225), .dinb(n32224), .dout(n32233));
  jor  g14971(.dina(n32233), .dinb(n32232), .dout(n32234));
  jand g14972(.dina(n32234), .dinb(n32231), .dout(n32235));
  jand g14973(.dina(n32232), .dinb(n31824), .dout(n32236));
  jand g14974(.dina(n31825), .dinb(n309), .dout(n32237));
  jand g14975(.dina(n32237), .dinb(n32227), .dout(n32238));
  jor  g14976(.dina(n32238), .dinb(n32236), .dout(n32239));
  jand g14977(.dina(n32239), .dinb(n289), .dout(n32240));
  jnot g14978(.din(n32239), .dout(n32241));
  jand g14979(.dina(n32241), .dinb(b52 ), .dout(n32242));
  jnot g14980(.din(n32242), .dout(n32243));
  jand g14981(.dina(n32235), .dinb(n288), .dout(n32244));
  jor  g14982(.dina(n32230), .dinb(n31833), .dout(n32245));
  jxor g14983(.dina(n32222), .dinb(n32221), .dout(n32246));
  jor  g14984(.dina(n32246), .dinb(n32232), .dout(n32247));
  jand g14985(.dina(n32247), .dinb(n32245), .dout(n32248));
  jand g14986(.dina(n32248), .dinb(n287), .dout(n32249));
  jor  g14987(.dina(n32230), .dinb(n31838), .dout(n32250));
  jxor g14988(.dina(n32219), .dinb(n32218), .dout(n32251));
  jor  g14989(.dina(n32251), .dinb(n32232), .dout(n32252));
  jand g14990(.dina(n32252), .dinb(n32250), .dout(n32253));
  jand g14991(.dina(n32253), .dinb(n286), .dout(n32254));
  jor  g14992(.dina(n32230), .dinb(n31843), .dout(n32255));
  jxor g14993(.dina(n32216), .dinb(n32215), .dout(n32256));
  jor  g14994(.dina(n32256), .dinb(n32232), .dout(n32257));
  jand g14995(.dina(n32257), .dinb(n32255), .dout(n32258));
  jand g14996(.dina(n32258), .dinb(n285), .dout(n32259));
  jor  g14997(.dina(n32230), .dinb(n31848), .dout(n32260));
  jxor g14998(.dina(n32213), .dinb(n32212), .dout(n32261));
  jor  g14999(.dina(n32261), .dinb(n32232), .dout(n32262));
  jand g15000(.dina(n32262), .dinb(n32260), .dout(n32263));
  jand g15001(.dina(n32263), .dinb(n284), .dout(n32264));
  jor  g15002(.dina(n32230), .dinb(n31853), .dout(n32265));
  jxor g15003(.dina(n32210), .dinb(n32209), .dout(n32266));
  jor  g15004(.dina(n32266), .dinb(n32232), .dout(n32267));
  jand g15005(.dina(n32267), .dinb(n32265), .dout(n32268));
  jand g15006(.dina(n32268), .dinb(n317), .dout(n32269));
  jor  g15007(.dina(n32230), .dinb(n31858), .dout(n32270));
  jxor g15008(.dina(n32207), .dinb(n32206), .dout(n32271));
  jor  g15009(.dina(n32271), .dinb(n32232), .dout(n32272));
  jand g15010(.dina(n32272), .dinb(n32270), .dout(n32273));
  jand g15011(.dina(n32273), .dinb(n316), .dout(n32274));
  jor  g15012(.dina(n32230), .dinb(n31863), .dout(n32275));
  jxor g15013(.dina(n32204), .dinb(n32203), .dout(n32276));
  jor  g15014(.dina(n32276), .dinb(n32232), .dout(n32277));
  jand g15015(.dina(n32277), .dinb(n32275), .dout(n32278));
  jand g15016(.dina(n32278), .dinb(n315), .dout(n32279));
  jor  g15017(.dina(n32230), .dinb(n31868), .dout(n32280));
  jxor g15018(.dina(n32201), .dinb(n32200), .dout(n32281));
  jor  g15019(.dina(n32281), .dinb(n32232), .dout(n32282));
  jand g15020(.dina(n32282), .dinb(n32280), .dout(n32283));
  jand g15021(.dina(n32283), .dinb(n283), .dout(n32284));
  jor  g15022(.dina(n32230), .dinb(n31873), .dout(n32285));
  jxor g15023(.dina(n32198), .dinb(n32197), .dout(n32286));
  jor  g15024(.dina(n32286), .dinb(n32232), .dout(n32287));
  jand g15025(.dina(n32287), .dinb(n32285), .dout(n32288));
  jand g15026(.dina(n32288), .dinb(n280), .dout(n32289));
  jor  g15027(.dina(n32230), .dinb(n31878), .dout(n32290));
  jxor g15028(.dina(n32195), .dinb(n32194), .dout(n32291));
  jor  g15029(.dina(n32291), .dinb(n32232), .dout(n32292));
  jand g15030(.dina(n32292), .dinb(n32290), .dout(n32293));
  jand g15031(.dina(n32293), .dinb(n279), .dout(n32294));
  jor  g15032(.dina(n32230), .dinb(n31883), .dout(n32295));
  jxor g15033(.dina(n32192), .dinb(n32191), .dout(n32296));
  jor  g15034(.dina(n32296), .dinb(n32232), .dout(n32297));
  jand g15035(.dina(n32297), .dinb(n32295), .dout(n32298));
  jand g15036(.dina(n32298), .dinb(n278), .dout(n32299));
  jor  g15037(.dina(n32230), .dinb(n31888), .dout(n32300));
  jxor g15038(.dina(n32189), .dinb(n32188), .dout(n32301));
  jor  g15039(.dina(n32301), .dinb(n32232), .dout(n32302));
  jand g15040(.dina(n32302), .dinb(n32300), .dout(n32303));
  jand g15041(.dina(n32303), .dinb(n277), .dout(n32304));
  jor  g15042(.dina(n32230), .dinb(n31893), .dout(n32305));
  jxor g15043(.dina(n32186), .dinb(n32185), .dout(n32306));
  jor  g15044(.dina(n32306), .dinb(n32232), .dout(n32307));
  jand g15045(.dina(n32307), .dinb(n32305), .dout(n32308));
  jand g15046(.dina(n32308), .dinb(n326), .dout(n32309));
  jor  g15047(.dina(n32230), .dinb(n31898), .dout(n32310));
  jxor g15048(.dina(n32183), .dinb(n32182), .dout(n32311));
  jor  g15049(.dina(n32311), .dinb(n32232), .dout(n32312));
  jand g15050(.dina(n32312), .dinb(n32310), .dout(n32313));
  jand g15051(.dina(n32313), .dinb(n325), .dout(n32314));
  jor  g15052(.dina(n32230), .dinb(n31903), .dout(n32315));
  jxor g15053(.dina(n32180), .dinb(n32179), .dout(n32316));
  jor  g15054(.dina(n32316), .dinb(n32232), .dout(n32317));
  jand g15055(.dina(n32317), .dinb(n32315), .dout(n32318));
  jand g15056(.dina(n32318), .dinb(n324), .dout(n32319));
  jor  g15057(.dina(n32230), .dinb(n31908), .dout(n32320));
  jxor g15058(.dina(n32177), .dinb(n32176), .dout(n32321));
  jor  g15059(.dina(n32321), .dinb(n32232), .dout(n32322));
  jand g15060(.dina(n32322), .dinb(n32320), .dout(n32323));
  jand g15061(.dina(n32323), .dinb(n276), .dout(n32324));
  jor  g15062(.dina(n32230), .dinb(n31913), .dout(n32325));
  jxor g15063(.dina(n32174), .dinb(n32173), .dout(n32326));
  jor  g15064(.dina(n32326), .dinb(n32232), .dout(n32327));
  jand g15065(.dina(n32327), .dinb(n32325), .dout(n32328));
  jand g15066(.dina(n32328), .dinb(n333), .dout(n32329));
  jor  g15067(.dina(n32230), .dinb(n31918), .dout(n32330));
  jxor g15068(.dina(n32171), .dinb(n32170), .dout(n32331));
  jor  g15069(.dina(n32331), .dinb(n32232), .dout(n32332));
  jand g15070(.dina(n32332), .dinb(n32330), .dout(n32333));
  jand g15071(.dina(n32333), .dinb(n332), .dout(n32334));
  jor  g15072(.dina(n32230), .dinb(n31923), .dout(n32335));
  jxor g15073(.dina(n32168), .dinb(n32167), .dout(n32336));
  jor  g15074(.dina(n32336), .dinb(n32232), .dout(n32337));
  jand g15075(.dina(n32337), .dinb(n32335), .dout(n32338));
  jand g15076(.dina(n32338), .dinb(n331), .dout(n32339));
  jor  g15077(.dina(n32230), .dinb(n31928), .dout(n32340));
  jxor g15078(.dina(n32165), .dinb(n32164), .dout(n32341));
  jor  g15079(.dina(n32341), .dinb(n32232), .dout(n32342));
  jand g15080(.dina(n32342), .dinb(n32340), .dout(n32343));
  jand g15081(.dina(n32343), .dinb(n275), .dout(n32344));
  jor  g15082(.dina(n32230), .dinb(n31933), .dout(n32345));
  jxor g15083(.dina(n32162), .dinb(n32161), .dout(n32346));
  jor  g15084(.dina(n32346), .dinb(n32232), .dout(n32347));
  jand g15085(.dina(n32347), .dinb(n32345), .dout(n32348));
  jand g15086(.dina(n32348), .dinb(n340), .dout(n32349));
  jor  g15087(.dina(n32230), .dinb(n31938), .dout(n32350));
  jxor g15088(.dina(n32159), .dinb(n32158), .dout(n32351));
  jor  g15089(.dina(n32351), .dinb(n32232), .dout(n32352));
  jand g15090(.dina(n32352), .dinb(n32350), .dout(n32353));
  jand g15091(.dina(n32353), .dinb(n339), .dout(n32354));
  jor  g15092(.dina(n32230), .dinb(n31943), .dout(n32355));
  jxor g15093(.dina(n32156), .dinb(n32155), .dout(n32356));
  jor  g15094(.dina(n32356), .dinb(n32232), .dout(n32357));
  jand g15095(.dina(n32357), .dinb(n32355), .dout(n32358));
  jand g15096(.dina(n32358), .dinb(n338), .dout(n32359));
  jor  g15097(.dina(n32230), .dinb(n31948), .dout(n32360));
  jxor g15098(.dina(n32153), .dinb(n32152), .dout(n32361));
  jor  g15099(.dina(n32361), .dinb(n32232), .dout(n32362));
  jand g15100(.dina(n32362), .dinb(n32360), .dout(n32363));
  jand g15101(.dina(n32363), .dinb(n271), .dout(n32364));
  jor  g15102(.dina(n32230), .dinb(n31953), .dout(n32365));
  jxor g15103(.dina(n32150), .dinb(n32149), .dout(n32366));
  jor  g15104(.dina(n32366), .dinb(n32232), .dout(n32367));
  jand g15105(.dina(n32367), .dinb(n32365), .dout(n32368));
  jand g15106(.dina(n32368), .dinb(n270), .dout(n32369));
  jor  g15107(.dina(n32230), .dinb(n31958), .dout(n32370));
  jxor g15108(.dina(n32147), .dinb(n32146), .dout(n32371));
  jor  g15109(.dina(n32371), .dinb(n32232), .dout(n32372));
  jand g15110(.dina(n32372), .dinb(n32370), .dout(n32373));
  jand g15111(.dina(n32373), .dinb(n269), .dout(n32374));
  jor  g15112(.dina(n32230), .dinb(n31963), .dout(n32375));
  jxor g15113(.dina(n32144), .dinb(n32143), .dout(n32376));
  jor  g15114(.dina(n32376), .dinb(n32232), .dout(n32377));
  jand g15115(.dina(n32377), .dinb(n32375), .dout(n32378));
  jand g15116(.dina(n32378), .dinb(n274), .dout(n32379));
  jor  g15117(.dina(n32230), .dinb(n31968), .dout(n32380));
  jxor g15118(.dina(n32141), .dinb(n32140), .dout(n32381));
  jor  g15119(.dina(n32381), .dinb(n32232), .dout(n32382));
  jand g15120(.dina(n32382), .dinb(n32380), .dout(n32383));
  jand g15121(.dina(n32383), .dinb(n268), .dout(n32384));
  jor  g15122(.dina(n32230), .dinb(n31973), .dout(n32385));
  jxor g15123(.dina(n32138), .dinb(n32137), .dout(n32386));
  jor  g15124(.dina(n32386), .dinb(n32232), .dout(n32387));
  jand g15125(.dina(n32387), .dinb(n32385), .dout(n32388));
  jand g15126(.dina(n32388), .dinb(n349), .dout(n32389));
  jor  g15127(.dina(n32230), .dinb(n31978), .dout(n32390));
  jxor g15128(.dina(n32135), .dinb(n32134), .dout(n32391));
  jor  g15129(.dina(n32391), .dinb(n32232), .dout(n32392));
  jand g15130(.dina(n32392), .dinb(n32390), .dout(n32393));
  jand g15131(.dina(n32393), .dinb(n348), .dout(n32394));
  jor  g15132(.dina(n32230), .dinb(n31983), .dout(n32395));
  jxor g15133(.dina(n32132), .dinb(n32131), .dout(n32396));
  jor  g15134(.dina(n32396), .dinb(n32232), .dout(n32397));
  jand g15135(.dina(n32397), .dinb(n32395), .dout(n32398));
  jand g15136(.dina(n32398), .dinb(n347), .dout(n32399));
  jor  g15137(.dina(n32230), .dinb(n31988), .dout(n32400));
  jxor g15138(.dina(n32129), .dinb(n32128), .dout(n32401));
  jor  g15139(.dina(n32401), .dinb(n32232), .dout(n32402));
  jand g15140(.dina(n32402), .dinb(n32400), .dout(n32403));
  jand g15141(.dina(n32403), .dinb(n267), .dout(n32404));
  jor  g15142(.dina(n32230), .dinb(n31993), .dout(n32405));
  jxor g15143(.dina(n32126), .dinb(n32125), .dout(n32406));
  jor  g15144(.dina(n32406), .dinb(n32232), .dout(n32407));
  jand g15145(.dina(n32407), .dinb(n32405), .dout(n32408));
  jand g15146(.dina(n32408), .dinb(n266), .dout(n32409));
  jor  g15147(.dina(n32230), .dinb(n31998), .dout(n32410));
  jxor g15148(.dina(n32123), .dinb(n32122), .dout(n32411));
  jor  g15149(.dina(n32411), .dinb(n32232), .dout(n32412));
  jand g15150(.dina(n32412), .dinb(n32410), .dout(n32413));
  jand g15151(.dina(n32413), .dinb(n356), .dout(n32414));
  jor  g15152(.dina(n32230), .dinb(n32003), .dout(n32415));
  jxor g15153(.dina(n32120), .dinb(n32119), .dout(n32416));
  jor  g15154(.dina(n32416), .dinb(n32232), .dout(n32417));
  jand g15155(.dina(n32417), .dinb(n32415), .dout(n32418));
  jand g15156(.dina(n32418), .dinb(n355), .dout(n32419));
  jor  g15157(.dina(n32230), .dinb(n32008), .dout(n32420));
  jxor g15158(.dina(n32117), .dinb(n32116), .dout(n32421));
  jor  g15159(.dina(n32421), .dinb(n32232), .dout(n32422));
  jand g15160(.dina(n32422), .dinb(n32420), .dout(n32423));
  jand g15161(.dina(n32423), .dinb(n364), .dout(n32424));
  jor  g15162(.dina(n32230), .dinb(n32013), .dout(n32425));
  jxor g15163(.dina(n32114), .dinb(n32113), .dout(n32426));
  jor  g15164(.dina(n32426), .dinb(n32232), .dout(n32427));
  jand g15165(.dina(n32427), .dinb(n32425), .dout(n32428));
  jand g15166(.dina(n32428), .dinb(n361), .dout(n32429));
  jor  g15167(.dina(n32230), .dinb(n32018), .dout(n32430));
  jxor g15168(.dina(n32111), .dinb(n32110), .dout(n32431));
  jor  g15169(.dina(n32431), .dinb(n32232), .dout(n32432));
  jand g15170(.dina(n32432), .dinb(n32430), .dout(n32433));
  jand g15171(.dina(n32433), .dinb(n360), .dout(n32434));
  jor  g15172(.dina(n32230), .dinb(n32023), .dout(n32435));
  jxor g15173(.dina(n32108), .dinb(n32107), .dout(n32436));
  jor  g15174(.dina(n32436), .dinb(n32232), .dout(n32437));
  jand g15175(.dina(n32437), .dinb(n32435), .dout(n32438));
  jand g15176(.dina(n32438), .dinb(n363), .dout(n32439));
  jor  g15177(.dina(n32230), .dinb(n32028), .dout(n32440));
  jxor g15178(.dina(n32105), .dinb(n32104), .dout(n32441));
  jor  g15179(.dina(n32441), .dinb(n32232), .dout(n32442));
  jand g15180(.dina(n32442), .dinb(n32440), .dout(n32443));
  jand g15181(.dina(n32443), .dinb(n359), .dout(n32444));
  jor  g15182(.dina(n32230), .dinb(n32033), .dout(n32445));
  jxor g15183(.dina(n32102), .dinb(n32101), .dout(n32446));
  jor  g15184(.dina(n32446), .dinb(n32232), .dout(n32447));
  jand g15185(.dina(n32447), .dinb(n32445), .dout(n32448));
  jand g15186(.dina(n32448), .dinb(n369), .dout(n32449));
  jor  g15187(.dina(n32230), .dinb(n32038), .dout(n32450));
  jxor g15188(.dina(n32099), .dinb(n32098), .dout(n32451));
  jor  g15189(.dina(n32451), .dinb(n32232), .dout(n32452));
  jand g15190(.dina(n32452), .dinb(n32450), .dout(n32453));
  jand g15191(.dina(n32453), .dinb(n368), .dout(n32454));
  jor  g15192(.dina(n32230), .dinb(n32043), .dout(n32455));
  jxor g15193(.dina(n32096), .dinb(n32095), .dout(n32456));
  jor  g15194(.dina(n32456), .dinb(n32232), .dout(n32457));
  jand g15195(.dina(n32457), .dinb(n32455), .dout(n32458));
  jand g15196(.dina(n32458), .dinb(n367), .dout(n32459));
  jor  g15197(.dina(n32230), .dinb(n32048), .dout(n32460));
  jxor g15198(.dina(n32093), .dinb(n32092), .dout(n32461));
  jor  g15199(.dina(n32461), .dinb(n32232), .dout(n32462));
  jand g15200(.dina(n32462), .dinb(n32460), .dout(n32463));
  jand g15201(.dina(n32463), .dinb(n265), .dout(n32464));
  jor  g15202(.dina(n32230), .dinb(n32053), .dout(n32465));
  jxor g15203(.dina(n32090), .dinb(n32089), .dout(n32466));
  jor  g15204(.dina(n32466), .dinb(n32232), .dout(n32467));
  jand g15205(.dina(n32467), .dinb(n32465), .dout(n32468));
  jand g15206(.dina(n32468), .dinb(n378), .dout(n32469));
  jor  g15207(.dina(n32230), .dinb(n32058), .dout(n32470));
  jxor g15208(.dina(n32087), .dinb(n32086), .dout(n32471));
  jor  g15209(.dina(n32471), .dinb(n32232), .dout(n32472));
  jand g15210(.dina(n32472), .dinb(n32470), .dout(n32473));
  jand g15211(.dina(n32473), .dinb(n377), .dout(n32474));
  jand g15212(.dina(n32232), .dinb(n32064), .dout(n32475));
  jnot g15213(.din(n32475), .dout(n32476));
  jxor g15214(.dina(n32084), .dinb(n32083), .dout(n32477));
  jor  g15215(.dina(n32477), .dinb(n32232), .dout(n32478));
  jand g15216(.dina(n32478), .dinb(n32476), .dout(n32479));
  jand g15217(.dina(n32479), .dinb(n376), .dout(n32480));
  jor  g15218(.dina(n32230), .dinb(n32072), .dout(n32481));
  jxor g15219(.dina(n32081), .dinb(n32080), .dout(n32482));
  jor  g15220(.dina(n32482), .dinb(n32232), .dout(n32483));
  jand g15221(.dina(n32483), .dinb(n32481), .dout(n32484));
  jand g15222(.dina(n32484), .dinb(n264), .dout(n32485));
  jor  g15223(.dina(n32230), .dinb(n32077), .dout(n32486));
  jxor g15224(.dina(n32078), .dinb(n12017), .dout(n32487));
  jand g15225(.dina(n32487), .dinb(n32230), .dout(n32488));
  jnot g15226(.din(n32488), .dout(n32489));
  jand g15227(.dina(n32489), .dinb(n32486), .dout(n32490));
  jnot g15228(.din(n32490), .dout(n32491));
  jand g15229(.dina(n32491), .dinb(n386), .dout(n32492));
  jnot g15230(.din(n12427), .dout(n32493));
  jnot g15231(.din(n31825), .dout(n32494));
  jnot g15232(.din(n31829), .dout(n32495));
  jnot g15233(.din(n31834), .dout(n32496));
  jnot g15234(.din(n31839), .dout(n32497));
  jnot g15235(.din(n31844), .dout(n32498));
  jnot g15236(.din(n31849), .dout(n32499));
  jnot g15237(.din(n31854), .dout(n32500));
  jnot g15238(.din(n31859), .dout(n32501));
  jnot g15239(.din(n31864), .dout(n32502));
  jnot g15240(.din(n31869), .dout(n32503));
  jnot g15241(.din(n31874), .dout(n32504));
  jnot g15242(.din(n31879), .dout(n32505));
  jnot g15243(.din(n31884), .dout(n32506));
  jnot g15244(.din(n31889), .dout(n32507));
  jnot g15245(.din(n31894), .dout(n32508));
  jnot g15246(.din(n31899), .dout(n32509));
  jnot g15247(.din(n31904), .dout(n32510));
  jnot g15248(.din(n31909), .dout(n32511));
  jnot g15249(.din(n31914), .dout(n32512));
  jnot g15250(.din(n31919), .dout(n32513));
  jnot g15251(.din(n31924), .dout(n32514));
  jnot g15252(.din(n31929), .dout(n32515));
  jnot g15253(.din(n31934), .dout(n32516));
  jnot g15254(.din(n31939), .dout(n32517));
  jnot g15255(.din(n31944), .dout(n32518));
  jnot g15256(.din(n31949), .dout(n32519));
  jnot g15257(.din(n31954), .dout(n32520));
  jnot g15258(.din(n31959), .dout(n32521));
  jnot g15259(.din(n31964), .dout(n32522));
  jnot g15260(.din(n31969), .dout(n32523));
  jnot g15261(.din(n31974), .dout(n32524));
  jnot g15262(.din(n31979), .dout(n32525));
  jnot g15263(.din(n31984), .dout(n32526));
  jnot g15264(.din(n31989), .dout(n32527));
  jnot g15265(.din(n31994), .dout(n32528));
  jnot g15266(.din(n31999), .dout(n32529));
  jnot g15267(.din(n32004), .dout(n32530));
  jnot g15268(.din(n32009), .dout(n32531));
  jnot g15269(.din(n32014), .dout(n32532));
  jnot g15270(.din(n32019), .dout(n32533));
  jnot g15271(.din(n32024), .dout(n32534));
  jnot g15272(.din(n32029), .dout(n32535));
  jnot g15273(.din(n32034), .dout(n32536));
  jnot g15274(.din(n32039), .dout(n32537));
  jnot g15275(.din(n32044), .dout(n32538));
  jnot g15276(.din(n32049), .dout(n32539));
  jnot g15277(.din(n32054), .dout(n32540));
  jnot g15278(.din(n32059), .dout(n32541));
  jnot g15279(.din(n32066), .dout(n32542));
  jnot g15280(.din(n32073), .dout(n32543));
  jnot g15281(.din(n32076), .dout(n32544));
  jxor g15282(.dina(n32077), .dinb(n259), .dout(n32545));
  jor  g15283(.dina(n32545), .dinb(n12016), .dout(n32546));
  jand g15284(.dina(n32546), .dinb(n32544), .dout(n32547));
  jnot g15285(.din(n32081), .dout(n32548));
  jor  g15286(.dina(n32548), .dinb(n32547), .dout(n32549));
  jand g15287(.dina(n32549), .dinb(n32543), .dout(n32550));
  jnot g15288(.din(n32084), .dout(n32551));
  jor  g15289(.dina(n32551), .dinb(n32550), .dout(n32552));
  jand g15290(.dina(n32552), .dinb(n32542), .dout(n32553));
  jnot g15291(.din(n32087), .dout(n32554));
  jor  g15292(.dina(n32554), .dinb(n32553), .dout(n32555));
  jand g15293(.dina(n32555), .dinb(n32541), .dout(n32556));
  jnot g15294(.din(n32090), .dout(n32557));
  jor  g15295(.dina(n32557), .dinb(n32556), .dout(n32558));
  jand g15296(.dina(n32558), .dinb(n32540), .dout(n32559));
  jnot g15297(.din(n32093), .dout(n32560));
  jor  g15298(.dina(n32560), .dinb(n32559), .dout(n32561));
  jand g15299(.dina(n32561), .dinb(n32539), .dout(n32562));
  jnot g15300(.din(n32096), .dout(n32563));
  jor  g15301(.dina(n32563), .dinb(n32562), .dout(n32564));
  jand g15302(.dina(n32564), .dinb(n32538), .dout(n32565));
  jnot g15303(.din(n32099), .dout(n32566));
  jor  g15304(.dina(n32566), .dinb(n32565), .dout(n32567));
  jand g15305(.dina(n32567), .dinb(n32537), .dout(n32568));
  jnot g15306(.din(n32102), .dout(n32569));
  jor  g15307(.dina(n32569), .dinb(n32568), .dout(n32570));
  jand g15308(.dina(n32570), .dinb(n32536), .dout(n32571));
  jnot g15309(.din(n32105), .dout(n32572));
  jor  g15310(.dina(n32572), .dinb(n32571), .dout(n32573));
  jand g15311(.dina(n32573), .dinb(n32535), .dout(n32574));
  jnot g15312(.din(n32108), .dout(n32575));
  jor  g15313(.dina(n32575), .dinb(n32574), .dout(n32576));
  jand g15314(.dina(n32576), .dinb(n32534), .dout(n32577));
  jnot g15315(.din(n32111), .dout(n32578));
  jor  g15316(.dina(n32578), .dinb(n32577), .dout(n32579));
  jand g15317(.dina(n32579), .dinb(n32533), .dout(n32580));
  jnot g15318(.din(n32114), .dout(n32581));
  jor  g15319(.dina(n32581), .dinb(n32580), .dout(n32582));
  jand g15320(.dina(n32582), .dinb(n32532), .dout(n32583));
  jnot g15321(.din(n32117), .dout(n32584));
  jor  g15322(.dina(n32584), .dinb(n32583), .dout(n32585));
  jand g15323(.dina(n32585), .dinb(n32531), .dout(n32586));
  jnot g15324(.din(n32120), .dout(n32587));
  jor  g15325(.dina(n32587), .dinb(n32586), .dout(n32588));
  jand g15326(.dina(n32588), .dinb(n32530), .dout(n32589));
  jnot g15327(.din(n32123), .dout(n32590));
  jor  g15328(.dina(n32590), .dinb(n32589), .dout(n32591));
  jand g15329(.dina(n32591), .dinb(n32529), .dout(n32592));
  jnot g15330(.din(n32126), .dout(n32593));
  jor  g15331(.dina(n32593), .dinb(n32592), .dout(n32594));
  jand g15332(.dina(n32594), .dinb(n32528), .dout(n32595));
  jnot g15333(.din(n32129), .dout(n32596));
  jor  g15334(.dina(n32596), .dinb(n32595), .dout(n32597));
  jand g15335(.dina(n32597), .dinb(n32527), .dout(n32598));
  jnot g15336(.din(n32132), .dout(n32599));
  jor  g15337(.dina(n32599), .dinb(n32598), .dout(n32600));
  jand g15338(.dina(n32600), .dinb(n32526), .dout(n32601));
  jnot g15339(.din(n32135), .dout(n32602));
  jor  g15340(.dina(n32602), .dinb(n32601), .dout(n32603));
  jand g15341(.dina(n32603), .dinb(n32525), .dout(n32604));
  jnot g15342(.din(n32138), .dout(n32605));
  jor  g15343(.dina(n32605), .dinb(n32604), .dout(n32606));
  jand g15344(.dina(n32606), .dinb(n32524), .dout(n32607));
  jnot g15345(.din(n32141), .dout(n32608));
  jor  g15346(.dina(n32608), .dinb(n32607), .dout(n32609));
  jand g15347(.dina(n32609), .dinb(n32523), .dout(n32610));
  jnot g15348(.din(n32144), .dout(n32611));
  jor  g15349(.dina(n32611), .dinb(n32610), .dout(n32612));
  jand g15350(.dina(n32612), .dinb(n32522), .dout(n32613));
  jnot g15351(.din(n32147), .dout(n32614));
  jor  g15352(.dina(n32614), .dinb(n32613), .dout(n32615));
  jand g15353(.dina(n32615), .dinb(n32521), .dout(n32616));
  jnot g15354(.din(n32150), .dout(n32617));
  jor  g15355(.dina(n32617), .dinb(n32616), .dout(n32618));
  jand g15356(.dina(n32618), .dinb(n32520), .dout(n32619));
  jnot g15357(.din(n32153), .dout(n32620));
  jor  g15358(.dina(n32620), .dinb(n32619), .dout(n32621));
  jand g15359(.dina(n32621), .dinb(n32519), .dout(n32622));
  jnot g15360(.din(n32156), .dout(n32623));
  jor  g15361(.dina(n32623), .dinb(n32622), .dout(n32624));
  jand g15362(.dina(n32624), .dinb(n32518), .dout(n32625));
  jnot g15363(.din(n32159), .dout(n32626));
  jor  g15364(.dina(n32626), .dinb(n32625), .dout(n32627));
  jand g15365(.dina(n32627), .dinb(n32517), .dout(n32628));
  jnot g15366(.din(n32162), .dout(n32629));
  jor  g15367(.dina(n32629), .dinb(n32628), .dout(n32630));
  jand g15368(.dina(n32630), .dinb(n32516), .dout(n32631));
  jnot g15369(.din(n32165), .dout(n32632));
  jor  g15370(.dina(n32632), .dinb(n32631), .dout(n32633));
  jand g15371(.dina(n32633), .dinb(n32515), .dout(n32634));
  jnot g15372(.din(n32168), .dout(n32635));
  jor  g15373(.dina(n32635), .dinb(n32634), .dout(n32636));
  jand g15374(.dina(n32636), .dinb(n32514), .dout(n32637));
  jnot g15375(.din(n32171), .dout(n32638));
  jor  g15376(.dina(n32638), .dinb(n32637), .dout(n32639));
  jand g15377(.dina(n32639), .dinb(n32513), .dout(n32640));
  jnot g15378(.din(n32174), .dout(n32641));
  jor  g15379(.dina(n32641), .dinb(n32640), .dout(n32642));
  jand g15380(.dina(n32642), .dinb(n32512), .dout(n32643));
  jnot g15381(.din(n32177), .dout(n32644));
  jor  g15382(.dina(n32644), .dinb(n32643), .dout(n32645));
  jand g15383(.dina(n32645), .dinb(n32511), .dout(n32646));
  jnot g15384(.din(n32180), .dout(n32647));
  jor  g15385(.dina(n32647), .dinb(n32646), .dout(n32648));
  jand g15386(.dina(n32648), .dinb(n32510), .dout(n32649));
  jnot g15387(.din(n32183), .dout(n32650));
  jor  g15388(.dina(n32650), .dinb(n32649), .dout(n32651));
  jand g15389(.dina(n32651), .dinb(n32509), .dout(n32652));
  jnot g15390(.din(n32186), .dout(n32653));
  jor  g15391(.dina(n32653), .dinb(n32652), .dout(n32654));
  jand g15392(.dina(n32654), .dinb(n32508), .dout(n32655));
  jnot g15393(.din(n32189), .dout(n32656));
  jor  g15394(.dina(n32656), .dinb(n32655), .dout(n32657));
  jand g15395(.dina(n32657), .dinb(n32507), .dout(n32658));
  jnot g15396(.din(n32192), .dout(n32659));
  jor  g15397(.dina(n32659), .dinb(n32658), .dout(n32660));
  jand g15398(.dina(n32660), .dinb(n32506), .dout(n32661));
  jnot g15399(.din(n32195), .dout(n32662));
  jor  g15400(.dina(n32662), .dinb(n32661), .dout(n32663));
  jand g15401(.dina(n32663), .dinb(n32505), .dout(n32664));
  jnot g15402(.din(n32198), .dout(n32665));
  jor  g15403(.dina(n32665), .dinb(n32664), .dout(n32666));
  jand g15404(.dina(n32666), .dinb(n32504), .dout(n32667));
  jnot g15405(.din(n32201), .dout(n32668));
  jor  g15406(.dina(n32668), .dinb(n32667), .dout(n32669));
  jand g15407(.dina(n32669), .dinb(n32503), .dout(n32670));
  jnot g15408(.din(n32204), .dout(n32671));
  jor  g15409(.dina(n32671), .dinb(n32670), .dout(n32672));
  jand g15410(.dina(n32672), .dinb(n32502), .dout(n32673));
  jnot g15411(.din(n32207), .dout(n32674));
  jor  g15412(.dina(n32674), .dinb(n32673), .dout(n32675));
  jand g15413(.dina(n32675), .dinb(n32501), .dout(n32676));
  jnot g15414(.din(n32210), .dout(n32677));
  jor  g15415(.dina(n32677), .dinb(n32676), .dout(n32678));
  jand g15416(.dina(n32678), .dinb(n32500), .dout(n32679));
  jnot g15417(.din(n32213), .dout(n32680));
  jor  g15418(.dina(n32680), .dinb(n32679), .dout(n32681));
  jand g15419(.dina(n32681), .dinb(n32499), .dout(n32682));
  jnot g15420(.din(n32216), .dout(n32683));
  jor  g15421(.dina(n32683), .dinb(n32682), .dout(n32684));
  jand g15422(.dina(n32684), .dinb(n32498), .dout(n32685));
  jnot g15423(.din(n32219), .dout(n32686));
  jor  g15424(.dina(n32686), .dinb(n32685), .dout(n32687));
  jand g15425(.dina(n32687), .dinb(n32497), .dout(n32688));
  jnot g15426(.din(n32222), .dout(n32689));
  jor  g15427(.dina(n32689), .dinb(n32688), .dout(n32690));
  jand g15428(.dina(n32690), .dinb(n32496), .dout(n32691));
  jnot g15429(.din(n32225), .dout(n32692));
  jor  g15430(.dina(n32692), .dinb(n32691), .dout(n32693));
  jand g15431(.dina(n32693), .dinb(n32495), .dout(n32694));
  jor  g15432(.dina(n32694), .dinb(n31827), .dout(n32695));
  jand g15433(.dina(n32695), .dinb(n32494), .dout(n32696));
  jor  g15434(.dina(n32696), .dinb(n32493), .dout(n32697));
  jand g15435(.dina(n32697), .dinb(a12 ), .dout(n32698));
  jnot g15436(.din(n12430), .dout(n32699));
  jor  g15437(.dina(n32696), .dinb(n32699), .dout(n32700));
  jnot g15438(.din(n32700), .dout(n32701));
  jor  g15439(.dina(n32701), .dinb(n32698), .dout(n32702));
  jand g15440(.dina(n32702), .dinb(n259), .dout(n32703));
  jand g15441(.dina(n32229), .dinb(n12427), .dout(n32704));
  jor  g15442(.dina(n32704), .dinb(n12015), .dout(n32705));
  jand g15443(.dina(n32700), .dinb(n32705), .dout(n32706));
  jxor g15444(.dina(n32706), .dinb(b1 ), .dout(n32707));
  jand g15445(.dina(n32707), .dinb(n12438), .dout(n32708));
  jor  g15446(.dina(n32708), .dinb(n32703), .dout(n32709));
  jxor g15447(.dina(n32490), .dinb(b2 ), .dout(n32710));
  jand g15448(.dina(n32710), .dinb(n32709), .dout(n32711));
  jor  g15449(.dina(n32711), .dinb(n32492), .dout(n32712));
  jxor g15450(.dina(n32484), .dinb(n264), .dout(n32713));
  jand g15451(.dina(n32713), .dinb(n32712), .dout(n32714));
  jor  g15452(.dina(n32714), .dinb(n32485), .dout(n32715));
  jxor g15453(.dina(n32479), .dinb(n376), .dout(n32716));
  jand g15454(.dina(n32716), .dinb(n32715), .dout(n32717));
  jor  g15455(.dina(n32717), .dinb(n32480), .dout(n32718));
  jxor g15456(.dina(n32473), .dinb(n377), .dout(n32719));
  jand g15457(.dina(n32719), .dinb(n32718), .dout(n32720));
  jor  g15458(.dina(n32720), .dinb(n32474), .dout(n32721));
  jxor g15459(.dina(n32468), .dinb(n378), .dout(n32722));
  jand g15460(.dina(n32722), .dinb(n32721), .dout(n32723));
  jor  g15461(.dina(n32723), .dinb(n32469), .dout(n32724));
  jxor g15462(.dina(n32463), .dinb(n265), .dout(n32725));
  jand g15463(.dina(n32725), .dinb(n32724), .dout(n32726));
  jor  g15464(.dina(n32726), .dinb(n32464), .dout(n32727));
  jxor g15465(.dina(n32458), .dinb(n367), .dout(n32728));
  jand g15466(.dina(n32728), .dinb(n32727), .dout(n32729));
  jor  g15467(.dina(n32729), .dinb(n32459), .dout(n32730));
  jxor g15468(.dina(n32453), .dinb(n368), .dout(n32731));
  jand g15469(.dina(n32731), .dinb(n32730), .dout(n32732));
  jor  g15470(.dina(n32732), .dinb(n32454), .dout(n32733));
  jxor g15471(.dina(n32448), .dinb(n369), .dout(n32734));
  jand g15472(.dina(n32734), .dinb(n32733), .dout(n32735));
  jor  g15473(.dina(n32735), .dinb(n32449), .dout(n32736));
  jxor g15474(.dina(n32443), .dinb(n359), .dout(n32737));
  jand g15475(.dina(n32737), .dinb(n32736), .dout(n32738));
  jor  g15476(.dina(n32738), .dinb(n32444), .dout(n32739));
  jxor g15477(.dina(n32438), .dinb(n363), .dout(n32740));
  jand g15478(.dina(n32740), .dinb(n32739), .dout(n32741));
  jor  g15479(.dina(n32741), .dinb(n32439), .dout(n32742));
  jxor g15480(.dina(n32433), .dinb(n360), .dout(n32743));
  jand g15481(.dina(n32743), .dinb(n32742), .dout(n32744));
  jor  g15482(.dina(n32744), .dinb(n32434), .dout(n32745));
  jxor g15483(.dina(n32428), .dinb(n361), .dout(n32746));
  jand g15484(.dina(n32746), .dinb(n32745), .dout(n32747));
  jor  g15485(.dina(n32747), .dinb(n32429), .dout(n32748));
  jxor g15486(.dina(n32423), .dinb(n364), .dout(n32749));
  jand g15487(.dina(n32749), .dinb(n32748), .dout(n32750));
  jor  g15488(.dina(n32750), .dinb(n32424), .dout(n32751));
  jxor g15489(.dina(n32418), .dinb(n355), .dout(n32752));
  jand g15490(.dina(n32752), .dinb(n32751), .dout(n32753));
  jor  g15491(.dina(n32753), .dinb(n32419), .dout(n32754));
  jxor g15492(.dina(n32413), .dinb(n356), .dout(n32755));
  jand g15493(.dina(n32755), .dinb(n32754), .dout(n32756));
  jor  g15494(.dina(n32756), .dinb(n32414), .dout(n32757));
  jxor g15495(.dina(n32408), .dinb(n266), .dout(n32758));
  jand g15496(.dina(n32758), .dinb(n32757), .dout(n32759));
  jor  g15497(.dina(n32759), .dinb(n32409), .dout(n32760));
  jxor g15498(.dina(n32403), .dinb(n267), .dout(n32761));
  jand g15499(.dina(n32761), .dinb(n32760), .dout(n32762));
  jor  g15500(.dina(n32762), .dinb(n32404), .dout(n32763));
  jxor g15501(.dina(n32398), .dinb(n347), .dout(n32764));
  jand g15502(.dina(n32764), .dinb(n32763), .dout(n32765));
  jor  g15503(.dina(n32765), .dinb(n32399), .dout(n32766));
  jxor g15504(.dina(n32393), .dinb(n348), .dout(n32767));
  jand g15505(.dina(n32767), .dinb(n32766), .dout(n32768));
  jor  g15506(.dina(n32768), .dinb(n32394), .dout(n32769));
  jxor g15507(.dina(n32388), .dinb(n349), .dout(n32770));
  jand g15508(.dina(n32770), .dinb(n32769), .dout(n32771));
  jor  g15509(.dina(n32771), .dinb(n32389), .dout(n32772));
  jxor g15510(.dina(n32383), .dinb(n268), .dout(n32773));
  jand g15511(.dina(n32773), .dinb(n32772), .dout(n32774));
  jor  g15512(.dina(n32774), .dinb(n32384), .dout(n32775));
  jxor g15513(.dina(n32378), .dinb(n274), .dout(n32776));
  jand g15514(.dina(n32776), .dinb(n32775), .dout(n32777));
  jor  g15515(.dina(n32777), .dinb(n32379), .dout(n32778));
  jxor g15516(.dina(n32373), .dinb(n269), .dout(n32779));
  jand g15517(.dina(n32779), .dinb(n32778), .dout(n32780));
  jor  g15518(.dina(n32780), .dinb(n32374), .dout(n32781));
  jxor g15519(.dina(n32368), .dinb(n270), .dout(n32782));
  jand g15520(.dina(n32782), .dinb(n32781), .dout(n32783));
  jor  g15521(.dina(n32783), .dinb(n32369), .dout(n32784));
  jxor g15522(.dina(n32363), .dinb(n271), .dout(n32785));
  jand g15523(.dina(n32785), .dinb(n32784), .dout(n32786));
  jor  g15524(.dina(n32786), .dinb(n32364), .dout(n32787));
  jxor g15525(.dina(n32358), .dinb(n338), .dout(n32788));
  jand g15526(.dina(n32788), .dinb(n32787), .dout(n32789));
  jor  g15527(.dina(n32789), .dinb(n32359), .dout(n32790));
  jxor g15528(.dina(n32353), .dinb(n339), .dout(n32791));
  jand g15529(.dina(n32791), .dinb(n32790), .dout(n32792));
  jor  g15530(.dina(n32792), .dinb(n32354), .dout(n32793));
  jxor g15531(.dina(n32348), .dinb(n340), .dout(n32794));
  jand g15532(.dina(n32794), .dinb(n32793), .dout(n32795));
  jor  g15533(.dina(n32795), .dinb(n32349), .dout(n32796));
  jxor g15534(.dina(n32343), .dinb(n275), .dout(n32797));
  jand g15535(.dina(n32797), .dinb(n32796), .dout(n32798));
  jor  g15536(.dina(n32798), .dinb(n32344), .dout(n32799));
  jxor g15537(.dina(n32338), .dinb(n331), .dout(n32800));
  jand g15538(.dina(n32800), .dinb(n32799), .dout(n32801));
  jor  g15539(.dina(n32801), .dinb(n32339), .dout(n32802));
  jxor g15540(.dina(n32333), .dinb(n332), .dout(n32803));
  jand g15541(.dina(n32803), .dinb(n32802), .dout(n32804));
  jor  g15542(.dina(n32804), .dinb(n32334), .dout(n32805));
  jxor g15543(.dina(n32328), .dinb(n333), .dout(n32806));
  jand g15544(.dina(n32806), .dinb(n32805), .dout(n32807));
  jor  g15545(.dina(n32807), .dinb(n32329), .dout(n32808));
  jxor g15546(.dina(n32323), .dinb(n276), .dout(n32809));
  jand g15547(.dina(n32809), .dinb(n32808), .dout(n32810));
  jor  g15548(.dina(n32810), .dinb(n32324), .dout(n32811));
  jxor g15549(.dina(n32318), .dinb(n324), .dout(n32812));
  jand g15550(.dina(n32812), .dinb(n32811), .dout(n32813));
  jor  g15551(.dina(n32813), .dinb(n32319), .dout(n32814));
  jxor g15552(.dina(n32313), .dinb(n325), .dout(n32815));
  jand g15553(.dina(n32815), .dinb(n32814), .dout(n32816));
  jor  g15554(.dina(n32816), .dinb(n32314), .dout(n32817));
  jxor g15555(.dina(n32308), .dinb(n326), .dout(n32818));
  jand g15556(.dina(n32818), .dinb(n32817), .dout(n32819));
  jor  g15557(.dina(n32819), .dinb(n32309), .dout(n32820));
  jxor g15558(.dina(n32303), .dinb(n277), .dout(n32821));
  jand g15559(.dina(n32821), .dinb(n32820), .dout(n32822));
  jor  g15560(.dina(n32822), .dinb(n32304), .dout(n32823));
  jxor g15561(.dina(n32298), .dinb(n278), .dout(n32824));
  jand g15562(.dina(n32824), .dinb(n32823), .dout(n32825));
  jor  g15563(.dina(n32825), .dinb(n32299), .dout(n32826));
  jxor g15564(.dina(n32293), .dinb(n279), .dout(n32827));
  jand g15565(.dina(n32827), .dinb(n32826), .dout(n32828));
  jor  g15566(.dina(n32828), .dinb(n32294), .dout(n32829));
  jxor g15567(.dina(n32288), .dinb(n280), .dout(n32830));
  jand g15568(.dina(n32830), .dinb(n32829), .dout(n32831));
  jor  g15569(.dina(n32831), .dinb(n32289), .dout(n32832));
  jxor g15570(.dina(n32283), .dinb(n283), .dout(n32833));
  jand g15571(.dina(n32833), .dinb(n32832), .dout(n32834));
  jor  g15572(.dina(n32834), .dinb(n32284), .dout(n32835));
  jxor g15573(.dina(n32278), .dinb(n315), .dout(n32836));
  jand g15574(.dina(n32836), .dinb(n32835), .dout(n32837));
  jor  g15575(.dina(n32837), .dinb(n32279), .dout(n32838));
  jxor g15576(.dina(n32273), .dinb(n316), .dout(n32839));
  jand g15577(.dina(n32839), .dinb(n32838), .dout(n32840));
  jor  g15578(.dina(n32840), .dinb(n32274), .dout(n32841));
  jxor g15579(.dina(n32268), .dinb(n317), .dout(n32842));
  jand g15580(.dina(n32842), .dinb(n32841), .dout(n32843));
  jor  g15581(.dina(n32843), .dinb(n32269), .dout(n32844));
  jxor g15582(.dina(n32263), .dinb(n284), .dout(n32845));
  jand g15583(.dina(n32845), .dinb(n32844), .dout(n32846));
  jor  g15584(.dina(n32846), .dinb(n32264), .dout(n32847));
  jxor g15585(.dina(n32258), .dinb(n285), .dout(n32848));
  jand g15586(.dina(n32848), .dinb(n32847), .dout(n32849));
  jor  g15587(.dina(n32849), .dinb(n32259), .dout(n32850));
  jxor g15588(.dina(n32253), .dinb(n286), .dout(n32851));
  jand g15589(.dina(n32851), .dinb(n32850), .dout(n32852));
  jor  g15590(.dina(n32852), .dinb(n32254), .dout(n32853));
  jxor g15591(.dina(n32248), .dinb(n287), .dout(n32854));
  jand g15592(.dina(n32854), .dinb(n32853), .dout(n32855));
  jor  g15593(.dina(n32855), .dinb(n32249), .dout(n32856));
  jxor g15594(.dina(n32235), .dinb(n288), .dout(n32857));
  jand g15595(.dina(n32857), .dinb(n32856), .dout(n32858));
  jor  g15596(.dina(n32858), .dinb(n32244), .dout(n32859));
  jand g15597(.dina(n32859), .dinb(n32243), .dout(n32860));
  jor  g15598(.dina(n32860), .dinb(n32240), .dout(n32861));
  jand g15599(.dina(n32861), .dinb(n308), .dout(n32862));
  jor  g15600(.dina(n32862), .dinb(n32235), .dout(n32863));
  jnot g15601(.din(n32862), .dout(n32864));
  jxor g15602(.dina(n32857), .dinb(n32856), .dout(n32865));
  jor  g15603(.dina(n32865), .dinb(n32864), .dout(n32866));
  jand g15604(.dina(n32866), .dinb(n32863), .dout(n32867));
  jand g15605(.dina(n32864), .dinb(n32239), .dout(n32868));
  jand g15606(.dina(n32859), .dinb(n32240), .dout(n32869));
  jor  g15607(.dina(n32869), .dinb(n32868), .dout(n32870));
  jand g15608(.dina(n32870), .dinb(n290), .dout(n32871));
  jnot g15609(.din(n32870), .dout(n32872));
  jand g15610(.dina(n32872), .dinb(b53 ), .dout(n32873));
  jnot g15611(.din(n32873), .dout(n32874));
  jand g15612(.dina(n32867), .dinb(n289), .dout(n32875));
  jor  g15613(.dina(n32862), .dinb(n32248), .dout(n32876));
  jxor g15614(.dina(n32854), .dinb(n32853), .dout(n32877));
  jor  g15615(.dina(n32877), .dinb(n32864), .dout(n32878));
  jand g15616(.dina(n32878), .dinb(n32876), .dout(n32879));
  jand g15617(.dina(n32879), .dinb(n288), .dout(n32880));
  jor  g15618(.dina(n32862), .dinb(n32253), .dout(n32881));
  jxor g15619(.dina(n32851), .dinb(n32850), .dout(n32882));
  jor  g15620(.dina(n32882), .dinb(n32864), .dout(n32883));
  jand g15621(.dina(n32883), .dinb(n32881), .dout(n32884));
  jand g15622(.dina(n32884), .dinb(n287), .dout(n32885));
  jor  g15623(.dina(n32862), .dinb(n32258), .dout(n32886));
  jxor g15624(.dina(n32848), .dinb(n32847), .dout(n32887));
  jor  g15625(.dina(n32887), .dinb(n32864), .dout(n32888));
  jand g15626(.dina(n32888), .dinb(n32886), .dout(n32889));
  jand g15627(.dina(n32889), .dinb(n286), .dout(n32890));
  jor  g15628(.dina(n32862), .dinb(n32263), .dout(n32891));
  jxor g15629(.dina(n32845), .dinb(n32844), .dout(n32892));
  jor  g15630(.dina(n32892), .dinb(n32864), .dout(n32893));
  jand g15631(.dina(n32893), .dinb(n32891), .dout(n32894));
  jand g15632(.dina(n32894), .dinb(n285), .dout(n32895));
  jor  g15633(.dina(n32862), .dinb(n32268), .dout(n32896));
  jxor g15634(.dina(n32842), .dinb(n32841), .dout(n32897));
  jor  g15635(.dina(n32897), .dinb(n32864), .dout(n32898));
  jand g15636(.dina(n32898), .dinb(n32896), .dout(n32899));
  jand g15637(.dina(n32899), .dinb(n284), .dout(n32900));
  jor  g15638(.dina(n32862), .dinb(n32273), .dout(n32901));
  jxor g15639(.dina(n32839), .dinb(n32838), .dout(n32902));
  jor  g15640(.dina(n32902), .dinb(n32864), .dout(n32903));
  jand g15641(.dina(n32903), .dinb(n32901), .dout(n32904));
  jand g15642(.dina(n32904), .dinb(n317), .dout(n32905));
  jor  g15643(.dina(n32862), .dinb(n32278), .dout(n32906));
  jxor g15644(.dina(n32836), .dinb(n32835), .dout(n32907));
  jor  g15645(.dina(n32907), .dinb(n32864), .dout(n32908));
  jand g15646(.dina(n32908), .dinb(n32906), .dout(n32909));
  jand g15647(.dina(n32909), .dinb(n316), .dout(n32910));
  jor  g15648(.dina(n32862), .dinb(n32283), .dout(n32911));
  jxor g15649(.dina(n32833), .dinb(n32832), .dout(n32912));
  jor  g15650(.dina(n32912), .dinb(n32864), .dout(n32913));
  jand g15651(.dina(n32913), .dinb(n32911), .dout(n32914));
  jand g15652(.dina(n32914), .dinb(n315), .dout(n32915));
  jor  g15653(.dina(n32862), .dinb(n32288), .dout(n32916));
  jxor g15654(.dina(n32830), .dinb(n32829), .dout(n32917));
  jor  g15655(.dina(n32917), .dinb(n32864), .dout(n32918));
  jand g15656(.dina(n32918), .dinb(n32916), .dout(n32919));
  jand g15657(.dina(n32919), .dinb(n283), .dout(n32920));
  jor  g15658(.dina(n32862), .dinb(n32293), .dout(n32921));
  jxor g15659(.dina(n32827), .dinb(n32826), .dout(n32922));
  jor  g15660(.dina(n32922), .dinb(n32864), .dout(n32923));
  jand g15661(.dina(n32923), .dinb(n32921), .dout(n32924));
  jand g15662(.dina(n32924), .dinb(n280), .dout(n32925));
  jor  g15663(.dina(n32862), .dinb(n32298), .dout(n32926));
  jxor g15664(.dina(n32824), .dinb(n32823), .dout(n32927));
  jor  g15665(.dina(n32927), .dinb(n32864), .dout(n32928));
  jand g15666(.dina(n32928), .dinb(n32926), .dout(n32929));
  jand g15667(.dina(n32929), .dinb(n279), .dout(n32930));
  jor  g15668(.dina(n32862), .dinb(n32303), .dout(n32931));
  jxor g15669(.dina(n32821), .dinb(n32820), .dout(n32932));
  jor  g15670(.dina(n32932), .dinb(n32864), .dout(n32933));
  jand g15671(.dina(n32933), .dinb(n32931), .dout(n32934));
  jand g15672(.dina(n32934), .dinb(n278), .dout(n32935));
  jor  g15673(.dina(n32862), .dinb(n32308), .dout(n32936));
  jxor g15674(.dina(n32818), .dinb(n32817), .dout(n32937));
  jor  g15675(.dina(n32937), .dinb(n32864), .dout(n32938));
  jand g15676(.dina(n32938), .dinb(n32936), .dout(n32939));
  jand g15677(.dina(n32939), .dinb(n277), .dout(n32940));
  jor  g15678(.dina(n32862), .dinb(n32313), .dout(n32941));
  jxor g15679(.dina(n32815), .dinb(n32814), .dout(n32942));
  jor  g15680(.dina(n32942), .dinb(n32864), .dout(n32943));
  jand g15681(.dina(n32943), .dinb(n32941), .dout(n32944));
  jand g15682(.dina(n32944), .dinb(n326), .dout(n32945));
  jor  g15683(.dina(n32862), .dinb(n32318), .dout(n32946));
  jxor g15684(.dina(n32812), .dinb(n32811), .dout(n32947));
  jor  g15685(.dina(n32947), .dinb(n32864), .dout(n32948));
  jand g15686(.dina(n32948), .dinb(n32946), .dout(n32949));
  jand g15687(.dina(n32949), .dinb(n325), .dout(n32950));
  jor  g15688(.dina(n32862), .dinb(n32323), .dout(n32951));
  jxor g15689(.dina(n32809), .dinb(n32808), .dout(n32952));
  jor  g15690(.dina(n32952), .dinb(n32864), .dout(n32953));
  jand g15691(.dina(n32953), .dinb(n32951), .dout(n32954));
  jand g15692(.dina(n32954), .dinb(n324), .dout(n32955));
  jor  g15693(.dina(n32862), .dinb(n32328), .dout(n32956));
  jxor g15694(.dina(n32806), .dinb(n32805), .dout(n32957));
  jor  g15695(.dina(n32957), .dinb(n32864), .dout(n32958));
  jand g15696(.dina(n32958), .dinb(n32956), .dout(n32959));
  jand g15697(.dina(n32959), .dinb(n276), .dout(n32960));
  jor  g15698(.dina(n32862), .dinb(n32333), .dout(n32961));
  jxor g15699(.dina(n32803), .dinb(n32802), .dout(n32962));
  jor  g15700(.dina(n32962), .dinb(n32864), .dout(n32963));
  jand g15701(.dina(n32963), .dinb(n32961), .dout(n32964));
  jand g15702(.dina(n32964), .dinb(n333), .dout(n32965));
  jor  g15703(.dina(n32862), .dinb(n32338), .dout(n32966));
  jxor g15704(.dina(n32800), .dinb(n32799), .dout(n32967));
  jor  g15705(.dina(n32967), .dinb(n32864), .dout(n32968));
  jand g15706(.dina(n32968), .dinb(n32966), .dout(n32969));
  jand g15707(.dina(n32969), .dinb(n332), .dout(n32970));
  jor  g15708(.dina(n32862), .dinb(n32343), .dout(n32971));
  jxor g15709(.dina(n32797), .dinb(n32796), .dout(n32972));
  jor  g15710(.dina(n32972), .dinb(n32864), .dout(n32973));
  jand g15711(.dina(n32973), .dinb(n32971), .dout(n32974));
  jand g15712(.dina(n32974), .dinb(n331), .dout(n32975));
  jor  g15713(.dina(n32862), .dinb(n32348), .dout(n32976));
  jxor g15714(.dina(n32794), .dinb(n32793), .dout(n32977));
  jor  g15715(.dina(n32977), .dinb(n32864), .dout(n32978));
  jand g15716(.dina(n32978), .dinb(n32976), .dout(n32979));
  jand g15717(.dina(n32979), .dinb(n275), .dout(n32980));
  jor  g15718(.dina(n32862), .dinb(n32353), .dout(n32981));
  jxor g15719(.dina(n32791), .dinb(n32790), .dout(n32982));
  jor  g15720(.dina(n32982), .dinb(n32864), .dout(n32983));
  jand g15721(.dina(n32983), .dinb(n32981), .dout(n32984));
  jand g15722(.dina(n32984), .dinb(n340), .dout(n32985));
  jor  g15723(.dina(n32862), .dinb(n32358), .dout(n32986));
  jxor g15724(.dina(n32788), .dinb(n32787), .dout(n32987));
  jor  g15725(.dina(n32987), .dinb(n32864), .dout(n32988));
  jand g15726(.dina(n32988), .dinb(n32986), .dout(n32989));
  jand g15727(.dina(n32989), .dinb(n339), .dout(n32990));
  jor  g15728(.dina(n32862), .dinb(n32363), .dout(n32991));
  jxor g15729(.dina(n32785), .dinb(n32784), .dout(n32992));
  jor  g15730(.dina(n32992), .dinb(n32864), .dout(n32993));
  jand g15731(.dina(n32993), .dinb(n32991), .dout(n32994));
  jand g15732(.dina(n32994), .dinb(n338), .dout(n32995));
  jor  g15733(.dina(n32862), .dinb(n32368), .dout(n32996));
  jxor g15734(.dina(n32782), .dinb(n32781), .dout(n32997));
  jor  g15735(.dina(n32997), .dinb(n32864), .dout(n32998));
  jand g15736(.dina(n32998), .dinb(n32996), .dout(n32999));
  jand g15737(.dina(n32999), .dinb(n271), .dout(n33000));
  jor  g15738(.dina(n32862), .dinb(n32373), .dout(n33001));
  jxor g15739(.dina(n32779), .dinb(n32778), .dout(n33002));
  jor  g15740(.dina(n33002), .dinb(n32864), .dout(n33003));
  jand g15741(.dina(n33003), .dinb(n33001), .dout(n33004));
  jand g15742(.dina(n33004), .dinb(n270), .dout(n33005));
  jor  g15743(.dina(n32862), .dinb(n32378), .dout(n33006));
  jxor g15744(.dina(n32776), .dinb(n32775), .dout(n33007));
  jor  g15745(.dina(n33007), .dinb(n32864), .dout(n33008));
  jand g15746(.dina(n33008), .dinb(n33006), .dout(n33009));
  jand g15747(.dina(n33009), .dinb(n269), .dout(n33010));
  jor  g15748(.dina(n32862), .dinb(n32383), .dout(n33011));
  jxor g15749(.dina(n32773), .dinb(n32772), .dout(n33012));
  jor  g15750(.dina(n33012), .dinb(n32864), .dout(n33013));
  jand g15751(.dina(n33013), .dinb(n33011), .dout(n33014));
  jand g15752(.dina(n33014), .dinb(n274), .dout(n33015));
  jor  g15753(.dina(n32862), .dinb(n32388), .dout(n33016));
  jxor g15754(.dina(n32770), .dinb(n32769), .dout(n33017));
  jor  g15755(.dina(n33017), .dinb(n32864), .dout(n33018));
  jand g15756(.dina(n33018), .dinb(n33016), .dout(n33019));
  jand g15757(.dina(n33019), .dinb(n268), .dout(n33020));
  jor  g15758(.dina(n32862), .dinb(n32393), .dout(n33021));
  jxor g15759(.dina(n32767), .dinb(n32766), .dout(n33022));
  jor  g15760(.dina(n33022), .dinb(n32864), .dout(n33023));
  jand g15761(.dina(n33023), .dinb(n33021), .dout(n33024));
  jand g15762(.dina(n33024), .dinb(n349), .dout(n33025));
  jor  g15763(.dina(n32862), .dinb(n32398), .dout(n33026));
  jxor g15764(.dina(n32764), .dinb(n32763), .dout(n33027));
  jor  g15765(.dina(n33027), .dinb(n32864), .dout(n33028));
  jand g15766(.dina(n33028), .dinb(n33026), .dout(n33029));
  jand g15767(.dina(n33029), .dinb(n348), .dout(n33030));
  jor  g15768(.dina(n32862), .dinb(n32403), .dout(n33031));
  jxor g15769(.dina(n32761), .dinb(n32760), .dout(n33032));
  jor  g15770(.dina(n33032), .dinb(n32864), .dout(n33033));
  jand g15771(.dina(n33033), .dinb(n33031), .dout(n33034));
  jand g15772(.dina(n33034), .dinb(n347), .dout(n33035));
  jor  g15773(.dina(n32862), .dinb(n32408), .dout(n33036));
  jxor g15774(.dina(n32758), .dinb(n32757), .dout(n33037));
  jor  g15775(.dina(n33037), .dinb(n32864), .dout(n33038));
  jand g15776(.dina(n33038), .dinb(n33036), .dout(n33039));
  jand g15777(.dina(n33039), .dinb(n267), .dout(n33040));
  jor  g15778(.dina(n32862), .dinb(n32413), .dout(n33041));
  jxor g15779(.dina(n32755), .dinb(n32754), .dout(n33042));
  jor  g15780(.dina(n33042), .dinb(n32864), .dout(n33043));
  jand g15781(.dina(n33043), .dinb(n33041), .dout(n33044));
  jand g15782(.dina(n33044), .dinb(n266), .dout(n33045));
  jor  g15783(.dina(n32862), .dinb(n32418), .dout(n33046));
  jxor g15784(.dina(n32752), .dinb(n32751), .dout(n33047));
  jor  g15785(.dina(n33047), .dinb(n32864), .dout(n33048));
  jand g15786(.dina(n33048), .dinb(n33046), .dout(n33049));
  jand g15787(.dina(n33049), .dinb(n356), .dout(n33050));
  jor  g15788(.dina(n32862), .dinb(n32423), .dout(n33051));
  jxor g15789(.dina(n32749), .dinb(n32748), .dout(n33052));
  jor  g15790(.dina(n33052), .dinb(n32864), .dout(n33053));
  jand g15791(.dina(n33053), .dinb(n33051), .dout(n33054));
  jand g15792(.dina(n33054), .dinb(n355), .dout(n33055));
  jor  g15793(.dina(n32862), .dinb(n32428), .dout(n33056));
  jxor g15794(.dina(n32746), .dinb(n32745), .dout(n33057));
  jor  g15795(.dina(n33057), .dinb(n32864), .dout(n33058));
  jand g15796(.dina(n33058), .dinb(n33056), .dout(n33059));
  jand g15797(.dina(n33059), .dinb(n364), .dout(n33060));
  jor  g15798(.dina(n32862), .dinb(n32433), .dout(n33061));
  jxor g15799(.dina(n32743), .dinb(n32742), .dout(n33062));
  jor  g15800(.dina(n33062), .dinb(n32864), .dout(n33063));
  jand g15801(.dina(n33063), .dinb(n33061), .dout(n33064));
  jand g15802(.dina(n33064), .dinb(n361), .dout(n33065));
  jor  g15803(.dina(n32862), .dinb(n32438), .dout(n33066));
  jxor g15804(.dina(n32740), .dinb(n32739), .dout(n33067));
  jor  g15805(.dina(n33067), .dinb(n32864), .dout(n33068));
  jand g15806(.dina(n33068), .dinb(n33066), .dout(n33069));
  jand g15807(.dina(n33069), .dinb(n360), .dout(n33070));
  jor  g15808(.dina(n32862), .dinb(n32443), .dout(n33071));
  jxor g15809(.dina(n32737), .dinb(n32736), .dout(n33072));
  jor  g15810(.dina(n33072), .dinb(n32864), .dout(n33073));
  jand g15811(.dina(n33073), .dinb(n33071), .dout(n33074));
  jand g15812(.dina(n33074), .dinb(n363), .dout(n33075));
  jor  g15813(.dina(n32862), .dinb(n32448), .dout(n33076));
  jxor g15814(.dina(n32734), .dinb(n32733), .dout(n33077));
  jor  g15815(.dina(n33077), .dinb(n32864), .dout(n33078));
  jand g15816(.dina(n33078), .dinb(n33076), .dout(n33079));
  jand g15817(.dina(n33079), .dinb(n359), .dout(n33080));
  jor  g15818(.dina(n32862), .dinb(n32453), .dout(n33081));
  jxor g15819(.dina(n32731), .dinb(n32730), .dout(n33082));
  jor  g15820(.dina(n33082), .dinb(n32864), .dout(n33083));
  jand g15821(.dina(n33083), .dinb(n33081), .dout(n33084));
  jand g15822(.dina(n33084), .dinb(n369), .dout(n33085));
  jor  g15823(.dina(n32862), .dinb(n32458), .dout(n33086));
  jxor g15824(.dina(n32728), .dinb(n32727), .dout(n33087));
  jor  g15825(.dina(n33087), .dinb(n32864), .dout(n33088));
  jand g15826(.dina(n33088), .dinb(n33086), .dout(n33089));
  jand g15827(.dina(n33089), .dinb(n368), .dout(n33090));
  jor  g15828(.dina(n32862), .dinb(n32463), .dout(n33091));
  jxor g15829(.dina(n32725), .dinb(n32724), .dout(n33092));
  jor  g15830(.dina(n33092), .dinb(n32864), .dout(n33093));
  jand g15831(.dina(n33093), .dinb(n33091), .dout(n33094));
  jand g15832(.dina(n33094), .dinb(n367), .dout(n33095));
  jor  g15833(.dina(n32862), .dinb(n32468), .dout(n33096));
  jxor g15834(.dina(n32722), .dinb(n32721), .dout(n33097));
  jor  g15835(.dina(n33097), .dinb(n32864), .dout(n33098));
  jand g15836(.dina(n33098), .dinb(n33096), .dout(n33099));
  jand g15837(.dina(n33099), .dinb(n265), .dout(n33100));
  jor  g15838(.dina(n32862), .dinb(n32473), .dout(n33101));
  jxor g15839(.dina(n32719), .dinb(n32718), .dout(n33102));
  jor  g15840(.dina(n33102), .dinb(n32864), .dout(n33103));
  jand g15841(.dina(n33103), .dinb(n33101), .dout(n33104));
  jand g15842(.dina(n33104), .dinb(n378), .dout(n33105));
  jor  g15843(.dina(n32862), .dinb(n32479), .dout(n33106));
  jxor g15844(.dina(n32716), .dinb(n32715), .dout(n33107));
  jor  g15845(.dina(n33107), .dinb(n32864), .dout(n33108));
  jand g15846(.dina(n33108), .dinb(n33106), .dout(n33109));
  jand g15847(.dina(n33109), .dinb(n377), .dout(n33110));
  jor  g15848(.dina(n32862), .dinb(n32484), .dout(n33111));
  jxor g15849(.dina(n32713), .dinb(n32712), .dout(n33112));
  jor  g15850(.dina(n33112), .dinb(n32864), .dout(n33113));
  jand g15851(.dina(n33113), .dinb(n33111), .dout(n33114));
  jand g15852(.dina(n33114), .dinb(n376), .dout(n33115));
  jor  g15853(.dina(n32862), .dinb(n32491), .dout(n33116));
  jxor g15854(.dina(n32710), .dinb(n32709), .dout(n33117));
  jor  g15855(.dina(n33117), .dinb(n32864), .dout(n33118));
  jand g15856(.dina(n33118), .dinb(n33116), .dout(n33119));
  jand g15857(.dina(n33119), .dinb(n264), .dout(n33120));
  jxor g15858(.dina(n32707), .dinb(n12438), .dout(n33121));
  jand g15859(.dina(n33121), .dinb(n32862), .dout(n33122));
  jnot g15860(.din(n33122), .dout(n33123));
  jor  g15861(.dina(n32862), .dinb(n32706), .dout(n33124));
  jand g15862(.dina(n33124), .dinb(n33123), .dout(n33125));
  jnot g15863(.din(n33125), .dout(n33126));
  jand g15864(.dina(n33126), .dinb(n386), .dout(n33127));
  jand g15865(.dina(n32862), .dinb(b0 ), .dout(n33128));
  jxor g15866(.dina(n33128), .dinb(a11 ), .dout(n33129));
  jand g15867(.dina(n33129), .dinb(n259), .dout(n33130));
  jxor g15868(.dina(n33128), .dinb(n12436), .dout(n33131));
  jxor g15869(.dina(n33131), .dinb(b1 ), .dout(n33132));
  jand g15870(.dina(n33132), .dinb(n12865), .dout(n33133));
  jor  g15871(.dina(n33133), .dinb(n33130), .dout(n33134));
  jxor g15872(.dina(n33125), .dinb(b2 ), .dout(n33135));
  jand g15873(.dina(n33135), .dinb(n33134), .dout(n33136));
  jor  g15874(.dina(n33136), .dinb(n33127), .dout(n33137));
  jxor g15875(.dina(n33119), .dinb(n264), .dout(n33138));
  jand g15876(.dina(n33138), .dinb(n33137), .dout(n33139));
  jor  g15877(.dina(n33139), .dinb(n33120), .dout(n33140));
  jxor g15878(.dina(n33114), .dinb(n376), .dout(n33141));
  jand g15879(.dina(n33141), .dinb(n33140), .dout(n33142));
  jor  g15880(.dina(n33142), .dinb(n33115), .dout(n33143));
  jxor g15881(.dina(n33109), .dinb(n377), .dout(n33144));
  jand g15882(.dina(n33144), .dinb(n33143), .dout(n33145));
  jor  g15883(.dina(n33145), .dinb(n33110), .dout(n33146));
  jxor g15884(.dina(n33104), .dinb(n378), .dout(n33147));
  jand g15885(.dina(n33147), .dinb(n33146), .dout(n33148));
  jor  g15886(.dina(n33148), .dinb(n33105), .dout(n33149));
  jxor g15887(.dina(n33099), .dinb(n265), .dout(n33150));
  jand g15888(.dina(n33150), .dinb(n33149), .dout(n33151));
  jor  g15889(.dina(n33151), .dinb(n33100), .dout(n33152));
  jxor g15890(.dina(n33094), .dinb(n367), .dout(n33153));
  jand g15891(.dina(n33153), .dinb(n33152), .dout(n33154));
  jor  g15892(.dina(n33154), .dinb(n33095), .dout(n33155));
  jxor g15893(.dina(n33089), .dinb(n368), .dout(n33156));
  jand g15894(.dina(n33156), .dinb(n33155), .dout(n33157));
  jor  g15895(.dina(n33157), .dinb(n33090), .dout(n33158));
  jxor g15896(.dina(n33084), .dinb(n369), .dout(n33159));
  jand g15897(.dina(n33159), .dinb(n33158), .dout(n33160));
  jor  g15898(.dina(n33160), .dinb(n33085), .dout(n33161));
  jxor g15899(.dina(n33079), .dinb(n359), .dout(n33162));
  jand g15900(.dina(n33162), .dinb(n33161), .dout(n33163));
  jor  g15901(.dina(n33163), .dinb(n33080), .dout(n33164));
  jxor g15902(.dina(n33074), .dinb(n363), .dout(n33165));
  jand g15903(.dina(n33165), .dinb(n33164), .dout(n33166));
  jor  g15904(.dina(n33166), .dinb(n33075), .dout(n33167));
  jxor g15905(.dina(n33069), .dinb(n360), .dout(n33168));
  jand g15906(.dina(n33168), .dinb(n33167), .dout(n33169));
  jor  g15907(.dina(n33169), .dinb(n33070), .dout(n33170));
  jxor g15908(.dina(n33064), .dinb(n361), .dout(n33171));
  jand g15909(.dina(n33171), .dinb(n33170), .dout(n33172));
  jor  g15910(.dina(n33172), .dinb(n33065), .dout(n33173));
  jxor g15911(.dina(n33059), .dinb(n364), .dout(n33174));
  jand g15912(.dina(n33174), .dinb(n33173), .dout(n33175));
  jor  g15913(.dina(n33175), .dinb(n33060), .dout(n33176));
  jxor g15914(.dina(n33054), .dinb(n355), .dout(n33177));
  jand g15915(.dina(n33177), .dinb(n33176), .dout(n33178));
  jor  g15916(.dina(n33178), .dinb(n33055), .dout(n33179));
  jxor g15917(.dina(n33049), .dinb(n356), .dout(n33180));
  jand g15918(.dina(n33180), .dinb(n33179), .dout(n33181));
  jor  g15919(.dina(n33181), .dinb(n33050), .dout(n33182));
  jxor g15920(.dina(n33044), .dinb(n266), .dout(n33183));
  jand g15921(.dina(n33183), .dinb(n33182), .dout(n33184));
  jor  g15922(.dina(n33184), .dinb(n33045), .dout(n33185));
  jxor g15923(.dina(n33039), .dinb(n267), .dout(n33186));
  jand g15924(.dina(n33186), .dinb(n33185), .dout(n33187));
  jor  g15925(.dina(n33187), .dinb(n33040), .dout(n33188));
  jxor g15926(.dina(n33034), .dinb(n347), .dout(n33189));
  jand g15927(.dina(n33189), .dinb(n33188), .dout(n33190));
  jor  g15928(.dina(n33190), .dinb(n33035), .dout(n33191));
  jxor g15929(.dina(n33029), .dinb(n348), .dout(n33192));
  jand g15930(.dina(n33192), .dinb(n33191), .dout(n33193));
  jor  g15931(.dina(n33193), .dinb(n33030), .dout(n33194));
  jxor g15932(.dina(n33024), .dinb(n349), .dout(n33195));
  jand g15933(.dina(n33195), .dinb(n33194), .dout(n33196));
  jor  g15934(.dina(n33196), .dinb(n33025), .dout(n33197));
  jxor g15935(.dina(n33019), .dinb(n268), .dout(n33198));
  jand g15936(.dina(n33198), .dinb(n33197), .dout(n33199));
  jor  g15937(.dina(n33199), .dinb(n33020), .dout(n33200));
  jxor g15938(.dina(n33014), .dinb(n274), .dout(n33201));
  jand g15939(.dina(n33201), .dinb(n33200), .dout(n33202));
  jor  g15940(.dina(n33202), .dinb(n33015), .dout(n33203));
  jxor g15941(.dina(n33009), .dinb(n269), .dout(n33204));
  jand g15942(.dina(n33204), .dinb(n33203), .dout(n33205));
  jor  g15943(.dina(n33205), .dinb(n33010), .dout(n33206));
  jxor g15944(.dina(n33004), .dinb(n270), .dout(n33207));
  jand g15945(.dina(n33207), .dinb(n33206), .dout(n33208));
  jor  g15946(.dina(n33208), .dinb(n33005), .dout(n33209));
  jxor g15947(.dina(n32999), .dinb(n271), .dout(n33210));
  jand g15948(.dina(n33210), .dinb(n33209), .dout(n33211));
  jor  g15949(.dina(n33211), .dinb(n33000), .dout(n33212));
  jxor g15950(.dina(n32994), .dinb(n338), .dout(n33213));
  jand g15951(.dina(n33213), .dinb(n33212), .dout(n33214));
  jor  g15952(.dina(n33214), .dinb(n32995), .dout(n33215));
  jxor g15953(.dina(n32989), .dinb(n339), .dout(n33216));
  jand g15954(.dina(n33216), .dinb(n33215), .dout(n33217));
  jor  g15955(.dina(n33217), .dinb(n32990), .dout(n33218));
  jxor g15956(.dina(n32984), .dinb(n340), .dout(n33219));
  jand g15957(.dina(n33219), .dinb(n33218), .dout(n33220));
  jor  g15958(.dina(n33220), .dinb(n32985), .dout(n33221));
  jxor g15959(.dina(n32979), .dinb(n275), .dout(n33222));
  jand g15960(.dina(n33222), .dinb(n33221), .dout(n33223));
  jor  g15961(.dina(n33223), .dinb(n32980), .dout(n33224));
  jxor g15962(.dina(n32974), .dinb(n331), .dout(n33225));
  jand g15963(.dina(n33225), .dinb(n33224), .dout(n33226));
  jor  g15964(.dina(n33226), .dinb(n32975), .dout(n33227));
  jxor g15965(.dina(n32969), .dinb(n332), .dout(n33228));
  jand g15966(.dina(n33228), .dinb(n33227), .dout(n33229));
  jor  g15967(.dina(n33229), .dinb(n32970), .dout(n33230));
  jxor g15968(.dina(n32964), .dinb(n333), .dout(n33231));
  jand g15969(.dina(n33231), .dinb(n33230), .dout(n33232));
  jor  g15970(.dina(n33232), .dinb(n32965), .dout(n33233));
  jxor g15971(.dina(n32959), .dinb(n276), .dout(n33234));
  jand g15972(.dina(n33234), .dinb(n33233), .dout(n33235));
  jor  g15973(.dina(n33235), .dinb(n32960), .dout(n33236));
  jxor g15974(.dina(n32954), .dinb(n324), .dout(n33237));
  jand g15975(.dina(n33237), .dinb(n33236), .dout(n33238));
  jor  g15976(.dina(n33238), .dinb(n32955), .dout(n33239));
  jxor g15977(.dina(n32949), .dinb(n325), .dout(n33240));
  jand g15978(.dina(n33240), .dinb(n33239), .dout(n33241));
  jor  g15979(.dina(n33241), .dinb(n32950), .dout(n33242));
  jxor g15980(.dina(n32944), .dinb(n326), .dout(n33243));
  jand g15981(.dina(n33243), .dinb(n33242), .dout(n33244));
  jor  g15982(.dina(n33244), .dinb(n32945), .dout(n33245));
  jxor g15983(.dina(n32939), .dinb(n277), .dout(n33246));
  jand g15984(.dina(n33246), .dinb(n33245), .dout(n33247));
  jor  g15985(.dina(n33247), .dinb(n32940), .dout(n33248));
  jxor g15986(.dina(n32934), .dinb(n278), .dout(n33249));
  jand g15987(.dina(n33249), .dinb(n33248), .dout(n33250));
  jor  g15988(.dina(n33250), .dinb(n32935), .dout(n33251));
  jxor g15989(.dina(n32929), .dinb(n279), .dout(n33252));
  jand g15990(.dina(n33252), .dinb(n33251), .dout(n33253));
  jor  g15991(.dina(n33253), .dinb(n32930), .dout(n33254));
  jxor g15992(.dina(n32924), .dinb(n280), .dout(n33255));
  jand g15993(.dina(n33255), .dinb(n33254), .dout(n33256));
  jor  g15994(.dina(n33256), .dinb(n32925), .dout(n33257));
  jxor g15995(.dina(n32919), .dinb(n283), .dout(n33258));
  jand g15996(.dina(n33258), .dinb(n33257), .dout(n33259));
  jor  g15997(.dina(n33259), .dinb(n32920), .dout(n33260));
  jxor g15998(.dina(n32914), .dinb(n315), .dout(n33261));
  jand g15999(.dina(n33261), .dinb(n33260), .dout(n33262));
  jor  g16000(.dina(n33262), .dinb(n32915), .dout(n33263));
  jxor g16001(.dina(n32909), .dinb(n316), .dout(n33264));
  jand g16002(.dina(n33264), .dinb(n33263), .dout(n33265));
  jor  g16003(.dina(n33265), .dinb(n32910), .dout(n33266));
  jxor g16004(.dina(n32904), .dinb(n317), .dout(n33267));
  jand g16005(.dina(n33267), .dinb(n33266), .dout(n33268));
  jor  g16006(.dina(n33268), .dinb(n32905), .dout(n33269));
  jxor g16007(.dina(n32899), .dinb(n284), .dout(n33270));
  jand g16008(.dina(n33270), .dinb(n33269), .dout(n33271));
  jor  g16009(.dina(n33271), .dinb(n32900), .dout(n33272));
  jxor g16010(.dina(n32894), .dinb(n285), .dout(n33273));
  jand g16011(.dina(n33273), .dinb(n33272), .dout(n33274));
  jor  g16012(.dina(n33274), .dinb(n32895), .dout(n33275));
  jxor g16013(.dina(n32889), .dinb(n286), .dout(n33276));
  jand g16014(.dina(n33276), .dinb(n33275), .dout(n33277));
  jor  g16015(.dina(n33277), .dinb(n32890), .dout(n33278));
  jxor g16016(.dina(n32884), .dinb(n287), .dout(n33279));
  jand g16017(.dina(n33279), .dinb(n33278), .dout(n33280));
  jor  g16018(.dina(n33280), .dinb(n32885), .dout(n33281));
  jxor g16019(.dina(n32879), .dinb(n288), .dout(n33282));
  jand g16020(.dina(n33282), .dinb(n33281), .dout(n33283));
  jor  g16021(.dina(n33283), .dinb(n32880), .dout(n33284));
  jxor g16022(.dina(n32867), .dinb(n289), .dout(n33285));
  jand g16023(.dina(n33285), .dinb(n33284), .dout(n33286));
  jor  g16024(.dina(n33286), .dinb(n32875), .dout(n33287));
  jand g16025(.dina(n33287), .dinb(n32874), .dout(n33288));
  jor  g16026(.dina(n33288), .dinb(n32871), .dout(n33289));
  jand g16027(.dina(n33289), .dinb(n307), .dout(n33290));
  jor  g16028(.dina(n33290), .dinb(n32867), .dout(n33291));
  jnot g16029(.din(n33290), .dout(n33292));
  jxor g16030(.dina(n33285), .dinb(n33284), .dout(n33293));
  jor  g16031(.dina(n33293), .dinb(n33292), .dout(n33294));
  jand g16032(.dina(n33294), .dinb(n33291), .dout(n33295));
  jand g16033(.dina(n33292), .dinb(n32870), .dout(n33296));
  jand g16034(.dina(n33287), .dinb(n32871), .dout(n33297));
  jor  g16035(.dina(n33297), .dinb(n33296), .dout(n33298));
  jand g16036(.dina(n33298), .dinb(n291), .dout(n33299));
  jnot g16037(.din(n33298), .dout(n33300));
  jand g16038(.dina(n33300), .dinb(b54 ), .dout(n33301));
  jnot g16039(.din(n33301), .dout(n33302));
  jand g16040(.dina(n33295), .dinb(n290), .dout(n33303));
  jor  g16041(.dina(n33290), .dinb(n32879), .dout(n33304));
  jxor g16042(.dina(n33282), .dinb(n33281), .dout(n33305));
  jor  g16043(.dina(n33305), .dinb(n33292), .dout(n33306));
  jand g16044(.dina(n33306), .dinb(n33304), .dout(n33307));
  jand g16045(.dina(n33307), .dinb(n289), .dout(n33308));
  jor  g16046(.dina(n33290), .dinb(n32884), .dout(n33309));
  jxor g16047(.dina(n33279), .dinb(n33278), .dout(n33310));
  jor  g16048(.dina(n33310), .dinb(n33292), .dout(n33311));
  jand g16049(.dina(n33311), .dinb(n33309), .dout(n33312));
  jand g16050(.dina(n33312), .dinb(n288), .dout(n33313));
  jor  g16051(.dina(n33290), .dinb(n32889), .dout(n33314));
  jxor g16052(.dina(n33276), .dinb(n33275), .dout(n33315));
  jor  g16053(.dina(n33315), .dinb(n33292), .dout(n33316));
  jand g16054(.dina(n33316), .dinb(n33314), .dout(n33317));
  jand g16055(.dina(n33317), .dinb(n287), .dout(n33318));
  jor  g16056(.dina(n33290), .dinb(n32894), .dout(n33319));
  jxor g16057(.dina(n33273), .dinb(n33272), .dout(n33320));
  jor  g16058(.dina(n33320), .dinb(n33292), .dout(n33321));
  jand g16059(.dina(n33321), .dinb(n33319), .dout(n33322));
  jand g16060(.dina(n33322), .dinb(n286), .dout(n33323));
  jor  g16061(.dina(n33290), .dinb(n32899), .dout(n33324));
  jxor g16062(.dina(n33270), .dinb(n33269), .dout(n33325));
  jor  g16063(.dina(n33325), .dinb(n33292), .dout(n33326));
  jand g16064(.dina(n33326), .dinb(n33324), .dout(n33327));
  jand g16065(.dina(n33327), .dinb(n285), .dout(n33328));
  jor  g16066(.dina(n33290), .dinb(n32904), .dout(n33329));
  jxor g16067(.dina(n33267), .dinb(n33266), .dout(n33330));
  jor  g16068(.dina(n33330), .dinb(n33292), .dout(n33331));
  jand g16069(.dina(n33331), .dinb(n33329), .dout(n33332));
  jand g16070(.dina(n33332), .dinb(n284), .dout(n33333));
  jor  g16071(.dina(n33290), .dinb(n32909), .dout(n33334));
  jxor g16072(.dina(n33264), .dinb(n33263), .dout(n33335));
  jor  g16073(.dina(n33335), .dinb(n33292), .dout(n33336));
  jand g16074(.dina(n33336), .dinb(n33334), .dout(n33337));
  jand g16075(.dina(n33337), .dinb(n317), .dout(n33338));
  jor  g16076(.dina(n33290), .dinb(n32914), .dout(n33339));
  jxor g16077(.dina(n33261), .dinb(n33260), .dout(n33340));
  jor  g16078(.dina(n33340), .dinb(n33292), .dout(n33341));
  jand g16079(.dina(n33341), .dinb(n33339), .dout(n33342));
  jand g16080(.dina(n33342), .dinb(n316), .dout(n33343));
  jor  g16081(.dina(n33290), .dinb(n32919), .dout(n33344));
  jxor g16082(.dina(n33258), .dinb(n33257), .dout(n33345));
  jor  g16083(.dina(n33345), .dinb(n33292), .dout(n33346));
  jand g16084(.dina(n33346), .dinb(n33344), .dout(n33347));
  jand g16085(.dina(n33347), .dinb(n315), .dout(n33348));
  jor  g16086(.dina(n33290), .dinb(n32924), .dout(n33349));
  jxor g16087(.dina(n33255), .dinb(n33254), .dout(n33350));
  jor  g16088(.dina(n33350), .dinb(n33292), .dout(n33351));
  jand g16089(.dina(n33351), .dinb(n33349), .dout(n33352));
  jand g16090(.dina(n33352), .dinb(n283), .dout(n33353));
  jor  g16091(.dina(n33290), .dinb(n32929), .dout(n33354));
  jxor g16092(.dina(n33252), .dinb(n33251), .dout(n33355));
  jor  g16093(.dina(n33355), .dinb(n33292), .dout(n33356));
  jand g16094(.dina(n33356), .dinb(n33354), .dout(n33357));
  jand g16095(.dina(n33357), .dinb(n280), .dout(n33358));
  jor  g16096(.dina(n33290), .dinb(n32934), .dout(n33359));
  jxor g16097(.dina(n33249), .dinb(n33248), .dout(n33360));
  jor  g16098(.dina(n33360), .dinb(n33292), .dout(n33361));
  jand g16099(.dina(n33361), .dinb(n33359), .dout(n33362));
  jand g16100(.dina(n33362), .dinb(n279), .dout(n33363));
  jor  g16101(.dina(n33290), .dinb(n32939), .dout(n33364));
  jxor g16102(.dina(n33246), .dinb(n33245), .dout(n33365));
  jor  g16103(.dina(n33365), .dinb(n33292), .dout(n33366));
  jand g16104(.dina(n33366), .dinb(n33364), .dout(n33367));
  jand g16105(.dina(n33367), .dinb(n278), .dout(n33368));
  jor  g16106(.dina(n33290), .dinb(n32944), .dout(n33369));
  jxor g16107(.dina(n33243), .dinb(n33242), .dout(n33370));
  jor  g16108(.dina(n33370), .dinb(n33292), .dout(n33371));
  jand g16109(.dina(n33371), .dinb(n33369), .dout(n33372));
  jand g16110(.dina(n33372), .dinb(n277), .dout(n33373));
  jor  g16111(.dina(n33290), .dinb(n32949), .dout(n33374));
  jxor g16112(.dina(n33240), .dinb(n33239), .dout(n33375));
  jor  g16113(.dina(n33375), .dinb(n33292), .dout(n33376));
  jand g16114(.dina(n33376), .dinb(n33374), .dout(n33377));
  jand g16115(.dina(n33377), .dinb(n326), .dout(n33378));
  jor  g16116(.dina(n33290), .dinb(n32954), .dout(n33379));
  jxor g16117(.dina(n33237), .dinb(n33236), .dout(n33380));
  jor  g16118(.dina(n33380), .dinb(n33292), .dout(n33381));
  jand g16119(.dina(n33381), .dinb(n33379), .dout(n33382));
  jand g16120(.dina(n33382), .dinb(n325), .dout(n33383));
  jor  g16121(.dina(n33290), .dinb(n32959), .dout(n33384));
  jxor g16122(.dina(n33234), .dinb(n33233), .dout(n33385));
  jor  g16123(.dina(n33385), .dinb(n33292), .dout(n33386));
  jand g16124(.dina(n33386), .dinb(n33384), .dout(n33387));
  jand g16125(.dina(n33387), .dinb(n324), .dout(n33388));
  jor  g16126(.dina(n33290), .dinb(n32964), .dout(n33389));
  jxor g16127(.dina(n33231), .dinb(n33230), .dout(n33390));
  jor  g16128(.dina(n33390), .dinb(n33292), .dout(n33391));
  jand g16129(.dina(n33391), .dinb(n33389), .dout(n33392));
  jand g16130(.dina(n33392), .dinb(n276), .dout(n33393));
  jor  g16131(.dina(n33290), .dinb(n32969), .dout(n33394));
  jxor g16132(.dina(n33228), .dinb(n33227), .dout(n33395));
  jor  g16133(.dina(n33395), .dinb(n33292), .dout(n33396));
  jand g16134(.dina(n33396), .dinb(n33394), .dout(n33397));
  jand g16135(.dina(n33397), .dinb(n333), .dout(n33398));
  jor  g16136(.dina(n33290), .dinb(n32974), .dout(n33399));
  jxor g16137(.dina(n33225), .dinb(n33224), .dout(n33400));
  jor  g16138(.dina(n33400), .dinb(n33292), .dout(n33401));
  jand g16139(.dina(n33401), .dinb(n33399), .dout(n33402));
  jand g16140(.dina(n33402), .dinb(n332), .dout(n33403));
  jor  g16141(.dina(n33290), .dinb(n32979), .dout(n33404));
  jxor g16142(.dina(n33222), .dinb(n33221), .dout(n33405));
  jor  g16143(.dina(n33405), .dinb(n33292), .dout(n33406));
  jand g16144(.dina(n33406), .dinb(n33404), .dout(n33407));
  jand g16145(.dina(n33407), .dinb(n331), .dout(n33408));
  jor  g16146(.dina(n33290), .dinb(n32984), .dout(n33409));
  jxor g16147(.dina(n33219), .dinb(n33218), .dout(n33410));
  jor  g16148(.dina(n33410), .dinb(n33292), .dout(n33411));
  jand g16149(.dina(n33411), .dinb(n33409), .dout(n33412));
  jand g16150(.dina(n33412), .dinb(n275), .dout(n33413));
  jor  g16151(.dina(n33290), .dinb(n32989), .dout(n33414));
  jxor g16152(.dina(n33216), .dinb(n33215), .dout(n33415));
  jor  g16153(.dina(n33415), .dinb(n33292), .dout(n33416));
  jand g16154(.dina(n33416), .dinb(n33414), .dout(n33417));
  jand g16155(.dina(n33417), .dinb(n340), .dout(n33418));
  jor  g16156(.dina(n33290), .dinb(n32994), .dout(n33419));
  jxor g16157(.dina(n33213), .dinb(n33212), .dout(n33420));
  jor  g16158(.dina(n33420), .dinb(n33292), .dout(n33421));
  jand g16159(.dina(n33421), .dinb(n33419), .dout(n33422));
  jand g16160(.dina(n33422), .dinb(n339), .dout(n33423));
  jor  g16161(.dina(n33290), .dinb(n32999), .dout(n33424));
  jxor g16162(.dina(n33210), .dinb(n33209), .dout(n33425));
  jor  g16163(.dina(n33425), .dinb(n33292), .dout(n33426));
  jand g16164(.dina(n33426), .dinb(n33424), .dout(n33427));
  jand g16165(.dina(n33427), .dinb(n338), .dout(n33428));
  jor  g16166(.dina(n33290), .dinb(n33004), .dout(n33429));
  jxor g16167(.dina(n33207), .dinb(n33206), .dout(n33430));
  jor  g16168(.dina(n33430), .dinb(n33292), .dout(n33431));
  jand g16169(.dina(n33431), .dinb(n33429), .dout(n33432));
  jand g16170(.dina(n33432), .dinb(n271), .dout(n33433));
  jor  g16171(.dina(n33290), .dinb(n33009), .dout(n33434));
  jxor g16172(.dina(n33204), .dinb(n33203), .dout(n33435));
  jor  g16173(.dina(n33435), .dinb(n33292), .dout(n33436));
  jand g16174(.dina(n33436), .dinb(n33434), .dout(n33437));
  jand g16175(.dina(n33437), .dinb(n270), .dout(n33438));
  jor  g16176(.dina(n33290), .dinb(n33014), .dout(n33439));
  jxor g16177(.dina(n33201), .dinb(n33200), .dout(n33440));
  jor  g16178(.dina(n33440), .dinb(n33292), .dout(n33441));
  jand g16179(.dina(n33441), .dinb(n33439), .dout(n33442));
  jand g16180(.dina(n33442), .dinb(n269), .dout(n33443));
  jor  g16181(.dina(n33290), .dinb(n33019), .dout(n33444));
  jxor g16182(.dina(n33198), .dinb(n33197), .dout(n33445));
  jor  g16183(.dina(n33445), .dinb(n33292), .dout(n33446));
  jand g16184(.dina(n33446), .dinb(n33444), .dout(n33447));
  jand g16185(.dina(n33447), .dinb(n274), .dout(n33448));
  jor  g16186(.dina(n33290), .dinb(n33024), .dout(n33449));
  jxor g16187(.dina(n33195), .dinb(n33194), .dout(n33450));
  jor  g16188(.dina(n33450), .dinb(n33292), .dout(n33451));
  jand g16189(.dina(n33451), .dinb(n33449), .dout(n33452));
  jand g16190(.dina(n33452), .dinb(n268), .dout(n33453));
  jor  g16191(.dina(n33290), .dinb(n33029), .dout(n33454));
  jxor g16192(.dina(n33192), .dinb(n33191), .dout(n33455));
  jor  g16193(.dina(n33455), .dinb(n33292), .dout(n33456));
  jand g16194(.dina(n33456), .dinb(n33454), .dout(n33457));
  jand g16195(.dina(n33457), .dinb(n349), .dout(n33458));
  jor  g16196(.dina(n33290), .dinb(n33034), .dout(n33459));
  jxor g16197(.dina(n33189), .dinb(n33188), .dout(n33460));
  jor  g16198(.dina(n33460), .dinb(n33292), .dout(n33461));
  jand g16199(.dina(n33461), .dinb(n33459), .dout(n33462));
  jand g16200(.dina(n33462), .dinb(n348), .dout(n33463));
  jor  g16201(.dina(n33290), .dinb(n33039), .dout(n33464));
  jxor g16202(.dina(n33186), .dinb(n33185), .dout(n33465));
  jor  g16203(.dina(n33465), .dinb(n33292), .dout(n33466));
  jand g16204(.dina(n33466), .dinb(n33464), .dout(n33467));
  jand g16205(.dina(n33467), .dinb(n347), .dout(n33468));
  jor  g16206(.dina(n33290), .dinb(n33044), .dout(n33469));
  jxor g16207(.dina(n33183), .dinb(n33182), .dout(n33470));
  jor  g16208(.dina(n33470), .dinb(n33292), .dout(n33471));
  jand g16209(.dina(n33471), .dinb(n33469), .dout(n33472));
  jand g16210(.dina(n33472), .dinb(n267), .dout(n33473));
  jor  g16211(.dina(n33290), .dinb(n33049), .dout(n33474));
  jxor g16212(.dina(n33180), .dinb(n33179), .dout(n33475));
  jor  g16213(.dina(n33475), .dinb(n33292), .dout(n33476));
  jand g16214(.dina(n33476), .dinb(n33474), .dout(n33477));
  jand g16215(.dina(n33477), .dinb(n266), .dout(n33478));
  jor  g16216(.dina(n33290), .dinb(n33054), .dout(n33479));
  jxor g16217(.dina(n33177), .dinb(n33176), .dout(n33480));
  jor  g16218(.dina(n33480), .dinb(n33292), .dout(n33481));
  jand g16219(.dina(n33481), .dinb(n33479), .dout(n33482));
  jand g16220(.dina(n33482), .dinb(n356), .dout(n33483));
  jor  g16221(.dina(n33290), .dinb(n33059), .dout(n33484));
  jxor g16222(.dina(n33174), .dinb(n33173), .dout(n33485));
  jor  g16223(.dina(n33485), .dinb(n33292), .dout(n33486));
  jand g16224(.dina(n33486), .dinb(n33484), .dout(n33487));
  jand g16225(.dina(n33487), .dinb(n355), .dout(n33488));
  jor  g16226(.dina(n33290), .dinb(n33064), .dout(n33489));
  jxor g16227(.dina(n33171), .dinb(n33170), .dout(n33490));
  jor  g16228(.dina(n33490), .dinb(n33292), .dout(n33491));
  jand g16229(.dina(n33491), .dinb(n33489), .dout(n33492));
  jand g16230(.dina(n33492), .dinb(n364), .dout(n33493));
  jor  g16231(.dina(n33290), .dinb(n33069), .dout(n33494));
  jxor g16232(.dina(n33168), .dinb(n33167), .dout(n33495));
  jor  g16233(.dina(n33495), .dinb(n33292), .dout(n33496));
  jand g16234(.dina(n33496), .dinb(n33494), .dout(n33497));
  jand g16235(.dina(n33497), .dinb(n361), .dout(n33498));
  jor  g16236(.dina(n33290), .dinb(n33074), .dout(n33499));
  jxor g16237(.dina(n33165), .dinb(n33164), .dout(n33500));
  jor  g16238(.dina(n33500), .dinb(n33292), .dout(n33501));
  jand g16239(.dina(n33501), .dinb(n33499), .dout(n33502));
  jand g16240(.dina(n33502), .dinb(n360), .dout(n33503));
  jor  g16241(.dina(n33290), .dinb(n33079), .dout(n33504));
  jxor g16242(.dina(n33162), .dinb(n33161), .dout(n33505));
  jor  g16243(.dina(n33505), .dinb(n33292), .dout(n33506));
  jand g16244(.dina(n33506), .dinb(n33504), .dout(n33507));
  jand g16245(.dina(n33507), .dinb(n363), .dout(n33508));
  jor  g16246(.dina(n33290), .dinb(n33084), .dout(n33509));
  jxor g16247(.dina(n33159), .dinb(n33158), .dout(n33510));
  jor  g16248(.dina(n33510), .dinb(n33292), .dout(n33511));
  jand g16249(.dina(n33511), .dinb(n33509), .dout(n33512));
  jand g16250(.dina(n33512), .dinb(n359), .dout(n33513));
  jor  g16251(.dina(n33290), .dinb(n33089), .dout(n33514));
  jxor g16252(.dina(n33156), .dinb(n33155), .dout(n33515));
  jor  g16253(.dina(n33515), .dinb(n33292), .dout(n33516));
  jand g16254(.dina(n33516), .dinb(n33514), .dout(n33517));
  jand g16255(.dina(n33517), .dinb(n369), .dout(n33518));
  jor  g16256(.dina(n33290), .dinb(n33094), .dout(n33519));
  jxor g16257(.dina(n33153), .dinb(n33152), .dout(n33520));
  jor  g16258(.dina(n33520), .dinb(n33292), .dout(n33521));
  jand g16259(.dina(n33521), .dinb(n33519), .dout(n33522));
  jand g16260(.dina(n33522), .dinb(n368), .dout(n33523));
  jor  g16261(.dina(n33290), .dinb(n33099), .dout(n33524));
  jxor g16262(.dina(n33150), .dinb(n33149), .dout(n33525));
  jor  g16263(.dina(n33525), .dinb(n33292), .dout(n33526));
  jand g16264(.dina(n33526), .dinb(n33524), .dout(n33527));
  jand g16265(.dina(n33527), .dinb(n367), .dout(n33528));
  jor  g16266(.dina(n33290), .dinb(n33104), .dout(n33529));
  jxor g16267(.dina(n33147), .dinb(n33146), .dout(n33530));
  jor  g16268(.dina(n33530), .dinb(n33292), .dout(n33531));
  jand g16269(.dina(n33531), .dinb(n33529), .dout(n33532));
  jand g16270(.dina(n33532), .dinb(n265), .dout(n33533));
  jor  g16271(.dina(n33290), .dinb(n33109), .dout(n33534));
  jxor g16272(.dina(n33144), .dinb(n33143), .dout(n33535));
  jor  g16273(.dina(n33535), .dinb(n33292), .dout(n33536));
  jand g16274(.dina(n33536), .dinb(n33534), .dout(n33537));
  jand g16275(.dina(n33537), .dinb(n378), .dout(n33538));
  jor  g16276(.dina(n33290), .dinb(n33114), .dout(n33539));
  jxor g16277(.dina(n33141), .dinb(n33140), .dout(n33540));
  jor  g16278(.dina(n33540), .dinb(n33292), .dout(n33541));
  jand g16279(.dina(n33541), .dinb(n33539), .dout(n33542));
  jand g16280(.dina(n33542), .dinb(n377), .dout(n33543));
  jor  g16281(.dina(n33290), .dinb(n33119), .dout(n33544));
  jxor g16282(.dina(n33138), .dinb(n33137), .dout(n33545));
  jor  g16283(.dina(n33545), .dinb(n33292), .dout(n33546));
  jand g16284(.dina(n33546), .dinb(n33544), .dout(n33547));
  jand g16285(.dina(n33547), .dinb(n376), .dout(n33548));
  jor  g16286(.dina(n33290), .dinb(n33126), .dout(n33549));
  jxor g16287(.dina(n33135), .dinb(n33134), .dout(n33550));
  jor  g16288(.dina(n33550), .dinb(n33292), .dout(n33551));
  jand g16289(.dina(n33551), .dinb(n33549), .dout(n33552));
  jand g16290(.dina(n33552), .dinb(n264), .dout(n33553));
  jxor g16291(.dina(n33132), .dinb(n12865), .dout(n33554));
  jand g16292(.dina(n33554), .dinb(n33290), .dout(n33555));
  jnot g16293(.din(n33555), .dout(n33556));
  jor  g16294(.dina(n33290), .dinb(n33131), .dout(n33557));
  jand g16295(.dina(n33557), .dinb(n33556), .dout(n33558));
  jnot g16296(.din(n33558), .dout(n33559));
  jand g16297(.dina(n33559), .dinb(n386), .dout(n33560));
  jand g16298(.dina(n33290), .dinb(b0 ), .dout(n33561));
  jxor g16299(.dina(n33561), .dinb(a10 ), .dout(n33562));
  jand g16300(.dina(n33562), .dinb(n259), .dout(n33563));
  jxor g16301(.dina(n33561), .dinb(n12863), .dout(n33564));
  jxor g16302(.dina(n33564), .dinb(b1 ), .dout(n33565));
  jand g16303(.dina(n33565), .dinb(n13302), .dout(n33566));
  jor  g16304(.dina(n33566), .dinb(n33563), .dout(n33567));
  jxor g16305(.dina(n33558), .dinb(b2 ), .dout(n33568));
  jand g16306(.dina(n33568), .dinb(n33567), .dout(n33569));
  jor  g16307(.dina(n33569), .dinb(n33560), .dout(n33570));
  jxor g16308(.dina(n33552), .dinb(n264), .dout(n33571));
  jand g16309(.dina(n33571), .dinb(n33570), .dout(n33572));
  jor  g16310(.dina(n33572), .dinb(n33553), .dout(n33573));
  jxor g16311(.dina(n33547), .dinb(n376), .dout(n33574));
  jand g16312(.dina(n33574), .dinb(n33573), .dout(n33575));
  jor  g16313(.dina(n33575), .dinb(n33548), .dout(n33576));
  jxor g16314(.dina(n33542), .dinb(n377), .dout(n33577));
  jand g16315(.dina(n33577), .dinb(n33576), .dout(n33578));
  jor  g16316(.dina(n33578), .dinb(n33543), .dout(n33579));
  jxor g16317(.dina(n33537), .dinb(n378), .dout(n33580));
  jand g16318(.dina(n33580), .dinb(n33579), .dout(n33581));
  jor  g16319(.dina(n33581), .dinb(n33538), .dout(n33582));
  jxor g16320(.dina(n33532), .dinb(n265), .dout(n33583));
  jand g16321(.dina(n33583), .dinb(n33582), .dout(n33584));
  jor  g16322(.dina(n33584), .dinb(n33533), .dout(n33585));
  jxor g16323(.dina(n33527), .dinb(n367), .dout(n33586));
  jand g16324(.dina(n33586), .dinb(n33585), .dout(n33587));
  jor  g16325(.dina(n33587), .dinb(n33528), .dout(n33588));
  jxor g16326(.dina(n33522), .dinb(n368), .dout(n33589));
  jand g16327(.dina(n33589), .dinb(n33588), .dout(n33590));
  jor  g16328(.dina(n33590), .dinb(n33523), .dout(n33591));
  jxor g16329(.dina(n33517), .dinb(n369), .dout(n33592));
  jand g16330(.dina(n33592), .dinb(n33591), .dout(n33593));
  jor  g16331(.dina(n33593), .dinb(n33518), .dout(n33594));
  jxor g16332(.dina(n33512), .dinb(n359), .dout(n33595));
  jand g16333(.dina(n33595), .dinb(n33594), .dout(n33596));
  jor  g16334(.dina(n33596), .dinb(n33513), .dout(n33597));
  jxor g16335(.dina(n33507), .dinb(n363), .dout(n33598));
  jand g16336(.dina(n33598), .dinb(n33597), .dout(n33599));
  jor  g16337(.dina(n33599), .dinb(n33508), .dout(n33600));
  jxor g16338(.dina(n33502), .dinb(n360), .dout(n33601));
  jand g16339(.dina(n33601), .dinb(n33600), .dout(n33602));
  jor  g16340(.dina(n33602), .dinb(n33503), .dout(n33603));
  jxor g16341(.dina(n33497), .dinb(n361), .dout(n33604));
  jand g16342(.dina(n33604), .dinb(n33603), .dout(n33605));
  jor  g16343(.dina(n33605), .dinb(n33498), .dout(n33606));
  jxor g16344(.dina(n33492), .dinb(n364), .dout(n33607));
  jand g16345(.dina(n33607), .dinb(n33606), .dout(n33608));
  jor  g16346(.dina(n33608), .dinb(n33493), .dout(n33609));
  jxor g16347(.dina(n33487), .dinb(n355), .dout(n33610));
  jand g16348(.dina(n33610), .dinb(n33609), .dout(n33611));
  jor  g16349(.dina(n33611), .dinb(n33488), .dout(n33612));
  jxor g16350(.dina(n33482), .dinb(n356), .dout(n33613));
  jand g16351(.dina(n33613), .dinb(n33612), .dout(n33614));
  jor  g16352(.dina(n33614), .dinb(n33483), .dout(n33615));
  jxor g16353(.dina(n33477), .dinb(n266), .dout(n33616));
  jand g16354(.dina(n33616), .dinb(n33615), .dout(n33617));
  jor  g16355(.dina(n33617), .dinb(n33478), .dout(n33618));
  jxor g16356(.dina(n33472), .dinb(n267), .dout(n33619));
  jand g16357(.dina(n33619), .dinb(n33618), .dout(n33620));
  jor  g16358(.dina(n33620), .dinb(n33473), .dout(n33621));
  jxor g16359(.dina(n33467), .dinb(n347), .dout(n33622));
  jand g16360(.dina(n33622), .dinb(n33621), .dout(n33623));
  jor  g16361(.dina(n33623), .dinb(n33468), .dout(n33624));
  jxor g16362(.dina(n33462), .dinb(n348), .dout(n33625));
  jand g16363(.dina(n33625), .dinb(n33624), .dout(n33626));
  jor  g16364(.dina(n33626), .dinb(n33463), .dout(n33627));
  jxor g16365(.dina(n33457), .dinb(n349), .dout(n33628));
  jand g16366(.dina(n33628), .dinb(n33627), .dout(n33629));
  jor  g16367(.dina(n33629), .dinb(n33458), .dout(n33630));
  jxor g16368(.dina(n33452), .dinb(n268), .dout(n33631));
  jand g16369(.dina(n33631), .dinb(n33630), .dout(n33632));
  jor  g16370(.dina(n33632), .dinb(n33453), .dout(n33633));
  jxor g16371(.dina(n33447), .dinb(n274), .dout(n33634));
  jand g16372(.dina(n33634), .dinb(n33633), .dout(n33635));
  jor  g16373(.dina(n33635), .dinb(n33448), .dout(n33636));
  jxor g16374(.dina(n33442), .dinb(n269), .dout(n33637));
  jand g16375(.dina(n33637), .dinb(n33636), .dout(n33638));
  jor  g16376(.dina(n33638), .dinb(n33443), .dout(n33639));
  jxor g16377(.dina(n33437), .dinb(n270), .dout(n33640));
  jand g16378(.dina(n33640), .dinb(n33639), .dout(n33641));
  jor  g16379(.dina(n33641), .dinb(n33438), .dout(n33642));
  jxor g16380(.dina(n33432), .dinb(n271), .dout(n33643));
  jand g16381(.dina(n33643), .dinb(n33642), .dout(n33644));
  jor  g16382(.dina(n33644), .dinb(n33433), .dout(n33645));
  jxor g16383(.dina(n33427), .dinb(n338), .dout(n33646));
  jand g16384(.dina(n33646), .dinb(n33645), .dout(n33647));
  jor  g16385(.dina(n33647), .dinb(n33428), .dout(n33648));
  jxor g16386(.dina(n33422), .dinb(n339), .dout(n33649));
  jand g16387(.dina(n33649), .dinb(n33648), .dout(n33650));
  jor  g16388(.dina(n33650), .dinb(n33423), .dout(n33651));
  jxor g16389(.dina(n33417), .dinb(n340), .dout(n33652));
  jand g16390(.dina(n33652), .dinb(n33651), .dout(n33653));
  jor  g16391(.dina(n33653), .dinb(n33418), .dout(n33654));
  jxor g16392(.dina(n33412), .dinb(n275), .dout(n33655));
  jand g16393(.dina(n33655), .dinb(n33654), .dout(n33656));
  jor  g16394(.dina(n33656), .dinb(n33413), .dout(n33657));
  jxor g16395(.dina(n33407), .dinb(n331), .dout(n33658));
  jand g16396(.dina(n33658), .dinb(n33657), .dout(n33659));
  jor  g16397(.dina(n33659), .dinb(n33408), .dout(n33660));
  jxor g16398(.dina(n33402), .dinb(n332), .dout(n33661));
  jand g16399(.dina(n33661), .dinb(n33660), .dout(n33662));
  jor  g16400(.dina(n33662), .dinb(n33403), .dout(n33663));
  jxor g16401(.dina(n33397), .dinb(n333), .dout(n33664));
  jand g16402(.dina(n33664), .dinb(n33663), .dout(n33665));
  jor  g16403(.dina(n33665), .dinb(n33398), .dout(n33666));
  jxor g16404(.dina(n33392), .dinb(n276), .dout(n33667));
  jand g16405(.dina(n33667), .dinb(n33666), .dout(n33668));
  jor  g16406(.dina(n33668), .dinb(n33393), .dout(n33669));
  jxor g16407(.dina(n33387), .dinb(n324), .dout(n33670));
  jand g16408(.dina(n33670), .dinb(n33669), .dout(n33671));
  jor  g16409(.dina(n33671), .dinb(n33388), .dout(n33672));
  jxor g16410(.dina(n33382), .dinb(n325), .dout(n33673));
  jand g16411(.dina(n33673), .dinb(n33672), .dout(n33674));
  jor  g16412(.dina(n33674), .dinb(n33383), .dout(n33675));
  jxor g16413(.dina(n33377), .dinb(n326), .dout(n33676));
  jand g16414(.dina(n33676), .dinb(n33675), .dout(n33677));
  jor  g16415(.dina(n33677), .dinb(n33378), .dout(n33678));
  jxor g16416(.dina(n33372), .dinb(n277), .dout(n33679));
  jand g16417(.dina(n33679), .dinb(n33678), .dout(n33680));
  jor  g16418(.dina(n33680), .dinb(n33373), .dout(n33681));
  jxor g16419(.dina(n33367), .dinb(n278), .dout(n33682));
  jand g16420(.dina(n33682), .dinb(n33681), .dout(n33683));
  jor  g16421(.dina(n33683), .dinb(n33368), .dout(n33684));
  jxor g16422(.dina(n33362), .dinb(n279), .dout(n33685));
  jand g16423(.dina(n33685), .dinb(n33684), .dout(n33686));
  jor  g16424(.dina(n33686), .dinb(n33363), .dout(n33687));
  jxor g16425(.dina(n33357), .dinb(n280), .dout(n33688));
  jand g16426(.dina(n33688), .dinb(n33687), .dout(n33689));
  jor  g16427(.dina(n33689), .dinb(n33358), .dout(n33690));
  jxor g16428(.dina(n33352), .dinb(n283), .dout(n33691));
  jand g16429(.dina(n33691), .dinb(n33690), .dout(n33692));
  jor  g16430(.dina(n33692), .dinb(n33353), .dout(n33693));
  jxor g16431(.dina(n33347), .dinb(n315), .dout(n33694));
  jand g16432(.dina(n33694), .dinb(n33693), .dout(n33695));
  jor  g16433(.dina(n33695), .dinb(n33348), .dout(n33696));
  jxor g16434(.dina(n33342), .dinb(n316), .dout(n33697));
  jand g16435(.dina(n33697), .dinb(n33696), .dout(n33698));
  jor  g16436(.dina(n33698), .dinb(n33343), .dout(n33699));
  jxor g16437(.dina(n33337), .dinb(n317), .dout(n33700));
  jand g16438(.dina(n33700), .dinb(n33699), .dout(n33701));
  jor  g16439(.dina(n33701), .dinb(n33338), .dout(n33702));
  jxor g16440(.dina(n33332), .dinb(n284), .dout(n33703));
  jand g16441(.dina(n33703), .dinb(n33702), .dout(n33704));
  jor  g16442(.dina(n33704), .dinb(n33333), .dout(n33705));
  jxor g16443(.dina(n33327), .dinb(n285), .dout(n33706));
  jand g16444(.dina(n33706), .dinb(n33705), .dout(n33707));
  jor  g16445(.dina(n33707), .dinb(n33328), .dout(n33708));
  jxor g16446(.dina(n33322), .dinb(n286), .dout(n33709));
  jand g16447(.dina(n33709), .dinb(n33708), .dout(n33710));
  jor  g16448(.dina(n33710), .dinb(n33323), .dout(n33711));
  jxor g16449(.dina(n33317), .dinb(n287), .dout(n33712));
  jand g16450(.dina(n33712), .dinb(n33711), .dout(n33713));
  jor  g16451(.dina(n33713), .dinb(n33318), .dout(n33714));
  jxor g16452(.dina(n33312), .dinb(n288), .dout(n33715));
  jand g16453(.dina(n33715), .dinb(n33714), .dout(n33716));
  jor  g16454(.dina(n33716), .dinb(n33313), .dout(n33717));
  jxor g16455(.dina(n33307), .dinb(n289), .dout(n33718));
  jand g16456(.dina(n33718), .dinb(n33717), .dout(n33719));
  jor  g16457(.dina(n33719), .dinb(n33308), .dout(n33720));
  jxor g16458(.dina(n33295), .dinb(n290), .dout(n33721));
  jand g16459(.dina(n33721), .dinb(n33720), .dout(n33722));
  jor  g16460(.dina(n33722), .dinb(n33303), .dout(n33723));
  jand g16461(.dina(n33723), .dinb(n33302), .dout(n33724));
  jor  g16462(.dina(n33724), .dinb(n33299), .dout(n33725));
  jand g16463(.dina(n33725), .dinb(n306), .dout(n33726));
  jor  g16464(.dina(n33726), .dinb(n33295), .dout(n33727));
  jnot g16465(.din(n33726), .dout(n33728));
  jxor g16466(.dina(n33721), .dinb(n33720), .dout(n33729));
  jor  g16467(.dina(n33729), .dinb(n33728), .dout(n33730));
  jand g16468(.dina(n33730), .dinb(n33727), .dout(n33731));
  jand g16469(.dina(n33728), .dinb(n33298), .dout(n33732));
  jand g16470(.dina(n33723), .dinb(n33299), .dout(n33733));
  jand g16471(.dina(n33733), .dinb(n306), .dout(n33734));
  jor  g16472(.dina(n33734), .dinb(n33732), .dout(n33735));
  jand g16473(.dina(n33735), .dinb(n306), .dout(n33736));
  jnot g16474(.din(n33735), .dout(n33737));
  jand g16475(.dina(n33737), .dinb(n292), .dout(n33738));
  jand g16476(.dina(n33298), .dinb(b55 ), .dout(n33739));
  jor  g16477(.dina(n33739), .dinb(n33738), .dout(n33740));
  jand g16478(.dina(n33731), .dinb(n291), .dout(n33741));
  jor  g16479(.dina(n33726), .dinb(n33307), .dout(n33742));
  jxor g16480(.dina(n33718), .dinb(n33717), .dout(n33743));
  jor  g16481(.dina(n33743), .dinb(n33728), .dout(n33744));
  jand g16482(.dina(n33744), .dinb(n33742), .dout(n33745));
  jand g16483(.dina(n33745), .dinb(n290), .dout(n33746));
  jor  g16484(.dina(n33726), .dinb(n33312), .dout(n33747));
  jxor g16485(.dina(n33715), .dinb(n33714), .dout(n33748));
  jor  g16486(.dina(n33748), .dinb(n33728), .dout(n33749));
  jand g16487(.dina(n33749), .dinb(n33747), .dout(n33750));
  jand g16488(.dina(n33750), .dinb(n289), .dout(n33751));
  jor  g16489(.dina(n33726), .dinb(n33317), .dout(n33752));
  jxor g16490(.dina(n33712), .dinb(n33711), .dout(n33753));
  jor  g16491(.dina(n33753), .dinb(n33728), .dout(n33754));
  jand g16492(.dina(n33754), .dinb(n33752), .dout(n33755));
  jand g16493(.dina(n33755), .dinb(n288), .dout(n33756));
  jor  g16494(.dina(n33726), .dinb(n33322), .dout(n33757));
  jxor g16495(.dina(n33709), .dinb(n33708), .dout(n33758));
  jor  g16496(.dina(n33758), .dinb(n33728), .dout(n33759));
  jand g16497(.dina(n33759), .dinb(n33757), .dout(n33760));
  jand g16498(.dina(n33760), .dinb(n287), .dout(n33761));
  jor  g16499(.dina(n33726), .dinb(n33327), .dout(n33762));
  jxor g16500(.dina(n33706), .dinb(n33705), .dout(n33763));
  jor  g16501(.dina(n33763), .dinb(n33728), .dout(n33764));
  jand g16502(.dina(n33764), .dinb(n33762), .dout(n33765));
  jand g16503(.dina(n33765), .dinb(n286), .dout(n33766));
  jor  g16504(.dina(n33726), .dinb(n33332), .dout(n33767));
  jxor g16505(.dina(n33703), .dinb(n33702), .dout(n33768));
  jor  g16506(.dina(n33768), .dinb(n33728), .dout(n33769));
  jand g16507(.dina(n33769), .dinb(n33767), .dout(n33770));
  jand g16508(.dina(n33770), .dinb(n285), .dout(n33771));
  jor  g16509(.dina(n33726), .dinb(n33337), .dout(n33772));
  jxor g16510(.dina(n33700), .dinb(n33699), .dout(n33773));
  jor  g16511(.dina(n33773), .dinb(n33728), .dout(n33774));
  jand g16512(.dina(n33774), .dinb(n33772), .dout(n33775));
  jand g16513(.dina(n33775), .dinb(n284), .dout(n33776));
  jor  g16514(.dina(n33726), .dinb(n33342), .dout(n33777));
  jxor g16515(.dina(n33697), .dinb(n33696), .dout(n33778));
  jor  g16516(.dina(n33778), .dinb(n33728), .dout(n33779));
  jand g16517(.dina(n33779), .dinb(n33777), .dout(n33780));
  jand g16518(.dina(n33780), .dinb(n317), .dout(n33781));
  jor  g16519(.dina(n33726), .dinb(n33347), .dout(n33782));
  jxor g16520(.dina(n33694), .dinb(n33693), .dout(n33783));
  jor  g16521(.dina(n33783), .dinb(n33728), .dout(n33784));
  jand g16522(.dina(n33784), .dinb(n33782), .dout(n33785));
  jand g16523(.dina(n33785), .dinb(n316), .dout(n33786));
  jor  g16524(.dina(n33726), .dinb(n33352), .dout(n33787));
  jxor g16525(.dina(n33691), .dinb(n33690), .dout(n33788));
  jor  g16526(.dina(n33788), .dinb(n33728), .dout(n33789));
  jand g16527(.dina(n33789), .dinb(n33787), .dout(n33790));
  jand g16528(.dina(n33790), .dinb(n315), .dout(n33791));
  jor  g16529(.dina(n33726), .dinb(n33357), .dout(n33792));
  jxor g16530(.dina(n33688), .dinb(n33687), .dout(n33793));
  jor  g16531(.dina(n33793), .dinb(n33728), .dout(n33794));
  jand g16532(.dina(n33794), .dinb(n33792), .dout(n33795));
  jand g16533(.dina(n33795), .dinb(n283), .dout(n33796));
  jor  g16534(.dina(n33726), .dinb(n33362), .dout(n33797));
  jxor g16535(.dina(n33685), .dinb(n33684), .dout(n33798));
  jor  g16536(.dina(n33798), .dinb(n33728), .dout(n33799));
  jand g16537(.dina(n33799), .dinb(n33797), .dout(n33800));
  jand g16538(.dina(n33800), .dinb(n280), .dout(n33801));
  jor  g16539(.dina(n33726), .dinb(n33367), .dout(n33802));
  jxor g16540(.dina(n33682), .dinb(n33681), .dout(n33803));
  jor  g16541(.dina(n33803), .dinb(n33728), .dout(n33804));
  jand g16542(.dina(n33804), .dinb(n33802), .dout(n33805));
  jand g16543(.dina(n33805), .dinb(n279), .dout(n33806));
  jor  g16544(.dina(n33726), .dinb(n33372), .dout(n33807));
  jxor g16545(.dina(n33679), .dinb(n33678), .dout(n33808));
  jor  g16546(.dina(n33808), .dinb(n33728), .dout(n33809));
  jand g16547(.dina(n33809), .dinb(n33807), .dout(n33810));
  jand g16548(.dina(n33810), .dinb(n278), .dout(n33811));
  jor  g16549(.dina(n33726), .dinb(n33377), .dout(n33812));
  jxor g16550(.dina(n33676), .dinb(n33675), .dout(n33813));
  jor  g16551(.dina(n33813), .dinb(n33728), .dout(n33814));
  jand g16552(.dina(n33814), .dinb(n33812), .dout(n33815));
  jand g16553(.dina(n33815), .dinb(n277), .dout(n33816));
  jor  g16554(.dina(n33726), .dinb(n33382), .dout(n33817));
  jxor g16555(.dina(n33673), .dinb(n33672), .dout(n33818));
  jor  g16556(.dina(n33818), .dinb(n33728), .dout(n33819));
  jand g16557(.dina(n33819), .dinb(n33817), .dout(n33820));
  jand g16558(.dina(n33820), .dinb(n326), .dout(n33821));
  jor  g16559(.dina(n33726), .dinb(n33387), .dout(n33822));
  jxor g16560(.dina(n33670), .dinb(n33669), .dout(n33823));
  jor  g16561(.dina(n33823), .dinb(n33728), .dout(n33824));
  jand g16562(.dina(n33824), .dinb(n33822), .dout(n33825));
  jand g16563(.dina(n33825), .dinb(n325), .dout(n33826));
  jor  g16564(.dina(n33726), .dinb(n33392), .dout(n33827));
  jxor g16565(.dina(n33667), .dinb(n33666), .dout(n33828));
  jor  g16566(.dina(n33828), .dinb(n33728), .dout(n33829));
  jand g16567(.dina(n33829), .dinb(n33827), .dout(n33830));
  jand g16568(.dina(n33830), .dinb(n324), .dout(n33831));
  jor  g16569(.dina(n33726), .dinb(n33397), .dout(n33832));
  jxor g16570(.dina(n33664), .dinb(n33663), .dout(n33833));
  jor  g16571(.dina(n33833), .dinb(n33728), .dout(n33834));
  jand g16572(.dina(n33834), .dinb(n33832), .dout(n33835));
  jand g16573(.dina(n33835), .dinb(n276), .dout(n33836));
  jor  g16574(.dina(n33726), .dinb(n33402), .dout(n33837));
  jxor g16575(.dina(n33661), .dinb(n33660), .dout(n33838));
  jor  g16576(.dina(n33838), .dinb(n33728), .dout(n33839));
  jand g16577(.dina(n33839), .dinb(n33837), .dout(n33840));
  jand g16578(.dina(n33840), .dinb(n333), .dout(n33841));
  jor  g16579(.dina(n33726), .dinb(n33407), .dout(n33842));
  jxor g16580(.dina(n33658), .dinb(n33657), .dout(n33843));
  jor  g16581(.dina(n33843), .dinb(n33728), .dout(n33844));
  jand g16582(.dina(n33844), .dinb(n33842), .dout(n33845));
  jand g16583(.dina(n33845), .dinb(n332), .dout(n33846));
  jor  g16584(.dina(n33726), .dinb(n33412), .dout(n33847));
  jxor g16585(.dina(n33655), .dinb(n33654), .dout(n33848));
  jor  g16586(.dina(n33848), .dinb(n33728), .dout(n33849));
  jand g16587(.dina(n33849), .dinb(n33847), .dout(n33850));
  jand g16588(.dina(n33850), .dinb(n331), .dout(n33851));
  jor  g16589(.dina(n33726), .dinb(n33417), .dout(n33852));
  jxor g16590(.dina(n33652), .dinb(n33651), .dout(n33853));
  jor  g16591(.dina(n33853), .dinb(n33728), .dout(n33854));
  jand g16592(.dina(n33854), .dinb(n33852), .dout(n33855));
  jand g16593(.dina(n33855), .dinb(n275), .dout(n33856));
  jor  g16594(.dina(n33726), .dinb(n33422), .dout(n33857));
  jxor g16595(.dina(n33649), .dinb(n33648), .dout(n33858));
  jor  g16596(.dina(n33858), .dinb(n33728), .dout(n33859));
  jand g16597(.dina(n33859), .dinb(n33857), .dout(n33860));
  jand g16598(.dina(n33860), .dinb(n340), .dout(n33861));
  jor  g16599(.dina(n33726), .dinb(n33427), .dout(n33862));
  jxor g16600(.dina(n33646), .dinb(n33645), .dout(n33863));
  jor  g16601(.dina(n33863), .dinb(n33728), .dout(n33864));
  jand g16602(.dina(n33864), .dinb(n33862), .dout(n33865));
  jand g16603(.dina(n33865), .dinb(n339), .dout(n33866));
  jor  g16604(.dina(n33726), .dinb(n33432), .dout(n33867));
  jxor g16605(.dina(n33643), .dinb(n33642), .dout(n33868));
  jor  g16606(.dina(n33868), .dinb(n33728), .dout(n33869));
  jand g16607(.dina(n33869), .dinb(n33867), .dout(n33870));
  jand g16608(.dina(n33870), .dinb(n338), .dout(n33871));
  jor  g16609(.dina(n33726), .dinb(n33437), .dout(n33872));
  jxor g16610(.dina(n33640), .dinb(n33639), .dout(n33873));
  jor  g16611(.dina(n33873), .dinb(n33728), .dout(n33874));
  jand g16612(.dina(n33874), .dinb(n33872), .dout(n33875));
  jand g16613(.dina(n33875), .dinb(n271), .dout(n33876));
  jor  g16614(.dina(n33726), .dinb(n33442), .dout(n33877));
  jxor g16615(.dina(n33637), .dinb(n33636), .dout(n33878));
  jor  g16616(.dina(n33878), .dinb(n33728), .dout(n33879));
  jand g16617(.dina(n33879), .dinb(n33877), .dout(n33880));
  jand g16618(.dina(n33880), .dinb(n270), .dout(n33881));
  jor  g16619(.dina(n33726), .dinb(n33447), .dout(n33882));
  jxor g16620(.dina(n33634), .dinb(n33633), .dout(n33883));
  jor  g16621(.dina(n33883), .dinb(n33728), .dout(n33884));
  jand g16622(.dina(n33884), .dinb(n33882), .dout(n33885));
  jand g16623(.dina(n33885), .dinb(n269), .dout(n33886));
  jor  g16624(.dina(n33726), .dinb(n33452), .dout(n33887));
  jxor g16625(.dina(n33631), .dinb(n33630), .dout(n33888));
  jor  g16626(.dina(n33888), .dinb(n33728), .dout(n33889));
  jand g16627(.dina(n33889), .dinb(n33887), .dout(n33890));
  jand g16628(.dina(n33890), .dinb(n274), .dout(n33891));
  jor  g16629(.dina(n33726), .dinb(n33457), .dout(n33892));
  jxor g16630(.dina(n33628), .dinb(n33627), .dout(n33893));
  jor  g16631(.dina(n33893), .dinb(n33728), .dout(n33894));
  jand g16632(.dina(n33894), .dinb(n33892), .dout(n33895));
  jand g16633(.dina(n33895), .dinb(n268), .dout(n33896));
  jor  g16634(.dina(n33726), .dinb(n33462), .dout(n33897));
  jxor g16635(.dina(n33625), .dinb(n33624), .dout(n33898));
  jor  g16636(.dina(n33898), .dinb(n33728), .dout(n33899));
  jand g16637(.dina(n33899), .dinb(n33897), .dout(n33900));
  jand g16638(.dina(n33900), .dinb(n349), .dout(n33901));
  jor  g16639(.dina(n33726), .dinb(n33467), .dout(n33902));
  jxor g16640(.dina(n33622), .dinb(n33621), .dout(n33903));
  jor  g16641(.dina(n33903), .dinb(n33728), .dout(n33904));
  jand g16642(.dina(n33904), .dinb(n33902), .dout(n33905));
  jand g16643(.dina(n33905), .dinb(n348), .dout(n33906));
  jor  g16644(.dina(n33726), .dinb(n33472), .dout(n33907));
  jxor g16645(.dina(n33619), .dinb(n33618), .dout(n33908));
  jor  g16646(.dina(n33908), .dinb(n33728), .dout(n33909));
  jand g16647(.dina(n33909), .dinb(n33907), .dout(n33910));
  jand g16648(.dina(n33910), .dinb(n347), .dout(n33911));
  jor  g16649(.dina(n33726), .dinb(n33477), .dout(n33912));
  jxor g16650(.dina(n33616), .dinb(n33615), .dout(n33913));
  jor  g16651(.dina(n33913), .dinb(n33728), .dout(n33914));
  jand g16652(.dina(n33914), .dinb(n33912), .dout(n33915));
  jand g16653(.dina(n33915), .dinb(n267), .dout(n33916));
  jor  g16654(.dina(n33726), .dinb(n33482), .dout(n33917));
  jxor g16655(.dina(n33613), .dinb(n33612), .dout(n33918));
  jor  g16656(.dina(n33918), .dinb(n33728), .dout(n33919));
  jand g16657(.dina(n33919), .dinb(n33917), .dout(n33920));
  jand g16658(.dina(n33920), .dinb(n266), .dout(n33921));
  jor  g16659(.dina(n33726), .dinb(n33487), .dout(n33922));
  jxor g16660(.dina(n33610), .dinb(n33609), .dout(n33923));
  jor  g16661(.dina(n33923), .dinb(n33728), .dout(n33924));
  jand g16662(.dina(n33924), .dinb(n33922), .dout(n33925));
  jand g16663(.dina(n33925), .dinb(n356), .dout(n33926));
  jor  g16664(.dina(n33726), .dinb(n33492), .dout(n33927));
  jxor g16665(.dina(n33607), .dinb(n33606), .dout(n33928));
  jor  g16666(.dina(n33928), .dinb(n33728), .dout(n33929));
  jand g16667(.dina(n33929), .dinb(n33927), .dout(n33930));
  jand g16668(.dina(n33930), .dinb(n355), .dout(n33931));
  jor  g16669(.dina(n33726), .dinb(n33497), .dout(n33932));
  jxor g16670(.dina(n33604), .dinb(n33603), .dout(n33933));
  jor  g16671(.dina(n33933), .dinb(n33728), .dout(n33934));
  jand g16672(.dina(n33934), .dinb(n33932), .dout(n33935));
  jand g16673(.dina(n33935), .dinb(n364), .dout(n33936));
  jor  g16674(.dina(n33726), .dinb(n33502), .dout(n33937));
  jxor g16675(.dina(n33601), .dinb(n33600), .dout(n33938));
  jor  g16676(.dina(n33938), .dinb(n33728), .dout(n33939));
  jand g16677(.dina(n33939), .dinb(n33937), .dout(n33940));
  jand g16678(.dina(n33940), .dinb(n361), .dout(n33941));
  jor  g16679(.dina(n33726), .dinb(n33507), .dout(n33942));
  jxor g16680(.dina(n33598), .dinb(n33597), .dout(n33943));
  jor  g16681(.dina(n33943), .dinb(n33728), .dout(n33944));
  jand g16682(.dina(n33944), .dinb(n33942), .dout(n33945));
  jand g16683(.dina(n33945), .dinb(n360), .dout(n33946));
  jor  g16684(.dina(n33726), .dinb(n33512), .dout(n33947));
  jxor g16685(.dina(n33595), .dinb(n33594), .dout(n33948));
  jor  g16686(.dina(n33948), .dinb(n33728), .dout(n33949));
  jand g16687(.dina(n33949), .dinb(n33947), .dout(n33950));
  jand g16688(.dina(n33950), .dinb(n363), .dout(n33951));
  jor  g16689(.dina(n33726), .dinb(n33517), .dout(n33952));
  jxor g16690(.dina(n33592), .dinb(n33591), .dout(n33953));
  jor  g16691(.dina(n33953), .dinb(n33728), .dout(n33954));
  jand g16692(.dina(n33954), .dinb(n33952), .dout(n33955));
  jand g16693(.dina(n33955), .dinb(n359), .dout(n33956));
  jor  g16694(.dina(n33726), .dinb(n33522), .dout(n33957));
  jxor g16695(.dina(n33589), .dinb(n33588), .dout(n33958));
  jor  g16696(.dina(n33958), .dinb(n33728), .dout(n33959));
  jand g16697(.dina(n33959), .dinb(n33957), .dout(n33960));
  jand g16698(.dina(n33960), .dinb(n369), .dout(n33961));
  jor  g16699(.dina(n33726), .dinb(n33527), .dout(n33962));
  jxor g16700(.dina(n33586), .dinb(n33585), .dout(n33963));
  jor  g16701(.dina(n33963), .dinb(n33728), .dout(n33964));
  jand g16702(.dina(n33964), .dinb(n33962), .dout(n33965));
  jand g16703(.dina(n33965), .dinb(n368), .dout(n33966));
  jor  g16704(.dina(n33726), .dinb(n33532), .dout(n33967));
  jxor g16705(.dina(n33583), .dinb(n33582), .dout(n33968));
  jor  g16706(.dina(n33968), .dinb(n33728), .dout(n33969));
  jand g16707(.dina(n33969), .dinb(n33967), .dout(n33970));
  jand g16708(.dina(n33970), .dinb(n367), .dout(n33971));
  jor  g16709(.dina(n33726), .dinb(n33537), .dout(n33972));
  jxor g16710(.dina(n33580), .dinb(n33579), .dout(n33973));
  jor  g16711(.dina(n33973), .dinb(n33728), .dout(n33974));
  jand g16712(.dina(n33974), .dinb(n33972), .dout(n33975));
  jand g16713(.dina(n33975), .dinb(n265), .dout(n33976));
  jor  g16714(.dina(n33726), .dinb(n33542), .dout(n33977));
  jxor g16715(.dina(n33577), .dinb(n33576), .dout(n33978));
  jor  g16716(.dina(n33978), .dinb(n33728), .dout(n33979));
  jand g16717(.dina(n33979), .dinb(n33977), .dout(n33980));
  jand g16718(.dina(n33980), .dinb(n378), .dout(n33981));
  jor  g16719(.dina(n33726), .dinb(n33547), .dout(n33982));
  jxor g16720(.dina(n33574), .dinb(n33573), .dout(n33983));
  jor  g16721(.dina(n33983), .dinb(n33728), .dout(n33984));
  jand g16722(.dina(n33984), .dinb(n33982), .dout(n33985));
  jand g16723(.dina(n33985), .dinb(n377), .dout(n33986));
  jor  g16724(.dina(n33726), .dinb(n33552), .dout(n33987));
  jxor g16725(.dina(n33571), .dinb(n33570), .dout(n33988));
  jor  g16726(.dina(n33988), .dinb(n33728), .dout(n33989));
  jand g16727(.dina(n33989), .dinb(n33987), .dout(n33990));
  jand g16728(.dina(n33990), .dinb(n376), .dout(n33991));
  jor  g16729(.dina(n33726), .dinb(n33559), .dout(n33992));
  jxor g16730(.dina(n33568), .dinb(n33567), .dout(n33993));
  jor  g16731(.dina(n33993), .dinb(n33728), .dout(n33994));
  jand g16732(.dina(n33994), .dinb(n33992), .dout(n33995));
  jand g16733(.dina(n33995), .dinb(n264), .dout(n33996));
  jor  g16734(.dina(n33726), .dinb(n33564), .dout(n33997));
  jxor g16735(.dina(n33565), .dinb(n13302), .dout(n33998));
  jand g16736(.dina(n33998), .dinb(n33726), .dout(n33999));
  jnot g16737(.din(n33999), .dout(n34000));
  jand g16738(.dina(n34000), .dinb(n33997), .dout(n34001));
  jnot g16739(.din(n34001), .dout(n34002));
  jand g16740(.dina(n34002), .dinb(n386), .dout(n34003));
  jnot g16741(.din(n13732), .dout(n34004));
  jnot g16742(.din(n33299), .dout(n34005));
  jnot g16743(.din(n33303), .dout(n34006));
  jnot g16744(.din(n33308), .dout(n34007));
  jnot g16745(.din(n33313), .dout(n34008));
  jnot g16746(.din(n33318), .dout(n34009));
  jnot g16747(.din(n33323), .dout(n34010));
  jnot g16748(.din(n33328), .dout(n34011));
  jnot g16749(.din(n33333), .dout(n34012));
  jnot g16750(.din(n33338), .dout(n34013));
  jnot g16751(.din(n33343), .dout(n34014));
  jnot g16752(.din(n33348), .dout(n34015));
  jnot g16753(.din(n33353), .dout(n34016));
  jnot g16754(.din(n33358), .dout(n34017));
  jnot g16755(.din(n33363), .dout(n34018));
  jnot g16756(.din(n33368), .dout(n34019));
  jnot g16757(.din(n33373), .dout(n34020));
  jnot g16758(.din(n33378), .dout(n34021));
  jnot g16759(.din(n33383), .dout(n34022));
  jnot g16760(.din(n33388), .dout(n34023));
  jnot g16761(.din(n33393), .dout(n34024));
  jnot g16762(.din(n33398), .dout(n34025));
  jnot g16763(.din(n33403), .dout(n34026));
  jnot g16764(.din(n33408), .dout(n34027));
  jnot g16765(.din(n33413), .dout(n34028));
  jnot g16766(.din(n33418), .dout(n34029));
  jnot g16767(.din(n33423), .dout(n34030));
  jnot g16768(.din(n33428), .dout(n34031));
  jnot g16769(.din(n33433), .dout(n34032));
  jnot g16770(.din(n33438), .dout(n34033));
  jnot g16771(.din(n33443), .dout(n34034));
  jnot g16772(.din(n33448), .dout(n34035));
  jnot g16773(.din(n33453), .dout(n34036));
  jnot g16774(.din(n33458), .dout(n34037));
  jnot g16775(.din(n33463), .dout(n34038));
  jnot g16776(.din(n33468), .dout(n34039));
  jnot g16777(.din(n33473), .dout(n34040));
  jnot g16778(.din(n33478), .dout(n34041));
  jnot g16779(.din(n33483), .dout(n34042));
  jnot g16780(.din(n33488), .dout(n34043));
  jnot g16781(.din(n33493), .dout(n34044));
  jnot g16782(.din(n33498), .dout(n34045));
  jnot g16783(.din(n33503), .dout(n34046));
  jnot g16784(.din(n33508), .dout(n34047));
  jnot g16785(.din(n33513), .dout(n34048));
  jnot g16786(.din(n33518), .dout(n34049));
  jnot g16787(.din(n33523), .dout(n34050));
  jnot g16788(.din(n33528), .dout(n34051));
  jnot g16789(.din(n33533), .dout(n34052));
  jnot g16790(.din(n33538), .dout(n34053));
  jnot g16791(.din(n33543), .dout(n34054));
  jnot g16792(.din(n33548), .dout(n34055));
  jnot g16793(.din(n33553), .dout(n34056));
  jnot g16794(.din(n33560), .dout(n34057));
  jnot g16795(.din(n33563), .dout(n34058));
  jxor g16796(.dina(n33564), .dinb(n259), .dout(n34059));
  jor  g16797(.dina(n34059), .dinb(n13301), .dout(n34060));
  jand g16798(.dina(n34060), .dinb(n34058), .dout(n34061));
  jnot g16799(.din(n33568), .dout(n34062));
  jor  g16800(.dina(n34062), .dinb(n34061), .dout(n34063));
  jand g16801(.dina(n34063), .dinb(n34057), .dout(n34064));
  jnot g16802(.din(n33571), .dout(n34065));
  jor  g16803(.dina(n34065), .dinb(n34064), .dout(n34066));
  jand g16804(.dina(n34066), .dinb(n34056), .dout(n34067));
  jnot g16805(.din(n33574), .dout(n34068));
  jor  g16806(.dina(n34068), .dinb(n34067), .dout(n34069));
  jand g16807(.dina(n34069), .dinb(n34055), .dout(n34070));
  jnot g16808(.din(n33577), .dout(n34071));
  jor  g16809(.dina(n34071), .dinb(n34070), .dout(n34072));
  jand g16810(.dina(n34072), .dinb(n34054), .dout(n34073));
  jnot g16811(.din(n33580), .dout(n34074));
  jor  g16812(.dina(n34074), .dinb(n34073), .dout(n34075));
  jand g16813(.dina(n34075), .dinb(n34053), .dout(n34076));
  jnot g16814(.din(n33583), .dout(n34077));
  jor  g16815(.dina(n34077), .dinb(n34076), .dout(n34078));
  jand g16816(.dina(n34078), .dinb(n34052), .dout(n34079));
  jnot g16817(.din(n33586), .dout(n34080));
  jor  g16818(.dina(n34080), .dinb(n34079), .dout(n34081));
  jand g16819(.dina(n34081), .dinb(n34051), .dout(n34082));
  jnot g16820(.din(n33589), .dout(n34083));
  jor  g16821(.dina(n34083), .dinb(n34082), .dout(n34084));
  jand g16822(.dina(n34084), .dinb(n34050), .dout(n34085));
  jnot g16823(.din(n33592), .dout(n34086));
  jor  g16824(.dina(n34086), .dinb(n34085), .dout(n34087));
  jand g16825(.dina(n34087), .dinb(n34049), .dout(n34088));
  jnot g16826(.din(n33595), .dout(n34089));
  jor  g16827(.dina(n34089), .dinb(n34088), .dout(n34090));
  jand g16828(.dina(n34090), .dinb(n34048), .dout(n34091));
  jnot g16829(.din(n33598), .dout(n34092));
  jor  g16830(.dina(n34092), .dinb(n34091), .dout(n34093));
  jand g16831(.dina(n34093), .dinb(n34047), .dout(n34094));
  jnot g16832(.din(n33601), .dout(n34095));
  jor  g16833(.dina(n34095), .dinb(n34094), .dout(n34096));
  jand g16834(.dina(n34096), .dinb(n34046), .dout(n34097));
  jnot g16835(.din(n33604), .dout(n34098));
  jor  g16836(.dina(n34098), .dinb(n34097), .dout(n34099));
  jand g16837(.dina(n34099), .dinb(n34045), .dout(n34100));
  jnot g16838(.din(n33607), .dout(n34101));
  jor  g16839(.dina(n34101), .dinb(n34100), .dout(n34102));
  jand g16840(.dina(n34102), .dinb(n34044), .dout(n34103));
  jnot g16841(.din(n33610), .dout(n34104));
  jor  g16842(.dina(n34104), .dinb(n34103), .dout(n34105));
  jand g16843(.dina(n34105), .dinb(n34043), .dout(n34106));
  jnot g16844(.din(n33613), .dout(n34107));
  jor  g16845(.dina(n34107), .dinb(n34106), .dout(n34108));
  jand g16846(.dina(n34108), .dinb(n34042), .dout(n34109));
  jnot g16847(.din(n33616), .dout(n34110));
  jor  g16848(.dina(n34110), .dinb(n34109), .dout(n34111));
  jand g16849(.dina(n34111), .dinb(n34041), .dout(n34112));
  jnot g16850(.din(n33619), .dout(n34113));
  jor  g16851(.dina(n34113), .dinb(n34112), .dout(n34114));
  jand g16852(.dina(n34114), .dinb(n34040), .dout(n34115));
  jnot g16853(.din(n33622), .dout(n34116));
  jor  g16854(.dina(n34116), .dinb(n34115), .dout(n34117));
  jand g16855(.dina(n34117), .dinb(n34039), .dout(n34118));
  jnot g16856(.din(n33625), .dout(n34119));
  jor  g16857(.dina(n34119), .dinb(n34118), .dout(n34120));
  jand g16858(.dina(n34120), .dinb(n34038), .dout(n34121));
  jnot g16859(.din(n33628), .dout(n34122));
  jor  g16860(.dina(n34122), .dinb(n34121), .dout(n34123));
  jand g16861(.dina(n34123), .dinb(n34037), .dout(n34124));
  jnot g16862(.din(n33631), .dout(n34125));
  jor  g16863(.dina(n34125), .dinb(n34124), .dout(n34126));
  jand g16864(.dina(n34126), .dinb(n34036), .dout(n34127));
  jnot g16865(.din(n33634), .dout(n34128));
  jor  g16866(.dina(n34128), .dinb(n34127), .dout(n34129));
  jand g16867(.dina(n34129), .dinb(n34035), .dout(n34130));
  jnot g16868(.din(n33637), .dout(n34131));
  jor  g16869(.dina(n34131), .dinb(n34130), .dout(n34132));
  jand g16870(.dina(n34132), .dinb(n34034), .dout(n34133));
  jnot g16871(.din(n33640), .dout(n34134));
  jor  g16872(.dina(n34134), .dinb(n34133), .dout(n34135));
  jand g16873(.dina(n34135), .dinb(n34033), .dout(n34136));
  jnot g16874(.din(n33643), .dout(n34137));
  jor  g16875(.dina(n34137), .dinb(n34136), .dout(n34138));
  jand g16876(.dina(n34138), .dinb(n34032), .dout(n34139));
  jnot g16877(.din(n33646), .dout(n34140));
  jor  g16878(.dina(n34140), .dinb(n34139), .dout(n34141));
  jand g16879(.dina(n34141), .dinb(n34031), .dout(n34142));
  jnot g16880(.din(n33649), .dout(n34143));
  jor  g16881(.dina(n34143), .dinb(n34142), .dout(n34144));
  jand g16882(.dina(n34144), .dinb(n34030), .dout(n34145));
  jnot g16883(.din(n33652), .dout(n34146));
  jor  g16884(.dina(n34146), .dinb(n34145), .dout(n34147));
  jand g16885(.dina(n34147), .dinb(n34029), .dout(n34148));
  jnot g16886(.din(n33655), .dout(n34149));
  jor  g16887(.dina(n34149), .dinb(n34148), .dout(n34150));
  jand g16888(.dina(n34150), .dinb(n34028), .dout(n34151));
  jnot g16889(.din(n33658), .dout(n34152));
  jor  g16890(.dina(n34152), .dinb(n34151), .dout(n34153));
  jand g16891(.dina(n34153), .dinb(n34027), .dout(n34154));
  jnot g16892(.din(n33661), .dout(n34155));
  jor  g16893(.dina(n34155), .dinb(n34154), .dout(n34156));
  jand g16894(.dina(n34156), .dinb(n34026), .dout(n34157));
  jnot g16895(.din(n33664), .dout(n34158));
  jor  g16896(.dina(n34158), .dinb(n34157), .dout(n34159));
  jand g16897(.dina(n34159), .dinb(n34025), .dout(n34160));
  jnot g16898(.din(n33667), .dout(n34161));
  jor  g16899(.dina(n34161), .dinb(n34160), .dout(n34162));
  jand g16900(.dina(n34162), .dinb(n34024), .dout(n34163));
  jnot g16901(.din(n33670), .dout(n34164));
  jor  g16902(.dina(n34164), .dinb(n34163), .dout(n34165));
  jand g16903(.dina(n34165), .dinb(n34023), .dout(n34166));
  jnot g16904(.din(n33673), .dout(n34167));
  jor  g16905(.dina(n34167), .dinb(n34166), .dout(n34168));
  jand g16906(.dina(n34168), .dinb(n34022), .dout(n34169));
  jnot g16907(.din(n33676), .dout(n34170));
  jor  g16908(.dina(n34170), .dinb(n34169), .dout(n34171));
  jand g16909(.dina(n34171), .dinb(n34021), .dout(n34172));
  jnot g16910(.din(n33679), .dout(n34173));
  jor  g16911(.dina(n34173), .dinb(n34172), .dout(n34174));
  jand g16912(.dina(n34174), .dinb(n34020), .dout(n34175));
  jnot g16913(.din(n33682), .dout(n34176));
  jor  g16914(.dina(n34176), .dinb(n34175), .dout(n34177));
  jand g16915(.dina(n34177), .dinb(n34019), .dout(n34178));
  jnot g16916(.din(n33685), .dout(n34179));
  jor  g16917(.dina(n34179), .dinb(n34178), .dout(n34180));
  jand g16918(.dina(n34180), .dinb(n34018), .dout(n34181));
  jnot g16919(.din(n33688), .dout(n34182));
  jor  g16920(.dina(n34182), .dinb(n34181), .dout(n34183));
  jand g16921(.dina(n34183), .dinb(n34017), .dout(n34184));
  jnot g16922(.din(n33691), .dout(n34185));
  jor  g16923(.dina(n34185), .dinb(n34184), .dout(n34186));
  jand g16924(.dina(n34186), .dinb(n34016), .dout(n34187));
  jnot g16925(.din(n33694), .dout(n34188));
  jor  g16926(.dina(n34188), .dinb(n34187), .dout(n34189));
  jand g16927(.dina(n34189), .dinb(n34015), .dout(n34190));
  jnot g16928(.din(n33697), .dout(n34191));
  jor  g16929(.dina(n34191), .dinb(n34190), .dout(n34192));
  jand g16930(.dina(n34192), .dinb(n34014), .dout(n34193));
  jnot g16931(.din(n33700), .dout(n34194));
  jor  g16932(.dina(n34194), .dinb(n34193), .dout(n34195));
  jand g16933(.dina(n34195), .dinb(n34013), .dout(n34196));
  jnot g16934(.din(n33703), .dout(n34197));
  jor  g16935(.dina(n34197), .dinb(n34196), .dout(n34198));
  jand g16936(.dina(n34198), .dinb(n34012), .dout(n34199));
  jnot g16937(.din(n33706), .dout(n34200));
  jor  g16938(.dina(n34200), .dinb(n34199), .dout(n34201));
  jand g16939(.dina(n34201), .dinb(n34011), .dout(n34202));
  jnot g16940(.din(n33709), .dout(n34203));
  jor  g16941(.dina(n34203), .dinb(n34202), .dout(n34204));
  jand g16942(.dina(n34204), .dinb(n34010), .dout(n34205));
  jnot g16943(.din(n33712), .dout(n34206));
  jor  g16944(.dina(n34206), .dinb(n34205), .dout(n34207));
  jand g16945(.dina(n34207), .dinb(n34009), .dout(n34208));
  jnot g16946(.din(n33715), .dout(n34209));
  jor  g16947(.dina(n34209), .dinb(n34208), .dout(n34210));
  jand g16948(.dina(n34210), .dinb(n34008), .dout(n34211));
  jnot g16949(.din(n33718), .dout(n34212));
  jor  g16950(.dina(n34212), .dinb(n34211), .dout(n34213));
  jand g16951(.dina(n34213), .dinb(n34007), .dout(n34214));
  jnot g16952(.din(n33721), .dout(n34215));
  jor  g16953(.dina(n34215), .dinb(n34214), .dout(n34216));
  jand g16954(.dina(n34216), .dinb(n34006), .dout(n34217));
  jor  g16955(.dina(n34217), .dinb(n33301), .dout(n34218));
  jand g16956(.dina(n34218), .dinb(n34005), .dout(n34219));
  jor  g16957(.dina(n34219), .dinb(n34004), .dout(n34220));
  jand g16958(.dina(n34220), .dinb(a9 ), .dout(n34221));
  jnot g16959(.din(n13735), .dout(n34222));
  jor  g16960(.dina(n34219), .dinb(n34222), .dout(n34223));
  jnot g16961(.din(n34223), .dout(n34224));
  jor  g16962(.dina(n34224), .dinb(n34221), .dout(n34225));
  jand g16963(.dina(n34225), .dinb(n259), .dout(n34226));
  jand g16964(.dina(n33725), .dinb(n13732), .dout(n34227));
  jor  g16965(.dina(n34227), .dinb(n13300), .dout(n34228));
  jand g16966(.dina(n34223), .dinb(n34228), .dout(n34229));
  jxor g16967(.dina(n34229), .dinb(b1 ), .dout(n34230));
  jand g16968(.dina(n34230), .dinb(n13743), .dout(n34231));
  jor  g16969(.dina(n34231), .dinb(n34226), .dout(n34232));
  jxor g16970(.dina(n34001), .dinb(b2 ), .dout(n34233));
  jand g16971(.dina(n34233), .dinb(n34232), .dout(n34234));
  jor  g16972(.dina(n34234), .dinb(n34003), .dout(n34235));
  jxor g16973(.dina(n33995), .dinb(n264), .dout(n34236));
  jand g16974(.dina(n34236), .dinb(n34235), .dout(n34237));
  jor  g16975(.dina(n34237), .dinb(n33996), .dout(n34238));
  jxor g16976(.dina(n33990), .dinb(n376), .dout(n34239));
  jand g16977(.dina(n34239), .dinb(n34238), .dout(n34240));
  jor  g16978(.dina(n34240), .dinb(n33991), .dout(n34241));
  jxor g16979(.dina(n33985), .dinb(n377), .dout(n34242));
  jand g16980(.dina(n34242), .dinb(n34241), .dout(n34243));
  jor  g16981(.dina(n34243), .dinb(n33986), .dout(n34244));
  jxor g16982(.dina(n33980), .dinb(n378), .dout(n34245));
  jand g16983(.dina(n34245), .dinb(n34244), .dout(n34246));
  jor  g16984(.dina(n34246), .dinb(n33981), .dout(n34247));
  jxor g16985(.dina(n33975), .dinb(n265), .dout(n34248));
  jand g16986(.dina(n34248), .dinb(n34247), .dout(n34249));
  jor  g16987(.dina(n34249), .dinb(n33976), .dout(n34250));
  jxor g16988(.dina(n33970), .dinb(n367), .dout(n34251));
  jand g16989(.dina(n34251), .dinb(n34250), .dout(n34252));
  jor  g16990(.dina(n34252), .dinb(n33971), .dout(n34253));
  jxor g16991(.dina(n33965), .dinb(n368), .dout(n34254));
  jand g16992(.dina(n34254), .dinb(n34253), .dout(n34255));
  jor  g16993(.dina(n34255), .dinb(n33966), .dout(n34256));
  jxor g16994(.dina(n33960), .dinb(n369), .dout(n34257));
  jand g16995(.dina(n34257), .dinb(n34256), .dout(n34258));
  jor  g16996(.dina(n34258), .dinb(n33961), .dout(n34259));
  jxor g16997(.dina(n33955), .dinb(n359), .dout(n34260));
  jand g16998(.dina(n34260), .dinb(n34259), .dout(n34261));
  jor  g16999(.dina(n34261), .dinb(n33956), .dout(n34262));
  jxor g17000(.dina(n33950), .dinb(n363), .dout(n34263));
  jand g17001(.dina(n34263), .dinb(n34262), .dout(n34264));
  jor  g17002(.dina(n34264), .dinb(n33951), .dout(n34265));
  jxor g17003(.dina(n33945), .dinb(n360), .dout(n34266));
  jand g17004(.dina(n34266), .dinb(n34265), .dout(n34267));
  jor  g17005(.dina(n34267), .dinb(n33946), .dout(n34268));
  jxor g17006(.dina(n33940), .dinb(n361), .dout(n34269));
  jand g17007(.dina(n34269), .dinb(n34268), .dout(n34270));
  jor  g17008(.dina(n34270), .dinb(n33941), .dout(n34271));
  jxor g17009(.dina(n33935), .dinb(n364), .dout(n34272));
  jand g17010(.dina(n34272), .dinb(n34271), .dout(n34273));
  jor  g17011(.dina(n34273), .dinb(n33936), .dout(n34274));
  jxor g17012(.dina(n33930), .dinb(n355), .dout(n34275));
  jand g17013(.dina(n34275), .dinb(n34274), .dout(n34276));
  jor  g17014(.dina(n34276), .dinb(n33931), .dout(n34277));
  jxor g17015(.dina(n33925), .dinb(n356), .dout(n34278));
  jand g17016(.dina(n34278), .dinb(n34277), .dout(n34279));
  jor  g17017(.dina(n34279), .dinb(n33926), .dout(n34280));
  jxor g17018(.dina(n33920), .dinb(n266), .dout(n34281));
  jand g17019(.dina(n34281), .dinb(n34280), .dout(n34282));
  jor  g17020(.dina(n34282), .dinb(n33921), .dout(n34283));
  jxor g17021(.dina(n33915), .dinb(n267), .dout(n34284));
  jand g17022(.dina(n34284), .dinb(n34283), .dout(n34285));
  jor  g17023(.dina(n34285), .dinb(n33916), .dout(n34286));
  jxor g17024(.dina(n33910), .dinb(n347), .dout(n34287));
  jand g17025(.dina(n34287), .dinb(n34286), .dout(n34288));
  jor  g17026(.dina(n34288), .dinb(n33911), .dout(n34289));
  jxor g17027(.dina(n33905), .dinb(n348), .dout(n34290));
  jand g17028(.dina(n34290), .dinb(n34289), .dout(n34291));
  jor  g17029(.dina(n34291), .dinb(n33906), .dout(n34292));
  jxor g17030(.dina(n33900), .dinb(n349), .dout(n34293));
  jand g17031(.dina(n34293), .dinb(n34292), .dout(n34294));
  jor  g17032(.dina(n34294), .dinb(n33901), .dout(n34295));
  jxor g17033(.dina(n33895), .dinb(n268), .dout(n34296));
  jand g17034(.dina(n34296), .dinb(n34295), .dout(n34297));
  jor  g17035(.dina(n34297), .dinb(n33896), .dout(n34298));
  jxor g17036(.dina(n33890), .dinb(n274), .dout(n34299));
  jand g17037(.dina(n34299), .dinb(n34298), .dout(n34300));
  jor  g17038(.dina(n34300), .dinb(n33891), .dout(n34301));
  jxor g17039(.dina(n33885), .dinb(n269), .dout(n34302));
  jand g17040(.dina(n34302), .dinb(n34301), .dout(n34303));
  jor  g17041(.dina(n34303), .dinb(n33886), .dout(n34304));
  jxor g17042(.dina(n33880), .dinb(n270), .dout(n34305));
  jand g17043(.dina(n34305), .dinb(n34304), .dout(n34306));
  jor  g17044(.dina(n34306), .dinb(n33881), .dout(n34307));
  jxor g17045(.dina(n33875), .dinb(n271), .dout(n34308));
  jand g17046(.dina(n34308), .dinb(n34307), .dout(n34309));
  jor  g17047(.dina(n34309), .dinb(n33876), .dout(n34310));
  jxor g17048(.dina(n33870), .dinb(n338), .dout(n34311));
  jand g17049(.dina(n34311), .dinb(n34310), .dout(n34312));
  jor  g17050(.dina(n34312), .dinb(n33871), .dout(n34313));
  jxor g17051(.dina(n33865), .dinb(n339), .dout(n34314));
  jand g17052(.dina(n34314), .dinb(n34313), .dout(n34315));
  jor  g17053(.dina(n34315), .dinb(n33866), .dout(n34316));
  jxor g17054(.dina(n33860), .dinb(n340), .dout(n34317));
  jand g17055(.dina(n34317), .dinb(n34316), .dout(n34318));
  jor  g17056(.dina(n34318), .dinb(n33861), .dout(n34319));
  jxor g17057(.dina(n33855), .dinb(n275), .dout(n34320));
  jand g17058(.dina(n34320), .dinb(n34319), .dout(n34321));
  jor  g17059(.dina(n34321), .dinb(n33856), .dout(n34322));
  jxor g17060(.dina(n33850), .dinb(n331), .dout(n34323));
  jand g17061(.dina(n34323), .dinb(n34322), .dout(n34324));
  jor  g17062(.dina(n34324), .dinb(n33851), .dout(n34325));
  jxor g17063(.dina(n33845), .dinb(n332), .dout(n34326));
  jand g17064(.dina(n34326), .dinb(n34325), .dout(n34327));
  jor  g17065(.dina(n34327), .dinb(n33846), .dout(n34328));
  jxor g17066(.dina(n33840), .dinb(n333), .dout(n34329));
  jand g17067(.dina(n34329), .dinb(n34328), .dout(n34330));
  jor  g17068(.dina(n34330), .dinb(n33841), .dout(n34331));
  jxor g17069(.dina(n33835), .dinb(n276), .dout(n34332));
  jand g17070(.dina(n34332), .dinb(n34331), .dout(n34333));
  jor  g17071(.dina(n34333), .dinb(n33836), .dout(n34334));
  jxor g17072(.dina(n33830), .dinb(n324), .dout(n34335));
  jand g17073(.dina(n34335), .dinb(n34334), .dout(n34336));
  jor  g17074(.dina(n34336), .dinb(n33831), .dout(n34337));
  jxor g17075(.dina(n33825), .dinb(n325), .dout(n34338));
  jand g17076(.dina(n34338), .dinb(n34337), .dout(n34339));
  jor  g17077(.dina(n34339), .dinb(n33826), .dout(n34340));
  jxor g17078(.dina(n33820), .dinb(n326), .dout(n34341));
  jand g17079(.dina(n34341), .dinb(n34340), .dout(n34342));
  jor  g17080(.dina(n34342), .dinb(n33821), .dout(n34343));
  jxor g17081(.dina(n33815), .dinb(n277), .dout(n34344));
  jand g17082(.dina(n34344), .dinb(n34343), .dout(n34345));
  jor  g17083(.dina(n34345), .dinb(n33816), .dout(n34346));
  jxor g17084(.dina(n33810), .dinb(n278), .dout(n34347));
  jand g17085(.dina(n34347), .dinb(n34346), .dout(n34348));
  jor  g17086(.dina(n34348), .dinb(n33811), .dout(n34349));
  jxor g17087(.dina(n33805), .dinb(n279), .dout(n34350));
  jand g17088(.dina(n34350), .dinb(n34349), .dout(n34351));
  jor  g17089(.dina(n34351), .dinb(n33806), .dout(n34352));
  jxor g17090(.dina(n33800), .dinb(n280), .dout(n34353));
  jand g17091(.dina(n34353), .dinb(n34352), .dout(n34354));
  jor  g17092(.dina(n34354), .dinb(n33801), .dout(n34355));
  jxor g17093(.dina(n33795), .dinb(n283), .dout(n34356));
  jand g17094(.dina(n34356), .dinb(n34355), .dout(n34357));
  jor  g17095(.dina(n34357), .dinb(n33796), .dout(n34358));
  jxor g17096(.dina(n33790), .dinb(n315), .dout(n34359));
  jand g17097(.dina(n34359), .dinb(n34358), .dout(n34360));
  jor  g17098(.dina(n34360), .dinb(n33791), .dout(n34361));
  jxor g17099(.dina(n33785), .dinb(n316), .dout(n34362));
  jand g17100(.dina(n34362), .dinb(n34361), .dout(n34363));
  jor  g17101(.dina(n34363), .dinb(n33786), .dout(n34364));
  jxor g17102(.dina(n33780), .dinb(n317), .dout(n34365));
  jand g17103(.dina(n34365), .dinb(n34364), .dout(n34366));
  jor  g17104(.dina(n34366), .dinb(n33781), .dout(n34367));
  jxor g17105(.dina(n33775), .dinb(n284), .dout(n34368));
  jand g17106(.dina(n34368), .dinb(n34367), .dout(n34369));
  jor  g17107(.dina(n34369), .dinb(n33776), .dout(n34370));
  jxor g17108(.dina(n33770), .dinb(n285), .dout(n34371));
  jand g17109(.dina(n34371), .dinb(n34370), .dout(n34372));
  jor  g17110(.dina(n34372), .dinb(n33771), .dout(n34373));
  jxor g17111(.dina(n33765), .dinb(n286), .dout(n34374));
  jand g17112(.dina(n34374), .dinb(n34373), .dout(n34375));
  jor  g17113(.dina(n34375), .dinb(n33766), .dout(n34376));
  jxor g17114(.dina(n33760), .dinb(n287), .dout(n34377));
  jand g17115(.dina(n34377), .dinb(n34376), .dout(n34378));
  jor  g17116(.dina(n34378), .dinb(n33761), .dout(n34379));
  jxor g17117(.dina(n33755), .dinb(n288), .dout(n34380));
  jand g17118(.dina(n34380), .dinb(n34379), .dout(n34381));
  jor  g17119(.dina(n34381), .dinb(n33756), .dout(n34382));
  jxor g17120(.dina(n33750), .dinb(n289), .dout(n34383));
  jand g17121(.dina(n34383), .dinb(n34382), .dout(n34384));
  jor  g17122(.dina(n34384), .dinb(n33751), .dout(n34385));
  jxor g17123(.dina(n33745), .dinb(n290), .dout(n34386));
  jand g17124(.dina(n34386), .dinb(n34385), .dout(n34387));
  jor  g17125(.dina(n34387), .dinb(n33746), .dout(n34388));
  jxor g17126(.dina(n33731), .dinb(n291), .dout(n34389));
  jand g17127(.dina(n34389), .dinb(n34388), .dout(n34390));
  jor  g17128(.dina(n34390), .dinb(n33741), .dout(n34391));
  jand g17129(.dina(n34391), .dinb(n305), .dout(n34392));
  jand g17130(.dina(n34392), .dinb(n33740), .dout(n34393));
  jor  g17131(.dina(n34393), .dinb(n33736), .dout(n34394));
  jor  g17132(.dina(n34394), .dinb(n33731), .dout(n34395));
  jnot g17133(.din(n34394), .dout(n34396));
  jxor g17134(.dina(n34389), .dinb(n34388), .dout(n34397));
  jor  g17135(.dina(n34397), .dinb(n34396), .dout(n34398));
  jand g17136(.dina(n34398), .dinb(n34395), .dout(n34399));
  jxor g17137(.dina(n34391), .dinb(n33740), .dout(n34400));
  jand g17138(.dina(n34400), .dinb(n306), .dout(n34401));
  jor  g17139(.dina(n34401), .dinb(n34396), .dout(n34402));
  jand g17140(.dina(n34402), .dinb(n33735), .dout(n34403));
  jand g17141(.dina(n34403), .dinb(n293), .dout(n34404));
  jxor g17142(.dina(n34403), .dinb(n293), .dout(n34405));
  jand g17143(.dina(n34399), .dinb(n292), .dout(n34406));
  jor  g17144(.dina(n34394), .dinb(n33745), .dout(n34407));
  jxor g17145(.dina(n34386), .dinb(n34385), .dout(n34408));
  jor  g17146(.dina(n34408), .dinb(n34396), .dout(n34409));
  jand g17147(.dina(n34409), .dinb(n34407), .dout(n34410));
  jand g17148(.dina(n34410), .dinb(n291), .dout(n34411));
  jor  g17149(.dina(n34394), .dinb(n33750), .dout(n34412));
  jxor g17150(.dina(n34383), .dinb(n34382), .dout(n34413));
  jor  g17151(.dina(n34413), .dinb(n34396), .dout(n34414));
  jand g17152(.dina(n34414), .dinb(n34412), .dout(n34415));
  jand g17153(.dina(n34415), .dinb(n290), .dout(n34416));
  jor  g17154(.dina(n34394), .dinb(n33755), .dout(n34417));
  jxor g17155(.dina(n34380), .dinb(n34379), .dout(n34418));
  jor  g17156(.dina(n34418), .dinb(n34396), .dout(n34419));
  jand g17157(.dina(n34419), .dinb(n34417), .dout(n34420));
  jand g17158(.dina(n34420), .dinb(n289), .dout(n34421));
  jor  g17159(.dina(n34394), .dinb(n33760), .dout(n34422));
  jxor g17160(.dina(n34377), .dinb(n34376), .dout(n34423));
  jor  g17161(.dina(n34423), .dinb(n34396), .dout(n34424));
  jand g17162(.dina(n34424), .dinb(n34422), .dout(n34425));
  jand g17163(.dina(n34425), .dinb(n288), .dout(n34426));
  jor  g17164(.dina(n34394), .dinb(n33765), .dout(n34427));
  jxor g17165(.dina(n34374), .dinb(n34373), .dout(n34428));
  jor  g17166(.dina(n34428), .dinb(n34396), .dout(n34429));
  jand g17167(.dina(n34429), .dinb(n34427), .dout(n34430));
  jand g17168(.dina(n34430), .dinb(n287), .dout(n34431));
  jor  g17169(.dina(n34394), .dinb(n33770), .dout(n34432));
  jxor g17170(.dina(n34371), .dinb(n34370), .dout(n34433));
  jor  g17171(.dina(n34433), .dinb(n34396), .dout(n34434));
  jand g17172(.dina(n34434), .dinb(n34432), .dout(n34435));
  jand g17173(.dina(n34435), .dinb(n286), .dout(n34436));
  jor  g17174(.dina(n34394), .dinb(n33775), .dout(n34437));
  jxor g17175(.dina(n34368), .dinb(n34367), .dout(n34438));
  jor  g17176(.dina(n34438), .dinb(n34396), .dout(n34439));
  jand g17177(.dina(n34439), .dinb(n34437), .dout(n34440));
  jand g17178(.dina(n34440), .dinb(n285), .dout(n34441));
  jor  g17179(.dina(n34394), .dinb(n33780), .dout(n34442));
  jxor g17180(.dina(n34365), .dinb(n34364), .dout(n34443));
  jor  g17181(.dina(n34443), .dinb(n34396), .dout(n34444));
  jand g17182(.dina(n34444), .dinb(n34442), .dout(n34445));
  jand g17183(.dina(n34445), .dinb(n284), .dout(n34446));
  jor  g17184(.dina(n34394), .dinb(n33785), .dout(n34447));
  jxor g17185(.dina(n34362), .dinb(n34361), .dout(n34448));
  jor  g17186(.dina(n34448), .dinb(n34396), .dout(n34449));
  jand g17187(.dina(n34449), .dinb(n34447), .dout(n34450));
  jand g17188(.dina(n34450), .dinb(n317), .dout(n34451));
  jor  g17189(.dina(n34394), .dinb(n33790), .dout(n34452));
  jxor g17190(.dina(n34359), .dinb(n34358), .dout(n34453));
  jor  g17191(.dina(n34453), .dinb(n34396), .dout(n34454));
  jand g17192(.dina(n34454), .dinb(n34452), .dout(n34455));
  jand g17193(.dina(n34455), .dinb(n316), .dout(n34456));
  jor  g17194(.dina(n34394), .dinb(n33795), .dout(n34457));
  jxor g17195(.dina(n34356), .dinb(n34355), .dout(n34458));
  jor  g17196(.dina(n34458), .dinb(n34396), .dout(n34459));
  jand g17197(.dina(n34459), .dinb(n34457), .dout(n34460));
  jand g17198(.dina(n34460), .dinb(n315), .dout(n34461));
  jor  g17199(.dina(n34394), .dinb(n33800), .dout(n34462));
  jxor g17200(.dina(n34353), .dinb(n34352), .dout(n34463));
  jor  g17201(.dina(n34463), .dinb(n34396), .dout(n34464));
  jand g17202(.dina(n34464), .dinb(n34462), .dout(n34465));
  jand g17203(.dina(n34465), .dinb(n283), .dout(n34466));
  jor  g17204(.dina(n34394), .dinb(n33805), .dout(n34467));
  jxor g17205(.dina(n34350), .dinb(n34349), .dout(n34468));
  jor  g17206(.dina(n34468), .dinb(n34396), .dout(n34469));
  jand g17207(.dina(n34469), .dinb(n34467), .dout(n34470));
  jand g17208(.dina(n34470), .dinb(n280), .dout(n34471));
  jor  g17209(.dina(n34394), .dinb(n33810), .dout(n34472));
  jxor g17210(.dina(n34347), .dinb(n34346), .dout(n34473));
  jor  g17211(.dina(n34473), .dinb(n34396), .dout(n34474));
  jand g17212(.dina(n34474), .dinb(n34472), .dout(n34475));
  jand g17213(.dina(n34475), .dinb(n279), .dout(n34476));
  jor  g17214(.dina(n34394), .dinb(n33815), .dout(n34477));
  jxor g17215(.dina(n34344), .dinb(n34343), .dout(n34478));
  jor  g17216(.dina(n34478), .dinb(n34396), .dout(n34479));
  jand g17217(.dina(n34479), .dinb(n34477), .dout(n34480));
  jand g17218(.dina(n34480), .dinb(n278), .dout(n34481));
  jor  g17219(.dina(n34394), .dinb(n33820), .dout(n34482));
  jxor g17220(.dina(n34341), .dinb(n34340), .dout(n34483));
  jor  g17221(.dina(n34483), .dinb(n34396), .dout(n34484));
  jand g17222(.dina(n34484), .dinb(n34482), .dout(n34485));
  jand g17223(.dina(n34485), .dinb(n277), .dout(n34486));
  jor  g17224(.dina(n34394), .dinb(n33825), .dout(n34487));
  jxor g17225(.dina(n34338), .dinb(n34337), .dout(n34488));
  jor  g17226(.dina(n34488), .dinb(n34396), .dout(n34489));
  jand g17227(.dina(n34489), .dinb(n34487), .dout(n34490));
  jand g17228(.dina(n34490), .dinb(n326), .dout(n34491));
  jor  g17229(.dina(n34394), .dinb(n33830), .dout(n34492));
  jxor g17230(.dina(n34335), .dinb(n34334), .dout(n34493));
  jor  g17231(.dina(n34493), .dinb(n34396), .dout(n34494));
  jand g17232(.dina(n34494), .dinb(n34492), .dout(n34495));
  jand g17233(.dina(n34495), .dinb(n325), .dout(n34496));
  jor  g17234(.dina(n34394), .dinb(n33835), .dout(n34497));
  jxor g17235(.dina(n34332), .dinb(n34331), .dout(n34498));
  jor  g17236(.dina(n34498), .dinb(n34396), .dout(n34499));
  jand g17237(.dina(n34499), .dinb(n34497), .dout(n34500));
  jand g17238(.dina(n34500), .dinb(n324), .dout(n34501));
  jor  g17239(.dina(n34394), .dinb(n33840), .dout(n34502));
  jxor g17240(.dina(n34329), .dinb(n34328), .dout(n34503));
  jor  g17241(.dina(n34503), .dinb(n34396), .dout(n34504));
  jand g17242(.dina(n34504), .dinb(n34502), .dout(n34505));
  jand g17243(.dina(n34505), .dinb(n276), .dout(n34506));
  jor  g17244(.dina(n34394), .dinb(n33845), .dout(n34507));
  jxor g17245(.dina(n34326), .dinb(n34325), .dout(n34508));
  jor  g17246(.dina(n34508), .dinb(n34396), .dout(n34509));
  jand g17247(.dina(n34509), .dinb(n34507), .dout(n34510));
  jand g17248(.dina(n34510), .dinb(n333), .dout(n34511));
  jor  g17249(.dina(n34394), .dinb(n33850), .dout(n34512));
  jxor g17250(.dina(n34323), .dinb(n34322), .dout(n34513));
  jor  g17251(.dina(n34513), .dinb(n34396), .dout(n34514));
  jand g17252(.dina(n34514), .dinb(n34512), .dout(n34515));
  jand g17253(.dina(n34515), .dinb(n332), .dout(n34516));
  jor  g17254(.dina(n34394), .dinb(n33855), .dout(n34517));
  jxor g17255(.dina(n34320), .dinb(n34319), .dout(n34518));
  jor  g17256(.dina(n34518), .dinb(n34396), .dout(n34519));
  jand g17257(.dina(n34519), .dinb(n34517), .dout(n34520));
  jand g17258(.dina(n34520), .dinb(n331), .dout(n34521));
  jor  g17259(.dina(n34394), .dinb(n33860), .dout(n34522));
  jxor g17260(.dina(n34317), .dinb(n34316), .dout(n34523));
  jor  g17261(.dina(n34523), .dinb(n34396), .dout(n34524));
  jand g17262(.dina(n34524), .dinb(n34522), .dout(n34525));
  jand g17263(.dina(n34525), .dinb(n275), .dout(n34526));
  jor  g17264(.dina(n34394), .dinb(n33865), .dout(n34527));
  jxor g17265(.dina(n34314), .dinb(n34313), .dout(n34528));
  jor  g17266(.dina(n34528), .dinb(n34396), .dout(n34529));
  jand g17267(.dina(n34529), .dinb(n34527), .dout(n34530));
  jand g17268(.dina(n34530), .dinb(n340), .dout(n34531));
  jor  g17269(.dina(n34394), .dinb(n33870), .dout(n34532));
  jxor g17270(.dina(n34311), .dinb(n34310), .dout(n34533));
  jor  g17271(.dina(n34533), .dinb(n34396), .dout(n34534));
  jand g17272(.dina(n34534), .dinb(n34532), .dout(n34535));
  jand g17273(.dina(n34535), .dinb(n339), .dout(n34536));
  jor  g17274(.dina(n34394), .dinb(n33875), .dout(n34537));
  jxor g17275(.dina(n34308), .dinb(n34307), .dout(n34538));
  jor  g17276(.dina(n34538), .dinb(n34396), .dout(n34539));
  jand g17277(.dina(n34539), .dinb(n34537), .dout(n34540));
  jand g17278(.dina(n34540), .dinb(n338), .dout(n34541));
  jor  g17279(.dina(n34394), .dinb(n33880), .dout(n34542));
  jxor g17280(.dina(n34305), .dinb(n34304), .dout(n34543));
  jor  g17281(.dina(n34543), .dinb(n34396), .dout(n34544));
  jand g17282(.dina(n34544), .dinb(n34542), .dout(n34545));
  jand g17283(.dina(n34545), .dinb(n271), .dout(n34546));
  jor  g17284(.dina(n34394), .dinb(n33885), .dout(n34547));
  jxor g17285(.dina(n34302), .dinb(n34301), .dout(n34548));
  jor  g17286(.dina(n34548), .dinb(n34396), .dout(n34549));
  jand g17287(.dina(n34549), .dinb(n34547), .dout(n34550));
  jand g17288(.dina(n34550), .dinb(n270), .dout(n34551));
  jor  g17289(.dina(n34394), .dinb(n33890), .dout(n34552));
  jxor g17290(.dina(n34299), .dinb(n34298), .dout(n34553));
  jor  g17291(.dina(n34553), .dinb(n34396), .dout(n34554));
  jand g17292(.dina(n34554), .dinb(n34552), .dout(n34555));
  jand g17293(.dina(n34555), .dinb(n269), .dout(n34556));
  jor  g17294(.dina(n34394), .dinb(n33895), .dout(n34557));
  jxor g17295(.dina(n34296), .dinb(n34295), .dout(n34558));
  jor  g17296(.dina(n34558), .dinb(n34396), .dout(n34559));
  jand g17297(.dina(n34559), .dinb(n34557), .dout(n34560));
  jand g17298(.dina(n34560), .dinb(n274), .dout(n34561));
  jor  g17299(.dina(n34394), .dinb(n33900), .dout(n34562));
  jxor g17300(.dina(n34293), .dinb(n34292), .dout(n34563));
  jor  g17301(.dina(n34563), .dinb(n34396), .dout(n34564));
  jand g17302(.dina(n34564), .dinb(n34562), .dout(n34565));
  jand g17303(.dina(n34565), .dinb(n268), .dout(n34566));
  jor  g17304(.dina(n34394), .dinb(n33905), .dout(n34567));
  jxor g17305(.dina(n34290), .dinb(n34289), .dout(n34568));
  jor  g17306(.dina(n34568), .dinb(n34396), .dout(n34569));
  jand g17307(.dina(n34569), .dinb(n34567), .dout(n34570));
  jand g17308(.dina(n34570), .dinb(n349), .dout(n34571));
  jor  g17309(.dina(n34394), .dinb(n33910), .dout(n34572));
  jxor g17310(.dina(n34287), .dinb(n34286), .dout(n34573));
  jor  g17311(.dina(n34573), .dinb(n34396), .dout(n34574));
  jand g17312(.dina(n34574), .dinb(n34572), .dout(n34575));
  jand g17313(.dina(n34575), .dinb(n348), .dout(n34576));
  jor  g17314(.dina(n34394), .dinb(n33915), .dout(n34577));
  jxor g17315(.dina(n34284), .dinb(n34283), .dout(n34578));
  jor  g17316(.dina(n34578), .dinb(n34396), .dout(n34579));
  jand g17317(.dina(n34579), .dinb(n34577), .dout(n34580));
  jand g17318(.dina(n34580), .dinb(n347), .dout(n34581));
  jor  g17319(.dina(n34394), .dinb(n33920), .dout(n34582));
  jxor g17320(.dina(n34281), .dinb(n34280), .dout(n34583));
  jor  g17321(.dina(n34583), .dinb(n34396), .dout(n34584));
  jand g17322(.dina(n34584), .dinb(n34582), .dout(n34585));
  jand g17323(.dina(n34585), .dinb(n267), .dout(n34586));
  jor  g17324(.dina(n34394), .dinb(n33925), .dout(n34587));
  jxor g17325(.dina(n34278), .dinb(n34277), .dout(n34588));
  jor  g17326(.dina(n34588), .dinb(n34396), .dout(n34589));
  jand g17327(.dina(n34589), .dinb(n34587), .dout(n34590));
  jand g17328(.dina(n34590), .dinb(n266), .dout(n34591));
  jor  g17329(.dina(n34394), .dinb(n33930), .dout(n34592));
  jxor g17330(.dina(n34275), .dinb(n34274), .dout(n34593));
  jor  g17331(.dina(n34593), .dinb(n34396), .dout(n34594));
  jand g17332(.dina(n34594), .dinb(n34592), .dout(n34595));
  jand g17333(.dina(n34595), .dinb(n356), .dout(n34596));
  jor  g17334(.dina(n34394), .dinb(n33935), .dout(n34597));
  jxor g17335(.dina(n34272), .dinb(n34271), .dout(n34598));
  jor  g17336(.dina(n34598), .dinb(n34396), .dout(n34599));
  jand g17337(.dina(n34599), .dinb(n34597), .dout(n34600));
  jand g17338(.dina(n34600), .dinb(n355), .dout(n34601));
  jor  g17339(.dina(n34394), .dinb(n33940), .dout(n34602));
  jxor g17340(.dina(n34269), .dinb(n34268), .dout(n34603));
  jor  g17341(.dina(n34603), .dinb(n34396), .dout(n34604));
  jand g17342(.dina(n34604), .dinb(n34602), .dout(n34605));
  jand g17343(.dina(n34605), .dinb(n364), .dout(n34606));
  jor  g17344(.dina(n34394), .dinb(n33945), .dout(n34607));
  jxor g17345(.dina(n34266), .dinb(n34265), .dout(n34608));
  jor  g17346(.dina(n34608), .dinb(n34396), .dout(n34609));
  jand g17347(.dina(n34609), .dinb(n34607), .dout(n34610));
  jand g17348(.dina(n34610), .dinb(n361), .dout(n34611));
  jor  g17349(.dina(n34394), .dinb(n33950), .dout(n34612));
  jxor g17350(.dina(n34263), .dinb(n34262), .dout(n34613));
  jor  g17351(.dina(n34613), .dinb(n34396), .dout(n34614));
  jand g17352(.dina(n34614), .dinb(n34612), .dout(n34615));
  jand g17353(.dina(n34615), .dinb(n360), .dout(n34616));
  jor  g17354(.dina(n34394), .dinb(n33955), .dout(n34617));
  jxor g17355(.dina(n34260), .dinb(n34259), .dout(n34618));
  jor  g17356(.dina(n34618), .dinb(n34396), .dout(n34619));
  jand g17357(.dina(n34619), .dinb(n34617), .dout(n34620));
  jand g17358(.dina(n34620), .dinb(n363), .dout(n34621));
  jor  g17359(.dina(n34394), .dinb(n33960), .dout(n34622));
  jxor g17360(.dina(n34257), .dinb(n34256), .dout(n34623));
  jor  g17361(.dina(n34623), .dinb(n34396), .dout(n34624));
  jand g17362(.dina(n34624), .dinb(n34622), .dout(n34625));
  jand g17363(.dina(n34625), .dinb(n359), .dout(n34626));
  jor  g17364(.dina(n34394), .dinb(n33965), .dout(n34627));
  jxor g17365(.dina(n34254), .dinb(n34253), .dout(n34628));
  jor  g17366(.dina(n34628), .dinb(n34396), .dout(n34629));
  jand g17367(.dina(n34629), .dinb(n34627), .dout(n34630));
  jand g17368(.dina(n34630), .dinb(n369), .dout(n34631));
  jor  g17369(.dina(n34394), .dinb(n33970), .dout(n34632));
  jxor g17370(.dina(n34251), .dinb(n34250), .dout(n34633));
  jor  g17371(.dina(n34633), .dinb(n34396), .dout(n34634));
  jand g17372(.dina(n34634), .dinb(n34632), .dout(n34635));
  jand g17373(.dina(n34635), .dinb(n368), .dout(n34636));
  jor  g17374(.dina(n34394), .dinb(n33975), .dout(n34637));
  jxor g17375(.dina(n34248), .dinb(n34247), .dout(n34638));
  jor  g17376(.dina(n34638), .dinb(n34396), .dout(n34639));
  jand g17377(.dina(n34639), .dinb(n34637), .dout(n34640));
  jand g17378(.dina(n34640), .dinb(n367), .dout(n34641));
  jor  g17379(.dina(n34394), .dinb(n33980), .dout(n34642));
  jxor g17380(.dina(n34245), .dinb(n34244), .dout(n34643));
  jor  g17381(.dina(n34643), .dinb(n34396), .dout(n34644));
  jand g17382(.dina(n34644), .dinb(n34642), .dout(n34645));
  jand g17383(.dina(n34645), .dinb(n265), .dout(n34646));
  jor  g17384(.dina(n34394), .dinb(n33985), .dout(n34647));
  jxor g17385(.dina(n34242), .dinb(n34241), .dout(n34648));
  jor  g17386(.dina(n34648), .dinb(n34396), .dout(n34649));
  jand g17387(.dina(n34649), .dinb(n34647), .dout(n34650));
  jand g17388(.dina(n34650), .dinb(n378), .dout(n34651));
  jor  g17389(.dina(n34394), .dinb(n33990), .dout(n34652));
  jxor g17390(.dina(n34239), .dinb(n34238), .dout(n34653));
  jor  g17391(.dina(n34653), .dinb(n34396), .dout(n34654));
  jand g17392(.dina(n34654), .dinb(n34652), .dout(n34655));
  jand g17393(.dina(n34655), .dinb(n377), .dout(n34656));
  jor  g17394(.dina(n34394), .dinb(n33995), .dout(n34657));
  jxor g17395(.dina(n34236), .dinb(n34235), .dout(n34658));
  jor  g17396(.dina(n34658), .dinb(n34396), .dout(n34659));
  jand g17397(.dina(n34659), .dinb(n34657), .dout(n34660));
  jand g17398(.dina(n34660), .dinb(n376), .dout(n34661));
  jor  g17399(.dina(n34394), .dinb(n34001), .dout(n34662));
  jxor g17400(.dina(n34233), .dinb(n34232), .dout(n34663));
  jnot g17401(.din(n34663), .dout(n34664));
  jor  g17402(.dina(n34664), .dinb(n34396), .dout(n34665));
  jand g17403(.dina(n34665), .dinb(n34662), .dout(n34666));
  jnot g17404(.din(n34666), .dout(n34667));
  jand g17405(.dina(n34667), .dinb(n264), .dout(n34668));
  jor  g17406(.dina(n34394), .dinb(n34225), .dout(n34669));
  jxor g17407(.dina(n34230), .dinb(n13743), .dout(n34670));
  jor  g17408(.dina(n34670), .dinb(n34396), .dout(n34671));
  jand g17409(.dina(n34671), .dinb(n34669), .dout(n34672));
  jand g17410(.dina(n34672), .dinb(n386), .dout(n34673));
  jand g17411(.dina(n34394), .dinb(b0 ), .dout(n34674));
  jxor g17412(.dina(n34674), .dinb(a8 ), .dout(n34675));
  jand g17413(.dina(n34675), .dinb(n259), .dout(n34676));
  jxor g17414(.dina(n34674), .dinb(n13741), .dout(n34677));
  jxor g17415(.dina(n34677), .dinb(b1 ), .dout(n34678));
  jand g17416(.dina(n34678), .dinb(n14205), .dout(n34679));
  jor  g17417(.dina(n34679), .dinb(n34676), .dout(n34680));
  jxor g17418(.dina(n34672), .dinb(n386), .dout(n34681));
  jand g17419(.dina(n34681), .dinb(n34680), .dout(n34682));
  jor  g17420(.dina(n34682), .dinb(n34673), .dout(n34683));
  jxor g17421(.dina(n34666), .dinb(b3 ), .dout(n34684));
  jand g17422(.dina(n34684), .dinb(n34683), .dout(n34685));
  jor  g17423(.dina(n34685), .dinb(n34668), .dout(n34686));
  jxor g17424(.dina(n34660), .dinb(n376), .dout(n34687));
  jand g17425(.dina(n34687), .dinb(n34686), .dout(n34688));
  jor  g17426(.dina(n34688), .dinb(n34661), .dout(n34689));
  jxor g17427(.dina(n34655), .dinb(n377), .dout(n34690));
  jand g17428(.dina(n34690), .dinb(n34689), .dout(n34691));
  jor  g17429(.dina(n34691), .dinb(n34656), .dout(n34692));
  jxor g17430(.dina(n34650), .dinb(n378), .dout(n34693));
  jand g17431(.dina(n34693), .dinb(n34692), .dout(n34694));
  jor  g17432(.dina(n34694), .dinb(n34651), .dout(n34695));
  jxor g17433(.dina(n34645), .dinb(n265), .dout(n34696));
  jand g17434(.dina(n34696), .dinb(n34695), .dout(n34697));
  jor  g17435(.dina(n34697), .dinb(n34646), .dout(n34698));
  jxor g17436(.dina(n34640), .dinb(n367), .dout(n34699));
  jand g17437(.dina(n34699), .dinb(n34698), .dout(n34700));
  jor  g17438(.dina(n34700), .dinb(n34641), .dout(n34701));
  jxor g17439(.dina(n34635), .dinb(n368), .dout(n34702));
  jand g17440(.dina(n34702), .dinb(n34701), .dout(n34703));
  jor  g17441(.dina(n34703), .dinb(n34636), .dout(n34704));
  jxor g17442(.dina(n34630), .dinb(n369), .dout(n34705));
  jand g17443(.dina(n34705), .dinb(n34704), .dout(n34706));
  jor  g17444(.dina(n34706), .dinb(n34631), .dout(n34707));
  jxor g17445(.dina(n34625), .dinb(n359), .dout(n34708));
  jand g17446(.dina(n34708), .dinb(n34707), .dout(n34709));
  jor  g17447(.dina(n34709), .dinb(n34626), .dout(n34710));
  jxor g17448(.dina(n34620), .dinb(n363), .dout(n34711));
  jand g17449(.dina(n34711), .dinb(n34710), .dout(n34712));
  jor  g17450(.dina(n34712), .dinb(n34621), .dout(n34713));
  jxor g17451(.dina(n34615), .dinb(n360), .dout(n34714));
  jand g17452(.dina(n34714), .dinb(n34713), .dout(n34715));
  jor  g17453(.dina(n34715), .dinb(n34616), .dout(n34716));
  jxor g17454(.dina(n34610), .dinb(n361), .dout(n34717));
  jand g17455(.dina(n34717), .dinb(n34716), .dout(n34718));
  jor  g17456(.dina(n34718), .dinb(n34611), .dout(n34719));
  jxor g17457(.dina(n34605), .dinb(n364), .dout(n34720));
  jand g17458(.dina(n34720), .dinb(n34719), .dout(n34721));
  jor  g17459(.dina(n34721), .dinb(n34606), .dout(n34722));
  jxor g17460(.dina(n34600), .dinb(n355), .dout(n34723));
  jand g17461(.dina(n34723), .dinb(n34722), .dout(n34724));
  jor  g17462(.dina(n34724), .dinb(n34601), .dout(n34725));
  jxor g17463(.dina(n34595), .dinb(n356), .dout(n34726));
  jand g17464(.dina(n34726), .dinb(n34725), .dout(n34727));
  jor  g17465(.dina(n34727), .dinb(n34596), .dout(n34728));
  jxor g17466(.dina(n34590), .dinb(n266), .dout(n34729));
  jand g17467(.dina(n34729), .dinb(n34728), .dout(n34730));
  jor  g17468(.dina(n34730), .dinb(n34591), .dout(n34731));
  jxor g17469(.dina(n34585), .dinb(n267), .dout(n34732));
  jand g17470(.dina(n34732), .dinb(n34731), .dout(n34733));
  jor  g17471(.dina(n34733), .dinb(n34586), .dout(n34734));
  jxor g17472(.dina(n34580), .dinb(n347), .dout(n34735));
  jand g17473(.dina(n34735), .dinb(n34734), .dout(n34736));
  jor  g17474(.dina(n34736), .dinb(n34581), .dout(n34737));
  jxor g17475(.dina(n34575), .dinb(n348), .dout(n34738));
  jand g17476(.dina(n34738), .dinb(n34737), .dout(n34739));
  jor  g17477(.dina(n34739), .dinb(n34576), .dout(n34740));
  jxor g17478(.dina(n34570), .dinb(n349), .dout(n34741));
  jand g17479(.dina(n34741), .dinb(n34740), .dout(n34742));
  jor  g17480(.dina(n34742), .dinb(n34571), .dout(n34743));
  jxor g17481(.dina(n34565), .dinb(n268), .dout(n34744));
  jand g17482(.dina(n34744), .dinb(n34743), .dout(n34745));
  jor  g17483(.dina(n34745), .dinb(n34566), .dout(n34746));
  jxor g17484(.dina(n34560), .dinb(n274), .dout(n34747));
  jand g17485(.dina(n34747), .dinb(n34746), .dout(n34748));
  jor  g17486(.dina(n34748), .dinb(n34561), .dout(n34749));
  jxor g17487(.dina(n34555), .dinb(n269), .dout(n34750));
  jand g17488(.dina(n34750), .dinb(n34749), .dout(n34751));
  jor  g17489(.dina(n34751), .dinb(n34556), .dout(n34752));
  jxor g17490(.dina(n34550), .dinb(n270), .dout(n34753));
  jand g17491(.dina(n34753), .dinb(n34752), .dout(n34754));
  jor  g17492(.dina(n34754), .dinb(n34551), .dout(n34755));
  jxor g17493(.dina(n34545), .dinb(n271), .dout(n34756));
  jand g17494(.dina(n34756), .dinb(n34755), .dout(n34757));
  jor  g17495(.dina(n34757), .dinb(n34546), .dout(n34758));
  jxor g17496(.dina(n34540), .dinb(n338), .dout(n34759));
  jand g17497(.dina(n34759), .dinb(n34758), .dout(n34760));
  jor  g17498(.dina(n34760), .dinb(n34541), .dout(n34761));
  jxor g17499(.dina(n34535), .dinb(n339), .dout(n34762));
  jand g17500(.dina(n34762), .dinb(n34761), .dout(n34763));
  jor  g17501(.dina(n34763), .dinb(n34536), .dout(n34764));
  jxor g17502(.dina(n34530), .dinb(n340), .dout(n34765));
  jand g17503(.dina(n34765), .dinb(n34764), .dout(n34766));
  jor  g17504(.dina(n34766), .dinb(n34531), .dout(n34767));
  jxor g17505(.dina(n34525), .dinb(n275), .dout(n34768));
  jand g17506(.dina(n34768), .dinb(n34767), .dout(n34769));
  jor  g17507(.dina(n34769), .dinb(n34526), .dout(n34770));
  jxor g17508(.dina(n34520), .dinb(n331), .dout(n34771));
  jand g17509(.dina(n34771), .dinb(n34770), .dout(n34772));
  jor  g17510(.dina(n34772), .dinb(n34521), .dout(n34773));
  jxor g17511(.dina(n34515), .dinb(n332), .dout(n34774));
  jand g17512(.dina(n34774), .dinb(n34773), .dout(n34775));
  jor  g17513(.dina(n34775), .dinb(n34516), .dout(n34776));
  jxor g17514(.dina(n34510), .dinb(n333), .dout(n34777));
  jand g17515(.dina(n34777), .dinb(n34776), .dout(n34778));
  jor  g17516(.dina(n34778), .dinb(n34511), .dout(n34779));
  jxor g17517(.dina(n34505), .dinb(n276), .dout(n34780));
  jand g17518(.dina(n34780), .dinb(n34779), .dout(n34781));
  jor  g17519(.dina(n34781), .dinb(n34506), .dout(n34782));
  jxor g17520(.dina(n34500), .dinb(n324), .dout(n34783));
  jand g17521(.dina(n34783), .dinb(n34782), .dout(n34784));
  jor  g17522(.dina(n34784), .dinb(n34501), .dout(n34785));
  jxor g17523(.dina(n34495), .dinb(n325), .dout(n34786));
  jand g17524(.dina(n34786), .dinb(n34785), .dout(n34787));
  jor  g17525(.dina(n34787), .dinb(n34496), .dout(n34788));
  jxor g17526(.dina(n34490), .dinb(n326), .dout(n34789));
  jand g17527(.dina(n34789), .dinb(n34788), .dout(n34790));
  jor  g17528(.dina(n34790), .dinb(n34491), .dout(n34791));
  jxor g17529(.dina(n34485), .dinb(n277), .dout(n34792));
  jand g17530(.dina(n34792), .dinb(n34791), .dout(n34793));
  jor  g17531(.dina(n34793), .dinb(n34486), .dout(n34794));
  jxor g17532(.dina(n34480), .dinb(n278), .dout(n34795));
  jand g17533(.dina(n34795), .dinb(n34794), .dout(n34796));
  jor  g17534(.dina(n34796), .dinb(n34481), .dout(n34797));
  jxor g17535(.dina(n34475), .dinb(n279), .dout(n34798));
  jand g17536(.dina(n34798), .dinb(n34797), .dout(n34799));
  jor  g17537(.dina(n34799), .dinb(n34476), .dout(n34800));
  jxor g17538(.dina(n34470), .dinb(n280), .dout(n34801));
  jand g17539(.dina(n34801), .dinb(n34800), .dout(n34802));
  jor  g17540(.dina(n34802), .dinb(n34471), .dout(n34803));
  jxor g17541(.dina(n34465), .dinb(n283), .dout(n34804));
  jand g17542(.dina(n34804), .dinb(n34803), .dout(n34805));
  jor  g17543(.dina(n34805), .dinb(n34466), .dout(n34806));
  jxor g17544(.dina(n34460), .dinb(n315), .dout(n34807));
  jand g17545(.dina(n34807), .dinb(n34806), .dout(n34808));
  jor  g17546(.dina(n34808), .dinb(n34461), .dout(n34809));
  jxor g17547(.dina(n34455), .dinb(n316), .dout(n34810));
  jand g17548(.dina(n34810), .dinb(n34809), .dout(n34811));
  jor  g17549(.dina(n34811), .dinb(n34456), .dout(n34812));
  jxor g17550(.dina(n34450), .dinb(n317), .dout(n34813));
  jand g17551(.dina(n34813), .dinb(n34812), .dout(n34814));
  jor  g17552(.dina(n34814), .dinb(n34451), .dout(n34815));
  jxor g17553(.dina(n34445), .dinb(n284), .dout(n34816));
  jand g17554(.dina(n34816), .dinb(n34815), .dout(n34817));
  jor  g17555(.dina(n34817), .dinb(n34446), .dout(n34818));
  jxor g17556(.dina(n34440), .dinb(n285), .dout(n34819));
  jand g17557(.dina(n34819), .dinb(n34818), .dout(n34820));
  jor  g17558(.dina(n34820), .dinb(n34441), .dout(n34821));
  jxor g17559(.dina(n34435), .dinb(n286), .dout(n34822));
  jand g17560(.dina(n34822), .dinb(n34821), .dout(n34823));
  jor  g17561(.dina(n34823), .dinb(n34436), .dout(n34824));
  jxor g17562(.dina(n34430), .dinb(n287), .dout(n34825));
  jand g17563(.dina(n34825), .dinb(n34824), .dout(n34826));
  jor  g17564(.dina(n34826), .dinb(n34431), .dout(n34827));
  jxor g17565(.dina(n34425), .dinb(n288), .dout(n34828));
  jand g17566(.dina(n34828), .dinb(n34827), .dout(n34829));
  jor  g17567(.dina(n34829), .dinb(n34426), .dout(n34830));
  jxor g17568(.dina(n34420), .dinb(n289), .dout(n34831));
  jand g17569(.dina(n34831), .dinb(n34830), .dout(n34832));
  jor  g17570(.dina(n34832), .dinb(n34421), .dout(n34833));
  jxor g17571(.dina(n34415), .dinb(n290), .dout(n34834));
  jand g17572(.dina(n34834), .dinb(n34833), .dout(n34835));
  jor  g17573(.dina(n34835), .dinb(n34416), .dout(n34836));
  jxor g17574(.dina(n34410), .dinb(n291), .dout(n34837));
  jand g17575(.dina(n34837), .dinb(n34836), .dout(n34838));
  jor  g17576(.dina(n34838), .dinb(n34411), .dout(n34839));
  jxor g17577(.dina(n34399), .dinb(n292), .dout(n34840));
  jand g17578(.dina(n34840), .dinb(n34839), .dout(n34841));
  jor  g17579(.dina(n34841), .dinb(n34406), .dout(n34842));
  jand g17580(.dina(n34842), .dinb(n34405), .dout(n34843));
  jor  g17581(.dina(n34843), .dinb(n34404), .dout(n34844));
  jand g17582(.dina(n34844), .dinb(n304), .dout(n34845));
  jor  g17583(.dina(n34845), .dinb(n34399), .dout(n34846));
  jnot g17584(.din(n34845), .dout(n34847));
  jxor g17585(.dina(n34840), .dinb(n34839), .dout(n34848));
  jor  g17586(.dina(n34848), .dinb(n34847), .dout(n34849));
  jand g17587(.dina(n34849), .dinb(n34846), .dout(n34850));
  jand g17588(.dina(n34847), .dinb(n34403), .dout(n34851));
  jand g17589(.dina(n34842), .dinb(n34404), .dout(n34852));
  jor  g17590(.dina(n34852), .dinb(n34851), .dout(n34853));
  jand g17591(.dina(n34853), .dinb(n294), .dout(n34854));
  jnot g17592(.din(n34853), .dout(n34855));
  jand g17593(.dina(n34855), .dinb(b57 ), .dout(n34856));
  jnot g17594(.din(n34856), .dout(n34857));
  jand g17595(.dina(n34850), .dinb(n293), .dout(n34858));
  jor  g17596(.dina(n34845), .dinb(n34410), .dout(n34859));
  jxor g17597(.dina(n34837), .dinb(n34836), .dout(n34860));
  jor  g17598(.dina(n34860), .dinb(n34847), .dout(n34861));
  jand g17599(.dina(n34861), .dinb(n34859), .dout(n34862));
  jand g17600(.dina(n34862), .dinb(n292), .dout(n34863));
  jor  g17601(.dina(n34845), .dinb(n34415), .dout(n34864));
  jxor g17602(.dina(n34834), .dinb(n34833), .dout(n34865));
  jor  g17603(.dina(n34865), .dinb(n34847), .dout(n34866));
  jand g17604(.dina(n34866), .dinb(n34864), .dout(n34867));
  jand g17605(.dina(n34867), .dinb(n291), .dout(n34868));
  jor  g17606(.dina(n34845), .dinb(n34420), .dout(n34869));
  jxor g17607(.dina(n34831), .dinb(n34830), .dout(n34870));
  jor  g17608(.dina(n34870), .dinb(n34847), .dout(n34871));
  jand g17609(.dina(n34871), .dinb(n34869), .dout(n34872));
  jand g17610(.dina(n34872), .dinb(n290), .dout(n34873));
  jor  g17611(.dina(n34845), .dinb(n34425), .dout(n34874));
  jxor g17612(.dina(n34828), .dinb(n34827), .dout(n34875));
  jor  g17613(.dina(n34875), .dinb(n34847), .dout(n34876));
  jand g17614(.dina(n34876), .dinb(n34874), .dout(n34877));
  jand g17615(.dina(n34877), .dinb(n289), .dout(n34878));
  jor  g17616(.dina(n34845), .dinb(n34430), .dout(n34879));
  jxor g17617(.dina(n34825), .dinb(n34824), .dout(n34880));
  jor  g17618(.dina(n34880), .dinb(n34847), .dout(n34881));
  jand g17619(.dina(n34881), .dinb(n34879), .dout(n34882));
  jand g17620(.dina(n34882), .dinb(n288), .dout(n34883));
  jor  g17621(.dina(n34845), .dinb(n34435), .dout(n34884));
  jxor g17622(.dina(n34822), .dinb(n34821), .dout(n34885));
  jor  g17623(.dina(n34885), .dinb(n34847), .dout(n34886));
  jand g17624(.dina(n34886), .dinb(n34884), .dout(n34887));
  jand g17625(.dina(n34887), .dinb(n287), .dout(n34888));
  jor  g17626(.dina(n34845), .dinb(n34440), .dout(n34889));
  jxor g17627(.dina(n34819), .dinb(n34818), .dout(n34890));
  jor  g17628(.dina(n34890), .dinb(n34847), .dout(n34891));
  jand g17629(.dina(n34891), .dinb(n34889), .dout(n34892));
  jand g17630(.dina(n34892), .dinb(n286), .dout(n34893));
  jor  g17631(.dina(n34845), .dinb(n34445), .dout(n34894));
  jxor g17632(.dina(n34816), .dinb(n34815), .dout(n34895));
  jor  g17633(.dina(n34895), .dinb(n34847), .dout(n34896));
  jand g17634(.dina(n34896), .dinb(n34894), .dout(n34897));
  jand g17635(.dina(n34897), .dinb(n285), .dout(n34898));
  jor  g17636(.dina(n34845), .dinb(n34450), .dout(n34899));
  jxor g17637(.dina(n34813), .dinb(n34812), .dout(n34900));
  jor  g17638(.dina(n34900), .dinb(n34847), .dout(n34901));
  jand g17639(.dina(n34901), .dinb(n34899), .dout(n34902));
  jand g17640(.dina(n34902), .dinb(n284), .dout(n34903));
  jor  g17641(.dina(n34845), .dinb(n34455), .dout(n34904));
  jxor g17642(.dina(n34810), .dinb(n34809), .dout(n34905));
  jor  g17643(.dina(n34905), .dinb(n34847), .dout(n34906));
  jand g17644(.dina(n34906), .dinb(n34904), .dout(n34907));
  jand g17645(.dina(n34907), .dinb(n317), .dout(n34908));
  jor  g17646(.dina(n34845), .dinb(n34460), .dout(n34909));
  jxor g17647(.dina(n34807), .dinb(n34806), .dout(n34910));
  jor  g17648(.dina(n34910), .dinb(n34847), .dout(n34911));
  jand g17649(.dina(n34911), .dinb(n34909), .dout(n34912));
  jand g17650(.dina(n34912), .dinb(n316), .dout(n34913));
  jor  g17651(.dina(n34845), .dinb(n34465), .dout(n34914));
  jxor g17652(.dina(n34804), .dinb(n34803), .dout(n34915));
  jor  g17653(.dina(n34915), .dinb(n34847), .dout(n34916));
  jand g17654(.dina(n34916), .dinb(n34914), .dout(n34917));
  jand g17655(.dina(n34917), .dinb(n315), .dout(n34918));
  jor  g17656(.dina(n34845), .dinb(n34470), .dout(n34919));
  jxor g17657(.dina(n34801), .dinb(n34800), .dout(n34920));
  jor  g17658(.dina(n34920), .dinb(n34847), .dout(n34921));
  jand g17659(.dina(n34921), .dinb(n34919), .dout(n34922));
  jand g17660(.dina(n34922), .dinb(n283), .dout(n34923));
  jor  g17661(.dina(n34845), .dinb(n34475), .dout(n34924));
  jxor g17662(.dina(n34798), .dinb(n34797), .dout(n34925));
  jor  g17663(.dina(n34925), .dinb(n34847), .dout(n34926));
  jand g17664(.dina(n34926), .dinb(n34924), .dout(n34927));
  jand g17665(.dina(n34927), .dinb(n280), .dout(n34928));
  jor  g17666(.dina(n34845), .dinb(n34480), .dout(n34929));
  jxor g17667(.dina(n34795), .dinb(n34794), .dout(n34930));
  jor  g17668(.dina(n34930), .dinb(n34847), .dout(n34931));
  jand g17669(.dina(n34931), .dinb(n34929), .dout(n34932));
  jand g17670(.dina(n34932), .dinb(n279), .dout(n34933));
  jor  g17671(.dina(n34845), .dinb(n34485), .dout(n34934));
  jxor g17672(.dina(n34792), .dinb(n34791), .dout(n34935));
  jor  g17673(.dina(n34935), .dinb(n34847), .dout(n34936));
  jand g17674(.dina(n34936), .dinb(n34934), .dout(n34937));
  jand g17675(.dina(n34937), .dinb(n278), .dout(n34938));
  jor  g17676(.dina(n34845), .dinb(n34490), .dout(n34939));
  jxor g17677(.dina(n34789), .dinb(n34788), .dout(n34940));
  jor  g17678(.dina(n34940), .dinb(n34847), .dout(n34941));
  jand g17679(.dina(n34941), .dinb(n34939), .dout(n34942));
  jand g17680(.dina(n34942), .dinb(n277), .dout(n34943));
  jor  g17681(.dina(n34845), .dinb(n34495), .dout(n34944));
  jxor g17682(.dina(n34786), .dinb(n34785), .dout(n34945));
  jor  g17683(.dina(n34945), .dinb(n34847), .dout(n34946));
  jand g17684(.dina(n34946), .dinb(n34944), .dout(n34947));
  jand g17685(.dina(n34947), .dinb(n326), .dout(n34948));
  jor  g17686(.dina(n34845), .dinb(n34500), .dout(n34949));
  jxor g17687(.dina(n34783), .dinb(n34782), .dout(n34950));
  jor  g17688(.dina(n34950), .dinb(n34847), .dout(n34951));
  jand g17689(.dina(n34951), .dinb(n34949), .dout(n34952));
  jand g17690(.dina(n34952), .dinb(n325), .dout(n34953));
  jor  g17691(.dina(n34845), .dinb(n34505), .dout(n34954));
  jxor g17692(.dina(n34780), .dinb(n34779), .dout(n34955));
  jor  g17693(.dina(n34955), .dinb(n34847), .dout(n34956));
  jand g17694(.dina(n34956), .dinb(n34954), .dout(n34957));
  jand g17695(.dina(n34957), .dinb(n324), .dout(n34958));
  jor  g17696(.dina(n34845), .dinb(n34510), .dout(n34959));
  jxor g17697(.dina(n34777), .dinb(n34776), .dout(n34960));
  jor  g17698(.dina(n34960), .dinb(n34847), .dout(n34961));
  jand g17699(.dina(n34961), .dinb(n34959), .dout(n34962));
  jand g17700(.dina(n34962), .dinb(n276), .dout(n34963));
  jor  g17701(.dina(n34845), .dinb(n34515), .dout(n34964));
  jxor g17702(.dina(n34774), .dinb(n34773), .dout(n34965));
  jor  g17703(.dina(n34965), .dinb(n34847), .dout(n34966));
  jand g17704(.dina(n34966), .dinb(n34964), .dout(n34967));
  jand g17705(.dina(n34967), .dinb(n333), .dout(n34968));
  jor  g17706(.dina(n34845), .dinb(n34520), .dout(n34969));
  jxor g17707(.dina(n34771), .dinb(n34770), .dout(n34970));
  jor  g17708(.dina(n34970), .dinb(n34847), .dout(n34971));
  jand g17709(.dina(n34971), .dinb(n34969), .dout(n34972));
  jand g17710(.dina(n34972), .dinb(n332), .dout(n34973));
  jor  g17711(.dina(n34845), .dinb(n34525), .dout(n34974));
  jxor g17712(.dina(n34768), .dinb(n34767), .dout(n34975));
  jor  g17713(.dina(n34975), .dinb(n34847), .dout(n34976));
  jand g17714(.dina(n34976), .dinb(n34974), .dout(n34977));
  jand g17715(.dina(n34977), .dinb(n331), .dout(n34978));
  jor  g17716(.dina(n34845), .dinb(n34530), .dout(n34979));
  jxor g17717(.dina(n34765), .dinb(n34764), .dout(n34980));
  jor  g17718(.dina(n34980), .dinb(n34847), .dout(n34981));
  jand g17719(.dina(n34981), .dinb(n34979), .dout(n34982));
  jand g17720(.dina(n34982), .dinb(n275), .dout(n34983));
  jor  g17721(.dina(n34845), .dinb(n34535), .dout(n34984));
  jxor g17722(.dina(n34762), .dinb(n34761), .dout(n34985));
  jor  g17723(.dina(n34985), .dinb(n34847), .dout(n34986));
  jand g17724(.dina(n34986), .dinb(n34984), .dout(n34987));
  jand g17725(.dina(n34987), .dinb(n340), .dout(n34988));
  jor  g17726(.dina(n34845), .dinb(n34540), .dout(n34989));
  jxor g17727(.dina(n34759), .dinb(n34758), .dout(n34990));
  jor  g17728(.dina(n34990), .dinb(n34847), .dout(n34991));
  jand g17729(.dina(n34991), .dinb(n34989), .dout(n34992));
  jand g17730(.dina(n34992), .dinb(n339), .dout(n34993));
  jor  g17731(.dina(n34845), .dinb(n34545), .dout(n34994));
  jxor g17732(.dina(n34756), .dinb(n34755), .dout(n34995));
  jor  g17733(.dina(n34995), .dinb(n34847), .dout(n34996));
  jand g17734(.dina(n34996), .dinb(n34994), .dout(n34997));
  jand g17735(.dina(n34997), .dinb(n338), .dout(n34998));
  jor  g17736(.dina(n34845), .dinb(n34550), .dout(n34999));
  jxor g17737(.dina(n34753), .dinb(n34752), .dout(n35000));
  jor  g17738(.dina(n35000), .dinb(n34847), .dout(n35001));
  jand g17739(.dina(n35001), .dinb(n34999), .dout(n35002));
  jand g17740(.dina(n35002), .dinb(n271), .dout(n35003));
  jor  g17741(.dina(n34845), .dinb(n34555), .dout(n35004));
  jxor g17742(.dina(n34750), .dinb(n34749), .dout(n35005));
  jor  g17743(.dina(n35005), .dinb(n34847), .dout(n35006));
  jand g17744(.dina(n35006), .dinb(n35004), .dout(n35007));
  jand g17745(.dina(n35007), .dinb(n270), .dout(n35008));
  jor  g17746(.dina(n34845), .dinb(n34560), .dout(n35009));
  jxor g17747(.dina(n34747), .dinb(n34746), .dout(n35010));
  jor  g17748(.dina(n35010), .dinb(n34847), .dout(n35011));
  jand g17749(.dina(n35011), .dinb(n35009), .dout(n35012));
  jand g17750(.dina(n35012), .dinb(n269), .dout(n35013));
  jor  g17751(.dina(n34845), .dinb(n34565), .dout(n35014));
  jxor g17752(.dina(n34744), .dinb(n34743), .dout(n35015));
  jor  g17753(.dina(n35015), .dinb(n34847), .dout(n35016));
  jand g17754(.dina(n35016), .dinb(n35014), .dout(n35017));
  jand g17755(.dina(n35017), .dinb(n274), .dout(n35018));
  jor  g17756(.dina(n34845), .dinb(n34570), .dout(n35019));
  jxor g17757(.dina(n34741), .dinb(n34740), .dout(n35020));
  jor  g17758(.dina(n35020), .dinb(n34847), .dout(n35021));
  jand g17759(.dina(n35021), .dinb(n35019), .dout(n35022));
  jand g17760(.dina(n35022), .dinb(n268), .dout(n35023));
  jor  g17761(.dina(n34845), .dinb(n34575), .dout(n35024));
  jxor g17762(.dina(n34738), .dinb(n34737), .dout(n35025));
  jor  g17763(.dina(n35025), .dinb(n34847), .dout(n35026));
  jand g17764(.dina(n35026), .dinb(n35024), .dout(n35027));
  jand g17765(.dina(n35027), .dinb(n349), .dout(n35028));
  jor  g17766(.dina(n34845), .dinb(n34580), .dout(n35029));
  jxor g17767(.dina(n34735), .dinb(n34734), .dout(n35030));
  jor  g17768(.dina(n35030), .dinb(n34847), .dout(n35031));
  jand g17769(.dina(n35031), .dinb(n35029), .dout(n35032));
  jand g17770(.dina(n35032), .dinb(n348), .dout(n35033));
  jor  g17771(.dina(n34845), .dinb(n34585), .dout(n35034));
  jxor g17772(.dina(n34732), .dinb(n34731), .dout(n35035));
  jor  g17773(.dina(n35035), .dinb(n34847), .dout(n35036));
  jand g17774(.dina(n35036), .dinb(n35034), .dout(n35037));
  jand g17775(.dina(n35037), .dinb(n347), .dout(n35038));
  jor  g17776(.dina(n34845), .dinb(n34590), .dout(n35039));
  jxor g17777(.dina(n34729), .dinb(n34728), .dout(n35040));
  jor  g17778(.dina(n35040), .dinb(n34847), .dout(n35041));
  jand g17779(.dina(n35041), .dinb(n35039), .dout(n35042));
  jand g17780(.dina(n35042), .dinb(n267), .dout(n35043));
  jor  g17781(.dina(n34845), .dinb(n34595), .dout(n35044));
  jxor g17782(.dina(n34726), .dinb(n34725), .dout(n35045));
  jor  g17783(.dina(n35045), .dinb(n34847), .dout(n35046));
  jand g17784(.dina(n35046), .dinb(n35044), .dout(n35047));
  jand g17785(.dina(n35047), .dinb(n266), .dout(n35048));
  jor  g17786(.dina(n34845), .dinb(n34600), .dout(n35049));
  jxor g17787(.dina(n34723), .dinb(n34722), .dout(n35050));
  jor  g17788(.dina(n35050), .dinb(n34847), .dout(n35051));
  jand g17789(.dina(n35051), .dinb(n35049), .dout(n35052));
  jand g17790(.dina(n35052), .dinb(n356), .dout(n35053));
  jor  g17791(.dina(n34845), .dinb(n34605), .dout(n35054));
  jxor g17792(.dina(n34720), .dinb(n34719), .dout(n35055));
  jor  g17793(.dina(n35055), .dinb(n34847), .dout(n35056));
  jand g17794(.dina(n35056), .dinb(n35054), .dout(n35057));
  jand g17795(.dina(n35057), .dinb(n355), .dout(n35058));
  jor  g17796(.dina(n34845), .dinb(n34610), .dout(n35059));
  jxor g17797(.dina(n34717), .dinb(n34716), .dout(n35060));
  jor  g17798(.dina(n35060), .dinb(n34847), .dout(n35061));
  jand g17799(.dina(n35061), .dinb(n35059), .dout(n35062));
  jand g17800(.dina(n35062), .dinb(n364), .dout(n35063));
  jor  g17801(.dina(n34845), .dinb(n34615), .dout(n35064));
  jxor g17802(.dina(n34714), .dinb(n34713), .dout(n35065));
  jor  g17803(.dina(n35065), .dinb(n34847), .dout(n35066));
  jand g17804(.dina(n35066), .dinb(n35064), .dout(n35067));
  jand g17805(.dina(n35067), .dinb(n361), .dout(n35068));
  jor  g17806(.dina(n34845), .dinb(n34620), .dout(n35069));
  jxor g17807(.dina(n34711), .dinb(n34710), .dout(n35070));
  jor  g17808(.dina(n35070), .dinb(n34847), .dout(n35071));
  jand g17809(.dina(n35071), .dinb(n35069), .dout(n35072));
  jand g17810(.dina(n35072), .dinb(n360), .dout(n35073));
  jor  g17811(.dina(n34845), .dinb(n34625), .dout(n35074));
  jxor g17812(.dina(n34708), .dinb(n34707), .dout(n35075));
  jor  g17813(.dina(n35075), .dinb(n34847), .dout(n35076));
  jand g17814(.dina(n35076), .dinb(n35074), .dout(n35077));
  jand g17815(.dina(n35077), .dinb(n363), .dout(n35078));
  jor  g17816(.dina(n34845), .dinb(n34630), .dout(n35079));
  jxor g17817(.dina(n34705), .dinb(n34704), .dout(n35080));
  jor  g17818(.dina(n35080), .dinb(n34847), .dout(n35081));
  jand g17819(.dina(n35081), .dinb(n35079), .dout(n35082));
  jand g17820(.dina(n35082), .dinb(n359), .dout(n35083));
  jor  g17821(.dina(n34845), .dinb(n34635), .dout(n35084));
  jxor g17822(.dina(n34702), .dinb(n34701), .dout(n35085));
  jor  g17823(.dina(n35085), .dinb(n34847), .dout(n35086));
  jand g17824(.dina(n35086), .dinb(n35084), .dout(n35087));
  jand g17825(.dina(n35087), .dinb(n369), .dout(n35088));
  jor  g17826(.dina(n34845), .dinb(n34640), .dout(n35089));
  jxor g17827(.dina(n34699), .dinb(n34698), .dout(n35090));
  jor  g17828(.dina(n35090), .dinb(n34847), .dout(n35091));
  jand g17829(.dina(n35091), .dinb(n35089), .dout(n35092));
  jand g17830(.dina(n35092), .dinb(n368), .dout(n35093));
  jor  g17831(.dina(n34845), .dinb(n34645), .dout(n35094));
  jxor g17832(.dina(n34696), .dinb(n34695), .dout(n35095));
  jor  g17833(.dina(n35095), .dinb(n34847), .dout(n35096));
  jand g17834(.dina(n35096), .dinb(n35094), .dout(n35097));
  jand g17835(.dina(n35097), .dinb(n367), .dout(n35098));
  jor  g17836(.dina(n34845), .dinb(n34650), .dout(n35099));
  jxor g17837(.dina(n34693), .dinb(n34692), .dout(n35100));
  jor  g17838(.dina(n35100), .dinb(n34847), .dout(n35101));
  jand g17839(.dina(n35101), .dinb(n35099), .dout(n35102));
  jand g17840(.dina(n35102), .dinb(n265), .dout(n35103));
  jor  g17841(.dina(n34845), .dinb(n34655), .dout(n35104));
  jxor g17842(.dina(n34690), .dinb(n34689), .dout(n35105));
  jor  g17843(.dina(n35105), .dinb(n34847), .dout(n35106));
  jand g17844(.dina(n35106), .dinb(n35104), .dout(n35107));
  jand g17845(.dina(n35107), .dinb(n378), .dout(n35108));
  jor  g17846(.dina(n34845), .dinb(n34660), .dout(n35109));
  jxor g17847(.dina(n34687), .dinb(n34686), .dout(n35110));
  jor  g17848(.dina(n35110), .dinb(n34847), .dout(n35111));
  jand g17849(.dina(n35111), .dinb(n35109), .dout(n35112));
  jand g17850(.dina(n35112), .dinb(n377), .dout(n35113));
  jand g17851(.dina(n34847), .dinb(n34666), .dout(n35114));
  jnot g17852(.din(n35114), .dout(n35115));
  jxor g17853(.dina(n34684), .dinb(n34683), .dout(n35116));
  jor  g17854(.dina(n35116), .dinb(n34847), .dout(n35117));
  jand g17855(.dina(n35117), .dinb(n35115), .dout(n35118));
  jand g17856(.dina(n35118), .dinb(n376), .dout(n35119));
  jor  g17857(.dina(n34845), .dinb(n34672), .dout(n35120));
  jxor g17858(.dina(n34681), .dinb(n34680), .dout(n35121));
  jor  g17859(.dina(n35121), .dinb(n34847), .dout(n35122));
  jand g17860(.dina(n35122), .dinb(n35120), .dout(n35123));
  jand g17861(.dina(n35123), .dinb(n264), .dout(n35124));
  jxor g17862(.dina(n34678), .dinb(n14205), .dout(n35125));
  jand g17863(.dina(n35125), .dinb(n34845), .dout(n35126));
  jnot g17864(.din(n35126), .dout(n35127));
  jor  g17865(.dina(n34845), .dinb(n34677), .dout(n35128));
  jand g17866(.dina(n35128), .dinb(n35127), .dout(n35129));
  jnot g17867(.din(n35129), .dout(n35130));
  jand g17868(.dina(n35130), .dinb(n386), .dout(n35131));
  jand g17869(.dina(n34845), .dinb(b0 ), .dout(n35132));
  jxor g17870(.dina(n35132), .dinb(a7 ), .dout(n35133));
  jand g17871(.dina(n35133), .dinb(n259), .dout(n35134));
  jxor g17872(.dina(n35132), .dinb(n14203), .dout(n35135));
  jxor g17873(.dina(n35135), .dinb(b1 ), .dout(n35136));
  jand g17874(.dina(n35136), .dinb(n14663), .dout(n35137));
  jor  g17875(.dina(n35137), .dinb(n35134), .dout(n35138));
  jxor g17876(.dina(n35129), .dinb(b2 ), .dout(n35139));
  jand g17877(.dina(n35139), .dinb(n35138), .dout(n35140));
  jor  g17878(.dina(n35140), .dinb(n35131), .dout(n35141));
  jxor g17879(.dina(n35123), .dinb(n264), .dout(n35142));
  jand g17880(.dina(n35142), .dinb(n35141), .dout(n35143));
  jor  g17881(.dina(n35143), .dinb(n35124), .dout(n35144));
  jxor g17882(.dina(n35118), .dinb(n376), .dout(n35145));
  jand g17883(.dina(n35145), .dinb(n35144), .dout(n35146));
  jor  g17884(.dina(n35146), .dinb(n35119), .dout(n35147));
  jxor g17885(.dina(n35112), .dinb(n377), .dout(n35148));
  jand g17886(.dina(n35148), .dinb(n35147), .dout(n35149));
  jor  g17887(.dina(n35149), .dinb(n35113), .dout(n35150));
  jxor g17888(.dina(n35107), .dinb(n378), .dout(n35151));
  jand g17889(.dina(n35151), .dinb(n35150), .dout(n35152));
  jor  g17890(.dina(n35152), .dinb(n35108), .dout(n35153));
  jxor g17891(.dina(n35102), .dinb(n265), .dout(n35154));
  jand g17892(.dina(n35154), .dinb(n35153), .dout(n35155));
  jor  g17893(.dina(n35155), .dinb(n35103), .dout(n35156));
  jxor g17894(.dina(n35097), .dinb(n367), .dout(n35157));
  jand g17895(.dina(n35157), .dinb(n35156), .dout(n35158));
  jor  g17896(.dina(n35158), .dinb(n35098), .dout(n35159));
  jxor g17897(.dina(n35092), .dinb(n368), .dout(n35160));
  jand g17898(.dina(n35160), .dinb(n35159), .dout(n35161));
  jor  g17899(.dina(n35161), .dinb(n35093), .dout(n35162));
  jxor g17900(.dina(n35087), .dinb(n369), .dout(n35163));
  jand g17901(.dina(n35163), .dinb(n35162), .dout(n35164));
  jor  g17902(.dina(n35164), .dinb(n35088), .dout(n35165));
  jxor g17903(.dina(n35082), .dinb(n359), .dout(n35166));
  jand g17904(.dina(n35166), .dinb(n35165), .dout(n35167));
  jor  g17905(.dina(n35167), .dinb(n35083), .dout(n35168));
  jxor g17906(.dina(n35077), .dinb(n363), .dout(n35169));
  jand g17907(.dina(n35169), .dinb(n35168), .dout(n35170));
  jor  g17908(.dina(n35170), .dinb(n35078), .dout(n35171));
  jxor g17909(.dina(n35072), .dinb(n360), .dout(n35172));
  jand g17910(.dina(n35172), .dinb(n35171), .dout(n35173));
  jor  g17911(.dina(n35173), .dinb(n35073), .dout(n35174));
  jxor g17912(.dina(n35067), .dinb(n361), .dout(n35175));
  jand g17913(.dina(n35175), .dinb(n35174), .dout(n35176));
  jor  g17914(.dina(n35176), .dinb(n35068), .dout(n35177));
  jxor g17915(.dina(n35062), .dinb(n364), .dout(n35178));
  jand g17916(.dina(n35178), .dinb(n35177), .dout(n35179));
  jor  g17917(.dina(n35179), .dinb(n35063), .dout(n35180));
  jxor g17918(.dina(n35057), .dinb(n355), .dout(n35181));
  jand g17919(.dina(n35181), .dinb(n35180), .dout(n35182));
  jor  g17920(.dina(n35182), .dinb(n35058), .dout(n35183));
  jxor g17921(.dina(n35052), .dinb(n356), .dout(n35184));
  jand g17922(.dina(n35184), .dinb(n35183), .dout(n35185));
  jor  g17923(.dina(n35185), .dinb(n35053), .dout(n35186));
  jxor g17924(.dina(n35047), .dinb(n266), .dout(n35187));
  jand g17925(.dina(n35187), .dinb(n35186), .dout(n35188));
  jor  g17926(.dina(n35188), .dinb(n35048), .dout(n35189));
  jxor g17927(.dina(n35042), .dinb(n267), .dout(n35190));
  jand g17928(.dina(n35190), .dinb(n35189), .dout(n35191));
  jor  g17929(.dina(n35191), .dinb(n35043), .dout(n35192));
  jxor g17930(.dina(n35037), .dinb(n347), .dout(n35193));
  jand g17931(.dina(n35193), .dinb(n35192), .dout(n35194));
  jor  g17932(.dina(n35194), .dinb(n35038), .dout(n35195));
  jxor g17933(.dina(n35032), .dinb(n348), .dout(n35196));
  jand g17934(.dina(n35196), .dinb(n35195), .dout(n35197));
  jor  g17935(.dina(n35197), .dinb(n35033), .dout(n35198));
  jxor g17936(.dina(n35027), .dinb(n349), .dout(n35199));
  jand g17937(.dina(n35199), .dinb(n35198), .dout(n35200));
  jor  g17938(.dina(n35200), .dinb(n35028), .dout(n35201));
  jxor g17939(.dina(n35022), .dinb(n268), .dout(n35202));
  jand g17940(.dina(n35202), .dinb(n35201), .dout(n35203));
  jor  g17941(.dina(n35203), .dinb(n35023), .dout(n35204));
  jxor g17942(.dina(n35017), .dinb(n274), .dout(n35205));
  jand g17943(.dina(n35205), .dinb(n35204), .dout(n35206));
  jor  g17944(.dina(n35206), .dinb(n35018), .dout(n35207));
  jxor g17945(.dina(n35012), .dinb(n269), .dout(n35208));
  jand g17946(.dina(n35208), .dinb(n35207), .dout(n35209));
  jor  g17947(.dina(n35209), .dinb(n35013), .dout(n35210));
  jxor g17948(.dina(n35007), .dinb(n270), .dout(n35211));
  jand g17949(.dina(n35211), .dinb(n35210), .dout(n35212));
  jor  g17950(.dina(n35212), .dinb(n35008), .dout(n35213));
  jxor g17951(.dina(n35002), .dinb(n271), .dout(n35214));
  jand g17952(.dina(n35214), .dinb(n35213), .dout(n35215));
  jor  g17953(.dina(n35215), .dinb(n35003), .dout(n35216));
  jxor g17954(.dina(n34997), .dinb(n338), .dout(n35217));
  jand g17955(.dina(n35217), .dinb(n35216), .dout(n35218));
  jor  g17956(.dina(n35218), .dinb(n34998), .dout(n35219));
  jxor g17957(.dina(n34992), .dinb(n339), .dout(n35220));
  jand g17958(.dina(n35220), .dinb(n35219), .dout(n35221));
  jor  g17959(.dina(n35221), .dinb(n34993), .dout(n35222));
  jxor g17960(.dina(n34987), .dinb(n340), .dout(n35223));
  jand g17961(.dina(n35223), .dinb(n35222), .dout(n35224));
  jor  g17962(.dina(n35224), .dinb(n34988), .dout(n35225));
  jxor g17963(.dina(n34982), .dinb(n275), .dout(n35226));
  jand g17964(.dina(n35226), .dinb(n35225), .dout(n35227));
  jor  g17965(.dina(n35227), .dinb(n34983), .dout(n35228));
  jxor g17966(.dina(n34977), .dinb(n331), .dout(n35229));
  jand g17967(.dina(n35229), .dinb(n35228), .dout(n35230));
  jor  g17968(.dina(n35230), .dinb(n34978), .dout(n35231));
  jxor g17969(.dina(n34972), .dinb(n332), .dout(n35232));
  jand g17970(.dina(n35232), .dinb(n35231), .dout(n35233));
  jor  g17971(.dina(n35233), .dinb(n34973), .dout(n35234));
  jxor g17972(.dina(n34967), .dinb(n333), .dout(n35235));
  jand g17973(.dina(n35235), .dinb(n35234), .dout(n35236));
  jor  g17974(.dina(n35236), .dinb(n34968), .dout(n35237));
  jxor g17975(.dina(n34962), .dinb(n276), .dout(n35238));
  jand g17976(.dina(n35238), .dinb(n35237), .dout(n35239));
  jor  g17977(.dina(n35239), .dinb(n34963), .dout(n35240));
  jxor g17978(.dina(n34957), .dinb(n324), .dout(n35241));
  jand g17979(.dina(n35241), .dinb(n35240), .dout(n35242));
  jor  g17980(.dina(n35242), .dinb(n34958), .dout(n35243));
  jxor g17981(.dina(n34952), .dinb(n325), .dout(n35244));
  jand g17982(.dina(n35244), .dinb(n35243), .dout(n35245));
  jor  g17983(.dina(n35245), .dinb(n34953), .dout(n35246));
  jxor g17984(.dina(n34947), .dinb(n326), .dout(n35247));
  jand g17985(.dina(n35247), .dinb(n35246), .dout(n35248));
  jor  g17986(.dina(n35248), .dinb(n34948), .dout(n35249));
  jxor g17987(.dina(n34942), .dinb(n277), .dout(n35250));
  jand g17988(.dina(n35250), .dinb(n35249), .dout(n35251));
  jor  g17989(.dina(n35251), .dinb(n34943), .dout(n35252));
  jxor g17990(.dina(n34937), .dinb(n278), .dout(n35253));
  jand g17991(.dina(n35253), .dinb(n35252), .dout(n35254));
  jor  g17992(.dina(n35254), .dinb(n34938), .dout(n35255));
  jxor g17993(.dina(n34932), .dinb(n279), .dout(n35256));
  jand g17994(.dina(n35256), .dinb(n35255), .dout(n35257));
  jor  g17995(.dina(n35257), .dinb(n34933), .dout(n35258));
  jxor g17996(.dina(n34927), .dinb(n280), .dout(n35259));
  jand g17997(.dina(n35259), .dinb(n35258), .dout(n35260));
  jor  g17998(.dina(n35260), .dinb(n34928), .dout(n35261));
  jxor g17999(.dina(n34922), .dinb(n283), .dout(n35262));
  jand g18000(.dina(n35262), .dinb(n35261), .dout(n35263));
  jor  g18001(.dina(n35263), .dinb(n34923), .dout(n35264));
  jxor g18002(.dina(n34917), .dinb(n315), .dout(n35265));
  jand g18003(.dina(n35265), .dinb(n35264), .dout(n35266));
  jor  g18004(.dina(n35266), .dinb(n34918), .dout(n35267));
  jxor g18005(.dina(n34912), .dinb(n316), .dout(n35268));
  jand g18006(.dina(n35268), .dinb(n35267), .dout(n35269));
  jor  g18007(.dina(n35269), .dinb(n34913), .dout(n35270));
  jxor g18008(.dina(n34907), .dinb(n317), .dout(n35271));
  jand g18009(.dina(n35271), .dinb(n35270), .dout(n35272));
  jor  g18010(.dina(n35272), .dinb(n34908), .dout(n35273));
  jxor g18011(.dina(n34902), .dinb(n284), .dout(n35274));
  jand g18012(.dina(n35274), .dinb(n35273), .dout(n35275));
  jor  g18013(.dina(n35275), .dinb(n34903), .dout(n35276));
  jxor g18014(.dina(n34897), .dinb(n285), .dout(n35277));
  jand g18015(.dina(n35277), .dinb(n35276), .dout(n35278));
  jor  g18016(.dina(n35278), .dinb(n34898), .dout(n35279));
  jxor g18017(.dina(n34892), .dinb(n286), .dout(n35280));
  jand g18018(.dina(n35280), .dinb(n35279), .dout(n35281));
  jor  g18019(.dina(n35281), .dinb(n34893), .dout(n35282));
  jxor g18020(.dina(n34887), .dinb(n287), .dout(n35283));
  jand g18021(.dina(n35283), .dinb(n35282), .dout(n35284));
  jor  g18022(.dina(n35284), .dinb(n34888), .dout(n35285));
  jxor g18023(.dina(n34882), .dinb(n288), .dout(n35286));
  jand g18024(.dina(n35286), .dinb(n35285), .dout(n35287));
  jor  g18025(.dina(n35287), .dinb(n34883), .dout(n35288));
  jxor g18026(.dina(n34877), .dinb(n289), .dout(n35289));
  jand g18027(.dina(n35289), .dinb(n35288), .dout(n35290));
  jor  g18028(.dina(n35290), .dinb(n34878), .dout(n35291));
  jxor g18029(.dina(n34872), .dinb(n290), .dout(n35292));
  jand g18030(.dina(n35292), .dinb(n35291), .dout(n35293));
  jor  g18031(.dina(n35293), .dinb(n34873), .dout(n35294));
  jxor g18032(.dina(n34867), .dinb(n291), .dout(n35295));
  jand g18033(.dina(n35295), .dinb(n35294), .dout(n35296));
  jor  g18034(.dina(n35296), .dinb(n34868), .dout(n35297));
  jxor g18035(.dina(n34862), .dinb(n292), .dout(n35298));
  jand g18036(.dina(n35298), .dinb(n35297), .dout(n35299));
  jor  g18037(.dina(n35299), .dinb(n34863), .dout(n35300));
  jxor g18038(.dina(n34850), .dinb(n293), .dout(n35301));
  jand g18039(.dina(n35301), .dinb(n35300), .dout(n35302));
  jor  g18040(.dina(n35302), .dinb(n34858), .dout(n35303));
  jand g18041(.dina(n35303), .dinb(n34857), .dout(n35304));
  jor  g18042(.dina(n35304), .dinb(n34854), .dout(n35305));
  jand g18043(.dina(n35305), .dinb(n303), .dout(n35306));
  jor  g18044(.dina(n35306), .dinb(n34850), .dout(n35307));
  jnot g18045(.din(n35306), .dout(n35308));
  jxor g18046(.dina(n35301), .dinb(n35300), .dout(n35309));
  jor  g18047(.dina(n35309), .dinb(n35308), .dout(n35310));
  jand g18048(.dina(n35310), .dinb(n35307), .dout(n35311));
  jand g18049(.dina(n35311), .dinb(n294), .dout(n35312));
  jor  g18050(.dina(n35306), .dinb(n34862), .dout(n35313));
  jxor g18051(.dina(n35298), .dinb(n35297), .dout(n35314));
  jor  g18052(.dina(n35314), .dinb(n35308), .dout(n35315));
  jand g18053(.dina(n35315), .dinb(n35313), .dout(n35316));
  jand g18054(.dina(n35316), .dinb(n293), .dout(n35317));
  jor  g18055(.dina(n35306), .dinb(n34867), .dout(n35318));
  jxor g18056(.dina(n35295), .dinb(n35294), .dout(n35319));
  jor  g18057(.dina(n35319), .dinb(n35308), .dout(n35320));
  jand g18058(.dina(n35320), .dinb(n35318), .dout(n35321));
  jand g18059(.dina(n35321), .dinb(n292), .dout(n35322));
  jor  g18060(.dina(n35306), .dinb(n34872), .dout(n35323));
  jxor g18061(.dina(n35292), .dinb(n35291), .dout(n35324));
  jor  g18062(.dina(n35324), .dinb(n35308), .dout(n35325));
  jand g18063(.dina(n35325), .dinb(n35323), .dout(n35326));
  jand g18064(.dina(n35326), .dinb(n291), .dout(n35327));
  jor  g18065(.dina(n35306), .dinb(n34877), .dout(n35328));
  jxor g18066(.dina(n35289), .dinb(n35288), .dout(n35329));
  jor  g18067(.dina(n35329), .dinb(n35308), .dout(n35330));
  jand g18068(.dina(n35330), .dinb(n35328), .dout(n35331));
  jand g18069(.dina(n35331), .dinb(n290), .dout(n35332));
  jor  g18070(.dina(n35306), .dinb(n34882), .dout(n35333));
  jxor g18071(.dina(n35286), .dinb(n35285), .dout(n35334));
  jor  g18072(.dina(n35334), .dinb(n35308), .dout(n35335));
  jand g18073(.dina(n35335), .dinb(n35333), .dout(n35336));
  jand g18074(.dina(n35336), .dinb(n289), .dout(n35337));
  jor  g18075(.dina(n35306), .dinb(n34887), .dout(n35338));
  jxor g18076(.dina(n35283), .dinb(n35282), .dout(n35339));
  jor  g18077(.dina(n35339), .dinb(n35308), .dout(n35340));
  jand g18078(.dina(n35340), .dinb(n35338), .dout(n35341));
  jand g18079(.dina(n35341), .dinb(n288), .dout(n35342));
  jor  g18080(.dina(n35306), .dinb(n34892), .dout(n35343));
  jxor g18081(.dina(n35280), .dinb(n35279), .dout(n35344));
  jor  g18082(.dina(n35344), .dinb(n35308), .dout(n35345));
  jand g18083(.dina(n35345), .dinb(n35343), .dout(n35346));
  jand g18084(.dina(n35346), .dinb(n287), .dout(n35347));
  jor  g18085(.dina(n35306), .dinb(n34897), .dout(n35348));
  jxor g18086(.dina(n35277), .dinb(n35276), .dout(n35349));
  jor  g18087(.dina(n35349), .dinb(n35308), .dout(n35350));
  jand g18088(.dina(n35350), .dinb(n35348), .dout(n35351));
  jand g18089(.dina(n35351), .dinb(n286), .dout(n35352));
  jor  g18090(.dina(n35306), .dinb(n34902), .dout(n35353));
  jxor g18091(.dina(n35274), .dinb(n35273), .dout(n35354));
  jor  g18092(.dina(n35354), .dinb(n35308), .dout(n35355));
  jand g18093(.dina(n35355), .dinb(n35353), .dout(n35356));
  jand g18094(.dina(n35356), .dinb(n285), .dout(n35357));
  jor  g18095(.dina(n35306), .dinb(n34907), .dout(n35358));
  jxor g18096(.dina(n35271), .dinb(n35270), .dout(n35359));
  jor  g18097(.dina(n35359), .dinb(n35308), .dout(n35360));
  jand g18098(.dina(n35360), .dinb(n35358), .dout(n35361));
  jand g18099(.dina(n35361), .dinb(n284), .dout(n35362));
  jor  g18100(.dina(n35306), .dinb(n34912), .dout(n35363));
  jxor g18101(.dina(n35268), .dinb(n35267), .dout(n35364));
  jor  g18102(.dina(n35364), .dinb(n35308), .dout(n35365));
  jand g18103(.dina(n35365), .dinb(n35363), .dout(n35366));
  jand g18104(.dina(n35366), .dinb(n317), .dout(n35367));
  jor  g18105(.dina(n35306), .dinb(n34917), .dout(n35368));
  jxor g18106(.dina(n35265), .dinb(n35264), .dout(n35369));
  jor  g18107(.dina(n35369), .dinb(n35308), .dout(n35370));
  jand g18108(.dina(n35370), .dinb(n35368), .dout(n35371));
  jand g18109(.dina(n35371), .dinb(n316), .dout(n35372));
  jor  g18110(.dina(n35306), .dinb(n34922), .dout(n35373));
  jxor g18111(.dina(n35262), .dinb(n35261), .dout(n35374));
  jor  g18112(.dina(n35374), .dinb(n35308), .dout(n35375));
  jand g18113(.dina(n35375), .dinb(n35373), .dout(n35376));
  jand g18114(.dina(n35376), .dinb(n315), .dout(n35377));
  jor  g18115(.dina(n35306), .dinb(n34927), .dout(n35378));
  jxor g18116(.dina(n35259), .dinb(n35258), .dout(n35379));
  jor  g18117(.dina(n35379), .dinb(n35308), .dout(n35380));
  jand g18118(.dina(n35380), .dinb(n35378), .dout(n35381));
  jand g18119(.dina(n35381), .dinb(n283), .dout(n35382));
  jor  g18120(.dina(n35306), .dinb(n34932), .dout(n35383));
  jxor g18121(.dina(n35256), .dinb(n35255), .dout(n35384));
  jor  g18122(.dina(n35384), .dinb(n35308), .dout(n35385));
  jand g18123(.dina(n35385), .dinb(n35383), .dout(n35386));
  jand g18124(.dina(n35386), .dinb(n280), .dout(n35387));
  jor  g18125(.dina(n35306), .dinb(n34937), .dout(n35388));
  jxor g18126(.dina(n35253), .dinb(n35252), .dout(n35389));
  jor  g18127(.dina(n35389), .dinb(n35308), .dout(n35390));
  jand g18128(.dina(n35390), .dinb(n35388), .dout(n35391));
  jand g18129(.dina(n35391), .dinb(n279), .dout(n35392));
  jor  g18130(.dina(n35306), .dinb(n34942), .dout(n35393));
  jxor g18131(.dina(n35250), .dinb(n35249), .dout(n35394));
  jor  g18132(.dina(n35394), .dinb(n35308), .dout(n35395));
  jand g18133(.dina(n35395), .dinb(n35393), .dout(n35396));
  jand g18134(.dina(n35396), .dinb(n278), .dout(n35397));
  jor  g18135(.dina(n35306), .dinb(n34947), .dout(n35398));
  jxor g18136(.dina(n35247), .dinb(n35246), .dout(n35399));
  jor  g18137(.dina(n35399), .dinb(n35308), .dout(n35400));
  jand g18138(.dina(n35400), .dinb(n35398), .dout(n35401));
  jand g18139(.dina(n35401), .dinb(n277), .dout(n35402));
  jor  g18140(.dina(n35306), .dinb(n34952), .dout(n35403));
  jxor g18141(.dina(n35244), .dinb(n35243), .dout(n35404));
  jor  g18142(.dina(n35404), .dinb(n35308), .dout(n35405));
  jand g18143(.dina(n35405), .dinb(n35403), .dout(n35406));
  jand g18144(.dina(n35406), .dinb(n326), .dout(n35407));
  jor  g18145(.dina(n35306), .dinb(n34957), .dout(n35408));
  jxor g18146(.dina(n35241), .dinb(n35240), .dout(n35409));
  jor  g18147(.dina(n35409), .dinb(n35308), .dout(n35410));
  jand g18148(.dina(n35410), .dinb(n35408), .dout(n35411));
  jand g18149(.dina(n35411), .dinb(n325), .dout(n35412));
  jor  g18150(.dina(n35306), .dinb(n34962), .dout(n35413));
  jxor g18151(.dina(n35238), .dinb(n35237), .dout(n35414));
  jor  g18152(.dina(n35414), .dinb(n35308), .dout(n35415));
  jand g18153(.dina(n35415), .dinb(n35413), .dout(n35416));
  jand g18154(.dina(n35416), .dinb(n324), .dout(n35417));
  jor  g18155(.dina(n35306), .dinb(n34967), .dout(n35418));
  jxor g18156(.dina(n35235), .dinb(n35234), .dout(n35419));
  jor  g18157(.dina(n35419), .dinb(n35308), .dout(n35420));
  jand g18158(.dina(n35420), .dinb(n35418), .dout(n35421));
  jand g18159(.dina(n35421), .dinb(n276), .dout(n35422));
  jor  g18160(.dina(n35306), .dinb(n34972), .dout(n35423));
  jxor g18161(.dina(n35232), .dinb(n35231), .dout(n35424));
  jor  g18162(.dina(n35424), .dinb(n35308), .dout(n35425));
  jand g18163(.dina(n35425), .dinb(n35423), .dout(n35426));
  jand g18164(.dina(n35426), .dinb(n333), .dout(n35427));
  jor  g18165(.dina(n35306), .dinb(n34977), .dout(n35428));
  jxor g18166(.dina(n35229), .dinb(n35228), .dout(n35429));
  jor  g18167(.dina(n35429), .dinb(n35308), .dout(n35430));
  jand g18168(.dina(n35430), .dinb(n35428), .dout(n35431));
  jand g18169(.dina(n35431), .dinb(n332), .dout(n35432));
  jor  g18170(.dina(n35306), .dinb(n34982), .dout(n35433));
  jxor g18171(.dina(n35226), .dinb(n35225), .dout(n35434));
  jor  g18172(.dina(n35434), .dinb(n35308), .dout(n35435));
  jand g18173(.dina(n35435), .dinb(n35433), .dout(n35436));
  jand g18174(.dina(n35436), .dinb(n331), .dout(n35437));
  jor  g18175(.dina(n35306), .dinb(n34987), .dout(n35438));
  jxor g18176(.dina(n35223), .dinb(n35222), .dout(n35439));
  jor  g18177(.dina(n35439), .dinb(n35308), .dout(n35440));
  jand g18178(.dina(n35440), .dinb(n35438), .dout(n35441));
  jand g18179(.dina(n35441), .dinb(n275), .dout(n35442));
  jor  g18180(.dina(n35306), .dinb(n34992), .dout(n35443));
  jxor g18181(.dina(n35220), .dinb(n35219), .dout(n35444));
  jor  g18182(.dina(n35444), .dinb(n35308), .dout(n35445));
  jand g18183(.dina(n35445), .dinb(n35443), .dout(n35446));
  jand g18184(.dina(n35446), .dinb(n340), .dout(n35447));
  jor  g18185(.dina(n35306), .dinb(n34997), .dout(n35448));
  jxor g18186(.dina(n35217), .dinb(n35216), .dout(n35449));
  jor  g18187(.dina(n35449), .dinb(n35308), .dout(n35450));
  jand g18188(.dina(n35450), .dinb(n35448), .dout(n35451));
  jand g18189(.dina(n35451), .dinb(n339), .dout(n35452));
  jor  g18190(.dina(n35306), .dinb(n35002), .dout(n35453));
  jxor g18191(.dina(n35214), .dinb(n35213), .dout(n35454));
  jor  g18192(.dina(n35454), .dinb(n35308), .dout(n35455));
  jand g18193(.dina(n35455), .dinb(n35453), .dout(n35456));
  jand g18194(.dina(n35456), .dinb(n338), .dout(n35457));
  jor  g18195(.dina(n35306), .dinb(n35007), .dout(n35458));
  jxor g18196(.dina(n35211), .dinb(n35210), .dout(n35459));
  jor  g18197(.dina(n35459), .dinb(n35308), .dout(n35460));
  jand g18198(.dina(n35460), .dinb(n35458), .dout(n35461));
  jand g18199(.dina(n35461), .dinb(n271), .dout(n35462));
  jor  g18200(.dina(n35306), .dinb(n35012), .dout(n35463));
  jxor g18201(.dina(n35208), .dinb(n35207), .dout(n35464));
  jor  g18202(.dina(n35464), .dinb(n35308), .dout(n35465));
  jand g18203(.dina(n35465), .dinb(n35463), .dout(n35466));
  jand g18204(.dina(n35466), .dinb(n270), .dout(n35467));
  jor  g18205(.dina(n35306), .dinb(n35017), .dout(n35468));
  jxor g18206(.dina(n35205), .dinb(n35204), .dout(n35469));
  jor  g18207(.dina(n35469), .dinb(n35308), .dout(n35470));
  jand g18208(.dina(n35470), .dinb(n35468), .dout(n35471));
  jand g18209(.dina(n35471), .dinb(n269), .dout(n35472));
  jor  g18210(.dina(n35306), .dinb(n35022), .dout(n35473));
  jxor g18211(.dina(n35202), .dinb(n35201), .dout(n35474));
  jor  g18212(.dina(n35474), .dinb(n35308), .dout(n35475));
  jand g18213(.dina(n35475), .dinb(n35473), .dout(n35476));
  jand g18214(.dina(n35476), .dinb(n274), .dout(n35477));
  jor  g18215(.dina(n35306), .dinb(n35027), .dout(n35478));
  jxor g18216(.dina(n35199), .dinb(n35198), .dout(n35479));
  jor  g18217(.dina(n35479), .dinb(n35308), .dout(n35480));
  jand g18218(.dina(n35480), .dinb(n35478), .dout(n35481));
  jand g18219(.dina(n35481), .dinb(n268), .dout(n35482));
  jor  g18220(.dina(n35306), .dinb(n35032), .dout(n35483));
  jxor g18221(.dina(n35196), .dinb(n35195), .dout(n35484));
  jor  g18222(.dina(n35484), .dinb(n35308), .dout(n35485));
  jand g18223(.dina(n35485), .dinb(n35483), .dout(n35486));
  jand g18224(.dina(n35486), .dinb(n349), .dout(n35487));
  jor  g18225(.dina(n35306), .dinb(n35037), .dout(n35488));
  jxor g18226(.dina(n35193), .dinb(n35192), .dout(n35489));
  jor  g18227(.dina(n35489), .dinb(n35308), .dout(n35490));
  jand g18228(.dina(n35490), .dinb(n35488), .dout(n35491));
  jand g18229(.dina(n35491), .dinb(n348), .dout(n35492));
  jor  g18230(.dina(n35306), .dinb(n35042), .dout(n35493));
  jxor g18231(.dina(n35190), .dinb(n35189), .dout(n35494));
  jor  g18232(.dina(n35494), .dinb(n35308), .dout(n35495));
  jand g18233(.dina(n35495), .dinb(n35493), .dout(n35496));
  jand g18234(.dina(n35496), .dinb(n347), .dout(n35497));
  jor  g18235(.dina(n35306), .dinb(n35047), .dout(n35498));
  jxor g18236(.dina(n35187), .dinb(n35186), .dout(n35499));
  jor  g18237(.dina(n35499), .dinb(n35308), .dout(n35500));
  jand g18238(.dina(n35500), .dinb(n35498), .dout(n35501));
  jand g18239(.dina(n35501), .dinb(n267), .dout(n35502));
  jor  g18240(.dina(n35306), .dinb(n35052), .dout(n35503));
  jxor g18241(.dina(n35184), .dinb(n35183), .dout(n35504));
  jor  g18242(.dina(n35504), .dinb(n35308), .dout(n35505));
  jand g18243(.dina(n35505), .dinb(n35503), .dout(n35506));
  jand g18244(.dina(n35506), .dinb(n266), .dout(n35507));
  jor  g18245(.dina(n35306), .dinb(n35057), .dout(n35508));
  jxor g18246(.dina(n35181), .dinb(n35180), .dout(n35509));
  jor  g18247(.dina(n35509), .dinb(n35308), .dout(n35510));
  jand g18248(.dina(n35510), .dinb(n35508), .dout(n35511));
  jand g18249(.dina(n35511), .dinb(n356), .dout(n35512));
  jor  g18250(.dina(n35306), .dinb(n35062), .dout(n35513));
  jxor g18251(.dina(n35178), .dinb(n35177), .dout(n35514));
  jor  g18252(.dina(n35514), .dinb(n35308), .dout(n35515));
  jand g18253(.dina(n35515), .dinb(n35513), .dout(n35516));
  jand g18254(.dina(n35516), .dinb(n355), .dout(n35517));
  jor  g18255(.dina(n35306), .dinb(n35067), .dout(n35518));
  jxor g18256(.dina(n35175), .dinb(n35174), .dout(n35519));
  jor  g18257(.dina(n35519), .dinb(n35308), .dout(n35520));
  jand g18258(.dina(n35520), .dinb(n35518), .dout(n35521));
  jand g18259(.dina(n35521), .dinb(n364), .dout(n35522));
  jor  g18260(.dina(n35306), .dinb(n35072), .dout(n35523));
  jxor g18261(.dina(n35172), .dinb(n35171), .dout(n35524));
  jor  g18262(.dina(n35524), .dinb(n35308), .dout(n35525));
  jand g18263(.dina(n35525), .dinb(n35523), .dout(n35526));
  jand g18264(.dina(n35526), .dinb(n361), .dout(n35527));
  jor  g18265(.dina(n35306), .dinb(n35077), .dout(n35528));
  jxor g18266(.dina(n35169), .dinb(n35168), .dout(n35529));
  jor  g18267(.dina(n35529), .dinb(n35308), .dout(n35530));
  jand g18268(.dina(n35530), .dinb(n35528), .dout(n35531));
  jand g18269(.dina(n35531), .dinb(n360), .dout(n35532));
  jor  g18270(.dina(n35306), .dinb(n35082), .dout(n35533));
  jxor g18271(.dina(n35166), .dinb(n35165), .dout(n35534));
  jor  g18272(.dina(n35534), .dinb(n35308), .dout(n35535));
  jand g18273(.dina(n35535), .dinb(n35533), .dout(n35536));
  jand g18274(.dina(n35536), .dinb(n363), .dout(n35537));
  jor  g18275(.dina(n35306), .dinb(n35087), .dout(n35538));
  jxor g18276(.dina(n35163), .dinb(n35162), .dout(n35539));
  jor  g18277(.dina(n35539), .dinb(n35308), .dout(n35540));
  jand g18278(.dina(n35540), .dinb(n35538), .dout(n35541));
  jand g18279(.dina(n35541), .dinb(n359), .dout(n35542));
  jor  g18280(.dina(n35306), .dinb(n35092), .dout(n35543));
  jxor g18281(.dina(n35160), .dinb(n35159), .dout(n35544));
  jor  g18282(.dina(n35544), .dinb(n35308), .dout(n35545));
  jand g18283(.dina(n35545), .dinb(n35543), .dout(n35546));
  jand g18284(.dina(n35546), .dinb(n369), .dout(n35547));
  jor  g18285(.dina(n35306), .dinb(n35097), .dout(n35548));
  jxor g18286(.dina(n35157), .dinb(n35156), .dout(n35549));
  jor  g18287(.dina(n35549), .dinb(n35308), .dout(n35550));
  jand g18288(.dina(n35550), .dinb(n35548), .dout(n35551));
  jand g18289(.dina(n35551), .dinb(n368), .dout(n35552));
  jor  g18290(.dina(n35306), .dinb(n35102), .dout(n35553));
  jxor g18291(.dina(n35154), .dinb(n35153), .dout(n35554));
  jor  g18292(.dina(n35554), .dinb(n35308), .dout(n35555));
  jand g18293(.dina(n35555), .dinb(n35553), .dout(n35556));
  jand g18294(.dina(n35556), .dinb(n367), .dout(n35557));
  jor  g18295(.dina(n35306), .dinb(n35107), .dout(n35558));
  jxor g18296(.dina(n35151), .dinb(n35150), .dout(n35559));
  jor  g18297(.dina(n35559), .dinb(n35308), .dout(n35560));
  jand g18298(.dina(n35560), .dinb(n35558), .dout(n35561));
  jand g18299(.dina(n35561), .dinb(n265), .dout(n35562));
  jor  g18300(.dina(n35306), .dinb(n35112), .dout(n35563));
  jxor g18301(.dina(n35148), .dinb(n35147), .dout(n35564));
  jor  g18302(.dina(n35564), .dinb(n35308), .dout(n35565));
  jand g18303(.dina(n35565), .dinb(n35563), .dout(n35566));
  jand g18304(.dina(n35566), .dinb(n378), .dout(n35567));
  jor  g18305(.dina(n35306), .dinb(n35118), .dout(n35568));
  jxor g18306(.dina(n35145), .dinb(n35144), .dout(n35569));
  jor  g18307(.dina(n35569), .dinb(n35308), .dout(n35570));
  jand g18308(.dina(n35570), .dinb(n35568), .dout(n35571));
  jand g18309(.dina(n35571), .dinb(n377), .dout(n35572));
  jor  g18310(.dina(n35306), .dinb(n35123), .dout(n35573));
  jxor g18311(.dina(n35142), .dinb(n35141), .dout(n35574));
  jor  g18312(.dina(n35574), .dinb(n35308), .dout(n35575));
  jand g18313(.dina(n35575), .dinb(n35573), .dout(n35576));
  jand g18314(.dina(n35576), .dinb(n376), .dout(n35577));
  jor  g18315(.dina(n35306), .dinb(n35130), .dout(n35578));
  jxor g18316(.dina(n35139), .dinb(n35138), .dout(n35579));
  jor  g18317(.dina(n35579), .dinb(n35308), .dout(n35580));
  jand g18318(.dina(n35580), .dinb(n35578), .dout(n35581));
  jand g18319(.dina(n35581), .dinb(n264), .dout(n35582));
  jxor g18320(.dina(n35136), .dinb(n14663), .dout(n35583));
  jand g18321(.dina(n35583), .dinb(n35306), .dout(n35584));
  jnot g18322(.din(n35584), .dout(n35585));
  jor  g18323(.dina(n35306), .dinb(n35135), .dout(n35586));
  jand g18324(.dina(n35586), .dinb(n35585), .dout(n35587));
  jnot g18325(.din(n35587), .dout(n35588));
  jand g18326(.dina(n35588), .dinb(n386), .dout(n35589));
  jnot g18327(.din(n15122), .dout(n35590));
  jnot g18328(.din(n34854), .dout(n35591));
  jnot g18329(.din(n34858), .dout(n35592));
  jnot g18330(.din(n34863), .dout(n35593));
  jnot g18331(.din(n34868), .dout(n35594));
  jnot g18332(.din(n34873), .dout(n35595));
  jnot g18333(.din(n34878), .dout(n35596));
  jnot g18334(.din(n34883), .dout(n35597));
  jnot g18335(.din(n34888), .dout(n35598));
  jnot g18336(.din(n34893), .dout(n35599));
  jnot g18337(.din(n34898), .dout(n35600));
  jnot g18338(.din(n34903), .dout(n35601));
  jnot g18339(.din(n34908), .dout(n35602));
  jnot g18340(.din(n34913), .dout(n35603));
  jnot g18341(.din(n34918), .dout(n35604));
  jnot g18342(.din(n34923), .dout(n35605));
  jnot g18343(.din(n34928), .dout(n35606));
  jnot g18344(.din(n34933), .dout(n35607));
  jnot g18345(.din(n34938), .dout(n35608));
  jnot g18346(.din(n34943), .dout(n35609));
  jnot g18347(.din(n34948), .dout(n35610));
  jnot g18348(.din(n34953), .dout(n35611));
  jnot g18349(.din(n34958), .dout(n35612));
  jnot g18350(.din(n34963), .dout(n35613));
  jnot g18351(.din(n34968), .dout(n35614));
  jnot g18352(.din(n34973), .dout(n35615));
  jnot g18353(.din(n34978), .dout(n35616));
  jnot g18354(.din(n34983), .dout(n35617));
  jnot g18355(.din(n34988), .dout(n35618));
  jnot g18356(.din(n34993), .dout(n35619));
  jnot g18357(.din(n34998), .dout(n35620));
  jnot g18358(.din(n35003), .dout(n35621));
  jnot g18359(.din(n35008), .dout(n35622));
  jnot g18360(.din(n35013), .dout(n35623));
  jnot g18361(.din(n35018), .dout(n35624));
  jnot g18362(.din(n35023), .dout(n35625));
  jnot g18363(.din(n35028), .dout(n35626));
  jnot g18364(.din(n35033), .dout(n35627));
  jnot g18365(.din(n35038), .dout(n35628));
  jnot g18366(.din(n35043), .dout(n35629));
  jnot g18367(.din(n35048), .dout(n35630));
  jnot g18368(.din(n35053), .dout(n35631));
  jnot g18369(.din(n35058), .dout(n35632));
  jnot g18370(.din(n35063), .dout(n35633));
  jnot g18371(.din(n35068), .dout(n35634));
  jnot g18372(.din(n35073), .dout(n35635));
  jnot g18373(.din(n35078), .dout(n35636));
  jnot g18374(.din(n35083), .dout(n35637));
  jnot g18375(.din(n35088), .dout(n35638));
  jnot g18376(.din(n35093), .dout(n35639));
  jnot g18377(.din(n35098), .dout(n35640));
  jnot g18378(.din(n35103), .dout(n35641));
  jnot g18379(.din(n35108), .dout(n35642));
  jnot g18380(.din(n35113), .dout(n35643));
  jnot g18381(.din(n35119), .dout(n35644));
  jnot g18382(.din(n35124), .dout(n35645));
  jnot g18383(.din(n35131), .dout(n35646));
  jnot g18384(.din(n35134), .dout(n35647));
  jxor g18385(.dina(n35135), .dinb(n259), .dout(n35648));
  jor  g18386(.dina(n35648), .dinb(n14662), .dout(n35649));
  jand g18387(.dina(n35649), .dinb(n35647), .dout(n35650));
  jnot g18388(.din(n35139), .dout(n35651));
  jor  g18389(.dina(n35651), .dinb(n35650), .dout(n35652));
  jand g18390(.dina(n35652), .dinb(n35646), .dout(n35653));
  jnot g18391(.din(n35142), .dout(n35654));
  jor  g18392(.dina(n35654), .dinb(n35653), .dout(n35655));
  jand g18393(.dina(n35655), .dinb(n35645), .dout(n35656));
  jnot g18394(.din(n35145), .dout(n35657));
  jor  g18395(.dina(n35657), .dinb(n35656), .dout(n35658));
  jand g18396(.dina(n35658), .dinb(n35644), .dout(n35659));
  jnot g18397(.din(n35148), .dout(n35660));
  jor  g18398(.dina(n35660), .dinb(n35659), .dout(n35661));
  jand g18399(.dina(n35661), .dinb(n35643), .dout(n35662));
  jnot g18400(.din(n35151), .dout(n35663));
  jor  g18401(.dina(n35663), .dinb(n35662), .dout(n35664));
  jand g18402(.dina(n35664), .dinb(n35642), .dout(n35665));
  jnot g18403(.din(n35154), .dout(n35666));
  jor  g18404(.dina(n35666), .dinb(n35665), .dout(n35667));
  jand g18405(.dina(n35667), .dinb(n35641), .dout(n35668));
  jnot g18406(.din(n35157), .dout(n35669));
  jor  g18407(.dina(n35669), .dinb(n35668), .dout(n35670));
  jand g18408(.dina(n35670), .dinb(n35640), .dout(n35671));
  jnot g18409(.din(n35160), .dout(n35672));
  jor  g18410(.dina(n35672), .dinb(n35671), .dout(n35673));
  jand g18411(.dina(n35673), .dinb(n35639), .dout(n35674));
  jnot g18412(.din(n35163), .dout(n35675));
  jor  g18413(.dina(n35675), .dinb(n35674), .dout(n35676));
  jand g18414(.dina(n35676), .dinb(n35638), .dout(n35677));
  jnot g18415(.din(n35166), .dout(n35678));
  jor  g18416(.dina(n35678), .dinb(n35677), .dout(n35679));
  jand g18417(.dina(n35679), .dinb(n35637), .dout(n35680));
  jnot g18418(.din(n35169), .dout(n35681));
  jor  g18419(.dina(n35681), .dinb(n35680), .dout(n35682));
  jand g18420(.dina(n35682), .dinb(n35636), .dout(n35683));
  jnot g18421(.din(n35172), .dout(n35684));
  jor  g18422(.dina(n35684), .dinb(n35683), .dout(n35685));
  jand g18423(.dina(n35685), .dinb(n35635), .dout(n35686));
  jnot g18424(.din(n35175), .dout(n35687));
  jor  g18425(.dina(n35687), .dinb(n35686), .dout(n35688));
  jand g18426(.dina(n35688), .dinb(n35634), .dout(n35689));
  jnot g18427(.din(n35178), .dout(n35690));
  jor  g18428(.dina(n35690), .dinb(n35689), .dout(n35691));
  jand g18429(.dina(n35691), .dinb(n35633), .dout(n35692));
  jnot g18430(.din(n35181), .dout(n35693));
  jor  g18431(.dina(n35693), .dinb(n35692), .dout(n35694));
  jand g18432(.dina(n35694), .dinb(n35632), .dout(n35695));
  jnot g18433(.din(n35184), .dout(n35696));
  jor  g18434(.dina(n35696), .dinb(n35695), .dout(n35697));
  jand g18435(.dina(n35697), .dinb(n35631), .dout(n35698));
  jnot g18436(.din(n35187), .dout(n35699));
  jor  g18437(.dina(n35699), .dinb(n35698), .dout(n35700));
  jand g18438(.dina(n35700), .dinb(n35630), .dout(n35701));
  jnot g18439(.din(n35190), .dout(n35702));
  jor  g18440(.dina(n35702), .dinb(n35701), .dout(n35703));
  jand g18441(.dina(n35703), .dinb(n35629), .dout(n35704));
  jnot g18442(.din(n35193), .dout(n35705));
  jor  g18443(.dina(n35705), .dinb(n35704), .dout(n35706));
  jand g18444(.dina(n35706), .dinb(n35628), .dout(n35707));
  jnot g18445(.din(n35196), .dout(n35708));
  jor  g18446(.dina(n35708), .dinb(n35707), .dout(n35709));
  jand g18447(.dina(n35709), .dinb(n35627), .dout(n35710));
  jnot g18448(.din(n35199), .dout(n35711));
  jor  g18449(.dina(n35711), .dinb(n35710), .dout(n35712));
  jand g18450(.dina(n35712), .dinb(n35626), .dout(n35713));
  jnot g18451(.din(n35202), .dout(n35714));
  jor  g18452(.dina(n35714), .dinb(n35713), .dout(n35715));
  jand g18453(.dina(n35715), .dinb(n35625), .dout(n35716));
  jnot g18454(.din(n35205), .dout(n35717));
  jor  g18455(.dina(n35717), .dinb(n35716), .dout(n35718));
  jand g18456(.dina(n35718), .dinb(n35624), .dout(n35719));
  jnot g18457(.din(n35208), .dout(n35720));
  jor  g18458(.dina(n35720), .dinb(n35719), .dout(n35721));
  jand g18459(.dina(n35721), .dinb(n35623), .dout(n35722));
  jnot g18460(.din(n35211), .dout(n35723));
  jor  g18461(.dina(n35723), .dinb(n35722), .dout(n35724));
  jand g18462(.dina(n35724), .dinb(n35622), .dout(n35725));
  jnot g18463(.din(n35214), .dout(n35726));
  jor  g18464(.dina(n35726), .dinb(n35725), .dout(n35727));
  jand g18465(.dina(n35727), .dinb(n35621), .dout(n35728));
  jnot g18466(.din(n35217), .dout(n35729));
  jor  g18467(.dina(n35729), .dinb(n35728), .dout(n35730));
  jand g18468(.dina(n35730), .dinb(n35620), .dout(n35731));
  jnot g18469(.din(n35220), .dout(n35732));
  jor  g18470(.dina(n35732), .dinb(n35731), .dout(n35733));
  jand g18471(.dina(n35733), .dinb(n35619), .dout(n35734));
  jnot g18472(.din(n35223), .dout(n35735));
  jor  g18473(.dina(n35735), .dinb(n35734), .dout(n35736));
  jand g18474(.dina(n35736), .dinb(n35618), .dout(n35737));
  jnot g18475(.din(n35226), .dout(n35738));
  jor  g18476(.dina(n35738), .dinb(n35737), .dout(n35739));
  jand g18477(.dina(n35739), .dinb(n35617), .dout(n35740));
  jnot g18478(.din(n35229), .dout(n35741));
  jor  g18479(.dina(n35741), .dinb(n35740), .dout(n35742));
  jand g18480(.dina(n35742), .dinb(n35616), .dout(n35743));
  jnot g18481(.din(n35232), .dout(n35744));
  jor  g18482(.dina(n35744), .dinb(n35743), .dout(n35745));
  jand g18483(.dina(n35745), .dinb(n35615), .dout(n35746));
  jnot g18484(.din(n35235), .dout(n35747));
  jor  g18485(.dina(n35747), .dinb(n35746), .dout(n35748));
  jand g18486(.dina(n35748), .dinb(n35614), .dout(n35749));
  jnot g18487(.din(n35238), .dout(n35750));
  jor  g18488(.dina(n35750), .dinb(n35749), .dout(n35751));
  jand g18489(.dina(n35751), .dinb(n35613), .dout(n35752));
  jnot g18490(.din(n35241), .dout(n35753));
  jor  g18491(.dina(n35753), .dinb(n35752), .dout(n35754));
  jand g18492(.dina(n35754), .dinb(n35612), .dout(n35755));
  jnot g18493(.din(n35244), .dout(n35756));
  jor  g18494(.dina(n35756), .dinb(n35755), .dout(n35757));
  jand g18495(.dina(n35757), .dinb(n35611), .dout(n35758));
  jnot g18496(.din(n35247), .dout(n35759));
  jor  g18497(.dina(n35759), .dinb(n35758), .dout(n35760));
  jand g18498(.dina(n35760), .dinb(n35610), .dout(n35761));
  jnot g18499(.din(n35250), .dout(n35762));
  jor  g18500(.dina(n35762), .dinb(n35761), .dout(n35763));
  jand g18501(.dina(n35763), .dinb(n35609), .dout(n35764));
  jnot g18502(.din(n35253), .dout(n35765));
  jor  g18503(.dina(n35765), .dinb(n35764), .dout(n35766));
  jand g18504(.dina(n35766), .dinb(n35608), .dout(n35767));
  jnot g18505(.din(n35256), .dout(n35768));
  jor  g18506(.dina(n35768), .dinb(n35767), .dout(n35769));
  jand g18507(.dina(n35769), .dinb(n35607), .dout(n35770));
  jnot g18508(.din(n35259), .dout(n35771));
  jor  g18509(.dina(n35771), .dinb(n35770), .dout(n35772));
  jand g18510(.dina(n35772), .dinb(n35606), .dout(n35773));
  jnot g18511(.din(n35262), .dout(n35774));
  jor  g18512(.dina(n35774), .dinb(n35773), .dout(n35775));
  jand g18513(.dina(n35775), .dinb(n35605), .dout(n35776));
  jnot g18514(.din(n35265), .dout(n35777));
  jor  g18515(.dina(n35777), .dinb(n35776), .dout(n35778));
  jand g18516(.dina(n35778), .dinb(n35604), .dout(n35779));
  jnot g18517(.din(n35268), .dout(n35780));
  jor  g18518(.dina(n35780), .dinb(n35779), .dout(n35781));
  jand g18519(.dina(n35781), .dinb(n35603), .dout(n35782));
  jnot g18520(.din(n35271), .dout(n35783));
  jor  g18521(.dina(n35783), .dinb(n35782), .dout(n35784));
  jand g18522(.dina(n35784), .dinb(n35602), .dout(n35785));
  jnot g18523(.din(n35274), .dout(n35786));
  jor  g18524(.dina(n35786), .dinb(n35785), .dout(n35787));
  jand g18525(.dina(n35787), .dinb(n35601), .dout(n35788));
  jnot g18526(.din(n35277), .dout(n35789));
  jor  g18527(.dina(n35789), .dinb(n35788), .dout(n35790));
  jand g18528(.dina(n35790), .dinb(n35600), .dout(n35791));
  jnot g18529(.din(n35280), .dout(n35792));
  jor  g18530(.dina(n35792), .dinb(n35791), .dout(n35793));
  jand g18531(.dina(n35793), .dinb(n35599), .dout(n35794));
  jnot g18532(.din(n35283), .dout(n35795));
  jor  g18533(.dina(n35795), .dinb(n35794), .dout(n35796));
  jand g18534(.dina(n35796), .dinb(n35598), .dout(n35797));
  jnot g18535(.din(n35286), .dout(n35798));
  jor  g18536(.dina(n35798), .dinb(n35797), .dout(n35799));
  jand g18537(.dina(n35799), .dinb(n35597), .dout(n35800));
  jnot g18538(.din(n35289), .dout(n35801));
  jor  g18539(.dina(n35801), .dinb(n35800), .dout(n35802));
  jand g18540(.dina(n35802), .dinb(n35596), .dout(n35803));
  jnot g18541(.din(n35292), .dout(n35804));
  jor  g18542(.dina(n35804), .dinb(n35803), .dout(n35805));
  jand g18543(.dina(n35805), .dinb(n35595), .dout(n35806));
  jnot g18544(.din(n35295), .dout(n35807));
  jor  g18545(.dina(n35807), .dinb(n35806), .dout(n35808));
  jand g18546(.dina(n35808), .dinb(n35594), .dout(n35809));
  jnot g18547(.din(n35298), .dout(n35810));
  jor  g18548(.dina(n35810), .dinb(n35809), .dout(n35811));
  jand g18549(.dina(n35811), .dinb(n35593), .dout(n35812));
  jnot g18550(.din(n35301), .dout(n35813));
  jor  g18551(.dina(n35813), .dinb(n35812), .dout(n35814));
  jand g18552(.dina(n35814), .dinb(n35592), .dout(n35815));
  jor  g18553(.dina(n35815), .dinb(n34856), .dout(n35816));
  jand g18554(.dina(n35816), .dinb(n35591), .dout(n35817));
  jor  g18555(.dina(n35817), .dinb(n35590), .dout(n35818));
  jand g18556(.dina(n35818), .dinb(a6 ), .dout(n35819));
  jnot g18557(.din(n15125), .dout(n35820));
  jor  g18558(.dina(n35817), .dinb(n35820), .dout(n35821));
  jnot g18559(.din(n35821), .dout(n35822));
  jor  g18560(.dina(n35822), .dinb(n35819), .dout(n35823));
  jand g18561(.dina(n35823), .dinb(n259), .dout(n35824));
  jand g18562(.dina(n35305), .dinb(n15122), .dout(n35825));
  jor  g18563(.dina(n35825), .dinb(n14661), .dout(n35826));
  jand g18564(.dina(n35821), .dinb(n35826), .dout(n35827));
  jxor g18565(.dina(n35827), .dinb(b1 ), .dout(n35828));
  jand g18566(.dina(n35828), .dinb(n15133), .dout(n35829));
  jor  g18567(.dina(n35829), .dinb(n35824), .dout(n35830));
  jxor g18568(.dina(n35587), .dinb(b2 ), .dout(n35831));
  jand g18569(.dina(n35831), .dinb(n35830), .dout(n35832));
  jor  g18570(.dina(n35832), .dinb(n35589), .dout(n35833));
  jxor g18571(.dina(n35581), .dinb(n264), .dout(n35834));
  jand g18572(.dina(n35834), .dinb(n35833), .dout(n35835));
  jor  g18573(.dina(n35835), .dinb(n35582), .dout(n35836));
  jxor g18574(.dina(n35576), .dinb(n376), .dout(n35837));
  jand g18575(.dina(n35837), .dinb(n35836), .dout(n35838));
  jor  g18576(.dina(n35838), .dinb(n35577), .dout(n35839));
  jxor g18577(.dina(n35571), .dinb(n377), .dout(n35840));
  jand g18578(.dina(n35840), .dinb(n35839), .dout(n35841));
  jor  g18579(.dina(n35841), .dinb(n35572), .dout(n35842));
  jxor g18580(.dina(n35566), .dinb(n378), .dout(n35843));
  jand g18581(.dina(n35843), .dinb(n35842), .dout(n35844));
  jor  g18582(.dina(n35844), .dinb(n35567), .dout(n35845));
  jxor g18583(.dina(n35561), .dinb(n265), .dout(n35846));
  jand g18584(.dina(n35846), .dinb(n35845), .dout(n35847));
  jor  g18585(.dina(n35847), .dinb(n35562), .dout(n35848));
  jxor g18586(.dina(n35556), .dinb(n367), .dout(n35849));
  jand g18587(.dina(n35849), .dinb(n35848), .dout(n35850));
  jor  g18588(.dina(n35850), .dinb(n35557), .dout(n35851));
  jxor g18589(.dina(n35551), .dinb(n368), .dout(n35852));
  jand g18590(.dina(n35852), .dinb(n35851), .dout(n35853));
  jor  g18591(.dina(n35853), .dinb(n35552), .dout(n35854));
  jxor g18592(.dina(n35546), .dinb(n369), .dout(n35855));
  jand g18593(.dina(n35855), .dinb(n35854), .dout(n35856));
  jor  g18594(.dina(n35856), .dinb(n35547), .dout(n35857));
  jxor g18595(.dina(n35541), .dinb(n359), .dout(n35858));
  jand g18596(.dina(n35858), .dinb(n35857), .dout(n35859));
  jor  g18597(.dina(n35859), .dinb(n35542), .dout(n35860));
  jxor g18598(.dina(n35536), .dinb(n363), .dout(n35861));
  jand g18599(.dina(n35861), .dinb(n35860), .dout(n35862));
  jor  g18600(.dina(n35862), .dinb(n35537), .dout(n35863));
  jxor g18601(.dina(n35531), .dinb(n360), .dout(n35864));
  jand g18602(.dina(n35864), .dinb(n35863), .dout(n35865));
  jor  g18603(.dina(n35865), .dinb(n35532), .dout(n35866));
  jxor g18604(.dina(n35526), .dinb(n361), .dout(n35867));
  jand g18605(.dina(n35867), .dinb(n35866), .dout(n35868));
  jor  g18606(.dina(n35868), .dinb(n35527), .dout(n35869));
  jxor g18607(.dina(n35521), .dinb(n364), .dout(n35870));
  jand g18608(.dina(n35870), .dinb(n35869), .dout(n35871));
  jor  g18609(.dina(n35871), .dinb(n35522), .dout(n35872));
  jxor g18610(.dina(n35516), .dinb(n355), .dout(n35873));
  jand g18611(.dina(n35873), .dinb(n35872), .dout(n35874));
  jor  g18612(.dina(n35874), .dinb(n35517), .dout(n35875));
  jxor g18613(.dina(n35511), .dinb(n356), .dout(n35876));
  jand g18614(.dina(n35876), .dinb(n35875), .dout(n35877));
  jor  g18615(.dina(n35877), .dinb(n35512), .dout(n35878));
  jxor g18616(.dina(n35506), .dinb(n266), .dout(n35879));
  jand g18617(.dina(n35879), .dinb(n35878), .dout(n35880));
  jor  g18618(.dina(n35880), .dinb(n35507), .dout(n35881));
  jxor g18619(.dina(n35501), .dinb(n267), .dout(n35882));
  jand g18620(.dina(n35882), .dinb(n35881), .dout(n35883));
  jor  g18621(.dina(n35883), .dinb(n35502), .dout(n35884));
  jxor g18622(.dina(n35496), .dinb(n347), .dout(n35885));
  jand g18623(.dina(n35885), .dinb(n35884), .dout(n35886));
  jor  g18624(.dina(n35886), .dinb(n35497), .dout(n35887));
  jxor g18625(.dina(n35491), .dinb(n348), .dout(n35888));
  jand g18626(.dina(n35888), .dinb(n35887), .dout(n35889));
  jor  g18627(.dina(n35889), .dinb(n35492), .dout(n35890));
  jxor g18628(.dina(n35486), .dinb(n349), .dout(n35891));
  jand g18629(.dina(n35891), .dinb(n35890), .dout(n35892));
  jor  g18630(.dina(n35892), .dinb(n35487), .dout(n35893));
  jxor g18631(.dina(n35481), .dinb(n268), .dout(n35894));
  jand g18632(.dina(n35894), .dinb(n35893), .dout(n35895));
  jor  g18633(.dina(n35895), .dinb(n35482), .dout(n35896));
  jxor g18634(.dina(n35476), .dinb(n274), .dout(n35897));
  jand g18635(.dina(n35897), .dinb(n35896), .dout(n35898));
  jor  g18636(.dina(n35898), .dinb(n35477), .dout(n35899));
  jxor g18637(.dina(n35471), .dinb(n269), .dout(n35900));
  jand g18638(.dina(n35900), .dinb(n35899), .dout(n35901));
  jor  g18639(.dina(n35901), .dinb(n35472), .dout(n35902));
  jxor g18640(.dina(n35466), .dinb(n270), .dout(n35903));
  jand g18641(.dina(n35903), .dinb(n35902), .dout(n35904));
  jor  g18642(.dina(n35904), .dinb(n35467), .dout(n35905));
  jxor g18643(.dina(n35461), .dinb(n271), .dout(n35906));
  jand g18644(.dina(n35906), .dinb(n35905), .dout(n35907));
  jor  g18645(.dina(n35907), .dinb(n35462), .dout(n35908));
  jxor g18646(.dina(n35456), .dinb(n338), .dout(n35909));
  jand g18647(.dina(n35909), .dinb(n35908), .dout(n35910));
  jor  g18648(.dina(n35910), .dinb(n35457), .dout(n35911));
  jxor g18649(.dina(n35451), .dinb(n339), .dout(n35912));
  jand g18650(.dina(n35912), .dinb(n35911), .dout(n35913));
  jor  g18651(.dina(n35913), .dinb(n35452), .dout(n35914));
  jxor g18652(.dina(n35446), .dinb(n340), .dout(n35915));
  jand g18653(.dina(n35915), .dinb(n35914), .dout(n35916));
  jor  g18654(.dina(n35916), .dinb(n35447), .dout(n35917));
  jxor g18655(.dina(n35441), .dinb(n275), .dout(n35918));
  jand g18656(.dina(n35918), .dinb(n35917), .dout(n35919));
  jor  g18657(.dina(n35919), .dinb(n35442), .dout(n35920));
  jxor g18658(.dina(n35436), .dinb(n331), .dout(n35921));
  jand g18659(.dina(n35921), .dinb(n35920), .dout(n35922));
  jor  g18660(.dina(n35922), .dinb(n35437), .dout(n35923));
  jxor g18661(.dina(n35431), .dinb(n332), .dout(n35924));
  jand g18662(.dina(n35924), .dinb(n35923), .dout(n35925));
  jor  g18663(.dina(n35925), .dinb(n35432), .dout(n35926));
  jxor g18664(.dina(n35426), .dinb(n333), .dout(n35927));
  jand g18665(.dina(n35927), .dinb(n35926), .dout(n35928));
  jor  g18666(.dina(n35928), .dinb(n35427), .dout(n35929));
  jxor g18667(.dina(n35421), .dinb(n276), .dout(n35930));
  jand g18668(.dina(n35930), .dinb(n35929), .dout(n35931));
  jor  g18669(.dina(n35931), .dinb(n35422), .dout(n35932));
  jxor g18670(.dina(n35416), .dinb(n324), .dout(n35933));
  jand g18671(.dina(n35933), .dinb(n35932), .dout(n35934));
  jor  g18672(.dina(n35934), .dinb(n35417), .dout(n35935));
  jxor g18673(.dina(n35411), .dinb(n325), .dout(n35936));
  jand g18674(.dina(n35936), .dinb(n35935), .dout(n35937));
  jor  g18675(.dina(n35937), .dinb(n35412), .dout(n35938));
  jxor g18676(.dina(n35406), .dinb(n326), .dout(n35939));
  jand g18677(.dina(n35939), .dinb(n35938), .dout(n35940));
  jor  g18678(.dina(n35940), .dinb(n35407), .dout(n35941));
  jxor g18679(.dina(n35401), .dinb(n277), .dout(n35942));
  jand g18680(.dina(n35942), .dinb(n35941), .dout(n35943));
  jor  g18681(.dina(n35943), .dinb(n35402), .dout(n35944));
  jxor g18682(.dina(n35396), .dinb(n278), .dout(n35945));
  jand g18683(.dina(n35945), .dinb(n35944), .dout(n35946));
  jor  g18684(.dina(n35946), .dinb(n35397), .dout(n35947));
  jxor g18685(.dina(n35391), .dinb(n279), .dout(n35948));
  jand g18686(.dina(n35948), .dinb(n35947), .dout(n35949));
  jor  g18687(.dina(n35949), .dinb(n35392), .dout(n35950));
  jxor g18688(.dina(n35386), .dinb(n280), .dout(n35951));
  jand g18689(.dina(n35951), .dinb(n35950), .dout(n35952));
  jor  g18690(.dina(n35952), .dinb(n35387), .dout(n35953));
  jxor g18691(.dina(n35381), .dinb(n283), .dout(n35954));
  jand g18692(.dina(n35954), .dinb(n35953), .dout(n35955));
  jor  g18693(.dina(n35955), .dinb(n35382), .dout(n35956));
  jxor g18694(.dina(n35376), .dinb(n315), .dout(n35957));
  jand g18695(.dina(n35957), .dinb(n35956), .dout(n35958));
  jor  g18696(.dina(n35958), .dinb(n35377), .dout(n35959));
  jxor g18697(.dina(n35371), .dinb(n316), .dout(n35960));
  jand g18698(.dina(n35960), .dinb(n35959), .dout(n35961));
  jor  g18699(.dina(n35961), .dinb(n35372), .dout(n35962));
  jxor g18700(.dina(n35366), .dinb(n317), .dout(n35963));
  jand g18701(.dina(n35963), .dinb(n35962), .dout(n35964));
  jor  g18702(.dina(n35964), .dinb(n35367), .dout(n35965));
  jxor g18703(.dina(n35361), .dinb(n284), .dout(n35966));
  jand g18704(.dina(n35966), .dinb(n35965), .dout(n35967));
  jor  g18705(.dina(n35967), .dinb(n35362), .dout(n35968));
  jxor g18706(.dina(n35356), .dinb(n285), .dout(n35969));
  jand g18707(.dina(n35969), .dinb(n35968), .dout(n35970));
  jor  g18708(.dina(n35970), .dinb(n35357), .dout(n35971));
  jxor g18709(.dina(n35351), .dinb(n286), .dout(n35972));
  jand g18710(.dina(n35972), .dinb(n35971), .dout(n35973));
  jor  g18711(.dina(n35973), .dinb(n35352), .dout(n35974));
  jxor g18712(.dina(n35346), .dinb(n287), .dout(n35975));
  jand g18713(.dina(n35975), .dinb(n35974), .dout(n35976));
  jor  g18714(.dina(n35976), .dinb(n35347), .dout(n35977));
  jxor g18715(.dina(n35341), .dinb(n288), .dout(n35978));
  jand g18716(.dina(n35978), .dinb(n35977), .dout(n35979));
  jor  g18717(.dina(n35979), .dinb(n35342), .dout(n35980));
  jxor g18718(.dina(n35336), .dinb(n289), .dout(n35981));
  jand g18719(.dina(n35981), .dinb(n35980), .dout(n35982));
  jor  g18720(.dina(n35982), .dinb(n35337), .dout(n35983));
  jxor g18721(.dina(n35331), .dinb(n290), .dout(n35984));
  jand g18722(.dina(n35984), .dinb(n35983), .dout(n35985));
  jor  g18723(.dina(n35985), .dinb(n35332), .dout(n35986));
  jxor g18724(.dina(n35326), .dinb(n291), .dout(n35987));
  jand g18725(.dina(n35987), .dinb(n35986), .dout(n35988));
  jor  g18726(.dina(n35988), .dinb(n35327), .dout(n35989));
  jxor g18727(.dina(n35321), .dinb(n292), .dout(n35990));
  jand g18728(.dina(n35990), .dinb(n35989), .dout(n35991));
  jor  g18729(.dina(n35991), .dinb(n35322), .dout(n35992));
  jxor g18730(.dina(n35316), .dinb(n293), .dout(n35993));
  jand g18731(.dina(n35993), .dinb(n35992), .dout(n35994));
  jor  g18732(.dina(n35994), .dinb(n35317), .dout(n35995));
  jxor g18733(.dina(n35311), .dinb(n294), .dout(n35996));
  jand g18734(.dina(n35996), .dinb(n35995), .dout(n35997));
  jor  g18735(.dina(n35997), .dinb(n35312), .dout(n35998));
  jand g18736(.dina(n35998), .dinb(n302), .dout(n35999));
  jand g18737(.dina(n35308), .dinb(n34853), .dout(n36000));
  jand g18738(.dina(n35303), .dinb(n34854), .dout(n36001));
  jand g18739(.dina(n36001), .dinb(n303), .dout(n36002));
  jor  g18740(.dina(n36002), .dinb(n36000), .dout(n36003));
  jand g18741(.dina(n36003), .dinb(n295), .dout(n36004));
  jand g18742(.dina(n34855), .dinb(b58 ), .dout(n36005));
  jor  g18743(.dina(n36005), .dinb(n36004), .dout(n36006));
  jnot g18744(.din(n36006), .dout(n36007));
  jand g18745(.dina(n36007), .dinb(n35999), .dout(n36008));
  jand g18746(.dina(n36004), .dinb(n302), .dout(n36009));
  jor  g18747(.dina(n36009), .dinb(n36008), .dout(n36010));
  jor  g18748(.dina(n36010), .dinb(n35311), .dout(n36011));
  jnot g18749(.din(n35312), .dout(n36012));
  jnot g18750(.din(n35317), .dout(n36013));
  jnot g18751(.din(n35322), .dout(n36014));
  jnot g18752(.din(n35327), .dout(n36015));
  jnot g18753(.din(n35332), .dout(n36016));
  jnot g18754(.din(n35337), .dout(n36017));
  jnot g18755(.din(n35342), .dout(n36018));
  jnot g18756(.din(n35347), .dout(n36019));
  jnot g18757(.din(n35352), .dout(n36020));
  jnot g18758(.din(n35357), .dout(n36021));
  jnot g18759(.din(n35362), .dout(n36022));
  jnot g18760(.din(n35367), .dout(n36023));
  jnot g18761(.din(n35372), .dout(n36024));
  jnot g18762(.din(n35377), .dout(n36025));
  jnot g18763(.din(n35382), .dout(n36026));
  jnot g18764(.din(n35387), .dout(n36027));
  jnot g18765(.din(n35392), .dout(n36028));
  jnot g18766(.din(n35397), .dout(n36029));
  jnot g18767(.din(n35402), .dout(n36030));
  jnot g18768(.din(n35407), .dout(n36031));
  jnot g18769(.din(n35412), .dout(n36032));
  jnot g18770(.din(n35417), .dout(n36033));
  jnot g18771(.din(n35422), .dout(n36034));
  jnot g18772(.din(n35427), .dout(n36035));
  jnot g18773(.din(n35432), .dout(n36036));
  jnot g18774(.din(n35437), .dout(n36037));
  jnot g18775(.din(n35442), .dout(n36038));
  jnot g18776(.din(n35447), .dout(n36039));
  jnot g18777(.din(n35452), .dout(n36040));
  jnot g18778(.din(n35457), .dout(n36041));
  jnot g18779(.din(n35462), .dout(n36042));
  jnot g18780(.din(n35467), .dout(n36043));
  jnot g18781(.din(n35472), .dout(n36044));
  jnot g18782(.din(n35477), .dout(n36045));
  jnot g18783(.din(n35482), .dout(n36046));
  jnot g18784(.din(n35487), .dout(n36047));
  jnot g18785(.din(n35492), .dout(n36048));
  jnot g18786(.din(n35497), .dout(n36049));
  jnot g18787(.din(n35502), .dout(n36050));
  jnot g18788(.din(n35507), .dout(n36051));
  jnot g18789(.din(n35512), .dout(n36052));
  jnot g18790(.din(n35517), .dout(n36053));
  jnot g18791(.din(n35522), .dout(n36054));
  jnot g18792(.din(n35527), .dout(n36055));
  jnot g18793(.din(n35532), .dout(n36056));
  jnot g18794(.din(n35537), .dout(n36057));
  jnot g18795(.din(n35542), .dout(n36058));
  jnot g18796(.din(n35547), .dout(n36059));
  jnot g18797(.din(n35552), .dout(n36060));
  jnot g18798(.din(n35557), .dout(n36061));
  jnot g18799(.din(n35562), .dout(n36062));
  jnot g18800(.din(n35567), .dout(n36063));
  jnot g18801(.din(n35572), .dout(n36064));
  jnot g18802(.din(n35577), .dout(n36065));
  jnot g18803(.din(n35582), .dout(n36066));
  jnot g18804(.din(n35589), .dout(n36067));
  jnot g18805(.din(n35824), .dout(n36068));
  jxor g18806(.dina(n35827), .dinb(n259), .dout(n36069));
  jor  g18807(.dina(n36069), .dinb(n15132), .dout(n36070));
  jand g18808(.dina(n36070), .dinb(n36068), .dout(n36071));
  jnot g18809(.din(n35831), .dout(n36072));
  jor  g18810(.dina(n36072), .dinb(n36071), .dout(n36073));
  jand g18811(.dina(n36073), .dinb(n36067), .dout(n36074));
  jnot g18812(.din(n35834), .dout(n36075));
  jor  g18813(.dina(n36075), .dinb(n36074), .dout(n36076));
  jand g18814(.dina(n36076), .dinb(n36066), .dout(n36077));
  jnot g18815(.din(n35837), .dout(n36078));
  jor  g18816(.dina(n36078), .dinb(n36077), .dout(n36079));
  jand g18817(.dina(n36079), .dinb(n36065), .dout(n36080));
  jnot g18818(.din(n35840), .dout(n36081));
  jor  g18819(.dina(n36081), .dinb(n36080), .dout(n36082));
  jand g18820(.dina(n36082), .dinb(n36064), .dout(n36083));
  jnot g18821(.din(n35843), .dout(n36084));
  jor  g18822(.dina(n36084), .dinb(n36083), .dout(n36085));
  jand g18823(.dina(n36085), .dinb(n36063), .dout(n36086));
  jnot g18824(.din(n35846), .dout(n36087));
  jor  g18825(.dina(n36087), .dinb(n36086), .dout(n36088));
  jand g18826(.dina(n36088), .dinb(n36062), .dout(n36089));
  jnot g18827(.din(n35849), .dout(n36090));
  jor  g18828(.dina(n36090), .dinb(n36089), .dout(n36091));
  jand g18829(.dina(n36091), .dinb(n36061), .dout(n36092));
  jnot g18830(.din(n35852), .dout(n36093));
  jor  g18831(.dina(n36093), .dinb(n36092), .dout(n36094));
  jand g18832(.dina(n36094), .dinb(n36060), .dout(n36095));
  jnot g18833(.din(n35855), .dout(n36096));
  jor  g18834(.dina(n36096), .dinb(n36095), .dout(n36097));
  jand g18835(.dina(n36097), .dinb(n36059), .dout(n36098));
  jnot g18836(.din(n35858), .dout(n36099));
  jor  g18837(.dina(n36099), .dinb(n36098), .dout(n36100));
  jand g18838(.dina(n36100), .dinb(n36058), .dout(n36101));
  jnot g18839(.din(n35861), .dout(n36102));
  jor  g18840(.dina(n36102), .dinb(n36101), .dout(n36103));
  jand g18841(.dina(n36103), .dinb(n36057), .dout(n36104));
  jnot g18842(.din(n35864), .dout(n36105));
  jor  g18843(.dina(n36105), .dinb(n36104), .dout(n36106));
  jand g18844(.dina(n36106), .dinb(n36056), .dout(n36107));
  jnot g18845(.din(n35867), .dout(n36108));
  jor  g18846(.dina(n36108), .dinb(n36107), .dout(n36109));
  jand g18847(.dina(n36109), .dinb(n36055), .dout(n36110));
  jnot g18848(.din(n35870), .dout(n36111));
  jor  g18849(.dina(n36111), .dinb(n36110), .dout(n36112));
  jand g18850(.dina(n36112), .dinb(n36054), .dout(n36113));
  jnot g18851(.din(n35873), .dout(n36114));
  jor  g18852(.dina(n36114), .dinb(n36113), .dout(n36115));
  jand g18853(.dina(n36115), .dinb(n36053), .dout(n36116));
  jnot g18854(.din(n35876), .dout(n36117));
  jor  g18855(.dina(n36117), .dinb(n36116), .dout(n36118));
  jand g18856(.dina(n36118), .dinb(n36052), .dout(n36119));
  jnot g18857(.din(n35879), .dout(n36120));
  jor  g18858(.dina(n36120), .dinb(n36119), .dout(n36121));
  jand g18859(.dina(n36121), .dinb(n36051), .dout(n36122));
  jnot g18860(.din(n35882), .dout(n36123));
  jor  g18861(.dina(n36123), .dinb(n36122), .dout(n36124));
  jand g18862(.dina(n36124), .dinb(n36050), .dout(n36125));
  jnot g18863(.din(n35885), .dout(n36126));
  jor  g18864(.dina(n36126), .dinb(n36125), .dout(n36127));
  jand g18865(.dina(n36127), .dinb(n36049), .dout(n36128));
  jnot g18866(.din(n35888), .dout(n36129));
  jor  g18867(.dina(n36129), .dinb(n36128), .dout(n36130));
  jand g18868(.dina(n36130), .dinb(n36048), .dout(n36131));
  jnot g18869(.din(n35891), .dout(n36132));
  jor  g18870(.dina(n36132), .dinb(n36131), .dout(n36133));
  jand g18871(.dina(n36133), .dinb(n36047), .dout(n36134));
  jnot g18872(.din(n35894), .dout(n36135));
  jor  g18873(.dina(n36135), .dinb(n36134), .dout(n36136));
  jand g18874(.dina(n36136), .dinb(n36046), .dout(n36137));
  jnot g18875(.din(n35897), .dout(n36138));
  jor  g18876(.dina(n36138), .dinb(n36137), .dout(n36139));
  jand g18877(.dina(n36139), .dinb(n36045), .dout(n36140));
  jnot g18878(.din(n35900), .dout(n36141));
  jor  g18879(.dina(n36141), .dinb(n36140), .dout(n36142));
  jand g18880(.dina(n36142), .dinb(n36044), .dout(n36143));
  jnot g18881(.din(n35903), .dout(n36144));
  jor  g18882(.dina(n36144), .dinb(n36143), .dout(n36145));
  jand g18883(.dina(n36145), .dinb(n36043), .dout(n36146));
  jnot g18884(.din(n35906), .dout(n36147));
  jor  g18885(.dina(n36147), .dinb(n36146), .dout(n36148));
  jand g18886(.dina(n36148), .dinb(n36042), .dout(n36149));
  jnot g18887(.din(n35909), .dout(n36150));
  jor  g18888(.dina(n36150), .dinb(n36149), .dout(n36151));
  jand g18889(.dina(n36151), .dinb(n36041), .dout(n36152));
  jnot g18890(.din(n35912), .dout(n36153));
  jor  g18891(.dina(n36153), .dinb(n36152), .dout(n36154));
  jand g18892(.dina(n36154), .dinb(n36040), .dout(n36155));
  jnot g18893(.din(n35915), .dout(n36156));
  jor  g18894(.dina(n36156), .dinb(n36155), .dout(n36157));
  jand g18895(.dina(n36157), .dinb(n36039), .dout(n36158));
  jnot g18896(.din(n35918), .dout(n36159));
  jor  g18897(.dina(n36159), .dinb(n36158), .dout(n36160));
  jand g18898(.dina(n36160), .dinb(n36038), .dout(n36161));
  jnot g18899(.din(n35921), .dout(n36162));
  jor  g18900(.dina(n36162), .dinb(n36161), .dout(n36163));
  jand g18901(.dina(n36163), .dinb(n36037), .dout(n36164));
  jnot g18902(.din(n35924), .dout(n36165));
  jor  g18903(.dina(n36165), .dinb(n36164), .dout(n36166));
  jand g18904(.dina(n36166), .dinb(n36036), .dout(n36167));
  jnot g18905(.din(n35927), .dout(n36168));
  jor  g18906(.dina(n36168), .dinb(n36167), .dout(n36169));
  jand g18907(.dina(n36169), .dinb(n36035), .dout(n36170));
  jnot g18908(.din(n35930), .dout(n36171));
  jor  g18909(.dina(n36171), .dinb(n36170), .dout(n36172));
  jand g18910(.dina(n36172), .dinb(n36034), .dout(n36173));
  jnot g18911(.din(n35933), .dout(n36174));
  jor  g18912(.dina(n36174), .dinb(n36173), .dout(n36175));
  jand g18913(.dina(n36175), .dinb(n36033), .dout(n36176));
  jnot g18914(.din(n35936), .dout(n36177));
  jor  g18915(.dina(n36177), .dinb(n36176), .dout(n36178));
  jand g18916(.dina(n36178), .dinb(n36032), .dout(n36179));
  jnot g18917(.din(n35939), .dout(n36180));
  jor  g18918(.dina(n36180), .dinb(n36179), .dout(n36181));
  jand g18919(.dina(n36181), .dinb(n36031), .dout(n36182));
  jnot g18920(.din(n35942), .dout(n36183));
  jor  g18921(.dina(n36183), .dinb(n36182), .dout(n36184));
  jand g18922(.dina(n36184), .dinb(n36030), .dout(n36185));
  jnot g18923(.din(n35945), .dout(n36186));
  jor  g18924(.dina(n36186), .dinb(n36185), .dout(n36187));
  jand g18925(.dina(n36187), .dinb(n36029), .dout(n36188));
  jnot g18926(.din(n35948), .dout(n36189));
  jor  g18927(.dina(n36189), .dinb(n36188), .dout(n36190));
  jand g18928(.dina(n36190), .dinb(n36028), .dout(n36191));
  jnot g18929(.din(n35951), .dout(n36192));
  jor  g18930(.dina(n36192), .dinb(n36191), .dout(n36193));
  jand g18931(.dina(n36193), .dinb(n36027), .dout(n36194));
  jnot g18932(.din(n35954), .dout(n36195));
  jor  g18933(.dina(n36195), .dinb(n36194), .dout(n36196));
  jand g18934(.dina(n36196), .dinb(n36026), .dout(n36197));
  jnot g18935(.din(n35957), .dout(n36198));
  jor  g18936(.dina(n36198), .dinb(n36197), .dout(n36199));
  jand g18937(.dina(n36199), .dinb(n36025), .dout(n36200));
  jnot g18938(.din(n35960), .dout(n36201));
  jor  g18939(.dina(n36201), .dinb(n36200), .dout(n36202));
  jand g18940(.dina(n36202), .dinb(n36024), .dout(n36203));
  jnot g18941(.din(n35963), .dout(n36204));
  jor  g18942(.dina(n36204), .dinb(n36203), .dout(n36205));
  jand g18943(.dina(n36205), .dinb(n36023), .dout(n36206));
  jnot g18944(.din(n35966), .dout(n36207));
  jor  g18945(.dina(n36207), .dinb(n36206), .dout(n36208));
  jand g18946(.dina(n36208), .dinb(n36022), .dout(n36209));
  jnot g18947(.din(n35969), .dout(n36210));
  jor  g18948(.dina(n36210), .dinb(n36209), .dout(n36211));
  jand g18949(.dina(n36211), .dinb(n36021), .dout(n36212));
  jnot g18950(.din(n35972), .dout(n36213));
  jor  g18951(.dina(n36213), .dinb(n36212), .dout(n36214));
  jand g18952(.dina(n36214), .dinb(n36020), .dout(n36215));
  jnot g18953(.din(n35975), .dout(n36216));
  jor  g18954(.dina(n36216), .dinb(n36215), .dout(n36217));
  jand g18955(.dina(n36217), .dinb(n36019), .dout(n36218));
  jnot g18956(.din(n35978), .dout(n36219));
  jor  g18957(.dina(n36219), .dinb(n36218), .dout(n36220));
  jand g18958(.dina(n36220), .dinb(n36018), .dout(n36221));
  jnot g18959(.din(n35981), .dout(n36222));
  jor  g18960(.dina(n36222), .dinb(n36221), .dout(n36223));
  jand g18961(.dina(n36223), .dinb(n36017), .dout(n36224));
  jnot g18962(.din(n35984), .dout(n36225));
  jor  g18963(.dina(n36225), .dinb(n36224), .dout(n36226));
  jand g18964(.dina(n36226), .dinb(n36016), .dout(n36227));
  jnot g18965(.din(n35987), .dout(n36228));
  jor  g18966(.dina(n36228), .dinb(n36227), .dout(n36229));
  jand g18967(.dina(n36229), .dinb(n36015), .dout(n36230));
  jnot g18968(.din(n35990), .dout(n36231));
  jor  g18969(.dina(n36231), .dinb(n36230), .dout(n36232));
  jand g18970(.dina(n36232), .dinb(n36014), .dout(n36233));
  jnot g18971(.din(n35993), .dout(n36234));
  jor  g18972(.dina(n36234), .dinb(n36233), .dout(n36235));
  jand g18973(.dina(n36235), .dinb(n36013), .dout(n36236));
  jnot g18974(.din(n35996), .dout(n36237));
  jor  g18975(.dina(n36237), .dinb(n36236), .dout(n36238));
  jand g18976(.dina(n36238), .dinb(n36012), .dout(n36239));
  jor  g18977(.dina(n36239), .dinb(n833), .dout(n36240));
  jor  g18978(.dina(n36006), .dinb(n36240), .dout(n36241));
  jnot g18979(.din(n36009), .dout(n36242));
  jand g18980(.dina(n36242), .dinb(n36241), .dout(n36243));
  jxor g18981(.dina(n35996), .dinb(n35995), .dout(n36244));
  jor  g18982(.dina(n36244), .dinb(n36243), .dout(n36245));
  jand g18983(.dina(n36245), .dinb(n36011), .dout(n36246));
  jand g18984(.dina(n35999), .dinb(n834), .dout(n36247));
  jnot g18985(.din(n36247), .dout(n36248));
  jand g18986(.dina(n36239), .dinb(n303), .dout(n36249));
  jnot g18987(.din(n36249), .dout(n36250));
  jand g18988(.dina(n36250), .dinb(n36003), .dout(n36251));
  jand g18989(.dina(n36251), .dinb(n36248), .dout(n36252));
  jand g18990(.dina(n36252), .dinb(n296), .dout(n36253));
  jand g18991(.dina(n36246), .dinb(n295), .dout(n36254));
  jor  g18992(.dina(n36010), .dinb(n35316), .dout(n36255));
  jxor g18993(.dina(n35993), .dinb(n35992), .dout(n36256));
  jor  g18994(.dina(n36256), .dinb(n36243), .dout(n36257));
  jand g18995(.dina(n36257), .dinb(n36255), .dout(n36258));
  jand g18996(.dina(n36258), .dinb(n294), .dout(n36259));
  jor  g18997(.dina(n36010), .dinb(n35321), .dout(n36260));
  jxor g18998(.dina(n35990), .dinb(n35989), .dout(n36261));
  jor  g18999(.dina(n36261), .dinb(n36243), .dout(n36262));
  jand g19000(.dina(n36262), .dinb(n36260), .dout(n36263));
  jand g19001(.dina(n36263), .dinb(n293), .dout(n36264));
  jor  g19002(.dina(n36010), .dinb(n35326), .dout(n36265));
  jxor g19003(.dina(n35987), .dinb(n35986), .dout(n36266));
  jor  g19004(.dina(n36266), .dinb(n36243), .dout(n36267));
  jand g19005(.dina(n36267), .dinb(n36265), .dout(n36268));
  jand g19006(.dina(n36268), .dinb(n292), .dout(n36269));
  jor  g19007(.dina(n36010), .dinb(n35331), .dout(n36270));
  jxor g19008(.dina(n35984), .dinb(n35983), .dout(n36271));
  jor  g19009(.dina(n36271), .dinb(n36243), .dout(n36272));
  jand g19010(.dina(n36272), .dinb(n36270), .dout(n36273));
  jand g19011(.dina(n36273), .dinb(n291), .dout(n36274));
  jor  g19012(.dina(n36010), .dinb(n35336), .dout(n36275));
  jxor g19013(.dina(n35981), .dinb(n35980), .dout(n36276));
  jor  g19014(.dina(n36276), .dinb(n36243), .dout(n36277));
  jand g19015(.dina(n36277), .dinb(n36275), .dout(n36278));
  jand g19016(.dina(n36278), .dinb(n290), .dout(n36279));
  jor  g19017(.dina(n36010), .dinb(n35341), .dout(n36280));
  jxor g19018(.dina(n35978), .dinb(n35977), .dout(n36281));
  jor  g19019(.dina(n36281), .dinb(n36243), .dout(n36282));
  jand g19020(.dina(n36282), .dinb(n36280), .dout(n36283));
  jand g19021(.dina(n36283), .dinb(n289), .dout(n36284));
  jor  g19022(.dina(n36010), .dinb(n35346), .dout(n36285));
  jxor g19023(.dina(n35975), .dinb(n35974), .dout(n36286));
  jor  g19024(.dina(n36286), .dinb(n36243), .dout(n36287));
  jand g19025(.dina(n36287), .dinb(n36285), .dout(n36288));
  jand g19026(.dina(n36288), .dinb(n288), .dout(n36289));
  jor  g19027(.dina(n36010), .dinb(n35351), .dout(n36290));
  jxor g19028(.dina(n35972), .dinb(n35971), .dout(n36291));
  jor  g19029(.dina(n36291), .dinb(n36243), .dout(n36292));
  jand g19030(.dina(n36292), .dinb(n36290), .dout(n36293));
  jand g19031(.dina(n36293), .dinb(n287), .dout(n36294));
  jor  g19032(.dina(n36010), .dinb(n35356), .dout(n36295));
  jxor g19033(.dina(n35969), .dinb(n35968), .dout(n36296));
  jor  g19034(.dina(n36296), .dinb(n36243), .dout(n36297));
  jand g19035(.dina(n36297), .dinb(n36295), .dout(n36298));
  jand g19036(.dina(n36298), .dinb(n286), .dout(n36299));
  jor  g19037(.dina(n36010), .dinb(n35361), .dout(n36300));
  jxor g19038(.dina(n35966), .dinb(n35965), .dout(n36301));
  jor  g19039(.dina(n36301), .dinb(n36243), .dout(n36302));
  jand g19040(.dina(n36302), .dinb(n36300), .dout(n36303));
  jand g19041(.dina(n36303), .dinb(n285), .dout(n36304));
  jor  g19042(.dina(n36010), .dinb(n35366), .dout(n36305));
  jxor g19043(.dina(n35963), .dinb(n35962), .dout(n36306));
  jor  g19044(.dina(n36306), .dinb(n36243), .dout(n36307));
  jand g19045(.dina(n36307), .dinb(n36305), .dout(n36308));
  jand g19046(.dina(n36308), .dinb(n284), .dout(n36309));
  jor  g19047(.dina(n36010), .dinb(n35371), .dout(n36310));
  jxor g19048(.dina(n35960), .dinb(n35959), .dout(n36311));
  jor  g19049(.dina(n36311), .dinb(n36243), .dout(n36312));
  jand g19050(.dina(n36312), .dinb(n36310), .dout(n36313));
  jand g19051(.dina(n36313), .dinb(n317), .dout(n36314));
  jor  g19052(.dina(n36010), .dinb(n35376), .dout(n36315));
  jxor g19053(.dina(n35957), .dinb(n35956), .dout(n36316));
  jor  g19054(.dina(n36316), .dinb(n36243), .dout(n36317));
  jand g19055(.dina(n36317), .dinb(n36315), .dout(n36318));
  jand g19056(.dina(n36318), .dinb(n316), .dout(n36319));
  jor  g19057(.dina(n36010), .dinb(n35381), .dout(n36320));
  jxor g19058(.dina(n35954), .dinb(n35953), .dout(n36321));
  jor  g19059(.dina(n36321), .dinb(n36243), .dout(n36322));
  jand g19060(.dina(n36322), .dinb(n36320), .dout(n36323));
  jand g19061(.dina(n36323), .dinb(n315), .dout(n36324));
  jor  g19062(.dina(n36010), .dinb(n35386), .dout(n36325));
  jxor g19063(.dina(n35951), .dinb(n35950), .dout(n36326));
  jor  g19064(.dina(n36326), .dinb(n36243), .dout(n36327));
  jand g19065(.dina(n36327), .dinb(n36325), .dout(n36328));
  jand g19066(.dina(n36328), .dinb(n283), .dout(n36329));
  jor  g19067(.dina(n36010), .dinb(n35391), .dout(n36330));
  jxor g19068(.dina(n35948), .dinb(n35947), .dout(n36331));
  jor  g19069(.dina(n36331), .dinb(n36243), .dout(n36332));
  jand g19070(.dina(n36332), .dinb(n36330), .dout(n36333));
  jand g19071(.dina(n36333), .dinb(n280), .dout(n36334));
  jor  g19072(.dina(n36010), .dinb(n35396), .dout(n36335));
  jxor g19073(.dina(n35945), .dinb(n35944), .dout(n36336));
  jor  g19074(.dina(n36336), .dinb(n36243), .dout(n36337));
  jand g19075(.dina(n36337), .dinb(n36335), .dout(n36338));
  jand g19076(.dina(n36338), .dinb(n279), .dout(n36339));
  jor  g19077(.dina(n36010), .dinb(n35401), .dout(n36340));
  jxor g19078(.dina(n35942), .dinb(n35941), .dout(n36341));
  jor  g19079(.dina(n36341), .dinb(n36243), .dout(n36342));
  jand g19080(.dina(n36342), .dinb(n36340), .dout(n36343));
  jand g19081(.dina(n36343), .dinb(n278), .dout(n36344));
  jor  g19082(.dina(n36010), .dinb(n35406), .dout(n36345));
  jxor g19083(.dina(n35939), .dinb(n35938), .dout(n36346));
  jor  g19084(.dina(n36346), .dinb(n36243), .dout(n36347));
  jand g19085(.dina(n36347), .dinb(n36345), .dout(n36348));
  jand g19086(.dina(n36348), .dinb(n277), .dout(n36349));
  jor  g19087(.dina(n36010), .dinb(n35411), .dout(n36350));
  jxor g19088(.dina(n35936), .dinb(n35935), .dout(n36351));
  jor  g19089(.dina(n36351), .dinb(n36243), .dout(n36352));
  jand g19090(.dina(n36352), .dinb(n36350), .dout(n36353));
  jand g19091(.dina(n36353), .dinb(n326), .dout(n36354));
  jor  g19092(.dina(n36010), .dinb(n35416), .dout(n36355));
  jxor g19093(.dina(n35933), .dinb(n35932), .dout(n36356));
  jor  g19094(.dina(n36356), .dinb(n36243), .dout(n36357));
  jand g19095(.dina(n36357), .dinb(n36355), .dout(n36358));
  jand g19096(.dina(n36358), .dinb(n325), .dout(n36359));
  jor  g19097(.dina(n36010), .dinb(n35421), .dout(n36360));
  jxor g19098(.dina(n35930), .dinb(n35929), .dout(n36361));
  jor  g19099(.dina(n36361), .dinb(n36243), .dout(n36362));
  jand g19100(.dina(n36362), .dinb(n36360), .dout(n36363));
  jand g19101(.dina(n36363), .dinb(n324), .dout(n36364));
  jor  g19102(.dina(n36010), .dinb(n35426), .dout(n36365));
  jxor g19103(.dina(n35927), .dinb(n35926), .dout(n36366));
  jor  g19104(.dina(n36366), .dinb(n36243), .dout(n36367));
  jand g19105(.dina(n36367), .dinb(n36365), .dout(n36368));
  jand g19106(.dina(n36368), .dinb(n276), .dout(n36369));
  jor  g19107(.dina(n36010), .dinb(n35431), .dout(n36370));
  jxor g19108(.dina(n35924), .dinb(n35923), .dout(n36371));
  jor  g19109(.dina(n36371), .dinb(n36243), .dout(n36372));
  jand g19110(.dina(n36372), .dinb(n36370), .dout(n36373));
  jand g19111(.dina(n36373), .dinb(n333), .dout(n36374));
  jor  g19112(.dina(n36010), .dinb(n35436), .dout(n36375));
  jxor g19113(.dina(n35921), .dinb(n35920), .dout(n36376));
  jor  g19114(.dina(n36376), .dinb(n36243), .dout(n36377));
  jand g19115(.dina(n36377), .dinb(n36375), .dout(n36378));
  jand g19116(.dina(n36378), .dinb(n332), .dout(n36379));
  jor  g19117(.dina(n36010), .dinb(n35441), .dout(n36380));
  jxor g19118(.dina(n35918), .dinb(n35917), .dout(n36381));
  jor  g19119(.dina(n36381), .dinb(n36243), .dout(n36382));
  jand g19120(.dina(n36382), .dinb(n36380), .dout(n36383));
  jand g19121(.dina(n36383), .dinb(n331), .dout(n36384));
  jor  g19122(.dina(n36010), .dinb(n35446), .dout(n36385));
  jxor g19123(.dina(n35915), .dinb(n35914), .dout(n36386));
  jor  g19124(.dina(n36386), .dinb(n36243), .dout(n36387));
  jand g19125(.dina(n36387), .dinb(n36385), .dout(n36388));
  jand g19126(.dina(n36388), .dinb(n275), .dout(n36389));
  jor  g19127(.dina(n36010), .dinb(n35451), .dout(n36390));
  jxor g19128(.dina(n35912), .dinb(n35911), .dout(n36391));
  jor  g19129(.dina(n36391), .dinb(n36243), .dout(n36392));
  jand g19130(.dina(n36392), .dinb(n36390), .dout(n36393));
  jand g19131(.dina(n36393), .dinb(n340), .dout(n36394));
  jor  g19132(.dina(n36010), .dinb(n35456), .dout(n36395));
  jxor g19133(.dina(n35909), .dinb(n35908), .dout(n36396));
  jor  g19134(.dina(n36396), .dinb(n36243), .dout(n36397));
  jand g19135(.dina(n36397), .dinb(n36395), .dout(n36398));
  jand g19136(.dina(n36398), .dinb(n339), .dout(n36399));
  jor  g19137(.dina(n36010), .dinb(n35461), .dout(n36400));
  jxor g19138(.dina(n35906), .dinb(n35905), .dout(n36401));
  jor  g19139(.dina(n36401), .dinb(n36243), .dout(n36402));
  jand g19140(.dina(n36402), .dinb(n36400), .dout(n36403));
  jand g19141(.dina(n36403), .dinb(n338), .dout(n36404));
  jor  g19142(.dina(n36010), .dinb(n35466), .dout(n36405));
  jxor g19143(.dina(n35903), .dinb(n35902), .dout(n36406));
  jor  g19144(.dina(n36406), .dinb(n36243), .dout(n36407));
  jand g19145(.dina(n36407), .dinb(n36405), .dout(n36408));
  jand g19146(.dina(n36408), .dinb(n271), .dout(n36409));
  jor  g19147(.dina(n36010), .dinb(n35471), .dout(n36410));
  jxor g19148(.dina(n35900), .dinb(n35899), .dout(n36411));
  jor  g19149(.dina(n36411), .dinb(n36243), .dout(n36412));
  jand g19150(.dina(n36412), .dinb(n36410), .dout(n36413));
  jand g19151(.dina(n36413), .dinb(n270), .dout(n36414));
  jor  g19152(.dina(n36010), .dinb(n35476), .dout(n36415));
  jxor g19153(.dina(n35897), .dinb(n35896), .dout(n36416));
  jor  g19154(.dina(n36416), .dinb(n36243), .dout(n36417));
  jand g19155(.dina(n36417), .dinb(n36415), .dout(n36418));
  jand g19156(.dina(n36418), .dinb(n269), .dout(n36419));
  jor  g19157(.dina(n36010), .dinb(n35481), .dout(n36420));
  jxor g19158(.dina(n35894), .dinb(n35893), .dout(n36421));
  jor  g19159(.dina(n36421), .dinb(n36243), .dout(n36422));
  jand g19160(.dina(n36422), .dinb(n36420), .dout(n36423));
  jand g19161(.dina(n36423), .dinb(n274), .dout(n36424));
  jor  g19162(.dina(n36010), .dinb(n35486), .dout(n36425));
  jxor g19163(.dina(n35891), .dinb(n35890), .dout(n36426));
  jor  g19164(.dina(n36426), .dinb(n36243), .dout(n36427));
  jand g19165(.dina(n36427), .dinb(n36425), .dout(n36428));
  jand g19166(.dina(n36428), .dinb(n268), .dout(n36429));
  jor  g19167(.dina(n36010), .dinb(n35491), .dout(n36430));
  jxor g19168(.dina(n35888), .dinb(n35887), .dout(n36431));
  jor  g19169(.dina(n36431), .dinb(n36243), .dout(n36432));
  jand g19170(.dina(n36432), .dinb(n36430), .dout(n36433));
  jand g19171(.dina(n36433), .dinb(n349), .dout(n36434));
  jor  g19172(.dina(n36010), .dinb(n35496), .dout(n36435));
  jxor g19173(.dina(n35885), .dinb(n35884), .dout(n36436));
  jor  g19174(.dina(n36436), .dinb(n36243), .dout(n36437));
  jand g19175(.dina(n36437), .dinb(n36435), .dout(n36438));
  jand g19176(.dina(n36438), .dinb(n348), .dout(n36439));
  jor  g19177(.dina(n36010), .dinb(n35501), .dout(n36440));
  jxor g19178(.dina(n35882), .dinb(n35881), .dout(n36441));
  jor  g19179(.dina(n36441), .dinb(n36243), .dout(n36442));
  jand g19180(.dina(n36442), .dinb(n36440), .dout(n36443));
  jand g19181(.dina(n36443), .dinb(n347), .dout(n36444));
  jor  g19182(.dina(n36010), .dinb(n35506), .dout(n36445));
  jxor g19183(.dina(n35879), .dinb(n35878), .dout(n36446));
  jor  g19184(.dina(n36446), .dinb(n36243), .dout(n36447));
  jand g19185(.dina(n36447), .dinb(n36445), .dout(n36448));
  jand g19186(.dina(n36448), .dinb(n267), .dout(n36449));
  jor  g19187(.dina(n36010), .dinb(n35511), .dout(n36450));
  jxor g19188(.dina(n35876), .dinb(n35875), .dout(n36451));
  jor  g19189(.dina(n36451), .dinb(n36243), .dout(n36452));
  jand g19190(.dina(n36452), .dinb(n36450), .dout(n36453));
  jand g19191(.dina(n36453), .dinb(n266), .dout(n36454));
  jor  g19192(.dina(n36010), .dinb(n35516), .dout(n36455));
  jxor g19193(.dina(n35873), .dinb(n35872), .dout(n36456));
  jor  g19194(.dina(n36456), .dinb(n36243), .dout(n36457));
  jand g19195(.dina(n36457), .dinb(n36455), .dout(n36458));
  jand g19196(.dina(n36458), .dinb(n356), .dout(n36459));
  jor  g19197(.dina(n36010), .dinb(n35521), .dout(n36460));
  jxor g19198(.dina(n35870), .dinb(n35869), .dout(n36461));
  jor  g19199(.dina(n36461), .dinb(n36243), .dout(n36462));
  jand g19200(.dina(n36462), .dinb(n36460), .dout(n36463));
  jand g19201(.dina(n36463), .dinb(n355), .dout(n36464));
  jor  g19202(.dina(n36010), .dinb(n35526), .dout(n36465));
  jxor g19203(.dina(n35867), .dinb(n35866), .dout(n36466));
  jor  g19204(.dina(n36466), .dinb(n36243), .dout(n36467));
  jand g19205(.dina(n36467), .dinb(n36465), .dout(n36468));
  jand g19206(.dina(n36468), .dinb(n364), .dout(n36469));
  jor  g19207(.dina(n36010), .dinb(n35531), .dout(n36470));
  jxor g19208(.dina(n35864), .dinb(n35863), .dout(n36471));
  jor  g19209(.dina(n36471), .dinb(n36243), .dout(n36472));
  jand g19210(.dina(n36472), .dinb(n36470), .dout(n36473));
  jand g19211(.dina(n36473), .dinb(n361), .dout(n36474));
  jor  g19212(.dina(n36010), .dinb(n35536), .dout(n36475));
  jxor g19213(.dina(n35861), .dinb(n35860), .dout(n36476));
  jor  g19214(.dina(n36476), .dinb(n36243), .dout(n36477));
  jand g19215(.dina(n36477), .dinb(n36475), .dout(n36478));
  jand g19216(.dina(n36478), .dinb(n360), .dout(n36479));
  jor  g19217(.dina(n36010), .dinb(n35541), .dout(n36480));
  jxor g19218(.dina(n35858), .dinb(n35857), .dout(n36481));
  jor  g19219(.dina(n36481), .dinb(n36243), .dout(n36482));
  jand g19220(.dina(n36482), .dinb(n36480), .dout(n36483));
  jand g19221(.dina(n36483), .dinb(n363), .dout(n36484));
  jor  g19222(.dina(n36010), .dinb(n35546), .dout(n36485));
  jxor g19223(.dina(n35855), .dinb(n35854), .dout(n36486));
  jor  g19224(.dina(n36486), .dinb(n36243), .dout(n36487));
  jand g19225(.dina(n36487), .dinb(n36485), .dout(n36488));
  jand g19226(.dina(n36488), .dinb(n359), .dout(n36489));
  jor  g19227(.dina(n36010), .dinb(n35551), .dout(n36490));
  jxor g19228(.dina(n35852), .dinb(n35851), .dout(n36491));
  jor  g19229(.dina(n36491), .dinb(n36243), .dout(n36492));
  jand g19230(.dina(n36492), .dinb(n36490), .dout(n36493));
  jand g19231(.dina(n36493), .dinb(n369), .dout(n36494));
  jor  g19232(.dina(n36010), .dinb(n35556), .dout(n36495));
  jxor g19233(.dina(n35849), .dinb(n35848), .dout(n36496));
  jor  g19234(.dina(n36496), .dinb(n36243), .dout(n36497));
  jand g19235(.dina(n36497), .dinb(n36495), .dout(n36498));
  jand g19236(.dina(n36498), .dinb(n368), .dout(n36499));
  jor  g19237(.dina(n36010), .dinb(n35561), .dout(n36500));
  jxor g19238(.dina(n35846), .dinb(n35845), .dout(n36501));
  jor  g19239(.dina(n36501), .dinb(n36243), .dout(n36502));
  jand g19240(.dina(n36502), .dinb(n36500), .dout(n36503));
  jand g19241(.dina(n36503), .dinb(n367), .dout(n36504));
  jor  g19242(.dina(n36010), .dinb(n35566), .dout(n36505));
  jxor g19243(.dina(n35843), .dinb(n35842), .dout(n36506));
  jor  g19244(.dina(n36506), .dinb(n36243), .dout(n36507));
  jand g19245(.dina(n36507), .dinb(n36505), .dout(n36508));
  jand g19246(.dina(n36508), .dinb(n265), .dout(n36509));
  jor  g19247(.dina(n36010), .dinb(n35571), .dout(n36510));
  jxor g19248(.dina(n35840), .dinb(n35839), .dout(n36511));
  jor  g19249(.dina(n36511), .dinb(n36243), .dout(n36512));
  jand g19250(.dina(n36512), .dinb(n36510), .dout(n36513));
  jand g19251(.dina(n36513), .dinb(n378), .dout(n36514));
  jor  g19252(.dina(n36010), .dinb(n35576), .dout(n36515));
  jxor g19253(.dina(n35837), .dinb(n35836), .dout(n36516));
  jor  g19254(.dina(n36516), .dinb(n36243), .dout(n36517));
  jand g19255(.dina(n36517), .dinb(n36515), .dout(n36518));
  jand g19256(.dina(n36518), .dinb(n377), .dout(n36519));
  jor  g19257(.dina(n36010), .dinb(n35581), .dout(n36520));
  jxor g19258(.dina(n35834), .dinb(n35833), .dout(n36521));
  jor  g19259(.dina(n36521), .dinb(n36243), .dout(n36522));
  jand g19260(.dina(n36522), .dinb(n36520), .dout(n36523));
  jand g19261(.dina(n36523), .dinb(n376), .dout(n36524));
  jor  g19262(.dina(n36010), .dinb(n35588), .dout(n36525));
  jxor g19263(.dina(n35831), .dinb(n35830), .dout(n36526));
  jor  g19264(.dina(n36526), .dinb(n36243), .dout(n36527));
  jand g19265(.dina(n36527), .dinb(n36525), .dout(n36528));
  jand g19266(.dina(n36528), .dinb(n264), .dout(n36529));
  jand g19267(.dina(n36069), .dinb(n15132), .dout(n36530));
  jor  g19268(.dina(n36243), .dinb(n35829), .dout(n36531));
  jor  g19269(.dina(n36531), .dinb(n36530), .dout(n36532));
  jand g19270(.dina(n36243), .dinb(n35823), .dout(n36533));
  jnot g19271(.din(n36533), .dout(n36534));
  jand g19272(.dina(n36534), .dinb(n36532), .dout(n36535));
  jnot g19273(.din(n36535), .dout(n36536));
  jand g19274(.dina(n36536), .dinb(n386), .dout(n36537));
  jand g19275(.dina(n36010), .dinb(b0 ), .dout(n36538));
  jxor g19276(.dina(n36538), .dinb(a5 ), .dout(n36539));
  jand g19277(.dina(n36539), .dinb(n259), .dout(n36540));
  jxor g19278(.dina(n36538), .dinb(n15131), .dout(n36541));
  jxor g19279(.dina(n36541), .dinb(b1 ), .dout(n36542));
  jand g19280(.dina(n36542), .dinb(n15614), .dout(n36543));
  jor  g19281(.dina(n36543), .dinb(n36540), .dout(n36544));
  jxor g19282(.dina(n36535), .dinb(b2 ), .dout(n36545));
  jand g19283(.dina(n36545), .dinb(n36544), .dout(n36546));
  jor  g19284(.dina(n36546), .dinb(n36537), .dout(n36547));
  jxor g19285(.dina(n36528), .dinb(n264), .dout(n36548));
  jand g19286(.dina(n36548), .dinb(n36547), .dout(n36549));
  jor  g19287(.dina(n36549), .dinb(n36529), .dout(n36550));
  jxor g19288(.dina(n36523), .dinb(n376), .dout(n36551));
  jand g19289(.dina(n36551), .dinb(n36550), .dout(n36552));
  jor  g19290(.dina(n36552), .dinb(n36524), .dout(n36553));
  jxor g19291(.dina(n36518), .dinb(n377), .dout(n36554));
  jand g19292(.dina(n36554), .dinb(n36553), .dout(n36555));
  jor  g19293(.dina(n36555), .dinb(n36519), .dout(n36556));
  jxor g19294(.dina(n36513), .dinb(n378), .dout(n36557));
  jand g19295(.dina(n36557), .dinb(n36556), .dout(n36558));
  jor  g19296(.dina(n36558), .dinb(n36514), .dout(n36559));
  jxor g19297(.dina(n36508), .dinb(n265), .dout(n36560));
  jand g19298(.dina(n36560), .dinb(n36559), .dout(n36561));
  jor  g19299(.dina(n36561), .dinb(n36509), .dout(n36562));
  jxor g19300(.dina(n36503), .dinb(n367), .dout(n36563));
  jand g19301(.dina(n36563), .dinb(n36562), .dout(n36564));
  jor  g19302(.dina(n36564), .dinb(n36504), .dout(n36565));
  jxor g19303(.dina(n36498), .dinb(n368), .dout(n36566));
  jand g19304(.dina(n36566), .dinb(n36565), .dout(n36567));
  jor  g19305(.dina(n36567), .dinb(n36499), .dout(n36568));
  jxor g19306(.dina(n36493), .dinb(n369), .dout(n36569));
  jand g19307(.dina(n36569), .dinb(n36568), .dout(n36570));
  jor  g19308(.dina(n36570), .dinb(n36494), .dout(n36571));
  jxor g19309(.dina(n36488), .dinb(n359), .dout(n36572));
  jand g19310(.dina(n36572), .dinb(n36571), .dout(n36573));
  jor  g19311(.dina(n36573), .dinb(n36489), .dout(n36574));
  jxor g19312(.dina(n36483), .dinb(n363), .dout(n36575));
  jand g19313(.dina(n36575), .dinb(n36574), .dout(n36576));
  jor  g19314(.dina(n36576), .dinb(n36484), .dout(n36577));
  jxor g19315(.dina(n36478), .dinb(n360), .dout(n36578));
  jand g19316(.dina(n36578), .dinb(n36577), .dout(n36579));
  jor  g19317(.dina(n36579), .dinb(n36479), .dout(n36580));
  jxor g19318(.dina(n36473), .dinb(n361), .dout(n36581));
  jand g19319(.dina(n36581), .dinb(n36580), .dout(n36582));
  jor  g19320(.dina(n36582), .dinb(n36474), .dout(n36583));
  jxor g19321(.dina(n36468), .dinb(n364), .dout(n36584));
  jand g19322(.dina(n36584), .dinb(n36583), .dout(n36585));
  jor  g19323(.dina(n36585), .dinb(n36469), .dout(n36586));
  jxor g19324(.dina(n36463), .dinb(n355), .dout(n36587));
  jand g19325(.dina(n36587), .dinb(n36586), .dout(n36588));
  jor  g19326(.dina(n36588), .dinb(n36464), .dout(n36589));
  jxor g19327(.dina(n36458), .dinb(n356), .dout(n36590));
  jand g19328(.dina(n36590), .dinb(n36589), .dout(n36591));
  jor  g19329(.dina(n36591), .dinb(n36459), .dout(n36592));
  jxor g19330(.dina(n36453), .dinb(n266), .dout(n36593));
  jand g19331(.dina(n36593), .dinb(n36592), .dout(n36594));
  jor  g19332(.dina(n36594), .dinb(n36454), .dout(n36595));
  jxor g19333(.dina(n36448), .dinb(n267), .dout(n36596));
  jand g19334(.dina(n36596), .dinb(n36595), .dout(n36597));
  jor  g19335(.dina(n36597), .dinb(n36449), .dout(n36598));
  jxor g19336(.dina(n36443), .dinb(n347), .dout(n36599));
  jand g19337(.dina(n36599), .dinb(n36598), .dout(n36600));
  jor  g19338(.dina(n36600), .dinb(n36444), .dout(n36601));
  jxor g19339(.dina(n36438), .dinb(n348), .dout(n36602));
  jand g19340(.dina(n36602), .dinb(n36601), .dout(n36603));
  jor  g19341(.dina(n36603), .dinb(n36439), .dout(n36604));
  jxor g19342(.dina(n36433), .dinb(n349), .dout(n36605));
  jand g19343(.dina(n36605), .dinb(n36604), .dout(n36606));
  jor  g19344(.dina(n36606), .dinb(n36434), .dout(n36607));
  jxor g19345(.dina(n36428), .dinb(n268), .dout(n36608));
  jand g19346(.dina(n36608), .dinb(n36607), .dout(n36609));
  jor  g19347(.dina(n36609), .dinb(n36429), .dout(n36610));
  jxor g19348(.dina(n36423), .dinb(n274), .dout(n36611));
  jand g19349(.dina(n36611), .dinb(n36610), .dout(n36612));
  jor  g19350(.dina(n36612), .dinb(n36424), .dout(n36613));
  jxor g19351(.dina(n36418), .dinb(n269), .dout(n36614));
  jand g19352(.dina(n36614), .dinb(n36613), .dout(n36615));
  jor  g19353(.dina(n36615), .dinb(n36419), .dout(n36616));
  jxor g19354(.dina(n36413), .dinb(n270), .dout(n36617));
  jand g19355(.dina(n36617), .dinb(n36616), .dout(n36618));
  jor  g19356(.dina(n36618), .dinb(n36414), .dout(n36619));
  jxor g19357(.dina(n36408), .dinb(n271), .dout(n36620));
  jand g19358(.dina(n36620), .dinb(n36619), .dout(n36621));
  jor  g19359(.dina(n36621), .dinb(n36409), .dout(n36622));
  jxor g19360(.dina(n36403), .dinb(n338), .dout(n36623));
  jand g19361(.dina(n36623), .dinb(n36622), .dout(n36624));
  jor  g19362(.dina(n36624), .dinb(n36404), .dout(n36625));
  jxor g19363(.dina(n36398), .dinb(n339), .dout(n36626));
  jand g19364(.dina(n36626), .dinb(n36625), .dout(n36627));
  jor  g19365(.dina(n36627), .dinb(n36399), .dout(n36628));
  jxor g19366(.dina(n36393), .dinb(n340), .dout(n36629));
  jand g19367(.dina(n36629), .dinb(n36628), .dout(n36630));
  jor  g19368(.dina(n36630), .dinb(n36394), .dout(n36631));
  jxor g19369(.dina(n36388), .dinb(n275), .dout(n36632));
  jand g19370(.dina(n36632), .dinb(n36631), .dout(n36633));
  jor  g19371(.dina(n36633), .dinb(n36389), .dout(n36634));
  jxor g19372(.dina(n36383), .dinb(n331), .dout(n36635));
  jand g19373(.dina(n36635), .dinb(n36634), .dout(n36636));
  jor  g19374(.dina(n36636), .dinb(n36384), .dout(n36637));
  jxor g19375(.dina(n36378), .dinb(n332), .dout(n36638));
  jand g19376(.dina(n36638), .dinb(n36637), .dout(n36639));
  jor  g19377(.dina(n36639), .dinb(n36379), .dout(n36640));
  jxor g19378(.dina(n36373), .dinb(n333), .dout(n36641));
  jand g19379(.dina(n36641), .dinb(n36640), .dout(n36642));
  jor  g19380(.dina(n36642), .dinb(n36374), .dout(n36643));
  jxor g19381(.dina(n36368), .dinb(n276), .dout(n36644));
  jand g19382(.dina(n36644), .dinb(n36643), .dout(n36645));
  jor  g19383(.dina(n36645), .dinb(n36369), .dout(n36646));
  jxor g19384(.dina(n36363), .dinb(n324), .dout(n36647));
  jand g19385(.dina(n36647), .dinb(n36646), .dout(n36648));
  jor  g19386(.dina(n36648), .dinb(n36364), .dout(n36649));
  jxor g19387(.dina(n36358), .dinb(n325), .dout(n36650));
  jand g19388(.dina(n36650), .dinb(n36649), .dout(n36651));
  jor  g19389(.dina(n36651), .dinb(n36359), .dout(n36652));
  jxor g19390(.dina(n36353), .dinb(n326), .dout(n36653));
  jand g19391(.dina(n36653), .dinb(n36652), .dout(n36654));
  jor  g19392(.dina(n36654), .dinb(n36354), .dout(n36655));
  jxor g19393(.dina(n36348), .dinb(n277), .dout(n36656));
  jand g19394(.dina(n36656), .dinb(n36655), .dout(n36657));
  jor  g19395(.dina(n36657), .dinb(n36349), .dout(n36658));
  jxor g19396(.dina(n36343), .dinb(n278), .dout(n36659));
  jand g19397(.dina(n36659), .dinb(n36658), .dout(n36660));
  jor  g19398(.dina(n36660), .dinb(n36344), .dout(n36661));
  jxor g19399(.dina(n36338), .dinb(n279), .dout(n36662));
  jand g19400(.dina(n36662), .dinb(n36661), .dout(n36663));
  jor  g19401(.dina(n36663), .dinb(n36339), .dout(n36664));
  jxor g19402(.dina(n36333), .dinb(n280), .dout(n36665));
  jand g19403(.dina(n36665), .dinb(n36664), .dout(n36666));
  jor  g19404(.dina(n36666), .dinb(n36334), .dout(n36667));
  jxor g19405(.dina(n36328), .dinb(n283), .dout(n36668));
  jand g19406(.dina(n36668), .dinb(n36667), .dout(n36669));
  jor  g19407(.dina(n36669), .dinb(n36329), .dout(n36670));
  jxor g19408(.dina(n36323), .dinb(n315), .dout(n36671));
  jand g19409(.dina(n36671), .dinb(n36670), .dout(n36672));
  jor  g19410(.dina(n36672), .dinb(n36324), .dout(n36673));
  jxor g19411(.dina(n36318), .dinb(n316), .dout(n36674));
  jand g19412(.dina(n36674), .dinb(n36673), .dout(n36675));
  jor  g19413(.dina(n36675), .dinb(n36319), .dout(n36676));
  jxor g19414(.dina(n36313), .dinb(n317), .dout(n36677));
  jand g19415(.dina(n36677), .dinb(n36676), .dout(n36678));
  jor  g19416(.dina(n36678), .dinb(n36314), .dout(n36679));
  jxor g19417(.dina(n36308), .dinb(n284), .dout(n36680));
  jand g19418(.dina(n36680), .dinb(n36679), .dout(n36681));
  jor  g19419(.dina(n36681), .dinb(n36309), .dout(n36682));
  jxor g19420(.dina(n36303), .dinb(n285), .dout(n36683));
  jand g19421(.dina(n36683), .dinb(n36682), .dout(n36684));
  jor  g19422(.dina(n36684), .dinb(n36304), .dout(n36685));
  jxor g19423(.dina(n36298), .dinb(n286), .dout(n36686));
  jand g19424(.dina(n36686), .dinb(n36685), .dout(n36687));
  jor  g19425(.dina(n36687), .dinb(n36299), .dout(n36688));
  jxor g19426(.dina(n36293), .dinb(n287), .dout(n36689));
  jand g19427(.dina(n36689), .dinb(n36688), .dout(n36690));
  jor  g19428(.dina(n36690), .dinb(n36294), .dout(n36691));
  jxor g19429(.dina(n36288), .dinb(n288), .dout(n36692));
  jand g19430(.dina(n36692), .dinb(n36691), .dout(n36693));
  jor  g19431(.dina(n36693), .dinb(n36289), .dout(n36694));
  jxor g19432(.dina(n36283), .dinb(n289), .dout(n36695));
  jand g19433(.dina(n36695), .dinb(n36694), .dout(n36696));
  jor  g19434(.dina(n36696), .dinb(n36284), .dout(n36697));
  jxor g19435(.dina(n36278), .dinb(n290), .dout(n36698));
  jand g19436(.dina(n36698), .dinb(n36697), .dout(n36699));
  jor  g19437(.dina(n36699), .dinb(n36279), .dout(n36700));
  jxor g19438(.dina(n36273), .dinb(n291), .dout(n36701));
  jand g19439(.dina(n36701), .dinb(n36700), .dout(n36702));
  jor  g19440(.dina(n36702), .dinb(n36274), .dout(n36703));
  jxor g19441(.dina(n36268), .dinb(n292), .dout(n36704));
  jand g19442(.dina(n36704), .dinb(n36703), .dout(n36705));
  jor  g19443(.dina(n36705), .dinb(n36269), .dout(n36706));
  jxor g19444(.dina(n36263), .dinb(n293), .dout(n36707));
  jand g19445(.dina(n36707), .dinb(n36706), .dout(n36708));
  jor  g19446(.dina(n36708), .dinb(n36264), .dout(n36709));
  jxor g19447(.dina(n36258), .dinb(n294), .dout(n36710));
  jand g19448(.dina(n36710), .dinb(n36709), .dout(n36711));
  jor  g19449(.dina(n36711), .dinb(n36259), .dout(n36712));
  jxor g19450(.dina(n36246), .dinb(n295), .dout(n36713));
  jand g19451(.dina(n36713), .dinb(n36712), .dout(n36714));
  jor  g19452(.dina(n36714), .dinb(n36254), .dout(n36715));
  jor  g19453(.dina(n36715), .dinb(n36253), .dout(n36716));
  jnot g19454(.din(n36252), .dout(n36717));
  jand g19455(.dina(n36717), .dinb(b59 ), .dout(n36718));
  jor  g19456(.dina(n36718), .dinb(n832), .dout(n36719));
  jnot g19457(.din(n36719), .dout(n36720));
  jand g19458(.dina(n36720), .dinb(n36716), .dout(n36721));
  jor  g19459(.dina(n36721), .dinb(n36246), .dout(n36722));
  jnot g19460(.din(n36721), .dout(n36723));
  jxor g19461(.dina(n36713), .dinb(n36712), .dout(n36724));
  jor  g19462(.dina(n36724), .dinb(n36723), .dout(n36725));
  jand g19463(.dina(n36725), .dinb(n36722), .dout(n36726));
  jand g19464(.dina(n36715), .dinb(n302), .dout(n36727));
  jor  g19465(.dina(n36727), .dinb(n36723), .dout(n36728));
  jand g19466(.dina(n36728), .dinb(n36252), .dout(n36729));
  jand g19467(.dina(n36729), .dinb(n297), .dout(n36730));
  jand g19468(.dina(n36726), .dinb(n296), .dout(n36731));
  jor  g19469(.dina(n36721), .dinb(n36258), .dout(n36732));
  jxor g19470(.dina(n36710), .dinb(n36709), .dout(n36733));
  jor  g19471(.dina(n36733), .dinb(n36723), .dout(n36734));
  jand g19472(.dina(n36734), .dinb(n36732), .dout(n36735));
  jand g19473(.dina(n36735), .dinb(n295), .dout(n36736));
  jor  g19474(.dina(n36721), .dinb(n36263), .dout(n36737));
  jxor g19475(.dina(n36707), .dinb(n36706), .dout(n36738));
  jor  g19476(.dina(n36738), .dinb(n36723), .dout(n36739));
  jand g19477(.dina(n36739), .dinb(n36737), .dout(n36740));
  jand g19478(.dina(n36740), .dinb(n294), .dout(n36741));
  jor  g19479(.dina(n36721), .dinb(n36268), .dout(n36742));
  jxor g19480(.dina(n36704), .dinb(n36703), .dout(n36743));
  jor  g19481(.dina(n36743), .dinb(n36723), .dout(n36744));
  jand g19482(.dina(n36744), .dinb(n36742), .dout(n36745));
  jand g19483(.dina(n36745), .dinb(n293), .dout(n36746));
  jor  g19484(.dina(n36721), .dinb(n36273), .dout(n36747));
  jxor g19485(.dina(n36701), .dinb(n36700), .dout(n36748));
  jor  g19486(.dina(n36748), .dinb(n36723), .dout(n36749));
  jand g19487(.dina(n36749), .dinb(n36747), .dout(n36750));
  jand g19488(.dina(n36750), .dinb(n292), .dout(n36751));
  jor  g19489(.dina(n36721), .dinb(n36278), .dout(n36752));
  jxor g19490(.dina(n36698), .dinb(n36697), .dout(n36753));
  jor  g19491(.dina(n36753), .dinb(n36723), .dout(n36754));
  jand g19492(.dina(n36754), .dinb(n36752), .dout(n36755));
  jand g19493(.dina(n36755), .dinb(n291), .dout(n36756));
  jor  g19494(.dina(n36721), .dinb(n36283), .dout(n36757));
  jxor g19495(.dina(n36695), .dinb(n36694), .dout(n36758));
  jor  g19496(.dina(n36758), .dinb(n36723), .dout(n36759));
  jand g19497(.dina(n36759), .dinb(n36757), .dout(n36760));
  jand g19498(.dina(n36760), .dinb(n290), .dout(n36761));
  jor  g19499(.dina(n36721), .dinb(n36288), .dout(n36762));
  jxor g19500(.dina(n36692), .dinb(n36691), .dout(n36763));
  jor  g19501(.dina(n36763), .dinb(n36723), .dout(n36764));
  jand g19502(.dina(n36764), .dinb(n36762), .dout(n36765));
  jand g19503(.dina(n36765), .dinb(n289), .dout(n36766));
  jor  g19504(.dina(n36721), .dinb(n36293), .dout(n36767));
  jxor g19505(.dina(n36689), .dinb(n36688), .dout(n36768));
  jor  g19506(.dina(n36768), .dinb(n36723), .dout(n36769));
  jand g19507(.dina(n36769), .dinb(n36767), .dout(n36770));
  jand g19508(.dina(n36770), .dinb(n288), .dout(n36771));
  jor  g19509(.dina(n36721), .dinb(n36298), .dout(n36772));
  jxor g19510(.dina(n36686), .dinb(n36685), .dout(n36773));
  jor  g19511(.dina(n36773), .dinb(n36723), .dout(n36774));
  jand g19512(.dina(n36774), .dinb(n36772), .dout(n36775));
  jand g19513(.dina(n36775), .dinb(n287), .dout(n36776));
  jor  g19514(.dina(n36721), .dinb(n36303), .dout(n36777));
  jxor g19515(.dina(n36683), .dinb(n36682), .dout(n36778));
  jor  g19516(.dina(n36778), .dinb(n36723), .dout(n36779));
  jand g19517(.dina(n36779), .dinb(n36777), .dout(n36780));
  jand g19518(.dina(n36780), .dinb(n286), .dout(n36781));
  jor  g19519(.dina(n36721), .dinb(n36308), .dout(n36782));
  jxor g19520(.dina(n36680), .dinb(n36679), .dout(n36783));
  jor  g19521(.dina(n36783), .dinb(n36723), .dout(n36784));
  jand g19522(.dina(n36784), .dinb(n36782), .dout(n36785));
  jand g19523(.dina(n36785), .dinb(n285), .dout(n36786));
  jor  g19524(.dina(n36721), .dinb(n36313), .dout(n36787));
  jxor g19525(.dina(n36677), .dinb(n36676), .dout(n36788));
  jor  g19526(.dina(n36788), .dinb(n36723), .dout(n36789));
  jand g19527(.dina(n36789), .dinb(n36787), .dout(n36790));
  jand g19528(.dina(n36790), .dinb(n284), .dout(n36791));
  jor  g19529(.dina(n36721), .dinb(n36318), .dout(n36792));
  jxor g19530(.dina(n36674), .dinb(n36673), .dout(n36793));
  jor  g19531(.dina(n36793), .dinb(n36723), .dout(n36794));
  jand g19532(.dina(n36794), .dinb(n36792), .dout(n36795));
  jand g19533(.dina(n36795), .dinb(n317), .dout(n36796));
  jor  g19534(.dina(n36721), .dinb(n36323), .dout(n36797));
  jxor g19535(.dina(n36671), .dinb(n36670), .dout(n36798));
  jor  g19536(.dina(n36798), .dinb(n36723), .dout(n36799));
  jand g19537(.dina(n36799), .dinb(n36797), .dout(n36800));
  jand g19538(.dina(n36800), .dinb(n316), .dout(n36801));
  jor  g19539(.dina(n36721), .dinb(n36328), .dout(n36802));
  jxor g19540(.dina(n36668), .dinb(n36667), .dout(n36803));
  jor  g19541(.dina(n36803), .dinb(n36723), .dout(n36804));
  jand g19542(.dina(n36804), .dinb(n36802), .dout(n36805));
  jand g19543(.dina(n36805), .dinb(n315), .dout(n36806));
  jor  g19544(.dina(n36721), .dinb(n36333), .dout(n36807));
  jxor g19545(.dina(n36665), .dinb(n36664), .dout(n36808));
  jor  g19546(.dina(n36808), .dinb(n36723), .dout(n36809));
  jand g19547(.dina(n36809), .dinb(n36807), .dout(n36810));
  jand g19548(.dina(n36810), .dinb(n283), .dout(n36811));
  jor  g19549(.dina(n36721), .dinb(n36338), .dout(n36812));
  jxor g19550(.dina(n36662), .dinb(n36661), .dout(n36813));
  jor  g19551(.dina(n36813), .dinb(n36723), .dout(n36814));
  jand g19552(.dina(n36814), .dinb(n36812), .dout(n36815));
  jand g19553(.dina(n36815), .dinb(n280), .dout(n36816));
  jor  g19554(.dina(n36721), .dinb(n36343), .dout(n36817));
  jxor g19555(.dina(n36659), .dinb(n36658), .dout(n36818));
  jor  g19556(.dina(n36818), .dinb(n36723), .dout(n36819));
  jand g19557(.dina(n36819), .dinb(n36817), .dout(n36820));
  jand g19558(.dina(n36820), .dinb(n279), .dout(n36821));
  jor  g19559(.dina(n36721), .dinb(n36348), .dout(n36822));
  jxor g19560(.dina(n36656), .dinb(n36655), .dout(n36823));
  jor  g19561(.dina(n36823), .dinb(n36723), .dout(n36824));
  jand g19562(.dina(n36824), .dinb(n36822), .dout(n36825));
  jand g19563(.dina(n36825), .dinb(n278), .dout(n36826));
  jor  g19564(.dina(n36721), .dinb(n36353), .dout(n36827));
  jxor g19565(.dina(n36653), .dinb(n36652), .dout(n36828));
  jor  g19566(.dina(n36828), .dinb(n36723), .dout(n36829));
  jand g19567(.dina(n36829), .dinb(n36827), .dout(n36830));
  jand g19568(.dina(n36830), .dinb(n277), .dout(n36831));
  jor  g19569(.dina(n36721), .dinb(n36358), .dout(n36832));
  jxor g19570(.dina(n36650), .dinb(n36649), .dout(n36833));
  jor  g19571(.dina(n36833), .dinb(n36723), .dout(n36834));
  jand g19572(.dina(n36834), .dinb(n36832), .dout(n36835));
  jand g19573(.dina(n36835), .dinb(n326), .dout(n36836));
  jor  g19574(.dina(n36721), .dinb(n36363), .dout(n36837));
  jxor g19575(.dina(n36647), .dinb(n36646), .dout(n36838));
  jor  g19576(.dina(n36838), .dinb(n36723), .dout(n36839));
  jand g19577(.dina(n36839), .dinb(n36837), .dout(n36840));
  jand g19578(.dina(n36840), .dinb(n325), .dout(n36841));
  jor  g19579(.dina(n36721), .dinb(n36368), .dout(n36842));
  jxor g19580(.dina(n36644), .dinb(n36643), .dout(n36843));
  jor  g19581(.dina(n36843), .dinb(n36723), .dout(n36844));
  jand g19582(.dina(n36844), .dinb(n36842), .dout(n36845));
  jand g19583(.dina(n36845), .dinb(n324), .dout(n36846));
  jor  g19584(.dina(n36721), .dinb(n36373), .dout(n36847));
  jxor g19585(.dina(n36641), .dinb(n36640), .dout(n36848));
  jor  g19586(.dina(n36848), .dinb(n36723), .dout(n36849));
  jand g19587(.dina(n36849), .dinb(n36847), .dout(n36850));
  jand g19588(.dina(n36850), .dinb(n276), .dout(n36851));
  jor  g19589(.dina(n36721), .dinb(n36378), .dout(n36852));
  jxor g19590(.dina(n36638), .dinb(n36637), .dout(n36853));
  jor  g19591(.dina(n36853), .dinb(n36723), .dout(n36854));
  jand g19592(.dina(n36854), .dinb(n36852), .dout(n36855));
  jand g19593(.dina(n36855), .dinb(n333), .dout(n36856));
  jor  g19594(.dina(n36721), .dinb(n36383), .dout(n36857));
  jxor g19595(.dina(n36635), .dinb(n36634), .dout(n36858));
  jor  g19596(.dina(n36858), .dinb(n36723), .dout(n36859));
  jand g19597(.dina(n36859), .dinb(n36857), .dout(n36860));
  jand g19598(.dina(n36860), .dinb(n332), .dout(n36861));
  jor  g19599(.dina(n36721), .dinb(n36388), .dout(n36862));
  jxor g19600(.dina(n36632), .dinb(n36631), .dout(n36863));
  jor  g19601(.dina(n36863), .dinb(n36723), .dout(n36864));
  jand g19602(.dina(n36864), .dinb(n36862), .dout(n36865));
  jand g19603(.dina(n36865), .dinb(n331), .dout(n36866));
  jor  g19604(.dina(n36721), .dinb(n36393), .dout(n36867));
  jxor g19605(.dina(n36629), .dinb(n36628), .dout(n36868));
  jor  g19606(.dina(n36868), .dinb(n36723), .dout(n36869));
  jand g19607(.dina(n36869), .dinb(n36867), .dout(n36870));
  jand g19608(.dina(n36870), .dinb(n275), .dout(n36871));
  jor  g19609(.dina(n36721), .dinb(n36398), .dout(n36872));
  jxor g19610(.dina(n36626), .dinb(n36625), .dout(n36873));
  jor  g19611(.dina(n36873), .dinb(n36723), .dout(n36874));
  jand g19612(.dina(n36874), .dinb(n36872), .dout(n36875));
  jand g19613(.dina(n36875), .dinb(n340), .dout(n36876));
  jor  g19614(.dina(n36721), .dinb(n36403), .dout(n36877));
  jxor g19615(.dina(n36623), .dinb(n36622), .dout(n36878));
  jor  g19616(.dina(n36878), .dinb(n36723), .dout(n36879));
  jand g19617(.dina(n36879), .dinb(n36877), .dout(n36880));
  jand g19618(.dina(n36880), .dinb(n339), .dout(n36881));
  jor  g19619(.dina(n36721), .dinb(n36408), .dout(n36882));
  jxor g19620(.dina(n36620), .dinb(n36619), .dout(n36883));
  jor  g19621(.dina(n36883), .dinb(n36723), .dout(n36884));
  jand g19622(.dina(n36884), .dinb(n36882), .dout(n36885));
  jand g19623(.dina(n36885), .dinb(n338), .dout(n36886));
  jor  g19624(.dina(n36721), .dinb(n36413), .dout(n36887));
  jxor g19625(.dina(n36617), .dinb(n36616), .dout(n36888));
  jor  g19626(.dina(n36888), .dinb(n36723), .dout(n36889));
  jand g19627(.dina(n36889), .dinb(n36887), .dout(n36890));
  jand g19628(.dina(n36890), .dinb(n271), .dout(n36891));
  jor  g19629(.dina(n36721), .dinb(n36418), .dout(n36892));
  jxor g19630(.dina(n36614), .dinb(n36613), .dout(n36893));
  jor  g19631(.dina(n36893), .dinb(n36723), .dout(n36894));
  jand g19632(.dina(n36894), .dinb(n36892), .dout(n36895));
  jand g19633(.dina(n36895), .dinb(n270), .dout(n36896));
  jor  g19634(.dina(n36721), .dinb(n36423), .dout(n36897));
  jxor g19635(.dina(n36611), .dinb(n36610), .dout(n36898));
  jor  g19636(.dina(n36898), .dinb(n36723), .dout(n36899));
  jand g19637(.dina(n36899), .dinb(n36897), .dout(n36900));
  jand g19638(.dina(n36900), .dinb(n269), .dout(n36901));
  jor  g19639(.dina(n36721), .dinb(n36428), .dout(n36902));
  jxor g19640(.dina(n36608), .dinb(n36607), .dout(n36903));
  jor  g19641(.dina(n36903), .dinb(n36723), .dout(n36904));
  jand g19642(.dina(n36904), .dinb(n36902), .dout(n36905));
  jand g19643(.dina(n36905), .dinb(n274), .dout(n36906));
  jor  g19644(.dina(n36721), .dinb(n36433), .dout(n36907));
  jxor g19645(.dina(n36605), .dinb(n36604), .dout(n36908));
  jor  g19646(.dina(n36908), .dinb(n36723), .dout(n36909));
  jand g19647(.dina(n36909), .dinb(n36907), .dout(n36910));
  jand g19648(.dina(n36910), .dinb(n268), .dout(n36911));
  jor  g19649(.dina(n36721), .dinb(n36438), .dout(n36912));
  jxor g19650(.dina(n36602), .dinb(n36601), .dout(n36913));
  jor  g19651(.dina(n36913), .dinb(n36723), .dout(n36914));
  jand g19652(.dina(n36914), .dinb(n36912), .dout(n36915));
  jand g19653(.dina(n36915), .dinb(n349), .dout(n36916));
  jor  g19654(.dina(n36721), .dinb(n36443), .dout(n36917));
  jxor g19655(.dina(n36599), .dinb(n36598), .dout(n36918));
  jor  g19656(.dina(n36918), .dinb(n36723), .dout(n36919));
  jand g19657(.dina(n36919), .dinb(n36917), .dout(n36920));
  jand g19658(.dina(n36920), .dinb(n348), .dout(n36921));
  jor  g19659(.dina(n36721), .dinb(n36448), .dout(n36922));
  jxor g19660(.dina(n36596), .dinb(n36595), .dout(n36923));
  jor  g19661(.dina(n36923), .dinb(n36723), .dout(n36924));
  jand g19662(.dina(n36924), .dinb(n36922), .dout(n36925));
  jand g19663(.dina(n36925), .dinb(n347), .dout(n36926));
  jor  g19664(.dina(n36721), .dinb(n36453), .dout(n36927));
  jxor g19665(.dina(n36593), .dinb(n36592), .dout(n36928));
  jor  g19666(.dina(n36928), .dinb(n36723), .dout(n36929));
  jand g19667(.dina(n36929), .dinb(n36927), .dout(n36930));
  jand g19668(.dina(n36930), .dinb(n267), .dout(n36931));
  jor  g19669(.dina(n36721), .dinb(n36458), .dout(n36932));
  jxor g19670(.dina(n36590), .dinb(n36589), .dout(n36933));
  jor  g19671(.dina(n36933), .dinb(n36723), .dout(n36934));
  jand g19672(.dina(n36934), .dinb(n36932), .dout(n36935));
  jand g19673(.dina(n36935), .dinb(n266), .dout(n36936));
  jor  g19674(.dina(n36721), .dinb(n36463), .dout(n36937));
  jxor g19675(.dina(n36587), .dinb(n36586), .dout(n36938));
  jor  g19676(.dina(n36938), .dinb(n36723), .dout(n36939));
  jand g19677(.dina(n36939), .dinb(n36937), .dout(n36940));
  jand g19678(.dina(n36940), .dinb(n356), .dout(n36941));
  jor  g19679(.dina(n36721), .dinb(n36468), .dout(n36942));
  jxor g19680(.dina(n36584), .dinb(n36583), .dout(n36943));
  jor  g19681(.dina(n36943), .dinb(n36723), .dout(n36944));
  jand g19682(.dina(n36944), .dinb(n36942), .dout(n36945));
  jand g19683(.dina(n36945), .dinb(n355), .dout(n36946));
  jor  g19684(.dina(n36721), .dinb(n36473), .dout(n36947));
  jxor g19685(.dina(n36581), .dinb(n36580), .dout(n36948));
  jor  g19686(.dina(n36948), .dinb(n36723), .dout(n36949));
  jand g19687(.dina(n36949), .dinb(n36947), .dout(n36950));
  jand g19688(.dina(n36950), .dinb(n364), .dout(n36951));
  jor  g19689(.dina(n36721), .dinb(n36478), .dout(n36952));
  jxor g19690(.dina(n36578), .dinb(n36577), .dout(n36953));
  jor  g19691(.dina(n36953), .dinb(n36723), .dout(n36954));
  jand g19692(.dina(n36954), .dinb(n36952), .dout(n36955));
  jand g19693(.dina(n36955), .dinb(n361), .dout(n36956));
  jor  g19694(.dina(n36721), .dinb(n36483), .dout(n36957));
  jxor g19695(.dina(n36575), .dinb(n36574), .dout(n36958));
  jor  g19696(.dina(n36958), .dinb(n36723), .dout(n36959));
  jand g19697(.dina(n36959), .dinb(n36957), .dout(n36960));
  jand g19698(.dina(n36960), .dinb(n360), .dout(n36961));
  jor  g19699(.dina(n36721), .dinb(n36488), .dout(n36962));
  jxor g19700(.dina(n36572), .dinb(n36571), .dout(n36963));
  jor  g19701(.dina(n36963), .dinb(n36723), .dout(n36964));
  jand g19702(.dina(n36964), .dinb(n36962), .dout(n36965));
  jand g19703(.dina(n36965), .dinb(n363), .dout(n36966));
  jor  g19704(.dina(n36721), .dinb(n36493), .dout(n36967));
  jxor g19705(.dina(n36569), .dinb(n36568), .dout(n36968));
  jor  g19706(.dina(n36968), .dinb(n36723), .dout(n36969));
  jand g19707(.dina(n36969), .dinb(n36967), .dout(n36970));
  jand g19708(.dina(n36970), .dinb(n359), .dout(n36971));
  jor  g19709(.dina(n36721), .dinb(n36498), .dout(n36972));
  jxor g19710(.dina(n36566), .dinb(n36565), .dout(n36973));
  jor  g19711(.dina(n36973), .dinb(n36723), .dout(n36974));
  jand g19712(.dina(n36974), .dinb(n36972), .dout(n36975));
  jand g19713(.dina(n36975), .dinb(n369), .dout(n36976));
  jor  g19714(.dina(n36721), .dinb(n36503), .dout(n36977));
  jxor g19715(.dina(n36563), .dinb(n36562), .dout(n36978));
  jor  g19716(.dina(n36978), .dinb(n36723), .dout(n36979));
  jand g19717(.dina(n36979), .dinb(n36977), .dout(n36980));
  jand g19718(.dina(n36980), .dinb(n368), .dout(n36981));
  jor  g19719(.dina(n36721), .dinb(n36508), .dout(n36982));
  jxor g19720(.dina(n36560), .dinb(n36559), .dout(n36983));
  jor  g19721(.dina(n36983), .dinb(n36723), .dout(n36984));
  jand g19722(.dina(n36984), .dinb(n36982), .dout(n36985));
  jand g19723(.dina(n36985), .dinb(n367), .dout(n36986));
  jor  g19724(.dina(n36721), .dinb(n36513), .dout(n36987));
  jxor g19725(.dina(n36557), .dinb(n36556), .dout(n36988));
  jor  g19726(.dina(n36988), .dinb(n36723), .dout(n36989));
  jand g19727(.dina(n36989), .dinb(n36987), .dout(n36990));
  jand g19728(.dina(n36990), .dinb(n265), .dout(n36991));
  jor  g19729(.dina(n36721), .dinb(n36518), .dout(n36992));
  jxor g19730(.dina(n36554), .dinb(n36553), .dout(n36993));
  jor  g19731(.dina(n36993), .dinb(n36723), .dout(n36994));
  jand g19732(.dina(n36994), .dinb(n36992), .dout(n36995));
  jand g19733(.dina(n36995), .dinb(n378), .dout(n36996));
  jor  g19734(.dina(n36721), .dinb(n36523), .dout(n36997));
  jxor g19735(.dina(n36551), .dinb(n36550), .dout(n36998));
  jor  g19736(.dina(n36998), .dinb(n36723), .dout(n36999));
  jand g19737(.dina(n36999), .dinb(n36997), .dout(n37000));
  jand g19738(.dina(n37000), .dinb(n377), .dout(n37001));
  jor  g19739(.dina(n36721), .dinb(n36528), .dout(n37002));
  jxor g19740(.dina(n36548), .dinb(n36547), .dout(n37003));
  jor  g19741(.dina(n37003), .dinb(n36723), .dout(n37004));
  jand g19742(.dina(n37004), .dinb(n37002), .dout(n37005));
  jand g19743(.dina(n37005), .dinb(n376), .dout(n37006));
  jor  g19744(.dina(n36721), .dinb(n36536), .dout(n37007));
  jxor g19745(.dina(n36545), .dinb(n36544), .dout(n37008));
  jor  g19746(.dina(n37008), .dinb(n36723), .dout(n37009));
  jand g19747(.dina(n37009), .dinb(n37007), .dout(n37010));
  jand g19748(.dina(n37010), .dinb(n264), .dout(n37011));
  jor  g19749(.dina(n36721), .dinb(n36541), .dout(n37012));
  jxor g19750(.dina(n36542), .dinb(n15614), .dout(n37013));
  jand g19751(.dina(n37013), .dinb(n36721), .dout(n37014));
  jnot g19752(.din(n37014), .dout(n37015));
  jand g19753(.dina(n37015), .dinb(n37012), .dout(n37016));
  jnot g19754(.din(n37016), .dout(n37017));
  jand g19755(.dina(n37017), .dinb(n386), .dout(n37018));
  jand g19756(.dina(n36721), .dinb(b0 ), .dout(n37019));
  jxor g19757(.dina(n37019), .dinb(a4 ), .dout(n37020));
  jand g19758(.dina(n37020), .dinb(n259), .dout(n37021));
  jxor g19759(.dina(n37019), .dinb(n15612), .dout(n37022));
  jxor g19760(.dina(n37022), .dinb(b1 ), .dout(n37023));
  jand g19761(.dina(n37023), .dinb(n16097), .dout(n37024));
  jor  g19762(.dina(n37024), .dinb(n37021), .dout(n37025));
  jxor g19763(.dina(n37016), .dinb(b2 ), .dout(n37026));
  jand g19764(.dina(n37026), .dinb(n37025), .dout(n37027));
  jor  g19765(.dina(n37027), .dinb(n37018), .dout(n37028));
  jxor g19766(.dina(n37010), .dinb(n264), .dout(n37029));
  jand g19767(.dina(n37029), .dinb(n37028), .dout(n37030));
  jor  g19768(.dina(n37030), .dinb(n37011), .dout(n37031));
  jxor g19769(.dina(n37005), .dinb(n376), .dout(n37032));
  jand g19770(.dina(n37032), .dinb(n37031), .dout(n37033));
  jor  g19771(.dina(n37033), .dinb(n37006), .dout(n37034));
  jxor g19772(.dina(n37000), .dinb(n377), .dout(n37035));
  jand g19773(.dina(n37035), .dinb(n37034), .dout(n37036));
  jor  g19774(.dina(n37036), .dinb(n37001), .dout(n37037));
  jxor g19775(.dina(n36995), .dinb(n378), .dout(n37038));
  jand g19776(.dina(n37038), .dinb(n37037), .dout(n37039));
  jor  g19777(.dina(n37039), .dinb(n36996), .dout(n37040));
  jxor g19778(.dina(n36990), .dinb(n265), .dout(n37041));
  jand g19779(.dina(n37041), .dinb(n37040), .dout(n37042));
  jor  g19780(.dina(n37042), .dinb(n36991), .dout(n37043));
  jxor g19781(.dina(n36985), .dinb(n367), .dout(n37044));
  jand g19782(.dina(n37044), .dinb(n37043), .dout(n37045));
  jor  g19783(.dina(n37045), .dinb(n36986), .dout(n37046));
  jxor g19784(.dina(n36980), .dinb(n368), .dout(n37047));
  jand g19785(.dina(n37047), .dinb(n37046), .dout(n37048));
  jor  g19786(.dina(n37048), .dinb(n36981), .dout(n37049));
  jxor g19787(.dina(n36975), .dinb(n369), .dout(n37050));
  jand g19788(.dina(n37050), .dinb(n37049), .dout(n37051));
  jor  g19789(.dina(n37051), .dinb(n36976), .dout(n37052));
  jxor g19790(.dina(n36970), .dinb(n359), .dout(n37053));
  jand g19791(.dina(n37053), .dinb(n37052), .dout(n37054));
  jor  g19792(.dina(n37054), .dinb(n36971), .dout(n37055));
  jxor g19793(.dina(n36965), .dinb(n363), .dout(n37056));
  jand g19794(.dina(n37056), .dinb(n37055), .dout(n37057));
  jor  g19795(.dina(n37057), .dinb(n36966), .dout(n37058));
  jxor g19796(.dina(n36960), .dinb(n360), .dout(n37059));
  jand g19797(.dina(n37059), .dinb(n37058), .dout(n37060));
  jor  g19798(.dina(n37060), .dinb(n36961), .dout(n37061));
  jxor g19799(.dina(n36955), .dinb(n361), .dout(n37062));
  jand g19800(.dina(n37062), .dinb(n37061), .dout(n37063));
  jor  g19801(.dina(n37063), .dinb(n36956), .dout(n37064));
  jxor g19802(.dina(n36950), .dinb(n364), .dout(n37065));
  jand g19803(.dina(n37065), .dinb(n37064), .dout(n37066));
  jor  g19804(.dina(n37066), .dinb(n36951), .dout(n37067));
  jxor g19805(.dina(n36945), .dinb(n355), .dout(n37068));
  jand g19806(.dina(n37068), .dinb(n37067), .dout(n37069));
  jor  g19807(.dina(n37069), .dinb(n36946), .dout(n37070));
  jxor g19808(.dina(n36940), .dinb(n356), .dout(n37071));
  jand g19809(.dina(n37071), .dinb(n37070), .dout(n37072));
  jor  g19810(.dina(n37072), .dinb(n36941), .dout(n37073));
  jxor g19811(.dina(n36935), .dinb(n266), .dout(n37074));
  jand g19812(.dina(n37074), .dinb(n37073), .dout(n37075));
  jor  g19813(.dina(n37075), .dinb(n36936), .dout(n37076));
  jxor g19814(.dina(n36930), .dinb(n267), .dout(n37077));
  jand g19815(.dina(n37077), .dinb(n37076), .dout(n37078));
  jor  g19816(.dina(n37078), .dinb(n36931), .dout(n37079));
  jxor g19817(.dina(n36925), .dinb(n347), .dout(n37080));
  jand g19818(.dina(n37080), .dinb(n37079), .dout(n37081));
  jor  g19819(.dina(n37081), .dinb(n36926), .dout(n37082));
  jxor g19820(.dina(n36920), .dinb(n348), .dout(n37083));
  jand g19821(.dina(n37083), .dinb(n37082), .dout(n37084));
  jor  g19822(.dina(n37084), .dinb(n36921), .dout(n37085));
  jxor g19823(.dina(n36915), .dinb(n349), .dout(n37086));
  jand g19824(.dina(n37086), .dinb(n37085), .dout(n37087));
  jor  g19825(.dina(n37087), .dinb(n36916), .dout(n37088));
  jxor g19826(.dina(n36910), .dinb(n268), .dout(n37089));
  jand g19827(.dina(n37089), .dinb(n37088), .dout(n37090));
  jor  g19828(.dina(n37090), .dinb(n36911), .dout(n37091));
  jxor g19829(.dina(n36905), .dinb(n274), .dout(n37092));
  jand g19830(.dina(n37092), .dinb(n37091), .dout(n37093));
  jor  g19831(.dina(n37093), .dinb(n36906), .dout(n37094));
  jxor g19832(.dina(n36900), .dinb(n269), .dout(n37095));
  jand g19833(.dina(n37095), .dinb(n37094), .dout(n37096));
  jor  g19834(.dina(n37096), .dinb(n36901), .dout(n37097));
  jxor g19835(.dina(n36895), .dinb(n270), .dout(n37098));
  jand g19836(.dina(n37098), .dinb(n37097), .dout(n37099));
  jor  g19837(.dina(n37099), .dinb(n36896), .dout(n37100));
  jxor g19838(.dina(n36890), .dinb(n271), .dout(n37101));
  jand g19839(.dina(n37101), .dinb(n37100), .dout(n37102));
  jor  g19840(.dina(n37102), .dinb(n36891), .dout(n37103));
  jxor g19841(.dina(n36885), .dinb(n338), .dout(n37104));
  jand g19842(.dina(n37104), .dinb(n37103), .dout(n37105));
  jor  g19843(.dina(n37105), .dinb(n36886), .dout(n37106));
  jxor g19844(.dina(n36880), .dinb(n339), .dout(n37107));
  jand g19845(.dina(n37107), .dinb(n37106), .dout(n37108));
  jor  g19846(.dina(n37108), .dinb(n36881), .dout(n37109));
  jxor g19847(.dina(n36875), .dinb(n340), .dout(n37110));
  jand g19848(.dina(n37110), .dinb(n37109), .dout(n37111));
  jor  g19849(.dina(n37111), .dinb(n36876), .dout(n37112));
  jxor g19850(.dina(n36870), .dinb(n275), .dout(n37113));
  jand g19851(.dina(n37113), .dinb(n37112), .dout(n37114));
  jor  g19852(.dina(n37114), .dinb(n36871), .dout(n37115));
  jxor g19853(.dina(n36865), .dinb(n331), .dout(n37116));
  jand g19854(.dina(n37116), .dinb(n37115), .dout(n37117));
  jor  g19855(.dina(n37117), .dinb(n36866), .dout(n37118));
  jxor g19856(.dina(n36860), .dinb(n332), .dout(n37119));
  jand g19857(.dina(n37119), .dinb(n37118), .dout(n37120));
  jor  g19858(.dina(n37120), .dinb(n36861), .dout(n37121));
  jxor g19859(.dina(n36855), .dinb(n333), .dout(n37122));
  jand g19860(.dina(n37122), .dinb(n37121), .dout(n37123));
  jor  g19861(.dina(n37123), .dinb(n36856), .dout(n37124));
  jxor g19862(.dina(n36850), .dinb(n276), .dout(n37125));
  jand g19863(.dina(n37125), .dinb(n37124), .dout(n37126));
  jor  g19864(.dina(n37126), .dinb(n36851), .dout(n37127));
  jxor g19865(.dina(n36845), .dinb(n324), .dout(n37128));
  jand g19866(.dina(n37128), .dinb(n37127), .dout(n37129));
  jor  g19867(.dina(n37129), .dinb(n36846), .dout(n37130));
  jxor g19868(.dina(n36840), .dinb(n325), .dout(n37131));
  jand g19869(.dina(n37131), .dinb(n37130), .dout(n37132));
  jor  g19870(.dina(n37132), .dinb(n36841), .dout(n37133));
  jxor g19871(.dina(n36835), .dinb(n326), .dout(n37134));
  jand g19872(.dina(n37134), .dinb(n37133), .dout(n37135));
  jor  g19873(.dina(n37135), .dinb(n36836), .dout(n37136));
  jxor g19874(.dina(n36830), .dinb(n277), .dout(n37137));
  jand g19875(.dina(n37137), .dinb(n37136), .dout(n37138));
  jor  g19876(.dina(n37138), .dinb(n36831), .dout(n37139));
  jxor g19877(.dina(n36825), .dinb(n278), .dout(n37140));
  jand g19878(.dina(n37140), .dinb(n37139), .dout(n37141));
  jor  g19879(.dina(n37141), .dinb(n36826), .dout(n37142));
  jxor g19880(.dina(n36820), .dinb(n279), .dout(n37143));
  jand g19881(.dina(n37143), .dinb(n37142), .dout(n37144));
  jor  g19882(.dina(n37144), .dinb(n36821), .dout(n37145));
  jxor g19883(.dina(n36815), .dinb(n280), .dout(n37146));
  jand g19884(.dina(n37146), .dinb(n37145), .dout(n37147));
  jor  g19885(.dina(n37147), .dinb(n36816), .dout(n37148));
  jxor g19886(.dina(n36810), .dinb(n283), .dout(n37149));
  jand g19887(.dina(n37149), .dinb(n37148), .dout(n37150));
  jor  g19888(.dina(n37150), .dinb(n36811), .dout(n37151));
  jxor g19889(.dina(n36805), .dinb(n315), .dout(n37152));
  jand g19890(.dina(n37152), .dinb(n37151), .dout(n37153));
  jor  g19891(.dina(n37153), .dinb(n36806), .dout(n37154));
  jxor g19892(.dina(n36800), .dinb(n316), .dout(n37155));
  jand g19893(.dina(n37155), .dinb(n37154), .dout(n37156));
  jor  g19894(.dina(n37156), .dinb(n36801), .dout(n37157));
  jxor g19895(.dina(n36795), .dinb(n317), .dout(n37158));
  jand g19896(.dina(n37158), .dinb(n37157), .dout(n37159));
  jor  g19897(.dina(n37159), .dinb(n36796), .dout(n37160));
  jxor g19898(.dina(n36790), .dinb(n284), .dout(n37161));
  jand g19899(.dina(n37161), .dinb(n37160), .dout(n37162));
  jor  g19900(.dina(n37162), .dinb(n36791), .dout(n37163));
  jxor g19901(.dina(n36785), .dinb(n285), .dout(n37164));
  jand g19902(.dina(n37164), .dinb(n37163), .dout(n37165));
  jor  g19903(.dina(n37165), .dinb(n36786), .dout(n37166));
  jxor g19904(.dina(n36780), .dinb(n286), .dout(n37167));
  jand g19905(.dina(n37167), .dinb(n37166), .dout(n37168));
  jor  g19906(.dina(n37168), .dinb(n36781), .dout(n37169));
  jxor g19907(.dina(n36775), .dinb(n287), .dout(n37170));
  jand g19908(.dina(n37170), .dinb(n37169), .dout(n37171));
  jor  g19909(.dina(n37171), .dinb(n36776), .dout(n37172));
  jxor g19910(.dina(n36770), .dinb(n288), .dout(n37173));
  jand g19911(.dina(n37173), .dinb(n37172), .dout(n37174));
  jor  g19912(.dina(n37174), .dinb(n36771), .dout(n37175));
  jxor g19913(.dina(n36765), .dinb(n289), .dout(n37176));
  jand g19914(.dina(n37176), .dinb(n37175), .dout(n37177));
  jor  g19915(.dina(n37177), .dinb(n36766), .dout(n37178));
  jxor g19916(.dina(n36760), .dinb(n290), .dout(n37179));
  jand g19917(.dina(n37179), .dinb(n37178), .dout(n37180));
  jor  g19918(.dina(n37180), .dinb(n36761), .dout(n37181));
  jxor g19919(.dina(n36755), .dinb(n291), .dout(n37182));
  jand g19920(.dina(n37182), .dinb(n37181), .dout(n37183));
  jor  g19921(.dina(n37183), .dinb(n36756), .dout(n37184));
  jxor g19922(.dina(n36750), .dinb(n292), .dout(n37185));
  jand g19923(.dina(n37185), .dinb(n37184), .dout(n37186));
  jor  g19924(.dina(n37186), .dinb(n36751), .dout(n37187));
  jxor g19925(.dina(n36745), .dinb(n293), .dout(n37188));
  jand g19926(.dina(n37188), .dinb(n37187), .dout(n37189));
  jor  g19927(.dina(n37189), .dinb(n36746), .dout(n37190));
  jxor g19928(.dina(n36740), .dinb(n294), .dout(n37191));
  jand g19929(.dina(n37191), .dinb(n37190), .dout(n37192));
  jor  g19930(.dina(n37192), .dinb(n36741), .dout(n37193));
  jxor g19931(.dina(n36735), .dinb(n295), .dout(n37194));
  jand g19932(.dina(n37194), .dinb(n37193), .dout(n37195));
  jor  g19933(.dina(n37195), .dinb(n36736), .dout(n37196));
  jxor g19934(.dina(n36726), .dinb(n296), .dout(n37197));
  jand g19935(.dina(n37197), .dinb(n37196), .dout(n37198));
  jor  g19936(.dina(n37198), .dinb(n36731), .dout(n37199));
  jor  g19937(.dina(n37199), .dinb(n36730), .dout(n37200));
  jnot g19938(.din(n36729), .dout(n37201));
  jand g19939(.dina(n37201), .dinb(b60 ), .dout(n37202));
  jor  g19940(.dina(n37202), .dinb(n831), .dout(n37203));
  jnot g19941(.din(n37203), .dout(n37204));
  jand g19942(.dina(n37204), .dinb(n37200), .dout(n37205));
  jor  g19943(.dina(n37205), .dinb(n36726), .dout(n37206));
  jnot g19944(.din(n37205), .dout(n37207));
  jxor g19945(.dina(n37197), .dinb(n37196), .dout(n37208));
  jor  g19946(.dina(n37208), .dinb(n37207), .dout(n37209));
  jand g19947(.dina(n37209), .dinb(n37206), .dout(n37210));
  jand g19948(.dina(n37210), .dinb(n297), .dout(n37211));
  jor  g19949(.dina(n37205), .dinb(n36735), .dout(n37212));
  jxor g19950(.dina(n37194), .dinb(n37193), .dout(n37213));
  jor  g19951(.dina(n37213), .dinb(n37207), .dout(n37214));
  jand g19952(.dina(n37214), .dinb(n37212), .dout(n37215));
  jand g19953(.dina(n37215), .dinb(n296), .dout(n37216));
  jor  g19954(.dina(n37205), .dinb(n36740), .dout(n37217));
  jxor g19955(.dina(n37191), .dinb(n37190), .dout(n37218));
  jor  g19956(.dina(n37218), .dinb(n37207), .dout(n37219));
  jand g19957(.dina(n37219), .dinb(n37217), .dout(n37220));
  jand g19958(.dina(n37220), .dinb(n295), .dout(n37221));
  jor  g19959(.dina(n37205), .dinb(n36745), .dout(n37222));
  jxor g19960(.dina(n37188), .dinb(n37187), .dout(n37223));
  jor  g19961(.dina(n37223), .dinb(n37207), .dout(n37224));
  jand g19962(.dina(n37224), .dinb(n37222), .dout(n37225));
  jand g19963(.dina(n37225), .dinb(n294), .dout(n37226));
  jor  g19964(.dina(n37205), .dinb(n36750), .dout(n37227));
  jxor g19965(.dina(n37185), .dinb(n37184), .dout(n37228));
  jor  g19966(.dina(n37228), .dinb(n37207), .dout(n37229));
  jand g19967(.dina(n37229), .dinb(n37227), .dout(n37230));
  jand g19968(.dina(n37230), .dinb(n293), .dout(n37231));
  jor  g19969(.dina(n37205), .dinb(n36755), .dout(n37232));
  jxor g19970(.dina(n37182), .dinb(n37181), .dout(n37233));
  jor  g19971(.dina(n37233), .dinb(n37207), .dout(n37234));
  jand g19972(.dina(n37234), .dinb(n37232), .dout(n37235));
  jand g19973(.dina(n37235), .dinb(n292), .dout(n37236));
  jor  g19974(.dina(n37205), .dinb(n36760), .dout(n37237));
  jxor g19975(.dina(n37179), .dinb(n37178), .dout(n37238));
  jor  g19976(.dina(n37238), .dinb(n37207), .dout(n37239));
  jand g19977(.dina(n37239), .dinb(n37237), .dout(n37240));
  jand g19978(.dina(n37240), .dinb(n291), .dout(n37241));
  jor  g19979(.dina(n37205), .dinb(n36765), .dout(n37242));
  jxor g19980(.dina(n37176), .dinb(n37175), .dout(n37243));
  jor  g19981(.dina(n37243), .dinb(n37207), .dout(n37244));
  jand g19982(.dina(n37244), .dinb(n37242), .dout(n37245));
  jand g19983(.dina(n37245), .dinb(n290), .dout(n37246));
  jor  g19984(.dina(n37205), .dinb(n36770), .dout(n37247));
  jxor g19985(.dina(n37173), .dinb(n37172), .dout(n37248));
  jor  g19986(.dina(n37248), .dinb(n37207), .dout(n37249));
  jand g19987(.dina(n37249), .dinb(n37247), .dout(n37250));
  jand g19988(.dina(n37250), .dinb(n289), .dout(n37251));
  jor  g19989(.dina(n37205), .dinb(n36775), .dout(n37252));
  jxor g19990(.dina(n37170), .dinb(n37169), .dout(n37253));
  jor  g19991(.dina(n37253), .dinb(n37207), .dout(n37254));
  jand g19992(.dina(n37254), .dinb(n37252), .dout(n37255));
  jand g19993(.dina(n37255), .dinb(n288), .dout(n37256));
  jor  g19994(.dina(n37205), .dinb(n36780), .dout(n37257));
  jxor g19995(.dina(n37167), .dinb(n37166), .dout(n37258));
  jor  g19996(.dina(n37258), .dinb(n37207), .dout(n37259));
  jand g19997(.dina(n37259), .dinb(n37257), .dout(n37260));
  jand g19998(.dina(n37260), .dinb(n287), .dout(n37261));
  jor  g19999(.dina(n37205), .dinb(n36785), .dout(n37262));
  jxor g20000(.dina(n37164), .dinb(n37163), .dout(n37263));
  jor  g20001(.dina(n37263), .dinb(n37207), .dout(n37264));
  jand g20002(.dina(n37264), .dinb(n37262), .dout(n37265));
  jand g20003(.dina(n37265), .dinb(n286), .dout(n37266));
  jor  g20004(.dina(n37205), .dinb(n36790), .dout(n37267));
  jxor g20005(.dina(n37161), .dinb(n37160), .dout(n37268));
  jor  g20006(.dina(n37268), .dinb(n37207), .dout(n37269));
  jand g20007(.dina(n37269), .dinb(n37267), .dout(n37270));
  jand g20008(.dina(n37270), .dinb(n285), .dout(n37271));
  jor  g20009(.dina(n37205), .dinb(n36795), .dout(n37272));
  jxor g20010(.dina(n37158), .dinb(n37157), .dout(n37273));
  jor  g20011(.dina(n37273), .dinb(n37207), .dout(n37274));
  jand g20012(.dina(n37274), .dinb(n37272), .dout(n37275));
  jand g20013(.dina(n37275), .dinb(n284), .dout(n37276));
  jor  g20014(.dina(n37205), .dinb(n36800), .dout(n37277));
  jxor g20015(.dina(n37155), .dinb(n37154), .dout(n37278));
  jor  g20016(.dina(n37278), .dinb(n37207), .dout(n37279));
  jand g20017(.dina(n37279), .dinb(n37277), .dout(n37280));
  jand g20018(.dina(n37280), .dinb(n317), .dout(n37281));
  jor  g20019(.dina(n37205), .dinb(n36805), .dout(n37282));
  jxor g20020(.dina(n37152), .dinb(n37151), .dout(n37283));
  jor  g20021(.dina(n37283), .dinb(n37207), .dout(n37284));
  jand g20022(.dina(n37284), .dinb(n37282), .dout(n37285));
  jand g20023(.dina(n37285), .dinb(n316), .dout(n37286));
  jor  g20024(.dina(n37205), .dinb(n36810), .dout(n37287));
  jxor g20025(.dina(n37149), .dinb(n37148), .dout(n37288));
  jor  g20026(.dina(n37288), .dinb(n37207), .dout(n37289));
  jand g20027(.dina(n37289), .dinb(n37287), .dout(n37290));
  jand g20028(.dina(n37290), .dinb(n315), .dout(n37291));
  jor  g20029(.dina(n37205), .dinb(n36815), .dout(n37292));
  jxor g20030(.dina(n37146), .dinb(n37145), .dout(n37293));
  jor  g20031(.dina(n37293), .dinb(n37207), .dout(n37294));
  jand g20032(.dina(n37294), .dinb(n37292), .dout(n37295));
  jand g20033(.dina(n37295), .dinb(n283), .dout(n37296));
  jor  g20034(.dina(n37205), .dinb(n36820), .dout(n37297));
  jxor g20035(.dina(n37143), .dinb(n37142), .dout(n37298));
  jor  g20036(.dina(n37298), .dinb(n37207), .dout(n37299));
  jand g20037(.dina(n37299), .dinb(n37297), .dout(n37300));
  jand g20038(.dina(n37300), .dinb(n280), .dout(n37301));
  jor  g20039(.dina(n37205), .dinb(n36825), .dout(n37302));
  jxor g20040(.dina(n37140), .dinb(n37139), .dout(n37303));
  jor  g20041(.dina(n37303), .dinb(n37207), .dout(n37304));
  jand g20042(.dina(n37304), .dinb(n37302), .dout(n37305));
  jand g20043(.dina(n37305), .dinb(n279), .dout(n37306));
  jor  g20044(.dina(n37205), .dinb(n36830), .dout(n37307));
  jxor g20045(.dina(n37137), .dinb(n37136), .dout(n37308));
  jor  g20046(.dina(n37308), .dinb(n37207), .dout(n37309));
  jand g20047(.dina(n37309), .dinb(n37307), .dout(n37310));
  jand g20048(.dina(n37310), .dinb(n278), .dout(n37311));
  jor  g20049(.dina(n37205), .dinb(n36835), .dout(n37312));
  jxor g20050(.dina(n37134), .dinb(n37133), .dout(n37313));
  jor  g20051(.dina(n37313), .dinb(n37207), .dout(n37314));
  jand g20052(.dina(n37314), .dinb(n37312), .dout(n37315));
  jand g20053(.dina(n37315), .dinb(n277), .dout(n37316));
  jor  g20054(.dina(n37205), .dinb(n36840), .dout(n37317));
  jxor g20055(.dina(n37131), .dinb(n37130), .dout(n37318));
  jor  g20056(.dina(n37318), .dinb(n37207), .dout(n37319));
  jand g20057(.dina(n37319), .dinb(n37317), .dout(n37320));
  jand g20058(.dina(n37320), .dinb(n326), .dout(n37321));
  jor  g20059(.dina(n37205), .dinb(n36845), .dout(n37322));
  jxor g20060(.dina(n37128), .dinb(n37127), .dout(n37323));
  jor  g20061(.dina(n37323), .dinb(n37207), .dout(n37324));
  jand g20062(.dina(n37324), .dinb(n37322), .dout(n37325));
  jand g20063(.dina(n37325), .dinb(n325), .dout(n37326));
  jor  g20064(.dina(n37205), .dinb(n36850), .dout(n37327));
  jxor g20065(.dina(n37125), .dinb(n37124), .dout(n37328));
  jor  g20066(.dina(n37328), .dinb(n37207), .dout(n37329));
  jand g20067(.dina(n37329), .dinb(n37327), .dout(n37330));
  jand g20068(.dina(n37330), .dinb(n324), .dout(n37331));
  jor  g20069(.dina(n37205), .dinb(n36855), .dout(n37332));
  jxor g20070(.dina(n37122), .dinb(n37121), .dout(n37333));
  jor  g20071(.dina(n37333), .dinb(n37207), .dout(n37334));
  jand g20072(.dina(n37334), .dinb(n37332), .dout(n37335));
  jand g20073(.dina(n37335), .dinb(n276), .dout(n37336));
  jor  g20074(.dina(n37205), .dinb(n36860), .dout(n37337));
  jxor g20075(.dina(n37119), .dinb(n37118), .dout(n37338));
  jor  g20076(.dina(n37338), .dinb(n37207), .dout(n37339));
  jand g20077(.dina(n37339), .dinb(n37337), .dout(n37340));
  jand g20078(.dina(n37340), .dinb(n333), .dout(n37341));
  jor  g20079(.dina(n37205), .dinb(n36865), .dout(n37342));
  jxor g20080(.dina(n37116), .dinb(n37115), .dout(n37343));
  jor  g20081(.dina(n37343), .dinb(n37207), .dout(n37344));
  jand g20082(.dina(n37344), .dinb(n37342), .dout(n37345));
  jand g20083(.dina(n37345), .dinb(n332), .dout(n37346));
  jor  g20084(.dina(n37205), .dinb(n36870), .dout(n37347));
  jxor g20085(.dina(n37113), .dinb(n37112), .dout(n37348));
  jor  g20086(.dina(n37348), .dinb(n37207), .dout(n37349));
  jand g20087(.dina(n37349), .dinb(n37347), .dout(n37350));
  jand g20088(.dina(n37350), .dinb(n331), .dout(n37351));
  jor  g20089(.dina(n37205), .dinb(n36875), .dout(n37352));
  jxor g20090(.dina(n37110), .dinb(n37109), .dout(n37353));
  jor  g20091(.dina(n37353), .dinb(n37207), .dout(n37354));
  jand g20092(.dina(n37354), .dinb(n37352), .dout(n37355));
  jand g20093(.dina(n37355), .dinb(n275), .dout(n37356));
  jor  g20094(.dina(n37205), .dinb(n36880), .dout(n37357));
  jxor g20095(.dina(n37107), .dinb(n37106), .dout(n37358));
  jor  g20096(.dina(n37358), .dinb(n37207), .dout(n37359));
  jand g20097(.dina(n37359), .dinb(n37357), .dout(n37360));
  jand g20098(.dina(n37360), .dinb(n340), .dout(n37361));
  jor  g20099(.dina(n37205), .dinb(n36885), .dout(n37362));
  jxor g20100(.dina(n37104), .dinb(n37103), .dout(n37363));
  jor  g20101(.dina(n37363), .dinb(n37207), .dout(n37364));
  jand g20102(.dina(n37364), .dinb(n37362), .dout(n37365));
  jand g20103(.dina(n37365), .dinb(n339), .dout(n37366));
  jor  g20104(.dina(n37205), .dinb(n36890), .dout(n37367));
  jxor g20105(.dina(n37101), .dinb(n37100), .dout(n37368));
  jor  g20106(.dina(n37368), .dinb(n37207), .dout(n37369));
  jand g20107(.dina(n37369), .dinb(n37367), .dout(n37370));
  jand g20108(.dina(n37370), .dinb(n338), .dout(n37371));
  jor  g20109(.dina(n37205), .dinb(n36895), .dout(n37372));
  jxor g20110(.dina(n37098), .dinb(n37097), .dout(n37373));
  jor  g20111(.dina(n37373), .dinb(n37207), .dout(n37374));
  jand g20112(.dina(n37374), .dinb(n37372), .dout(n37375));
  jand g20113(.dina(n37375), .dinb(n271), .dout(n37376));
  jor  g20114(.dina(n37205), .dinb(n36900), .dout(n37377));
  jxor g20115(.dina(n37095), .dinb(n37094), .dout(n37378));
  jor  g20116(.dina(n37378), .dinb(n37207), .dout(n37379));
  jand g20117(.dina(n37379), .dinb(n37377), .dout(n37380));
  jand g20118(.dina(n37380), .dinb(n270), .dout(n37381));
  jor  g20119(.dina(n37205), .dinb(n36905), .dout(n37382));
  jxor g20120(.dina(n37092), .dinb(n37091), .dout(n37383));
  jor  g20121(.dina(n37383), .dinb(n37207), .dout(n37384));
  jand g20122(.dina(n37384), .dinb(n37382), .dout(n37385));
  jand g20123(.dina(n37385), .dinb(n269), .dout(n37386));
  jor  g20124(.dina(n37205), .dinb(n36910), .dout(n37387));
  jxor g20125(.dina(n37089), .dinb(n37088), .dout(n37388));
  jor  g20126(.dina(n37388), .dinb(n37207), .dout(n37389));
  jand g20127(.dina(n37389), .dinb(n37387), .dout(n37390));
  jand g20128(.dina(n37390), .dinb(n274), .dout(n37391));
  jor  g20129(.dina(n37205), .dinb(n36915), .dout(n37392));
  jxor g20130(.dina(n37086), .dinb(n37085), .dout(n37393));
  jor  g20131(.dina(n37393), .dinb(n37207), .dout(n37394));
  jand g20132(.dina(n37394), .dinb(n37392), .dout(n37395));
  jand g20133(.dina(n37395), .dinb(n268), .dout(n37396));
  jor  g20134(.dina(n37205), .dinb(n36920), .dout(n37397));
  jxor g20135(.dina(n37083), .dinb(n37082), .dout(n37398));
  jor  g20136(.dina(n37398), .dinb(n37207), .dout(n37399));
  jand g20137(.dina(n37399), .dinb(n37397), .dout(n37400));
  jand g20138(.dina(n37400), .dinb(n349), .dout(n37401));
  jor  g20139(.dina(n37205), .dinb(n36925), .dout(n37402));
  jxor g20140(.dina(n37080), .dinb(n37079), .dout(n37403));
  jor  g20141(.dina(n37403), .dinb(n37207), .dout(n37404));
  jand g20142(.dina(n37404), .dinb(n37402), .dout(n37405));
  jand g20143(.dina(n37405), .dinb(n348), .dout(n37406));
  jor  g20144(.dina(n37205), .dinb(n36930), .dout(n37407));
  jxor g20145(.dina(n37077), .dinb(n37076), .dout(n37408));
  jor  g20146(.dina(n37408), .dinb(n37207), .dout(n37409));
  jand g20147(.dina(n37409), .dinb(n37407), .dout(n37410));
  jand g20148(.dina(n37410), .dinb(n347), .dout(n37411));
  jor  g20149(.dina(n37205), .dinb(n36935), .dout(n37412));
  jxor g20150(.dina(n37074), .dinb(n37073), .dout(n37413));
  jor  g20151(.dina(n37413), .dinb(n37207), .dout(n37414));
  jand g20152(.dina(n37414), .dinb(n37412), .dout(n37415));
  jand g20153(.dina(n37415), .dinb(n267), .dout(n37416));
  jor  g20154(.dina(n37205), .dinb(n36940), .dout(n37417));
  jxor g20155(.dina(n37071), .dinb(n37070), .dout(n37418));
  jor  g20156(.dina(n37418), .dinb(n37207), .dout(n37419));
  jand g20157(.dina(n37419), .dinb(n37417), .dout(n37420));
  jand g20158(.dina(n37420), .dinb(n266), .dout(n37421));
  jor  g20159(.dina(n37205), .dinb(n36945), .dout(n37422));
  jxor g20160(.dina(n37068), .dinb(n37067), .dout(n37423));
  jor  g20161(.dina(n37423), .dinb(n37207), .dout(n37424));
  jand g20162(.dina(n37424), .dinb(n37422), .dout(n37425));
  jand g20163(.dina(n37425), .dinb(n356), .dout(n37426));
  jor  g20164(.dina(n37205), .dinb(n36950), .dout(n37427));
  jxor g20165(.dina(n37065), .dinb(n37064), .dout(n37428));
  jor  g20166(.dina(n37428), .dinb(n37207), .dout(n37429));
  jand g20167(.dina(n37429), .dinb(n37427), .dout(n37430));
  jand g20168(.dina(n37430), .dinb(n355), .dout(n37431));
  jor  g20169(.dina(n37205), .dinb(n36955), .dout(n37432));
  jxor g20170(.dina(n37062), .dinb(n37061), .dout(n37433));
  jor  g20171(.dina(n37433), .dinb(n37207), .dout(n37434));
  jand g20172(.dina(n37434), .dinb(n37432), .dout(n37435));
  jand g20173(.dina(n37435), .dinb(n364), .dout(n37436));
  jor  g20174(.dina(n37205), .dinb(n36960), .dout(n37437));
  jxor g20175(.dina(n37059), .dinb(n37058), .dout(n37438));
  jor  g20176(.dina(n37438), .dinb(n37207), .dout(n37439));
  jand g20177(.dina(n37439), .dinb(n37437), .dout(n37440));
  jand g20178(.dina(n37440), .dinb(n361), .dout(n37441));
  jor  g20179(.dina(n37205), .dinb(n36965), .dout(n37442));
  jxor g20180(.dina(n37056), .dinb(n37055), .dout(n37443));
  jor  g20181(.dina(n37443), .dinb(n37207), .dout(n37444));
  jand g20182(.dina(n37444), .dinb(n37442), .dout(n37445));
  jand g20183(.dina(n37445), .dinb(n360), .dout(n37446));
  jor  g20184(.dina(n37205), .dinb(n36970), .dout(n37447));
  jxor g20185(.dina(n37053), .dinb(n37052), .dout(n37448));
  jor  g20186(.dina(n37448), .dinb(n37207), .dout(n37449));
  jand g20187(.dina(n37449), .dinb(n37447), .dout(n37450));
  jand g20188(.dina(n37450), .dinb(n363), .dout(n37451));
  jor  g20189(.dina(n37205), .dinb(n36975), .dout(n37452));
  jxor g20190(.dina(n37050), .dinb(n37049), .dout(n37453));
  jor  g20191(.dina(n37453), .dinb(n37207), .dout(n37454));
  jand g20192(.dina(n37454), .dinb(n37452), .dout(n37455));
  jand g20193(.dina(n37455), .dinb(n359), .dout(n37456));
  jor  g20194(.dina(n37205), .dinb(n36980), .dout(n37457));
  jxor g20195(.dina(n37047), .dinb(n37046), .dout(n37458));
  jor  g20196(.dina(n37458), .dinb(n37207), .dout(n37459));
  jand g20197(.dina(n37459), .dinb(n37457), .dout(n37460));
  jand g20198(.dina(n37460), .dinb(n369), .dout(n37461));
  jor  g20199(.dina(n37205), .dinb(n36985), .dout(n37462));
  jxor g20200(.dina(n37044), .dinb(n37043), .dout(n37463));
  jor  g20201(.dina(n37463), .dinb(n37207), .dout(n37464));
  jand g20202(.dina(n37464), .dinb(n37462), .dout(n37465));
  jand g20203(.dina(n37465), .dinb(n368), .dout(n37466));
  jor  g20204(.dina(n37205), .dinb(n36990), .dout(n37467));
  jxor g20205(.dina(n37041), .dinb(n37040), .dout(n37468));
  jor  g20206(.dina(n37468), .dinb(n37207), .dout(n37469));
  jand g20207(.dina(n37469), .dinb(n37467), .dout(n37470));
  jand g20208(.dina(n37470), .dinb(n367), .dout(n37471));
  jor  g20209(.dina(n37205), .dinb(n36995), .dout(n37472));
  jxor g20210(.dina(n37038), .dinb(n37037), .dout(n37473));
  jor  g20211(.dina(n37473), .dinb(n37207), .dout(n37474));
  jand g20212(.dina(n37474), .dinb(n37472), .dout(n37475));
  jand g20213(.dina(n37475), .dinb(n265), .dout(n37476));
  jor  g20214(.dina(n37205), .dinb(n37000), .dout(n37477));
  jxor g20215(.dina(n37035), .dinb(n37034), .dout(n37478));
  jor  g20216(.dina(n37478), .dinb(n37207), .dout(n37479));
  jand g20217(.dina(n37479), .dinb(n37477), .dout(n37480));
  jand g20218(.dina(n37480), .dinb(n378), .dout(n37481));
  jor  g20219(.dina(n37205), .dinb(n37005), .dout(n37482));
  jxor g20220(.dina(n37032), .dinb(n37031), .dout(n37483));
  jor  g20221(.dina(n37483), .dinb(n37207), .dout(n37484));
  jand g20222(.dina(n37484), .dinb(n37482), .dout(n37485));
  jand g20223(.dina(n37485), .dinb(n377), .dout(n37486));
  jor  g20224(.dina(n37205), .dinb(n37010), .dout(n37487));
  jxor g20225(.dina(n37029), .dinb(n37028), .dout(n37488));
  jor  g20226(.dina(n37488), .dinb(n37207), .dout(n37489));
  jand g20227(.dina(n37489), .dinb(n37487), .dout(n37490));
  jand g20228(.dina(n37490), .dinb(n376), .dout(n37491));
  jor  g20229(.dina(n37205), .dinb(n37017), .dout(n37492));
  jxor g20230(.dina(n37026), .dinb(n37025), .dout(n37493));
  jor  g20231(.dina(n37493), .dinb(n37207), .dout(n37494));
  jand g20232(.dina(n37494), .dinb(n37492), .dout(n37495));
  jand g20233(.dina(n37495), .dinb(n264), .dout(n37496));
  jor  g20234(.dina(n37205), .dinb(n37022), .dout(n37497));
  jxor g20235(.dina(n37023), .dinb(n16097), .dout(n37498));
  jand g20236(.dina(n37498), .dinb(n37205), .dout(n37499));
  jnot g20237(.din(n37499), .dout(n37500));
  jand g20238(.dina(n37500), .dinb(n37497), .dout(n37501));
  jor  g20239(.dina(n37501), .dinb(b2 ), .dout(n37502));
  jnot g20240(.din(n37502), .dout(n37503));
  jand g20241(.dina(n37205), .dinb(b0 ), .dout(n37504));
  jxor g20242(.dina(n37504), .dinb(a3 ), .dout(n37505));
  jand g20243(.dina(n37505), .dinb(n259), .dout(n37506));
  jxor g20244(.dina(n37504), .dinb(n16095), .dout(n37507));
  jxor g20245(.dina(n37507), .dinb(b1 ), .dout(n37508));
  jand g20246(.dina(n37508), .dinb(n16587), .dout(n37509));
  jor  g20247(.dina(n37509), .dinb(n37506), .dout(n37510));
  jxor g20248(.dina(n37501), .dinb(b2 ), .dout(n37511));
  jand g20249(.dina(n37511), .dinb(n37510), .dout(n37512));
  jor  g20250(.dina(n37512), .dinb(n37503), .dout(n37513));
  jxor g20251(.dina(n37495), .dinb(n264), .dout(n37514));
  jand g20252(.dina(n37514), .dinb(n37513), .dout(n37515));
  jor  g20253(.dina(n37515), .dinb(n37496), .dout(n37516));
  jxor g20254(.dina(n37490), .dinb(n376), .dout(n37517));
  jand g20255(.dina(n37517), .dinb(n37516), .dout(n37518));
  jor  g20256(.dina(n37518), .dinb(n37491), .dout(n37519));
  jxor g20257(.dina(n37485), .dinb(n377), .dout(n37520));
  jand g20258(.dina(n37520), .dinb(n37519), .dout(n37521));
  jor  g20259(.dina(n37521), .dinb(n37486), .dout(n37522));
  jxor g20260(.dina(n37480), .dinb(n378), .dout(n37523));
  jand g20261(.dina(n37523), .dinb(n37522), .dout(n37524));
  jor  g20262(.dina(n37524), .dinb(n37481), .dout(n37525));
  jxor g20263(.dina(n37475), .dinb(n265), .dout(n37526));
  jand g20264(.dina(n37526), .dinb(n37525), .dout(n37527));
  jor  g20265(.dina(n37527), .dinb(n37476), .dout(n37528));
  jxor g20266(.dina(n37470), .dinb(n367), .dout(n37529));
  jand g20267(.dina(n37529), .dinb(n37528), .dout(n37530));
  jor  g20268(.dina(n37530), .dinb(n37471), .dout(n37531));
  jxor g20269(.dina(n37465), .dinb(n368), .dout(n37532));
  jand g20270(.dina(n37532), .dinb(n37531), .dout(n37533));
  jor  g20271(.dina(n37533), .dinb(n37466), .dout(n37534));
  jxor g20272(.dina(n37460), .dinb(n369), .dout(n37535));
  jand g20273(.dina(n37535), .dinb(n37534), .dout(n37536));
  jor  g20274(.dina(n37536), .dinb(n37461), .dout(n37537));
  jxor g20275(.dina(n37455), .dinb(n359), .dout(n37538));
  jand g20276(.dina(n37538), .dinb(n37537), .dout(n37539));
  jor  g20277(.dina(n37539), .dinb(n37456), .dout(n37540));
  jxor g20278(.dina(n37450), .dinb(n363), .dout(n37541));
  jand g20279(.dina(n37541), .dinb(n37540), .dout(n37542));
  jor  g20280(.dina(n37542), .dinb(n37451), .dout(n37543));
  jxor g20281(.dina(n37445), .dinb(n360), .dout(n37544));
  jand g20282(.dina(n37544), .dinb(n37543), .dout(n37545));
  jor  g20283(.dina(n37545), .dinb(n37446), .dout(n37546));
  jxor g20284(.dina(n37440), .dinb(n361), .dout(n37547));
  jand g20285(.dina(n37547), .dinb(n37546), .dout(n37548));
  jor  g20286(.dina(n37548), .dinb(n37441), .dout(n37549));
  jxor g20287(.dina(n37435), .dinb(n364), .dout(n37550));
  jand g20288(.dina(n37550), .dinb(n37549), .dout(n37551));
  jor  g20289(.dina(n37551), .dinb(n37436), .dout(n37552));
  jxor g20290(.dina(n37430), .dinb(n355), .dout(n37553));
  jand g20291(.dina(n37553), .dinb(n37552), .dout(n37554));
  jor  g20292(.dina(n37554), .dinb(n37431), .dout(n37555));
  jxor g20293(.dina(n37425), .dinb(n356), .dout(n37556));
  jand g20294(.dina(n37556), .dinb(n37555), .dout(n37557));
  jor  g20295(.dina(n37557), .dinb(n37426), .dout(n37558));
  jxor g20296(.dina(n37420), .dinb(n266), .dout(n37559));
  jand g20297(.dina(n37559), .dinb(n37558), .dout(n37560));
  jor  g20298(.dina(n37560), .dinb(n37421), .dout(n37561));
  jxor g20299(.dina(n37415), .dinb(n267), .dout(n37562));
  jand g20300(.dina(n37562), .dinb(n37561), .dout(n37563));
  jor  g20301(.dina(n37563), .dinb(n37416), .dout(n37564));
  jxor g20302(.dina(n37410), .dinb(n347), .dout(n37565));
  jand g20303(.dina(n37565), .dinb(n37564), .dout(n37566));
  jor  g20304(.dina(n37566), .dinb(n37411), .dout(n37567));
  jxor g20305(.dina(n37405), .dinb(n348), .dout(n37568));
  jand g20306(.dina(n37568), .dinb(n37567), .dout(n37569));
  jor  g20307(.dina(n37569), .dinb(n37406), .dout(n37570));
  jxor g20308(.dina(n37400), .dinb(n349), .dout(n37571));
  jand g20309(.dina(n37571), .dinb(n37570), .dout(n37572));
  jor  g20310(.dina(n37572), .dinb(n37401), .dout(n37573));
  jxor g20311(.dina(n37395), .dinb(n268), .dout(n37574));
  jand g20312(.dina(n37574), .dinb(n37573), .dout(n37575));
  jor  g20313(.dina(n37575), .dinb(n37396), .dout(n37576));
  jxor g20314(.dina(n37390), .dinb(n274), .dout(n37577));
  jand g20315(.dina(n37577), .dinb(n37576), .dout(n37578));
  jor  g20316(.dina(n37578), .dinb(n37391), .dout(n37579));
  jxor g20317(.dina(n37385), .dinb(n269), .dout(n37580));
  jand g20318(.dina(n37580), .dinb(n37579), .dout(n37581));
  jor  g20319(.dina(n37581), .dinb(n37386), .dout(n37582));
  jxor g20320(.dina(n37380), .dinb(n270), .dout(n37583));
  jand g20321(.dina(n37583), .dinb(n37582), .dout(n37584));
  jor  g20322(.dina(n37584), .dinb(n37381), .dout(n37585));
  jxor g20323(.dina(n37375), .dinb(n271), .dout(n37586));
  jand g20324(.dina(n37586), .dinb(n37585), .dout(n37587));
  jor  g20325(.dina(n37587), .dinb(n37376), .dout(n37588));
  jxor g20326(.dina(n37370), .dinb(n338), .dout(n37589));
  jand g20327(.dina(n37589), .dinb(n37588), .dout(n37590));
  jor  g20328(.dina(n37590), .dinb(n37371), .dout(n37591));
  jxor g20329(.dina(n37365), .dinb(n339), .dout(n37592));
  jand g20330(.dina(n37592), .dinb(n37591), .dout(n37593));
  jor  g20331(.dina(n37593), .dinb(n37366), .dout(n37594));
  jxor g20332(.dina(n37360), .dinb(n340), .dout(n37595));
  jand g20333(.dina(n37595), .dinb(n37594), .dout(n37596));
  jor  g20334(.dina(n37596), .dinb(n37361), .dout(n37597));
  jxor g20335(.dina(n37355), .dinb(n275), .dout(n37598));
  jand g20336(.dina(n37598), .dinb(n37597), .dout(n37599));
  jor  g20337(.dina(n37599), .dinb(n37356), .dout(n37600));
  jxor g20338(.dina(n37350), .dinb(n331), .dout(n37601));
  jand g20339(.dina(n37601), .dinb(n37600), .dout(n37602));
  jor  g20340(.dina(n37602), .dinb(n37351), .dout(n37603));
  jxor g20341(.dina(n37345), .dinb(n332), .dout(n37604));
  jand g20342(.dina(n37604), .dinb(n37603), .dout(n37605));
  jor  g20343(.dina(n37605), .dinb(n37346), .dout(n37606));
  jxor g20344(.dina(n37340), .dinb(n333), .dout(n37607));
  jand g20345(.dina(n37607), .dinb(n37606), .dout(n37608));
  jor  g20346(.dina(n37608), .dinb(n37341), .dout(n37609));
  jxor g20347(.dina(n37335), .dinb(n276), .dout(n37610));
  jand g20348(.dina(n37610), .dinb(n37609), .dout(n37611));
  jor  g20349(.dina(n37611), .dinb(n37336), .dout(n37612));
  jxor g20350(.dina(n37330), .dinb(n324), .dout(n37613));
  jand g20351(.dina(n37613), .dinb(n37612), .dout(n37614));
  jor  g20352(.dina(n37614), .dinb(n37331), .dout(n37615));
  jxor g20353(.dina(n37325), .dinb(n325), .dout(n37616));
  jand g20354(.dina(n37616), .dinb(n37615), .dout(n37617));
  jor  g20355(.dina(n37617), .dinb(n37326), .dout(n37618));
  jxor g20356(.dina(n37320), .dinb(n326), .dout(n37619));
  jand g20357(.dina(n37619), .dinb(n37618), .dout(n37620));
  jor  g20358(.dina(n37620), .dinb(n37321), .dout(n37621));
  jxor g20359(.dina(n37315), .dinb(n277), .dout(n37622));
  jand g20360(.dina(n37622), .dinb(n37621), .dout(n37623));
  jor  g20361(.dina(n37623), .dinb(n37316), .dout(n37624));
  jxor g20362(.dina(n37310), .dinb(n278), .dout(n37625));
  jand g20363(.dina(n37625), .dinb(n37624), .dout(n37626));
  jor  g20364(.dina(n37626), .dinb(n37311), .dout(n37627));
  jxor g20365(.dina(n37305), .dinb(n279), .dout(n37628));
  jand g20366(.dina(n37628), .dinb(n37627), .dout(n37629));
  jor  g20367(.dina(n37629), .dinb(n37306), .dout(n37630));
  jxor g20368(.dina(n37300), .dinb(n280), .dout(n37631));
  jand g20369(.dina(n37631), .dinb(n37630), .dout(n37632));
  jor  g20370(.dina(n37632), .dinb(n37301), .dout(n37633));
  jxor g20371(.dina(n37295), .dinb(n283), .dout(n37634));
  jand g20372(.dina(n37634), .dinb(n37633), .dout(n37635));
  jor  g20373(.dina(n37635), .dinb(n37296), .dout(n37636));
  jxor g20374(.dina(n37290), .dinb(n315), .dout(n37637));
  jand g20375(.dina(n37637), .dinb(n37636), .dout(n37638));
  jor  g20376(.dina(n37638), .dinb(n37291), .dout(n37639));
  jxor g20377(.dina(n37285), .dinb(n316), .dout(n37640));
  jand g20378(.dina(n37640), .dinb(n37639), .dout(n37641));
  jor  g20379(.dina(n37641), .dinb(n37286), .dout(n37642));
  jxor g20380(.dina(n37280), .dinb(n317), .dout(n37643));
  jand g20381(.dina(n37643), .dinb(n37642), .dout(n37644));
  jor  g20382(.dina(n37644), .dinb(n37281), .dout(n37645));
  jxor g20383(.dina(n37275), .dinb(n284), .dout(n37646));
  jand g20384(.dina(n37646), .dinb(n37645), .dout(n37647));
  jor  g20385(.dina(n37647), .dinb(n37276), .dout(n37648));
  jxor g20386(.dina(n37270), .dinb(n285), .dout(n37649));
  jand g20387(.dina(n37649), .dinb(n37648), .dout(n37650));
  jor  g20388(.dina(n37650), .dinb(n37271), .dout(n37651));
  jxor g20389(.dina(n37265), .dinb(n286), .dout(n37652));
  jand g20390(.dina(n37652), .dinb(n37651), .dout(n37653));
  jor  g20391(.dina(n37653), .dinb(n37266), .dout(n37654));
  jxor g20392(.dina(n37260), .dinb(n287), .dout(n37655));
  jand g20393(.dina(n37655), .dinb(n37654), .dout(n37656));
  jor  g20394(.dina(n37656), .dinb(n37261), .dout(n37657));
  jxor g20395(.dina(n37255), .dinb(n288), .dout(n37658));
  jand g20396(.dina(n37658), .dinb(n37657), .dout(n37659));
  jor  g20397(.dina(n37659), .dinb(n37256), .dout(n37660));
  jxor g20398(.dina(n37250), .dinb(n289), .dout(n37661));
  jand g20399(.dina(n37661), .dinb(n37660), .dout(n37662));
  jor  g20400(.dina(n37662), .dinb(n37251), .dout(n37663));
  jxor g20401(.dina(n37245), .dinb(n290), .dout(n37664));
  jand g20402(.dina(n37664), .dinb(n37663), .dout(n37665));
  jor  g20403(.dina(n37665), .dinb(n37246), .dout(n37666));
  jxor g20404(.dina(n37240), .dinb(n291), .dout(n37667));
  jand g20405(.dina(n37667), .dinb(n37666), .dout(n37668));
  jor  g20406(.dina(n37668), .dinb(n37241), .dout(n37669));
  jxor g20407(.dina(n37235), .dinb(n292), .dout(n37670));
  jand g20408(.dina(n37670), .dinb(n37669), .dout(n37671));
  jor  g20409(.dina(n37671), .dinb(n37236), .dout(n37672));
  jxor g20410(.dina(n37230), .dinb(n293), .dout(n37673));
  jand g20411(.dina(n37673), .dinb(n37672), .dout(n37674));
  jor  g20412(.dina(n37674), .dinb(n37231), .dout(n37675));
  jxor g20413(.dina(n37225), .dinb(n294), .dout(n37676));
  jand g20414(.dina(n37676), .dinb(n37675), .dout(n37677));
  jor  g20415(.dina(n37677), .dinb(n37226), .dout(n37678));
  jxor g20416(.dina(n37220), .dinb(n295), .dout(n37679));
  jand g20417(.dina(n37679), .dinb(n37678), .dout(n37680));
  jor  g20418(.dina(n37680), .dinb(n37221), .dout(n37681));
  jxor g20419(.dina(n37215), .dinb(n296), .dout(n37682));
  jand g20420(.dina(n37682), .dinb(n37681), .dout(n37683));
  jor  g20421(.dina(n37683), .dinb(n37216), .dout(n37684));
  jxor g20422(.dina(n37210), .dinb(n297), .dout(n37685));
  jand g20423(.dina(n37685), .dinb(n37684), .dout(n37686));
  jor  g20424(.dina(n37686), .dinb(n37211), .dout(n37687));
  jand g20425(.dina(n37199), .dinb(n301), .dout(n37688));
  jor  g20426(.dina(n37688), .dinb(n37207), .dout(n37689));
  jand g20427(.dina(n37689), .dinb(n36729), .dout(n37690));
  jand g20428(.dina(n37690), .dinb(n300), .dout(n37691));
  jand g20429(.dina(n37691), .dinb(n37687), .dout(n37692));
  jnot g20430(.din(n37211), .dout(n37693));
  jnot g20431(.din(n37216), .dout(n37694));
  jnot g20432(.din(n37221), .dout(n37695));
  jnot g20433(.din(n37226), .dout(n37696));
  jnot g20434(.din(n37231), .dout(n37697));
  jnot g20435(.din(n37236), .dout(n37698));
  jnot g20436(.din(n37241), .dout(n37699));
  jnot g20437(.din(n37246), .dout(n37700));
  jnot g20438(.din(n37251), .dout(n37701));
  jnot g20439(.din(n37256), .dout(n37702));
  jnot g20440(.din(n37261), .dout(n37703));
  jnot g20441(.din(n37266), .dout(n37704));
  jnot g20442(.din(n37271), .dout(n37705));
  jnot g20443(.din(n37276), .dout(n37706));
  jnot g20444(.din(n37281), .dout(n37707));
  jnot g20445(.din(n37286), .dout(n37708));
  jnot g20446(.din(n37291), .dout(n37709));
  jnot g20447(.din(n37296), .dout(n37710));
  jnot g20448(.din(n37301), .dout(n37711));
  jnot g20449(.din(n37306), .dout(n37712));
  jnot g20450(.din(n37311), .dout(n37713));
  jnot g20451(.din(n37316), .dout(n37714));
  jnot g20452(.din(n37321), .dout(n37715));
  jnot g20453(.din(n37326), .dout(n37716));
  jnot g20454(.din(n37331), .dout(n37717));
  jnot g20455(.din(n37336), .dout(n37718));
  jnot g20456(.din(n37341), .dout(n37719));
  jnot g20457(.din(n37346), .dout(n37720));
  jnot g20458(.din(n37351), .dout(n37721));
  jnot g20459(.din(n37356), .dout(n37722));
  jnot g20460(.din(n37361), .dout(n37723));
  jnot g20461(.din(n37366), .dout(n37724));
  jnot g20462(.din(n37371), .dout(n37725));
  jnot g20463(.din(n37376), .dout(n37726));
  jnot g20464(.din(n37381), .dout(n37727));
  jnot g20465(.din(n37386), .dout(n37728));
  jnot g20466(.din(n37391), .dout(n37729));
  jnot g20467(.din(n37396), .dout(n37730));
  jnot g20468(.din(n37401), .dout(n37731));
  jnot g20469(.din(n37406), .dout(n37732));
  jnot g20470(.din(n37411), .dout(n37733));
  jnot g20471(.din(n37416), .dout(n37734));
  jnot g20472(.din(n37421), .dout(n37735));
  jnot g20473(.din(n37426), .dout(n37736));
  jnot g20474(.din(n37431), .dout(n37737));
  jnot g20475(.din(n37436), .dout(n37738));
  jnot g20476(.din(n37441), .dout(n37739));
  jnot g20477(.din(n37446), .dout(n37740));
  jnot g20478(.din(n37451), .dout(n37741));
  jnot g20479(.din(n37456), .dout(n37742));
  jnot g20480(.din(n37461), .dout(n37743));
  jnot g20481(.din(n37466), .dout(n37744));
  jnot g20482(.din(n37471), .dout(n37745));
  jnot g20483(.din(n37476), .dout(n37746));
  jnot g20484(.din(n37481), .dout(n37747));
  jnot g20485(.din(n37486), .dout(n37748));
  jnot g20486(.din(n37491), .dout(n37749));
  jnot g20487(.din(n37496), .dout(n37750));
  jnot g20488(.din(n37506), .dout(n37751));
  jxor g20489(.dina(n37507), .dinb(n259), .dout(n37752));
  jor  g20490(.dina(n37752), .dinb(n16586), .dout(n37753));
  jand g20491(.dina(n37753), .dinb(n37751), .dout(n37754));
  jnot g20492(.din(n37511), .dout(n37755));
  jor  g20493(.dina(n37755), .dinb(n37754), .dout(n37756));
  jand g20494(.dina(n37756), .dinb(n37502), .dout(n37757));
  jnot g20495(.din(n37514), .dout(n37758));
  jor  g20496(.dina(n37758), .dinb(n37757), .dout(n37759));
  jand g20497(.dina(n37759), .dinb(n37750), .dout(n37760));
  jnot g20498(.din(n37517), .dout(n37761));
  jor  g20499(.dina(n37761), .dinb(n37760), .dout(n37762));
  jand g20500(.dina(n37762), .dinb(n37749), .dout(n37763));
  jnot g20501(.din(n37520), .dout(n37764));
  jor  g20502(.dina(n37764), .dinb(n37763), .dout(n37765));
  jand g20503(.dina(n37765), .dinb(n37748), .dout(n37766));
  jnot g20504(.din(n37523), .dout(n37767));
  jor  g20505(.dina(n37767), .dinb(n37766), .dout(n37768));
  jand g20506(.dina(n37768), .dinb(n37747), .dout(n37769));
  jnot g20507(.din(n37526), .dout(n37770));
  jor  g20508(.dina(n37770), .dinb(n37769), .dout(n37771));
  jand g20509(.dina(n37771), .dinb(n37746), .dout(n37772));
  jnot g20510(.din(n37529), .dout(n37773));
  jor  g20511(.dina(n37773), .dinb(n37772), .dout(n37774));
  jand g20512(.dina(n37774), .dinb(n37745), .dout(n37775));
  jnot g20513(.din(n37532), .dout(n37776));
  jor  g20514(.dina(n37776), .dinb(n37775), .dout(n37777));
  jand g20515(.dina(n37777), .dinb(n37744), .dout(n37778));
  jnot g20516(.din(n37535), .dout(n37779));
  jor  g20517(.dina(n37779), .dinb(n37778), .dout(n37780));
  jand g20518(.dina(n37780), .dinb(n37743), .dout(n37781));
  jnot g20519(.din(n37538), .dout(n37782));
  jor  g20520(.dina(n37782), .dinb(n37781), .dout(n37783));
  jand g20521(.dina(n37783), .dinb(n37742), .dout(n37784));
  jnot g20522(.din(n37541), .dout(n37785));
  jor  g20523(.dina(n37785), .dinb(n37784), .dout(n37786));
  jand g20524(.dina(n37786), .dinb(n37741), .dout(n37787));
  jnot g20525(.din(n37544), .dout(n37788));
  jor  g20526(.dina(n37788), .dinb(n37787), .dout(n37789));
  jand g20527(.dina(n37789), .dinb(n37740), .dout(n37790));
  jnot g20528(.din(n37547), .dout(n37791));
  jor  g20529(.dina(n37791), .dinb(n37790), .dout(n37792));
  jand g20530(.dina(n37792), .dinb(n37739), .dout(n37793));
  jnot g20531(.din(n37550), .dout(n37794));
  jor  g20532(.dina(n37794), .dinb(n37793), .dout(n37795));
  jand g20533(.dina(n37795), .dinb(n37738), .dout(n37796));
  jnot g20534(.din(n37553), .dout(n37797));
  jor  g20535(.dina(n37797), .dinb(n37796), .dout(n37798));
  jand g20536(.dina(n37798), .dinb(n37737), .dout(n37799));
  jnot g20537(.din(n37556), .dout(n37800));
  jor  g20538(.dina(n37800), .dinb(n37799), .dout(n37801));
  jand g20539(.dina(n37801), .dinb(n37736), .dout(n37802));
  jnot g20540(.din(n37559), .dout(n37803));
  jor  g20541(.dina(n37803), .dinb(n37802), .dout(n37804));
  jand g20542(.dina(n37804), .dinb(n37735), .dout(n37805));
  jnot g20543(.din(n37562), .dout(n37806));
  jor  g20544(.dina(n37806), .dinb(n37805), .dout(n37807));
  jand g20545(.dina(n37807), .dinb(n37734), .dout(n37808));
  jnot g20546(.din(n37565), .dout(n37809));
  jor  g20547(.dina(n37809), .dinb(n37808), .dout(n37810));
  jand g20548(.dina(n37810), .dinb(n37733), .dout(n37811));
  jnot g20549(.din(n37568), .dout(n37812));
  jor  g20550(.dina(n37812), .dinb(n37811), .dout(n37813));
  jand g20551(.dina(n37813), .dinb(n37732), .dout(n37814));
  jnot g20552(.din(n37571), .dout(n37815));
  jor  g20553(.dina(n37815), .dinb(n37814), .dout(n37816));
  jand g20554(.dina(n37816), .dinb(n37731), .dout(n37817));
  jnot g20555(.din(n37574), .dout(n37818));
  jor  g20556(.dina(n37818), .dinb(n37817), .dout(n37819));
  jand g20557(.dina(n37819), .dinb(n37730), .dout(n37820));
  jnot g20558(.din(n37577), .dout(n37821));
  jor  g20559(.dina(n37821), .dinb(n37820), .dout(n37822));
  jand g20560(.dina(n37822), .dinb(n37729), .dout(n37823));
  jnot g20561(.din(n37580), .dout(n37824));
  jor  g20562(.dina(n37824), .dinb(n37823), .dout(n37825));
  jand g20563(.dina(n37825), .dinb(n37728), .dout(n37826));
  jnot g20564(.din(n37583), .dout(n37827));
  jor  g20565(.dina(n37827), .dinb(n37826), .dout(n37828));
  jand g20566(.dina(n37828), .dinb(n37727), .dout(n37829));
  jnot g20567(.din(n37586), .dout(n37830));
  jor  g20568(.dina(n37830), .dinb(n37829), .dout(n37831));
  jand g20569(.dina(n37831), .dinb(n37726), .dout(n37832));
  jnot g20570(.din(n37589), .dout(n37833));
  jor  g20571(.dina(n37833), .dinb(n37832), .dout(n37834));
  jand g20572(.dina(n37834), .dinb(n37725), .dout(n37835));
  jnot g20573(.din(n37592), .dout(n37836));
  jor  g20574(.dina(n37836), .dinb(n37835), .dout(n37837));
  jand g20575(.dina(n37837), .dinb(n37724), .dout(n37838));
  jnot g20576(.din(n37595), .dout(n37839));
  jor  g20577(.dina(n37839), .dinb(n37838), .dout(n37840));
  jand g20578(.dina(n37840), .dinb(n37723), .dout(n37841));
  jnot g20579(.din(n37598), .dout(n37842));
  jor  g20580(.dina(n37842), .dinb(n37841), .dout(n37843));
  jand g20581(.dina(n37843), .dinb(n37722), .dout(n37844));
  jnot g20582(.din(n37601), .dout(n37845));
  jor  g20583(.dina(n37845), .dinb(n37844), .dout(n37846));
  jand g20584(.dina(n37846), .dinb(n37721), .dout(n37847));
  jnot g20585(.din(n37604), .dout(n37848));
  jor  g20586(.dina(n37848), .dinb(n37847), .dout(n37849));
  jand g20587(.dina(n37849), .dinb(n37720), .dout(n37850));
  jnot g20588(.din(n37607), .dout(n37851));
  jor  g20589(.dina(n37851), .dinb(n37850), .dout(n37852));
  jand g20590(.dina(n37852), .dinb(n37719), .dout(n37853));
  jnot g20591(.din(n37610), .dout(n37854));
  jor  g20592(.dina(n37854), .dinb(n37853), .dout(n37855));
  jand g20593(.dina(n37855), .dinb(n37718), .dout(n37856));
  jnot g20594(.din(n37613), .dout(n37857));
  jor  g20595(.dina(n37857), .dinb(n37856), .dout(n37858));
  jand g20596(.dina(n37858), .dinb(n37717), .dout(n37859));
  jnot g20597(.din(n37616), .dout(n37860));
  jor  g20598(.dina(n37860), .dinb(n37859), .dout(n37861));
  jand g20599(.dina(n37861), .dinb(n37716), .dout(n37862));
  jnot g20600(.din(n37619), .dout(n37863));
  jor  g20601(.dina(n37863), .dinb(n37862), .dout(n37864));
  jand g20602(.dina(n37864), .dinb(n37715), .dout(n37865));
  jnot g20603(.din(n37622), .dout(n37866));
  jor  g20604(.dina(n37866), .dinb(n37865), .dout(n37867));
  jand g20605(.dina(n37867), .dinb(n37714), .dout(n37868));
  jnot g20606(.din(n37625), .dout(n37869));
  jor  g20607(.dina(n37869), .dinb(n37868), .dout(n37870));
  jand g20608(.dina(n37870), .dinb(n37713), .dout(n37871));
  jnot g20609(.din(n37628), .dout(n37872));
  jor  g20610(.dina(n37872), .dinb(n37871), .dout(n37873));
  jand g20611(.dina(n37873), .dinb(n37712), .dout(n37874));
  jnot g20612(.din(n37631), .dout(n37875));
  jor  g20613(.dina(n37875), .dinb(n37874), .dout(n37876));
  jand g20614(.dina(n37876), .dinb(n37711), .dout(n37877));
  jnot g20615(.din(n37634), .dout(n37878));
  jor  g20616(.dina(n37878), .dinb(n37877), .dout(n37879));
  jand g20617(.dina(n37879), .dinb(n37710), .dout(n37880));
  jnot g20618(.din(n37637), .dout(n37881));
  jor  g20619(.dina(n37881), .dinb(n37880), .dout(n37882));
  jand g20620(.dina(n37882), .dinb(n37709), .dout(n37883));
  jnot g20621(.din(n37640), .dout(n37884));
  jor  g20622(.dina(n37884), .dinb(n37883), .dout(n37885));
  jand g20623(.dina(n37885), .dinb(n37708), .dout(n37886));
  jnot g20624(.din(n37643), .dout(n37887));
  jor  g20625(.dina(n37887), .dinb(n37886), .dout(n37888));
  jand g20626(.dina(n37888), .dinb(n37707), .dout(n37889));
  jnot g20627(.din(n37646), .dout(n37890));
  jor  g20628(.dina(n37890), .dinb(n37889), .dout(n37891));
  jand g20629(.dina(n37891), .dinb(n37706), .dout(n37892));
  jnot g20630(.din(n37649), .dout(n37893));
  jor  g20631(.dina(n37893), .dinb(n37892), .dout(n37894));
  jand g20632(.dina(n37894), .dinb(n37705), .dout(n37895));
  jnot g20633(.din(n37652), .dout(n37896));
  jor  g20634(.dina(n37896), .dinb(n37895), .dout(n37897));
  jand g20635(.dina(n37897), .dinb(n37704), .dout(n37898));
  jnot g20636(.din(n37655), .dout(n37899));
  jor  g20637(.dina(n37899), .dinb(n37898), .dout(n37900));
  jand g20638(.dina(n37900), .dinb(n37703), .dout(n37901));
  jnot g20639(.din(n37658), .dout(n37902));
  jor  g20640(.dina(n37902), .dinb(n37901), .dout(n37903));
  jand g20641(.dina(n37903), .dinb(n37702), .dout(n37904));
  jnot g20642(.din(n37661), .dout(n37905));
  jor  g20643(.dina(n37905), .dinb(n37904), .dout(n37906));
  jand g20644(.dina(n37906), .dinb(n37701), .dout(n37907));
  jnot g20645(.din(n37664), .dout(n37908));
  jor  g20646(.dina(n37908), .dinb(n37907), .dout(n37909));
  jand g20647(.dina(n37909), .dinb(n37700), .dout(n37910));
  jnot g20648(.din(n37667), .dout(n37911));
  jor  g20649(.dina(n37911), .dinb(n37910), .dout(n37912));
  jand g20650(.dina(n37912), .dinb(n37699), .dout(n37913));
  jnot g20651(.din(n37670), .dout(n37914));
  jor  g20652(.dina(n37914), .dinb(n37913), .dout(n37915));
  jand g20653(.dina(n37915), .dinb(n37698), .dout(n37916));
  jnot g20654(.din(n37673), .dout(n37917));
  jor  g20655(.dina(n37917), .dinb(n37916), .dout(n37918));
  jand g20656(.dina(n37918), .dinb(n37697), .dout(n37919));
  jnot g20657(.din(n37676), .dout(n37920));
  jor  g20658(.dina(n37920), .dinb(n37919), .dout(n37921));
  jand g20659(.dina(n37921), .dinb(n37696), .dout(n37922));
  jnot g20660(.din(n37679), .dout(n37923));
  jor  g20661(.dina(n37923), .dinb(n37922), .dout(n37924));
  jand g20662(.dina(n37924), .dinb(n37695), .dout(n37925));
  jnot g20663(.din(n37682), .dout(n37926));
  jor  g20664(.dina(n37926), .dinb(n37925), .dout(n37927));
  jand g20665(.dina(n37927), .dinb(n37694), .dout(n37928));
  jnot g20666(.din(n37685), .dout(n37929));
  jor  g20667(.dina(n37929), .dinb(n37928), .dout(n37930));
  jand g20668(.dina(n37930), .dinb(n37693), .dout(n37931));
  jor  g20669(.dina(n37931), .dinb(n830), .dout(n37932));
  jand g20670(.dina(n36729), .dinb(n831), .dout(n37933));
  jand g20671(.dina(n37933), .dinb(n37932), .dout(n37934));
  jor  g20672(.dina(n37934), .dinb(n37692), .dout(n37935));
  jand g20673(.dina(n37935), .dinb(n298), .dout(n37936));
  jor  g20674(.dina(n37690), .dinb(n257), .dout(n37937));
  jand g20675(.dina(n37687), .dinb(n299), .dout(n37938));
  jor  g20676(.dina(n37938), .dinb(n37691), .dout(n37939));
  jand g20677(.dina(n37939), .dinb(n37937), .dout(n37940));
  jor  g20678(.dina(n37940), .dinb(n37210), .dout(n37941));
  jnot g20679(.din(n37937), .dout(n37942));
  jnot g20680(.din(n37691), .dout(n37943));
  jand g20681(.dina(n37932), .dinb(n37943), .dout(n37944));
  jor  g20682(.dina(n37944), .dinb(n37942), .dout(n37945));
  jxor g20683(.dina(n37685), .dinb(n37684), .dout(n37946));
  jor  g20684(.dina(n37946), .dinb(n37945), .dout(n37947));
  jand g20685(.dina(n37947), .dinb(n37941), .dout(n37948));
  jand g20686(.dina(n37948), .dinb(n257), .dout(n37949));
  jor  g20687(.dina(n37940), .dinb(n37215), .dout(n37950));
  jxor g20688(.dina(n37682), .dinb(n37681), .dout(n37951));
  jor  g20689(.dina(n37951), .dinb(n37945), .dout(n37952));
  jand g20690(.dina(n37952), .dinb(n37950), .dout(n37953));
  jand g20691(.dina(n37953), .dinb(n297), .dout(n37954));
  jor  g20692(.dina(n37940), .dinb(n37220), .dout(n37955));
  jxor g20693(.dina(n37679), .dinb(n37678), .dout(n37956));
  jor  g20694(.dina(n37956), .dinb(n37945), .dout(n37957));
  jand g20695(.dina(n37957), .dinb(n37955), .dout(n37958));
  jand g20696(.dina(n37958), .dinb(n296), .dout(n37959));
  jor  g20697(.dina(n37940), .dinb(n37225), .dout(n37960));
  jxor g20698(.dina(n37676), .dinb(n37675), .dout(n37961));
  jor  g20699(.dina(n37961), .dinb(n37945), .dout(n37962));
  jand g20700(.dina(n37962), .dinb(n37960), .dout(n37963));
  jand g20701(.dina(n37963), .dinb(n295), .dout(n37964));
  jor  g20702(.dina(n37940), .dinb(n37230), .dout(n37965));
  jxor g20703(.dina(n37673), .dinb(n37672), .dout(n37966));
  jor  g20704(.dina(n37966), .dinb(n37945), .dout(n37967));
  jand g20705(.dina(n37967), .dinb(n37965), .dout(n37968));
  jand g20706(.dina(n37968), .dinb(n294), .dout(n37969));
  jor  g20707(.dina(n37940), .dinb(n37235), .dout(n37970));
  jxor g20708(.dina(n37670), .dinb(n37669), .dout(n37971));
  jor  g20709(.dina(n37971), .dinb(n37945), .dout(n37972));
  jand g20710(.dina(n37972), .dinb(n37970), .dout(n37973));
  jand g20711(.dina(n37973), .dinb(n293), .dout(n37974));
  jor  g20712(.dina(n37940), .dinb(n37240), .dout(n37975));
  jxor g20713(.dina(n37667), .dinb(n37666), .dout(n37976));
  jor  g20714(.dina(n37976), .dinb(n37945), .dout(n37977));
  jand g20715(.dina(n37977), .dinb(n37975), .dout(n37978));
  jand g20716(.dina(n37978), .dinb(n292), .dout(n37979));
  jor  g20717(.dina(n37940), .dinb(n37245), .dout(n37980));
  jxor g20718(.dina(n37664), .dinb(n37663), .dout(n37981));
  jor  g20719(.dina(n37981), .dinb(n37945), .dout(n37982));
  jand g20720(.dina(n37982), .dinb(n37980), .dout(n37983));
  jand g20721(.dina(n37983), .dinb(n291), .dout(n37984));
  jor  g20722(.dina(n37940), .dinb(n37250), .dout(n37985));
  jxor g20723(.dina(n37661), .dinb(n37660), .dout(n37986));
  jor  g20724(.dina(n37986), .dinb(n37945), .dout(n37987));
  jand g20725(.dina(n37987), .dinb(n37985), .dout(n37988));
  jand g20726(.dina(n37988), .dinb(n290), .dout(n37989));
  jor  g20727(.dina(n37940), .dinb(n37255), .dout(n37990));
  jxor g20728(.dina(n37658), .dinb(n37657), .dout(n37991));
  jor  g20729(.dina(n37991), .dinb(n37945), .dout(n37992));
  jand g20730(.dina(n37992), .dinb(n37990), .dout(n37993));
  jand g20731(.dina(n37993), .dinb(n289), .dout(n37994));
  jor  g20732(.dina(n37940), .dinb(n37260), .dout(n37995));
  jxor g20733(.dina(n37655), .dinb(n37654), .dout(n37996));
  jor  g20734(.dina(n37996), .dinb(n37945), .dout(n37997));
  jand g20735(.dina(n37997), .dinb(n37995), .dout(n37998));
  jand g20736(.dina(n37998), .dinb(n288), .dout(n37999));
  jor  g20737(.dina(n37940), .dinb(n37265), .dout(n38000));
  jxor g20738(.dina(n37652), .dinb(n37651), .dout(n38001));
  jor  g20739(.dina(n38001), .dinb(n37945), .dout(n38002));
  jand g20740(.dina(n38002), .dinb(n38000), .dout(n38003));
  jand g20741(.dina(n38003), .dinb(n287), .dout(n38004));
  jor  g20742(.dina(n37940), .dinb(n37270), .dout(n38005));
  jxor g20743(.dina(n37649), .dinb(n37648), .dout(n38006));
  jor  g20744(.dina(n38006), .dinb(n37945), .dout(n38007));
  jand g20745(.dina(n38007), .dinb(n38005), .dout(n38008));
  jand g20746(.dina(n38008), .dinb(n286), .dout(n38009));
  jor  g20747(.dina(n37940), .dinb(n37275), .dout(n38010));
  jxor g20748(.dina(n37646), .dinb(n37645), .dout(n38011));
  jor  g20749(.dina(n38011), .dinb(n37945), .dout(n38012));
  jand g20750(.dina(n38012), .dinb(n38010), .dout(n38013));
  jand g20751(.dina(n38013), .dinb(n285), .dout(n38014));
  jor  g20752(.dina(n37940), .dinb(n37280), .dout(n38015));
  jxor g20753(.dina(n37643), .dinb(n37642), .dout(n38016));
  jor  g20754(.dina(n38016), .dinb(n37945), .dout(n38017));
  jand g20755(.dina(n38017), .dinb(n38015), .dout(n38018));
  jand g20756(.dina(n38018), .dinb(n284), .dout(n38019));
  jor  g20757(.dina(n37940), .dinb(n37285), .dout(n38020));
  jxor g20758(.dina(n37640), .dinb(n37639), .dout(n38021));
  jor  g20759(.dina(n38021), .dinb(n37945), .dout(n38022));
  jand g20760(.dina(n38022), .dinb(n38020), .dout(n38023));
  jand g20761(.dina(n38023), .dinb(n317), .dout(n38024));
  jor  g20762(.dina(n37940), .dinb(n37290), .dout(n38025));
  jxor g20763(.dina(n37637), .dinb(n37636), .dout(n38026));
  jor  g20764(.dina(n38026), .dinb(n37945), .dout(n38027));
  jand g20765(.dina(n38027), .dinb(n38025), .dout(n38028));
  jand g20766(.dina(n38028), .dinb(n316), .dout(n38029));
  jor  g20767(.dina(n37940), .dinb(n37295), .dout(n38030));
  jxor g20768(.dina(n37634), .dinb(n37633), .dout(n38031));
  jor  g20769(.dina(n38031), .dinb(n37945), .dout(n38032));
  jand g20770(.dina(n38032), .dinb(n38030), .dout(n38033));
  jand g20771(.dina(n38033), .dinb(n315), .dout(n38034));
  jor  g20772(.dina(n37940), .dinb(n37300), .dout(n38035));
  jxor g20773(.dina(n37631), .dinb(n37630), .dout(n38036));
  jor  g20774(.dina(n38036), .dinb(n37945), .dout(n38037));
  jand g20775(.dina(n38037), .dinb(n38035), .dout(n38038));
  jand g20776(.dina(n38038), .dinb(n283), .dout(n38039));
  jor  g20777(.dina(n37940), .dinb(n37305), .dout(n38040));
  jxor g20778(.dina(n37628), .dinb(n37627), .dout(n38041));
  jor  g20779(.dina(n38041), .dinb(n37945), .dout(n38042));
  jand g20780(.dina(n38042), .dinb(n38040), .dout(n38043));
  jand g20781(.dina(n38043), .dinb(n280), .dout(n38044));
  jor  g20782(.dina(n37940), .dinb(n37310), .dout(n38045));
  jxor g20783(.dina(n37625), .dinb(n37624), .dout(n38046));
  jor  g20784(.dina(n38046), .dinb(n37945), .dout(n38047));
  jand g20785(.dina(n38047), .dinb(n38045), .dout(n38048));
  jand g20786(.dina(n38048), .dinb(n279), .dout(n38049));
  jor  g20787(.dina(n37940), .dinb(n37315), .dout(n38050));
  jxor g20788(.dina(n37622), .dinb(n37621), .dout(n38051));
  jor  g20789(.dina(n38051), .dinb(n37945), .dout(n38052));
  jand g20790(.dina(n38052), .dinb(n38050), .dout(n38053));
  jand g20791(.dina(n38053), .dinb(n278), .dout(n38054));
  jor  g20792(.dina(n37940), .dinb(n37320), .dout(n38055));
  jxor g20793(.dina(n37619), .dinb(n37618), .dout(n38056));
  jor  g20794(.dina(n38056), .dinb(n37945), .dout(n38057));
  jand g20795(.dina(n38057), .dinb(n38055), .dout(n38058));
  jand g20796(.dina(n38058), .dinb(n277), .dout(n38059));
  jor  g20797(.dina(n37940), .dinb(n37325), .dout(n38060));
  jxor g20798(.dina(n37616), .dinb(n37615), .dout(n38061));
  jor  g20799(.dina(n38061), .dinb(n37945), .dout(n38062));
  jand g20800(.dina(n38062), .dinb(n38060), .dout(n38063));
  jand g20801(.dina(n38063), .dinb(n326), .dout(n38064));
  jor  g20802(.dina(n37940), .dinb(n37330), .dout(n38065));
  jxor g20803(.dina(n37613), .dinb(n37612), .dout(n38066));
  jor  g20804(.dina(n38066), .dinb(n37945), .dout(n38067));
  jand g20805(.dina(n38067), .dinb(n38065), .dout(n38068));
  jand g20806(.dina(n38068), .dinb(n325), .dout(n38069));
  jor  g20807(.dina(n37940), .dinb(n37335), .dout(n38070));
  jxor g20808(.dina(n37610), .dinb(n37609), .dout(n38071));
  jor  g20809(.dina(n38071), .dinb(n37945), .dout(n38072));
  jand g20810(.dina(n38072), .dinb(n38070), .dout(n38073));
  jand g20811(.dina(n38073), .dinb(n324), .dout(n38074));
  jor  g20812(.dina(n37940), .dinb(n37340), .dout(n38075));
  jxor g20813(.dina(n37607), .dinb(n37606), .dout(n38076));
  jor  g20814(.dina(n38076), .dinb(n37945), .dout(n38077));
  jand g20815(.dina(n38077), .dinb(n38075), .dout(n38078));
  jand g20816(.dina(n38078), .dinb(n276), .dout(n38079));
  jor  g20817(.dina(n37940), .dinb(n37345), .dout(n38080));
  jxor g20818(.dina(n37604), .dinb(n37603), .dout(n38081));
  jor  g20819(.dina(n38081), .dinb(n37945), .dout(n38082));
  jand g20820(.dina(n38082), .dinb(n38080), .dout(n38083));
  jand g20821(.dina(n38083), .dinb(n333), .dout(n38084));
  jor  g20822(.dina(n37940), .dinb(n37350), .dout(n38085));
  jxor g20823(.dina(n37601), .dinb(n37600), .dout(n38086));
  jor  g20824(.dina(n38086), .dinb(n37945), .dout(n38087));
  jand g20825(.dina(n38087), .dinb(n38085), .dout(n38088));
  jand g20826(.dina(n38088), .dinb(n332), .dout(n38089));
  jor  g20827(.dina(n37940), .dinb(n37355), .dout(n38090));
  jxor g20828(.dina(n37598), .dinb(n37597), .dout(n38091));
  jor  g20829(.dina(n38091), .dinb(n37945), .dout(n38092));
  jand g20830(.dina(n38092), .dinb(n38090), .dout(n38093));
  jand g20831(.dina(n38093), .dinb(n331), .dout(n38094));
  jor  g20832(.dina(n37940), .dinb(n37360), .dout(n38095));
  jxor g20833(.dina(n37595), .dinb(n37594), .dout(n38096));
  jor  g20834(.dina(n38096), .dinb(n37945), .dout(n38097));
  jand g20835(.dina(n38097), .dinb(n38095), .dout(n38098));
  jand g20836(.dina(n38098), .dinb(n275), .dout(n38099));
  jor  g20837(.dina(n37940), .dinb(n37365), .dout(n38100));
  jxor g20838(.dina(n37592), .dinb(n37591), .dout(n38101));
  jor  g20839(.dina(n38101), .dinb(n37945), .dout(n38102));
  jand g20840(.dina(n38102), .dinb(n38100), .dout(n38103));
  jand g20841(.dina(n38103), .dinb(n340), .dout(n38104));
  jor  g20842(.dina(n37940), .dinb(n37370), .dout(n38105));
  jxor g20843(.dina(n37589), .dinb(n37588), .dout(n38106));
  jor  g20844(.dina(n38106), .dinb(n37945), .dout(n38107));
  jand g20845(.dina(n38107), .dinb(n38105), .dout(n38108));
  jand g20846(.dina(n38108), .dinb(n339), .dout(n38109));
  jor  g20847(.dina(n37940), .dinb(n37375), .dout(n38110));
  jxor g20848(.dina(n37586), .dinb(n37585), .dout(n38111));
  jor  g20849(.dina(n38111), .dinb(n37945), .dout(n38112));
  jand g20850(.dina(n38112), .dinb(n38110), .dout(n38113));
  jand g20851(.dina(n38113), .dinb(n338), .dout(n38114));
  jor  g20852(.dina(n37940), .dinb(n37380), .dout(n38115));
  jxor g20853(.dina(n37583), .dinb(n37582), .dout(n38116));
  jor  g20854(.dina(n38116), .dinb(n37945), .dout(n38117));
  jand g20855(.dina(n38117), .dinb(n38115), .dout(n38118));
  jand g20856(.dina(n38118), .dinb(n271), .dout(n38119));
  jor  g20857(.dina(n37940), .dinb(n37385), .dout(n38120));
  jxor g20858(.dina(n37580), .dinb(n37579), .dout(n38121));
  jor  g20859(.dina(n38121), .dinb(n37945), .dout(n38122));
  jand g20860(.dina(n38122), .dinb(n38120), .dout(n38123));
  jand g20861(.dina(n38123), .dinb(n270), .dout(n38124));
  jor  g20862(.dina(n37940), .dinb(n37390), .dout(n38125));
  jxor g20863(.dina(n37577), .dinb(n37576), .dout(n38126));
  jor  g20864(.dina(n38126), .dinb(n37945), .dout(n38127));
  jand g20865(.dina(n38127), .dinb(n38125), .dout(n38128));
  jand g20866(.dina(n38128), .dinb(n269), .dout(n38129));
  jor  g20867(.dina(n37940), .dinb(n37395), .dout(n38130));
  jxor g20868(.dina(n37574), .dinb(n37573), .dout(n38131));
  jor  g20869(.dina(n38131), .dinb(n37945), .dout(n38132));
  jand g20870(.dina(n38132), .dinb(n38130), .dout(n38133));
  jand g20871(.dina(n38133), .dinb(n274), .dout(n38134));
  jor  g20872(.dina(n37940), .dinb(n37400), .dout(n38135));
  jxor g20873(.dina(n37571), .dinb(n37570), .dout(n38136));
  jor  g20874(.dina(n38136), .dinb(n37945), .dout(n38137));
  jand g20875(.dina(n38137), .dinb(n38135), .dout(n38138));
  jand g20876(.dina(n38138), .dinb(n268), .dout(n38139));
  jor  g20877(.dina(n37940), .dinb(n37405), .dout(n38140));
  jxor g20878(.dina(n37568), .dinb(n37567), .dout(n38141));
  jor  g20879(.dina(n38141), .dinb(n37945), .dout(n38142));
  jand g20880(.dina(n38142), .dinb(n38140), .dout(n38143));
  jand g20881(.dina(n38143), .dinb(n349), .dout(n38144));
  jor  g20882(.dina(n37940), .dinb(n37410), .dout(n38145));
  jxor g20883(.dina(n37565), .dinb(n37564), .dout(n38146));
  jor  g20884(.dina(n38146), .dinb(n37945), .dout(n38147));
  jand g20885(.dina(n38147), .dinb(n38145), .dout(n38148));
  jand g20886(.dina(n38148), .dinb(n348), .dout(n38149));
  jor  g20887(.dina(n37940), .dinb(n37415), .dout(n38150));
  jxor g20888(.dina(n37562), .dinb(n37561), .dout(n38151));
  jor  g20889(.dina(n38151), .dinb(n37945), .dout(n38152));
  jand g20890(.dina(n38152), .dinb(n38150), .dout(n38153));
  jand g20891(.dina(n38153), .dinb(n347), .dout(n38154));
  jor  g20892(.dina(n37940), .dinb(n37420), .dout(n38155));
  jxor g20893(.dina(n37559), .dinb(n37558), .dout(n38156));
  jor  g20894(.dina(n38156), .dinb(n37945), .dout(n38157));
  jand g20895(.dina(n38157), .dinb(n38155), .dout(n38158));
  jand g20896(.dina(n38158), .dinb(n267), .dout(n38159));
  jor  g20897(.dina(n37940), .dinb(n37425), .dout(n38160));
  jxor g20898(.dina(n37556), .dinb(n37555), .dout(n38161));
  jor  g20899(.dina(n38161), .dinb(n37945), .dout(n38162));
  jand g20900(.dina(n38162), .dinb(n38160), .dout(n38163));
  jand g20901(.dina(n38163), .dinb(n266), .dout(n38164));
  jor  g20902(.dina(n37940), .dinb(n37430), .dout(n38165));
  jxor g20903(.dina(n37553), .dinb(n37552), .dout(n38166));
  jor  g20904(.dina(n38166), .dinb(n37945), .dout(n38167));
  jand g20905(.dina(n38167), .dinb(n38165), .dout(n38168));
  jand g20906(.dina(n38168), .dinb(n356), .dout(n38169));
  jor  g20907(.dina(n37940), .dinb(n37435), .dout(n38170));
  jxor g20908(.dina(n37550), .dinb(n37549), .dout(n38171));
  jor  g20909(.dina(n38171), .dinb(n37945), .dout(n38172));
  jand g20910(.dina(n38172), .dinb(n38170), .dout(n38173));
  jand g20911(.dina(n38173), .dinb(n355), .dout(n38174));
  jor  g20912(.dina(n37940), .dinb(n37440), .dout(n38175));
  jxor g20913(.dina(n37547), .dinb(n37546), .dout(n38176));
  jor  g20914(.dina(n38176), .dinb(n37945), .dout(n38177));
  jand g20915(.dina(n38177), .dinb(n38175), .dout(n38178));
  jand g20916(.dina(n38178), .dinb(n364), .dout(n38179));
  jor  g20917(.dina(n37940), .dinb(n37445), .dout(n38180));
  jxor g20918(.dina(n37544), .dinb(n37543), .dout(n38181));
  jor  g20919(.dina(n38181), .dinb(n37945), .dout(n38182));
  jand g20920(.dina(n38182), .dinb(n38180), .dout(n38183));
  jand g20921(.dina(n38183), .dinb(n361), .dout(n38184));
  jor  g20922(.dina(n37940), .dinb(n37450), .dout(n38185));
  jxor g20923(.dina(n37541), .dinb(n37540), .dout(n38186));
  jor  g20924(.dina(n38186), .dinb(n37945), .dout(n38187));
  jand g20925(.dina(n38187), .dinb(n38185), .dout(n38188));
  jand g20926(.dina(n38188), .dinb(n360), .dout(n38189));
  jor  g20927(.dina(n37940), .dinb(n37455), .dout(n38190));
  jxor g20928(.dina(n37538), .dinb(n37537), .dout(n38191));
  jor  g20929(.dina(n38191), .dinb(n37945), .dout(n38192));
  jand g20930(.dina(n38192), .dinb(n38190), .dout(n38193));
  jand g20931(.dina(n38193), .dinb(n363), .dout(n38194));
  jor  g20932(.dina(n37940), .dinb(n37460), .dout(n38195));
  jxor g20933(.dina(n37535), .dinb(n37534), .dout(n38196));
  jor  g20934(.dina(n38196), .dinb(n37945), .dout(n38197));
  jand g20935(.dina(n38197), .dinb(n38195), .dout(n38198));
  jand g20936(.dina(n38198), .dinb(n359), .dout(n38199));
  jor  g20937(.dina(n37940), .dinb(n37465), .dout(n38200));
  jxor g20938(.dina(n37532), .dinb(n37531), .dout(n38201));
  jor  g20939(.dina(n38201), .dinb(n37945), .dout(n38202));
  jand g20940(.dina(n38202), .dinb(n38200), .dout(n38203));
  jand g20941(.dina(n38203), .dinb(n369), .dout(n38204));
  jor  g20942(.dina(n37940), .dinb(n37470), .dout(n38205));
  jxor g20943(.dina(n37529), .dinb(n37528), .dout(n38206));
  jor  g20944(.dina(n38206), .dinb(n37945), .dout(n38207));
  jand g20945(.dina(n38207), .dinb(n38205), .dout(n38208));
  jand g20946(.dina(n38208), .dinb(n368), .dout(n38209));
  jor  g20947(.dina(n37940), .dinb(n37475), .dout(n38210));
  jxor g20948(.dina(n37526), .dinb(n37525), .dout(n38211));
  jor  g20949(.dina(n38211), .dinb(n37945), .dout(n38212));
  jand g20950(.dina(n38212), .dinb(n38210), .dout(n38213));
  jand g20951(.dina(n38213), .dinb(n367), .dout(n38214));
  jor  g20952(.dina(n37940), .dinb(n37480), .dout(n38215));
  jxor g20953(.dina(n37523), .dinb(n37522), .dout(n38216));
  jor  g20954(.dina(n38216), .dinb(n37945), .dout(n38217));
  jand g20955(.dina(n38217), .dinb(n38215), .dout(n38218));
  jand g20956(.dina(n38218), .dinb(n265), .dout(n38219));
  jor  g20957(.dina(n37940), .dinb(n37485), .dout(n38220));
  jxor g20958(.dina(n37520), .dinb(n37519), .dout(n38221));
  jor  g20959(.dina(n38221), .dinb(n37945), .dout(n38222));
  jand g20960(.dina(n38222), .dinb(n38220), .dout(n38223));
  jand g20961(.dina(n38223), .dinb(n378), .dout(n38224));
  jor  g20962(.dina(n37940), .dinb(n37490), .dout(n38225));
  jxor g20963(.dina(n37517), .dinb(n37516), .dout(n38226));
  jor  g20964(.dina(n38226), .dinb(n37945), .dout(n38227));
  jand g20965(.dina(n38227), .dinb(n38225), .dout(n38228));
  jand g20966(.dina(n38228), .dinb(n377), .dout(n38229));
  jor  g20967(.dina(n37940), .dinb(n37495), .dout(n38230));
  jxor g20968(.dina(n37514), .dinb(n37513), .dout(n38231));
  jor  g20969(.dina(n38231), .dinb(n37945), .dout(n38232));
  jand g20970(.dina(n38232), .dinb(n38230), .dout(n38233));
  jand g20971(.dina(n38233), .dinb(n376), .dout(n38234));
  jand g20972(.dina(n37945), .dinb(n37501), .dout(n38235));
  jnot g20973(.din(n38235), .dout(n38236));
  jxor g20974(.dina(n37511), .dinb(n37510), .dout(n38237));
  jor  g20975(.dina(n38237), .dinb(n37945), .dout(n38238));
  jand g20976(.dina(n38238), .dinb(n38236), .dout(n38239));
  jand g20977(.dina(n38239), .dinb(n264), .dout(n38240));
  jxor g20978(.dina(n37508), .dinb(n16587), .dout(n38241));
  jand g20979(.dina(n38241), .dinb(n37940), .dout(n38242));
  jand g20980(.dina(n37945), .dinb(n37505), .dout(n38243));
  jor  g20981(.dina(n38243), .dinb(n38242), .dout(n38244));
  jand g20982(.dina(n38244), .dinb(n386), .dout(n38245));
  jor  g20983(.dina(n37945), .dinb(n17822), .dout(n38246));
  jand g20984(.dina(n38246), .dinb(a2 ), .dout(n38247));
  jor  g20985(.dina(n37945), .dinb(n16587), .dout(n38248));
  jnot g20986(.din(n38248), .dout(n38249));
  jor  g20987(.dina(n38249), .dinb(n38247), .dout(n38250));
  jand g20988(.dina(n38250), .dinb(n259), .dout(n38251));
  jand g20989(.dina(n37940), .dinb(b0 ), .dout(n38252));
  jor  g20990(.dina(n38252), .dinb(n16585), .dout(n38253));
  jand g20991(.dina(n38248), .dinb(n38253), .dout(n38254));
  jxor g20992(.dina(n38254), .dinb(b1 ), .dout(n38255));
  jand g20993(.dina(n38255), .dinb(n17079), .dout(n38256));
  jor  g20994(.dina(n38256), .dinb(n38251), .dout(n38257));
  jxor g20995(.dina(n38244), .dinb(n386), .dout(n38258));
  jand g20996(.dina(n38258), .dinb(n38257), .dout(n38259));
  jor  g20997(.dina(n38259), .dinb(n38245), .dout(n38260));
  jxor g20998(.dina(n38239), .dinb(n264), .dout(n38261));
  jand g20999(.dina(n38261), .dinb(n38260), .dout(n38262));
  jor  g21000(.dina(n38262), .dinb(n38240), .dout(n38263));
  jxor g21001(.dina(n38233), .dinb(n376), .dout(n38264));
  jand g21002(.dina(n38264), .dinb(n38263), .dout(n38265));
  jor  g21003(.dina(n38265), .dinb(n38234), .dout(n38266));
  jxor g21004(.dina(n38228), .dinb(n377), .dout(n38267));
  jand g21005(.dina(n38267), .dinb(n38266), .dout(n38268));
  jor  g21006(.dina(n38268), .dinb(n38229), .dout(n38269));
  jxor g21007(.dina(n38223), .dinb(n378), .dout(n38270));
  jand g21008(.dina(n38270), .dinb(n38269), .dout(n38271));
  jor  g21009(.dina(n38271), .dinb(n38224), .dout(n38272));
  jxor g21010(.dina(n38218), .dinb(n265), .dout(n38273));
  jand g21011(.dina(n38273), .dinb(n38272), .dout(n38274));
  jor  g21012(.dina(n38274), .dinb(n38219), .dout(n38275));
  jxor g21013(.dina(n38213), .dinb(n367), .dout(n38276));
  jand g21014(.dina(n38276), .dinb(n38275), .dout(n38277));
  jor  g21015(.dina(n38277), .dinb(n38214), .dout(n38278));
  jxor g21016(.dina(n38208), .dinb(n368), .dout(n38279));
  jand g21017(.dina(n38279), .dinb(n38278), .dout(n38280));
  jor  g21018(.dina(n38280), .dinb(n38209), .dout(n38281));
  jxor g21019(.dina(n38203), .dinb(n369), .dout(n38282));
  jand g21020(.dina(n38282), .dinb(n38281), .dout(n38283));
  jor  g21021(.dina(n38283), .dinb(n38204), .dout(n38284));
  jxor g21022(.dina(n38198), .dinb(n359), .dout(n38285));
  jand g21023(.dina(n38285), .dinb(n38284), .dout(n38286));
  jor  g21024(.dina(n38286), .dinb(n38199), .dout(n38287));
  jxor g21025(.dina(n38193), .dinb(n363), .dout(n38288));
  jand g21026(.dina(n38288), .dinb(n38287), .dout(n38289));
  jor  g21027(.dina(n38289), .dinb(n38194), .dout(n38290));
  jxor g21028(.dina(n38188), .dinb(n360), .dout(n38291));
  jand g21029(.dina(n38291), .dinb(n38290), .dout(n38292));
  jor  g21030(.dina(n38292), .dinb(n38189), .dout(n38293));
  jxor g21031(.dina(n38183), .dinb(n361), .dout(n38294));
  jand g21032(.dina(n38294), .dinb(n38293), .dout(n38295));
  jor  g21033(.dina(n38295), .dinb(n38184), .dout(n38296));
  jxor g21034(.dina(n38178), .dinb(n364), .dout(n38297));
  jand g21035(.dina(n38297), .dinb(n38296), .dout(n38298));
  jor  g21036(.dina(n38298), .dinb(n38179), .dout(n38299));
  jxor g21037(.dina(n38173), .dinb(n355), .dout(n38300));
  jand g21038(.dina(n38300), .dinb(n38299), .dout(n38301));
  jor  g21039(.dina(n38301), .dinb(n38174), .dout(n38302));
  jxor g21040(.dina(n38168), .dinb(n356), .dout(n38303));
  jand g21041(.dina(n38303), .dinb(n38302), .dout(n38304));
  jor  g21042(.dina(n38304), .dinb(n38169), .dout(n38305));
  jxor g21043(.dina(n38163), .dinb(n266), .dout(n38306));
  jand g21044(.dina(n38306), .dinb(n38305), .dout(n38307));
  jor  g21045(.dina(n38307), .dinb(n38164), .dout(n38308));
  jxor g21046(.dina(n38158), .dinb(n267), .dout(n38309));
  jand g21047(.dina(n38309), .dinb(n38308), .dout(n38310));
  jor  g21048(.dina(n38310), .dinb(n38159), .dout(n38311));
  jxor g21049(.dina(n38153), .dinb(n347), .dout(n38312));
  jand g21050(.dina(n38312), .dinb(n38311), .dout(n38313));
  jor  g21051(.dina(n38313), .dinb(n38154), .dout(n38314));
  jxor g21052(.dina(n38148), .dinb(n348), .dout(n38315));
  jand g21053(.dina(n38315), .dinb(n38314), .dout(n38316));
  jor  g21054(.dina(n38316), .dinb(n38149), .dout(n38317));
  jxor g21055(.dina(n38143), .dinb(n349), .dout(n38318));
  jand g21056(.dina(n38318), .dinb(n38317), .dout(n38319));
  jor  g21057(.dina(n38319), .dinb(n38144), .dout(n38320));
  jxor g21058(.dina(n38138), .dinb(n268), .dout(n38321));
  jand g21059(.dina(n38321), .dinb(n38320), .dout(n38322));
  jor  g21060(.dina(n38322), .dinb(n38139), .dout(n38323));
  jxor g21061(.dina(n38133), .dinb(n274), .dout(n38324));
  jand g21062(.dina(n38324), .dinb(n38323), .dout(n38325));
  jor  g21063(.dina(n38325), .dinb(n38134), .dout(n38326));
  jxor g21064(.dina(n38128), .dinb(n269), .dout(n38327));
  jand g21065(.dina(n38327), .dinb(n38326), .dout(n38328));
  jor  g21066(.dina(n38328), .dinb(n38129), .dout(n38329));
  jxor g21067(.dina(n38123), .dinb(n270), .dout(n38330));
  jand g21068(.dina(n38330), .dinb(n38329), .dout(n38331));
  jor  g21069(.dina(n38331), .dinb(n38124), .dout(n38332));
  jxor g21070(.dina(n38118), .dinb(n271), .dout(n38333));
  jand g21071(.dina(n38333), .dinb(n38332), .dout(n38334));
  jor  g21072(.dina(n38334), .dinb(n38119), .dout(n38335));
  jxor g21073(.dina(n38113), .dinb(n338), .dout(n38336));
  jand g21074(.dina(n38336), .dinb(n38335), .dout(n38337));
  jor  g21075(.dina(n38337), .dinb(n38114), .dout(n38338));
  jxor g21076(.dina(n38108), .dinb(n339), .dout(n38339));
  jand g21077(.dina(n38339), .dinb(n38338), .dout(n38340));
  jor  g21078(.dina(n38340), .dinb(n38109), .dout(n38341));
  jxor g21079(.dina(n38103), .dinb(n340), .dout(n38342));
  jand g21080(.dina(n38342), .dinb(n38341), .dout(n38343));
  jor  g21081(.dina(n38343), .dinb(n38104), .dout(n38344));
  jxor g21082(.dina(n38098), .dinb(n275), .dout(n38345));
  jand g21083(.dina(n38345), .dinb(n38344), .dout(n38346));
  jor  g21084(.dina(n38346), .dinb(n38099), .dout(n38347));
  jxor g21085(.dina(n38093), .dinb(n331), .dout(n38348));
  jand g21086(.dina(n38348), .dinb(n38347), .dout(n38349));
  jor  g21087(.dina(n38349), .dinb(n38094), .dout(n38350));
  jxor g21088(.dina(n38088), .dinb(n332), .dout(n38351));
  jand g21089(.dina(n38351), .dinb(n38350), .dout(n38352));
  jor  g21090(.dina(n38352), .dinb(n38089), .dout(n38353));
  jxor g21091(.dina(n38083), .dinb(n333), .dout(n38354));
  jand g21092(.dina(n38354), .dinb(n38353), .dout(n38355));
  jor  g21093(.dina(n38355), .dinb(n38084), .dout(n38356));
  jxor g21094(.dina(n38078), .dinb(n276), .dout(n38357));
  jand g21095(.dina(n38357), .dinb(n38356), .dout(n38358));
  jor  g21096(.dina(n38358), .dinb(n38079), .dout(n38359));
  jxor g21097(.dina(n38073), .dinb(n324), .dout(n38360));
  jand g21098(.dina(n38360), .dinb(n38359), .dout(n38361));
  jor  g21099(.dina(n38361), .dinb(n38074), .dout(n38362));
  jxor g21100(.dina(n38068), .dinb(n325), .dout(n38363));
  jand g21101(.dina(n38363), .dinb(n38362), .dout(n38364));
  jor  g21102(.dina(n38364), .dinb(n38069), .dout(n38365));
  jxor g21103(.dina(n38063), .dinb(n326), .dout(n38366));
  jand g21104(.dina(n38366), .dinb(n38365), .dout(n38367));
  jor  g21105(.dina(n38367), .dinb(n38064), .dout(n38368));
  jxor g21106(.dina(n38058), .dinb(n277), .dout(n38369));
  jand g21107(.dina(n38369), .dinb(n38368), .dout(n38370));
  jor  g21108(.dina(n38370), .dinb(n38059), .dout(n38371));
  jxor g21109(.dina(n38053), .dinb(n278), .dout(n38372));
  jand g21110(.dina(n38372), .dinb(n38371), .dout(n38373));
  jor  g21111(.dina(n38373), .dinb(n38054), .dout(n38374));
  jxor g21112(.dina(n38048), .dinb(n279), .dout(n38375));
  jand g21113(.dina(n38375), .dinb(n38374), .dout(n38376));
  jor  g21114(.dina(n38376), .dinb(n38049), .dout(n38377));
  jxor g21115(.dina(n38043), .dinb(n280), .dout(n38378));
  jand g21116(.dina(n38378), .dinb(n38377), .dout(n38379));
  jor  g21117(.dina(n38379), .dinb(n38044), .dout(n38380));
  jxor g21118(.dina(n38038), .dinb(n283), .dout(n38381));
  jand g21119(.dina(n38381), .dinb(n38380), .dout(n38382));
  jor  g21120(.dina(n38382), .dinb(n38039), .dout(n38383));
  jxor g21121(.dina(n38033), .dinb(n315), .dout(n38384));
  jand g21122(.dina(n38384), .dinb(n38383), .dout(n38385));
  jor  g21123(.dina(n38385), .dinb(n38034), .dout(n38386));
  jxor g21124(.dina(n38028), .dinb(n316), .dout(n38387));
  jand g21125(.dina(n38387), .dinb(n38386), .dout(n38388));
  jor  g21126(.dina(n38388), .dinb(n38029), .dout(n38389));
  jxor g21127(.dina(n38023), .dinb(n317), .dout(n38390));
  jand g21128(.dina(n38390), .dinb(n38389), .dout(n38391));
  jor  g21129(.dina(n38391), .dinb(n38024), .dout(n38392));
  jxor g21130(.dina(n38018), .dinb(n284), .dout(n38393));
  jand g21131(.dina(n38393), .dinb(n38392), .dout(n38394));
  jor  g21132(.dina(n38394), .dinb(n38019), .dout(n38395));
  jxor g21133(.dina(n38013), .dinb(n285), .dout(n38396));
  jand g21134(.dina(n38396), .dinb(n38395), .dout(n38397));
  jor  g21135(.dina(n38397), .dinb(n38014), .dout(n38398));
  jxor g21136(.dina(n38008), .dinb(n286), .dout(n38399));
  jand g21137(.dina(n38399), .dinb(n38398), .dout(n38400));
  jor  g21138(.dina(n38400), .dinb(n38009), .dout(n38401));
  jxor g21139(.dina(n38003), .dinb(n287), .dout(n38402));
  jand g21140(.dina(n38402), .dinb(n38401), .dout(n38403));
  jor  g21141(.dina(n38403), .dinb(n38004), .dout(n38404));
  jxor g21142(.dina(n37998), .dinb(n288), .dout(n38405));
  jand g21143(.dina(n38405), .dinb(n38404), .dout(n38406));
  jor  g21144(.dina(n38406), .dinb(n37999), .dout(n38407));
  jxor g21145(.dina(n37993), .dinb(n289), .dout(n38408));
  jand g21146(.dina(n38408), .dinb(n38407), .dout(n38409));
  jor  g21147(.dina(n38409), .dinb(n37994), .dout(n38410));
  jxor g21148(.dina(n37988), .dinb(n290), .dout(n38411));
  jand g21149(.dina(n38411), .dinb(n38410), .dout(n38412));
  jor  g21150(.dina(n38412), .dinb(n37989), .dout(n38413));
  jxor g21151(.dina(n37983), .dinb(n291), .dout(n38414));
  jand g21152(.dina(n38414), .dinb(n38413), .dout(n38415));
  jor  g21153(.dina(n38415), .dinb(n37984), .dout(n38416));
  jxor g21154(.dina(n37978), .dinb(n292), .dout(n38417));
  jand g21155(.dina(n38417), .dinb(n38416), .dout(n38418));
  jor  g21156(.dina(n38418), .dinb(n37979), .dout(n38419));
  jxor g21157(.dina(n37973), .dinb(n293), .dout(n38420));
  jand g21158(.dina(n38420), .dinb(n38419), .dout(n38421));
  jor  g21159(.dina(n38421), .dinb(n37974), .dout(n38422));
  jxor g21160(.dina(n37968), .dinb(n294), .dout(n38423));
  jand g21161(.dina(n38423), .dinb(n38422), .dout(n38424));
  jor  g21162(.dina(n38424), .dinb(n37969), .dout(n38425));
  jxor g21163(.dina(n37963), .dinb(n295), .dout(n38426));
  jand g21164(.dina(n38426), .dinb(n38425), .dout(n38427));
  jor  g21165(.dina(n38427), .dinb(n37964), .dout(n38428));
  jxor g21166(.dina(n37958), .dinb(n296), .dout(n38429));
  jand g21167(.dina(n38429), .dinb(n38428), .dout(n38430));
  jor  g21168(.dina(n38430), .dinb(n37959), .dout(n38431));
  jxor g21169(.dina(n37953), .dinb(n297), .dout(n38432));
  jand g21170(.dina(n38432), .dinb(n38431), .dout(n38433));
  jor  g21171(.dina(n38433), .dinb(n37954), .dout(n38434));
  jxor g21172(.dina(n37948), .dinb(n257), .dout(n38435));
  jand g21173(.dina(n38435), .dinb(n38434), .dout(n38436));
  jor  g21174(.dina(n38436), .dinb(n37949), .dout(n38437));
  jor  g21175(.dina(n38437), .dinb(n37936), .dout(n38438));
  jnot g21176(.din(n37935), .dout(n38439));
  jand g21177(.dina(n38439), .dinb(b62 ), .dout(n38440));
  jor  g21178(.dina(n38440), .dinb(b63 ), .dout(n38441));
  jnot g21179(.din(n38441), .dout(n38442));
  jand g21180(.dina(n38442), .dinb(n38438), .dout(n38443));
  jnot g21181(.din(n38443), .dout(n38444));
  jand g21182(.dina(n38437), .dinb(n299), .dout(n38445));
  jor  g21183(.dina(n38445), .dinb(n38444), .dout(n38446));
  jand g21184(.dina(n38446), .dinb(n37935), .dout(n38447));
  jand g21185(.dina(n38447), .dinb(n256), .dout(n38448));
  jand g21186(.dina(n38439), .dinb(b63 ), .dout(n38449));
  jnot g21187(.din(n38449), .dout(n38450));
  jor  g21188(.dina(n38443), .dinb(n37948), .dout(n38451));
  jxor g21189(.dina(n38435), .dinb(n38434), .dout(n38452));
  jor  g21190(.dina(n38452), .dinb(n38444), .dout(n38453));
  jand g21191(.dina(n38453), .dinb(n38451), .dout(n38454));
  jand g21192(.dina(n38454), .dinb(n298), .dout(n38455));
  jor  g21193(.dina(n38443), .dinb(n37953), .dout(n38456));
  jxor g21194(.dina(n38432), .dinb(n38431), .dout(n38457));
  jor  g21195(.dina(n38457), .dinb(n38444), .dout(n38458));
  jand g21196(.dina(n38458), .dinb(n38456), .dout(n38459));
  jand g21197(.dina(n38459), .dinb(n257), .dout(n38460));
  jor  g21198(.dina(n38443), .dinb(n37958), .dout(n38461));
  jxor g21199(.dina(n38429), .dinb(n38428), .dout(n38462));
  jor  g21200(.dina(n38462), .dinb(n38444), .dout(n38463));
  jand g21201(.dina(n38463), .dinb(n38461), .dout(n38464));
  jand g21202(.dina(n38464), .dinb(n297), .dout(n38465));
  jor  g21203(.dina(n38443), .dinb(n37963), .dout(n38466));
  jxor g21204(.dina(n38426), .dinb(n38425), .dout(n38467));
  jor  g21205(.dina(n38467), .dinb(n38444), .dout(n38468));
  jand g21206(.dina(n38468), .dinb(n38466), .dout(n38469));
  jand g21207(.dina(n38469), .dinb(n296), .dout(n38470));
  jor  g21208(.dina(n38443), .dinb(n37968), .dout(n38471));
  jxor g21209(.dina(n38423), .dinb(n38422), .dout(n38472));
  jor  g21210(.dina(n38472), .dinb(n38444), .dout(n38473));
  jand g21211(.dina(n38473), .dinb(n38471), .dout(n38474));
  jand g21212(.dina(n38474), .dinb(n295), .dout(n38475));
  jor  g21213(.dina(n38443), .dinb(n37973), .dout(n38476));
  jxor g21214(.dina(n38420), .dinb(n38419), .dout(n38477));
  jor  g21215(.dina(n38477), .dinb(n38444), .dout(n38478));
  jand g21216(.dina(n38478), .dinb(n38476), .dout(n38479));
  jand g21217(.dina(n38479), .dinb(n294), .dout(n38480));
  jor  g21218(.dina(n38443), .dinb(n37978), .dout(n38481));
  jxor g21219(.dina(n38417), .dinb(n38416), .dout(n38482));
  jor  g21220(.dina(n38482), .dinb(n38444), .dout(n38483));
  jand g21221(.dina(n38483), .dinb(n38481), .dout(n38484));
  jand g21222(.dina(n38484), .dinb(n293), .dout(n38485));
  jor  g21223(.dina(n38443), .dinb(n37983), .dout(n38486));
  jxor g21224(.dina(n38414), .dinb(n38413), .dout(n38487));
  jor  g21225(.dina(n38487), .dinb(n38444), .dout(n38488));
  jand g21226(.dina(n38488), .dinb(n38486), .dout(n38489));
  jand g21227(.dina(n38489), .dinb(n292), .dout(n38490));
  jor  g21228(.dina(n38443), .dinb(n37988), .dout(n38491));
  jxor g21229(.dina(n38411), .dinb(n38410), .dout(n38492));
  jor  g21230(.dina(n38492), .dinb(n38444), .dout(n38493));
  jand g21231(.dina(n38493), .dinb(n38491), .dout(n38494));
  jand g21232(.dina(n38494), .dinb(n291), .dout(n38495));
  jor  g21233(.dina(n38443), .dinb(n37993), .dout(n38496));
  jxor g21234(.dina(n38408), .dinb(n38407), .dout(n38497));
  jor  g21235(.dina(n38497), .dinb(n38444), .dout(n38498));
  jand g21236(.dina(n38498), .dinb(n38496), .dout(n38499));
  jand g21237(.dina(n38499), .dinb(n290), .dout(n38500));
  jor  g21238(.dina(n38443), .dinb(n37998), .dout(n38501));
  jxor g21239(.dina(n38405), .dinb(n38404), .dout(n38502));
  jor  g21240(.dina(n38502), .dinb(n38444), .dout(n38503));
  jand g21241(.dina(n38503), .dinb(n38501), .dout(n38504));
  jand g21242(.dina(n38504), .dinb(n289), .dout(n38505));
  jor  g21243(.dina(n38443), .dinb(n38003), .dout(n38506));
  jxor g21244(.dina(n38402), .dinb(n38401), .dout(n38507));
  jor  g21245(.dina(n38507), .dinb(n38444), .dout(n38508));
  jand g21246(.dina(n38508), .dinb(n38506), .dout(n38509));
  jand g21247(.dina(n38509), .dinb(n288), .dout(n38510));
  jor  g21248(.dina(n38443), .dinb(n38008), .dout(n38511));
  jxor g21249(.dina(n38399), .dinb(n38398), .dout(n38512));
  jor  g21250(.dina(n38512), .dinb(n38444), .dout(n38513));
  jand g21251(.dina(n38513), .dinb(n38511), .dout(n38514));
  jand g21252(.dina(n38514), .dinb(n287), .dout(n38515));
  jor  g21253(.dina(n38443), .dinb(n38013), .dout(n38516));
  jxor g21254(.dina(n38396), .dinb(n38395), .dout(n38517));
  jor  g21255(.dina(n38517), .dinb(n38444), .dout(n38518));
  jand g21256(.dina(n38518), .dinb(n38516), .dout(n38519));
  jand g21257(.dina(n38519), .dinb(n286), .dout(n38520));
  jor  g21258(.dina(n38443), .dinb(n38018), .dout(n38521));
  jxor g21259(.dina(n38393), .dinb(n38392), .dout(n38522));
  jor  g21260(.dina(n38522), .dinb(n38444), .dout(n38523));
  jand g21261(.dina(n38523), .dinb(n38521), .dout(n38524));
  jand g21262(.dina(n38524), .dinb(n285), .dout(n38525));
  jor  g21263(.dina(n38443), .dinb(n38023), .dout(n38526));
  jxor g21264(.dina(n38390), .dinb(n38389), .dout(n38527));
  jor  g21265(.dina(n38527), .dinb(n38444), .dout(n38528));
  jand g21266(.dina(n38528), .dinb(n38526), .dout(n38529));
  jand g21267(.dina(n38529), .dinb(n284), .dout(n38530));
  jor  g21268(.dina(n38443), .dinb(n38028), .dout(n38531));
  jxor g21269(.dina(n38387), .dinb(n38386), .dout(n38532));
  jor  g21270(.dina(n38532), .dinb(n38444), .dout(n38533));
  jand g21271(.dina(n38533), .dinb(n38531), .dout(n38534));
  jand g21272(.dina(n38534), .dinb(n317), .dout(n38535));
  jor  g21273(.dina(n38443), .dinb(n38033), .dout(n38536));
  jxor g21274(.dina(n38384), .dinb(n38383), .dout(n38537));
  jor  g21275(.dina(n38537), .dinb(n38444), .dout(n38538));
  jand g21276(.dina(n38538), .dinb(n38536), .dout(n38539));
  jand g21277(.dina(n38539), .dinb(n316), .dout(n38540));
  jor  g21278(.dina(n38443), .dinb(n38038), .dout(n38541));
  jxor g21279(.dina(n38381), .dinb(n38380), .dout(n38542));
  jor  g21280(.dina(n38542), .dinb(n38444), .dout(n38543));
  jand g21281(.dina(n38543), .dinb(n38541), .dout(n38544));
  jand g21282(.dina(n38544), .dinb(n315), .dout(n38545));
  jor  g21283(.dina(n38443), .dinb(n38043), .dout(n38546));
  jxor g21284(.dina(n38378), .dinb(n38377), .dout(n38547));
  jor  g21285(.dina(n38547), .dinb(n38444), .dout(n38548));
  jand g21286(.dina(n38548), .dinb(n38546), .dout(n38549));
  jand g21287(.dina(n38549), .dinb(n283), .dout(n38550));
  jor  g21288(.dina(n38443), .dinb(n38048), .dout(n38551));
  jxor g21289(.dina(n38375), .dinb(n38374), .dout(n38552));
  jor  g21290(.dina(n38552), .dinb(n38444), .dout(n38553));
  jand g21291(.dina(n38553), .dinb(n38551), .dout(n38554));
  jand g21292(.dina(n38554), .dinb(n280), .dout(n38555));
  jor  g21293(.dina(n38443), .dinb(n38053), .dout(n38556));
  jxor g21294(.dina(n38372), .dinb(n38371), .dout(n38557));
  jor  g21295(.dina(n38557), .dinb(n38444), .dout(n38558));
  jand g21296(.dina(n38558), .dinb(n38556), .dout(n38559));
  jand g21297(.dina(n38559), .dinb(n279), .dout(n38560));
  jor  g21298(.dina(n38443), .dinb(n38058), .dout(n38561));
  jxor g21299(.dina(n38369), .dinb(n38368), .dout(n38562));
  jor  g21300(.dina(n38562), .dinb(n38444), .dout(n38563));
  jand g21301(.dina(n38563), .dinb(n38561), .dout(n38564));
  jand g21302(.dina(n38564), .dinb(n278), .dout(n38565));
  jor  g21303(.dina(n38443), .dinb(n38063), .dout(n38566));
  jxor g21304(.dina(n38366), .dinb(n38365), .dout(n38567));
  jor  g21305(.dina(n38567), .dinb(n38444), .dout(n38568));
  jand g21306(.dina(n38568), .dinb(n38566), .dout(n38569));
  jand g21307(.dina(n38569), .dinb(n277), .dout(n38570));
  jor  g21308(.dina(n38443), .dinb(n38068), .dout(n38571));
  jxor g21309(.dina(n38363), .dinb(n38362), .dout(n38572));
  jor  g21310(.dina(n38572), .dinb(n38444), .dout(n38573));
  jand g21311(.dina(n38573), .dinb(n38571), .dout(n38574));
  jand g21312(.dina(n38574), .dinb(n326), .dout(n38575));
  jor  g21313(.dina(n38443), .dinb(n38073), .dout(n38576));
  jxor g21314(.dina(n38360), .dinb(n38359), .dout(n38577));
  jor  g21315(.dina(n38577), .dinb(n38444), .dout(n38578));
  jand g21316(.dina(n38578), .dinb(n38576), .dout(n38579));
  jand g21317(.dina(n38579), .dinb(n325), .dout(n38580));
  jor  g21318(.dina(n38443), .dinb(n38078), .dout(n38581));
  jxor g21319(.dina(n38357), .dinb(n38356), .dout(n38582));
  jor  g21320(.dina(n38582), .dinb(n38444), .dout(n38583));
  jand g21321(.dina(n38583), .dinb(n38581), .dout(n38584));
  jand g21322(.dina(n38584), .dinb(n324), .dout(n38585));
  jor  g21323(.dina(n38443), .dinb(n38083), .dout(n38586));
  jxor g21324(.dina(n38354), .dinb(n38353), .dout(n38587));
  jor  g21325(.dina(n38587), .dinb(n38444), .dout(n38588));
  jand g21326(.dina(n38588), .dinb(n38586), .dout(n38589));
  jand g21327(.dina(n38589), .dinb(n276), .dout(n38590));
  jor  g21328(.dina(n38443), .dinb(n38088), .dout(n38591));
  jxor g21329(.dina(n38351), .dinb(n38350), .dout(n38592));
  jor  g21330(.dina(n38592), .dinb(n38444), .dout(n38593));
  jand g21331(.dina(n38593), .dinb(n38591), .dout(n38594));
  jand g21332(.dina(n38594), .dinb(n333), .dout(n38595));
  jor  g21333(.dina(n38443), .dinb(n38093), .dout(n38596));
  jxor g21334(.dina(n38348), .dinb(n38347), .dout(n38597));
  jor  g21335(.dina(n38597), .dinb(n38444), .dout(n38598));
  jand g21336(.dina(n38598), .dinb(n38596), .dout(n38599));
  jand g21337(.dina(n38599), .dinb(n332), .dout(n38600));
  jor  g21338(.dina(n38443), .dinb(n38098), .dout(n38601));
  jxor g21339(.dina(n38345), .dinb(n38344), .dout(n38602));
  jor  g21340(.dina(n38602), .dinb(n38444), .dout(n38603));
  jand g21341(.dina(n38603), .dinb(n38601), .dout(n38604));
  jand g21342(.dina(n38604), .dinb(n331), .dout(n38605));
  jor  g21343(.dina(n38443), .dinb(n38103), .dout(n38606));
  jxor g21344(.dina(n38342), .dinb(n38341), .dout(n38607));
  jor  g21345(.dina(n38607), .dinb(n38444), .dout(n38608));
  jand g21346(.dina(n38608), .dinb(n38606), .dout(n38609));
  jand g21347(.dina(n38609), .dinb(n275), .dout(n38610));
  jor  g21348(.dina(n38443), .dinb(n38108), .dout(n38611));
  jxor g21349(.dina(n38339), .dinb(n38338), .dout(n38612));
  jor  g21350(.dina(n38612), .dinb(n38444), .dout(n38613));
  jand g21351(.dina(n38613), .dinb(n38611), .dout(n38614));
  jand g21352(.dina(n38614), .dinb(n340), .dout(n38615));
  jor  g21353(.dina(n38443), .dinb(n38113), .dout(n38616));
  jxor g21354(.dina(n38336), .dinb(n38335), .dout(n38617));
  jor  g21355(.dina(n38617), .dinb(n38444), .dout(n38618));
  jand g21356(.dina(n38618), .dinb(n38616), .dout(n38619));
  jand g21357(.dina(n38619), .dinb(n339), .dout(n38620));
  jor  g21358(.dina(n38443), .dinb(n38118), .dout(n38621));
  jxor g21359(.dina(n38333), .dinb(n38332), .dout(n38622));
  jor  g21360(.dina(n38622), .dinb(n38444), .dout(n38623));
  jand g21361(.dina(n38623), .dinb(n38621), .dout(n38624));
  jand g21362(.dina(n38624), .dinb(n338), .dout(n38625));
  jor  g21363(.dina(n38443), .dinb(n38123), .dout(n38626));
  jxor g21364(.dina(n38330), .dinb(n38329), .dout(n38627));
  jor  g21365(.dina(n38627), .dinb(n38444), .dout(n38628));
  jand g21366(.dina(n38628), .dinb(n38626), .dout(n38629));
  jand g21367(.dina(n38629), .dinb(n271), .dout(n38630));
  jor  g21368(.dina(n38443), .dinb(n38128), .dout(n38631));
  jxor g21369(.dina(n38327), .dinb(n38326), .dout(n38632));
  jor  g21370(.dina(n38632), .dinb(n38444), .dout(n38633));
  jand g21371(.dina(n38633), .dinb(n38631), .dout(n38634));
  jand g21372(.dina(n38634), .dinb(n270), .dout(n38635));
  jor  g21373(.dina(n38443), .dinb(n38133), .dout(n38636));
  jxor g21374(.dina(n38324), .dinb(n38323), .dout(n38637));
  jor  g21375(.dina(n38637), .dinb(n38444), .dout(n38638));
  jand g21376(.dina(n38638), .dinb(n38636), .dout(n38639));
  jand g21377(.dina(n38639), .dinb(n269), .dout(n38640));
  jor  g21378(.dina(n38443), .dinb(n38138), .dout(n38641));
  jxor g21379(.dina(n38321), .dinb(n38320), .dout(n38642));
  jor  g21380(.dina(n38642), .dinb(n38444), .dout(n38643));
  jand g21381(.dina(n38643), .dinb(n38641), .dout(n38644));
  jand g21382(.dina(n38644), .dinb(n274), .dout(n38645));
  jor  g21383(.dina(n38443), .dinb(n38143), .dout(n38646));
  jxor g21384(.dina(n38318), .dinb(n38317), .dout(n38647));
  jor  g21385(.dina(n38647), .dinb(n38444), .dout(n38648));
  jand g21386(.dina(n38648), .dinb(n38646), .dout(n38649));
  jand g21387(.dina(n38649), .dinb(n268), .dout(n38650));
  jor  g21388(.dina(n38443), .dinb(n38148), .dout(n38651));
  jxor g21389(.dina(n38315), .dinb(n38314), .dout(n38652));
  jor  g21390(.dina(n38652), .dinb(n38444), .dout(n38653));
  jand g21391(.dina(n38653), .dinb(n38651), .dout(n38654));
  jand g21392(.dina(n38654), .dinb(n349), .dout(n38655));
  jor  g21393(.dina(n38443), .dinb(n38153), .dout(n38656));
  jxor g21394(.dina(n38312), .dinb(n38311), .dout(n38657));
  jor  g21395(.dina(n38657), .dinb(n38444), .dout(n38658));
  jand g21396(.dina(n38658), .dinb(n38656), .dout(n38659));
  jand g21397(.dina(n38659), .dinb(n348), .dout(n38660));
  jor  g21398(.dina(n38443), .dinb(n38158), .dout(n38661));
  jxor g21399(.dina(n38309), .dinb(n38308), .dout(n38662));
  jor  g21400(.dina(n38662), .dinb(n38444), .dout(n38663));
  jand g21401(.dina(n38663), .dinb(n38661), .dout(n38664));
  jand g21402(.dina(n38664), .dinb(n347), .dout(n38665));
  jor  g21403(.dina(n38443), .dinb(n38163), .dout(n38666));
  jxor g21404(.dina(n38306), .dinb(n38305), .dout(n38667));
  jor  g21405(.dina(n38667), .dinb(n38444), .dout(n38668));
  jand g21406(.dina(n38668), .dinb(n38666), .dout(n38669));
  jand g21407(.dina(n38669), .dinb(n267), .dout(n38670));
  jor  g21408(.dina(n38443), .dinb(n38168), .dout(n38671));
  jxor g21409(.dina(n38303), .dinb(n38302), .dout(n38672));
  jor  g21410(.dina(n38672), .dinb(n38444), .dout(n38673));
  jand g21411(.dina(n38673), .dinb(n38671), .dout(n38674));
  jand g21412(.dina(n38674), .dinb(n266), .dout(n38675));
  jor  g21413(.dina(n38443), .dinb(n38173), .dout(n38676));
  jxor g21414(.dina(n38300), .dinb(n38299), .dout(n38677));
  jor  g21415(.dina(n38677), .dinb(n38444), .dout(n38678));
  jand g21416(.dina(n38678), .dinb(n38676), .dout(n38679));
  jand g21417(.dina(n38679), .dinb(n356), .dout(n38680));
  jor  g21418(.dina(n38443), .dinb(n38178), .dout(n38681));
  jxor g21419(.dina(n38297), .dinb(n38296), .dout(n38682));
  jor  g21420(.dina(n38682), .dinb(n38444), .dout(n38683));
  jand g21421(.dina(n38683), .dinb(n38681), .dout(n38684));
  jand g21422(.dina(n38684), .dinb(n355), .dout(n38685));
  jor  g21423(.dina(n38443), .dinb(n38183), .dout(n38686));
  jxor g21424(.dina(n38294), .dinb(n38293), .dout(n38687));
  jor  g21425(.dina(n38687), .dinb(n38444), .dout(n38688));
  jand g21426(.dina(n38688), .dinb(n38686), .dout(n38689));
  jand g21427(.dina(n38689), .dinb(n364), .dout(n38690));
  jor  g21428(.dina(n38443), .dinb(n38188), .dout(n38691));
  jxor g21429(.dina(n38291), .dinb(n38290), .dout(n38692));
  jor  g21430(.dina(n38692), .dinb(n38444), .dout(n38693));
  jand g21431(.dina(n38693), .dinb(n38691), .dout(n38694));
  jand g21432(.dina(n38694), .dinb(n361), .dout(n38695));
  jor  g21433(.dina(n38443), .dinb(n38193), .dout(n38696));
  jxor g21434(.dina(n38288), .dinb(n38287), .dout(n38697));
  jor  g21435(.dina(n38697), .dinb(n38444), .dout(n38698));
  jand g21436(.dina(n38698), .dinb(n38696), .dout(n38699));
  jand g21437(.dina(n38699), .dinb(n360), .dout(n38700));
  jor  g21438(.dina(n38443), .dinb(n38198), .dout(n38701));
  jxor g21439(.dina(n38285), .dinb(n38284), .dout(n38702));
  jor  g21440(.dina(n38702), .dinb(n38444), .dout(n38703));
  jand g21441(.dina(n38703), .dinb(n38701), .dout(n38704));
  jand g21442(.dina(n38704), .dinb(n363), .dout(n38705));
  jor  g21443(.dina(n38443), .dinb(n38203), .dout(n38706));
  jxor g21444(.dina(n38282), .dinb(n38281), .dout(n38707));
  jor  g21445(.dina(n38707), .dinb(n38444), .dout(n38708));
  jand g21446(.dina(n38708), .dinb(n38706), .dout(n38709));
  jand g21447(.dina(n38709), .dinb(n359), .dout(n38710));
  jor  g21448(.dina(n38443), .dinb(n38208), .dout(n38711));
  jxor g21449(.dina(n38279), .dinb(n38278), .dout(n38712));
  jor  g21450(.dina(n38712), .dinb(n38444), .dout(n38713));
  jand g21451(.dina(n38713), .dinb(n38711), .dout(n38714));
  jand g21452(.dina(n38714), .dinb(n369), .dout(n38715));
  jor  g21453(.dina(n38443), .dinb(n38213), .dout(n38716));
  jxor g21454(.dina(n38276), .dinb(n38275), .dout(n38717));
  jor  g21455(.dina(n38717), .dinb(n38444), .dout(n38718));
  jand g21456(.dina(n38718), .dinb(n38716), .dout(n38719));
  jand g21457(.dina(n38719), .dinb(n368), .dout(n38720));
  jor  g21458(.dina(n38443), .dinb(n38218), .dout(n38721));
  jxor g21459(.dina(n38273), .dinb(n38272), .dout(n38722));
  jor  g21460(.dina(n38722), .dinb(n38444), .dout(n38723));
  jand g21461(.dina(n38723), .dinb(n38721), .dout(n38724));
  jand g21462(.dina(n38724), .dinb(n367), .dout(n38725));
  jor  g21463(.dina(n38443), .dinb(n38223), .dout(n38726));
  jxor g21464(.dina(n38270), .dinb(n38269), .dout(n38727));
  jor  g21465(.dina(n38727), .dinb(n38444), .dout(n38728));
  jand g21466(.dina(n38728), .dinb(n38726), .dout(n38729));
  jand g21467(.dina(n38729), .dinb(n265), .dout(n38730));
  jor  g21468(.dina(n38443), .dinb(n38228), .dout(n38731));
  jxor g21469(.dina(n38267), .dinb(n38266), .dout(n38732));
  jor  g21470(.dina(n38732), .dinb(n38444), .dout(n38733));
  jand g21471(.dina(n38733), .dinb(n38731), .dout(n38734));
  jand g21472(.dina(n38734), .dinb(n378), .dout(n38735));
  jor  g21473(.dina(n38443), .dinb(n38233), .dout(n38736));
  jxor g21474(.dina(n38264), .dinb(n38263), .dout(n38737));
  jor  g21475(.dina(n38737), .dinb(n38444), .dout(n38738));
  jand g21476(.dina(n38738), .dinb(n38736), .dout(n38739));
  jand g21477(.dina(n38739), .dinb(n377), .dout(n38740));
  jor  g21478(.dina(n38443), .dinb(n38239), .dout(n38741));
  jxor g21479(.dina(n38261), .dinb(n38260), .dout(n38742));
  jor  g21480(.dina(n38742), .dinb(n38444), .dout(n38743));
  jand g21481(.dina(n38743), .dinb(n38741), .dout(n38744));
  jand g21482(.dina(n38744), .dinb(n376), .dout(n38745));
  jor  g21483(.dina(n38443), .dinb(n38244), .dout(n38746));
  jxor g21484(.dina(n38258), .dinb(n38257), .dout(n38747));
  jor  g21485(.dina(n38747), .dinb(n38444), .dout(n38748));
  jand g21486(.dina(n38748), .dinb(n38746), .dout(n38749));
  jand g21487(.dina(n38749), .dinb(n264), .dout(n38750));
  jor  g21488(.dina(n38443), .dinb(n38254), .dout(n38751));
  jxor g21489(.dina(n38255), .dinb(n17079), .dout(n38752));
  jand g21490(.dina(n38752), .dinb(n38443), .dout(n38753));
  jnot g21491(.din(n38753), .dout(n38754));
  jand g21492(.dina(n38754), .dinb(n38751), .dout(n38755));
  jor  g21493(.dina(n38755), .dinb(b2 ), .dout(n38756));
  jnot g21494(.din(n38756), .dout(n38757));
  jand g21495(.dina(n38443), .dinb(b0 ), .dout(n38758));
  jxor g21496(.dina(n38758), .dinb(a1 ), .dout(n38759));
  jand g21497(.dina(n38759), .dinb(n259), .dout(n38760));
  jxor g21498(.dina(n38758), .dinb(n17077), .dout(n38761));
  jxor g21499(.dina(n38761), .dinb(b1 ), .dout(n38762));
  jand g21500(.dina(n38762), .dinb(n17823), .dout(n38763));
  jor  g21501(.dina(n38763), .dinb(n38760), .dout(n38764));
  jxor g21502(.dina(n38755), .dinb(b2 ), .dout(n38765));
  jand g21503(.dina(n38765), .dinb(n38764), .dout(n38766));
  jor  g21504(.dina(n38766), .dinb(n38757), .dout(n38767));
  jxor g21505(.dina(n38749), .dinb(n264), .dout(n38768));
  jand g21506(.dina(n38768), .dinb(n38767), .dout(n38769));
  jor  g21507(.dina(n38769), .dinb(n38750), .dout(n38770));
  jxor g21508(.dina(n38744), .dinb(n376), .dout(n38771));
  jand g21509(.dina(n38771), .dinb(n38770), .dout(n38772));
  jor  g21510(.dina(n38772), .dinb(n38745), .dout(n38773));
  jxor g21511(.dina(n38739), .dinb(n377), .dout(n38774));
  jand g21512(.dina(n38774), .dinb(n38773), .dout(n38775));
  jor  g21513(.dina(n38775), .dinb(n38740), .dout(n38776));
  jxor g21514(.dina(n38734), .dinb(n378), .dout(n38777));
  jand g21515(.dina(n38777), .dinb(n38776), .dout(n38778));
  jor  g21516(.dina(n38778), .dinb(n38735), .dout(n38779));
  jxor g21517(.dina(n38729), .dinb(n265), .dout(n38780));
  jand g21518(.dina(n38780), .dinb(n38779), .dout(n38781));
  jor  g21519(.dina(n38781), .dinb(n38730), .dout(n38782));
  jxor g21520(.dina(n38724), .dinb(n367), .dout(n38783));
  jand g21521(.dina(n38783), .dinb(n38782), .dout(n38784));
  jor  g21522(.dina(n38784), .dinb(n38725), .dout(n38785));
  jxor g21523(.dina(n38719), .dinb(n368), .dout(n38786));
  jand g21524(.dina(n38786), .dinb(n38785), .dout(n38787));
  jor  g21525(.dina(n38787), .dinb(n38720), .dout(n38788));
  jxor g21526(.dina(n38714), .dinb(n369), .dout(n38789));
  jand g21527(.dina(n38789), .dinb(n38788), .dout(n38790));
  jor  g21528(.dina(n38790), .dinb(n38715), .dout(n38791));
  jxor g21529(.dina(n38709), .dinb(n359), .dout(n38792));
  jand g21530(.dina(n38792), .dinb(n38791), .dout(n38793));
  jor  g21531(.dina(n38793), .dinb(n38710), .dout(n38794));
  jxor g21532(.dina(n38704), .dinb(n363), .dout(n38795));
  jand g21533(.dina(n38795), .dinb(n38794), .dout(n38796));
  jor  g21534(.dina(n38796), .dinb(n38705), .dout(n38797));
  jxor g21535(.dina(n38699), .dinb(n360), .dout(n38798));
  jand g21536(.dina(n38798), .dinb(n38797), .dout(n38799));
  jor  g21537(.dina(n38799), .dinb(n38700), .dout(n38800));
  jxor g21538(.dina(n38694), .dinb(n361), .dout(n38801));
  jand g21539(.dina(n38801), .dinb(n38800), .dout(n38802));
  jor  g21540(.dina(n38802), .dinb(n38695), .dout(n38803));
  jxor g21541(.dina(n38689), .dinb(n364), .dout(n38804));
  jand g21542(.dina(n38804), .dinb(n38803), .dout(n38805));
  jor  g21543(.dina(n38805), .dinb(n38690), .dout(n38806));
  jxor g21544(.dina(n38684), .dinb(n355), .dout(n38807));
  jand g21545(.dina(n38807), .dinb(n38806), .dout(n38808));
  jor  g21546(.dina(n38808), .dinb(n38685), .dout(n38809));
  jxor g21547(.dina(n38679), .dinb(n356), .dout(n38810));
  jand g21548(.dina(n38810), .dinb(n38809), .dout(n38811));
  jor  g21549(.dina(n38811), .dinb(n38680), .dout(n38812));
  jxor g21550(.dina(n38674), .dinb(n266), .dout(n38813));
  jand g21551(.dina(n38813), .dinb(n38812), .dout(n38814));
  jor  g21552(.dina(n38814), .dinb(n38675), .dout(n38815));
  jxor g21553(.dina(n38669), .dinb(n267), .dout(n38816));
  jand g21554(.dina(n38816), .dinb(n38815), .dout(n38817));
  jor  g21555(.dina(n38817), .dinb(n38670), .dout(n38818));
  jxor g21556(.dina(n38664), .dinb(n347), .dout(n38819));
  jand g21557(.dina(n38819), .dinb(n38818), .dout(n38820));
  jor  g21558(.dina(n38820), .dinb(n38665), .dout(n38821));
  jxor g21559(.dina(n38659), .dinb(n348), .dout(n38822));
  jand g21560(.dina(n38822), .dinb(n38821), .dout(n38823));
  jor  g21561(.dina(n38823), .dinb(n38660), .dout(n38824));
  jxor g21562(.dina(n38654), .dinb(n349), .dout(n38825));
  jand g21563(.dina(n38825), .dinb(n38824), .dout(n38826));
  jor  g21564(.dina(n38826), .dinb(n38655), .dout(n38827));
  jxor g21565(.dina(n38649), .dinb(n268), .dout(n38828));
  jand g21566(.dina(n38828), .dinb(n38827), .dout(n38829));
  jor  g21567(.dina(n38829), .dinb(n38650), .dout(n38830));
  jxor g21568(.dina(n38644), .dinb(n274), .dout(n38831));
  jand g21569(.dina(n38831), .dinb(n38830), .dout(n38832));
  jor  g21570(.dina(n38832), .dinb(n38645), .dout(n38833));
  jxor g21571(.dina(n38639), .dinb(n269), .dout(n38834));
  jand g21572(.dina(n38834), .dinb(n38833), .dout(n38835));
  jor  g21573(.dina(n38835), .dinb(n38640), .dout(n38836));
  jxor g21574(.dina(n38634), .dinb(n270), .dout(n38837));
  jand g21575(.dina(n38837), .dinb(n38836), .dout(n38838));
  jor  g21576(.dina(n38838), .dinb(n38635), .dout(n38839));
  jxor g21577(.dina(n38629), .dinb(n271), .dout(n38840));
  jand g21578(.dina(n38840), .dinb(n38839), .dout(n38841));
  jor  g21579(.dina(n38841), .dinb(n38630), .dout(n38842));
  jxor g21580(.dina(n38624), .dinb(n338), .dout(n38843));
  jand g21581(.dina(n38843), .dinb(n38842), .dout(n38844));
  jor  g21582(.dina(n38844), .dinb(n38625), .dout(n38845));
  jxor g21583(.dina(n38619), .dinb(n339), .dout(n38846));
  jand g21584(.dina(n38846), .dinb(n38845), .dout(n38847));
  jor  g21585(.dina(n38847), .dinb(n38620), .dout(n38848));
  jxor g21586(.dina(n38614), .dinb(n340), .dout(n38849));
  jand g21587(.dina(n38849), .dinb(n38848), .dout(n38850));
  jor  g21588(.dina(n38850), .dinb(n38615), .dout(n38851));
  jxor g21589(.dina(n38609), .dinb(n275), .dout(n38852));
  jand g21590(.dina(n38852), .dinb(n38851), .dout(n38853));
  jor  g21591(.dina(n38853), .dinb(n38610), .dout(n38854));
  jxor g21592(.dina(n38604), .dinb(n331), .dout(n38855));
  jand g21593(.dina(n38855), .dinb(n38854), .dout(n38856));
  jor  g21594(.dina(n38856), .dinb(n38605), .dout(n38857));
  jxor g21595(.dina(n38599), .dinb(n332), .dout(n38858));
  jand g21596(.dina(n38858), .dinb(n38857), .dout(n38859));
  jor  g21597(.dina(n38859), .dinb(n38600), .dout(n38860));
  jxor g21598(.dina(n38594), .dinb(n333), .dout(n38861));
  jand g21599(.dina(n38861), .dinb(n38860), .dout(n38862));
  jor  g21600(.dina(n38862), .dinb(n38595), .dout(n38863));
  jxor g21601(.dina(n38589), .dinb(n276), .dout(n38864));
  jand g21602(.dina(n38864), .dinb(n38863), .dout(n38865));
  jor  g21603(.dina(n38865), .dinb(n38590), .dout(n38866));
  jxor g21604(.dina(n38584), .dinb(n324), .dout(n38867));
  jand g21605(.dina(n38867), .dinb(n38866), .dout(n38868));
  jor  g21606(.dina(n38868), .dinb(n38585), .dout(n38869));
  jxor g21607(.dina(n38579), .dinb(n325), .dout(n38870));
  jand g21608(.dina(n38870), .dinb(n38869), .dout(n38871));
  jor  g21609(.dina(n38871), .dinb(n38580), .dout(n38872));
  jxor g21610(.dina(n38574), .dinb(n326), .dout(n38873));
  jand g21611(.dina(n38873), .dinb(n38872), .dout(n38874));
  jor  g21612(.dina(n38874), .dinb(n38575), .dout(n38875));
  jxor g21613(.dina(n38569), .dinb(n277), .dout(n38876));
  jand g21614(.dina(n38876), .dinb(n38875), .dout(n38877));
  jor  g21615(.dina(n38877), .dinb(n38570), .dout(n38878));
  jxor g21616(.dina(n38564), .dinb(n278), .dout(n38879));
  jand g21617(.dina(n38879), .dinb(n38878), .dout(n38880));
  jor  g21618(.dina(n38880), .dinb(n38565), .dout(n38881));
  jxor g21619(.dina(n38559), .dinb(n279), .dout(n38882));
  jand g21620(.dina(n38882), .dinb(n38881), .dout(n38883));
  jor  g21621(.dina(n38883), .dinb(n38560), .dout(n38884));
  jxor g21622(.dina(n38554), .dinb(n280), .dout(n38885));
  jand g21623(.dina(n38885), .dinb(n38884), .dout(n38886));
  jor  g21624(.dina(n38886), .dinb(n38555), .dout(n38887));
  jxor g21625(.dina(n38549), .dinb(n283), .dout(n38888));
  jand g21626(.dina(n38888), .dinb(n38887), .dout(n38889));
  jor  g21627(.dina(n38889), .dinb(n38550), .dout(n38890));
  jxor g21628(.dina(n38544), .dinb(n315), .dout(n38891));
  jand g21629(.dina(n38891), .dinb(n38890), .dout(n38892));
  jor  g21630(.dina(n38892), .dinb(n38545), .dout(n38893));
  jxor g21631(.dina(n38539), .dinb(n316), .dout(n38894));
  jand g21632(.dina(n38894), .dinb(n38893), .dout(n38895));
  jor  g21633(.dina(n38895), .dinb(n38540), .dout(n38896));
  jxor g21634(.dina(n38534), .dinb(n317), .dout(n38897));
  jand g21635(.dina(n38897), .dinb(n38896), .dout(n38898));
  jor  g21636(.dina(n38898), .dinb(n38535), .dout(n38899));
  jxor g21637(.dina(n38529), .dinb(n284), .dout(n38900));
  jand g21638(.dina(n38900), .dinb(n38899), .dout(n38901));
  jor  g21639(.dina(n38901), .dinb(n38530), .dout(n38902));
  jxor g21640(.dina(n38524), .dinb(n285), .dout(n38903));
  jand g21641(.dina(n38903), .dinb(n38902), .dout(n38904));
  jor  g21642(.dina(n38904), .dinb(n38525), .dout(n38905));
  jxor g21643(.dina(n38519), .dinb(n286), .dout(n38906));
  jand g21644(.dina(n38906), .dinb(n38905), .dout(n38907));
  jor  g21645(.dina(n38907), .dinb(n38520), .dout(n38908));
  jxor g21646(.dina(n38514), .dinb(n287), .dout(n38909));
  jand g21647(.dina(n38909), .dinb(n38908), .dout(n38910));
  jor  g21648(.dina(n38910), .dinb(n38515), .dout(n38911));
  jxor g21649(.dina(n38509), .dinb(n288), .dout(n38912));
  jand g21650(.dina(n38912), .dinb(n38911), .dout(n38913));
  jor  g21651(.dina(n38913), .dinb(n38510), .dout(n38914));
  jxor g21652(.dina(n38504), .dinb(n289), .dout(n38915));
  jand g21653(.dina(n38915), .dinb(n38914), .dout(n38916));
  jor  g21654(.dina(n38916), .dinb(n38505), .dout(n38917));
  jxor g21655(.dina(n38499), .dinb(n290), .dout(n38918));
  jand g21656(.dina(n38918), .dinb(n38917), .dout(n38919));
  jor  g21657(.dina(n38919), .dinb(n38500), .dout(n38920));
  jxor g21658(.dina(n38494), .dinb(n291), .dout(n38921));
  jand g21659(.dina(n38921), .dinb(n38920), .dout(n38922));
  jor  g21660(.dina(n38922), .dinb(n38495), .dout(n38923));
  jxor g21661(.dina(n38489), .dinb(n292), .dout(n38924));
  jand g21662(.dina(n38924), .dinb(n38923), .dout(n38925));
  jor  g21663(.dina(n38925), .dinb(n38490), .dout(n38926));
  jxor g21664(.dina(n38484), .dinb(n293), .dout(n38927));
  jand g21665(.dina(n38927), .dinb(n38926), .dout(n38928));
  jor  g21666(.dina(n38928), .dinb(n38485), .dout(n38929));
  jxor g21667(.dina(n38479), .dinb(n294), .dout(n38930));
  jand g21668(.dina(n38930), .dinb(n38929), .dout(n38931));
  jor  g21669(.dina(n38931), .dinb(n38480), .dout(n38932));
  jxor g21670(.dina(n38474), .dinb(n295), .dout(n38933));
  jand g21671(.dina(n38933), .dinb(n38932), .dout(n38934));
  jor  g21672(.dina(n38934), .dinb(n38475), .dout(n38935));
  jxor g21673(.dina(n38469), .dinb(n296), .dout(n38936));
  jand g21674(.dina(n38936), .dinb(n38935), .dout(n38937));
  jor  g21675(.dina(n38937), .dinb(n38470), .dout(n38938));
  jxor g21676(.dina(n38464), .dinb(n297), .dout(n38939));
  jand g21677(.dina(n38939), .dinb(n38938), .dout(n38940));
  jor  g21678(.dina(n38940), .dinb(n38465), .dout(n38941));
  jxor g21679(.dina(n38459), .dinb(n257), .dout(n38942));
  jand g21680(.dina(n38942), .dinb(n38941), .dout(n38943));
  jor  g21681(.dina(n38943), .dinb(n38460), .dout(n38944));
  jxor g21682(.dina(n38454), .dinb(n298), .dout(n38945));
  jand g21683(.dina(n38945), .dinb(n38944), .dout(n38946));
  jor  g21684(.dina(n38946), .dinb(n38455), .dout(n38947));
  jand g21685(.dina(n38947), .dinb(n38450), .dout(n38948));
  jor  g21686(.dina(n38948), .dinb(n38448), .dout(n38949));
  jand g21687(.dina(n38949), .dinb(b0 ), .dout(n38950));
  jxor g21688(.dina(n38950), .dinb(a0 ), .dout(remainder0 ));
  jnot g21689(.din(n38448), .dout(n38952));
  jnot g21690(.din(n38455), .dout(n38953));
  jnot g21691(.din(n38460), .dout(n38954));
  jnot g21692(.din(n38465), .dout(n38955));
  jnot g21693(.din(n38470), .dout(n38956));
  jnot g21694(.din(n38475), .dout(n38957));
  jnot g21695(.din(n38480), .dout(n38958));
  jnot g21696(.din(n38485), .dout(n38959));
  jnot g21697(.din(n38490), .dout(n38960));
  jnot g21698(.din(n38495), .dout(n38961));
  jnot g21699(.din(n38500), .dout(n38962));
  jnot g21700(.din(n38505), .dout(n38963));
  jnot g21701(.din(n38510), .dout(n38964));
  jnot g21702(.din(n38515), .dout(n38965));
  jnot g21703(.din(n38520), .dout(n38966));
  jnot g21704(.din(n38525), .dout(n38967));
  jnot g21705(.din(n38530), .dout(n38968));
  jnot g21706(.din(n38535), .dout(n38969));
  jnot g21707(.din(n38540), .dout(n38970));
  jnot g21708(.din(n38545), .dout(n38971));
  jnot g21709(.din(n38550), .dout(n38972));
  jnot g21710(.din(n38555), .dout(n38973));
  jnot g21711(.din(n38560), .dout(n38974));
  jnot g21712(.din(n38565), .dout(n38975));
  jnot g21713(.din(n38570), .dout(n38976));
  jnot g21714(.din(n38575), .dout(n38977));
  jnot g21715(.din(n38580), .dout(n38978));
  jnot g21716(.din(n38585), .dout(n38979));
  jnot g21717(.din(n38590), .dout(n38980));
  jnot g21718(.din(n38595), .dout(n38981));
  jnot g21719(.din(n38600), .dout(n38982));
  jnot g21720(.din(n38605), .dout(n38983));
  jnot g21721(.din(n38610), .dout(n38984));
  jnot g21722(.din(n38615), .dout(n38985));
  jnot g21723(.din(n38620), .dout(n38986));
  jnot g21724(.din(n38625), .dout(n38987));
  jnot g21725(.din(n38630), .dout(n38988));
  jnot g21726(.din(n38635), .dout(n38989));
  jnot g21727(.din(n38640), .dout(n38990));
  jnot g21728(.din(n38645), .dout(n38991));
  jnot g21729(.din(n38650), .dout(n38992));
  jnot g21730(.din(n38655), .dout(n38993));
  jnot g21731(.din(n38660), .dout(n38994));
  jnot g21732(.din(n38665), .dout(n38995));
  jnot g21733(.din(n38670), .dout(n38996));
  jnot g21734(.din(n38675), .dout(n38997));
  jnot g21735(.din(n38680), .dout(n38998));
  jnot g21736(.din(n38685), .dout(n38999));
  jnot g21737(.din(n38690), .dout(n39000));
  jnot g21738(.din(n38695), .dout(n39001));
  jnot g21739(.din(n38700), .dout(n39002));
  jnot g21740(.din(n38705), .dout(n39003));
  jnot g21741(.din(n38710), .dout(n39004));
  jnot g21742(.din(n38715), .dout(n39005));
  jnot g21743(.din(n38720), .dout(n39006));
  jnot g21744(.din(n38725), .dout(n39007));
  jnot g21745(.din(n38730), .dout(n39008));
  jnot g21746(.din(n38735), .dout(n39009));
  jnot g21747(.din(n38740), .dout(n39010));
  jnot g21748(.din(n38745), .dout(n39011));
  jnot g21749(.din(n38750), .dout(n39012));
  jor  g21750(.dina(n38761), .dinb(b1 ), .dout(n39013));
  jnot g21751(.din(n17823), .dout(n39014));
  jxor g21752(.dina(n38761), .dinb(n259), .dout(n39015));
  jor  g21753(.dina(n39015), .dinb(n39014), .dout(n39016));
  jand g21754(.dina(n39016), .dinb(n39013), .dout(n39017));
  jxor g21755(.dina(n38755), .dinb(n386), .dout(n39018));
  jor  g21756(.dina(n39018), .dinb(n39017), .dout(n39019));
  jand g21757(.dina(n39019), .dinb(n38756), .dout(n39020));
  jnot g21758(.din(n38768), .dout(n39021));
  jor  g21759(.dina(n39021), .dinb(n39020), .dout(n39022));
  jand g21760(.dina(n39022), .dinb(n39012), .dout(n39023));
  jnot g21761(.din(n38771), .dout(n39024));
  jor  g21762(.dina(n39024), .dinb(n39023), .dout(n39025));
  jand g21763(.dina(n39025), .dinb(n39011), .dout(n39026));
  jnot g21764(.din(n38774), .dout(n39027));
  jor  g21765(.dina(n39027), .dinb(n39026), .dout(n39028));
  jand g21766(.dina(n39028), .dinb(n39010), .dout(n39029));
  jnot g21767(.din(n38777), .dout(n39030));
  jor  g21768(.dina(n39030), .dinb(n39029), .dout(n39031));
  jand g21769(.dina(n39031), .dinb(n39009), .dout(n39032));
  jnot g21770(.din(n38780), .dout(n39033));
  jor  g21771(.dina(n39033), .dinb(n39032), .dout(n39034));
  jand g21772(.dina(n39034), .dinb(n39008), .dout(n39035));
  jnot g21773(.din(n38783), .dout(n39036));
  jor  g21774(.dina(n39036), .dinb(n39035), .dout(n39037));
  jand g21775(.dina(n39037), .dinb(n39007), .dout(n39038));
  jnot g21776(.din(n38786), .dout(n39039));
  jor  g21777(.dina(n39039), .dinb(n39038), .dout(n39040));
  jand g21778(.dina(n39040), .dinb(n39006), .dout(n39041));
  jnot g21779(.din(n38789), .dout(n39042));
  jor  g21780(.dina(n39042), .dinb(n39041), .dout(n39043));
  jand g21781(.dina(n39043), .dinb(n39005), .dout(n39044));
  jnot g21782(.din(n38792), .dout(n39045));
  jor  g21783(.dina(n39045), .dinb(n39044), .dout(n39046));
  jand g21784(.dina(n39046), .dinb(n39004), .dout(n39047));
  jnot g21785(.din(n38795), .dout(n39048));
  jor  g21786(.dina(n39048), .dinb(n39047), .dout(n39049));
  jand g21787(.dina(n39049), .dinb(n39003), .dout(n39050));
  jnot g21788(.din(n38798), .dout(n39051));
  jor  g21789(.dina(n39051), .dinb(n39050), .dout(n39052));
  jand g21790(.dina(n39052), .dinb(n39002), .dout(n39053));
  jnot g21791(.din(n38801), .dout(n39054));
  jor  g21792(.dina(n39054), .dinb(n39053), .dout(n39055));
  jand g21793(.dina(n39055), .dinb(n39001), .dout(n39056));
  jnot g21794(.din(n38804), .dout(n39057));
  jor  g21795(.dina(n39057), .dinb(n39056), .dout(n39058));
  jand g21796(.dina(n39058), .dinb(n39000), .dout(n39059));
  jnot g21797(.din(n38807), .dout(n39060));
  jor  g21798(.dina(n39060), .dinb(n39059), .dout(n39061));
  jand g21799(.dina(n39061), .dinb(n38999), .dout(n39062));
  jnot g21800(.din(n38810), .dout(n39063));
  jor  g21801(.dina(n39063), .dinb(n39062), .dout(n39064));
  jand g21802(.dina(n39064), .dinb(n38998), .dout(n39065));
  jnot g21803(.din(n38813), .dout(n39066));
  jor  g21804(.dina(n39066), .dinb(n39065), .dout(n39067));
  jand g21805(.dina(n39067), .dinb(n38997), .dout(n39068));
  jnot g21806(.din(n38816), .dout(n39069));
  jor  g21807(.dina(n39069), .dinb(n39068), .dout(n39070));
  jand g21808(.dina(n39070), .dinb(n38996), .dout(n39071));
  jnot g21809(.din(n38819), .dout(n39072));
  jor  g21810(.dina(n39072), .dinb(n39071), .dout(n39073));
  jand g21811(.dina(n39073), .dinb(n38995), .dout(n39074));
  jnot g21812(.din(n38822), .dout(n39075));
  jor  g21813(.dina(n39075), .dinb(n39074), .dout(n39076));
  jand g21814(.dina(n39076), .dinb(n38994), .dout(n39077));
  jnot g21815(.din(n38825), .dout(n39078));
  jor  g21816(.dina(n39078), .dinb(n39077), .dout(n39079));
  jand g21817(.dina(n39079), .dinb(n38993), .dout(n39080));
  jnot g21818(.din(n38828), .dout(n39081));
  jor  g21819(.dina(n39081), .dinb(n39080), .dout(n39082));
  jand g21820(.dina(n39082), .dinb(n38992), .dout(n39083));
  jnot g21821(.din(n38831), .dout(n39084));
  jor  g21822(.dina(n39084), .dinb(n39083), .dout(n39085));
  jand g21823(.dina(n39085), .dinb(n38991), .dout(n39086));
  jnot g21824(.din(n38834), .dout(n39087));
  jor  g21825(.dina(n39087), .dinb(n39086), .dout(n39088));
  jand g21826(.dina(n39088), .dinb(n38990), .dout(n39089));
  jnot g21827(.din(n38837), .dout(n39090));
  jor  g21828(.dina(n39090), .dinb(n39089), .dout(n39091));
  jand g21829(.dina(n39091), .dinb(n38989), .dout(n39092));
  jnot g21830(.din(n38840), .dout(n39093));
  jor  g21831(.dina(n39093), .dinb(n39092), .dout(n39094));
  jand g21832(.dina(n39094), .dinb(n38988), .dout(n39095));
  jnot g21833(.din(n38843), .dout(n39096));
  jor  g21834(.dina(n39096), .dinb(n39095), .dout(n39097));
  jand g21835(.dina(n39097), .dinb(n38987), .dout(n39098));
  jnot g21836(.din(n38846), .dout(n39099));
  jor  g21837(.dina(n39099), .dinb(n39098), .dout(n39100));
  jand g21838(.dina(n39100), .dinb(n38986), .dout(n39101));
  jnot g21839(.din(n38849), .dout(n39102));
  jor  g21840(.dina(n39102), .dinb(n39101), .dout(n39103));
  jand g21841(.dina(n39103), .dinb(n38985), .dout(n39104));
  jnot g21842(.din(n38852), .dout(n39105));
  jor  g21843(.dina(n39105), .dinb(n39104), .dout(n39106));
  jand g21844(.dina(n39106), .dinb(n38984), .dout(n39107));
  jnot g21845(.din(n38855), .dout(n39108));
  jor  g21846(.dina(n39108), .dinb(n39107), .dout(n39109));
  jand g21847(.dina(n39109), .dinb(n38983), .dout(n39110));
  jnot g21848(.din(n38858), .dout(n39111));
  jor  g21849(.dina(n39111), .dinb(n39110), .dout(n39112));
  jand g21850(.dina(n39112), .dinb(n38982), .dout(n39113));
  jnot g21851(.din(n38861), .dout(n39114));
  jor  g21852(.dina(n39114), .dinb(n39113), .dout(n39115));
  jand g21853(.dina(n39115), .dinb(n38981), .dout(n39116));
  jnot g21854(.din(n38864), .dout(n39117));
  jor  g21855(.dina(n39117), .dinb(n39116), .dout(n39118));
  jand g21856(.dina(n39118), .dinb(n38980), .dout(n39119));
  jnot g21857(.din(n38867), .dout(n39120));
  jor  g21858(.dina(n39120), .dinb(n39119), .dout(n39121));
  jand g21859(.dina(n39121), .dinb(n38979), .dout(n39122));
  jnot g21860(.din(n38870), .dout(n39123));
  jor  g21861(.dina(n39123), .dinb(n39122), .dout(n39124));
  jand g21862(.dina(n39124), .dinb(n38978), .dout(n39125));
  jnot g21863(.din(n38873), .dout(n39126));
  jor  g21864(.dina(n39126), .dinb(n39125), .dout(n39127));
  jand g21865(.dina(n39127), .dinb(n38977), .dout(n39128));
  jnot g21866(.din(n38876), .dout(n39129));
  jor  g21867(.dina(n39129), .dinb(n39128), .dout(n39130));
  jand g21868(.dina(n39130), .dinb(n38976), .dout(n39131));
  jnot g21869(.din(n38879), .dout(n39132));
  jor  g21870(.dina(n39132), .dinb(n39131), .dout(n39133));
  jand g21871(.dina(n39133), .dinb(n38975), .dout(n39134));
  jnot g21872(.din(n38882), .dout(n39135));
  jor  g21873(.dina(n39135), .dinb(n39134), .dout(n39136));
  jand g21874(.dina(n39136), .dinb(n38974), .dout(n39137));
  jnot g21875(.din(n38885), .dout(n39138));
  jor  g21876(.dina(n39138), .dinb(n39137), .dout(n39139));
  jand g21877(.dina(n39139), .dinb(n38973), .dout(n39140));
  jnot g21878(.din(n38888), .dout(n39141));
  jor  g21879(.dina(n39141), .dinb(n39140), .dout(n39142));
  jand g21880(.dina(n39142), .dinb(n38972), .dout(n39143));
  jnot g21881(.din(n38891), .dout(n39144));
  jor  g21882(.dina(n39144), .dinb(n39143), .dout(n39145));
  jand g21883(.dina(n39145), .dinb(n38971), .dout(n39146));
  jnot g21884(.din(n38894), .dout(n39147));
  jor  g21885(.dina(n39147), .dinb(n39146), .dout(n39148));
  jand g21886(.dina(n39148), .dinb(n38970), .dout(n39149));
  jnot g21887(.din(n38897), .dout(n39150));
  jor  g21888(.dina(n39150), .dinb(n39149), .dout(n39151));
  jand g21889(.dina(n39151), .dinb(n38969), .dout(n39152));
  jnot g21890(.din(n38900), .dout(n39153));
  jor  g21891(.dina(n39153), .dinb(n39152), .dout(n39154));
  jand g21892(.dina(n39154), .dinb(n38968), .dout(n39155));
  jnot g21893(.din(n38903), .dout(n39156));
  jor  g21894(.dina(n39156), .dinb(n39155), .dout(n39157));
  jand g21895(.dina(n39157), .dinb(n38967), .dout(n39158));
  jnot g21896(.din(n38906), .dout(n39159));
  jor  g21897(.dina(n39159), .dinb(n39158), .dout(n39160));
  jand g21898(.dina(n39160), .dinb(n38966), .dout(n39161));
  jnot g21899(.din(n38909), .dout(n39162));
  jor  g21900(.dina(n39162), .dinb(n39161), .dout(n39163));
  jand g21901(.dina(n39163), .dinb(n38965), .dout(n39164));
  jnot g21902(.din(n38912), .dout(n39165));
  jor  g21903(.dina(n39165), .dinb(n39164), .dout(n39166));
  jand g21904(.dina(n39166), .dinb(n38964), .dout(n39167));
  jnot g21905(.din(n38915), .dout(n39168));
  jor  g21906(.dina(n39168), .dinb(n39167), .dout(n39169));
  jand g21907(.dina(n39169), .dinb(n38963), .dout(n39170));
  jnot g21908(.din(n38918), .dout(n39171));
  jor  g21909(.dina(n39171), .dinb(n39170), .dout(n39172));
  jand g21910(.dina(n39172), .dinb(n38962), .dout(n39173));
  jnot g21911(.din(n38921), .dout(n39174));
  jor  g21912(.dina(n39174), .dinb(n39173), .dout(n39175));
  jand g21913(.dina(n39175), .dinb(n38961), .dout(n39176));
  jnot g21914(.din(n38924), .dout(n39177));
  jor  g21915(.dina(n39177), .dinb(n39176), .dout(n39178));
  jand g21916(.dina(n39178), .dinb(n38960), .dout(n39179));
  jnot g21917(.din(n38927), .dout(n39180));
  jor  g21918(.dina(n39180), .dinb(n39179), .dout(n39181));
  jand g21919(.dina(n39181), .dinb(n38959), .dout(n39182));
  jnot g21920(.din(n38930), .dout(n39183));
  jor  g21921(.dina(n39183), .dinb(n39182), .dout(n39184));
  jand g21922(.dina(n39184), .dinb(n38958), .dout(n39185));
  jnot g21923(.din(n38933), .dout(n39186));
  jor  g21924(.dina(n39186), .dinb(n39185), .dout(n39187));
  jand g21925(.dina(n39187), .dinb(n38957), .dout(n39188));
  jnot g21926(.din(n38936), .dout(n39189));
  jor  g21927(.dina(n39189), .dinb(n39188), .dout(n39190));
  jand g21928(.dina(n39190), .dinb(n38956), .dout(n39191));
  jnot g21929(.din(n38939), .dout(n39192));
  jor  g21930(.dina(n39192), .dinb(n39191), .dout(n39193));
  jand g21931(.dina(n39193), .dinb(n38955), .dout(n39194));
  jnot g21932(.din(n38942), .dout(n39195));
  jor  g21933(.dina(n39195), .dinb(n39194), .dout(n39196));
  jand g21934(.dina(n39196), .dinb(n38954), .dout(n39197));
  jnot g21935(.din(n38945), .dout(n39198));
  jor  g21936(.dina(n39198), .dinb(n39197), .dout(n39199));
  jand g21937(.dina(n39199), .dinb(n38953), .dout(n39200));
  jor  g21938(.dina(n39200), .dinb(n38449), .dout(n39201));
  jand g21939(.dina(n39201), .dinb(n38952), .dout(n39202));
  jand g21940(.dina(n39202), .dinb(n38759), .dout(n39203));
  jxor g21941(.dina(n38762), .dinb(n17823), .dout(n39204));
  jand g21942(.dina(n39204), .dinb(n38949), .dout(n39205));
  jor  g21943(.dina(n39205), .dinb(n39203), .dout(remainder1 ));
  jnot g21944(.din(n38755), .dout(n39207));
  jor  g21945(.dina(n38949), .dinb(n39207), .dout(n39208));
  jxor g21946(.dina(n38765), .dinb(n38764), .dout(n39209));
  jor  g21947(.dina(n39209), .dinb(n39202), .dout(n39210));
  jand g21948(.dina(n39210), .dinb(n39208), .dout(remainder2 ));
  jor  g21949(.dina(n38949), .dinb(n38749), .dout(n39212));
  jxor g21950(.dina(n38768), .dinb(n38767), .dout(n39213));
  jor  g21951(.dina(n39213), .dinb(n39202), .dout(n39214));
  jand g21952(.dina(n39214), .dinb(n39212), .dout(remainder3 ));
  jor  g21953(.dina(n38949), .dinb(n38744), .dout(n39216));
  jxor g21954(.dina(n38771), .dinb(n38770), .dout(n39217));
  jor  g21955(.dina(n39217), .dinb(n39202), .dout(n39218));
  jand g21956(.dina(n39218), .dinb(n39216), .dout(remainder4 ));
  jor  g21957(.dina(n38949), .dinb(n38739), .dout(n39220));
  jxor g21958(.dina(n38774), .dinb(n38773), .dout(n39221));
  jor  g21959(.dina(n39221), .dinb(n39202), .dout(n39222));
  jand g21960(.dina(n39222), .dinb(n39220), .dout(remainder5 ));
  jor  g21961(.dina(n38949), .dinb(n38734), .dout(n39224));
  jxor g21962(.dina(n38777), .dinb(n38776), .dout(n39225));
  jor  g21963(.dina(n39225), .dinb(n39202), .dout(n39226));
  jand g21964(.dina(n39226), .dinb(n39224), .dout(remainder6 ));
  jor  g21965(.dina(n38949), .dinb(n38729), .dout(n39228));
  jxor g21966(.dina(n38780), .dinb(n38779), .dout(n39229));
  jor  g21967(.dina(n39229), .dinb(n39202), .dout(n39230));
  jand g21968(.dina(n39230), .dinb(n39228), .dout(remainder7 ));
  jor  g21969(.dina(n38949), .dinb(n38724), .dout(n39232));
  jxor g21970(.dina(n38783), .dinb(n38782), .dout(n39233));
  jor  g21971(.dina(n39233), .dinb(n39202), .dout(n39234));
  jand g21972(.dina(n39234), .dinb(n39232), .dout(remainder8 ));
  jor  g21973(.dina(n38949), .dinb(n38719), .dout(n39236));
  jxor g21974(.dina(n38786), .dinb(n38785), .dout(n39237));
  jor  g21975(.dina(n39237), .dinb(n39202), .dout(n39238));
  jand g21976(.dina(n39238), .dinb(n39236), .dout(remainder9 ));
  jor  g21977(.dina(n38949), .dinb(n38714), .dout(n39240));
  jxor g21978(.dina(n38789), .dinb(n38788), .dout(n39241));
  jor  g21979(.dina(n39241), .dinb(n39202), .dout(n39242));
  jand g21980(.dina(n39242), .dinb(n39240), .dout(remainder10 ));
  jor  g21981(.dina(n38949), .dinb(n38709), .dout(n39244));
  jxor g21982(.dina(n38792), .dinb(n38791), .dout(n39245));
  jor  g21983(.dina(n39245), .dinb(n39202), .dout(n39246));
  jand g21984(.dina(n39246), .dinb(n39244), .dout(remainder11 ));
  jor  g21985(.dina(n38949), .dinb(n38704), .dout(n39248));
  jxor g21986(.dina(n38795), .dinb(n38794), .dout(n39249));
  jor  g21987(.dina(n39249), .dinb(n39202), .dout(n39250));
  jand g21988(.dina(n39250), .dinb(n39248), .dout(remainder12 ));
  jor  g21989(.dina(n38949), .dinb(n38699), .dout(n39252));
  jxor g21990(.dina(n38798), .dinb(n38797), .dout(n39253));
  jor  g21991(.dina(n39253), .dinb(n39202), .dout(n39254));
  jand g21992(.dina(n39254), .dinb(n39252), .dout(remainder13 ));
  jor  g21993(.dina(n38949), .dinb(n38694), .dout(n39256));
  jxor g21994(.dina(n38801), .dinb(n38800), .dout(n39257));
  jor  g21995(.dina(n39257), .dinb(n39202), .dout(n39258));
  jand g21996(.dina(n39258), .dinb(n39256), .dout(remainder14 ));
  jor  g21997(.dina(n38949), .dinb(n38689), .dout(n39260));
  jxor g21998(.dina(n38804), .dinb(n38803), .dout(n39261));
  jor  g21999(.dina(n39261), .dinb(n39202), .dout(n39262));
  jand g22000(.dina(n39262), .dinb(n39260), .dout(remainder15 ));
  jor  g22001(.dina(n38949), .dinb(n38684), .dout(n39264));
  jxor g22002(.dina(n38807), .dinb(n38806), .dout(n39265));
  jor  g22003(.dina(n39265), .dinb(n39202), .dout(n39266));
  jand g22004(.dina(n39266), .dinb(n39264), .dout(remainder16 ));
  jor  g22005(.dina(n38949), .dinb(n38679), .dout(n39268));
  jxor g22006(.dina(n38810), .dinb(n38809), .dout(n39269));
  jor  g22007(.dina(n39269), .dinb(n39202), .dout(n39270));
  jand g22008(.dina(n39270), .dinb(n39268), .dout(remainder17 ));
  jor  g22009(.dina(n38949), .dinb(n38674), .dout(n39272));
  jxor g22010(.dina(n38813), .dinb(n38812), .dout(n39273));
  jor  g22011(.dina(n39273), .dinb(n39202), .dout(n39274));
  jand g22012(.dina(n39274), .dinb(n39272), .dout(remainder18 ));
  jor  g22013(.dina(n38949), .dinb(n38669), .dout(n39276));
  jxor g22014(.dina(n38816), .dinb(n38815), .dout(n39277));
  jor  g22015(.dina(n39277), .dinb(n39202), .dout(n39278));
  jand g22016(.dina(n39278), .dinb(n39276), .dout(remainder19 ));
  jor  g22017(.dina(n38949), .dinb(n38664), .dout(n39280));
  jxor g22018(.dina(n38819), .dinb(n38818), .dout(n39281));
  jor  g22019(.dina(n39281), .dinb(n39202), .dout(n39282));
  jand g22020(.dina(n39282), .dinb(n39280), .dout(remainder20 ));
  jor  g22021(.dina(n38949), .dinb(n38659), .dout(n39284));
  jxor g22022(.dina(n38822), .dinb(n38821), .dout(n39285));
  jor  g22023(.dina(n39285), .dinb(n39202), .dout(n39286));
  jand g22024(.dina(n39286), .dinb(n39284), .dout(remainder21 ));
  jor  g22025(.dina(n38949), .dinb(n38654), .dout(n39288));
  jxor g22026(.dina(n38825), .dinb(n38824), .dout(n39289));
  jor  g22027(.dina(n39289), .dinb(n39202), .dout(n39290));
  jand g22028(.dina(n39290), .dinb(n39288), .dout(remainder22 ));
  jor  g22029(.dina(n38949), .dinb(n38649), .dout(n39292));
  jxor g22030(.dina(n38828), .dinb(n38827), .dout(n39293));
  jor  g22031(.dina(n39293), .dinb(n39202), .dout(n39294));
  jand g22032(.dina(n39294), .dinb(n39292), .dout(remainder23 ));
  jor  g22033(.dina(n38949), .dinb(n38644), .dout(n39296));
  jxor g22034(.dina(n38831), .dinb(n38830), .dout(n39297));
  jor  g22035(.dina(n39297), .dinb(n39202), .dout(n39298));
  jand g22036(.dina(n39298), .dinb(n39296), .dout(remainder24 ));
  jor  g22037(.dina(n38949), .dinb(n38639), .dout(n39300));
  jxor g22038(.dina(n38834), .dinb(n38833), .dout(n39301));
  jor  g22039(.dina(n39301), .dinb(n39202), .dout(n39302));
  jand g22040(.dina(n39302), .dinb(n39300), .dout(remainder25 ));
  jor  g22041(.dina(n38949), .dinb(n38634), .dout(n39304));
  jxor g22042(.dina(n38837), .dinb(n38836), .dout(n39305));
  jor  g22043(.dina(n39305), .dinb(n39202), .dout(n39306));
  jand g22044(.dina(n39306), .dinb(n39304), .dout(remainder26 ));
  jor  g22045(.dina(n38949), .dinb(n38629), .dout(n39308));
  jxor g22046(.dina(n38840), .dinb(n38839), .dout(n39309));
  jor  g22047(.dina(n39309), .dinb(n39202), .dout(n39310));
  jand g22048(.dina(n39310), .dinb(n39308), .dout(remainder27 ));
  jor  g22049(.dina(n38949), .dinb(n38624), .dout(n39312));
  jxor g22050(.dina(n38843), .dinb(n38842), .dout(n39313));
  jor  g22051(.dina(n39313), .dinb(n39202), .dout(n39314));
  jand g22052(.dina(n39314), .dinb(n39312), .dout(remainder28 ));
  jor  g22053(.dina(n38949), .dinb(n38619), .dout(n39316));
  jxor g22054(.dina(n38846), .dinb(n38845), .dout(n39317));
  jor  g22055(.dina(n39317), .dinb(n39202), .dout(n39318));
  jand g22056(.dina(n39318), .dinb(n39316), .dout(remainder29 ));
  jor  g22057(.dina(n38949), .dinb(n38614), .dout(n39320));
  jxor g22058(.dina(n38849), .dinb(n38848), .dout(n39321));
  jor  g22059(.dina(n39321), .dinb(n39202), .dout(n39322));
  jand g22060(.dina(n39322), .dinb(n39320), .dout(remainder30 ));
  jor  g22061(.dina(n38949), .dinb(n38609), .dout(n39324));
  jxor g22062(.dina(n38852), .dinb(n38851), .dout(n39325));
  jor  g22063(.dina(n39325), .dinb(n39202), .dout(n39326));
  jand g22064(.dina(n39326), .dinb(n39324), .dout(remainder31 ));
  jor  g22065(.dina(n38949), .dinb(n38604), .dout(n39328));
  jxor g22066(.dina(n38855), .dinb(n38854), .dout(n39329));
  jor  g22067(.dina(n39329), .dinb(n39202), .dout(n39330));
  jand g22068(.dina(n39330), .dinb(n39328), .dout(remainder32 ));
  jor  g22069(.dina(n38949), .dinb(n38599), .dout(n39332));
  jxor g22070(.dina(n38858), .dinb(n38857), .dout(n39333));
  jor  g22071(.dina(n39333), .dinb(n39202), .dout(n39334));
  jand g22072(.dina(n39334), .dinb(n39332), .dout(remainder33 ));
  jor  g22073(.dina(n38949), .dinb(n38594), .dout(n39336));
  jxor g22074(.dina(n38861), .dinb(n38860), .dout(n39337));
  jor  g22075(.dina(n39337), .dinb(n39202), .dout(n39338));
  jand g22076(.dina(n39338), .dinb(n39336), .dout(remainder34 ));
  jor  g22077(.dina(n38949), .dinb(n38589), .dout(n39340));
  jxor g22078(.dina(n38864), .dinb(n38863), .dout(n39341));
  jor  g22079(.dina(n39341), .dinb(n39202), .dout(n39342));
  jand g22080(.dina(n39342), .dinb(n39340), .dout(remainder35 ));
  jor  g22081(.dina(n38949), .dinb(n38584), .dout(n39344));
  jxor g22082(.dina(n38867), .dinb(n38866), .dout(n39345));
  jor  g22083(.dina(n39345), .dinb(n39202), .dout(n39346));
  jand g22084(.dina(n39346), .dinb(n39344), .dout(remainder36 ));
  jor  g22085(.dina(n38949), .dinb(n38579), .dout(n39348));
  jxor g22086(.dina(n38870), .dinb(n38869), .dout(n39349));
  jor  g22087(.dina(n39349), .dinb(n39202), .dout(n39350));
  jand g22088(.dina(n39350), .dinb(n39348), .dout(remainder37 ));
  jor  g22089(.dina(n38949), .dinb(n38574), .dout(n39352));
  jxor g22090(.dina(n38873), .dinb(n38872), .dout(n39353));
  jor  g22091(.dina(n39353), .dinb(n39202), .dout(n39354));
  jand g22092(.dina(n39354), .dinb(n39352), .dout(remainder38 ));
  jor  g22093(.dina(n38949), .dinb(n38569), .dout(n39356));
  jxor g22094(.dina(n38876), .dinb(n38875), .dout(n39357));
  jor  g22095(.dina(n39357), .dinb(n39202), .dout(n39358));
  jand g22096(.dina(n39358), .dinb(n39356), .dout(remainder39 ));
  jor  g22097(.dina(n38949), .dinb(n38564), .dout(n39360));
  jxor g22098(.dina(n38879), .dinb(n38878), .dout(n39361));
  jor  g22099(.dina(n39361), .dinb(n39202), .dout(n39362));
  jand g22100(.dina(n39362), .dinb(n39360), .dout(remainder40 ));
  jor  g22101(.dina(n38949), .dinb(n38559), .dout(n39364));
  jxor g22102(.dina(n38882), .dinb(n38881), .dout(n39365));
  jor  g22103(.dina(n39365), .dinb(n39202), .dout(n39366));
  jand g22104(.dina(n39366), .dinb(n39364), .dout(remainder41 ));
  jor  g22105(.dina(n38949), .dinb(n38554), .dout(n39368));
  jxor g22106(.dina(n38885), .dinb(n38884), .dout(n39369));
  jor  g22107(.dina(n39369), .dinb(n39202), .dout(n39370));
  jand g22108(.dina(n39370), .dinb(n39368), .dout(remainder42 ));
  jor  g22109(.dina(n38949), .dinb(n38549), .dout(n39372));
  jxor g22110(.dina(n38888), .dinb(n38887), .dout(n39373));
  jor  g22111(.dina(n39373), .dinb(n39202), .dout(n39374));
  jand g22112(.dina(n39374), .dinb(n39372), .dout(remainder43 ));
  jor  g22113(.dina(n38949), .dinb(n38544), .dout(n39376));
  jxor g22114(.dina(n38891), .dinb(n38890), .dout(n39377));
  jor  g22115(.dina(n39377), .dinb(n39202), .dout(n39378));
  jand g22116(.dina(n39378), .dinb(n39376), .dout(remainder44 ));
  jor  g22117(.dina(n38949), .dinb(n38539), .dout(n39380));
  jxor g22118(.dina(n38894), .dinb(n38893), .dout(n39381));
  jor  g22119(.dina(n39381), .dinb(n39202), .dout(n39382));
  jand g22120(.dina(n39382), .dinb(n39380), .dout(remainder45 ));
  jor  g22121(.dina(n38949), .dinb(n38534), .dout(n39384));
  jxor g22122(.dina(n38897), .dinb(n38896), .dout(n39385));
  jor  g22123(.dina(n39385), .dinb(n39202), .dout(n39386));
  jand g22124(.dina(n39386), .dinb(n39384), .dout(remainder46 ));
  jor  g22125(.dina(n38949), .dinb(n38529), .dout(n39388));
  jxor g22126(.dina(n38900), .dinb(n38899), .dout(n39389));
  jor  g22127(.dina(n39389), .dinb(n39202), .dout(n39390));
  jand g22128(.dina(n39390), .dinb(n39388), .dout(remainder47 ));
  jor  g22129(.dina(n38949), .dinb(n38524), .dout(n39392));
  jxor g22130(.dina(n38903), .dinb(n38902), .dout(n39393));
  jor  g22131(.dina(n39393), .dinb(n39202), .dout(n39394));
  jand g22132(.dina(n39394), .dinb(n39392), .dout(remainder48 ));
  jor  g22133(.dina(n38949), .dinb(n38519), .dout(n39396));
  jxor g22134(.dina(n38906), .dinb(n38905), .dout(n39397));
  jor  g22135(.dina(n39397), .dinb(n39202), .dout(n39398));
  jand g22136(.dina(n39398), .dinb(n39396), .dout(remainder49 ));
  jor  g22137(.dina(n38949), .dinb(n38514), .dout(n39400));
  jxor g22138(.dina(n38909), .dinb(n38908), .dout(n39401));
  jor  g22139(.dina(n39401), .dinb(n39202), .dout(n39402));
  jand g22140(.dina(n39402), .dinb(n39400), .dout(remainder50 ));
  jor  g22141(.dina(n38949), .dinb(n38509), .dout(n39404));
  jxor g22142(.dina(n38912), .dinb(n38911), .dout(n39405));
  jor  g22143(.dina(n39405), .dinb(n39202), .dout(n39406));
  jand g22144(.dina(n39406), .dinb(n39404), .dout(remainder51 ));
  jor  g22145(.dina(n38949), .dinb(n38504), .dout(n39408));
  jxor g22146(.dina(n38915), .dinb(n38914), .dout(n39409));
  jor  g22147(.dina(n39409), .dinb(n39202), .dout(n39410));
  jand g22148(.dina(n39410), .dinb(n39408), .dout(remainder52 ));
  jor  g22149(.dina(n38949), .dinb(n38499), .dout(n39412));
  jxor g22150(.dina(n38918), .dinb(n38917), .dout(n39413));
  jor  g22151(.dina(n39413), .dinb(n39202), .dout(n39414));
  jand g22152(.dina(n39414), .dinb(n39412), .dout(remainder53 ));
  jor  g22153(.dina(n38949), .dinb(n38494), .dout(n39416));
  jxor g22154(.dina(n38921), .dinb(n38920), .dout(n39417));
  jor  g22155(.dina(n39417), .dinb(n39202), .dout(n39418));
  jand g22156(.dina(n39418), .dinb(n39416), .dout(remainder54 ));
  jor  g22157(.dina(n38949), .dinb(n38489), .dout(n39420));
  jxor g22158(.dina(n38924), .dinb(n38923), .dout(n39421));
  jor  g22159(.dina(n39421), .dinb(n39202), .dout(n39422));
  jand g22160(.dina(n39422), .dinb(n39420), .dout(remainder55 ));
  jor  g22161(.dina(n38949), .dinb(n38484), .dout(n39424));
  jxor g22162(.dina(n38927), .dinb(n38926), .dout(n39425));
  jor  g22163(.dina(n39425), .dinb(n39202), .dout(n39426));
  jand g22164(.dina(n39426), .dinb(n39424), .dout(remainder56 ));
  jor  g22165(.dina(n38949), .dinb(n38479), .dout(n39428));
  jxor g22166(.dina(n38930), .dinb(n38929), .dout(n39429));
  jor  g22167(.dina(n39429), .dinb(n39202), .dout(n39430));
  jand g22168(.dina(n39430), .dinb(n39428), .dout(remainder57 ));
  jor  g22169(.dina(n38949), .dinb(n38474), .dout(n39432));
  jxor g22170(.dina(n38933), .dinb(n38932), .dout(n39433));
  jor  g22171(.dina(n39433), .dinb(n39202), .dout(n39434));
  jand g22172(.dina(n39434), .dinb(n39432), .dout(remainder58 ));
  jor  g22173(.dina(n38949), .dinb(n38469), .dout(n39436));
  jxor g22174(.dina(n38936), .dinb(n38935), .dout(n39437));
  jor  g22175(.dina(n39437), .dinb(n39202), .dout(n39438));
  jand g22176(.dina(n39438), .dinb(n39436), .dout(remainder59 ));
  jor  g22177(.dina(n38949), .dinb(n38464), .dout(n39440));
  jxor g22178(.dina(n38939), .dinb(n38938), .dout(n39441));
  jor  g22179(.dina(n39441), .dinb(n39202), .dout(n39442));
  jand g22180(.dina(n39442), .dinb(n39440), .dout(remainder60 ));
  jor  g22181(.dina(n38949), .dinb(n38459), .dout(n39444));
  jxor g22182(.dina(n38942), .dinb(n38941), .dout(n39445));
  jor  g22183(.dina(n39445), .dinb(n39202), .dout(n39446));
  jand g22184(.dina(n39446), .dinb(n39444), .dout(remainder61 ));
  jor  g22185(.dina(n38949), .dinb(n38454), .dout(n39448));
  jxor g22186(.dina(n38945), .dinb(n38944), .dout(n39449));
  jor  g22187(.dina(n39449), .dinb(n39202), .dout(n39450));
  jand g22188(.dina(n39450), .dinb(n39448), .dout(remainder62 ));
  jand g22189(.dina(n39202), .dinb(n38447), .dout(n39452));
  jand g22190(.dina(n38947), .dinb(n38448), .dout(n39453));
  jor  g22191(.dina(n39453), .dinb(n39452), .dout(remainder63 ));
endmodule


