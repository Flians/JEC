/*

c5315:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jdff: 3497
	jand: 606
	jor: 486

Summary:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jdff: 3497
	jand: 606
	jor: 486

The maximum logic level gap of any gate:
	c5315: 22
*/

module gf_c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[1:0] w_G1_2;
	wire[2:0] w_G4_0;
	wire[1:0] w_G11_0;
	wire[1:0] w_G14_0;
	wire[1:0] w_G17_0;
	wire[1:0] w_G20_0;
	wire[1:0] w_G37_0;
	wire[1:0] w_G40_0;
	wire[1:0] w_G43_0;
	wire[1:0] w_G46_0;
	wire[1:0] w_G49_0;
	wire[2:0] w_G54_0;
	wire[1:0] w_G61_0;
	wire[1:0] w_G64_0;
	wire[1:0] w_G67_0;
	wire[1:0] w_G70_0;
	wire[1:0] w_G73_0;
	wire[1:0] w_G76_0;
	wire[1:0] w_G91_0;
	wire[1:0] w_G100_0;
	wire[1:0] w_G103_0;
	wire[1:0] w_G106_0;
	wire[1:0] w_G109_0;
	wire[1:0] w_G123_0;
	wire[2:0] w_G137_0;
	wire[2:0] w_G137_1;
	wire[2:0] w_G137_2;
	wire[2:0] w_G137_3;
	wire[2:0] w_G137_4;
	wire[2:0] w_G137_5;
	wire[2:0] w_G137_6;
	wire[2:0] w_G137_7;
	wire[2:0] w_G137_8;
	wire[1:0] w_G137_9;
	wire[2:0] w_G141_0;
	wire[2:0] w_G141_1;
	wire[2:0] w_G141_2;
	wire[1:0] w_G146_0;
	wire[1:0] w_G149_0;
	wire[1:0] w_G152_0;
	wire[1:0] w_G155_0;
	wire[1:0] w_G158_0;
	wire[1:0] w_G161_0;
	wire[1:0] w_G164_0;
	wire[1:0] w_G167_0;
	wire[1:0] w_G170_0;
	wire[1:0] w_G173_0;
	wire[1:0] w_G182_0;
	wire[1:0] w_G185_0;
	wire[1:0] w_G188_0;
	wire[1:0] w_G191_0;
	wire[1:0] w_G194_0;
	wire[1:0] w_G197_0;
	wire[1:0] w_G200_0;
	wire[1:0] w_G203_0;
	wire[2:0] w_G206_0;
	wire[2:0] w_G206_1;
	wire[2:0] w_G210_0;
	wire[2:0] w_G210_1;
	wire[1:0] w_G210_2;
	wire[2:0] w_G218_0;
	wire[2:0] w_G218_1;
	wire[1:0] w_G218_2;
	wire[2:0] w_G226_0;
	wire[2:0] w_G226_1;
	wire[1:0] w_G226_2;
	wire[2:0] w_G234_0;
	wire[2:0] w_G234_1;
	wire[1:0] w_G234_2;
	wire[2:0] w_G242_0;
	wire[1:0] w_G242_1;
	wire[1:0] w_G245_0;
	wire[2:0] w_G248_0;
	wire[2:0] w_G248_1;
	wire[2:0] w_G248_2;
	wire[2:0] w_G248_3;
	wire[2:0] w_G248_4;
	wire[2:0] w_G248_5;
	wire[2:0] w_G251_0;
	wire[2:0] w_G251_1;
	wire[2:0] w_G251_2;
	wire[2:0] w_G251_3;
	wire[2:0] w_G251_4;
	wire[1:0] w_G251_5;
	wire[2:0] w_G254_0;
	wire[1:0] w_G254_1;
	wire[2:0] w_G257_0;
	wire[2:0] w_G257_1;
	wire[1:0] w_G257_2;
	wire[2:0] w_G265_0;
	wire[2:0] w_G265_1;
	wire[2:0] w_G273_0;
	wire[2:0] w_G273_1;
	wire[1:0] w_G273_2;
	wire[2:0] w_G281_0;
	wire[2:0] w_G281_1;
	wire[1:0] w_G281_2;
	wire[1:0] w_G289_0;
	wire[2:0] w_G293_0;
	wire[2:0] w_G299_0;
	wire[2:0] w_G302_0;
	wire[2:0] w_G308_0;
	wire[2:0] w_G308_1;
	wire[2:0] w_G316_0;
	wire[1:0] w_G316_1;
	wire[2:0] w_G324_0;
	wire[2:0] w_G324_1;
	wire[1:0] w_G331_0;
	wire[2:0] w_G332_0;
	wire[2:0] w_G332_1;
	wire[2:0] w_G332_2;
	wire[2:0] w_G332_3;
	wire[2:0] w_G335_0;
	wire[1:0] w_G338_0;
	wire[2:0] w_G341_0;
	wire[2:0] w_G341_1;
	wire[2:0] w_G341_2;
	wire[1:0] w_G348_0;
	wire[2:0] w_G351_0;
	wire[2:0] w_G351_1;
	wire[2:0] w_G351_2;
	wire[1:0] w_G358_0;
	wire[2:0] w_G361_0;
	wire[1:0] w_G361_1;
	wire[1:0] w_G366_0;
	wire[1:0] w_G369_0;
	wire[2:0] w_G374_0;
	wire[2:0] w_G374_1;
	wire[2:0] w_G389_0;
	wire[2:0] w_G389_1;
	wire[2:0] w_G400_0;
	wire[2:0] w_G400_1;
	wire[2:0] w_G411_0;
	wire[2:0] w_G411_1;
	wire[1:0] w_G411_2;
	wire[2:0] w_G422_0;
	wire[1:0] w_G422_1;
	wire[2:0] w_G435_0;
	wire[2:0] w_G435_1;
	wire[2:0] w_G446_0;
	wire[2:0] w_G446_1;
	wire[2:0] w_G457_0;
	wire[2:0] w_G457_1;
	wire[2:0] w_G468_0;
	wire[2:0] w_G468_1;
	wire[2:0] w_G479_0;
	wire[2:0] w_G490_0;
	wire[1:0] w_G490_1;
	wire[2:0] w_G503_0;
	wire[2:0] w_G503_1;
	wire[1:0] w_G503_2;
	wire[2:0] w_G514_0;
	wire[2:0] w_G514_1;
	wire[1:0] w_G514_2;
	wire[2:0] w_G523_0;
	wire[2:0] w_G523_1;
	wire[2:0] w_G534_0;
	wire[2:0] w_G534_1;
	wire[1:0] w_G534_2;
	wire[2:0] w_G545_0;
	wire[2:0] w_G549_0;
	wire[1:0] w_G552_0;
	wire[1:0] w_G559_0;
	wire[1:0] w_G562_0;
	wire[2:0] w_G1497_0;
	wire[2:0] w_G1689_0;
	wire[2:0] w_G1689_1;
	wire[2:0] w_G1689_2;
	wire[2:0] w_G1689_3;
	wire[2:0] w_G1689_4;
	wire[1:0] w_G1689_5;
	wire[2:0] w_G1690_0;
	wire[1:0] w_G1690_1;
	wire[2:0] w_G1691_0;
	wire[2:0] w_G1691_1;
	wire[2:0] w_G1691_2;
	wire[2:0] w_G1691_3;
	wire[2:0] w_G1691_4;
	wire[1:0] w_G1691_5;
	wire[2:0] w_G1694_0;
	wire[1:0] w_G1694_1;
	wire[2:0] w_G2174_0;
	wire[2:0] w_G2358_0;
	wire[2:0] w_G2358_1;
	wire[2:0] w_G2358_2;
	wire[1:0] w_G3173_0;
	wire[2:0] w_G3546_0;
	wire[2:0] w_G3546_1;
	wire[2:0] w_G3546_2;
	wire[2:0] w_G3546_3;
	wire[2:0] w_G3546_4;
	wire[1:0] w_G3546_5;
	wire[2:0] w_G3548_0;
	wire[2:0] w_G3548_1;
	wire[2:0] w_G3548_2;
	wire[2:0] w_G3548_3;
	wire[2:0] w_G3548_4;
	wire[1:0] w_G3552_0;
	wire[1:0] w_G3717_0;
	wire[2:0] w_G3724_0;
	wire[2:0] w_G4087_0;
	wire[2:0] w_G4087_1;
	wire[2:0] w_G4087_2;
	wire[2:0] w_G4087_3;
	wire[2:0] w_G4087_4;
	wire[2:0] w_G4088_0;
	wire[2:0] w_G4088_1;
	wire[2:0] w_G4088_2;
	wire[2:0] w_G4088_3;
	wire[2:0] w_G4088_4;
	wire[2:0] w_G4088_5;
	wire[2:0] w_G4088_6;
	wire[2:0] w_G4088_7;
	wire[2:0] w_G4088_8;
	wire[2:0] w_G4088_9;
	wire[2:0] w_G4089_0;
	wire[2:0] w_G4089_1;
	wire[2:0] w_G4089_2;
	wire[2:0] w_G4089_3;
	wire[2:0] w_G4089_4;
	wire[2:0] w_G4089_5;
	wire[2:0] w_G4089_6;
	wire[2:0] w_G4089_7;
	wire[2:0] w_G4089_8;
	wire[2:0] w_G4089_9;
	wire[2:0] w_G4090_0;
	wire[2:0] w_G4090_1;
	wire[2:0] w_G4090_2;
	wire[2:0] w_G4090_3;
	wire[2:0] w_G4090_4;
	wire[2:0] w_G4091_0;
	wire[2:0] w_G4091_1;
	wire[2:0] w_G4091_2;
	wire[2:0] w_G4091_3;
	wire[2:0] w_G4091_4;
	wire[2:0] w_G4091_5;
	wire[1:0] w_G4091_6;
	wire[2:0] w_G4092_0;
	wire[2:0] w_G4092_1;
	wire[2:0] w_G4092_2;
	wire[2:0] w_G4092_3;
	wire[2:0] w_G4092_4;
	wire[2:0] w_G4092_5;
	wire[2:0] w_G4092_6;
	wire[2:0] w_G4092_7;
	wire[2:0] w_G4092_8;
	wire[2:0] w_G4092_9;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire[2:0] w_G809_0;
	wire[2:0] w_G809_1;
	wire[2:0] w_G809_2;
	wire[1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G623_0;
	wire G623_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G998_0;
	wire G998_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G865_0;
	wire G865_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire[1:0] w_n316_0;
	wire[1:0] w_n318_0;
	wire[2:0] w_n326_0;
	wire[2:0] w_n326_1;
	wire[1:0] w_n326_2;
	wire[1:0] w_n333_0;
	wire[1:0] w_n336_0;
	wire[1:0] w_n361_0;
	wire[1:0] w_n365_0;
	wire[2:0] w_n366_0;
	wire[2:0] w_n366_1;
	wire[2:0] w_n369_0;
	wire[2:0] w_n369_1;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[2:0] w_n374_0;
	wire[1:0] w_n374_1;
	wire[2:0] w_n375_0;
	wire[2:0] w_n375_1;
	wire[2:0] w_n375_2;
	wire[2:0] w_n375_3;
	wire[2:0] w_n375_4;
	wire[2:0] w_n377_0;
	wire[1:0] w_n377_1;
	wire[2:0] w_n378_0;
	wire[2:0] w_n378_1;
	wire[2:0] w_n378_2;
	wire[2:0] w_n378_3;
	wire[2:0] w_n378_4;
	wire[1:0] w_n386_0;
	wire[2:0] w_n387_0;
	wire[1:0] w_n387_1;
	wire[2:0] w_n389_0;
	wire[1:0] w_n389_1;
	wire[1:0] w_n397_0;
	wire[1:0] w_n401_0;
	wire[2:0] w_n402_0;
	wire[2:0] w_n406_0;
	wire[2:0] w_n406_1;
	wire[2:0] w_n406_2;
	wire[2:0] w_n406_3;
	wire[2:0] w_n406_4;
	wire[1:0] w_n406_5;
	wire[2:0] w_n408_0;
	wire[2:0] w_n408_1;
	wire[2:0] w_n408_2;
	wire[2:0] w_n408_3;
	wire[2:0] w_n408_4;
	wire[2:0] w_n408_5;
	wire[2:0] w_n412_0;
	wire[1:0] w_n414_0;
	wire[1:0] w_n415_0;
	wire[2:0] w_n423_0;
	wire[2:0] w_n425_0;
	wire[2:0] w_n428_0;
	wire[1:0] w_n428_1;
	wire[1:0] w_n429_0;
	wire[2:0] w_n433_0;
	wire[2:0] w_n435_0;
	wire[2:0] w_n435_1;
	wire[1:0] w_n435_2;
	wire[1:0] w_n437_0;
	wire[1:0] w_n445_0;
	wire[2:0] w_n449_0;
	wire[2:0] w_n449_1;
	wire[2:0] w_n451_0;
	wire[1:0] w_n459_0;
	wire[2:0] w_n460_0;
	wire[2:0] w_n460_1;
	wire[2:0] w_n462_0;
	wire[1:0] w_n470_0;
	wire[2:0] w_n471_0;
	wire[2:0] w_n471_1;
	wire[2:0] w_n473_0;
	wire[1:0] w_n473_1;
	wire[1:0] w_n481_0;
	wire[2:0] w_n483_0;
	wire[2:0] w_n483_1;
	wire[1:0] w_n483_2;
	wire[2:0] w_n485_0;
	wire[1:0] w_n485_1;
	wire[1:0] w_n493_0;
	wire[2:0] w_n494_0;
	wire[2:0] w_n494_1;
	wire[2:0] w_n496_0;
	wire[1:0] w_n496_1;
	wire[1:0] w_n504_0;
	wire[2:0] w_n507_0;
	wire[2:0] w_n507_1;
	wire[2:0] w_n509_0;
	wire[1:0] w_n517_0;
	wire[2:0] w_n518_0;
	wire[2:0] w_n518_1;
	wire[2:0] w_n520_0;
	wire[1:0] w_n528_0;
	wire[2:0] w_n530_0;
	wire[2:0] w_n530_1;
	wire[2:0] w_n532_0;
	wire[1:0] w_n532_1;
	wire[1:0] w_n540_0;
	wire[1:0] w_n543_0;
	wire[2:0] w_n551_0;
	wire[2:0] w_n556_0;
	wire[2:0] w_n556_1;
	wire[2:0] w_n556_2;
	wire[2:0] w_n556_3;
	wire[2:0] w_n556_4;
	wire[2:0] w_n556_5;
	wire[2:0] w_n556_6;
	wire[2:0] w_n556_7;
	wire[1:0] w_n556_8;
	wire[1:0] w_n557_0;
	wire[1:0] w_n559_0;
	wire[2:0] w_n560_0;
	wire[2:0] w_n561_0;
	wire[1:0] w_n561_1;
	wire[1:0] w_n562_0;
	wire[1:0] w_n564_0;
	wire[2:0] w_n565_0;
	wire[2:0] w_n566_0;
	wire[2:0] w_n567_0;
	wire[1:0] w_n569_0;
	wire[1:0] w_n571_0;
	wire[2:0] w_n572_0;
	wire[2:0] w_n573_0;
	wire[2:0] w_n574_0;
	wire[2:0] w_n578_0;
	wire[1:0] w_n578_1;
	wire[2:0] w_n579_0;
	wire[1:0] w_n579_1;
	wire[1:0] w_n581_0;
	wire[2:0] w_n586_0;
	wire[1:0] w_n586_1;
	wire[1:0] w_n587_0;
	wire[2:0] w_n588_0;
	wire[1:0] w_n588_1;
	wire[2:0] w_n591_0;
	wire[1:0] w_n591_1;
	wire[2:0] w_n592_0;
	wire[2:0] w_n596_0;
	wire[1:0] w_n596_1;
	wire[2:0] w_n597_0;
	wire[2:0] w_n601_0;
	wire[1:0] w_n601_1;
	wire[2:0] w_n602_0;
	wire[1:0] w_n603_0;
	wire[2:0] w_n607_0;
	wire[1:0] w_n607_1;
	wire[2:0] w_n608_0;
	wire[2:0] w_n609_0;
	wire[2:0] w_n611_0;
	wire[2:0] w_n613_0;
	wire[2:0] w_n613_1;
	wire[2:0] w_n613_2;
	wire[2:0] w_n613_3;
	wire[2:0] w_n613_4;
	wire[2:0] w_n613_5;
	wire[2:0] w_n617_0;
	wire[1:0] w_n617_1;
	wire[2:0] w_n618_0;
	wire[2:0] w_n619_0;
	wire[2:0] w_n619_1;
	wire[2:0] w_n620_0;
	wire[1:0] w_n620_1;
	wire[1:0] w_n621_0;
	wire[1:0] w_n623_0;
	wire[2:0] w_n624_0;
	wire[1:0] w_n625_0;
	wire[2:0] w_n627_0;
	wire[1:0] w_n627_1;
	wire[2:0] w_n628_0;
	wire[1:0] w_n631_0;
	wire[1:0] w_n632_0;
	wire[2:0] w_n635_0;
	wire[1:0] w_n635_1;
	wire[2:0] w_n636_0;
	wire[2:0] w_n637_0;
	wire[1:0] w_n638_0;
	wire[2:0] w_n639_0;
	wire[1:0] w_n640_0;
	wire[2:0] w_n641_0;
	wire[2:0] w_n641_1;
	wire[2:0] w_n644_0;
	wire[2:0] w_n648_0;
	wire[1:0] w_n648_1;
	wire[1:0] w_n649_0;
	wire[1:0] w_n650_0;
	wire[2:0] w_n653_0;
	wire[2:0] w_n654_0;
	wire[2:0] w_n654_1;
	wire[2:0] w_n654_2;
	wire[2:0] w_n658_0;
	wire[1:0] w_n658_1;
	wire[1:0] w_n659_0;
	wire[2:0] w_n660_0;
	wire[1:0] w_n660_1;
	wire[1:0] w_n661_0;
	wire[1:0] w_n670_0;
	wire[1:0] w_n680_0;
	wire[2:0] w_n682_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n685_0;
	wire[1:0] w_n686_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n692_0;
	wire[2:0] w_n694_0;
	wire[2:0] w_n695_0;
	wire[2:0] w_n699_0;
	wire[1:0] w_n701_0;
	wire[2:0] w_n703_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n709_0;
	wire[1:0] w_n710_0;
	wire[1:0] w_n711_0;
	wire[2:0] w_n713_0;
	wire[2:0] w_n715_0;
	wire[1:0] w_n717_0;
	wire[1:0] w_n719_0;
	wire[1:0] w_n720_0;
	wire[1:0] w_n721_0;
	wire[1:0] w_n722_0;
	wire[2:0] w_n725_0;
	wire[1:0] w_n726_0;
	wire[1:0] w_n728_0;
	wire[2:0] w_n733_0;
	wire[2:0] w_n735_0;
	wire[2:0] w_n737_0;
	wire[1:0] w_n737_1;
	wire[1:0] w_n738_0;
	wire[2:0] w_n742_0;
	wire[1:0] w_n745_0;
	wire[2:0] w_n746_0;
	wire[1:0] w_n747_0;
	wire[2:0] w_n749_0;
	wire[2:0] w_n749_1;
	wire[2:0] w_n749_2;
	wire[2:0] w_n749_3;
	wire[2:0] w_n749_4;
	wire[2:0] w_n749_5;
	wire[2:0] w_n749_6;
	wire[2:0] w_n749_7;
	wire[2:0] w_n749_8;
	wire[2:0] w_n749_9;
	wire[2:0] w_n749_10;
	wire[2:0] w_n749_11;
	wire[2:0] w_n749_12;
	wire[1:0] w_n749_13;
	wire[2:0] w_n750_0;
	wire[2:0] w_n750_1;
	wire[2:0] w_n750_2;
	wire[2:0] w_n750_3;
	wire[2:0] w_n750_4;
	wire[2:0] w_n750_5;
	wire[2:0] w_n750_6;
	wire[2:0] w_n750_7;
	wire[2:0] w_n750_8;
	wire[2:0] w_n753_0;
	wire[1:0] w_n753_1;
	wire[1:0] w_n755_0;
	wire[2:0] w_n763_0;
	wire[1:0] w_n767_0;
	wire[1:0] w_n779_0;
	wire[2:0] w_n786_0;
	wire[2:0] w_n788_0;
	wire[2:0] w_n790_0;
	wire[2:0] w_n792_0;
	wire[2:0] w_n795_0;
	wire[1:0] w_n795_1;
	wire[2:0] w_n797_0;
	wire[2:0] w_n797_1;
	wire[2:0] w_n797_2;
	wire[2:0] w_n797_3;
	wire[2:0] w_n797_4;
	wire[2:0] w_n797_5;
	wire[2:0] w_n797_6;
	wire[2:0] w_n797_7;
	wire[2:0] w_n797_8;
	wire[1:0] w_n797_9;
	wire[2:0] w_n798_0;
	wire[1:0] w_n798_1;
	wire[2:0] w_n800_0;
	wire[2:0] w_n800_1;
	wire[2:0] w_n800_2;
	wire[2:0] w_n800_3;
	wire[1:0] w_n800_4;
	wire[2:0] w_n801_0;
	wire[1:0] w_n801_1;
	wire[2:0] w_n814_0;
	wire[2:0] w_n819_0;
	wire[1:0] w_n821_0;
	wire[1:0] w_n824_0;
	wire[1:0] w_n827_0;
	wire[1:0] w_n836_0;
	wire[1:0] w_n847_0;
	wire[2:0] w_n852_0;
	wire[2:0] w_n852_1;
	wire[2:0] w_n852_2;
	wire[2:0] w_n852_3;
	wire[2:0] w_n852_4;
	wire[2:0] w_n852_5;
	wire[2:0] w_n852_6;
	wire[2:0] w_n852_7;
	wire[2:0] w_n852_8;
	wire[1:0] w_n852_9;
	wire[2:0] w_n854_0;
	wire[2:0] w_n854_1;
	wire[2:0] w_n854_2;
	wire[2:0] w_n854_3;
	wire[1:0] w_n854_4;
	wire[2:0] w_n865_0;
	wire[1:0] w_n867_0;
	wire[1:0] w_n868_0;
	wire[1:0] w_n870_0;
	wire[1:0] w_n871_0;
	wire[1:0] w_n880_0;
	wire[1:0] w_n890_0;
	wire[1:0] w_n901_0;
	wire[2:0] w_n923_0;
	wire[1:0] w_n935_0;
	wire[2:0] w_n938_0;
	wire[2:0] w_n940_0;
	wire[1:0] w_n940_1;
	wire[1:0] w_n944_0;
	wire[1:0] w_n949_0;
	wire[1:0] w_n953_0;
	wire[2:0] w_n954_0;
	wire[1:0] w_n957_0;
	wire[1:0] w_n962_0;
	wire[1:0] w_n964_0;
	wire[1:0] w_n969_0;
	wire[2:0] w_n977_0;
	wire[1:0] w_n981_0;
	wire[1:0] w_n986_0;
	wire[1:0] w_n989_0;
	wire[2:0] w_n993_0;
	wire[2:0] w_n993_1;
	wire[2:0] w_n993_2;
	wire[2:0] w_n993_3;
	wire[2:0] w_n993_4;
	wire[2:0] w_n994_0;
	wire[2:0] w_n994_1;
	wire[2:0] w_n994_2;
	wire[2:0] w_n994_3;
	wire[1:0] w_n994_4;
	wire[2:0] w_n996_0;
	wire[2:0] w_n996_1;
	wire[2:0] w_n996_2;
	wire[2:0] w_n996_3;
	wire[1:0] w_n996_4;
	wire[2:0] w_n999_0;
	wire[2:0] w_n999_1;
	wire[2:0] w_n999_2;
	wire[2:0] w_n999_3;
	wire[2:0] w_n1007_0;
	wire[2:0] w_n1007_1;
	wire[2:0] w_n1007_2;
	wire[2:0] w_n1007_3;
	wire[2:0] w_n1008_0;
	wire[2:0] w_n1008_1;
	wire[2:0] w_n1008_2;
	wire[2:0] w_n1008_3;
	wire[2:0] w_n1008_4;
	wire[2:0] w_n1012_0;
	wire[2:0] w_n1012_1;
	wire[2:0] w_n1012_2;
	wire[2:0] w_n1012_3;
	wire[1:0] w_n1012_4;
	wire[2:0] w_n1014_0;
	wire[2:0] w_n1014_1;
	wire[2:0] w_n1014_2;
	wire[2:0] w_n1014_3;
	wire[1:0] w_n1014_4;
	wire[2:0] w_n1019_0;
	wire[1:0] w_n1019_1;
	wire[2:0] w_n1021_0;
	wire[1:0] w_n1021_1;
	wire[2:0] w_n1030_0;
	wire[1:0] w_n1030_1;
	wire[2:0] w_n1032_0;
	wire[1:0] w_n1032_1;
	wire[2:0] w_n1041_0;
	wire[1:0] w_n1041_1;
	wire[2:0] w_n1043_0;
	wire[1:0] w_n1043_1;
	wire[2:0] w_n1052_0;
	wire[1:0] w_n1052_1;
	wire[2:0] w_n1054_0;
	wire[1:0] w_n1054_1;
	wire[1:0] w_n1177_0;
	wire[1:0] w_n1179_0;
	wire[2:0] w_n1196_0;
	wire[2:0] w_n1196_1;
	wire[2:0] w_n1201_0;
	wire[2:0] w_n1205_0;
	wire[2:0] w_n1205_1;
	wire[2:0] w_n1213_0;
	wire[2:0] w_n1213_1;
	wire[2:0] w_n1236_0;
	wire[2:0] w_n1236_1;
	wire[2:0] w_n1251_0;
	wire[2:0] w_n1251_1;
	wire[2:0] w_n1279_0;
	wire[1:0] w_n1279_1;
	wire[2:0] w_n1297_0;
	wire[1:0] w_n1297_1;
	wire[2:0] w_n1299_0;
	wire[1:0] w_n1299_1;
	wire[2:0] w_n1410_0;
	wire[2:0] w_n1412_0;
	wire[1:0] w_n1416_0;
	wire[1:0] w_n1422_0;
	wire[1:0] w_n1425_0;
	wire[1:0] w_n1428_0;
	wire[1:0] w_n1429_0;
	wire[1:0] w_n1451_0;
	wire[1:0] w_n1503_0;
	wire[1:0] w_n1504_0;
	wire[1:0] w_n1592_0;
	wire[1:0] w_n1593_0;
	wire[1:0] w_n1596_0;
	wire[1:0] w_n1599_0;
	wire[1:0] w_n1603_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1609_0;
	wire[2:0] w_n1611_0;
	wire[1:0] w_n1613_0;
	wire[1:0] w_n1615_0;
	wire[1:0] w_n1618_0;
	wire[1:0] w_n1633_0;
	wire[1:0] w_n1637_0;
	wire[1:0] w_n1643_0;
	wire[1:0] w_n1652_0;
	wire[1:0] w_n1665_0;
	wire[2:0] w_n1674_0;
	wire[1:0] w_n1675_0;
	wire[2:0] w_n1679_0;
	wire[1:0] w_n1680_0;
	wire[1:0] w_n1694_0;
	wire[1:0] w_n1695_0;
	wire[1:0] w_n1698_0;
	wire w_dff_B_1XDqtN614_1;
	wire w_dff_B_NWXNKUrM1_0;
	wire w_dff_B_DGe8f2Ly5_1;
	wire w_dff_B_02uGgqTc3_1;
	wire w_dff_B_8mCnqYH29_2;
	wire w_dff_B_WU1X1XVA1_1;
	wire w_dff_B_cWl4mArx2_1;
	wire w_dff_B_ymTIAQl32_0;
	wire w_dff_B_evs6UKxu5_1;
	wire w_dff_B_4hxtTxcj6_0;
	wire w_dff_A_aTDcNNYc3_0;
	wire w_dff_A_6TXUEXf09_0;
	wire w_dff_A_UMdNmIRg8_0;
	wire w_dff_A_NY7cL5aH0_0;
	wire w_dff_A_CTZAlmyf1_1;
	wire w_dff_A_VNgfi1wZ6_1;
	wire w_dff_A_5VzWEKJm9_1;
	wire w_dff_A_nCk6XHLC6_1;
	wire w_dff_B_uVFbPRHM4_1;
	wire w_dff_B_ct9crCYT1_0;
	wire w_dff_B_t7LjX50Y3_1;
	wire w_dff_B_YVG9Lfyh4_1;
	wire w_dff_A_QYFEgyJ75_1;
	wire w_dff_A_rtIH0M167_1;
	wire w_dff_A_3YClfHk96_1;
	wire w_dff_A_Z7jBtOZN9_1;
	wire w_dff_A_E051C3Hs2_2;
	wire w_dff_A_P9uuXgGt3_2;
	wire w_dff_A_jqXwJ04v1_2;
	wire w_dff_A_NDNz4G301_2;
	wire w_dff_B_QLc7tfjg4_2;
	wire w_dff_B_yxUZZkK22_2;
	wire w_dff_B_ejixAcWz8_2;
	wire w_dff_B_LnBv0cEL0_2;
	wire w_dff_B_ZpYFQVyI0_2;
	wire w_dff_B_dL1fOSbo0_2;
	wire w_dff_B_42FdxOi56_1;
	wire w_dff_B_nYAXIFgQ6_1;
	wire w_dff_A_wuoPVNGL9_0;
	wire w_dff_A_1WsWmMIa4_0;
	wire w_dff_A_Q3QhfmJ97_0;
	wire w_dff_A_N2EbYwlV9_0;
	wire w_dff_A_I23wfQs24_0;
	wire w_dff_B_SrbdkDKe1_0;
	wire w_dff_B_CLpfSep24_0;
	wire w_dff_B_VLthB9qI7_0;
	wire w_dff_B_pXxDp6Gp4_0;
	wire w_dff_B_W0hYXjTc2_0;
	wire w_dff_B_2gpE8J2N2_0;
	wire w_dff_B_vGuJ81Mt1_0;
	wire w_dff_B_qGsbcCoP7_0;
	wire w_dff_B_I3EXTdrl5_0;
	wire w_dff_B_sdoMaWUL3_0;
	wire w_dff_B_h0oYGuxO9_0;
	wire w_dff_B_PsD8Npqn0_0;
	wire w_dff_B_FCir2w6a8_0;
	wire w_dff_B_Y5xQJbdQ2_0;
	wire w_dff_B_UoJE27xX2_0;
	wire w_dff_B_r7vsXoro3_0;
	wire w_dff_B_LDQicVIw5_0;
	wire w_dff_B_zZKmTWFN9_0;
	wire w_dff_B_wHakUf6M9_0;
	wire w_dff_B_hLiWu55m5_0;
	wire w_dff_B_VjAzt5NF2_0;
	wire w_dff_B_2QD7IzGH6_0;
	wire w_dff_B_e9C2TA1l0_0;
	wire w_dff_B_pCqoakHu4_1;
	wire w_dff_B_TFXHJJCi8_1;
	wire w_dff_B_1f6Bj5Ek6_1;
	wire w_dff_B_xuXpjySI2_1;
	wire w_dff_B_thoFfn6c7_1;
	wire w_dff_B_rNexfRzB6_1;
	wire w_dff_B_7yMBzruG2_1;
	wire w_dff_B_wbZMDG4q2_1;
	wire w_dff_B_aBxZBdJR1_1;
	wire w_dff_B_pwN17cui4_1;
	wire w_dff_B_iITFd7oW1_1;
	wire w_dff_B_REj9hCEs1_1;
	wire w_dff_B_2NVMryv08_1;
	wire w_dff_B_1J9G3Uuu6_1;
	wire w_dff_B_8tTiHC1z2_1;
	wire w_dff_B_2mbvwedk1_1;
	wire w_dff_B_8D4Cehdn5_1;
	wire w_dff_B_MJIvSDTw3_1;
	wire w_dff_B_qQYNLmVd5_1;
	wire w_dff_B_LriefBrK7_1;
	wire w_dff_B_OAH3sFTR3_1;
	wire w_dff_B_PwyMtHtu2_1;
	wire w_dff_B_Kvi4Oh500_1;
	wire w_dff_B_L3pEp55h8_1;
	wire w_dff_B_BvbV19yi7_1;
	wire w_dff_B_zOxoHVXV3_1;
	wire w_dff_B_PqIQVwuk4_1;
	wire w_dff_B_siH4tvwf9_1;
	wire w_dff_B_uHiqWlh60_1;
	wire w_dff_B_rMnhefMo1_0;
	wire w_dff_B_DIwzV3yi0_0;
	wire w_dff_B_mzplZVB74_0;
	wire w_dff_B_P3URP6Jn0_0;
	wire w_dff_B_WejOFSqx6_0;
	wire w_dff_B_Tah9espN4_0;
	wire w_dff_B_uT0vOAA74_0;
	wire w_dff_B_lrFqCve71_0;
	wire w_dff_B_04iIw3AU5_0;
	wire w_dff_B_VGzPUyC36_0;
	wire w_dff_B_bYh6fuTv8_0;
	wire w_dff_B_RZOzaCt11_1;
	wire w_dff_B_LVbo2nxR3_1;
	wire w_dff_B_YZS4p8r72_1;
	wire w_dff_B_OZuyXFgh3_0;
	wire w_dff_B_TZeEagoR7_0;
	wire w_dff_B_RNGNwtdz4_0;
	wire w_dff_B_NrS56NpP3_0;
	wire w_dff_B_UfNREkOv9_0;
	wire w_dff_B_3M7YxRyR4_0;
	wire w_dff_B_2Jfz7Zt00_0;
	wire w_dff_B_4UOLOE5W6_0;
	wire w_dff_B_q2lMszzI4_0;
	wire w_dff_B_TotN7z2m8_0;
	wire w_dff_B_hqeALvmp3_0;
	wire w_dff_B_IFuUqoQf6_0;
	wire w_dff_B_tXLsthCU3_0;
	wire w_dff_B_WQB4AGs89_0;
	wire w_dff_B_5mZAup1X2_0;
	wire w_dff_B_baGPJQFF2_0;
	wire w_dff_B_TSxWOlHm2_1;
	wire w_dff_A_y0fqPlcu6_0;
	wire w_dff_A_sbO4wRnm7_0;
	wire w_dff_A_7fY6GrcM0_0;
	wire w_dff_A_XvKYeoGL6_0;
	wire w_dff_A_lfP0Vq4G8_0;
	wire w_dff_A_XGsL5Nx21_0;
	wire w_dff_A_i5zeMe8m5_0;
	wire w_dff_B_UkuSXVZ87_0;
	wire w_dff_B_nvvzkRGz5_0;
	wire w_dff_B_mOfkBuob3_0;
	wire w_dff_B_fVx42glE8_0;
	wire w_dff_B_pwUFTuat9_0;
	wire w_dff_B_A7VEBaJA1_0;
	wire w_dff_B_hpv8jVYK1_0;
	wire w_dff_B_xIKTjiuK4_0;
	wire w_dff_B_I5o47Je97_0;
	wire w_dff_B_9apthTB20_0;
	wire w_dff_B_GC6dFs5Q2_0;
	wire w_dff_B_ZZA6qjNH5_0;
	wire w_dff_B_ljwCGGod1_0;
	wire w_dff_B_jRLIr8sL6_0;
	wire w_dff_B_vsXxz3Ng1_0;
	wire w_dff_B_PWB45Tqz8_1;
	wire w_dff_B_Y8Qdl6VR9_1;
	wire w_dff_B_ZPONdbT25_0;
	wire w_dff_B_48vW2mRd5_0;
	wire w_dff_B_6R72KguM9_0;
	wire w_dff_B_FR9HuwVd8_0;
	wire w_dff_B_V6Eikr194_0;
	wire w_dff_B_7rlcIVMq2_0;
	wire w_dff_B_FglxMB1B0_0;
	wire w_dff_B_y7Lshb6E1_0;
	wire w_dff_B_0aXLOIpJ1_0;
	wire w_dff_B_1WBtCBOx5_0;
	wire w_dff_B_OGsxnyeT8_0;
	wire w_dff_B_gvGwydth1_0;
	wire w_dff_B_D13BJunD9_0;
	wire w_dff_B_8s8YOFXV9_1;
	wire w_dff_B_PgOL7VEo2_0;
	wire w_dff_B_E3OnIGUU0_0;
	wire w_dff_B_eiIB6mQO3_0;
	wire w_dff_B_UlwlA0fX1_0;
	wire w_dff_B_B2REas4L4_0;
	wire w_dff_B_HlK88dhT0_0;
	wire w_dff_B_kpM6Du0e2_0;
	wire w_dff_B_ZQYkGd7d7_0;
	wire w_dff_B_oH8U7Bho9_0;
	wire w_dff_B_q6YpXPcs4_0;
	wire w_dff_B_DlVTVJYc3_0;
	wire w_dff_B_y0Ay3AzT5_0;
	wire w_dff_B_3Jkd2jMy3_0;
	wire w_dff_B_TocnJ47N6_0;
	wire w_dff_B_kyKZDjEP3_1;
	wire w_dff_B_8WwbDecL4_1;
	wire w_dff_B_66V6EbF32_1;
	wire w_dff_A_OzL5O6s65_0;
	wire w_dff_A_mSNHzLrI6_2;
	wire w_dff_A_AHqMAjRY7_2;
	wire w_dff_B_P7G6dOCY0_1;
	wire w_dff_B_iDUut8Ig3_1;
	wire w_dff_B_HlHw4r4Z8_1;
	wire w_dff_B_mAETDW4n0_1;
	wire w_dff_B_Ss7mZ6oL8_1;
	wire w_dff_B_6SRlSjqt5_1;
	wire w_dff_B_KHObKrTC0_1;
	wire w_dff_B_TCJLlppF8_1;
	wire w_dff_B_aav5VX5B9_1;
	wire w_dff_B_avB97Oq41_1;
	wire w_dff_B_shrUwFB68_1;
	wire w_dff_B_nMke7Iym7_1;
	wire w_dff_B_9cgTWemn0_1;
	wire w_dff_B_z0ktVAng5_1;
	wire w_dff_B_0rAy1vbr2_1;
	wire w_dff_A_p1TMc0sP2_0;
	wire w_dff_A_o7YhbvWz6_0;
	wire w_dff_A_kC6bmOQa3_0;
	wire w_dff_A_3TdTeVSQ9_0;
	wire w_dff_A_gt2pzEm99_0;
	wire w_dff_A_Ph7CHpmE9_0;
	wire w_dff_A_fjg75LeW8_0;
	wire w_dff_A_EjKLw5jY3_0;
	wire w_dff_B_MLk6KA3G8_1;
	wire w_dff_B_ZZuCoweL7_1;
	wire w_dff_B_Qscbnwhp2_1;
	wire w_dff_B_plH4Uu8A8_1;
	wire w_dff_B_6qR45CO72_1;
	wire w_dff_B_V0UDLpRB9_1;
	wire w_dff_B_ZaiO6gz98_1;
	wire w_dff_B_JZMAV0XQ6_1;
	wire w_dff_B_WfXQttZa4_1;
	wire w_dff_B_Y2CBN6gi9_1;
	wire w_dff_B_lAYgpfSH5_1;
	wire w_dff_B_dtzgPbxY0_1;
	wire w_dff_B_3IJSS4FF6_1;
	wire w_dff_B_WO2QjJZx1_1;
	wire w_dff_B_WtjqIDdJ3_0;
	wire w_dff_B_Wk9Y8kd14_1;
	wire w_dff_B_wptY5y6H0_1;
	wire w_dff_B_I0MucakO7_1;
	wire w_dff_B_naT1y9Xs0_1;
	wire w_dff_B_RzAhAgK08_1;
	wire w_dff_B_eyWrL4c61_1;
	wire w_dff_B_eknu4SOh1_1;
	wire w_dff_B_VPfWt4Ou7_1;
	wire w_dff_B_9O0tHRuR8_1;
	wire w_dff_B_2PdW1mX86_1;
	wire w_dff_B_pxtOYEPZ7_1;
	wire w_dff_B_vdVDT8fO7_1;
	wire w_dff_B_nzWmdS5U0_0;
	wire w_dff_B_nh0Zbccj3_0;
	wire w_dff_B_zlEUIu1y4_0;
	wire w_dff_B_FXJ24YZv4_0;
	wire w_dff_B_JshCWRao6_0;
	wire w_dff_B_RooTn53j1_0;
	wire w_dff_B_7hba4mDo1_0;
	wire w_dff_B_Tdyjeyzi3_0;
	wire w_dff_B_cpcPuiuM3_0;
	wire w_dff_B_jnCmFogt4_0;
	wire w_dff_B_a20HcxR97_0;
	wire w_dff_B_xm2v5N5I8_0;
	wire w_dff_B_zX9qkJnc3_0;
	wire w_dff_B_ePcFd7uz4_0;
	wire w_dff_B_6TYDbxhT4_1;
	wire w_dff_B_9HSbRjVc2_1;
	wire w_dff_B_rdYUYjWb3_1;
	wire w_dff_A_yuVUJRug6_2;
	wire w_dff_A_P2s8uA8u4_2;
	wire w_dff_B_dlYx2j1Q4_0;
	wire w_dff_B_sNuZ5cFE9_0;
	wire w_dff_B_HoCY4SA79_0;
	wire w_dff_B_RlwrtYV62_0;
	wire w_dff_B_5Yy2qkgE2_0;
	wire w_dff_B_fsvYl8F98_0;
	wire w_dff_B_U8RIMQyq1_0;
	wire w_dff_B_S68Ih2m87_0;
	wire w_dff_B_eBnMiTXi9_0;
	wire w_dff_B_rZQAnHAz7_0;
	wire w_dff_B_xVAPP0WQ9_0;
	wire w_dff_B_obB8VCKb3_0;
	wire w_dff_B_OQ2cJw1E0_0;
	wire w_dff_B_yyBZyRr94_0;
	wire w_dff_B_Hci9Zji85_0;
	wire w_dff_B_b3hbbYEy1_1;
	wire w_dff_B_XMnLS7YG8_0;
	wire w_dff_B_UO0V1KFA6_0;
	wire w_dff_B_QIpU5tY40_0;
	wire w_dff_B_At0f5HrN7_0;
	wire w_dff_B_0oCccyPS5_0;
	wire w_dff_B_EPKsemQA7_0;
	wire w_dff_B_jHDUVhod8_0;
	wire w_dff_B_CkjCoHxC9_0;
	wire w_dff_B_3Y0GYcFm4_0;
	wire w_dff_B_UdI0GnYB9_0;
	wire w_dff_B_rmEus8dW7_0;
	wire w_dff_B_Suvoinvj4_0;
	wire w_dff_B_YpGI6jln1_0;
	wire w_dff_A_rEkd99D39_0;
	wire w_dff_A_HGhebhM94_0;
	wire w_dff_A_MwSGsGmt7_0;
	wire w_dff_A_kcapujoy5_1;
	wire w_dff_A_zIehUUja3_1;
	wire w_dff_A_1dzGRIFT0_1;
	wire w_dff_A_X5yVBLaX7_1;
	wire w_dff_A_ALTtceVh9_1;
	wire w_dff_A_xD53gBXo1_1;
	wire w_dff_A_ZHlsjuj38_1;
	wire w_dff_A_kkwRc1Fa1_0;
	wire w_dff_A_9JDF0wyn4_0;
	wire w_dff_A_LJznGtt23_0;
	wire w_dff_A_LFhCZYSH3_0;
	wire w_dff_A_ULX69nvB6_0;
	wire w_dff_A_UPrmTDyU9_1;
	wire w_dff_A_89LOEPJJ0_1;
	wire w_dff_A_l6gYRpAo7_1;
	wire w_dff_A_7cuavIbH0_1;
	wire w_dff_A_fG87pw2R0_1;
	wire w_dff_A_2lyjNTof5_1;
	wire w_dff_A_JdFhaelb0_1;
	wire w_dff_B_2fsWrDcZ2_0;
	wire w_dff_B_dHBPR1nd2_0;
	wire w_dff_B_7jUGA8E67_0;
	wire w_dff_B_9elJXMvt8_0;
	wire w_dff_B_DsHfFmhI8_0;
	wire w_dff_B_WSXC1QKs9_0;
	wire w_dff_B_aps5827G2_0;
	wire w_dff_B_4SatGGgD4_0;
	wire w_dff_B_Q1Aglej13_0;
	wire w_dff_B_brgsmrrX9_0;
	wire w_dff_B_Bk8tETIl3_0;
	wire w_dff_B_Y7YB1tXd4_0;
	wire w_dff_B_PvQKJ1lH9_1;
	wire w_dff_A_LHTlblFS7_2;
	wire w_dff_A_QgzC8xx93_2;
	wire w_dff_A_CbUuo9Gv3_2;
	wire w_dff_B_Js8RLDsD4_0;
	wire w_dff_B_Drjgelto1_0;
	wire w_dff_B_CMJUo9XR2_0;
	wire w_dff_B_0pHUcuBP5_0;
	wire w_dff_B_GDpbnEjJ8_0;
	wire w_dff_B_Zhve6e8w0_0;
	wire w_dff_B_KnwXlI7I8_0;
	wire w_dff_B_uymMJo6F5_0;
	wire w_dff_B_FYTBqWQe6_0;
	wire w_dff_B_3fMqkkZ20_0;
	wire w_dff_B_C3lzjKps7_0;
	wire w_dff_B_c6InWFUx7_0;
	wire w_dff_B_Sq6Y1wZs9_0;
	wire w_dff_A_kM4Ok63H1_0;
	wire w_dff_A_F2Q6BTQG0_0;
	wire w_dff_A_fhl7roYl2_1;
	wire w_dff_B_ybdAiMZK7_1;
	wire w_dff_B_DwjsQlGf0_1;
	wire w_dff_B_cAQLgNRl4_1;
	wire w_dff_B_HsSKzZDF1_1;
	wire w_dff_B_CeNcjF2b4_1;
	wire w_dff_B_ACwUTcPA8_1;
	wire w_dff_B_FToaxKG98_1;
	wire w_dff_B_Z4wexT3S3_1;
	wire w_dff_B_8iD17oYr0_1;
	wire w_dff_B_sBPiagre0_1;
	wire w_dff_B_m7meNjhp8_1;
	wire w_dff_B_2FbThkxa8_1;
	wire w_dff_B_lwChKyxl1_1;
	wire w_dff_B_37WBQKT70_1;
	wire w_dff_B_8tWgp4Jh7_1;
	wire w_dff_B_Fsu4cCZy0_1;
	wire w_dff_B_ILpdYLST9_1;
	wire w_dff_B_1Okr1deu8_1;
	wire w_dff_B_z0fjnVN23_1;
	wire w_dff_B_pYOdEXAk3_1;
	wire w_dff_B_v3MvVb3h3_1;
	wire w_dff_B_d8Kx8qZ75_1;
	wire w_dff_B_LvCcI1oo8_1;
	wire w_dff_B_Wi9RNXN35_1;
	wire w_dff_B_fl36zeOT7_1;
	wire w_dff_B_5thsbeGK3_1;
	wire w_dff_B_qDKTk91n6_1;
	wire w_dff_B_QcRAS6s42_1;
	wire w_dff_B_yLHma9SI5_1;
	wire w_dff_B_GkyL48KR9_1;
	wire w_dff_B_A7uZoiyP5_1;
	wire w_dff_B_FnpRua1h8_1;
	wire w_dff_B_6H7jaLad3_1;
	wire w_dff_B_DCt5fdP63_1;
	wire w_dff_B_TUFBbBAt5_1;
	wire w_dff_B_zXGAUlEA6_1;
	wire w_dff_B_MbKSQnhm4_1;
	wire w_dff_B_KVmAjwlj9_1;
	wire w_dff_B_XWUq6Fah9_1;
	wire w_dff_B_jP5Ik2EJ0_1;
	wire w_dff_B_tMHefNiG9_1;
	wire w_dff_B_It6OdICZ9_1;
	wire w_dff_B_AjcHYoEb5_1;
	wire w_dff_B_eluNYSm06_1;
	wire w_dff_B_nhvyUovY4_0;
	wire w_dff_B_wOyIj7qj3_0;
	wire w_dff_B_rQqkwRhB6_0;
	wire w_dff_B_65aqk9292_0;
	wire w_dff_B_xjmPbzyC7_0;
	wire w_dff_B_g4VSIKkr6_0;
	wire w_dff_B_P0QGvQNP1_1;
	wire w_dff_B_KtEtKJji2_1;
	wire w_dff_B_BJbGIzEY5_1;
	wire w_dff_B_xxdvb4ew8_1;
	wire w_dff_B_JYWRbbI97_1;
	wire w_dff_B_GYlf9tmp0_0;
	wire w_dff_B_QaQDSJFo4_0;
	wire w_dff_B_T0qrOHgi4_0;
	wire w_dff_B_IlgMwBIO6_0;
	wire w_dff_B_YAgN0rkF8_0;
	wire w_dff_B_L4m7v8lK9_0;
	wire w_dff_B_iOqssW0V2_0;
	wire w_dff_B_D5ri3bxJ3_0;
	wire w_dff_B_pXI7YmXC2_0;
	wire w_dff_B_wzyJFi5n6_0;
	wire w_dff_B_X3rX3h1N3_0;
	wire w_dff_B_WBQU4sIr8_0;
	wire w_dff_B_i1xdznr45_0;
	wire w_dff_A_PIcgelcc1_0;
	wire w_dff_A_NwuXZuxK5_1;
	wire w_dff_A_vHywm2w90_1;
	wire w_dff_A_iE53cuUi2_1;
	wire w_dff_A_KRGFQMvu0_1;
	wire w_dff_A_Q5q0762m9_1;
	wire w_dff_A_9gFfPl351_1;
	wire w_dff_B_Rn4WCP9Z0_1;
	wire w_dff_B_geuXO1e88_1;
	wire w_dff_B_OtJa7mWN0_1;
	wire w_dff_B_6JElo9hD4_1;
	wire w_dff_B_6eKDnRiu8_1;
	wire w_dff_B_LZtyHhp22_1;
	wire w_dff_B_b0KXPMBY7_1;
	wire w_dff_B_1h6ymRVb5_1;
	wire w_dff_B_Aj3s74Qr4_0;
	wire w_dff_B_4CZvdFqP8_0;
	wire w_dff_B_zV1xcR2g4_0;
	wire w_dff_B_gT4N4AbX2_0;
	wire w_dff_B_EI8qdsfc3_0;
	wire w_dff_B_88nphrFP2_0;
	wire w_dff_B_8s4KVCS63_0;
	wire w_dff_B_mqpqi7DM5_0;
	wire w_dff_A_394idVPZ4_1;
	wire w_dff_A_kjJ1EEFO9_1;
	wire w_dff_A_JjLejf5U9_1;
	wire w_dff_A_0JDJpoad9_1;
	wire w_dff_A_r8xWbjbI8_2;
	wire w_dff_A_My38uOGv8_0;
	wire w_dff_A_dH68NgwT8_0;
	wire w_dff_A_FA9GbpNf2_1;
	wire w_dff_A_Exb9jyy65_1;
	wire w_dff_B_lb1qM44B4_0;
	wire w_dff_B_Ryn9RK0i8_0;
	wire w_dff_B_UJqb6P6u9_0;
	wire w_dff_B_WmlnOgTz8_0;
	wire w_dff_B_8wM9d6928_0;
	wire w_dff_B_VHvu3BTi2_0;
	wire w_dff_B_gVy0gIJY5_0;
	wire w_dff_B_DTqzfii80_0;
	wire w_dff_B_bitBGjAr2_0;
	wire w_dff_B_EvUtjhT30_0;
	wire w_dff_B_BFFTF91n5_0;
	wire w_dff_B_6dxuLh870_0;
	wire w_dff_B_3qN4cbYf0_1;
	wire w_dff_B_XBy4Vuwp3_1;
	wire w_dff_B_QnOTtXCy1_1;
	wire w_dff_B_ApErmMJk6_1;
	wire w_dff_B_nEVJ6oVV3_1;
	wire w_dff_B_QLOQPG8i0_1;
	wire w_dff_B_9pOpdXtw3_1;
	wire w_dff_B_ZeJDghyp9_1;
	wire w_dff_B_tgDCCe2M3_1;
	wire w_dff_B_beOOIN0R0_1;
	wire w_dff_B_s7MYspbX0_1;
	wire w_dff_B_5z9KsX4z9_1;
	wire w_dff_A_JcH5yEVp0_0;
	wire w_dff_A_YKVLwzCi9_0;
	wire w_dff_A_Qc9LS6Lr6_0;
	wire w_dff_A_u255Ju3h1_0;
	wire w_dff_A_QOxkxB1I3_0;
	wire w_dff_B_DaxcvxvW4_0;
	wire w_dff_B_QEMgVGea6_0;
	wire w_dff_B_loUNumSK5_0;
	wire w_dff_B_ZzPWaRZK7_0;
	wire w_dff_B_G3mwbcmp7_0;
	wire w_dff_B_Q5f7ILYP8_0;
	wire w_dff_B_HQhAEU7Z2_0;
	wire w_dff_B_Ux9JRKrS5_0;
	wire w_dff_B_WsIEIQma6_0;
	wire w_dff_B_OdClI2C52_0;
	wire w_dff_B_abBQ0BRH3_0;
	wire w_dff_B_wX6OIxDw5_0;
	wire w_dff_B_1oUwOJya1_0;
	wire w_dff_A_ANLfMAZe9_0;
	wire w_dff_A_PHmYnQ426_0;
	wire w_dff_A_CNn93fsX2_1;
	wire w_dff_B_MPOcCkTp6_1;
	wire w_dff_B_2fYVIv2c2_1;
	wire w_dff_B_cDVfxSgn1_1;
	wire w_dff_B_8rzkGeZV9_1;
	wire w_dff_B_tQ91bYHC3_1;
	wire w_dff_B_cG1SKwuA2_1;
	wire w_dff_B_QKEJEcGo1_1;
	wire w_dff_B_FUjWWtXH5_1;
	wire w_dff_B_b7l7TUX85_1;
	wire w_dff_B_hwfvK0fe6_0;
	wire w_dff_B_w0DLYHA09_0;
	wire w_dff_B_1vKv8XKJ5_0;
	wire w_dff_B_SVYZF8wu0_0;
	wire w_dff_B_hN8odqwb6_0;
	wire w_dff_B_2YSxb2fz8_0;
	wire w_dff_A_JzCI1fDH0_0;
	wire w_dff_A_1MQZQAK70_0;
	wire w_dff_A_G6xBS8gp1_0;
	wire w_dff_A_LjcwLS5f1_0;
	wire w_dff_A_qib1nwvv2_0;
	wire w_dff_A_0VV33D722_0;
	wire w_dff_A_bKVOydk43_0;
	wire w_dff_B_v1bO5mI78_1;
	wire w_dff_B_9J5Yro5B3_1;
	wire w_dff_B_ieXzWPEE4_1;
	wire w_dff_B_wzNgKGVX6_1;
	wire w_dff_B_ne0AMC961_1;
	wire w_dff_B_4pA0ScO27_1;
	wire w_dff_B_aFAcwiUP0_1;
	wire w_dff_B_LCvqKDej3_1;
	wire w_dff_B_Zx0NJew23_1;
	wire w_dff_B_SzOYvOBJ6_1;
	wire w_dff_B_qip4DymN3_1;
	wire w_dff_B_8DhUfWxj1_1;
	wire w_dff_B_C5ATztjV6_1;
	wire w_dff_B_7xJhnG052_1;
	wire w_dff_B_ZPgOoydR5_1;
	wire w_dff_B_V7or1dHo8_1;
	wire w_dff_B_DMam5gA08_1;
	wire w_dff_B_1JZQHkVQ8_1;
	wire w_dff_B_m9XErvMi0_1;
	wire w_dff_B_MMnb1Wq13_1;
	wire w_dff_B_WTKqezxX2_1;
	wire w_dff_B_KEnsGmEz5_1;
	wire w_dff_B_qWpozdUN2_1;
	wire w_dff_B_emT5n7H64_1;
	wire w_dff_B_CFBEcHnW3_1;
	wire w_dff_B_uZlHwleW0_1;
	wire w_dff_B_cN5UFef44_1;
	wire w_dff_B_3gDUGkFP6_1;
	wire w_dff_B_GeuIZe7S9_0;
	wire w_dff_B_SKf02YKw3_0;
	wire w_dff_B_gHwkZVsd2_0;
	wire w_dff_B_EBkLG0Sg0_0;
	wire w_dff_B_w1UVBfmU1_0;
	wire w_dff_B_xnvLp0aB6_0;
	wire w_dff_B_b2vb30T19_0;
	wire w_dff_B_KO2DtA1o8_0;
	wire w_dff_B_rzXwiNao3_0;
	wire w_dff_B_aimPF6Yl5_0;
	wire w_dff_B_fs01Md6z6_0;
	wire w_dff_B_BzKjiF2z6_0;
	wire w_dff_B_tCHeFHea9_0;
	wire w_dff_B_45hcvCJ00_0;
	wire w_dff_B_7p2bQJV08_0;
	wire w_dff_B_FSaM279M7_0;
	wire w_dff_B_5ZDP9ftx9_1;
	wire w_dff_B_0fADwkXw9_1;
	wire w_dff_B_g6dH3Znt0_1;
	wire w_dff_B_lSSq5HWT9_1;
	wire w_dff_B_4GYBegJO0_1;
	wire w_dff_B_FuCfEokb2_1;
	wire w_dff_B_MOZGd3nc5_1;
	wire w_dff_B_KqV8IN1E0_1;
	wire w_dff_B_c9rVHgUN5_1;
	wire w_dff_A_xbbYYgWi3_0;
	wire w_dff_A_rsMdykz66_0;
	wire w_dff_A_SfEJBOaA0_0;
	wire w_dff_A_Q15o28yw6_0;
	wire w_dff_A_TGo1IMHy8_0;
	wire w_dff_A_4UL1BwAG7_0;
	wire w_dff_A_iu4QtZnr1_0;
	wire w_dff_A_pPSMOaFR4_0;
	wire w_dff_A_GK6LHLhs1_0;
	wire w_dff_A_p0MWBDBZ0_0;
	wire w_dff_A_jcFJtrsX8_0;
	wire w_dff_B_FT0M63c13_2;
	wire w_dff_B_LmrubnDT9_2;
	wire w_dff_B_XrQQAS405_2;
	wire w_dff_B_MH6DOu3F7_2;
	wire w_dff_B_xmNcrysp8_2;
	wire w_dff_A_c0gJlOqo4_0;
	wire w_dff_A_PnqvxPzc0_0;
	wire w_dff_A_7B7hsHaq2_0;
	wire w_dff_A_VBhZXm0p8_0;
	wire w_dff_A_miGwPmJY7_0;
	wire w_dff_A_2KYoFuJn0_0;
	wire w_dff_A_5wGTqp6I1_0;
	wire w_dff_A_dmkHZ2qv4_0;
	wire w_dff_A_oiBMTlRc5_0;
	wire w_dff_A_jpdcUoa39_0;
	wire w_dff_A_cinRNd2W2_0;
	wire w_dff_B_hCGCbvbn5_1;
	wire w_dff_B_HdAI6Y7T4_1;
	wire w_dff_B_2YvGSUPm0_1;
	wire w_dff_B_XYwVKQL19_1;
	wire w_dff_B_DKZt5hg95_1;
	wire w_dff_B_5F4cHltd1_0;
	wire w_dff_B_k4bFRORr8_0;
	wire w_dff_B_HLQ2XLlh4_0;
	wire w_dff_B_uXwQUzK48_0;
	wire w_dff_B_BzKGYPfc6_0;
	wire w_dff_A_L8qNNPTz3_0;
	wire w_dff_A_XYykHfUK1_0;
	wire w_dff_B_GLcQe6Os9_1;
	wire w_dff_B_IjWP77AJ0_1;
	wire w_dff_B_YwVVYjAq7_1;
	wire w_dff_B_1lWxf8dv3_1;
	wire w_dff_B_rZrAkUxI5_1;
	wire w_dff_B_3tDQzPvF4_1;
	wire w_dff_B_n66KbUP66_1;
	wire w_dff_B_NkSbuJrO0_1;
	wire w_dff_B_UVobcjTu0_1;
	wire w_dff_B_fPO83u4t8_1;
	wire w_dff_B_QbdKbOSC0_1;
	wire w_dff_B_gVUlk6Jo7_1;
	wire w_dff_B_0lZz5DDD5_1;
	wire w_dff_B_L30WRLTa1_1;
	wire w_dff_B_A94QpvrG7_1;
	wire w_dff_B_N4D3wLzj6_1;
	wire w_dff_B_7UY5i46H8_1;
	wire w_dff_B_fMhhPfwW0_1;
	wire w_dff_B_IlR4EslL7_1;
	wire w_dff_B_DrAd6EK05_1;
	wire w_dff_B_9knjpEj62_1;
	wire w_dff_B_Qz8uHCUV4_0;
	wire w_dff_B_QDvttSih6_0;
	wire w_dff_B_1wbw8wJY6_0;
	wire w_dff_B_AfiNB8fZ2_0;
	wire w_dff_B_MG0o2Qo24_0;
	wire w_dff_B_IWeYiSDd6_0;
	wire w_dff_B_5qv22RKN8_0;
	wire w_dff_B_GwwHDRTv8_0;
	wire w_dff_B_1YIloZ8U6_0;
	wire w_dff_B_NZifnjeV3_0;
	wire w_dff_B_vYBVypmd4_0;
	wire w_dff_B_KjRmi9ya0_0;
	wire w_dff_B_ccO3gIBX2_0;
	wire w_dff_B_xzfbcL2i0_0;
	wire w_dff_B_G05FjTiQ9_0;
	wire w_dff_B_7KI8fp1b4_0;
	wire w_dff_B_TfPXlL9x9_0;
	wire w_dff_B_38VjsrQn8_0;
	wire w_dff_B_czTqUtTy6_0;
	wire w_dff_B_TcphjBEB3_0;
	wire w_dff_B_uPb3CPjh2_0;
	wire w_dff_B_u4rw8Rgz0_1;
	wire w_dff_B_Ra935SOO5_1;
	wire w_dff_B_cEyVO6YC9_0;
	wire w_dff_B_xpsMYQWM6_0;
	wire w_dff_B_JuhiCCYr2_0;
	wire w_dff_B_qFhmG7bL7_0;
	wire w_dff_B_QzSkQ6Ak8_0;
	wire w_dff_B_fKiclD4E7_0;
	wire w_dff_B_62nVizES5_0;
	wire w_dff_B_BqAnvREk8_0;
	wire w_dff_B_ks4pwvVr8_0;
	wire w_dff_B_zqX8sWj22_0;
	wire w_dff_B_QEUynro25_0;
	wire w_dff_B_VucP6jzv4_0;
	wire w_dff_B_a4Q4fBzU3_0;
	wire w_dff_B_c9lb9DbS0_0;
	wire w_dff_B_QACwt3cS3_0;
	wire w_dff_B_hY2ktPb48_0;
	wire w_dff_B_oAW1pntw0_0;
	wire w_dff_B_qQshgjp18_0;
	wire w_dff_B_UaN4cfuL3_0;
	wire w_dff_B_DAHkaWdf2_0;
	wire w_dff_B_uqs01sJ80_1;
	wire w_dff_B_KCaiDqnp0_1;
	wire w_dff_B_69LiQYJu4_0;
	wire w_dff_B_fqIW3bFR4_0;
	wire w_dff_B_wOMXoJY60_0;
	wire w_dff_B_aUOW9rYY7_0;
	wire w_dff_B_EHHoNx5I6_0;
	wire w_dff_B_Wf6AqbXm9_0;
	wire w_dff_B_jutsZBvQ0_0;
	wire w_dff_B_0v1Dyp9T7_0;
	wire w_dff_B_rcDig1ys9_0;
	wire w_dff_B_QmnjDsoR4_0;
	wire w_dff_B_PpgskbsT6_0;
	wire w_dff_B_Myx8Pffw1_0;
	wire w_dff_B_qGj7Qvvm7_0;
	wire w_dff_B_GNMiNKJC0_0;
	wire w_dff_B_UDIbEXSU4_0;
	wire w_dff_B_WVOelZyV9_0;
	wire w_dff_B_1R4rIOX53_0;
	wire w_dff_B_6dQTneQC5_0;
	wire w_dff_B_IV3JDKjo5_0;
	wire w_dff_B_hnqC9Wmu9_0;
	wire w_dff_B_hm6V1Wnr4_1;
	wire w_dff_B_OWmEd2mP0_0;
	wire w_dff_B_hj10rN1A3_0;
	wire w_dff_B_oBefjrpf0_0;
	wire w_dff_B_TO8PTPjT1_0;
	wire w_dff_B_LhOTchzw1_0;
	wire w_dff_B_BkCZ02jQ4_0;
	wire w_dff_B_V4HvfDVr6_0;
	wire w_dff_B_TNujeIGZ0_0;
	wire w_dff_B_v7k8lmsA5_0;
	wire w_dff_B_nGBsGt7N0_0;
	wire w_dff_B_lrfQuAcZ7_0;
	wire w_dff_B_KLt5u9AE4_0;
	wire w_dff_B_e7fmj5O26_0;
	wire w_dff_B_z52kPYiP3_0;
	wire w_dff_B_sLD9yEMq8_0;
	wire w_dff_B_60rfgGGJ6_0;
	wire w_dff_B_YqnqiXvc0_0;
	wire w_dff_B_Wr43gGI56_0;
	wire w_dff_B_6tvoiiKt9_0;
	wire w_dff_B_xIPwIWEz4_1;
	wire w_dff_B_euO5JJwY7_1;
	wire w_dff_B_6YQPmrv72_1;
	wire w_dff_B_gWcJGIq66_0;
	wire w_dff_B_IAwTJ3XL7_0;
	wire w_dff_B_q2hityIo8_0;
	wire w_dff_B_7jLilQQb2_0;
	wire w_dff_B_dAjVjDeS6_0;
	wire w_dff_B_xzrmSwrU6_0;
	wire w_dff_B_HcsDbYQR9_0;
	wire w_dff_B_yRcSlln43_0;
	wire w_dff_B_2pOQFaYC7_0;
	wire w_dff_B_UO99Msyj3_0;
	wire w_dff_B_2s5Dp15B0_0;
	wire w_dff_B_vTtu1iVF2_0;
	wire w_dff_B_6eV0mzNp9_0;
	wire w_dff_B_bRjX76MI7_0;
	wire w_dff_B_iLxVazOV3_0;
	wire w_dff_B_H0r8ToYp6_0;
	wire w_dff_B_T8LeiYVU3_0;
	wire w_dff_B_G64iDjM79_0;
	wire w_dff_B_pQoMNivd5_0;
	wire w_dff_B_9PryGx0C4_0;
	wire w_dff_B_mO2zrwY48_1;
	wire w_dff_B_bodC3ZIz1_1;
	wire w_dff_B_UXK7apd76_0;
	wire w_dff_B_adkpNogp9_0;
	wire w_dff_B_kTgAz6n64_0;
	wire w_dff_B_LtrCHKnv5_0;
	wire w_dff_B_XTQDDthb0_0;
	wire w_dff_B_V5aBo9AX3_0;
	wire w_dff_B_etyq1JQu7_0;
	wire w_dff_B_iUrlhMZ51_0;
	wire w_dff_B_y0hQiWpe2_0;
	wire w_dff_B_wutJfm3E8_0;
	wire w_dff_B_aIMHjenc7_0;
	wire w_dff_B_fONAimIc1_0;
	wire w_dff_B_zeplCKIF0_0;
	wire w_dff_B_FrhCLHKb5_0;
	wire w_dff_B_gCPQXe5a1_0;
	wire w_dff_B_uAy1IlF57_0;
	wire w_dff_B_kD783my76_0;
	wire w_dff_B_4DerBogf4_0;
	wire w_dff_B_7nGbBVgL3_0;
	wire w_dff_B_fSABNbnM3_0;
	wire w_dff_B_5OLRqP5N6_1;
	wire w_dff_B_dZ9GkMBf3_0;
	wire w_dff_B_9dSPemVe7_0;
	wire w_dff_B_qyBGboWp9_0;
	wire w_dff_B_ROktWTfw4_0;
	wire w_dff_B_qVXjMkcK7_0;
	wire w_dff_B_q1dhFLJr8_0;
	wire w_dff_B_6jKirput2_0;
	wire w_dff_B_07j5ZC1S3_0;
	wire w_dff_B_ZxQWxorr6_0;
	wire w_dff_B_UGROEVBm4_0;
	wire w_dff_B_FsFLOcxn6_0;
	wire w_dff_B_9i6DTtca6_0;
	wire w_dff_B_Uct4yhOZ9_0;
	wire w_dff_B_911KCZeX7_0;
	wire w_dff_B_9T6epfvs1_0;
	wire w_dff_B_0cZr8IVw2_0;
	wire w_dff_B_1A5EE5ey4_0;
	wire w_dff_B_sYnGfNlc2_0;
	wire w_dff_B_3gu5XD3k4_0;
	wire w_dff_B_7meUkI0u9_1;
	wire w_dff_B_jp45zAfo8_1;
	wire w_dff_B_2v01HJmp0_1;
	wire w_dff_B_TDMGOcA01_0;
	wire w_dff_B_LGAgcm9p9_0;
	wire w_dff_B_Ch9jmSvg4_0;
	wire w_dff_B_aMVLQMCi1_0;
	wire w_dff_B_ipVPKn0K3_0;
	wire w_dff_B_7n6S5Bru3_0;
	wire w_dff_B_pibtBhVE9_0;
	wire w_dff_B_94kI7B865_0;
	wire w_dff_B_F3OXVLc20_0;
	wire w_dff_B_ZDwl5qtR0_0;
	wire w_dff_B_IrzLVC3D6_0;
	wire w_dff_B_qE8bZEgv9_0;
	wire w_dff_B_P8ZLFqVY3_0;
	wire w_dff_B_e9EC6BW10_0;
	wire w_dff_B_4psK4a7V2_0;
	wire w_dff_B_izuzLfvx0_0;
	wire w_dff_B_EkczzdOU3_0;
	wire w_dff_B_G0EZjB2W9_0;
	wire w_dff_B_AWnJyqHo5_1;
	wire w_dff_B_K6LR4AuM9_1;
	wire w_dff_B_E6w3HOae8_1;
	wire w_dff_A_gbXeYHvc4_0;
	wire w_dff_A_AOg5Gn541_0;
	wire w_dff_A_Ml7TkT2B2_0;
	wire w_dff_A_WcF6UrZo9_0;
	wire w_dff_A_Tvcmhn8o9_0;
	wire w_dff_A_ivUFOrEV2_0;
	wire w_dff_A_NTmV4l3H9_1;
	wire w_dff_A_zjkof0W22_0;
	wire w_dff_A_RCBIsjoV0_0;
	wire w_dff_A_WjxIsejb9_0;
	wire w_dff_A_iU8dCjJT9_0;
	wire w_dff_A_FA9bbewr7_1;
	wire w_dff_A_jF0uhBbI8_1;
	wire w_dff_A_ZPuicIJu9_0;
	wire w_dff_A_L9DBkmu36_0;
	wire w_dff_A_PKx2ksOL4_0;
	wire w_dff_A_mvxhc2rT6_0;
	wire w_dff_A_B1rvDeUY7_0;
	wire w_dff_A_xKN9JgQ47_0;
	wire w_dff_A_YvJlGhkA9_1;
	wire w_dff_B_tpHjaZk99_0;
	wire w_dff_B_cNw2JI3f9_0;
	wire w_dff_B_Qmi3bZFr2_0;
	wire w_dff_B_e6NDENEr4_0;
	wire w_dff_B_CarBhQgQ1_0;
	wire w_dff_B_o6eCxcjT9_0;
	wire w_dff_B_0DlEfZDK9_0;
	wire w_dff_B_kiATk3UA4_0;
	wire w_dff_B_kcchts2Z2_0;
	wire w_dff_B_3qg3vMfd6_0;
	wire w_dff_B_yf1GRtxK2_0;
	wire w_dff_B_6FhekFqE8_0;
	wire w_dff_B_20dEYXXm0_0;
	wire w_dff_B_B9wMvP9S5_0;
	wire w_dff_B_hUnmoUaW2_0;
	wire w_dff_B_NYOrrIvv7_0;
	wire w_dff_B_pDBKcYpv3_0;
	wire w_dff_B_Ml0byOD53_0;
	wire w_dff_B_7juUKr1R2_0;
	wire w_dff_B_RrZERRcd2_1;
	wire w_dff_B_dy17jKP27_1;
	wire w_dff_B_NN8ODGRh3_1;
	wire w_dff_B_XmPbZfZG9_1;
	wire w_dff_B_o05U0mQu7_1;
	wire w_dff_B_YZHheBjb5_1;
	wire w_dff_B_OLjlaJPK5_1;
	wire w_dff_B_vyZbQ8gT1_1;
	wire w_dff_B_wouDNh8N6_1;
	wire w_dff_B_DoSch3yf7_1;
	wire w_dff_B_RJC5Adxi6_1;
	wire w_dff_B_QwMpfBiy3_1;
	wire w_dff_B_9oldovLf3_1;
	wire w_dff_B_B3uUZbeY6_1;
	wire w_dff_B_BOVlg43r4_1;
	wire w_dff_B_Gyfxcz5j5_1;
	wire w_dff_B_2t2ERVPV8_1;
	wire w_dff_B_blXfLzAg4_1;
	wire w_dff_B_RkdtCZS46_1;
	wire w_dff_B_4HwUVt8K3_1;
	wire w_dff_B_sHmOrsaS5_1;
	wire w_dff_B_fOOBOERz1_1;
	wire w_dff_B_7cptEJjy1_1;
	wire w_dff_B_yqsMho1u5_1;
	wire w_dff_B_ffg94stE7_1;
	wire w_dff_B_xR4NIlIh8_1;
	wire w_dff_B_RBoZkkFK0_1;
	wire w_dff_B_krzhbRS92_1;
	wire w_dff_B_Iye6Ecwo1_1;
	wire w_dff_B_DZLXNBib9_1;
	wire w_dff_B_Gml0mgvj3_1;
	wire w_dff_B_LjvRrO8y4_1;
	wire w_dff_B_xaCtBOEk5_1;
	wire w_dff_B_vNn6kkaM3_1;
	wire w_dff_B_WpYX64Gj6_1;
	wire w_dff_B_JMefzPri5_1;
	wire w_dff_B_2Z3tpeZB3_1;
	wire w_dff_B_K2ojCJ1l3_1;
	wire w_dff_B_V4kzJ57b9_1;
	wire w_dff_B_pl9hiy5V5_1;
	wire w_dff_B_2xEXa9Lg2_1;
	wire w_dff_B_nrRPA6hl1_1;
	wire w_dff_A_EGN9FuvV8_0;
	wire w_dff_A_M0L6Ldl49_2;
	wire w_dff_A_ikw8tFQf0_0;
	wire w_dff_A_THe3ti0z9_0;
	wire w_dff_A_pZ4xnjMO7_1;
	wire w_dff_A_0WmIePRO0_0;
	wire w_dff_A_quVqaCYT7_0;
	wire w_dff_A_LQdcHjuO1_0;
	wire w_dff_A_NhLnp8g58_0;
	wire w_dff_A_nedQqdSK4_0;
	wire w_dff_A_45gEDq8A8_0;
	wire w_dff_A_PDC8W0kX8_0;
	wire w_dff_A_ezaybMgx1_0;
	wire w_dff_A_KwK6V8yu7_0;
	wire w_dff_A_knwgzp2Z0_0;
	wire w_dff_A_MuefKJ1V5_0;
	wire w_dff_A_GYu0ObsI3_1;
	wire w_dff_A_3jKFTcgm2_1;
	wire w_dff_A_wah9tYab7_1;
	wire w_dff_A_MgODUluG2_1;
	wire w_dff_B_lVjrjxam5_3;
	wire w_dff_B_xKL7xCJi0_3;
	wire w_dff_B_EAPQsA3u5_3;
	wire w_dff_B_GNwySFt44_3;
	wire w_dff_B_bSoTJuYO5_3;
	wire w_dff_B_NPn9aIMq5_3;
	wire w_dff_B_snxe0hOv7_3;
	wire w_dff_B_D4re5cxl9_3;
	wire w_dff_B_mVgp88tn7_3;
	wire w_dff_A_vqLHpnx04_0;
	wire w_dff_B_1kgEqDhl6_0;
	wire w_dff_B_Bl42KRDz0_0;
	wire w_dff_B_tnYgqKKr0_0;
	wire w_dff_B_yj2pBBtj0_0;
	wire w_dff_B_evfSjFA60_0;
	wire w_dff_B_5Dr8PS0c4_0;
	wire w_dff_B_lOtE5Dxo0_0;
	wire w_dff_B_UNWoYuVY6_0;
	wire w_dff_B_uWvhuz0m4_0;
	wire w_dff_B_mdTfyy6N0_0;
	wire w_dff_B_PoXiGYQX7_0;
	wire w_dff_B_hMWuKB3c7_0;
	wire w_dff_B_sAlOrGG95_0;
	wire w_dff_B_2G67SzrQ2_0;
	wire w_dff_B_Ta3ZJzoP6_0;
	wire w_dff_B_ZHL8Q97O5_0;
	wire w_dff_B_sAVEzkxK1_0;
	wire w_dff_B_XSJFcWbz3_0;
	wire w_dff_B_QGk5GiZJ1_1;
	wire w_dff_B_orhWyvos4_1;
	wire w_dff_B_LBJurNfu5_1;
	wire w_dff_A_jSks2Rud7_0;
	wire w_dff_A_XLBgMlmK4_0;
	wire w_dff_A_Ea0dKlLg2_0;
	wire w_dff_A_zRPifxMd7_0;
	wire w_dff_A_S6lmztv56_0;
	wire w_dff_A_dgPqd10H5_0;
	wire w_dff_A_LTUJUBnO9_1;
	wire w_dff_B_p4yWtnyB7_1;
	wire w_dff_B_WQkQyFdP6_1;
	wire w_dff_B_4lWuZyOJ7_1;
	wire w_dff_B_kJQ3Yeru5_1;
	wire w_dff_B_IOYW8IEU2_1;
	wire w_dff_B_QDj30bRT2_1;
	wire w_dff_B_wZB3cbBV1_1;
	wire w_dff_B_ArPgHb7L5_1;
	wire w_dff_B_8VZKDMGW1_1;
	wire w_dff_B_ty52Xt5r4_1;
	wire w_dff_B_oEGnkt1Y0_1;
	wire w_dff_B_RYh6DWOm4_0;
	wire w_dff_B_R9p2FXyb6_0;
	wire w_dff_B_UTLi8MrO5_0;
	wire w_dff_B_wkiCQYnH1_0;
	wire w_dff_B_PGKwaFuX5_0;
	wire w_dff_B_DGBkJHNe4_0;
	wire w_dff_B_Z4JsXH4x2_0;
	wire w_dff_A_s1FilO8V2_1;
	wire w_dff_A_Apmot8Vw3_1;
	wire w_dff_A_IC9Kw6aN7_1;
	wire w_dff_A_lFtRrneu6_1;
	wire w_dff_A_WnRpMoNw1_1;
	wire w_dff_B_76XzOmlq6_1;
	wire w_dff_B_0aVmP3li7_1;
	wire w_dff_B_MRe0avuu7_1;
	wire w_dff_B_GXYEBK7E6_1;
	wire w_dff_B_nLG1eGJV1_1;
	wire w_dff_B_UILrsiJX5_1;
	wire w_dff_A_WYo4t0Ao5_0;
	wire w_dff_A_AbwhbL5y8_0;
	wire w_dff_A_rc7LdPML3_0;
	wire w_dff_A_55ySoC9q4_0;
	wire w_dff_A_9WetyqJg1_1;
	wire w_dff_A_2iyUexrb4_1;
	wire w_dff_B_myvVPbSd7_1;
	wire w_dff_B_GlPdXiY42_1;
	wire w_dff_B_aMu63uXL3_1;
	wire w_dff_B_YM5TZrGh1_1;
	wire w_dff_B_3f3TY8vL6_1;
	wire w_dff_B_L8PaIB0r9_1;
	wire w_dff_B_FIwAXgMv5_1;
	wire w_dff_B_2GX8UCpz5_1;
	wire w_dff_B_WINLHToP6_1;
	wire w_dff_B_8SWCRkgH0_1;
	wire w_dff_B_rLIXuRet4_1;
	wire w_dff_B_SeHfmNLb1_1;
	wire w_dff_B_n9LEvZSr3_1;
	wire w_dff_B_8DioIkAS1_1;
	wire w_dff_B_EzH0H0Dj1_1;
	wire w_dff_B_sORWbYPy7_1;
	wire w_dff_B_4TDqEHkO5_1;
	wire w_dff_B_mm87ihes8_1;
	wire w_dff_B_VkGZTCwZ0_1;
	wire w_dff_B_02ECiP6D3_1;
	wire w_dff_B_cIiDLppA7_1;
	wire w_dff_B_8jBPDOJG1_1;
	wire w_dff_B_tneGJfTT2_1;
	wire w_dff_B_TMR7AuPx0_1;
	wire w_dff_B_KzbH4jb70_1;
	wire w_dff_B_L68SKDEG0_1;
	wire w_dff_B_gzxYdMJX9_1;
	wire w_dff_B_ws94ad5S2_1;
	wire w_dff_B_Z5UuduDE7_1;
	wire w_dff_B_lbRTFf7C9_1;
	wire w_dff_B_1l9XPtdR6_1;
	wire w_dff_B_XgoKzcAF1_1;
	wire w_dff_B_Z4VfJ3uk9_1;
	wire w_dff_B_SuvowPje4_1;
	wire w_dff_B_M3qIf25O9_1;
	wire w_dff_B_WKfF4zB30_0;
	wire w_dff_B_S4fAFmOo6_0;
	wire w_dff_B_9MYWyWhf2_0;
	wire w_dff_B_OUB5DwPz1_0;
	wire w_dff_B_iRXoc1t62_0;
	wire w_dff_B_YdoE0Sty7_0;
	wire w_dff_B_V7IvcMX07_0;
	wire w_dff_B_oIpz3zf67_0;
	wire w_dff_B_VrvEw4Un4_0;
	wire w_dff_B_AMlJ6zkX7_0;
	wire w_dff_B_auJqx8k39_1;
	wire w_dff_B_Z5FXd1Xe2_1;
	wire w_dff_B_AOJviqIu3_1;
	wire w_dff_B_PeZZZXUX1_1;
	wire w_dff_B_4FJdQSby2_1;
	wire w_dff_B_vCCl4NZP7_1;
	wire w_dff_B_NhUoNeKe9_1;
	wire w_dff_B_U0qnV3rS4_1;
	wire w_dff_B_q3yblBT83_1;
	wire w_dff_B_6pLzhFzy3_1;
	wire w_dff_B_PYmBybxC3_1;
	wire w_dff_B_Gt6mEJbL1_1;
	wire w_dff_B_Zy2FpPAN4_1;
	wire w_dff_B_ouss8ttY5_1;
	wire w_dff_B_KtJt2y784_1;
	wire w_dff_B_6KR0qW3n2_0;
	wire w_dff_B_P1tojrHZ4_0;
	wire w_dff_B_wMnlK9Bc6_0;
	wire w_dff_B_x10XzrrB6_0;
	wire w_dff_B_xI8VjsDx1_0;
	wire w_dff_B_0Zf1eCYS9_0;
	wire w_dff_B_71UCjA3L0_0;
	wire w_dff_B_bjU1o1PW6_0;
	wire w_dff_B_Q6MOeho38_0;
	wire w_dff_B_O4NrzNrM6_0;
	wire w_dff_B_nC3ScYUk1_0;
	wire w_dff_B_OIO3nJy82_0;
	wire w_dff_B_tuPQzDkg2_0;
	wire w_dff_B_ne1VmxbK3_0;
	wire w_dff_B_yqEFetps2_0;
	wire w_dff_B_Civl0PfK2_0;
	wire w_dff_B_ppCAZ6H29_0;
	wire w_dff_B_cNpLALwU9_0;
	wire w_dff_B_j5DK7ZyH8_0;
	wire w_dff_B_MTWm3H7E2_1;
	wire w_dff_B_MyNQdqJ97_1;
	wire w_dff_B_tmwvDAz70_1;
	wire w_dff_B_4BFDwHec1_1;
	wire w_dff_B_LPquafu73_1;
	wire w_dff_B_2JSczoHV2_1;
	wire w_dff_B_paZagDH31_1;
	wire w_dff_B_acv8bJlo5_1;
	wire w_dff_B_zE3SP0cj1_1;
	wire w_dff_B_drglUFN87_1;
	wire w_dff_B_pwSHXP8X2_1;
	wire w_dff_B_oMreKgB77_1;
	wire w_dff_B_ENz6bOd40_1;
	wire w_dff_B_2hUhRn792_1;
	wire w_dff_B_55ngfZWA2_1;
	wire w_dff_B_EBtMAoV48_1;
	wire w_dff_B_bArBZE0s8_1;
	wire w_dff_B_UwkZLPuQ0_1;
	wire w_dff_B_8c3WVdlW9_1;
	wire w_dff_B_6i5RmBAb4_1;
	wire w_dff_B_Urhfa7Ty2_1;
	wire w_dff_B_2eHnOBm39_1;
	wire w_dff_B_J0pQXekf9_1;
	wire w_dff_B_g2lPKBsA1_1;
	wire w_dff_B_S2egDuPP7_1;
	wire w_dff_B_3sYPQFlP3_1;
	wire w_dff_B_fxewUeBb5_1;
	wire w_dff_B_HLuv4sqU8_1;
	wire w_dff_A_gzOtYmBM1_0;
	wire w_dff_A_gS3Eofon3_0;
	wire w_dff_A_P2eVeULF3_0;
	wire w_dff_A_nn4ttwY30_0;
	wire w_dff_A_4rwhmoIk3_0;
	wire w_dff_A_gXwNeGG20_0;
	wire w_dff_A_BDFNMZel4_0;
	wire w_dff_A_LPflsroB5_0;
	wire w_dff_A_To32fPpX3_0;
	wire w_dff_A_2eqtmcpk1_0;
	wire w_dff_A_XR3oOArB3_1;
	wire w_dff_A_G7amS7XX3_0;
	wire w_dff_A_pbfR3EOA6_0;
	wire w_dff_A_BbXgFDnt3_0;
	wire w_dff_A_O0QeAVG97_0;
	wire w_dff_A_depvRx9i3_0;
	wire w_dff_A_x9nhREvs5_0;
	wire w_dff_A_IWURhLYv1_1;
	wire w_dff_A_gACeJiaX0_1;
	wire w_dff_A_syYjlyYb9_1;
	wire w_dff_A_rtE8NXtz0_1;
	wire w_dff_A_Ypq6KGFq9_1;
	wire w_dff_A_Tpl2WCYT4_1;
	wire w_dff_A_2ZM4WqgQ8_1;
	wire w_dff_B_2ZLJ7NYe7_0;
	wire w_dff_B_uBTTkax61_0;
	wire w_dff_B_oCnSXvnh7_0;
	wire w_dff_B_v1hnzv5y0_0;
	wire w_dff_B_LlDicOws2_0;
	wire w_dff_B_07lxF3nb9_0;
	wire w_dff_B_6Cb1L1au1_0;
	wire w_dff_B_mAskDXiv5_0;
	wire w_dff_B_Xu8XUfAu2_0;
	wire w_dff_B_0ZEJd4oe8_0;
	wire w_dff_B_7ISTpVOO4_0;
	wire w_dff_B_Wl5DfmZW0_0;
	wire w_dff_B_8UJhFz3S7_0;
	wire w_dff_B_7e9tf7xK5_0;
	wire w_dff_B_ct5tzXPR4_0;
	wire w_dff_B_uOohp7LV9_0;
	wire w_dff_B_UYuDaZAK2_0;
	wire w_dff_B_rvhzNEDX1_0;
	wire w_dff_B_FNMQBBlP1_0;
	wire w_dff_B_ooJGcptk8_1;
	wire w_dff_B_9CqpIqcP7_1;
	wire w_dff_B_vIhROdJC9_1;
	wire w_dff_B_O0o0c5Bu4_1;
	wire w_dff_B_hvggMN5O5_1;
	wire w_dff_B_RusAHTLs7_1;
	wire w_dff_B_tMxI4zBR4_1;
	wire w_dff_B_rSccarmi8_1;
	wire w_dff_B_r0OYv9tN8_1;
	wire w_dff_B_g39610bw8_1;
	wire w_dff_B_6uiVvotc0_1;
	wire w_dff_B_5f4B6GHy7_1;
	wire w_dff_B_QW6eZToC4_1;
	wire w_dff_B_zBUb8bse1_1;
	wire w_dff_B_b9b6f4gL0_1;
	wire w_dff_B_3D7jzu8O1_1;
	wire w_dff_B_NQuquT6l6_0;
	wire w_dff_B_NxCGFaZD2_0;
	wire w_dff_B_etRqYYem7_0;
	wire w_dff_B_Des77N1z8_0;
	wire w_dff_B_tqeZaejH9_0;
	wire w_dff_B_OPvJpz5I7_0;
	wire w_dff_B_nlz3gFFR6_0;
	wire w_dff_B_7WiQ2i248_0;
	wire w_dff_B_IE3mTKN15_0;
	wire w_dff_B_ihkLqLvt3_0;
	wire w_dff_B_9BEy8dXA3_0;
	wire w_dff_B_zoa86Shm5_0;
	wire w_dff_B_4xUKJLD13_0;
	wire w_dff_B_6f5qogMe0_0;
	wire w_dff_A_HRL9jvSt8_0;
	wire w_dff_A_JgzjklZa3_2;
	wire w_dff_A_o4xpqt266_2;
	wire w_dff_A_TuZO65Nc5_0;
	wire w_dff_A_mohINigu2_0;
	wire w_dff_A_GoHp2ciy6_0;
	wire w_dff_A_X7HYLeqh9_0;
	wire w_dff_A_VSkI485R4_0;
	wire w_dff_A_67Cq9LhJ9_0;
	wire w_dff_A_cdyTpUGQ7_0;
	wire w_dff_A_A7G5W8cI1_0;
	wire w_dff_A_X5ele9mj2_0;
	wire w_dff_A_vMs6C9cH4_1;
	wire w_dff_A_nRJ4LMDu5_1;
	wire w_dff_B_B6msR1jS2_3;
	wire w_dff_B_IBMPP6gy4_3;
	wire w_dff_B_WRqTiJIW3_3;
	wire w_dff_B_39zhnG930_3;
	wire w_dff_B_YLTODweL4_3;
	wire w_dff_B_JiPs2Uey3_3;
	wire w_dff_B_tcAAeZDE9_3;
	wire w_dff_B_ErmE05f45_3;
	wire w_dff_B_iD6VkauB9_3;
	wire w_dff_B_bCwz9kcY5_3;
	wire w_dff_B_ilgOphnQ3_3;
	wire w_dff_B_amnl6vVa9_0;
	wire w_dff_B_UgiRTvBr2_0;
	wire w_dff_B_6dnbct4N1_0;
	wire w_dff_B_bHUa4NyD8_0;
	wire w_dff_B_jMgib4gx2_0;
	wire w_dff_B_GsWcKexc1_0;
	wire w_dff_B_yOalO2bq8_0;
	wire w_dff_B_qgMjZx972_0;
	wire w_dff_B_NrmhjzzI0_0;
	wire w_dff_B_EA9YhuCd8_0;
	wire w_dff_B_dlEDUn5B4_0;
	wire w_dff_B_O4dvStjK1_0;
	wire w_dff_B_mlEKmy3i0_0;
	wire w_dff_B_14vUnwef5_0;
	wire w_dff_B_BkagvVka9_0;
	wire w_dff_B_MVrJ394e1_0;
	wire w_dff_B_sLrBGO7P3_0;
	wire w_dff_B_WYnrzB081_0;
	wire w_dff_B_cefAZnSV1_0;
	wire w_dff_B_VXfN6Rxl6_0;
	wire w_dff_B_WPf0VP3U1_0;
	wire w_dff_B_QbfSDge96_0;
	wire w_dff_B_tsAkeTqc0_0;
	wire w_dff_B_ICqstP6q0_0;
	wire w_dff_B_Rt9wbP2j2_0;
	wire w_dff_B_TIVDoktD9_0;
	wire w_dff_B_ajr3RozC7_0;
	wire w_dff_B_4rw2JdVK8_0;
	wire w_dff_B_ku1WFQUH9_0;
	wire w_dff_B_LWtLpZwX1_0;
	wire w_dff_B_SVQGD7k93_0;
	wire w_dff_B_QnczFIBi2_0;
	wire w_dff_B_DMV76sid3_0;
	wire w_dff_B_shEHb3tA0_0;
	wire w_dff_B_5MBjdzIM7_1;
	wire w_dff_B_WOsrwc1U7_1;
	wire w_dff_B_R8Mb56158_1;
	wire w_dff_B_RcASiONo7_1;
	wire w_dff_B_QyonVpYp2_1;
	wire w_dff_B_pdZk2Oli6_1;
	wire w_dff_B_H5v8wQ9J8_1;
	wire w_dff_B_GxQiWWLU4_1;
	wire w_dff_B_qWF2oG3R3_1;
	wire w_dff_B_ENOlmBFP4_1;
	wire w_dff_B_D5AQM6tC9_1;
	wire w_dff_B_fjmZhyw96_1;
	wire w_dff_B_2LjtTI2E8_1;
	wire w_dff_B_4JCscMMW8_1;
	wire w_dff_B_JeoGxJYG0_1;
	wire w_dff_B_IkB6CCCa3_1;
	wire w_dff_B_KzMwOGDP0_1;
	wire w_dff_B_C4opgz5m0_1;
	wire w_dff_B_SfarNTi77_1;
	wire w_dff_B_AH4fPRSj2_1;
	wire w_dff_B_MF4eaZkD4_1;
	wire w_dff_B_MSftF2H93_1;
	wire w_dff_B_EEzYRZkM4_1;
	wire w_dff_A_RHfzNSPg1_1;
	wire w_dff_A_rystDuU95_1;
	wire w_dff_A_zbA8LNwf7_1;
	wire w_dff_A_5VbY4wKc4_1;
	wire w_dff_A_ZzkiHjCq1_1;
	wire w_dff_A_VIeei1bg2_1;
	wire w_dff_A_i1Jer8HA9_1;
	wire w_dff_A_vKxGeqiP9_1;
	wire w_dff_A_9ms7kQtp6_1;
	wire w_dff_A_DOF0jgwQ0_1;
	wire w_dff_A_9bemO3lg7_1;
	wire w_dff_A_cOifCqaX4_1;
	wire w_dff_A_4GGle7XC4_1;
	wire w_dff_A_rW7yqhoM0_1;
	wire w_dff_A_9uD4KlcF1_2;
	wire w_dff_A_eriU6EEM6_2;
	wire w_dff_A_PM4ciDnd2_2;
	wire w_dff_A_zhNNRsm78_2;
	wire w_dff_A_C9Tsq5js6_2;
	wire w_dff_A_yRGbStaz4_2;
	wire w_dff_A_YrGbzQji2_2;
	wire w_dff_A_JOxejTlT8_2;
	wire w_dff_A_ixhmkYSC6_2;
	wire w_dff_A_fW8OGSka8_2;
	wire w_dff_B_zJcJ2KQI2_1;
	wire w_dff_B_5MYgQLxb5_1;
	wire w_dff_B_NddqbPXm3_1;
	wire w_dff_B_9Tgjv4SM2_1;
	wire w_dff_B_9IuPFjWc3_1;
	wire w_dff_B_f6Jh1WVy9_1;
	wire w_dff_B_UydghEbs2_1;
	wire w_dff_B_UNhxR9L72_1;
	wire w_dff_B_shbRryZK9_1;
	wire w_dff_B_aM4m7D2d8_1;
	wire w_dff_B_iluRJHjN2_1;
	wire w_dff_B_czxlWPxq3_1;
	wire w_dff_B_sndVJQE01_1;
	wire w_dff_B_1VemC9UF1_1;
	wire w_dff_B_GsPBGEDN6_1;
	wire w_dff_B_NUxOlpXU9_1;
	wire w_dff_B_rZ3P8Ezx8_1;
	wire w_dff_B_2hqh731n3_1;
	wire w_dff_B_B0nDGpt26_1;
	wire w_dff_B_nPaF7WtD1_1;
	wire w_dff_B_FGZyo1Ue0_1;
	wire w_dff_B_IcnpIemx3_1;
	wire w_dff_B_HgvF8hE49_1;
	wire w_dff_A_GgUroV2W1_1;
	wire w_dff_A_jVSXcdB16_1;
	wire w_dff_A_CJWeJFSh3_1;
	wire w_dff_A_Tirp1Pd82_1;
	wire w_dff_A_LG0FfJmp8_1;
	wire w_dff_A_Du1CZ2Xa5_1;
	wire w_dff_A_0iMtQxWI2_1;
	wire w_dff_A_OkZGQjhi2_1;
	wire w_dff_A_yzQhIqpR5_1;
	wire w_dff_A_s9dsHqFi9_1;
	wire w_dff_A_MWVJ7jpg3_1;
	wire w_dff_A_UFcy6zM52_1;
	wire w_dff_A_eR5qvQQc5_1;
	wire w_dff_A_E2vII9n89_1;
	wire w_dff_A_j6gsq6um5_2;
	wire w_dff_A_upXRwyB17_2;
	wire w_dff_A_KBLre0CC9_2;
	wire w_dff_A_Ee7j38Og1_2;
	wire w_dff_A_eM0UDtrK2_2;
	wire w_dff_A_GErvG4gT4_2;
	wire w_dff_A_e9wGZ5i35_2;
	wire w_dff_A_irKNyDSR9_2;
	wire w_dff_A_v4Ji4mre7_2;
	wire w_dff_A_w3eUXdrG5_2;
	wire w_dff_B_nyYvB2tj6_1;
	wire w_dff_B_xy3ImAAq3_1;
	wire w_dff_B_2oyRlj3a4_1;
	wire w_dff_B_iVNGJi6z1_1;
	wire w_dff_B_eC6dIvtR0_1;
	wire w_dff_B_BLm1o4kV1_1;
	wire w_dff_B_dJ4bMt2e9_1;
	wire w_dff_B_eT8mCMpY8_1;
	wire w_dff_B_4BHqEVxU3_1;
	wire w_dff_B_K8PIzCKL6_1;
	wire w_dff_B_wKEkvZPw4_1;
	wire w_dff_B_4zNlqT5V6_1;
	wire w_dff_B_AKd0NSDS6_1;
	wire w_dff_B_OXG23iN70_1;
	wire w_dff_B_XuTEtqXe2_1;
	wire w_dff_B_uy8rerwp8_1;
	wire w_dff_B_Ulx3NKyY5_1;
	wire w_dff_B_8ZOx98qG7_1;
	wire w_dff_B_IUuIk5yZ6_1;
	wire w_dff_B_UyIHkBuD5_1;
	wire w_dff_B_mnr5EtXf9_1;
	wire w_dff_B_Y2Qk5IFA0_1;
	wire w_dff_B_xFRH1E7d1_1;
	wire w_dff_B_UCyxkDuz9_1;
	wire w_dff_B_IEpbaqTd3_1;
	wire w_dff_B_aUeayiQz7_1;
	wire w_dff_B_sxQEjlpR4_1;
	wire w_dff_B_SuZgzeC56_1;
	wire w_dff_B_FmqYyeU43_1;
	wire w_dff_B_HaorQlKU5_1;
	wire w_dff_B_woz3DQCA1_1;
	wire w_dff_B_d5Gs0Tdi7_1;
	wire w_dff_B_wFSc6V042_1;
	wire w_dff_B_GE4vzV4B0_1;
	wire w_dff_B_Ik53PXFx7_1;
	wire w_dff_B_plbUrMv81_1;
	wire w_dff_B_RmVWAyyF7_1;
	wire w_dff_B_yw8HwcB69_1;
	wire w_dff_B_WxCQHscR9_1;
	wire w_dff_B_hEb9Ov7e2_1;
	wire w_dff_B_aiHHvdUR5_1;
	wire w_dff_B_w0UPXMMj5_1;
	wire w_dff_B_BB80w2h76_1;
	wire w_dff_B_S1TlZL3Q5_1;
	wire w_dff_B_OyrKFmYT7_1;
	wire w_dff_B_SHDFiHai4_1;
	wire w_dff_B_r4nl3ba44_1;
	wire w_dff_B_1R4LT2rQ8_1;
	wire w_dff_B_y6LL5sP02_1;
	wire w_dff_B_d7VdmAkg5_1;
	wire w_dff_B_CKTWOprv3_1;
	wire w_dff_B_HmYxEVDQ9_1;
	wire w_dff_B_PrCjGr6S1_1;
	wire w_dff_B_6hw44P118_1;
	wire w_dff_B_qOaxueCp3_1;
	wire w_dff_B_wYx89UmX7_1;
	wire w_dff_B_3ghB2Ggm3_1;
	wire w_dff_B_5yEehwxw9_1;
	wire w_dff_B_enloygGK2_1;
	wire w_dff_B_7RHKiZSp3_1;
	wire w_dff_B_mkvQskNg2_1;
	wire w_dff_B_wQ5qyDNm1_1;
	wire w_dff_B_2dFyI4c60_1;
	wire w_dff_B_D6l5Yjcy1_1;
	wire w_dff_B_cjjzdCiv1_1;
	wire w_dff_B_YWc2PxDc3_1;
	wire w_dff_B_aqcr2WXc9_1;
	wire w_dff_B_5wark3kh5_1;
	wire w_dff_B_FG9q5yje3_1;
	wire w_dff_B_RzXeeNyg4_1;
	wire w_dff_B_HVfQU3664_1;
	wire w_dff_B_gfY1tcdS5_1;
	wire w_dff_B_Yv3NyAhq8_1;
	wire w_dff_B_JN1TonOg3_1;
	wire w_dff_B_7z5hVVUh6_1;
	wire w_dff_B_R0q1cWjx6_1;
	wire w_dff_B_F0Pbj0uN5_1;
	wire w_dff_B_IZTA4Esk5_1;
	wire w_dff_B_lKE4yU3v2_1;
	wire w_dff_B_VTghs1Pl6_1;
	wire w_dff_B_Gb7dGKxX2_1;
	wire w_dff_B_lBuFHirz3_1;
	wire w_dff_B_wjcyD9Pv7_1;
	wire w_dff_B_4aH8sZ125_1;
	wire w_dff_B_Q1RHRg5T0_1;
	wire w_dff_B_qjpJX1UX7_1;
	wire w_dff_B_ugSKk3lK5_1;
	wire w_dff_B_mVGjxRFb1_1;
	wire w_dff_B_UhhF2aeY9_1;
	wire w_dff_B_qck1SFfG3_1;
	wire w_dff_B_Ywku2r8g2_0;
	wire w_dff_B_fRU7VHFG1_0;
	wire w_dff_B_rQdDj2eA7_0;
	wire w_dff_B_CdO5itrP2_0;
	wire w_dff_B_3DfPf54M9_0;
	wire w_dff_B_mq5e2Zzx6_0;
	wire w_dff_B_9Sia1E4D3_0;
	wire w_dff_B_QDndUrLm7_0;
	wire w_dff_B_ABFe8TIy3_0;
	wire w_dff_B_jzHHyC1G5_0;
	wire w_dff_B_nZuCHGPA4_0;
	wire w_dff_B_uxJvCPl38_0;
	wire w_dff_B_Z8XCAVaB1_0;
	wire w_dff_B_ouBIezaM0_0;
	wire w_dff_B_7Mx015AW6_0;
	wire w_dff_B_SItuqPlM5_0;
	wire w_dff_B_ZVYJLPdy5_0;
	wire w_dff_B_zNNL6OLI0_0;
	wire w_dff_B_11Y5fuYu3_0;
	wire w_dff_B_wZ4qtbJV6_0;
	wire w_dff_B_B6ZabqjA5_0;
	wire w_dff_B_iYc4xeuz8_0;
	wire w_dff_B_YUSImXH81_0;
	wire w_dff_B_fuor0P728_0;
	wire w_dff_B_vnyppdtj0_0;
	wire w_dff_B_hDjk5vER8_0;
	wire w_dff_B_rBb9Fa5m0_0;
	wire w_dff_B_z22eYMUi6_0;
	wire w_dff_B_0i2kTdtc2_1;
	wire w_dff_B_NO5SrzkV7_0;
	wire w_dff_A_UpHFzeke5_0;
	wire w_dff_A_7wxXQokn0_0;
	wire w_dff_B_b8J3pfmx8_0;
	wire w_dff_B_SFlZDlf13_0;
	wire w_dff_B_8TqIhvGq3_0;
	wire w_dff_B_J1AkRO136_1;
	wire w_dff_B_ib2IL73b4_1;
	wire w_dff_B_p1RAyhWe0_1;
	wire w_dff_B_ZqKnkvmN1_1;
	wire w_dff_B_ojDaT3h42_1;
	wire w_dff_B_W3Dv9XHm7_0;
	wire w_dff_B_lb2sWyLx1_0;
	wire w_dff_A_cssLASeX9_0;
	wire w_dff_B_GELGpxoG6_1;
	wire w_dff_A_yiq9g2aP7_2;
	wire w_dff_A_AB6PTBb39_2;
	wire w_dff_A_QIqXiJiq1_0;
	wire w_dff_A_lgyLa82g0_0;
	wire w_dff_A_e0HmERPy0_0;
	wire w_dff_A_OHwws77V4_0;
	wire w_dff_A_f4Qd0c5u7_1;
	wire w_dff_B_K8LUhpwg3_3;
	wire w_dff_B_Pns1XHaU6_3;
	wire w_dff_A_77FCiIJy7_0;
	wire w_dff_B_y7USFW1T9_1;
	wire w_dff_A_XjBaWqj13_0;
	wire w_dff_B_u8AEOMbS8_1;
	wire w_dff_B_v6bKkAAY4_1;
	wire w_dff_B_nfYiIvAu1_1;
	wire w_dff_A_drZdhkdz7_2;
	wire w_dff_A_7DptGaxU0_2;
	wire w_dff_A_Rd9Qk2go1_2;
	wire w_dff_A_8Hfju6PD7_2;
	wire w_dff_A_tG9trZYe2_2;
	wire w_dff_A_0RBPngsx4_2;
	wire w_dff_A_tv11bPYw0_2;
	wire w_dff_A_dUIBOcCW1_2;
	wire w_dff_A_zmpyFrKI5_2;
	wire w_dff_A_Ae76oq8l4_1;
	wire w_dff_A_RA4bUFWW9_1;
	wire w_dff_A_4yHa4Zxk5_1;
	wire w_dff_A_CJXrbhge1_1;
	wire w_dff_A_xmPDzEJ46_1;
	wire w_dff_A_y6WFFCKg1_1;
	wire w_dff_A_Dwcuz1Mt6_1;
	wire w_dff_A_fkiZc9bO0_1;
	wire w_dff_A_9NadUDZn9_1;
	wire w_dff_A_YMMn1aJu8_1;
	wire w_dff_B_ZiixEKxx1_1;
	wire w_dff_B_ZsMevCQX5_1;
	wire w_dff_B_JKDdWWuv9_1;
	wire w_dff_B_kwom3u9N4_1;
	wire w_dff_B_GKmUyL8K8_1;
	wire w_dff_B_bDlfFRgC2_1;
	wire w_dff_B_2FUUdo6f3_1;
	wire w_dff_A_NA9Df6H68_1;
	wire w_dff_B_9zmzvveo6_1;
	wire w_dff_B_N2ElJB7k8_1;
	wire w_dff_B_vucXC8zj6_1;
	wire w_dff_B_okWyP26V2_1;
	wire w_dff_B_IN16bStA5_1;
	wire w_dff_B_chb4fUGz8_1;
	wire w_dff_B_wsuO4F6W8_1;
	wire w_dff_A_CvaPLRfG1_1;
	wire w_dff_A_eUZQ0gCo5_1;
	wire w_dff_A_hxGff9QT8_0;
	wire w_dff_A_l2d0QREj0_0;
	wire w_dff_A_AL4TBzB66_0;
	wire w_dff_A_oND0CmAJ6_1;
	wire w_dff_A_EEJ6wBEC7_1;
	wire w_dff_A_TaBuKhQ45_1;
	wire w_dff_A_Zmmqp0qp7_1;
	wire w_dff_A_0XMBlSB18_2;
	wire w_dff_B_piuNxwIg6_3;
	wire w_dff_B_brFdKLeN3_3;
	wire w_dff_B_lwwr2A2p8_3;
	wire w_dff_B_sUQf3Mlt0_3;
	wire w_dff_B_aSEUAJJ42_3;
	wire w_dff_B_cDJVJztp5_3;
	wire w_dff_B_EVhQzDYu4_3;
	wire w_dff_B_faHhOZgZ0_3;
	wire w_dff_B_kD7cOaV19_3;
	wire w_dff_B_9csyNqWX5_3;
	wire w_dff_A_TL0ht9Jp2_0;
	wire w_dff_B_A7oqnMQB8_0;
	wire w_dff_B_HiDGTUnB7_0;
	wire w_dff_A_b30ZD7DE2_0;
	wire w_dff_A_QuYbWtTq1_0;
	wire w_dff_A_jTuHUfu36_0;
	wire w_dff_A_PyNPhz278_0;
	wire w_dff_A_LuUV5yCQ1_2;
	wire w_dff_A_uLWTeDtJ1_2;
	wire w_dff_B_oSMEsVHY2_1;
	wire w_dff_A_PzJQwF4I3_0;
	wire w_dff_A_uvSGRqJ13_0;
	wire w_dff_B_HPmUIL054_2;
	wire w_dff_B_9fwOs6c77_2;
	wire w_dff_B_Thd5Vae35_2;
	wire w_dff_B_eDjis2yY9_2;
	wire w_dff_B_Qw7943Sf2_2;
	wire w_dff_B_SSx1WpRp3_2;
	wire w_dff_B_Ao5tScGk0_2;
	wire w_dff_B_pJL1NtXi5_2;
	wire w_dff_B_8R5WqX8z9_2;
	wire w_dff_B_fB6juIMr0_2;
	wire w_dff_B_aFYCOJbS2_2;
	wire w_dff_B_XDInrnuN8_2;
	wire w_dff_B_HaRs99yT4_2;
	wire w_dff_B_VnWqcvaT1_2;
	wire w_dff_B_vFv4DzFa8_2;
	wire w_dff_B_KnMLcJqJ3_2;
	wire w_dff_B_etcTJXVC3_2;
	wire w_dff_B_enkNTEp98_2;
	wire w_dff_B_gHLFmskD2_2;
	wire w_dff_B_TovuJMhW8_2;
	wire w_dff_B_fa94FOAF1_2;
	wire w_dff_B_ZTGF89tH2_2;
	wire w_dff_B_L8UPxx8e1_2;
	wire w_dff_B_PPiahgxs9_2;
	wire w_dff_B_F2zmgtPn2_2;
	wire w_dff_B_N8xjebfb1_2;
	wire w_dff_A_tFCKOFNL4_1;
	wire w_dff_A_IlZsEDUK1_0;
	wire w_dff_A_CEcT4a6e9_0;
	wire w_dff_A_4VV4GkaV1_0;
	wire w_dff_A_2PBcT4QF6_0;
	wire w_dff_A_svF7vANG6_0;
	wire w_dff_A_xHISj5mx7_0;
	wire w_dff_A_BMspYHVI9_0;
	wire w_dff_A_lnoOPcSL4_0;
	wire w_dff_A_c6YR15Kn0_0;
	wire w_dff_A_FdUmNxvz7_0;
	wire w_dff_A_14FSDXLG3_0;
	wire w_dff_A_DxmdopC61_0;
	wire w_dff_A_q56tQ0zC5_0;
	wire w_dff_A_4GaniFXN0_0;
	wire w_dff_A_Bs74xH8Y3_0;
	wire w_dff_A_M2SiTpMy0_0;
	wire w_dff_A_9UBehGnl5_0;
	wire w_dff_A_Q94LseRR7_0;
	wire w_dff_A_2hKHFtfk7_0;
	wire w_dff_A_CWJCZpaH4_0;
	wire w_dff_A_ls03wzJm9_0;
	wire w_dff_A_RdMGEhjR3_0;
	wire w_dff_A_7XceqW1U3_0;
	wire w_dff_A_LO1GnWZF9_0;
	wire w_dff_A_W9PKCXPe5_0;
	wire w_dff_A_6oc6LFNX4_0;
	wire w_dff_A_54vrj7St8_0;
	wire w_dff_A_Bir94Gwe0_1;
	wire w_dff_A_adTFoNZk7_0;
	wire w_dff_A_eBaIsSic1_0;
	wire w_dff_A_8RzHka1B2_0;
	wire w_dff_A_y9ZXT5La9_0;
	wire w_dff_A_WuxbsWnc9_0;
	wire w_dff_A_QZ4T2PjB9_0;
	wire w_dff_A_soBDb5fj5_0;
	wire w_dff_A_jh2zniJb6_0;
	wire w_dff_A_F0lzzu2m0_0;
	wire w_dff_A_FQCsMyot8_0;
	wire w_dff_A_buoWIpoR5_0;
	wire w_dff_A_HmLMOibi4_0;
	wire w_dff_A_uxw6RwgI6_0;
	wire w_dff_A_qehoy7UX7_0;
	wire w_dff_A_tpqGvAKw7_0;
	wire w_dff_A_YoZ5tzuC2_0;
	wire w_dff_A_Hjm9D9fg0_0;
	wire w_dff_A_BoDHA4QK7_0;
	wire w_dff_A_ovB82ksM3_0;
	wire w_dff_A_nzWHdgM34_0;
	wire w_dff_A_Xtpe54Fi3_0;
	wire w_dff_A_QtOT82I86_0;
	wire w_dff_A_PKMcqa5r9_0;
	wire w_dff_A_2Z02vyXc3_0;
	wire w_dff_A_1aBOBSgY5_0;
	wire w_dff_A_6ElIMykj1_0;
	wire w_dff_A_VFKfeA661_0;
	wire w_dff_A_H773dteS1_1;
	wire w_dff_A_Wrb6XQ9M3_0;
	wire w_dff_A_gjolEoZm8_0;
	wire w_dff_A_cDiMoD0l6_0;
	wire w_dff_A_pVAc7uwU2_0;
	wire w_dff_A_LSTP7cjW7_0;
	wire w_dff_A_sqniW66f4_0;
	wire w_dff_A_6dTVZnDz5_0;
	wire w_dff_A_NbDrMkrj4_0;
	wire w_dff_A_Xte8DpDg1_0;
	wire w_dff_A_qbbP2Bre2_0;
	wire w_dff_A_Js5nZOvU1_0;
	wire w_dff_A_QfOule055_0;
	wire w_dff_A_wXdDOOIp2_0;
	wire w_dff_A_5cRvcW8U0_0;
	wire w_dff_A_eSnQq50H8_0;
	wire w_dff_A_u36tr0Uk9_0;
	wire w_dff_A_LyD1bGZw7_0;
	wire w_dff_A_9ZGrWXR51_0;
	wire w_dff_A_IezzxeHx2_0;
	wire w_dff_A_gTe6RvbS9_0;
	wire w_dff_A_nsvwWbP60_0;
	wire w_dff_A_ePmEMqIg2_0;
	wire w_dff_A_eCCmkl9E7_0;
	wire w_dff_A_LAdfQCgz7_0;
	wire w_dff_A_x3SHnhVE1_0;
	wire w_dff_A_MjbNilE46_0;
	wire w_dff_A_8g2vocKL1_0;
	wire w_dff_A_H1rIXdYd7_1;
	wire w_dff_A_GXWBBTVX5_0;
	wire w_dff_A_XpN5hJdD3_0;
	wire w_dff_A_m7DBhqto6_0;
	wire w_dff_A_7aWAnjDg8_0;
	wire w_dff_A_wSEwcVj96_0;
	wire w_dff_A_w9lVZ12u0_0;
	wire w_dff_A_MPHbYqjQ9_0;
	wire w_dff_A_JznfRGiE9_0;
	wire w_dff_A_pyKXWd1D1_0;
	wire w_dff_A_ZD85smjf6_0;
	wire w_dff_A_GW7ScZib9_0;
	wire w_dff_A_Uug7XAZ92_0;
	wire w_dff_A_nKbHBH6W0_0;
	wire w_dff_A_zxN7p3io2_0;
	wire w_dff_A_mpS3mQ7V7_0;
	wire w_dff_A_O8nC4jad7_0;
	wire w_dff_A_YHcjhaOu1_0;
	wire w_dff_A_ndtwybAt6_0;
	wire w_dff_A_b8kuF6Xe6_0;
	wire w_dff_A_Mwrz6Mvt2_0;
	wire w_dff_A_DuFWqoLP1_0;
	wire w_dff_A_mcOIk3Fx2_0;
	wire w_dff_A_5DZM0TFf2_0;
	wire w_dff_A_7iyGSHtR8_0;
	wire w_dff_A_TajBF7E89_0;
	wire w_dff_A_MNmoIlqo7_0;
	wire w_dff_A_QA8TyQ3f3_1;
	wire w_dff_A_QBROjjOd0_0;
	wire w_dff_A_c9iPnlNf3_0;
	wire w_dff_A_s4LwXeps4_0;
	wire w_dff_A_4JoHyEzQ7_0;
	wire w_dff_A_9z6bFZaj2_0;
	wire w_dff_A_7OVFCuU01_0;
	wire w_dff_A_7TwucoQR3_0;
	wire w_dff_A_58Um3fd75_0;
	wire w_dff_A_LkdHHjQe9_0;
	wire w_dff_A_mVil7j4e0_0;
	wire w_dff_A_o2CqpAva4_0;
	wire w_dff_A_mjBr6zl40_0;
	wire w_dff_A_ryB8kxCI7_0;
	wire w_dff_A_qBtYsWeu9_0;
	wire w_dff_A_5UHIoTlL9_0;
	wire w_dff_A_JJL6Zjyo9_0;
	wire w_dff_A_s7bcHlga8_0;
	wire w_dff_A_S2Taeel45_0;
	wire w_dff_A_ByNIFjWL6_0;
	wire w_dff_A_Qwf1AUPT8_0;
	wire w_dff_A_z9w1kiHo4_0;
	wire w_dff_A_NpZ04Uab0_0;
	wire w_dff_A_KNT9MsG93_0;
	wire w_dff_A_ibWsWtvQ8_0;
	wire w_dff_A_7780QqlZ4_0;
	wire w_dff_A_SyA7bhbB9_0;
	wire w_dff_A_HCUTE1hH8_1;
	wire w_dff_A_D2th1dxC8_0;
	wire w_dff_A_zQc6KNTr9_0;
	wire w_dff_A_WFdFNGRX2_0;
	wire w_dff_A_u17W9g6y4_0;
	wire w_dff_A_zNnRUM9D8_0;
	wire w_dff_A_84A0Ie8H4_0;
	wire w_dff_A_dLbxZUUK2_0;
	wire w_dff_A_899P7Vdo1_0;
	wire w_dff_A_K275nXcx4_0;
	wire w_dff_A_56RexwDu0_0;
	wire w_dff_A_SWxtiXqn4_0;
	wire w_dff_A_PQ6AwPzD4_0;
	wire w_dff_A_mR56OXx80_0;
	wire w_dff_A_43qxwe5n4_0;
	wire w_dff_A_lM4cQxuK8_0;
	wire w_dff_A_P02dXyHs2_0;
	wire w_dff_A_gPnPbhlk2_0;
	wire w_dff_A_pjPlahOv5_0;
	wire w_dff_A_sd4yuauN4_0;
	wire w_dff_A_pMGsOJDe5_0;
	wire w_dff_A_WIdxZpcC7_0;
	wire w_dff_A_7edUgzrp8_0;
	wire w_dff_A_eGFurfib8_0;
	wire w_dff_A_cnAalqim5_0;
	wire w_dff_A_s8XYea018_0;
	wire w_dff_A_SgELGMm62_0;
	wire w_dff_A_B5zaQhi98_1;
	wire w_dff_A_kw8rr8Nl7_0;
	wire w_dff_A_KYBBMnJJ6_0;
	wire w_dff_A_aHi9xvcF3_0;
	wire w_dff_A_roJLgMVP1_0;
	wire w_dff_A_3JDIISQ00_0;
	wire w_dff_A_1cM70qXy2_0;
	wire w_dff_A_SytAfQnO7_0;
	wire w_dff_A_oX47xxQO7_0;
	wire w_dff_A_Dl72Iv3P9_0;
	wire w_dff_A_R5giQd9G7_0;
	wire w_dff_A_RRJqQEfR2_0;
	wire w_dff_A_U31w5LeJ4_0;
	wire w_dff_A_wELXTeHb9_0;
	wire w_dff_A_McTbMLZN9_0;
	wire w_dff_A_XtRoVTfS9_0;
	wire w_dff_A_qYN43HMH4_0;
	wire w_dff_A_Zds1RHDK6_0;
	wire w_dff_A_2Ywc9JdV4_0;
	wire w_dff_A_sdLUWOH84_0;
	wire w_dff_A_cT8CFlQB5_0;
	wire w_dff_A_yJ8iasqj9_0;
	wire w_dff_A_VqBUACDa0_0;
	wire w_dff_A_2tZH7ec25_0;
	wire w_dff_A_skYbwueA9_0;
	wire w_dff_A_dr2oqWfh1_0;
	wire w_dff_A_BubwsMNS6_0;
	wire w_dff_A_wsRicFXl5_1;
	wire w_dff_A_lMMs7hJv3_0;
	wire w_dff_A_4tkXWEsA3_0;
	wire w_dff_A_DfnJXHkz0_0;
	wire w_dff_A_whsLhFcA3_0;
	wire w_dff_A_5OYSFGq80_0;
	wire w_dff_A_NnUSuJHM0_0;
	wire w_dff_A_7DCEQMkB8_0;
	wire w_dff_A_htuo9FSx2_0;
	wire w_dff_A_k97GJOOY8_0;
	wire w_dff_A_i9basHgR1_0;
	wire w_dff_A_Q1JFKpPs7_0;
	wire w_dff_A_ufocaaEK6_0;
	wire w_dff_A_WEbBZDyb9_0;
	wire w_dff_A_xRzkgRa43_0;
	wire w_dff_A_votJOWvl2_0;
	wire w_dff_A_BkKx0VBP8_0;
	wire w_dff_A_RHncwQeX4_0;
	wire w_dff_A_wK8pW0BO6_0;
	wire w_dff_A_IirWNDv19_0;
	wire w_dff_A_8WJSC0E14_0;
	wire w_dff_A_5CoaPKEU5_0;
	wire w_dff_A_xp6pNGAQ7_0;
	wire w_dff_A_VDwXIE4E5_0;
	wire w_dff_A_RO5r0N2e7_0;
	wire w_dff_A_6xRw4hWc7_0;
	wire w_dff_A_Ke9X6fvb2_0;
	wire w_dff_A_5wc4wnAA5_1;
	wire w_dff_A_2qNRjnX37_0;
	wire w_dff_A_c1bnQw2Z8_0;
	wire w_dff_A_86uySLNB7_0;
	wire w_dff_A_Q5jBzqUI3_0;
	wire w_dff_A_ueIqyRhO2_0;
	wire w_dff_A_S6ZOIxqh7_0;
	wire w_dff_A_Z4aiqFLt1_0;
	wire w_dff_A_Rnt4wmwV6_0;
	wire w_dff_A_Zjg07G7H0_0;
	wire w_dff_A_BAbJkfWu6_0;
	wire w_dff_A_N71oDIZv2_0;
	wire w_dff_A_gTcxvjPt7_0;
	wire w_dff_A_51cDu1Xn7_0;
	wire w_dff_A_UidG5YXB7_0;
	wire w_dff_A_7DMLheaJ2_0;
	wire w_dff_A_9Y6AxvSH9_0;
	wire w_dff_A_6WHusuzJ2_0;
	wire w_dff_A_63aDm5KU0_0;
	wire w_dff_A_Uct3V7rS5_0;
	wire w_dff_A_vStka29A1_0;
	wire w_dff_A_WHgyj6Ee1_0;
	wire w_dff_A_0RG0TIzb9_0;
	wire w_dff_A_kQjhXkOH3_0;
	wire w_dff_A_UaIFjqUD1_0;
	wire w_dff_A_S8sqmpI97_0;
	wire w_dff_A_4uwWC8Qm6_0;
	wire w_dff_A_iFcdHZpN8_1;
	wire w_dff_A_Mx1X726q8_0;
	wire w_dff_A_iPviCIs37_0;
	wire w_dff_A_7eI7kD5X9_0;
	wire w_dff_A_1pBmZcdT4_0;
	wire w_dff_A_ai3mTQ3z0_0;
	wire w_dff_A_kdGJnj6t1_0;
	wire w_dff_A_ECnEZZwQ9_0;
	wire w_dff_A_MMDbtLqk1_0;
	wire w_dff_A_ePWq3UBc0_0;
	wire w_dff_A_5oqBe5EH2_0;
	wire w_dff_A_6t9HqlM23_0;
	wire w_dff_A_07OyTkp68_0;
	wire w_dff_A_co11kp2N7_0;
	wire w_dff_A_bcLdXrdQ7_0;
	wire w_dff_A_9WLKyMj34_0;
	wire w_dff_A_nsxR5qEy0_0;
	wire w_dff_A_GWJhRBhU5_0;
	wire w_dff_A_iIfeIdj21_0;
	wire w_dff_A_0kLKVHac6_0;
	wire w_dff_A_3IeRq1wj9_0;
	wire w_dff_A_F1Xq0dlN9_0;
	wire w_dff_A_n7TI19Rg7_0;
	wire w_dff_A_bREk1lkZ4_0;
	wire w_dff_A_RGwOJmSC2_0;
	wire w_dff_A_Bztaqpdq6_0;
	wire w_dff_A_hOzwgkhi2_0;
	wire w_dff_A_6Sa7Xvf97_1;
	wire w_dff_A_Uf2jSV5b7_0;
	wire w_dff_A_rZfsHOJt3_0;
	wire w_dff_A_RpUp8Alr6_0;
	wire w_dff_A_SFJlVtsc9_0;
	wire w_dff_A_KehKZ3l47_0;
	wire w_dff_A_PzvtLay25_0;
	wire w_dff_A_210zCSDV5_0;
	wire w_dff_A_SZfDYcQl6_0;
	wire w_dff_A_RPdSk9mK4_0;
	wire w_dff_A_naZQSBVL9_0;
	wire w_dff_A_uetRDmOr3_0;
	wire w_dff_A_NBEnAyvh3_0;
	wire w_dff_A_VW0juebU2_0;
	wire w_dff_A_ts3Kubfk9_0;
	wire w_dff_A_id7yic8Z6_0;
	wire w_dff_A_TFTHJbxc8_0;
	wire w_dff_A_emAsT7vR0_0;
	wire w_dff_A_3ALw9M8d9_0;
	wire w_dff_A_KmpkTfpE0_0;
	wire w_dff_A_qfEDelqT2_0;
	wire w_dff_A_6BCkUk5Y0_0;
	wire w_dff_A_XMjGGtsr5_0;
	wire w_dff_A_hD3yCD5v0_0;
	wire w_dff_A_jNVRaYYi8_0;
	wire w_dff_A_l75UpMBg1_0;
	wire w_dff_A_6Aq8FD5u4_0;
	wire w_dff_A_aWb3Bder3_1;
	wire w_dff_A_37qidPkF0_0;
	wire w_dff_A_Q6fFJPZb4_0;
	wire w_dff_A_uRyH7K3K9_0;
	wire w_dff_A_4NRPImzl0_0;
	wire w_dff_A_BRWbNyB77_0;
	wire w_dff_A_XWy7JglP7_0;
	wire w_dff_A_61JnoIBW2_0;
	wire w_dff_A_ZCJvXGZe1_0;
	wire w_dff_A_1q4FCxbs0_0;
	wire w_dff_A_eA0dgkzs4_0;
	wire w_dff_A_YRIjOYI94_0;
	wire w_dff_A_zTNwIrWC7_0;
	wire w_dff_A_kmrbAwfV0_0;
	wire w_dff_A_Ox8EP8me8_0;
	wire w_dff_A_sndsVV9d8_0;
	wire w_dff_A_O5KbiIx65_0;
	wire w_dff_A_aLKeHqcp8_0;
	wire w_dff_A_nR60EwYh4_0;
	wire w_dff_A_RIjzj0jG8_0;
	wire w_dff_A_yVTjbZxL4_0;
	wire w_dff_A_lNo6GqT56_0;
	wire w_dff_A_qYjj9DpR2_0;
	wire w_dff_A_n629pjA98_0;
	wire w_dff_A_dSWu2JMH3_0;
	wire w_dff_A_IuCpVn6p1_0;
	wire w_dff_A_24FkzvG86_0;
	wire w_dff_A_EJSBV4R46_2;
	wire w_dff_A_TIELi39v9_0;
	wire w_dff_A_GVghg9bM9_0;
	wire w_dff_A_SDmsdrjL1_0;
	wire w_dff_A_aKCiX8WE3_0;
	wire w_dff_A_Pwk7GOeq1_0;
	wire w_dff_A_ttDfJGRe8_0;
	wire w_dff_A_o9ORt5Of5_0;
	wire w_dff_A_PTjsbeIh6_0;
	wire w_dff_A_Ke32ivLL0_0;
	wire w_dff_A_DOM2kqXq7_0;
	wire w_dff_A_MQZhC69F6_0;
	wire w_dff_A_HalNvWIm0_0;
	wire w_dff_A_Ggisu0AC2_0;
	wire w_dff_A_FF7QhOBt5_0;
	wire w_dff_A_4oIQ4CII8_0;
	wire w_dff_A_5o70XSRu5_0;
	wire w_dff_A_6NclDxdl4_0;
	wire w_dff_A_x1pekYJs3_0;
	wire w_dff_A_NtouRkLw1_0;
	wire w_dff_A_kpY8J51a4_0;
	wire w_dff_A_6Vpx65ZK3_0;
	wire w_dff_A_TS2hjwmc2_0;
	wire w_dff_A_ZGNjP5nh3_0;
	wire w_dff_A_pIyMq1T61_0;
	wire w_dff_A_psfa3IAA7_0;
	wire w_dff_A_Qz3g3XdO7_0;
	wire w_dff_A_C0wtGoAE3_1;
	wire w_dff_A_2h0KxOym5_0;
	wire w_dff_A_OWrkQTk52_0;
	wire w_dff_A_AlY58BUz8_0;
	wire w_dff_A_ht2SxEAa9_0;
	wire w_dff_A_G8akYSOr8_0;
	wire w_dff_A_4QQeJKHz5_0;
	wire w_dff_A_7OrlUbxO2_0;
	wire w_dff_A_XK02slre7_0;
	wire w_dff_A_CTDGqpaF6_0;
	wire w_dff_A_KzwYXyOC3_0;
	wire w_dff_A_7GQrzYxo1_0;
	wire w_dff_A_4azZmAGj3_0;
	wire w_dff_A_VIUP5geH9_0;
	wire w_dff_A_a1kw8kaT5_0;
	wire w_dff_A_qrAtofiT7_0;
	wire w_dff_A_1eeGagY18_0;
	wire w_dff_A_OE1VORvO6_0;
	wire w_dff_A_RkzhPTIv2_0;
	wire w_dff_A_tEab5lgN4_0;
	wire w_dff_A_tMXXNwq55_0;
	wire w_dff_A_wRTpQvsx3_0;
	wire w_dff_A_Wo3NGruI6_0;
	wire w_dff_A_UwlsSxj38_0;
	wire w_dff_A_HRvzKhzK6_0;
	wire w_dff_A_7FtUQ8he6_0;
	wire w_dff_A_e1gUUK8D8_0;
	wire w_dff_A_ZcBak8Wz0_1;
	wire w_dff_A_d6Zmd3nD4_0;
	wire w_dff_A_V6mA00sq6_0;
	wire w_dff_A_WUdKXxqu6_0;
	wire w_dff_A_53xY64Mt6_0;
	wire w_dff_A_vnmyTlvZ1_0;
	wire w_dff_A_T4Ly5fbj3_0;
	wire w_dff_A_9MWoWyTM4_0;
	wire w_dff_A_oHiwbgD08_0;
	wire w_dff_A_66mEnOOU3_0;
	wire w_dff_A_7p4kKu1b7_0;
	wire w_dff_A_LY0ED1MY8_0;
	wire w_dff_A_P5siTwNL5_0;
	wire w_dff_A_GJIPEppz7_0;
	wire w_dff_A_OE62B7CQ3_0;
	wire w_dff_A_XJidZEOv9_0;
	wire w_dff_A_TGSrF0Bo2_0;
	wire w_dff_A_wBHJ4t5C7_0;
	wire w_dff_A_QUJtWDbP0_0;
	wire w_dff_A_WrGC2sDE4_0;
	wire w_dff_A_CeFX0CnR4_0;
	wire w_dff_A_75vGWjBU8_0;
	wire w_dff_A_1S16eqBq7_0;
	wire w_dff_A_cry6awpr7_0;
	wire w_dff_A_Ni5dg4iN7_0;
	wire w_dff_A_IRJ1jwDa5_0;
	wire w_dff_A_q7VcqtXf2_0;
	wire w_dff_A_11gMwd6c1_1;
	wire w_dff_A_DgSuzRmG0_0;
	wire w_dff_A_w0iVHi3J9_0;
	wire w_dff_A_GT5xiU5F3_0;
	wire w_dff_A_MyiXWURi6_0;
	wire w_dff_A_YzaojHkK1_0;
	wire w_dff_A_HVNic8zf5_0;
	wire w_dff_A_oYJ2F1f43_0;
	wire w_dff_A_E2hWJkdu2_0;
	wire w_dff_A_4kt8yL2l0_0;
	wire w_dff_A_idHBsHLM5_0;
	wire w_dff_A_5eWmLYEj9_0;
	wire w_dff_A_HEnZeIni7_0;
	wire w_dff_A_iJ242T1M6_0;
	wire w_dff_A_sYliSE2D2_0;
	wire w_dff_A_8csViICh1_0;
	wire w_dff_A_ucVAyJuO7_0;
	wire w_dff_A_uEBK0OSV7_0;
	wire w_dff_A_eDAbYZIk2_0;
	wire w_dff_A_EUz0yJH81_0;
	wire w_dff_A_X6D4NQWF5_0;
	wire w_dff_A_Jq7iJYdi3_0;
	wire w_dff_A_Yjc51a5W8_0;
	wire w_dff_A_kWey6ZCY1_0;
	wire w_dff_A_aIATRkWV5_0;
	wire w_dff_A_JnfrM3eY5_0;
	wire w_dff_A_b0kcHwIx9_0;
	wire w_dff_A_Yhp1kSkX5_1;
	wire w_dff_A_4755lNO00_0;
	wire w_dff_A_eJ6AB6SP3_0;
	wire w_dff_A_jIxzoZVo2_0;
	wire w_dff_A_31G2phhd7_0;
	wire w_dff_A_DhUeKY8a0_0;
	wire w_dff_A_FADsnsv75_0;
	wire w_dff_A_nVlY46uf7_0;
	wire w_dff_A_2P1Z4ldK9_0;
	wire w_dff_A_HjlgrXy65_0;
	wire w_dff_A_IR4yVBWR5_0;
	wire w_dff_A_TwUAFyaG0_0;
	wire w_dff_A_hp0ZPgsW7_0;
	wire w_dff_A_CzJUzp0U8_0;
	wire w_dff_A_y3DPTehL1_0;
	wire w_dff_A_8LL1JtOT2_0;
	wire w_dff_A_nKeFnkHY4_0;
	wire w_dff_A_JzsBgQVP9_0;
	wire w_dff_A_aeXoUm8T5_0;
	wire w_dff_A_oONrYMeZ5_0;
	wire w_dff_A_mfi7YCDQ4_0;
	wire w_dff_A_6S7CztCU1_0;
	wire w_dff_A_exCZ1ihX1_0;
	wire w_dff_A_rskND1Rz4_0;
	wire w_dff_A_uin5GKpW9_0;
	wire w_dff_A_JRV5moa65_0;
	wire w_dff_A_gJJjhMvl0_0;
	wire w_dff_A_yO5mAeIh3_2;
	wire w_dff_A_RjRfhNgA7_0;
	wire w_dff_A_8GFNQy1I5_0;
	wire w_dff_A_wVLADo1z7_0;
	wire w_dff_A_8q1uKPao5_0;
	wire w_dff_A_Ks2GVdeT5_0;
	wire w_dff_A_1a5rZWHF6_0;
	wire w_dff_A_iswYPrAg8_0;
	wire w_dff_A_jzWxOYOT5_0;
	wire w_dff_A_nPgekng83_0;
	wire w_dff_A_tEMX9oRN9_0;
	wire w_dff_A_TI09GShc2_0;
	wire w_dff_A_PL6kwVX03_0;
	wire w_dff_A_WCvWDdPG7_0;
	wire w_dff_A_1OhX25aX6_0;
	wire w_dff_A_rNtBoynd0_0;
	wire w_dff_A_3D7ljEMI2_0;
	wire w_dff_A_LvzGJYUi9_0;
	wire w_dff_A_eIkqh5s40_0;
	wire w_dff_A_JbH58zZu9_0;
	wire w_dff_A_kGzAnvD47_0;
	wire w_dff_A_jOtCDVt65_0;
	wire w_dff_A_utL2w7AN0_0;
	wire w_dff_A_m7qFaZLq5_0;
	wire w_dff_A_gVm80JcI8_0;
	wire w_dff_A_aHFy5ff96_0;
	wire w_dff_A_DSGeUlm45_0;
	wire w_dff_A_exStBqkQ5_2;
	wire w_dff_A_wuWBSvkX1_0;
	wire w_dff_A_sWU2c14H7_0;
	wire w_dff_A_ifKrietX1_0;
	wire w_dff_A_CBMKM7pt5_0;
	wire w_dff_A_cKNcyqqd6_0;
	wire w_dff_A_YzAeThHe1_0;
	wire w_dff_A_XCg6C0rR1_0;
	wire w_dff_A_Y2cdZ01X2_0;
	wire w_dff_A_P4Ckavm71_0;
	wire w_dff_A_IPLI65ef5_0;
	wire w_dff_A_abzK3VH78_0;
	wire w_dff_A_LPDUQsau6_0;
	wire w_dff_A_0J3DAQz32_0;
	wire w_dff_A_3xCap0Mj8_0;
	wire w_dff_A_lBXDLFVS9_0;
	wire w_dff_A_CQ46U00c2_0;
	wire w_dff_A_Y7L5ftOy9_0;
	wire w_dff_A_VtWdf7Dz6_0;
	wire w_dff_A_aaYvH3vo7_0;
	wire w_dff_A_etZ9ZXnN3_0;
	wire w_dff_A_fqB1lQAs3_0;
	wire w_dff_A_SF599VBN1_0;
	wire w_dff_A_vDBYVT3T9_0;
	wire w_dff_A_IXVxdoHg8_0;
	wire w_dff_A_LER4ChrA4_0;
	wire w_dff_A_TqMoaJk03_2;
	wire w_dff_A_wX0tWmqN4_0;
	wire w_dff_A_tax51nS43_0;
	wire w_dff_A_iHRLFPRF5_0;
	wire w_dff_A_rOfsVARI3_0;
	wire w_dff_A_xy8qDcDh8_0;
	wire w_dff_A_kwydTDlu0_0;
	wire w_dff_A_KZK8FBHa9_0;
	wire w_dff_A_BKOrgFgS3_0;
	wire w_dff_A_K8oGeYbo5_0;
	wire w_dff_A_F0YoVC4q5_0;
	wire w_dff_A_Eyrjf1Aa7_0;
	wire w_dff_A_dvyRq3G07_0;
	wire w_dff_A_CCSbbp4O5_0;
	wire w_dff_A_kpI7ahMl0_0;
	wire w_dff_A_0f30fpFz1_0;
	wire w_dff_A_Rw0Qhv6R7_0;
	wire w_dff_A_8cxXHgb43_0;
	wire w_dff_A_GTWRWzMJ1_0;
	wire w_dff_A_kNfBVaqN5_0;
	wire w_dff_A_jYZljm1K3_0;
	wire w_dff_A_tN44kCaU6_0;
	wire w_dff_A_7xzm6zBw3_0;
	wire w_dff_A_Y80qzSBW2_0;
	wire w_dff_A_jTF1pupG7_0;
	wire w_dff_A_9CvpmEld7_0;
	wire w_dff_A_X7F1HKYL4_1;
	wire w_dff_A_uolmimfa7_0;
	wire w_dff_A_N9AqXNZj4_0;
	wire w_dff_A_eYsRJPwR2_0;
	wire w_dff_A_ullLoJye8_0;
	wire w_dff_A_W5SJSUET1_0;
	wire w_dff_A_oN66D3234_0;
	wire w_dff_A_njo6NJt84_0;
	wire w_dff_A_TwGOlEDQ3_0;
	wire w_dff_A_05yKt7xE7_0;
	wire w_dff_A_nWhjeQUn1_0;
	wire w_dff_A_0k5yljyq4_0;
	wire w_dff_A_joeKOMa00_0;
	wire w_dff_A_1W5ct2YD4_0;
	wire w_dff_A_jgrFbjJM0_0;
	wire w_dff_A_2svmAVov8_0;
	wire w_dff_A_fymio6HD2_0;
	wire w_dff_A_2y5WtJwj2_0;
	wire w_dff_A_rapHXvm16_0;
	wire w_dff_A_UV1gxB2A0_0;
	wire w_dff_A_Qb1y4N3U2_0;
	wire w_dff_A_yE9pNrb00_0;
	wire w_dff_A_bC9yovAL8_0;
	wire w_dff_A_SRGktNGU7_0;
	wire w_dff_A_gGXfGeiv4_0;
	wire w_dff_A_HyNuPhMA7_0;
	wire w_dff_A_TKuoKSCW6_1;
	wire w_dff_A_kZTx9DQi5_0;
	wire w_dff_A_XAMLZK897_0;
	wire w_dff_A_Q0KDuIQD5_0;
	wire w_dff_A_7HskTq8i1_0;
	wire w_dff_A_p0dUaPYs2_0;
	wire w_dff_A_dPB2mbSR9_0;
	wire w_dff_A_6DoRZaxf7_0;
	wire w_dff_A_KtB1YAE87_0;
	wire w_dff_A_8r1zBTMk4_0;
	wire w_dff_A_ZvjI8cll1_0;
	wire w_dff_A_V4Vrc5Gq4_0;
	wire w_dff_A_oZ86eTmZ4_0;
	wire w_dff_A_lCenTC5v2_0;
	wire w_dff_A_m0rGnH2a3_0;
	wire w_dff_A_ZuHOqMvl8_0;
	wire w_dff_A_PaIkXcRc8_0;
	wire w_dff_A_XiLAzX2v0_0;
	wire w_dff_A_W3C6j8an3_0;
	wire w_dff_A_oTAmvKeV6_0;
	wire w_dff_A_Fdx07G1M3_0;
	wire w_dff_A_pP7Lof4f8_0;
	wire w_dff_A_TUK6L97F4_0;
	wire w_dff_A_1oJ631Nj6_0;
	wire w_dff_A_UBYY5Txl7_0;
	wire w_dff_A_KoPsLqfG6_0;
	wire w_dff_A_nl539tiC9_0;
	wire w_dff_A_lxqjMQZT1_0;
	wire w_dff_A_K6wpGJWd3_1;
	wire w_dff_A_svZrmNcT1_0;
	wire w_dff_A_9glUybEI4_0;
	wire w_dff_A_YCiEjFmB0_0;
	wire w_dff_A_x8QmaDmv5_0;
	wire w_dff_A_h1tcUOTL7_0;
	wire w_dff_A_kdTQgwsB1_0;
	wire w_dff_A_DRN1mrgV8_0;
	wire w_dff_A_nmj3gwya5_0;
	wire w_dff_A_VGMn8EBD2_0;
	wire w_dff_A_4vSHMUWt7_0;
	wire w_dff_A_ZVqvWqnY1_0;
	wire w_dff_A_AizFZySo8_0;
	wire w_dff_A_qRzsO6K48_0;
	wire w_dff_A_84LrDuoC8_0;
	wire w_dff_A_pcbL62Am2_0;
	wire w_dff_A_3Z9WgCgd0_0;
	wire w_dff_A_BYPa2LIP9_0;
	wire w_dff_A_kmWpum7a4_0;
	wire w_dff_A_HnPGqevu0_0;
	wire w_dff_A_bdGU1SC37_0;
	wire w_dff_A_tjOBBkxe5_0;
	wire w_dff_A_iloMe4C68_0;
	wire w_dff_A_8iAIhAUm1_0;
	wire w_dff_A_veLfxbv81_0;
	wire w_dff_A_5BeclRPt5_0;
	wire w_dff_A_rldhZ6m63_0;
	wire w_dff_A_5F3MKZkd9_0;
	wire w_dff_A_7l1xJPxg8_1;
	wire w_dff_A_3BtInpLT1_0;
	wire w_dff_A_Dxpbdw9F3_0;
	wire w_dff_A_BSbxc1X46_0;
	wire w_dff_A_J6W2mOVq3_0;
	wire w_dff_A_x0c4WEPB3_0;
	wire w_dff_A_Btim2EmK9_0;
	wire w_dff_A_Rm9xGRml6_0;
	wire w_dff_A_3KwY0D8P4_0;
	wire w_dff_A_Bj9mIC140_0;
	wire w_dff_A_A8tdTRLX4_0;
	wire w_dff_A_l0UNyCUa6_0;
	wire w_dff_A_VP4EwxVk1_0;
	wire w_dff_A_di23gKqp9_0;
	wire w_dff_A_y8tQFYT21_0;
	wire w_dff_A_LvUPQXoD7_0;
	wire w_dff_A_ZqL753SO0_0;
	wire w_dff_A_0ekW3pl70_0;
	wire w_dff_A_u4EQxJVr5_0;
	wire w_dff_A_C7UhureO5_0;
	wire w_dff_A_6yTXDHJQ2_0;
	wire w_dff_A_8uEaIVUC2_0;
	wire w_dff_A_3grzfB785_0;
	wire w_dff_A_UQLSSYID3_0;
	wire w_dff_A_qP045btj2_0;
	wire w_dff_A_NGwoo8C80_0;
	wire w_dff_A_MskSZxQV0_0;
	wire w_dff_A_7fWrvqMH1_0;
	wire w_dff_A_2dIO24Jj4_1;
	wire w_dff_A_JZFRN4bg2_0;
	wire w_dff_A_hBEiWT7E1_0;
	wire w_dff_A_05KovSCo7_0;
	wire w_dff_A_C4E5evo04_0;
	wire w_dff_A_TuXHF67f6_0;
	wire w_dff_A_jmsVYBMe5_0;
	wire w_dff_A_WkZyNZYE1_0;
	wire w_dff_A_GKzmejjr5_0;
	wire w_dff_A_3yjqPXRu3_0;
	wire w_dff_A_wa3LCTQR6_0;
	wire w_dff_A_Op8uBwhR6_0;
	wire w_dff_A_b3ZWdLmK3_0;
	wire w_dff_A_y1CmGoI21_0;
	wire w_dff_A_XN3l33IS4_0;
	wire w_dff_A_trz5VlK68_0;
	wire w_dff_A_n7EYXIdz7_0;
	wire w_dff_A_9QOtFYE66_0;
	wire w_dff_A_L7AYeuKv3_0;
	wire w_dff_A_RBeo2VRm9_0;
	wire w_dff_A_J3hIDXpq7_0;
	wire w_dff_A_i7wMwufA7_0;
	wire w_dff_A_xPbSj6o89_0;
	wire w_dff_A_QmYk2Xnp1_0;
	wire w_dff_A_nGDtdNpn7_0;
	wire w_dff_A_BvFAkxhV2_0;
	wire w_dff_A_1jMbOY4l0_0;
	wire w_dff_A_H6KQgU2i4_0;
	wire w_dff_A_lRm1ZvdP4_1;
	wire w_dff_A_fidZ2kb52_0;
	wire w_dff_A_kInfo4lD6_0;
	wire w_dff_A_KMjoz2Vx1_0;
	wire w_dff_A_JmxLcGv83_0;
	wire w_dff_A_ui9jUVXr9_0;
	wire w_dff_A_DN2FgIAM8_0;
	wire w_dff_A_RZdDCcOz3_0;
	wire w_dff_A_hbdCbXy21_0;
	wire w_dff_A_M8Z17VPj6_0;
	wire w_dff_A_SYOPsecX8_0;
	wire w_dff_A_XKu1PCda4_0;
	wire w_dff_A_8OmycR1V2_0;
	wire w_dff_A_TxCas6dB8_0;
	wire w_dff_A_N0gzojVw9_0;
	wire w_dff_A_kh8NhTMo8_0;
	wire w_dff_A_rwR7Xe3H1_0;
	wire w_dff_A_yI90uVPX5_0;
	wire w_dff_A_b6jvVOdI6_0;
	wire w_dff_A_dhe6uz7V4_0;
	wire w_dff_A_H3gmHbEy4_0;
	wire w_dff_A_yMtsPDPo7_0;
	wire w_dff_A_DoxEIe4l3_0;
	wire w_dff_A_yxT7KSTO6_0;
	wire w_dff_A_0fe5NYxD3_0;
	wire w_dff_A_zdwmYmkE7_0;
	wire w_dff_A_SsdBe5ct7_0;
	wire w_dff_A_jKZjYG0l5_0;
	wire w_dff_A_VRuQeKNr1_1;
	wire w_dff_A_9dRG4BhY4_0;
	wire w_dff_A_kCDmO6Y39_0;
	wire w_dff_A_iq4yiSHG1_0;
	wire w_dff_A_pd17vWUi1_0;
	wire w_dff_A_rLhQvUlX8_0;
	wire w_dff_A_d4qsAZCa0_0;
	wire w_dff_A_oP7jJvD27_0;
	wire w_dff_A_J5JPQTd18_0;
	wire w_dff_A_Z0qnVw5v6_0;
	wire w_dff_A_HeVKRGNY5_0;
	wire w_dff_A_jLrRvOig5_0;
	wire w_dff_A_0yv65RKl1_0;
	wire w_dff_A_vflgsjhW7_0;
	wire w_dff_A_sP3kGwxG9_0;
	wire w_dff_A_CR8lprwe6_0;
	wire w_dff_A_fYFJzdR15_0;
	wire w_dff_A_OZ7OF0x22_0;
	wire w_dff_A_ic9h4GPH4_0;
	wire w_dff_A_dmeUYhbd6_0;
	wire w_dff_A_ZTWK0T7B8_0;
	wire w_dff_A_DKGHJwYl9_0;
	wire w_dff_A_xEoJ4PH74_0;
	wire w_dff_A_7xLa8arg7_0;
	wire w_dff_A_cuiR6SJb7_0;
	wire w_dff_A_w7kXvGwR3_0;
	wire w_dff_A_FWpDfBEp2_0;
	wire w_dff_A_gg3PgASV0_2;
	wire w_dff_A_aR4I8e2K2_0;
	wire w_dff_A_Ie7QgcyS2_0;
	wire w_dff_A_CRtd59Gh5_0;
	wire w_dff_A_8nY0sgGo7_0;
	wire w_dff_A_AfSjFJ1y3_0;
	wire w_dff_A_b1p62XoN6_0;
	wire w_dff_A_0t3v89To7_0;
	wire w_dff_A_aWMnwsv82_0;
	wire w_dff_A_IPp4htNW4_0;
	wire w_dff_A_ayhWAWw79_0;
	wire w_dff_A_iFtYWRGX8_0;
	wire w_dff_A_nfQuiThr9_0;
	wire w_dff_A_r03sexoY6_0;
	wire w_dff_A_pkSq7Xgv3_0;
	wire w_dff_A_9Va8nnXD6_0;
	wire w_dff_A_MdlN1K6W7_0;
	wire w_dff_A_27y9WcvV6_0;
	wire w_dff_A_Im5N1SSr6_0;
	wire w_dff_A_1Rp6iL4m3_0;
	wire w_dff_A_iYkgZ1bF0_0;
	wire w_dff_A_ZNMqHimi9_0;
	wire w_dff_A_RHpnLfV68_0;
	wire w_dff_A_uPLTWHaV8_0;
	wire w_dff_A_5Eeh20Wr7_0;
	wire w_dff_A_yuNhCNJz3_2;
	wire w_dff_A_WvrD45bc8_0;
	wire w_dff_A_5H6WQno93_0;
	wire w_dff_A_ivQAUMxH8_0;
	wire w_dff_A_bQjt1a1G0_0;
	wire w_dff_A_GSt8cXHT4_0;
	wire w_dff_A_uMkgMiZf3_0;
	wire w_dff_A_MzDnONN47_0;
	wire w_dff_A_a6Pot5A36_0;
	wire w_dff_A_KAZbcTXc0_0;
	wire w_dff_A_5MWOhsnT4_0;
	wire w_dff_A_so1wG80E3_0;
	wire w_dff_A_47Tc0aO99_0;
	wire w_dff_A_DiPs3LSX3_0;
	wire w_dff_A_fzQQPQQr6_0;
	wire w_dff_A_NbxfKrOW2_0;
	wire w_dff_A_gB4h6JBI1_0;
	wire w_dff_A_cEwu8iz73_0;
	wire w_dff_A_L7zAtZmE4_0;
	wire w_dff_A_dkg99LSj6_0;
	wire w_dff_A_qjWZ4vUH3_0;
	wire w_dff_A_vTcdfKT48_0;
	wire w_dff_A_jwgxTFxz7_0;
	wire w_dff_A_RYfOJeG11_0;
	wire w_dff_A_EFLsrP0x4_0;
	wire w_dff_A_m703jvyh6_0;
	wire w_dff_A_kHDc557D8_1;
	wire w_dff_A_tHQUoPYV4_0;
	wire w_dff_A_JWnk32uO1_0;
	wire w_dff_A_6yfjsOLV6_0;
	wire w_dff_A_RE9UljRM3_0;
	wire w_dff_A_xPAN24Gg7_0;
	wire w_dff_A_fRXrni0X7_0;
	wire w_dff_A_JD4p8yJT9_0;
	wire w_dff_A_UkgFFqRz4_0;
	wire w_dff_A_2fkSJ1ds0_0;
	wire w_dff_A_sfopnZ7L9_0;
	wire w_dff_A_mDvVVJk68_0;
	wire w_dff_A_OxXF5fDc3_0;
	wire w_dff_A_68sPz6aE4_0;
	wire w_dff_A_poE1YTcD5_0;
	wire w_dff_A_JsQkrAfx1_0;
	wire w_dff_A_U9Ahwjuy5_0;
	wire w_dff_A_JsEbNU8Q7_0;
	wire w_dff_A_9kUhDqqt2_0;
	wire w_dff_A_AFMP7DaI7_0;
	wire w_dff_A_SCLIygbe4_0;
	wire w_dff_A_pEaPMiuy1_0;
	wire w_dff_A_bEsuk1930_0;
	wire w_dff_A_TcJnLONY7_0;
	wire w_dff_A_UD2G7XuA8_0;
	wire w_dff_A_r7uy8L3S1_0;
	wire w_dff_A_rOjpEODb0_0;
	wire w_dff_A_lzxLPuzi5_0;
	wire w_dff_A_GL80qaD07_1;
	wire w_dff_A_kWakDpog6_0;
	wire w_dff_A_Vo1PcdKq3_0;
	wire w_dff_A_lR0QA30s2_0;
	wire w_dff_A_vGJS5vWd8_0;
	wire w_dff_A_ZHIt9AMD1_0;
	wire w_dff_A_qEYSLesI6_0;
	wire w_dff_A_23jqGqgc6_0;
	wire w_dff_A_40ITOBCG8_0;
	wire w_dff_A_RhIRWPRt6_0;
	wire w_dff_A_9rvfiyRD6_0;
	wire w_dff_A_3yITJfY47_0;
	wire w_dff_A_nHpMnFic5_0;
	wire w_dff_A_IKOeYurh5_0;
	wire w_dff_A_blXyaCrD7_0;
	wire w_dff_A_dL4X1qm12_0;
	wire w_dff_A_j9OeQzmB7_0;
	wire w_dff_A_OQoWEMgG1_0;
	wire w_dff_A_V5NDIerF7_0;
	wire w_dff_A_TKmN7Ysz0_0;
	wire w_dff_A_2k7ESiSz6_0;
	wire w_dff_A_whASYpX52_0;
	wire w_dff_A_sWXcdNLY3_0;
	wire w_dff_A_7PvL0IXM7_0;
	wire w_dff_A_d60VyGJu2_0;
	wire w_dff_A_VZlvfsq45_0;
	wire w_dff_A_JhRE7CG32_0;
	wire w_dff_A_I4saYtgB8_0;
	wire w_dff_A_DSogMvSP0_1;
	wire w_dff_A_C4gJVj634_0;
	wire w_dff_A_dx9VHOy94_0;
	wire w_dff_A_CGBEwkDY2_0;
	wire w_dff_A_m0ldYnrN3_0;
	wire w_dff_A_tOL6xVWu9_0;
	wire w_dff_A_rpw6DQMo7_0;
	wire w_dff_A_857cWHrX9_0;
	wire w_dff_A_Xic6uetH5_0;
	wire w_dff_A_ZNXKv3sL5_0;
	wire w_dff_A_OX3jQDPM7_0;
	wire w_dff_A_Y4R5hK3X2_0;
	wire w_dff_A_YECpAPEX6_0;
	wire w_dff_A_Z5tanN8y8_0;
	wire w_dff_A_SEbXML8t1_0;
	wire w_dff_A_kiILA36z4_0;
	wire w_dff_A_dduyINLq4_0;
	wire w_dff_A_yh9MxF8o9_0;
	wire w_dff_A_fSJicmTz9_0;
	wire w_dff_A_hU4Mgo6l2_0;
	wire w_dff_A_Ecj0khgj6_0;
	wire w_dff_A_YdIz7Gjr0_0;
	wire w_dff_A_d4UBJGGz6_0;
	wire w_dff_A_lBds5kpI7_0;
	wire w_dff_A_oyPXV0ai1_0;
	wire w_dff_A_sHd6jvbM1_0;
	wire w_dff_A_e3O8wnjN1_0;
	wire w_dff_A_13metCxG7_0;
	wire w_dff_A_icCkjrtN9_1;
	wire w_dff_A_19iUWqEI7_0;
	wire w_dff_A_JnRpjgjB5_0;
	wire w_dff_A_Rawa0EVo0_0;
	wire w_dff_A_zZsP4AEc1_0;
	wire w_dff_A_RbIpnAqe4_0;
	wire w_dff_A_BTU9xes56_0;
	wire w_dff_A_y2nK58US2_0;
	wire w_dff_A_O8WNIf8A1_0;
	wire w_dff_A_OCtkCjLF7_0;
	wire w_dff_A_M7MSGmvC2_0;
	wire w_dff_A_Yn9lY7Bv8_0;
	wire w_dff_A_fvxQu5hT4_0;
	wire w_dff_A_HKulKoja1_0;
	wire w_dff_A_tBJlzOuX6_0;
	wire w_dff_A_xHdlANjI3_0;
	wire w_dff_A_KhBIWZB19_0;
	wire w_dff_A_XHIJn5oW8_0;
	wire w_dff_A_BWzNvPEo9_0;
	wire w_dff_A_mK02EGtM5_0;
	wire w_dff_A_AAp6yyvL6_0;
	wire w_dff_A_JVPlbqT78_0;
	wire w_dff_A_b2uXC3is0_0;
	wire w_dff_A_YnxnsBmf6_0;
	wire w_dff_A_EjOPzYaz8_0;
	wire w_dff_A_Q5HRcTLO0_0;
	wire w_dff_A_NSEEvzcA4_0;
	wire w_dff_A_Juz5QEP89_0;
	wire w_dff_A_fys1SLwP5_1;
	wire w_dff_A_03AV6cOF7_0;
	wire w_dff_A_YNtWI2A51_0;
	wire w_dff_A_n0hVXxYY0_0;
	wire w_dff_A_6oHBMrwI7_0;
	wire w_dff_A_yViWC5cv3_0;
	wire w_dff_A_iSnmxgFp8_0;
	wire w_dff_A_yUeI6QGd8_0;
	wire w_dff_A_f5lYtiih3_0;
	wire w_dff_A_XCjfE83U0_0;
	wire w_dff_A_jttIpTwo5_0;
	wire w_dff_A_sQOSlP209_0;
	wire w_dff_A_ZaPRMZIa9_0;
	wire w_dff_A_dhrTnkyF2_0;
	wire w_dff_A_mlgafr6e8_0;
	wire w_dff_A_TI1mhfOY5_0;
	wire w_dff_A_eeH0C1ff1_0;
	wire w_dff_A_Tie7n15P6_0;
	wire w_dff_A_zHTmS7JN2_0;
	wire w_dff_A_JawBmFkl7_0;
	wire w_dff_A_nV7evQ6t1_0;
	wire w_dff_A_m7gYe2MG0_0;
	wire w_dff_A_hh9qEkVP6_0;
	wire w_dff_A_wvsdtkKl5_0;
	wire w_dff_A_vWk6R8zK2_0;
	wire w_dff_A_q1qOcbL21_0;
	wire w_dff_A_pjZozWlJ0_0;
	wire w_dff_A_kqgBN8412_0;
	wire w_dff_A_ugDvOh8h3_1;
	wire w_dff_A_hsZh9E3t1_0;
	wire w_dff_A_Ic0JfziH3_0;
	wire w_dff_A_bueculMr9_0;
	wire w_dff_A_iVmqxflh9_0;
	wire w_dff_A_zx7i1Ip78_0;
	wire w_dff_A_vqDgRTU94_0;
	wire w_dff_A_uYPb1Vht7_0;
	wire w_dff_A_hg3tWgNL8_0;
	wire w_dff_A_nQHuPJJa7_0;
	wire w_dff_A_KerKxsGh9_0;
	wire w_dff_A_GvDcWhrR9_0;
	wire w_dff_A_HALWxpLy7_0;
	wire w_dff_A_SD9aFa6x9_0;
	wire w_dff_A_LVOW0u2p2_0;
	wire w_dff_A_akyrYSbX9_0;
	wire w_dff_A_nGWzfI9f7_0;
	wire w_dff_A_J3WM7dtJ3_0;
	wire w_dff_A_RHOYpTgT5_0;
	wire w_dff_A_oo7IHECP7_0;
	wire w_dff_A_ydeQ5ayO5_0;
	wire w_dff_A_hZYUJVo60_0;
	wire w_dff_A_EsKHFbn93_0;
	wire w_dff_A_ssxZdoPJ9_0;
	wire w_dff_A_7X0MkftL8_0;
	wire w_dff_A_YtbrXaaO6_0;
	wire w_dff_A_f5apguHw2_0;
	wire w_dff_A_1oUSV6XM4_2;
	wire w_dff_A_nC0NXBua2_0;
	wire w_dff_A_ZQbu3un66_0;
	wire w_dff_A_CXKX5Dup2_0;
	wire w_dff_A_BKwKrpvP4_0;
	wire w_dff_A_4QXByxUV8_0;
	wire w_dff_A_BQEhQaQ47_0;
	wire w_dff_A_TZB0iEli7_0;
	wire w_dff_A_0nHBNFlf5_0;
	wire w_dff_A_8DkTLxmb9_0;
	wire w_dff_A_ufmbZPiW9_0;
	wire w_dff_A_njwkmYS01_0;
	wire w_dff_A_WANDuyqQ2_0;
	wire w_dff_A_zNyzGZ896_0;
	wire w_dff_A_iSUqzAb20_0;
	wire w_dff_A_1hIRuFMn4_0;
	wire w_dff_A_kirutSCW2_0;
	wire w_dff_A_XnZSXl2U4_0;
	wire w_dff_A_qReVuPGl6_0;
	wire w_dff_A_zOtnA8He2_0;
	wire w_dff_A_Bi5hURtT2_0;
	wire w_dff_A_9VEz5i4k0_0;
	wire w_dff_A_LQbAxgAT1_0;
	wire w_dff_A_QGLXUlOm7_0;
	wire w_dff_A_Z3ftPUiG7_2;
	wire w_dff_A_zrVz5la56_0;
	wire w_dff_A_bCStDZfy2_0;
	wire w_dff_A_Ra7FCRXm2_0;
	wire w_dff_A_7n7Jb1vb1_0;
	wire w_dff_A_lUVkydTd9_0;
	wire w_dff_A_s24DJm9f7_0;
	wire w_dff_A_HpQvrubS3_0;
	wire w_dff_A_8Ao1vih75_0;
	wire w_dff_A_EWiY3Q5b1_0;
	wire w_dff_A_odf1XUXH9_0;
	wire w_dff_A_i4hdn9WJ7_0;
	wire w_dff_A_VNFg8XVd8_0;
	wire w_dff_A_gRbGBBeR8_0;
	wire w_dff_A_PXEivqZw7_0;
	wire w_dff_A_FudwoYCP4_0;
	wire w_dff_A_myuVa9p54_0;
	wire w_dff_A_NO1QizLD5_0;
	wire w_dff_A_NwC58MJ06_0;
	wire w_dff_A_LpCHxOlX5_0;
	wire w_dff_A_QWjWVOXW1_0;
	wire w_dff_A_jHdqJ5y54_0;
	wire w_dff_A_Y7kUXdtv0_0;
	wire w_dff_A_O29KIGL57_0;
	wire w_dff_A_3bTGddH80_2;
	wire w_dff_A_HCmD40Ox0_0;
	wire w_dff_A_ds1O7zvS3_0;
	wire w_dff_A_8pNByWip8_0;
	wire w_dff_A_KYO7g1q22_0;
	wire w_dff_A_8cNRoMUS5_0;
	wire w_dff_A_uJb5aO7c0_0;
	wire w_dff_A_x1vViBng8_0;
	wire w_dff_A_1uY6diiv4_0;
	wire w_dff_A_eAMttTla5_0;
	wire w_dff_A_OfXwfuHb9_0;
	wire w_dff_A_gWMkCEob1_0;
	wire w_dff_A_oF59FTBX1_0;
	wire w_dff_A_NDELbzed2_0;
	wire w_dff_A_ymAq8dQA9_0;
	wire w_dff_A_WlU1xGcq3_0;
	wire w_dff_A_NfW3AOru4_0;
	wire w_dff_A_8Dz2EDTB9_0;
	wire w_dff_A_uBZOwhgZ3_0;
	wire w_dff_A_uPz3MWrE4_0;
	wire w_dff_A_uyJTFp7l6_0;
	wire w_dff_A_BXQ9Qi7n6_0;
	wire w_dff_A_Ym7FKmPV3_0;
	wire w_dff_A_NtDooD8A4_0;
	wire w_dff_A_a4NcGCQI4_2;
	wire w_dff_A_QKnPcnPn2_0;
	wire w_dff_A_Hao5ODkW2_0;
	wire w_dff_A_EcaA0shY7_0;
	wire w_dff_A_ZAwsnKGm4_0;
	wire w_dff_A_OxrKGEvZ3_0;
	wire w_dff_A_NOStlwC57_0;
	wire w_dff_A_9YIZJniB0_0;
	wire w_dff_A_yG9z7hDW0_0;
	wire w_dff_A_Q9KC1zNf3_0;
	wire w_dff_A_OSNP0dIS0_0;
	wire w_dff_A_yVb18zSB1_0;
	wire w_dff_A_MDeFogBm4_0;
	wire w_dff_A_4TGxZztf4_0;
	wire w_dff_A_dURurCjF6_0;
	wire w_dff_A_MB8IZYMQ1_0;
	wire w_dff_A_vjfKkrUX7_0;
	wire w_dff_A_yQwX7LmR1_0;
	wire w_dff_A_ImnVyFQH6_0;
	wire w_dff_A_pcj3Bf2f3_0;
	wire w_dff_A_dO4I6j6B6_0;
	wire w_dff_A_ZXNNfepP5_0;
	wire w_dff_A_nMfCKEhz9_0;
	wire w_dff_A_cisNgDn53_0;
	wire w_dff_A_lfGETm8V7_0;
	wire w_dff_A_InPKo1G29_2;
	wire w_dff_A_RwKtsVDd3_0;
	wire w_dff_A_TVtmQzl49_0;
	wire w_dff_A_uTmujb7u3_0;
	wire w_dff_A_wPBheNWZ1_0;
	wire w_dff_A_uTPbD6A49_0;
	wire w_dff_A_XO7BKUc82_0;
	wire w_dff_A_oGIhk7Qj5_0;
	wire w_dff_A_ZGZuUFTI9_0;
	wire w_dff_A_WfTViwob2_0;
	wire w_dff_A_DTvmW2dO8_0;
	wire w_dff_A_CPf2djyN7_0;
	wire w_dff_A_V5iusUgI1_0;
	wire w_dff_A_pxZ1f6pi0_0;
	wire w_dff_A_9ICQSLOh2_0;
	wire w_dff_A_1sTci4oT5_0;
	wire w_dff_A_ra3nyH0h2_0;
	wire w_dff_A_oyCfNH146_0;
	wire w_dff_A_zPiRrCQN5_0;
	wire w_dff_A_FsaLbdMq2_0;
	wire w_dff_A_9lY6IMdd1_0;
	wire w_dff_A_n6aSC5Pb0_0;
	wire w_dff_A_5Y76D0cZ2_0;
	wire w_dff_A_eXrdnHUC7_2;
	wire w_dff_A_u1sMo46g2_0;
	wire w_dff_A_RJYXGLdr0_0;
	wire w_dff_A_FC7ANpav9_0;
	wire w_dff_A_C4p3N5fD4_0;
	wire w_dff_A_OVkOGZZK8_0;
	wire w_dff_A_4Xb0k8sk7_0;
	wire w_dff_A_y4KY4Ro38_0;
	wire w_dff_A_oydTkysa7_0;
	wire w_dff_A_1OC6eWBv6_0;
	wire w_dff_A_8FBFMwdL0_0;
	wire w_dff_A_OUrSPaBO9_0;
	wire w_dff_A_avoKFPxF5_0;
	wire w_dff_A_p3HQEiET6_0;
	wire w_dff_A_Y0mOjRHp2_0;
	wire w_dff_A_xfR59igd6_0;
	wire w_dff_A_Q0dzHYlW1_0;
	wire w_dff_A_LyjDufMW5_0;
	wire w_dff_A_wM3WlXOf4_0;
	wire w_dff_A_UEQdPovE5_0;
	wire w_dff_A_XYofgA0K5_0;
	wire w_dff_A_qIgnYrt85_0;
	wire w_dff_A_MVFrvlp67_0;
	wire w_dff_A_GOXYE6495_2;
	wire w_dff_A_rrgAvDCo1_0;
	wire w_dff_A_abmdGtit6_0;
	wire w_dff_A_ePLLtNQT8_0;
	wire w_dff_A_fiByJLgb2_0;
	wire w_dff_A_1YU481FK8_0;
	wire w_dff_A_ShF32XcK9_0;
	wire w_dff_A_5dwbqAYk4_0;
	wire w_dff_A_OypP6riD4_0;
	wire w_dff_A_UTTrFT1U0_0;
	wire w_dff_A_N3aA6p2m1_0;
	wire w_dff_A_lvY1EtVy5_0;
	wire w_dff_A_6o4csVod0_0;
	wire w_dff_A_G1GFN9IS1_0;
	wire w_dff_A_TIljWDqV9_0;
	wire w_dff_A_fOszQBqM9_0;
	wire w_dff_A_peONeGsp4_0;
	wire w_dff_A_1QSxXp7N7_0;
	wire w_dff_A_iXLeS8WU8_0;
	wire w_dff_A_O8wjXCpb9_0;
	wire w_dff_A_rFGLQ1Lb2_0;
	wire w_dff_A_bN2Cbh5L4_0;
	wire w_dff_A_n5YAR0C05_0;
	wire w_dff_A_59IPRAJR0_2;
	wire w_dff_A_pM1DUbWl9_0;
	wire w_dff_A_L8T2dIff8_0;
	wire w_dff_A_BnICfQy90_0;
	wire w_dff_A_aRN2JmoO8_0;
	wire w_dff_A_j54jGt0z4_0;
	wire w_dff_A_zGD3TdRE6_0;
	wire w_dff_A_d6iSFEJg3_0;
	wire w_dff_A_6Xb0cQX82_0;
	wire w_dff_A_SqzJMgv70_0;
	wire w_dff_A_MTH5LWoJ7_0;
	wire w_dff_A_YFehd9rc3_0;
	wire w_dff_A_q6UiJCbA5_0;
	wire w_dff_A_NLG1sG239_0;
	wire w_dff_A_GJNI5DAO8_0;
	wire w_dff_A_uz3Te3mx6_0;
	wire w_dff_A_I9rOEXAD0_0;
	wire w_dff_A_P8K2jCqv9_0;
	wire w_dff_A_M0u9Bkms3_0;
	wire w_dff_A_rLTcttWG4_0;
	wire w_dff_A_hhWKcooo7_0;
	wire w_dff_A_dHxLZpSh1_0;
	wire w_dff_A_MqvG8nK23_0;
	wire w_dff_A_mkTkpc2K4_2;
	wire w_dff_A_BxVuoL1y7_0;
	wire w_dff_A_bqeudy5n0_0;
	wire w_dff_A_CdCkLa7D5_0;
	wire w_dff_A_ZsCv6uyj3_0;
	wire w_dff_A_1idQKwMK6_0;
	wire w_dff_A_HzLMPAOj1_0;
	wire w_dff_A_TEuTX86W1_0;
	wire w_dff_A_rBjjsj4U8_0;
	wire w_dff_A_YOusoUNe5_0;
	wire w_dff_A_AfEyve3F0_0;
	wire w_dff_A_jHbabJfW1_0;
	wire w_dff_A_NwNF5n1l2_0;
	wire w_dff_A_z1a9tGqO4_0;
	wire w_dff_A_iXv1nSAS2_0;
	wire w_dff_A_iDc2sWM92_0;
	wire w_dff_A_QowlBAUQ5_0;
	wire w_dff_A_YJBpxGXv4_0;
	wire w_dff_A_NyZzKhCF1_0;
	wire w_dff_A_FRdV0Z5a2_0;
	wire w_dff_A_kiJeiQer6_2;
	wire w_dff_A_UoJuqcDo4_0;
	wire w_dff_A_qSCHkV0l4_0;
	wire w_dff_A_ZImzSTMT4_0;
	wire w_dff_A_XJWHgbw74_0;
	wire w_dff_A_efk9w5E78_0;
	wire w_dff_A_vpuqTvCW6_0;
	wire w_dff_A_3RPdVmKu5_0;
	wire w_dff_A_nfN0EqsT1_0;
	wire w_dff_A_EcRKQ7Eb1_0;
	wire w_dff_A_12o9XDQz3_0;
	wire w_dff_A_tIJq6nDZ2_0;
	wire w_dff_A_3zzxky5u6_0;
	wire w_dff_A_1iX5lI5n9_0;
	wire w_dff_A_XhDmHjHt3_0;
	wire w_dff_A_eznnZOei5_0;
	wire w_dff_A_wXsQ7jNt0_0;
	wire w_dff_A_4uSpfTKP6_0;
	wire w_dff_A_tMcjrITX7_0;
	wire w_dff_A_1Y5z3GHA5_2;
	wire w_dff_A_6mKFJZtH4_0;
	wire w_dff_A_SClSIx3D4_0;
	wire w_dff_A_mO3TAI7N9_0;
	wire w_dff_A_BsXMaR2q6_0;
	wire w_dff_A_wyyUYXBi0_0;
	wire w_dff_A_1K3U7Dog4_0;
	wire w_dff_A_Zkpdexlu9_0;
	wire w_dff_A_bgTExiT65_0;
	wire w_dff_A_39LV0Tle6_0;
	wire w_dff_A_YAEenahu5_0;
	wire w_dff_A_QZqQ3MDU8_0;
	wire w_dff_A_ysQvKkY57_0;
	wire w_dff_A_Qo3YxnXS4_0;
	wire w_dff_A_rW1A6dMn7_0;
	wire w_dff_A_gtzFmx681_0;
	wire w_dff_A_fe9XJN7P3_0;
	wire w_dff_A_1RVBZJEC9_2;
	wire w_dff_A_lg3O4dSr0_0;
	wire w_dff_A_PyMsVnxY7_0;
	wire w_dff_A_tjNuhyl60_0;
	wire w_dff_A_Bc6Pi9S97_0;
	wire w_dff_A_DHpRZK6A6_0;
	wire w_dff_A_8VtVH8Zc9_0;
	wire w_dff_A_tMm9O2NF4_0;
	wire w_dff_A_tk5gZflL7_0;
	wire w_dff_A_zMzcfgqZ6_0;
	wire w_dff_A_g6DLGaA93_0;
	wire w_dff_A_9zgSJVXK9_0;
	wire w_dff_A_y11EIFcp0_0;
	wire w_dff_A_gW4fRWOh3_0;
	wire w_dff_A_eo7xhwDm5_0;
	wire w_dff_A_S1PPWCCf4_0;
	wire w_dff_A_OqjykQxo0_0;
	wire w_dff_A_Ix4GRr790_0;
	wire w_dff_A_6f5g0anK1_2;
	wire w_dff_A_38CuFKku4_0;
	wire w_dff_A_SzKK9Fja5_0;
	wire w_dff_A_mmkQvEi36_0;
	wire w_dff_A_rqeZYy1E6_0;
	wire w_dff_A_T099VD2t0_0;
	wire w_dff_A_TWZOUUEW6_0;
	wire w_dff_A_fJZqshVa5_0;
	wire w_dff_A_MwaSSTyt6_0;
	wire w_dff_A_KLBo8KOs1_0;
	wire w_dff_A_tGUpexzz3_0;
	wire w_dff_A_c8KBWf9d8_0;
	wire w_dff_A_tFSk4fLO9_0;
	wire w_dff_A_uVeofMBM9_0;
	wire w_dff_A_iJPTT4OC1_0;
	wire w_dff_A_KugvriIB1_0;
	wire w_dff_A_NUMpbhzy4_0;
	wire w_dff_A_Wdrk0HfE8_0;
	wire w_dff_A_gMde8Pq87_2;
	wire w_dff_A_mUELzTNT7_0;
	wire w_dff_A_EEbaj8fe6_0;
	wire w_dff_A_lbS2m6tv1_0;
	wire w_dff_A_yjByoIOU9_0;
	wire w_dff_A_tmQ5SDGO2_0;
	wire w_dff_A_M7a6ZIA49_0;
	wire w_dff_A_aCwq3sVQ4_0;
	wire w_dff_A_6gz6ynCf5_0;
	wire w_dff_A_MUyoWCGW4_0;
	wire w_dff_A_ba10qmmZ2_0;
	wire w_dff_A_lvd94Pe93_0;
	wire w_dff_A_misKMs3Y2_0;
	wire w_dff_A_NYuERfdE4_0;
	wire w_dff_A_xm2H86XY3_0;
	wire w_dff_A_jdEkR0ve4_0;
	wire w_dff_A_snxzDqXo5_0;
	wire w_dff_A_jl9DVvEN6_1;
	wire w_dff_A_zmXuPf7S1_0;
	wire w_dff_A_B9T7G3PS5_0;
	wire w_dff_A_eiicRrsq4_0;
	wire w_dff_A_AXlfZhwq4_0;
	wire w_dff_A_vUYvSS6t9_0;
	wire w_dff_A_xD0wl7nN6_0;
	wire w_dff_A_jluNa5RS8_0;
	wire w_dff_A_6WXl4seo8_0;
	wire w_dff_A_TIM5BsFK4_0;
	wire w_dff_A_lu6Xl9b30_0;
	wire w_dff_A_ddVIOdPE8_0;
	wire w_dff_A_oZ1LAy2l3_0;
	wire w_dff_A_NxvexjAB3_0;
	wire w_dff_A_2Dx8xmxM2_0;
	wire w_dff_A_OLFFV1fO6_0;
	wire w_dff_A_MagLAuyn3_0;
	wire w_dff_A_i04Fd4Iv1_0;
	wire w_dff_A_hFhS8SEb8_0;
	wire w_dff_A_vMBXWVcX1_0;
	wire w_dff_A_sw7Bi2oV4_0;
	wire w_dff_A_vYiPlc5d7_0;
	wire w_dff_A_YqVRDqit3_0;
	wire w_dff_A_9BfOiUdX0_1;
	wire w_dff_A_svXeqnba4_0;
	wire w_dff_A_XsK7Yd838_0;
	wire w_dff_A_pexPtVeX2_0;
	wire w_dff_A_Bz761Y1V6_0;
	wire w_dff_A_0nTzUGia5_0;
	wire w_dff_A_Z34NABgk1_0;
	wire w_dff_A_20tJYRad7_0;
	wire w_dff_A_ghTPUouy1_0;
	wire w_dff_A_iOmxQnJb5_0;
	wire w_dff_A_Vnydl0Od7_0;
	wire w_dff_A_bmTpO0vX7_0;
	wire w_dff_A_mfa69Sig2_0;
	wire w_dff_A_EUFshqh56_0;
	wire w_dff_A_7VTg7RxP4_0;
	wire w_dff_A_gv9A0ZLZ1_0;
	wire w_dff_A_3Yth2iJE9_0;
	wire w_dff_A_c9c0t3Hh7_0;
	wire w_dff_A_D9F6MfN13_0;
	wire w_dff_A_VFbQQQC16_0;
	wire w_dff_A_PDpvrrDB6_0;
	wire w_dff_A_iUwMaq9k0_0;
	wire w_dff_A_nNBaGDLA8_0;
	wire w_dff_A_SAvAS5ac4_2;
	wire w_dff_A_0ZmKSFZq0_0;
	wire w_dff_A_Su4B4ZxA6_0;
	wire w_dff_A_tEpm2T1x9_0;
	wire w_dff_A_yaQLeFVI3_0;
	wire w_dff_A_SgJ4JHkq2_0;
	wire w_dff_A_qmvuXtsa6_0;
	wire w_dff_A_uAOCnff88_0;
	wire w_dff_A_e7AYugUu0_0;
	wire w_dff_A_bELKA3yD0_0;
	wire w_dff_A_xYqzNEyw7_0;
	wire w_dff_A_LqrRWkdQ1_0;
	wire w_dff_A_v4tDnsaq1_0;
	wire w_dff_A_1lamenRD4_0;
	wire w_dff_A_GkJoW1s90_2;
	wire w_dff_A_kHHxi3Eg5_0;
	wire w_dff_A_tWAHHwad8_0;
	wire w_dff_A_yRaoE6ub6_0;
	wire w_dff_A_QSB2vzVF0_0;
	wire w_dff_A_CR2oVjbp0_0;
	wire w_dff_A_pqyknbbY7_0;
	wire w_dff_A_AMzYwiJV6_0;
	wire w_dff_A_RnIMg0oD0_0;
	wire w_dff_A_95iPqvg70_0;
	wire w_dff_A_zNjTUnoR9_0;
	wire w_dff_A_vrUoWyx38_0;
	wire w_dff_A_r8nApT5A3_0;
	wire w_dff_A_Np0KkK0m3_0;
	wire w_dff_A_lGedkKfI9_0;
	wire w_dff_A_SEr1vClL9_2;
	wire w_dff_A_lD8JTnvG5_0;
	wire w_dff_A_sCHPlANe3_0;
	wire w_dff_A_iYkt8Cqv1_0;
	wire w_dff_A_cMRybDRq1_0;
	wire w_dff_A_2X7E52Sn6_0;
	wire w_dff_A_a0qmWvzK5_0;
	wire w_dff_A_mbANAgzG8_0;
	wire w_dff_A_ICFyReGj3_0;
	wire w_dff_A_rsWZvl7p4_0;
	wire w_dff_A_1obtUJJx0_0;
	wire w_dff_A_UyrFTC8R9_0;
	wire w_dff_A_egFEADV73_0;
	wire w_dff_A_tWd3LFVg6_0;
	wire w_dff_A_FP0rTFvM2_2;
	wire w_dff_A_FCe3qd0e1_0;
	wire w_dff_A_eRd5USvR9_0;
	wire w_dff_A_E8eSqdeW2_0;
	wire w_dff_A_kGiw5Vi43_0;
	wire w_dff_A_Gh4X3QHl7_0;
	wire w_dff_A_ZzrmXXHP1_0;
	wire w_dff_A_uBmhPkcc7_0;
	wire w_dff_A_PgWNlTPo2_0;
	wire w_dff_A_ik9mDEgu2_0;
	wire w_dff_A_AZEL8e0W7_0;
	wire w_dff_A_SQfEEdu85_0;
	wire w_dff_A_0UCpNHT47_0;
	wire w_dff_A_rfYQQaAQ3_0;
	wire w_dff_A_y6aTy7GM3_0;
	wire w_dff_A_VYShTGcq8_1;
	wire w_dff_A_xyW8xbEx9_0;
	wire w_dff_A_WCff8LI80_0;
	wire w_dff_A_Fw1PBLGG1_0;
	wire w_dff_A_40glEXYn3_0;
	wire w_dff_A_EUyf9Bfa4_0;
	wire w_dff_A_4EGNw5dr6_0;
	wire w_dff_A_7n38dQYW1_0;
	wire w_dff_A_xxKOFpVR4_0;
	wire w_dff_A_K0lIoeYy9_0;
	wire w_dff_A_IWT87sXT8_0;
	wire w_dff_A_nKDkwGaY3_0;
	wire w_dff_A_zCMl7dFs7_0;
	wire w_dff_A_OC11v3q14_0;
	wire w_dff_A_Jr3knpH14_0;
	wire w_dff_A_uiFkqbSb7_0;
	wire w_dff_A_e8F93ljk0_0;
	wire w_dff_A_OdXzH4895_0;
	wire w_dff_A_bMx2MXwA4_0;
	wire w_dff_A_GsjzM8tQ4_0;
	wire w_dff_A_UAv8zeNK0_1;
	wire w_dff_A_ls6mhGSr5_0;
	wire w_dff_A_4ocDkuqr3_0;
	wire w_dff_A_bUbhWxaa5_0;
	wire w_dff_A_ESFZwOak5_0;
	wire w_dff_A_evMm0Wyl8_0;
	wire w_dff_A_cqcqpeiv9_0;
	wire w_dff_A_3dtCgJOa6_0;
	wire w_dff_A_hLjg8dKo5_0;
	wire w_dff_A_xFTgryao0_0;
	wire w_dff_A_htkS74VD0_0;
	wire w_dff_A_RvdXaJ2C8_0;
	wire w_dff_A_fNsojorH1_0;
	wire w_dff_A_zjiM5xx56_0;
	wire w_dff_A_nRxtJe0P7_0;
	wire w_dff_A_IgwmqSnl4_1;
	wire w_dff_A_CVw9f9ZQ0_0;
	wire w_dff_A_kgvT1LDn1_0;
	wire w_dff_A_QsJHV1aW7_0;
	wire w_dff_A_aWkJYRAU2_0;
	wire w_dff_A_eC2gi2Dt8_0;
	wire w_dff_A_s59l3sbf2_0;
	wire w_dff_A_DRdD1hxp6_0;
	wire w_dff_A_6XBHXxyY9_0;
	wire w_dff_A_zWnInFWt9_0;
	wire w_dff_A_cJmTzp6k2_0;
	wire w_dff_A_v9fxuwNP4_0;
	wire w_dff_A_TagAa3n83_0;
	wire w_dff_A_texKzv0j4_0;
	wire w_dff_A_jsGW8a3P6_0;
	wire w_dff_A_rRSyD1XI1_0;
	wire w_dff_A_K4sjGOlI5_0;
	wire w_dff_A_elshjJ2a6_0;
	wire w_dff_A_b7Uj8T3n5_1;
	wire w_dff_A_Q5Bl4VHM5_0;
	wire w_dff_A_F6Fyb4PK9_0;
	wire w_dff_A_ORhDGbi24_0;
	wire w_dff_A_yIg9xb0S5_0;
	wire w_dff_A_VuKjo45b0_0;
	wire w_dff_A_aFvmcpgY1_0;
	wire w_dff_A_RrmLO3lS0_0;
	wire w_dff_A_FbwFgVBz2_0;
	wire w_dff_A_B8YhUJlE8_0;
	wire w_dff_A_O7wYAVdt7_2;
	wire w_dff_A_cJ1xjnVx9_0;
	wire w_dff_A_O5aBwdkq7_0;
	wire w_dff_A_MUpUZpCL0_0;
	wire w_dff_A_melqquDJ0_0;
	wire w_dff_A_k0NN3Ywp3_0;
	wire w_dff_A_G7tl7YLo8_0;
	wire w_dff_A_Bkgeuktz1_0;
	wire w_dff_A_t2lJX0nL8_0;
	wire w_dff_A_dKmiRRz30_0;
	wire w_dff_A_6SCb69Xz2_0;
	wire w_dff_A_Ryq8wyXX4_0;
	wire w_dff_A_UNqPTvZZ1_0;
	wire w_dff_A_8AKhhv408_0;
	wire w_dff_A_TjtWKR5k2_1;
	wire w_dff_A_6O1ncbqr8_0;
	wire w_dff_A_Z8S8p4Et6_0;
	wire w_dff_A_C8sX4F7e2_0;
	wire w_dff_A_AbcY5CPb6_0;
	wire w_dff_A_cXmOX0607_0;
	wire w_dff_A_1mje5fvU4_0;
	wire w_dff_A_7OsreSFE6_0;
	wire w_dff_A_DG1LGQhe9_0;
	wire w_dff_A_4jxs10DW8_0;
	wire w_dff_A_EKGmmqRE8_0;
	wire w_dff_A_H3Ie7GYo3_0;
	wire w_dff_A_5v8gAEv80_0;
	wire w_dff_A_ICQfSecU6_1;
	wire w_dff_A_HBq5g8BD2_0;
	wire w_dff_A_UurNwGC50_0;
	wire w_dff_A_BMfZRL0S7_0;
	wire w_dff_A_zXAtMbVa4_0;
	wire w_dff_A_lNRIbo8S5_0;
	wire w_dff_A_mLd0LmI91_0;
	wire w_dff_A_G7go82SA9_0;
	wire w_dff_A_XMX7SZIL3_0;
	wire w_dff_A_bfLltZk06_0;
	wire w_dff_A_eWJlX53v9_0;
	wire w_dff_A_VCaEGqlS3_0;
	wire w_dff_A_R1gMeFM25_0;
	wire w_dff_A_VpNYpXeO6_0;
	wire w_dff_A_DX7YKSnO2_1;
	wire w_dff_A_V1ipFKI50_0;
	wire w_dff_A_71wCERyd5_0;
	wire w_dff_A_Qk0UTxZ88_0;
	wire w_dff_A_bKMqDHhF2_0;
	wire w_dff_A_9JDT9cUL6_0;
	wire w_dff_A_733b8GSb6_0;
	wire w_dff_A_5MfQFAFV6_0;
	wire w_dff_A_ZfBiNJ3K1_0;
	wire w_dff_A_ifCqtWTi1_0;
	wire w_dff_A_mpvxJe0J1_0;
	wire w_dff_A_T6zbLVaV4_0;
	wire w_dff_A_xH5JX65S8_0;
	wire w_dff_A_XOZeyNdL8_0;
	wire w_dff_A_h8iynxhB5_0;
	wire w_dff_A_bVecHrRU9_0;
	wire w_dff_A_YcIv6Ant5_2;
	wire w_dff_A_LvCLKEHe6_0;
	wire w_dff_A_p7Vu2e9s1_0;
	wire w_dff_A_LCsMit8Q6_0;
	wire w_dff_A_GjJmMtvB5_0;
	wire w_dff_A_1AE6zYd27_0;
	wire w_dff_A_hvEwHQYS9_0;
	wire w_dff_A_2uN7VHXT1_0;
	wire w_dff_A_gla9WPjz3_0;
	wire w_dff_A_tfKgofmr3_0;
	wire w_dff_A_HdoQgVSL0_0;
	wire w_dff_A_IckMEeNR6_0;
	wire w_dff_A_YYKl1Pk89_0;
	wire w_dff_A_8s3ojIhh0_0;
	wire w_dff_A_zejxgGKu4_1;
	wire w_dff_A_Swr7ePZR6_0;
	wire w_dff_A_lxhTkNBZ7_0;
	wire w_dff_A_7LmGl7iO2_0;
	wire w_dff_A_3kEi4fWn7_0;
	wire w_dff_A_NqsgGsBB6_0;
	wire w_dff_A_vKsavxpf8_0;
	wire w_dff_A_cC5lB1vs8_0;
	wire w_dff_A_YZ7eOhAK6_0;
	wire w_dff_A_CdxDHFtJ8_0;
	wire w_dff_A_pD1sp2v62_0;
	wire w_dff_A_T9d2ZPJ94_0;
	wire w_dff_A_ToOisfaa0_0;
	wire w_dff_A_GJ5SWN8q8_1;
	wire w_dff_A_BAhmKwth2_0;
	wire w_dff_A_GiN9TrU71_0;
	wire w_dff_A_uzZ4rg3E6_0;
	wire w_dff_A_n2wEUx6e6_0;
	wire w_dff_A_oikmc1Of0_0;
	wire w_dff_A_LtPMtd7i4_0;
	wire w_dff_A_ilgVdTpA3_0;
	wire w_dff_A_Q79gbO417_0;
	wire w_dff_A_tnGp9QKG4_0;
	wire w_dff_A_dCZ14Seu2_0;
	wire w_dff_A_tyhJ43JA8_0;
	wire w_dff_A_N9Y2z3J89_0;
	wire w_dff_A_Lm0zIVvd0_0;
	wire w_dff_A_Tr4PIag82_0;
	wire w_dff_A_Mw7p5bZZ9_1;
	wire w_dff_A_riPvdVm94_0;
	wire w_dff_A_96hsr8m75_0;
	wire w_dff_A_UDPQ0TMp0_0;
	wire w_dff_A_NVelT6201_0;
	wire w_dff_A_zNyBUt6x9_0;
	wire w_dff_A_QZloL7CX6_0;
	wire w_dff_A_kIMkhQaN1_0;
	wire w_dff_A_rOJqvXHS1_0;
	wire w_dff_A_Jx62Wi8y3_0;
	wire w_dff_A_kyo4D9q72_0;
	wire w_dff_A_Xd1Dq2hO6_0;
	wire w_dff_A_bU2asTuS1_0;
	wire w_dff_A_EL2eZkGB1_0;
	wire w_dff_A_0W3XIyY75_0;
	wire w_dff_A_Cbga3JiT6_0;
	wire w_dff_A_tYluNs5U4_1;
	wire w_dff_A_AkfcQQ514_0;
	wire w_dff_A_VOK4Vf6D5_0;
	wire w_dff_A_UfUGh8qC2_0;
	wire w_dff_A_lfufGkjl8_0;
	wire w_dff_A_k1MVLzG81_0;
	wire w_dff_A_ZDMPVXmH9_0;
	wire w_dff_A_Z18riH2b9_0;
	wire w_dff_A_bxd1OX6V3_0;
	wire w_dff_A_A7s0WCXi5_0;
	wire w_dff_A_1hb5tI9c0_0;
	wire w_dff_A_WruQ7unO2_0;
	wire w_dff_A_AG1Yefvt4_0;
	wire w_dff_A_Js2Iwlbi9_0;
	wire w_dff_A_SDeLTR803_0;
	wire w_dff_A_lxbpSUFO1_0;
	wire w_dff_A_VZhTkJ8A9_0;
	wire w_dff_A_VCOqhx971_1;
	wire w_dff_A_DSsVtlGx1_0;
	wire w_dff_A_bvgUWODH4_0;
	wire w_dff_A_wx7f1ws41_0;
	wire w_dff_A_lll9M0gF2_0;
	wire w_dff_A_VDnvuVfq4_0;
	wire w_dff_A_B7n5shkg1_0;
	wire w_dff_A_rIVw8x059_0;
	wire w_dff_A_kc5eWfPe8_0;
	wire w_dff_A_GruaQll22_0;
	wire w_dff_A_GomFKmbj6_0;
	wire w_dff_A_nIofH8gm5_0;
	wire w_dff_A_Qkga69BT1_0;
	wire w_dff_A_Zs6yYYrq1_0;
	wire w_dff_A_6mdw8nKD8_0;
	wire w_dff_A_zjPEDVJY6_0;
	wire w_dff_A_gisvbRPS4_0;
	wire w_dff_A_wMQj2HOW1_0;
	wire w_dff_A_ZeDwIcdB4_0;
	wire w_dff_A_w5QIYCX30_0;
	wire w_dff_A_LwGy0wKt8_1;
	wire w_dff_A_UMWbK1I59_0;
	wire w_dff_A_wOpQxbba9_0;
	wire w_dff_A_H628PjGa7_0;
	wire w_dff_A_5dcQwNL23_0;
	wire w_dff_A_RI9xOgm12_0;
	wire w_dff_A_6mZPKRnS4_0;
	wire w_dff_A_byCsdSYY1_0;
	wire w_dff_A_RE8xx5Y86_0;
	wire w_dff_A_Gz7OPc0w6_0;
	wire w_dff_A_Ey6ZTc9l3_0;
	wire w_dff_A_5pYGop5e6_0;
	wire w_dff_A_USPkTnw22_0;
	wire w_dff_A_8hLPYmK71_0;
	wire w_dff_A_qNgihvDH8_0;
	wire w_dff_A_Xjdwz6K91_0;
	wire w_dff_A_3OgcdmYG1_0;
	wire w_dff_A_PYPhHZgk5_0;
	wire w_dff_A_42ToleIv4_0;
	wire w_dff_A_FSDJereM4_2;
	wire w_dff_A_HHiqvebf1_0;
	wire w_dff_A_dJUBUOwU3_0;
	wire w_dff_A_lub9GHR85_0;
	wire w_dff_A_JOpDG86Z1_0;
	wire w_dff_A_dLcHtqtE8_0;
	wire w_dff_A_R51BVZxY1_0;
	wire w_dff_A_WF5LyqbK8_0;
	wire w_dff_A_5ltDjXuT8_2;
	wire w_dff_A_9elRzTD92_0;
	wire w_dff_A_13r5drHY0_0;
	wire w_dff_A_tKUZ6f0L6_0;
	wire w_dff_A_ShtN6qJE5_0;
	wire w_dff_A_u0euAwMQ6_0;
	wire w_dff_A_nB7mZ6QU1_0;
	wire w_dff_A_09IHvNaL4_2;
	wire w_dff_A_0z5KShPv8_0;
	wire w_dff_A_wdlBjPRD8_0;
	wire w_dff_A_avpExcFZ4_0;
	wire w_dff_A_ZRN1OL2a7_0;
	wire w_dff_A_jzCJoAw88_0;
	wire w_dff_A_9kWVhh6m3_0;
	wire w_dff_A_rfuAabCB2_0;
	wire w_dff_A_iPLSuyM16_0;
	wire w_dff_A_I5lE0ZMI8_0;
	wire w_dff_A_jId4hxGS5_0;
	wire w_dff_A_GD0IxNRl0_0;
	wire w_dff_A_SWMAgAUJ9_2;
	wire w_dff_A_X8hPznN83_0;
	wire w_dff_A_t7Y1YB2L2_0;
	wire w_dff_A_gRc20hDv8_0;
	wire w_dff_A_ZqvBhCuH3_0;
	wire w_dff_A_jjchhgrc3_0;
	wire w_dff_A_2Df1oeOe4_0;
	wire w_dff_A_0X8yqpJ23_0;
	wire w_dff_A_JglzB5JZ1_0;
	wire w_dff_A_vtKLSkfV0_0;
	wire w_dff_A_iAdslHC67_0;
	wire w_dff_A_Vs5YWyeM5_0;
	wire w_dff_A_Z13qQidg2_2;
	wire w_dff_A_iaw37lKi0_0;
	wire w_dff_A_PJIlZVhL5_0;
	wire w_dff_A_nPVp7hgW5_0;
	wire w_dff_A_Msx2FQCk2_0;
	wire w_dff_A_OnEzG93A8_0;
	wire w_dff_A_686Kjme78_0;
	wire w_dff_A_zC53FGcG8_0;
	wire w_dff_A_NZTKntos3_2;
	wire w_dff_A_E6caPdRQ5_0;
	wire w_dff_A_UFV7DIaL8_0;
	wire w_dff_A_1TEYMkQF2_0;
	wire w_dff_A_jshwYzZa9_0;
	wire w_dff_A_h08DBtkS3_0;
	wire w_dff_A_HJmdpaXa5_0;
	wire w_dff_A_aZfPtXqN0_0;
	wire w_dff_A_daZ8IuUb1_0;
	wire w_dff_A_qtJUbwCW9_2;
	wire w_dff_A_OQdHWbEG0_0;
	wire w_dff_A_ld4v8GRD8_0;
	wire w_dff_A_BvsGC0n13_0;
	wire w_dff_A_v46Juft24_0;
	wire w_dff_A_jv2rH8Mi2_0;
	wire w_dff_A_ZEUcR0DH0_0;
	wire w_dff_A_vksXmgQj2_0;
	wire w_dff_A_XeOilhG90_0;
	wire w_dff_A_gjWOBSJW8_0;
	wire w_dff_A_8sHvb8cP2_0;
	wire w_dff_A_0IUNpq9e5_2;
	wire w_dff_A_qjBO1FYl0_0;
	wire w_dff_A_lyixb6jW9_0;
	wire w_dff_A_BEnYyW0t0_0;
	wire w_dff_A_MV8PkqOu3_0;
	wire w_dff_A_ALKN8NLc6_0;
	wire w_dff_A_J35WFDl26_0;
	wire w_dff_A_9Y82Ca4a4_0;
	wire w_dff_A_pfcEfYFX1_0;
	wire w_dff_A_hxEKEWhE7_0;
	wire w_dff_A_7okTC8Yv1_2;
	wire w_dff_A_UdOHfssJ2_0;
	wire w_dff_A_wUyKTX7H2_0;
	wire w_dff_A_136G7pCc2_0;
	wire w_dff_A_6xN0F4Ky9_0;
	wire w_dff_A_El1yBSPs2_0;
	wire w_dff_A_jc0Nd6Ch7_0;
	wire w_dff_A_N7VnJMEt4_0;
	wire w_dff_A_la5HpM0d0_2;
	wire w_dff_A_uhU1qVvX1_0;
	wire w_dff_A_ld8Okegi0_0;
	wire w_dff_A_rwPsz4Vu7_0;
	wire w_dff_A_MvUyKAxC6_0;
	wire w_dff_A_b47ixkoL5_0;
	wire w_dff_A_x6MDbt6g2_0;
	wire w_dff_A_d4v70wGJ5_0;
	wire w_dff_A_TZiQctQs4_0;
	wire w_dff_A_K4sCI48D9_2;
	wire w_dff_A_uK49aPco9_0;
	wire w_dff_A_bPgwSsLQ7_0;
	wire w_dff_A_4DRn44Wr6_0;
	wire w_dff_A_zp1xJMM23_0;
	wire w_dff_A_1MHXBTZU7_0;
	wire w_dff_A_xTISa4Gm6_0;
	wire w_dff_A_pEwuXo406_0;
	wire w_dff_A_rrLmQzxn5_0;
	wire w_dff_A_Lf5p5ICS0_0;
	wire w_dff_A_mzwdSda61_0;
	wire w_dff_A_aqlIY8yf5_2;
	wire w_dff_A_DFSNL7144_0;
	wire w_dff_A_rmPsxOxx1_0;
	wire w_dff_A_amVKJrEN7_0;
	wire w_dff_A_oxQn4gGd5_0;
	wire w_dff_A_7eb8C3BA7_0;
	wire w_dff_A_t4oGr6SV6_0;
	wire w_dff_A_xRwmHPoW1_0;
	wire w_dff_A_bNr40E0a0_0;
	wire w_dff_A_ZOWXptlU5_0;
	wire w_dff_A_eXtTYCE04_2;
	wire w_dff_A_vLQhPHQD5_0;
	wire w_dff_A_MscugdSa8_0;
	wire w_dff_A_NLAFOEsr3_0;
	wire w_dff_A_84gJBveH0_0;
	wire w_dff_A_loWyxih61_0;
	wire w_dff_A_DPlg8d4j7_0;
	wire w_dff_A_vEcDfA282_2;
	wire w_dff_A_hjGNh0Ov3_0;
	wire w_dff_A_yICnxMbu7_0;
	wire w_dff_A_J4t0CWys9_0;
	wire w_dff_A_85X6aOHD4_0;
	wire w_dff_A_q0fHmOFP9_0;
	wire w_dff_A_hh8VPUhr5_0;
	wire w_dff_A_zd9X5JB64_0;
	wire w_dff_A_82lGhO7J4_0;
	wire w_dff_A_DN1txea69_0;
	wire w_dff_A_b47UtnYZ5_2;
	wire w_dff_A_RNg2sWhJ3_0;
	wire w_dff_A_bTnVNkDb6_0;
	wire w_dff_A_PRX7tc082_0;
	wire w_dff_A_L689P2z35_0;
	wire w_dff_A_6LTlPDZi0_0;
	wire w_dff_A_xBqalnDu3_0;
	wire w_dff_A_Jtl3DNmx6_0;
	wire w_dff_A_W5aAhiir0_0;
	wire w_dff_A_XwjwO0SP4_0;
	wire w_dff_A_TjGCcada8_2;
	wire w_dff_A_lNidFfVa1_0;
	wire w_dff_A_HnHEaCUI1_0;
	wire w_dff_A_XwUVbQzP7_0;
	wire w_dff_A_CnVd3AWM2_0;
	wire w_dff_A_3sCpdZ7t4_0;
	wire w_dff_A_EwaKgt3w8_0;
	wire w_dff_A_4JjTPkhD2_0;
	wire w_dff_A_r0clN1f40_0;
	wire w_dff_A_CNem8CWd3_2;
	wire w_dff_A_On70pndX7_0;
	wire w_dff_A_hrWcbxEX9_0;
	wire w_dff_A_D6qH2stF1_0;
	wire w_dff_A_uGb9sllM2_0;
	wire w_dff_A_r64SKWGI5_0;
	wire w_dff_A_rqUWwm8M5_2;
	wire w_dff_A_RVgwCXR00_0;
	wire w_dff_A_7YlJ9mEM7_0;
	wire w_dff_A_eKUg72am9_0;
	wire w_dff_A_5YzybX6G4_0;
	wire w_dff_A_YANTPxk09_0;
	wire w_dff_A_tYg2fACr8_0;
	wire w_dff_A_GNYJi9ud8_0;
	wire w_dff_A_73A43DHf0_0;
	wire w_dff_A_AdDZzCPb6_0;
	wire w_dff_A_Wj8inUZF4_2;
	wire w_dff_A_m1ysEKYC5_0;
	wire w_dff_A_TerU8ija8_0;
	wire w_dff_A_fSESxPlQ3_0;
	wire w_dff_A_hAhKblHz6_0;
	wire w_dff_A_YhryUOm46_0;
	wire w_dff_A_rakfXR4h6_0;
	wire w_dff_A_89qsdqi22_0;
	wire w_dff_A_bH1RFDNj6_0;
	wire w_dff_A_HnHM054f8_0;
	wire w_dff_A_8GjDZDev4_2;
	wire w_dff_A_OUJpiErG8_0;
	wire w_dff_A_eK4G8LO80_0;
	wire w_dff_A_iHvmmtZ78_0;
	wire w_dff_A_PmvazPgh1_0;
	wire w_dff_A_6CL4psut4_0;
	wire w_dff_A_ugJeT2CF6_0;
	wire w_dff_A_UEELVarc9_0;
	wire w_dff_A_nV8OGsFS9_0;
	wire w_dff_A_TaBL4Brs2_2;
	wire w_dff_A_aX8uaQA84_0;
	wire w_dff_A_hGewjCFE3_0;
	wire w_dff_A_RUnnaiW58_0;
	wire w_dff_A_t3nFALht1_0;
	wire w_dff_A_YoPMJSqe7_0;
	wire w_dff_A_l25XVDb49_0;
	wire w_dff_A_8tn0NyFO1_2;
	wire w_dff_A_i4HuO8CL5_0;
	wire w_dff_A_n3XQRd0k8_0;
	wire w_dff_A_27NPS7526_0;
	wire w_dff_A_R4cvzddh6_0;
	wire w_dff_A_g50MpUcu0_0;
	wire w_dff_A_p0MuONXz7_0;
	wire w_dff_A_lngJ7pm18_0;
	wire w_dff_A_wsb8YRE63_0;
	wire w_dff_A_04KwKPAI3_0;
	wire w_dff_A_qGyy1NWt1_1;
	wire w_dff_A_9udiq8sW3_0;
	wire w_dff_A_TeoSuiwr3_0;
	wire w_dff_A_ThNxRt8K2_0;
	wire w_dff_A_QN73JLJy3_0;
	wire w_dff_A_IUXEYW0j0_0;
	wire w_dff_A_AUdd2RtT1_0;
	wire w_dff_A_EVE9Od673_1;
	wire w_dff_A_IBGsDboQ8_0;
	wire w_dff_A_V5Kd3ZdL7_0;
	wire w_dff_A_P6oYNQt77_0;
	wire w_dff_A_WAYN5J1M7_0;
	wire w_dff_A_EIHCPb6O5_0;
	wire w_dff_A_n8bX5quK9_0;
	wire w_dff_A_D04dZ3iq8_0;
	wire w_dff_A_vpYvFGV21_1;
	wire w_dff_A_7d1GtTVh1_0;
	wire w_dff_A_g1BN4ShE0_0;
	wire w_dff_A_mHCZCoet1_0;
	wire w_dff_A_hR5TQsUY8_0;
	wire w_dff_A_YszCFn920_0;
	wire w_dff_A_UsZQS2zR0_0;
	wire w_dff_A_CpoHOeGU4_1;
	wire w_dff_A_40UM4Gm46_0;
	wire w_dff_A_Gn1N5gGs0_0;
	wire w_dff_A_aTlV2qug6_0;
	wire w_dff_A_6LA6kV310_0;
	wire w_dff_A_vIdbinNX7_0;
	wire w_dff_A_Y0LvZxw86_0;
	wire w_dff_A_og5PqnC33_0;
	wire w_dff_A_tquKRHqe5_0;
	wire w_dff_A_7AvzbBGl1_0;
	wire w_dff_A_NrDadm585_0;
	wire w_dff_A_zEMcQFle9_0;
	wire w_dff_A_HFgIIjdN5_2;
	wire w_dff_A_ooiQQtaX5_0;
	wire w_dff_A_1qbW3D1c9_0;
	wire w_dff_A_G3PhFWIu5_0;
	wire w_dff_A_cG5ObuCm2_0;
	wire w_dff_A_v6BqUteU5_0;
	wire w_dff_A_kiQ5mfNK6_0;
	wire w_dff_A_NQN3EwPf8_0;
	wire w_dff_A_WsOyHbMF3_0;
	wire w_dff_A_lEq7x3RI4_0;
	wire w_dff_A_coaJiB730_0;
	wire w_dff_A_e1piiQAt9_0;
	wire w_dff_A_G3wm3Dk56_0;
	wire w_dff_A_iXpnZ5X21_0;
	wire w_dff_A_cq8gQ2nO1_0;
	wire w_dff_A_pwfMFyjE5_0;
	wire w_dff_A_bz3TO0ZZ9_0;
	wire w_dff_A_TarUmmSU2_1;
	wire w_dff_A_LCwyfpbh4_0;
	wire w_dff_A_BbQD3Zps0_0;
	wire w_dff_A_GRlkehMQ9_0;
	wire w_dff_A_YfJci39l0_0;
	wire w_dff_A_FGag6nlK5_0;
	wire w_dff_A_bx1a0Rhg8_1;
	wire w_dff_A_qDFT43pG4_0;
	wire w_dff_A_4gLWta1w7_0;
	wire w_dff_A_K2ccRX827_0;
	wire w_dff_A_quagDw2X3_0;
	wire w_dff_A_YQJEdmnT2_0;
	wire w_dff_A_ax7oc2fh9_0;
	wire w_dff_A_XNWDjkFu4_0;
	wire w_dff_A_jlqeiFKW9_0;
	wire w_dff_A_mmpAPBTa5_1;
	wire w_dff_A_0KVkXGpU7_0;
	wire w_dff_A_cciaEVbv3_0;
	wire w_dff_A_ujBfOO7C9_0;
	wire w_dff_A_yNfjHOCH1_0;
	wire w_dff_A_p4NjGlo98_0;
	wire w_dff_A_phV0KFNN6_0;
	wire w_dff_A_2o5mNUNN0_1;
	wire w_dff_A_xbvKmbTE9_0;
	wire w_dff_A_f6RXQBsj0_0;
	wire w_dff_A_7i8SECPA4_0;
	wire w_dff_A_fLEa04VA1_0;
	wire w_dff_A_U9mEhFMP1_0;
	wire w_dff_A_SiaW7h2d5_0;
	wire w_dff_A_LIXYn4HD6_0;
	wire w_dff_A_d8ELLy8O1_0;
	wire w_dff_A_dkTqBuXF4_0;
	wire w_dff_A_dkFs5zUM9_2;
	wire w_dff_A_9KNRyLUd4_0;
	wire w_dff_A_06QcdIBx6_0;
	wire w_dff_A_GsRwyzkb8_0;
	wire w_dff_A_xn8VXQlt9_2;
	wire w_dff_A_rMDzb1GG3_0;
	wire w_dff_A_QLjD2Cn63_0;
	wire w_dff_A_ThgarqCR8_2;
	wire w_dff_A_qysuLA4i7_0;
	wire w_dff_A_yDzih88r6_0;
	wire w_dff_A_FcZtCV8G2_0;
	wire w_dff_A_iLcxeVf72_2;
	wire w_dff_A_f5FTN0vF7_0;
	wire w_dff_A_tQEcwiIb0_0;
	wire w_dff_A_B8Yf720Y3_0;
	wire w_dff_A_VciU7eAY5_2;
	wire w_dff_A_T84PciTu9_0;
	wire w_dff_A_9JuzTgrz0_0;
	wire w_dff_A_9NOqxWAq6_0;
	wire w_dff_A_VaDNWgO74_0;
	wire w_dff_A_iVCTOc7f1_2;
	wire w_dff_A_EIppLBGv6_0;
	wire w_dff_A_tG2R1g567_0;
	wire w_dff_A_Hb80b2Iz1_0;
	wire w_dff_A_QaYaxUiX3_2;
	wire w_dff_A_3MJ5qlH03_0;
	wire w_dff_A_faciHVZ36_0;
	wire w_dff_A_db1yODmM4_0;
	wire w_dff_A_ukNOl0VY4_2;
	wire w_dff_A_7YO21lXD0_0;
	wire w_dff_A_ubVsCTJd9_0;
	wire w_dff_A_cdz5R05I0_0;
	wire w_dff_A_zJeWIyi92_0;
	wire w_dff_A_OlaI97sX7_2;
	wire w_dff_A_S58ioXd06_0;
	wire w_dff_A_7JwnNXlg0_0;
	wire w_dff_A_hA4dvUqD0_0;
	wire w_dff_A_TBsLnPUK2_2;
	wire w_dff_A_RgdYOw2L6_0;
	wire w_dff_A_iCXl4u621_0;
	wire w_dff_A_dzvMNPTC6_2;
	wire w_dff_A_B3NYq2Fm8_0;
	wire w_dff_A_cTWeL9db5_0;
	wire w_dff_A_NOl4MacD3_2;
	wire w_dff_A_MbvSoAG75_0;
	wire w_dff_A_Udi9HLES1_2;
	wire w_dff_A_WL61JqNm2_0;
	wire w_dff_A_UrviIedY4_0;
	wire w_dff_A_rrSdEsv22_0;
	wire w_dff_A_CXlZvC9V9_2;
	wire w_dff_A_ig96CRdK0_0;
	wire w_dff_A_SWrQAXbD7_0;
	wire w_dff_A_jSG9y9fp6_2;
	wire w_dff_A_59OFn7UG6_0;
	wire w_dff_A_FIXTm6cC6_0;
	wire w_dff_A_xHbVfs0P9_2;
	wire w_dff_A_WA0UNGcW0_0;
	wire w_dff_A_2QiH6WY53_0;
	wire w_dff_A_YSK6IrZh6_2;
	wire w_dff_A_JLlRlcw25_0;
	wire w_dff_A_cr7Vl9ua8_0;
	wire w_dff_A_iMYy5M7z7_0;
	wire w_dff_A_75L5Xd0x9_0;
	wire w_dff_A_FsBNdA3J3_0;
	wire w_dff_A_vmfcvb7t4_2;
	wire w_dff_A_ZQ3ej7MJ4_0;
	wire w_dff_A_m9uFebf27_0;
	wire w_dff_A_8opvLAEc3_0;
	wire w_dff_A_CzW6VcWB6_0;
	wire w_dff_A_8ZbA5KkE6_0;
	wire w_dff_A_RE0tB8YO4_2;
	wire w_dff_A_pwFU8BN14_2;
	jnot g0000(.din(w_G545_0[2]),.dout(w_dff_A_H1rIXdYd7_1),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(w_G366_0[1]),.dout(w_dff_A_HCUTE1hH8_1),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(w_dff_A_wsRicFXl5_1),.clk(gclk));
	jnot g0005(.din(w_G338_0[1]),.dout(w_dff_A_6Sa7Xvf97_1),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(w_dff_A_EJSBV4R46_2),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(w_dff_A_C0wtGoAE3_1),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(w_dff_A_ZcBak8Wz0_1),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(w_dff_A_11gMwd6c1_1),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(w_dff_A_Yhp1kSkX5_1),.clk(gclk));
	jand g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(w_dff_A_yO5mAeIh3_2),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_1XDqtN614_1),.dout(w_dff_A_exStBqkQ5_2),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jor g0016(.dina(w_dff_B_NWXNKUrM1_0),.dinb(w_n316_0[1]),.dout(w_dff_A_TqMoaJk03_2),.clk(gclk));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(w_dff_A_X7F1HKYL4_1),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jor g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_),.clk(gclk));
	jor g0022(.dina(w_G809_3[1]),.dinb(w_dff_B_DGe8f2Ly5_1),.dout(w_dff_A_gg3PgASV0_2),.clk(gclk));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jor g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330),.clk(gclk));
	jor g0030(.dina(n330),.dinb(w_dff_B_02uGgqTc3_1),.dout(w_dff_A_1oUSV6XM4_2),.clk(gclk));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jor g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336),.clk(gclk));
	jor g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(w_dff_A_Z3ftPUiG7_2),.clk(gclk));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jor g0038(.dina(w_G809_2[1]),.dinb(w_dff_B_WU1X1XVA1_1),.dout(w_dff_A_a4NcGCQI4_2),.clk(gclk));
	jand g0039(.dina(w_n326_1[2]),.dinb(G24),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jor g0041(.dina(w_dff_B_ymTIAQl32_0),.dinb(w_G809_2[0]),.dout(n342),.clk(gclk));
	jor g0042(.dina(n342),.dinb(w_dff_B_cWl4mArx2_1),.dout(n343),.clk(gclk));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(w_dff_A_InPKo1G29_2),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(G26),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jor g0046(.dina(w_dff_B_4hxtTxcj6_0),.dinb(w_G809_1[2]),.dout(n347),.clk(gclk));
	jor g0047(.dina(n347),.dinb(w_dff_B_evs6UKxu5_1),.dout(n348),.clk(gclk));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(w_dff_A_eXrdnHUC7_2),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(G79),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jor g0051(.dina(w_dff_B_ct9crCYT1_0),.dinb(w_G809_1[1]),.dout(n352),.clk(gclk));
	jor g0052(.dina(n352),.dinb(w_dff_B_uVFbPRHM4_1),.dout(n353),.clk(gclk));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(w_dff_A_GOXYE6495_2),.clk(gclk));
	jand g0054(.dina(w_G2358_0[2]),.dinb(G80),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_n326_0[2]),.dinb(G82),.dout(n356),.clk(gclk));
	jor g0056(.dina(n356),.dinb(w_G809_1[0]),.dout(n357),.clk(gclk));
	jor g0057(.dina(n357),.dinb(w_dff_B_YVG9Lfyh4_1),.dout(n358),.clk(gclk));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(w_dff_A_59IPRAJR0_2),.clk(gclk));
	jand g0059(.dina(w_G3552_0[1]),.dinb(w_G514_2[1]),.dout(n360),.clk(gclk));
	jnot g0060(.din(w_G514_2[0]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G3546_5[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(n362),.dinb(w_n361_0[1]),.dout(n363),.clk(gclk));
	jor g0063(.dina(n363),.dinb(n360),.dout(n364),.clk(gclk));
	jnot g0064(.din(n364),.dout(n365),.clk(gclk));
	jnot g0065(.din(w_G251_5[1]),.dout(n366),.clk(gclk));
	jnot g0066(.din(w_G361_1[1]),.dout(n367),.clk(gclk));
	jand g0067(.dina(n367),.dinb(w_n366_1[2]),.dout(n368),.clk(gclk));
	jnot g0068(.din(w_G248_5[2]),.dout(n369),.clk(gclk));
	jand g0069(.dina(w_G361_1[0]),.dinb(w_n369_1[2]),.dout(n370),.clk(gclk));
	jor g0070(.dina(n370),.dinb(n368),.dout(n371),.clk(gclk));
	jnot g0071(.din(w_n371_0[1]),.dout(n372),.clk(gclk));
	jand g0072(.dina(w_n372_0[1]),.dinb(w_n365_0[1]),.dout(n373),.clk(gclk));
	jnot g0073(.din(w_G351_2[2]),.dout(n374),.clk(gclk));
	jnot g0074(.din(G3550),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_n375_4[2]),.dinb(w_n374_1[1]),.dout(n376),.clk(gclk));
	jnot g0076(.din(w_G534_2[1]),.dout(n377),.clk(gclk));
	jnot g0077(.din(w_G3552_0[0]),.dout(n378),.clk(gclk));
	jand g0078(.dina(w_n378_4[2]),.dinb(w_G351_2[1]),.dout(n379),.clk(gclk));
	jor g0079(.dina(n379),.dinb(w_n377_1[1]),.dout(n380),.clk(gclk));
	jor g0080(.dina(n380),.dinb(n376),.dout(n381),.clk(gclk));
	jand g0081(.dina(w_G3546_5[0]),.dinb(w_G351_2[0]),.dout(n382),.clk(gclk));
	jand g0082(.dina(w_G3548_4[2]),.dinb(w_n374_1[0]),.dout(n383),.clk(gclk));
	jor g0083(.dina(n383),.dinb(n382),.dout(n384),.clk(gclk));
	jor g0084(.dina(n384),.dinb(w_G534_2[0]),.dout(n385),.clk(gclk));
	jand g0085(.dina(n385),.dinb(n381),.dout(n386),.clk(gclk));
	jnot g0086(.din(w_G341_2[2]),.dout(n387),.clk(gclk));
	jand g0087(.dina(w_n375_4[1]),.dinb(w_n387_1[1]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G523_1[2]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n378_4[1]),.dinb(w_G341_2[1]),.dout(n390),.clk(gclk));
	jor g0090(.dina(n390),.dinb(w_n389_1[1]),.dout(n391),.clk(gclk));
	jor g0091(.dina(n391),.dinb(n388),.dout(n392),.clk(gclk));
	jand g0092(.dina(w_G3546_4[2]),.dinb(w_G341_2[0]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3548_4[1]),.dinb(w_n387_1[0]),.dout(n394),.clk(gclk));
	jor g0094(.dina(n394),.dinb(n393),.dout(n395),.clk(gclk));
	jor g0095(.dina(n395),.dinb(w_G523_1[1]),.dout(n396),.clk(gclk));
	jand g0096(.dina(n396),.dinb(n392),.dout(n397),.clk(gclk));
	jand g0097(.dina(w_n397_0[1]),.dinb(w_n386_0[1]),.dout(n398),.clk(gclk));
	jand g0098(.dina(n398),.dinb(n373),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G316_1[1]),.dinb(w_G248_5[1]),.dout(n400),.clk(gclk));
	jnot g0100(.din(w_G490_1[1]),.dout(n401),.clk(gclk));
	jnot g0101(.din(w_G316_1[0]),.dout(n402),.clk(gclk));
	jand g0102(.dina(w_n402_0[2]),.dinb(w_G251_5[0]),.dout(n403),.clk(gclk));
	jor g0103(.dina(n403),.dinb(w_n401_0[1]),.dout(n404),.clk(gclk));
	jor g0104(.dina(n404),.dinb(n400),.dout(n405),.clk(gclk));
	jnot g0105(.din(w_G254_1[1]),.dout(n406),.clk(gclk));
	jand g0106(.dina(w_n402_0[1]),.dinb(w_n406_5[1]),.dout(n407),.clk(gclk));
	jnot g0107(.din(w_G242_1[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_G316_0[2]),.dinb(w_n408_5[2]),.dout(n409),.clk(gclk));
	jor g0109(.dina(n409),.dinb(n407),.dout(n410),.clk(gclk));
	jor g0110(.dina(n410),.dinb(w_G490_1[0]),.dout(n411),.clk(gclk));
	jand g0111(.dina(n411),.dinb(n405),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G308_1[2]),.dinb(w_G248_5[0]),.dout(n413),.clk(gclk));
	jnot g0113(.din(w_G479_0[2]),.dout(n414),.clk(gclk));
	jnot g0114(.din(w_G308_1[1]),.dout(n415),.clk(gclk));
	jand g0115(.dina(w_n415_0[1]),.dinb(w_G251_4[2]),.dout(n416),.clk(gclk));
	jor g0116(.dina(n416),.dinb(w_n414_0[1]),.dout(n417),.clk(gclk));
	jor g0117(.dina(n417),.dinb(n413),.dout(n418),.clk(gclk));
	jand g0118(.dina(w_n415_0[0]),.dinb(w_n406_5[0]),.dout(n419),.clk(gclk));
	jand g0119(.dina(w_G308_1[0]),.dinb(w_n408_5[1]),.dout(n420),.clk(gclk));
	jor g0120(.dina(n420),.dinb(n419),.dout(n421),.clk(gclk));
	jor g0121(.dina(n421),.dinb(w_G479_0[1]),.dout(n422),.clk(gclk));
	jand g0122(.dina(n422),.dinb(n418),.dout(n423),.clk(gclk));
	jand g0123(.dina(w_n423_0[2]),.dinb(w_n412_0[2]),.dout(n424),.clk(gclk));
	jnot g0124(.din(w_G293_0[2]),.dout(n425),.clk(gclk));
	jand g0125(.dina(w_n425_0[2]),.dinb(w_n406_4[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_G293_0[1]),.dinb(w_n408_5[0]),.dout(n427),.clk(gclk));
	jor g0127(.dina(n427),.dinb(n426),.dout(n428),.clk(gclk));
	jnot g0128(.din(w_G302_0[2]),.dout(n429),.clk(gclk));
	jand g0129(.dina(w_n429_0[1]),.dinb(w_n366_1[1]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G302_0[1]),.dinb(w_n369_1[1]),.dout(n431),.clk(gclk));
	jor g0131(.dina(n431),.dinb(n430),.dout(n432),.clk(gclk));
	jnot g0132(.din(n432),.dout(n433),.clk(gclk));
	jand g0133(.dina(w_n433_0[2]),.dinb(w_n428_1[1]),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G324_1[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n375_4[0]),.dinb(w_n435_2[1]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G503_2[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n378_4[0]),.dinb(w_G324_1[1]),.dout(n438),.clk(gclk));
	jor g0138(.dina(n438),.dinb(w_n437_0[1]),.dout(n439),.clk(gclk));
	jor g0139(.dina(n439),.dinb(n436),.dout(n440),.clk(gclk));
	jand g0140(.dina(w_G3546_4[1]),.dinb(w_G324_1[0]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3548_4[0]),.dinb(w_n435_2[0]),.dout(n442),.clk(gclk));
	jor g0142(.dina(n442),.dinb(n441),.dout(n443),.clk(gclk));
	jor g0143(.dina(n443),.dinb(w_G503_2[0]),.dout(n444),.clk(gclk));
	jand g0144(.dina(n444),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(n434),.dout(n446),.clk(gclk));
	jand g0146(.dina(n446),.dinb(n424),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(n399),.dout(w_dff_A_mkTkpc2K4_2),.clk(gclk));
	jnot g0148(.din(w_G210_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n375_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G457_1[2]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n378_3[2]),.dinb(w_G210_2[0]),.dout(n452),.clk(gclk));
	jor g0152(.dina(n452),.dinb(w_n451_0[2]),.dout(n453),.clk(gclk));
	jor g0153(.dina(n453),.dinb(n450),.dout(n454),.clk(gclk));
	jand g0154(.dina(w_G3546_4[0]),.dinb(w_G210_1[2]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n456),.clk(gclk));
	jor g0156(.dina(n456),.dinb(n455),.dout(n457),.clk(gclk));
	jor g0157(.dina(n457),.dinb(w_G457_1[1]),.dout(n458),.clk(gclk));
	jand g0158(.dina(n458),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n375_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n378_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jor g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464),.clk(gclk));
	jor g0164(.dina(n464),.dinb(n461),.dout(n465),.clk(gclk));
	jand g0165(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n467),.clk(gclk));
	jor g0167(.dina(n467),.dinb(n466),.dout(n468),.clk(gclk));
	jor g0168(.dina(n468),.dinb(w_G435_1[1]),.dout(n469),.clk(gclk));
	jand g0169(.dina(n469),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G273_2[1]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n375_3[0]),.dinb(w_n471_1[2]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G411_2[1]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n378_3[0]),.dinb(w_G273_2[0]),.dout(n474),.clk(gclk));
	jor g0174(.dina(n474),.dinb(w_n473_1[1]),.dout(n475),.clk(gclk));
	jor g0175(.dina(n475),.dinb(n472),.dout(n476),.clk(gclk));
	jand g0176(.dina(w_G3546_3[1]),.dinb(w_G273_1[2]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3548_3[0]),.dinb(w_n471_1[1]),.dout(n478),.clk(gclk));
	jor g0178(.dina(n478),.dinb(n477),.dout(n479),.clk(gclk));
	jor g0179(.dina(n479),.dinb(w_G411_2[0]),.dout(n480),.clk(gclk));
	jand g0180(.dina(n480),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jnot g0182(.din(w_G265_1[2]),.dout(n483),.clk(gclk));
	jand g0183(.dina(w_n375_2[2]),.dinb(w_n483_2[1]),.dout(n484),.clk(gclk));
	jnot g0184(.din(w_G400_1[2]),.dout(n485),.clk(gclk));
	jand g0185(.dina(w_n378_2[2]),.dinb(w_G265_1[1]),.dout(n486),.clk(gclk));
	jor g0186(.dina(n486),.dinb(w_n485_1[1]),.dout(n487),.clk(gclk));
	jor g0187(.dina(n487),.dinb(n484),.dout(n488),.clk(gclk));
	jand g0188(.dina(w_G3546_3[0]),.dinb(w_G265_1[0]),.dout(n489),.clk(gclk));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n483_2[0]),.dout(n490),.clk(gclk));
	jor g0190(.dina(n490),.dinb(n489),.dout(n491),.clk(gclk));
	jor g0191(.dina(n491),.dinb(w_G400_1[1]),.dout(n492),.clk(gclk));
	jand g0192(.dina(n492),.dinb(n488),.dout(n493),.clk(gclk));
	jnot g0193(.din(w_G226_2[1]),.dout(n494),.clk(gclk));
	jand g0194(.dina(w_n375_2[1]),.dinb(w_n494_1[2]),.dout(n495),.clk(gclk));
	jnot g0195(.din(w_G422_1[1]),.dout(n496),.clk(gclk));
	jand g0196(.dina(w_n378_2[1]),.dinb(w_G226_2[0]),.dout(n497),.clk(gclk));
	jor g0197(.dina(n497),.dinb(w_n496_1[1]),.dout(n498),.clk(gclk));
	jor g0198(.dina(n498),.dinb(n495),.dout(n499),.clk(gclk));
	jand g0199(.dina(w_G3546_2[2]),.dinb(w_G226_1[2]),.dout(n500),.clk(gclk));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n494_1[1]),.dout(n501),.clk(gclk));
	jor g0201(.dina(n501),.dinb(n500),.dout(n502),.clk(gclk));
	jor g0202(.dina(n502),.dinb(w_G422_1[0]),.dout(n503),.clk(gclk));
	jand g0203(.dina(n503),.dinb(n499),.dout(n504),.clk(gclk));
	jand g0204(.dina(w_n504_0[1]),.dinb(w_n493_0[1]),.dout(n505),.clk(gclk));
	jand g0205(.dina(n505),.dinb(n482),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[1]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n375_2[0]),.dinb(w_n507_1[2]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n378_2[0]),.dinb(w_G218_2[0]),.dout(n510),.clk(gclk));
	jor g0210(.dina(n510),.dinb(w_n509_0[2]),.dout(n511),.clk(gclk));
	jor g0211(.dina(n511),.dinb(n508),.dout(n512),.clk(gclk));
	jand g0212(.dina(w_G3546_2[1]),.dinb(w_G218_1[2]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3548_2[0]),.dinb(w_n507_1[1]),.dout(n514),.clk(gclk));
	jor g0214(.dina(n514),.dinb(n513),.dout(n515),.clk(gclk));
	jor g0215(.dina(n515),.dinb(w_G468_1[1]),.dout(n516),.clk(gclk));
	jand g0216(.dina(n516),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G257_2[1]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_n375_1[2]),.dinb(w_n518_1[2]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G389_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_n378_1[2]),.dinb(w_G257_2[0]),.dout(n521),.clk(gclk));
	jor g0221(.dina(n521),.dinb(w_n520_0[2]),.dout(n522),.clk(gclk));
	jor g0222(.dina(n522),.dinb(n519),.dout(n523),.clk(gclk));
	jand g0223(.dina(w_G3546_2[0]),.dinb(w_G257_1[2]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_G3548_1[2]),.dinb(w_n518_1[1]),.dout(n525),.clk(gclk));
	jor g0225(.dina(n525),.dinb(n524),.dout(n526),.clk(gclk));
	jor g0226(.dina(n526),.dinb(w_G389_1[1]),.dout(n527),.clk(gclk));
	jand g0227(.dina(n527),.dinb(n523),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[1]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G281_2[1]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n375_1[1]),.dinb(w_n530_1[2]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G374_1[2]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n378_1[1]),.dinb(w_G281_2[0]),.dout(n533),.clk(gclk));
	jor g0233(.dina(n533),.dinb(w_n532_1[1]),.dout(n534),.clk(gclk));
	jor g0234(.dina(n534),.dinb(n531),.dout(n535),.clk(gclk));
	jand g0235(.dina(w_G3546_1[2]),.dinb(w_G281_1[2]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3548_1[1]),.dinb(w_n530_1[1]),.dout(n537),.clk(gclk));
	jor g0237(.dina(n537),.dinb(n536),.dout(n538),.clk(gclk));
	jor g0238(.dina(n538),.dinb(w_G374_1[1]),.dout(n539),.clk(gclk));
	jand g0239(.dina(n539),.dinb(n535),.dout(n540),.clk(gclk));
	jand g0240(.dina(w_G248_4[2]),.dinb(w_G206_1[2]),.dout(n541),.clk(gclk));
	jnot g0241(.din(w_G446_1[2]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G206_1[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_G251_4[1]),.dinb(w_n543_0[1]),.dout(n544),.clk(gclk));
	jor g0244(.dina(n544),.dinb(n542),.dout(n545),.clk(gclk));
	jor g0245(.dina(n545),.dinb(n541),.dout(n546),.clk(gclk));
	jand g0246(.dina(w_n406_4[1]),.dinb(w_n543_0[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_n408_4[2]),.dinb(w_G206_1[0]),.dout(n548),.clk(gclk));
	jor g0248(.dina(n548),.dinb(n547),.dout(n549),.clk(gclk));
	jor g0249(.dina(n549),.dinb(w_G446_1[1]),.dout(n550),.clk(gclk));
	jand g0250(.dina(n550),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[2]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(n506),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_n459_0[1]),.dout(w_dff_A_kiJeiQer6_2),.clk(gclk));
	jnot g0255(.din(w_G335_0[2]),.dout(n556),.clk(gclk));
	jand g0256(.dina(w_n556_8[1]),.dinb(w_n530_1[0]),.dout(n557),.clk(gclk));
	jnot g0257(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jor g0258(.dina(w_n556_8[0]),.dinb(G288),.dout(n559),.clk(gclk));
	jand g0259(.dina(w_n559_0[1]),.dinb(n558),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_0[2]),.dinb(w_G374_1[0]),.dout(n561),.clk(gclk));
	jand g0261(.dina(w_n556_7[2]),.dinb(w_n471_1[0]),.dout(n562),.clk(gclk));
	jnot g0262(.din(w_n562_0[1]),.dout(n563),.clk(gclk));
	jor g0263(.dina(w_n556_7[1]),.dinb(G280),.dout(n564),.clk(gclk));
	jand g0264(.dina(w_n564_0[1]),.dinb(n563),.dout(n565),.clk(gclk));
	jxor g0265(.dina(w_n565_0[2]),.dinb(w_G411_1[2]),.dout(n566),.clk(gclk));
	jand g0266(.dina(w_n566_0[2]),.dinb(w_n561_1[1]),.dout(n567),.clk(gclk));
	jnot g0267(.din(w_n567_0[2]),.dout(n568),.clk(gclk));
	jand g0268(.dina(w_n556_7[0]),.dinb(w_n483_1[2]),.dout(n569),.clk(gclk));
	jnot g0269(.din(w_n569_0[1]),.dout(n570),.clk(gclk));
	jor g0270(.dina(w_n556_6[2]),.dinb(G272),.dout(n571),.clk(gclk));
	jand g0271(.dina(w_n571_0[1]),.dinb(n570),.dout(n572),.clk(gclk));
	jxor g0272(.dina(w_n572_0[2]),.dinb(w_G400_1[0]),.dout(n573),.clk(gclk));
	jnot g0273(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jand g0274(.dina(w_n556_6[1]),.dinb(w_n518_1[0]),.dout(n575),.clk(gclk));
	jnot g0275(.din(n575),.dout(n576),.clk(gclk));
	jor g0276(.dina(w_n556_6[0]),.dinb(G264),.dout(n577),.clk(gclk));
	jand g0277(.dina(n577),.dinb(n576),.dout(n578),.clk(gclk));
	jxor g0278(.dina(w_n578_1[1]),.dinb(w_n520_0[1]),.dout(n579),.clk(gclk));
	jor g0279(.dina(w_n579_1[1]),.dinb(w_n574_0[2]),.dout(n580),.clk(gclk));
	jor g0280(.dina(n580),.dinb(n568),.dout(n581),.clk(gclk));
	jnot g0281(.din(w_n581_0[1]),.dout(n582),.clk(gclk));
	jand g0282(.dina(w_n556_5[2]),.dinb(w_n460_1[0]),.dout(n583),.clk(gclk));
	jnot g0283(.din(n583),.dout(n584),.clk(gclk));
	jor g0284(.dina(w_n556_5[1]),.dinb(G241),.dout(n585),.clk(gclk));
	jand g0285(.dina(n585),.dinb(n584),.dout(n586),.clk(gclk));
	jxor g0286(.dina(w_n586_1[1]),.dinb(w_G435_1[0]),.dout(n587),.clk(gclk));
	jand g0287(.dina(w_n587_0[1]),.dinb(n582),.dout(n588),.clk(gclk));
	jor g0288(.dina(w_G335_0[1]),.dinb(w_G206_0[2]),.dout(n589),.clk(gclk));
	jor g0289(.dina(w_n556_5[0]),.dinb(G209),.dout(n590),.clk(gclk));
	jand g0290(.dina(n590),.dinb(n589),.dout(n591),.clk(gclk));
	jxor g0291(.dina(w_n591_1[1]),.dinb(w_G446_1[0]),.dout(n592),.clk(gclk));
	jand g0292(.dina(w_n556_4[2]),.dinb(w_n494_1[0]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jor g0294(.dina(w_n556_4[1]),.dinb(G233),.dout(n595),.clk(gclk));
	jand g0295(.dina(n595),.dinb(n594),.dout(n596),.clk(gclk));
	jxor g0296(.dina(w_n596_1[1]),.dinb(w_n496_1[0]),.dout(n597),.clk(gclk));
	jand g0297(.dina(w_n556_4[0]),.dinb(w_n507_1[0]),.dout(n598),.clk(gclk));
	jnot g0298(.din(n598),.dout(n599),.clk(gclk));
	jor g0299(.dina(w_n556_3[2]),.dinb(G225),.dout(n600),.clk(gclk));
	jand g0300(.dina(n600),.dinb(n599),.dout(n601),.clk(gclk));
	jxor g0301(.dina(w_n601_1[1]),.dinb(w_n509_0[1]),.dout(n602),.clk(gclk));
	jor g0302(.dina(w_n602_0[2]),.dinb(w_n597_0[2]),.dout(n603),.clk(gclk));
	jand g0303(.dina(w_n556_3[1]),.dinb(w_n449_1[0]),.dout(n604),.clk(gclk));
	jnot g0304(.din(n604),.dout(n605),.clk(gclk));
	jor g0305(.dina(w_n556_3[0]),.dinb(G217),.dout(n606),.clk(gclk));
	jand g0306(.dina(n606),.dinb(n605),.dout(n607),.clk(gclk));
	jxor g0307(.dina(w_n607_1[1]),.dinb(w_n451_0[1]),.dout(n608),.clk(gclk));
	jor g0308(.dina(w_n608_0[2]),.dinb(w_n603_0[1]),.dout(n609),.clk(gclk));
	jnot g0309(.din(w_n609_0[2]),.dout(n610),.clk(gclk));
	jand g0310(.dina(n610),.dinb(w_n592_0[2]),.dout(n611),.clk(gclk));
	jand g0311(.dina(w_n611_0[2]),.dinb(w_n588_1[1]),.dout(w_dff_A_1Y5z3GHA5_2),.clk(gclk));
	jnot g0312(.din(w_G332_3[2]),.dout(n613),.clk(gclk));
	jand g0313(.dina(w_n613_5[2]),.dinb(w_n435_1[2]),.dout(n614),.clk(gclk));
	jnot g0314(.din(n614),.dout(n615),.clk(gclk));
	jor g0315(.dina(w_n613_5[1]),.dinb(w_G331_0[1]),.dout(n616),.clk(gclk));
	jand g0316(.dina(n616),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_G503_1[2]),.dout(n618),.clk(gclk));
	jor g0318(.dina(w_G338_0[0]),.dinb(w_n613_5[0]),.dout(n619),.clk(gclk));
	jxor g0319(.dina(w_n619_1[2]),.dinb(w_G514_1[2]),.dout(n620),.clk(gclk));
	jor g0320(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n621),.clk(gclk));
	jor g0321(.dina(w_G348_0[0]),.dinb(w_n613_4[2]),.dout(n622),.clk(gclk));
	jand g0322(.dina(n622),.dinb(w_n621_0[1]),.dout(n623),.clk(gclk));
	jxor g0323(.dina(w_n623_0[1]),.dinb(w_G523_1[0]),.dout(n624),.clk(gclk));
	jor g0324(.dina(w_G351_1[2]),.dinb(w_G332_3[0]),.dout(n625),.clk(gclk));
	jor g0325(.dina(w_G358_0[0]),.dinb(w_n613_4[1]),.dout(n626),.clk(gclk));
	jand g0326(.dina(n626),.dinb(w_n625_0[1]),.dout(n627),.clk(gclk));
	jor g0327(.dina(w_n627_1[1]),.dinb(w_G534_1[2]),.dout(n628),.clk(gclk));
	jnot g0328(.din(w_n625_0[0]),.dout(n629),.clk(gclk));
	jand g0329(.dina(w_G612_0),.dinb(w_G332_2[2]),.dout(n630),.clk(gclk));
	jor g0330(.dina(n630),.dinb(n629),.dout(n631),.clk(gclk));
	jor g0331(.dina(w_n631_0[1]),.dinb(w_n377_1[0]),.dout(n632),.clk(gclk));
	jor g0332(.dina(w_G361_0[2]),.dinb(w_G332_2[1]),.dout(n633),.clk(gclk));
	jor g0333(.dina(w_G366_0[0]),.dinb(w_n613_4[0]),.dout(n634),.clk(gclk));
	jand g0334(.dina(n634),.dinb(n633),.dout(n635),.clk(gclk));
	jnot g0335(.din(w_n635_1[1]),.dout(n636),.clk(gclk));
	jand g0336(.dina(w_n636_0[2]),.dinb(w_n632_0[1]),.dout(n637),.clk(gclk));
	jand g0337(.dina(w_n637_0[2]),.dinb(w_n628_0[2]),.dout(n638),.clk(gclk));
	jand g0338(.dina(w_n638_0[1]),.dinb(w_n624_0[2]),.dout(n639),.clk(gclk));
	jand g0339(.dina(w_n639_0[2]),.dinb(w_n620_1[1]),.dout(n640),.clk(gclk));
	jand g0340(.dina(w_n640_0[1]),.dinb(w_n618_0[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n613_3[2]),.dinb(w_n425_0[1]),.dout(n642),.clk(gclk));
	jand g0342(.dina(w_G332_2[0]),.dinb(w_G593_0),.dout(n643),.clk(gclk));
	jor g0343(.dina(n643),.dinb(n642),.dout(n644),.clk(gclk));
	jand g0344(.dina(w_n613_3[1]),.dinb(w_n429_0[0]),.dout(n645),.clk(gclk));
	jnot g0345(.din(n645),.dout(n646),.clk(gclk));
	jor g0346(.dina(w_n613_3[0]),.dinb(G307),.dout(n647),.clk(gclk));
	jand g0347(.dina(n647),.dinb(n646),.dout(n648),.clk(gclk));
	jnot g0348(.din(w_n648_1[1]),.dout(n649),.clk(gclk));
	jand g0349(.dina(w_n649_0[1]),.dinb(w_n644_0[2]),.dout(n650),.clk(gclk));
	jor g0350(.dina(w_G332_1[2]),.dinb(w_G308_0[2]),.dout(n651),.clk(gclk));
	jor g0351(.dina(w_n613_2[2]),.dinb(G315),.dout(n652),.clk(gclk));
	jand g0352(.dina(n652),.dinb(n651),.dout(n653),.clk(gclk));
	jxor g0353(.dina(w_n653_0[2]),.dinb(w_G479_0[0]),.dout(n654),.clk(gclk));
	jand g0354(.dina(w_n613_2[1]),.dinb(w_n402_0[0]),.dout(n655),.clk(gclk));
	jnot g0355(.din(n655),.dout(n656),.clk(gclk));
	jor g0356(.dina(w_n613_2[0]),.dinb(G323),.dout(n657),.clk(gclk));
	jand g0357(.dina(n657),.dinb(n656),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_n658_1[1]),.dinb(w_G490_0[2]),.dout(n659),.clk(gclk));
	jand g0359(.dina(w_n659_0[1]),.dinb(w_n654_2[2]),.dout(n660),.clk(gclk));
	jand g0360(.dina(w_n660_1[1]),.dinb(w_n650_0[1]),.dout(n661),.clk(gclk));
	jand g0361(.dina(w_n661_0[1]),.dinb(w_n641_1[2]),.dout(w_dff_A_1RVBZJEC9_2),.clk(gclk));
	jxor g0362(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G302_0[0]),.dinb(w_n425_0[0]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(n663),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G369_0[1]),.dinb(w_G361_0[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(n666),.dinb(w_n435_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n668),.clk(gclk));
	jxor g0368(.dina(n668),.dinb(n667),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n665),.dout(n670),.clk(gclk));
	jnot g0370(.din(w_n670_0[1]),.dout(w_dff_A_jl9DVvEN6_1),.clk(gclk));
	jxor g0371(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n672),.clk(gclk));
	jxor g0372(.dina(w_G273_1[1]),.dinb(w_n483_1[1]),.dout(n673),.clk(gclk));
	jxor g0373(.dina(n673),.dinb(n672),.dout(n674),.clk(gclk));
	jxor g0374(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n675),.clk(gclk));
	jxor g0375(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n676),.clk(gclk));
	jxor g0376(.dina(n676),.dinb(n675),.dout(n677),.clk(gclk));
	jxor g0377(.dina(w_G210_1[1]),.dinb(w_G206_0[1]),.dout(n678),.clk(gclk));
	jxor g0378(.dina(n678),.dinb(n677),.dout(n679),.clk(gclk));
	jxor g0379(.dina(n679),.dinb(n674),.dout(n680),.clk(gclk));
	jnot g0380(.din(w_n680_0[1]),.dout(w_dff_A_9BfOiUdX0_1),.clk(gclk));
	jand g0381(.dina(w_n586_1[0]),.dinb(w_G435_0[2]),.dout(n682),.clk(gclk));
	jnot g0382(.din(w_n586_0[2]),.dout(n683),.clk(gclk));
	jand g0383(.dina(n683),.dinb(w_n462_0[1]),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n684_0[1]),.dout(n685),.clk(gclk));
	jand g0385(.dina(w_n578_1[0]),.dinb(w_G389_1[0]),.dout(n686),.clk(gclk));
	jor g0386(.dina(w_n578_0[2]),.dinb(w_G389_0[2]),.dout(n687),.clk(gclk));
	jnot g0387(.din(w_n571_0[0]),.dout(n688),.clk(gclk));
	jor g0388(.dina(n688),.dinb(w_n569_0[0]),.dout(n689),.clk(gclk));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n485_1[0]),.dout(n690),.clk(gclk));
	jnot g0390(.din(w_n690_0[1]),.dout(n691),.clk(gclk));
	jand g0391(.dina(w_n560_0[1]),.dinb(w_G374_0[2]),.dout(n692),.clk(gclk));
	jor g0392(.dina(w_n565_0[1]),.dinb(w_G411_1[1]),.dout(n693),.clk(gclk));
	jand g0393(.dina(n693),.dinb(w_n692_0[1]),.dout(n694),.clk(gclk));
	jand g0394(.dina(w_n565_0[0]),.dinb(w_G411_1[0]),.dout(n695),.clk(gclk));
	jand g0395(.dina(w_n572_0[1]),.dinb(w_G400_0[2]),.dout(n696),.clk(gclk));
	jor g0396(.dina(n696),.dinb(w_n695_0[2]),.dout(n697),.clk(gclk));
	jor g0397(.dina(n697),.dinb(w_n694_0[2]),.dout(n698),.clk(gclk));
	jand g0398(.dina(n698),.dinb(n691),.dout(n699),.clk(gclk));
	jand g0399(.dina(w_n699_0[2]),.dinb(w_n687_0[1]),.dout(n700),.clk(gclk));
	jor g0400(.dina(n700),.dinb(w_n686_0[1]),.dout(n701),.clk(gclk));
	jand g0401(.dina(w_n701_0[1]),.dinb(w_n685_0[1]),.dout(n702),.clk(gclk));
	jor g0402(.dina(n702),.dinb(w_n682_0[2]),.dout(n703),.clk(gclk));
	jand g0403(.dina(w_n703_0[2]),.dinb(w_n611_0[1]),.dout(n704),.clk(gclk));
	jand g0404(.dina(w_n591_1[0]),.dinb(w_G446_0[2]),.dout(n705),.clk(gclk));
	jor g0405(.dina(w_n591_0[2]),.dinb(w_G446_0[1]),.dout(n706),.clk(gclk));
	jand g0406(.dina(w_n607_1[0]),.dinb(w_G457_1[0]),.dout(n707),.clk(gclk));
	jor g0407(.dina(w_n607_0[2]),.dinb(w_G457_0[2]),.dout(n708),.clk(gclk));
	jand g0408(.dina(w_n601_1[0]),.dinb(w_G468_1[0]),.dout(n709),.clk(gclk));
	jand g0409(.dina(w_n596_1[0]),.dinb(w_G422_0[2]),.dout(n710),.clk(gclk));
	jor g0410(.dina(w_n601_0[2]),.dinb(w_G468_0[2]),.dout(n711),.clk(gclk));
	jand g0411(.dina(w_n711_0[1]),.dinb(w_n710_0[1]),.dout(n712),.clk(gclk));
	jor g0412(.dina(n712),.dinb(w_n709_0[1]),.dout(n713),.clk(gclk));
	jand g0413(.dina(w_n713_0[2]),.dinb(n708),.dout(n714),.clk(gclk));
	jor g0414(.dina(n714),.dinb(n707),.dout(n715),.clk(gclk));
	jand g0415(.dina(w_n715_0[2]),.dinb(n706),.dout(n716),.clk(gclk));
	jor g0416(.dina(n716),.dinb(n705),.dout(n717),.clk(gclk));
	jor g0417(.dina(w_n717_0[1]),.dinb(w_n704_0[1]),.dout(w_dff_A_SAvAS5ac4_2),.clk(gclk));
	jand g0418(.dina(w_n617_1[0]),.dinb(w_G503_1[1]),.dout(n719),.clk(gclk));
	jor g0419(.dina(w_n617_0[2]),.dinb(w_G503_1[0]),.dout(n720),.clk(gclk));
	jor g0420(.dina(w_n619_1[1]),.dinb(w_G514_1[1]),.dout(n721),.clk(gclk));
	jand g0421(.dina(w_n619_1[0]),.dinb(w_G514_1[0]),.dout(n722),.clk(gclk));
	jnot g0422(.din(w_n621_0[0]),.dout(n723),.clk(gclk));
	jand g0423(.dina(w_G599_0),.dinb(w_G332_1[1]),.dout(n724),.clk(gclk));
	jor g0424(.dina(n724),.dinb(n723),.dout(n725),.clk(gclk));
	jand g0425(.dina(w_n725_0[2]),.dinb(w_n389_1[0]),.dout(n726),.clk(gclk));
	jnot g0426(.din(w_n726_0[1]),.dout(n727),.clk(gclk));
	jand g0427(.dina(w_n635_1[0]),.dinb(w_n628_0[1]),.dout(n728),.clk(gclk));
	jand g0428(.dina(w_n623_0[0]),.dinb(w_G523_0[2]),.dout(n729),.clk(gclk));
	jand g0429(.dina(w_n627_1[0]),.dinb(w_G534_1[1]),.dout(n730),.clk(gclk));
	jor g0430(.dina(n730),.dinb(n729),.dout(n731),.clk(gclk));
	jor g0431(.dina(n731),.dinb(w_n728_0[1]),.dout(n732),.clk(gclk));
	jand g0432(.dina(n732),.dinb(w_dff_B_oSMEsVHY2_1),.dout(n733),.clk(gclk));
	jor g0433(.dina(w_n733_0[2]),.dinb(w_n722_0[1]),.dout(n734),.clk(gclk));
	jand g0434(.dina(n734),.dinb(w_n721_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[2]),.dinb(w_n720_0[1]),.dout(n736),.clk(gclk));
	jor g0436(.dina(n736),.dinb(w_n719_0[1]),.dout(n737),.clk(gclk));
	jand g0437(.dina(w_n737_1[1]),.dinb(w_n660_1[0]),.dout(n738),.clk(gclk));
	jnot g0438(.din(w_n650_0[0]),.dout(n739),.clk(gclk));
	jnot g0439(.din(w_n653_0[1]),.dout(n740),.clk(gclk));
	jor g0440(.dina(n740),.dinb(w_n414_0[0]),.dout(n741),.clk(gclk));
	jand g0441(.dina(w_n658_1[0]),.dinb(w_G490_0[1]),.dout(n742),.clk(gclk));
	jand g0442(.dina(w_n742_0[2]),.dinb(w_n654_2[1]),.dout(n743),.clk(gclk));
	jnot g0443(.din(n743),.dout(n744),.clk(gclk));
	jand g0444(.dina(n744),.dinb(n741),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_n745_0[1]),.dout(n746),.clk(gclk));
	jor g0446(.dina(w_n746_0[2]),.dinb(w_dff_B_nYAXIFgQ6_1),.dout(n747),.clk(gclk));
	jor g0447(.dina(w_n747_0[1]),.dinb(w_n738_0[1]),.dout(w_dff_A_GkJoW1s90_2),.clk(gclk));
	jnot g0448(.din(w_G4091_6[1]),.dout(n749),.clk(gclk));
	jand g0449(.dina(w_G4092_9[2]),.dinb(w_n749_13[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n750_8[2]),.dinb(G131),.dout(n751),.clk(gclk));
	jnot g0451(.din(n751),.dout(n752),.clk(gclk));
	jnot g0452(.din(w_G54_0[2]),.dout(n753),.clk(gclk));
	jxor g0453(.dina(w_n635_0[2]),.dinb(w_n753_1[1]),.dout(n754),.clk(gclk));
	jnot g0454(.din(n754),.dout(n755),.clk(gclk));
	jand g0455(.dina(w_n755_0[1]),.dinb(w_G4091_6[0]),.dout(n756),.clk(gclk));
	jand g0456(.dina(w_n372_0[0]),.dinb(w_n749_13[0]),.dout(n757),.clk(gclk));
	jor g0457(.dina(n757),.dinb(w_G4092_9[1]),.dout(n758),.clk(gclk));
	jor g0458(.dina(n758),.dinb(n756),.dout(n759),.clk(gclk));
	jand g0459(.dina(n759),.dinb(n752),.dout(G822_fa_),.clk(gclk));
	jand g0460(.dina(w_n750_8[1]),.dinb(G129),.dout(n761),.clk(gclk));
	jnot g0461(.din(n761),.dout(n762),.clk(gclk));
	jxor g0462(.dina(w_n627_0[2]),.dinb(w_G534_1[0]),.dout(n763),.clk(gclk));
	jnot g0463(.din(w_n763_0[2]),.dout(n764),.clk(gclk));
	jand g0464(.dina(n764),.dinb(w_n635_0[1]),.dout(n765),.clk(gclk));
	jor g0465(.dina(n765),.dinb(w_n638_0[0]),.dout(n766),.clk(gclk));
	jnot g0466(.din(n766),.dout(n767),.clk(gclk));
	jand g0467(.dina(w_n767_0[1]),.dinb(w_n753_1[0]),.dout(n768),.clk(gclk));
	jand g0468(.dina(w_n763_0[1]),.dinb(w_G54_0[1]),.dout(n769),.clk(gclk));
	jor g0469(.dina(w_dff_B_mqpqi7DM5_0),.dinb(n768),.dout(n770),.clk(gclk));
	jand g0470(.dina(n770),.dinb(w_G4091_5[2]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n386_0[0]),.dinb(w_n749_12[2]),.dout(n772),.clk(gclk));
	jor g0472(.dina(n772),.dinb(w_G4092_9[0]),.dout(n773),.clk(gclk));
	jor g0473(.dina(w_dff_B_gT4N4AbX2_0),.dinb(n771),.dout(n774),.clk(gclk));
	jand g0474(.dina(n774),.dinb(w_dff_B_1h6ymRVb5_1),.dout(G838_fa_),.clk(gclk));
	jand g0475(.dina(w_n750_8[0]),.dinb(G117),.dout(n776),.clk(gclk));
	jnot g0476(.din(n776),.dout(n777),.clk(gclk));
	jxor g0477(.dina(w_n561_1[0]),.dinb(w_G4_0[2]),.dout(n778),.clk(gclk));
	jnot g0478(.din(n778),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n779_0[1]),.dinb(w_G4091_5[1]),.dout(n780),.clk(gclk));
	jand g0480(.dina(w_n540_0[0]),.dinb(w_n749_12[1]),.dout(n781),.clk(gclk));
	jor g0481(.dina(n781),.dinb(w_G4092_8[2]),.dout(n782),.clk(gclk));
	jor g0482(.dina(n782),.dinb(n780),.dout(n783),.clk(gclk));
	jand g0483(.dina(n783),.dinb(n777),.dout(G861_fa_),.clk(gclk));
	jand g0484(.dina(w_n641_1[1]),.dinb(w_G54_0[0]),.dout(n785),.clk(gclk));
	jor g0485(.dina(w_dff_B_6f5qogMe0_0),.dinb(w_n737_1[0]),.dout(n786),.clk(gclk));
	jand g0486(.dina(w_n786_0[2]),.dinb(w_n660_0[2]),.dout(n787),.clk(gclk));
	jor g0487(.dina(n787),.dinb(w_n746_0[1]),.dout(n788),.clk(gclk));
	jnot g0488(.din(w_n788_0[2]),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n644_0[1]),.dout(n790),.clk(gclk));
	jxor g0490(.dina(w_n648_1[0]),.dinb(w_n790_0[2]),.dout(n791),.clk(gclk));
	jnot g0491(.din(n791),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_n792_0[2]),.dinb(n789),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n788_0[1]),.dinb(w_n790_0[1]),.dout(n794),.clk(gclk));
	jor g0494(.dina(w_dff_B_4xUKJLD13_0),.dinb(n793),.dout(n795),.clk(gclk));
	jnot g0495(.din(w_n795_1[1]),.dout(G623_fa_),.clk(gclk));
	jnot g0496(.din(w_G4088_9[2]),.dout(n797),.clk(gclk));
	jnot g0497(.din(w_G861_0),.dout(n798),.clk(gclk));
	jor g0498(.dina(w_n798_1[1]),.dinb(w_n797_9[1]),.dout(n799),.clk(gclk));
	jnot g0499(.din(w_G4087_4[2]),.dout(n800),.clk(gclk));
	jnot g0500(.din(w_G822_0),.dout(n801),.clk(gclk));
	jor g0501(.dina(w_n801_1[1]),.dinb(w_G4088_9[1]),.dout(n802),.clk(gclk));
	jand g0502(.dina(n802),.dinb(w_n800_4[1]),.dout(n803),.clk(gclk));
	jand g0503(.dina(w_dff_B_h0oYGuxO9_0),.dinb(n799),.dout(n804),.clk(gclk));
	jor g0504(.dina(w_n797_9[0]),.dinb(w_G61_0[1]),.dout(n805),.clk(gclk));
	jor g0505(.dina(w_G4088_9[0]),.dinb(w_G11_0[1]),.dout(n806),.clk(gclk));
	jand g0506(.dina(n806),.dinb(w_G4087_4[1]),.dout(n807),.clk(gclk));
	jand g0507(.dina(n807),.dinb(n805),.dout(n808),.clk(gclk));
	jor g0508(.dina(w_dff_B_sdoMaWUL3_0),.dinb(n804),.dout(w_dff_A_O7wYAVdt7_2),.clk(gclk));
	jand g0509(.dina(w_n750_7[2]),.dinb(G52),.dout(n810),.clk(gclk));
	jnot g0510(.din(n810),.dout(n811),.clk(gclk));
	jnot g0511(.din(w_n721_0[0]),.dout(n812),.clk(gclk));
	jnot g0512(.din(w_n722_0[0]),.dout(n813),.clk(gclk));
	jand g0513(.dina(w_n631_0[0]),.dinb(w_n377_0[2]),.dout(n814),.clk(gclk));
	jor g0514(.dina(w_n636_0[1]),.dinb(w_n814_0[2]),.dout(n815),.clk(gclk));
	jor g0515(.dina(w_n725_0[1]),.dinb(w_n389_0[2]),.dout(n816),.clk(gclk));
	jand g0516(.dina(w_n632_0[0]),.dinb(n816),.dout(n817),.clk(gclk));
	jand g0517(.dina(n817),.dinb(n815),.dout(n818),.clk(gclk));
	jor g0518(.dina(n818),.dinb(w_n726_0[0]),.dout(n819),.clk(gclk));
	jand g0519(.dina(w_n819_0[2]),.dinb(w_dff_B_wsuO4F6W8_1),.dout(n820),.clk(gclk));
	jor g0520(.dina(n820),.dinb(w_dff_B_okWyP26V2_1),.dout(n821),.clk(gclk));
	jnot g0521(.din(w_n620_1[0]),.dout(n822),.clk(gclk));
	jnot g0522(.din(w_n639_0[1]),.dout(n823),.clk(gclk));
	jor g0523(.dina(n823),.dinb(w_n753_0[2]),.dout(n824),.clk(gclk));
	jor g0524(.dina(w_n824_0[1]),.dinb(w_dff_B_JYWRbbI97_1),.dout(n825),.clk(gclk));
	jand g0525(.dina(n825),.dinb(w_n821_0[1]),.dout(n826),.clk(gclk));
	jxor g0526(.dina(n826),.dinb(w_n618_0[1]),.dout(n827),.clk(gclk));
	jand g0527(.dina(w_n827_0[1]),.dinb(w_G4091_5[0]),.dout(n828),.clk(gclk));
	jand g0528(.dina(w_n445_0[0]),.dinb(w_n749_12[0]),.dout(n829),.clk(gclk));
	jor g0529(.dina(n829),.dinb(w_G4092_8[1]),.dout(n830),.clk(gclk));
	jor g0530(.dina(w_dff_B_g4VSIKkr6_0),.dinb(n828),.dout(n831),.clk(gclk));
	jand g0531(.dina(n831),.dinb(w_dff_B_eluNYSm06_1),.dout(G832_fa_),.clk(gclk));
	jand g0532(.dina(w_n750_7[1]),.dinb(G130),.dout(n833),.clk(gclk));
	jnot g0533(.din(n833),.dout(n834),.clk(gclk));
	jand g0534(.dina(w_n824_0[0]),.dinb(w_n819_0[1]),.dout(n835),.clk(gclk));
	jxor g0535(.dina(n835),.dinb(w_n620_0[2]),.dout(n836),.clk(gclk));
	jand g0536(.dina(w_n836_0[1]),.dinb(w_G4091_4[2]),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_n365_0[0]),.dinb(w_n749_11[2]),.dout(n838),.clk(gclk));
	jor g0538(.dina(n838),.dinb(w_G4092_8[0]),.dout(n839),.clk(gclk));
	jor g0539(.dina(w_dff_B_2YSxb2fz8_0),.dinb(n837),.dout(n840),.clk(gclk));
	jand g0540(.dina(n840),.dinb(w_dff_B_b7l7TUX85_1),.dout(G834_fa_),.clk(gclk));
	jand g0541(.dina(w_n750_7[0]),.dinb(G119),.dout(n842),.clk(gclk));
	jnot g0542(.din(n842),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n397_0[0]),.dinb(w_n749_11[1]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_n637_0[1]),.dinb(w_n753_0[1]),.dout(n845),.clk(gclk));
	jor g0545(.dina(n845),.dinb(w_n814_0[1]),.dout(n846),.clk(gclk));
	jxor g0546(.dina(n846),.dinb(w_n624_0[1]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_0[1]),.dinb(w_G4091_4[1]),.dout(n848),.clk(gclk));
	jor g0548(.dina(n848),.dinb(w_G4092_7[2]),.dout(n849),.clk(gclk));
	jor g0549(.dina(n849),.dinb(w_dff_B_5z9KsX4z9_1),.dout(n850),.clk(gclk));
	jand g0550(.dina(n850),.dinb(w_dff_B_ZeJDghyp9_1),.dout(G836_fa_),.clk(gclk));
	jnot g0551(.din(w_G4089_9[2]),.dout(n852),.clk(gclk));
	jor g0552(.dina(w_n798_1[0]),.dinb(w_n852_9[1]),.dout(n853),.clk(gclk));
	jnot g0553(.din(w_G4090_4[2]),.dout(n854),.clk(gclk));
	jor g0554(.dina(w_n801_1[0]),.dinb(w_G4089_9[1]),.dout(n855),.clk(gclk));
	jand g0555(.dina(n855),.dinb(w_n854_4[1]),.dout(n856),.clk(gclk));
	jand g0556(.dina(w_dff_B_2QD7IzGH6_0),.dinb(n853),.dout(n857),.clk(gclk));
	jor g0557(.dina(w_n852_9[0]),.dinb(w_G61_0[0]),.dout(n858),.clk(gclk));
	jor g0558(.dina(w_G4089_9[0]),.dinb(w_G11_0[0]),.dout(n859),.clk(gclk));
	jand g0559(.dina(n859),.dinb(w_G4090_4[1]),.dout(n860),.clk(gclk));
	jand g0560(.dina(n860),.dinb(n858),.dout(n861),.clk(gclk));
	jor g0561(.dina(w_dff_B_VjAzt5NF2_0),.dinb(n857),.dout(w_dff_A_YcIv6Ant5_2),.clk(gclk));
	jand g0562(.dina(w_n750_6[2]),.dinb(G122),.dout(n863),.clk(gclk));
	jnot g0563(.din(n863),.dout(n864),.clk(gclk));
	jnot g0564(.din(w_n587_0[0]),.dout(n865),.clk(gclk));
	jnot g0565(.din(w_n579_1[0]),.dout(n866),.clk(gclk));
	jand g0566(.dina(w_n567_0[1]),.dinb(w_G4_0[1]),.dout(n867),.clk(gclk));
	jand g0567(.dina(w_n867_0[1]),.dinb(w_n573_0[1]),.dout(n868),.clk(gclk));
	jand g0568(.dina(w_n868_0[1]),.dinb(n866),.dout(n869),.clk(gclk));
	jor g0569(.dina(n869),.dinb(w_n701_0[0]),.dout(n870),.clk(gclk));
	jxor g0570(.dina(w_n870_0[1]),.dinb(w_n865_0[2]),.dout(n871),.clk(gclk));
	jand g0571(.dina(w_n871_0[1]),.dinb(w_G4091_4[0]),.dout(n872),.clk(gclk));
	jand g0572(.dina(w_n470_0[0]),.dinb(w_n749_11[0]),.dout(n873),.clk(gclk));
	jor g0573(.dina(n873),.dinb(w_G4092_7[1]),.dout(n874),.clk(gclk));
	jor g0574(.dina(n874),.dinb(n872),.dout(n875),.clk(gclk));
	jand g0575(.dina(n875),.dinb(n864),.dout(G871_fa_),.clk(gclk));
	jand g0576(.dina(w_n750_6[1]),.dinb(G128),.dout(n877),.clk(gclk));
	jnot g0577(.din(n877),.dout(n878),.clk(gclk));
	jor g0578(.dina(w_n868_0[0]),.dinb(w_n699_0[1]),.dout(n879),.clk(gclk));
	jxor g0579(.dina(n879),.dinb(w_n579_0[2]),.dout(n880),.clk(gclk));
	jand g0580(.dina(w_n880_0[1]),.dinb(w_G4091_3[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n528_0[0]),.dinb(w_n749_10[2]),.dout(n882),.clk(gclk));
	jor g0582(.dina(n882),.dinb(w_G4092_7[0]),.dout(n883),.clk(gclk));
	jor g0583(.dina(n883),.dinb(n881),.dout(n884),.clk(gclk));
	jand g0584(.dina(n884),.dinb(n878),.dout(G873_fa_),.clk(gclk));
	jand g0585(.dina(w_n750_6[0]),.dinb(G127),.dout(n886),.clk(gclk));
	jnot g0586(.din(n886),.dout(n887),.clk(gclk));
	jor g0587(.dina(w_n694_0[1]),.dinb(w_n695_0[1]),.dout(n888),.clk(gclk));
	jor g0588(.dina(n888),.dinb(w_n867_0[0]),.dout(n889),.clk(gclk));
	jxor g0589(.dina(n889),.dinb(w_n574_0[1]),.dout(n890),.clk(gclk));
	jand g0590(.dina(w_n890_0[1]),.dinb(w_G4091_3[1]),.dout(n891),.clk(gclk));
	jand g0591(.dina(w_n493_0[0]),.dinb(w_n749_10[1]),.dout(n892),.clk(gclk));
	jor g0592(.dina(n892),.dinb(w_G4092_6[2]),.dout(n893),.clk(gclk));
	jor g0593(.dina(n893),.dinb(n891),.dout(n894),.clk(gclk));
	jand g0594(.dina(n894),.dinb(n887),.dout(G875_fa_),.clk(gclk));
	jand g0595(.dina(w_n750_5[2]),.dinb(G126),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jnot g0597(.din(w_n566_0[1]),.dout(n898),.clk(gclk));
	jand g0598(.dina(w_n561_0[2]),.dinb(w_G4_0[0]),.dout(n899),.clk(gclk));
	jor g0599(.dina(n899),.dinb(w_n692_0[0]),.dout(n900),.clk(gclk));
	jxor g0600(.dina(n900),.dinb(n898),.dout(n901),.clk(gclk));
	jand g0601(.dina(w_n901_0[1]),.dinb(w_G4091_3[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_n481_0[0]),.dinb(w_n749_10[0]),.dout(n903),.clk(gclk));
	jor g0603(.dina(n903),.dinb(w_G4092_6[1]),.dout(n904),.clk(gclk));
	jor g0604(.dina(n904),.dinb(n902),.dout(n905),.clk(gclk));
	jand g0605(.dina(n905),.dinb(n897),.dout(G877_fa_),.clk(gclk));
	jnot g0606(.din(w_G331_0[0]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_n619_0[2]),.dout(n908),.clk(gclk));
	jand g0608(.dina(n908),.dinb(n907),.dout(n909),.clk(gclk));
	jand g0609(.dina(w_n619_0[1]),.dinb(w_n617_0[1]),.dout(n910),.clk(gclk));
	jor g0610(.dina(n910),.dinb(n909),.dout(n911),.clk(gclk));
	jxor g0611(.dina(n911),.dinb(w_n792_0[1]),.dout(n912),.clk(gclk));
	jor g0612(.dina(w_G369_0[0]),.dinb(w_G332_1[0]),.dout(n913),.clk(gclk));
	jor g0613(.dina(G372),.dinb(w_n613_1[2]),.dout(n914),.clk(gclk));
	jand g0614(.dina(n914),.dinb(n913),.dout(n915),.clk(gclk));
	jxor g0615(.dina(n915),.dinb(w_n636_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n627_0[1]),.dinb(w_n725_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(w_n658_0[2]),.dinb(w_n653_0[0]),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_dff_B_IjWP77AJ0_1),.dout(n919),.clk(gclk));
	jxor g0619(.dina(n919),.dinb(w_dff_B_GLcQe6Os9_1),.dout(n920),.clk(gclk));
	jxor g0620(.dina(n920),.dinb(n912),.dout(G998_fa_),.clk(gclk));
	jnot g0621(.din(w_n564_0[0]),.dout(n922),.clk(gclk));
	jor g0622(.dina(n922),.dinb(w_n562_0[0]),.dout(n923),.clk(gclk));
	jxor g0623(.dina(w_n578_0[1]),.dinb(w_n923_0[2]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n572_0[0]),.dinb(w_n560_0[0]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jor g0626(.dina(w_G335_0[0]),.dinb(w_G289_0[0]),.dout(n927),.clk(gclk));
	jor g0627(.dina(w_n556_2[2]),.dinb(G292),.dout(n928),.clk(gclk));
	jand g0628(.dina(n928),.dinb(n927),.dout(n929),.clk(gclk));
	jxor g0629(.dina(n929),.dinb(w_n591_0[1]),.dout(n930),.clk(gclk));
	jxor g0630(.dina(w_n596_0[2]),.dinb(w_n586_0[1]),.dout(n931),.clk(gclk));
	jxor g0631(.dina(w_n607_0[1]),.dinb(w_n601_0[1]),.dout(n932),.clk(gclk));
	jxor g0632(.dina(n932),.dinb(n931),.dout(n933),.clk(gclk));
	jxor g0633(.dina(n933),.dinb(n930),.dout(n934),.clk(gclk));
	jxor g0634(.dina(n934),.dinb(n926),.dout(n935),.clk(gclk));
	jnot g0635(.din(w_n935_0[1]),.dout(w_dff_A_LwGy0wKt8_1),.clk(gclk));
	jnot g0636(.din(w_n592_0[1]),.dout(n937),.clk(gclk));
	jnot g0637(.din(w_n715_0[1]),.dout(n938),.clk(gclk));
	jor g0638(.dina(w_n870_0[0]),.dinb(w_n682_0[1]),.dout(n939),.clk(gclk));
	jand g0639(.dina(n939),.dinb(w_n685_0[0]),.dout(n940),.clk(gclk));
	jnot g0640(.din(w_n940_1[1]),.dout(n941),.clk(gclk));
	jor g0641(.dina(n941),.dinb(w_n609_0[1]),.dout(n942),.clk(gclk));
	jand g0642(.dina(n942),.dinb(w_n938_0[2]),.dout(n943),.clk(gclk));
	jxor g0643(.dina(n943),.dinb(n937),.dout(n944),.clk(gclk));
	jnot g0644(.din(w_n944_0[1]),.dout(n945),.clk(gclk));
	jnot g0645(.din(w_n603_0[0]),.dout(n946),.clk(gclk));
	jand g0646(.dina(w_n940_1[0]),.dinb(n946),.dout(n947),.clk(gclk));
	jor g0647(.dina(n947),.dinb(w_n713_0[1]),.dout(n948),.clk(gclk));
	jxor g0648(.dina(n948),.dinb(w_n608_0[1]),.dout(n949),.clk(gclk));
	jand g0649(.dina(w_n949_0[1]),.dinb(n945),.dout(n950),.clk(gclk));
	jnot g0650(.din(w_n602_0[1]),.dout(n951),.clk(gclk));
	jnot g0651(.din(w_n596_0[1]),.dout(n952),.clk(gclk));
	jand g0652(.dina(n952),.dinb(w_n496_0[2]),.dout(n953),.clk(gclk));
	jnot g0653(.din(w_n953_0[1]),.dout(n954),.clk(gclk));
	jor g0654(.dina(w_n940_0[2]),.dinb(w_n710_0[0]),.dout(n955),.clk(gclk));
	jand g0655(.dina(n955),.dinb(w_n954_0[2]),.dout(n956),.clk(gclk));
	jxor g0656(.dina(n956),.dinb(n951),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n957_0[1]),.dout(n958),.clk(gclk));
	jand g0658(.dina(w_n890_0[0]),.dinb(w_n779_0[0]),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(w_n901_0[0]),.dout(n960),.clk(gclk));
	jand g0660(.dina(n960),.dinb(w_n871_0[0]),.dout(n961),.clk(gclk));
	jnot g0661(.din(w_n597_0[1]),.dout(n962),.clk(gclk));
	jxor g0662(.dina(w_n940_0[1]),.dinb(w_n962_0[1]),.dout(n963),.clk(gclk));
	jnot g0663(.din(n963),.dout(n964),.clk(gclk));
	jand g0664(.dina(w_n964_0[1]),.dinb(w_n880_0[0]),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(n961),.dout(n966),.clk(gclk));
	jand g0666(.dina(n966),.dinb(n958),.dout(n967),.clk(gclk));
	jand g0667(.dina(w_dff_B_e9C2TA1l0_0),.dinb(n950),.dout(w_dff_A_FSDJereM4_2),.clk(gclk));
	jxor g0668(.dina(w_n788_0[0]),.dinb(w_n649_0[0]),.dout(n969),.clk(gclk));
	jnot g0669(.din(w_n969_0[1]),.dout(n970),.clk(gclk));
	jand g0670(.dina(n970),.dinb(w_n755_0[0]),.dout(n971),.clk(gclk));
	jand g0671(.dina(w_n836_0[0]),.dinb(w_G623_0),.dout(n972),.clk(gclk));
	jand g0672(.dina(n972),.dinb(w_dff_B_7yMBzruG2_1),.dout(n973),.clk(gclk));
	jand g0673(.dina(w_n827_0[0]),.dinb(w_n763_0[0]),.dout(n974),.clk(gclk));
	jand g0674(.dina(n974),.dinb(w_n847_0[0]),.dout(n975),.clk(gclk));
	jnot g0675(.din(w_n658_0[1]),.dout(n976),.clk(gclk));
	jand g0676(.dina(n976),.dinb(w_n401_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(w_n977_0[2]),.dinb(w_n654_2[0]),.dout(n978),.clk(gclk));
	jor g0678(.dina(w_n977_0[1]),.dinb(w_n654_1[2]),.dout(n979),.clk(gclk));
	jnot g0679(.din(n979),.dout(n980),.clk(gclk));
	jor g0680(.dina(w_n786_0[1]),.dinb(w_n742_0[1]),.dout(n981),.clk(gclk));
	jand g0681(.dina(w_n981_0[1]),.dinb(w_dff_B_KtJt2y784_1),.dout(n982),.clk(gclk));
	jnot g0682(.din(w_n981_0[0]),.dout(n983),.clk(gclk));
	jand g0683(.dina(n983),.dinb(w_n654_1[1]),.dout(n984),.clk(gclk));
	jor g0684(.dina(n984),.dinb(w_dff_B_6pLzhFzy3_1),.dout(n985),.clk(gclk));
	jor g0685(.dina(n985),.dinb(w_dff_B_q3yblBT83_1),.dout(n986),.clk(gclk));
	jnot g0686(.din(w_n986_0[1]),.dout(n987),.clk(gclk));
	jnot g0687(.din(w_n659_0[0]),.dout(n988),.clk(gclk));
	jxor g0688(.dina(w_n786_0[0]),.dinb(w_dff_B_UILrsiJX5_1),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_n989_0[1]),.dinb(n987),.dout(n990),.clk(gclk));
	jand g0690(.dina(n990),.dinb(w_dff_B_thoFfn6c7_1),.dout(n991),.clk(gclk));
	jand g0691(.dina(n991),.dinb(n973),.dout(w_dff_A_5ltDjXuT8_2),.clk(gclk));
	jnot g0692(.din(w_G1689_5[1]),.dout(n993),.clk(gclk));
	jand g0693(.dina(w_G1690_1[1]),.dinb(w_n993_4[2]),.dout(n994),.clk(gclk));
	jand g0694(.dina(w_n994_4[1]),.dinb(w_G182_0[1]),.dout(n995),.clk(gclk));
	jand g0695(.dina(w_G1690_1[0]),.dinb(w_G1689_5[0]),.dout(n996),.clk(gclk));
	jand g0696(.dina(w_n996_4[1]),.dinb(w_G185_0[1]),.dout(n997),.clk(gclk));
	jor g0697(.dina(w_n798_0[2]),.dinb(w_n993_4[1]),.dout(n998),.clk(gclk));
	jnot g0698(.din(w_G1690_0[2]),.dout(n999),.clk(gclk));
	jor g0699(.dina(w_n801_0[2]),.dinb(w_G1689_4[2]),.dout(n1000),.clk(gclk));
	jand g0700(.dina(n1000),.dinb(w_n999_3[2]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_dff_B_rMnhefMo1_0),.dinb(n998),.dout(n1002),.clk(gclk));
	jor g0702(.dina(n1002),.dinb(w_dff_B_uHiqWlh60_1),.dout(n1003),.clk(gclk));
	jor g0703(.dina(n1003),.dinb(w_dff_B_MJIvSDTw3_1),.dout(n1004),.clk(gclk));
	jand g0704(.dina(n1004),.dinb(w_G137_9[1]),.dout(w_dff_A_09IHvNaL4_2),.clk(gclk));
	jor g0705(.dina(w_n801_0[1]),.dinb(w_G1691_5[1]),.dout(n1006),.clk(gclk));
	jnot g0706(.din(w_G1694_1[1]),.dout(n1007),.clk(gclk));
	jnot g0707(.din(w_G1691_5[0]),.dout(n1008),.clk(gclk));
	jor g0708(.dina(w_n798_0[1]),.dinb(w_n1008_4[2]),.dout(n1009),.clk(gclk));
	jand g0709(.dina(n1009),.dinb(w_n1007_3[2]),.dout(n1010),.clk(gclk));
	jand g0710(.dina(n1010),.dinb(w_dff_B_YZS4p8r72_1),.dout(n1011),.clk(gclk));
	jand g0711(.dina(w_G1694_1[0]),.dinb(w_G1691_4[2]),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_4[1]),.dinb(w_G185_0[0]),.dout(n1013),.clk(gclk));
	jand g0713(.dina(w_G1694_0[2]),.dinb(w_n1008_4[1]),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_4[1]),.dinb(w_G182_0[0]),.dout(n1015),.clk(gclk));
	jor g0715(.dina(n1015),.dinb(n1013),.dout(n1016),.clk(gclk));
	jor g0716(.dina(w_dff_B_bYh6fuTv8_0),.dinb(n1011),.dout(n1017),.clk(gclk));
	jand g0717(.dina(n1017),.dinb(w_G137_9[0]),.dout(w_dff_A_SWMAgAUJ9_2),.clk(gclk));
	jnot g0718(.din(w_G871_0),.dout(n1019),.clk(gclk));
	jor g0719(.dina(w_n1019_1[1]),.dinb(w_n797_8[2]),.dout(n1020),.clk(gclk));
	jnot g0720(.din(w_G832_0),.dout(n1021),.clk(gclk));
	jor g0721(.dina(w_n1021_1[1]),.dinb(w_G4088_8[2]),.dout(n1022),.clk(gclk));
	jand g0722(.dina(n1022),.dinb(w_n800_4[0]),.dout(n1023),.clk(gclk));
	jand g0723(.dina(n1023),.dinb(w_dff_B_TSxWOlHm2_1),.dout(n1024),.clk(gclk));
	jor g0724(.dina(w_n797_8[1]),.dinb(w_G37_0[1]),.dout(n1025),.clk(gclk));
	jor g0725(.dina(w_G4088_8[1]),.dinb(w_G43_0[1]),.dout(n1026),.clk(gclk));
	jand g0726(.dina(n1026),.dinb(w_G4087_4[0]),.dout(n1027),.clk(gclk));
	jand g0727(.dina(n1027),.dinb(n1025),.dout(n1028),.clk(gclk));
	jor g0728(.dina(w_dff_B_baGPJQFF2_0),.dinb(n1024),.dout(w_dff_A_Z13qQidg2_2),.clk(gclk));
	jnot g0729(.din(w_G873_0),.dout(n1030),.clk(gclk));
	jor g0730(.dina(w_n1030_1[1]),.dinb(w_n797_8[0]),.dout(n1031),.clk(gclk));
	jnot g0731(.din(w_G834_0),.dout(n1032),.clk(gclk));
	jor g0732(.dina(w_n1032_1[1]),.dinb(w_G4088_8[0]),.dout(n1033),.clk(gclk));
	jand g0733(.dina(n1033),.dinb(w_n800_3[2]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(n1034),.dinb(w_dff_B_Y8Qdl6VR9_1),.dout(n1035),.clk(gclk));
	jor g0735(.dina(w_n797_7[2]),.dinb(w_G20_0[1]),.dout(n1036),.clk(gclk));
	jor g0736(.dina(w_G4088_7[2]),.dinb(w_G76_0[1]),.dout(n1037),.clk(gclk));
	jand g0737(.dina(n1037),.dinb(w_G4087_3[2]),.dout(n1038),.clk(gclk));
	jand g0738(.dina(n1038),.dinb(n1036),.dout(n1039),.clk(gclk));
	jor g0739(.dina(w_dff_B_vsXxz3Ng1_0),.dinb(n1035),.dout(w_dff_A_NZTKntos3_2),.clk(gclk));
	jnot g0740(.din(w_G836_0),.dout(n1041),.clk(gclk));
	jor g0741(.dina(w_n1041_1[1]),.dinb(w_G4088_7[1]),.dout(n1042),.clk(gclk));
	jnot g0742(.din(w_G875_0),.dout(n1043),.clk(gclk));
	jor g0743(.dina(w_n1043_1[1]),.dinb(w_n797_7[1]),.dout(n1044),.clk(gclk));
	jand g0744(.dina(n1044),.dinb(w_n800_3[1]),.dout(n1045),.clk(gclk));
	jand g0745(.dina(n1045),.dinb(w_dff_B_8s8YOFXV9_1),.dout(n1046),.clk(gclk));
	jor g0746(.dina(w_n797_7[0]),.dinb(w_G17_0[1]),.dout(n1047),.clk(gclk));
	jor g0747(.dina(w_G4088_7[0]),.dinb(w_G73_0[1]),.dout(n1048),.clk(gclk));
	jand g0748(.dina(n1048),.dinb(w_G4087_3[1]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(n1049),.dinb(n1047),.dout(n1050),.clk(gclk));
	jor g0750(.dina(w_dff_B_D13BJunD9_0),.dinb(n1046),.dout(w_dff_A_qtJUbwCW9_2),.clk(gclk));
	jnot g0751(.din(w_G877_0),.dout(n1052),.clk(gclk));
	jor g0752(.dina(w_n1052_1[1]),.dinb(w_n797_6[2]),.dout(n1053),.clk(gclk));
	jnot g0753(.din(w_G838_0),.dout(n1054),.clk(gclk));
	jor g0754(.dina(w_n1054_1[1]),.dinb(w_G4088_6[2]),.dout(n1055),.clk(gclk));
	jand g0755(.dina(n1055),.dinb(w_n800_3[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(n1056),.dinb(w_dff_B_66V6EbF32_1),.dout(n1057),.clk(gclk));
	jor g0757(.dina(w_n797_6[1]),.dinb(w_G70_0[1]),.dout(n1058),.clk(gclk));
	jor g0758(.dina(w_G4088_6[1]),.dinb(w_G67_0[1]),.dout(n1059),.clk(gclk));
	jand g0759(.dina(n1059),.dinb(w_G4087_3[0]),.dout(n1060),.clk(gclk));
	jand g0760(.dina(n1060),.dinb(n1058),.dout(n1061),.clk(gclk));
	jor g0761(.dina(w_dff_B_TocnJ47N6_0),.dinb(n1057),.dout(w_dff_A_0IUNpq9e5_2),.clk(gclk));
	jor g0762(.dina(w_G4089_8[2]),.dinb(w_G43_0[0]),.dout(n1063),.clk(gclk));
	jor g0763(.dina(w_n852_8[2]),.dinb(w_G37_0[0]),.dout(n1064),.clk(gclk));
	jand g0764(.dina(n1064),.dinb(w_G4090_4[0]),.dout(n1065),.clk(gclk));
	jand g0765(.dina(n1065),.dinb(n1063),.dout(n1066),.clk(gclk));
	jor g0766(.dina(w_n1021_1[0]),.dinb(w_G4089_8[1]),.dout(n1067),.clk(gclk));
	jor g0767(.dina(w_n1019_1[0]),.dinb(w_n852_8[1]),.dout(n1068),.clk(gclk));
	jand g0768(.dina(n1068),.dinb(n1067),.dout(n1069),.clk(gclk));
	jand g0769(.dina(n1069),.dinb(w_n854_4[0]),.dout(n1070),.clk(gclk));
	jor g0770(.dina(n1070),.dinb(w_dff_B_0rAy1vbr2_1),.dout(w_dff_A_7okTC8Yv1_2),.clk(gclk));
	jor g0771(.dina(w_G4089_8[0]),.dinb(w_G76_0[0]),.dout(n1072),.clk(gclk));
	jor g0772(.dina(w_n852_8[0]),.dinb(w_G20_0[0]),.dout(n1073),.clk(gclk));
	jand g0773(.dina(n1073),.dinb(w_G4090_3[2]),.dout(n1074),.clk(gclk));
	jand g0774(.dina(n1074),.dinb(n1072),.dout(n1075),.clk(gclk));
	jor g0775(.dina(w_n1032_1[0]),.dinb(w_G4089_7[2]),.dout(n1076),.clk(gclk));
	jor g0776(.dina(w_n1030_1[0]),.dinb(w_n852_7[2]),.dout(n1077),.clk(gclk));
	jand g0777(.dina(w_dff_B_WtjqIDdJ3_0),.dinb(n1076),.dout(n1078),.clk(gclk));
	jand g0778(.dina(n1078),.dinb(w_n854_3[2]),.dout(n1079),.clk(gclk));
	jor g0779(.dina(n1079),.dinb(w_dff_B_WO2QjJZx1_1),.dout(w_dff_A_la5HpM0d0_2),.clk(gclk));
	jor g0780(.dina(w_G4089_7[1]),.dinb(w_G73_0[0]),.dout(n1081),.clk(gclk));
	jor g0781(.dina(w_n852_7[1]),.dinb(w_G17_0[0]),.dout(n1082),.clk(gclk));
	jand g0782(.dina(n1082),.dinb(w_G4090_3[1]),.dout(n1083),.clk(gclk));
	jand g0783(.dina(n1083),.dinb(n1081),.dout(n1084),.clk(gclk));
	jor g0784(.dina(w_n1043_1[0]),.dinb(w_n852_7[0]),.dout(n1085),.clk(gclk));
	jor g0785(.dina(w_n1041_1[0]),.dinb(w_G4089_7[0]),.dout(n1086),.clk(gclk));
	jand g0786(.dina(n1086),.dinb(n1085),.dout(n1087),.clk(gclk));
	jand g0787(.dina(n1087),.dinb(w_n854_3[1]),.dout(n1088),.clk(gclk));
	jor g0788(.dina(n1088),.dinb(w_dff_B_vdVDT8fO7_1),.dout(w_dff_A_K4sCI48D9_2),.clk(gclk));
	jor g0789(.dina(w_n1052_1[0]),.dinb(w_n852_6[2]),.dout(n1090),.clk(gclk));
	jor g0790(.dina(w_n1054_1[0]),.dinb(w_G4089_6[2]),.dout(n1091),.clk(gclk));
	jand g0791(.dina(n1091),.dinb(w_n854_3[0]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(n1092),.dinb(w_dff_B_rdYUYjWb3_1),.dout(n1093),.clk(gclk));
	jor g0793(.dina(w_n852_6[1]),.dinb(w_G70_0[0]),.dout(n1094),.clk(gclk));
	jor g0794(.dina(w_G4089_6[1]),.dinb(w_G67_0[0]),.dout(n1095),.clk(gclk));
	jand g0795(.dina(n1095),.dinb(w_G4090_3[0]),.dout(n1096),.clk(gclk));
	jand g0796(.dina(n1096),.dinb(n1094),.dout(n1097),.clk(gclk));
	jor g0797(.dina(w_dff_B_ePcFd7uz4_0),.dinb(n1093),.dout(w_dff_A_aqlIY8yf5_2),.clk(gclk));
	jor g0798(.dina(w_n1021_0[2]),.dinb(w_G1689_4[1]),.dout(n1099),.clk(gclk));
	jor g0799(.dina(w_n1019_0[2]),.dinb(w_n993_4[0]),.dout(n1100),.clk(gclk));
	jand g0800(.dina(n1100),.dinb(w_n999_3[1]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(n1101),.dinb(w_dff_B_b3hbbYEy1_1),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n994_4[0]),.dinb(w_G200_0[1]),.dout(n1103),.clk(gclk));
	jand g0803(.dina(w_n996_4[0]),.dinb(w_G170_0[1]),.dout(n1104),.clk(gclk));
	jor g0804(.dina(n1104),.dinb(n1103),.dout(n1105),.clk(gclk));
	jor g0805(.dina(w_dff_B_Hci9Zji85_0),.dinb(n1102),.dout(n1106),.clk(gclk));
	jand g0806(.dina(n1106),.dinb(w_G137_8[2]),.dout(w_dff_A_eXtTYCE04_2),.clk(gclk));
	jor g0807(.dina(w_n1054_0[2]),.dinb(w_G1689_4[0]),.dout(n1108),.clk(gclk));
	jor g0808(.dina(w_n1052_0[2]),.dinb(w_n993_3[2]),.dout(n1109),.clk(gclk));
	jand g0809(.dina(n1109),.dinb(w_n999_3[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(w_dff_B_YpGI6jln1_0),.dinb(n1108),.dout(n1111),.clk(gclk));
	jand g0811(.dina(w_n994_3[2]),.dinb(w_G188_0[1]),.dout(n1112),.clk(gclk));
	jand g0812(.dina(w_n996_3[2]),.dinb(w_G158_0[1]),.dout(n1113),.clk(gclk));
	jor g0813(.dina(n1113),.dinb(n1112),.dout(n1114),.clk(gclk));
	jor g0814(.dina(w_dff_B_Suvoinvj4_0),.dinb(n1111),.dout(n1115),.clk(gclk));
	jand g0815(.dina(n1115),.dinb(w_G137_8[1]),.dout(w_dff_A_vEcDfA282_2),.clk(gclk));
	jor g0816(.dina(w_n1041_0[2]),.dinb(w_G1689_3[2]),.dout(n1117),.clk(gclk));
	jor g0817(.dina(w_n1043_0[2]),.dinb(w_n993_3[1]),.dout(n1118),.clk(gclk));
	jand g0818(.dina(n1118),.dinb(w_n999_2[2]),.dout(n1119),.clk(gclk));
	jand g0819(.dina(n1119),.dinb(w_dff_B_PvQKJ1lH9_1),.dout(n1120),.clk(gclk));
	jand g0820(.dina(w_n994_3[1]),.dinb(w_G155_0[1]),.dout(n1121),.clk(gclk));
	jand g0821(.dina(w_n996_3[1]),.dinb(w_G152_0[1]),.dout(n1122),.clk(gclk));
	jor g0822(.dina(n1122),.dinb(n1121),.dout(n1123),.clk(gclk));
	jor g0823(.dina(w_dff_B_Y7YB1tXd4_0),.dinb(n1120),.dout(n1124),.clk(gclk));
	jand g0824(.dina(n1124),.dinb(w_G137_8[0]),.dout(w_dff_A_b47UtnYZ5_2),.clk(gclk));
	jor g0825(.dina(w_n1032_0[2]),.dinb(w_G1689_3[1]),.dout(n1126),.clk(gclk));
	jor g0826(.dina(w_n1030_0[2]),.dinb(w_n993_3[0]),.dout(n1127),.clk(gclk));
	jand g0827(.dina(n1127),.dinb(w_n999_2[1]),.dout(n1128),.clk(gclk));
	jand g0828(.dina(n1128),.dinb(n1126),.dout(n1129),.clk(gclk));
	jand g0829(.dina(w_n994_3[0]),.dinb(w_G149_0[1]),.dout(n1130),.clk(gclk));
	jand g0830(.dina(w_n996_3[0]),.dinb(w_G146_0[1]),.dout(n1131),.clk(gclk));
	jor g0831(.dina(n1131),.dinb(n1130),.dout(n1132),.clk(gclk));
	jor g0832(.dina(w_dff_B_Sq6Y1wZs9_0),.dinb(n1129),.dout(n1133),.clk(gclk));
	jand g0833(.dina(n1133),.dinb(w_G137_7[2]),.dout(w_dff_A_TjGCcada8_2),.clk(gclk));
	jand g0834(.dina(w_n1014_4[0]),.dinb(w_G200_0[0]),.dout(n1135),.clk(gclk));
	jand g0835(.dina(w_n1012_4[0]),.dinb(w_G170_0[0]),.dout(n1136),.clk(gclk));
	jor g0836(.dina(w_n1019_0[1]),.dinb(w_n1008_4[0]),.dout(n1137),.clk(gclk));
	jor g0837(.dina(w_n1021_0[1]),.dinb(w_G1691_4[1]),.dout(n1138),.clk(gclk));
	jand g0838(.dina(n1138),.dinb(n1137),.dout(n1139),.clk(gclk));
	jand g0839(.dina(n1139),.dinb(w_n1007_3[1]),.dout(n1140),.clk(gclk));
	jor g0840(.dina(n1140),.dinb(w_dff_B_DCt5fdP63_1),.dout(n1141),.clk(gclk));
	jor g0841(.dina(n1141),.dinb(w_dff_B_ILpdYLST9_1),.dout(n1142),.clk(gclk));
	jand g0842(.dina(n1142),.dinb(w_G137_7[1]),.dout(w_dff_A_CNem8CWd3_2),.clk(gclk));
	jor g0843(.dina(w_n1054_0[1]),.dinb(w_G1691_4[0]),.dout(n1144),.clk(gclk));
	jor g0844(.dina(w_n1052_0[1]),.dinb(w_n1008_3[2]),.dout(n1145),.clk(gclk));
	jand g0845(.dina(n1145),.dinb(w_n1007_3[0]),.dout(n1146),.clk(gclk));
	jand g0846(.dina(w_dff_B_i1xdznr45_0),.dinb(n1144),.dout(n1147),.clk(gclk));
	jand g0847(.dina(w_n1014_3[2]),.dinb(w_G188_0[0]),.dout(n1148),.clk(gclk));
	jand g0848(.dina(w_n1012_3[2]),.dinb(w_G158_0[0]),.dout(n1149),.clk(gclk));
	jor g0849(.dina(n1149),.dinb(n1148),.dout(n1150),.clk(gclk));
	jor g0850(.dina(w_dff_B_WBQU4sIr8_0),.dinb(n1147),.dout(n1151),.clk(gclk));
	jand g0851(.dina(n1151),.dinb(w_G137_7[0]),.dout(w_dff_A_rqUWwm8M5_2),.clk(gclk));
	jor g0852(.dina(w_n1041_0[1]),.dinb(w_G1691_3[2]),.dout(n1153),.clk(gclk));
	jor g0853(.dina(w_n1043_0[1]),.dinb(w_n1008_3[1]),.dout(n1154),.clk(gclk));
	jand g0854(.dina(n1154),.dinb(w_n1007_2[2]),.dout(n1155),.clk(gclk));
	jand g0855(.dina(n1155),.dinb(w_dff_B_3qN4cbYf0_1),.dout(n1156),.clk(gclk));
	jand g0856(.dina(w_n1014_3[1]),.dinb(w_G155_0[0]),.dout(n1157),.clk(gclk));
	jand g0857(.dina(w_n1012_3[1]),.dinb(w_G152_0[0]),.dout(n1158),.clk(gclk));
	jor g0858(.dina(n1158),.dinb(n1157),.dout(n1159),.clk(gclk));
	jor g0859(.dina(w_dff_B_6dxuLh870_0),.dinb(n1156),.dout(n1160),.clk(gclk));
	jand g0860(.dina(n1160),.dinb(w_G137_6[2]),.dout(w_dff_A_Wj8inUZF4_2),.clk(gclk));
	jor g0861(.dina(w_n1032_0[1]),.dinb(w_G1691_3[1]),.dout(n1162),.clk(gclk));
	jor g0862(.dina(w_n1030_0[1]),.dinb(w_n1008_3[0]),.dout(n1163),.clk(gclk));
	jand g0863(.dina(n1163),.dinb(w_n1007_2[1]),.dout(n1164),.clk(gclk));
	jand g0864(.dina(n1164),.dinb(n1162),.dout(n1165),.clk(gclk));
	jand g0865(.dina(w_n1014_3[0]),.dinb(w_G149_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n1012_3[0]),.dinb(w_G146_0[0]),.dout(n1167),.clk(gclk));
	jor g0867(.dina(n1167),.dinb(n1166),.dout(n1168),.clk(gclk));
	jor g0868(.dina(w_dff_B_1oUwOJya1_0),.dinb(n1165),.dout(n1169),.clk(gclk));
	jand g0869(.dina(n1169),.dinb(w_G137_6[1]),.dout(w_dff_A_8GjDZDev4_2),.clk(gclk));
	jnot g0870(.din(G135),.dout(n1171),.clk(gclk));
	jnot g0871(.din(G4115),.dout(n1172),.clk(gclk));
	jor g0872(.dina(n1172),.dinb(n1171),.dout(n1173),.clk(gclk));
	jnot g0873(.din(w_n428_1[0]),.dout(n1174),.clk(gclk));
	jor g0874(.dina(n1174),.dinb(w_G3724_0[2]),.dout(n1175),.clk(gclk));
	jnot g0875(.din(w_G3717_0[1]),.dout(n1176),.clk(gclk));
	jnot g0876(.din(w_G3724_0[1]),.dout(n1177),.clk(gclk));
	jxor g0877(.dina(w_n790_0[0]),.dinb(w_dff_B_XYwVKQL19_1),.dout(n1178),.clk(gclk));
	jnot g0878(.din(n1178),.dout(n1179),.clk(gclk));
	jor g0879(.dina(w_n1179_0[1]),.dinb(w_n1177_0[1]),.dout(n1180),.clk(gclk));
	jand g0880(.dina(n1180),.dinb(w_dff_B_c9rVHgUN5_1),.dout(n1181),.clk(gclk));
	jand g0881(.dina(n1181),.dinb(w_dff_B_g6dH3Znt0_1),.dout(n1182),.clk(gclk));
	jor g0882(.dina(w_n795_1[0]),.dinb(w_n1177_0[0]),.dout(n1183),.clk(gclk));
	jor g0883(.dina(w_G3724_0[0]),.dinb(w_G123_0[1]),.dout(n1184),.clk(gclk));
	jand g0884(.dina(n1184),.dinb(w_G3717_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(w_dff_B_FSaM279M7_0),.dinb(n1183),.dout(n1186),.clk(gclk));
	jor g0886(.dina(n1186),.dinb(w_dff_B_3gDUGkFP6_1),.dout(n1187),.clk(gclk));
	jand g0887(.dina(n1187),.dinb(w_dff_B_1JZQHkVQ8_1),.dout(w_dff_A_TaBL4Brs2_2),.clk(gclk));
	jxor g0888(.dina(w_n1179_0[0]),.dinb(w_n795_0[2]),.dout(w_dff_A_8tn0NyFO1_2),.clk(gclk));
	jand g0889(.dina(w_n750_5[1]),.dinb(w_G123_0[0]),.dout(n1190),.clk(gclk));
	jor g0890(.dina(w_n795_0[1]),.dinb(w_n749_9[2]),.dout(n1191),.clk(gclk));
	jand g0891(.dina(w_n428_0[2]),.dinb(w_n749_9[1]),.dout(n1192),.clk(gclk));
	jor g0892(.dina(n1192),.dinb(w_G4092_6[0]),.dout(n1193),.clk(gclk));
	jnot g0893(.din(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_dff_B_zoa86Shm5_0),.dinb(n1191),.dout(n1195),.clk(gclk));
	jor g0895(.dina(n1195),.dinb(w_dff_B_3D7jzu8O1_1),.dout(n1196),.clk(gclk));
	jnot g0896(.din(w_n1196_1[2]),.dout(w_dff_A_qGyy1NWt1_1),.clk(gclk));
	jand g0897(.dina(w_n750_5[0]),.dinb(G121),.dout(n1198),.clk(gclk));
	jand g0898(.dina(w_n433_0[1]),.dinb(w_n749_9[0]),.dout(n1199),.clk(gclk));
	jnot g0899(.din(n1199),.dout(n1200),.clk(gclk));
	jnot g0900(.din(w_G4092_5[2]),.dout(n1201),.clk(gclk));
	jor g0901(.dina(w_n969_0[0]),.dinb(w_n749_8[2]),.dout(n1202),.clk(gclk));
	jand g0902(.dina(n1202),.dinb(w_n1201_0[2]),.dout(n1203),.clk(gclk));
	jand g0903(.dina(n1203),.dinb(w_dff_B_HLuv4sqU8_1),.dout(n1204),.clk(gclk));
	jor g0904(.dina(n1204),.dinb(w_dff_B_bArBZE0s8_1),.dout(n1205),.clk(gclk));
	jnot g0905(.din(w_n1205_1[2]),.dout(w_dff_A_EVE9Od673_1),.clk(gclk));
	jand g0906(.dina(w_n750_4[2]),.dinb(G116),.dout(n1207),.clk(gclk));
	jor g0907(.dina(w_n986_0[0]),.dinb(w_n749_8[1]),.dout(n1208),.clk(gclk));
	jand g0908(.dina(w_n423_0[1]),.dinb(w_n749_8[0]),.dout(n1209),.clk(gclk));
	jor g0909(.dina(n1209),.dinb(w_G4092_5[1]),.dout(n1210),.clk(gclk));
	jnot g0910(.din(n1210),.dout(n1211),.clk(gclk));
	jand g0911(.dina(w_dff_B_AMlJ6zkX7_0),.dinb(n1208),.dout(n1212),.clk(gclk));
	jor g0912(.dina(n1212),.dinb(w_dff_B_M3qIf25O9_1),.dout(n1213),.clk(gclk));
	jnot g0913(.din(w_n1213_1[2]),.dout(w_dff_A_vpYvFGV21_1),.clk(gclk));
	jand g0914(.dina(w_n750_4[1]),.dinb(G112),.dout(n1215),.clk(gclk));
	jnot g0915(.din(n1215),.dout(n1216),.clk(gclk));
	jand g0916(.dina(w_n989_0[0]),.dinb(w_G4091_2[2]),.dout(n1217),.clk(gclk));
	jand g0917(.dina(w_n412_0[1]),.dinb(w_n749_7[2]),.dout(n1218),.clk(gclk));
	jor g0918(.dina(n1218),.dinb(w_G4092_5[0]),.dout(n1219),.clk(gclk));
	jor g0919(.dina(w_dff_B_Z4JsXH4x2_0),.dinb(n1217),.dout(n1220),.clk(gclk));
	jand g0920(.dina(n1220),.dinb(w_dff_B_oEGnkt1Y0_1),.dout(G830_fa_),.clk(gclk));
	jand g0921(.dina(w_n680_0[0]),.dinb(w_G245_0[0]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(n1222),.dinb(w_n935_0[0]),.dout(n1223),.clk(gclk));
	jnot g0923(.din(w_G998_0),.dout(n1224),.clk(gclk));
	jand g0924(.dina(w_n318_0[0]),.dinb(w_G601_0),.dout(n1225),.clk(gclk));
	jand g0925(.dina(n1225),.dinb(w_G559_0[0]),.dout(n1226),.clk(gclk));
	jand g0926(.dina(w_dff_B_BzKGYPfc6_0),.dinb(w_n670_0[0]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_dff_B_uXwQUzK48_0),.dinb(n1224),.dout(n1228),.clk(gclk));
	jand g0928(.dina(n1228),.dinb(w_dff_B_DKZt5hg95_1),.dout(w_dff_A_HFgIIjdN5_2),.clk(gclk));
	jand g0929(.dina(w_n750_4[0]),.dinb(G115),.dout(n1230),.clk(gclk));
	jand g0930(.dina(w_n551_0[1]),.dinb(w_n749_7[1]),.dout(n1231),.clk(gclk));
	jnot g0931(.din(n1231),.dout(n1232),.clk(gclk));
	jor g0932(.dina(w_n944_0[0]),.dinb(w_n749_7[0]),.dout(n1233),.clk(gclk));
	jand g0933(.dina(n1233),.dinb(w_n1201_0[1]),.dout(n1234),.clk(gclk));
	jand g0934(.dina(n1234),.dinb(n1232),.dout(n1235),.clk(gclk));
	jor g0935(.dina(n1235),.dinb(n1230),.dout(n1236),.clk(gclk));
	jnot g0936(.din(w_n1236_1[2]),.dout(w_dff_A_TarUmmSU2_1),.clk(gclk));
	jand g0937(.dina(w_n750_3[2]),.dinb(G114),.dout(n1238),.clk(gclk));
	jnot g0938(.din(n1238),.dout(n1239),.clk(gclk));
	jand g0939(.dina(w_n949_0[0]),.dinb(w_G4091_2[1]),.dout(n1240),.clk(gclk));
	jand g0940(.dina(w_n459_0[0]),.dinb(w_n749_6[2]),.dout(n1241),.clk(gclk));
	jor g0941(.dina(n1241),.dinb(w_G4092_4[2]),.dout(n1242),.clk(gclk));
	jor g0942(.dina(n1242),.dinb(n1240),.dout(n1243),.clk(gclk));
	jand g0943(.dina(n1243),.dinb(n1239),.dout(G865_fa_),.clk(gclk));
	jand g0944(.dina(w_n750_3[1]),.dinb(G53),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n517_0[0]),.dinb(w_n749_6[1]),.dout(n1246),.clk(gclk));
	jnot g0946(.din(n1246),.dout(n1247),.clk(gclk));
	jor g0947(.dina(w_n957_0[0]),.dinb(w_n749_6[0]),.dout(n1248),.clk(gclk));
	jand g0948(.dina(n1248),.dinb(w_n1201_0[0]),.dout(n1249),.clk(gclk));
	jand g0949(.dina(n1249),.dinb(n1247),.dout(n1250),.clk(gclk));
	jor g0950(.dina(n1250),.dinb(n1245),.dout(n1251),.clk(gclk));
	jnot g0951(.din(w_n1251_1[2]),.dout(w_dff_A_mmpAPBTa5_1),.clk(gclk));
	jand g0952(.dina(w_n750_3[0]),.dinb(G113),.dout(n1253),.clk(gclk));
	jnot g0953(.din(n1253),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n964_0[0]),.dinb(w_G4091_2[0]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n504_0[0]),.dinb(w_n749_5[2]),.dout(n1256),.clk(gclk));
	jor g0956(.dina(n1256),.dinb(w_G4092_4[1]),.dout(n1257),.clk(gclk));
	jor g0957(.dina(n1257),.dinb(n1255),.dout(n1258),.clk(gclk));
	jand g0958(.dina(n1258),.dinb(n1254),.dout(G869_fa_),.clk(gclk));
	jor g0959(.dina(w_G4089_6[0]),.dinb(w_G109_0[1]),.dout(n1260),.clk(gclk));
	jor g0960(.dina(w_n852_6[0]),.dinb(w_G106_0[1]),.dout(n1261),.clk(gclk));
	jand g0961(.dina(n1261),.dinb(w_G4090_2[2]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(n1262),.dinb(n1260),.dout(n1263),.clk(gclk));
	jor g0963(.dina(w_n1236_1[1]),.dinb(w_n852_5[2]),.dout(n1264),.clk(gclk));
	jor g0964(.dina(w_n1196_1[1]),.dinb(w_G4089_5[2]),.dout(n1265),.clk(gclk));
	jand g0965(.dina(n1265),.dinb(w_n854_2[2]),.dout(n1266),.clk(gclk));
	jand g0966(.dina(n1266),.dinb(n1264),.dout(n1267),.clk(gclk));
	jor g0967(.dina(n1267),.dinb(w_dff_B_9knjpEj62_1),.dout(w_dff_A_dkFs5zUM9_2),.clk(gclk));
	jor g0968(.dina(w_n1196_1[0]),.dinb(w_G4088_6[0]),.dout(n1269),.clk(gclk));
	jor g0969(.dina(w_n1236_1[0]),.dinb(w_n797_6[0]),.dout(n1270),.clk(gclk));
	jand g0970(.dina(n1270),.dinb(w_n800_2[2]),.dout(n1271),.clk(gclk));
	jand g0971(.dina(n1271),.dinb(w_dff_B_Ra935SOO5_1),.dout(n1272),.clk(gclk));
	jor g0972(.dina(w_n797_5[2]),.dinb(w_G106_0[0]),.dout(n1273),.clk(gclk));
	jor g0973(.dina(w_G4088_5[2]),.dinb(w_G109_0[0]),.dout(n1274),.clk(gclk));
	jand g0974(.dina(n1274),.dinb(w_G4087_2[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(n1275),.dinb(n1273),.dout(n1276),.clk(gclk));
	jor g0976(.dina(w_dff_B_uPb3CPjh2_0),.dinb(n1272),.dout(w_dff_A_xn8VXQlt9_2),.clk(gclk));
	jor g0977(.dina(w_n1205_1[1]),.dinb(w_G4088_5[1]),.dout(n1278),.clk(gclk));
	jnot g0978(.din(w_G865_0),.dout(n1279),.clk(gclk));
	jor g0979(.dina(w_n1279_1[1]),.dinb(w_n797_5[1]),.dout(n1280),.clk(gclk));
	jand g0980(.dina(n1280),.dinb(w_n800_2[1]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(n1281),.dinb(w_dff_B_KCaiDqnp0_1),.dout(n1282),.clk(gclk));
	jor g0982(.dina(w_n797_5[0]),.dinb(w_G49_0[1]),.dout(n1283),.clk(gclk));
	jor g0983(.dina(w_G4088_5[0]),.dinb(w_G46_0[1]),.dout(n1284),.clk(gclk));
	jand g0984(.dina(n1284),.dinb(w_G4087_2[1]),.dout(n1285),.clk(gclk));
	jand g0985(.dina(n1285),.dinb(n1283),.dout(n1286),.clk(gclk));
	jor g0986(.dina(w_dff_B_DAHkaWdf2_0),.dinb(n1282),.dout(w_dff_A_ThgarqCR8_2),.clk(gclk));
	jor g0987(.dina(w_n1213_1[1]),.dinb(w_G4088_4[2]),.dout(n1288),.clk(gclk));
	jor g0988(.dina(w_n1251_1[1]),.dinb(w_n797_4[2]),.dout(n1289),.clk(gclk));
	jand g0989(.dina(n1289),.dinb(w_n800_2[0]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(n1290),.dinb(w_dff_B_hm6V1Wnr4_1),.dout(n1291),.clk(gclk));
	jor g0991(.dina(w_n797_4[1]),.dinb(w_G103_0[1]),.dout(n1292),.clk(gclk));
	jor g0992(.dina(w_G4088_4[1]),.dinb(w_G100_0[1]),.dout(n1293),.clk(gclk));
	jand g0993(.dina(n1293),.dinb(w_G4087_2[0]),.dout(n1294),.clk(gclk));
	jand g0994(.dina(n1294),.dinb(n1292),.dout(n1295),.clk(gclk));
	jor g0995(.dina(w_dff_B_hnqC9Wmu9_0),.dinb(n1291),.dout(w_dff_A_iLcxeVf72_2),.clk(gclk));
	jnot g0996(.din(w_G830_0),.dout(n1297),.clk(gclk));
	jor g0997(.dina(w_n1297_1[1]),.dinb(w_G4088_4[0]),.dout(n1298),.clk(gclk));
	jnot g0998(.din(w_G869_0),.dout(n1299),.clk(gclk));
	jor g0999(.dina(w_n1299_1[1]),.dinb(w_n797_4[0]),.dout(n1300),.clk(gclk));
	jand g1000(.dina(n1300),.dinb(w_n800_1[2]),.dout(n1301),.clk(gclk));
	jand g1001(.dina(n1301),.dinb(w_dff_B_6YQPmrv72_1),.dout(n1302),.clk(gclk));
	jor g1002(.dina(w_n797_3[2]),.dinb(w_G40_0[1]),.dout(n1303),.clk(gclk));
	jor g1003(.dina(w_G4088_3[2]),.dinb(w_G91_0[1]),.dout(n1304),.clk(gclk));
	jand g1004(.dina(n1304),.dinb(w_G4087_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(n1305),.dinb(n1303),.dout(n1306),.clk(gclk));
	jor g1006(.dina(w_dff_B_6tvoiiKt9_0),.dinb(n1302),.dout(w_dff_A_VciU7eAY5_2),.clk(gclk));
	jor g1007(.dina(w_n1205_1[0]),.dinb(w_G4089_5[1]),.dout(n1308),.clk(gclk));
	jor g1008(.dina(w_n1279_1[0]),.dinb(w_n852_5[1]),.dout(n1309),.clk(gclk));
	jand g1009(.dina(n1309),.dinb(w_n854_2[1]),.dout(n1310),.clk(gclk));
	jand g1010(.dina(n1310),.dinb(w_dff_B_bodC3ZIz1_1),.dout(n1311),.clk(gclk));
	jor g1011(.dina(w_n852_5[0]),.dinb(w_G49_0[0]),.dout(n1312),.clk(gclk));
	jor g1012(.dina(w_G4089_5[0]),.dinb(w_G46_0[0]),.dout(n1313),.clk(gclk));
	jand g1013(.dina(n1313),.dinb(w_G4090_2[1]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(n1314),.dinb(n1312),.dout(n1315),.clk(gclk));
	jor g1015(.dina(w_dff_B_9PryGx0C4_0),.dinb(n1311),.dout(w_dff_A_iVCTOc7f1_2),.clk(gclk));
	jor g1016(.dina(w_n1213_1[0]),.dinb(w_G4089_4[2]),.dout(n1317),.clk(gclk));
	jor g1017(.dina(w_n1251_1[0]),.dinb(w_n852_4[2]),.dout(n1318),.clk(gclk));
	jand g1018(.dina(n1318),.dinb(w_n854_2[0]),.dout(n1319),.clk(gclk));
	jand g1019(.dina(n1319),.dinb(w_dff_B_5OLRqP5N6_1),.dout(n1320),.clk(gclk));
	jor g1020(.dina(w_n852_4[1]),.dinb(w_G103_0[0]),.dout(n1321),.clk(gclk));
	jor g1021(.dina(w_G4089_4[1]),.dinb(w_G100_0[0]),.dout(n1322),.clk(gclk));
	jand g1022(.dina(n1322),.dinb(w_G4090_2[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(n1323),.dinb(n1321),.dout(n1324),.clk(gclk));
	jor g1024(.dina(w_dff_B_fSABNbnM3_0),.dinb(n1320),.dout(w_dff_A_QaYaxUiX3_2),.clk(gclk));
	jor g1025(.dina(w_n1297_1[0]),.dinb(w_G4089_4[0]),.dout(n1326),.clk(gclk));
	jor g1026(.dina(w_n1299_1[0]),.dinb(w_n852_4[0]),.dout(n1327),.clk(gclk));
	jand g1027(.dina(n1327),.dinb(w_n854_1[2]),.dout(n1328),.clk(gclk));
	jand g1028(.dina(n1328),.dinb(w_dff_B_2v01HJmp0_1),.dout(n1329),.clk(gclk));
	jor g1029(.dina(w_n852_3[2]),.dinb(w_G40_0[0]),.dout(n1330),.clk(gclk));
	jor g1030(.dina(w_G4089_3[2]),.dinb(w_G91_0[0]),.dout(n1331),.clk(gclk));
	jand g1031(.dina(n1331),.dinb(w_G4090_1[2]),.dout(n1332),.clk(gclk));
	jand g1032(.dina(n1332),.dinb(n1330),.dout(n1333),.clk(gclk));
	jor g1033(.dina(w_dff_B_3gu5XD3k4_0),.dinb(n1329),.dout(w_dff_A_ukNOl0VY4_2),.clk(gclk));
	jor g1034(.dina(w_n1297_0[2]),.dinb(w_G1689_3[0]),.dout(n1335),.clk(gclk));
	jor g1035(.dina(w_n1299_0[2]),.dinb(w_n993_2[2]),.dout(n1336),.clk(gclk));
	jand g1036(.dina(n1336),.dinb(w_n999_2[0]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(n1337),.dinb(w_dff_B_E6w3HOae8_1),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n994_2[2]),.dinb(w_G203_0[1]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n996_2[2]),.dinb(w_G173_0[1]),.dout(n1340),.clk(gclk));
	jor g1040(.dina(n1340),.dinb(n1339),.dout(n1341),.clk(gclk));
	jor g1041(.dina(w_dff_B_G0EZjB2W9_0),.dinb(n1338),.dout(n1342),.clk(gclk));
	jand g1042(.dina(n1342),.dinb(w_G137_6[0]),.dout(w_dff_A_OlaI97sX7_2),.clk(gclk));
	jor g1043(.dina(w_n1251_0[2]),.dinb(w_n993_2[1]),.dout(n1344),.clk(gclk));
	jor g1044(.dina(w_n1213_0[2]),.dinb(w_G1689_2[2]),.dout(n1345),.clk(gclk));
	jand g1045(.dina(n1345),.dinb(w_n999_1[2]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(n1346),.dinb(w_dff_B_RrZERRcd2_1),.dout(n1347),.clk(gclk));
	jand g1047(.dina(w_n994_2[1]),.dinb(w_G197_0[1]),.dout(n1348),.clk(gclk));
	jand g1048(.dina(w_n996_2[1]),.dinb(w_G167_0[1]),.dout(n1349),.clk(gclk));
	jor g1049(.dina(n1349),.dinb(n1348),.dout(n1350),.clk(gclk));
	jor g1050(.dina(w_dff_B_7juUKr1R2_0),.dinb(n1347),.dout(n1351),.clk(gclk));
	jand g1051(.dina(n1351),.dinb(w_G137_5[2]),.dout(w_dff_A_TBsLnPUK2_2),.clk(gclk));
	jand g1052(.dina(w_n994_2[0]),.dinb(w_G194_0[1]),.dout(n1353),.clk(gclk));
	jand g1053(.dina(w_n996_2[0]),.dinb(w_G164_0[1]),.dout(n1354),.clk(gclk));
	jor g1054(.dina(n1354),.dinb(n1353),.dout(n1355),.clk(gclk));
	jor g1055(.dina(w_n1205_0[2]),.dinb(w_G1689_2[1]),.dout(n1356),.clk(gclk));
	jor g1056(.dina(w_n1279_0[2]),.dinb(w_n993_2[0]),.dout(n1357),.clk(gclk));
	jand g1057(.dina(n1357),.dinb(w_dff_B_sHmOrsaS5_1),.dout(n1358),.clk(gclk));
	jand g1058(.dina(n1358),.dinb(w_n999_1[1]),.dout(n1359),.clk(gclk));
	jor g1059(.dina(n1359),.dinb(w_dff_B_4HwUVt8K3_1),.dout(n1360),.clk(gclk));
	jand g1060(.dina(n1360),.dinb(w_G137_5[1]),.dout(w_dff_A_dzvMNPTC6_2),.clk(gclk));
	jand g1061(.dina(w_n994_1[2]),.dinb(w_G191_0[1]),.dout(n1362),.clk(gclk));
	jand g1062(.dina(w_n996_1[2]),.dinb(w_G161_0[1]),.dout(n1363),.clk(gclk));
	jor g1063(.dina(n1363),.dinb(n1362),.dout(n1364),.clk(gclk));
	jor g1064(.dina(w_n1196_0[2]),.dinb(w_G1689_2[0]),.dout(n1365),.clk(gclk));
	jor g1065(.dina(w_n1236_0[2]),.dinb(w_n993_1[2]),.dout(n1366),.clk(gclk));
	jand g1066(.dina(n1366),.dinb(w_dff_B_nrRPA6hl1_1),.dout(n1367),.clk(gclk));
	jand g1067(.dina(n1367),.dinb(w_n999_1[0]),.dout(n1368),.clk(gclk));
	jor g1068(.dina(n1368),.dinb(w_dff_B_2xEXa9Lg2_1),.dout(n1369),.clk(gclk));
	jand g1069(.dina(n1369),.dinb(w_G137_5[0]),.dout(w_dff_A_NOl4MacD3_2),.clk(gclk));
	jor g1070(.dina(w_n1297_0[1]),.dinb(w_G1691_3[0]),.dout(n1371),.clk(gclk));
	jor g1071(.dina(w_n1299_0[1]),.dinb(w_n1008_2[2]),.dout(n1372),.clk(gclk));
	jand g1072(.dina(n1372),.dinb(w_n1007_2[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(n1373),.dinb(w_dff_B_LBJurNfu5_1),.dout(n1374),.clk(gclk));
	jand g1074(.dina(w_n1014_2[2]),.dinb(w_G203_0[0]),.dout(n1375),.clk(gclk));
	jand g1075(.dina(w_n1012_2[2]),.dinb(w_G173_0[0]),.dout(n1376),.clk(gclk));
	jor g1076(.dina(n1376),.dinb(n1375),.dout(n1377),.clk(gclk));
	jor g1077(.dina(w_dff_B_XSJFcWbz3_0),.dinb(n1374),.dout(n1378),.clk(gclk));
	jand g1078(.dina(n1378),.dinb(w_G137_4[2]),.dout(w_dff_A_Udi9HLES1_2),.clk(gclk));
	jand g1079(.dina(w_n1014_2[1]),.dinb(w_G197_0[0]),.dout(n1380),.clk(gclk));
	jand g1080(.dina(w_n1012_2[1]),.dinb(w_G167_0[0]),.dout(n1381),.clk(gclk));
	jor g1081(.dina(n1381),.dinb(n1380),.dout(n1382),.clk(gclk));
	jor g1082(.dina(w_n1213_0[1]),.dinb(w_G1691_2[2]),.dout(n1383),.clk(gclk));
	jor g1083(.dina(w_n1251_0[1]),.dinb(w_n1008_2[1]),.dout(n1384),.clk(gclk));
	jand g1084(.dina(n1384),.dinb(n1383),.dout(n1385),.clk(gclk));
	jand g1085(.dina(n1385),.dinb(w_n1007_1[2]),.dout(n1386),.clk(gclk));
	jor g1086(.dina(n1386),.dinb(w_dff_B_VkGZTCwZ0_1),.dout(n1387),.clk(gclk));
	jand g1087(.dina(n1387),.dinb(w_G137_4[1]),.dout(w_dff_A_CXlZvC9V9_2),.clk(gclk));
	jor g1088(.dina(w_n1205_0[1]),.dinb(w_G1691_2[1]),.dout(n1389),.clk(gclk));
	jor g1089(.dina(w_n1279_0[1]),.dinb(w_n1008_2[0]),.dout(n1390),.clk(gclk));
	jand g1090(.dina(n1390),.dinb(w_n1007_1[1]),.dout(n1391),.clk(gclk));
	jand g1091(.dina(n1391),.dinb(w_dff_B_MyNQdqJ97_1),.dout(n1392),.clk(gclk));
	jand g1092(.dina(w_n1014_2[0]),.dinb(w_G194_0[0]),.dout(n1393),.clk(gclk));
	jand g1093(.dina(w_n1012_2[0]),.dinb(w_G164_0[0]),.dout(n1394),.clk(gclk));
	jor g1094(.dina(n1394),.dinb(n1393),.dout(n1395),.clk(gclk));
	jor g1095(.dina(w_dff_B_j5DK7ZyH8_0),.dinb(n1392),.dout(n1396),.clk(gclk));
	jand g1096(.dina(n1396),.dinb(w_G137_4[0]),.dout(w_dff_A_jSG9y9fp6_2),.clk(gclk));
	jor g1097(.dina(w_n1236_0[1]),.dinb(w_n1008_1[2]),.dout(n1398),.clk(gclk));
	jor g1098(.dina(w_n1196_0[1]),.dinb(w_G1691_2[0]),.dout(n1399),.clk(gclk));
	jand g1099(.dina(n1399),.dinb(w_n1007_1[0]),.dout(n1400),.clk(gclk));
	jand g1100(.dina(n1400),.dinb(n1398),.dout(n1401),.clk(gclk));
	jand g1101(.dina(w_n1014_1[2]),.dinb(w_G191_0[0]),.dout(n1402),.clk(gclk));
	jand g1102(.dina(w_n1012_1[2]),.dinb(w_G161_0[0]),.dout(n1403),.clk(gclk));
	jor g1103(.dina(n1403),.dinb(n1402),.dout(n1404),.clk(gclk));
	jor g1104(.dina(w_dff_B_FNMQBBlP1_0),.dinb(n1401),.dout(n1405),.clk(gclk));
	jand g1105(.dina(n1405),.dinb(w_G137_3[2]),.dout(w_dff_A_xHbVfs0P9_2),.clk(gclk));
	jand g1106(.dina(w_n746_0[0]),.dinb(w_n648_0[2]),.dout(n1407),.clk(gclk));
	jxor g1107(.dina(w_n977_0[0]),.dinb(w_n654_1[0]),.dout(n1408),.clk(gclk));
	jxor g1108(.dina(n1408),.dinb(w_n644_0[0]),.dout(n1409),.clk(gclk));
	jxor g1109(.dina(w_dff_B_HiDGTUnB7_0),.dinb(n1407),.dout(n1410),.clk(gclk));
	jor g1110(.dina(w_n1410_0[2]),.dinb(w_n737_0[2]),.dout(n1411),.clk(gclk));
	jnot g1111(.din(w_G2174_0[2]),.dout(n1412),.clk(gclk));
	jnot g1112(.din(w_n719_0[0]),.dout(n1413),.clk(gclk));
	jnot g1113(.din(w_n720_0[0]),.dout(n1414),.clk(gclk));
	jor g1114(.dina(w_n821_0[0]),.dinb(w_dff_B_2FUUdo6f3_1),.dout(n1415),.clk(gclk));
	jand g1115(.dina(n1415),.dinb(w_dff_B_kwom3u9N4_1),.dout(n1416),.clk(gclk));
	jxor g1116(.dina(w_n742_0[0]),.dinb(w_n654_0[2]),.dout(n1417),.clk(gclk));
	jxor g1117(.dina(n1417),.dinb(w_n792_0[0]),.dout(n1418),.clk(gclk));
	jnot g1118(.din(w_n660_0[1]),.dout(n1419),.clk(gclk));
	jand g1119(.dina(w_n745_0[0]),.dinb(w_n648_0[1]),.dout(n1420),.clk(gclk));
	jand g1120(.dina(n1420),.dinb(n1419),.dout(n1421),.clk(gclk));
	jxor g1121(.dina(n1421),.dinb(w_dff_B_nfYiIvAu1_1),.dout(n1422),.clk(gclk));
	jor g1122(.dina(w_n1422_0[1]),.dinb(w_n1416_0[1]),.dout(n1423),.clk(gclk));
	jand g1123(.dina(n1423),.dinb(w_n1412_0[2]),.dout(n1424),.clk(gclk));
	jand g1124(.dina(n1424),.dinb(w_dff_B_y7USFW1T9_1),.dout(n1425),.clk(gclk));
	jnot g1125(.din(w_n1425_0[1]),.dout(n1426),.clk(gclk));
	jnot g1126(.din(w_n641_1[0]),.dout(n1427),.clk(gclk));
	jand g1127(.dina(w_n1416_0[0]),.dinb(w_dff_B_GELGpxoG6_1),.dout(n1428),.clk(gclk));
	jor g1128(.dina(w_n1428_0[1]),.dinb(w_n1422_0[0]),.dout(n1429),.clk(gclk));
	jnot g1129(.din(w_n1429_0[1]),.dout(n1430),.clk(gclk));
	jnot g1130(.din(w_n1410_0[1]),.dout(n1431),.clk(gclk));
	jand g1131(.dina(w_n1428_0[0]),.dinb(n1431),.dout(n1432),.clk(gclk));
	jor g1132(.dina(n1432),.dinb(w_n1412_0[1]),.dout(n1433),.clk(gclk));
	jor g1133(.dina(n1433),.dinb(n1430),.dout(n1434),.clk(gclk));
	jand g1134(.dina(n1434),.dinb(n1426),.dout(n1435),.clk(gclk));
	jor g1135(.dina(w_n728_0[0]),.dinb(w_n637_0[0]),.dout(n1436),.clk(gclk));
	jxor g1136(.dina(w_dff_B_lb2sWyLx1_0),.dinb(w_n733_0[1]),.dout(n1437),.clk(gclk));
	jxor g1137(.dina(w_dff_B_W3Dv9XHm7_0),.dinb(w_n735_0[1]),.dout(n1438),.clk(gclk));
	jor g1138(.dina(n1438),.dinb(w_G2174_0[1]),.dout(n1439),.clk(gclk));
	jor g1139(.dina(w_n735_0[0]),.dinb(w_n640_0[0]),.dout(n1440),.clk(gclk));
	jor g1140(.dina(w_n819_0[0]),.dinb(w_n628_0[0]),.dout(n1441),.clk(gclk));
	jor g1141(.dina(w_n733_0[0]),.dinb(w_n814_0[0]),.dout(n1442),.clk(gclk));
	jor g1142(.dina(n1442),.dinb(w_n639_0[0]),.dout(n1443),.clk(gclk));
	jand g1143(.dina(n1443),.dinb(w_dff_B_ojDaT3h42_1),.dout(n1444),.clk(gclk));
	jxor g1144(.dina(n1444),.dinb(n1440),.dout(n1445),.clk(gclk));
	jor g1145(.dina(n1445),.dinb(w_n1412_0[0]),.dout(n1446),.clk(gclk));
	jand g1146(.dina(n1446),.dinb(w_dff_B_ZqKnkvmN1_1),.dout(n1447),.clk(gclk));
	jxor g1147(.dina(w_n620_0[1]),.dinb(w_n618_0[0]),.dout(n1448),.clk(gclk));
	jxor g1148(.dina(w_n767_0[0]),.dinb(w_n624_0[0]),.dout(n1449),.clk(gclk));
	jxor g1149(.dina(n1449),.dinb(w_dff_B_p1RAyhWe0_1),.dout(n1450),.clk(gclk));
	jxor g1150(.dina(w_dff_B_8TqIhvGq3_0),.dinb(n1447),.dout(n1451),.clk(gclk));
	jnot g1151(.din(w_n1451_0[1]),.dout(n1452),.clk(gclk));
	jand g1152(.dina(w_dff_B_NO5SrzkV7_0),.dinb(n1435),.dout(n1453),.clk(gclk));
	jor g1153(.dina(w_n737_0[1]),.dinb(w_n641_0[2]),.dout(n1454),.clk(gclk));
	jor g1154(.dina(n1454),.dinb(w_n1410_0[0]),.dout(n1455),.clk(gclk));
	jand g1155(.dina(n1455),.dinb(w_G2174_0[0]),.dout(n1456),.clk(gclk));
	jand g1156(.dina(n1456),.dinb(w_n1429_0[0]),.dout(n1457),.clk(gclk));
	jor g1157(.dina(n1457),.dinb(w_n1425_0[0]),.dout(n1458),.clk(gclk));
	jand g1158(.dina(w_n1451_0[0]),.dinb(n1458),.dout(n1459),.clk(gclk));
	jor g1159(.dina(n1459),.dinb(w_n749_5[1]),.dout(n1460),.clk(gclk));
	jor g1160(.dina(n1460),.dinb(w_dff_B_0i2kTdtc2_1),.dout(n1461),.clk(gclk));
	jand g1161(.dina(w_G351_1[0]),.dinb(w_G248_4[1]),.dout(n1462),.clk(gclk));
	jand g1162(.dina(w_n374_0[2]),.dinb(w_G251_4[0]),.dout(n1463),.clk(gclk));
	jor g1163(.dina(n1463),.dinb(w_n377_0[1]),.dout(n1464),.clk(gclk));
	jor g1164(.dina(n1464),.dinb(n1462),.dout(n1465),.clk(gclk));
	jand g1165(.dina(w_n374_0[1]),.dinb(w_n406_4[0]),.dout(n1466),.clk(gclk));
	jand g1166(.dina(w_G351_0[2]),.dinb(w_n408_4[1]),.dout(n1467),.clk(gclk));
	jor g1167(.dina(n1467),.dinb(n1466),.dout(n1468),.clk(gclk));
	jor g1168(.dina(n1468),.dinb(w_G534_0[2]),.dout(n1469),.clk(gclk));
	jand g1169(.dina(n1469),.dinb(n1465),.dout(n1470),.clk(gclk));
	jand g1170(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1471),.clk(gclk));
	jand g1171(.dina(w_n387_0[2]),.dinb(w_G251_3[2]),.dout(n1472),.clk(gclk));
	jor g1172(.dina(n1472),.dinb(w_n389_0[1]),.dout(n1473),.clk(gclk));
	jor g1173(.dina(n1473),.dinb(n1471),.dout(n1474),.clk(gclk));
	jand g1174(.dina(w_n387_0[1]),.dinb(w_n406_3[2]),.dout(n1475),.clk(gclk));
	jand g1175(.dina(w_G341_0[2]),.dinb(w_n408_4[0]),.dout(n1476),.clk(gclk));
	jor g1176(.dina(n1476),.dinb(n1475),.dout(n1477),.clk(gclk));
	jor g1177(.dina(n1477),.dinb(w_G523_0[1]),.dout(n1478),.clk(gclk));
	jand g1178(.dina(n1478),.dinb(n1474),.dout(n1479),.clk(gclk));
	jxor g1179(.dina(n1479),.dinb(n1470),.dout(n1480),.clk(gclk));
	jor g1180(.dina(w_n435_1[0]),.dinb(w_n369_1[0]),.dout(n1481),.clk(gclk));
	jor g1181(.dina(w_G324_0[2]),.dinb(w_n366_1[0]),.dout(n1482),.clk(gclk));
	jand g1182(.dina(n1482),.dinb(w_G503_0[2]),.dout(n1483),.clk(gclk));
	jand g1183(.dina(n1483),.dinb(n1481),.dout(n1484),.clk(gclk));
	jor g1184(.dina(w_G324_0[1]),.dinb(w_G254_1[0]),.dout(n1485),.clk(gclk));
	jor g1185(.dina(w_n435_0[2]),.dinb(w_G242_1[0]),.dout(n1486),.clk(gclk));
	jand g1186(.dina(n1486),.dinb(n1485),.dout(n1487),.clk(gclk));
	jand g1187(.dina(n1487),.dinb(w_n437_0[0]),.dout(n1488),.clk(gclk));
	jor g1188(.dina(n1488),.dinb(n1484),.dout(n1489),.clk(gclk));
	jor g1189(.dina(w_G514_0[2]),.dinb(w_n408_3[2]),.dout(n1490),.clk(gclk));
	jor g1190(.dina(w_n361_0[0]),.dinb(w_G248_3[2]),.dout(n1491),.clk(gclk));
	jand g1191(.dina(n1491),.dinb(n1490),.dout(n1492),.clk(gclk));
	jxor g1192(.dina(n1492),.dinb(w_n371_0[0]),.dout(n1493),.clk(gclk));
	jxor g1193(.dina(n1493),.dinb(n1489),.dout(n1494),.clk(gclk));
	jxor g1194(.dina(n1494),.dinb(n1480),.dout(n1495),.clk(gclk));
	jxor g1195(.dina(w_n433_0[0]),.dinb(w_n428_0[1]),.dout(n1496),.clk(gclk));
	jxor g1196(.dina(w_n423_0[0]),.dinb(w_n412_0[0]),.dout(n1497),.clk(gclk));
	jxor g1197(.dina(n1497),.dinb(n1496),.dout(n1498),.clk(gclk));
	jxor g1198(.dina(n1498),.dinb(n1495),.dout(n1499),.clk(gclk));
	jand g1199(.dina(n1499),.dinb(w_n749_5[0]),.dout(n1500),.clk(gclk));
	jnot g1200(.din(n1500),.dout(n1501),.clk(gclk));
	jand g1201(.dina(w_dff_B_z22eYMUi6_0),.dinb(n1461),.dout(n1502),.clk(gclk));
	jor g1202(.dina(n1502),.dinb(w_G4092_4[0]),.dout(n1503),.clk(gclk));
	jnot g1203(.din(w_n750_2[2]),.dout(n1504),.clk(gclk));
	jor g1204(.dina(w_n1504_0[1]),.dinb(G120),.dout(n1505),.clk(gclk));
	jand g1205(.dina(w_dff_B_sLrBGO7P3_0),.dinb(w_n1503_0[1]),.dout(w_dff_A_YSK6IrZh6_2),.clk(gclk));
	jand g1206(.dina(w_G273_1[0]),.dinb(w_G248_3[1]),.dout(n1507),.clk(gclk));
	jand g1207(.dina(w_n471_0[2]),.dinb(w_G251_3[1]),.dout(n1508),.clk(gclk));
	jor g1208(.dina(n1508),.dinb(w_n473_1[0]),.dout(n1509),.clk(gclk));
	jor g1209(.dina(n1509),.dinb(n1507),.dout(n1510),.clk(gclk));
	jand g1210(.dina(w_n471_0[1]),.dinb(w_n406_3[1]),.dout(n1511),.clk(gclk));
	jand g1211(.dina(w_G273_0[2]),.dinb(w_n408_3[1]),.dout(n1512),.clk(gclk));
	jor g1212(.dina(n1512),.dinb(n1511),.dout(n1513),.clk(gclk));
	jor g1213(.dina(n1513),.dinb(w_G411_0[2]),.dout(n1514),.clk(gclk));
	jand g1214(.dina(n1514),.dinb(n1510),.dout(n1515),.clk(gclk));
	jand g1215(.dina(w_G281_1[0]),.dinb(w_G248_3[0]),.dout(n1516),.clk(gclk));
	jand g1216(.dina(w_n530_0[2]),.dinb(w_G251_3[0]),.dout(n1517),.clk(gclk));
	jor g1217(.dina(n1517),.dinb(w_n532_1[0]),.dout(n1518),.clk(gclk));
	jor g1218(.dina(n1518),.dinb(n1516),.dout(n1519),.clk(gclk));
	jand g1219(.dina(w_n530_0[1]),.dinb(w_n406_3[0]),.dout(n1520),.clk(gclk));
	jand g1220(.dina(w_G281_0[2]),.dinb(w_n408_3[0]),.dout(n1521),.clk(gclk));
	jor g1221(.dina(n1521),.dinb(n1520),.dout(n1522),.clk(gclk));
	jor g1222(.dina(n1522),.dinb(w_G374_0[1]),.dout(n1523),.clk(gclk));
	jand g1223(.dina(n1523),.dinb(n1519),.dout(n1524),.clk(gclk));
	jxor g1224(.dina(n1524),.dinb(n1515),.dout(n1525),.clk(gclk));
	jor g1225(.dina(w_n483_1[0]),.dinb(w_n369_0[2]),.dout(n1526),.clk(gclk));
	jor g1226(.dina(w_G265_0[2]),.dinb(w_n366_0[2]),.dout(n1527),.clk(gclk));
	jand g1227(.dina(n1527),.dinb(w_G400_0[1]),.dout(n1528),.clk(gclk));
	jand g1228(.dina(n1528),.dinb(n1526),.dout(n1529),.clk(gclk));
	jor g1229(.dina(w_G265_0[1]),.dinb(w_G254_0[2]),.dout(n1530),.clk(gclk));
	jor g1230(.dina(w_n483_0[2]),.dinb(w_G242_0[2]),.dout(n1531),.clk(gclk));
	jand g1231(.dina(n1531),.dinb(n1530),.dout(n1532),.clk(gclk));
	jand g1232(.dina(n1532),.dinb(w_n485_0[2]),.dout(n1533),.clk(gclk));
	jor g1233(.dina(n1533),.dinb(n1529),.dout(n1534),.clk(gclk));
	jand g1234(.dina(w_G257_1[0]),.dinb(w_G248_2[2]),.dout(n1535),.clk(gclk));
	jand g1235(.dina(w_n518_0[2]),.dinb(w_G251_2[2]),.dout(n1536),.clk(gclk));
	jor g1236(.dina(n1536),.dinb(w_n520_0[0]),.dout(n1537),.clk(gclk));
	jor g1237(.dina(n1537),.dinb(n1535),.dout(n1538),.clk(gclk));
	jand g1238(.dina(w_n518_0[1]),.dinb(w_n406_2[2]),.dout(n1539),.clk(gclk));
	jand g1239(.dina(w_G257_0[2]),.dinb(w_n408_2[2]),.dout(n1540),.clk(gclk));
	jor g1240(.dina(n1540),.dinb(n1539),.dout(n1541),.clk(gclk));
	jor g1241(.dina(n1541),.dinb(w_G389_0[1]),.dout(n1542),.clk(gclk));
	jand g1242(.dina(n1542),.dinb(n1538),.dout(n1543),.clk(gclk));
	jand g1243(.dina(w_G248_2[1]),.dinb(w_G234_1[0]),.dout(n1544),.clk(gclk));
	jand g1244(.dina(w_G251_2[1]),.dinb(w_n460_0[2]),.dout(n1545),.clk(gclk));
	jor g1245(.dina(n1545),.dinb(w_n462_0[0]),.dout(n1546),.clk(gclk));
	jor g1246(.dina(n1546),.dinb(n1544),.dout(n1547),.clk(gclk));
	jand g1247(.dina(w_n406_2[1]),.dinb(w_n460_0[1]),.dout(n1548),.clk(gclk));
	jand g1248(.dina(w_n408_2[1]),.dinb(w_G234_0[2]),.dout(n1549),.clk(gclk));
	jor g1249(.dina(n1549),.dinb(n1548),.dout(n1550),.clk(gclk));
	jor g1250(.dina(n1550),.dinb(w_G435_0[1]),.dout(n1551),.clk(gclk));
	jand g1251(.dina(n1551),.dinb(n1547),.dout(n1552),.clk(gclk));
	jxor g1252(.dina(n1552),.dinb(n1543),.dout(n1553),.clk(gclk));
	jxor g1253(.dina(n1553),.dinb(n1534),.dout(n1554),.clk(gclk));
	jxor g1254(.dina(n1554),.dinb(n1525),.dout(n1555),.clk(gclk));
	jand g1255(.dina(w_G248_2[0]),.dinb(w_G226_1[0]),.dout(n1556),.clk(gclk));
	jand g1256(.dina(w_G251_2[0]),.dinb(w_n494_0[2]),.dout(n1557),.clk(gclk));
	jor g1257(.dina(n1557),.dinb(w_n496_0[1]),.dout(n1558),.clk(gclk));
	jor g1258(.dina(n1558),.dinb(n1556),.dout(n1559),.clk(gclk));
	jand g1259(.dina(w_n406_2[0]),.dinb(w_n494_0[1]),.dout(n1560),.clk(gclk));
	jand g1260(.dina(w_n408_2[0]),.dinb(w_G226_0[2]),.dout(n1561),.clk(gclk));
	jor g1261(.dina(n1561),.dinb(n1560),.dout(n1562),.clk(gclk));
	jor g1262(.dina(n1562),.dinb(w_G422_0[1]),.dout(n1563),.clk(gclk));
	jand g1263(.dina(n1563),.dinb(n1559),.dout(n1564),.clk(gclk));
	jxor g1264(.dina(n1564),.dinb(w_n551_0[0]),.dout(n1565),.clk(gclk));
	jor g1265(.dina(w_n369_0[1]),.dinb(w_n507_0[2]),.dout(n1566),.clk(gclk));
	jor g1266(.dina(w_n366_0[1]),.dinb(w_G218_1[0]),.dout(n1567),.clk(gclk));
	jand g1267(.dina(n1567),.dinb(w_G468_0[1]),.dout(n1568),.clk(gclk));
	jand g1268(.dina(n1568),.dinb(n1566),.dout(n1569),.clk(gclk));
	jor g1269(.dina(w_G254_0[1]),.dinb(w_G218_0[2]),.dout(n1570),.clk(gclk));
	jor g1270(.dina(w_G242_0[1]),.dinb(w_n507_0[1]),.dout(n1571),.clk(gclk));
	jand g1271(.dina(n1571),.dinb(n1570),.dout(n1572),.clk(gclk));
	jand g1272(.dina(n1572),.dinb(w_n509_0[0]),.dout(n1573),.clk(gclk));
	jor g1273(.dina(n1573),.dinb(n1569),.dout(n1574),.clk(gclk));
	jand g1274(.dina(w_G248_1[2]),.dinb(w_G210_1[0]),.dout(n1575),.clk(gclk));
	jand g1275(.dina(w_G251_1[2]),.dinb(w_n449_0[2]),.dout(n1576),.clk(gclk));
	jor g1276(.dina(n1576),.dinb(w_n451_0[0]),.dout(n1577),.clk(gclk));
	jor g1277(.dina(n1577),.dinb(n1575),.dout(n1578),.clk(gclk));
	jand g1278(.dina(w_n406_1[2]),.dinb(w_n449_0[1]),.dout(n1579),.clk(gclk));
	jand g1279(.dina(w_n408_1[2]),.dinb(w_G210_0[2]),.dout(n1580),.clk(gclk));
	jor g1280(.dina(n1580),.dinb(n1579),.dout(n1581),.clk(gclk));
	jor g1281(.dina(n1581),.dinb(w_G457_0[1]),.dout(n1582),.clk(gclk));
	jand g1282(.dina(n1582),.dinb(n1578),.dout(n1583),.clk(gclk));
	jxor g1283(.dina(n1583),.dinb(n1574),.dout(n1584),.clk(gclk));
	jxor g1284(.dina(n1584),.dinb(n1565),.dout(n1585),.clk(gclk));
	jxor g1285(.dina(n1585),.dinb(n1555),.dout(n1586),.clk(gclk));
	jand g1286(.dina(n1586),.dinb(w_n749_4[2]),.dout(n1587),.clk(gclk));
	jnot g1287(.din(n1587),.dout(n1588),.clk(gclk));
	jand g1288(.dina(w_n573_0[0]),.dinb(w_n567_0[0]),.dout(n1589),.clk(gclk));
	jor g1289(.dina(n1589),.dinb(w_n699_0[0]),.dout(n1590),.clk(gclk));
	jnot g1290(.din(w_n559_0[0]),.dout(n1591),.clk(gclk));
	jor g1291(.dina(n1591),.dinb(w_n557_0[0]),.dout(n1592),.clk(gclk));
	jand g1292(.dina(w_n1592_0[1]),.dinb(w_n532_0[2]),.dout(n1593),.clk(gclk));
	jnot g1293(.din(w_n1593_0[1]),.dout(n1594),.clk(gclk));
	jor g1294(.dina(w_n695_0[0]),.dinb(n1594),.dout(n1595),.clk(gclk));
	jand g1295(.dina(w_n923_0[1]),.dinb(w_n473_0[2]),.dout(n1596),.clk(gclk));
	jor g1296(.dina(w_n1596_0[1]),.dinb(w_n1593_0[0]),.dout(n1597),.clk(gclk));
	jand g1297(.dina(n1597),.dinb(n1595),.dout(n1598),.clk(gclk));
	jxor g1298(.dina(n1598),.dinb(n1590),.dout(n1599),.clk(gclk));
	jnot g1299(.din(w_n1599_0[1]),.dout(n1600),.clk(gclk));
	jnot g1300(.din(w_n686_0[0]),.dout(n1601),.clk(gclk));
	jnot g1301(.din(w_n687_0[0]),.dout(n1602),.clk(gclk));
	jor g1302(.dina(w_n1592_0[0]),.dinb(w_n532_0[1]),.dout(n1603),.clk(gclk));
	jor g1303(.dina(w_n1596_0[0]),.dinb(w_n1603_0[1]),.dout(n1604),.clk(gclk));
	jor g1304(.dina(w_n923_0[0]),.dinb(w_n473_0[1]),.dout(n1605),.clk(gclk));
	jor g1305(.dina(w_n689_0[0]),.dinb(w_n485_0[1]),.dout(n1606),.clk(gclk));
	jand g1306(.dina(n1606),.dinb(w_n1605_0[1]),.dout(n1607),.clk(gclk));
	jand g1307(.dina(n1607),.dinb(n1604),.dout(n1608),.clk(gclk));
	jor g1308(.dina(n1608),.dinb(w_n690_0[0]),.dout(n1609),.clk(gclk));
	jor g1309(.dina(w_n1609_0[1]),.dinb(n1602),.dout(n1610),.clk(gclk));
	jand g1310(.dina(n1610),.dinb(n1601),.dout(n1611),.clk(gclk));
	jand g1311(.dina(w_n1611_0[2]),.dinb(w_n581_0[0]),.dout(n1612),.clk(gclk));
	jxor g1312(.dina(w_n566_0[0]),.dinb(w_n561_0[1]),.dout(n1613),.clk(gclk));
	jxor g1313(.dina(w_n1613_0[1]),.dinb(w_n865_0[1]),.dout(n1614),.clk(gclk));
	jxor g1314(.dina(n1614),.dinb(n1612),.dout(n1615),.clk(gclk));
	jnot g1315(.din(w_n1615_0[1]),.dout(n1616),.clk(gclk));
	jand g1316(.dina(n1616),.dinb(n1600),.dout(n1617),.clk(gclk));
	jnot g1317(.din(w_G1497_0[2]),.dout(n1618),.clk(gclk));
	jand g1318(.dina(w_n1615_0[0]),.dinb(w_n1599_0[0]),.dout(n1619),.clk(gclk));
	jor g1319(.dina(n1619),.dinb(w_n1618_0[1]),.dout(n1620),.clk(gclk));
	jor g1320(.dina(n1620),.dinb(n1617),.dout(n1621),.clk(gclk));
	jand g1321(.dina(w_n1605_0[0]),.dinb(w_n1603_0[0]),.dout(n1622),.clk(gclk));
	jor g1322(.dina(n1622),.dinb(w_n694_0[0]),.dout(n1623),.clk(gclk));
	jxor g1323(.dina(w_n1613_0[0]),.dinb(w_n1609_0[0]),.dout(n1624),.clk(gclk));
	jxor g1324(.dina(n1624),.dinb(n1623),.dout(n1625),.clk(gclk));
	jxor g1325(.dina(w_n1611_0[1]),.dinb(w_n865_0[0]),.dout(n1626),.clk(gclk));
	jxor g1326(.dina(n1626),.dinb(n1625),.dout(n1627),.clk(gclk));
	jor g1327(.dina(n1627),.dinb(w_G1497_0[1]),.dout(n1628),.clk(gclk));
	jand g1328(.dina(n1628),.dinb(n1621),.dout(n1629),.clk(gclk));
	jxor g1329(.dina(w_n579_0[1]),.dinb(w_n574_0[0]),.dout(n1630),.clk(gclk));
	jxor g1330(.dina(n1630),.dinb(n1629),.dout(n1631),.clk(gclk));
	jnot g1331(.din(w_n709_0[0]),.dout(n1632),.clk(gclk));
	jand g1332(.dina(n1632),.dinb(w_n953_0[0]),.dout(n1633),.clk(gclk));
	jand g1333(.dina(w_n711_0[0]),.dinb(w_n954_0[1]),.dout(n1634),.clk(gclk));
	jor g1334(.dina(n1634),.dinb(w_n1633_0[1]),.dout(n1635),.clk(gclk));
	jxor g1335(.dina(w_n608_0[0]),.dinb(w_n592_0[0]),.dout(n1636),.clk(gclk));
	jxor g1336(.dina(n1636),.dinb(w_n602_0[0]),.dout(n1637),.clk(gclk));
	jxor g1337(.dina(w_n1637_0[1]),.dinb(n1635),.dout(n1638),.clk(gclk));
	jor g1338(.dina(w_n938_0[1]),.dinb(w_n597_0[0]),.dout(n1639),.clk(gclk));
	jand g1339(.dina(w_n609_0[0]),.dinb(w_n962_0[0]),.dout(n1640),.clk(gclk));
	jor g1340(.dina(n1640),.dinb(w_n715_0[0]),.dout(n1641),.clk(gclk));
	jand g1341(.dina(n1641),.dinb(n1639),.dout(n1642),.clk(gclk));
	jxor g1342(.dina(n1642),.dinb(n1638),.dout(n1643),.clk(gclk));
	jand g1343(.dina(w_n1643_0[1]),.dinb(w_n703_0[1]),.dout(n1644),.clk(gclk));
	jnot g1344(.din(w_n682_0[0]),.dout(n1645),.clk(gclk));
	jor g1345(.dina(w_n1611_0[0]),.dinb(w_n684_0[0]),.dout(n1646),.clk(gclk));
	jand g1346(.dina(n1646),.dinb(n1645),.dout(n1647),.clk(gclk));
	jand g1347(.dina(w_n713_0[0]),.dinb(w_n954_0[0]),.dout(n1648),.clk(gclk));
	jor g1348(.dina(n1648),.dinb(w_n1633_0[0]),.dout(n1649),.clk(gclk));
	jxor g1349(.dina(n1649),.dinb(w_n938_0[0]),.dout(n1650),.clk(gclk));
	jxor g1350(.dina(n1650),.dinb(w_n1637_0[0]),.dout(n1651),.clk(gclk));
	jand g1351(.dina(n1651),.dinb(n1647),.dout(n1652),.clk(gclk));
	jor g1352(.dina(w_n1652_0[1]),.dinb(n1644),.dout(n1653),.clk(gclk));
	jor g1353(.dina(n1653),.dinb(w_G1497_0[0]),.dout(n1654),.clk(gclk));
	jnot g1354(.din(w_n588_1[0]),.dout(n1655),.clk(gclk));
	jand g1355(.dina(w_n1652_0[0]),.dinb(n1655),.dout(n1656),.clk(gclk));
	jor g1356(.dina(w_n703_0[0]),.dinb(w_n588_0[2]),.dout(n1657),.clk(gclk));
	jand g1357(.dina(n1657),.dinb(w_n1643_0[0]),.dout(n1658),.clk(gclk));
	jor g1358(.dina(n1658),.dinb(n1656),.dout(n1659),.clk(gclk));
	jor g1359(.dina(n1659),.dinb(w_n1618_0[0]),.dout(n1660),.clk(gclk));
	jand g1360(.dina(n1660),.dinb(n1654),.dout(n1661),.clk(gclk));
	jxor g1361(.dina(n1661),.dinb(n1631),.dout(n1662),.clk(gclk));
	jor g1362(.dina(n1662),.dinb(w_n749_4[1]),.dout(n1663),.clk(gclk));
	jand g1363(.dina(n1663),.dinb(n1588),.dout(n1664),.clk(gclk));
	jor g1364(.dina(n1664),.dinb(w_G4092_3[2]),.dout(n1665),.clk(gclk));
	jor g1365(.dina(w_n1504_0[0]),.dinb(G118),.dout(n1666),.clk(gclk));
	jand g1366(.dina(w_dff_B_shEHb3tA0_0),.dinb(w_n1665_0[1]),.dout(w_dff_A_vmfcvb7t4_2),.clk(gclk));
	jor g1367(.dina(w_G4088_3[1]),.dinb(w_G14_0[1]),.dout(n1668),.clk(gclk));
	jor g1368(.dina(w_n797_3[1]),.dinb(w_G64_0[1]),.dout(n1669),.clk(gclk));
	jand g1369(.dina(n1669),.dinb(w_G4087_1[1]),.dout(n1670),.clk(gclk));
	jand g1370(.dina(n1670),.dinb(n1668),.dout(n1671),.clk(gclk));
	jand g1371(.dina(w_G4092_3[1]),.dinb(G97),.dout(n1672),.clk(gclk));
	jnot g1372(.din(n1672),.dout(n1673),.clk(gclk));
	jand g1373(.dina(n1673),.dinb(w_n1665_0[0]),.dout(n1674),.clk(gclk));
	jnot g1374(.din(w_n1674_0[2]),.dout(n1675),.clk(gclk));
	jor g1375(.dina(w_n1675_0[1]),.dinb(w_n797_3[0]),.dout(n1676),.clk(gclk));
	jand g1376(.dina(w_G4092_3[0]),.dinb(G94),.dout(n1677),.clk(gclk));
	jnot g1377(.din(n1677),.dout(n1678),.clk(gclk));
	jand g1378(.dina(w_dff_B_11Y5fuYu3_0),.dinb(w_n1503_0[0]),.dout(n1679),.clk(gclk));
	jnot g1379(.din(w_n1679_0[2]),.dout(n1680),.clk(gclk));
	jor g1380(.dina(w_n1680_0[1]),.dinb(w_G4088_3[0]),.dout(n1681),.clk(gclk));
	jand g1381(.dina(n1681),.dinb(w_n800_1[1]),.dout(n1682),.clk(gclk));
	jand g1382(.dina(n1682),.dinb(w_dff_B_EEzYRZkM4_1),.dout(n1683),.clk(gclk));
	jor g1383(.dina(n1683),.dinb(w_dff_B_MSftF2H93_1),.dout(w_dff_A_RE0tB8YO4_2),.clk(gclk));
	jor g1384(.dina(w_G4089_3[1]),.dinb(w_G14_0[0]),.dout(n1685),.clk(gclk));
	jor g1385(.dina(w_n852_3[1]),.dinb(w_G64_0[0]),.dout(n1686),.clk(gclk));
	jand g1386(.dina(n1686),.dinb(w_G4090_1[1]),.dout(n1687),.clk(gclk));
	jand g1387(.dina(n1687),.dinb(n1685),.dout(n1688),.clk(gclk));
	jor g1388(.dina(w_n1675_0[0]),.dinb(w_n852_3[0]),.dout(n1689),.clk(gclk));
	jor g1389(.dina(w_n1680_0[0]),.dinb(w_G4089_3[0]),.dout(n1690),.clk(gclk));
	jand g1390(.dina(n1690),.dinb(w_n854_1[1]),.dout(n1691),.clk(gclk));
	jand g1391(.dina(n1691),.dinb(w_dff_B_HgvF8hE49_1),.dout(n1692),.clk(gclk));
	jor g1392(.dina(n1692),.dinb(w_dff_B_IcnpIemx3_1),.dout(w_dff_A_pwFU8BN14_2),.clk(gclk));
	jnot g1393(.din(w_G137_3[1]),.dout(n1694),.clk(gclk));
	jnot g1394(.din(G179),.dout(n1695),.clk(gclk));
	jnot g1395(.din(w_n996_1[1]),.dout(n1696),.clk(gclk));
	jor g1396(.dina(n1696),.dinb(w_n1695_0[1]),.dout(n1697),.clk(gclk));
	jnot g1397(.din(G176),.dout(n1698),.clk(gclk));
	jnot g1398(.din(w_n994_1[1]),.dout(n1699),.clk(gclk));
	jor g1399(.dina(n1699),.dinb(w_n1698_0[1]),.dout(n1700),.clk(gclk));
	jand g1400(.dina(w_n1674_0[1]),.dinb(w_G1689_1[2]),.dout(n1701),.clk(gclk));
	jand g1401(.dina(w_n1679_0[1]),.dinb(w_n993_1[1]),.dout(n1702),.clk(gclk));
	jor g1402(.dina(n1702),.dinb(w_G1690_0[1]),.dout(n1703),.clk(gclk));
	jor g1403(.dina(n1703),.dinb(w_dff_B_OyrKFmYT7_1),.dout(n1704),.clk(gclk));
	jand g1404(.dina(n1704),.dinb(w_dff_B_S1TlZL3Q5_1),.dout(n1705),.clk(gclk));
	jand g1405(.dina(n1705),.dinb(w_dff_B_xFRH1E7d1_1),.dout(n1706),.clk(gclk));
	jor g1406(.dina(n1706),.dinb(w_n1694_0[1]),.dout(G658),.clk(gclk));
	jnot g1407(.din(w_n1012_1[1]),.dout(n1708),.clk(gclk));
	jor g1408(.dina(n1708),.dinb(w_n1695_0[0]),.dout(n1709),.clk(gclk));
	jnot g1409(.din(w_n1014_1[1]),.dout(n1710),.clk(gclk));
	jor g1410(.dina(n1710),.dinb(w_n1698_0[0]),.dout(n1711),.clk(gclk));
	jand g1411(.dina(w_n1674_0[0]),.dinb(w_G1691_1[2]),.dout(n1712),.clk(gclk));
	jand g1412(.dina(w_n1679_0[0]),.dinb(w_n1008_1[1]),.dout(n1713),.clk(gclk));
	jor g1413(.dina(n1713),.dinb(w_G1694_0[1]),.dout(n1714),.clk(gclk));
	jor g1414(.dina(n1714),.dinb(w_dff_B_qck1SFfG3_1),.dout(n1715),.clk(gclk));
	jand g1415(.dina(n1715),.dinb(w_dff_B_UhhF2aeY9_1),.dout(n1716),.clk(gclk));
	jand g1416(.dina(n1716),.dinb(w_dff_B_5wark3kh5_1),.dout(n1717),.clk(gclk));
	jor g1417(.dina(n1717),.dinb(w_n1694_0[0]),.dout(G690),.clk(gclk));
	jdff g1418(.din(w_G141_1[0]),.dout(w_dff_A_tFCKOFNL4_1));
	jdff g1419(.din(w_G293_0[0]),.dout(w_dff_A_Bir94Gwe0_1));
	jdff g1420(.din(w_G3173_0[0]),.dout(w_dff_A_H773dteS1_1));
	jnot g1421(.din(w_G545_0[1]),.dout(w_dff_A_5wc4wnAA5_1),.clk(gclk));
	jnot g1422(.din(w_G545_0[0]),.dout(w_dff_A_iFcdHZpN8_1),.clk(gclk));
	jdff g1423(.din(w_G137_3[0]),.dout(w_dff_A_TKuoKSCW6_1));
	jdff g1424(.din(w_G141_0[2]),.dout(w_dff_A_K6wpGJWd3_1));
	jdff g1425(.din(w_G1_2[0]),.dout(w_dff_A_7l1xJPxg8_1));
	jdff g1426(.din(w_G549_0[1]),.dout(w_dff_A_2dIO24Jj4_1));
	jdff g1427(.din(w_G299_0[1]),.dout(w_dff_A_lRm1ZvdP4_1));
	jnot g1428(.din(w_G549_0[0]),.dout(w_dff_A_VRuQeKNr1_1),.clk(gclk));
	jdff g1429(.din(w_G1_1[2]),.dout(w_dff_A_kHDc557D8_1));
	jdff g1430(.din(w_G1_1[1]),.dout(w_dff_A_GL80qaD07_1));
	jdff g1431(.din(w_G1_1[0]),.dout(w_dff_A_DSogMvSP0_1));
	jdff g1432(.din(w_G1_0[2]),.dout(w_dff_A_icCkjrtN9_1));
	jdff g1433(.din(w_G299_0[0]),.dout(w_dff_A_fys1SLwP5_1));
	jor g1434(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(w_dff_A_3bTGddH80_2),.clk(gclk));
	jand g1435(.dina(w_n661_0[0]),.dinb(w_n641_0[1]),.dout(w_dff_A_6f5g0anK1_2),.clk(gclk));
	jand g1436(.dina(w_n611_0[0]),.dinb(w_n588_0[1]),.dout(w_dff_A_gMde8Pq87_2),.clk(gclk));
	jor g1437(.dina(w_n717_0[0]),.dinb(w_n704_0[0]),.dout(w_dff_A_SEr1vClL9_2),.clk(gclk));
	jor g1438(.dina(w_n747_0[0]),.dinb(w_n738_0[0]),.dout(w_dff_A_FP0rTFvM2_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_G4_0[1]),.doutc(w_G4_0[2]),.din(G4));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(G11));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(G14));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(G17));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(G20));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(G37));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(G40));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(G43));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(G46));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(G49));
	jspl3 jspl3_w_G54_0(.douta(w_G54_0[0]),.doutb(w_G54_0[1]),.doutc(w_G54_0[2]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(G61));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(G64));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(G67));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(G70));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(G73));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(G76));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(G91));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(G100));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(G103));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(G106));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(G109));
	jspl jspl_w_G123_0(.douta(w_G123_0[0]),.doutb(w_G123_0[1]),.din(G123));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_x9nhREvs5_0),.doutb(w_dff_A_2ZM4WqgQ8_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_dH68NgwT8_0),.doutb(w_dff_A_Exb9jyy65_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_G137_3[2]),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_dff_A_2eqtmcpk1_0),.doutb(w_dff_A_XR3oOArB3_1),.doutc(w_G137_4[2]),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_dff_A_vqLHpnx04_0),.doutb(w_G137_5[1]),.doutc(w_G137_5[2]),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_xKN9JgQ47_0),.doutb(w_dff_A_YvJlGhkA9_1),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_0JDJpoad9_1),.doutc(w_dff_A_r8xWbjbI8_2),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_G137_8[0]),.doutb(w_G137_8[1]),.doutc(w_dff_A_CbUuo9Gv3_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_G137_9[0]),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_Z7jBtOZN9_1),.doutc(w_dff_A_NDNz4G301_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_NY7cL5aH0_0),.doutb(w_dff_A_nCk6XHLC6_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(G146));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(G149));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(G152));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(G155));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(G158));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(G161));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(G164));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(G167));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(G170));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(G173));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(G182));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(G185));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(G188));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(G191));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(G194));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(G197));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(G200));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(G203));
	jspl3 jspl3_w_G206_0(.douta(w_G206_0[0]),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G206_1(.douta(w_G206_1[0]),.doutb(w_G206_1[1]),.doutc(w_G206_1[2]),.din(w_G206_0[0]));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_G210_0[2]),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_G210_1[1]),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl jspl_w_G210_2(.douta(w_G210_2[0]),.doutb(w_G210_2[1]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_G218_1[0]),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl jspl_w_G218_2(.douta(w_G218_2[0]),.doutb(w_G218_2[1]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_G226_0[2]),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_G226_1[0]),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl jspl_w_G226_2(.douta(w_G226_2[0]),.doutb(w_G226_2[1]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_G234_0[2]),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_G234_2[0]),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_G242_0[1]),.doutc(w_G242_0[2]),.din(G242));
	jspl jspl_w_G242_1(.douta(w_G242_1[0]),.doutb(w_G242_1[1]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_G245_0[0]),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_G248_3[2]),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl3 jspl3_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.doutc(w_G248_5[2]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_G251_0[1]),.doutc(w_G251_0[2]),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_G251_1[0]),.doutb(w_G251_1[1]),.doutc(w_G251_1[2]),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_G251_4[1]),.doutc(w_G251_4[2]),.din(w_G251_1[0]));
	jspl jspl_w_G251_5(.douta(w_G251_5[0]),.doutb(w_G251_5[1]),.din(w_G251_1[1]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl jspl_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_G257_0[2]),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_G257_1[0]),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl jspl_w_G257_2(.douta(w_G257_2[0]),.doutb(w_G257_2[1]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_G265_0[2]),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_G265_1[1]),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_G273_0[2]),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_G273_1[1]),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl jspl_w_G273_2(.douta(w_G273_2[0]),.doutb(w_G273_2[1]),.din(w_G273_0[1]));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_G281_0[2]),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_G281_2[0]),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_G289_0[0]),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_G293_0[1]),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_G302_0[0]),.doutb(w_G302_0[1]),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_G308_1[0]),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_G316_0[2]),.din(G316));
	jspl jspl_w_G316_1(.douta(w_G316_1[0]),.doutb(w_G316_1[1]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_G324_0[1]),.doutc(w_G324_0[2]),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_G324_1[1]),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_G331_0[1]),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_G332_1[1]),.doutc(w_G332_1[2]),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_G332_2[0]),.doutb(w_G332_2[1]),.doutc(w_G332_2[2]),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_G332_3[0]),.doutb(w_G332_3[1]),.doutc(w_G332_3[2]),.din(w_G332_0[2]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl jspl_w_G338_0(.douta(w_G338_0[0]),.doutb(w_G338_0[1]),.din(G338));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_G341_0[2]),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_G341_2[1]),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_G348_0[0]),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_G351_0[2]),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_G351_1[0]),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_G351_2[1]),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_G358_0[0]),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_G361_0[1]),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G361_1(.douta(w_G361_1[0]),.doutb(w_G361_1[1]),.din(w_G361_0[0]));
	jspl jspl_w_G366_0(.douta(w_G366_0[0]),.doutb(w_G366_0[1]),.din(G366));
	jspl jspl_w_G369_0(.douta(w_G369_0[0]),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_G374_0[0]),.doutb(w_G374_0[1]),.doutc(w_G374_0[2]),.din(G374));
	jspl3 jspl3_w_G374_1(.douta(w_G374_1[0]),.doutb(w_G374_1[1]),.doutc(w_G374_1[2]),.din(w_G374_0[0]));
	jspl3 jspl3_w_G389_0(.douta(w_G389_0[0]),.doutb(w_G389_0[1]),.doutc(w_G389_0[2]),.din(G389));
	jspl3 jspl3_w_G389_1(.douta(w_G389_1[0]),.doutb(w_G389_1[1]),.doutc(w_G389_1[2]),.din(w_G389_0[0]));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_G400_0[1]),.doutc(w_G400_0[2]),.din(G400));
	jspl3 jspl3_w_G400_1(.douta(w_G400_1[0]),.doutb(w_G400_1[1]),.doutc(w_G400_1[2]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_G411_0[0]),.doutb(w_G411_0[1]),.doutc(w_G411_0[2]),.din(G411));
	jspl3 jspl3_w_G411_1(.douta(w_G411_1[0]),.doutb(w_G411_1[1]),.doutc(w_G411_1[2]),.din(w_G411_0[0]));
	jspl jspl_w_G411_2(.douta(w_G411_2[0]),.doutb(w_G411_2[1]),.din(w_G411_0[1]));
	jspl3 jspl3_w_G422_0(.douta(w_G422_0[0]),.doutb(w_G422_0[1]),.doutc(w_G422_0[2]),.din(G422));
	jspl jspl_w_G422_1(.douta(w_G422_1[0]),.doutb(w_G422_1[1]),.din(w_G422_0[0]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_G435_0[1]),.doutc(w_G435_0[2]),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_G435_1[0]),.doutb(w_G435_1[1]),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_G446_0[1]),.doutc(w_G446_0[2]),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_G446_1[0]),.doutb(w_G446_1[1]),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_G457_0[0]),.doutb(w_G457_0[1]),.doutc(w_G457_0[2]),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_G457_1[0]),.doutb(w_G457_1[1]),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_G468_0[1]),.doutc(w_G468_0[2]),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_G468_1[0]),.doutb(w_G468_1[1]),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_G479_0[0]),.doutb(w_G479_0[1]),.doutc(w_G479_0[2]),.din(G479));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_G490_0[1]),.doutc(w_G490_0[2]),.din(G490));
	jspl jspl_w_G490_1(.douta(w_G490_1[0]),.doutb(w_G490_1[1]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_G503_0[0]),.doutb(w_G503_0[1]),.doutc(w_G503_0[2]),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_G503_1[0]),.doutb(w_G503_1[1]),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl jspl_w_G503_2(.douta(w_G503_2[0]),.doutb(w_G503_2[1]),.din(w_G503_0[1]));
	jspl3 jspl3_w_G514_0(.douta(w_G514_0[0]),.doutb(w_G514_0[1]),.doutc(w_G514_0[2]),.din(G514));
	jspl3 jspl3_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.doutc(w_G514_1[2]),.din(w_G514_0[0]));
	jspl jspl_w_G514_2(.douta(w_G514_2[0]),.doutb(w_G514_2[1]),.din(w_G514_0[1]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_G523_0[1]),.doutc(w_G523_0[2]),.din(G523));
	jspl3 jspl3_w_G523_1(.douta(w_G523_1[0]),.doutb(w_G523_1[1]),.doutc(w_G523_1[2]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_G534_0[0]),.doutb(w_G534_0[1]),.doutc(w_G534_0[2]),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_G534_1[0]),.doutb(w_G534_1[1]),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl jspl_w_G534_2(.douta(w_G534_2[0]),.doutb(w_G534_2[1]),.din(w_G534_0[1]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_dff_A_XYykHfUK1_0),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_G1497_0[0]),.doutb(w_G1497_0[1]),.doutc(w_G1497_0[2]),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_G1689_0[1]),.doutc(w_G1689_0[2]),.din(G1689));
	jspl3 jspl3_w_G1689_1(.douta(w_G1689_1[0]),.doutb(w_G1689_1[1]),.doutc(w_G1689_1[2]),.din(w_G1689_0[0]));
	jspl3 jspl3_w_G1689_2(.douta(w_dff_A_EGN9FuvV8_0),.doutb(w_G1689_2[1]),.doutc(w_dff_A_M0L6Ldl49_2),.din(w_G1689_0[1]));
	jspl3 jspl3_w_G1689_3(.douta(w_dff_A_iU8dCjJT9_0),.doutb(w_dff_A_jF0uhBbI8_1),.doutc(w_G1689_3[2]),.din(w_G1689_0[2]));
	jspl3 jspl3_w_G1689_4(.douta(w_dff_A_ULX69nvB6_0),.doutb(w_dff_A_JdFhaelb0_1),.doutc(w_G1689_4[2]),.din(w_G1689_1[0]));
	jspl jspl_w_G1689_5(.douta(w_G1689_5[0]),.doutb(w_G1689_5[1]),.din(w_G1689_1[1]));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_G1690_0[1]),.doutc(w_G1690_0[2]),.din(G1690));
	jspl jspl_w_G1690_1(.douta(w_G1690_1[0]),.doutb(w_G1690_1[1]),.din(w_G1690_0[0]));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_G1691_0[1]),.doutc(w_G1691_0[2]),.din(G1691));
	jspl3 jspl3_w_G1691_1(.douta(w_G1691_1[0]),.doutb(w_G1691_1[1]),.doutc(w_G1691_1[2]),.din(w_G1691_0[0]));
	jspl3 jspl3_w_G1691_2(.douta(w_dff_A_HRL9jvSt8_0),.doutb(w_G1691_2[1]),.doutc(w_dff_A_JgzjklZa3_2),.din(w_G1691_0[1]));
	jspl3 jspl3_w_G1691_3(.douta(w_dff_A_55ySoC9q4_0),.doutb(w_dff_A_2iyUexrb4_1),.doutc(w_G1691_3[2]),.din(w_G1691_0[2]));
	jspl3 jspl3_w_G1691_4(.douta(w_G1691_4[0]),.doutb(w_G1691_4[1]),.doutc(w_G1691_4[2]),.din(w_G1691_1[0]));
	jspl jspl_w_G1691_5(.douta(w_G1691_5[0]),.doutb(w_G1691_5[1]),.din(w_G1691_1[1]));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_G1694_0[1]),.doutc(w_G1694_0[2]),.din(G1694));
	jspl jspl_w_G1694_1(.douta(w_G1694_1[0]),.doutb(w_G1694_1[1]),.din(w_G1694_0[0]));
	jspl3 jspl3_w_G2174_0(.douta(w_G2174_0[0]),.doutb(w_G2174_0[1]),.doutc(w_G2174_0[2]),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_G2358_2[0]),.doutb(w_G2358_2[1]),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(G3548));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_G3717_0[0]),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_G3724_0[0]),.doutb(w_G3724_0[1]),.doutc(w_G3724_0[2]),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_G4087_0[1]),.doutc(w_G4087_0[2]),.din(G4087));
	jspl3 jspl3_w_G4087_1(.douta(w_G4087_1[0]),.doutb(w_G4087_1[1]),.doutc(w_G4087_1[2]),.din(w_G4087_0[0]));
	jspl3 jspl3_w_G4087_2(.douta(w_G4087_2[0]),.doutb(w_G4087_2[1]),.doutc(w_G4087_2[2]),.din(w_G4087_0[1]));
	jspl3 jspl3_w_G4087_3(.douta(w_G4087_3[0]),.doutb(w_G4087_3[1]),.doutc(w_G4087_3[2]),.din(w_G4087_0[2]));
	jspl3 jspl3_w_G4087_4(.douta(w_G4087_4[0]),.doutb(w_G4087_4[1]),.doutc(w_G4087_4[2]),.din(w_G4087_1[0]));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_G4088_0[2]),.din(G4088));
	jspl3 jspl3_w_G4088_1(.douta(w_G4088_1[0]),.doutb(w_G4088_1[1]),.doutc(w_G4088_1[2]),.din(w_G4088_0[0]));
	jspl3 jspl3_w_G4088_2(.douta(w_G4088_2[0]),.doutb(w_G4088_2[1]),.doutc(w_G4088_2[2]),.din(w_G4088_0[1]));
	jspl3 jspl3_w_G4088_3(.douta(w_G4088_3[0]),.doutb(w_G4088_3[1]),.doutc(w_G4088_3[2]),.din(w_G4088_0[2]));
	jspl3 jspl3_w_G4088_4(.douta(w_G4088_4[0]),.doutb(w_G4088_4[1]),.doutc(w_G4088_4[2]),.din(w_G4088_1[0]));
	jspl3 jspl3_w_G4088_5(.douta(w_G4088_5[0]),.doutb(w_G4088_5[1]),.doutc(w_G4088_5[2]),.din(w_G4088_1[1]));
	jspl3 jspl3_w_G4088_6(.douta(w_G4088_6[0]),.doutb(w_G4088_6[1]),.doutc(w_G4088_6[2]),.din(w_G4088_1[2]));
	jspl3 jspl3_w_G4088_7(.douta(w_G4088_7[0]),.doutb(w_G4088_7[1]),.doutc(w_G4088_7[2]),.din(w_G4088_2[0]));
	jspl3 jspl3_w_G4088_8(.douta(w_G4088_8[0]),.doutb(w_G4088_8[1]),.doutc(w_G4088_8[2]),.din(w_G4088_2[1]));
	jspl3 jspl3_w_G4088_9(.douta(w_G4088_9[0]),.doutb(w_G4088_9[1]),.doutc(w_G4088_9[2]),.din(w_G4088_2[2]));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_G4089_0[2]),.din(G4089));
	jspl3 jspl3_w_G4089_1(.douta(w_G4089_1[0]),.doutb(w_G4089_1[1]),.doutc(w_G4089_1[2]),.din(w_G4089_0[0]));
	jspl3 jspl3_w_G4089_2(.douta(w_G4089_2[0]),.doutb(w_G4089_2[1]),.doutc(w_G4089_2[2]),.din(w_G4089_0[1]));
	jspl3 jspl3_w_G4089_3(.douta(w_G4089_3[0]),.doutb(w_G4089_3[1]),.doutc(w_G4089_3[2]),.din(w_G4089_0[2]));
	jspl3 jspl3_w_G4089_4(.douta(w_G4089_4[0]),.doutb(w_G4089_4[1]),.doutc(w_G4089_4[2]),.din(w_G4089_1[0]));
	jspl3 jspl3_w_G4089_5(.douta(w_G4089_5[0]),.doutb(w_G4089_5[1]),.doutc(w_G4089_5[2]),.din(w_G4089_1[1]));
	jspl3 jspl3_w_G4089_6(.douta(w_G4089_6[0]),.doutb(w_G4089_6[1]),.doutc(w_G4089_6[2]),.din(w_G4089_1[2]));
	jspl3 jspl3_w_G4089_7(.douta(w_G4089_7[0]),.doutb(w_G4089_7[1]),.doutc(w_G4089_7[2]),.din(w_G4089_2[0]));
	jspl3 jspl3_w_G4089_8(.douta(w_G4089_8[0]),.doutb(w_G4089_8[1]),.doutc(w_G4089_8[2]),.din(w_G4089_2[1]));
	jspl3 jspl3_w_G4089_9(.douta(w_G4089_9[0]),.doutb(w_G4089_9[1]),.doutc(w_G4089_9[2]),.din(w_G4089_2[2]));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_G4090_0[1]),.doutc(w_G4090_0[2]),.din(G4090));
	jspl3 jspl3_w_G4090_1(.douta(w_G4090_1[0]),.doutb(w_G4090_1[1]),.doutc(w_G4090_1[2]),.din(w_G4090_0[0]));
	jspl3 jspl3_w_G4090_2(.douta(w_G4090_2[0]),.doutb(w_G4090_2[1]),.doutc(w_G4090_2[2]),.din(w_G4090_0[1]));
	jspl3 jspl3_w_G4090_3(.douta(w_G4090_3[0]),.doutb(w_G4090_3[1]),.doutc(w_G4090_3[2]),.din(w_G4090_0[2]));
	jspl3 jspl3_w_G4090_4(.douta(w_G4090_4[0]),.doutb(w_G4090_4[1]),.doutc(w_G4090_4[2]),.din(w_G4090_1[0]));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_G4091_0[1]),.doutc(w_G4091_0[2]),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_G4091_1[0]),.doutb(w_G4091_1[1]),.doutc(w_G4091_1[2]),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_G4091_2[0]),.doutb(w_G4091_2[1]),.doutc(w_G4091_2[2]),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4091_3(.douta(w_G4091_3[0]),.doutb(w_G4091_3[1]),.doutc(w_G4091_3[2]),.din(w_G4091_0[2]));
	jspl3 jspl3_w_G4091_4(.douta(w_G4091_4[0]),.doutb(w_G4091_4[1]),.doutc(w_G4091_4[2]),.din(w_G4091_1[0]));
	jspl3 jspl3_w_G4091_5(.douta(w_G4091_5[0]),.doutb(w_G4091_5[1]),.doutc(w_G4091_5[2]),.din(w_G4091_1[1]));
	jspl jspl_w_G4091_6(.douta(w_G4091_6[0]),.doutb(w_G4091_6[1]),.din(w_G4091_1[2]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_G4092_0[1]),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_G4092_1[0]),.doutb(w_G4092_1[1]),.doutc(w_G4092_1[2]),.din(w_G4092_0[0]));
	jspl3 jspl3_w_G4092_2(.douta(w_G4092_2[0]),.doutb(w_G4092_2[1]),.doutc(w_G4092_2[2]),.din(w_G4092_0[1]));
	jspl3 jspl3_w_G4092_3(.douta(w_G4092_3[0]),.doutb(w_G4092_3[1]),.doutc(w_G4092_3[2]),.din(w_G4092_0[2]));
	jspl3 jspl3_w_G4092_4(.douta(w_G4092_4[0]),.doutb(w_G4092_4[1]),.doutc(w_G4092_4[2]),.din(w_G4092_1[0]));
	jspl3 jspl3_w_G4092_5(.douta(w_G4092_5[0]),.doutb(w_G4092_5[1]),.doutc(w_G4092_5[2]),.din(w_G4092_1[1]));
	jspl3 jspl3_w_G4092_6(.douta(w_G4092_6[0]),.doutb(w_G4092_6[1]),.doutc(w_G4092_6[2]),.din(w_G4092_1[2]));
	jspl3 jspl3_w_G4092_7(.douta(w_G4092_7[0]),.doutb(w_G4092_7[1]),.doutc(w_G4092_7[2]),.din(w_G4092_2[0]));
	jspl3 jspl3_w_G4092_8(.douta(w_G4092_8[0]),.doutb(w_G4092_8[1]),.doutc(w_G4092_8[2]),.din(w_G4092_2[1]));
	jspl3 jspl3_w_G4092_9(.douta(w_G4092_9[0]),.doutb(w_G4092_9[1]),.doutc(w_G4092_9[2]),.din(w_G4092_2[2]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(w_dff_A_QA8TyQ3f3_1),.din(G599_fa_));
	jspl jspl_w_G601_0(.douta(w_G601_0),.doutb(w_dff_A_B5zaQhi98_1),.din(G601_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(w_dff_A_aWb3Bder3_1),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_G809_1[0]),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_G809_2[2]),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_G809_3[0]),.doutb(w_G809_3[1]),.doutc(w_dff_A_yuNhCNJz3_2),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(w_dff_A_ugDvOh8h3_1),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(w_dff_A_VYShTGcq8_1),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(w_dff_A_UAv8zeNK0_1),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(w_dff_A_IgwmqSnl4_1),.din(G861_fa_));
	jspl jspl_w_G623_0(.douta(w_G623_0),.doutb(w_dff_A_b7Uj8T3n5_1),.din(G623_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(w_dff_A_TjtWKR5k2_1),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(w_dff_A_ICQfSecU6_1),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(w_dff_A_DX7YKSnO2_1),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(w_dff_A_zejxgGKu4_1),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(w_dff_A_GJ5SWN8q8_1),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(w_dff_A_Mw7p5bZZ9_1),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(w_dff_A_tYluNs5U4_1),.din(G877_fa_));
	jspl jspl_w_G998_0(.douta(w_G998_0),.doutb(w_dff_A_VCOqhx971_1),.din(G998_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(w_dff_A_CpoHOeGU4_1),.din(G830_fa_));
	jspl jspl_w_G865_0(.douta(w_G865_0),.doutb(w_dff_A_bx1a0Rhg8_1),.din(G865_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(w_dff_A_2o5mNUNN0_1),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(w_dff_B_8mCnqYH29_2));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.doutc(w_n369_0[2]),.din(n369));
	jspl3 jspl3_w_n369_1(.douta(w_n369_1[0]),.doutb(w_n369_1[1]),.doutc(w_n369_1[2]),.din(w_n369_0[0]));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl3 jspl3_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.doutc(w_n374_0[2]),.din(n374));
	jspl jspl_w_n374_1(.douta(w_n374_1[0]),.doutb(w_n374_1[1]),.din(w_n374_0[0]));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl3 jspl3_w_n375_1(.douta(w_n375_1[0]),.doutb(w_n375_1[1]),.doutc(w_n375_1[2]),.din(w_n375_0[0]));
	jspl3 jspl3_w_n375_2(.douta(w_n375_2[0]),.doutb(w_n375_2[1]),.doutc(w_n375_2[2]),.din(w_n375_0[1]));
	jspl3 jspl3_w_n375_3(.douta(w_n375_3[0]),.doutb(w_n375_3[1]),.doutc(w_n375_3[2]),.din(w_n375_0[2]));
	jspl3 jspl3_w_n375_4(.douta(w_n375_4[0]),.doutb(w_n375_4[1]),.doutc(w_n375_4[2]),.din(w_n375_1[0]));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_n377_0[2]),.din(n377));
	jspl jspl_w_n377_1(.douta(w_n377_1[0]),.doutb(w_n377_1[1]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.doutc(w_n378_0[2]),.din(n378));
	jspl3 jspl3_w_n378_1(.douta(w_n378_1[0]),.doutb(w_n378_1[1]),.doutc(w_n378_1[2]),.din(w_n378_0[0]));
	jspl3 jspl3_w_n378_2(.douta(w_n378_2[0]),.doutb(w_n378_2[1]),.doutc(w_n378_2[2]),.din(w_n378_0[1]));
	jspl3 jspl3_w_n378_3(.douta(w_n378_3[0]),.doutb(w_n378_3[1]),.doutc(w_n378_3[2]),.din(w_n378_0[2]));
	jspl3 jspl3_w_n378_4(.douta(w_n378_4[0]),.doutb(w_n378_4[1]),.doutc(w_n378_4[2]),.din(w_n378_1[0]));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_n389_0[2]),.din(n389));
	jspl jspl_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.din(w_n389_0[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.din(n401));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.doutc(w_n406_0[2]),.din(n406));
	jspl3 jspl3_w_n406_1(.douta(w_n406_1[0]),.doutb(w_n406_1[1]),.doutc(w_n406_1[2]),.din(w_n406_0[0]));
	jspl3 jspl3_w_n406_2(.douta(w_n406_2[0]),.doutb(w_n406_2[1]),.doutc(w_n406_2[2]),.din(w_n406_0[1]));
	jspl3 jspl3_w_n406_3(.douta(w_n406_3[0]),.doutb(w_n406_3[1]),.doutc(w_n406_3[2]),.din(w_n406_0[2]));
	jspl3 jspl3_w_n406_4(.douta(w_n406_4[0]),.doutb(w_n406_4[1]),.doutc(w_n406_4[2]),.din(w_n406_1[0]));
	jspl jspl_w_n406_5(.douta(w_n406_5[0]),.doutb(w_n406_5[1]),.din(w_n406_1[1]));
	jspl3 jspl3_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.doutc(w_n408_0[2]),.din(n408));
	jspl3 jspl3_w_n408_1(.douta(w_n408_1[0]),.doutb(w_n408_1[1]),.doutc(w_n408_1[2]),.din(w_n408_0[0]));
	jspl3 jspl3_w_n408_2(.douta(w_n408_2[0]),.doutb(w_n408_2[1]),.doutc(w_n408_2[2]),.din(w_n408_0[1]));
	jspl3 jspl3_w_n408_3(.douta(w_n408_3[0]),.doutb(w_n408_3[1]),.doutc(w_n408_3[2]),.din(w_n408_0[2]));
	jspl3 jspl3_w_n408_4(.douta(w_n408_4[0]),.doutb(w_n408_4[1]),.doutc(w_n408_4[2]),.din(w_n408_1[0]));
	jspl3 jspl3_w_n408_5(.douta(w_n408_5[0]),.doutb(w_n408_5[1]),.doutc(w_n408_5[2]),.din(w_n408_1[1]));
	jspl3 jspl3_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.doutc(w_n412_0[2]),.din(n412));
	jspl jspl_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.din(n414));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl3 jspl3_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.doutc(w_n423_0[2]),.din(n423));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_n425_0[2]),.din(n425));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.doutc(w_n428_0[2]),.din(n428));
	jspl jspl_w_n428_1(.douta(w_n428_1[0]),.doutb(w_n428_1[1]),.din(w_n428_0[0]));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl3 jspl3_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.doutc(w_n433_0[2]),.din(n433));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl jspl_w_n435_2(.douta(w_n435_2[0]),.doutb(w_n435_2[1]),.din(w_n435_0[1]));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_n451_0[1]),.doutc(w_n451_0[2]),.din(n451));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl3 jspl3_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.doutc(w_n471_1[2]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.doutc(w_n473_0[2]),.din(n473));
	jspl jspl_w_n473_1(.douta(w_n473_1[0]),.doutb(w_n473_1[1]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.doutc(w_n483_0[2]),.din(n483));
	jspl3 jspl3_w_n483_1(.douta(w_n483_1[0]),.doutb(w_n483_1[1]),.doutc(w_n483_1[2]),.din(w_n483_0[0]));
	jspl jspl_w_n483_2(.douta(w_n483_2[0]),.doutb(w_n483_2[1]),.din(w_n483_0[1]));
	jspl3 jspl3_w_n485_0(.douta(w_n485_0[0]),.doutb(w_n485_0[1]),.doutc(w_n485_0[2]),.din(n485));
	jspl jspl_w_n485_1(.douta(w_n485_1[0]),.doutb(w_n485_1[1]),.din(w_n485_0[0]));
	jspl jspl_w_n493_0(.douta(w_n493_0[0]),.doutb(w_n493_0[1]),.din(n493));
	jspl3 jspl3_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.doutc(w_n494_0[2]),.din(n494));
	jspl3 jspl3_w_n494_1(.douta(w_n494_1[0]),.doutb(w_n494_1[1]),.doutc(w_n494_1[2]),.din(w_n494_0[0]));
	jspl3 jspl3_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.doutc(w_n496_0[2]),.din(n496));
	jspl jspl_w_n496_1(.douta(w_n496_1[0]),.doutb(w_n496_1[1]),.din(w_n496_0[0]));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl3 jspl3_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.doutc(w_n509_0[2]),.din(n509));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl3 jspl3_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.doutc(w_n518_1[2]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.doutc(w_n520_0[2]),.din(n520));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl3 jspl3_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.doutc(w_n530_1[2]),.din(w_n530_0[0]));
	jspl3 jspl3_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.doutc(w_n532_0[2]),.din(n532));
	jspl jspl_w_n532_1(.douta(w_n532_1[0]),.doutb(w_n532_1[1]),.din(w_n532_0[0]));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.doutc(w_n551_0[2]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl3 jspl3_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.doutc(w_n556_5[2]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n556_6(.douta(w_n556_6[0]),.doutb(w_n556_6[1]),.doutc(w_n556_6[2]),.din(w_n556_1[2]));
	jspl3 jspl3_w_n556_7(.douta(w_n556_7[0]),.doutb(w_n556_7[1]),.doutc(w_n556_7[2]),.din(w_n556_2[0]));
	jspl jspl_w_n556_8(.douta(w_n556_8[0]),.doutb(w_n556_8[1]),.din(w_n556_2[1]));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_n559_0[1]),.din(n559));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n561_1(.douta(w_n561_1[0]),.doutb(w_n561_1[1]),.din(w_n561_0[0]));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_n564_0[1]),.din(n564));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.din(n569));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.doutc(w_n578_0[2]),.din(n578));
	jspl jspl_w_n578_1(.douta(w_n578_1[0]),.doutb(w_n578_1[1]),.din(w_n578_0[0]));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.doutc(w_n579_0[2]),.din(n579));
	jspl jspl_w_n579_1(.douta(w_n579_1[0]),.doutb(w_n579_1[1]),.din(w_n579_0[0]));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n586_1(.douta(w_n586_1[0]),.doutb(w_n586_1[1]),.din(w_n586_0[0]));
	jspl jspl_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.din(n587));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.doutc(w_n591_0[2]),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.doutc(w_n592_0[2]),.din(n592));
	jspl3 jspl3_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl jspl_w_n596_1(.douta(w_n596_1[0]),.doutb(w_n596_1[1]),.din(w_n596_0[0]));
	jspl3 jspl3_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.doutc(w_n597_0[2]),.din(n597));
	jspl3 jspl3_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.doutc(w_n601_0[2]),.din(n601));
	jspl jspl_w_n601_1(.douta(w_n601_1[0]),.doutb(w_n601_1[1]),.din(w_n601_0[0]));
	jspl3 jspl3_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.doutc(w_n602_0[2]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n607_1(.douta(w_n607_1[0]),.doutb(w_n607_1[1]),.din(w_n607_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.doutc(w_n608_0[2]),.din(n608));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n611_0(.douta(w_n611_0[0]),.doutb(w_n611_0[1]),.doutc(w_n611_0[2]),.din(n611));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.doutc(w_n613_1[2]),.din(w_n613_0[0]));
	jspl3 jspl3_w_n613_2(.douta(w_n613_2[0]),.doutb(w_n613_2[1]),.doutc(w_n613_2[2]),.din(w_n613_0[1]));
	jspl3 jspl3_w_n613_3(.douta(w_n613_3[0]),.doutb(w_n613_3[1]),.doutc(w_n613_3[2]),.din(w_n613_0[2]));
	jspl3 jspl3_w_n613_4(.douta(w_n613_4[0]),.doutb(w_n613_4[1]),.doutc(w_n613_4[2]),.din(w_n613_1[0]));
	jspl3 jspl3_w_n613_5(.douta(w_n613_5[0]),.doutb(w_n613_5[1]),.doutc(w_n613_5[2]),.din(w_n613_1[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n619_1(.douta(w_n619_1[0]),.doutb(w_n619_1[1]),.doutc(w_n619_1[2]),.din(w_n619_0[0]));
	jspl3 jspl3_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.doutc(w_n620_0[2]),.din(n620));
	jspl jspl_w_n620_1(.douta(w_n620_1[0]),.doutb(w_n620_1[1]),.din(w_n620_0[0]));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.din(n621));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_dff_A_OHwws77V4_0),.doutb(w_dff_A_f4Qd0c5u7_1),.doutc(w_n624_0[2]),.din(w_dff_B_Pns1XHaU6_3));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.din(n625));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl jspl_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.doutc(w_n628_0[2]),.din(n628));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n635_1(.douta(w_n635_1[0]),.doutb(w_n635_1[1]),.din(w_n635_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.doutc(w_n637_0[2]),.din(n637));
	jspl jspl_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.din(n638));
	jspl3 jspl3_w_n639_0(.douta(w_dff_A_lgyLa82g0_0),.doutb(w_n639_0[1]),.doutc(w_n639_0[2]),.din(n639));
	jspl jspl_w_n640_0(.douta(w_dff_A_QIqXiJiq1_0),.doutb(w_n640_0[1]),.din(n640));
	jspl3 jspl3_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.doutc(w_dff_A_AB6PTBb39_2),.din(n641));
	jspl3 jspl3_w_n641_1(.douta(w_n641_1[0]),.doutb(w_n641_1[1]),.doutc(w_n641_1[2]),.din(w_n641_0[0]));
	jspl3 jspl3_w_n644_0(.douta(w_dff_A_PyNPhz278_0),.doutb(w_n644_0[1]),.doutc(w_dff_A_uLWTeDtJ1_2),.din(n644));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.doutc(w_n648_0[2]),.din(n648));
	jspl jspl_w_n648_1(.douta(w_n648_1[0]),.doutb(w_n648_1[1]),.din(w_n648_0[0]));
	jspl jspl_w_n649_0(.douta(w_dff_A_To32fPpX3_0),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n653_0(.douta(w_n653_0[0]),.doutb(w_n653_0[1]),.doutc(w_n653_0[2]),.din(n653));
	jspl3 jspl3_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.doutc(w_n654_0[2]),.din(n654));
	jspl3 jspl3_w_n654_1(.douta(w_n654_1[0]),.doutb(w_n654_1[1]),.doutc(w_n654_1[2]),.din(w_n654_0[0]));
	jspl3 jspl3_w_n654_2(.douta(w_n654_2[0]),.doutb(w_n654_2[1]),.doutc(w_n654_2[2]),.din(w_n654_0[1]));
	jspl3 jspl3_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.doutc(w_n658_0[2]),.din(n658));
	jspl jspl_w_n658_1(.douta(w_n658_1[0]),.doutb(w_n658_1[1]),.din(w_n658_0[0]));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_n660_0[2]),.din(n660));
	jspl jspl_w_n660_1(.douta(w_dff_A_I23wfQs24_0),.doutb(w_n660_1[1]),.din(w_n660_0[0]));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(w_dff_B_yxUZZkK22_2));
	jspl jspl_w_n670_0(.douta(w_n670_0[0]),.doutb(w_n670_0[1]),.din(n670));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl3 jspl3_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.doutc(w_n682_0[2]),.din(n682));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.din(n692));
	jspl3 jspl3_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.doutc(w_n694_0[2]),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.doutc(w_n695_0[2]),.din(n695));
	jspl3 jspl3_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.doutc(w_n699_0[2]),.din(n699));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(n709));
	jspl jspl_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl3 jspl3_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.doutc(w_n713_0[2]),.din(n713));
	jspl3 jspl3_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.doutc(w_n715_0[2]),.din(n715));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(w_dff_B_LnBv0cEL0_2));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(n719));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(n721));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl3 jspl3_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.doutc(w_n725_0[2]),.din(n725));
	jspl jspl_w_n726_0(.douta(w_dff_A_uvSGRqJ13_0),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.doutc(w_n733_0[2]),.din(n733));
	jspl3 jspl3_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.doutc(w_n735_0[2]),.din(n735));
	jspl3 jspl3_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl jspl_w_n737_1(.douta(w_n737_1[0]),.doutb(w_n737_1[1]),.din(w_n737_0[0]));
	jspl jspl_w_n738_0(.douta(w_n738_0[0]),.doutb(w_n738_0[1]),.din(n738));
	jspl3 jspl3_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.doutc(w_n742_0[2]),.din(n742));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.doutc(w_n746_0[2]),.din(n746));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(w_dff_B_dL1fOSbo0_2));
	jspl3 jspl3_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.doutc(w_n749_0[2]),.din(n749));
	jspl3 jspl3_w_n749_1(.douta(w_n749_1[0]),.doutb(w_n749_1[1]),.doutc(w_n749_1[2]),.din(w_n749_0[0]));
	jspl3 jspl3_w_n749_2(.douta(w_n749_2[0]),.doutb(w_n749_2[1]),.doutc(w_n749_2[2]),.din(w_n749_0[1]));
	jspl3 jspl3_w_n749_3(.douta(w_n749_3[0]),.doutb(w_n749_3[1]),.doutc(w_n749_3[2]),.din(w_n749_0[2]));
	jspl3 jspl3_w_n749_4(.douta(w_n749_4[0]),.doutb(w_n749_4[1]),.doutc(w_n749_4[2]),.din(w_n749_1[0]));
	jspl3 jspl3_w_n749_5(.douta(w_n749_5[0]),.doutb(w_n749_5[1]),.doutc(w_n749_5[2]),.din(w_n749_1[1]));
	jspl3 jspl3_w_n749_6(.douta(w_n749_6[0]),.doutb(w_n749_6[1]),.doutc(w_n749_6[2]),.din(w_n749_1[2]));
	jspl3 jspl3_w_n749_7(.douta(w_n749_7[0]),.doutb(w_n749_7[1]),.doutc(w_n749_7[2]),.din(w_n749_2[0]));
	jspl3 jspl3_w_n749_8(.douta(w_n749_8[0]),.doutb(w_n749_8[1]),.doutc(w_n749_8[2]),.din(w_n749_2[1]));
	jspl3 jspl3_w_n749_9(.douta(w_n749_9[0]),.doutb(w_n749_9[1]),.doutc(w_n749_9[2]),.din(w_n749_2[2]));
	jspl3 jspl3_w_n749_10(.douta(w_n749_10[0]),.doutb(w_n749_10[1]),.doutc(w_n749_10[2]),.din(w_n749_3[0]));
	jspl3 jspl3_w_n749_11(.douta(w_n749_11[0]),.doutb(w_n749_11[1]),.doutc(w_n749_11[2]),.din(w_n749_3[1]));
	jspl3 jspl3_w_n749_12(.douta(w_n749_12[0]),.doutb(w_n749_12[1]),.doutc(w_n749_12[2]),.din(w_n749_3[2]));
	jspl jspl_w_n749_13(.douta(w_n749_13[0]),.doutb(w_n749_13[1]),.din(w_n749_4[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.doutc(w_n750_0[2]),.din(n750));
	jspl3 jspl3_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.doutc(w_n750_1[2]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n750_2(.douta(w_n750_2[0]),.doutb(w_n750_2[1]),.doutc(w_n750_2[2]),.din(w_n750_0[1]));
	jspl3 jspl3_w_n750_3(.douta(w_n750_3[0]),.doutb(w_n750_3[1]),.doutc(w_n750_3[2]),.din(w_n750_0[2]));
	jspl3 jspl3_w_n750_4(.douta(w_n750_4[0]),.doutb(w_n750_4[1]),.doutc(w_n750_4[2]),.din(w_n750_1[0]));
	jspl3 jspl3_w_n750_5(.douta(w_n750_5[0]),.doutb(w_n750_5[1]),.doutc(w_n750_5[2]),.din(w_n750_1[1]));
	jspl3 jspl3_w_n750_6(.douta(w_n750_6[0]),.doutb(w_n750_6[1]),.doutc(w_n750_6[2]),.din(w_n750_1[2]));
	jspl3 jspl3_w_n750_7(.douta(w_n750_7[0]),.doutb(w_n750_7[1]),.doutc(w_n750_7[2]),.din(w_n750_2[0]));
	jspl3 jspl3_w_n750_8(.douta(w_n750_8[0]),.doutb(w_n750_8[1]),.doutc(w_n750_8[2]),.din(w_n750_2[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.doutc(w_n753_0[2]),.din(n753));
	jspl jspl_w_n753_1(.douta(w_n753_1[0]),.doutb(w_n753_1[1]),.din(w_n753_0[0]));
	jspl jspl_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.din(n755));
	jspl3 jspl3_w_n763_0(.douta(w_n763_0[0]),.doutb(w_n763_0[1]),.doutc(w_n763_0[2]),.din(n763));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.din(n779));
	jspl3 jspl3_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.doutc(w_n786_0[2]),.din(n786));
	jspl3 jspl3_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.doutc(w_n788_0[2]),.din(n788));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_dff_A_YMMn1aJu8_1),.doutc(w_n790_0[2]),.din(n790));
	jspl3 jspl3_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.doutc(w_dff_A_zmpyFrKI5_2),.din(n792));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_n797_1[1]),.doutc(w_n797_1[2]),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_n797_2[2]),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_n797_3[0]),.doutb(w_n797_3[1]),.doutc(w_n797_3[2]),.din(w_n797_0[2]));
	jspl3 jspl3_w_n797_4(.douta(w_n797_4[0]),.doutb(w_n797_4[1]),.doutc(w_n797_4[2]),.din(w_n797_1[0]));
	jspl3 jspl3_w_n797_5(.douta(w_n797_5[0]),.doutb(w_n797_5[1]),.doutc(w_n797_5[2]),.din(w_n797_1[1]));
	jspl3 jspl3_w_n797_6(.douta(w_n797_6[0]),.doutb(w_n797_6[1]),.doutc(w_n797_6[2]),.din(w_n797_1[2]));
	jspl3 jspl3_w_n797_7(.douta(w_n797_7[0]),.doutb(w_n797_7[1]),.doutc(w_n797_7[2]),.din(w_n797_2[0]));
	jspl3 jspl3_w_n797_8(.douta(w_n797_8[0]),.doutb(w_n797_8[1]),.doutc(w_n797_8[2]),.din(w_n797_2[1]));
	jspl jspl_w_n797_9(.douta(w_n797_9[0]),.doutb(w_n797_9[1]),.din(w_n797_2[2]));
	jspl3 jspl3_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.doutc(w_n798_0[2]),.din(n798));
	jspl jspl_w_n798_1(.douta(w_n798_1[0]),.doutb(w_n798_1[1]),.din(w_n798_0[0]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.doutc(w_n800_0[2]),.din(n800));
	jspl3 jspl3_w_n800_1(.douta(w_n800_1[0]),.doutb(w_dff_A_rW7yqhoM0_1),.doutc(w_dff_A_fW8OGSka8_2),.din(w_n800_0[0]));
	jspl3 jspl3_w_n800_2(.douta(w_n800_2[0]),.doutb(w_n800_2[1]),.doutc(w_n800_2[2]),.din(w_n800_0[1]));
	jspl3 jspl3_w_n800_3(.douta(w_dff_A_OzL5O6s65_0),.doutb(w_n800_3[1]),.doutc(w_dff_A_AHqMAjRY7_2),.din(w_n800_0[2]));
	jspl jspl_w_n800_4(.douta(w_dff_A_i5zeMe8m5_0),.doutb(w_n800_4[1]),.din(w_n800_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl jspl_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n814_0(.douta(w_dff_A_AL4TBzB66_0),.doutb(w_dff_A_EEJ6wBEC7_1),.doutc(w_n814_0[2]),.din(n814));
	jspl3 jspl3_w_n819_0(.douta(w_n819_0[0]),.doutb(w_dff_A_eUZQ0gCo5_1),.doutc(w_n819_0[2]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_dff_A_NA9Df6H68_1),.din(n821));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n836_0(.douta(w_dff_A_bKVOydk43_0),.doutb(w_n836_0[1]),.din(n836));
	jspl jspl_w_n847_0(.douta(w_dff_A_QOxkxB1I3_0),.doutb(w_n847_0[1]),.din(n847));
	jspl3 jspl3_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.doutc(w_n852_0[2]),.din(n852));
	jspl3 jspl3_w_n852_1(.douta(w_n852_1[0]),.doutb(w_n852_1[1]),.doutc(w_n852_1[2]),.din(w_n852_0[0]));
	jspl3 jspl3_w_n852_2(.douta(w_n852_2[0]),.doutb(w_n852_2[1]),.doutc(w_n852_2[2]),.din(w_n852_0[1]));
	jspl3 jspl3_w_n852_3(.douta(w_n852_3[0]),.doutb(w_n852_3[1]),.doutc(w_n852_3[2]),.din(w_n852_0[2]));
	jspl3 jspl3_w_n852_4(.douta(w_n852_4[0]),.doutb(w_n852_4[1]),.doutc(w_n852_4[2]),.din(w_n852_1[0]));
	jspl3 jspl3_w_n852_5(.douta(w_n852_5[0]),.doutb(w_n852_5[1]),.doutc(w_n852_5[2]),.din(w_n852_1[1]));
	jspl3 jspl3_w_n852_6(.douta(w_n852_6[0]),.doutb(w_n852_6[1]),.doutc(w_n852_6[2]),.din(w_n852_1[2]));
	jspl3 jspl3_w_n852_7(.douta(w_n852_7[0]),.doutb(w_n852_7[1]),.doutc(w_n852_7[2]),.din(w_n852_2[0]));
	jspl3 jspl3_w_n852_8(.douta(w_n852_8[0]),.doutb(w_n852_8[1]),.doutc(w_n852_8[2]),.din(w_n852_2[1]));
	jspl jspl_w_n852_9(.douta(w_n852_9[0]),.doutb(w_n852_9[1]),.din(w_n852_2[2]));
	jspl3 jspl3_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.doutc(w_n854_0[2]),.din(n854));
	jspl3 jspl3_w_n854_1(.douta(w_n854_1[0]),.doutb(w_dff_A_E2vII9n89_1),.doutc(w_dff_A_w3eUXdrG5_2),.din(w_n854_0[0]));
	jspl3 jspl3_w_n854_2(.douta(w_n854_2[0]),.doutb(w_n854_2[1]),.doutc(w_n854_2[2]),.din(w_n854_0[1]));
	jspl3 jspl3_w_n854_3(.douta(w_n854_3[0]),.doutb(w_n854_3[1]),.doutc(w_dff_A_P2s8uA8u4_2),.din(w_n854_0[2]));
	jspl jspl_w_n854_4(.douta(w_dff_A_EjKLw5jY3_0),.doutb(w_n854_4[1]),.din(w_n854_1[0]));
	jspl3 jspl3_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.doutc(w_n865_0[2]),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n868_0(.douta(w_n868_0[0]),.doutb(w_n868_0[1]),.din(n868));
	jspl jspl_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.din(n870));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl jspl_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.din(n880));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(n890));
	jspl jspl_w_n901_0(.douta(w_n901_0[0]),.doutb(w_n901_0[1]),.din(n901));
	jspl3 jspl3_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.doutc(w_n923_0[2]),.din(n923));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl3 jspl3_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.doutc(w_n938_0[2]),.din(n938));
	jspl3 jspl3_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.doutc(w_n940_0[2]),.din(n940));
	jspl jspl_w_n940_1(.douta(w_n940_1[0]),.doutb(w_n940_1[1]),.din(w_n940_0[0]));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(n944));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(n949));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl3 jspl3_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.doutc(w_n954_0[2]),.din(n954));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl3 jspl3_w_n977_0(.douta(w_n977_0[0]),.doutb(w_n977_0[1]),.doutc(w_n977_0[2]),.din(n977));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_dff_A_WnRpMoNw1_1),.din(n989));
	jspl3 jspl3_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.doutc(w_n993_0[2]),.din(n993));
	jspl3 jspl3_w_n993_1(.douta(w_n993_1[0]),.doutb(w_n993_1[1]),.doutc(w_n993_1[2]),.din(w_n993_0[0]));
	jspl3 jspl3_w_n993_2(.douta(w_n993_2[0]),.doutb(w_n993_2[1]),.doutc(w_n993_2[2]),.din(w_n993_0[1]));
	jspl3 jspl3_w_n993_3(.douta(w_dff_A_F2Q6BTQG0_0),.doutb(w_dff_A_fhl7roYl2_1),.doutc(w_n993_3[2]),.din(w_n993_0[2]));
	jspl3 jspl3_w_n993_4(.douta(w_n993_4[0]),.doutb(w_n993_4[1]),.doutc(w_n993_4[2]),.din(w_n993_1[0]));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n994_1(.douta(w_n994_1[0]),.doutb(w_n994_1[1]),.doutc(w_n994_1[2]),.din(w_n994_0[0]));
	jspl3 jspl3_w_n994_2(.douta(w_n994_2[0]),.doutb(w_n994_2[1]),.doutc(w_n994_2[2]),.din(w_n994_0[1]));
	jspl3 jspl3_w_n994_3(.douta(w_n994_3[0]),.doutb(w_n994_3[1]),.doutc(w_n994_3[2]),.din(w_n994_0[2]));
	jspl jspl_w_n994_4(.douta(w_n994_4[0]),.doutb(w_n994_4[1]),.din(w_n994_1[0]));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl3 jspl3_w_n996_1(.douta(w_n996_1[0]),.doutb(w_n996_1[1]),.doutc(w_n996_1[2]),.din(w_n996_0[0]));
	jspl3 jspl3_w_n996_2(.douta(w_n996_2[0]),.doutb(w_n996_2[1]),.doutc(w_n996_2[2]),.din(w_n996_0[1]));
	jspl3 jspl3_w_n996_3(.douta(w_n996_3[0]),.doutb(w_n996_3[1]),.doutc(w_n996_3[2]),.din(w_n996_0[2]));
	jspl jspl_w_n996_4(.douta(w_n996_4[0]),.doutb(w_n996_4[1]),.din(w_n996_1[0]));
	jspl3 jspl3_w_n999_0(.douta(w_dff_A_MuefKJ1V5_0),.doutb(w_dff_A_MgODUluG2_1),.doutc(w_n999_0[2]),.din(w_dff_B_mVgp88tn7_3));
	jspl3 jspl3_w_n999_1(.douta(w_dff_A_THe3ti0z9_0),.doutb(w_dff_A_pZ4xnjMO7_1),.doutc(w_n999_1[2]),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_dff_A_ivUFOrEV2_0),.doutb(w_dff_A_NTmV4l3H9_1),.doutc(w_n999_2[2]),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_dff_A_MwSGsGmt7_0),.doutb(w_dff_A_ZHlsjuj38_1),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl3 jspl3_w_n1007_0(.douta(w_dff_A_X5ele9mj2_0),.doutb(w_dff_A_nRJ4LMDu5_1),.doutc(w_n1007_0[2]),.din(w_dff_B_ilgOphnQ3_3));
	jspl3 jspl3_w_n1007_1(.douta(w_n1007_1[0]),.doutb(w_n1007_1[1]),.doutc(w_dff_A_o4xpqt266_2),.din(w_n1007_0[0]));
	jspl3 jspl3_w_n1007_2(.douta(w_dff_A_dgPqd10H5_0),.doutb(w_dff_A_LTUJUBnO9_1),.doutc(w_n1007_2[2]),.din(w_n1007_0[1]));
	jspl3 jspl3_w_n1007_3(.douta(w_dff_A_PIcgelcc1_0),.doutb(w_dff_A_9gFfPl351_1),.doutc(w_n1007_3[2]),.din(w_n1007_0[2]));
	jspl3 jspl3_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.doutc(w_n1008_0[2]),.din(n1008));
	jspl3 jspl3_w_n1008_1(.douta(w_n1008_1[0]),.doutb(w_n1008_1[1]),.doutc(w_n1008_1[2]),.din(w_n1008_0[0]));
	jspl3 jspl3_w_n1008_2(.douta(w_n1008_2[0]),.doutb(w_n1008_2[1]),.doutc(w_n1008_2[2]),.din(w_n1008_0[1]));
	jspl3 jspl3_w_n1008_3(.douta(w_dff_A_PHmYnQ426_0),.doutb(w_dff_A_CNn93fsX2_1),.doutc(w_n1008_3[2]),.din(w_n1008_0[2]));
	jspl3 jspl3_w_n1008_4(.douta(w_n1008_4[0]),.doutb(w_n1008_4[1]),.doutc(w_n1008_4[2]),.din(w_n1008_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl3 jspl3_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.doutc(w_n1012_1[2]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1012_2(.douta(w_n1012_2[0]),.doutb(w_n1012_2[1]),.doutc(w_n1012_2[2]),.din(w_n1012_0[1]));
	jspl3 jspl3_w_n1012_3(.douta(w_n1012_3[0]),.doutb(w_n1012_3[1]),.doutc(w_n1012_3[2]),.din(w_n1012_0[2]));
	jspl jspl_w_n1012_4(.douta(w_n1012_4[0]),.doutb(w_n1012_4[1]),.din(w_n1012_1[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl3 jspl3_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.doutc(w_n1014_1[2]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1014_2(.douta(w_n1014_2[0]),.doutb(w_n1014_2[1]),.doutc(w_n1014_2[2]),.din(w_n1014_0[1]));
	jspl3 jspl3_w_n1014_3(.douta(w_n1014_3[0]),.doutb(w_n1014_3[1]),.doutc(w_n1014_3[2]),.din(w_n1014_0[2]));
	jspl jspl_w_n1014_4(.douta(w_n1014_4[0]),.doutb(w_n1014_4[1]),.din(w_n1014_1[0]));
	jspl3 jspl3_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.doutc(w_n1019_0[2]),.din(n1019));
	jspl jspl_w_n1019_1(.douta(w_n1019_1[0]),.doutb(w_n1019_1[1]),.din(w_n1019_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl3 jspl3_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.doutc(w_n1043_0[2]),.din(n1043));
	jspl jspl_w_n1043_1(.douta(w_n1043_1[0]),.doutb(w_n1043_1[1]),.din(w_n1043_0[0]));
	jspl3 jspl3_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.doutc(w_n1052_0[2]),.din(n1052));
	jspl jspl_w_n1052_1(.douta(w_n1052_1[0]),.doutb(w_n1052_1[1]),.din(w_n1052_0[0]));
	jspl3 jspl3_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.doutc(w_n1054_0[2]),.din(n1054));
	jspl jspl_w_n1054_1(.douta(w_n1054_1[0]),.doutb(w_n1054_1[1]),.din(w_n1054_0[0]));
	jspl jspl_w_n1177_0(.douta(w_dff_A_jcFJtrsX8_0),.doutb(w_n1177_0[1]),.din(w_dff_B_xmNcrysp8_2));
	jspl jspl_w_n1179_0(.douta(w_dff_A_cinRNd2W2_0),.doutb(w_n1179_0[1]),.din(n1179));
	jspl3 jspl3_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.doutc(w_n1196_0[2]),.din(n1196));
	jspl3 jspl3_w_n1196_1(.douta(w_n1196_1[0]),.doutb(w_n1196_1[1]),.doutc(w_n1196_1[2]),.din(w_n1196_0[0]));
	jspl3 jspl3_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.doutc(w_n1201_0[2]),.din(n1201));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.doutc(w_n1213_0[2]),.din(n1213));
	jspl3 jspl3_w_n1213_1(.douta(w_n1213_1[0]),.doutb(w_n1213_1[1]),.doutc(w_n1213_1[2]),.din(w_n1213_0[0]));
	jspl3 jspl3_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.doutc(w_n1236_0[2]),.din(n1236));
	jspl3 jspl3_w_n1236_1(.douta(w_n1236_1[0]),.doutb(w_n1236_1[1]),.doutc(w_n1236_1[2]),.din(w_n1236_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl3 jspl3_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.doutc(w_n1251_1[2]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.doutc(w_n1279_0[2]),.din(n1279));
	jspl jspl_w_n1279_1(.douta(w_n1279_1[0]),.doutb(w_n1279_1[1]),.din(w_n1279_0[0]));
	jspl3 jspl3_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.doutc(w_n1297_0[2]),.din(n1297));
	jspl jspl_w_n1297_1(.douta(w_n1297_1[0]),.doutb(w_n1297_1[1]),.din(w_n1297_0[0]));
	jspl3 jspl3_w_n1299_0(.douta(w_n1299_0[0]),.doutb(w_n1299_0[1]),.doutc(w_n1299_0[2]),.din(n1299));
	jspl jspl_w_n1299_1(.douta(w_n1299_1[0]),.doutb(w_n1299_1[1]),.din(w_n1299_0[0]));
	jspl3 jspl3_w_n1410_0(.douta(w_dff_A_TL0ht9Jp2_0),.doutb(w_n1410_0[1]),.doutc(w_n1410_0[2]),.din(n1410));
	jspl3 jspl3_w_n1412_0(.douta(w_n1412_0[0]),.doutb(w_dff_A_Zmmqp0qp7_1),.doutc(w_dff_A_0XMBlSB18_2),.din(w_dff_B_9csyNqWX5_3));
	jspl jspl_w_n1416_0(.douta(w_n1416_0[0]),.doutb(w_n1416_0[1]),.din(n1416));
	jspl jspl_w_n1422_0(.douta(w_dff_A_XjBaWqj13_0),.doutb(w_n1422_0[1]),.din(n1422));
	jspl jspl_w_n1425_0(.douta(w_dff_A_77FCiIJy7_0),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(n1428));
	jspl jspl_w_n1429_0(.douta(w_dff_A_cssLASeX9_0),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1451_0(.douta(w_dff_A_7wxXQokn0_0),.doutb(w_n1451_0[1]),.din(n1451));
	jspl jspl_w_n1503_0(.douta(w_n1503_0[0]),.doutb(w_n1503_0[1]),.din(n1503));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1592_0(.douta(w_n1592_0[0]),.doutb(w_n1592_0[1]),.din(n1592));
	jspl jspl_w_n1593_0(.douta(w_n1593_0[0]),.doutb(w_n1593_0[1]),.din(n1593));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_n1603_0[1]),.din(n1603));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl3 jspl3_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.doutc(w_n1611_0[2]),.din(n1611));
	jspl jspl_w_n1613_0(.douta(w_n1613_0[0]),.doutb(w_n1613_0[1]),.din(n1613));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(n1615));
	jspl jspl_w_n1618_0(.douta(w_n1618_0[0]),.doutb(w_n1618_0[1]),.din(n1618));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(n1633));
	jspl jspl_w_n1637_0(.douta(w_n1637_0[0]),.doutb(w_n1637_0[1]),.din(n1637));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(n1643));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_n1652_0[1]),.din(n1652));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl3 jspl3_w_n1674_0(.douta(w_n1674_0[0]),.doutb(w_n1674_0[1]),.doutc(w_n1674_0[2]),.din(n1674));
	jspl jspl_w_n1675_0(.douta(w_n1675_0[0]),.doutb(w_n1675_0[1]),.din(n1675));
	jspl3 jspl3_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.doutc(w_n1679_0[2]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(w_dff_B_N8xjebfb1_2));
	jspl jspl_w_n1695_0(.douta(w_n1695_0[0]),.doutb(w_n1695_0[1]),.din(n1695));
	jspl jspl_w_n1698_0(.douta(w_n1698_0[0]),.doutb(w_n1698_0[1]),.din(n1698));
	jdff dff_B_1XDqtN614_1(.din(G136),.dout(w_dff_B_1XDqtN614_1),.clk(gclk));
	jdff dff_B_NWXNKUrM1_0(.din(G2824),.dout(w_dff_B_NWXNKUrM1_0),.clk(gclk));
	jdff dff_B_DGe8f2Ly5_1(.din(n320),.dout(w_dff_B_DGe8f2Ly5_1),.clk(gclk));
	jdff dff_B_02uGgqTc3_1(.din(n327),.dout(w_dff_B_02uGgqTc3_1),.clk(gclk));
	jdff dff_B_8mCnqYH29_2(.din(n333),.dout(w_dff_B_8mCnqYH29_2),.clk(gclk));
	jdff dff_B_WU1X1XVA1_1(.din(n338),.dout(w_dff_B_WU1X1XVA1_1),.clk(gclk));
	jdff dff_B_cWl4mArx2_1(.din(n340),.dout(w_dff_B_cWl4mArx2_1),.clk(gclk));
	jdff dff_B_ymTIAQl32_0(.din(n341),.dout(w_dff_B_ymTIAQl32_0),.clk(gclk));
	jdff dff_B_evs6UKxu5_1(.din(n345),.dout(w_dff_B_evs6UKxu5_1),.clk(gclk));
	jdff dff_B_4hxtTxcj6_0(.din(n346),.dout(w_dff_B_4hxtTxcj6_0),.clk(gclk));
	jdff dff_A_aTDcNNYc3_0(.dout(w_G141_2[0]),.din(w_dff_A_aTDcNNYc3_0),.clk(gclk));
	jdff dff_A_6TXUEXf09_0(.dout(w_dff_A_aTDcNNYc3_0),.din(w_dff_A_6TXUEXf09_0),.clk(gclk));
	jdff dff_A_UMdNmIRg8_0(.dout(w_dff_A_6TXUEXf09_0),.din(w_dff_A_UMdNmIRg8_0),.clk(gclk));
	jdff dff_A_NY7cL5aH0_0(.dout(w_dff_A_UMdNmIRg8_0),.din(w_dff_A_NY7cL5aH0_0),.clk(gclk));
	jdff dff_A_CTZAlmyf1_1(.dout(w_G141_2[1]),.din(w_dff_A_CTZAlmyf1_1),.clk(gclk));
	jdff dff_A_VNgfi1wZ6_1(.dout(w_dff_A_CTZAlmyf1_1),.din(w_dff_A_VNgfi1wZ6_1),.clk(gclk));
	jdff dff_A_5VzWEKJm9_1(.dout(w_dff_A_VNgfi1wZ6_1),.din(w_dff_A_5VzWEKJm9_1),.clk(gclk));
	jdff dff_A_nCk6XHLC6_1(.dout(w_dff_A_5VzWEKJm9_1),.din(w_dff_A_nCk6XHLC6_1),.clk(gclk));
	jdff dff_B_uVFbPRHM4_1(.din(n350),.dout(w_dff_B_uVFbPRHM4_1),.clk(gclk));
	jdff dff_B_ct9crCYT1_0(.din(n351),.dout(w_dff_B_ct9crCYT1_0),.clk(gclk));
	jdff dff_B_t7LjX50Y3_1(.din(n355),.dout(w_dff_B_t7LjX50Y3_1),.clk(gclk));
	jdff dff_B_YVG9Lfyh4_1(.din(w_dff_B_t7LjX50Y3_1),.dout(w_dff_B_YVG9Lfyh4_1),.clk(gclk));
	jdff dff_A_QYFEgyJ75_1(.dout(w_G141_1[1]),.din(w_dff_A_QYFEgyJ75_1),.clk(gclk));
	jdff dff_A_rtIH0M167_1(.dout(w_dff_A_QYFEgyJ75_1),.din(w_dff_A_rtIH0M167_1),.clk(gclk));
	jdff dff_A_3YClfHk96_1(.dout(w_dff_A_rtIH0M167_1),.din(w_dff_A_3YClfHk96_1),.clk(gclk));
	jdff dff_A_Z7jBtOZN9_1(.dout(w_dff_A_3YClfHk96_1),.din(w_dff_A_Z7jBtOZN9_1),.clk(gclk));
	jdff dff_A_E051C3Hs2_2(.dout(w_G141_1[2]),.din(w_dff_A_E051C3Hs2_2),.clk(gclk));
	jdff dff_A_P9uuXgGt3_2(.dout(w_dff_A_E051C3Hs2_2),.din(w_dff_A_P9uuXgGt3_2),.clk(gclk));
	jdff dff_A_jqXwJ04v1_2(.dout(w_dff_A_P9uuXgGt3_2),.din(w_dff_A_jqXwJ04v1_2),.clk(gclk));
	jdff dff_A_NDNz4G301_2(.dout(w_dff_A_jqXwJ04v1_2),.din(w_dff_A_NDNz4G301_2),.clk(gclk));
	jdff dff_B_QLc7tfjg4_2(.din(n661),.dout(w_dff_B_QLc7tfjg4_2),.clk(gclk));
	jdff dff_B_yxUZZkK22_2(.din(w_dff_B_QLc7tfjg4_2),.dout(w_dff_B_yxUZZkK22_2),.clk(gclk));
	jdff dff_B_ejixAcWz8_2(.din(n717),.dout(w_dff_B_ejixAcWz8_2),.clk(gclk));
	jdff dff_B_LnBv0cEL0_2(.din(w_dff_B_ejixAcWz8_2),.dout(w_dff_B_LnBv0cEL0_2),.clk(gclk));
	jdff dff_B_ZpYFQVyI0_2(.din(n747),.dout(w_dff_B_ZpYFQVyI0_2),.clk(gclk));
	jdff dff_B_dL1fOSbo0_2(.din(w_dff_B_ZpYFQVyI0_2),.dout(w_dff_B_dL1fOSbo0_2),.clk(gclk));
	jdff dff_B_42FdxOi56_1(.din(n739),.dout(w_dff_B_42FdxOi56_1),.clk(gclk));
	jdff dff_B_nYAXIFgQ6_1(.din(w_dff_B_42FdxOi56_1),.dout(w_dff_B_nYAXIFgQ6_1),.clk(gclk));
	jdff dff_A_wuoPVNGL9_0(.dout(w_n660_1[0]),.din(w_dff_A_wuoPVNGL9_0),.clk(gclk));
	jdff dff_A_1WsWmMIa4_0(.dout(w_dff_A_wuoPVNGL9_0),.din(w_dff_A_1WsWmMIa4_0),.clk(gclk));
	jdff dff_A_Q3QhfmJ97_0(.dout(w_dff_A_1WsWmMIa4_0),.din(w_dff_A_Q3QhfmJ97_0),.clk(gclk));
	jdff dff_A_N2EbYwlV9_0(.dout(w_dff_A_Q3QhfmJ97_0),.din(w_dff_A_N2EbYwlV9_0),.clk(gclk));
	jdff dff_A_I23wfQs24_0(.dout(w_dff_A_N2EbYwlV9_0),.din(w_dff_A_I23wfQs24_0),.clk(gclk));
	jdff dff_B_SrbdkDKe1_0(.din(n808),.dout(w_dff_B_SrbdkDKe1_0),.clk(gclk));
	jdff dff_B_CLpfSep24_0(.din(w_dff_B_SrbdkDKe1_0),.dout(w_dff_B_CLpfSep24_0),.clk(gclk));
	jdff dff_B_VLthB9qI7_0(.din(w_dff_B_CLpfSep24_0),.dout(w_dff_B_VLthB9qI7_0),.clk(gclk));
	jdff dff_B_pXxDp6Gp4_0(.din(w_dff_B_VLthB9qI7_0),.dout(w_dff_B_pXxDp6Gp4_0),.clk(gclk));
	jdff dff_B_W0hYXjTc2_0(.din(w_dff_B_pXxDp6Gp4_0),.dout(w_dff_B_W0hYXjTc2_0),.clk(gclk));
	jdff dff_B_2gpE8J2N2_0(.din(w_dff_B_W0hYXjTc2_0),.dout(w_dff_B_2gpE8J2N2_0),.clk(gclk));
	jdff dff_B_vGuJ81Mt1_0(.din(w_dff_B_2gpE8J2N2_0),.dout(w_dff_B_vGuJ81Mt1_0),.clk(gclk));
	jdff dff_B_qGsbcCoP7_0(.din(w_dff_B_vGuJ81Mt1_0),.dout(w_dff_B_qGsbcCoP7_0),.clk(gclk));
	jdff dff_B_I3EXTdrl5_0(.din(w_dff_B_qGsbcCoP7_0),.dout(w_dff_B_I3EXTdrl5_0),.clk(gclk));
	jdff dff_B_sdoMaWUL3_0(.din(w_dff_B_I3EXTdrl5_0),.dout(w_dff_B_sdoMaWUL3_0),.clk(gclk));
	jdff dff_B_h0oYGuxO9_0(.din(n803),.dout(w_dff_B_h0oYGuxO9_0),.clk(gclk));
	jdff dff_B_PsD8Npqn0_0(.din(n861),.dout(w_dff_B_PsD8Npqn0_0),.clk(gclk));
	jdff dff_B_FCir2w6a8_0(.din(w_dff_B_PsD8Npqn0_0),.dout(w_dff_B_FCir2w6a8_0),.clk(gclk));
	jdff dff_B_Y5xQJbdQ2_0(.din(w_dff_B_FCir2w6a8_0),.dout(w_dff_B_Y5xQJbdQ2_0),.clk(gclk));
	jdff dff_B_UoJE27xX2_0(.din(w_dff_B_Y5xQJbdQ2_0),.dout(w_dff_B_UoJE27xX2_0),.clk(gclk));
	jdff dff_B_r7vsXoro3_0(.din(w_dff_B_UoJE27xX2_0),.dout(w_dff_B_r7vsXoro3_0),.clk(gclk));
	jdff dff_B_LDQicVIw5_0(.din(w_dff_B_r7vsXoro3_0),.dout(w_dff_B_LDQicVIw5_0),.clk(gclk));
	jdff dff_B_zZKmTWFN9_0(.din(w_dff_B_LDQicVIw5_0),.dout(w_dff_B_zZKmTWFN9_0),.clk(gclk));
	jdff dff_B_wHakUf6M9_0(.din(w_dff_B_zZKmTWFN9_0),.dout(w_dff_B_wHakUf6M9_0),.clk(gclk));
	jdff dff_B_hLiWu55m5_0(.din(w_dff_B_wHakUf6M9_0),.dout(w_dff_B_hLiWu55m5_0),.clk(gclk));
	jdff dff_B_VjAzt5NF2_0(.din(w_dff_B_hLiWu55m5_0),.dout(w_dff_B_VjAzt5NF2_0),.clk(gclk));
	jdff dff_B_2QD7IzGH6_0(.din(n856),.dout(w_dff_B_2QD7IzGH6_0),.clk(gclk));
	jdff dff_B_e9C2TA1l0_0(.din(n967),.dout(w_dff_B_e9C2TA1l0_0),.clk(gclk));
	jdff dff_B_pCqoakHu4_1(.din(n975),.dout(w_dff_B_pCqoakHu4_1),.clk(gclk));
	jdff dff_B_TFXHJJCi8_1(.din(w_dff_B_pCqoakHu4_1),.dout(w_dff_B_TFXHJJCi8_1),.clk(gclk));
	jdff dff_B_1f6Bj5Ek6_1(.din(w_dff_B_TFXHJJCi8_1),.dout(w_dff_B_1f6Bj5Ek6_1),.clk(gclk));
	jdff dff_B_xuXpjySI2_1(.din(w_dff_B_1f6Bj5Ek6_1),.dout(w_dff_B_xuXpjySI2_1),.clk(gclk));
	jdff dff_B_thoFfn6c7_1(.din(w_dff_B_xuXpjySI2_1),.dout(w_dff_B_thoFfn6c7_1),.clk(gclk));
	jdff dff_B_rNexfRzB6_1(.din(n971),.dout(w_dff_B_rNexfRzB6_1),.clk(gclk));
	jdff dff_B_7yMBzruG2_1(.din(w_dff_B_rNexfRzB6_1),.dout(w_dff_B_7yMBzruG2_1),.clk(gclk));
	jdff dff_B_wbZMDG4q2_1(.din(n995),.dout(w_dff_B_wbZMDG4q2_1),.clk(gclk));
	jdff dff_B_aBxZBdJR1_1(.din(w_dff_B_wbZMDG4q2_1),.dout(w_dff_B_aBxZBdJR1_1),.clk(gclk));
	jdff dff_B_pwN17cui4_1(.din(w_dff_B_aBxZBdJR1_1),.dout(w_dff_B_pwN17cui4_1),.clk(gclk));
	jdff dff_B_iITFd7oW1_1(.din(w_dff_B_pwN17cui4_1),.dout(w_dff_B_iITFd7oW1_1),.clk(gclk));
	jdff dff_B_REj9hCEs1_1(.din(w_dff_B_iITFd7oW1_1),.dout(w_dff_B_REj9hCEs1_1),.clk(gclk));
	jdff dff_B_2NVMryv08_1(.din(w_dff_B_REj9hCEs1_1),.dout(w_dff_B_2NVMryv08_1),.clk(gclk));
	jdff dff_B_1J9G3Uuu6_1(.din(w_dff_B_2NVMryv08_1),.dout(w_dff_B_1J9G3Uuu6_1),.clk(gclk));
	jdff dff_B_8tTiHC1z2_1(.din(w_dff_B_1J9G3Uuu6_1),.dout(w_dff_B_8tTiHC1z2_1),.clk(gclk));
	jdff dff_B_2mbvwedk1_1(.din(w_dff_B_8tTiHC1z2_1),.dout(w_dff_B_2mbvwedk1_1),.clk(gclk));
	jdff dff_B_8D4Cehdn5_1(.din(w_dff_B_2mbvwedk1_1),.dout(w_dff_B_8D4Cehdn5_1),.clk(gclk));
	jdff dff_B_MJIvSDTw3_1(.din(w_dff_B_8D4Cehdn5_1),.dout(w_dff_B_MJIvSDTw3_1),.clk(gclk));
	jdff dff_B_qQYNLmVd5_1(.din(n997),.dout(w_dff_B_qQYNLmVd5_1),.clk(gclk));
	jdff dff_B_LriefBrK7_1(.din(w_dff_B_qQYNLmVd5_1),.dout(w_dff_B_LriefBrK7_1),.clk(gclk));
	jdff dff_B_OAH3sFTR3_1(.din(w_dff_B_LriefBrK7_1),.dout(w_dff_B_OAH3sFTR3_1),.clk(gclk));
	jdff dff_B_PwyMtHtu2_1(.din(w_dff_B_OAH3sFTR3_1),.dout(w_dff_B_PwyMtHtu2_1),.clk(gclk));
	jdff dff_B_Kvi4Oh500_1(.din(w_dff_B_PwyMtHtu2_1),.dout(w_dff_B_Kvi4Oh500_1),.clk(gclk));
	jdff dff_B_L3pEp55h8_1(.din(w_dff_B_Kvi4Oh500_1),.dout(w_dff_B_L3pEp55h8_1),.clk(gclk));
	jdff dff_B_BvbV19yi7_1(.din(w_dff_B_L3pEp55h8_1),.dout(w_dff_B_BvbV19yi7_1),.clk(gclk));
	jdff dff_B_zOxoHVXV3_1(.din(w_dff_B_BvbV19yi7_1),.dout(w_dff_B_zOxoHVXV3_1),.clk(gclk));
	jdff dff_B_PqIQVwuk4_1(.din(w_dff_B_zOxoHVXV3_1),.dout(w_dff_B_PqIQVwuk4_1),.clk(gclk));
	jdff dff_B_siH4tvwf9_1(.din(w_dff_B_PqIQVwuk4_1),.dout(w_dff_B_siH4tvwf9_1),.clk(gclk));
	jdff dff_B_uHiqWlh60_1(.din(w_dff_B_siH4tvwf9_1),.dout(w_dff_B_uHiqWlh60_1),.clk(gclk));
	jdff dff_B_rMnhefMo1_0(.din(n1001),.dout(w_dff_B_rMnhefMo1_0),.clk(gclk));
	jdff dff_B_DIwzV3yi0_0(.din(n1016),.dout(w_dff_B_DIwzV3yi0_0),.clk(gclk));
	jdff dff_B_mzplZVB74_0(.din(w_dff_B_DIwzV3yi0_0),.dout(w_dff_B_mzplZVB74_0),.clk(gclk));
	jdff dff_B_P3URP6Jn0_0(.din(w_dff_B_mzplZVB74_0),.dout(w_dff_B_P3URP6Jn0_0),.clk(gclk));
	jdff dff_B_WejOFSqx6_0(.din(w_dff_B_P3URP6Jn0_0),.dout(w_dff_B_WejOFSqx6_0),.clk(gclk));
	jdff dff_B_Tah9espN4_0(.din(w_dff_B_WejOFSqx6_0),.dout(w_dff_B_Tah9espN4_0),.clk(gclk));
	jdff dff_B_uT0vOAA74_0(.din(w_dff_B_Tah9espN4_0),.dout(w_dff_B_uT0vOAA74_0),.clk(gclk));
	jdff dff_B_lrFqCve71_0(.din(w_dff_B_uT0vOAA74_0),.dout(w_dff_B_lrFqCve71_0),.clk(gclk));
	jdff dff_B_04iIw3AU5_0(.din(w_dff_B_lrFqCve71_0),.dout(w_dff_B_04iIw3AU5_0),.clk(gclk));
	jdff dff_B_VGzPUyC36_0(.din(w_dff_B_04iIw3AU5_0),.dout(w_dff_B_VGzPUyC36_0),.clk(gclk));
	jdff dff_B_bYh6fuTv8_0(.din(w_dff_B_VGzPUyC36_0),.dout(w_dff_B_bYh6fuTv8_0),.clk(gclk));
	jdff dff_B_RZOzaCt11_1(.din(n1006),.dout(w_dff_B_RZOzaCt11_1),.clk(gclk));
	jdff dff_B_LVbo2nxR3_1(.din(w_dff_B_RZOzaCt11_1),.dout(w_dff_B_LVbo2nxR3_1),.clk(gclk));
	jdff dff_B_YZS4p8r72_1(.din(w_dff_B_LVbo2nxR3_1),.dout(w_dff_B_YZS4p8r72_1),.clk(gclk));
	jdff dff_B_OZuyXFgh3_0(.din(n1028),.dout(w_dff_B_OZuyXFgh3_0),.clk(gclk));
	jdff dff_B_TZeEagoR7_0(.din(w_dff_B_OZuyXFgh3_0),.dout(w_dff_B_TZeEagoR7_0),.clk(gclk));
	jdff dff_B_RNGNwtdz4_0(.din(w_dff_B_TZeEagoR7_0),.dout(w_dff_B_RNGNwtdz4_0),.clk(gclk));
	jdff dff_B_NrS56NpP3_0(.din(w_dff_B_RNGNwtdz4_0),.dout(w_dff_B_NrS56NpP3_0),.clk(gclk));
	jdff dff_B_UfNREkOv9_0(.din(w_dff_B_NrS56NpP3_0),.dout(w_dff_B_UfNREkOv9_0),.clk(gclk));
	jdff dff_B_3M7YxRyR4_0(.din(w_dff_B_UfNREkOv9_0),.dout(w_dff_B_3M7YxRyR4_0),.clk(gclk));
	jdff dff_B_2Jfz7Zt00_0(.din(w_dff_B_3M7YxRyR4_0),.dout(w_dff_B_2Jfz7Zt00_0),.clk(gclk));
	jdff dff_B_4UOLOE5W6_0(.din(w_dff_B_2Jfz7Zt00_0),.dout(w_dff_B_4UOLOE5W6_0),.clk(gclk));
	jdff dff_B_q2lMszzI4_0(.din(w_dff_B_4UOLOE5W6_0),.dout(w_dff_B_q2lMszzI4_0),.clk(gclk));
	jdff dff_B_TotN7z2m8_0(.din(w_dff_B_q2lMszzI4_0),.dout(w_dff_B_TotN7z2m8_0),.clk(gclk));
	jdff dff_B_hqeALvmp3_0(.din(w_dff_B_TotN7z2m8_0),.dout(w_dff_B_hqeALvmp3_0),.clk(gclk));
	jdff dff_B_IFuUqoQf6_0(.din(w_dff_B_hqeALvmp3_0),.dout(w_dff_B_IFuUqoQf6_0),.clk(gclk));
	jdff dff_B_tXLsthCU3_0(.din(w_dff_B_IFuUqoQf6_0),.dout(w_dff_B_tXLsthCU3_0),.clk(gclk));
	jdff dff_B_WQB4AGs89_0(.din(w_dff_B_tXLsthCU3_0),.dout(w_dff_B_WQB4AGs89_0),.clk(gclk));
	jdff dff_B_5mZAup1X2_0(.din(w_dff_B_WQB4AGs89_0),.dout(w_dff_B_5mZAup1X2_0),.clk(gclk));
	jdff dff_B_baGPJQFF2_0(.din(w_dff_B_5mZAup1X2_0),.dout(w_dff_B_baGPJQFF2_0),.clk(gclk));
	jdff dff_B_TSxWOlHm2_1(.din(n1020),.dout(w_dff_B_TSxWOlHm2_1),.clk(gclk));
	jdff dff_A_y0fqPlcu6_0(.dout(w_n800_4[0]),.din(w_dff_A_y0fqPlcu6_0),.clk(gclk));
	jdff dff_A_sbO4wRnm7_0(.dout(w_dff_A_y0fqPlcu6_0),.din(w_dff_A_sbO4wRnm7_0),.clk(gclk));
	jdff dff_A_7fY6GrcM0_0(.dout(w_dff_A_sbO4wRnm7_0),.din(w_dff_A_7fY6GrcM0_0),.clk(gclk));
	jdff dff_A_XvKYeoGL6_0(.dout(w_dff_A_7fY6GrcM0_0),.din(w_dff_A_XvKYeoGL6_0),.clk(gclk));
	jdff dff_A_lfP0Vq4G8_0(.dout(w_dff_A_XvKYeoGL6_0),.din(w_dff_A_lfP0Vq4G8_0),.clk(gclk));
	jdff dff_A_XGsL5Nx21_0(.dout(w_dff_A_lfP0Vq4G8_0),.din(w_dff_A_XGsL5Nx21_0),.clk(gclk));
	jdff dff_A_i5zeMe8m5_0(.dout(w_dff_A_XGsL5Nx21_0),.din(w_dff_A_i5zeMe8m5_0),.clk(gclk));
	jdff dff_B_UkuSXVZ87_0(.din(n1039),.dout(w_dff_B_UkuSXVZ87_0),.clk(gclk));
	jdff dff_B_nvvzkRGz5_0(.din(w_dff_B_UkuSXVZ87_0),.dout(w_dff_B_nvvzkRGz5_0),.clk(gclk));
	jdff dff_B_mOfkBuob3_0(.din(w_dff_B_nvvzkRGz5_0),.dout(w_dff_B_mOfkBuob3_0),.clk(gclk));
	jdff dff_B_fVx42glE8_0(.din(w_dff_B_mOfkBuob3_0),.dout(w_dff_B_fVx42glE8_0),.clk(gclk));
	jdff dff_B_pwUFTuat9_0(.din(w_dff_B_fVx42glE8_0),.dout(w_dff_B_pwUFTuat9_0),.clk(gclk));
	jdff dff_B_A7VEBaJA1_0(.din(w_dff_B_pwUFTuat9_0),.dout(w_dff_B_A7VEBaJA1_0),.clk(gclk));
	jdff dff_B_hpv8jVYK1_0(.din(w_dff_B_A7VEBaJA1_0),.dout(w_dff_B_hpv8jVYK1_0),.clk(gclk));
	jdff dff_B_xIKTjiuK4_0(.din(w_dff_B_hpv8jVYK1_0),.dout(w_dff_B_xIKTjiuK4_0),.clk(gclk));
	jdff dff_B_I5o47Je97_0(.din(w_dff_B_xIKTjiuK4_0),.dout(w_dff_B_I5o47Je97_0),.clk(gclk));
	jdff dff_B_9apthTB20_0(.din(w_dff_B_I5o47Je97_0),.dout(w_dff_B_9apthTB20_0),.clk(gclk));
	jdff dff_B_GC6dFs5Q2_0(.din(w_dff_B_9apthTB20_0),.dout(w_dff_B_GC6dFs5Q2_0),.clk(gclk));
	jdff dff_B_ZZA6qjNH5_0(.din(w_dff_B_GC6dFs5Q2_0),.dout(w_dff_B_ZZA6qjNH5_0),.clk(gclk));
	jdff dff_B_ljwCGGod1_0(.din(w_dff_B_ZZA6qjNH5_0),.dout(w_dff_B_ljwCGGod1_0),.clk(gclk));
	jdff dff_B_jRLIr8sL6_0(.din(w_dff_B_ljwCGGod1_0),.dout(w_dff_B_jRLIr8sL6_0),.clk(gclk));
	jdff dff_B_vsXxz3Ng1_0(.din(w_dff_B_jRLIr8sL6_0),.dout(w_dff_B_vsXxz3Ng1_0),.clk(gclk));
	jdff dff_B_PWB45Tqz8_1(.din(n1031),.dout(w_dff_B_PWB45Tqz8_1),.clk(gclk));
	jdff dff_B_Y8Qdl6VR9_1(.din(w_dff_B_PWB45Tqz8_1),.dout(w_dff_B_Y8Qdl6VR9_1),.clk(gclk));
	jdff dff_B_ZPONdbT25_0(.din(n1050),.dout(w_dff_B_ZPONdbT25_0),.clk(gclk));
	jdff dff_B_48vW2mRd5_0(.din(w_dff_B_ZPONdbT25_0),.dout(w_dff_B_48vW2mRd5_0),.clk(gclk));
	jdff dff_B_6R72KguM9_0(.din(w_dff_B_48vW2mRd5_0),.dout(w_dff_B_6R72KguM9_0),.clk(gclk));
	jdff dff_B_FR9HuwVd8_0(.din(w_dff_B_6R72KguM9_0),.dout(w_dff_B_FR9HuwVd8_0),.clk(gclk));
	jdff dff_B_V6Eikr194_0(.din(w_dff_B_FR9HuwVd8_0),.dout(w_dff_B_V6Eikr194_0),.clk(gclk));
	jdff dff_B_7rlcIVMq2_0(.din(w_dff_B_V6Eikr194_0),.dout(w_dff_B_7rlcIVMq2_0),.clk(gclk));
	jdff dff_B_FglxMB1B0_0(.din(w_dff_B_7rlcIVMq2_0),.dout(w_dff_B_FglxMB1B0_0),.clk(gclk));
	jdff dff_B_y7Lshb6E1_0(.din(w_dff_B_FglxMB1B0_0),.dout(w_dff_B_y7Lshb6E1_0),.clk(gclk));
	jdff dff_B_0aXLOIpJ1_0(.din(w_dff_B_y7Lshb6E1_0),.dout(w_dff_B_0aXLOIpJ1_0),.clk(gclk));
	jdff dff_B_1WBtCBOx5_0(.din(w_dff_B_0aXLOIpJ1_0),.dout(w_dff_B_1WBtCBOx5_0),.clk(gclk));
	jdff dff_B_OGsxnyeT8_0(.din(w_dff_B_1WBtCBOx5_0),.dout(w_dff_B_OGsxnyeT8_0),.clk(gclk));
	jdff dff_B_gvGwydth1_0(.din(w_dff_B_OGsxnyeT8_0),.dout(w_dff_B_gvGwydth1_0),.clk(gclk));
	jdff dff_B_D13BJunD9_0(.din(w_dff_B_gvGwydth1_0),.dout(w_dff_B_D13BJunD9_0),.clk(gclk));
	jdff dff_B_8s8YOFXV9_1(.din(n1042),.dout(w_dff_B_8s8YOFXV9_1),.clk(gclk));
	jdff dff_B_PgOL7VEo2_0(.din(n1061),.dout(w_dff_B_PgOL7VEo2_0),.clk(gclk));
	jdff dff_B_E3OnIGUU0_0(.din(w_dff_B_PgOL7VEo2_0),.dout(w_dff_B_E3OnIGUU0_0),.clk(gclk));
	jdff dff_B_eiIB6mQO3_0(.din(w_dff_B_E3OnIGUU0_0),.dout(w_dff_B_eiIB6mQO3_0),.clk(gclk));
	jdff dff_B_UlwlA0fX1_0(.din(w_dff_B_eiIB6mQO3_0),.dout(w_dff_B_UlwlA0fX1_0),.clk(gclk));
	jdff dff_B_B2REas4L4_0(.din(w_dff_B_UlwlA0fX1_0),.dout(w_dff_B_B2REas4L4_0),.clk(gclk));
	jdff dff_B_HlK88dhT0_0(.din(w_dff_B_B2REas4L4_0),.dout(w_dff_B_HlK88dhT0_0),.clk(gclk));
	jdff dff_B_kpM6Du0e2_0(.din(w_dff_B_HlK88dhT0_0),.dout(w_dff_B_kpM6Du0e2_0),.clk(gclk));
	jdff dff_B_ZQYkGd7d7_0(.din(w_dff_B_kpM6Du0e2_0),.dout(w_dff_B_ZQYkGd7d7_0),.clk(gclk));
	jdff dff_B_oH8U7Bho9_0(.din(w_dff_B_ZQYkGd7d7_0),.dout(w_dff_B_oH8U7Bho9_0),.clk(gclk));
	jdff dff_B_q6YpXPcs4_0(.din(w_dff_B_oH8U7Bho9_0),.dout(w_dff_B_q6YpXPcs4_0),.clk(gclk));
	jdff dff_B_DlVTVJYc3_0(.din(w_dff_B_q6YpXPcs4_0),.dout(w_dff_B_DlVTVJYc3_0),.clk(gclk));
	jdff dff_B_y0Ay3AzT5_0(.din(w_dff_B_DlVTVJYc3_0),.dout(w_dff_B_y0Ay3AzT5_0),.clk(gclk));
	jdff dff_B_3Jkd2jMy3_0(.din(w_dff_B_y0Ay3AzT5_0),.dout(w_dff_B_3Jkd2jMy3_0),.clk(gclk));
	jdff dff_B_TocnJ47N6_0(.din(w_dff_B_3Jkd2jMy3_0),.dout(w_dff_B_TocnJ47N6_0),.clk(gclk));
	jdff dff_B_kyKZDjEP3_1(.din(n1053),.dout(w_dff_B_kyKZDjEP3_1),.clk(gclk));
	jdff dff_B_8WwbDecL4_1(.din(w_dff_B_kyKZDjEP3_1),.dout(w_dff_B_8WwbDecL4_1),.clk(gclk));
	jdff dff_B_66V6EbF32_1(.din(w_dff_B_8WwbDecL4_1),.dout(w_dff_B_66V6EbF32_1),.clk(gclk));
	jdff dff_A_OzL5O6s65_0(.dout(w_n800_3[0]),.din(w_dff_A_OzL5O6s65_0),.clk(gclk));
	jdff dff_A_mSNHzLrI6_2(.dout(w_n800_3[2]),.din(w_dff_A_mSNHzLrI6_2),.clk(gclk));
	jdff dff_A_AHqMAjRY7_2(.dout(w_dff_A_mSNHzLrI6_2),.din(w_dff_A_AHqMAjRY7_2),.clk(gclk));
	jdff dff_B_P7G6dOCY0_1(.din(n1066),.dout(w_dff_B_P7G6dOCY0_1),.clk(gclk));
	jdff dff_B_iDUut8Ig3_1(.din(w_dff_B_P7G6dOCY0_1),.dout(w_dff_B_iDUut8Ig3_1),.clk(gclk));
	jdff dff_B_HlHw4r4Z8_1(.din(w_dff_B_iDUut8Ig3_1),.dout(w_dff_B_HlHw4r4Z8_1),.clk(gclk));
	jdff dff_B_mAETDW4n0_1(.din(w_dff_B_HlHw4r4Z8_1),.dout(w_dff_B_mAETDW4n0_1),.clk(gclk));
	jdff dff_B_Ss7mZ6oL8_1(.din(w_dff_B_mAETDW4n0_1),.dout(w_dff_B_Ss7mZ6oL8_1),.clk(gclk));
	jdff dff_B_6SRlSjqt5_1(.din(w_dff_B_Ss7mZ6oL8_1),.dout(w_dff_B_6SRlSjqt5_1),.clk(gclk));
	jdff dff_B_KHObKrTC0_1(.din(w_dff_B_6SRlSjqt5_1),.dout(w_dff_B_KHObKrTC0_1),.clk(gclk));
	jdff dff_B_TCJLlppF8_1(.din(w_dff_B_KHObKrTC0_1),.dout(w_dff_B_TCJLlppF8_1),.clk(gclk));
	jdff dff_B_aav5VX5B9_1(.din(w_dff_B_TCJLlppF8_1),.dout(w_dff_B_aav5VX5B9_1),.clk(gclk));
	jdff dff_B_avB97Oq41_1(.din(w_dff_B_aav5VX5B9_1),.dout(w_dff_B_avB97Oq41_1),.clk(gclk));
	jdff dff_B_shrUwFB68_1(.din(w_dff_B_avB97Oq41_1),.dout(w_dff_B_shrUwFB68_1),.clk(gclk));
	jdff dff_B_nMke7Iym7_1(.din(w_dff_B_shrUwFB68_1),.dout(w_dff_B_nMke7Iym7_1),.clk(gclk));
	jdff dff_B_9cgTWemn0_1(.din(w_dff_B_nMke7Iym7_1),.dout(w_dff_B_9cgTWemn0_1),.clk(gclk));
	jdff dff_B_z0ktVAng5_1(.din(w_dff_B_9cgTWemn0_1),.dout(w_dff_B_z0ktVAng5_1),.clk(gclk));
	jdff dff_B_0rAy1vbr2_1(.din(w_dff_B_z0ktVAng5_1),.dout(w_dff_B_0rAy1vbr2_1),.clk(gclk));
	jdff dff_A_p1TMc0sP2_0(.dout(w_n854_4[0]),.din(w_dff_A_p1TMc0sP2_0),.clk(gclk));
	jdff dff_A_o7YhbvWz6_0(.dout(w_dff_A_p1TMc0sP2_0),.din(w_dff_A_o7YhbvWz6_0),.clk(gclk));
	jdff dff_A_kC6bmOQa3_0(.dout(w_dff_A_o7YhbvWz6_0),.din(w_dff_A_kC6bmOQa3_0),.clk(gclk));
	jdff dff_A_3TdTeVSQ9_0(.dout(w_dff_A_kC6bmOQa3_0),.din(w_dff_A_3TdTeVSQ9_0),.clk(gclk));
	jdff dff_A_gt2pzEm99_0(.dout(w_dff_A_3TdTeVSQ9_0),.din(w_dff_A_gt2pzEm99_0),.clk(gclk));
	jdff dff_A_Ph7CHpmE9_0(.dout(w_dff_A_gt2pzEm99_0),.din(w_dff_A_Ph7CHpmE9_0),.clk(gclk));
	jdff dff_A_fjg75LeW8_0(.dout(w_dff_A_Ph7CHpmE9_0),.din(w_dff_A_fjg75LeW8_0),.clk(gclk));
	jdff dff_A_EjKLw5jY3_0(.dout(w_dff_A_fjg75LeW8_0),.din(w_dff_A_EjKLw5jY3_0),.clk(gclk));
	jdff dff_B_MLk6KA3G8_1(.din(n1075),.dout(w_dff_B_MLk6KA3G8_1),.clk(gclk));
	jdff dff_B_ZZuCoweL7_1(.din(w_dff_B_MLk6KA3G8_1),.dout(w_dff_B_ZZuCoweL7_1),.clk(gclk));
	jdff dff_B_Qscbnwhp2_1(.din(w_dff_B_ZZuCoweL7_1),.dout(w_dff_B_Qscbnwhp2_1),.clk(gclk));
	jdff dff_B_plH4Uu8A8_1(.din(w_dff_B_Qscbnwhp2_1),.dout(w_dff_B_plH4Uu8A8_1),.clk(gclk));
	jdff dff_B_6qR45CO72_1(.din(w_dff_B_plH4Uu8A8_1),.dout(w_dff_B_6qR45CO72_1),.clk(gclk));
	jdff dff_B_V0UDLpRB9_1(.din(w_dff_B_6qR45CO72_1),.dout(w_dff_B_V0UDLpRB9_1),.clk(gclk));
	jdff dff_B_ZaiO6gz98_1(.din(w_dff_B_V0UDLpRB9_1),.dout(w_dff_B_ZaiO6gz98_1),.clk(gclk));
	jdff dff_B_JZMAV0XQ6_1(.din(w_dff_B_ZaiO6gz98_1),.dout(w_dff_B_JZMAV0XQ6_1),.clk(gclk));
	jdff dff_B_WfXQttZa4_1(.din(w_dff_B_JZMAV0XQ6_1),.dout(w_dff_B_WfXQttZa4_1),.clk(gclk));
	jdff dff_B_Y2CBN6gi9_1(.din(w_dff_B_WfXQttZa4_1),.dout(w_dff_B_Y2CBN6gi9_1),.clk(gclk));
	jdff dff_B_lAYgpfSH5_1(.din(w_dff_B_Y2CBN6gi9_1),.dout(w_dff_B_lAYgpfSH5_1),.clk(gclk));
	jdff dff_B_dtzgPbxY0_1(.din(w_dff_B_lAYgpfSH5_1),.dout(w_dff_B_dtzgPbxY0_1),.clk(gclk));
	jdff dff_B_3IJSS4FF6_1(.din(w_dff_B_dtzgPbxY0_1),.dout(w_dff_B_3IJSS4FF6_1),.clk(gclk));
	jdff dff_B_WO2QjJZx1_1(.din(w_dff_B_3IJSS4FF6_1),.dout(w_dff_B_WO2QjJZx1_1),.clk(gclk));
	jdff dff_B_WtjqIDdJ3_0(.din(n1077),.dout(w_dff_B_WtjqIDdJ3_0),.clk(gclk));
	jdff dff_B_Wk9Y8kd14_1(.din(n1084),.dout(w_dff_B_Wk9Y8kd14_1),.clk(gclk));
	jdff dff_B_wptY5y6H0_1(.din(w_dff_B_Wk9Y8kd14_1),.dout(w_dff_B_wptY5y6H0_1),.clk(gclk));
	jdff dff_B_I0MucakO7_1(.din(w_dff_B_wptY5y6H0_1),.dout(w_dff_B_I0MucakO7_1),.clk(gclk));
	jdff dff_B_naT1y9Xs0_1(.din(w_dff_B_I0MucakO7_1),.dout(w_dff_B_naT1y9Xs0_1),.clk(gclk));
	jdff dff_B_RzAhAgK08_1(.din(w_dff_B_naT1y9Xs0_1),.dout(w_dff_B_RzAhAgK08_1),.clk(gclk));
	jdff dff_B_eyWrL4c61_1(.din(w_dff_B_RzAhAgK08_1),.dout(w_dff_B_eyWrL4c61_1),.clk(gclk));
	jdff dff_B_eknu4SOh1_1(.din(w_dff_B_eyWrL4c61_1),.dout(w_dff_B_eknu4SOh1_1),.clk(gclk));
	jdff dff_B_VPfWt4Ou7_1(.din(w_dff_B_eknu4SOh1_1),.dout(w_dff_B_VPfWt4Ou7_1),.clk(gclk));
	jdff dff_B_9O0tHRuR8_1(.din(w_dff_B_VPfWt4Ou7_1),.dout(w_dff_B_9O0tHRuR8_1),.clk(gclk));
	jdff dff_B_2PdW1mX86_1(.din(w_dff_B_9O0tHRuR8_1),.dout(w_dff_B_2PdW1mX86_1),.clk(gclk));
	jdff dff_B_pxtOYEPZ7_1(.din(w_dff_B_2PdW1mX86_1),.dout(w_dff_B_pxtOYEPZ7_1),.clk(gclk));
	jdff dff_B_vdVDT8fO7_1(.din(w_dff_B_pxtOYEPZ7_1),.dout(w_dff_B_vdVDT8fO7_1),.clk(gclk));
	jdff dff_B_nzWmdS5U0_0(.din(n1097),.dout(w_dff_B_nzWmdS5U0_0),.clk(gclk));
	jdff dff_B_nh0Zbccj3_0(.din(w_dff_B_nzWmdS5U0_0),.dout(w_dff_B_nh0Zbccj3_0),.clk(gclk));
	jdff dff_B_zlEUIu1y4_0(.din(w_dff_B_nh0Zbccj3_0),.dout(w_dff_B_zlEUIu1y4_0),.clk(gclk));
	jdff dff_B_FXJ24YZv4_0(.din(w_dff_B_zlEUIu1y4_0),.dout(w_dff_B_FXJ24YZv4_0),.clk(gclk));
	jdff dff_B_JshCWRao6_0(.din(w_dff_B_FXJ24YZv4_0),.dout(w_dff_B_JshCWRao6_0),.clk(gclk));
	jdff dff_B_RooTn53j1_0(.din(w_dff_B_JshCWRao6_0),.dout(w_dff_B_RooTn53j1_0),.clk(gclk));
	jdff dff_B_7hba4mDo1_0(.din(w_dff_B_RooTn53j1_0),.dout(w_dff_B_7hba4mDo1_0),.clk(gclk));
	jdff dff_B_Tdyjeyzi3_0(.din(w_dff_B_7hba4mDo1_0),.dout(w_dff_B_Tdyjeyzi3_0),.clk(gclk));
	jdff dff_B_cpcPuiuM3_0(.din(w_dff_B_Tdyjeyzi3_0),.dout(w_dff_B_cpcPuiuM3_0),.clk(gclk));
	jdff dff_B_jnCmFogt4_0(.din(w_dff_B_cpcPuiuM3_0),.dout(w_dff_B_jnCmFogt4_0),.clk(gclk));
	jdff dff_B_a20HcxR97_0(.din(w_dff_B_jnCmFogt4_0),.dout(w_dff_B_a20HcxR97_0),.clk(gclk));
	jdff dff_B_xm2v5N5I8_0(.din(w_dff_B_a20HcxR97_0),.dout(w_dff_B_xm2v5N5I8_0),.clk(gclk));
	jdff dff_B_zX9qkJnc3_0(.din(w_dff_B_xm2v5N5I8_0),.dout(w_dff_B_zX9qkJnc3_0),.clk(gclk));
	jdff dff_B_ePcFd7uz4_0(.din(w_dff_B_zX9qkJnc3_0),.dout(w_dff_B_ePcFd7uz4_0),.clk(gclk));
	jdff dff_B_6TYDbxhT4_1(.din(n1090),.dout(w_dff_B_6TYDbxhT4_1),.clk(gclk));
	jdff dff_B_9HSbRjVc2_1(.din(w_dff_B_6TYDbxhT4_1),.dout(w_dff_B_9HSbRjVc2_1),.clk(gclk));
	jdff dff_B_rdYUYjWb3_1(.din(w_dff_B_9HSbRjVc2_1),.dout(w_dff_B_rdYUYjWb3_1),.clk(gclk));
	jdff dff_A_yuVUJRug6_2(.dout(w_n854_3[2]),.din(w_dff_A_yuVUJRug6_2),.clk(gclk));
	jdff dff_A_P2s8uA8u4_2(.dout(w_dff_A_yuVUJRug6_2),.din(w_dff_A_P2s8uA8u4_2),.clk(gclk));
	jdff dff_B_dlYx2j1Q4_0(.din(n1105),.dout(w_dff_B_dlYx2j1Q4_0),.clk(gclk));
	jdff dff_B_sNuZ5cFE9_0(.din(w_dff_B_dlYx2j1Q4_0),.dout(w_dff_B_sNuZ5cFE9_0),.clk(gclk));
	jdff dff_B_HoCY4SA79_0(.din(w_dff_B_sNuZ5cFE9_0),.dout(w_dff_B_HoCY4SA79_0),.clk(gclk));
	jdff dff_B_RlwrtYV62_0(.din(w_dff_B_HoCY4SA79_0),.dout(w_dff_B_RlwrtYV62_0),.clk(gclk));
	jdff dff_B_5Yy2qkgE2_0(.din(w_dff_B_RlwrtYV62_0),.dout(w_dff_B_5Yy2qkgE2_0),.clk(gclk));
	jdff dff_B_fsvYl8F98_0(.din(w_dff_B_5Yy2qkgE2_0),.dout(w_dff_B_fsvYl8F98_0),.clk(gclk));
	jdff dff_B_U8RIMQyq1_0(.din(w_dff_B_fsvYl8F98_0),.dout(w_dff_B_U8RIMQyq1_0),.clk(gclk));
	jdff dff_B_S68Ih2m87_0(.din(w_dff_B_U8RIMQyq1_0),.dout(w_dff_B_S68Ih2m87_0),.clk(gclk));
	jdff dff_B_eBnMiTXi9_0(.din(w_dff_B_S68Ih2m87_0),.dout(w_dff_B_eBnMiTXi9_0),.clk(gclk));
	jdff dff_B_rZQAnHAz7_0(.din(w_dff_B_eBnMiTXi9_0),.dout(w_dff_B_rZQAnHAz7_0),.clk(gclk));
	jdff dff_B_xVAPP0WQ9_0(.din(w_dff_B_rZQAnHAz7_0),.dout(w_dff_B_xVAPP0WQ9_0),.clk(gclk));
	jdff dff_B_obB8VCKb3_0(.din(w_dff_B_xVAPP0WQ9_0),.dout(w_dff_B_obB8VCKb3_0),.clk(gclk));
	jdff dff_B_OQ2cJw1E0_0(.din(w_dff_B_obB8VCKb3_0),.dout(w_dff_B_OQ2cJw1E0_0),.clk(gclk));
	jdff dff_B_yyBZyRr94_0(.din(w_dff_B_OQ2cJw1E0_0),.dout(w_dff_B_yyBZyRr94_0),.clk(gclk));
	jdff dff_B_Hci9Zji85_0(.din(w_dff_B_yyBZyRr94_0),.dout(w_dff_B_Hci9Zji85_0),.clk(gclk));
	jdff dff_B_b3hbbYEy1_1(.din(n1099),.dout(w_dff_B_b3hbbYEy1_1),.clk(gclk));
	jdff dff_B_XMnLS7YG8_0(.din(n1114),.dout(w_dff_B_XMnLS7YG8_0),.clk(gclk));
	jdff dff_B_UO0V1KFA6_0(.din(w_dff_B_XMnLS7YG8_0),.dout(w_dff_B_UO0V1KFA6_0),.clk(gclk));
	jdff dff_B_QIpU5tY40_0(.din(w_dff_B_UO0V1KFA6_0),.dout(w_dff_B_QIpU5tY40_0),.clk(gclk));
	jdff dff_B_At0f5HrN7_0(.din(w_dff_B_QIpU5tY40_0),.dout(w_dff_B_At0f5HrN7_0),.clk(gclk));
	jdff dff_B_0oCccyPS5_0(.din(w_dff_B_At0f5HrN7_0),.dout(w_dff_B_0oCccyPS5_0),.clk(gclk));
	jdff dff_B_EPKsemQA7_0(.din(w_dff_B_0oCccyPS5_0),.dout(w_dff_B_EPKsemQA7_0),.clk(gclk));
	jdff dff_B_jHDUVhod8_0(.din(w_dff_B_EPKsemQA7_0),.dout(w_dff_B_jHDUVhod8_0),.clk(gclk));
	jdff dff_B_CkjCoHxC9_0(.din(w_dff_B_jHDUVhod8_0),.dout(w_dff_B_CkjCoHxC9_0),.clk(gclk));
	jdff dff_B_3Y0GYcFm4_0(.din(w_dff_B_CkjCoHxC9_0),.dout(w_dff_B_3Y0GYcFm4_0),.clk(gclk));
	jdff dff_B_UdI0GnYB9_0(.din(w_dff_B_3Y0GYcFm4_0),.dout(w_dff_B_UdI0GnYB9_0),.clk(gclk));
	jdff dff_B_rmEus8dW7_0(.din(w_dff_B_UdI0GnYB9_0),.dout(w_dff_B_rmEus8dW7_0),.clk(gclk));
	jdff dff_B_Suvoinvj4_0(.din(w_dff_B_rmEus8dW7_0),.dout(w_dff_B_Suvoinvj4_0),.clk(gclk));
	jdff dff_B_YpGI6jln1_0(.din(n1110),.dout(w_dff_B_YpGI6jln1_0),.clk(gclk));
	jdff dff_A_rEkd99D39_0(.dout(w_n999_3[0]),.din(w_dff_A_rEkd99D39_0),.clk(gclk));
	jdff dff_A_HGhebhM94_0(.dout(w_dff_A_rEkd99D39_0),.din(w_dff_A_HGhebhM94_0),.clk(gclk));
	jdff dff_A_MwSGsGmt7_0(.dout(w_dff_A_HGhebhM94_0),.din(w_dff_A_MwSGsGmt7_0),.clk(gclk));
	jdff dff_A_kcapujoy5_1(.dout(w_n999_3[1]),.din(w_dff_A_kcapujoy5_1),.clk(gclk));
	jdff dff_A_zIehUUja3_1(.dout(w_dff_A_kcapujoy5_1),.din(w_dff_A_zIehUUja3_1),.clk(gclk));
	jdff dff_A_1dzGRIFT0_1(.dout(w_dff_A_zIehUUja3_1),.din(w_dff_A_1dzGRIFT0_1),.clk(gclk));
	jdff dff_A_X5yVBLaX7_1(.dout(w_dff_A_1dzGRIFT0_1),.din(w_dff_A_X5yVBLaX7_1),.clk(gclk));
	jdff dff_A_ALTtceVh9_1(.dout(w_dff_A_X5yVBLaX7_1),.din(w_dff_A_ALTtceVh9_1),.clk(gclk));
	jdff dff_A_xD53gBXo1_1(.dout(w_dff_A_ALTtceVh9_1),.din(w_dff_A_xD53gBXo1_1),.clk(gclk));
	jdff dff_A_ZHlsjuj38_1(.dout(w_dff_A_xD53gBXo1_1),.din(w_dff_A_ZHlsjuj38_1),.clk(gclk));
	jdff dff_A_kkwRc1Fa1_0(.dout(w_G1689_4[0]),.din(w_dff_A_kkwRc1Fa1_0),.clk(gclk));
	jdff dff_A_9JDF0wyn4_0(.dout(w_dff_A_kkwRc1Fa1_0),.din(w_dff_A_9JDF0wyn4_0),.clk(gclk));
	jdff dff_A_LJznGtt23_0(.dout(w_dff_A_9JDF0wyn4_0),.din(w_dff_A_LJznGtt23_0),.clk(gclk));
	jdff dff_A_LFhCZYSH3_0(.dout(w_dff_A_LJznGtt23_0),.din(w_dff_A_LFhCZYSH3_0),.clk(gclk));
	jdff dff_A_ULX69nvB6_0(.dout(w_dff_A_LFhCZYSH3_0),.din(w_dff_A_ULX69nvB6_0),.clk(gclk));
	jdff dff_A_UPrmTDyU9_1(.dout(w_G1689_4[1]),.din(w_dff_A_UPrmTDyU9_1),.clk(gclk));
	jdff dff_A_89LOEPJJ0_1(.dout(w_dff_A_UPrmTDyU9_1),.din(w_dff_A_89LOEPJJ0_1),.clk(gclk));
	jdff dff_A_l6gYRpAo7_1(.dout(w_dff_A_89LOEPJJ0_1),.din(w_dff_A_l6gYRpAo7_1),.clk(gclk));
	jdff dff_A_7cuavIbH0_1(.dout(w_dff_A_l6gYRpAo7_1),.din(w_dff_A_7cuavIbH0_1),.clk(gclk));
	jdff dff_A_fG87pw2R0_1(.dout(w_dff_A_7cuavIbH0_1),.din(w_dff_A_fG87pw2R0_1),.clk(gclk));
	jdff dff_A_2lyjNTof5_1(.dout(w_dff_A_fG87pw2R0_1),.din(w_dff_A_2lyjNTof5_1),.clk(gclk));
	jdff dff_A_JdFhaelb0_1(.dout(w_dff_A_2lyjNTof5_1),.din(w_dff_A_JdFhaelb0_1),.clk(gclk));
	jdff dff_B_2fsWrDcZ2_0(.din(n1123),.dout(w_dff_B_2fsWrDcZ2_0),.clk(gclk));
	jdff dff_B_dHBPR1nd2_0(.din(w_dff_B_2fsWrDcZ2_0),.dout(w_dff_B_dHBPR1nd2_0),.clk(gclk));
	jdff dff_B_7jUGA8E67_0(.din(w_dff_B_dHBPR1nd2_0),.dout(w_dff_B_7jUGA8E67_0),.clk(gclk));
	jdff dff_B_9elJXMvt8_0(.din(w_dff_B_7jUGA8E67_0),.dout(w_dff_B_9elJXMvt8_0),.clk(gclk));
	jdff dff_B_DsHfFmhI8_0(.din(w_dff_B_9elJXMvt8_0),.dout(w_dff_B_DsHfFmhI8_0),.clk(gclk));
	jdff dff_B_WSXC1QKs9_0(.din(w_dff_B_DsHfFmhI8_0),.dout(w_dff_B_WSXC1QKs9_0),.clk(gclk));
	jdff dff_B_aps5827G2_0(.din(w_dff_B_WSXC1QKs9_0),.dout(w_dff_B_aps5827G2_0),.clk(gclk));
	jdff dff_B_4SatGGgD4_0(.din(w_dff_B_aps5827G2_0),.dout(w_dff_B_4SatGGgD4_0),.clk(gclk));
	jdff dff_B_Q1Aglej13_0(.din(w_dff_B_4SatGGgD4_0),.dout(w_dff_B_Q1Aglej13_0),.clk(gclk));
	jdff dff_B_brgsmrrX9_0(.din(w_dff_B_Q1Aglej13_0),.dout(w_dff_B_brgsmrrX9_0),.clk(gclk));
	jdff dff_B_Bk8tETIl3_0(.din(w_dff_B_brgsmrrX9_0),.dout(w_dff_B_Bk8tETIl3_0),.clk(gclk));
	jdff dff_B_Y7YB1tXd4_0(.din(w_dff_B_Bk8tETIl3_0),.dout(w_dff_B_Y7YB1tXd4_0),.clk(gclk));
	jdff dff_B_PvQKJ1lH9_1(.din(n1117),.dout(w_dff_B_PvQKJ1lH9_1),.clk(gclk));
	jdff dff_A_LHTlblFS7_2(.dout(w_G137_8[2]),.din(w_dff_A_LHTlblFS7_2),.clk(gclk));
	jdff dff_A_QgzC8xx93_2(.dout(w_dff_A_LHTlblFS7_2),.din(w_dff_A_QgzC8xx93_2),.clk(gclk));
	jdff dff_A_CbUuo9Gv3_2(.dout(w_dff_A_QgzC8xx93_2),.din(w_dff_A_CbUuo9Gv3_2),.clk(gclk));
	jdff dff_B_Js8RLDsD4_0(.din(n1132),.dout(w_dff_B_Js8RLDsD4_0),.clk(gclk));
	jdff dff_B_Drjgelto1_0(.din(w_dff_B_Js8RLDsD4_0),.dout(w_dff_B_Drjgelto1_0),.clk(gclk));
	jdff dff_B_CMJUo9XR2_0(.din(w_dff_B_Drjgelto1_0),.dout(w_dff_B_CMJUo9XR2_0),.clk(gclk));
	jdff dff_B_0pHUcuBP5_0(.din(w_dff_B_CMJUo9XR2_0),.dout(w_dff_B_0pHUcuBP5_0),.clk(gclk));
	jdff dff_B_GDpbnEjJ8_0(.din(w_dff_B_0pHUcuBP5_0),.dout(w_dff_B_GDpbnEjJ8_0),.clk(gclk));
	jdff dff_B_Zhve6e8w0_0(.din(w_dff_B_GDpbnEjJ8_0),.dout(w_dff_B_Zhve6e8w0_0),.clk(gclk));
	jdff dff_B_KnwXlI7I8_0(.din(w_dff_B_Zhve6e8w0_0),.dout(w_dff_B_KnwXlI7I8_0),.clk(gclk));
	jdff dff_B_uymMJo6F5_0(.din(w_dff_B_KnwXlI7I8_0),.dout(w_dff_B_uymMJo6F5_0),.clk(gclk));
	jdff dff_B_FYTBqWQe6_0(.din(w_dff_B_uymMJo6F5_0),.dout(w_dff_B_FYTBqWQe6_0),.clk(gclk));
	jdff dff_B_3fMqkkZ20_0(.din(w_dff_B_FYTBqWQe6_0),.dout(w_dff_B_3fMqkkZ20_0),.clk(gclk));
	jdff dff_B_C3lzjKps7_0(.din(w_dff_B_3fMqkkZ20_0),.dout(w_dff_B_C3lzjKps7_0),.clk(gclk));
	jdff dff_B_c6InWFUx7_0(.din(w_dff_B_C3lzjKps7_0),.dout(w_dff_B_c6InWFUx7_0),.clk(gclk));
	jdff dff_B_Sq6Y1wZs9_0(.din(w_dff_B_c6InWFUx7_0),.dout(w_dff_B_Sq6Y1wZs9_0),.clk(gclk));
	jdff dff_A_kM4Ok63H1_0(.dout(w_n993_3[0]),.din(w_dff_A_kM4Ok63H1_0),.clk(gclk));
	jdff dff_A_F2Q6BTQG0_0(.dout(w_dff_A_kM4Ok63H1_0),.din(w_dff_A_F2Q6BTQG0_0),.clk(gclk));
	jdff dff_A_fhl7roYl2_1(.dout(w_n993_3[1]),.din(w_dff_A_fhl7roYl2_1),.clk(gclk));
	jdff dff_B_ybdAiMZK7_1(.din(n1135),.dout(w_dff_B_ybdAiMZK7_1),.clk(gclk));
	jdff dff_B_DwjsQlGf0_1(.din(w_dff_B_ybdAiMZK7_1),.dout(w_dff_B_DwjsQlGf0_1),.clk(gclk));
	jdff dff_B_cAQLgNRl4_1(.din(w_dff_B_DwjsQlGf0_1),.dout(w_dff_B_cAQLgNRl4_1),.clk(gclk));
	jdff dff_B_HsSKzZDF1_1(.din(w_dff_B_cAQLgNRl4_1),.dout(w_dff_B_HsSKzZDF1_1),.clk(gclk));
	jdff dff_B_CeNcjF2b4_1(.din(w_dff_B_HsSKzZDF1_1),.dout(w_dff_B_CeNcjF2b4_1),.clk(gclk));
	jdff dff_B_ACwUTcPA8_1(.din(w_dff_B_CeNcjF2b4_1),.dout(w_dff_B_ACwUTcPA8_1),.clk(gclk));
	jdff dff_B_FToaxKG98_1(.din(w_dff_B_ACwUTcPA8_1),.dout(w_dff_B_FToaxKG98_1),.clk(gclk));
	jdff dff_B_Z4wexT3S3_1(.din(w_dff_B_FToaxKG98_1),.dout(w_dff_B_Z4wexT3S3_1),.clk(gclk));
	jdff dff_B_8iD17oYr0_1(.din(w_dff_B_Z4wexT3S3_1),.dout(w_dff_B_8iD17oYr0_1),.clk(gclk));
	jdff dff_B_sBPiagre0_1(.din(w_dff_B_8iD17oYr0_1),.dout(w_dff_B_sBPiagre0_1),.clk(gclk));
	jdff dff_B_m7meNjhp8_1(.din(w_dff_B_sBPiagre0_1),.dout(w_dff_B_m7meNjhp8_1),.clk(gclk));
	jdff dff_B_2FbThkxa8_1(.din(w_dff_B_m7meNjhp8_1),.dout(w_dff_B_2FbThkxa8_1),.clk(gclk));
	jdff dff_B_lwChKyxl1_1(.din(w_dff_B_2FbThkxa8_1),.dout(w_dff_B_lwChKyxl1_1),.clk(gclk));
	jdff dff_B_37WBQKT70_1(.din(w_dff_B_lwChKyxl1_1),.dout(w_dff_B_37WBQKT70_1),.clk(gclk));
	jdff dff_B_8tWgp4Jh7_1(.din(w_dff_B_37WBQKT70_1),.dout(w_dff_B_8tWgp4Jh7_1),.clk(gclk));
	jdff dff_B_Fsu4cCZy0_1(.din(w_dff_B_8tWgp4Jh7_1),.dout(w_dff_B_Fsu4cCZy0_1),.clk(gclk));
	jdff dff_B_ILpdYLST9_1(.din(w_dff_B_Fsu4cCZy0_1),.dout(w_dff_B_ILpdYLST9_1),.clk(gclk));
	jdff dff_B_1Okr1deu8_1(.din(n1136),.dout(w_dff_B_1Okr1deu8_1),.clk(gclk));
	jdff dff_B_z0fjnVN23_1(.din(w_dff_B_1Okr1deu8_1),.dout(w_dff_B_z0fjnVN23_1),.clk(gclk));
	jdff dff_B_pYOdEXAk3_1(.din(w_dff_B_z0fjnVN23_1),.dout(w_dff_B_pYOdEXAk3_1),.clk(gclk));
	jdff dff_B_v3MvVb3h3_1(.din(w_dff_B_pYOdEXAk3_1),.dout(w_dff_B_v3MvVb3h3_1),.clk(gclk));
	jdff dff_B_d8Kx8qZ75_1(.din(w_dff_B_v3MvVb3h3_1),.dout(w_dff_B_d8Kx8qZ75_1),.clk(gclk));
	jdff dff_B_LvCcI1oo8_1(.din(w_dff_B_d8Kx8qZ75_1),.dout(w_dff_B_LvCcI1oo8_1),.clk(gclk));
	jdff dff_B_Wi9RNXN35_1(.din(w_dff_B_LvCcI1oo8_1),.dout(w_dff_B_Wi9RNXN35_1),.clk(gclk));
	jdff dff_B_fl36zeOT7_1(.din(w_dff_B_Wi9RNXN35_1),.dout(w_dff_B_fl36zeOT7_1),.clk(gclk));
	jdff dff_B_5thsbeGK3_1(.din(w_dff_B_fl36zeOT7_1),.dout(w_dff_B_5thsbeGK3_1),.clk(gclk));
	jdff dff_B_qDKTk91n6_1(.din(w_dff_B_5thsbeGK3_1),.dout(w_dff_B_qDKTk91n6_1),.clk(gclk));
	jdff dff_B_QcRAS6s42_1(.din(w_dff_B_qDKTk91n6_1),.dout(w_dff_B_QcRAS6s42_1),.clk(gclk));
	jdff dff_B_yLHma9SI5_1(.din(w_dff_B_QcRAS6s42_1),.dout(w_dff_B_yLHma9SI5_1),.clk(gclk));
	jdff dff_B_GkyL48KR9_1(.din(w_dff_B_yLHma9SI5_1),.dout(w_dff_B_GkyL48KR9_1),.clk(gclk));
	jdff dff_B_A7uZoiyP5_1(.din(w_dff_B_GkyL48KR9_1),.dout(w_dff_B_A7uZoiyP5_1),.clk(gclk));
	jdff dff_B_FnpRua1h8_1(.din(w_dff_B_A7uZoiyP5_1),.dout(w_dff_B_FnpRua1h8_1),.clk(gclk));
	jdff dff_B_6H7jaLad3_1(.din(w_dff_B_FnpRua1h8_1),.dout(w_dff_B_6H7jaLad3_1),.clk(gclk));
	jdff dff_B_DCt5fdP63_1(.din(w_dff_B_6H7jaLad3_1),.dout(w_dff_B_DCt5fdP63_1),.clk(gclk));
	jdff dff_B_TUFBbBAt5_1(.din(n811),.dout(w_dff_B_TUFBbBAt5_1),.clk(gclk));
	jdff dff_B_zXGAUlEA6_1(.din(w_dff_B_TUFBbBAt5_1),.dout(w_dff_B_zXGAUlEA6_1),.clk(gclk));
	jdff dff_B_MbKSQnhm4_1(.din(w_dff_B_zXGAUlEA6_1),.dout(w_dff_B_MbKSQnhm4_1),.clk(gclk));
	jdff dff_B_KVmAjwlj9_1(.din(w_dff_B_MbKSQnhm4_1),.dout(w_dff_B_KVmAjwlj9_1),.clk(gclk));
	jdff dff_B_XWUq6Fah9_1(.din(w_dff_B_KVmAjwlj9_1),.dout(w_dff_B_XWUq6Fah9_1),.clk(gclk));
	jdff dff_B_jP5Ik2EJ0_1(.din(w_dff_B_XWUq6Fah9_1),.dout(w_dff_B_jP5Ik2EJ0_1),.clk(gclk));
	jdff dff_B_tMHefNiG9_1(.din(w_dff_B_jP5Ik2EJ0_1),.dout(w_dff_B_tMHefNiG9_1),.clk(gclk));
	jdff dff_B_It6OdICZ9_1(.din(w_dff_B_tMHefNiG9_1),.dout(w_dff_B_It6OdICZ9_1),.clk(gclk));
	jdff dff_B_AjcHYoEb5_1(.din(w_dff_B_It6OdICZ9_1),.dout(w_dff_B_AjcHYoEb5_1),.clk(gclk));
	jdff dff_B_eluNYSm06_1(.din(w_dff_B_AjcHYoEb5_1),.dout(w_dff_B_eluNYSm06_1),.clk(gclk));
	jdff dff_B_nhvyUovY4_0(.din(n830),.dout(w_dff_B_nhvyUovY4_0),.clk(gclk));
	jdff dff_B_wOyIj7qj3_0(.din(w_dff_B_nhvyUovY4_0),.dout(w_dff_B_wOyIj7qj3_0),.clk(gclk));
	jdff dff_B_rQqkwRhB6_0(.din(w_dff_B_wOyIj7qj3_0),.dout(w_dff_B_rQqkwRhB6_0),.clk(gclk));
	jdff dff_B_65aqk9292_0(.din(w_dff_B_rQqkwRhB6_0),.dout(w_dff_B_65aqk9292_0),.clk(gclk));
	jdff dff_B_xjmPbzyC7_0(.din(w_dff_B_65aqk9292_0),.dout(w_dff_B_xjmPbzyC7_0),.clk(gclk));
	jdff dff_B_g4VSIKkr6_0(.din(w_dff_B_xjmPbzyC7_0),.dout(w_dff_B_g4VSIKkr6_0),.clk(gclk));
	jdff dff_B_P0QGvQNP1_1(.din(n822),.dout(w_dff_B_P0QGvQNP1_1),.clk(gclk));
	jdff dff_B_KtEtKJji2_1(.din(w_dff_B_P0QGvQNP1_1),.dout(w_dff_B_KtEtKJji2_1),.clk(gclk));
	jdff dff_B_BJbGIzEY5_1(.din(w_dff_B_KtEtKJji2_1),.dout(w_dff_B_BJbGIzEY5_1),.clk(gclk));
	jdff dff_B_xxdvb4ew8_1(.din(w_dff_B_BJbGIzEY5_1),.dout(w_dff_B_xxdvb4ew8_1),.clk(gclk));
	jdff dff_B_JYWRbbI97_1(.din(w_dff_B_xxdvb4ew8_1),.dout(w_dff_B_JYWRbbI97_1),.clk(gclk));
	jdff dff_B_GYlf9tmp0_0(.din(n1150),.dout(w_dff_B_GYlf9tmp0_0),.clk(gclk));
	jdff dff_B_QaQDSJFo4_0(.din(w_dff_B_GYlf9tmp0_0),.dout(w_dff_B_QaQDSJFo4_0),.clk(gclk));
	jdff dff_B_T0qrOHgi4_0(.din(w_dff_B_QaQDSJFo4_0),.dout(w_dff_B_T0qrOHgi4_0),.clk(gclk));
	jdff dff_B_IlgMwBIO6_0(.din(w_dff_B_T0qrOHgi4_0),.dout(w_dff_B_IlgMwBIO6_0),.clk(gclk));
	jdff dff_B_YAgN0rkF8_0(.din(w_dff_B_IlgMwBIO6_0),.dout(w_dff_B_YAgN0rkF8_0),.clk(gclk));
	jdff dff_B_L4m7v8lK9_0(.din(w_dff_B_YAgN0rkF8_0),.dout(w_dff_B_L4m7v8lK9_0),.clk(gclk));
	jdff dff_B_iOqssW0V2_0(.din(w_dff_B_L4m7v8lK9_0),.dout(w_dff_B_iOqssW0V2_0),.clk(gclk));
	jdff dff_B_D5ri3bxJ3_0(.din(w_dff_B_iOqssW0V2_0),.dout(w_dff_B_D5ri3bxJ3_0),.clk(gclk));
	jdff dff_B_pXI7YmXC2_0(.din(w_dff_B_D5ri3bxJ3_0),.dout(w_dff_B_pXI7YmXC2_0),.clk(gclk));
	jdff dff_B_wzyJFi5n6_0(.din(w_dff_B_pXI7YmXC2_0),.dout(w_dff_B_wzyJFi5n6_0),.clk(gclk));
	jdff dff_B_X3rX3h1N3_0(.din(w_dff_B_wzyJFi5n6_0),.dout(w_dff_B_X3rX3h1N3_0),.clk(gclk));
	jdff dff_B_WBQU4sIr8_0(.din(w_dff_B_X3rX3h1N3_0),.dout(w_dff_B_WBQU4sIr8_0),.clk(gclk));
	jdff dff_B_i1xdznr45_0(.din(n1146),.dout(w_dff_B_i1xdznr45_0),.clk(gclk));
	jdff dff_A_PIcgelcc1_0(.dout(w_n1007_3[0]),.din(w_dff_A_PIcgelcc1_0),.clk(gclk));
	jdff dff_A_NwuXZuxK5_1(.dout(w_n1007_3[1]),.din(w_dff_A_NwuXZuxK5_1),.clk(gclk));
	jdff dff_A_vHywm2w90_1(.dout(w_dff_A_NwuXZuxK5_1),.din(w_dff_A_vHywm2w90_1),.clk(gclk));
	jdff dff_A_iE53cuUi2_1(.dout(w_dff_A_vHywm2w90_1),.din(w_dff_A_iE53cuUi2_1),.clk(gclk));
	jdff dff_A_KRGFQMvu0_1(.dout(w_dff_A_iE53cuUi2_1),.din(w_dff_A_KRGFQMvu0_1),.clk(gclk));
	jdff dff_A_Q5q0762m9_1(.dout(w_dff_A_KRGFQMvu0_1),.din(w_dff_A_Q5q0762m9_1),.clk(gclk));
	jdff dff_A_9gFfPl351_1(.dout(w_dff_A_Q5q0762m9_1),.din(w_dff_A_9gFfPl351_1),.clk(gclk));
	jdff dff_B_Rn4WCP9Z0_1(.din(n762),.dout(w_dff_B_Rn4WCP9Z0_1),.clk(gclk));
	jdff dff_B_geuXO1e88_1(.din(w_dff_B_Rn4WCP9Z0_1),.dout(w_dff_B_geuXO1e88_1),.clk(gclk));
	jdff dff_B_OtJa7mWN0_1(.din(w_dff_B_geuXO1e88_1),.dout(w_dff_B_OtJa7mWN0_1),.clk(gclk));
	jdff dff_B_6JElo9hD4_1(.din(w_dff_B_OtJa7mWN0_1),.dout(w_dff_B_6JElo9hD4_1),.clk(gclk));
	jdff dff_B_6eKDnRiu8_1(.din(w_dff_B_6JElo9hD4_1),.dout(w_dff_B_6eKDnRiu8_1),.clk(gclk));
	jdff dff_B_LZtyHhp22_1(.din(w_dff_B_6eKDnRiu8_1),.dout(w_dff_B_LZtyHhp22_1),.clk(gclk));
	jdff dff_B_b0KXPMBY7_1(.din(w_dff_B_LZtyHhp22_1),.dout(w_dff_B_b0KXPMBY7_1),.clk(gclk));
	jdff dff_B_1h6ymRVb5_1(.din(w_dff_B_b0KXPMBY7_1),.dout(w_dff_B_1h6ymRVb5_1),.clk(gclk));
	jdff dff_B_Aj3s74Qr4_0(.din(n773),.dout(w_dff_B_Aj3s74Qr4_0),.clk(gclk));
	jdff dff_B_4CZvdFqP8_0(.din(w_dff_B_Aj3s74Qr4_0),.dout(w_dff_B_4CZvdFqP8_0),.clk(gclk));
	jdff dff_B_zV1xcR2g4_0(.din(w_dff_B_4CZvdFqP8_0),.dout(w_dff_B_zV1xcR2g4_0),.clk(gclk));
	jdff dff_B_gT4N4AbX2_0(.din(w_dff_B_zV1xcR2g4_0),.dout(w_dff_B_gT4N4AbX2_0),.clk(gclk));
	jdff dff_B_EI8qdsfc3_0(.din(n769),.dout(w_dff_B_EI8qdsfc3_0),.clk(gclk));
	jdff dff_B_88nphrFP2_0(.din(w_dff_B_EI8qdsfc3_0),.dout(w_dff_B_88nphrFP2_0),.clk(gclk));
	jdff dff_B_8s4KVCS63_0(.din(w_dff_B_88nphrFP2_0),.dout(w_dff_B_8s4KVCS63_0),.clk(gclk));
	jdff dff_B_mqpqi7DM5_0(.din(w_dff_B_8s4KVCS63_0),.dout(w_dff_B_mqpqi7DM5_0),.clk(gclk));
	jdff dff_A_394idVPZ4_1(.dout(w_G137_7[1]),.din(w_dff_A_394idVPZ4_1),.clk(gclk));
	jdff dff_A_kjJ1EEFO9_1(.dout(w_dff_A_394idVPZ4_1),.din(w_dff_A_kjJ1EEFO9_1),.clk(gclk));
	jdff dff_A_JjLejf5U9_1(.dout(w_dff_A_kjJ1EEFO9_1),.din(w_dff_A_JjLejf5U9_1),.clk(gclk));
	jdff dff_A_0JDJpoad9_1(.dout(w_dff_A_JjLejf5U9_1),.din(w_dff_A_0JDJpoad9_1),.clk(gclk));
	jdff dff_A_r8xWbjbI8_2(.dout(w_G137_7[2]),.din(w_dff_A_r8xWbjbI8_2),.clk(gclk));
	jdff dff_A_My38uOGv8_0(.dout(w_G137_2[0]),.din(w_dff_A_My38uOGv8_0),.clk(gclk));
	jdff dff_A_dH68NgwT8_0(.dout(w_dff_A_My38uOGv8_0),.din(w_dff_A_dH68NgwT8_0),.clk(gclk));
	jdff dff_A_FA9GbpNf2_1(.dout(w_G137_2[1]),.din(w_dff_A_FA9GbpNf2_1),.clk(gclk));
	jdff dff_A_Exb9jyy65_1(.dout(w_dff_A_FA9GbpNf2_1),.din(w_dff_A_Exb9jyy65_1),.clk(gclk));
	jdff dff_B_lb1qM44B4_0(.din(n1159),.dout(w_dff_B_lb1qM44B4_0),.clk(gclk));
	jdff dff_B_Ryn9RK0i8_0(.din(w_dff_B_lb1qM44B4_0),.dout(w_dff_B_Ryn9RK0i8_0),.clk(gclk));
	jdff dff_B_UJqb6P6u9_0(.din(w_dff_B_Ryn9RK0i8_0),.dout(w_dff_B_UJqb6P6u9_0),.clk(gclk));
	jdff dff_B_WmlnOgTz8_0(.din(w_dff_B_UJqb6P6u9_0),.dout(w_dff_B_WmlnOgTz8_0),.clk(gclk));
	jdff dff_B_8wM9d6928_0(.din(w_dff_B_WmlnOgTz8_0),.dout(w_dff_B_8wM9d6928_0),.clk(gclk));
	jdff dff_B_VHvu3BTi2_0(.din(w_dff_B_8wM9d6928_0),.dout(w_dff_B_VHvu3BTi2_0),.clk(gclk));
	jdff dff_B_gVy0gIJY5_0(.din(w_dff_B_VHvu3BTi2_0),.dout(w_dff_B_gVy0gIJY5_0),.clk(gclk));
	jdff dff_B_DTqzfii80_0(.din(w_dff_B_gVy0gIJY5_0),.dout(w_dff_B_DTqzfii80_0),.clk(gclk));
	jdff dff_B_bitBGjAr2_0(.din(w_dff_B_DTqzfii80_0),.dout(w_dff_B_bitBGjAr2_0),.clk(gclk));
	jdff dff_B_EvUtjhT30_0(.din(w_dff_B_bitBGjAr2_0),.dout(w_dff_B_EvUtjhT30_0),.clk(gclk));
	jdff dff_B_BFFTF91n5_0(.din(w_dff_B_EvUtjhT30_0),.dout(w_dff_B_BFFTF91n5_0),.clk(gclk));
	jdff dff_B_6dxuLh870_0(.din(w_dff_B_BFFTF91n5_0),.dout(w_dff_B_6dxuLh870_0),.clk(gclk));
	jdff dff_B_3qN4cbYf0_1(.din(n1153),.dout(w_dff_B_3qN4cbYf0_1),.clk(gclk));
	jdff dff_B_XBy4Vuwp3_1(.din(n843),.dout(w_dff_B_XBy4Vuwp3_1),.clk(gclk));
	jdff dff_B_QnOTtXCy1_1(.din(w_dff_B_XBy4Vuwp3_1),.dout(w_dff_B_QnOTtXCy1_1),.clk(gclk));
	jdff dff_B_ApErmMJk6_1(.din(w_dff_B_QnOTtXCy1_1),.dout(w_dff_B_ApErmMJk6_1),.clk(gclk));
	jdff dff_B_nEVJ6oVV3_1(.din(w_dff_B_ApErmMJk6_1),.dout(w_dff_B_nEVJ6oVV3_1),.clk(gclk));
	jdff dff_B_QLOQPG8i0_1(.din(w_dff_B_nEVJ6oVV3_1),.dout(w_dff_B_QLOQPG8i0_1),.clk(gclk));
	jdff dff_B_9pOpdXtw3_1(.din(w_dff_B_QLOQPG8i0_1),.dout(w_dff_B_9pOpdXtw3_1),.clk(gclk));
	jdff dff_B_ZeJDghyp9_1(.din(w_dff_B_9pOpdXtw3_1),.dout(w_dff_B_ZeJDghyp9_1),.clk(gclk));
	jdff dff_B_tgDCCe2M3_1(.din(n844),.dout(w_dff_B_tgDCCe2M3_1),.clk(gclk));
	jdff dff_B_beOOIN0R0_1(.din(w_dff_B_tgDCCe2M3_1),.dout(w_dff_B_beOOIN0R0_1),.clk(gclk));
	jdff dff_B_s7MYspbX0_1(.din(w_dff_B_beOOIN0R0_1),.dout(w_dff_B_s7MYspbX0_1),.clk(gclk));
	jdff dff_B_5z9KsX4z9_1(.din(w_dff_B_s7MYspbX0_1),.dout(w_dff_B_5z9KsX4z9_1),.clk(gclk));
	jdff dff_A_JcH5yEVp0_0(.dout(w_n847_0[0]),.din(w_dff_A_JcH5yEVp0_0),.clk(gclk));
	jdff dff_A_YKVLwzCi9_0(.dout(w_dff_A_JcH5yEVp0_0),.din(w_dff_A_YKVLwzCi9_0),.clk(gclk));
	jdff dff_A_Qc9LS6Lr6_0(.dout(w_dff_A_YKVLwzCi9_0),.din(w_dff_A_Qc9LS6Lr6_0),.clk(gclk));
	jdff dff_A_u255Ju3h1_0(.dout(w_dff_A_Qc9LS6Lr6_0),.din(w_dff_A_u255Ju3h1_0),.clk(gclk));
	jdff dff_A_QOxkxB1I3_0(.dout(w_dff_A_u255Ju3h1_0),.din(w_dff_A_QOxkxB1I3_0),.clk(gclk));
	jdff dff_B_DaxcvxvW4_0(.din(n1168),.dout(w_dff_B_DaxcvxvW4_0),.clk(gclk));
	jdff dff_B_QEMgVGea6_0(.din(w_dff_B_DaxcvxvW4_0),.dout(w_dff_B_QEMgVGea6_0),.clk(gclk));
	jdff dff_B_loUNumSK5_0(.din(w_dff_B_QEMgVGea6_0),.dout(w_dff_B_loUNumSK5_0),.clk(gclk));
	jdff dff_B_ZzPWaRZK7_0(.din(w_dff_B_loUNumSK5_0),.dout(w_dff_B_ZzPWaRZK7_0),.clk(gclk));
	jdff dff_B_G3mwbcmp7_0(.din(w_dff_B_ZzPWaRZK7_0),.dout(w_dff_B_G3mwbcmp7_0),.clk(gclk));
	jdff dff_B_Q5f7ILYP8_0(.din(w_dff_B_G3mwbcmp7_0),.dout(w_dff_B_Q5f7ILYP8_0),.clk(gclk));
	jdff dff_B_HQhAEU7Z2_0(.din(w_dff_B_Q5f7ILYP8_0),.dout(w_dff_B_HQhAEU7Z2_0),.clk(gclk));
	jdff dff_B_Ux9JRKrS5_0(.din(w_dff_B_HQhAEU7Z2_0),.dout(w_dff_B_Ux9JRKrS5_0),.clk(gclk));
	jdff dff_B_WsIEIQma6_0(.din(w_dff_B_Ux9JRKrS5_0),.dout(w_dff_B_WsIEIQma6_0),.clk(gclk));
	jdff dff_B_OdClI2C52_0(.din(w_dff_B_WsIEIQma6_0),.dout(w_dff_B_OdClI2C52_0),.clk(gclk));
	jdff dff_B_abBQ0BRH3_0(.din(w_dff_B_OdClI2C52_0),.dout(w_dff_B_abBQ0BRH3_0),.clk(gclk));
	jdff dff_B_wX6OIxDw5_0(.din(w_dff_B_abBQ0BRH3_0),.dout(w_dff_B_wX6OIxDw5_0),.clk(gclk));
	jdff dff_B_1oUwOJya1_0(.din(w_dff_B_wX6OIxDw5_0),.dout(w_dff_B_1oUwOJya1_0),.clk(gclk));
	jdff dff_A_ANLfMAZe9_0(.dout(w_n1008_3[0]),.din(w_dff_A_ANLfMAZe9_0),.clk(gclk));
	jdff dff_A_PHmYnQ426_0(.dout(w_dff_A_ANLfMAZe9_0),.din(w_dff_A_PHmYnQ426_0),.clk(gclk));
	jdff dff_A_CNn93fsX2_1(.dout(w_n1008_3[1]),.din(w_dff_A_CNn93fsX2_1),.clk(gclk));
	jdff dff_B_MPOcCkTp6_1(.din(n834),.dout(w_dff_B_MPOcCkTp6_1),.clk(gclk));
	jdff dff_B_2fYVIv2c2_1(.din(w_dff_B_MPOcCkTp6_1),.dout(w_dff_B_2fYVIv2c2_1),.clk(gclk));
	jdff dff_B_cDVfxSgn1_1(.din(w_dff_B_2fYVIv2c2_1),.dout(w_dff_B_cDVfxSgn1_1),.clk(gclk));
	jdff dff_B_8rzkGeZV9_1(.din(w_dff_B_cDVfxSgn1_1),.dout(w_dff_B_8rzkGeZV9_1),.clk(gclk));
	jdff dff_B_tQ91bYHC3_1(.din(w_dff_B_8rzkGeZV9_1),.dout(w_dff_B_tQ91bYHC3_1),.clk(gclk));
	jdff dff_B_cG1SKwuA2_1(.din(w_dff_B_tQ91bYHC3_1),.dout(w_dff_B_cG1SKwuA2_1),.clk(gclk));
	jdff dff_B_QKEJEcGo1_1(.din(w_dff_B_cG1SKwuA2_1),.dout(w_dff_B_QKEJEcGo1_1),.clk(gclk));
	jdff dff_B_FUjWWtXH5_1(.din(w_dff_B_QKEJEcGo1_1),.dout(w_dff_B_FUjWWtXH5_1),.clk(gclk));
	jdff dff_B_b7l7TUX85_1(.din(w_dff_B_FUjWWtXH5_1),.dout(w_dff_B_b7l7TUX85_1),.clk(gclk));
	jdff dff_B_hwfvK0fe6_0(.din(n839),.dout(w_dff_B_hwfvK0fe6_0),.clk(gclk));
	jdff dff_B_w0DLYHA09_0(.din(w_dff_B_hwfvK0fe6_0),.dout(w_dff_B_w0DLYHA09_0),.clk(gclk));
	jdff dff_B_1vKv8XKJ5_0(.din(w_dff_B_w0DLYHA09_0),.dout(w_dff_B_1vKv8XKJ5_0),.clk(gclk));
	jdff dff_B_SVYZF8wu0_0(.din(w_dff_B_1vKv8XKJ5_0),.dout(w_dff_B_SVYZF8wu0_0),.clk(gclk));
	jdff dff_B_hN8odqwb6_0(.din(w_dff_B_SVYZF8wu0_0),.dout(w_dff_B_hN8odqwb6_0),.clk(gclk));
	jdff dff_B_2YSxb2fz8_0(.din(w_dff_B_hN8odqwb6_0),.dout(w_dff_B_2YSxb2fz8_0),.clk(gclk));
	jdff dff_A_JzCI1fDH0_0(.dout(w_n836_0[0]),.din(w_dff_A_JzCI1fDH0_0),.clk(gclk));
	jdff dff_A_1MQZQAK70_0(.dout(w_dff_A_JzCI1fDH0_0),.din(w_dff_A_1MQZQAK70_0),.clk(gclk));
	jdff dff_A_G6xBS8gp1_0(.dout(w_dff_A_1MQZQAK70_0),.din(w_dff_A_G6xBS8gp1_0),.clk(gclk));
	jdff dff_A_LjcwLS5f1_0(.dout(w_dff_A_G6xBS8gp1_0),.din(w_dff_A_LjcwLS5f1_0),.clk(gclk));
	jdff dff_A_qib1nwvv2_0(.dout(w_dff_A_LjcwLS5f1_0),.din(w_dff_A_qib1nwvv2_0),.clk(gclk));
	jdff dff_A_0VV33D722_0(.dout(w_dff_A_qib1nwvv2_0),.din(w_dff_A_0VV33D722_0),.clk(gclk));
	jdff dff_A_bKVOydk43_0(.dout(w_dff_A_0VV33D722_0),.din(w_dff_A_bKVOydk43_0),.clk(gclk));
	jdff dff_B_v1bO5mI78_1(.din(n1173),.dout(w_dff_B_v1bO5mI78_1),.clk(gclk));
	jdff dff_B_9J5Yro5B3_1(.din(w_dff_B_v1bO5mI78_1),.dout(w_dff_B_9J5Yro5B3_1),.clk(gclk));
	jdff dff_B_ieXzWPEE4_1(.din(w_dff_B_9J5Yro5B3_1),.dout(w_dff_B_ieXzWPEE4_1),.clk(gclk));
	jdff dff_B_wzNgKGVX6_1(.din(w_dff_B_ieXzWPEE4_1),.dout(w_dff_B_wzNgKGVX6_1),.clk(gclk));
	jdff dff_B_ne0AMC961_1(.din(w_dff_B_wzNgKGVX6_1),.dout(w_dff_B_ne0AMC961_1),.clk(gclk));
	jdff dff_B_4pA0ScO27_1(.din(w_dff_B_ne0AMC961_1),.dout(w_dff_B_4pA0ScO27_1),.clk(gclk));
	jdff dff_B_aFAcwiUP0_1(.din(w_dff_B_4pA0ScO27_1),.dout(w_dff_B_aFAcwiUP0_1),.clk(gclk));
	jdff dff_B_LCvqKDej3_1(.din(w_dff_B_aFAcwiUP0_1),.dout(w_dff_B_LCvqKDej3_1),.clk(gclk));
	jdff dff_B_Zx0NJew23_1(.din(w_dff_B_LCvqKDej3_1),.dout(w_dff_B_Zx0NJew23_1),.clk(gclk));
	jdff dff_B_SzOYvOBJ6_1(.din(w_dff_B_Zx0NJew23_1),.dout(w_dff_B_SzOYvOBJ6_1),.clk(gclk));
	jdff dff_B_qip4DymN3_1(.din(w_dff_B_SzOYvOBJ6_1),.dout(w_dff_B_qip4DymN3_1),.clk(gclk));
	jdff dff_B_8DhUfWxj1_1(.din(w_dff_B_qip4DymN3_1),.dout(w_dff_B_8DhUfWxj1_1),.clk(gclk));
	jdff dff_B_C5ATztjV6_1(.din(w_dff_B_8DhUfWxj1_1),.dout(w_dff_B_C5ATztjV6_1),.clk(gclk));
	jdff dff_B_7xJhnG052_1(.din(w_dff_B_C5ATztjV6_1),.dout(w_dff_B_7xJhnG052_1),.clk(gclk));
	jdff dff_B_ZPgOoydR5_1(.din(w_dff_B_7xJhnG052_1),.dout(w_dff_B_ZPgOoydR5_1),.clk(gclk));
	jdff dff_B_V7or1dHo8_1(.din(w_dff_B_ZPgOoydR5_1),.dout(w_dff_B_V7or1dHo8_1),.clk(gclk));
	jdff dff_B_DMam5gA08_1(.din(w_dff_B_V7or1dHo8_1),.dout(w_dff_B_DMam5gA08_1),.clk(gclk));
	jdff dff_B_1JZQHkVQ8_1(.din(w_dff_B_DMam5gA08_1),.dout(w_dff_B_1JZQHkVQ8_1),.clk(gclk));
	jdff dff_B_m9XErvMi0_1(.din(n1182),.dout(w_dff_B_m9XErvMi0_1),.clk(gclk));
	jdff dff_B_MMnb1Wq13_1(.din(w_dff_B_m9XErvMi0_1),.dout(w_dff_B_MMnb1Wq13_1),.clk(gclk));
	jdff dff_B_WTKqezxX2_1(.din(w_dff_B_MMnb1Wq13_1),.dout(w_dff_B_WTKqezxX2_1),.clk(gclk));
	jdff dff_B_KEnsGmEz5_1(.din(w_dff_B_WTKqezxX2_1),.dout(w_dff_B_KEnsGmEz5_1),.clk(gclk));
	jdff dff_B_qWpozdUN2_1(.din(w_dff_B_KEnsGmEz5_1),.dout(w_dff_B_qWpozdUN2_1),.clk(gclk));
	jdff dff_B_emT5n7H64_1(.din(w_dff_B_qWpozdUN2_1),.dout(w_dff_B_emT5n7H64_1),.clk(gclk));
	jdff dff_B_CFBEcHnW3_1(.din(w_dff_B_emT5n7H64_1),.dout(w_dff_B_CFBEcHnW3_1),.clk(gclk));
	jdff dff_B_uZlHwleW0_1(.din(w_dff_B_CFBEcHnW3_1),.dout(w_dff_B_uZlHwleW0_1),.clk(gclk));
	jdff dff_B_cN5UFef44_1(.din(w_dff_B_uZlHwleW0_1),.dout(w_dff_B_cN5UFef44_1),.clk(gclk));
	jdff dff_B_3gDUGkFP6_1(.din(w_dff_B_cN5UFef44_1),.dout(w_dff_B_3gDUGkFP6_1),.clk(gclk));
	jdff dff_B_GeuIZe7S9_0(.din(n1185),.dout(w_dff_B_GeuIZe7S9_0),.clk(gclk));
	jdff dff_B_SKf02YKw3_0(.din(w_dff_B_GeuIZe7S9_0),.dout(w_dff_B_SKf02YKw3_0),.clk(gclk));
	jdff dff_B_gHwkZVsd2_0(.din(w_dff_B_SKf02YKw3_0),.dout(w_dff_B_gHwkZVsd2_0),.clk(gclk));
	jdff dff_B_EBkLG0Sg0_0(.din(w_dff_B_gHwkZVsd2_0),.dout(w_dff_B_EBkLG0Sg0_0),.clk(gclk));
	jdff dff_B_w1UVBfmU1_0(.din(w_dff_B_EBkLG0Sg0_0),.dout(w_dff_B_w1UVBfmU1_0),.clk(gclk));
	jdff dff_B_xnvLp0aB6_0(.din(w_dff_B_w1UVBfmU1_0),.dout(w_dff_B_xnvLp0aB6_0),.clk(gclk));
	jdff dff_B_b2vb30T19_0(.din(w_dff_B_xnvLp0aB6_0),.dout(w_dff_B_b2vb30T19_0),.clk(gclk));
	jdff dff_B_KO2DtA1o8_0(.din(w_dff_B_b2vb30T19_0),.dout(w_dff_B_KO2DtA1o8_0),.clk(gclk));
	jdff dff_B_rzXwiNao3_0(.din(w_dff_B_KO2DtA1o8_0),.dout(w_dff_B_rzXwiNao3_0),.clk(gclk));
	jdff dff_B_aimPF6Yl5_0(.din(w_dff_B_rzXwiNao3_0),.dout(w_dff_B_aimPF6Yl5_0),.clk(gclk));
	jdff dff_B_fs01Md6z6_0(.din(w_dff_B_aimPF6Yl5_0),.dout(w_dff_B_fs01Md6z6_0),.clk(gclk));
	jdff dff_B_BzKjiF2z6_0(.din(w_dff_B_fs01Md6z6_0),.dout(w_dff_B_BzKjiF2z6_0),.clk(gclk));
	jdff dff_B_tCHeFHea9_0(.din(w_dff_B_BzKjiF2z6_0),.dout(w_dff_B_tCHeFHea9_0),.clk(gclk));
	jdff dff_B_45hcvCJ00_0(.din(w_dff_B_tCHeFHea9_0),.dout(w_dff_B_45hcvCJ00_0),.clk(gclk));
	jdff dff_B_7p2bQJV08_0(.din(w_dff_B_45hcvCJ00_0),.dout(w_dff_B_7p2bQJV08_0),.clk(gclk));
	jdff dff_B_FSaM279M7_0(.din(w_dff_B_7p2bQJV08_0),.dout(w_dff_B_FSaM279M7_0),.clk(gclk));
	jdff dff_B_5ZDP9ftx9_1(.din(n1175),.dout(w_dff_B_5ZDP9ftx9_1),.clk(gclk));
	jdff dff_B_0fADwkXw9_1(.din(w_dff_B_5ZDP9ftx9_1),.dout(w_dff_B_0fADwkXw9_1),.clk(gclk));
	jdff dff_B_g6dH3Znt0_1(.din(w_dff_B_0fADwkXw9_1),.dout(w_dff_B_g6dH3Znt0_1),.clk(gclk));
	jdff dff_B_lSSq5HWT9_1(.din(n1176),.dout(w_dff_B_lSSq5HWT9_1),.clk(gclk));
	jdff dff_B_4GYBegJO0_1(.din(w_dff_B_lSSq5HWT9_1),.dout(w_dff_B_4GYBegJO0_1),.clk(gclk));
	jdff dff_B_FuCfEokb2_1(.din(w_dff_B_4GYBegJO0_1),.dout(w_dff_B_FuCfEokb2_1),.clk(gclk));
	jdff dff_B_MOZGd3nc5_1(.din(w_dff_B_FuCfEokb2_1),.dout(w_dff_B_MOZGd3nc5_1),.clk(gclk));
	jdff dff_B_KqV8IN1E0_1(.din(w_dff_B_MOZGd3nc5_1),.dout(w_dff_B_KqV8IN1E0_1),.clk(gclk));
	jdff dff_B_c9rVHgUN5_1(.din(w_dff_B_KqV8IN1E0_1),.dout(w_dff_B_c9rVHgUN5_1),.clk(gclk));
	jdff dff_A_xbbYYgWi3_0(.dout(w_n1177_0[0]),.din(w_dff_A_xbbYYgWi3_0),.clk(gclk));
	jdff dff_A_rsMdykz66_0(.dout(w_dff_A_xbbYYgWi3_0),.din(w_dff_A_rsMdykz66_0),.clk(gclk));
	jdff dff_A_SfEJBOaA0_0(.dout(w_dff_A_rsMdykz66_0),.din(w_dff_A_SfEJBOaA0_0),.clk(gclk));
	jdff dff_A_Q15o28yw6_0(.dout(w_dff_A_SfEJBOaA0_0),.din(w_dff_A_Q15o28yw6_0),.clk(gclk));
	jdff dff_A_TGo1IMHy8_0(.dout(w_dff_A_Q15o28yw6_0),.din(w_dff_A_TGo1IMHy8_0),.clk(gclk));
	jdff dff_A_4UL1BwAG7_0(.dout(w_dff_A_TGo1IMHy8_0),.din(w_dff_A_4UL1BwAG7_0),.clk(gclk));
	jdff dff_A_iu4QtZnr1_0(.dout(w_dff_A_4UL1BwAG7_0),.din(w_dff_A_iu4QtZnr1_0),.clk(gclk));
	jdff dff_A_pPSMOaFR4_0(.dout(w_dff_A_iu4QtZnr1_0),.din(w_dff_A_pPSMOaFR4_0),.clk(gclk));
	jdff dff_A_GK6LHLhs1_0(.dout(w_dff_A_pPSMOaFR4_0),.din(w_dff_A_GK6LHLhs1_0),.clk(gclk));
	jdff dff_A_p0MWBDBZ0_0(.dout(w_dff_A_GK6LHLhs1_0),.din(w_dff_A_p0MWBDBZ0_0),.clk(gclk));
	jdff dff_A_jcFJtrsX8_0(.dout(w_dff_A_p0MWBDBZ0_0),.din(w_dff_A_jcFJtrsX8_0),.clk(gclk));
	jdff dff_B_FT0M63c13_2(.din(n1177),.dout(w_dff_B_FT0M63c13_2),.clk(gclk));
	jdff dff_B_LmrubnDT9_2(.din(w_dff_B_FT0M63c13_2),.dout(w_dff_B_LmrubnDT9_2),.clk(gclk));
	jdff dff_B_XrQQAS405_2(.din(w_dff_B_LmrubnDT9_2),.dout(w_dff_B_XrQQAS405_2),.clk(gclk));
	jdff dff_B_MH6DOu3F7_2(.din(w_dff_B_XrQQAS405_2),.dout(w_dff_B_MH6DOu3F7_2),.clk(gclk));
	jdff dff_B_xmNcrysp8_2(.din(w_dff_B_MH6DOu3F7_2),.dout(w_dff_B_xmNcrysp8_2),.clk(gclk));
	jdff dff_A_c0gJlOqo4_0(.dout(w_n1179_0[0]),.din(w_dff_A_c0gJlOqo4_0),.clk(gclk));
	jdff dff_A_PnqvxPzc0_0(.dout(w_dff_A_c0gJlOqo4_0),.din(w_dff_A_PnqvxPzc0_0),.clk(gclk));
	jdff dff_A_7B7hsHaq2_0(.dout(w_dff_A_PnqvxPzc0_0),.din(w_dff_A_7B7hsHaq2_0),.clk(gclk));
	jdff dff_A_VBhZXm0p8_0(.dout(w_dff_A_7B7hsHaq2_0),.din(w_dff_A_VBhZXm0p8_0),.clk(gclk));
	jdff dff_A_miGwPmJY7_0(.dout(w_dff_A_VBhZXm0p8_0),.din(w_dff_A_miGwPmJY7_0),.clk(gclk));
	jdff dff_A_2KYoFuJn0_0(.dout(w_dff_A_miGwPmJY7_0),.din(w_dff_A_2KYoFuJn0_0),.clk(gclk));
	jdff dff_A_5wGTqp6I1_0(.dout(w_dff_A_2KYoFuJn0_0),.din(w_dff_A_5wGTqp6I1_0),.clk(gclk));
	jdff dff_A_dmkHZ2qv4_0(.dout(w_dff_A_5wGTqp6I1_0),.din(w_dff_A_dmkHZ2qv4_0),.clk(gclk));
	jdff dff_A_oiBMTlRc5_0(.dout(w_dff_A_dmkHZ2qv4_0),.din(w_dff_A_oiBMTlRc5_0),.clk(gclk));
	jdff dff_A_jpdcUoa39_0(.dout(w_dff_A_oiBMTlRc5_0),.din(w_dff_A_jpdcUoa39_0),.clk(gclk));
	jdff dff_A_cinRNd2W2_0(.dout(w_dff_A_jpdcUoa39_0),.din(w_dff_A_cinRNd2W2_0),.clk(gclk));
	jdff dff_B_hCGCbvbn5_1(.din(G132),.dout(w_dff_B_hCGCbvbn5_1),.clk(gclk));
	jdff dff_B_HdAI6Y7T4_1(.din(w_dff_B_hCGCbvbn5_1),.dout(w_dff_B_HdAI6Y7T4_1),.clk(gclk));
	jdff dff_B_2YvGSUPm0_1(.din(w_dff_B_HdAI6Y7T4_1),.dout(w_dff_B_2YvGSUPm0_1),.clk(gclk));
	jdff dff_B_XYwVKQL19_1(.din(w_dff_B_2YvGSUPm0_1),.dout(w_dff_B_XYwVKQL19_1),.clk(gclk));
	jdff dff_B_DKZt5hg95_1(.din(n1223),.dout(w_dff_B_DKZt5hg95_1),.clk(gclk));
	jdff dff_B_5F4cHltd1_0(.din(n1227),.dout(w_dff_B_5F4cHltd1_0),.clk(gclk));
	jdff dff_B_k4bFRORr8_0(.din(w_dff_B_5F4cHltd1_0),.dout(w_dff_B_k4bFRORr8_0),.clk(gclk));
	jdff dff_B_HLQ2XLlh4_0(.din(w_dff_B_k4bFRORr8_0),.dout(w_dff_B_HLQ2XLlh4_0),.clk(gclk));
	jdff dff_B_uXwQUzK48_0(.din(w_dff_B_HLQ2XLlh4_0),.dout(w_dff_B_uXwQUzK48_0),.clk(gclk));
	jdff dff_B_BzKGYPfc6_0(.din(n1226),.dout(w_dff_B_BzKGYPfc6_0),.clk(gclk));
	jdff dff_A_L8qNNPTz3_0(.dout(w_G559_0[0]),.din(w_dff_A_L8qNNPTz3_0),.clk(gclk));
	jdff dff_A_XYykHfUK1_0(.dout(w_dff_A_L8qNNPTz3_0),.din(w_dff_A_XYykHfUK1_0),.clk(gclk));
	jdff dff_B_GLcQe6Os9_1(.din(n916),.dout(w_dff_B_GLcQe6Os9_1),.clk(gclk));
	jdff dff_B_IjWP77AJ0_1(.din(n917),.dout(w_dff_B_IjWP77AJ0_1),.clk(gclk));
	jdff dff_B_YwVVYjAq7_1(.din(n1263),.dout(w_dff_B_YwVVYjAq7_1),.clk(gclk));
	jdff dff_B_1lWxf8dv3_1(.din(w_dff_B_YwVVYjAq7_1),.dout(w_dff_B_1lWxf8dv3_1),.clk(gclk));
	jdff dff_B_rZrAkUxI5_1(.din(w_dff_B_1lWxf8dv3_1),.dout(w_dff_B_rZrAkUxI5_1),.clk(gclk));
	jdff dff_B_3tDQzPvF4_1(.din(w_dff_B_rZrAkUxI5_1),.dout(w_dff_B_3tDQzPvF4_1),.clk(gclk));
	jdff dff_B_n66KbUP66_1(.din(w_dff_B_3tDQzPvF4_1),.dout(w_dff_B_n66KbUP66_1),.clk(gclk));
	jdff dff_B_NkSbuJrO0_1(.din(w_dff_B_n66KbUP66_1),.dout(w_dff_B_NkSbuJrO0_1),.clk(gclk));
	jdff dff_B_UVobcjTu0_1(.din(w_dff_B_NkSbuJrO0_1),.dout(w_dff_B_UVobcjTu0_1),.clk(gclk));
	jdff dff_B_fPO83u4t8_1(.din(w_dff_B_UVobcjTu0_1),.dout(w_dff_B_fPO83u4t8_1),.clk(gclk));
	jdff dff_B_QbdKbOSC0_1(.din(w_dff_B_fPO83u4t8_1),.dout(w_dff_B_QbdKbOSC0_1),.clk(gclk));
	jdff dff_B_gVUlk6Jo7_1(.din(w_dff_B_QbdKbOSC0_1),.dout(w_dff_B_gVUlk6Jo7_1),.clk(gclk));
	jdff dff_B_0lZz5DDD5_1(.din(w_dff_B_gVUlk6Jo7_1),.dout(w_dff_B_0lZz5DDD5_1),.clk(gclk));
	jdff dff_B_L30WRLTa1_1(.din(w_dff_B_0lZz5DDD5_1),.dout(w_dff_B_L30WRLTa1_1),.clk(gclk));
	jdff dff_B_A94QpvrG7_1(.din(w_dff_B_L30WRLTa1_1),.dout(w_dff_B_A94QpvrG7_1),.clk(gclk));
	jdff dff_B_N4D3wLzj6_1(.din(w_dff_B_A94QpvrG7_1),.dout(w_dff_B_N4D3wLzj6_1),.clk(gclk));
	jdff dff_B_7UY5i46H8_1(.din(w_dff_B_N4D3wLzj6_1),.dout(w_dff_B_7UY5i46H8_1),.clk(gclk));
	jdff dff_B_fMhhPfwW0_1(.din(w_dff_B_7UY5i46H8_1),.dout(w_dff_B_fMhhPfwW0_1),.clk(gclk));
	jdff dff_B_IlR4EslL7_1(.din(w_dff_B_fMhhPfwW0_1),.dout(w_dff_B_IlR4EslL7_1),.clk(gclk));
	jdff dff_B_DrAd6EK05_1(.din(w_dff_B_IlR4EslL7_1),.dout(w_dff_B_DrAd6EK05_1),.clk(gclk));
	jdff dff_B_9knjpEj62_1(.din(w_dff_B_DrAd6EK05_1),.dout(w_dff_B_9knjpEj62_1),.clk(gclk));
	jdff dff_B_Qz8uHCUV4_0(.din(n1276),.dout(w_dff_B_Qz8uHCUV4_0),.clk(gclk));
	jdff dff_B_QDvttSih6_0(.din(w_dff_B_Qz8uHCUV4_0),.dout(w_dff_B_QDvttSih6_0),.clk(gclk));
	jdff dff_B_1wbw8wJY6_0(.din(w_dff_B_QDvttSih6_0),.dout(w_dff_B_1wbw8wJY6_0),.clk(gclk));
	jdff dff_B_AfiNB8fZ2_0(.din(w_dff_B_1wbw8wJY6_0),.dout(w_dff_B_AfiNB8fZ2_0),.clk(gclk));
	jdff dff_B_MG0o2Qo24_0(.din(w_dff_B_AfiNB8fZ2_0),.dout(w_dff_B_MG0o2Qo24_0),.clk(gclk));
	jdff dff_B_IWeYiSDd6_0(.din(w_dff_B_MG0o2Qo24_0),.dout(w_dff_B_IWeYiSDd6_0),.clk(gclk));
	jdff dff_B_5qv22RKN8_0(.din(w_dff_B_IWeYiSDd6_0),.dout(w_dff_B_5qv22RKN8_0),.clk(gclk));
	jdff dff_B_GwwHDRTv8_0(.din(w_dff_B_5qv22RKN8_0),.dout(w_dff_B_GwwHDRTv8_0),.clk(gclk));
	jdff dff_B_1YIloZ8U6_0(.din(w_dff_B_GwwHDRTv8_0),.dout(w_dff_B_1YIloZ8U6_0),.clk(gclk));
	jdff dff_B_NZifnjeV3_0(.din(w_dff_B_1YIloZ8U6_0),.dout(w_dff_B_NZifnjeV3_0),.clk(gclk));
	jdff dff_B_vYBVypmd4_0(.din(w_dff_B_NZifnjeV3_0),.dout(w_dff_B_vYBVypmd4_0),.clk(gclk));
	jdff dff_B_KjRmi9ya0_0(.din(w_dff_B_vYBVypmd4_0),.dout(w_dff_B_KjRmi9ya0_0),.clk(gclk));
	jdff dff_B_ccO3gIBX2_0(.din(w_dff_B_KjRmi9ya0_0),.dout(w_dff_B_ccO3gIBX2_0),.clk(gclk));
	jdff dff_B_xzfbcL2i0_0(.din(w_dff_B_ccO3gIBX2_0),.dout(w_dff_B_xzfbcL2i0_0),.clk(gclk));
	jdff dff_B_G05FjTiQ9_0(.din(w_dff_B_xzfbcL2i0_0),.dout(w_dff_B_G05FjTiQ9_0),.clk(gclk));
	jdff dff_B_7KI8fp1b4_0(.din(w_dff_B_G05FjTiQ9_0),.dout(w_dff_B_7KI8fp1b4_0),.clk(gclk));
	jdff dff_B_TfPXlL9x9_0(.din(w_dff_B_7KI8fp1b4_0),.dout(w_dff_B_TfPXlL9x9_0),.clk(gclk));
	jdff dff_B_38VjsrQn8_0(.din(w_dff_B_TfPXlL9x9_0),.dout(w_dff_B_38VjsrQn8_0),.clk(gclk));
	jdff dff_B_czTqUtTy6_0(.din(w_dff_B_38VjsrQn8_0),.dout(w_dff_B_czTqUtTy6_0),.clk(gclk));
	jdff dff_B_TcphjBEB3_0(.din(w_dff_B_czTqUtTy6_0),.dout(w_dff_B_TcphjBEB3_0),.clk(gclk));
	jdff dff_B_uPb3CPjh2_0(.din(w_dff_B_TcphjBEB3_0),.dout(w_dff_B_uPb3CPjh2_0),.clk(gclk));
	jdff dff_B_u4rw8Rgz0_1(.din(n1269),.dout(w_dff_B_u4rw8Rgz0_1),.clk(gclk));
	jdff dff_B_Ra935SOO5_1(.din(w_dff_B_u4rw8Rgz0_1),.dout(w_dff_B_Ra935SOO5_1),.clk(gclk));
	jdff dff_B_cEyVO6YC9_0(.din(n1286),.dout(w_dff_B_cEyVO6YC9_0),.clk(gclk));
	jdff dff_B_xpsMYQWM6_0(.din(w_dff_B_cEyVO6YC9_0),.dout(w_dff_B_xpsMYQWM6_0),.clk(gclk));
	jdff dff_B_JuhiCCYr2_0(.din(w_dff_B_xpsMYQWM6_0),.dout(w_dff_B_JuhiCCYr2_0),.clk(gclk));
	jdff dff_B_qFhmG7bL7_0(.din(w_dff_B_JuhiCCYr2_0),.dout(w_dff_B_qFhmG7bL7_0),.clk(gclk));
	jdff dff_B_QzSkQ6Ak8_0(.din(w_dff_B_qFhmG7bL7_0),.dout(w_dff_B_QzSkQ6Ak8_0),.clk(gclk));
	jdff dff_B_fKiclD4E7_0(.din(w_dff_B_QzSkQ6Ak8_0),.dout(w_dff_B_fKiclD4E7_0),.clk(gclk));
	jdff dff_B_62nVizES5_0(.din(w_dff_B_fKiclD4E7_0),.dout(w_dff_B_62nVizES5_0),.clk(gclk));
	jdff dff_B_BqAnvREk8_0(.din(w_dff_B_62nVizES5_0),.dout(w_dff_B_BqAnvREk8_0),.clk(gclk));
	jdff dff_B_ks4pwvVr8_0(.din(w_dff_B_BqAnvREk8_0),.dout(w_dff_B_ks4pwvVr8_0),.clk(gclk));
	jdff dff_B_zqX8sWj22_0(.din(w_dff_B_ks4pwvVr8_0),.dout(w_dff_B_zqX8sWj22_0),.clk(gclk));
	jdff dff_B_QEUynro25_0(.din(w_dff_B_zqX8sWj22_0),.dout(w_dff_B_QEUynro25_0),.clk(gclk));
	jdff dff_B_VucP6jzv4_0(.din(w_dff_B_QEUynro25_0),.dout(w_dff_B_VucP6jzv4_0),.clk(gclk));
	jdff dff_B_a4Q4fBzU3_0(.din(w_dff_B_VucP6jzv4_0),.dout(w_dff_B_a4Q4fBzU3_0),.clk(gclk));
	jdff dff_B_c9lb9DbS0_0(.din(w_dff_B_a4Q4fBzU3_0),.dout(w_dff_B_c9lb9DbS0_0),.clk(gclk));
	jdff dff_B_QACwt3cS3_0(.din(w_dff_B_c9lb9DbS0_0),.dout(w_dff_B_QACwt3cS3_0),.clk(gclk));
	jdff dff_B_hY2ktPb48_0(.din(w_dff_B_QACwt3cS3_0),.dout(w_dff_B_hY2ktPb48_0),.clk(gclk));
	jdff dff_B_oAW1pntw0_0(.din(w_dff_B_hY2ktPb48_0),.dout(w_dff_B_oAW1pntw0_0),.clk(gclk));
	jdff dff_B_qQshgjp18_0(.din(w_dff_B_oAW1pntw0_0),.dout(w_dff_B_qQshgjp18_0),.clk(gclk));
	jdff dff_B_UaN4cfuL3_0(.din(w_dff_B_qQshgjp18_0),.dout(w_dff_B_UaN4cfuL3_0),.clk(gclk));
	jdff dff_B_DAHkaWdf2_0(.din(w_dff_B_UaN4cfuL3_0),.dout(w_dff_B_DAHkaWdf2_0),.clk(gclk));
	jdff dff_B_uqs01sJ80_1(.din(n1278),.dout(w_dff_B_uqs01sJ80_1),.clk(gclk));
	jdff dff_B_KCaiDqnp0_1(.din(w_dff_B_uqs01sJ80_1),.dout(w_dff_B_KCaiDqnp0_1),.clk(gclk));
	jdff dff_B_69LiQYJu4_0(.din(n1295),.dout(w_dff_B_69LiQYJu4_0),.clk(gclk));
	jdff dff_B_fqIW3bFR4_0(.din(w_dff_B_69LiQYJu4_0),.dout(w_dff_B_fqIW3bFR4_0),.clk(gclk));
	jdff dff_B_wOMXoJY60_0(.din(w_dff_B_fqIW3bFR4_0),.dout(w_dff_B_wOMXoJY60_0),.clk(gclk));
	jdff dff_B_aUOW9rYY7_0(.din(w_dff_B_wOMXoJY60_0),.dout(w_dff_B_aUOW9rYY7_0),.clk(gclk));
	jdff dff_B_EHHoNx5I6_0(.din(w_dff_B_aUOW9rYY7_0),.dout(w_dff_B_EHHoNx5I6_0),.clk(gclk));
	jdff dff_B_Wf6AqbXm9_0(.din(w_dff_B_EHHoNx5I6_0),.dout(w_dff_B_Wf6AqbXm9_0),.clk(gclk));
	jdff dff_B_jutsZBvQ0_0(.din(w_dff_B_Wf6AqbXm9_0),.dout(w_dff_B_jutsZBvQ0_0),.clk(gclk));
	jdff dff_B_0v1Dyp9T7_0(.din(w_dff_B_jutsZBvQ0_0),.dout(w_dff_B_0v1Dyp9T7_0),.clk(gclk));
	jdff dff_B_rcDig1ys9_0(.din(w_dff_B_0v1Dyp9T7_0),.dout(w_dff_B_rcDig1ys9_0),.clk(gclk));
	jdff dff_B_QmnjDsoR4_0(.din(w_dff_B_rcDig1ys9_0),.dout(w_dff_B_QmnjDsoR4_0),.clk(gclk));
	jdff dff_B_PpgskbsT6_0(.din(w_dff_B_QmnjDsoR4_0),.dout(w_dff_B_PpgskbsT6_0),.clk(gclk));
	jdff dff_B_Myx8Pffw1_0(.din(w_dff_B_PpgskbsT6_0),.dout(w_dff_B_Myx8Pffw1_0),.clk(gclk));
	jdff dff_B_qGj7Qvvm7_0(.din(w_dff_B_Myx8Pffw1_0),.dout(w_dff_B_qGj7Qvvm7_0),.clk(gclk));
	jdff dff_B_GNMiNKJC0_0(.din(w_dff_B_qGj7Qvvm7_0),.dout(w_dff_B_GNMiNKJC0_0),.clk(gclk));
	jdff dff_B_UDIbEXSU4_0(.din(w_dff_B_GNMiNKJC0_0),.dout(w_dff_B_UDIbEXSU4_0),.clk(gclk));
	jdff dff_B_WVOelZyV9_0(.din(w_dff_B_UDIbEXSU4_0),.dout(w_dff_B_WVOelZyV9_0),.clk(gclk));
	jdff dff_B_1R4rIOX53_0(.din(w_dff_B_WVOelZyV9_0),.dout(w_dff_B_1R4rIOX53_0),.clk(gclk));
	jdff dff_B_6dQTneQC5_0(.din(w_dff_B_1R4rIOX53_0),.dout(w_dff_B_6dQTneQC5_0),.clk(gclk));
	jdff dff_B_IV3JDKjo5_0(.din(w_dff_B_6dQTneQC5_0),.dout(w_dff_B_IV3JDKjo5_0),.clk(gclk));
	jdff dff_B_hnqC9Wmu9_0(.din(w_dff_B_IV3JDKjo5_0),.dout(w_dff_B_hnqC9Wmu9_0),.clk(gclk));
	jdff dff_B_hm6V1Wnr4_1(.din(n1288),.dout(w_dff_B_hm6V1Wnr4_1),.clk(gclk));
	jdff dff_B_OWmEd2mP0_0(.din(n1306),.dout(w_dff_B_OWmEd2mP0_0),.clk(gclk));
	jdff dff_B_hj10rN1A3_0(.din(w_dff_B_OWmEd2mP0_0),.dout(w_dff_B_hj10rN1A3_0),.clk(gclk));
	jdff dff_B_oBefjrpf0_0(.din(w_dff_B_hj10rN1A3_0),.dout(w_dff_B_oBefjrpf0_0),.clk(gclk));
	jdff dff_B_TO8PTPjT1_0(.din(w_dff_B_oBefjrpf0_0),.dout(w_dff_B_TO8PTPjT1_0),.clk(gclk));
	jdff dff_B_LhOTchzw1_0(.din(w_dff_B_TO8PTPjT1_0),.dout(w_dff_B_LhOTchzw1_0),.clk(gclk));
	jdff dff_B_BkCZ02jQ4_0(.din(w_dff_B_LhOTchzw1_0),.dout(w_dff_B_BkCZ02jQ4_0),.clk(gclk));
	jdff dff_B_V4HvfDVr6_0(.din(w_dff_B_BkCZ02jQ4_0),.dout(w_dff_B_V4HvfDVr6_0),.clk(gclk));
	jdff dff_B_TNujeIGZ0_0(.din(w_dff_B_V4HvfDVr6_0),.dout(w_dff_B_TNujeIGZ0_0),.clk(gclk));
	jdff dff_B_v7k8lmsA5_0(.din(w_dff_B_TNujeIGZ0_0),.dout(w_dff_B_v7k8lmsA5_0),.clk(gclk));
	jdff dff_B_nGBsGt7N0_0(.din(w_dff_B_v7k8lmsA5_0),.dout(w_dff_B_nGBsGt7N0_0),.clk(gclk));
	jdff dff_B_lrfQuAcZ7_0(.din(w_dff_B_nGBsGt7N0_0),.dout(w_dff_B_lrfQuAcZ7_0),.clk(gclk));
	jdff dff_B_KLt5u9AE4_0(.din(w_dff_B_lrfQuAcZ7_0),.dout(w_dff_B_KLt5u9AE4_0),.clk(gclk));
	jdff dff_B_e7fmj5O26_0(.din(w_dff_B_KLt5u9AE4_0),.dout(w_dff_B_e7fmj5O26_0),.clk(gclk));
	jdff dff_B_z52kPYiP3_0(.din(w_dff_B_e7fmj5O26_0),.dout(w_dff_B_z52kPYiP3_0),.clk(gclk));
	jdff dff_B_sLD9yEMq8_0(.din(w_dff_B_z52kPYiP3_0),.dout(w_dff_B_sLD9yEMq8_0),.clk(gclk));
	jdff dff_B_60rfgGGJ6_0(.din(w_dff_B_sLD9yEMq8_0),.dout(w_dff_B_60rfgGGJ6_0),.clk(gclk));
	jdff dff_B_YqnqiXvc0_0(.din(w_dff_B_60rfgGGJ6_0),.dout(w_dff_B_YqnqiXvc0_0),.clk(gclk));
	jdff dff_B_Wr43gGI56_0(.din(w_dff_B_YqnqiXvc0_0),.dout(w_dff_B_Wr43gGI56_0),.clk(gclk));
	jdff dff_B_6tvoiiKt9_0(.din(w_dff_B_Wr43gGI56_0),.dout(w_dff_B_6tvoiiKt9_0),.clk(gclk));
	jdff dff_B_xIPwIWEz4_1(.din(n1298),.dout(w_dff_B_xIPwIWEz4_1),.clk(gclk));
	jdff dff_B_euO5JJwY7_1(.din(w_dff_B_xIPwIWEz4_1),.dout(w_dff_B_euO5JJwY7_1),.clk(gclk));
	jdff dff_B_6YQPmrv72_1(.din(w_dff_B_euO5JJwY7_1),.dout(w_dff_B_6YQPmrv72_1),.clk(gclk));
	jdff dff_B_gWcJGIq66_0(.din(n1315),.dout(w_dff_B_gWcJGIq66_0),.clk(gclk));
	jdff dff_B_IAwTJ3XL7_0(.din(w_dff_B_gWcJGIq66_0),.dout(w_dff_B_IAwTJ3XL7_0),.clk(gclk));
	jdff dff_B_q2hityIo8_0(.din(w_dff_B_IAwTJ3XL7_0),.dout(w_dff_B_q2hityIo8_0),.clk(gclk));
	jdff dff_B_7jLilQQb2_0(.din(w_dff_B_q2hityIo8_0),.dout(w_dff_B_7jLilQQb2_0),.clk(gclk));
	jdff dff_B_dAjVjDeS6_0(.din(w_dff_B_7jLilQQb2_0),.dout(w_dff_B_dAjVjDeS6_0),.clk(gclk));
	jdff dff_B_xzrmSwrU6_0(.din(w_dff_B_dAjVjDeS6_0),.dout(w_dff_B_xzrmSwrU6_0),.clk(gclk));
	jdff dff_B_HcsDbYQR9_0(.din(w_dff_B_xzrmSwrU6_0),.dout(w_dff_B_HcsDbYQR9_0),.clk(gclk));
	jdff dff_B_yRcSlln43_0(.din(w_dff_B_HcsDbYQR9_0),.dout(w_dff_B_yRcSlln43_0),.clk(gclk));
	jdff dff_B_2pOQFaYC7_0(.din(w_dff_B_yRcSlln43_0),.dout(w_dff_B_2pOQFaYC7_0),.clk(gclk));
	jdff dff_B_UO99Msyj3_0(.din(w_dff_B_2pOQFaYC7_0),.dout(w_dff_B_UO99Msyj3_0),.clk(gclk));
	jdff dff_B_2s5Dp15B0_0(.din(w_dff_B_UO99Msyj3_0),.dout(w_dff_B_2s5Dp15B0_0),.clk(gclk));
	jdff dff_B_vTtu1iVF2_0(.din(w_dff_B_2s5Dp15B0_0),.dout(w_dff_B_vTtu1iVF2_0),.clk(gclk));
	jdff dff_B_6eV0mzNp9_0(.din(w_dff_B_vTtu1iVF2_0),.dout(w_dff_B_6eV0mzNp9_0),.clk(gclk));
	jdff dff_B_bRjX76MI7_0(.din(w_dff_B_6eV0mzNp9_0),.dout(w_dff_B_bRjX76MI7_0),.clk(gclk));
	jdff dff_B_iLxVazOV3_0(.din(w_dff_B_bRjX76MI7_0),.dout(w_dff_B_iLxVazOV3_0),.clk(gclk));
	jdff dff_B_H0r8ToYp6_0(.din(w_dff_B_iLxVazOV3_0),.dout(w_dff_B_H0r8ToYp6_0),.clk(gclk));
	jdff dff_B_T8LeiYVU3_0(.din(w_dff_B_H0r8ToYp6_0),.dout(w_dff_B_T8LeiYVU3_0),.clk(gclk));
	jdff dff_B_G64iDjM79_0(.din(w_dff_B_T8LeiYVU3_0),.dout(w_dff_B_G64iDjM79_0),.clk(gclk));
	jdff dff_B_pQoMNivd5_0(.din(w_dff_B_G64iDjM79_0),.dout(w_dff_B_pQoMNivd5_0),.clk(gclk));
	jdff dff_B_9PryGx0C4_0(.din(w_dff_B_pQoMNivd5_0),.dout(w_dff_B_9PryGx0C4_0),.clk(gclk));
	jdff dff_B_mO2zrwY48_1(.din(n1308),.dout(w_dff_B_mO2zrwY48_1),.clk(gclk));
	jdff dff_B_bodC3ZIz1_1(.din(w_dff_B_mO2zrwY48_1),.dout(w_dff_B_bodC3ZIz1_1),.clk(gclk));
	jdff dff_B_UXK7apd76_0(.din(n1324),.dout(w_dff_B_UXK7apd76_0),.clk(gclk));
	jdff dff_B_adkpNogp9_0(.din(w_dff_B_UXK7apd76_0),.dout(w_dff_B_adkpNogp9_0),.clk(gclk));
	jdff dff_B_kTgAz6n64_0(.din(w_dff_B_adkpNogp9_0),.dout(w_dff_B_kTgAz6n64_0),.clk(gclk));
	jdff dff_B_LtrCHKnv5_0(.din(w_dff_B_kTgAz6n64_0),.dout(w_dff_B_LtrCHKnv5_0),.clk(gclk));
	jdff dff_B_XTQDDthb0_0(.din(w_dff_B_LtrCHKnv5_0),.dout(w_dff_B_XTQDDthb0_0),.clk(gclk));
	jdff dff_B_V5aBo9AX3_0(.din(w_dff_B_XTQDDthb0_0),.dout(w_dff_B_V5aBo9AX3_0),.clk(gclk));
	jdff dff_B_etyq1JQu7_0(.din(w_dff_B_V5aBo9AX3_0),.dout(w_dff_B_etyq1JQu7_0),.clk(gclk));
	jdff dff_B_iUrlhMZ51_0(.din(w_dff_B_etyq1JQu7_0),.dout(w_dff_B_iUrlhMZ51_0),.clk(gclk));
	jdff dff_B_y0hQiWpe2_0(.din(w_dff_B_iUrlhMZ51_0),.dout(w_dff_B_y0hQiWpe2_0),.clk(gclk));
	jdff dff_B_wutJfm3E8_0(.din(w_dff_B_y0hQiWpe2_0),.dout(w_dff_B_wutJfm3E8_0),.clk(gclk));
	jdff dff_B_aIMHjenc7_0(.din(w_dff_B_wutJfm3E8_0),.dout(w_dff_B_aIMHjenc7_0),.clk(gclk));
	jdff dff_B_fONAimIc1_0(.din(w_dff_B_aIMHjenc7_0),.dout(w_dff_B_fONAimIc1_0),.clk(gclk));
	jdff dff_B_zeplCKIF0_0(.din(w_dff_B_fONAimIc1_0),.dout(w_dff_B_zeplCKIF0_0),.clk(gclk));
	jdff dff_B_FrhCLHKb5_0(.din(w_dff_B_zeplCKIF0_0),.dout(w_dff_B_FrhCLHKb5_0),.clk(gclk));
	jdff dff_B_gCPQXe5a1_0(.din(w_dff_B_FrhCLHKb5_0),.dout(w_dff_B_gCPQXe5a1_0),.clk(gclk));
	jdff dff_B_uAy1IlF57_0(.din(w_dff_B_gCPQXe5a1_0),.dout(w_dff_B_uAy1IlF57_0),.clk(gclk));
	jdff dff_B_kD783my76_0(.din(w_dff_B_uAy1IlF57_0),.dout(w_dff_B_kD783my76_0),.clk(gclk));
	jdff dff_B_4DerBogf4_0(.din(w_dff_B_kD783my76_0),.dout(w_dff_B_4DerBogf4_0),.clk(gclk));
	jdff dff_B_7nGbBVgL3_0(.din(w_dff_B_4DerBogf4_0),.dout(w_dff_B_7nGbBVgL3_0),.clk(gclk));
	jdff dff_B_fSABNbnM3_0(.din(w_dff_B_7nGbBVgL3_0),.dout(w_dff_B_fSABNbnM3_0),.clk(gclk));
	jdff dff_B_5OLRqP5N6_1(.din(n1317),.dout(w_dff_B_5OLRqP5N6_1),.clk(gclk));
	jdff dff_B_dZ9GkMBf3_0(.din(n1333),.dout(w_dff_B_dZ9GkMBf3_0),.clk(gclk));
	jdff dff_B_9dSPemVe7_0(.din(w_dff_B_dZ9GkMBf3_0),.dout(w_dff_B_9dSPemVe7_0),.clk(gclk));
	jdff dff_B_qyBGboWp9_0(.din(w_dff_B_9dSPemVe7_0),.dout(w_dff_B_qyBGboWp9_0),.clk(gclk));
	jdff dff_B_ROktWTfw4_0(.din(w_dff_B_qyBGboWp9_0),.dout(w_dff_B_ROktWTfw4_0),.clk(gclk));
	jdff dff_B_qVXjMkcK7_0(.din(w_dff_B_ROktWTfw4_0),.dout(w_dff_B_qVXjMkcK7_0),.clk(gclk));
	jdff dff_B_q1dhFLJr8_0(.din(w_dff_B_qVXjMkcK7_0),.dout(w_dff_B_q1dhFLJr8_0),.clk(gclk));
	jdff dff_B_6jKirput2_0(.din(w_dff_B_q1dhFLJr8_0),.dout(w_dff_B_6jKirput2_0),.clk(gclk));
	jdff dff_B_07j5ZC1S3_0(.din(w_dff_B_6jKirput2_0),.dout(w_dff_B_07j5ZC1S3_0),.clk(gclk));
	jdff dff_B_ZxQWxorr6_0(.din(w_dff_B_07j5ZC1S3_0),.dout(w_dff_B_ZxQWxorr6_0),.clk(gclk));
	jdff dff_B_UGROEVBm4_0(.din(w_dff_B_ZxQWxorr6_0),.dout(w_dff_B_UGROEVBm4_0),.clk(gclk));
	jdff dff_B_FsFLOcxn6_0(.din(w_dff_B_UGROEVBm4_0),.dout(w_dff_B_FsFLOcxn6_0),.clk(gclk));
	jdff dff_B_9i6DTtca6_0(.din(w_dff_B_FsFLOcxn6_0),.dout(w_dff_B_9i6DTtca6_0),.clk(gclk));
	jdff dff_B_Uct4yhOZ9_0(.din(w_dff_B_9i6DTtca6_0),.dout(w_dff_B_Uct4yhOZ9_0),.clk(gclk));
	jdff dff_B_911KCZeX7_0(.din(w_dff_B_Uct4yhOZ9_0),.dout(w_dff_B_911KCZeX7_0),.clk(gclk));
	jdff dff_B_9T6epfvs1_0(.din(w_dff_B_911KCZeX7_0),.dout(w_dff_B_9T6epfvs1_0),.clk(gclk));
	jdff dff_B_0cZr8IVw2_0(.din(w_dff_B_9T6epfvs1_0),.dout(w_dff_B_0cZr8IVw2_0),.clk(gclk));
	jdff dff_B_1A5EE5ey4_0(.din(w_dff_B_0cZr8IVw2_0),.dout(w_dff_B_1A5EE5ey4_0),.clk(gclk));
	jdff dff_B_sYnGfNlc2_0(.din(w_dff_B_1A5EE5ey4_0),.dout(w_dff_B_sYnGfNlc2_0),.clk(gclk));
	jdff dff_B_3gu5XD3k4_0(.din(w_dff_B_sYnGfNlc2_0),.dout(w_dff_B_3gu5XD3k4_0),.clk(gclk));
	jdff dff_B_7meUkI0u9_1(.din(n1326),.dout(w_dff_B_7meUkI0u9_1),.clk(gclk));
	jdff dff_B_jp45zAfo8_1(.din(w_dff_B_7meUkI0u9_1),.dout(w_dff_B_jp45zAfo8_1),.clk(gclk));
	jdff dff_B_2v01HJmp0_1(.din(w_dff_B_jp45zAfo8_1),.dout(w_dff_B_2v01HJmp0_1),.clk(gclk));
	jdff dff_B_TDMGOcA01_0(.din(n1341),.dout(w_dff_B_TDMGOcA01_0),.clk(gclk));
	jdff dff_B_LGAgcm9p9_0(.din(w_dff_B_TDMGOcA01_0),.dout(w_dff_B_LGAgcm9p9_0),.clk(gclk));
	jdff dff_B_Ch9jmSvg4_0(.din(w_dff_B_LGAgcm9p9_0),.dout(w_dff_B_Ch9jmSvg4_0),.clk(gclk));
	jdff dff_B_aMVLQMCi1_0(.din(w_dff_B_Ch9jmSvg4_0),.dout(w_dff_B_aMVLQMCi1_0),.clk(gclk));
	jdff dff_B_ipVPKn0K3_0(.din(w_dff_B_aMVLQMCi1_0),.dout(w_dff_B_ipVPKn0K3_0),.clk(gclk));
	jdff dff_B_7n6S5Bru3_0(.din(w_dff_B_ipVPKn0K3_0),.dout(w_dff_B_7n6S5Bru3_0),.clk(gclk));
	jdff dff_B_pibtBhVE9_0(.din(w_dff_B_7n6S5Bru3_0),.dout(w_dff_B_pibtBhVE9_0),.clk(gclk));
	jdff dff_B_94kI7B865_0(.din(w_dff_B_pibtBhVE9_0),.dout(w_dff_B_94kI7B865_0),.clk(gclk));
	jdff dff_B_F3OXVLc20_0(.din(w_dff_B_94kI7B865_0),.dout(w_dff_B_F3OXVLc20_0),.clk(gclk));
	jdff dff_B_ZDwl5qtR0_0(.din(w_dff_B_F3OXVLc20_0),.dout(w_dff_B_ZDwl5qtR0_0),.clk(gclk));
	jdff dff_B_IrzLVC3D6_0(.din(w_dff_B_ZDwl5qtR0_0),.dout(w_dff_B_IrzLVC3D6_0),.clk(gclk));
	jdff dff_B_qE8bZEgv9_0(.din(w_dff_B_IrzLVC3D6_0),.dout(w_dff_B_qE8bZEgv9_0),.clk(gclk));
	jdff dff_B_P8ZLFqVY3_0(.din(w_dff_B_qE8bZEgv9_0),.dout(w_dff_B_P8ZLFqVY3_0),.clk(gclk));
	jdff dff_B_e9EC6BW10_0(.din(w_dff_B_P8ZLFqVY3_0),.dout(w_dff_B_e9EC6BW10_0),.clk(gclk));
	jdff dff_B_4psK4a7V2_0(.din(w_dff_B_e9EC6BW10_0),.dout(w_dff_B_4psK4a7V2_0),.clk(gclk));
	jdff dff_B_izuzLfvx0_0(.din(w_dff_B_4psK4a7V2_0),.dout(w_dff_B_izuzLfvx0_0),.clk(gclk));
	jdff dff_B_EkczzdOU3_0(.din(w_dff_B_izuzLfvx0_0),.dout(w_dff_B_EkczzdOU3_0),.clk(gclk));
	jdff dff_B_G0EZjB2W9_0(.din(w_dff_B_EkczzdOU3_0),.dout(w_dff_B_G0EZjB2W9_0),.clk(gclk));
	jdff dff_B_AWnJyqHo5_1(.din(n1335),.dout(w_dff_B_AWnJyqHo5_1),.clk(gclk));
	jdff dff_B_K6LR4AuM9_1(.din(w_dff_B_AWnJyqHo5_1),.dout(w_dff_B_K6LR4AuM9_1),.clk(gclk));
	jdff dff_B_E6w3HOae8_1(.din(w_dff_B_K6LR4AuM9_1),.dout(w_dff_B_E6w3HOae8_1),.clk(gclk));
	jdff dff_A_gbXeYHvc4_0(.dout(w_n999_2[0]),.din(w_dff_A_gbXeYHvc4_0),.clk(gclk));
	jdff dff_A_AOg5Gn541_0(.dout(w_dff_A_gbXeYHvc4_0),.din(w_dff_A_AOg5Gn541_0),.clk(gclk));
	jdff dff_A_Ml7TkT2B2_0(.dout(w_dff_A_AOg5Gn541_0),.din(w_dff_A_Ml7TkT2B2_0),.clk(gclk));
	jdff dff_A_WcF6UrZo9_0(.dout(w_dff_A_Ml7TkT2B2_0),.din(w_dff_A_WcF6UrZo9_0),.clk(gclk));
	jdff dff_A_Tvcmhn8o9_0(.dout(w_dff_A_WcF6UrZo9_0),.din(w_dff_A_Tvcmhn8o9_0),.clk(gclk));
	jdff dff_A_ivUFOrEV2_0(.dout(w_dff_A_Tvcmhn8o9_0),.din(w_dff_A_ivUFOrEV2_0),.clk(gclk));
	jdff dff_A_NTmV4l3H9_1(.dout(w_n999_2[1]),.din(w_dff_A_NTmV4l3H9_1),.clk(gclk));
	jdff dff_A_zjkof0W22_0(.dout(w_G1689_3[0]),.din(w_dff_A_zjkof0W22_0),.clk(gclk));
	jdff dff_A_RCBIsjoV0_0(.dout(w_dff_A_zjkof0W22_0),.din(w_dff_A_RCBIsjoV0_0),.clk(gclk));
	jdff dff_A_WjxIsejb9_0(.dout(w_dff_A_RCBIsjoV0_0),.din(w_dff_A_WjxIsejb9_0),.clk(gclk));
	jdff dff_A_iU8dCjJT9_0(.dout(w_dff_A_WjxIsejb9_0),.din(w_dff_A_iU8dCjJT9_0),.clk(gclk));
	jdff dff_A_FA9bbewr7_1(.dout(w_G1689_3[1]),.din(w_dff_A_FA9bbewr7_1),.clk(gclk));
	jdff dff_A_jF0uhBbI8_1(.dout(w_dff_A_FA9bbewr7_1),.din(w_dff_A_jF0uhBbI8_1),.clk(gclk));
	jdff dff_A_ZPuicIJu9_0(.dout(w_G137_6[0]),.din(w_dff_A_ZPuicIJu9_0),.clk(gclk));
	jdff dff_A_L9DBkmu36_0(.dout(w_dff_A_ZPuicIJu9_0),.din(w_dff_A_L9DBkmu36_0),.clk(gclk));
	jdff dff_A_PKx2ksOL4_0(.dout(w_dff_A_L9DBkmu36_0),.din(w_dff_A_PKx2ksOL4_0),.clk(gclk));
	jdff dff_A_mvxhc2rT6_0(.dout(w_dff_A_PKx2ksOL4_0),.din(w_dff_A_mvxhc2rT6_0),.clk(gclk));
	jdff dff_A_B1rvDeUY7_0(.dout(w_dff_A_mvxhc2rT6_0),.din(w_dff_A_B1rvDeUY7_0),.clk(gclk));
	jdff dff_A_xKN9JgQ47_0(.dout(w_dff_A_B1rvDeUY7_0),.din(w_dff_A_xKN9JgQ47_0),.clk(gclk));
	jdff dff_A_YvJlGhkA9_1(.dout(w_G137_6[1]),.din(w_dff_A_YvJlGhkA9_1),.clk(gclk));
	jdff dff_B_tpHjaZk99_0(.din(n1350),.dout(w_dff_B_tpHjaZk99_0),.clk(gclk));
	jdff dff_B_cNw2JI3f9_0(.din(w_dff_B_tpHjaZk99_0),.dout(w_dff_B_cNw2JI3f9_0),.clk(gclk));
	jdff dff_B_Qmi3bZFr2_0(.din(w_dff_B_cNw2JI3f9_0),.dout(w_dff_B_Qmi3bZFr2_0),.clk(gclk));
	jdff dff_B_e6NDENEr4_0(.din(w_dff_B_Qmi3bZFr2_0),.dout(w_dff_B_e6NDENEr4_0),.clk(gclk));
	jdff dff_B_CarBhQgQ1_0(.din(w_dff_B_e6NDENEr4_0),.dout(w_dff_B_CarBhQgQ1_0),.clk(gclk));
	jdff dff_B_o6eCxcjT9_0(.din(w_dff_B_CarBhQgQ1_0),.dout(w_dff_B_o6eCxcjT9_0),.clk(gclk));
	jdff dff_B_0DlEfZDK9_0(.din(w_dff_B_o6eCxcjT9_0),.dout(w_dff_B_0DlEfZDK9_0),.clk(gclk));
	jdff dff_B_kiATk3UA4_0(.din(w_dff_B_0DlEfZDK9_0),.dout(w_dff_B_kiATk3UA4_0),.clk(gclk));
	jdff dff_B_kcchts2Z2_0(.din(w_dff_B_kiATk3UA4_0),.dout(w_dff_B_kcchts2Z2_0),.clk(gclk));
	jdff dff_B_3qg3vMfd6_0(.din(w_dff_B_kcchts2Z2_0),.dout(w_dff_B_3qg3vMfd6_0),.clk(gclk));
	jdff dff_B_yf1GRtxK2_0(.din(w_dff_B_3qg3vMfd6_0),.dout(w_dff_B_yf1GRtxK2_0),.clk(gclk));
	jdff dff_B_6FhekFqE8_0(.din(w_dff_B_yf1GRtxK2_0),.dout(w_dff_B_6FhekFqE8_0),.clk(gclk));
	jdff dff_B_20dEYXXm0_0(.din(w_dff_B_6FhekFqE8_0),.dout(w_dff_B_20dEYXXm0_0),.clk(gclk));
	jdff dff_B_B9wMvP9S5_0(.din(w_dff_B_20dEYXXm0_0),.dout(w_dff_B_B9wMvP9S5_0),.clk(gclk));
	jdff dff_B_hUnmoUaW2_0(.din(w_dff_B_B9wMvP9S5_0),.dout(w_dff_B_hUnmoUaW2_0),.clk(gclk));
	jdff dff_B_NYOrrIvv7_0(.din(w_dff_B_hUnmoUaW2_0),.dout(w_dff_B_NYOrrIvv7_0),.clk(gclk));
	jdff dff_B_pDBKcYpv3_0(.din(w_dff_B_NYOrrIvv7_0),.dout(w_dff_B_pDBKcYpv3_0),.clk(gclk));
	jdff dff_B_Ml0byOD53_0(.din(w_dff_B_pDBKcYpv3_0),.dout(w_dff_B_Ml0byOD53_0),.clk(gclk));
	jdff dff_B_7juUKr1R2_0(.din(w_dff_B_Ml0byOD53_0),.dout(w_dff_B_7juUKr1R2_0),.clk(gclk));
	jdff dff_B_RrZERRcd2_1(.din(n1344),.dout(w_dff_B_RrZERRcd2_1),.clk(gclk));
	jdff dff_B_dy17jKP27_1(.din(n1355),.dout(w_dff_B_dy17jKP27_1),.clk(gclk));
	jdff dff_B_NN8ODGRh3_1(.din(w_dff_B_dy17jKP27_1),.dout(w_dff_B_NN8ODGRh3_1),.clk(gclk));
	jdff dff_B_XmPbZfZG9_1(.din(w_dff_B_NN8ODGRh3_1),.dout(w_dff_B_XmPbZfZG9_1),.clk(gclk));
	jdff dff_B_o05U0mQu7_1(.din(w_dff_B_XmPbZfZG9_1),.dout(w_dff_B_o05U0mQu7_1),.clk(gclk));
	jdff dff_B_YZHheBjb5_1(.din(w_dff_B_o05U0mQu7_1),.dout(w_dff_B_YZHheBjb5_1),.clk(gclk));
	jdff dff_B_OLjlaJPK5_1(.din(w_dff_B_YZHheBjb5_1),.dout(w_dff_B_OLjlaJPK5_1),.clk(gclk));
	jdff dff_B_vyZbQ8gT1_1(.din(w_dff_B_OLjlaJPK5_1),.dout(w_dff_B_vyZbQ8gT1_1),.clk(gclk));
	jdff dff_B_wouDNh8N6_1(.din(w_dff_B_vyZbQ8gT1_1),.dout(w_dff_B_wouDNh8N6_1),.clk(gclk));
	jdff dff_B_DoSch3yf7_1(.din(w_dff_B_wouDNh8N6_1),.dout(w_dff_B_DoSch3yf7_1),.clk(gclk));
	jdff dff_B_RJC5Adxi6_1(.din(w_dff_B_DoSch3yf7_1),.dout(w_dff_B_RJC5Adxi6_1),.clk(gclk));
	jdff dff_B_QwMpfBiy3_1(.din(w_dff_B_RJC5Adxi6_1),.dout(w_dff_B_QwMpfBiy3_1),.clk(gclk));
	jdff dff_B_9oldovLf3_1(.din(w_dff_B_QwMpfBiy3_1),.dout(w_dff_B_9oldovLf3_1),.clk(gclk));
	jdff dff_B_B3uUZbeY6_1(.din(w_dff_B_9oldovLf3_1),.dout(w_dff_B_B3uUZbeY6_1),.clk(gclk));
	jdff dff_B_BOVlg43r4_1(.din(w_dff_B_B3uUZbeY6_1),.dout(w_dff_B_BOVlg43r4_1),.clk(gclk));
	jdff dff_B_Gyfxcz5j5_1(.din(w_dff_B_BOVlg43r4_1),.dout(w_dff_B_Gyfxcz5j5_1),.clk(gclk));
	jdff dff_B_2t2ERVPV8_1(.din(w_dff_B_Gyfxcz5j5_1),.dout(w_dff_B_2t2ERVPV8_1),.clk(gclk));
	jdff dff_B_blXfLzAg4_1(.din(w_dff_B_2t2ERVPV8_1),.dout(w_dff_B_blXfLzAg4_1),.clk(gclk));
	jdff dff_B_RkdtCZS46_1(.din(w_dff_B_blXfLzAg4_1),.dout(w_dff_B_RkdtCZS46_1),.clk(gclk));
	jdff dff_B_4HwUVt8K3_1(.din(w_dff_B_RkdtCZS46_1),.dout(w_dff_B_4HwUVt8K3_1),.clk(gclk));
	jdff dff_B_sHmOrsaS5_1(.din(n1356),.dout(w_dff_B_sHmOrsaS5_1),.clk(gclk));
	jdff dff_B_fOOBOERz1_1(.din(n1364),.dout(w_dff_B_fOOBOERz1_1),.clk(gclk));
	jdff dff_B_7cptEJjy1_1(.din(w_dff_B_fOOBOERz1_1),.dout(w_dff_B_7cptEJjy1_1),.clk(gclk));
	jdff dff_B_yqsMho1u5_1(.din(w_dff_B_7cptEJjy1_1),.dout(w_dff_B_yqsMho1u5_1),.clk(gclk));
	jdff dff_B_ffg94stE7_1(.din(w_dff_B_yqsMho1u5_1),.dout(w_dff_B_ffg94stE7_1),.clk(gclk));
	jdff dff_B_xR4NIlIh8_1(.din(w_dff_B_ffg94stE7_1),.dout(w_dff_B_xR4NIlIh8_1),.clk(gclk));
	jdff dff_B_RBoZkkFK0_1(.din(w_dff_B_xR4NIlIh8_1),.dout(w_dff_B_RBoZkkFK0_1),.clk(gclk));
	jdff dff_B_krzhbRS92_1(.din(w_dff_B_RBoZkkFK0_1),.dout(w_dff_B_krzhbRS92_1),.clk(gclk));
	jdff dff_B_Iye6Ecwo1_1(.din(w_dff_B_krzhbRS92_1),.dout(w_dff_B_Iye6Ecwo1_1),.clk(gclk));
	jdff dff_B_DZLXNBib9_1(.din(w_dff_B_Iye6Ecwo1_1),.dout(w_dff_B_DZLXNBib9_1),.clk(gclk));
	jdff dff_B_Gml0mgvj3_1(.din(w_dff_B_DZLXNBib9_1),.dout(w_dff_B_Gml0mgvj3_1),.clk(gclk));
	jdff dff_B_LjvRrO8y4_1(.din(w_dff_B_Gml0mgvj3_1),.dout(w_dff_B_LjvRrO8y4_1),.clk(gclk));
	jdff dff_B_xaCtBOEk5_1(.din(w_dff_B_LjvRrO8y4_1),.dout(w_dff_B_xaCtBOEk5_1),.clk(gclk));
	jdff dff_B_vNn6kkaM3_1(.din(w_dff_B_xaCtBOEk5_1),.dout(w_dff_B_vNn6kkaM3_1),.clk(gclk));
	jdff dff_B_WpYX64Gj6_1(.din(w_dff_B_vNn6kkaM3_1),.dout(w_dff_B_WpYX64Gj6_1),.clk(gclk));
	jdff dff_B_JMefzPri5_1(.din(w_dff_B_WpYX64Gj6_1),.dout(w_dff_B_JMefzPri5_1),.clk(gclk));
	jdff dff_B_2Z3tpeZB3_1(.din(w_dff_B_JMefzPri5_1),.dout(w_dff_B_2Z3tpeZB3_1),.clk(gclk));
	jdff dff_B_K2ojCJ1l3_1(.din(w_dff_B_2Z3tpeZB3_1),.dout(w_dff_B_K2ojCJ1l3_1),.clk(gclk));
	jdff dff_B_V4kzJ57b9_1(.din(w_dff_B_K2ojCJ1l3_1),.dout(w_dff_B_V4kzJ57b9_1),.clk(gclk));
	jdff dff_B_pl9hiy5V5_1(.din(w_dff_B_V4kzJ57b9_1),.dout(w_dff_B_pl9hiy5V5_1),.clk(gclk));
	jdff dff_B_2xEXa9Lg2_1(.din(w_dff_B_pl9hiy5V5_1),.dout(w_dff_B_2xEXa9Lg2_1),.clk(gclk));
	jdff dff_B_nrRPA6hl1_1(.din(n1365),.dout(w_dff_B_nrRPA6hl1_1),.clk(gclk));
	jdff dff_A_EGN9FuvV8_0(.dout(w_G1689_2[0]),.din(w_dff_A_EGN9FuvV8_0),.clk(gclk));
	jdff dff_A_M0L6Ldl49_2(.dout(w_G1689_2[2]),.din(w_dff_A_M0L6Ldl49_2),.clk(gclk));
	jdff dff_A_ikw8tFQf0_0(.dout(w_n999_1[0]),.din(w_dff_A_ikw8tFQf0_0),.clk(gclk));
	jdff dff_A_THe3ti0z9_0(.dout(w_dff_A_ikw8tFQf0_0),.din(w_dff_A_THe3ti0z9_0),.clk(gclk));
	jdff dff_A_pZ4xnjMO7_1(.dout(w_n999_1[1]),.din(w_dff_A_pZ4xnjMO7_1),.clk(gclk));
	jdff dff_A_0WmIePRO0_0(.dout(w_n999_0[0]),.din(w_dff_A_0WmIePRO0_0),.clk(gclk));
	jdff dff_A_quVqaCYT7_0(.dout(w_dff_A_0WmIePRO0_0),.din(w_dff_A_quVqaCYT7_0),.clk(gclk));
	jdff dff_A_LQdcHjuO1_0(.dout(w_dff_A_quVqaCYT7_0),.din(w_dff_A_LQdcHjuO1_0),.clk(gclk));
	jdff dff_A_NhLnp8g58_0(.dout(w_dff_A_LQdcHjuO1_0),.din(w_dff_A_NhLnp8g58_0),.clk(gclk));
	jdff dff_A_nedQqdSK4_0(.dout(w_dff_A_NhLnp8g58_0),.din(w_dff_A_nedQqdSK4_0),.clk(gclk));
	jdff dff_A_45gEDq8A8_0(.dout(w_dff_A_nedQqdSK4_0),.din(w_dff_A_45gEDq8A8_0),.clk(gclk));
	jdff dff_A_PDC8W0kX8_0(.dout(w_dff_A_45gEDq8A8_0),.din(w_dff_A_PDC8W0kX8_0),.clk(gclk));
	jdff dff_A_ezaybMgx1_0(.dout(w_dff_A_PDC8W0kX8_0),.din(w_dff_A_ezaybMgx1_0),.clk(gclk));
	jdff dff_A_KwK6V8yu7_0(.dout(w_dff_A_ezaybMgx1_0),.din(w_dff_A_KwK6V8yu7_0),.clk(gclk));
	jdff dff_A_knwgzp2Z0_0(.dout(w_dff_A_KwK6V8yu7_0),.din(w_dff_A_knwgzp2Z0_0),.clk(gclk));
	jdff dff_A_MuefKJ1V5_0(.dout(w_dff_A_knwgzp2Z0_0),.din(w_dff_A_MuefKJ1V5_0),.clk(gclk));
	jdff dff_A_GYu0ObsI3_1(.dout(w_n999_0[1]),.din(w_dff_A_GYu0ObsI3_1),.clk(gclk));
	jdff dff_A_3jKFTcgm2_1(.dout(w_dff_A_GYu0ObsI3_1),.din(w_dff_A_3jKFTcgm2_1),.clk(gclk));
	jdff dff_A_wah9tYab7_1(.dout(w_dff_A_3jKFTcgm2_1),.din(w_dff_A_wah9tYab7_1),.clk(gclk));
	jdff dff_A_MgODUluG2_1(.dout(w_dff_A_wah9tYab7_1),.din(w_dff_A_MgODUluG2_1),.clk(gclk));
	jdff dff_B_lVjrjxam5_3(.din(n999),.dout(w_dff_B_lVjrjxam5_3),.clk(gclk));
	jdff dff_B_xKL7xCJi0_3(.din(w_dff_B_lVjrjxam5_3),.dout(w_dff_B_xKL7xCJi0_3),.clk(gclk));
	jdff dff_B_EAPQsA3u5_3(.din(w_dff_B_xKL7xCJi0_3),.dout(w_dff_B_EAPQsA3u5_3),.clk(gclk));
	jdff dff_B_GNwySFt44_3(.din(w_dff_B_EAPQsA3u5_3),.dout(w_dff_B_GNwySFt44_3),.clk(gclk));
	jdff dff_B_bSoTJuYO5_3(.din(w_dff_B_GNwySFt44_3),.dout(w_dff_B_bSoTJuYO5_3),.clk(gclk));
	jdff dff_B_NPn9aIMq5_3(.din(w_dff_B_bSoTJuYO5_3),.dout(w_dff_B_NPn9aIMq5_3),.clk(gclk));
	jdff dff_B_snxe0hOv7_3(.din(w_dff_B_NPn9aIMq5_3),.dout(w_dff_B_snxe0hOv7_3),.clk(gclk));
	jdff dff_B_D4re5cxl9_3(.din(w_dff_B_snxe0hOv7_3),.dout(w_dff_B_D4re5cxl9_3),.clk(gclk));
	jdff dff_B_mVgp88tn7_3(.din(w_dff_B_D4re5cxl9_3),.dout(w_dff_B_mVgp88tn7_3),.clk(gclk));
	jdff dff_A_vqLHpnx04_0(.dout(w_G137_5[0]),.din(w_dff_A_vqLHpnx04_0),.clk(gclk));
	jdff dff_B_1kgEqDhl6_0(.din(n1377),.dout(w_dff_B_1kgEqDhl6_0),.clk(gclk));
	jdff dff_B_Bl42KRDz0_0(.din(w_dff_B_1kgEqDhl6_0),.dout(w_dff_B_Bl42KRDz0_0),.clk(gclk));
	jdff dff_B_tnYgqKKr0_0(.din(w_dff_B_Bl42KRDz0_0),.dout(w_dff_B_tnYgqKKr0_0),.clk(gclk));
	jdff dff_B_yj2pBBtj0_0(.din(w_dff_B_tnYgqKKr0_0),.dout(w_dff_B_yj2pBBtj0_0),.clk(gclk));
	jdff dff_B_evfSjFA60_0(.din(w_dff_B_yj2pBBtj0_0),.dout(w_dff_B_evfSjFA60_0),.clk(gclk));
	jdff dff_B_5Dr8PS0c4_0(.din(w_dff_B_evfSjFA60_0),.dout(w_dff_B_5Dr8PS0c4_0),.clk(gclk));
	jdff dff_B_lOtE5Dxo0_0(.din(w_dff_B_5Dr8PS0c4_0),.dout(w_dff_B_lOtE5Dxo0_0),.clk(gclk));
	jdff dff_B_UNWoYuVY6_0(.din(w_dff_B_lOtE5Dxo0_0),.dout(w_dff_B_UNWoYuVY6_0),.clk(gclk));
	jdff dff_B_uWvhuz0m4_0(.din(w_dff_B_UNWoYuVY6_0),.dout(w_dff_B_uWvhuz0m4_0),.clk(gclk));
	jdff dff_B_mdTfyy6N0_0(.din(w_dff_B_uWvhuz0m4_0),.dout(w_dff_B_mdTfyy6N0_0),.clk(gclk));
	jdff dff_B_PoXiGYQX7_0(.din(w_dff_B_mdTfyy6N0_0),.dout(w_dff_B_PoXiGYQX7_0),.clk(gclk));
	jdff dff_B_hMWuKB3c7_0(.din(w_dff_B_PoXiGYQX7_0),.dout(w_dff_B_hMWuKB3c7_0),.clk(gclk));
	jdff dff_B_sAlOrGG95_0(.din(w_dff_B_hMWuKB3c7_0),.dout(w_dff_B_sAlOrGG95_0),.clk(gclk));
	jdff dff_B_2G67SzrQ2_0(.din(w_dff_B_sAlOrGG95_0),.dout(w_dff_B_2G67SzrQ2_0),.clk(gclk));
	jdff dff_B_Ta3ZJzoP6_0(.din(w_dff_B_2G67SzrQ2_0),.dout(w_dff_B_Ta3ZJzoP6_0),.clk(gclk));
	jdff dff_B_ZHL8Q97O5_0(.din(w_dff_B_Ta3ZJzoP6_0),.dout(w_dff_B_ZHL8Q97O5_0),.clk(gclk));
	jdff dff_B_sAVEzkxK1_0(.din(w_dff_B_ZHL8Q97O5_0),.dout(w_dff_B_sAVEzkxK1_0),.clk(gclk));
	jdff dff_B_XSJFcWbz3_0(.din(w_dff_B_sAVEzkxK1_0),.dout(w_dff_B_XSJFcWbz3_0),.clk(gclk));
	jdff dff_B_QGk5GiZJ1_1(.din(n1371),.dout(w_dff_B_QGk5GiZJ1_1),.clk(gclk));
	jdff dff_B_orhWyvos4_1(.din(w_dff_B_QGk5GiZJ1_1),.dout(w_dff_B_orhWyvos4_1),.clk(gclk));
	jdff dff_B_LBJurNfu5_1(.din(w_dff_B_orhWyvos4_1),.dout(w_dff_B_LBJurNfu5_1),.clk(gclk));
	jdff dff_A_jSks2Rud7_0(.dout(w_n1007_2[0]),.din(w_dff_A_jSks2Rud7_0),.clk(gclk));
	jdff dff_A_XLBgMlmK4_0(.dout(w_dff_A_jSks2Rud7_0),.din(w_dff_A_XLBgMlmK4_0),.clk(gclk));
	jdff dff_A_Ea0dKlLg2_0(.dout(w_dff_A_XLBgMlmK4_0),.din(w_dff_A_Ea0dKlLg2_0),.clk(gclk));
	jdff dff_A_zRPifxMd7_0(.dout(w_dff_A_Ea0dKlLg2_0),.din(w_dff_A_zRPifxMd7_0),.clk(gclk));
	jdff dff_A_S6lmztv56_0(.dout(w_dff_A_zRPifxMd7_0),.din(w_dff_A_S6lmztv56_0),.clk(gclk));
	jdff dff_A_dgPqd10H5_0(.dout(w_dff_A_S6lmztv56_0),.din(w_dff_A_dgPqd10H5_0),.clk(gclk));
	jdff dff_A_LTUJUBnO9_1(.dout(w_n1007_2[1]),.din(w_dff_A_LTUJUBnO9_1),.clk(gclk));
	jdff dff_B_p4yWtnyB7_1(.din(n1216),.dout(w_dff_B_p4yWtnyB7_1),.clk(gclk));
	jdff dff_B_WQkQyFdP6_1(.din(w_dff_B_p4yWtnyB7_1),.dout(w_dff_B_WQkQyFdP6_1),.clk(gclk));
	jdff dff_B_4lWuZyOJ7_1(.din(w_dff_B_WQkQyFdP6_1),.dout(w_dff_B_4lWuZyOJ7_1),.clk(gclk));
	jdff dff_B_kJQ3Yeru5_1(.din(w_dff_B_4lWuZyOJ7_1),.dout(w_dff_B_kJQ3Yeru5_1),.clk(gclk));
	jdff dff_B_IOYW8IEU2_1(.din(w_dff_B_kJQ3Yeru5_1),.dout(w_dff_B_IOYW8IEU2_1),.clk(gclk));
	jdff dff_B_QDj30bRT2_1(.din(w_dff_B_IOYW8IEU2_1),.dout(w_dff_B_QDj30bRT2_1),.clk(gclk));
	jdff dff_B_wZB3cbBV1_1(.din(w_dff_B_QDj30bRT2_1),.dout(w_dff_B_wZB3cbBV1_1),.clk(gclk));
	jdff dff_B_ArPgHb7L5_1(.din(w_dff_B_wZB3cbBV1_1),.dout(w_dff_B_ArPgHb7L5_1),.clk(gclk));
	jdff dff_B_8VZKDMGW1_1(.din(w_dff_B_ArPgHb7L5_1),.dout(w_dff_B_8VZKDMGW1_1),.clk(gclk));
	jdff dff_B_ty52Xt5r4_1(.din(w_dff_B_8VZKDMGW1_1),.dout(w_dff_B_ty52Xt5r4_1),.clk(gclk));
	jdff dff_B_oEGnkt1Y0_1(.din(w_dff_B_ty52Xt5r4_1),.dout(w_dff_B_oEGnkt1Y0_1),.clk(gclk));
	jdff dff_B_RYh6DWOm4_0(.din(n1219),.dout(w_dff_B_RYh6DWOm4_0),.clk(gclk));
	jdff dff_B_R9p2FXyb6_0(.din(w_dff_B_RYh6DWOm4_0),.dout(w_dff_B_R9p2FXyb6_0),.clk(gclk));
	jdff dff_B_UTLi8MrO5_0(.din(w_dff_B_R9p2FXyb6_0),.dout(w_dff_B_UTLi8MrO5_0),.clk(gclk));
	jdff dff_B_wkiCQYnH1_0(.din(w_dff_B_UTLi8MrO5_0),.dout(w_dff_B_wkiCQYnH1_0),.clk(gclk));
	jdff dff_B_PGKwaFuX5_0(.din(w_dff_B_wkiCQYnH1_0),.dout(w_dff_B_PGKwaFuX5_0),.clk(gclk));
	jdff dff_B_DGBkJHNe4_0(.din(w_dff_B_PGKwaFuX5_0),.dout(w_dff_B_DGBkJHNe4_0),.clk(gclk));
	jdff dff_B_Z4JsXH4x2_0(.din(w_dff_B_DGBkJHNe4_0),.dout(w_dff_B_Z4JsXH4x2_0),.clk(gclk));
	jdff dff_A_s1FilO8V2_1(.dout(w_n989_0[1]),.din(w_dff_A_s1FilO8V2_1),.clk(gclk));
	jdff dff_A_Apmot8Vw3_1(.dout(w_dff_A_s1FilO8V2_1),.din(w_dff_A_Apmot8Vw3_1),.clk(gclk));
	jdff dff_A_IC9Kw6aN7_1(.dout(w_dff_A_Apmot8Vw3_1),.din(w_dff_A_IC9Kw6aN7_1),.clk(gclk));
	jdff dff_A_lFtRrneu6_1(.dout(w_dff_A_IC9Kw6aN7_1),.din(w_dff_A_lFtRrneu6_1),.clk(gclk));
	jdff dff_A_WnRpMoNw1_1(.dout(w_dff_A_lFtRrneu6_1),.din(w_dff_A_WnRpMoNw1_1),.clk(gclk));
	jdff dff_B_76XzOmlq6_1(.din(n988),.dout(w_dff_B_76XzOmlq6_1),.clk(gclk));
	jdff dff_B_0aVmP3li7_1(.din(w_dff_B_76XzOmlq6_1),.dout(w_dff_B_0aVmP3li7_1),.clk(gclk));
	jdff dff_B_MRe0avuu7_1(.din(w_dff_B_0aVmP3li7_1),.dout(w_dff_B_MRe0avuu7_1),.clk(gclk));
	jdff dff_B_GXYEBK7E6_1(.din(w_dff_B_MRe0avuu7_1),.dout(w_dff_B_GXYEBK7E6_1),.clk(gclk));
	jdff dff_B_nLG1eGJV1_1(.din(w_dff_B_GXYEBK7E6_1),.dout(w_dff_B_nLG1eGJV1_1),.clk(gclk));
	jdff dff_B_UILrsiJX5_1(.din(w_dff_B_nLG1eGJV1_1),.dout(w_dff_B_UILrsiJX5_1),.clk(gclk));
	jdff dff_A_WYo4t0Ao5_0(.dout(w_G1691_3[0]),.din(w_dff_A_WYo4t0Ao5_0),.clk(gclk));
	jdff dff_A_AbwhbL5y8_0(.dout(w_dff_A_WYo4t0Ao5_0),.din(w_dff_A_AbwhbL5y8_0),.clk(gclk));
	jdff dff_A_rc7LdPML3_0(.dout(w_dff_A_AbwhbL5y8_0),.din(w_dff_A_rc7LdPML3_0),.clk(gclk));
	jdff dff_A_55ySoC9q4_0(.dout(w_dff_A_rc7LdPML3_0),.din(w_dff_A_55ySoC9q4_0),.clk(gclk));
	jdff dff_A_9WetyqJg1_1(.dout(w_G1691_3[1]),.din(w_dff_A_9WetyqJg1_1),.clk(gclk));
	jdff dff_A_2iyUexrb4_1(.dout(w_dff_A_9WetyqJg1_1),.din(w_dff_A_2iyUexrb4_1),.clk(gclk));
	jdff dff_B_myvVPbSd7_1(.din(n1382),.dout(w_dff_B_myvVPbSd7_1),.clk(gclk));
	jdff dff_B_GlPdXiY42_1(.din(w_dff_B_myvVPbSd7_1),.dout(w_dff_B_GlPdXiY42_1),.clk(gclk));
	jdff dff_B_aMu63uXL3_1(.din(w_dff_B_GlPdXiY42_1),.dout(w_dff_B_aMu63uXL3_1),.clk(gclk));
	jdff dff_B_YM5TZrGh1_1(.din(w_dff_B_aMu63uXL3_1),.dout(w_dff_B_YM5TZrGh1_1),.clk(gclk));
	jdff dff_B_3f3TY8vL6_1(.din(w_dff_B_YM5TZrGh1_1),.dout(w_dff_B_3f3TY8vL6_1),.clk(gclk));
	jdff dff_B_L8PaIB0r9_1(.din(w_dff_B_3f3TY8vL6_1),.dout(w_dff_B_L8PaIB0r9_1),.clk(gclk));
	jdff dff_B_FIwAXgMv5_1(.din(w_dff_B_L8PaIB0r9_1),.dout(w_dff_B_FIwAXgMv5_1),.clk(gclk));
	jdff dff_B_2GX8UCpz5_1(.din(w_dff_B_FIwAXgMv5_1),.dout(w_dff_B_2GX8UCpz5_1),.clk(gclk));
	jdff dff_B_WINLHToP6_1(.din(w_dff_B_2GX8UCpz5_1),.dout(w_dff_B_WINLHToP6_1),.clk(gclk));
	jdff dff_B_8SWCRkgH0_1(.din(w_dff_B_WINLHToP6_1),.dout(w_dff_B_8SWCRkgH0_1),.clk(gclk));
	jdff dff_B_rLIXuRet4_1(.din(w_dff_B_8SWCRkgH0_1),.dout(w_dff_B_rLIXuRet4_1),.clk(gclk));
	jdff dff_B_SeHfmNLb1_1(.din(w_dff_B_rLIXuRet4_1),.dout(w_dff_B_SeHfmNLb1_1),.clk(gclk));
	jdff dff_B_n9LEvZSr3_1(.din(w_dff_B_SeHfmNLb1_1),.dout(w_dff_B_n9LEvZSr3_1),.clk(gclk));
	jdff dff_B_8DioIkAS1_1(.din(w_dff_B_n9LEvZSr3_1),.dout(w_dff_B_8DioIkAS1_1),.clk(gclk));
	jdff dff_B_EzH0H0Dj1_1(.din(w_dff_B_8DioIkAS1_1),.dout(w_dff_B_EzH0H0Dj1_1),.clk(gclk));
	jdff dff_B_sORWbYPy7_1(.din(w_dff_B_EzH0H0Dj1_1),.dout(w_dff_B_sORWbYPy7_1),.clk(gclk));
	jdff dff_B_4TDqEHkO5_1(.din(w_dff_B_sORWbYPy7_1),.dout(w_dff_B_4TDqEHkO5_1),.clk(gclk));
	jdff dff_B_mm87ihes8_1(.din(w_dff_B_4TDqEHkO5_1),.dout(w_dff_B_mm87ihes8_1),.clk(gclk));
	jdff dff_B_VkGZTCwZ0_1(.din(w_dff_B_mm87ihes8_1),.dout(w_dff_B_VkGZTCwZ0_1),.clk(gclk));
	jdff dff_B_02ECiP6D3_1(.din(n1207),.dout(w_dff_B_02ECiP6D3_1),.clk(gclk));
	jdff dff_B_cIiDLppA7_1(.din(w_dff_B_02ECiP6D3_1),.dout(w_dff_B_cIiDLppA7_1),.clk(gclk));
	jdff dff_B_8jBPDOJG1_1(.din(w_dff_B_cIiDLppA7_1),.dout(w_dff_B_8jBPDOJG1_1),.clk(gclk));
	jdff dff_B_tneGJfTT2_1(.din(w_dff_B_8jBPDOJG1_1),.dout(w_dff_B_tneGJfTT2_1),.clk(gclk));
	jdff dff_B_TMR7AuPx0_1(.din(w_dff_B_tneGJfTT2_1),.dout(w_dff_B_TMR7AuPx0_1),.clk(gclk));
	jdff dff_B_KzbH4jb70_1(.din(w_dff_B_TMR7AuPx0_1),.dout(w_dff_B_KzbH4jb70_1),.clk(gclk));
	jdff dff_B_L68SKDEG0_1(.din(w_dff_B_KzbH4jb70_1),.dout(w_dff_B_L68SKDEG0_1),.clk(gclk));
	jdff dff_B_gzxYdMJX9_1(.din(w_dff_B_L68SKDEG0_1),.dout(w_dff_B_gzxYdMJX9_1),.clk(gclk));
	jdff dff_B_ws94ad5S2_1(.din(w_dff_B_gzxYdMJX9_1),.dout(w_dff_B_ws94ad5S2_1),.clk(gclk));
	jdff dff_B_Z5UuduDE7_1(.din(w_dff_B_ws94ad5S2_1),.dout(w_dff_B_Z5UuduDE7_1),.clk(gclk));
	jdff dff_B_lbRTFf7C9_1(.din(w_dff_B_Z5UuduDE7_1),.dout(w_dff_B_lbRTFf7C9_1),.clk(gclk));
	jdff dff_B_1l9XPtdR6_1(.din(w_dff_B_lbRTFf7C9_1),.dout(w_dff_B_1l9XPtdR6_1),.clk(gclk));
	jdff dff_B_XgoKzcAF1_1(.din(w_dff_B_1l9XPtdR6_1),.dout(w_dff_B_XgoKzcAF1_1),.clk(gclk));
	jdff dff_B_Z4VfJ3uk9_1(.din(w_dff_B_XgoKzcAF1_1),.dout(w_dff_B_Z4VfJ3uk9_1),.clk(gclk));
	jdff dff_B_SuvowPje4_1(.din(w_dff_B_Z4VfJ3uk9_1),.dout(w_dff_B_SuvowPje4_1),.clk(gclk));
	jdff dff_B_M3qIf25O9_1(.din(w_dff_B_SuvowPje4_1),.dout(w_dff_B_M3qIf25O9_1),.clk(gclk));
	jdff dff_B_WKfF4zB30_0(.din(n1211),.dout(w_dff_B_WKfF4zB30_0),.clk(gclk));
	jdff dff_B_S4fAFmOo6_0(.din(w_dff_B_WKfF4zB30_0),.dout(w_dff_B_S4fAFmOo6_0),.clk(gclk));
	jdff dff_B_9MYWyWhf2_0(.din(w_dff_B_S4fAFmOo6_0),.dout(w_dff_B_9MYWyWhf2_0),.clk(gclk));
	jdff dff_B_OUB5DwPz1_0(.din(w_dff_B_9MYWyWhf2_0),.dout(w_dff_B_OUB5DwPz1_0),.clk(gclk));
	jdff dff_B_iRXoc1t62_0(.din(w_dff_B_OUB5DwPz1_0),.dout(w_dff_B_iRXoc1t62_0),.clk(gclk));
	jdff dff_B_YdoE0Sty7_0(.din(w_dff_B_iRXoc1t62_0),.dout(w_dff_B_YdoE0Sty7_0),.clk(gclk));
	jdff dff_B_V7IvcMX07_0(.din(w_dff_B_YdoE0Sty7_0),.dout(w_dff_B_V7IvcMX07_0),.clk(gclk));
	jdff dff_B_oIpz3zf67_0(.din(w_dff_B_V7IvcMX07_0),.dout(w_dff_B_oIpz3zf67_0),.clk(gclk));
	jdff dff_B_VrvEw4Un4_0(.din(w_dff_B_oIpz3zf67_0),.dout(w_dff_B_VrvEw4Un4_0),.clk(gclk));
	jdff dff_B_AMlJ6zkX7_0(.din(w_dff_B_VrvEw4Un4_0),.dout(w_dff_B_AMlJ6zkX7_0),.clk(gclk));
	jdff dff_B_auJqx8k39_1(.din(n978),.dout(w_dff_B_auJqx8k39_1),.clk(gclk));
	jdff dff_B_Z5FXd1Xe2_1(.din(w_dff_B_auJqx8k39_1),.dout(w_dff_B_Z5FXd1Xe2_1),.clk(gclk));
	jdff dff_B_AOJviqIu3_1(.din(w_dff_B_Z5FXd1Xe2_1),.dout(w_dff_B_AOJviqIu3_1),.clk(gclk));
	jdff dff_B_PeZZZXUX1_1(.din(w_dff_B_AOJviqIu3_1),.dout(w_dff_B_PeZZZXUX1_1),.clk(gclk));
	jdff dff_B_4FJdQSby2_1(.din(w_dff_B_PeZZZXUX1_1),.dout(w_dff_B_4FJdQSby2_1),.clk(gclk));
	jdff dff_B_vCCl4NZP7_1(.din(w_dff_B_4FJdQSby2_1),.dout(w_dff_B_vCCl4NZP7_1),.clk(gclk));
	jdff dff_B_NhUoNeKe9_1(.din(w_dff_B_vCCl4NZP7_1),.dout(w_dff_B_NhUoNeKe9_1),.clk(gclk));
	jdff dff_B_U0qnV3rS4_1(.din(w_dff_B_NhUoNeKe9_1),.dout(w_dff_B_U0qnV3rS4_1),.clk(gclk));
	jdff dff_B_q3yblBT83_1(.din(w_dff_B_U0qnV3rS4_1),.dout(w_dff_B_q3yblBT83_1),.clk(gclk));
	jdff dff_B_6pLzhFzy3_1(.din(n982),.dout(w_dff_B_6pLzhFzy3_1),.clk(gclk));
	jdff dff_B_PYmBybxC3_1(.din(n980),.dout(w_dff_B_PYmBybxC3_1),.clk(gclk));
	jdff dff_B_Gt6mEJbL1_1(.din(w_dff_B_PYmBybxC3_1),.dout(w_dff_B_Gt6mEJbL1_1),.clk(gclk));
	jdff dff_B_Zy2FpPAN4_1(.din(w_dff_B_Gt6mEJbL1_1),.dout(w_dff_B_Zy2FpPAN4_1),.clk(gclk));
	jdff dff_B_ouss8ttY5_1(.din(w_dff_B_Zy2FpPAN4_1),.dout(w_dff_B_ouss8ttY5_1),.clk(gclk));
	jdff dff_B_KtJt2y784_1(.din(w_dff_B_ouss8ttY5_1),.dout(w_dff_B_KtJt2y784_1),.clk(gclk));
	jdff dff_B_6KR0qW3n2_0(.din(n1395),.dout(w_dff_B_6KR0qW3n2_0),.clk(gclk));
	jdff dff_B_P1tojrHZ4_0(.din(w_dff_B_6KR0qW3n2_0),.dout(w_dff_B_P1tojrHZ4_0),.clk(gclk));
	jdff dff_B_wMnlK9Bc6_0(.din(w_dff_B_P1tojrHZ4_0),.dout(w_dff_B_wMnlK9Bc6_0),.clk(gclk));
	jdff dff_B_x10XzrrB6_0(.din(w_dff_B_wMnlK9Bc6_0),.dout(w_dff_B_x10XzrrB6_0),.clk(gclk));
	jdff dff_B_xI8VjsDx1_0(.din(w_dff_B_x10XzrrB6_0),.dout(w_dff_B_xI8VjsDx1_0),.clk(gclk));
	jdff dff_B_0Zf1eCYS9_0(.din(w_dff_B_xI8VjsDx1_0),.dout(w_dff_B_0Zf1eCYS9_0),.clk(gclk));
	jdff dff_B_71UCjA3L0_0(.din(w_dff_B_0Zf1eCYS9_0),.dout(w_dff_B_71UCjA3L0_0),.clk(gclk));
	jdff dff_B_bjU1o1PW6_0(.din(w_dff_B_71UCjA3L0_0),.dout(w_dff_B_bjU1o1PW6_0),.clk(gclk));
	jdff dff_B_Q6MOeho38_0(.din(w_dff_B_bjU1o1PW6_0),.dout(w_dff_B_Q6MOeho38_0),.clk(gclk));
	jdff dff_B_O4NrzNrM6_0(.din(w_dff_B_Q6MOeho38_0),.dout(w_dff_B_O4NrzNrM6_0),.clk(gclk));
	jdff dff_B_nC3ScYUk1_0(.din(w_dff_B_O4NrzNrM6_0),.dout(w_dff_B_nC3ScYUk1_0),.clk(gclk));
	jdff dff_B_OIO3nJy82_0(.din(w_dff_B_nC3ScYUk1_0),.dout(w_dff_B_OIO3nJy82_0),.clk(gclk));
	jdff dff_B_tuPQzDkg2_0(.din(w_dff_B_OIO3nJy82_0),.dout(w_dff_B_tuPQzDkg2_0),.clk(gclk));
	jdff dff_B_ne1VmxbK3_0(.din(w_dff_B_tuPQzDkg2_0),.dout(w_dff_B_ne1VmxbK3_0),.clk(gclk));
	jdff dff_B_yqEFetps2_0(.din(w_dff_B_ne1VmxbK3_0),.dout(w_dff_B_yqEFetps2_0),.clk(gclk));
	jdff dff_B_Civl0PfK2_0(.din(w_dff_B_yqEFetps2_0),.dout(w_dff_B_Civl0PfK2_0),.clk(gclk));
	jdff dff_B_ppCAZ6H29_0(.din(w_dff_B_Civl0PfK2_0),.dout(w_dff_B_ppCAZ6H29_0),.clk(gclk));
	jdff dff_B_cNpLALwU9_0(.din(w_dff_B_ppCAZ6H29_0),.dout(w_dff_B_cNpLALwU9_0),.clk(gclk));
	jdff dff_B_j5DK7ZyH8_0(.din(w_dff_B_cNpLALwU9_0),.dout(w_dff_B_j5DK7ZyH8_0),.clk(gclk));
	jdff dff_B_MTWm3H7E2_1(.din(n1389),.dout(w_dff_B_MTWm3H7E2_1),.clk(gclk));
	jdff dff_B_MyNQdqJ97_1(.din(w_dff_B_MTWm3H7E2_1),.dout(w_dff_B_MyNQdqJ97_1),.clk(gclk));
	jdff dff_B_tmwvDAz70_1(.din(n1198),.dout(w_dff_B_tmwvDAz70_1),.clk(gclk));
	jdff dff_B_4BFDwHec1_1(.din(w_dff_B_tmwvDAz70_1),.dout(w_dff_B_4BFDwHec1_1),.clk(gclk));
	jdff dff_B_LPquafu73_1(.din(w_dff_B_4BFDwHec1_1),.dout(w_dff_B_LPquafu73_1),.clk(gclk));
	jdff dff_B_2JSczoHV2_1(.din(w_dff_B_LPquafu73_1),.dout(w_dff_B_2JSczoHV2_1),.clk(gclk));
	jdff dff_B_paZagDH31_1(.din(w_dff_B_2JSczoHV2_1),.dout(w_dff_B_paZagDH31_1),.clk(gclk));
	jdff dff_B_acv8bJlo5_1(.din(w_dff_B_paZagDH31_1),.dout(w_dff_B_acv8bJlo5_1),.clk(gclk));
	jdff dff_B_zE3SP0cj1_1(.din(w_dff_B_acv8bJlo5_1),.dout(w_dff_B_zE3SP0cj1_1),.clk(gclk));
	jdff dff_B_drglUFN87_1(.din(w_dff_B_zE3SP0cj1_1),.dout(w_dff_B_drglUFN87_1),.clk(gclk));
	jdff dff_B_pwSHXP8X2_1(.din(w_dff_B_drglUFN87_1),.dout(w_dff_B_pwSHXP8X2_1),.clk(gclk));
	jdff dff_B_oMreKgB77_1(.din(w_dff_B_pwSHXP8X2_1),.dout(w_dff_B_oMreKgB77_1),.clk(gclk));
	jdff dff_B_ENz6bOd40_1(.din(w_dff_B_oMreKgB77_1),.dout(w_dff_B_ENz6bOd40_1),.clk(gclk));
	jdff dff_B_2hUhRn792_1(.din(w_dff_B_ENz6bOd40_1),.dout(w_dff_B_2hUhRn792_1),.clk(gclk));
	jdff dff_B_55ngfZWA2_1(.din(w_dff_B_2hUhRn792_1),.dout(w_dff_B_55ngfZWA2_1),.clk(gclk));
	jdff dff_B_EBtMAoV48_1(.din(w_dff_B_55ngfZWA2_1),.dout(w_dff_B_EBtMAoV48_1),.clk(gclk));
	jdff dff_B_bArBZE0s8_1(.din(w_dff_B_EBtMAoV48_1),.dout(w_dff_B_bArBZE0s8_1),.clk(gclk));
	jdff dff_B_UwkZLPuQ0_1(.din(n1200),.dout(w_dff_B_UwkZLPuQ0_1),.clk(gclk));
	jdff dff_B_8c3WVdlW9_1(.din(w_dff_B_UwkZLPuQ0_1),.dout(w_dff_B_8c3WVdlW9_1),.clk(gclk));
	jdff dff_B_6i5RmBAb4_1(.din(w_dff_B_8c3WVdlW9_1),.dout(w_dff_B_6i5RmBAb4_1),.clk(gclk));
	jdff dff_B_Urhfa7Ty2_1(.din(w_dff_B_6i5RmBAb4_1),.dout(w_dff_B_Urhfa7Ty2_1),.clk(gclk));
	jdff dff_B_2eHnOBm39_1(.din(w_dff_B_Urhfa7Ty2_1),.dout(w_dff_B_2eHnOBm39_1),.clk(gclk));
	jdff dff_B_J0pQXekf9_1(.din(w_dff_B_2eHnOBm39_1),.dout(w_dff_B_J0pQXekf9_1),.clk(gclk));
	jdff dff_B_g2lPKBsA1_1(.din(w_dff_B_J0pQXekf9_1),.dout(w_dff_B_g2lPKBsA1_1),.clk(gclk));
	jdff dff_B_S2egDuPP7_1(.din(w_dff_B_g2lPKBsA1_1),.dout(w_dff_B_S2egDuPP7_1),.clk(gclk));
	jdff dff_B_3sYPQFlP3_1(.din(w_dff_B_S2egDuPP7_1),.dout(w_dff_B_3sYPQFlP3_1),.clk(gclk));
	jdff dff_B_fxewUeBb5_1(.din(w_dff_B_3sYPQFlP3_1),.dout(w_dff_B_fxewUeBb5_1),.clk(gclk));
	jdff dff_B_HLuv4sqU8_1(.din(w_dff_B_fxewUeBb5_1),.dout(w_dff_B_HLuv4sqU8_1),.clk(gclk));
	jdff dff_A_gzOtYmBM1_0(.dout(w_n649_0[0]),.din(w_dff_A_gzOtYmBM1_0),.clk(gclk));
	jdff dff_A_gS3Eofon3_0(.dout(w_dff_A_gzOtYmBM1_0),.din(w_dff_A_gS3Eofon3_0),.clk(gclk));
	jdff dff_A_P2eVeULF3_0(.dout(w_dff_A_gS3Eofon3_0),.din(w_dff_A_P2eVeULF3_0),.clk(gclk));
	jdff dff_A_nn4ttwY30_0(.dout(w_dff_A_P2eVeULF3_0),.din(w_dff_A_nn4ttwY30_0),.clk(gclk));
	jdff dff_A_4rwhmoIk3_0(.dout(w_dff_A_nn4ttwY30_0),.din(w_dff_A_4rwhmoIk3_0),.clk(gclk));
	jdff dff_A_gXwNeGG20_0(.dout(w_dff_A_4rwhmoIk3_0),.din(w_dff_A_gXwNeGG20_0),.clk(gclk));
	jdff dff_A_BDFNMZel4_0(.dout(w_dff_A_gXwNeGG20_0),.din(w_dff_A_BDFNMZel4_0),.clk(gclk));
	jdff dff_A_LPflsroB5_0(.dout(w_dff_A_BDFNMZel4_0),.din(w_dff_A_LPflsroB5_0),.clk(gclk));
	jdff dff_A_To32fPpX3_0(.dout(w_dff_A_LPflsroB5_0),.din(w_dff_A_To32fPpX3_0),.clk(gclk));
	jdff dff_A_2eqtmcpk1_0(.dout(w_G137_4[0]),.din(w_dff_A_2eqtmcpk1_0),.clk(gclk));
	jdff dff_A_XR3oOArB3_1(.dout(w_G137_4[1]),.din(w_dff_A_XR3oOArB3_1),.clk(gclk));
	jdff dff_A_G7amS7XX3_0(.dout(w_G137_1[0]),.din(w_dff_A_G7amS7XX3_0),.clk(gclk));
	jdff dff_A_pbfR3EOA6_0(.dout(w_dff_A_G7amS7XX3_0),.din(w_dff_A_pbfR3EOA6_0),.clk(gclk));
	jdff dff_A_BbXgFDnt3_0(.dout(w_dff_A_pbfR3EOA6_0),.din(w_dff_A_BbXgFDnt3_0),.clk(gclk));
	jdff dff_A_O0QeAVG97_0(.dout(w_dff_A_BbXgFDnt3_0),.din(w_dff_A_O0QeAVG97_0),.clk(gclk));
	jdff dff_A_depvRx9i3_0(.dout(w_dff_A_O0QeAVG97_0),.din(w_dff_A_depvRx9i3_0),.clk(gclk));
	jdff dff_A_x9nhREvs5_0(.dout(w_dff_A_depvRx9i3_0),.din(w_dff_A_x9nhREvs5_0),.clk(gclk));
	jdff dff_A_IWURhLYv1_1(.dout(w_G137_1[1]),.din(w_dff_A_IWURhLYv1_1),.clk(gclk));
	jdff dff_A_gACeJiaX0_1(.dout(w_dff_A_IWURhLYv1_1),.din(w_dff_A_gACeJiaX0_1),.clk(gclk));
	jdff dff_A_syYjlyYb9_1(.dout(w_dff_A_gACeJiaX0_1),.din(w_dff_A_syYjlyYb9_1),.clk(gclk));
	jdff dff_A_rtE8NXtz0_1(.dout(w_dff_A_syYjlyYb9_1),.din(w_dff_A_rtE8NXtz0_1),.clk(gclk));
	jdff dff_A_Ypq6KGFq9_1(.dout(w_dff_A_rtE8NXtz0_1),.din(w_dff_A_Ypq6KGFq9_1),.clk(gclk));
	jdff dff_A_Tpl2WCYT4_1(.dout(w_dff_A_Ypq6KGFq9_1),.din(w_dff_A_Tpl2WCYT4_1),.clk(gclk));
	jdff dff_A_2ZM4WqgQ8_1(.dout(w_dff_A_Tpl2WCYT4_1),.din(w_dff_A_2ZM4WqgQ8_1),.clk(gclk));
	jdff dff_B_2ZLJ7NYe7_0(.din(n1404),.dout(w_dff_B_2ZLJ7NYe7_0),.clk(gclk));
	jdff dff_B_uBTTkax61_0(.din(w_dff_B_2ZLJ7NYe7_0),.dout(w_dff_B_uBTTkax61_0),.clk(gclk));
	jdff dff_B_oCnSXvnh7_0(.din(w_dff_B_uBTTkax61_0),.dout(w_dff_B_oCnSXvnh7_0),.clk(gclk));
	jdff dff_B_v1hnzv5y0_0(.din(w_dff_B_oCnSXvnh7_0),.dout(w_dff_B_v1hnzv5y0_0),.clk(gclk));
	jdff dff_B_LlDicOws2_0(.din(w_dff_B_v1hnzv5y0_0),.dout(w_dff_B_LlDicOws2_0),.clk(gclk));
	jdff dff_B_07lxF3nb9_0(.din(w_dff_B_LlDicOws2_0),.dout(w_dff_B_07lxF3nb9_0),.clk(gclk));
	jdff dff_B_6Cb1L1au1_0(.din(w_dff_B_07lxF3nb9_0),.dout(w_dff_B_6Cb1L1au1_0),.clk(gclk));
	jdff dff_B_mAskDXiv5_0(.din(w_dff_B_6Cb1L1au1_0),.dout(w_dff_B_mAskDXiv5_0),.clk(gclk));
	jdff dff_B_Xu8XUfAu2_0(.din(w_dff_B_mAskDXiv5_0),.dout(w_dff_B_Xu8XUfAu2_0),.clk(gclk));
	jdff dff_B_0ZEJd4oe8_0(.din(w_dff_B_Xu8XUfAu2_0),.dout(w_dff_B_0ZEJd4oe8_0),.clk(gclk));
	jdff dff_B_7ISTpVOO4_0(.din(w_dff_B_0ZEJd4oe8_0),.dout(w_dff_B_7ISTpVOO4_0),.clk(gclk));
	jdff dff_B_Wl5DfmZW0_0(.din(w_dff_B_7ISTpVOO4_0),.dout(w_dff_B_Wl5DfmZW0_0),.clk(gclk));
	jdff dff_B_8UJhFz3S7_0(.din(w_dff_B_Wl5DfmZW0_0),.dout(w_dff_B_8UJhFz3S7_0),.clk(gclk));
	jdff dff_B_7e9tf7xK5_0(.din(w_dff_B_8UJhFz3S7_0),.dout(w_dff_B_7e9tf7xK5_0),.clk(gclk));
	jdff dff_B_ct5tzXPR4_0(.din(w_dff_B_7e9tf7xK5_0),.dout(w_dff_B_ct5tzXPR4_0),.clk(gclk));
	jdff dff_B_uOohp7LV9_0(.din(w_dff_B_ct5tzXPR4_0),.dout(w_dff_B_uOohp7LV9_0),.clk(gclk));
	jdff dff_B_UYuDaZAK2_0(.din(w_dff_B_uOohp7LV9_0),.dout(w_dff_B_UYuDaZAK2_0),.clk(gclk));
	jdff dff_B_rvhzNEDX1_0(.din(w_dff_B_UYuDaZAK2_0),.dout(w_dff_B_rvhzNEDX1_0),.clk(gclk));
	jdff dff_B_FNMQBBlP1_0(.din(w_dff_B_rvhzNEDX1_0),.dout(w_dff_B_FNMQBBlP1_0),.clk(gclk));
	jdff dff_B_ooJGcptk8_1(.din(n1190),.dout(w_dff_B_ooJGcptk8_1),.clk(gclk));
	jdff dff_B_9CqpIqcP7_1(.din(w_dff_B_ooJGcptk8_1),.dout(w_dff_B_9CqpIqcP7_1),.clk(gclk));
	jdff dff_B_vIhROdJC9_1(.din(w_dff_B_9CqpIqcP7_1),.dout(w_dff_B_vIhROdJC9_1),.clk(gclk));
	jdff dff_B_O0o0c5Bu4_1(.din(w_dff_B_vIhROdJC9_1),.dout(w_dff_B_O0o0c5Bu4_1),.clk(gclk));
	jdff dff_B_hvggMN5O5_1(.din(w_dff_B_O0o0c5Bu4_1),.dout(w_dff_B_hvggMN5O5_1),.clk(gclk));
	jdff dff_B_RusAHTLs7_1(.din(w_dff_B_hvggMN5O5_1),.dout(w_dff_B_RusAHTLs7_1),.clk(gclk));
	jdff dff_B_tMxI4zBR4_1(.din(w_dff_B_RusAHTLs7_1),.dout(w_dff_B_tMxI4zBR4_1),.clk(gclk));
	jdff dff_B_rSccarmi8_1(.din(w_dff_B_tMxI4zBR4_1),.dout(w_dff_B_rSccarmi8_1),.clk(gclk));
	jdff dff_B_r0OYv9tN8_1(.din(w_dff_B_rSccarmi8_1),.dout(w_dff_B_r0OYv9tN8_1),.clk(gclk));
	jdff dff_B_g39610bw8_1(.din(w_dff_B_r0OYv9tN8_1),.dout(w_dff_B_g39610bw8_1),.clk(gclk));
	jdff dff_B_6uiVvotc0_1(.din(w_dff_B_g39610bw8_1),.dout(w_dff_B_6uiVvotc0_1),.clk(gclk));
	jdff dff_B_5f4B6GHy7_1(.din(w_dff_B_6uiVvotc0_1),.dout(w_dff_B_5f4B6GHy7_1),.clk(gclk));
	jdff dff_B_QW6eZToC4_1(.din(w_dff_B_5f4B6GHy7_1),.dout(w_dff_B_QW6eZToC4_1),.clk(gclk));
	jdff dff_B_zBUb8bse1_1(.din(w_dff_B_QW6eZToC4_1),.dout(w_dff_B_zBUb8bse1_1),.clk(gclk));
	jdff dff_B_b9b6f4gL0_1(.din(w_dff_B_zBUb8bse1_1),.dout(w_dff_B_b9b6f4gL0_1),.clk(gclk));
	jdff dff_B_3D7jzu8O1_1(.din(w_dff_B_b9b6f4gL0_1),.dout(w_dff_B_3D7jzu8O1_1),.clk(gclk));
	jdff dff_B_NQuquT6l6_0(.din(n1194),.dout(w_dff_B_NQuquT6l6_0),.clk(gclk));
	jdff dff_B_NxCGFaZD2_0(.din(w_dff_B_NQuquT6l6_0),.dout(w_dff_B_NxCGFaZD2_0),.clk(gclk));
	jdff dff_B_etRqYYem7_0(.din(w_dff_B_NxCGFaZD2_0),.dout(w_dff_B_etRqYYem7_0),.clk(gclk));
	jdff dff_B_Des77N1z8_0(.din(w_dff_B_etRqYYem7_0),.dout(w_dff_B_Des77N1z8_0),.clk(gclk));
	jdff dff_B_tqeZaejH9_0(.din(w_dff_B_Des77N1z8_0),.dout(w_dff_B_tqeZaejH9_0),.clk(gclk));
	jdff dff_B_OPvJpz5I7_0(.din(w_dff_B_tqeZaejH9_0),.dout(w_dff_B_OPvJpz5I7_0),.clk(gclk));
	jdff dff_B_nlz3gFFR6_0(.din(w_dff_B_OPvJpz5I7_0),.dout(w_dff_B_nlz3gFFR6_0),.clk(gclk));
	jdff dff_B_7WiQ2i248_0(.din(w_dff_B_nlz3gFFR6_0),.dout(w_dff_B_7WiQ2i248_0),.clk(gclk));
	jdff dff_B_IE3mTKN15_0(.din(w_dff_B_7WiQ2i248_0),.dout(w_dff_B_IE3mTKN15_0),.clk(gclk));
	jdff dff_B_ihkLqLvt3_0(.din(w_dff_B_IE3mTKN15_0),.dout(w_dff_B_ihkLqLvt3_0),.clk(gclk));
	jdff dff_B_9BEy8dXA3_0(.din(w_dff_B_ihkLqLvt3_0),.dout(w_dff_B_9BEy8dXA3_0),.clk(gclk));
	jdff dff_B_zoa86Shm5_0(.din(w_dff_B_9BEy8dXA3_0),.dout(w_dff_B_zoa86Shm5_0),.clk(gclk));
	jdff dff_B_4xUKJLD13_0(.din(n794),.dout(w_dff_B_4xUKJLD13_0),.clk(gclk));
	jdff dff_B_6f5qogMe0_0(.din(n785),.dout(w_dff_B_6f5qogMe0_0),.clk(gclk));
	jdff dff_A_HRL9jvSt8_0(.dout(w_G1691_2[0]),.din(w_dff_A_HRL9jvSt8_0),.clk(gclk));
	jdff dff_A_JgzjklZa3_2(.dout(w_G1691_2[2]),.din(w_dff_A_JgzjklZa3_2),.clk(gclk));
	jdff dff_A_o4xpqt266_2(.dout(w_n1007_1[2]),.din(w_dff_A_o4xpqt266_2),.clk(gclk));
	jdff dff_A_TuZO65Nc5_0(.dout(w_n1007_0[0]),.din(w_dff_A_TuZO65Nc5_0),.clk(gclk));
	jdff dff_A_mohINigu2_0(.dout(w_dff_A_TuZO65Nc5_0),.din(w_dff_A_mohINigu2_0),.clk(gclk));
	jdff dff_A_GoHp2ciy6_0(.dout(w_dff_A_mohINigu2_0),.din(w_dff_A_GoHp2ciy6_0),.clk(gclk));
	jdff dff_A_X7HYLeqh9_0(.dout(w_dff_A_GoHp2ciy6_0),.din(w_dff_A_X7HYLeqh9_0),.clk(gclk));
	jdff dff_A_VSkI485R4_0(.dout(w_dff_A_X7HYLeqh9_0),.din(w_dff_A_VSkI485R4_0),.clk(gclk));
	jdff dff_A_67Cq9LhJ9_0(.dout(w_dff_A_VSkI485R4_0),.din(w_dff_A_67Cq9LhJ9_0),.clk(gclk));
	jdff dff_A_cdyTpUGQ7_0(.dout(w_dff_A_67Cq9LhJ9_0),.din(w_dff_A_cdyTpUGQ7_0),.clk(gclk));
	jdff dff_A_A7G5W8cI1_0(.dout(w_dff_A_cdyTpUGQ7_0),.din(w_dff_A_A7G5W8cI1_0),.clk(gclk));
	jdff dff_A_X5ele9mj2_0(.dout(w_dff_A_A7G5W8cI1_0),.din(w_dff_A_X5ele9mj2_0),.clk(gclk));
	jdff dff_A_vMs6C9cH4_1(.dout(w_n1007_0[1]),.din(w_dff_A_vMs6C9cH4_1),.clk(gclk));
	jdff dff_A_nRJ4LMDu5_1(.dout(w_dff_A_vMs6C9cH4_1),.din(w_dff_A_nRJ4LMDu5_1),.clk(gclk));
	jdff dff_B_B6msR1jS2_3(.din(n1007),.dout(w_dff_B_B6msR1jS2_3),.clk(gclk));
	jdff dff_B_IBMPP6gy4_3(.din(w_dff_B_B6msR1jS2_3),.dout(w_dff_B_IBMPP6gy4_3),.clk(gclk));
	jdff dff_B_WRqTiJIW3_3(.din(w_dff_B_IBMPP6gy4_3),.dout(w_dff_B_WRqTiJIW3_3),.clk(gclk));
	jdff dff_B_39zhnG930_3(.din(w_dff_B_WRqTiJIW3_3),.dout(w_dff_B_39zhnG930_3),.clk(gclk));
	jdff dff_B_YLTODweL4_3(.din(w_dff_B_39zhnG930_3),.dout(w_dff_B_YLTODweL4_3),.clk(gclk));
	jdff dff_B_JiPs2Uey3_3(.din(w_dff_B_YLTODweL4_3),.dout(w_dff_B_JiPs2Uey3_3),.clk(gclk));
	jdff dff_B_tcAAeZDE9_3(.din(w_dff_B_JiPs2Uey3_3),.dout(w_dff_B_tcAAeZDE9_3),.clk(gclk));
	jdff dff_B_ErmE05f45_3(.din(w_dff_B_tcAAeZDE9_3),.dout(w_dff_B_ErmE05f45_3),.clk(gclk));
	jdff dff_B_iD6VkauB9_3(.din(w_dff_B_ErmE05f45_3),.dout(w_dff_B_iD6VkauB9_3),.clk(gclk));
	jdff dff_B_bCwz9kcY5_3(.din(w_dff_B_iD6VkauB9_3),.dout(w_dff_B_bCwz9kcY5_3),.clk(gclk));
	jdff dff_B_ilgOphnQ3_3(.din(w_dff_B_bCwz9kcY5_3),.dout(w_dff_B_ilgOphnQ3_3),.clk(gclk));
	jdff dff_B_amnl6vVa9_0(.din(n1505),.dout(w_dff_B_amnl6vVa9_0),.clk(gclk));
	jdff dff_B_UgiRTvBr2_0(.din(w_dff_B_amnl6vVa9_0),.dout(w_dff_B_UgiRTvBr2_0),.clk(gclk));
	jdff dff_B_6dnbct4N1_0(.din(w_dff_B_UgiRTvBr2_0),.dout(w_dff_B_6dnbct4N1_0),.clk(gclk));
	jdff dff_B_bHUa4NyD8_0(.din(w_dff_B_6dnbct4N1_0),.dout(w_dff_B_bHUa4NyD8_0),.clk(gclk));
	jdff dff_B_jMgib4gx2_0(.din(w_dff_B_bHUa4NyD8_0),.dout(w_dff_B_jMgib4gx2_0),.clk(gclk));
	jdff dff_B_GsWcKexc1_0(.din(w_dff_B_jMgib4gx2_0),.dout(w_dff_B_GsWcKexc1_0),.clk(gclk));
	jdff dff_B_yOalO2bq8_0(.din(w_dff_B_GsWcKexc1_0),.dout(w_dff_B_yOalO2bq8_0),.clk(gclk));
	jdff dff_B_qgMjZx972_0(.din(w_dff_B_yOalO2bq8_0),.dout(w_dff_B_qgMjZx972_0),.clk(gclk));
	jdff dff_B_NrmhjzzI0_0(.din(w_dff_B_qgMjZx972_0),.dout(w_dff_B_NrmhjzzI0_0),.clk(gclk));
	jdff dff_B_EA9YhuCd8_0(.din(w_dff_B_NrmhjzzI0_0),.dout(w_dff_B_EA9YhuCd8_0),.clk(gclk));
	jdff dff_B_dlEDUn5B4_0(.din(w_dff_B_EA9YhuCd8_0),.dout(w_dff_B_dlEDUn5B4_0),.clk(gclk));
	jdff dff_B_O4dvStjK1_0(.din(w_dff_B_dlEDUn5B4_0),.dout(w_dff_B_O4dvStjK1_0),.clk(gclk));
	jdff dff_B_mlEKmy3i0_0(.din(w_dff_B_O4dvStjK1_0),.dout(w_dff_B_mlEKmy3i0_0),.clk(gclk));
	jdff dff_B_14vUnwef5_0(.din(w_dff_B_mlEKmy3i0_0),.dout(w_dff_B_14vUnwef5_0),.clk(gclk));
	jdff dff_B_BkagvVka9_0(.din(w_dff_B_14vUnwef5_0),.dout(w_dff_B_BkagvVka9_0),.clk(gclk));
	jdff dff_B_MVrJ394e1_0(.din(w_dff_B_BkagvVka9_0),.dout(w_dff_B_MVrJ394e1_0),.clk(gclk));
	jdff dff_B_sLrBGO7P3_0(.din(w_dff_B_MVrJ394e1_0),.dout(w_dff_B_sLrBGO7P3_0),.clk(gclk));
	jdff dff_B_WYnrzB081_0(.din(n1666),.dout(w_dff_B_WYnrzB081_0),.clk(gclk));
	jdff dff_B_cefAZnSV1_0(.din(w_dff_B_WYnrzB081_0),.dout(w_dff_B_cefAZnSV1_0),.clk(gclk));
	jdff dff_B_VXfN6Rxl6_0(.din(w_dff_B_cefAZnSV1_0),.dout(w_dff_B_VXfN6Rxl6_0),.clk(gclk));
	jdff dff_B_WPf0VP3U1_0(.din(w_dff_B_VXfN6Rxl6_0),.dout(w_dff_B_WPf0VP3U1_0),.clk(gclk));
	jdff dff_B_QbfSDge96_0(.din(w_dff_B_WPf0VP3U1_0),.dout(w_dff_B_QbfSDge96_0),.clk(gclk));
	jdff dff_B_tsAkeTqc0_0(.din(w_dff_B_QbfSDge96_0),.dout(w_dff_B_tsAkeTqc0_0),.clk(gclk));
	jdff dff_B_ICqstP6q0_0(.din(w_dff_B_tsAkeTqc0_0),.dout(w_dff_B_ICqstP6q0_0),.clk(gclk));
	jdff dff_B_Rt9wbP2j2_0(.din(w_dff_B_ICqstP6q0_0),.dout(w_dff_B_Rt9wbP2j2_0),.clk(gclk));
	jdff dff_B_TIVDoktD9_0(.din(w_dff_B_Rt9wbP2j2_0),.dout(w_dff_B_TIVDoktD9_0),.clk(gclk));
	jdff dff_B_ajr3RozC7_0(.din(w_dff_B_TIVDoktD9_0),.dout(w_dff_B_ajr3RozC7_0),.clk(gclk));
	jdff dff_B_4rw2JdVK8_0(.din(w_dff_B_ajr3RozC7_0),.dout(w_dff_B_4rw2JdVK8_0),.clk(gclk));
	jdff dff_B_ku1WFQUH9_0(.din(w_dff_B_4rw2JdVK8_0),.dout(w_dff_B_ku1WFQUH9_0),.clk(gclk));
	jdff dff_B_LWtLpZwX1_0(.din(w_dff_B_ku1WFQUH9_0),.dout(w_dff_B_LWtLpZwX1_0),.clk(gclk));
	jdff dff_B_SVQGD7k93_0(.din(w_dff_B_LWtLpZwX1_0),.dout(w_dff_B_SVQGD7k93_0),.clk(gclk));
	jdff dff_B_QnczFIBi2_0(.din(w_dff_B_SVQGD7k93_0),.dout(w_dff_B_QnczFIBi2_0),.clk(gclk));
	jdff dff_B_DMV76sid3_0(.din(w_dff_B_QnczFIBi2_0),.dout(w_dff_B_DMV76sid3_0),.clk(gclk));
	jdff dff_B_shEHb3tA0_0(.din(w_dff_B_DMV76sid3_0),.dout(w_dff_B_shEHb3tA0_0),.clk(gclk));
	jdff dff_B_5MBjdzIM7_1(.din(n1671),.dout(w_dff_B_5MBjdzIM7_1),.clk(gclk));
	jdff dff_B_WOsrwc1U7_1(.din(w_dff_B_5MBjdzIM7_1),.dout(w_dff_B_WOsrwc1U7_1),.clk(gclk));
	jdff dff_B_R8Mb56158_1(.din(w_dff_B_WOsrwc1U7_1),.dout(w_dff_B_R8Mb56158_1),.clk(gclk));
	jdff dff_B_RcASiONo7_1(.din(w_dff_B_R8Mb56158_1),.dout(w_dff_B_RcASiONo7_1),.clk(gclk));
	jdff dff_B_QyonVpYp2_1(.din(w_dff_B_RcASiONo7_1),.dout(w_dff_B_QyonVpYp2_1),.clk(gclk));
	jdff dff_B_pdZk2Oli6_1(.din(w_dff_B_QyonVpYp2_1),.dout(w_dff_B_pdZk2Oli6_1),.clk(gclk));
	jdff dff_B_H5v8wQ9J8_1(.din(w_dff_B_pdZk2Oli6_1),.dout(w_dff_B_H5v8wQ9J8_1),.clk(gclk));
	jdff dff_B_GxQiWWLU4_1(.din(w_dff_B_H5v8wQ9J8_1),.dout(w_dff_B_GxQiWWLU4_1),.clk(gclk));
	jdff dff_B_qWF2oG3R3_1(.din(w_dff_B_GxQiWWLU4_1),.dout(w_dff_B_qWF2oG3R3_1),.clk(gclk));
	jdff dff_B_ENOlmBFP4_1(.din(w_dff_B_qWF2oG3R3_1),.dout(w_dff_B_ENOlmBFP4_1),.clk(gclk));
	jdff dff_B_D5AQM6tC9_1(.din(w_dff_B_ENOlmBFP4_1),.dout(w_dff_B_D5AQM6tC9_1),.clk(gclk));
	jdff dff_B_fjmZhyw96_1(.din(w_dff_B_D5AQM6tC9_1),.dout(w_dff_B_fjmZhyw96_1),.clk(gclk));
	jdff dff_B_2LjtTI2E8_1(.din(w_dff_B_fjmZhyw96_1),.dout(w_dff_B_2LjtTI2E8_1),.clk(gclk));
	jdff dff_B_4JCscMMW8_1(.din(w_dff_B_2LjtTI2E8_1),.dout(w_dff_B_4JCscMMW8_1),.clk(gclk));
	jdff dff_B_JeoGxJYG0_1(.din(w_dff_B_4JCscMMW8_1),.dout(w_dff_B_JeoGxJYG0_1),.clk(gclk));
	jdff dff_B_IkB6CCCa3_1(.din(w_dff_B_JeoGxJYG0_1),.dout(w_dff_B_IkB6CCCa3_1),.clk(gclk));
	jdff dff_B_KzMwOGDP0_1(.din(w_dff_B_IkB6CCCa3_1),.dout(w_dff_B_KzMwOGDP0_1),.clk(gclk));
	jdff dff_B_C4opgz5m0_1(.din(w_dff_B_KzMwOGDP0_1),.dout(w_dff_B_C4opgz5m0_1),.clk(gclk));
	jdff dff_B_SfarNTi77_1(.din(w_dff_B_C4opgz5m0_1),.dout(w_dff_B_SfarNTi77_1),.clk(gclk));
	jdff dff_B_AH4fPRSj2_1(.din(w_dff_B_SfarNTi77_1),.dout(w_dff_B_AH4fPRSj2_1),.clk(gclk));
	jdff dff_B_MF4eaZkD4_1(.din(w_dff_B_AH4fPRSj2_1),.dout(w_dff_B_MF4eaZkD4_1),.clk(gclk));
	jdff dff_B_MSftF2H93_1(.din(w_dff_B_MF4eaZkD4_1),.dout(w_dff_B_MSftF2H93_1),.clk(gclk));
	jdff dff_B_EEzYRZkM4_1(.din(n1676),.dout(w_dff_B_EEzYRZkM4_1),.clk(gclk));
	jdff dff_A_RHfzNSPg1_1(.dout(w_n800_1[1]),.din(w_dff_A_RHfzNSPg1_1),.clk(gclk));
	jdff dff_A_rystDuU95_1(.dout(w_dff_A_RHfzNSPg1_1),.din(w_dff_A_rystDuU95_1),.clk(gclk));
	jdff dff_A_zbA8LNwf7_1(.dout(w_dff_A_rystDuU95_1),.din(w_dff_A_zbA8LNwf7_1),.clk(gclk));
	jdff dff_A_5VbY4wKc4_1(.dout(w_dff_A_zbA8LNwf7_1),.din(w_dff_A_5VbY4wKc4_1),.clk(gclk));
	jdff dff_A_ZzkiHjCq1_1(.dout(w_dff_A_5VbY4wKc4_1),.din(w_dff_A_ZzkiHjCq1_1),.clk(gclk));
	jdff dff_A_VIeei1bg2_1(.dout(w_dff_A_ZzkiHjCq1_1),.din(w_dff_A_VIeei1bg2_1),.clk(gclk));
	jdff dff_A_i1Jer8HA9_1(.dout(w_dff_A_VIeei1bg2_1),.din(w_dff_A_i1Jer8HA9_1),.clk(gclk));
	jdff dff_A_vKxGeqiP9_1(.dout(w_dff_A_i1Jer8HA9_1),.din(w_dff_A_vKxGeqiP9_1),.clk(gclk));
	jdff dff_A_9ms7kQtp6_1(.dout(w_dff_A_vKxGeqiP9_1),.din(w_dff_A_9ms7kQtp6_1),.clk(gclk));
	jdff dff_A_DOF0jgwQ0_1(.dout(w_dff_A_9ms7kQtp6_1),.din(w_dff_A_DOF0jgwQ0_1),.clk(gclk));
	jdff dff_A_9bemO3lg7_1(.dout(w_dff_A_DOF0jgwQ0_1),.din(w_dff_A_9bemO3lg7_1),.clk(gclk));
	jdff dff_A_cOifCqaX4_1(.dout(w_dff_A_9bemO3lg7_1),.din(w_dff_A_cOifCqaX4_1),.clk(gclk));
	jdff dff_A_4GGle7XC4_1(.dout(w_dff_A_cOifCqaX4_1),.din(w_dff_A_4GGle7XC4_1),.clk(gclk));
	jdff dff_A_rW7yqhoM0_1(.dout(w_dff_A_4GGle7XC4_1),.din(w_dff_A_rW7yqhoM0_1),.clk(gclk));
	jdff dff_A_9uD4KlcF1_2(.dout(w_n800_1[2]),.din(w_dff_A_9uD4KlcF1_2),.clk(gclk));
	jdff dff_A_eriU6EEM6_2(.dout(w_dff_A_9uD4KlcF1_2),.din(w_dff_A_eriU6EEM6_2),.clk(gclk));
	jdff dff_A_PM4ciDnd2_2(.dout(w_dff_A_eriU6EEM6_2),.din(w_dff_A_PM4ciDnd2_2),.clk(gclk));
	jdff dff_A_zhNNRsm78_2(.dout(w_dff_A_PM4ciDnd2_2),.din(w_dff_A_zhNNRsm78_2),.clk(gclk));
	jdff dff_A_C9Tsq5js6_2(.dout(w_dff_A_zhNNRsm78_2),.din(w_dff_A_C9Tsq5js6_2),.clk(gclk));
	jdff dff_A_yRGbStaz4_2(.dout(w_dff_A_C9Tsq5js6_2),.din(w_dff_A_yRGbStaz4_2),.clk(gclk));
	jdff dff_A_YrGbzQji2_2(.dout(w_dff_A_yRGbStaz4_2),.din(w_dff_A_YrGbzQji2_2),.clk(gclk));
	jdff dff_A_JOxejTlT8_2(.dout(w_dff_A_YrGbzQji2_2),.din(w_dff_A_JOxejTlT8_2),.clk(gclk));
	jdff dff_A_ixhmkYSC6_2(.dout(w_dff_A_JOxejTlT8_2),.din(w_dff_A_ixhmkYSC6_2),.clk(gclk));
	jdff dff_A_fW8OGSka8_2(.dout(w_dff_A_ixhmkYSC6_2),.din(w_dff_A_fW8OGSka8_2),.clk(gclk));
	jdff dff_B_zJcJ2KQI2_1(.din(n1688),.dout(w_dff_B_zJcJ2KQI2_1),.clk(gclk));
	jdff dff_B_5MYgQLxb5_1(.din(w_dff_B_zJcJ2KQI2_1),.dout(w_dff_B_5MYgQLxb5_1),.clk(gclk));
	jdff dff_B_NddqbPXm3_1(.din(w_dff_B_5MYgQLxb5_1),.dout(w_dff_B_NddqbPXm3_1),.clk(gclk));
	jdff dff_B_9Tgjv4SM2_1(.din(w_dff_B_NddqbPXm3_1),.dout(w_dff_B_9Tgjv4SM2_1),.clk(gclk));
	jdff dff_B_9IuPFjWc3_1(.din(w_dff_B_9Tgjv4SM2_1),.dout(w_dff_B_9IuPFjWc3_1),.clk(gclk));
	jdff dff_B_f6Jh1WVy9_1(.din(w_dff_B_9IuPFjWc3_1),.dout(w_dff_B_f6Jh1WVy9_1),.clk(gclk));
	jdff dff_B_UydghEbs2_1(.din(w_dff_B_f6Jh1WVy9_1),.dout(w_dff_B_UydghEbs2_1),.clk(gclk));
	jdff dff_B_UNhxR9L72_1(.din(w_dff_B_UydghEbs2_1),.dout(w_dff_B_UNhxR9L72_1),.clk(gclk));
	jdff dff_B_shbRryZK9_1(.din(w_dff_B_UNhxR9L72_1),.dout(w_dff_B_shbRryZK9_1),.clk(gclk));
	jdff dff_B_aM4m7D2d8_1(.din(w_dff_B_shbRryZK9_1),.dout(w_dff_B_aM4m7D2d8_1),.clk(gclk));
	jdff dff_B_iluRJHjN2_1(.din(w_dff_B_aM4m7D2d8_1),.dout(w_dff_B_iluRJHjN2_1),.clk(gclk));
	jdff dff_B_czxlWPxq3_1(.din(w_dff_B_iluRJHjN2_1),.dout(w_dff_B_czxlWPxq3_1),.clk(gclk));
	jdff dff_B_sndVJQE01_1(.din(w_dff_B_czxlWPxq3_1),.dout(w_dff_B_sndVJQE01_1),.clk(gclk));
	jdff dff_B_1VemC9UF1_1(.din(w_dff_B_sndVJQE01_1),.dout(w_dff_B_1VemC9UF1_1),.clk(gclk));
	jdff dff_B_GsPBGEDN6_1(.din(w_dff_B_1VemC9UF1_1),.dout(w_dff_B_GsPBGEDN6_1),.clk(gclk));
	jdff dff_B_NUxOlpXU9_1(.din(w_dff_B_GsPBGEDN6_1),.dout(w_dff_B_NUxOlpXU9_1),.clk(gclk));
	jdff dff_B_rZ3P8Ezx8_1(.din(w_dff_B_NUxOlpXU9_1),.dout(w_dff_B_rZ3P8Ezx8_1),.clk(gclk));
	jdff dff_B_2hqh731n3_1(.din(w_dff_B_rZ3P8Ezx8_1),.dout(w_dff_B_2hqh731n3_1),.clk(gclk));
	jdff dff_B_B0nDGpt26_1(.din(w_dff_B_2hqh731n3_1),.dout(w_dff_B_B0nDGpt26_1),.clk(gclk));
	jdff dff_B_nPaF7WtD1_1(.din(w_dff_B_B0nDGpt26_1),.dout(w_dff_B_nPaF7WtD1_1),.clk(gclk));
	jdff dff_B_FGZyo1Ue0_1(.din(w_dff_B_nPaF7WtD1_1),.dout(w_dff_B_FGZyo1Ue0_1),.clk(gclk));
	jdff dff_B_IcnpIemx3_1(.din(w_dff_B_FGZyo1Ue0_1),.dout(w_dff_B_IcnpIemx3_1),.clk(gclk));
	jdff dff_B_HgvF8hE49_1(.din(n1689),.dout(w_dff_B_HgvF8hE49_1),.clk(gclk));
	jdff dff_A_GgUroV2W1_1(.dout(w_n854_1[1]),.din(w_dff_A_GgUroV2W1_1),.clk(gclk));
	jdff dff_A_jVSXcdB16_1(.dout(w_dff_A_GgUroV2W1_1),.din(w_dff_A_jVSXcdB16_1),.clk(gclk));
	jdff dff_A_CJWeJFSh3_1(.dout(w_dff_A_jVSXcdB16_1),.din(w_dff_A_CJWeJFSh3_1),.clk(gclk));
	jdff dff_A_Tirp1Pd82_1(.dout(w_dff_A_CJWeJFSh3_1),.din(w_dff_A_Tirp1Pd82_1),.clk(gclk));
	jdff dff_A_LG0FfJmp8_1(.dout(w_dff_A_Tirp1Pd82_1),.din(w_dff_A_LG0FfJmp8_1),.clk(gclk));
	jdff dff_A_Du1CZ2Xa5_1(.dout(w_dff_A_LG0FfJmp8_1),.din(w_dff_A_Du1CZ2Xa5_1),.clk(gclk));
	jdff dff_A_0iMtQxWI2_1(.dout(w_dff_A_Du1CZ2Xa5_1),.din(w_dff_A_0iMtQxWI2_1),.clk(gclk));
	jdff dff_A_OkZGQjhi2_1(.dout(w_dff_A_0iMtQxWI2_1),.din(w_dff_A_OkZGQjhi2_1),.clk(gclk));
	jdff dff_A_yzQhIqpR5_1(.dout(w_dff_A_OkZGQjhi2_1),.din(w_dff_A_yzQhIqpR5_1),.clk(gclk));
	jdff dff_A_s9dsHqFi9_1(.dout(w_dff_A_yzQhIqpR5_1),.din(w_dff_A_s9dsHqFi9_1),.clk(gclk));
	jdff dff_A_MWVJ7jpg3_1(.dout(w_dff_A_s9dsHqFi9_1),.din(w_dff_A_MWVJ7jpg3_1),.clk(gclk));
	jdff dff_A_UFcy6zM52_1(.dout(w_dff_A_MWVJ7jpg3_1),.din(w_dff_A_UFcy6zM52_1),.clk(gclk));
	jdff dff_A_eR5qvQQc5_1(.dout(w_dff_A_UFcy6zM52_1),.din(w_dff_A_eR5qvQQc5_1),.clk(gclk));
	jdff dff_A_E2vII9n89_1(.dout(w_dff_A_eR5qvQQc5_1),.din(w_dff_A_E2vII9n89_1),.clk(gclk));
	jdff dff_A_j6gsq6um5_2(.dout(w_n854_1[2]),.din(w_dff_A_j6gsq6um5_2),.clk(gclk));
	jdff dff_A_upXRwyB17_2(.dout(w_dff_A_j6gsq6um5_2),.din(w_dff_A_upXRwyB17_2),.clk(gclk));
	jdff dff_A_KBLre0CC9_2(.dout(w_dff_A_upXRwyB17_2),.din(w_dff_A_KBLre0CC9_2),.clk(gclk));
	jdff dff_A_Ee7j38Og1_2(.dout(w_dff_A_KBLre0CC9_2),.din(w_dff_A_Ee7j38Og1_2),.clk(gclk));
	jdff dff_A_eM0UDtrK2_2(.dout(w_dff_A_Ee7j38Og1_2),.din(w_dff_A_eM0UDtrK2_2),.clk(gclk));
	jdff dff_A_GErvG4gT4_2(.dout(w_dff_A_eM0UDtrK2_2),.din(w_dff_A_GErvG4gT4_2),.clk(gclk));
	jdff dff_A_e9wGZ5i35_2(.dout(w_dff_A_GErvG4gT4_2),.din(w_dff_A_e9wGZ5i35_2),.clk(gclk));
	jdff dff_A_irKNyDSR9_2(.dout(w_dff_A_e9wGZ5i35_2),.din(w_dff_A_irKNyDSR9_2),.clk(gclk));
	jdff dff_A_v4Ji4mre7_2(.dout(w_dff_A_irKNyDSR9_2),.din(w_dff_A_v4Ji4mre7_2),.clk(gclk));
	jdff dff_A_w3eUXdrG5_2(.dout(w_dff_A_v4Ji4mre7_2),.din(w_dff_A_w3eUXdrG5_2),.clk(gclk));
	jdff dff_B_nyYvB2tj6_1(.din(n1697),.dout(w_dff_B_nyYvB2tj6_1),.clk(gclk));
	jdff dff_B_xy3ImAAq3_1(.din(w_dff_B_nyYvB2tj6_1),.dout(w_dff_B_xy3ImAAq3_1),.clk(gclk));
	jdff dff_B_2oyRlj3a4_1(.din(w_dff_B_xy3ImAAq3_1),.dout(w_dff_B_2oyRlj3a4_1),.clk(gclk));
	jdff dff_B_iVNGJi6z1_1(.din(w_dff_B_2oyRlj3a4_1),.dout(w_dff_B_iVNGJi6z1_1),.clk(gclk));
	jdff dff_B_eC6dIvtR0_1(.din(w_dff_B_iVNGJi6z1_1),.dout(w_dff_B_eC6dIvtR0_1),.clk(gclk));
	jdff dff_B_BLm1o4kV1_1(.din(w_dff_B_eC6dIvtR0_1),.dout(w_dff_B_BLm1o4kV1_1),.clk(gclk));
	jdff dff_B_dJ4bMt2e9_1(.din(w_dff_B_BLm1o4kV1_1),.dout(w_dff_B_dJ4bMt2e9_1),.clk(gclk));
	jdff dff_B_eT8mCMpY8_1(.din(w_dff_B_dJ4bMt2e9_1),.dout(w_dff_B_eT8mCMpY8_1),.clk(gclk));
	jdff dff_B_4BHqEVxU3_1(.din(w_dff_B_eT8mCMpY8_1),.dout(w_dff_B_4BHqEVxU3_1),.clk(gclk));
	jdff dff_B_K8PIzCKL6_1(.din(w_dff_B_4BHqEVxU3_1),.dout(w_dff_B_K8PIzCKL6_1),.clk(gclk));
	jdff dff_B_wKEkvZPw4_1(.din(w_dff_B_K8PIzCKL6_1),.dout(w_dff_B_wKEkvZPw4_1),.clk(gclk));
	jdff dff_B_4zNlqT5V6_1(.din(w_dff_B_wKEkvZPw4_1),.dout(w_dff_B_4zNlqT5V6_1),.clk(gclk));
	jdff dff_B_AKd0NSDS6_1(.din(w_dff_B_4zNlqT5V6_1),.dout(w_dff_B_AKd0NSDS6_1),.clk(gclk));
	jdff dff_B_OXG23iN70_1(.din(w_dff_B_AKd0NSDS6_1),.dout(w_dff_B_OXG23iN70_1),.clk(gclk));
	jdff dff_B_XuTEtqXe2_1(.din(w_dff_B_OXG23iN70_1),.dout(w_dff_B_XuTEtqXe2_1),.clk(gclk));
	jdff dff_B_uy8rerwp8_1(.din(w_dff_B_XuTEtqXe2_1),.dout(w_dff_B_uy8rerwp8_1),.clk(gclk));
	jdff dff_B_Ulx3NKyY5_1(.din(w_dff_B_uy8rerwp8_1),.dout(w_dff_B_Ulx3NKyY5_1),.clk(gclk));
	jdff dff_B_8ZOx98qG7_1(.din(w_dff_B_Ulx3NKyY5_1),.dout(w_dff_B_8ZOx98qG7_1),.clk(gclk));
	jdff dff_B_IUuIk5yZ6_1(.din(w_dff_B_8ZOx98qG7_1),.dout(w_dff_B_IUuIk5yZ6_1),.clk(gclk));
	jdff dff_B_UyIHkBuD5_1(.din(w_dff_B_IUuIk5yZ6_1),.dout(w_dff_B_UyIHkBuD5_1),.clk(gclk));
	jdff dff_B_mnr5EtXf9_1(.din(w_dff_B_UyIHkBuD5_1),.dout(w_dff_B_mnr5EtXf9_1),.clk(gclk));
	jdff dff_B_Y2Qk5IFA0_1(.din(w_dff_B_mnr5EtXf9_1),.dout(w_dff_B_Y2Qk5IFA0_1),.clk(gclk));
	jdff dff_B_xFRH1E7d1_1(.din(w_dff_B_Y2Qk5IFA0_1),.dout(w_dff_B_xFRH1E7d1_1),.clk(gclk));
	jdff dff_B_UCyxkDuz9_1(.din(n1700),.dout(w_dff_B_UCyxkDuz9_1),.clk(gclk));
	jdff dff_B_IEpbaqTd3_1(.din(w_dff_B_UCyxkDuz9_1),.dout(w_dff_B_IEpbaqTd3_1),.clk(gclk));
	jdff dff_B_aUeayiQz7_1(.din(w_dff_B_IEpbaqTd3_1),.dout(w_dff_B_aUeayiQz7_1),.clk(gclk));
	jdff dff_B_sxQEjlpR4_1(.din(w_dff_B_aUeayiQz7_1),.dout(w_dff_B_sxQEjlpR4_1),.clk(gclk));
	jdff dff_B_SuZgzeC56_1(.din(w_dff_B_sxQEjlpR4_1),.dout(w_dff_B_SuZgzeC56_1),.clk(gclk));
	jdff dff_B_FmqYyeU43_1(.din(w_dff_B_SuZgzeC56_1),.dout(w_dff_B_FmqYyeU43_1),.clk(gclk));
	jdff dff_B_HaorQlKU5_1(.din(w_dff_B_FmqYyeU43_1),.dout(w_dff_B_HaorQlKU5_1),.clk(gclk));
	jdff dff_B_woz3DQCA1_1(.din(w_dff_B_HaorQlKU5_1),.dout(w_dff_B_woz3DQCA1_1),.clk(gclk));
	jdff dff_B_d5Gs0Tdi7_1(.din(w_dff_B_woz3DQCA1_1),.dout(w_dff_B_d5Gs0Tdi7_1),.clk(gclk));
	jdff dff_B_wFSc6V042_1(.din(w_dff_B_d5Gs0Tdi7_1),.dout(w_dff_B_wFSc6V042_1),.clk(gclk));
	jdff dff_B_GE4vzV4B0_1(.din(w_dff_B_wFSc6V042_1),.dout(w_dff_B_GE4vzV4B0_1),.clk(gclk));
	jdff dff_B_Ik53PXFx7_1(.din(w_dff_B_GE4vzV4B0_1),.dout(w_dff_B_Ik53PXFx7_1),.clk(gclk));
	jdff dff_B_plbUrMv81_1(.din(w_dff_B_Ik53PXFx7_1),.dout(w_dff_B_plbUrMv81_1),.clk(gclk));
	jdff dff_B_RmVWAyyF7_1(.din(w_dff_B_plbUrMv81_1),.dout(w_dff_B_RmVWAyyF7_1),.clk(gclk));
	jdff dff_B_yw8HwcB69_1(.din(w_dff_B_RmVWAyyF7_1),.dout(w_dff_B_yw8HwcB69_1),.clk(gclk));
	jdff dff_B_WxCQHscR9_1(.din(w_dff_B_yw8HwcB69_1),.dout(w_dff_B_WxCQHscR9_1),.clk(gclk));
	jdff dff_B_hEb9Ov7e2_1(.din(w_dff_B_WxCQHscR9_1),.dout(w_dff_B_hEb9Ov7e2_1),.clk(gclk));
	jdff dff_B_aiHHvdUR5_1(.din(w_dff_B_hEb9Ov7e2_1),.dout(w_dff_B_aiHHvdUR5_1),.clk(gclk));
	jdff dff_B_w0UPXMMj5_1(.din(w_dff_B_aiHHvdUR5_1),.dout(w_dff_B_w0UPXMMj5_1),.clk(gclk));
	jdff dff_B_BB80w2h76_1(.din(w_dff_B_w0UPXMMj5_1),.dout(w_dff_B_BB80w2h76_1),.clk(gclk));
	jdff dff_B_S1TlZL3Q5_1(.din(w_dff_B_BB80w2h76_1),.dout(w_dff_B_S1TlZL3Q5_1),.clk(gclk));
	jdff dff_B_OyrKFmYT7_1(.din(n1701),.dout(w_dff_B_OyrKFmYT7_1),.clk(gclk));
	jdff dff_B_SHDFiHai4_1(.din(n1709),.dout(w_dff_B_SHDFiHai4_1),.clk(gclk));
	jdff dff_B_r4nl3ba44_1(.din(w_dff_B_SHDFiHai4_1),.dout(w_dff_B_r4nl3ba44_1),.clk(gclk));
	jdff dff_B_1R4LT2rQ8_1(.din(w_dff_B_r4nl3ba44_1),.dout(w_dff_B_1R4LT2rQ8_1),.clk(gclk));
	jdff dff_B_y6LL5sP02_1(.din(w_dff_B_1R4LT2rQ8_1),.dout(w_dff_B_y6LL5sP02_1),.clk(gclk));
	jdff dff_B_d7VdmAkg5_1(.din(w_dff_B_y6LL5sP02_1),.dout(w_dff_B_d7VdmAkg5_1),.clk(gclk));
	jdff dff_B_CKTWOprv3_1(.din(w_dff_B_d7VdmAkg5_1),.dout(w_dff_B_CKTWOprv3_1),.clk(gclk));
	jdff dff_B_HmYxEVDQ9_1(.din(w_dff_B_CKTWOprv3_1),.dout(w_dff_B_HmYxEVDQ9_1),.clk(gclk));
	jdff dff_B_PrCjGr6S1_1(.din(w_dff_B_HmYxEVDQ9_1),.dout(w_dff_B_PrCjGr6S1_1),.clk(gclk));
	jdff dff_B_6hw44P118_1(.din(w_dff_B_PrCjGr6S1_1),.dout(w_dff_B_6hw44P118_1),.clk(gclk));
	jdff dff_B_qOaxueCp3_1(.din(w_dff_B_6hw44P118_1),.dout(w_dff_B_qOaxueCp3_1),.clk(gclk));
	jdff dff_B_wYx89UmX7_1(.din(w_dff_B_qOaxueCp3_1),.dout(w_dff_B_wYx89UmX7_1),.clk(gclk));
	jdff dff_B_3ghB2Ggm3_1(.din(w_dff_B_wYx89UmX7_1),.dout(w_dff_B_3ghB2Ggm3_1),.clk(gclk));
	jdff dff_B_5yEehwxw9_1(.din(w_dff_B_3ghB2Ggm3_1),.dout(w_dff_B_5yEehwxw9_1),.clk(gclk));
	jdff dff_B_enloygGK2_1(.din(w_dff_B_5yEehwxw9_1),.dout(w_dff_B_enloygGK2_1),.clk(gclk));
	jdff dff_B_7RHKiZSp3_1(.din(w_dff_B_enloygGK2_1),.dout(w_dff_B_7RHKiZSp3_1),.clk(gclk));
	jdff dff_B_mkvQskNg2_1(.din(w_dff_B_7RHKiZSp3_1),.dout(w_dff_B_mkvQskNg2_1),.clk(gclk));
	jdff dff_B_wQ5qyDNm1_1(.din(w_dff_B_mkvQskNg2_1),.dout(w_dff_B_wQ5qyDNm1_1),.clk(gclk));
	jdff dff_B_2dFyI4c60_1(.din(w_dff_B_wQ5qyDNm1_1),.dout(w_dff_B_2dFyI4c60_1),.clk(gclk));
	jdff dff_B_D6l5Yjcy1_1(.din(w_dff_B_2dFyI4c60_1),.dout(w_dff_B_D6l5Yjcy1_1),.clk(gclk));
	jdff dff_B_cjjzdCiv1_1(.din(w_dff_B_D6l5Yjcy1_1),.dout(w_dff_B_cjjzdCiv1_1),.clk(gclk));
	jdff dff_B_YWc2PxDc3_1(.din(w_dff_B_cjjzdCiv1_1),.dout(w_dff_B_YWc2PxDc3_1),.clk(gclk));
	jdff dff_B_aqcr2WXc9_1(.din(w_dff_B_YWc2PxDc3_1),.dout(w_dff_B_aqcr2WXc9_1),.clk(gclk));
	jdff dff_B_5wark3kh5_1(.din(w_dff_B_aqcr2WXc9_1),.dout(w_dff_B_5wark3kh5_1),.clk(gclk));
	jdff dff_B_FG9q5yje3_1(.din(n1711),.dout(w_dff_B_FG9q5yje3_1),.clk(gclk));
	jdff dff_B_RzXeeNyg4_1(.din(w_dff_B_FG9q5yje3_1),.dout(w_dff_B_RzXeeNyg4_1),.clk(gclk));
	jdff dff_B_HVfQU3664_1(.din(w_dff_B_RzXeeNyg4_1),.dout(w_dff_B_HVfQU3664_1),.clk(gclk));
	jdff dff_B_gfY1tcdS5_1(.din(w_dff_B_HVfQU3664_1),.dout(w_dff_B_gfY1tcdS5_1),.clk(gclk));
	jdff dff_B_Yv3NyAhq8_1(.din(w_dff_B_gfY1tcdS5_1),.dout(w_dff_B_Yv3NyAhq8_1),.clk(gclk));
	jdff dff_B_JN1TonOg3_1(.din(w_dff_B_Yv3NyAhq8_1),.dout(w_dff_B_JN1TonOg3_1),.clk(gclk));
	jdff dff_B_7z5hVVUh6_1(.din(w_dff_B_JN1TonOg3_1),.dout(w_dff_B_7z5hVVUh6_1),.clk(gclk));
	jdff dff_B_R0q1cWjx6_1(.din(w_dff_B_7z5hVVUh6_1),.dout(w_dff_B_R0q1cWjx6_1),.clk(gclk));
	jdff dff_B_F0Pbj0uN5_1(.din(w_dff_B_R0q1cWjx6_1),.dout(w_dff_B_F0Pbj0uN5_1),.clk(gclk));
	jdff dff_B_IZTA4Esk5_1(.din(w_dff_B_F0Pbj0uN5_1),.dout(w_dff_B_IZTA4Esk5_1),.clk(gclk));
	jdff dff_B_lKE4yU3v2_1(.din(w_dff_B_IZTA4Esk5_1),.dout(w_dff_B_lKE4yU3v2_1),.clk(gclk));
	jdff dff_B_VTghs1Pl6_1(.din(w_dff_B_lKE4yU3v2_1),.dout(w_dff_B_VTghs1Pl6_1),.clk(gclk));
	jdff dff_B_Gb7dGKxX2_1(.din(w_dff_B_VTghs1Pl6_1),.dout(w_dff_B_Gb7dGKxX2_1),.clk(gclk));
	jdff dff_B_lBuFHirz3_1(.din(w_dff_B_Gb7dGKxX2_1),.dout(w_dff_B_lBuFHirz3_1),.clk(gclk));
	jdff dff_B_wjcyD9Pv7_1(.din(w_dff_B_lBuFHirz3_1),.dout(w_dff_B_wjcyD9Pv7_1),.clk(gclk));
	jdff dff_B_4aH8sZ125_1(.din(w_dff_B_wjcyD9Pv7_1),.dout(w_dff_B_4aH8sZ125_1),.clk(gclk));
	jdff dff_B_Q1RHRg5T0_1(.din(w_dff_B_4aH8sZ125_1),.dout(w_dff_B_Q1RHRg5T0_1),.clk(gclk));
	jdff dff_B_qjpJX1UX7_1(.din(w_dff_B_Q1RHRg5T0_1),.dout(w_dff_B_qjpJX1UX7_1),.clk(gclk));
	jdff dff_B_ugSKk3lK5_1(.din(w_dff_B_qjpJX1UX7_1),.dout(w_dff_B_ugSKk3lK5_1),.clk(gclk));
	jdff dff_B_mVGjxRFb1_1(.din(w_dff_B_ugSKk3lK5_1),.dout(w_dff_B_mVGjxRFb1_1),.clk(gclk));
	jdff dff_B_UhhF2aeY9_1(.din(w_dff_B_mVGjxRFb1_1),.dout(w_dff_B_UhhF2aeY9_1),.clk(gclk));
	jdff dff_B_qck1SFfG3_1(.din(n1712),.dout(w_dff_B_qck1SFfG3_1),.clk(gclk));
	jdff dff_B_Ywku2r8g2_0(.din(n1678),.dout(w_dff_B_Ywku2r8g2_0),.clk(gclk));
	jdff dff_B_fRU7VHFG1_0(.din(w_dff_B_Ywku2r8g2_0),.dout(w_dff_B_fRU7VHFG1_0),.clk(gclk));
	jdff dff_B_rQdDj2eA7_0(.din(w_dff_B_fRU7VHFG1_0),.dout(w_dff_B_rQdDj2eA7_0),.clk(gclk));
	jdff dff_B_CdO5itrP2_0(.din(w_dff_B_rQdDj2eA7_0),.dout(w_dff_B_CdO5itrP2_0),.clk(gclk));
	jdff dff_B_3DfPf54M9_0(.din(w_dff_B_CdO5itrP2_0),.dout(w_dff_B_3DfPf54M9_0),.clk(gclk));
	jdff dff_B_mq5e2Zzx6_0(.din(w_dff_B_3DfPf54M9_0),.dout(w_dff_B_mq5e2Zzx6_0),.clk(gclk));
	jdff dff_B_9Sia1E4D3_0(.din(w_dff_B_mq5e2Zzx6_0),.dout(w_dff_B_9Sia1E4D3_0),.clk(gclk));
	jdff dff_B_QDndUrLm7_0(.din(w_dff_B_9Sia1E4D3_0),.dout(w_dff_B_QDndUrLm7_0),.clk(gclk));
	jdff dff_B_ABFe8TIy3_0(.din(w_dff_B_QDndUrLm7_0),.dout(w_dff_B_ABFe8TIy3_0),.clk(gclk));
	jdff dff_B_jzHHyC1G5_0(.din(w_dff_B_ABFe8TIy3_0),.dout(w_dff_B_jzHHyC1G5_0),.clk(gclk));
	jdff dff_B_nZuCHGPA4_0(.din(w_dff_B_jzHHyC1G5_0),.dout(w_dff_B_nZuCHGPA4_0),.clk(gclk));
	jdff dff_B_uxJvCPl38_0(.din(w_dff_B_nZuCHGPA4_0),.dout(w_dff_B_uxJvCPl38_0),.clk(gclk));
	jdff dff_B_Z8XCAVaB1_0(.din(w_dff_B_uxJvCPl38_0),.dout(w_dff_B_Z8XCAVaB1_0),.clk(gclk));
	jdff dff_B_ouBIezaM0_0(.din(w_dff_B_Z8XCAVaB1_0),.dout(w_dff_B_ouBIezaM0_0),.clk(gclk));
	jdff dff_B_7Mx015AW6_0(.din(w_dff_B_ouBIezaM0_0),.dout(w_dff_B_7Mx015AW6_0),.clk(gclk));
	jdff dff_B_SItuqPlM5_0(.din(w_dff_B_7Mx015AW6_0),.dout(w_dff_B_SItuqPlM5_0),.clk(gclk));
	jdff dff_B_ZVYJLPdy5_0(.din(w_dff_B_SItuqPlM5_0),.dout(w_dff_B_ZVYJLPdy5_0),.clk(gclk));
	jdff dff_B_zNNL6OLI0_0(.din(w_dff_B_ZVYJLPdy5_0),.dout(w_dff_B_zNNL6OLI0_0),.clk(gclk));
	jdff dff_B_11Y5fuYu3_0(.din(w_dff_B_zNNL6OLI0_0),.dout(w_dff_B_11Y5fuYu3_0),.clk(gclk));
	jdff dff_B_wZ4qtbJV6_0(.din(n1501),.dout(w_dff_B_wZ4qtbJV6_0),.clk(gclk));
	jdff dff_B_B6ZabqjA5_0(.din(w_dff_B_wZ4qtbJV6_0),.dout(w_dff_B_B6ZabqjA5_0),.clk(gclk));
	jdff dff_B_iYc4xeuz8_0(.din(w_dff_B_B6ZabqjA5_0),.dout(w_dff_B_iYc4xeuz8_0),.clk(gclk));
	jdff dff_B_YUSImXH81_0(.din(w_dff_B_iYc4xeuz8_0),.dout(w_dff_B_YUSImXH81_0),.clk(gclk));
	jdff dff_B_fuor0P728_0(.din(w_dff_B_YUSImXH81_0),.dout(w_dff_B_fuor0P728_0),.clk(gclk));
	jdff dff_B_vnyppdtj0_0(.din(w_dff_B_fuor0P728_0),.dout(w_dff_B_vnyppdtj0_0),.clk(gclk));
	jdff dff_B_hDjk5vER8_0(.din(w_dff_B_vnyppdtj0_0),.dout(w_dff_B_hDjk5vER8_0),.clk(gclk));
	jdff dff_B_rBb9Fa5m0_0(.din(w_dff_B_hDjk5vER8_0),.dout(w_dff_B_rBb9Fa5m0_0),.clk(gclk));
	jdff dff_B_z22eYMUi6_0(.din(w_dff_B_rBb9Fa5m0_0),.dout(w_dff_B_z22eYMUi6_0),.clk(gclk));
	jdff dff_B_0i2kTdtc2_1(.din(n1453),.dout(w_dff_B_0i2kTdtc2_1),.clk(gclk));
	jdff dff_B_NO5SrzkV7_0(.din(n1452),.dout(w_dff_B_NO5SrzkV7_0),.clk(gclk));
	jdff dff_A_UpHFzeke5_0(.dout(w_n1451_0[0]),.din(w_dff_A_UpHFzeke5_0),.clk(gclk));
	jdff dff_A_7wxXQokn0_0(.dout(w_dff_A_UpHFzeke5_0),.din(w_dff_A_7wxXQokn0_0),.clk(gclk));
	jdff dff_B_b8J3pfmx8_0(.din(n1450),.dout(w_dff_B_b8J3pfmx8_0),.clk(gclk));
	jdff dff_B_SFlZDlf13_0(.din(w_dff_B_b8J3pfmx8_0),.dout(w_dff_B_SFlZDlf13_0),.clk(gclk));
	jdff dff_B_8TqIhvGq3_0(.din(w_dff_B_SFlZDlf13_0),.dout(w_dff_B_8TqIhvGq3_0),.clk(gclk));
	jdff dff_B_J1AkRO136_1(.din(n1448),.dout(w_dff_B_J1AkRO136_1),.clk(gclk));
	jdff dff_B_ib2IL73b4_1(.din(w_dff_B_J1AkRO136_1),.dout(w_dff_B_ib2IL73b4_1),.clk(gclk));
	jdff dff_B_p1RAyhWe0_1(.din(w_dff_B_ib2IL73b4_1),.dout(w_dff_B_p1RAyhWe0_1),.clk(gclk));
	jdff dff_B_ZqKnkvmN1_1(.din(n1439),.dout(w_dff_B_ZqKnkvmN1_1),.clk(gclk));
	jdff dff_B_ojDaT3h42_1(.din(n1441),.dout(w_dff_B_ojDaT3h42_1),.clk(gclk));
	jdff dff_B_W3Dv9XHm7_0(.din(n1437),.dout(w_dff_B_W3Dv9XHm7_0),.clk(gclk));
	jdff dff_B_lb2sWyLx1_0(.din(n1436),.dout(w_dff_B_lb2sWyLx1_0),.clk(gclk));
	jdff dff_A_cssLASeX9_0(.dout(w_n1429_0[0]),.din(w_dff_A_cssLASeX9_0),.clk(gclk));
	jdff dff_B_GELGpxoG6_1(.din(n1427),.dout(w_dff_B_GELGpxoG6_1),.clk(gclk));
	jdff dff_A_yiq9g2aP7_2(.dout(w_n641_0[2]),.din(w_dff_A_yiq9g2aP7_2),.clk(gclk));
	jdff dff_A_AB6PTBb39_2(.dout(w_dff_A_yiq9g2aP7_2),.din(w_dff_A_AB6PTBb39_2),.clk(gclk));
	jdff dff_A_QIqXiJiq1_0(.dout(w_n640_0[0]),.din(w_dff_A_QIqXiJiq1_0),.clk(gclk));
	jdff dff_A_lgyLa82g0_0(.dout(w_n639_0[0]),.din(w_dff_A_lgyLa82g0_0),.clk(gclk));
	jdff dff_A_e0HmERPy0_0(.dout(w_n624_0[0]),.din(w_dff_A_e0HmERPy0_0),.clk(gclk));
	jdff dff_A_OHwws77V4_0(.dout(w_dff_A_e0HmERPy0_0),.din(w_dff_A_OHwws77V4_0),.clk(gclk));
	jdff dff_A_f4Qd0c5u7_1(.dout(w_n624_0[1]),.din(w_dff_A_f4Qd0c5u7_1),.clk(gclk));
	jdff dff_B_K8LUhpwg3_3(.din(n624),.dout(w_dff_B_K8LUhpwg3_3),.clk(gclk));
	jdff dff_B_Pns1XHaU6_3(.din(w_dff_B_K8LUhpwg3_3),.dout(w_dff_B_Pns1XHaU6_3),.clk(gclk));
	jdff dff_A_77FCiIJy7_0(.dout(w_n1425_0[0]),.din(w_dff_A_77FCiIJy7_0),.clk(gclk));
	jdff dff_B_y7USFW1T9_1(.din(n1411),.dout(w_dff_B_y7USFW1T9_1),.clk(gclk));
	jdff dff_A_XjBaWqj13_0(.dout(w_n1422_0[0]),.din(w_dff_A_XjBaWqj13_0),.clk(gclk));
	jdff dff_B_u8AEOMbS8_1(.din(n1418),.dout(w_dff_B_u8AEOMbS8_1),.clk(gclk));
	jdff dff_B_v6bKkAAY4_1(.din(w_dff_B_u8AEOMbS8_1),.dout(w_dff_B_v6bKkAAY4_1),.clk(gclk));
	jdff dff_B_nfYiIvAu1_1(.din(w_dff_B_v6bKkAAY4_1),.dout(w_dff_B_nfYiIvAu1_1),.clk(gclk));
	jdff dff_A_drZdhkdz7_2(.dout(w_n792_0[2]),.din(w_dff_A_drZdhkdz7_2),.clk(gclk));
	jdff dff_A_7DptGaxU0_2(.dout(w_dff_A_drZdhkdz7_2),.din(w_dff_A_7DptGaxU0_2),.clk(gclk));
	jdff dff_A_Rd9Qk2go1_2(.dout(w_dff_A_7DptGaxU0_2),.din(w_dff_A_Rd9Qk2go1_2),.clk(gclk));
	jdff dff_A_8Hfju6PD7_2(.dout(w_dff_A_Rd9Qk2go1_2),.din(w_dff_A_8Hfju6PD7_2),.clk(gclk));
	jdff dff_A_tG9trZYe2_2(.dout(w_dff_A_8Hfju6PD7_2),.din(w_dff_A_tG9trZYe2_2),.clk(gclk));
	jdff dff_A_0RBPngsx4_2(.dout(w_dff_A_tG9trZYe2_2),.din(w_dff_A_0RBPngsx4_2),.clk(gclk));
	jdff dff_A_tv11bPYw0_2(.dout(w_dff_A_0RBPngsx4_2),.din(w_dff_A_tv11bPYw0_2),.clk(gclk));
	jdff dff_A_dUIBOcCW1_2(.dout(w_dff_A_tv11bPYw0_2),.din(w_dff_A_dUIBOcCW1_2),.clk(gclk));
	jdff dff_A_zmpyFrKI5_2(.dout(w_dff_A_dUIBOcCW1_2),.din(w_dff_A_zmpyFrKI5_2),.clk(gclk));
	jdff dff_A_Ae76oq8l4_1(.dout(w_n790_0[1]),.din(w_dff_A_Ae76oq8l4_1),.clk(gclk));
	jdff dff_A_RA4bUFWW9_1(.dout(w_dff_A_Ae76oq8l4_1),.din(w_dff_A_RA4bUFWW9_1),.clk(gclk));
	jdff dff_A_4yHa4Zxk5_1(.dout(w_dff_A_RA4bUFWW9_1),.din(w_dff_A_4yHa4Zxk5_1),.clk(gclk));
	jdff dff_A_CJXrbhge1_1(.dout(w_dff_A_4yHa4Zxk5_1),.din(w_dff_A_CJXrbhge1_1),.clk(gclk));
	jdff dff_A_xmPDzEJ46_1(.dout(w_dff_A_CJXrbhge1_1),.din(w_dff_A_xmPDzEJ46_1),.clk(gclk));
	jdff dff_A_y6WFFCKg1_1(.dout(w_dff_A_xmPDzEJ46_1),.din(w_dff_A_y6WFFCKg1_1),.clk(gclk));
	jdff dff_A_Dwcuz1Mt6_1(.dout(w_dff_A_y6WFFCKg1_1),.din(w_dff_A_Dwcuz1Mt6_1),.clk(gclk));
	jdff dff_A_fkiZc9bO0_1(.dout(w_dff_A_Dwcuz1Mt6_1),.din(w_dff_A_fkiZc9bO0_1),.clk(gclk));
	jdff dff_A_9NadUDZn9_1(.dout(w_dff_A_fkiZc9bO0_1),.din(w_dff_A_9NadUDZn9_1),.clk(gclk));
	jdff dff_A_YMMn1aJu8_1(.dout(w_dff_A_9NadUDZn9_1),.din(w_dff_A_YMMn1aJu8_1),.clk(gclk));
	jdff dff_B_ZiixEKxx1_1(.din(n1413),.dout(w_dff_B_ZiixEKxx1_1),.clk(gclk));
	jdff dff_B_ZsMevCQX5_1(.din(w_dff_B_ZiixEKxx1_1),.dout(w_dff_B_ZsMevCQX5_1),.clk(gclk));
	jdff dff_B_JKDdWWuv9_1(.din(w_dff_B_ZsMevCQX5_1),.dout(w_dff_B_JKDdWWuv9_1),.clk(gclk));
	jdff dff_B_kwom3u9N4_1(.din(w_dff_B_JKDdWWuv9_1),.dout(w_dff_B_kwom3u9N4_1),.clk(gclk));
	jdff dff_B_GKmUyL8K8_1(.din(n1414),.dout(w_dff_B_GKmUyL8K8_1),.clk(gclk));
	jdff dff_B_bDlfFRgC2_1(.din(w_dff_B_GKmUyL8K8_1),.dout(w_dff_B_bDlfFRgC2_1),.clk(gclk));
	jdff dff_B_2FUUdo6f3_1(.din(w_dff_B_bDlfFRgC2_1),.dout(w_dff_B_2FUUdo6f3_1),.clk(gclk));
	jdff dff_A_NA9Df6H68_1(.dout(w_n821_0[1]),.din(w_dff_A_NA9Df6H68_1),.clk(gclk));
	jdff dff_B_9zmzvveo6_1(.din(n812),.dout(w_dff_B_9zmzvveo6_1),.clk(gclk));
	jdff dff_B_N2ElJB7k8_1(.din(w_dff_B_9zmzvveo6_1),.dout(w_dff_B_N2ElJB7k8_1),.clk(gclk));
	jdff dff_B_vucXC8zj6_1(.din(w_dff_B_N2ElJB7k8_1),.dout(w_dff_B_vucXC8zj6_1),.clk(gclk));
	jdff dff_B_okWyP26V2_1(.din(w_dff_B_vucXC8zj6_1),.dout(w_dff_B_okWyP26V2_1),.clk(gclk));
	jdff dff_B_IN16bStA5_1(.din(n813),.dout(w_dff_B_IN16bStA5_1),.clk(gclk));
	jdff dff_B_chb4fUGz8_1(.din(w_dff_B_IN16bStA5_1),.dout(w_dff_B_chb4fUGz8_1),.clk(gclk));
	jdff dff_B_wsuO4F6W8_1(.din(w_dff_B_chb4fUGz8_1),.dout(w_dff_B_wsuO4F6W8_1),.clk(gclk));
	jdff dff_A_CvaPLRfG1_1(.dout(w_n819_0[1]),.din(w_dff_A_CvaPLRfG1_1),.clk(gclk));
	jdff dff_A_eUZQ0gCo5_1(.dout(w_dff_A_CvaPLRfG1_1),.din(w_dff_A_eUZQ0gCo5_1),.clk(gclk));
	jdff dff_A_hxGff9QT8_0(.dout(w_n814_0[0]),.din(w_dff_A_hxGff9QT8_0),.clk(gclk));
	jdff dff_A_l2d0QREj0_0(.dout(w_dff_A_hxGff9QT8_0),.din(w_dff_A_l2d0QREj0_0),.clk(gclk));
	jdff dff_A_AL4TBzB66_0(.dout(w_dff_A_l2d0QREj0_0),.din(w_dff_A_AL4TBzB66_0),.clk(gclk));
	jdff dff_A_oND0CmAJ6_1(.dout(w_n814_0[1]),.din(w_dff_A_oND0CmAJ6_1),.clk(gclk));
	jdff dff_A_EEJ6wBEC7_1(.dout(w_dff_A_oND0CmAJ6_1),.din(w_dff_A_EEJ6wBEC7_1),.clk(gclk));
	jdff dff_A_TaBuKhQ45_1(.dout(w_n1412_0[1]),.din(w_dff_A_TaBuKhQ45_1),.clk(gclk));
	jdff dff_A_Zmmqp0qp7_1(.dout(w_dff_A_TaBuKhQ45_1),.din(w_dff_A_Zmmqp0qp7_1),.clk(gclk));
	jdff dff_A_0XMBlSB18_2(.dout(w_n1412_0[2]),.din(w_dff_A_0XMBlSB18_2),.clk(gclk));
	jdff dff_B_piuNxwIg6_3(.din(n1412),.dout(w_dff_B_piuNxwIg6_3),.clk(gclk));
	jdff dff_B_brFdKLeN3_3(.din(w_dff_B_piuNxwIg6_3),.dout(w_dff_B_brFdKLeN3_3),.clk(gclk));
	jdff dff_B_lwwr2A2p8_3(.din(w_dff_B_brFdKLeN3_3),.dout(w_dff_B_lwwr2A2p8_3),.clk(gclk));
	jdff dff_B_sUQf3Mlt0_3(.din(w_dff_B_lwwr2A2p8_3),.dout(w_dff_B_sUQf3Mlt0_3),.clk(gclk));
	jdff dff_B_aSEUAJJ42_3(.din(w_dff_B_sUQf3Mlt0_3),.dout(w_dff_B_aSEUAJJ42_3),.clk(gclk));
	jdff dff_B_cDJVJztp5_3(.din(w_dff_B_aSEUAJJ42_3),.dout(w_dff_B_cDJVJztp5_3),.clk(gclk));
	jdff dff_B_EVhQzDYu4_3(.din(w_dff_B_cDJVJztp5_3),.dout(w_dff_B_EVhQzDYu4_3),.clk(gclk));
	jdff dff_B_faHhOZgZ0_3(.din(w_dff_B_EVhQzDYu4_3),.dout(w_dff_B_faHhOZgZ0_3),.clk(gclk));
	jdff dff_B_kD7cOaV19_3(.din(w_dff_B_faHhOZgZ0_3),.dout(w_dff_B_kD7cOaV19_3),.clk(gclk));
	jdff dff_B_9csyNqWX5_3(.din(w_dff_B_kD7cOaV19_3),.dout(w_dff_B_9csyNqWX5_3),.clk(gclk));
	jdff dff_A_TL0ht9Jp2_0(.dout(w_n1410_0[0]),.din(w_dff_A_TL0ht9Jp2_0),.clk(gclk));
	jdff dff_B_A7oqnMQB8_0(.din(n1409),.dout(w_dff_B_A7oqnMQB8_0),.clk(gclk));
	jdff dff_B_HiDGTUnB7_0(.din(w_dff_B_A7oqnMQB8_0),.dout(w_dff_B_HiDGTUnB7_0),.clk(gclk));
	jdff dff_A_b30ZD7DE2_0(.dout(w_n644_0[0]),.din(w_dff_A_b30ZD7DE2_0),.clk(gclk));
	jdff dff_A_QuYbWtTq1_0(.dout(w_dff_A_b30ZD7DE2_0),.din(w_dff_A_QuYbWtTq1_0),.clk(gclk));
	jdff dff_A_jTuHUfu36_0(.dout(w_dff_A_QuYbWtTq1_0),.din(w_dff_A_jTuHUfu36_0),.clk(gclk));
	jdff dff_A_PyNPhz278_0(.dout(w_dff_A_jTuHUfu36_0),.din(w_dff_A_PyNPhz278_0),.clk(gclk));
	jdff dff_A_LuUV5yCQ1_2(.dout(w_n644_0[2]),.din(w_dff_A_LuUV5yCQ1_2),.clk(gclk));
	jdff dff_A_uLWTeDtJ1_2(.dout(w_dff_A_LuUV5yCQ1_2),.din(w_dff_A_uLWTeDtJ1_2),.clk(gclk));
	jdff dff_B_oSMEsVHY2_1(.din(n727),.dout(w_dff_B_oSMEsVHY2_1),.clk(gclk));
	jdff dff_A_PzJQwF4I3_0(.dout(w_n726_0[0]),.din(w_dff_A_PzJQwF4I3_0),.clk(gclk));
	jdff dff_A_uvSGRqJ13_0(.dout(w_dff_A_PzJQwF4I3_0),.din(w_dff_A_uvSGRqJ13_0),.clk(gclk));
	jdff dff_B_HPmUIL054_2(.din(n1694),.dout(w_dff_B_HPmUIL054_2),.clk(gclk));
	jdff dff_B_9fwOs6c77_2(.din(w_dff_B_HPmUIL054_2),.dout(w_dff_B_9fwOs6c77_2),.clk(gclk));
	jdff dff_B_Thd5Vae35_2(.din(w_dff_B_9fwOs6c77_2),.dout(w_dff_B_Thd5Vae35_2),.clk(gclk));
	jdff dff_B_eDjis2yY9_2(.din(w_dff_B_Thd5Vae35_2),.dout(w_dff_B_eDjis2yY9_2),.clk(gclk));
	jdff dff_B_Qw7943Sf2_2(.din(w_dff_B_eDjis2yY9_2),.dout(w_dff_B_Qw7943Sf2_2),.clk(gclk));
	jdff dff_B_SSx1WpRp3_2(.din(w_dff_B_Qw7943Sf2_2),.dout(w_dff_B_SSx1WpRp3_2),.clk(gclk));
	jdff dff_B_Ao5tScGk0_2(.din(w_dff_B_SSx1WpRp3_2),.dout(w_dff_B_Ao5tScGk0_2),.clk(gclk));
	jdff dff_B_pJL1NtXi5_2(.din(w_dff_B_Ao5tScGk0_2),.dout(w_dff_B_pJL1NtXi5_2),.clk(gclk));
	jdff dff_B_8R5WqX8z9_2(.din(w_dff_B_pJL1NtXi5_2),.dout(w_dff_B_8R5WqX8z9_2),.clk(gclk));
	jdff dff_B_fB6juIMr0_2(.din(w_dff_B_8R5WqX8z9_2),.dout(w_dff_B_fB6juIMr0_2),.clk(gclk));
	jdff dff_B_aFYCOJbS2_2(.din(w_dff_B_fB6juIMr0_2),.dout(w_dff_B_aFYCOJbS2_2),.clk(gclk));
	jdff dff_B_XDInrnuN8_2(.din(w_dff_B_aFYCOJbS2_2),.dout(w_dff_B_XDInrnuN8_2),.clk(gclk));
	jdff dff_B_HaRs99yT4_2(.din(w_dff_B_XDInrnuN8_2),.dout(w_dff_B_HaRs99yT4_2),.clk(gclk));
	jdff dff_B_VnWqcvaT1_2(.din(w_dff_B_HaRs99yT4_2),.dout(w_dff_B_VnWqcvaT1_2),.clk(gclk));
	jdff dff_B_vFv4DzFa8_2(.din(w_dff_B_VnWqcvaT1_2),.dout(w_dff_B_vFv4DzFa8_2),.clk(gclk));
	jdff dff_B_KnMLcJqJ3_2(.din(w_dff_B_vFv4DzFa8_2),.dout(w_dff_B_KnMLcJqJ3_2),.clk(gclk));
	jdff dff_B_etcTJXVC3_2(.din(w_dff_B_KnMLcJqJ3_2),.dout(w_dff_B_etcTJXVC3_2),.clk(gclk));
	jdff dff_B_enkNTEp98_2(.din(w_dff_B_etcTJXVC3_2),.dout(w_dff_B_enkNTEp98_2),.clk(gclk));
	jdff dff_B_gHLFmskD2_2(.din(w_dff_B_enkNTEp98_2),.dout(w_dff_B_gHLFmskD2_2),.clk(gclk));
	jdff dff_B_TovuJMhW8_2(.din(w_dff_B_gHLFmskD2_2),.dout(w_dff_B_TovuJMhW8_2),.clk(gclk));
	jdff dff_B_fa94FOAF1_2(.din(w_dff_B_TovuJMhW8_2),.dout(w_dff_B_fa94FOAF1_2),.clk(gclk));
	jdff dff_B_ZTGF89tH2_2(.din(w_dff_B_fa94FOAF1_2),.dout(w_dff_B_ZTGF89tH2_2),.clk(gclk));
	jdff dff_B_L8UPxx8e1_2(.din(w_dff_B_ZTGF89tH2_2),.dout(w_dff_B_L8UPxx8e1_2),.clk(gclk));
	jdff dff_B_PPiahgxs9_2(.din(w_dff_B_L8UPxx8e1_2),.dout(w_dff_B_PPiahgxs9_2),.clk(gclk));
	jdff dff_B_F2zmgtPn2_2(.din(w_dff_B_PPiahgxs9_2),.dout(w_dff_B_F2zmgtPn2_2),.clk(gclk));
	jdff dff_B_N8xjebfb1_2(.din(w_dff_B_F2zmgtPn2_2),.dout(w_dff_B_N8xjebfb1_2),.clk(gclk));
	jdff dff_A_tFCKOFNL4_1(.dout(w_dff_A_IlZsEDUK1_0),.din(w_dff_A_tFCKOFNL4_1),.clk(gclk));
	jdff dff_A_IlZsEDUK1_0(.dout(w_dff_A_CEcT4a6e9_0),.din(w_dff_A_IlZsEDUK1_0),.clk(gclk));
	jdff dff_A_CEcT4a6e9_0(.dout(w_dff_A_4VV4GkaV1_0),.din(w_dff_A_CEcT4a6e9_0),.clk(gclk));
	jdff dff_A_4VV4GkaV1_0(.dout(w_dff_A_2PBcT4QF6_0),.din(w_dff_A_4VV4GkaV1_0),.clk(gclk));
	jdff dff_A_2PBcT4QF6_0(.dout(w_dff_A_svF7vANG6_0),.din(w_dff_A_2PBcT4QF6_0),.clk(gclk));
	jdff dff_A_svF7vANG6_0(.dout(w_dff_A_xHISj5mx7_0),.din(w_dff_A_svF7vANG6_0),.clk(gclk));
	jdff dff_A_xHISj5mx7_0(.dout(w_dff_A_BMspYHVI9_0),.din(w_dff_A_xHISj5mx7_0),.clk(gclk));
	jdff dff_A_BMspYHVI9_0(.dout(w_dff_A_lnoOPcSL4_0),.din(w_dff_A_BMspYHVI9_0),.clk(gclk));
	jdff dff_A_lnoOPcSL4_0(.dout(w_dff_A_c6YR15Kn0_0),.din(w_dff_A_lnoOPcSL4_0),.clk(gclk));
	jdff dff_A_c6YR15Kn0_0(.dout(w_dff_A_FdUmNxvz7_0),.din(w_dff_A_c6YR15Kn0_0),.clk(gclk));
	jdff dff_A_FdUmNxvz7_0(.dout(w_dff_A_14FSDXLG3_0),.din(w_dff_A_FdUmNxvz7_0),.clk(gclk));
	jdff dff_A_14FSDXLG3_0(.dout(w_dff_A_DxmdopC61_0),.din(w_dff_A_14FSDXLG3_0),.clk(gclk));
	jdff dff_A_DxmdopC61_0(.dout(w_dff_A_q56tQ0zC5_0),.din(w_dff_A_DxmdopC61_0),.clk(gclk));
	jdff dff_A_q56tQ0zC5_0(.dout(w_dff_A_4GaniFXN0_0),.din(w_dff_A_q56tQ0zC5_0),.clk(gclk));
	jdff dff_A_4GaniFXN0_0(.dout(w_dff_A_Bs74xH8Y3_0),.din(w_dff_A_4GaniFXN0_0),.clk(gclk));
	jdff dff_A_Bs74xH8Y3_0(.dout(w_dff_A_M2SiTpMy0_0),.din(w_dff_A_Bs74xH8Y3_0),.clk(gclk));
	jdff dff_A_M2SiTpMy0_0(.dout(w_dff_A_9UBehGnl5_0),.din(w_dff_A_M2SiTpMy0_0),.clk(gclk));
	jdff dff_A_9UBehGnl5_0(.dout(w_dff_A_Q94LseRR7_0),.din(w_dff_A_9UBehGnl5_0),.clk(gclk));
	jdff dff_A_Q94LseRR7_0(.dout(w_dff_A_2hKHFtfk7_0),.din(w_dff_A_Q94LseRR7_0),.clk(gclk));
	jdff dff_A_2hKHFtfk7_0(.dout(w_dff_A_CWJCZpaH4_0),.din(w_dff_A_2hKHFtfk7_0),.clk(gclk));
	jdff dff_A_CWJCZpaH4_0(.dout(w_dff_A_ls03wzJm9_0),.din(w_dff_A_CWJCZpaH4_0),.clk(gclk));
	jdff dff_A_ls03wzJm9_0(.dout(w_dff_A_RdMGEhjR3_0),.din(w_dff_A_ls03wzJm9_0),.clk(gclk));
	jdff dff_A_RdMGEhjR3_0(.dout(w_dff_A_7XceqW1U3_0),.din(w_dff_A_RdMGEhjR3_0),.clk(gclk));
	jdff dff_A_7XceqW1U3_0(.dout(w_dff_A_LO1GnWZF9_0),.din(w_dff_A_7XceqW1U3_0),.clk(gclk));
	jdff dff_A_LO1GnWZF9_0(.dout(w_dff_A_W9PKCXPe5_0),.din(w_dff_A_LO1GnWZF9_0),.clk(gclk));
	jdff dff_A_W9PKCXPe5_0(.dout(w_dff_A_6oc6LFNX4_0),.din(w_dff_A_W9PKCXPe5_0),.clk(gclk));
	jdff dff_A_6oc6LFNX4_0(.dout(w_dff_A_54vrj7St8_0),.din(w_dff_A_6oc6LFNX4_0),.clk(gclk));
	jdff dff_A_54vrj7St8_0(.dout(G144),.din(w_dff_A_54vrj7St8_0),.clk(gclk));
	jdff dff_A_Bir94Gwe0_1(.dout(w_dff_A_adTFoNZk7_0),.din(w_dff_A_Bir94Gwe0_1),.clk(gclk));
	jdff dff_A_adTFoNZk7_0(.dout(w_dff_A_eBaIsSic1_0),.din(w_dff_A_adTFoNZk7_0),.clk(gclk));
	jdff dff_A_eBaIsSic1_0(.dout(w_dff_A_8RzHka1B2_0),.din(w_dff_A_eBaIsSic1_0),.clk(gclk));
	jdff dff_A_8RzHka1B2_0(.dout(w_dff_A_y9ZXT5La9_0),.din(w_dff_A_8RzHka1B2_0),.clk(gclk));
	jdff dff_A_y9ZXT5La9_0(.dout(w_dff_A_WuxbsWnc9_0),.din(w_dff_A_y9ZXT5La9_0),.clk(gclk));
	jdff dff_A_WuxbsWnc9_0(.dout(w_dff_A_QZ4T2PjB9_0),.din(w_dff_A_WuxbsWnc9_0),.clk(gclk));
	jdff dff_A_QZ4T2PjB9_0(.dout(w_dff_A_soBDb5fj5_0),.din(w_dff_A_QZ4T2PjB9_0),.clk(gclk));
	jdff dff_A_soBDb5fj5_0(.dout(w_dff_A_jh2zniJb6_0),.din(w_dff_A_soBDb5fj5_0),.clk(gclk));
	jdff dff_A_jh2zniJb6_0(.dout(w_dff_A_F0lzzu2m0_0),.din(w_dff_A_jh2zniJb6_0),.clk(gclk));
	jdff dff_A_F0lzzu2m0_0(.dout(w_dff_A_FQCsMyot8_0),.din(w_dff_A_F0lzzu2m0_0),.clk(gclk));
	jdff dff_A_FQCsMyot8_0(.dout(w_dff_A_buoWIpoR5_0),.din(w_dff_A_FQCsMyot8_0),.clk(gclk));
	jdff dff_A_buoWIpoR5_0(.dout(w_dff_A_HmLMOibi4_0),.din(w_dff_A_buoWIpoR5_0),.clk(gclk));
	jdff dff_A_HmLMOibi4_0(.dout(w_dff_A_uxw6RwgI6_0),.din(w_dff_A_HmLMOibi4_0),.clk(gclk));
	jdff dff_A_uxw6RwgI6_0(.dout(w_dff_A_qehoy7UX7_0),.din(w_dff_A_uxw6RwgI6_0),.clk(gclk));
	jdff dff_A_qehoy7UX7_0(.dout(w_dff_A_tpqGvAKw7_0),.din(w_dff_A_qehoy7UX7_0),.clk(gclk));
	jdff dff_A_tpqGvAKw7_0(.dout(w_dff_A_YoZ5tzuC2_0),.din(w_dff_A_tpqGvAKw7_0),.clk(gclk));
	jdff dff_A_YoZ5tzuC2_0(.dout(w_dff_A_Hjm9D9fg0_0),.din(w_dff_A_YoZ5tzuC2_0),.clk(gclk));
	jdff dff_A_Hjm9D9fg0_0(.dout(w_dff_A_BoDHA4QK7_0),.din(w_dff_A_Hjm9D9fg0_0),.clk(gclk));
	jdff dff_A_BoDHA4QK7_0(.dout(w_dff_A_ovB82ksM3_0),.din(w_dff_A_BoDHA4QK7_0),.clk(gclk));
	jdff dff_A_ovB82ksM3_0(.dout(w_dff_A_nzWHdgM34_0),.din(w_dff_A_ovB82ksM3_0),.clk(gclk));
	jdff dff_A_nzWHdgM34_0(.dout(w_dff_A_Xtpe54Fi3_0),.din(w_dff_A_nzWHdgM34_0),.clk(gclk));
	jdff dff_A_Xtpe54Fi3_0(.dout(w_dff_A_QtOT82I86_0),.din(w_dff_A_Xtpe54Fi3_0),.clk(gclk));
	jdff dff_A_QtOT82I86_0(.dout(w_dff_A_PKMcqa5r9_0),.din(w_dff_A_QtOT82I86_0),.clk(gclk));
	jdff dff_A_PKMcqa5r9_0(.dout(w_dff_A_2Z02vyXc3_0),.din(w_dff_A_PKMcqa5r9_0),.clk(gclk));
	jdff dff_A_2Z02vyXc3_0(.dout(w_dff_A_1aBOBSgY5_0),.din(w_dff_A_2Z02vyXc3_0),.clk(gclk));
	jdff dff_A_1aBOBSgY5_0(.dout(w_dff_A_6ElIMykj1_0),.din(w_dff_A_1aBOBSgY5_0),.clk(gclk));
	jdff dff_A_6ElIMykj1_0(.dout(w_dff_A_VFKfeA661_0),.din(w_dff_A_6ElIMykj1_0),.clk(gclk));
	jdff dff_A_VFKfeA661_0(.dout(G298),.din(w_dff_A_VFKfeA661_0),.clk(gclk));
	jdff dff_A_H773dteS1_1(.dout(w_dff_A_Wrb6XQ9M3_0),.din(w_dff_A_H773dteS1_1),.clk(gclk));
	jdff dff_A_Wrb6XQ9M3_0(.dout(w_dff_A_gjolEoZm8_0),.din(w_dff_A_Wrb6XQ9M3_0),.clk(gclk));
	jdff dff_A_gjolEoZm8_0(.dout(w_dff_A_cDiMoD0l6_0),.din(w_dff_A_gjolEoZm8_0),.clk(gclk));
	jdff dff_A_cDiMoD0l6_0(.dout(w_dff_A_pVAc7uwU2_0),.din(w_dff_A_cDiMoD0l6_0),.clk(gclk));
	jdff dff_A_pVAc7uwU2_0(.dout(w_dff_A_LSTP7cjW7_0),.din(w_dff_A_pVAc7uwU2_0),.clk(gclk));
	jdff dff_A_LSTP7cjW7_0(.dout(w_dff_A_sqniW66f4_0),.din(w_dff_A_LSTP7cjW7_0),.clk(gclk));
	jdff dff_A_sqniW66f4_0(.dout(w_dff_A_6dTVZnDz5_0),.din(w_dff_A_sqniW66f4_0),.clk(gclk));
	jdff dff_A_6dTVZnDz5_0(.dout(w_dff_A_NbDrMkrj4_0),.din(w_dff_A_6dTVZnDz5_0),.clk(gclk));
	jdff dff_A_NbDrMkrj4_0(.dout(w_dff_A_Xte8DpDg1_0),.din(w_dff_A_NbDrMkrj4_0),.clk(gclk));
	jdff dff_A_Xte8DpDg1_0(.dout(w_dff_A_qbbP2Bre2_0),.din(w_dff_A_Xte8DpDg1_0),.clk(gclk));
	jdff dff_A_qbbP2Bre2_0(.dout(w_dff_A_Js5nZOvU1_0),.din(w_dff_A_qbbP2Bre2_0),.clk(gclk));
	jdff dff_A_Js5nZOvU1_0(.dout(w_dff_A_QfOule055_0),.din(w_dff_A_Js5nZOvU1_0),.clk(gclk));
	jdff dff_A_QfOule055_0(.dout(w_dff_A_wXdDOOIp2_0),.din(w_dff_A_QfOule055_0),.clk(gclk));
	jdff dff_A_wXdDOOIp2_0(.dout(w_dff_A_5cRvcW8U0_0),.din(w_dff_A_wXdDOOIp2_0),.clk(gclk));
	jdff dff_A_5cRvcW8U0_0(.dout(w_dff_A_eSnQq50H8_0),.din(w_dff_A_5cRvcW8U0_0),.clk(gclk));
	jdff dff_A_eSnQq50H8_0(.dout(w_dff_A_u36tr0Uk9_0),.din(w_dff_A_eSnQq50H8_0),.clk(gclk));
	jdff dff_A_u36tr0Uk9_0(.dout(w_dff_A_LyD1bGZw7_0),.din(w_dff_A_u36tr0Uk9_0),.clk(gclk));
	jdff dff_A_LyD1bGZw7_0(.dout(w_dff_A_9ZGrWXR51_0),.din(w_dff_A_LyD1bGZw7_0),.clk(gclk));
	jdff dff_A_9ZGrWXR51_0(.dout(w_dff_A_IezzxeHx2_0),.din(w_dff_A_9ZGrWXR51_0),.clk(gclk));
	jdff dff_A_IezzxeHx2_0(.dout(w_dff_A_gTe6RvbS9_0),.din(w_dff_A_IezzxeHx2_0),.clk(gclk));
	jdff dff_A_gTe6RvbS9_0(.dout(w_dff_A_nsvwWbP60_0),.din(w_dff_A_gTe6RvbS9_0),.clk(gclk));
	jdff dff_A_nsvwWbP60_0(.dout(w_dff_A_ePmEMqIg2_0),.din(w_dff_A_nsvwWbP60_0),.clk(gclk));
	jdff dff_A_ePmEMqIg2_0(.dout(w_dff_A_eCCmkl9E7_0),.din(w_dff_A_ePmEMqIg2_0),.clk(gclk));
	jdff dff_A_eCCmkl9E7_0(.dout(w_dff_A_LAdfQCgz7_0),.din(w_dff_A_eCCmkl9E7_0),.clk(gclk));
	jdff dff_A_LAdfQCgz7_0(.dout(w_dff_A_x3SHnhVE1_0),.din(w_dff_A_LAdfQCgz7_0),.clk(gclk));
	jdff dff_A_x3SHnhVE1_0(.dout(w_dff_A_MjbNilE46_0),.din(w_dff_A_x3SHnhVE1_0),.clk(gclk));
	jdff dff_A_MjbNilE46_0(.dout(w_dff_A_8g2vocKL1_0),.din(w_dff_A_MjbNilE46_0),.clk(gclk));
	jdff dff_A_8g2vocKL1_0(.dout(G973),.din(w_dff_A_8g2vocKL1_0),.clk(gclk));
	jdff dff_A_H1rIXdYd7_1(.dout(w_dff_A_GXWBBTVX5_0),.din(w_dff_A_H1rIXdYd7_1),.clk(gclk));
	jdff dff_A_GXWBBTVX5_0(.dout(w_dff_A_XpN5hJdD3_0),.din(w_dff_A_GXWBBTVX5_0),.clk(gclk));
	jdff dff_A_XpN5hJdD3_0(.dout(w_dff_A_m7DBhqto6_0),.din(w_dff_A_XpN5hJdD3_0),.clk(gclk));
	jdff dff_A_m7DBhqto6_0(.dout(w_dff_A_7aWAnjDg8_0),.din(w_dff_A_m7DBhqto6_0),.clk(gclk));
	jdff dff_A_7aWAnjDg8_0(.dout(w_dff_A_wSEwcVj96_0),.din(w_dff_A_7aWAnjDg8_0),.clk(gclk));
	jdff dff_A_wSEwcVj96_0(.dout(w_dff_A_w9lVZ12u0_0),.din(w_dff_A_wSEwcVj96_0),.clk(gclk));
	jdff dff_A_w9lVZ12u0_0(.dout(w_dff_A_MPHbYqjQ9_0),.din(w_dff_A_w9lVZ12u0_0),.clk(gclk));
	jdff dff_A_MPHbYqjQ9_0(.dout(w_dff_A_JznfRGiE9_0),.din(w_dff_A_MPHbYqjQ9_0),.clk(gclk));
	jdff dff_A_JznfRGiE9_0(.dout(w_dff_A_pyKXWd1D1_0),.din(w_dff_A_JznfRGiE9_0),.clk(gclk));
	jdff dff_A_pyKXWd1D1_0(.dout(w_dff_A_ZD85smjf6_0),.din(w_dff_A_pyKXWd1D1_0),.clk(gclk));
	jdff dff_A_ZD85smjf6_0(.dout(w_dff_A_GW7ScZib9_0),.din(w_dff_A_ZD85smjf6_0),.clk(gclk));
	jdff dff_A_GW7ScZib9_0(.dout(w_dff_A_Uug7XAZ92_0),.din(w_dff_A_GW7ScZib9_0),.clk(gclk));
	jdff dff_A_Uug7XAZ92_0(.dout(w_dff_A_nKbHBH6W0_0),.din(w_dff_A_Uug7XAZ92_0),.clk(gclk));
	jdff dff_A_nKbHBH6W0_0(.dout(w_dff_A_zxN7p3io2_0),.din(w_dff_A_nKbHBH6W0_0),.clk(gclk));
	jdff dff_A_zxN7p3io2_0(.dout(w_dff_A_mpS3mQ7V7_0),.din(w_dff_A_zxN7p3io2_0),.clk(gclk));
	jdff dff_A_mpS3mQ7V7_0(.dout(w_dff_A_O8nC4jad7_0),.din(w_dff_A_mpS3mQ7V7_0),.clk(gclk));
	jdff dff_A_O8nC4jad7_0(.dout(w_dff_A_YHcjhaOu1_0),.din(w_dff_A_O8nC4jad7_0),.clk(gclk));
	jdff dff_A_YHcjhaOu1_0(.dout(w_dff_A_ndtwybAt6_0),.din(w_dff_A_YHcjhaOu1_0),.clk(gclk));
	jdff dff_A_ndtwybAt6_0(.dout(w_dff_A_b8kuF6Xe6_0),.din(w_dff_A_ndtwybAt6_0),.clk(gclk));
	jdff dff_A_b8kuF6Xe6_0(.dout(w_dff_A_Mwrz6Mvt2_0),.din(w_dff_A_b8kuF6Xe6_0),.clk(gclk));
	jdff dff_A_Mwrz6Mvt2_0(.dout(w_dff_A_DuFWqoLP1_0),.din(w_dff_A_Mwrz6Mvt2_0),.clk(gclk));
	jdff dff_A_DuFWqoLP1_0(.dout(w_dff_A_mcOIk3Fx2_0),.din(w_dff_A_DuFWqoLP1_0),.clk(gclk));
	jdff dff_A_mcOIk3Fx2_0(.dout(w_dff_A_5DZM0TFf2_0),.din(w_dff_A_mcOIk3Fx2_0),.clk(gclk));
	jdff dff_A_5DZM0TFf2_0(.dout(w_dff_A_7iyGSHtR8_0),.din(w_dff_A_5DZM0TFf2_0),.clk(gclk));
	jdff dff_A_7iyGSHtR8_0(.dout(w_dff_A_TajBF7E89_0),.din(w_dff_A_7iyGSHtR8_0),.clk(gclk));
	jdff dff_A_TajBF7E89_0(.dout(w_dff_A_MNmoIlqo7_0),.din(w_dff_A_TajBF7E89_0),.clk(gclk));
	jdff dff_A_MNmoIlqo7_0(.dout(G594),.din(w_dff_A_MNmoIlqo7_0),.clk(gclk));
	jdff dff_A_QA8TyQ3f3_1(.dout(w_dff_A_QBROjjOd0_0),.din(w_dff_A_QA8TyQ3f3_1),.clk(gclk));
	jdff dff_A_QBROjjOd0_0(.dout(w_dff_A_c9iPnlNf3_0),.din(w_dff_A_QBROjjOd0_0),.clk(gclk));
	jdff dff_A_c9iPnlNf3_0(.dout(w_dff_A_s4LwXeps4_0),.din(w_dff_A_c9iPnlNf3_0),.clk(gclk));
	jdff dff_A_s4LwXeps4_0(.dout(w_dff_A_4JoHyEzQ7_0),.din(w_dff_A_s4LwXeps4_0),.clk(gclk));
	jdff dff_A_4JoHyEzQ7_0(.dout(w_dff_A_9z6bFZaj2_0),.din(w_dff_A_4JoHyEzQ7_0),.clk(gclk));
	jdff dff_A_9z6bFZaj2_0(.dout(w_dff_A_7OVFCuU01_0),.din(w_dff_A_9z6bFZaj2_0),.clk(gclk));
	jdff dff_A_7OVFCuU01_0(.dout(w_dff_A_7TwucoQR3_0),.din(w_dff_A_7OVFCuU01_0),.clk(gclk));
	jdff dff_A_7TwucoQR3_0(.dout(w_dff_A_58Um3fd75_0),.din(w_dff_A_7TwucoQR3_0),.clk(gclk));
	jdff dff_A_58Um3fd75_0(.dout(w_dff_A_LkdHHjQe9_0),.din(w_dff_A_58Um3fd75_0),.clk(gclk));
	jdff dff_A_LkdHHjQe9_0(.dout(w_dff_A_mVil7j4e0_0),.din(w_dff_A_LkdHHjQe9_0),.clk(gclk));
	jdff dff_A_mVil7j4e0_0(.dout(w_dff_A_o2CqpAva4_0),.din(w_dff_A_mVil7j4e0_0),.clk(gclk));
	jdff dff_A_o2CqpAva4_0(.dout(w_dff_A_mjBr6zl40_0),.din(w_dff_A_o2CqpAva4_0),.clk(gclk));
	jdff dff_A_mjBr6zl40_0(.dout(w_dff_A_ryB8kxCI7_0),.din(w_dff_A_mjBr6zl40_0),.clk(gclk));
	jdff dff_A_ryB8kxCI7_0(.dout(w_dff_A_qBtYsWeu9_0),.din(w_dff_A_ryB8kxCI7_0),.clk(gclk));
	jdff dff_A_qBtYsWeu9_0(.dout(w_dff_A_5UHIoTlL9_0),.din(w_dff_A_qBtYsWeu9_0),.clk(gclk));
	jdff dff_A_5UHIoTlL9_0(.dout(w_dff_A_JJL6Zjyo9_0),.din(w_dff_A_5UHIoTlL9_0),.clk(gclk));
	jdff dff_A_JJL6Zjyo9_0(.dout(w_dff_A_s7bcHlga8_0),.din(w_dff_A_JJL6Zjyo9_0),.clk(gclk));
	jdff dff_A_s7bcHlga8_0(.dout(w_dff_A_S2Taeel45_0),.din(w_dff_A_s7bcHlga8_0),.clk(gclk));
	jdff dff_A_S2Taeel45_0(.dout(w_dff_A_ByNIFjWL6_0),.din(w_dff_A_S2Taeel45_0),.clk(gclk));
	jdff dff_A_ByNIFjWL6_0(.dout(w_dff_A_Qwf1AUPT8_0),.din(w_dff_A_ByNIFjWL6_0),.clk(gclk));
	jdff dff_A_Qwf1AUPT8_0(.dout(w_dff_A_z9w1kiHo4_0),.din(w_dff_A_Qwf1AUPT8_0),.clk(gclk));
	jdff dff_A_z9w1kiHo4_0(.dout(w_dff_A_NpZ04Uab0_0),.din(w_dff_A_z9w1kiHo4_0),.clk(gclk));
	jdff dff_A_NpZ04Uab0_0(.dout(w_dff_A_KNT9MsG93_0),.din(w_dff_A_NpZ04Uab0_0),.clk(gclk));
	jdff dff_A_KNT9MsG93_0(.dout(w_dff_A_ibWsWtvQ8_0),.din(w_dff_A_KNT9MsG93_0),.clk(gclk));
	jdff dff_A_ibWsWtvQ8_0(.dout(w_dff_A_7780QqlZ4_0),.din(w_dff_A_ibWsWtvQ8_0),.clk(gclk));
	jdff dff_A_7780QqlZ4_0(.dout(w_dff_A_SyA7bhbB9_0),.din(w_dff_A_7780QqlZ4_0),.clk(gclk));
	jdff dff_A_SyA7bhbB9_0(.dout(G599),.din(w_dff_A_SyA7bhbB9_0),.clk(gclk));
	jdff dff_A_HCUTE1hH8_1(.dout(w_dff_A_D2th1dxC8_0),.din(w_dff_A_HCUTE1hH8_1),.clk(gclk));
	jdff dff_A_D2th1dxC8_0(.dout(w_dff_A_zQc6KNTr9_0),.din(w_dff_A_D2th1dxC8_0),.clk(gclk));
	jdff dff_A_zQc6KNTr9_0(.dout(w_dff_A_WFdFNGRX2_0),.din(w_dff_A_zQc6KNTr9_0),.clk(gclk));
	jdff dff_A_WFdFNGRX2_0(.dout(w_dff_A_u17W9g6y4_0),.din(w_dff_A_WFdFNGRX2_0),.clk(gclk));
	jdff dff_A_u17W9g6y4_0(.dout(w_dff_A_zNnRUM9D8_0),.din(w_dff_A_u17W9g6y4_0),.clk(gclk));
	jdff dff_A_zNnRUM9D8_0(.dout(w_dff_A_84A0Ie8H4_0),.din(w_dff_A_zNnRUM9D8_0),.clk(gclk));
	jdff dff_A_84A0Ie8H4_0(.dout(w_dff_A_dLbxZUUK2_0),.din(w_dff_A_84A0Ie8H4_0),.clk(gclk));
	jdff dff_A_dLbxZUUK2_0(.dout(w_dff_A_899P7Vdo1_0),.din(w_dff_A_dLbxZUUK2_0),.clk(gclk));
	jdff dff_A_899P7Vdo1_0(.dout(w_dff_A_K275nXcx4_0),.din(w_dff_A_899P7Vdo1_0),.clk(gclk));
	jdff dff_A_K275nXcx4_0(.dout(w_dff_A_56RexwDu0_0),.din(w_dff_A_K275nXcx4_0),.clk(gclk));
	jdff dff_A_56RexwDu0_0(.dout(w_dff_A_SWxtiXqn4_0),.din(w_dff_A_56RexwDu0_0),.clk(gclk));
	jdff dff_A_SWxtiXqn4_0(.dout(w_dff_A_PQ6AwPzD4_0),.din(w_dff_A_SWxtiXqn4_0),.clk(gclk));
	jdff dff_A_PQ6AwPzD4_0(.dout(w_dff_A_mR56OXx80_0),.din(w_dff_A_PQ6AwPzD4_0),.clk(gclk));
	jdff dff_A_mR56OXx80_0(.dout(w_dff_A_43qxwe5n4_0),.din(w_dff_A_mR56OXx80_0),.clk(gclk));
	jdff dff_A_43qxwe5n4_0(.dout(w_dff_A_lM4cQxuK8_0),.din(w_dff_A_43qxwe5n4_0),.clk(gclk));
	jdff dff_A_lM4cQxuK8_0(.dout(w_dff_A_P02dXyHs2_0),.din(w_dff_A_lM4cQxuK8_0),.clk(gclk));
	jdff dff_A_P02dXyHs2_0(.dout(w_dff_A_gPnPbhlk2_0),.din(w_dff_A_P02dXyHs2_0),.clk(gclk));
	jdff dff_A_gPnPbhlk2_0(.dout(w_dff_A_pjPlahOv5_0),.din(w_dff_A_gPnPbhlk2_0),.clk(gclk));
	jdff dff_A_pjPlahOv5_0(.dout(w_dff_A_sd4yuauN4_0),.din(w_dff_A_pjPlahOv5_0),.clk(gclk));
	jdff dff_A_sd4yuauN4_0(.dout(w_dff_A_pMGsOJDe5_0),.din(w_dff_A_sd4yuauN4_0),.clk(gclk));
	jdff dff_A_pMGsOJDe5_0(.dout(w_dff_A_WIdxZpcC7_0),.din(w_dff_A_pMGsOJDe5_0),.clk(gclk));
	jdff dff_A_WIdxZpcC7_0(.dout(w_dff_A_7edUgzrp8_0),.din(w_dff_A_WIdxZpcC7_0),.clk(gclk));
	jdff dff_A_7edUgzrp8_0(.dout(w_dff_A_eGFurfib8_0),.din(w_dff_A_7edUgzrp8_0),.clk(gclk));
	jdff dff_A_eGFurfib8_0(.dout(w_dff_A_cnAalqim5_0),.din(w_dff_A_eGFurfib8_0),.clk(gclk));
	jdff dff_A_cnAalqim5_0(.dout(w_dff_A_s8XYea018_0),.din(w_dff_A_cnAalqim5_0),.clk(gclk));
	jdff dff_A_s8XYea018_0(.dout(w_dff_A_SgELGMm62_0),.din(w_dff_A_s8XYea018_0),.clk(gclk));
	jdff dff_A_SgELGMm62_0(.dout(G600),.din(w_dff_A_SgELGMm62_0),.clk(gclk));
	jdff dff_A_B5zaQhi98_1(.dout(w_dff_A_kw8rr8Nl7_0),.din(w_dff_A_B5zaQhi98_1),.clk(gclk));
	jdff dff_A_kw8rr8Nl7_0(.dout(w_dff_A_KYBBMnJJ6_0),.din(w_dff_A_kw8rr8Nl7_0),.clk(gclk));
	jdff dff_A_KYBBMnJJ6_0(.dout(w_dff_A_aHi9xvcF3_0),.din(w_dff_A_KYBBMnJJ6_0),.clk(gclk));
	jdff dff_A_aHi9xvcF3_0(.dout(w_dff_A_roJLgMVP1_0),.din(w_dff_A_aHi9xvcF3_0),.clk(gclk));
	jdff dff_A_roJLgMVP1_0(.dout(w_dff_A_3JDIISQ00_0),.din(w_dff_A_roJLgMVP1_0),.clk(gclk));
	jdff dff_A_3JDIISQ00_0(.dout(w_dff_A_1cM70qXy2_0),.din(w_dff_A_3JDIISQ00_0),.clk(gclk));
	jdff dff_A_1cM70qXy2_0(.dout(w_dff_A_SytAfQnO7_0),.din(w_dff_A_1cM70qXy2_0),.clk(gclk));
	jdff dff_A_SytAfQnO7_0(.dout(w_dff_A_oX47xxQO7_0),.din(w_dff_A_SytAfQnO7_0),.clk(gclk));
	jdff dff_A_oX47xxQO7_0(.dout(w_dff_A_Dl72Iv3P9_0),.din(w_dff_A_oX47xxQO7_0),.clk(gclk));
	jdff dff_A_Dl72Iv3P9_0(.dout(w_dff_A_R5giQd9G7_0),.din(w_dff_A_Dl72Iv3P9_0),.clk(gclk));
	jdff dff_A_R5giQd9G7_0(.dout(w_dff_A_RRJqQEfR2_0),.din(w_dff_A_R5giQd9G7_0),.clk(gclk));
	jdff dff_A_RRJqQEfR2_0(.dout(w_dff_A_U31w5LeJ4_0),.din(w_dff_A_RRJqQEfR2_0),.clk(gclk));
	jdff dff_A_U31w5LeJ4_0(.dout(w_dff_A_wELXTeHb9_0),.din(w_dff_A_U31w5LeJ4_0),.clk(gclk));
	jdff dff_A_wELXTeHb9_0(.dout(w_dff_A_McTbMLZN9_0),.din(w_dff_A_wELXTeHb9_0),.clk(gclk));
	jdff dff_A_McTbMLZN9_0(.dout(w_dff_A_XtRoVTfS9_0),.din(w_dff_A_McTbMLZN9_0),.clk(gclk));
	jdff dff_A_XtRoVTfS9_0(.dout(w_dff_A_qYN43HMH4_0),.din(w_dff_A_XtRoVTfS9_0),.clk(gclk));
	jdff dff_A_qYN43HMH4_0(.dout(w_dff_A_Zds1RHDK6_0),.din(w_dff_A_qYN43HMH4_0),.clk(gclk));
	jdff dff_A_Zds1RHDK6_0(.dout(w_dff_A_2Ywc9JdV4_0),.din(w_dff_A_Zds1RHDK6_0),.clk(gclk));
	jdff dff_A_2Ywc9JdV4_0(.dout(w_dff_A_sdLUWOH84_0),.din(w_dff_A_2Ywc9JdV4_0),.clk(gclk));
	jdff dff_A_sdLUWOH84_0(.dout(w_dff_A_cT8CFlQB5_0),.din(w_dff_A_sdLUWOH84_0),.clk(gclk));
	jdff dff_A_cT8CFlQB5_0(.dout(w_dff_A_yJ8iasqj9_0),.din(w_dff_A_cT8CFlQB5_0),.clk(gclk));
	jdff dff_A_yJ8iasqj9_0(.dout(w_dff_A_VqBUACDa0_0),.din(w_dff_A_yJ8iasqj9_0),.clk(gclk));
	jdff dff_A_VqBUACDa0_0(.dout(w_dff_A_2tZH7ec25_0),.din(w_dff_A_VqBUACDa0_0),.clk(gclk));
	jdff dff_A_2tZH7ec25_0(.dout(w_dff_A_skYbwueA9_0),.din(w_dff_A_2tZH7ec25_0),.clk(gclk));
	jdff dff_A_skYbwueA9_0(.dout(w_dff_A_dr2oqWfh1_0),.din(w_dff_A_skYbwueA9_0),.clk(gclk));
	jdff dff_A_dr2oqWfh1_0(.dout(w_dff_A_BubwsMNS6_0),.din(w_dff_A_dr2oqWfh1_0),.clk(gclk));
	jdff dff_A_BubwsMNS6_0(.dout(G601),.din(w_dff_A_BubwsMNS6_0),.clk(gclk));
	jdff dff_A_wsRicFXl5_1(.dout(w_dff_A_lMMs7hJv3_0),.din(w_dff_A_wsRicFXl5_1),.clk(gclk));
	jdff dff_A_lMMs7hJv3_0(.dout(w_dff_A_4tkXWEsA3_0),.din(w_dff_A_lMMs7hJv3_0),.clk(gclk));
	jdff dff_A_4tkXWEsA3_0(.dout(w_dff_A_DfnJXHkz0_0),.din(w_dff_A_4tkXWEsA3_0),.clk(gclk));
	jdff dff_A_DfnJXHkz0_0(.dout(w_dff_A_whsLhFcA3_0),.din(w_dff_A_DfnJXHkz0_0),.clk(gclk));
	jdff dff_A_whsLhFcA3_0(.dout(w_dff_A_5OYSFGq80_0),.din(w_dff_A_whsLhFcA3_0),.clk(gclk));
	jdff dff_A_5OYSFGq80_0(.dout(w_dff_A_NnUSuJHM0_0),.din(w_dff_A_5OYSFGq80_0),.clk(gclk));
	jdff dff_A_NnUSuJHM0_0(.dout(w_dff_A_7DCEQMkB8_0),.din(w_dff_A_NnUSuJHM0_0),.clk(gclk));
	jdff dff_A_7DCEQMkB8_0(.dout(w_dff_A_htuo9FSx2_0),.din(w_dff_A_7DCEQMkB8_0),.clk(gclk));
	jdff dff_A_htuo9FSx2_0(.dout(w_dff_A_k97GJOOY8_0),.din(w_dff_A_htuo9FSx2_0),.clk(gclk));
	jdff dff_A_k97GJOOY8_0(.dout(w_dff_A_i9basHgR1_0),.din(w_dff_A_k97GJOOY8_0),.clk(gclk));
	jdff dff_A_i9basHgR1_0(.dout(w_dff_A_Q1JFKpPs7_0),.din(w_dff_A_i9basHgR1_0),.clk(gclk));
	jdff dff_A_Q1JFKpPs7_0(.dout(w_dff_A_ufocaaEK6_0),.din(w_dff_A_Q1JFKpPs7_0),.clk(gclk));
	jdff dff_A_ufocaaEK6_0(.dout(w_dff_A_WEbBZDyb9_0),.din(w_dff_A_ufocaaEK6_0),.clk(gclk));
	jdff dff_A_WEbBZDyb9_0(.dout(w_dff_A_xRzkgRa43_0),.din(w_dff_A_WEbBZDyb9_0),.clk(gclk));
	jdff dff_A_xRzkgRa43_0(.dout(w_dff_A_votJOWvl2_0),.din(w_dff_A_xRzkgRa43_0),.clk(gclk));
	jdff dff_A_votJOWvl2_0(.dout(w_dff_A_BkKx0VBP8_0),.din(w_dff_A_votJOWvl2_0),.clk(gclk));
	jdff dff_A_BkKx0VBP8_0(.dout(w_dff_A_RHncwQeX4_0),.din(w_dff_A_BkKx0VBP8_0),.clk(gclk));
	jdff dff_A_RHncwQeX4_0(.dout(w_dff_A_wK8pW0BO6_0),.din(w_dff_A_RHncwQeX4_0),.clk(gclk));
	jdff dff_A_wK8pW0BO6_0(.dout(w_dff_A_IirWNDv19_0),.din(w_dff_A_wK8pW0BO6_0),.clk(gclk));
	jdff dff_A_IirWNDv19_0(.dout(w_dff_A_8WJSC0E14_0),.din(w_dff_A_IirWNDv19_0),.clk(gclk));
	jdff dff_A_8WJSC0E14_0(.dout(w_dff_A_5CoaPKEU5_0),.din(w_dff_A_8WJSC0E14_0),.clk(gclk));
	jdff dff_A_5CoaPKEU5_0(.dout(w_dff_A_xp6pNGAQ7_0),.din(w_dff_A_5CoaPKEU5_0),.clk(gclk));
	jdff dff_A_xp6pNGAQ7_0(.dout(w_dff_A_VDwXIE4E5_0),.din(w_dff_A_xp6pNGAQ7_0),.clk(gclk));
	jdff dff_A_VDwXIE4E5_0(.dout(w_dff_A_RO5r0N2e7_0),.din(w_dff_A_VDwXIE4E5_0),.clk(gclk));
	jdff dff_A_RO5r0N2e7_0(.dout(w_dff_A_6xRw4hWc7_0),.din(w_dff_A_RO5r0N2e7_0),.clk(gclk));
	jdff dff_A_6xRw4hWc7_0(.dout(w_dff_A_Ke9X6fvb2_0),.din(w_dff_A_6xRw4hWc7_0),.clk(gclk));
	jdff dff_A_Ke9X6fvb2_0(.dout(G602),.din(w_dff_A_Ke9X6fvb2_0),.clk(gclk));
	jdff dff_A_5wc4wnAA5_1(.dout(w_dff_A_2qNRjnX37_0),.din(w_dff_A_5wc4wnAA5_1),.clk(gclk));
	jdff dff_A_2qNRjnX37_0(.dout(w_dff_A_c1bnQw2Z8_0),.din(w_dff_A_2qNRjnX37_0),.clk(gclk));
	jdff dff_A_c1bnQw2Z8_0(.dout(w_dff_A_86uySLNB7_0),.din(w_dff_A_c1bnQw2Z8_0),.clk(gclk));
	jdff dff_A_86uySLNB7_0(.dout(w_dff_A_Q5jBzqUI3_0),.din(w_dff_A_86uySLNB7_0),.clk(gclk));
	jdff dff_A_Q5jBzqUI3_0(.dout(w_dff_A_ueIqyRhO2_0),.din(w_dff_A_Q5jBzqUI3_0),.clk(gclk));
	jdff dff_A_ueIqyRhO2_0(.dout(w_dff_A_S6ZOIxqh7_0),.din(w_dff_A_ueIqyRhO2_0),.clk(gclk));
	jdff dff_A_S6ZOIxqh7_0(.dout(w_dff_A_Z4aiqFLt1_0),.din(w_dff_A_S6ZOIxqh7_0),.clk(gclk));
	jdff dff_A_Z4aiqFLt1_0(.dout(w_dff_A_Rnt4wmwV6_0),.din(w_dff_A_Z4aiqFLt1_0),.clk(gclk));
	jdff dff_A_Rnt4wmwV6_0(.dout(w_dff_A_Zjg07G7H0_0),.din(w_dff_A_Rnt4wmwV6_0),.clk(gclk));
	jdff dff_A_Zjg07G7H0_0(.dout(w_dff_A_BAbJkfWu6_0),.din(w_dff_A_Zjg07G7H0_0),.clk(gclk));
	jdff dff_A_BAbJkfWu6_0(.dout(w_dff_A_N71oDIZv2_0),.din(w_dff_A_BAbJkfWu6_0),.clk(gclk));
	jdff dff_A_N71oDIZv2_0(.dout(w_dff_A_gTcxvjPt7_0),.din(w_dff_A_N71oDIZv2_0),.clk(gclk));
	jdff dff_A_gTcxvjPt7_0(.dout(w_dff_A_51cDu1Xn7_0),.din(w_dff_A_gTcxvjPt7_0),.clk(gclk));
	jdff dff_A_51cDu1Xn7_0(.dout(w_dff_A_UidG5YXB7_0),.din(w_dff_A_51cDu1Xn7_0),.clk(gclk));
	jdff dff_A_UidG5YXB7_0(.dout(w_dff_A_7DMLheaJ2_0),.din(w_dff_A_UidG5YXB7_0),.clk(gclk));
	jdff dff_A_7DMLheaJ2_0(.dout(w_dff_A_9Y6AxvSH9_0),.din(w_dff_A_7DMLheaJ2_0),.clk(gclk));
	jdff dff_A_9Y6AxvSH9_0(.dout(w_dff_A_6WHusuzJ2_0),.din(w_dff_A_9Y6AxvSH9_0),.clk(gclk));
	jdff dff_A_6WHusuzJ2_0(.dout(w_dff_A_63aDm5KU0_0),.din(w_dff_A_6WHusuzJ2_0),.clk(gclk));
	jdff dff_A_63aDm5KU0_0(.dout(w_dff_A_Uct3V7rS5_0),.din(w_dff_A_63aDm5KU0_0),.clk(gclk));
	jdff dff_A_Uct3V7rS5_0(.dout(w_dff_A_vStka29A1_0),.din(w_dff_A_Uct3V7rS5_0),.clk(gclk));
	jdff dff_A_vStka29A1_0(.dout(w_dff_A_WHgyj6Ee1_0),.din(w_dff_A_vStka29A1_0),.clk(gclk));
	jdff dff_A_WHgyj6Ee1_0(.dout(w_dff_A_0RG0TIzb9_0),.din(w_dff_A_WHgyj6Ee1_0),.clk(gclk));
	jdff dff_A_0RG0TIzb9_0(.dout(w_dff_A_kQjhXkOH3_0),.din(w_dff_A_0RG0TIzb9_0),.clk(gclk));
	jdff dff_A_kQjhXkOH3_0(.dout(w_dff_A_UaIFjqUD1_0),.din(w_dff_A_kQjhXkOH3_0),.clk(gclk));
	jdff dff_A_UaIFjqUD1_0(.dout(w_dff_A_S8sqmpI97_0),.din(w_dff_A_UaIFjqUD1_0),.clk(gclk));
	jdff dff_A_S8sqmpI97_0(.dout(w_dff_A_4uwWC8Qm6_0),.din(w_dff_A_S8sqmpI97_0),.clk(gclk));
	jdff dff_A_4uwWC8Qm6_0(.dout(G603),.din(w_dff_A_4uwWC8Qm6_0),.clk(gclk));
	jdff dff_A_iFcdHZpN8_1(.dout(w_dff_A_Mx1X726q8_0),.din(w_dff_A_iFcdHZpN8_1),.clk(gclk));
	jdff dff_A_Mx1X726q8_0(.dout(w_dff_A_iPviCIs37_0),.din(w_dff_A_Mx1X726q8_0),.clk(gclk));
	jdff dff_A_iPviCIs37_0(.dout(w_dff_A_7eI7kD5X9_0),.din(w_dff_A_iPviCIs37_0),.clk(gclk));
	jdff dff_A_7eI7kD5X9_0(.dout(w_dff_A_1pBmZcdT4_0),.din(w_dff_A_7eI7kD5X9_0),.clk(gclk));
	jdff dff_A_1pBmZcdT4_0(.dout(w_dff_A_ai3mTQ3z0_0),.din(w_dff_A_1pBmZcdT4_0),.clk(gclk));
	jdff dff_A_ai3mTQ3z0_0(.dout(w_dff_A_kdGJnj6t1_0),.din(w_dff_A_ai3mTQ3z0_0),.clk(gclk));
	jdff dff_A_kdGJnj6t1_0(.dout(w_dff_A_ECnEZZwQ9_0),.din(w_dff_A_kdGJnj6t1_0),.clk(gclk));
	jdff dff_A_ECnEZZwQ9_0(.dout(w_dff_A_MMDbtLqk1_0),.din(w_dff_A_ECnEZZwQ9_0),.clk(gclk));
	jdff dff_A_MMDbtLqk1_0(.dout(w_dff_A_ePWq3UBc0_0),.din(w_dff_A_MMDbtLqk1_0),.clk(gclk));
	jdff dff_A_ePWq3UBc0_0(.dout(w_dff_A_5oqBe5EH2_0),.din(w_dff_A_ePWq3UBc0_0),.clk(gclk));
	jdff dff_A_5oqBe5EH2_0(.dout(w_dff_A_6t9HqlM23_0),.din(w_dff_A_5oqBe5EH2_0),.clk(gclk));
	jdff dff_A_6t9HqlM23_0(.dout(w_dff_A_07OyTkp68_0),.din(w_dff_A_6t9HqlM23_0),.clk(gclk));
	jdff dff_A_07OyTkp68_0(.dout(w_dff_A_co11kp2N7_0),.din(w_dff_A_07OyTkp68_0),.clk(gclk));
	jdff dff_A_co11kp2N7_0(.dout(w_dff_A_bcLdXrdQ7_0),.din(w_dff_A_co11kp2N7_0),.clk(gclk));
	jdff dff_A_bcLdXrdQ7_0(.dout(w_dff_A_9WLKyMj34_0),.din(w_dff_A_bcLdXrdQ7_0),.clk(gclk));
	jdff dff_A_9WLKyMj34_0(.dout(w_dff_A_nsxR5qEy0_0),.din(w_dff_A_9WLKyMj34_0),.clk(gclk));
	jdff dff_A_nsxR5qEy0_0(.dout(w_dff_A_GWJhRBhU5_0),.din(w_dff_A_nsxR5qEy0_0),.clk(gclk));
	jdff dff_A_GWJhRBhU5_0(.dout(w_dff_A_iIfeIdj21_0),.din(w_dff_A_GWJhRBhU5_0),.clk(gclk));
	jdff dff_A_iIfeIdj21_0(.dout(w_dff_A_0kLKVHac6_0),.din(w_dff_A_iIfeIdj21_0),.clk(gclk));
	jdff dff_A_0kLKVHac6_0(.dout(w_dff_A_3IeRq1wj9_0),.din(w_dff_A_0kLKVHac6_0),.clk(gclk));
	jdff dff_A_3IeRq1wj9_0(.dout(w_dff_A_F1Xq0dlN9_0),.din(w_dff_A_3IeRq1wj9_0),.clk(gclk));
	jdff dff_A_F1Xq0dlN9_0(.dout(w_dff_A_n7TI19Rg7_0),.din(w_dff_A_F1Xq0dlN9_0),.clk(gclk));
	jdff dff_A_n7TI19Rg7_0(.dout(w_dff_A_bREk1lkZ4_0),.din(w_dff_A_n7TI19Rg7_0),.clk(gclk));
	jdff dff_A_bREk1lkZ4_0(.dout(w_dff_A_RGwOJmSC2_0),.din(w_dff_A_bREk1lkZ4_0),.clk(gclk));
	jdff dff_A_RGwOJmSC2_0(.dout(w_dff_A_Bztaqpdq6_0),.din(w_dff_A_RGwOJmSC2_0),.clk(gclk));
	jdff dff_A_Bztaqpdq6_0(.dout(w_dff_A_hOzwgkhi2_0),.din(w_dff_A_Bztaqpdq6_0),.clk(gclk));
	jdff dff_A_hOzwgkhi2_0(.dout(G604),.din(w_dff_A_hOzwgkhi2_0),.clk(gclk));
	jdff dff_A_6Sa7Xvf97_1(.dout(w_dff_A_Uf2jSV5b7_0),.din(w_dff_A_6Sa7Xvf97_1),.clk(gclk));
	jdff dff_A_Uf2jSV5b7_0(.dout(w_dff_A_rZfsHOJt3_0),.din(w_dff_A_Uf2jSV5b7_0),.clk(gclk));
	jdff dff_A_rZfsHOJt3_0(.dout(w_dff_A_RpUp8Alr6_0),.din(w_dff_A_rZfsHOJt3_0),.clk(gclk));
	jdff dff_A_RpUp8Alr6_0(.dout(w_dff_A_SFJlVtsc9_0),.din(w_dff_A_RpUp8Alr6_0),.clk(gclk));
	jdff dff_A_SFJlVtsc9_0(.dout(w_dff_A_KehKZ3l47_0),.din(w_dff_A_SFJlVtsc9_0),.clk(gclk));
	jdff dff_A_KehKZ3l47_0(.dout(w_dff_A_PzvtLay25_0),.din(w_dff_A_KehKZ3l47_0),.clk(gclk));
	jdff dff_A_PzvtLay25_0(.dout(w_dff_A_210zCSDV5_0),.din(w_dff_A_PzvtLay25_0),.clk(gclk));
	jdff dff_A_210zCSDV5_0(.dout(w_dff_A_SZfDYcQl6_0),.din(w_dff_A_210zCSDV5_0),.clk(gclk));
	jdff dff_A_SZfDYcQl6_0(.dout(w_dff_A_RPdSk9mK4_0),.din(w_dff_A_SZfDYcQl6_0),.clk(gclk));
	jdff dff_A_RPdSk9mK4_0(.dout(w_dff_A_naZQSBVL9_0),.din(w_dff_A_RPdSk9mK4_0),.clk(gclk));
	jdff dff_A_naZQSBVL9_0(.dout(w_dff_A_uetRDmOr3_0),.din(w_dff_A_naZQSBVL9_0),.clk(gclk));
	jdff dff_A_uetRDmOr3_0(.dout(w_dff_A_NBEnAyvh3_0),.din(w_dff_A_uetRDmOr3_0),.clk(gclk));
	jdff dff_A_NBEnAyvh3_0(.dout(w_dff_A_VW0juebU2_0),.din(w_dff_A_NBEnAyvh3_0),.clk(gclk));
	jdff dff_A_VW0juebU2_0(.dout(w_dff_A_ts3Kubfk9_0),.din(w_dff_A_VW0juebU2_0),.clk(gclk));
	jdff dff_A_ts3Kubfk9_0(.dout(w_dff_A_id7yic8Z6_0),.din(w_dff_A_ts3Kubfk9_0),.clk(gclk));
	jdff dff_A_id7yic8Z6_0(.dout(w_dff_A_TFTHJbxc8_0),.din(w_dff_A_id7yic8Z6_0),.clk(gclk));
	jdff dff_A_TFTHJbxc8_0(.dout(w_dff_A_emAsT7vR0_0),.din(w_dff_A_TFTHJbxc8_0),.clk(gclk));
	jdff dff_A_emAsT7vR0_0(.dout(w_dff_A_3ALw9M8d9_0),.din(w_dff_A_emAsT7vR0_0),.clk(gclk));
	jdff dff_A_3ALw9M8d9_0(.dout(w_dff_A_KmpkTfpE0_0),.din(w_dff_A_3ALw9M8d9_0),.clk(gclk));
	jdff dff_A_KmpkTfpE0_0(.dout(w_dff_A_qfEDelqT2_0),.din(w_dff_A_KmpkTfpE0_0),.clk(gclk));
	jdff dff_A_qfEDelqT2_0(.dout(w_dff_A_6BCkUk5Y0_0),.din(w_dff_A_qfEDelqT2_0),.clk(gclk));
	jdff dff_A_6BCkUk5Y0_0(.dout(w_dff_A_XMjGGtsr5_0),.din(w_dff_A_6BCkUk5Y0_0),.clk(gclk));
	jdff dff_A_XMjGGtsr5_0(.dout(w_dff_A_hD3yCD5v0_0),.din(w_dff_A_XMjGGtsr5_0),.clk(gclk));
	jdff dff_A_hD3yCD5v0_0(.dout(w_dff_A_jNVRaYYi8_0),.din(w_dff_A_hD3yCD5v0_0),.clk(gclk));
	jdff dff_A_jNVRaYYi8_0(.dout(w_dff_A_l75UpMBg1_0),.din(w_dff_A_jNVRaYYi8_0),.clk(gclk));
	jdff dff_A_l75UpMBg1_0(.dout(w_dff_A_6Aq8FD5u4_0),.din(w_dff_A_l75UpMBg1_0),.clk(gclk));
	jdff dff_A_6Aq8FD5u4_0(.dout(G611),.din(w_dff_A_6Aq8FD5u4_0),.clk(gclk));
	jdff dff_A_aWb3Bder3_1(.dout(w_dff_A_37qidPkF0_0),.din(w_dff_A_aWb3Bder3_1),.clk(gclk));
	jdff dff_A_37qidPkF0_0(.dout(w_dff_A_Q6fFJPZb4_0),.din(w_dff_A_37qidPkF0_0),.clk(gclk));
	jdff dff_A_Q6fFJPZb4_0(.dout(w_dff_A_uRyH7K3K9_0),.din(w_dff_A_Q6fFJPZb4_0),.clk(gclk));
	jdff dff_A_uRyH7K3K9_0(.dout(w_dff_A_4NRPImzl0_0),.din(w_dff_A_uRyH7K3K9_0),.clk(gclk));
	jdff dff_A_4NRPImzl0_0(.dout(w_dff_A_BRWbNyB77_0),.din(w_dff_A_4NRPImzl0_0),.clk(gclk));
	jdff dff_A_BRWbNyB77_0(.dout(w_dff_A_XWy7JglP7_0),.din(w_dff_A_BRWbNyB77_0),.clk(gclk));
	jdff dff_A_XWy7JglP7_0(.dout(w_dff_A_61JnoIBW2_0),.din(w_dff_A_XWy7JglP7_0),.clk(gclk));
	jdff dff_A_61JnoIBW2_0(.dout(w_dff_A_ZCJvXGZe1_0),.din(w_dff_A_61JnoIBW2_0),.clk(gclk));
	jdff dff_A_ZCJvXGZe1_0(.dout(w_dff_A_1q4FCxbs0_0),.din(w_dff_A_ZCJvXGZe1_0),.clk(gclk));
	jdff dff_A_1q4FCxbs0_0(.dout(w_dff_A_eA0dgkzs4_0),.din(w_dff_A_1q4FCxbs0_0),.clk(gclk));
	jdff dff_A_eA0dgkzs4_0(.dout(w_dff_A_YRIjOYI94_0),.din(w_dff_A_eA0dgkzs4_0),.clk(gclk));
	jdff dff_A_YRIjOYI94_0(.dout(w_dff_A_zTNwIrWC7_0),.din(w_dff_A_YRIjOYI94_0),.clk(gclk));
	jdff dff_A_zTNwIrWC7_0(.dout(w_dff_A_kmrbAwfV0_0),.din(w_dff_A_zTNwIrWC7_0),.clk(gclk));
	jdff dff_A_kmrbAwfV0_0(.dout(w_dff_A_Ox8EP8me8_0),.din(w_dff_A_kmrbAwfV0_0),.clk(gclk));
	jdff dff_A_Ox8EP8me8_0(.dout(w_dff_A_sndsVV9d8_0),.din(w_dff_A_Ox8EP8me8_0),.clk(gclk));
	jdff dff_A_sndsVV9d8_0(.dout(w_dff_A_O5KbiIx65_0),.din(w_dff_A_sndsVV9d8_0),.clk(gclk));
	jdff dff_A_O5KbiIx65_0(.dout(w_dff_A_aLKeHqcp8_0),.din(w_dff_A_O5KbiIx65_0),.clk(gclk));
	jdff dff_A_aLKeHqcp8_0(.dout(w_dff_A_nR60EwYh4_0),.din(w_dff_A_aLKeHqcp8_0),.clk(gclk));
	jdff dff_A_nR60EwYh4_0(.dout(w_dff_A_RIjzj0jG8_0),.din(w_dff_A_nR60EwYh4_0),.clk(gclk));
	jdff dff_A_RIjzj0jG8_0(.dout(w_dff_A_yVTjbZxL4_0),.din(w_dff_A_RIjzj0jG8_0),.clk(gclk));
	jdff dff_A_yVTjbZxL4_0(.dout(w_dff_A_lNo6GqT56_0),.din(w_dff_A_yVTjbZxL4_0),.clk(gclk));
	jdff dff_A_lNo6GqT56_0(.dout(w_dff_A_qYjj9DpR2_0),.din(w_dff_A_lNo6GqT56_0),.clk(gclk));
	jdff dff_A_qYjj9DpR2_0(.dout(w_dff_A_n629pjA98_0),.din(w_dff_A_qYjj9DpR2_0),.clk(gclk));
	jdff dff_A_n629pjA98_0(.dout(w_dff_A_dSWu2JMH3_0),.din(w_dff_A_n629pjA98_0),.clk(gclk));
	jdff dff_A_dSWu2JMH3_0(.dout(w_dff_A_IuCpVn6p1_0),.din(w_dff_A_dSWu2JMH3_0),.clk(gclk));
	jdff dff_A_IuCpVn6p1_0(.dout(w_dff_A_24FkzvG86_0),.din(w_dff_A_IuCpVn6p1_0),.clk(gclk));
	jdff dff_A_24FkzvG86_0(.dout(G612),.din(w_dff_A_24FkzvG86_0),.clk(gclk));
	jdff dff_A_EJSBV4R46_2(.dout(w_dff_A_TIELi39v9_0),.din(w_dff_A_EJSBV4R46_2),.clk(gclk));
	jdff dff_A_TIELi39v9_0(.dout(w_dff_A_GVghg9bM9_0),.din(w_dff_A_TIELi39v9_0),.clk(gclk));
	jdff dff_A_GVghg9bM9_0(.dout(w_dff_A_SDmsdrjL1_0),.din(w_dff_A_GVghg9bM9_0),.clk(gclk));
	jdff dff_A_SDmsdrjL1_0(.dout(w_dff_A_aKCiX8WE3_0),.din(w_dff_A_SDmsdrjL1_0),.clk(gclk));
	jdff dff_A_aKCiX8WE3_0(.dout(w_dff_A_Pwk7GOeq1_0),.din(w_dff_A_aKCiX8WE3_0),.clk(gclk));
	jdff dff_A_Pwk7GOeq1_0(.dout(w_dff_A_ttDfJGRe8_0),.din(w_dff_A_Pwk7GOeq1_0),.clk(gclk));
	jdff dff_A_ttDfJGRe8_0(.dout(w_dff_A_o9ORt5Of5_0),.din(w_dff_A_ttDfJGRe8_0),.clk(gclk));
	jdff dff_A_o9ORt5Of5_0(.dout(w_dff_A_PTjsbeIh6_0),.din(w_dff_A_o9ORt5Of5_0),.clk(gclk));
	jdff dff_A_PTjsbeIh6_0(.dout(w_dff_A_Ke32ivLL0_0),.din(w_dff_A_PTjsbeIh6_0),.clk(gclk));
	jdff dff_A_Ke32ivLL0_0(.dout(w_dff_A_DOM2kqXq7_0),.din(w_dff_A_Ke32ivLL0_0),.clk(gclk));
	jdff dff_A_DOM2kqXq7_0(.dout(w_dff_A_MQZhC69F6_0),.din(w_dff_A_DOM2kqXq7_0),.clk(gclk));
	jdff dff_A_MQZhC69F6_0(.dout(w_dff_A_HalNvWIm0_0),.din(w_dff_A_MQZhC69F6_0),.clk(gclk));
	jdff dff_A_HalNvWIm0_0(.dout(w_dff_A_Ggisu0AC2_0),.din(w_dff_A_HalNvWIm0_0),.clk(gclk));
	jdff dff_A_Ggisu0AC2_0(.dout(w_dff_A_FF7QhOBt5_0),.din(w_dff_A_Ggisu0AC2_0),.clk(gclk));
	jdff dff_A_FF7QhOBt5_0(.dout(w_dff_A_4oIQ4CII8_0),.din(w_dff_A_FF7QhOBt5_0),.clk(gclk));
	jdff dff_A_4oIQ4CII8_0(.dout(w_dff_A_5o70XSRu5_0),.din(w_dff_A_4oIQ4CII8_0),.clk(gclk));
	jdff dff_A_5o70XSRu5_0(.dout(w_dff_A_6NclDxdl4_0),.din(w_dff_A_5o70XSRu5_0),.clk(gclk));
	jdff dff_A_6NclDxdl4_0(.dout(w_dff_A_x1pekYJs3_0),.din(w_dff_A_6NclDxdl4_0),.clk(gclk));
	jdff dff_A_x1pekYJs3_0(.dout(w_dff_A_NtouRkLw1_0),.din(w_dff_A_x1pekYJs3_0),.clk(gclk));
	jdff dff_A_NtouRkLw1_0(.dout(w_dff_A_kpY8J51a4_0),.din(w_dff_A_NtouRkLw1_0),.clk(gclk));
	jdff dff_A_kpY8J51a4_0(.dout(w_dff_A_6Vpx65ZK3_0),.din(w_dff_A_kpY8J51a4_0),.clk(gclk));
	jdff dff_A_6Vpx65ZK3_0(.dout(w_dff_A_TS2hjwmc2_0),.din(w_dff_A_6Vpx65ZK3_0),.clk(gclk));
	jdff dff_A_TS2hjwmc2_0(.dout(w_dff_A_ZGNjP5nh3_0),.din(w_dff_A_TS2hjwmc2_0),.clk(gclk));
	jdff dff_A_ZGNjP5nh3_0(.dout(w_dff_A_pIyMq1T61_0),.din(w_dff_A_ZGNjP5nh3_0),.clk(gclk));
	jdff dff_A_pIyMq1T61_0(.dout(w_dff_A_psfa3IAA7_0),.din(w_dff_A_pIyMq1T61_0),.clk(gclk));
	jdff dff_A_psfa3IAA7_0(.dout(w_dff_A_Qz3g3XdO7_0),.din(w_dff_A_psfa3IAA7_0),.clk(gclk));
	jdff dff_A_Qz3g3XdO7_0(.dout(G810),.din(w_dff_A_Qz3g3XdO7_0),.clk(gclk));
	jdff dff_A_C0wtGoAE3_1(.dout(w_dff_A_2h0KxOym5_0),.din(w_dff_A_C0wtGoAE3_1),.clk(gclk));
	jdff dff_A_2h0KxOym5_0(.dout(w_dff_A_OWrkQTk52_0),.din(w_dff_A_2h0KxOym5_0),.clk(gclk));
	jdff dff_A_OWrkQTk52_0(.dout(w_dff_A_AlY58BUz8_0),.din(w_dff_A_OWrkQTk52_0),.clk(gclk));
	jdff dff_A_AlY58BUz8_0(.dout(w_dff_A_ht2SxEAa9_0),.din(w_dff_A_AlY58BUz8_0),.clk(gclk));
	jdff dff_A_ht2SxEAa9_0(.dout(w_dff_A_G8akYSOr8_0),.din(w_dff_A_ht2SxEAa9_0),.clk(gclk));
	jdff dff_A_G8akYSOr8_0(.dout(w_dff_A_4QQeJKHz5_0),.din(w_dff_A_G8akYSOr8_0),.clk(gclk));
	jdff dff_A_4QQeJKHz5_0(.dout(w_dff_A_7OrlUbxO2_0),.din(w_dff_A_4QQeJKHz5_0),.clk(gclk));
	jdff dff_A_7OrlUbxO2_0(.dout(w_dff_A_XK02slre7_0),.din(w_dff_A_7OrlUbxO2_0),.clk(gclk));
	jdff dff_A_XK02slre7_0(.dout(w_dff_A_CTDGqpaF6_0),.din(w_dff_A_XK02slre7_0),.clk(gclk));
	jdff dff_A_CTDGqpaF6_0(.dout(w_dff_A_KzwYXyOC3_0),.din(w_dff_A_CTDGqpaF6_0),.clk(gclk));
	jdff dff_A_KzwYXyOC3_0(.dout(w_dff_A_7GQrzYxo1_0),.din(w_dff_A_KzwYXyOC3_0),.clk(gclk));
	jdff dff_A_7GQrzYxo1_0(.dout(w_dff_A_4azZmAGj3_0),.din(w_dff_A_7GQrzYxo1_0),.clk(gclk));
	jdff dff_A_4azZmAGj3_0(.dout(w_dff_A_VIUP5geH9_0),.din(w_dff_A_4azZmAGj3_0),.clk(gclk));
	jdff dff_A_VIUP5geH9_0(.dout(w_dff_A_a1kw8kaT5_0),.din(w_dff_A_VIUP5geH9_0),.clk(gclk));
	jdff dff_A_a1kw8kaT5_0(.dout(w_dff_A_qrAtofiT7_0),.din(w_dff_A_a1kw8kaT5_0),.clk(gclk));
	jdff dff_A_qrAtofiT7_0(.dout(w_dff_A_1eeGagY18_0),.din(w_dff_A_qrAtofiT7_0),.clk(gclk));
	jdff dff_A_1eeGagY18_0(.dout(w_dff_A_OE1VORvO6_0),.din(w_dff_A_1eeGagY18_0),.clk(gclk));
	jdff dff_A_OE1VORvO6_0(.dout(w_dff_A_RkzhPTIv2_0),.din(w_dff_A_OE1VORvO6_0),.clk(gclk));
	jdff dff_A_RkzhPTIv2_0(.dout(w_dff_A_tEab5lgN4_0),.din(w_dff_A_RkzhPTIv2_0),.clk(gclk));
	jdff dff_A_tEab5lgN4_0(.dout(w_dff_A_tMXXNwq55_0),.din(w_dff_A_tEab5lgN4_0),.clk(gclk));
	jdff dff_A_tMXXNwq55_0(.dout(w_dff_A_wRTpQvsx3_0),.din(w_dff_A_tMXXNwq55_0),.clk(gclk));
	jdff dff_A_wRTpQvsx3_0(.dout(w_dff_A_Wo3NGruI6_0),.din(w_dff_A_wRTpQvsx3_0),.clk(gclk));
	jdff dff_A_Wo3NGruI6_0(.dout(w_dff_A_UwlsSxj38_0),.din(w_dff_A_Wo3NGruI6_0),.clk(gclk));
	jdff dff_A_UwlsSxj38_0(.dout(w_dff_A_HRvzKhzK6_0),.din(w_dff_A_UwlsSxj38_0),.clk(gclk));
	jdff dff_A_HRvzKhzK6_0(.dout(w_dff_A_7FtUQ8he6_0),.din(w_dff_A_HRvzKhzK6_0),.clk(gclk));
	jdff dff_A_7FtUQ8he6_0(.dout(w_dff_A_e1gUUK8D8_0),.din(w_dff_A_7FtUQ8he6_0),.clk(gclk));
	jdff dff_A_e1gUUK8D8_0(.dout(G848),.din(w_dff_A_e1gUUK8D8_0),.clk(gclk));
	jdff dff_A_ZcBak8Wz0_1(.dout(w_dff_A_d6Zmd3nD4_0),.din(w_dff_A_ZcBak8Wz0_1),.clk(gclk));
	jdff dff_A_d6Zmd3nD4_0(.dout(w_dff_A_V6mA00sq6_0),.din(w_dff_A_d6Zmd3nD4_0),.clk(gclk));
	jdff dff_A_V6mA00sq6_0(.dout(w_dff_A_WUdKXxqu6_0),.din(w_dff_A_V6mA00sq6_0),.clk(gclk));
	jdff dff_A_WUdKXxqu6_0(.dout(w_dff_A_53xY64Mt6_0),.din(w_dff_A_WUdKXxqu6_0),.clk(gclk));
	jdff dff_A_53xY64Mt6_0(.dout(w_dff_A_vnmyTlvZ1_0),.din(w_dff_A_53xY64Mt6_0),.clk(gclk));
	jdff dff_A_vnmyTlvZ1_0(.dout(w_dff_A_T4Ly5fbj3_0),.din(w_dff_A_vnmyTlvZ1_0),.clk(gclk));
	jdff dff_A_T4Ly5fbj3_0(.dout(w_dff_A_9MWoWyTM4_0),.din(w_dff_A_T4Ly5fbj3_0),.clk(gclk));
	jdff dff_A_9MWoWyTM4_0(.dout(w_dff_A_oHiwbgD08_0),.din(w_dff_A_9MWoWyTM4_0),.clk(gclk));
	jdff dff_A_oHiwbgD08_0(.dout(w_dff_A_66mEnOOU3_0),.din(w_dff_A_oHiwbgD08_0),.clk(gclk));
	jdff dff_A_66mEnOOU3_0(.dout(w_dff_A_7p4kKu1b7_0),.din(w_dff_A_66mEnOOU3_0),.clk(gclk));
	jdff dff_A_7p4kKu1b7_0(.dout(w_dff_A_LY0ED1MY8_0),.din(w_dff_A_7p4kKu1b7_0),.clk(gclk));
	jdff dff_A_LY0ED1MY8_0(.dout(w_dff_A_P5siTwNL5_0),.din(w_dff_A_LY0ED1MY8_0),.clk(gclk));
	jdff dff_A_P5siTwNL5_0(.dout(w_dff_A_GJIPEppz7_0),.din(w_dff_A_P5siTwNL5_0),.clk(gclk));
	jdff dff_A_GJIPEppz7_0(.dout(w_dff_A_OE62B7CQ3_0),.din(w_dff_A_GJIPEppz7_0),.clk(gclk));
	jdff dff_A_OE62B7CQ3_0(.dout(w_dff_A_XJidZEOv9_0),.din(w_dff_A_OE62B7CQ3_0),.clk(gclk));
	jdff dff_A_XJidZEOv9_0(.dout(w_dff_A_TGSrF0Bo2_0),.din(w_dff_A_XJidZEOv9_0),.clk(gclk));
	jdff dff_A_TGSrF0Bo2_0(.dout(w_dff_A_wBHJ4t5C7_0),.din(w_dff_A_TGSrF0Bo2_0),.clk(gclk));
	jdff dff_A_wBHJ4t5C7_0(.dout(w_dff_A_QUJtWDbP0_0),.din(w_dff_A_wBHJ4t5C7_0),.clk(gclk));
	jdff dff_A_QUJtWDbP0_0(.dout(w_dff_A_WrGC2sDE4_0),.din(w_dff_A_QUJtWDbP0_0),.clk(gclk));
	jdff dff_A_WrGC2sDE4_0(.dout(w_dff_A_CeFX0CnR4_0),.din(w_dff_A_WrGC2sDE4_0),.clk(gclk));
	jdff dff_A_CeFX0CnR4_0(.dout(w_dff_A_75vGWjBU8_0),.din(w_dff_A_CeFX0CnR4_0),.clk(gclk));
	jdff dff_A_75vGWjBU8_0(.dout(w_dff_A_1S16eqBq7_0),.din(w_dff_A_75vGWjBU8_0),.clk(gclk));
	jdff dff_A_1S16eqBq7_0(.dout(w_dff_A_cry6awpr7_0),.din(w_dff_A_1S16eqBq7_0),.clk(gclk));
	jdff dff_A_cry6awpr7_0(.dout(w_dff_A_Ni5dg4iN7_0),.din(w_dff_A_cry6awpr7_0),.clk(gclk));
	jdff dff_A_Ni5dg4iN7_0(.dout(w_dff_A_IRJ1jwDa5_0),.din(w_dff_A_Ni5dg4iN7_0),.clk(gclk));
	jdff dff_A_IRJ1jwDa5_0(.dout(w_dff_A_q7VcqtXf2_0),.din(w_dff_A_IRJ1jwDa5_0),.clk(gclk));
	jdff dff_A_q7VcqtXf2_0(.dout(G849),.din(w_dff_A_q7VcqtXf2_0),.clk(gclk));
	jdff dff_A_11gMwd6c1_1(.dout(w_dff_A_DgSuzRmG0_0),.din(w_dff_A_11gMwd6c1_1),.clk(gclk));
	jdff dff_A_DgSuzRmG0_0(.dout(w_dff_A_w0iVHi3J9_0),.din(w_dff_A_DgSuzRmG0_0),.clk(gclk));
	jdff dff_A_w0iVHi3J9_0(.dout(w_dff_A_GT5xiU5F3_0),.din(w_dff_A_w0iVHi3J9_0),.clk(gclk));
	jdff dff_A_GT5xiU5F3_0(.dout(w_dff_A_MyiXWURi6_0),.din(w_dff_A_GT5xiU5F3_0),.clk(gclk));
	jdff dff_A_MyiXWURi6_0(.dout(w_dff_A_YzaojHkK1_0),.din(w_dff_A_MyiXWURi6_0),.clk(gclk));
	jdff dff_A_YzaojHkK1_0(.dout(w_dff_A_HVNic8zf5_0),.din(w_dff_A_YzaojHkK1_0),.clk(gclk));
	jdff dff_A_HVNic8zf5_0(.dout(w_dff_A_oYJ2F1f43_0),.din(w_dff_A_HVNic8zf5_0),.clk(gclk));
	jdff dff_A_oYJ2F1f43_0(.dout(w_dff_A_E2hWJkdu2_0),.din(w_dff_A_oYJ2F1f43_0),.clk(gclk));
	jdff dff_A_E2hWJkdu2_0(.dout(w_dff_A_4kt8yL2l0_0),.din(w_dff_A_E2hWJkdu2_0),.clk(gclk));
	jdff dff_A_4kt8yL2l0_0(.dout(w_dff_A_idHBsHLM5_0),.din(w_dff_A_4kt8yL2l0_0),.clk(gclk));
	jdff dff_A_idHBsHLM5_0(.dout(w_dff_A_5eWmLYEj9_0),.din(w_dff_A_idHBsHLM5_0),.clk(gclk));
	jdff dff_A_5eWmLYEj9_0(.dout(w_dff_A_HEnZeIni7_0),.din(w_dff_A_5eWmLYEj9_0),.clk(gclk));
	jdff dff_A_HEnZeIni7_0(.dout(w_dff_A_iJ242T1M6_0),.din(w_dff_A_HEnZeIni7_0),.clk(gclk));
	jdff dff_A_iJ242T1M6_0(.dout(w_dff_A_sYliSE2D2_0),.din(w_dff_A_iJ242T1M6_0),.clk(gclk));
	jdff dff_A_sYliSE2D2_0(.dout(w_dff_A_8csViICh1_0),.din(w_dff_A_sYliSE2D2_0),.clk(gclk));
	jdff dff_A_8csViICh1_0(.dout(w_dff_A_ucVAyJuO7_0),.din(w_dff_A_8csViICh1_0),.clk(gclk));
	jdff dff_A_ucVAyJuO7_0(.dout(w_dff_A_uEBK0OSV7_0),.din(w_dff_A_ucVAyJuO7_0),.clk(gclk));
	jdff dff_A_uEBK0OSV7_0(.dout(w_dff_A_eDAbYZIk2_0),.din(w_dff_A_uEBK0OSV7_0),.clk(gclk));
	jdff dff_A_eDAbYZIk2_0(.dout(w_dff_A_EUz0yJH81_0),.din(w_dff_A_eDAbYZIk2_0),.clk(gclk));
	jdff dff_A_EUz0yJH81_0(.dout(w_dff_A_X6D4NQWF5_0),.din(w_dff_A_EUz0yJH81_0),.clk(gclk));
	jdff dff_A_X6D4NQWF5_0(.dout(w_dff_A_Jq7iJYdi3_0),.din(w_dff_A_X6D4NQWF5_0),.clk(gclk));
	jdff dff_A_Jq7iJYdi3_0(.dout(w_dff_A_Yjc51a5W8_0),.din(w_dff_A_Jq7iJYdi3_0),.clk(gclk));
	jdff dff_A_Yjc51a5W8_0(.dout(w_dff_A_kWey6ZCY1_0),.din(w_dff_A_Yjc51a5W8_0),.clk(gclk));
	jdff dff_A_kWey6ZCY1_0(.dout(w_dff_A_aIATRkWV5_0),.din(w_dff_A_kWey6ZCY1_0),.clk(gclk));
	jdff dff_A_aIATRkWV5_0(.dout(w_dff_A_JnfrM3eY5_0),.din(w_dff_A_aIATRkWV5_0),.clk(gclk));
	jdff dff_A_JnfrM3eY5_0(.dout(w_dff_A_b0kcHwIx9_0),.din(w_dff_A_JnfrM3eY5_0),.clk(gclk));
	jdff dff_A_b0kcHwIx9_0(.dout(G850),.din(w_dff_A_b0kcHwIx9_0),.clk(gclk));
	jdff dff_A_Yhp1kSkX5_1(.dout(w_dff_A_4755lNO00_0),.din(w_dff_A_Yhp1kSkX5_1),.clk(gclk));
	jdff dff_A_4755lNO00_0(.dout(w_dff_A_eJ6AB6SP3_0),.din(w_dff_A_4755lNO00_0),.clk(gclk));
	jdff dff_A_eJ6AB6SP3_0(.dout(w_dff_A_jIxzoZVo2_0),.din(w_dff_A_eJ6AB6SP3_0),.clk(gclk));
	jdff dff_A_jIxzoZVo2_0(.dout(w_dff_A_31G2phhd7_0),.din(w_dff_A_jIxzoZVo2_0),.clk(gclk));
	jdff dff_A_31G2phhd7_0(.dout(w_dff_A_DhUeKY8a0_0),.din(w_dff_A_31G2phhd7_0),.clk(gclk));
	jdff dff_A_DhUeKY8a0_0(.dout(w_dff_A_FADsnsv75_0),.din(w_dff_A_DhUeKY8a0_0),.clk(gclk));
	jdff dff_A_FADsnsv75_0(.dout(w_dff_A_nVlY46uf7_0),.din(w_dff_A_FADsnsv75_0),.clk(gclk));
	jdff dff_A_nVlY46uf7_0(.dout(w_dff_A_2P1Z4ldK9_0),.din(w_dff_A_nVlY46uf7_0),.clk(gclk));
	jdff dff_A_2P1Z4ldK9_0(.dout(w_dff_A_HjlgrXy65_0),.din(w_dff_A_2P1Z4ldK9_0),.clk(gclk));
	jdff dff_A_HjlgrXy65_0(.dout(w_dff_A_IR4yVBWR5_0),.din(w_dff_A_HjlgrXy65_0),.clk(gclk));
	jdff dff_A_IR4yVBWR5_0(.dout(w_dff_A_TwUAFyaG0_0),.din(w_dff_A_IR4yVBWR5_0),.clk(gclk));
	jdff dff_A_TwUAFyaG0_0(.dout(w_dff_A_hp0ZPgsW7_0),.din(w_dff_A_TwUAFyaG0_0),.clk(gclk));
	jdff dff_A_hp0ZPgsW7_0(.dout(w_dff_A_CzJUzp0U8_0),.din(w_dff_A_hp0ZPgsW7_0),.clk(gclk));
	jdff dff_A_CzJUzp0U8_0(.dout(w_dff_A_y3DPTehL1_0),.din(w_dff_A_CzJUzp0U8_0),.clk(gclk));
	jdff dff_A_y3DPTehL1_0(.dout(w_dff_A_8LL1JtOT2_0),.din(w_dff_A_y3DPTehL1_0),.clk(gclk));
	jdff dff_A_8LL1JtOT2_0(.dout(w_dff_A_nKeFnkHY4_0),.din(w_dff_A_8LL1JtOT2_0),.clk(gclk));
	jdff dff_A_nKeFnkHY4_0(.dout(w_dff_A_JzsBgQVP9_0),.din(w_dff_A_nKeFnkHY4_0),.clk(gclk));
	jdff dff_A_JzsBgQVP9_0(.dout(w_dff_A_aeXoUm8T5_0),.din(w_dff_A_JzsBgQVP9_0),.clk(gclk));
	jdff dff_A_aeXoUm8T5_0(.dout(w_dff_A_oONrYMeZ5_0),.din(w_dff_A_aeXoUm8T5_0),.clk(gclk));
	jdff dff_A_oONrYMeZ5_0(.dout(w_dff_A_mfi7YCDQ4_0),.din(w_dff_A_oONrYMeZ5_0),.clk(gclk));
	jdff dff_A_mfi7YCDQ4_0(.dout(w_dff_A_6S7CztCU1_0),.din(w_dff_A_mfi7YCDQ4_0),.clk(gclk));
	jdff dff_A_6S7CztCU1_0(.dout(w_dff_A_exCZ1ihX1_0),.din(w_dff_A_6S7CztCU1_0),.clk(gclk));
	jdff dff_A_exCZ1ihX1_0(.dout(w_dff_A_rskND1Rz4_0),.din(w_dff_A_exCZ1ihX1_0),.clk(gclk));
	jdff dff_A_rskND1Rz4_0(.dout(w_dff_A_uin5GKpW9_0),.din(w_dff_A_rskND1Rz4_0),.clk(gclk));
	jdff dff_A_uin5GKpW9_0(.dout(w_dff_A_JRV5moa65_0),.din(w_dff_A_uin5GKpW9_0),.clk(gclk));
	jdff dff_A_JRV5moa65_0(.dout(w_dff_A_gJJjhMvl0_0),.din(w_dff_A_JRV5moa65_0),.clk(gclk));
	jdff dff_A_gJJjhMvl0_0(.dout(G851),.din(w_dff_A_gJJjhMvl0_0),.clk(gclk));
	jdff dff_A_yO5mAeIh3_2(.dout(w_dff_A_RjRfhNgA7_0),.din(w_dff_A_yO5mAeIh3_2),.clk(gclk));
	jdff dff_A_RjRfhNgA7_0(.dout(w_dff_A_8GFNQy1I5_0),.din(w_dff_A_RjRfhNgA7_0),.clk(gclk));
	jdff dff_A_8GFNQy1I5_0(.dout(w_dff_A_wVLADo1z7_0),.din(w_dff_A_8GFNQy1I5_0),.clk(gclk));
	jdff dff_A_wVLADo1z7_0(.dout(w_dff_A_8q1uKPao5_0),.din(w_dff_A_wVLADo1z7_0),.clk(gclk));
	jdff dff_A_8q1uKPao5_0(.dout(w_dff_A_Ks2GVdeT5_0),.din(w_dff_A_8q1uKPao5_0),.clk(gclk));
	jdff dff_A_Ks2GVdeT5_0(.dout(w_dff_A_1a5rZWHF6_0),.din(w_dff_A_Ks2GVdeT5_0),.clk(gclk));
	jdff dff_A_1a5rZWHF6_0(.dout(w_dff_A_iswYPrAg8_0),.din(w_dff_A_1a5rZWHF6_0),.clk(gclk));
	jdff dff_A_iswYPrAg8_0(.dout(w_dff_A_jzWxOYOT5_0),.din(w_dff_A_iswYPrAg8_0),.clk(gclk));
	jdff dff_A_jzWxOYOT5_0(.dout(w_dff_A_nPgekng83_0),.din(w_dff_A_jzWxOYOT5_0),.clk(gclk));
	jdff dff_A_nPgekng83_0(.dout(w_dff_A_tEMX9oRN9_0),.din(w_dff_A_nPgekng83_0),.clk(gclk));
	jdff dff_A_tEMX9oRN9_0(.dout(w_dff_A_TI09GShc2_0),.din(w_dff_A_tEMX9oRN9_0),.clk(gclk));
	jdff dff_A_TI09GShc2_0(.dout(w_dff_A_PL6kwVX03_0),.din(w_dff_A_TI09GShc2_0),.clk(gclk));
	jdff dff_A_PL6kwVX03_0(.dout(w_dff_A_WCvWDdPG7_0),.din(w_dff_A_PL6kwVX03_0),.clk(gclk));
	jdff dff_A_WCvWDdPG7_0(.dout(w_dff_A_1OhX25aX6_0),.din(w_dff_A_WCvWDdPG7_0),.clk(gclk));
	jdff dff_A_1OhX25aX6_0(.dout(w_dff_A_rNtBoynd0_0),.din(w_dff_A_1OhX25aX6_0),.clk(gclk));
	jdff dff_A_rNtBoynd0_0(.dout(w_dff_A_3D7ljEMI2_0),.din(w_dff_A_rNtBoynd0_0),.clk(gclk));
	jdff dff_A_3D7ljEMI2_0(.dout(w_dff_A_LvzGJYUi9_0),.din(w_dff_A_3D7ljEMI2_0),.clk(gclk));
	jdff dff_A_LvzGJYUi9_0(.dout(w_dff_A_eIkqh5s40_0),.din(w_dff_A_LvzGJYUi9_0),.clk(gclk));
	jdff dff_A_eIkqh5s40_0(.dout(w_dff_A_JbH58zZu9_0),.din(w_dff_A_eIkqh5s40_0),.clk(gclk));
	jdff dff_A_JbH58zZu9_0(.dout(w_dff_A_kGzAnvD47_0),.din(w_dff_A_JbH58zZu9_0),.clk(gclk));
	jdff dff_A_kGzAnvD47_0(.dout(w_dff_A_jOtCDVt65_0),.din(w_dff_A_kGzAnvD47_0),.clk(gclk));
	jdff dff_A_jOtCDVt65_0(.dout(w_dff_A_utL2w7AN0_0),.din(w_dff_A_jOtCDVt65_0),.clk(gclk));
	jdff dff_A_utL2w7AN0_0(.dout(w_dff_A_m7qFaZLq5_0),.din(w_dff_A_utL2w7AN0_0),.clk(gclk));
	jdff dff_A_m7qFaZLq5_0(.dout(w_dff_A_gVm80JcI8_0),.din(w_dff_A_m7qFaZLq5_0),.clk(gclk));
	jdff dff_A_gVm80JcI8_0(.dout(w_dff_A_aHFy5ff96_0),.din(w_dff_A_gVm80JcI8_0),.clk(gclk));
	jdff dff_A_aHFy5ff96_0(.dout(w_dff_A_DSGeUlm45_0),.din(w_dff_A_aHFy5ff96_0),.clk(gclk));
	jdff dff_A_DSGeUlm45_0(.dout(G634),.din(w_dff_A_DSGeUlm45_0),.clk(gclk));
	jdff dff_A_exStBqkQ5_2(.dout(w_dff_A_wuWBSvkX1_0),.din(w_dff_A_exStBqkQ5_2),.clk(gclk));
	jdff dff_A_wuWBSvkX1_0(.dout(w_dff_A_sWU2c14H7_0),.din(w_dff_A_wuWBSvkX1_0),.clk(gclk));
	jdff dff_A_sWU2c14H7_0(.dout(w_dff_A_ifKrietX1_0),.din(w_dff_A_sWU2c14H7_0),.clk(gclk));
	jdff dff_A_ifKrietX1_0(.dout(w_dff_A_CBMKM7pt5_0),.din(w_dff_A_ifKrietX1_0),.clk(gclk));
	jdff dff_A_CBMKM7pt5_0(.dout(w_dff_A_cKNcyqqd6_0),.din(w_dff_A_CBMKM7pt5_0),.clk(gclk));
	jdff dff_A_cKNcyqqd6_0(.dout(w_dff_A_YzAeThHe1_0),.din(w_dff_A_cKNcyqqd6_0),.clk(gclk));
	jdff dff_A_YzAeThHe1_0(.dout(w_dff_A_XCg6C0rR1_0),.din(w_dff_A_YzAeThHe1_0),.clk(gclk));
	jdff dff_A_XCg6C0rR1_0(.dout(w_dff_A_Y2cdZ01X2_0),.din(w_dff_A_XCg6C0rR1_0),.clk(gclk));
	jdff dff_A_Y2cdZ01X2_0(.dout(w_dff_A_P4Ckavm71_0),.din(w_dff_A_Y2cdZ01X2_0),.clk(gclk));
	jdff dff_A_P4Ckavm71_0(.dout(w_dff_A_IPLI65ef5_0),.din(w_dff_A_P4Ckavm71_0),.clk(gclk));
	jdff dff_A_IPLI65ef5_0(.dout(w_dff_A_abzK3VH78_0),.din(w_dff_A_IPLI65ef5_0),.clk(gclk));
	jdff dff_A_abzK3VH78_0(.dout(w_dff_A_LPDUQsau6_0),.din(w_dff_A_abzK3VH78_0),.clk(gclk));
	jdff dff_A_LPDUQsau6_0(.dout(w_dff_A_0J3DAQz32_0),.din(w_dff_A_LPDUQsau6_0),.clk(gclk));
	jdff dff_A_0J3DAQz32_0(.dout(w_dff_A_3xCap0Mj8_0),.din(w_dff_A_0J3DAQz32_0),.clk(gclk));
	jdff dff_A_3xCap0Mj8_0(.dout(w_dff_A_lBXDLFVS9_0),.din(w_dff_A_3xCap0Mj8_0),.clk(gclk));
	jdff dff_A_lBXDLFVS9_0(.dout(w_dff_A_CQ46U00c2_0),.din(w_dff_A_lBXDLFVS9_0),.clk(gclk));
	jdff dff_A_CQ46U00c2_0(.dout(w_dff_A_Y7L5ftOy9_0),.din(w_dff_A_CQ46U00c2_0),.clk(gclk));
	jdff dff_A_Y7L5ftOy9_0(.dout(w_dff_A_VtWdf7Dz6_0),.din(w_dff_A_Y7L5ftOy9_0),.clk(gclk));
	jdff dff_A_VtWdf7Dz6_0(.dout(w_dff_A_aaYvH3vo7_0),.din(w_dff_A_VtWdf7Dz6_0),.clk(gclk));
	jdff dff_A_aaYvH3vo7_0(.dout(w_dff_A_etZ9ZXnN3_0),.din(w_dff_A_aaYvH3vo7_0),.clk(gclk));
	jdff dff_A_etZ9ZXnN3_0(.dout(w_dff_A_fqB1lQAs3_0),.din(w_dff_A_etZ9ZXnN3_0),.clk(gclk));
	jdff dff_A_fqB1lQAs3_0(.dout(w_dff_A_SF599VBN1_0),.din(w_dff_A_fqB1lQAs3_0),.clk(gclk));
	jdff dff_A_SF599VBN1_0(.dout(w_dff_A_vDBYVT3T9_0),.din(w_dff_A_SF599VBN1_0),.clk(gclk));
	jdff dff_A_vDBYVT3T9_0(.dout(w_dff_A_IXVxdoHg8_0),.din(w_dff_A_vDBYVT3T9_0),.clk(gclk));
	jdff dff_A_IXVxdoHg8_0(.dout(w_dff_A_LER4ChrA4_0),.din(w_dff_A_IXVxdoHg8_0),.clk(gclk));
	jdff dff_A_LER4ChrA4_0(.dout(G815),.din(w_dff_A_LER4ChrA4_0),.clk(gclk));
	jdff dff_A_TqMoaJk03_2(.dout(w_dff_A_wX0tWmqN4_0),.din(w_dff_A_TqMoaJk03_2),.clk(gclk));
	jdff dff_A_wX0tWmqN4_0(.dout(w_dff_A_tax51nS43_0),.din(w_dff_A_wX0tWmqN4_0),.clk(gclk));
	jdff dff_A_tax51nS43_0(.dout(w_dff_A_iHRLFPRF5_0),.din(w_dff_A_tax51nS43_0),.clk(gclk));
	jdff dff_A_iHRLFPRF5_0(.dout(w_dff_A_rOfsVARI3_0),.din(w_dff_A_iHRLFPRF5_0),.clk(gclk));
	jdff dff_A_rOfsVARI3_0(.dout(w_dff_A_xy8qDcDh8_0),.din(w_dff_A_rOfsVARI3_0),.clk(gclk));
	jdff dff_A_xy8qDcDh8_0(.dout(w_dff_A_kwydTDlu0_0),.din(w_dff_A_xy8qDcDh8_0),.clk(gclk));
	jdff dff_A_kwydTDlu0_0(.dout(w_dff_A_KZK8FBHa9_0),.din(w_dff_A_kwydTDlu0_0),.clk(gclk));
	jdff dff_A_KZK8FBHa9_0(.dout(w_dff_A_BKOrgFgS3_0),.din(w_dff_A_KZK8FBHa9_0),.clk(gclk));
	jdff dff_A_BKOrgFgS3_0(.dout(w_dff_A_K8oGeYbo5_0),.din(w_dff_A_BKOrgFgS3_0),.clk(gclk));
	jdff dff_A_K8oGeYbo5_0(.dout(w_dff_A_F0YoVC4q5_0),.din(w_dff_A_K8oGeYbo5_0),.clk(gclk));
	jdff dff_A_F0YoVC4q5_0(.dout(w_dff_A_Eyrjf1Aa7_0),.din(w_dff_A_F0YoVC4q5_0),.clk(gclk));
	jdff dff_A_Eyrjf1Aa7_0(.dout(w_dff_A_dvyRq3G07_0),.din(w_dff_A_Eyrjf1Aa7_0),.clk(gclk));
	jdff dff_A_dvyRq3G07_0(.dout(w_dff_A_CCSbbp4O5_0),.din(w_dff_A_dvyRq3G07_0),.clk(gclk));
	jdff dff_A_CCSbbp4O5_0(.dout(w_dff_A_kpI7ahMl0_0),.din(w_dff_A_CCSbbp4O5_0),.clk(gclk));
	jdff dff_A_kpI7ahMl0_0(.dout(w_dff_A_0f30fpFz1_0),.din(w_dff_A_kpI7ahMl0_0),.clk(gclk));
	jdff dff_A_0f30fpFz1_0(.dout(w_dff_A_Rw0Qhv6R7_0),.din(w_dff_A_0f30fpFz1_0),.clk(gclk));
	jdff dff_A_Rw0Qhv6R7_0(.dout(w_dff_A_8cxXHgb43_0),.din(w_dff_A_Rw0Qhv6R7_0),.clk(gclk));
	jdff dff_A_8cxXHgb43_0(.dout(w_dff_A_GTWRWzMJ1_0),.din(w_dff_A_8cxXHgb43_0),.clk(gclk));
	jdff dff_A_GTWRWzMJ1_0(.dout(w_dff_A_kNfBVaqN5_0),.din(w_dff_A_GTWRWzMJ1_0),.clk(gclk));
	jdff dff_A_kNfBVaqN5_0(.dout(w_dff_A_jYZljm1K3_0),.din(w_dff_A_kNfBVaqN5_0),.clk(gclk));
	jdff dff_A_jYZljm1K3_0(.dout(w_dff_A_tN44kCaU6_0),.din(w_dff_A_jYZljm1K3_0),.clk(gclk));
	jdff dff_A_tN44kCaU6_0(.dout(w_dff_A_7xzm6zBw3_0),.din(w_dff_A_tN44kCaU6_0),.clk(gclk));
	jdff dff_A_7xzm6zBw3_0(.dout(w_dff_A_Y80qzSBW2_0),.din(w_dff_A_7xzm6zBw3_0),.clk(gclk));
	jdff dff_A_Y80qzSBW2_0(.dout(w_dff_A_jTF1pupG7_0),.din(w_dff_A_Y80qzSBW2_0),.clk(gclk));
	jdff dff_A_jTF1pupG7_0(.dout(w_dff_A_9CvpmEld7_0),.din(w_dff_A_jTF1pupG7_0),.clk(gclk));
	jdff dff_A_9CvpmEld7_0(.dout(G845),.din(w_dff_A_9CvpmEld7_0),.clk(gclk));
	jdff dff_A_X7F1HKYL4_1(.dout(w_dff_A_uolmimfa7_0),.din(w_dff_A_X7F1HKYL4_1),.clk(gclk));
	jdff dff_A_uolmimfa7_0(.dout(w_dff_A_N9AqXNZj4_0),.din(w_dff_A_uolmimfa7_0),.clk(gclk));
	jdff dff_A_N9AqXNZj4_0(.dout(w_dff_A_eYsRJPwR2_0),.din(w_dff_A_N9AqXNZj4_0),.clk(gclk));
	jdff dff_A_eYsRJPwR2_0(.dout(w_dff_A_ullLoJye8_0),.din(w_dff_A_eYsRJPwR2_0),.clk(gclk));
	jdff dff_A_ullLoJye8_0(.dout(w_dff_A_W5SJSUET1_0),.din(w_dff_A_ullLoJye8_0),.clk(gclk));
	jdff dff_A_W5SJSUET1_0(.dout(w_dff_A_oN66D3234_0),.din(w_dff_A_W5SJSUET1_0),.clk(gclk));
	jdff dff_A_oN66D3234_0(.dout(w_dff_A_njo6NJt84_0),.din(w_dff_A_oN66D3234_0),.clk(gclk));
	jdff dff_A_njo6NJt84_0(.dout(w_dff_A_TwGOlEDQ3_0),.din(w_dff_A_njo6NJt84_0),.clk(gclk));
	jdff dff_A_TwGOlEDQ3_0(.dout(w_dff_A_05yKt7xE7_0),.din(w_dff_A_TwGOlEDQ3_0),.clk(gclk));
	jdff dff_A_05yKt7xE7_0(.dout(w_dff_A_nWhjeQUn1_0),.din(w_dff_A_05yKt7xE7_0),.clk(gclk));
	jdff dff_A_nWhjeQUn1_0(.dout(w_dff_A_0k5yljyq4_0),.din(w_dff_A_nWhjeQUn1_0),.clk(gclk));
	jdff dff_A_0k5yljyq4_0(.dout(w_dff_A_joeKOMa00_0),.din(w_dff_A_0k5yljyq4_0),.clk(gclk));
	jdff dff_A_joeKOMa00_0(.dout(w_dff_A_1W5ct2YD4_0),.din(w_dff_A_joeKOMa00_0),.clk(gclk));
	jdff dff_A_1W5ct2YD4_0(.dout(w_dff_A_jgrFbjJM0_0),.din(w_dff_A_1W5ct2YD4_0),.clk(gclk));
	jdff dff_A_jgrFbjJM0_0(.dout(w_dff_A_2svmAVov8_0),.din(w_dff_A_jgrFbjJM0_0),.clk(gclk));
	jdff dff_A_2svmAVov8_0(.dout(w_dff_A_fymio6HD2_0),.din(w_dff_A_2svmAVov8_0),.clk(gclk));
	jdff dff_A_fymio6HD2_0(.dout(w_dff_A_2y5WtJwj2_0),.din(w_dff_A_fymio6HD2_0),.clk(gclk));
	jdff dff_A_2y5WtJwj2_0(.dout(w_dff_A_rapHXvm16_0),.din(w_dff_A_2y5WtJwj2_0),.clk(gclk));
	jdff dff_A_rapHXvm16_0(.dout(w_dff_A_UV1gxB2A0_0),.din(w_dff_A_rapHXvm16_0),.clk(gclk));
	jdff dff_A_UV1gxB2A0_0(.dout(w_dff_A_Qb1y4N3U2_0),.din(w_dff_A_UV1gxB2A0_0),.clk(gclk));
	jdff dff_A_Qb1y4N3U2_0(.dout(w_dff_A_yE9pNrb00_0),.din(w_dff_A_Qb1y4N3U2_0),.clk(gclk));
	jdff dff_A_yE9pNrb00_0(.dout(w_dff_A_bC9yovAL8_0),.din(w_dff_A_yE9pNrb00_0),.clk(gclk));
	jdff dff_A_bC9yovAL8_0(.dout(w_dff_A_SRGktNGU7_0),.din(w_dff_A_bC9yovAL8_0),.clk(gclk));
	jdff dff_A_SRGktNGU7_0(.dout(w_dff_A_gGXfGeiv4_0),.din(w_dff_A_SRGktNGU7_0),.clk(gclk));
	jdff dff_A_gGXfGeiv4_0(.dout(w_dff_A_HyNuPhMA7_0),.din(w_dff_A_gGXfGeiv4_0),.clk(gclk));
	jdff dff_A_HyNuPhMA7_0(.dout(G847),.din(w_dff_A_HyNuPhMA7_0),.clk(gclk));
	jdff dff_A_TKuoKSCW6_1(.dout(w_dff_A_kZTx9DQi5_0),.din(w_dff_A_TKuoKSCW6_1),.clk(gclk));
	jdff dff_A_kZTx9DQi5_0(.dout(w_dff_A_XAMLZK897_0),.din(w_dff_A_kZTx9DQi5_0),.clk(gclk));
	jdff dff_A_XAMLZK897_0(.dout(w_dff_A_Q0KDuIQD5_0),.din(w_dff_A_XAMLZK897_0),.clk(gclk));
	jdff dff_A_Q0KDuIQD5_0(.dout(w_dff_A_7HskTq8i1_0),.din(w_dff_A_Q0KDuIQD5_0),.clk(gclk));
	jdff dff_A_7HskTq8i1_0(.dout(w_dff_A_p0dUaPYs2_0),.din(w_dff_A_7HskTq8i1_0),.clk(gclk));
	jdff dff_A_p0dUaPYs2_0(.dout(w_dff_A_dPB2mbSR9_0),.din(w_dff_A_p0dUaPYs2_0),.clk(gclk));
	jdff dff_A_dPB2mbSR9_0(.dout(w_dff_A_6DoRZaxf7_0),.din(w_dff_A_dPB2mbSR9_0),.clk(gclk));
	jdff dff_A_6DoRZaxf7_0(.dout(w_dff_A_KtB1YAE87_0),.din(w_dff_A_6DoRZaxf7_0),.clk(gclk));
	jdff dff_A_KtB1YAE87_0(.dout(w_dff_A_8r1zBTMk4_0),.din(w_dff_A_KtB1YAE87_0),.clk(gclk));
	jdff dff_A_8r1zBTMk4_0(.dout(w_dff_A_ZvjI8cll1_0),.din(w_dff_A_8r1zBTMk4_0),.clk(gclk));
	jdff dff_A_ZvjI8cll1_0(.dout(w_dff_A_V4Vrc5Gq4_0),.din(w_dff_A_ZvjI8cll1_0),.clk(gclk));
	jdff dff_A_V4Vrc5Gq4_0(.dout(w_dff_A_oZ86eTmZ4_0),.din(w_dff_A_V4Vrc5Gq4_0),.clk(gclk));
	jdff dff_A_oZ86eTmZ4_0(.dout(w_dff_A_lCenTC5v2_0),.din(w_dff_A_oZ86eTmZ4_0),.clk(gclk));
	jdff dff_A_lCenTC5v2_0(.dout(w_dff_A_m0rGnH2a3_0),.din(w_dff_A_lCenTC5v2_0),.clk(gclk));
	jdff dff_A_m0rGnH2a3_0(.dout(w_dff_A_ZuHOqMvl8_0),.din(w_dff_A_m0rGnH2a3_0),.clk(gclk));
	jdff dff_A_ZuHOqMvl8_0(.dout(w_dff_A_PaIkXcRc8_0),.din(w_dff_A_ZuHOqMvl8_0),.clk(gclk));
	jdff dff_A_PaIkXcRc8_0(.dout(w_dff_A_XiLAzX2v0_0),.din(w_dff_A_PaIkXcRc8_0),.clk(gclk));
	jdff dff_A_XiLAzX2v0_0(.dout(w_dff_A_W3C6j8an3_0),.din(w_dff_A_XiLAzX2v0_0),.clk(gclk));
	jdff dff_A_W3C6j8an3_0(.dout(w_dff_A_oTAmvKeV6_0),.din(w_dff_A_W3C6j8an3_0),.clk(gclk));
	jdff dff_A_oTAmvKeV6_0(.dout(w_dff_A_Fdx07G1M3_0),.din(w_dff_A_oTAmvKeV6_0),.clk(gclk));
	jdff dff_A_Fdx07G1M3_0(.dout(w_dff_A_pP7Lof4f8_0),.din(w_dff_A_Fdx07G1M3_0),.clk(gclk));
	jdff dff_A_pP7Lof4f8_0(.dout(w_dff_A_TUK6L97F4_0),.din(w_dff_A_pP7Lof4f8_0),.clk(gclk));
	jdff dff_A_TUK6L97F4_0(.dout(w_dff_A_1oJ631Nj6_0),.din(w_dff_A_TUK6L97F4_0),.clk(gclk));
	jdff dff_A_1oJ631Nj6_0(.dout(w_dff_A_UBYY5Txl7_0),.din(w_dff_A_1oJ631Nj6_0),.clk(gclk));
	jdff dff_A_UBYY5Txl7_0(.dout(w_dff_A_KoPsLqfG6_0),.din(w_dff_A_UBYY5Txl7_0),.clk(gclk));
	jdff dff_A_KoPsLqfG6_0(.dout(w_dff_A_nl539tiC9_0),.din(w_dff_A_KoPsLqfG6_0),.clk(gclk));
	jdff dff_A_nl539tiC9_0(.dout(w_dff_A_lxqjMQZT1_0),.din(w_dff_A_nl539tiC9_0),.clk(gclk));
	jdff dff_A_lxqjMQZT1_0(.dout(G926),.din(w_dff_A_lxqjMQZT1_0),.clk(gclk));
	jdff dff_A_K6wpGJWd3_1(.dout(w_dff_A_svZrmNcT1_0),.din(w_dff_A_K6wpGJWd3_1),.clk(gclk));
	jdff dff_A_svZrmNcT1_0(.dout(w_dff_A_9glUybEI4_0),.din(w_dff_A_svZrmNcT1_0),.clk(gclk));
	jdff dff_A_9glUybEI4_0(.dout(w_dff_A_YCiEjFmB0_0),.din(w_dff_A_9glUybEI4_0),.clk(gclk));
	jdff dff_A_YCiEjFmB0_0(.dout(w_dff_A_x8QmaDmv5_0),.din(w_dff_A_YCiEjFmB0_0),.clk(gclk));
	jdff dff_A_x8QmaDmv5_0(.dout(w_dff_A_h1tcUOTL7_0),.din(w_dff_A_x8QmaDmv5_0),.clk(gclk));
	jdff dff_A_h1tcUOTL7_0(.dout(w_dff_A_kdTQgwsB1_0),.din(w_dff_A_h1tcUOTL7_0),.clk(gclk));
	jdff dff_A_kdTQgwsB1_0(.dout(w_dff_A_DRN1mrgV8_0),.din(w_dff_A_kdTQgwsB1_0),.clk(gclk));
	jdff dff_A_DRN1mrgV8_0(.dout(w_dff_A_nmj3gwya5_0),.din(w_dff_A_DRN1mrgV8_0),.clk(gclk));
	jdff dff_A_nmj3gwya5_0(.dout(w_dff_A_VGMn8EBD2_0),.din(w_dff_A_nmj3gwya5_0),.clk(gclk));
	jdff dff_A_VGMn8EBD2_0(.dout(w_dff_A_4vSHMUWt7_0),.din(w_dff_A_VGMn8EBD2_0),.clk(gclk));
	jdff dff_A_4vSHMUWt7_0(.dout(w_dff_A_ZVqvWqnY1_0),.din(w_dff_A_4vSHMUWt7_0),.clk(gclk));
	jdff dff_A_ZVqvWqnY1_0(.dout(w_dff_A_AizFZySo8_0),.din(w_dff_A_ZVqvWqnY1_0),.clk(gclk));
	jdff dff_A_AizFZySo8_0(.dout(w_dff_A_qRzsO6K48_0),.din(w_dff_A_AizFZySo8_0),.clk(gclk));
	jdff dff_A_qRzsO6K48_0(.dout(w_dff_A_84LrDuoC8_0),.din(w_dff_A_qRzsO6K48_0),.clk(gclk));
	jdff dff_A_84LrDuoC8_0(.dout(w_dff_A_pcbL62Am2_0),.din(w_dff_A_84LrDuoC8_0),.clk(gclk));
	jdff dff_A_pcbL62Am2_0(.dout(w_dff_A_3Z9WgCgd0_0),.din(w_dff_A_pcbL62Am2_0),.clk(gclk));
	jdff dff_A_3Z9WgCgd0_0(.dout(w_dff_A_BYPa2LIP9_0),.din(w_dff_A_3Z9WgCgd0_0),.clk(gclk));
	jdff dff_A_BYPa2LIP9_0(.dout(w_dff_A_kmWpum7a4_0),.din(w_dff_A_BYPa2LIP9_0),.clk(gclk));
	jdff dff_A_kmWpum7a4_0(.dout(w_dff_A_HnPGqevu0_0),.din(w_dff_A_kmWpum7a4_0),.clk(gclk));
	jdff dff_A_HnPGqevu0_0(.dout(w_dff_A_bdGU1SC37_0),.din(w_dff_A_HnPGqevu0_0),.clk(gclk));
	jdff dff_A_bdGU1SC37_0(.dout(w_dff_A_tjOBBkxe5_0),.din(w_dff_A_bdGU1SC37_0),.clk(gclk));
	jdff dff_A_tjOBBkxe5_0(.dout(w_dff_A_iloMe4C68_0),.din(w_dff_A_tjOBBkxe5_0),.clk(gclk));
	jdff dff_A_iloMe4C68_0(.dout(w_dff_A_8iAIhAUm1_0),.din(w_dff_A_iloMe4C68_0),.clk(gclk));
	jdff dff_A_8iAIhAUm1_0(.dout(w_dff_A_veLfxbv81_0),.din(w_dff_A_8iAIhAUm1_0),.clk(gclk));
	jdff dff_A_veLfxbv81_0(.dout(w_dff_A_5BeclRPt5_0),.din(w_dff_A_veLfxbv81_0),.clk(gclk));
	jdff dff_A_5BeclRPt5_0(.dout(w_dff_A_rldhZ6m63_0),.din(w_dff_A_5BeclRPt5_0),.clk(gclk));
	jdff dff_A_rldhZ6m63_0(.dout(w_dff_A_5F3MKZkd9_0),.din(w_dff_A_rldhZ6m63_0),.clk(gclk));
	jdff dff_A_5F3MKZkd9_0(.dout(G923),.din(w_dff_A_5F3MKZkd9_0),.clk(gclk));
	jdff dff_A_7l1xJPxg8_1(.dout(w_dff_A_3BtInpLT1_0),.din(w_dff_A_7l1xJPxg8_1),.clk(gclk));
	jdff dff_A_3BtInpLT1_0(.dout(w_dff_A_Dxpbdw9F3_0),.din(w_dff_A_3BtInpLT1_0),.clk(gclk));
	jdff dff_A_Dxpbdw9F3_0(.dout(w_dff_A_BSbxc1X46_0),.din(w_dff_A_Dxpbdw9F3_0),.clk(gclk));
	jdff dff_A_BSbxc1X46_0(.dout(w_dff_A_J6W2mOVq3_0),.din(w_dff_A_BSbxc1X46_0),.clk(gclk));
	jdff dff_A_J6W2mOVq3_0(.dout(w_dff_A_x0c4WEPB3_0),.din(w_dff_A_J6W2mOVq3_0),.clk(gclk));
	jdff dff_A_x0c4WEPB3_0(.dout(w_dff_A_Btim2EmK9_0),.din(w_dff_A_x0c4WEPB3_0),.clk(gclk));
	jdff dff_A_Btim2EmK9_0(.dout(w_dff_A_Rm9xGRml6_0),.din(w_dff_A_Btim2EmK9_0),.clk(gclk));
	jdff dff_A_Rm9xGRml6_0(.dout(w_dff_A_3KwY0D8P4_0),.din(w_dff_A_Rm9xGRml6_0),.clk(gclk));
	jdff dff_A_3KwY0D8P4_0(.dout(w_dff_A_Bj9mIC140_0),.din(w_dff_A_3KwY0D8P4_0),.clk(gclk));
	jdff dff_A_Bj9mIC140_0(.dout(w_dff_A_A8tdTRLX4_0),.din(w_dff_A_Bj9mIC140_0),.clk(gclk));
	jdff dff_A_A8tdTRLX4_0(.dout(w_dff_A_l0UNyCUa6_0),.din(w_dff_A_A8tdTRLX4_0),.clk(gclk));
	jdff dff_A_l0UNyCUa6_0(.dout(w_dff_A_VP4EwxVk1_0),.din(w_dff_A_l0UNyCUa6_0),.clk(gclk));
	jdff dff_A_VP4EwxVk1_0(.dout(w_dff_A_di23gKqp9_0),.din(w_dff_A_VP4EwxVk1_0),.clk(gclk));
	jdff dff_A_di23gKqp9_0(.dout(w_dff_A_y8tQFYT21_0),.din(w_dff_A_di23gKqp9_0),.clk(gclk));
	jdff dff_A_y8tQFYT21_0(.dout(w_dff_A_LvUPQXoD7_0),.din(w_dff_A_y8tQFYT21_0),.clk(gclk));
	jdff dff_A_LvUPQXoD7_0(.dout(w_dff_A_ZqL753SO0_0),.din(w_dff_A_LvUPQXoD7_0),.clk(gclk));
	jdff dff_A_ZqL753SO0_0(.dout(w_dff_A_0ekW3pl70_0),.din(w_dff_A_ZqL753SO0_0),.clk(gclk));
	jdff dff_A_0ekW3pl70_0(.dout(w_dff_A_u4EQxJVr5_0),.din(w_dff_A_0ekW3pl70_0),.clk(gclk));
	jdff dff_A_u4EQxJVr5_0(.dout(w_dff_A_C7UhureO5_0),.din(w_dff_A_u4EQxJVr5_0),.clk(gclk));
	jdff dff_A_C7UhureO5_0(.dout(w_dff_A_6yTXDHJQ2_0),.din(w_dff_A_C7UhureO5_0),.clk(gclk));
	jdff dff_A_6yTXDHJQ2_0(.dout(w_dff_A_8uEaIVUC2_0),.din(w_dff_A_6yTXDHJQ2_0),.clk(gclk));
	jdff dff_A_8uEaIVUC2_0(.dout(w_dff_A_3grzfB785_0),.din(w_dff_A_8uEaIVUC2_0),.clk(gclk));
	jdff dff_A_3grzfB785_0(.dout(w_dff_A_UQLSSYID3_0),.din(w_dff_A_3grzfB785_0),.clk(gclk));
	jdff dff_A_UQLSSYID3_0(.dout(w_dff_A_qP045btj2_0),.din(w_dff_A_UQLSSYID3_0),.clk(gclk));
	jdff dff_A_qP045btj2_0(.dout(w_dff_A_NGwoo8C80_0),.din(w_dff_A_qP045btj2_0),.clk(gclk));
	jdff dff_A_NGwoo8C80_0(.dout(w_dff_A_MskSZxQV0_0),.din(w_dff_A_NGwoo8C80_0),.clk(gclk));
	jdff dff_A_MskSZxQV0_0(.dout(w_dff_A_7fWrvqMH1_0),.din(w_dff_A_MskSZxQV0_0),.clk(gclk));
	jdff dff_A_7fWrvqMH1_0(.dout(G921),.din(w_dff_A_7fWrvqMH1_0),.clk(gclk));
	jdff dff_A_2dIO24Jj4_1(.dout(w_dff_A_JZFRN4bg2_0),.din(w_dff_A_2dIO24Jj4_1),.clk(gclk));
	jdff dff_A_JZFRN4bg2_0(.dout(w_dff_A_hBEiWT7E1_0),.din(w_dff_A_JZFRN4bg2_0),.clk(gclk));
	jdff dff_A_hBEiWT7E1_0(.dout(w_dff_A_05KovSCo7_0),.din(w_dff_A_hBEiWT7E1_0),.clk(gclk));
	jdff dff_A_05KovSCo7_0(.dout(w_dff_A_C4E5evo04_0),.din(w_dff_A_05KovSCo7_0),.clk(gclk));
	jdff dff_A_C4E5evo04_0(.dout(w_dff_A_TuXHF67f6_0),.din(w_dff_A_C4E5evo04_0),.clk(gclk));
	jdff dff_A_TuXHF67f6_0(.dout(w_dff_A_jmsVYBMe5_0),.din(w_dff_A_TuXHF67f6_0),.clk(gclk));
	jdff dff_A_jmsVYBMe5_0(.dout(w_dff_A_WkZyNZYE1_0),.din(w_dff_A_jmsVYBMe5_0),.clk(gclk));
	jdff dff_A_WkZyNZYE1_0(.dout(w_dff_A_GKzmejjr5_0),.din(w_dff_A_WkZyNZYE1_0),.clk(gclk));
	jdff dff_A_GKzmejjr5_0(.dout(w_dff_A_3yjqPXRu3_0),.din(w_dff_A_GKzmejjr5_0),.clk(gclk));
	jdff dff_A_3yjqPXRu3_0(.dout(w_dff_A_wa3LCTQR6_0),.din(w_dff_A_3yjqPXRu3_0),.clk(gclk));
	jdff dff_A_wa3LCTQR6_0(.dout(w_dff_A_Op8uBwhR6_0),.din(w_dff_A_wa3LCTQR6_0),.clk(gclk));
	jdff dff_A_Op8uBwhR6_0(.dout(w_dff_A_b3ZWdLmK3_0),.din(w_dff_A_Op8uBwhR6_0),.clk(gclk));
	jdff dff_A_b3ZWdLmK3_0(.dout(w_dff_A_y1CmGoI21_0),.din(w_dff_A_b3ZWdLmK3_0),.clk(gclk));
	jdff dff_A_y1CmGoI21_0(.dout(w_dff_A_XN3l33IS4_0),.din(w_dff_A_y1CmGoI21_0),.clk(gclk));
	jdff dff_A_XN3l33IS4_0(.dout(w_dff_A_trz5VlK68_0),.din(w_dff_A_XN3l33IS4_0),.clk(gclk));
	jdff dff_A_trz5VlK68_0(.dout(w_dff_A_n7EYXIdz7_0),.din(w_dff_A_trz5VlK68_0),.clk(gclk));
	jdff dff_A_n7EYXIdz7_0(.dout(w_dff_A_9QOtFYE66_0),.din(w_dff_A_n7EYXIdz7_0),.clk(gclk));
	jdff dff_A_9QOtFYE66_0(.dout(w_dff_A_L7AYeuKv3_0),.din(w_dff_A_9QOtFYE66_0),.clk(gclk));
	jdff dff_A_L7AYeuKv3_0(.dout(w_dff_A_RBeo2VRm9_0),.din(w_dff_A_L7AYeuKv3_0),.clk(gclk));
	jdff dff_A_RBeo2VRm9_0(.dout(w_dff_A_J3hIDXpq7_0),.din(w_dff_A_RBeo2VRm9_0),.clk(gclk));
	jdff dff_A_J3hIDXpq7_0(.dout(w_dff_A_i7wMwufA7_0),.din(w_dff_A_J3hIDXpq7_0),.clk(gclk));
	jdff dff_A_i7wMwufA7_0(.dout(w_dff_A_xPbSj6o89_0),.din(w_dff_A_i7wMwufA7_0),.clk(gclk));
	jdff dff_A_xPbSj6o89_0(.dout(w_dff_A_QmYk2Xnp1_0),.din(w_dff_A_xPbSj6o89_0),.clk(gclk));
	jdff dff_A_QmYk2Xnp1_0(.dout(w_dff_A_nGDtdNpn7_0),.din(w_dff_A_QmYk2Xnp1_0),.clk(gclk));
	jdff dff_A_nGDtdNpn7_0(.dout(w_dff_A_BvFAkxhV2_0),.din(w_dff_A_nGDtdNpn7_0),.clk(gclk));
	jdff dff_A_BvFAkxhV2_0(.dout(w_dff_A_1jMbOY4l0_0),.din(w_dff_A_BvFAkxhV2_0),.clk(gclk));
	jdff dff_A_1jMbOY4l0_0(.dout(w_dff_A_H6KQgU2i4_0),.din(w_dff_A_1jMbOY4l0_0),.clk(gclk));
	jdff dff_A_H6KQgU2i4_0(.dout(G892),.din(w_dff_A_H6KQgU2i4_0),.clk(gclk));
	jdff dff_A_lRm1ZvdP4_1(.dout(w_dff_A_fidZ2kb52_0),.din(w_dff_A_lRm1ZvdP4_1),.clk(gclk));
	jdff dff_A_fidZ2kb52_0(.dout(w_dff_A_kInfo4lD6_0),.din(w_dff_A_fidZ2kb52_0),.clk(gclk));
	jdff dff_A_kInfo4lD6_0(.dout(w_dff_A_KMjoz2Vx1_0),.din(w_dff_A_kInfo4lD6_0),.clk(gclk));
	jdff dff_A_KMjoz2Vx1_0(.dout(w_dff_A_JmxLcGv83_0),.din(w_dff_A_KMjoz2Vx1_0),.clk(gclk));
	jdff dff_A_JmxLcGv83_0(.dout(w_dff_A_ui9jUVXr9_0),.din(w_dff_A_JmxLcGv83_0),.clk(gclk));
	jdff dff_A_ui9jUVXr9_0(.dout(w_dff_A_DN2FgIAM8_0),.din(w_dff_A_ui9jUVXr9_0),.clk(gclk));
	jdff dff_A_DN2FgIAM8_0(.dout(w_dff_A_RZdDCcOz3_0),.din(w_dff_A_DN2FgIAM8_0),.clk(gclk));
	jdff dff_A_RZdDCcOz3_0(.dout(w_dff_A_hbdCbXy21_0),.din(w_dff_A_RZdDCcOz3_0),.clk(gclk));
	jdff dff_A_hbdCbXy21_0(.dout(w_dff_A_M8Z17VPj6_0),.din(w_dff_A_hbdCbXy21_0),.clk(gclk));
	jdff dff_A_M8Z17VPj6_0(.dout(w_dff_A_SYOPsecX8_0),.din(w_dff_A_M8Z17VPj6_0),.clk(gclk));
	jdff dff_A_SYOPsecX8_0(.dout(w_dff_A_XKu1PCda4_0),.din(w_dff_A_SYOPsecX8_0),.clk(gclk));
	jdff dff_A_XKu1PCda4_0(.dout(w_dff_A_8OmycR1V2_0),.din(w_dff_A_XKu1PCda4_0),.clk(gclk));
	jdff dff_A_8OmycR1V2_0(.dout(w_dff_A_TxCas6dB8_0),.din(w_dff_A_8OmycR1V2_0),.clk(gclk));
	jdff dff_A_TxCas6dB8_0(.dout(w_dff_A_N0gzojVw9_0),.din(w_dff_A_TxCas6dB8_0),.clk(gclk));
	jdff dff_A_N0gzojVw9_0(.dout(w_dff_A_kh8NhTMo8_0),.din(w_dff_A_N0gzojVw9_0),.clk(gclk));
	jdff dff_A_kh8NhTMo8_0(.dout(w_dff_A_rwR7Xe3H1_0),.din(w_dff_A_kh8NhTMo8_0),.clk(gclk));
	jdff dff_A_rwR7Xe3H1_0(.dout(w_dff_A_yI90uVPX5_0),.din(w_dff_A_rwR7Xe3H1_0),.clk(gclk));
	jdff dff_A_yI90uVPX5_0(.dout(w_dff_A_b6jvVOdI6_0),.din(w_dff_A_yI90uVPX5_0),.clk(gclk));
	jdff dff_A_b6jvVOdI6_0(.dout(w_dff_A_dhe6uz7V4_0),.din(w_dff_A_b6jvVOdI6_0),.clk(gclk));
	jdff dff_A_dhe6uz7V4_0(.dout(w_dff_A_H3gmHbEy4_0),.din(w_dff_A_dhe6uz7V4_0),.clk(gclk));
	jdff dff_A_H3gmHbEy4_0(.dout(w_dff_A_yMtsPDPo7_0),.din(w_dff_A_H3gmHbEy4_0),.clk(gclk));
	jdff dff_A_yMtsPDPo7_0(.dout(w_dff_A_DoxEIe4l3_0),.din(w_dff_A_yMtsPDPo7_0),.clk(gclk));
	jdff dff_A_DoxEIe4l3_0(.dout(w_dff_A_yxT7KSTO6_0),.din(w_dff_A_DoxEIe4l3_0),.clk(gclk));
	jdff dff_A_yxT7KSTO6_0(.dout(w_dff_A_0fe5NYxD3_0),.din(w_dff_A_yxT7KSTO6_0),.clk(gclk));
	jdff dff_A_0fe5NYxD3_0(.dout(w_dff_A_zdwmYmkE7_0),.din(w_dff_A_0fe5NYxD3_0),.clk(gclk));
	jdff dff_A_zdwmYmkE7_0(.dout(w_dff_A_SsdBe5ct7_0),.din(w_dff_A_zdwmYmkE7_0),.clk(gclk));
	jdff dff_A_SsdBe5ct7_0(.dout(w_dff_A_jKZjYG0l5_0),.din(w_dff_A_SsdBe5ct7_0),.clk(gclk));
	jdff dff_A_jKZjYG0l5_0(.dout(G887),.din(w_dff_A_jKZjYG0l5_0),.clk(gclk));
	jdff dff_A_VRuQeKNr1_1(.dout(w_dff_A_9dRG4BhY4_0),.din(w_dff_A_VRuQeKNr1_1),.clk(gclk));
	jdff dff_A_9dRG4BhY4_0(.dout(w_dff_A_kCDmO6Y39_0),.din(w_dff_A_9dRG4BhY4_0),.clk(gclk));
	jdff dff_A_kCDmO6Y39_0(.dout(w_dff_A_iq4yiSHG1_0),.din(w_dff_A_kCDmO6Y39_0),.clk(gclk));
	jdff dff_A_iq4yiSHG1_0(.dout(w_dff_A_pd17vWUi1_0),.din(w_dff_A_iq4yiSHG1_0),.clk(gclk));
	jdff dff_A_pd17vWUi1_0(.dout(w_dff_A_rLhQvUlX8_0),.din(w_dff_A_pd17vWUi1_0),.clk(gclk));
	jdff dff_A_rLhQvUlX8_0(.dout(w_dff_A_d4qsAZCa0_0),.din(w_dff_A_rLhQvUlX8_0),.clk(gclk));
	jdff dff_A_d4qsAZCa0_0(.dout(w_dff_A_oP7jJvD27_0),.din(w_dff_A_d4qsAZCa0_0),.clk(gclk));
	jdff dff_A_oP7jJvD27_0(.dout(w_dff_A_J5JPQTd18_0),.din(w_dff_A_oP7jJvD27_0),.clk(gclk));
	jdff dff_A_J5JPQTd18_0(.dout(w_dff_A_Z0qnVw5v6_0),.din(w_dff_A_J5JPQTd18_0),.clk(gclk));
	jdff dff_A_Z0qnVw5v6_0(.dout(w_dff_A_HeVKRGNY5_0),.din(w_dff_A_Z0qnVw5v6_0),.clk(gclk));
	jdff dff_A_HeVKRGNY5_0(.dout(w_dff_A_jLrRvOig5_0),.din(w_dff_A_HeVKRGNY5_0),.clk(gclk));
	jdff dff_A_jLrRvOig5_0(.dout(w_dff_A_0yv65RKl1_0),.din(w_dff_A_jLrRvOig5_0),.clk(gclk));
	jdff dff_A_0yv65RKl1_0(.dout(w_dff_A_vflgsjhW7_0),.din(w_dff_A_0yv65RKl1_0),.clk(gclk));
	jdff dff_A_vflgsjhW7_0(.dout(w_dff_A_sP3kGwxG9_0),.din(w_dff_A_vflgsjhW7_0),.clk(gclk));
	jdff dff_A_sP3kGwxG9_0(.dout(w_dff_A_CR8lprwe6_0),.din(w_dff_A_sP3kGwxG9_0),.clk(gclk));
	jdff dff_A_CR8lprwe6_0(.dout(w_dff_A_fYFJzdR15_0),.din(w_dff_A_CR8lprwe6_0),.clk(gclk));
	jdff dff_A_fYFJzdR15_0(.dout(w_dff_A_OZ7OF0x22_0),.din(w_dff_A_fYFJzdR15_0),.clk(gclk));
	jdff dff_A_OZ7OF0x22_0(.dout(w_dff_A_ic9h4GPH4_0),.din(w_dff_A_OZ7OF0x22_0),.clk(gclk));
	jdff dff_A_ic9h4GPH4_0(.dout(w_dff_A_dmeUYhbd6_0),.din(w_dff_A_ic9h4GPH4_0),.clk(gclk));
	jdff dff_A_dmeUYhbd6_0(.dout(w_dff_A_ZTWK0T7B8_0),.din(w_dff_A_dmeUYhbd6_0),.clk(gclk));
	jdff dff_A_ZTWK0T7B8_0(.dout(w_dff_A_DKGHJwYl9_0),.din(w_dff_A_ZTWK0T7B8_0),.clk(gclk));
	jdff dff_A_DKGHJwYl9_0(.dout(w_dff_A_xEoJ4PH74_0),.din(w_dff_A_DKGHJwYl9_0),.clk(gclk));
	jdff dff_A_xEoJ4PH74_0(.dout(w_dff_A_7xLa8arg7_0),.din(w_dff_A_xEoJ4PH74_0),.clk(gclk));
	jdff dff_A_7xLa8arg7_0(.dout(w_dff_A_cuiR6SJb7_0),.din(w_dff_A_7xLa8arg7_0),.clk(gclk));
	jdff dff_A_cuiR6SJb7_0(.dout(w_dff_A_w7kXvGwR3_0),.din(w_dff_A_cuiR6SJb7_0),.clk(gclk));
	jdff dff_A_w7kXvGwR3_0(.dout(w_dff_A_FWpDfBEp2_0),.din(w_dff_A_w7kXvGwR3_0),.clk(gclk));
	jdff dff_A_FWpDfBEp2_0(.dout(G606),.din(w_dff_A_FWpDfBEp2_0),.clk(gclk));
	jdff dff_A_gg3PgASV0_2(.dout(w_dff_A_aR4I8e2K2_0),.din(w_dff_A_gg3PgASV0_2),.clk(gclk));
	jdff dff_A_aR4I8e2K2_0(.dout(w_dff_A_Ie7QgcyS2_0),.din(w_dff_A_aR4I8e2K2_0),.clk(gclk));
	jdff dff_A_Ie7QgcyS2_0(.dout(w_dff_A_CRtd59Gh5_0),.din(w_dff_A_Ie7QgcyS2_0),.clk(gclk));
	jdff dff_A_CRtd59Gh5_0(.dout(w_dff_A_8nY0sgGo7_0),.din(w_dff_A_CRtd59Gh5_0),.clk(gclk));
	jdff dff_A_8nY0sgGo7_0(.dout(w_dff_A_AfSjFJ1y3_0),.din(w_dff_A_8nY0sgGo7_0),.clk(gclk));
	jdff dff_A_AfSjFJ1y3_0(.dout(w_dff_A_b1p62XoN6_0),.din(w_dff_A_AfSjFJ1y3_0),.clk(gclk));
	jdff dff_A_b1p62XoN6_0(.dout(w_dff_A_0t3v89To7_0),.din(w_dff_A_b1p62XoN6_0),.clk(gclk));
	jdff dff_A_0t3v89To7_0(.dout(w_dff_A_aWMnwsv82_0),.din(w_dff_A_0t3v89To7_0),.clk(gclk));
	jdff dff_A_aWMnwsv82_0(.dout(w_dff_A_IPp4htNW4_0),.din(w_dff_A_aWMnwsv82_0),.clk(gclk));
	jdff dff_A_IPp4htNW4_0(.dout(w_dff_A_ayhWAWw79_0),.din(w_dff_A_IPp4htNW4_0),.clk(gclk));
	jdff dff_A_ayhWAWw79_0(.dout(w_dff_A_iFtYWRGX8_0),.din(w_dff_A_ayhWAWw79_0),.clk(gclk));
	jdff dff_A_iFtYWRGX8_0(.dout(w_dff_A_nfQuiThr9_0),.din(w_dff_A_iFtYWRGX8_0),.clk(gclk));
	jdff dff_A_nfQuiThr9_0(.dout(w_dff_A_r03sexoY6_0),.din(w_dff_A_nfQuiThr9_0),.clk(gclk));
	jdff dff_A_r03sexoY6_0(.dout(w_dff_A_pkSq7Xgv3_0),.din(w_dff_A_r03sexoY6_0),.clk(gclk));
	jdff dff_A_pkSq7Xgv3_0(.dout(w_dff_A_9Va8nnXD6_0),.din(w_dff_A_pkSq7Xgv3_0),.clk(gclk));
	jdff dff_A_9Va8nnXD6_0(.dout(w_dff_A_MdlN1K6W7_0),.din(w_dff_A_9Va8nnXD6_0),.clk(gclk));
	jdff dff_A_MdlN1K6W7_0(.dout(w_dff_A_27y9WcvV6_0),.din(w_dff_A_MdlN1K6W7_0),.clk(gclk));
	jdff dff_A_27y9WcvV6_0(.dout(w_dff_A_Im5N1SSr6_0),.din(w_dff_A_27y9WcvV6_0),.clk(gclk));
	jdff dff_A_Im5N1SSr6_0(.dout(w_dff_A_1Rp6iL4m3_0),.din(w_dff_A_Im5N1SSr6_0),.clk(gclk));
	jdff dff_A_1Rp6iL4m3_0(.dout(w_dff_A_iYkgZ1bF0_0),.din(w_dff_A_1Rp6iL4m3_0),.clk(gclk));
	jdff dff_A_iYkgZ1bF0_0(.dout(w_dff_A_ZNMqHimi9_0),.din(w_dff_A_iYkgZ1bF0_0),.clk(gclk));
	jdff dff_A_ZNMqHimi9_0(.dout(w_dff_A_RHpnLfV68_0),.din(w_dff_A_ZNMqHimi9_0),.clk(gclk));
	jdff dff_A_RHpnLfV68_0(.dout(w_dff_A_uPLTWHaV8_0),.din(w_dff_A_RHpnLfV68_0),.clk(gclk));
	jdff dff_A_uPLTWHaV8_0(.dout(w_dff_A_5Eeh20Wr7_0),.din(w_dff_A_uPLTWHaV8_0),.clk(gclk));
	jdff dff_A_5Eeh20Wr7_0(.dout(G656),.din(w_dff_A_5Eeh20Wr7_0),.clk(gclk));
	jdff dff_A_yuNhCNJz3_2(.dout(w_dff_A_WvrD45bc8_0),.din(w_dff_A_yuNhCNJz3_2),.clk(gclk));
	jdff dff_A_WvrD45bc8_0(.dout(w_dff_A_5H6WQno93_0),.din(w_dff_A_WvrD45bc8_0),.clk(gclk));
	jdff dff_A_5H6WQno93_0(.dout(w_dff_A_ivQAUMxH8_0),.din(w_dff_A_5H6WQno93_0),.clk(gclk));
	jdff dff_A_ivQAUMxH8_0(.dout(w_dff_A_bQjt1a1G0_0),.din(w_dff_A_ivQAUMxH8_0),.clk(gclk));
	jdff dff_A_bQjt1a1G0_0(.dout(w_dff_A_GSt8cXHT4_0),.din(w_dff_A_bQjt1a1G0_0),.clk(gclk));
	jdff dff_A_GSt8cXHT4_0(.dout(w_dff_A_uMkgMiZf3_0),.din(w_dff_A_GSt8cXHT4_0),.clk(gclk));
	jdff dff_A_uMkgMiZf3_0(.dout(w_dff_A_MzDnONN47_0),.din(w_dff_A_uMkgMiZf3_0),.clk(gclk));
	jdff dff_A_MzDnONN47_0(.dout(w_dff_A_a6Pot5A36_0),.din(w_dff_A_MzDnONN47_0),.clk(gclk));
	jdff dff_A_a6Pot5A36_0(.dout(w_dff_A_KAZbcTXc0_0),.din(w_dff_A_a6Pot5A36_0),.clk(gclk));
	jdff dff_A_KAZbcTXc0_0(.dout(w_dff_A_5MWOhsnT4_0),.din(w_dff_A_KAZbcTXc0_0),.clk(gclk));
	jdff dff_A_5MWOhsnT4_0(.dout(w_dff_A_so1wG80E3_0),.din(w_dff_A_5MWOhsnT4_0),.clk(gclk));
	jdff dff_A_so1wG80E3_0(.dout(w_dff_A_47Tc0aO99_0),.din(w_dff_A_so1wG80E3_0),.clk(gclk));
	jdff dff_A_47Tc0aO99_0(.dout(w_dff_A_DiPs3LSX3_0),.din(w_dff_A_47Tc0aO99_0),.clk(gclk));
	jdff dff_A_DiPs3LSX3_0(.dout(w_dff_A_fzQQPQQr6_0),.din(w_dff_A_DiPs3LSX3_0),.clk(gclk));
	jdff dff_A_fzQQPQQr6_0(.dout(w_dff_A_NbxfKrOW2_0),.din(w_dff_A_fzQQPQQr6_0),.clk(gclk));
	jdff dff_A_NbxfKrOW2_0(.dout(w_dff_A_gB4h6JBI1_0),.din(w_dff_A_NbxfKrOW2_0),.clk(gclk));
	jdff dff_A_gB4h6JBI1_0(.dout(w_dff_A_cEwu8iz73_0),.din(w_dff_A_gB4h6JBI1_0),.clk(gclk));
	jdff dff_A_cEwu8iz73_0(.dout(w_dff_A_L7zAtZmE4_0),.din(w_dff_A_cEwu8iz73_0),.clk(gclk));
	jdff dff_A_L7zAtZmE4_0(.dout(w_dff_A_dkg99LSj6_0),.din(w_dff_A_L7zAtZmE4_0),.clk(gclk));
	jdff dff_A_dkg99LSj6_0(.dout(w_dff_A_qjWZ4vUH3_0),.din(w_dff_A_dkg99LSj6_0),.clk(gclk));
	jdff dff_A_qjWZ4vUH3_0(.dout(w_dff_A_vTcdfKT48_0),.din(w_dff_A_qjWZ4vUH3_0),.clk(gclk));
	jdff dff_A_vTcdfKT48_0(.dout(w_dff_A_jwgxTFxz7_0),.din(w_dff_A_vTcdfKT48_0),.clk(gclk));
	jdff dff_A_jwgxTFxz7_0(.dout(w_dff_A_RYfOJeG11_0),.din(w_dff_A_jwgxTFxz7_0),.clk(gclk));
	jdff dff_A_RYfOJeG11_0(.dout(w_dff_A_EFLsrP0x4_0),.din(w_dff_A_RYfOJeG11_0),.clk(gclk));
	jdff dff_A_EFLsrP0x4_0(.dout(w_dff_A_m703jvyh6_0),.din(w_dff_A_EFLsrP0x4_0),.clk(gclk));
	jdff dff_A_m703jvyh6_0(.dout(G809),.din(w_dff_A_m703jvyh6_0),.clk(gclk));
	jdff dff_A_kHDc557D8_1(.dout(w_dff_A_tHQUoPYV4_0),.din(w_dff_A_kHDc557D8_1),.clk(gclk));
	jdff dff_A_tHQUoPYV4_0(.dout(w_dff_A_JWnk32uO1_0),.din(w_dff_A_tHQUoPYV4_0),.clk(gclk));
	jdff dff_A_JWnk32uO1_0(.dout(w_dff_A_6yfjsOLV6_0),.din(w_dff_A_JWnk32uO1_0),.clk(gclk));
	jdff dff_A_6yfjsOLV6_0(.dout(w_dff_A_RE9UljRM3_0),.din(w_dff_A_6yfjsOLV6_0),.clk(gclk));
	jdff dff_A_RE9UljRM3_0(.dout(w_dff_A_xPAN24Gg7_0),.din(w_dff_A_RE9UljRM3_0),.clk(gclk));
	jdff dff_A_xPAN24Gg7_0(.dout(w_dff_A_fRXrni0X7_0),.din(w_dff_A_xPAN24Gg7_0),.clk(gclk));
	jdff dff_A_fRXrni0X7_0(.dout(w_dff_A_JD4p8yJT9_0),.din(w_dff_A_fRXrni0X7_0),.clk(gclk));
	jdff dff_A_JD4p8yJT9_0(.dout(w_dff_A_UkgFFqRz4_0),.din(w_dff_A_JD4p8yJT9_0),.clk(gclk));
	jdff dff_A_UkgFFqRz4_0(.dout(w_dff_A_2fkSJ1ds0_0),.din(w_dff_A_UkgFFqRz4_0),.clk(gclk));
	jdff dff_A_2fkSJ1ds0_0(.dout(w_dff_A_sfopnZ7L9_0),.din(w_dff_A_2fkSJ1ds0_0),.clk(gclk));
	jdff dff_A_sfopnZ7L9_0(.dout(w_dff_A_mDvVVJk68_0),.din(w_dff_A_sfopnZ7L9_0),.clk(gclk));
	jdff dff_A_mDvVVJk68_0(.dout(w_dff_A_OxXF5fDc3_0),.din(w_dff_A_mDvVVJk68_0),.clk(gclk));
	jdff dff_A_OxXF5fDc3_0(.dout(w_dff_A_68sPz6aE4_0),.din(w_dff_A_OxXF5fDc3_0),.clk(gclk));
	jdff dff_A_68sPz6aE4_0(.dout(w_dff_A_poE1YTcD5_0),.din(w_dff_A_68sPz6aE4_0),.clk(gclk));
	jdff dff_A_poE1YTcD5_0(.dout(w_dff_A_JsQkrAfx1_0),.din(w_dff_A_poE1YTcD5_0),.clk(gclk));
	jdff dff_A_JsQkrAfx1_0(.dout(w_dff_A_U9Ahwjuy5_0),.din(w_dff_A_JsQkrAfx1_0),.clk(gclk));
	jdff dff_A_U9Ahwjuy5_0(.dout(w_dff_A_JsEbNU8Q7_0),.din(w_dff_A_U9Ahwjuy5_0),.clk(gclk));
	jdff dff_A_JsEbNU8Q7_0(.dout(w_dff_A_9kUhDqqt2_0),.din(w_dff_A_JsEbNU8Q7_0),.clk(gclk));
	jdff dff_A_9kUhDqqt2_0(.dout(w_dff_A_AFMP7DaI7_0),.din(w_dff_A_9kUhDqqt2_0),.clk(gclk));
	jdff dff_A_AFMP7DaI7_0(.dout(w_dff_A_SCLIygbe4_0),.din(w_dff_A_AFMP7DaI7_0),.clk(gclk));
	jdff dff_A_SCLIygbe4_0(.dout(w_dff_A_pEaPMiuy1_0),.din(w_dff_A_SCLIygbe4_0),.clk(gclk));
	jdff dff_A_pEaPMiuy1_0(.dout(w_dff_A_bEsuk1930_0),.din(w_dff_A_pEaPMiuy1_0),.clk(gclk));
	jdff dff_A_bEsuk1930_0(.dout(w_dff_A_TcJnLONY7_0),.din(w_dff_A_bEsuk1930_0),.clk(gclk));
	jdff dff_A_TcJnLONY7_0(.dout(w_dff_A_UD2G7XuA8_0),.din(w_dff_A_TcJnLONY7_0),.clk(gclk));
	jdff dff_A_UD2G7XuA8_0(.dout(w_dff_A_r7uy8L3S1_0),.din(w_dff_A_UD2G7XuA8_0),.clk(gclk));
	jdff dff_A_r7uy8L3S1_0(.dout(w_dff_A_rOjpEODb0_0),.din(w_dff_A_r7uy8L3S1_0),.clk(gclk));
	jdff dff_A_rOjpEODb0_0(.dout(w_dff_A_lzxLPuzi5_0),.din(w_dff_A_rOjpEODb0_0),.clk(gclk));
	jdff dff_A_lzxLPuzi5_0(.dout(G993),.din(w_dff_A_lzxLPuzi5_0),.clk(gclk));
	jdff dff_A_GL80qaD07_1(.dout(w_dff_A_kWakDpog6_0),.din(w_dff_A_GL80qaD07_1),.clk(gclk));
	jdff dff_A_kWakDpog6_0(.dout(w_dff_A_Vo1PcdKq3_0),.din(w_dff_A_kWakDpog6_0),.clk(gclk));
	jdff dff_A_Vo1PcdKq3_0(.dout(w_dff_A_lR0QA30s2_0),.din(w_dff_A_Vo1PcdKq3_0),.clk(gclk));
	jdff dff_A_lR0QA30s2_0(.dout(w_dff_A_vGJS5vWd8_0),.din(w_dff_A_lR0QA30s2_0),.clk(gclk));
	jdff dff_A_vGJS5vWd8_0(.dout(w_dff_A_ZHIt9AMD1_0),.din(w_dff_A_vGJS5vWd8_0),.clk(gclk));
	jdff dff_A_ZHIt9AMD1_0(.dout(w_dff_A_qEYSLesI6_0),.din(w_dff_A_ZHIt9AMD1_0),.clk(gclk));
	jdff dff_A_qEYSLesI6_0(.dout(w_dff_A_23jqGqgc6_0),.din(w_dff_A_qEYSLesI6_0),.clk(gclk));
	jdff dff_A_23jqGqgc6_0(.dout(w_dff_A_40ITOBCG8_0),.din(w_dff_A_23jqGqgc6_0),.clk(gclk));
	jdff dff_A_40ITOBCG8_0(.dout(w_dff_A_RhIRWPRt6_0),.din(w_dff_A_40ITOBCG8_0),.clk(gclk));
	jdff dff_A_RhIRWPRt6_0(.dout(w_dff_A_9rvfiyRD6_0),.din(w_dff_A_RhIRWPRt6_0),.clk(gclk));
	jdff dff_A_9rvfiyRD6_0(.dout(w_dff_A_3yITJfY47_0),.din(w_dff_A_9rvfiyRD6_0),.clk(gclk));
	jdff dff_A_3yITJfY47_0(.dout(w_dff_A_nHpMnFic5_0),.din(w_dff_A_3yITJfY47_0),.clk(gclk));
	jdff dff_A_nHpMnFic5_0(.dout(w_dff_A_IKOeYurh5_0),.din(w_dff_A_nHpMnFic5_0),.clk(gclk));
	jdff dff_A_IKOeYurh5_0(.dout(w_dff_A_blXyaCrD7_0),.din(w_dff_A_IKOeYurh5_0),.clk(gclk));
	jdff dff_A_blXyaCrD7_0(.dout(w_dff_A_dL4X1qm12_0),.din(w_dff_A_blXyaCrD7_0),.clk(gclk));
	jdff dff_A_dL4X1qm12_0(.dout(w_dff_A_j9OeQzmB7_0),.din(w_dff_A_dL4X1qm12_0),.clk(gclk));
	jdff dff_A_j9OeQzmB7_0(.dout(w_dff_A_OQoWEMgG1_0),.din(w_dff_A_j9OeQzmB7_0),.clk(gclk));
	jdff dff_A_OQoWEMgG1_0(.dout(w_dff_A_V5NDIerF7_0),.din(w_dff_A_OQoWEMgG1_0),.clk(gclk));
	jdff dff_A_V5NDIerF7_0(.dout(w_dff_A_TKmN7Ysz0_0),.din(w_dff_A_V5NDIerF7_0),.clk(gclk));
	jdff dff_A_TKmN7Ysz0_0(.dout(w_dff_A_2k7ESiSz6_0),.din(w_dff_A_TKmN7Ysz0_0),.clk(gclk));
	jdff dff_A_2k7ESiSz6_0(.dout(w_dff_A_whASYpX52_0),.din(w_dff_A_2k7ESiSz6_0),.clk(gclk));
	jdff dff_A_whASYpX52_0(.dout(w_dff_A_sWXcdNLY3_0),.din(w_dff_A_whASYpX52_0),.clk(gclk));
	jdff dff_A_sWXcdNLY3_0(.dout(w_dff_A_7PvL0IXM7_0),.din(w_dff_A_sWXcdNLY3_0),.clk(gclk));
	jdff dff_A_7PvL0IXM7_0(.dout(w_dff_A_d60VyGJu2_0),.din(w_dff_A_7PvL0IXM7_0),.clk(gclk));
	jdff dff_A_d60VyGJu2_0(.dout(w_dff_A_VZlvfsq45_0),.din(w_dff_A_d60VyGJu2_0),.clk(gclk));
	jdff dff_A_VZlvfsq45_0(.dout(w_dff_A_JhRE7CG32_0),.din(w_dff_A_VZlvfsq45_0),.clk(gclk));
	jdff dff_A_JhRE7CG32_0(.dout(w_dff_A_I4saYtgB8_0),.din(w_dff_A_JhRE7CG32_0),.clk(gclk));
	jdff dff_A_I4saYtgB8_0(.dout(G978),.din(w_dff_A_I4saYtgB8_0),.clk(gclk));
	jdff dff_A_DSogMvSP0_1(.dout(w_dff_A_C4gJVj634_0),.din(w_dff_A_DSogMvSP0_1),.clk(gclk));
	jdff dff_A_C4gJVj634_0(.dout(w_dff_A_dx9VHOy94_0),.din(w_dff_A_C4gJVj634_0),.clk(gclk));
	jdff dff_A_dx9VHOy94_0(.dout(w_dff_A_CGBEwkDY2_0),.din(w_dff_A_dx9VHOy94_0),.clk(gclk));
	jdff dff_A_CGBEwkDY2_0(.dout(w_dff_A_m0ldYnrN3_0),.din(w_dff_A_CGBEwkDY2_0),.clk(gclk));
	jdff dff_A_m0ldYnrN3_0(.dout(w_dff_A_tOL6xVWu9_0),.din(w_dff_A_m0ldYnrN3_0),.clk(gclk));
	jdff dff_A_tOL6xVWu9_0(.dout(w_dff_A_rpw6DQMo7_0),.din(w_dff_A_tOL6xVWu9_0),.clk(gclk));
	jdff dff_A_rpw6DQMo7_0(.dout(w_dff_A_857cWHrX9_0),.din(w_dff_A_rpw6DQMo7_0),.clk(gclk));
	jdff dff_A_857cWHrX9_0(.dout(w_dff_A_Xic6uetH5_0),.din(w_dff_A_857cWHrX9_0),.clk(gclk));
	jdff dff_A_Xic6uetH5_0(.dout(w_dff_A_ZNXKv3sL5_0),.din(w_dff_A_Xic6uetH5_0),.clk(gclk));
	jdff dff_A_ZNXKv3sL5_0(.dout(w_dff_A_OX3jQDPM7_0),.din(w_dff_A_ZNXKv3sL5_0),.clk(gclk));
	jdff dff_A_OX3jQDPM7_0(.dout(w_dff_A_Y4R5hK3X2_0),.din(w_dff_A_OX3jQDPM7_0),.clk(gclk));
	jdff dff_A_Y4R5hK3X2_0(.dout(w_dff_A_YECpAPEX6_0),.din(w_dff_A_Y4R5hK3X2_0),.clk(gclk));
	jdff dff_A_YECpAPEX6_0(.dout(w_dff_A_Z5tanN8y8_0),.din(w_dff_A_YECpAPEX6_0),.clk(gclk));
	jdff dff_A_Z5tanN8y8_0(.dout(w_dff_A_SEbXML8t1_0),.din(w_dff_A_Z5tanN8y8_0),.clk(gclk));
	jdff dff_A_SEbXML8t1_0(.dout(w_dff_A_kiILA36z4_0),.din(w_dff_A_SEbXML8t1_0),.clk(gclk));
	jdff dff_A_kiILA36z4_0(.dout(w_dff_A_dduyINLq4_0),.din(w_dff_A_kiILA36z4_0),.clk(gclk));
	jdff dff_A_dduyINLq4_0(.dout(w_dff_A_yh9MxF8o9_0),.din(w_dff_A_dduyINLq4_0),.clk(gclk));
	jdff dff_A_yh9MxF8o9_0(.dout(w_dff_A_fSJicmTz9_0),.din(w_dff_A_yh9MxF8o9_0),.clk(gclk));
	jdff dff_A_fSJicmTz9_0(.dout(w_dff_A_hU4Mgo6l2_0),.din(w_dff_A_fSJicmTz9_0),.clk(gclk));
	jdff dff_A_hU4Mgo6l2_0(.dout(w_dff_A_Ecj0khgj6_0),.din(w_dff_A_hU4Mgo6l2_0),.clk(gclk));
	jdff dff_A_Ecj0khgj6_0(.dout(w_dff_A_YdIz7Gjr0_0),.din(w_dff_A_Ecj0khgj6_0),.clk(gclk));
	jdff dff_A_YdIz7Gjr0_0(.dout(w_dff_A_d4UBJGGz6_0),.din(w_dff_A_YdIz7Gjr0_0),.clk(gclk));
	jdff dff_A_d4UBJGGz6_0(.dout(w_dff_A_lBds5kpI7_0),.din(w_dff_A_d4UBJGGz6_0),.clk(gclk));
	jdff dff_A_lBds5kpI7_0(.dout(w_dff_A_oyPXV0ai1_0),.din(w_dff_A_lBds5kpI7_0),.clk(gclk));
	jdff dff_A_oyPXV0ai1_0(.dout(w_dff_A_sHd6jvbM1_0),.din(w_dff_A_oyPXV0ai1_0),.clk(gclk));
	jdff dff_A_sHd6jvbM1_0(.dout(w_dff_A_e3O8wnjN1_0),.din(w_dff_A_sHd6jvbM1_0),.clk(gclk));
	jdff dff_A_e3O8wnjN1_0(.dout(w_dff_A_13metCxG7_0),.din(w_dff_A_e3O8wnjN1_0),.clk(gclk));
	jdff dff_A_13metCxG7_0(.dout(G949),.din(w_dff_A_13metCxG7_0),.clk(gclk));
	jdff dff_A_icCkjrtN9_1(.dout(w_dff_A_19iUWqEI7_0),.din(w_dff_A_icCkjrtN9_1),.clk(gclk));
	jdff dff_A_19iUWqEI7_0(.dout(w_dff_A_JnRpjgjB5_0),.din(w_dff_A_19iUWqEI7_0),.clk(gclk));
	jdff dff_A_JnRpjgjB5_0(.dout(w_dff_A_Rawa0EVo0_0),.din(w_dff_A_JnRpjgjB5_0),.clk(gclk));
	jdff dff_A_Rawa0EVo0_0(.dout(w_dff_A_zZsP4AEc1_0),.din(w_dff_A_Rawa0EVo0_0),.clk(gclk));
	jdff dff_A_zZsP4AEc1_0(.dout(w_dff_A_RbIpnAqe4_0),.din(w_dff_A_zZsP4AEc1_0),.clk(gclk));
	jdff dff_A_RbIpnAqe4_0(.dout(w_dff_A_BTU9xes56_0),.din(w_dff_A_RbIpnAqe4_0),.clk(gclk));
	jdff dff_A_BTU9xes56_0(.dout(w_dff_A_y2nK58US2_0),.din(w_dff_A_BTU9xes56_0),.clk(gclk));
	jdff dff_A_y2nK58US2_0(.dout(w_dff_A_O8WNIf8A1_0),.din(w_dff_A_y2nK58US2_0),.clk(gclk));
	jdff dff_A_O8WNIf8A1_0(.dout(w_dff_A_OCtkCjLF7_0),.din(w_dff_A_O8WNIf8A1_0),.clk(gclk));
	jdff dff_A_OCtkCjLF7_0(.dout(w_dff_A_M7MSGmvC2_0),.din(w_dff_A_OCtkCjLF7_0),.clk(gclk));
	jdff dff_A_M7MSGmvC2_0(.dout(w_dff_A_Yn9lY7Bv8_0),.din(w_dff_A_M7MSGmvC2_0),.clk(gclk));
	jdff dff_A_Yn9lY7Bv8_0(.dout(w_dff_A_fvxQu5hT4_0),.din(w_dff_A_Yn9lY7Bv8_0),.clk(gclk));
	jdff dff_A_fvxQu5hT4_0(.dout(w_dff_A_HKulKoja1_0),.din(w_dff_A_fvxQu5hT4_0),.clk(gclk));
	jdff dff_A_HKulKoja1_0(.dout(w_dff_A_tBJlzOuX6_0),.din(w_dff_A_HKulKoja1_0),.clk(gclk));
	jdff dff_A_tBJlzOuX6_0(.dout(w_dff_A_xHdlANjI3_0),.din(w_dff_A_tBJlzOuX6_0),.clk(gclk));
	jdff dff_A_xHdlANjI3_0(.dout(w_dff_A_KhBIWZB19_0),.din(w_dff_A_xHdlANjI3_0),.clk(gclk));
	jdff dff_A_KhBIWZB19_0(.dout(w_dff_A_XHIJn5oW8_0),.din(w_dff_A_KhBIWZB19_0),.clk(gclk));
	jdff dff_A_XHIJn5oW8_0(.dout(w_dff_A_BWzNvPEo9_0),.din(w_dff_A_XHIJn5oW8_0),.clk(gclk));
	jdff dff_A_BWzNvPEo9_0(.dout(w_dff_A_mK02EGtM5_0),.din(w_dff_A_BWzNvPEo9_0),.clk(gclk));
	jdff dff_A_mK02EGtM5_0(.dout(w_dff_A_AAp6yyvL6_0),.din(w_dff_A_mK02EGtM5_0),.clk(gclk));
	jdff dff_A_AAp6yyvL6_0(.dout(w_dff_A_JVPlbqT78_0),.din(w_dff_A_AAp6yyvL6_0),.clk(gclk));
	jdff dff_A_JVPlbqT78_0(.dout(w_dff_A_b2uXC3is0_0),.din(w_dff_A_JVPlbqT78_0),.clk(gclk));
	jdff dff_A_b2uXC3is0_0(.dout(w_dff_A_YnxnsBmf6_0),.din(w_dff_A_b2uXC3is0_0),.clk(gclk));
	jdff dff_A_YnxnsBmf6_0(.dout(w_dff_A_EjOPzYaz8_0),.din(w_dff_A_YnxnsBmf6_0),.clk(gclk));
	jdff dff_A_EjOPzYaz8_0(.dout(w_dff_A_Q5HRcTLO0_0),.din(w_dff_A_EjOPzYaz8_0),.clk(gclk));
	jdff dff_A_Q5HRcTLO0_0(.dout(w_dff_A_NSEEvzcA4_0),.din(w_dff_A_Q5HRcTLO0_0),.clk(gclk));
	jdff dff_A_NSEEvzcA4_0(.dout(w_dff_A_Juz5QEP89_0),.din(w_dff_A_NSEEvzcA4_0),.clk(gclk));
	jdff dff_A_Juz5QEP89_0(.dout(G939),.din(w_dff_A_Juz5QEP89_0),.clk(gclk));
	jdff dff_A_fys1SLwP5_1(.dout(w_dff_A_03AV6cOF7_0),.din(w_dff_A_fys1SLwP5_1),.clk(gclk));
	jdff dff_A_03AV6cOF7_0(.dout(w_dff_A_YNtWI2A51_0),.din(w_dff_A_03AV6cOF7_0),.clk(gclk));
	jdff dff_A_YNtWI2A51_0(.dout(w_dff_A_n0hVXxYY0_0),.din(w_dff_A_YNtWI2A51_0),.clk(gclk));
	jdff dff_A_n0hVXxYY0_0(.dout(w_dff_A_6oHBMrwI7_0),.din(w_dff_A_n0hVXxYY0_0),.clk(gclk));
	jdff dff_A_6oHBMrwI7_0(.dout(w_dff_A_yViWC5cv3_0),.din(w_dff_A_6oHBMrwI7_0),.clk(gclk));
	jdff dff_A_yViWC5cv3_0(.dout(w_dff_A_iSnmxgFp8_0),.din(w_dff_A_yViWC5cv3_0),.clk(gclk));
	jdff dff_A_iSnmxgFp8_0(.dout(w_dff_A_yUeI6QGd8_0),.din(w_dff_A_iSnmxgFp8_0),.clk(gclk));
	jdff dff_A_yUeI6QGd8_0(.dout(w_dff_A_f5lYtiih3_0),.din(w_dff_A_yUeI6QGd8_0),.clk(gclk));
	jdff dff_A_f5lYtiih3_0(.dout(w_dff_A_XCjfE83U0_0),.din(w_dff_A_f5lYtiih3_0),.clk(gclk));
	jdff dff_A_XCjfE83U0_0(.dout(w_dff_A_jttIpTwo5_0),.din(w_dff_A_XCjfE83U0_0),.clk(gclk));
	jdff dff_A_jttIpTwo5_0(.dout(w_dff_A_sQOSlP209_0),.din(w_dff_A_jttIpTwo5_0),.clk(gclk));
	jdff dff_A_sQOSlP209_0(.dout(w_dff_A_ZaPRMZIa9_0),.din(w_dff_A_sQOSlP209_0),.clk(gclk));
	jdff dff_A_ZaPRMZIa9_0(.dout(w_dff_A_dhrTnkyF2_0),.din(w_dff_A_ZaPRMZIa9_0),.clk(gclk));
	jdff dff_A_dhrTnkyF2_0(.dout(w_dff_A_mlgafr6e8_0),.din(w_dff_A_dhrTnkyF2_0),.clk(gclk));
	jdff dff_A_mlgafr6e8_0(.dout(w_dff_A_TI1mhfOY5_0),.din(w_dff_A_mlgafr6e8_0),.clk(gclk));
	jdff dff_A_TI1mhfOY5_0(.dout(w_dff_A_eeH0C1ff1_0),.din(w_dff_A_TI1mhfOY5_0),.clk(gclk));
	jdff dff_A_eeH0C1ff1_0(.dout(w_dff_A_Tie7n15P6_0),.din(w_dff_A_eeH0C1ff1_0),.clk(gclk));
	jdff dff_A_Tie7n15P6_0(.dout(w_dff_A_zHTmS7JN2_0),.din(w_dff_A_Tie7n15P6_0),.clk(gclk));
	jdff dff_A_zHTmS7JN2_0(.dout(w_dff_A_JawBmFkl7_0),.din(w_dff_A_zHTmS7JN2_0),.clk(gclk));
	jdff dff_A_JawBmFkl7_0(.dout(w_dff_A_nV7evQ6t1_0),.din(w_dff_A_JawBmFkl7_0),.clk(gclk));
	jdff dff_A_nV7evQ6t1_0(.dout(w_dff_A_m7gYe2MG0_0),.din(w_dff_A_nV7evQ6t1_0),.clk(gclk));
	jdff dff_A_m7gYe2MG0_0(.dout(w_dff_A_hh9qEkVP6_0),.din(w_dff_A_m7gYe2MG0_0),.clk(gclk));
	jdff dff_A_hh9qEkVP6_0(.dout(w_dff_A_wvsdtkKl5_0),.din(w_dff_A_hh9qEkVP6_0),.clk(gclk));
	jdff dff_A_wvsdtkKl5_0(.dout(w_dff_A_vWk6R8zK2_0),.din(w_dff_A_wvsdtkKl5_0),.clk(gclk));
	jdff dff_A_vWk6R8zK2_0(.dout(w_dff_A_q1qOcbL21_0),.din(w_dff_A_vWk6R8zK2_0),.clk(gclk));
	jdff dff_A_q1qOcbL21_0(.dout(w_dff_A_pjZozWlJ0_0),.din(w_dff_A_q1qOcbL21_0),.clk(gclk));
	jdff dff_A_pjZozWlJ0_0(.dout(w_dff_A_kqgBN8412_0),.din(w_dff_A_pjZozWlJ0_0),.clk(gclk));
	jdff dff_A_kqgBN8412_0(.dout(G889),.din(w_dff_A_kqgBN8412_0),.clk(gclk));
	jdff dff_A_ugDvOh8h3_1(.dout(w_dff_A_hsZh9E3t1_0),.din(w_dff_A_ugDvOh8h3_1),.clk(gclk));
	jdff dff_A_hsZh9E3t1_0(.dout(w_dff_A_Ic0JfziH3_0),.din(w_dff_A_hsZh9E3t1_0),.clk(gclk));
	jdff dff_A_Ic0JfziH3_0(.dout(w_dff_A_bueculMr9_0),.din(w_dff_A_Ic0JfziH3_0),.clk(gclk));
	jdff dff_A_bueculMr9_0(.dout(w_dff_A_iVmqxflh9_0),.din(w_dff_A_bueculMr9_0),.clk(gclk));
	jdff dff_A_iVmqxflh9_0(.dout(w_dff_A_zx7i1Ip78_0),.din(w_dff_A_iVmqxflh9_0),.clk(gclk));
	jdff dff_A_zx7i1Ip78_0(.dout(w_dff_A_vqDgRTU94_0),.din(w_dff_A_zx7i1Ip78_0),.clk(gclk));
	jdff dff_A_vqDgRTU94_0(.dout(w_dff_A_uYPb1Vht7_0),.din(w_dff_A_vqDgRTU94_0),.clk(gclk));
	jdff dff_A_uYPb1Vht7_0(.dout(w_dff_A_hg3tWgNL8_0),.din(w_dff_A_uYPb1Vht7_0),.clk(gclk));
	jdff dff_A_hg3tWgNL8_0(.dout(w_dff_A_nQHuPJJa7_0),.din(w_dff_A_hg3tWgNL8_0),.clk(gclk));
	jdff dff_A_nQHuPJJa7_0(.dout(w_dff_A_KerKxsGh9_0),.din(w_dff_A_nQHuPJJa7_0),.clk(gclk));
	jdff dff_A_KerKxsGh9_0(.dout(w_dff_A_GvDcWhrR9_0),.din(w_dff_A_KerKxsGh9_0),.clk(gclk));
	jdff dff_A_GvDcWhrR9_0(.dout(w_dff_A_HALWxpLy7_0),.din(w_dff_A_GvDcWhrR9_0),.clk(gclk));
	jdff dff_A_HALWxpLy7_0(.dout(w_dff_A_SD9aFa6x9_0),.din(w_dff_A_HALWxpLy7_0),.clk(gclk));
	jdff dff_A_SD9aFa6x9_0(.dout(w_dff_A_LVOW0u2p2_0),.din(w_dff_A_SD9aFa6x9_0),.clk(gclk));
	jdff dff_A_LVOW0u2p2_0(.dout(w_dff_A_akyrYSbX9_0),.din(w_dff_A_LVOW0u2p2_0),.clk(gclk));
	jdff dff_A_akyrYSbX9_0(.dout(w_dff_A_nGWzfI9f7_0),.din(w_dff_A_akyrYSbX9_0),.clk(gclk));
	jdff dff_A_nGWzfI9f7_0(.dout(w_dff_A_J3WM7dtJ3_0),.din(w_dff_A_nGWzfI9f7_0),.clk(gclk));
	jdff dff_A_J3WM7dtJ3_0(.dout(w_dff_A_RHOYpTgT5_0),.din(w_dff_A_J3WM7dtJ3_0),.clk(gclk));
	jdff dff_A_RHOYpTgT5_0(.dout(w_dff_A_oo7IHECP7_0),.din(w_dff_A_RHOYpTgT5_0),.clk(gclk));
	jdff dff_A_oo7IHECP7_0(.dout(w_dff_A_ydeQ5ayO5_0),.din(w_dff_A_oo7IHECP7_0),.clk(gclk));
	jdff dff_A_ydeQ5ayO5_0(.dout(w_dff_A_hZYUJVo60_0),.din(w_dff_A_ydeQ5ayO5_0),.clk(gclk));
	jdff dff_A_hZYUJVo60_0(.dout(w_dff_A_EsKHFbn93_0),.din(w_dff_A_hZYUJVo60_0),.clk(gclk));
	jdff dff_A_EsKHFbn93_0(.dout(w_dff_A_ssxZdoPJ9_0),.din(w_dff_A_EsKHFbn93_0),.clk(gclk));
	jdff dff_A_ssxZdoPJ9_0(.dout(w_dff_A_7X0MkftL8_0),.din(w_dff_A_ssxZdoPJ9_0),.clk(gclk));
	jdff dff_A_7X0MkftL8_0(.dout(w_dff_A_YtbrXaaO6_0),.din(w_dff_A_7X0MkftL8_0),.clk(gclk));
	jdff dff_A_YtbrXaaO6_0(.dout(w_dff_A_f5apguHw2_0),.din(w_dff_A_YtbrXaaO6_0),.clk(gclk));
	jdff dff_A_f5apguHw2_0(.dout(G593),.din(w_dff_A_f5apguHw2_0),.clk(gclk));
	jdff dff_A_1oUSV6XM4_2(.dout(w_dff_A_nC0NXBua2_0),.din(w_dff_A_1oUSV6XM4_2),.clk(gclk));
	jdff dff_A_nC0NXBua2_0(.dout(w_dff_A_ZQbu3un66_0),.din(w_dff_A_nC0NXBua2_0),.clk(gclk));
	jdff dff_A_ZQbu3un66_0(.dout(w_dff_A_CXKX5Dup2_0),.din(w_dff_A_ZQbu3un66_0),.clk(gclk));
	jdff dff_A_CXKX5Dup2_0(.dout(w_dff_A_BKwKrpvP4_0),.din(w_dff_A_CXKX5Dup2_0),.clk(gclk));
	jdff dff_A_BKwKrpvP4_0(.dout(w_dff_A_4QXByxUV8_0),.din(w_dff_A_BKwKrpvP4_0),.clk(gclk));
	jdff dff_A_4QXByxUV8_0(.dout(w_dff_A_BQEhQaQ47_0),.din(w_dff_A_4QXByxUV8_0),.clk(gclk));
	jdff dff_A_BQEhQaQ47_0(.dout(w_dff_A_TZB0iEli7_0),.din(w_dff_A_BQEhQaQ47_0),.clk(gclk));
	jdff dff_A_TZB0iEli7_0(.dout(w_dff_A_0nHBNFlf5_0),.din(w_dff_A_TZB0iEli7_0),.clk(gclk));
	jdff dff_A_0nHBNFlf5_0(.dout(w_dff_A_8DkTLxmb9_0),.din(w_dff_A_0nHBNFlf5_0),.clk(gclk));
	jdff dff_A_8DkTLxmb9_0(.dout(w_dff_A_ufmbZPiW9_0),.din(w_dff_A_8DkTLxmb9_0),.clk(gclk));
	jdff dff_A_ufmbZPiW9_0(.dout(w_dff_A_njwkmYS01_0),.din(w_dff_A_ufmbZPiW9_0),.clk(gclk));
	jdff dff_A_njwkmYS01_0(.dout(w_dff_A_WANDuyqQ2_0),.din(w_dff_A_njwkmYS01_0),.clk(gclk));
	jdff dff_A_WANDuyqQ2_0(.dout(w_dff_A_zNyzGZ896_0),.din(w_dff_A_WANDuyqQ2_0),.clk(gclk));
	jdff dff_A_zNyzGZ896_0(.dout(w_dff_A_iSUqzAb20_0),.din(w_dff_A_zNyzGZ896_0),.clk(gclk));
	jdff dff_A_iSUqzAb20_0(.dout(w_dff_A_1hIRuFMn4_0),.din(w_dff_A_iSUqzAb20_0),.clk(gclk));
	jdff dff_A_1hIRuFMn4_0(.dout(w_dff_A_kirutSCW2_0),.din(w_dff_A_1hIRuFMn4_0),.clk(gclk));
	jdff dff_A_kirutSCW2_0(.dout(w_dff_A_XnZSXl2U4_0),.din(w_dff_A_kirutSCW2_0),.clk(gclk));
	jdff dff_A_XnZSXl2U4_0(.dout(w_dff_A_qReVuPGl6_0),.din(w_dff_A_XnZSXl2U4_0),.clk(gclk));
	jdff dff_A_qReVuPGl6_0(.dout(w_dff_A_zOtnA8He2_0),.din(w_dff_A_qReVuPGl6_0),.clk(gclk));
	jdff dff_A_zOtnA8He2_0(.dout(w_dff_A_Bi5hURtT2_0),.din(w_dff_A_zOtnA8He2_0),.clk(gclk));
	jdff dff_A_Bi5hURtT2_0(.dout(w_dff_A_9VEz5i4k0_0),.din(w_dff_A_Bi5hURtT2_0),.clk(gclk));
	jdff dff_A_9VEz5i4k0_0(.dout(w_dff_A_LQbAxgAT1_0),.din(w_dff_A_9VEz5i4k0_0),.clk(gclk));
	jdff dff_A_LQbAxgAT1_0(.dout(w_dff_A_QGLXUlOm7_0),.din(w_dff_A_LQbAxgAT1_0),.clk(gclk));
	jdff dff_A_QGLXUlOm7_0(.dout(G636),.din(w_dff_A_QGLXUlOm7_0),.clk(gclk));
	jdff dff_A_Z3ftPUiG7_2(.dout(w_dff_A_zrVz5la56_0),.din(w_dff_A_Z3ftPUiG7_2),.clk(gclk));
	jdff dff_A_zrVz5la56_0(.dout(w_dff_A_bCStDZfy2_0),.din(w_dff_A_zrVz5la56_0),.clk(gclk));
	jdff dff_A_bCStDZfy2_0(.dout(w_dff_A_Ra7FCRXm2_0),.din(w_dff_A_bCStDZfy2_0),.clk(gclk));
	jdff dff_A_Ra7FCRXm2_0(.dout(w_dff_A_7n7Jb1vb1_0),.din(w_dff_A_Ra7FCRXm2_0),.clk(gclk));
	jdff dff_A_7n7Jb1vb1_0(.dout(w_dff_A_lUVkydTd9_0),.din(w_dff_A_7n7Jb1vb1_0),.clk(gclk));
	jdff dff_A_lUVkydTd9_0(.dout(w_dff_A_s24DJm9f7_0),.din(w_dff_A_lUVkydTd9_0),.clk(gclk));
	jdff dff_A_s24DJm9f7_0(.dout(w_dff_A_HpQvrubS3_0),.din(w_dff_A_s24DJm9f7_0),.clk(gclk));
	jdff dff_A_HpQvrubS3_0(.dout(w_dff_A_8Ao1vih75_0),.din(w_dff_A_HpQvrubS3_0),.clk(gclk));
	jdff dff_A_8Ao1vih75_0(.dout(w_dff_A_EWiY3Q5b1_0),.din(w_dff_A_8Ao1vih75_0),.clk(gclk));
	jdff dff_A_EWiY3Q5b1_0(.dout(w_dff_A_odf1XUXH9_0),.din(w_dff_A_EWiY3Q5b1_0),.clk(gclk));
	jdff dff_A_odf1XUXH9_0(.dout(w_dff_A_i4hdn9WJ7_0),.din(w_dff_A_odf1XUXH9_0),.clk(gclk));
	jdff dff_A_i4hdn9WJ7_0(.dout(w_dff_A_VNFg8XVd8_0),.din(w_dff_A_i4hdn9WJ7_0),.clk(gclk));
	jdff dff_A_VNFg8XVd8_0(.dout(w_dff_A_gRbGBBeR8_0),.din(w_dff_A_VNFg8XVd8_0),.clk(gclk));
	jdff dff_A_gRbGBBeR8_0(.dout(w_dff_A_PXEivqZw7_0),.din(w_dff_A_gRbGBBeR8_0),.clk(gclk));
	jdff dff_A_PXEivqZw7_0(.dout(w_dff_A_FudwoYCP4_0),.din(w_dff_A_PXEivqZw7_0),.clk(gclk));
	jdff dff_A_FudwoYCP4_0(.dout(w_dff_A_myuVa9p54_0),.din(w_dff_A_FudwoYCP4_0),.clk(gclk));
	jdff dff_A_myuVa9p54_0(.dout(w_dff_A_NO1QizLD5_0),.din(w_dff_A_myuVa9p54_0),.clk(gclk));
	jdff dff_A_NO1QizLD5_0(.dout(w_dff_A_NwC58MJ06_0),.din(w_dff_A_NO1QizLD5_0),.clk(gclk));
	jdff dff_A_NwC58MJ06_0(.dout(w_dff_A_LpCHxOlX5_0),.din(w_dff_A_NwC58MJ06_0),.clk(gclk));
	jdff dff_A_LpCHxOlX5_0(.dout(w_dff_A_QWjWVOXW1_0),.din(w_dff_A_LpCHxOlX5_0),.clk(gclk));
	jdff dff_A_QWjWVOXW1_0(.dout(w_dff_A_jHdqJ5y54_0),.din(w_dff_A_QWjWVOXW1_0),.clk(gclk));
	jdff dff_A_jHdqJ5y54_0(.dout(w_dff_A_Y7kUXdtv0_0),.din(w_dff_A_jHdqJ5y54_0),.clk(gclk));
	jdff dff_A_Y7kUXdtv0_0(.dout(w_dff_A_O29KIGL57_0),.din(w_dff_A_Y7kUXdtv0_0),.clk(gclk));
	jdff dff_A_O29KIGL57_0(.dout(G704),.din(w_dff_A_O29KIGL57_0),.clk(gclk));
	jdff dff_A_3bTGddH80_2(.dout(w_dff_A_HCmD40Ox0_0),.din(w_dff_A_3bTGddH80_2),.clk(gclk));
	jdff dff_A_HCmD40Ox0_0(.dout(w_dff_A_ds1O7zvS3_0),.din(w_dff_A_HCmD40Ox0_0),.clk(gclk));
	jdff dff_A_ds1O7zvS3_0(.dout(w_dff_A_8pNByWip8_0),.din(w_dff_A_ds1O7zvS3_0),.clk(gclk));
	jdff dff_A_8pNByWip8_0(.dout(w_dff_A_KYO7g1q22_0),.din(w_dff_A_8pNByWip8_0),.clk(gclk));
	jdff dff_A_KYO7g1q22_0(.dout(w_dff_A_8cNRoMUS5_0),.din(w_dff_A_KYO7g1q22_0),.clk(gclk));
	jdff dff_A_8cNRoMUS5_0(.dout(w_dff_A_uJb5aO7c0_0),.din(w_dff_A_8cNRoMUS5_0),.clk(gclk));
	jdff dff_A_uJb5aO7c0_0(.dout(w_dff_A_x1vViBng8_0),.din(w_dff_A_uJb5aO7c0_0),.clk(gclk));
	jdff dff_A_x1vViBng8_0(.dout(w_dff_A_1uY6diiv4_0),.din(w_dff_A_x1vViBng8_0),.clk(gclk));
	jdff dff_A_1uY6diiv4_0(.dout(w_dff_A_eAMttTla5_0),.din(w_dff_A_1uY6diiv4_0),.clk(gclk));
	jdff dff_A_eAMttTla5_0(.dout(w_dff_A_OfXwfuHb9_0),.din(w_dff_A_eAMttTla5_0),.clk(gclk));
	jdff dff_A_OfXwfuHb9_0(.dout(w_dff_A_gWMkCEob1_0),.din(w_dff_A_OfXwfuHb9_0),.clk(gclk));
	jdff dff_A_gWMkCEob1_0(.dout(w_dff_A_oF59FTBX1_0),.din(w_dff_A_gWMkCEob1_0),.clk(gclk));
	jdff dff_A_oF59FTBX1_0(.dout(w_dff_A_NDELbzed2_0),.din(w_dff_A_oF59FTBX1_0),.clk(gclk));
	jdff dff_A_NDELbzed2_0(.dout(w_dff_A_ymAq8dQA9_0),.din(w_dff_A_NDELbzed2_0),.clk(gclk));
	jdff dff_A_ymAq8dQA9_0(.dout(w_dff_A_WlU1xGcq3_0),.din(w_dff_A_ymAq8dQA9_0),.clk(gclk));
	jdff dff_A_WlU1xGcq3_0(.dout(w_dff_A_NfW3AOru4_0),.din(w_dff_A_WlU1xGcq3_0),.clk(gclk));
	jdff dff_A_NfW3AOru4_0(.dout(w_dff_A_8Dz2EDTB9_0),.din(w_dff_A_NfW3AOru4_0),.clk(gclk));
	jdff dff_A_8Dz2EDTB9_0(.dout(w_dff_A_uBZOwhgZ3_0),.din(w_dff_A_8Dz2EDTB9_0),.clk(gclk));
	jdff dff_A_uBZOwhgZ3_0(.dout(w_dff_A_uPz3MWrE4_0),.din(w_dff_A_uBZOwhgZ3_0),.clk(gclk));
	jdff dff_A_uPz3MWrE4_0(.dout(w_dff_A_uyJTFp7l6_0),.din(w_dff_A_uPz3MWrE4_0),.clk(gclk));
	jdff dff_A_uyJTFp7l6_0(.dout(w_dff_A_BXQ9Qi7n6_0),.din(w_dff_A_uyJTFp7l6_0),.clk(gclk));
	jdff dff_A_BXQ9Qi7n6_0(.dout(w_dff_A_Ym7FKmPV3_0),.din(w_dff_A_BXQ9Qi7n6_0),.clk(gclk));
	jdff dff_A_Ym7FKmPV3_0(.dout(w_dff_A_NtDooD8A4_0),.din(w_dff_A_Ym7FKmPV3_0),.clk(gclk));
	jdff dff_A_NtDooD8A4_0(.dout(G717),.din(w_dff_A_NtDooD8A4_0),.clk(gclk));
	jdff dff_A_a4NcGCQI4_2(.dout(w_dff_A_QKnPcnPn2_0),.din(w_dff_A_a4NcGCQI4_2),.clk(gclk));
	jdff dff_A_QKnPcnPn2_0(.dout(w_dff_A_Hao5ODkW2_0),.din(w_dff_A_QKnPcnPn2_0),.clk(gclk));
	jdff dff_A_Hao5ODkW2_0(.dout(w_dff_A_EcaA0shY7_0),.din(w_dff_A_Hao5ODkW2_0),.clk(gclk));
	jdff dff_A_EcaA0shY7_0(.dout(w_dff_A_ZAwsnKGm4_0),.din(w_dff_A_EcaA0shY7_0),.clk(gclk));
	jdff dff_A_ZAwsnKGm4_0(.dout(w_dff_A_OxrKGEvZ3_0),.din(w_dff_A_ZAwsnKGm4_0),.clk(gclk));
	jdff dff_A_OxrKGEvZ3_0(.dout(w_dff_A_NOStlwC57_0),.din(w_dff_A_OxrKGEvZ3_0),.clk(gclk));
	jdff dff_A_NOStlwC57_0(.dout(w_dff_A_9YIZJniB0_0),.din(w_dff_A_NOStlwC57_0),.clk(gclk));
	jdff dff_A_9YIZJniB0_0(.dout(w_dff_A_yG9z7hDW0_0),.din(w_dff_A_9YIZJniB0_0),.clk(gclk));
	jdff dff_A_yG9z7hDW0_0(.dout(w_dff_A_Q9KC1zNf3_0),.din(w_dff_A_yG9z7hDW0_0),.clk(gclk));
	jdff dff_A_Q9KC1zNf3_0(.dout(w_dff_A_OSNP0dIS0_0),.din(w_dff_A_Q9KC1zNf3_0),.clk(gclk));
	jdff dff_A_OSNP0dIS0_0(.dout(w_dff_A_yVb18zSB1_0),.din(w_dff_A_OSNP0dIS0_0),.clk(gclk));
	jdff dff_A_yVb18zSB1_0(.dout(w_dff_A_MDeFogBm4_0),.din(w_dff_A_yVb18zSB1_0),.clk(gclk));
	jdff dff_A_MDeFogBm4_0(.dout(w_dff_A_4TGxZztf4_0),.din(w_dff_A_MDeFogBm4_0),.clk(gclk));
	jdff dff_A_4TGxZztf4_0(.dout(w_dff_A_dURurCjF6_0),.din(w_dff_A_4TGxZztf4_0),.clk(gclk));
	jdff dff_A_dURurCjF6_0(.dout(w_dff_A_MB8IZYMQ1_0),.din(w_dff_A_dURurCjF6_0),.clk(gclk));
	jdff dff_A_MB8IZYMQ1_0(.dout(w_dff_A_vjfKkrUX7_0),.din(w_dff_A_MB8IZYMQ1_0),.clk(gclk));
	jdff dff_A_vjfKkrUX7_0(.dout(w_dff_A_yQwX7LmR1_0),.din(w_dff_A_vjfKkrUX7_0),.clk(gclk));
	jdff dff_A_yQwX7LmR1_0(.dout(w_dff_A_ImnVyFQH6_0),.din(w_dff_A_yQwX7LmR1_0),.clk(gclk));
	jdff dff_A_ImnVyFQH6_0(.dout(w_dff_A_pcj3Bf2f3_0),.din(w_dff_A_ImnVyFQH6_0),.clk(gclk));
	jdff dff_A_pcj3Bf2f3_0(.dout(w_dff_A_dO4I6j6B6_0),.din(w_dff_A_pcj3Bf2f3_0),.clk(gclk));
	jdff dff_A_dO4I6j6B6_0(.dout(w_dff_A_ZXNNfepP5_0),.din(w_dff_A_dO4I6j6B6_0),.clk(gclk));
	jdff dff_A_ZXNNfepP5_0(.dout(w_dff_A_nMfCKEhz9_0),.din(w_dff_A_ZXNNfepP5_0),.clk(gclk));
	jdff dff_A_nMfCKEhz9_0(.dout(w_dff_A_cisNgDn53_0),.din(w_dff_A_nMfCKEhz9_0),.clk(gclk));
	jdff dff_A_cisNgDn53_0(.dout(w_dff_A_lfGETm8V7_0),.din(w_dff_A_cisNgDn53_0),.clk(gclk));
	jdff dff_A_lfGETm8V7_0(.dout(G820),.din(w_dff_A_lfGETm8V7_0),.clk(gclk));
	jdff dff_A_InPKo1G29_2(.dout(w_dff_A_RwKtsVDd3_0),.din(w_dff_A_InPKo1G29_2),.clk(gclk));
	jdff dff_A_RwKtsVDd3_0(.dout(w_dff_A_TVtmQzl49_0),.din(w_dff_A_RwKtsVDd3_0),.clk(gclk));
	jdff dff_A_TVtmQzl49_0(.dout(w_dff_A_uTmujb7u3_0),.din(w_dff_A_TVtmQzl49_0),.clk(gclk));
	jdff dff_A_uTmujb7u3_0(.dout(w_dff_A_wPBheNWZ1_0),.din(w_dff_A_uTmujb7u3_0),.clk(gclk));
	jdff dff_A_wPBheNWZ1_0(.dout(w_dff_A_uTPbD6A49_0),.din(w_dff_A_wPBheNWZ1_0),.clk(gclk));
	jdff dff_A_uTPbD6A49_0(.dout(w_dff_A_XO7BKUc82_0),.din(w_dff_A_uTPbD6A49_0),.clk(gclk));
	jdff dff_A_XO7BKUc82_0(.dout(w_dff_A_oGIhk7Qj5_0),.din(w_dff_A_XO7BKUc82_0),.clk(gclk));
	jdff dff_A_oGIhk7Qj5_0(.dout(w_dff_A_ZGZuUFTI9_0),.din(w_dff_A_oGIhk7Qj5_0),.clk(gclk));
	jdff dff_A_ZGZuUFTI9_0(.dout(w_dff_A_WfTViwob2_0),.din(w_dff_A_ZGZuUFTI9_0),.clk(gclk));
	jdff dff_A_WfTViwob2_0(.dout(w_dff_A_DTvmW2dO8_0),.din(w_dff_A_WfTViwob2_0),.clk(gclk));
	jdff dff_A_DTvmW2dO8_0(.dout(w_dff_A_CPf2djyN7_0),.din(w_dff_A_DTvmW2dO8_0),.clk(gclk));
	jdff dff_A_CPf2djyN7_0(.dout(w_dff_A_V5iusUgI1_0),.din(w_dff_A_CPf2djyN7_0),.clk(gclk));
	jdff dff_A_V5iusUgI1_0(.dout(w_dff_A_pxZ1f6pi0_0),.din(w_dff_A_V5iusUgI1_0),.clk(gclk));
	jdff dff_A_pxZ1f6pi0_0(.dout(w_dff_A_9ICQSLOh2_0),.din(w_dff_A_pxZ1f6pi0_0),.clk(gclk));
	jdff dff_A_9ICQSLOh2_0(.dout(w_dff_A_1sTci4oT5_0),.din(w_dff_A_9ICQSLOh2_0),.clk(gclk));
	jdff dff_A_1sTci4oT5_0(.dout(w_dff_A_ra3nyH0h2_0),.din(w_dff_A_1sTci4oT5_0),.clk(gclk));
	jdff dff_A_ra3nyH0h2_0(.dout(w_dff_A_oyCfNH146_0),.din(w_dff_A_ra3nyH0h2_0),.clk(gclk));
	jdff dff_A_oyCfNH146_0(.dout(w_dff_A_zPiRrCQN5_0),.din(w_dff_A_oyCfNH146_0),.clk(gclk));
	jdff dff_A_zPiRrCQN5_0(.dout(w_dff_A_FsaLbdMq2_0),.din(w_dff_A_zPiRrCQN5_0),.clk(gclk));
	jdff dff_A_FsaLbdMq2_0(.dout(w_dff_A_9lY6IMdd1_0),.din(w_dff_A_FsaLbdMq2_0),.clk(gclk));
	jdff dff_A_9lY6IMdd1_0(.dout(w_dff_A_n6aSC5Pb0_0),.din(w_dff_A_9lY6IMdd1_0),.clk(gclk));
	jdff dff_A_n6aSC5Pb0_0(.dout(w_dff_A_5Y76D0cZ2_0),.din(w_dff_A_n6aSC5Pb0_0),.clk(gclk));
	jdff dff_A_5Y76D0cZ2_0(.dout(G639),.din(w_dff_A_5Y76D0cZ2_0),.clk(gclk));
	jdff dff_A_eXrdnHUC7_2(.dout(w_dff_A_u1sMo46g2_0),.din(w_dff_A_eXrdnHUC7_2),.clk(gclk));
	jdff dff_A_u1sMo46g2_0(.dout(w_dff_A_RJYXGLdr0_0),.din(w_dff_A_u1sMo46g2_0),.clk(gclk));
	jdff dff_A_RJYXGLdr0_0(.dout(w_dff_A_FC7ANpav9_0),.din(w_dff_A_RJYXGLdr0_0),.clk(gclk));
	jdff dff_A_FC7ANpav9_0(.dout(w_dff_A_C4p3N5fD4_0),.din(w_dff_A_FC7ANpav9_0),.clk(gclk));
	jdff dff_A_C4p3N5fD4_0(.dout(w_dff_A_OVkOGZZK8_0),.din(w_dff_A_C4p3N5fD4_0),.clk(gclk));
	jdff dff_A_OVkOGZZK8_0(.dout(w_dff_A_4Xb0k8sk7_0),.din(w_dff_A_OVkOGZZK8_0),.clk(gclk));
	jdff dff_A_4Xb0k8sk7_0(.dout(w_dff_A_y4KY4Ro38_0),.din(w_dff_A_4Xb0k8sk7_0),.clk(gclk));
	jdff dff_A_y4KY4Ro38_0(.dout(w_dff_A_oydTkysa7_0),.din(w_dff_A_y4KY4Ro38_0),.clk(gclk));
	jdff dff_A_oydTkysa7_0(.dout(w_dff_A_1OC6eWBv6_0),.din(w_dff_A_oydTkysa7_0),.clk(gclk));
	jdff dff_A_1OC6eWBv6_0(.dout(w_dff_A_8FBFMwdL0_0),.din(w_dff_A_1OC6eWBv6_0),.clk(gclk));
	jdff dff_A_8FBFMwdL0_0(.dout(w_dff_A_OUrSPaBO9_0),.din(w_dff_A_8FBFMwdL0_0),.clk(gclk));
	jdff dff_A_OUrSPaBO9_0(.dout(w_dff_A_avoKFPxF5_0),.din(w_dff_A_OUrSPaBO9_0),.clk(gclk));
	jdff dff_A_avoKFPxF5_0(.dout(w_dff_A_p3HQEiET6_0),.din(w_dff_A_avoKFPxF5_0),.clk(gclk));
	jdff dff_A_p3HQEiET6_0(.dout(w_dff_A_Y0mOjRHp2_0),.din(w_dff_A_p3HQEiET6_0),.clk(gclk));
	jdff dff_A_Y0mOjRHp2_0(.dout(w_dff_A_xfR59igd6_0),.din(w_dff_A_Y0mOjRHp2_0),.clk(gclk));
	jdff dff_A_xfR59igd6_0(.dout(w_dff_A_Q0dzHYlW1_0),.din(w_dff_A_xfR59igd6_0),.clk(gclk));
	jdff dff_A_Q0dzHYlW1_0(.dout(w_dff_A_LyjDufMW5_0),.din(w_dff_A_Q0dzHYlW1_0),.clk(gclk));
	jdff dff_A_LyjDufMW5_0(.dout(w_dff_A_wM3WlXOf4_0),.din(w_dff_A_LyjDufMW5_0),.clk(gclk));
	jdff dff_A_wM3WlXOf4_0(.dout(w_dff_A_UEQdPovE5_0),.din(w_dff_A_wM3WlXOf4_0),.clk(gclk));
	jdff dff_A_UEQdPovE5_0(.dout(w_dff_A_XYofgA0K5_0),.din(w_dff_A_UEQdPovE5_0),.clk(gclk));
	jdff dff_A_XYofgA0K5_0(.dout(w_dff_A_qIgnYrt85_0),.din(w_dff_A_XYofgA0K5_0),.clk(gclk));
	jdff dff_A_qIgnYrt85_0(.dout(w_dff_A_MVFrvlp67_0),.din(w_dff_A_qIgnYrt85_0),.clk(gclk));
	jdff dff_A_MVFrvlp67_0(.dout(G673),.din(w_dff_A_MVFrvlp67_0),.clk(gclk));
	jdff dff_A_GOXYE6495_2(.dout(w_dff_A_rrgAvDCo1_0),.din(w_dff_A_GOXYE6495_2),.clk(gclk));
	jdff dff_A_rrgAvDCo1_0(.dout(w_dff_A_abmdGtit6_0),.din(w_dff_A_rrgAvDCo1_0),.clk(gclk));
	jdff dff_A_abmdGtit6_0(.dout(w_dff_A_ePLLtNQT8_0),.din(w_dff_A_abmdGtit6_0),.clk(gclk));
	jdff dff_A_ePLLtNQT8_0(.dout(w_dff_A_fiByJLgb2_0),.din(w_dff_A_ePLLtNQT8_0),.clk(gclk));
	jdff dff_A_fiByJLgb2_0(.dout(w_dff_A_1YU481FK8_0),.din(w_dff_A_fiByJLgb2_0),.clk(gclk));
	jdff dff_A_1YU481FK8_0(.dout(w_dff_A_ShF32XcK9_0),.din(w_dff_A_1YU481FK8_0),.clk(gclk));
	jdff dff_A_ShF32XcK9_0(.dout(w_dff_A_5dwbqAYk4_0),.din(w_dff_A_ShF32XcK9_0),.clk(gclk));
	jdff dff_A_5dwbqAYk4_0(.dout(w_dff_A_OypP6riD4_0),.din(w_dff_A_5dwbqAYk4_0),.clk(gclk));
	jdff dff_A_OypP6riD4_0(.dout(w_dff_A_UTTrFT1U0_0),.din(w_dff_A_OypP6riD4_0),.clk(gclk));
	jdff dff_A_UTTrFT1U0_0(.dout(w_dff_A_N3aA6p2m1_0),.din(w_dff_A_UTTrFT1U0_0),.clk(gclk));
	jdff dff_A_N3aA6p2m1_0(.dout(w_dff_A_lvY1EtVy5_0),.din(w_dff_A_N3aA6p2m1_0),.clk(gclk));
	jdff dff_A_lvY1EtVy5_0(.dout(w_dff_A_6o4csVod0_0),.din(w_dff_A_lvY1EtVy5_0),.clk(gclk));
	jdff dff_A_6o4csVod0_0(.dout(w_dff_A_G1GFN9IS1_0),.din(w_dff_A_6o4csVod0_0),.clk(gclk));
	jdff dff_A_G1GFN9IS1_0(.dout(w_dff_A_TIljWDqV9_0),.din(w_dff_A_G1GFN9IS1_0),.clk(gclk));
	jdff dff_A_TIljWDqV9_0(.dout(w_dff_A_fOszQBqM9_0),.din(w_dff_A_TIljWDqV9_0),.clk(gclk));
	jdff dff_A_fOszQBqM9_0(.dout(w_dff_A_peONeGsp4_0),.din(w_dff_A_fOszQBqM9_0),.clk(gclk));
	jdff dff_A_peONeGsp4_0(.dout(w_dff_A_1QSxXp7N7_0),.din(w_dff_A_peONeGsp4_0),.clk(gclk));
	jdff dff_A_1QSxXp7N7_0(.dout(w_dff_A_iXLeS8WU8_0),.din(w_dff_A_1QSxXp7N7_0),.clk(gclk));
	jdff dff_A_iXLeS8WU8_0(.dout(w_dff_A_O8wjXCpb9_0),.din(w_dff_A_iXLeS8WU8_0),.clk(gclk));
	jdff dff_A_O8wjXCpb9_0(.dout(w_dff_A_rFGLQ1Lb2_0),.din(w_dff_A_O8wjXCpb9_0),.clk(gclk));
	jdff dff_A_rFGLQ1Lb2_0(.dout(w_dff_A_bN2Cbh5L4_0),.din(w_dff_A_rFGLQ1Lb2_0),.clk(gclk));
	jdff dff_A_bN2Cbh5L4_0(.dout(w_dff_A_n5YAR0C05_0),.din(w_dff_A_bN2Cbh5L4_0),.clk(gclk));
	jdff dff_A_n5YAR0C05_0(.dout(G707),.din(w_dff_A_n5YAR0C05_0),.clk(gclk));
	jdff dff_A_59IPRAJR0_2(.dout(w_dff_A_pM1DUbWl9_0),.din(w_dff_A_59IPRAJR0_2),.clk(gclk));
	jdff dff_A_pM1DUbWl9_0(.dout(w_dff_A_L8T2dIff8_0),.din(w_dff_A_pM1DUbWl9_0),.clk(gclk));
	jdff dff_A_L8T2dIff8_0(.dout(w_dff_A_BnICfQy90_0),.din(w_dff_A_L8T2dIff8_0),.clk(gclk));
	jdff dff_A_BnICfQy90_0(.dout(w_dff_A_aRN2JmoO8_0),.din(w_dff_A_BnICfQy90_0),.clk(gclk));
	jdff dff_A_aRN2JmoO8_0(.dout(w_dff_A_j54jGt0z4_0),.din(w_dff_A_aRN2JmoO8_0),.clk(gclk));
	jdff dff_A_j54jGt0z4_0(.dout(w_dff_A_zGD3TdRE6_0),.din(w_dff_A_j54jGt0z4_0),.clk(gclk));
	jdff dff_A_zGD3TdRE6_0(.dout(w_dff_A_d6iSFEJg3_0),.din(w_dff_A_zGD3TdRE6_0),.clk(gclk));
	jdff dff_A_d6iSFEJg3_0(.dout(w_dff_A_6Xb0cQX82_0),.din(w_dff_A_d6iSFEJg3_0),.clk(gclk));
	jdff dff_A_6Xb0cQX82_0(.dout(w_dff_A_SqzJMgv70_0),.din(w_dff_A_6Xb0cQX82_0),.clk(gclk));
	jdff dff_A_SqzJMgv70_0(.dout(w_dff_A_MTH5LWoJ7_0),.din(w_dff_A_SqzJMgv70_0),.clk(gclk));
	jdff dff_A_MTH5LWoJ7_0(.dout(w_dff_A_YFehd9rc3_0),.din(w_dff_A_MTH5LWoJ7_0),.clk(gclk));
	jdff dff_A_YFehd9rc3_0(.dout(w_dff_A_q6UiJCbA5_0),.din(w_dff_A_YFehd9rc3_0),.clk(gclk));
	jdff dff_A_q6UiJCbA5_0(.dout(w_dff_A_NLG1sG239_0),.din(w_dff_A_q6UiJCbA5_0),.clk(gclk));
	jdff dff_A_NLG1sG239_0(.dout(w_dff_A_GJNI5DAO8_0),.din(w_dff_A_NLG1sG239_0),.clk(gclk));
	jdff dff_A_GJNI5DAO8_0(.dout(w_dff_A_uz3Te3mx6_0),.din(w_dff_A_GJNI5DAO8_0),.clk(gclk));
	jdff dff_A_uz3Te3mx6_0(.dout(w_dff_A_I9rOEXAD0_0),.din(w_dff_A_uz3Te3mx6_0),.clk(gclk));
	jdff dff_A_I9rOEXAD0_0(.dout(w_dff_A_P8K2jCqv9_0),.din(w_dff_A_I9rOEXAD0_0),.clk(gclk));
	jdff dff_A_P8K2jCqv9_0(.dout(w_dff_A_M0u9Bkms3_0),.din(w_dff_A_P8K2jCqv9_0),.clk(gclk));
	jdff dff_A_M0u9Bkms3_0(.dout(w_dff_A_rLTcttWG4_0),.din(w_dff_A_M0u9Bkms3_0),.clk(gclk));
	jdff dff_A_rLTcttWG4_0(.dout(w_dff_A_hhWKcooo7_0),.din(w_dff_A_rLTcttWG4_0),.clk(gclk));
	jdff dff_A_hhWKcooo7_0(.dout(w_dff_A_dHxLZpSh1_0),.din(w_dff_A_hhWKcooo7_0),.clk(gclk));
	jdff dff_A_dHxLZpSh1_0(.dout(w_dff_A_MqvG8nK23_0),.din(w_dff_A_dHxLZpSh1_0),.clk(gclk));
	jdff dff_A_MqvG8nK23_0(.dout(G715),.din(w_dff_A_MqvG8nK23_0),.clk(gclk));
	jdff dff_A_mkTkpc2K4_2(.dout(w_dff_A_BxVuoL1y7_0),.din(w_dff_A_mkTkpc2K4_2),.clk(gclk));
	jdff dff_A_BxVuoL1y7_0(.dout(w_dff_A_bqeudy5n0_0),.din(w_dff_A_BxVuoL1y7_0),.clk(gclk));
	jdff dff_A_bqeudy5n0_0(.dout(w_dff_A_CdCkLa7D5_0),.din(w_dff_A_bqeudy5n0_0),.clk(gclk));
	jdff dff_A_CdCkLa7D5_0(.dout(w_dff_A_ZsCv6uyj3_0),.din(w_dff_A_CdCkLa7D5_0),.clk(gclk));
	jdff dff_A_ZsCv6uyj3_0(.dout(w_dff_A_1idQKwMK6_0),.din(w_dff_A_ZsCv6uyj3_0),.clk(gclk));
	jdff dff_A_1idQKwMK6_0(.dout(w_dff_A_HzLMPAOj1_0),.din(w_dff_A_1idQKwMK6_0),.clk(gclk));
	jdff dff_A_HzLMPAOj1_0(.dout(w_dff_A_TEuTX86W1_0),.din(w_dff_A_HzLMPAOj1_0),.clk(gclk));
	jdff dff_A_TEuTX86W1_0(.dout(w_dff_A_rBjjsj4U8_0),.din(w_dff_A_TEuTX86W1_0),.clk(gclk));
	jdff dff_A_rBjjsj4U8_0(.dout(w_dff_A_YOusoUNe5_0),.din(w_dff_A_rBjjsj4U8_0),.clk(gclk));
	jdff dff_A_YOusoUNe5_0(.dout(w_dff_A_AfEyve3F0_0),.din(w_dff_A_YOusoUNe5_0),.clk(gclk));
	jdff dff_A_AfEyve3F0_0(.dout(w_dff_A_jHbabJfW1_0),.din(w_dff_A_AfEyve3F0_0),.clk(gclk));
	jdff dff_A_jHbabJfW1_0(.dout(w_dff_A_NwNF5n1l2_0),.din(w_dff_A_jHbabJfW1_0),.clk(gclk));
	jdff dff_A_NwNF5n1l2_0(.dout(w_dff_A_z1a9tGqO4_0),.din(w_dff_A_NwNF5n1l2_0),.clk(gclk));
	jdff dff_A_z1a9tGqO4_0(.dout(w_dff_A_iXv1nSAS2_0),.din(w_dff_A_z1a9tGqO4_0),.clk(gclk));
	jdff dff_A_iXv1nSAS2_0(.dout(w_dff_A_iDc2sWM92_0),.din(w_dff_A_iXv1nSAS2_0),.clk(gclk));
	jdff dff_A_iDc2sWM92_0(.dout(w_dff_A_QowlBAUQ5_0),.din(w_dff_A_iDc2sWM92_0),.clk(gclk));
	jdff dff_A_QowlBAUQ5_0(.dout(w_dff_A_YJBpxGXv4_0),.din(w_dff_A_QowlBAUQ5_0),.clk(gclk));
	jdff dff_A_YJBpxGXv4_0(.dout(w_dff_A_NyZzKhCF1_0),.din(w_dff_A_YJBpxGXv4_0),.clk(gclk));
	jdff dff_A_NyZzKhCF1_0(.dout(w_dff_A_FRdV0Z5a2_0),.din(w_dff_A_NyZzKhCF1_0),.clk(gclk));
	jdff dff_A_FRdV0Z5a2_0(.dout(G598),.din(w_dff_A_FRdV0Z5a2_0),.clk(gclk));
	jdff dff_A_kiJeiQer6_2(.dout(w_dff_A_UoJuqcDo4_0),.din(w_dff_A_kiJeiQer6_2),.clk(gclk));
	jdff dff_A_UoJuqcDo4_0(.dout(w_dff_A_qSCHkV0l4_0),.din(w_dff_A_UoJuqcDo4_0),.clk(gclk));
	jdff dff_A_qSCHkV0l4_0(.dout(w_dff_A_ZImzSTMT4_0),.din(w_dff_A_qSCHkV0l4_0),.clk(gclk));
	jdff dff_A_ZImzSTMT4_0(.dout(w_dff_A_XJWHgbw74_0),.din(w_dff_A_ZImzSTMT4_0),.clk(gclk));
	jdff dff_A_XJWHgbw74_0(.dout(w_dff_A_efk9w5E78_0),.din(w_dff_A_XJWHgbw74_0),.clk(gclk));
	jdff dff_A_efk9w5E78_0(.dout(w_dff_A_vpuqTvCW6_0),.din(w_dff_A_efk9w5E78_0),.clk(gclk));
	jdff dff_A_vpuqTvCW6_0(.dout(w_dff_A_3RPdVmKu5_0),.din(w_dff_A_vpuqTvCW6_0),.clk(gclk));
	jdff dff_A_3RPdVmKu5_0(.dout(w_dff_A_nfN0EqsT1_0),.din(w_dff_A_3RPdVmKu5_0),.clk(gclk));
	jdff dff_A_nfN0EqsT1_0(.dout(w_dff_A_EcRKQ7Eb1_0),.din(w_dff_A_nfN0EqsT1_0),.clk(gclk));
	jdff dff_A_EcRKQ7Eb1_0(.dout(w_dff_A_12o9XDQz3_0),.din(w_dff_A_EcRKQ7Eb1_0),.clk(gclk));
	jdff dff_A_12o9XDQz3_0(.dout(w_dff_A_tIJq6nDZ2_0),.din(w_dff_A_12o9XDQz3_0),.clk(gclk));
	jdff dff_A_tIJq6nDZ2_0(.dout(w_dff_A_3zzxky5u6_0),.din(w_dff_A_tIJq6nDZ2_0),.clk(gclk));
	jdff dff_A_3zzxky5u6_0(.dout(w_dff_A_1iX5lI5n9_0),.din(w_dff_A_3zzxky5u6_0),.clk(gclk));
	jdff dff_A_1iX5lI5n9_0(.dout(w_dff_A_XhDmHjHt3_0),.din(w_dff_A_1iX5lI5n9_0),.clk(gclk));
	jdff dff_A_XhDmHjHt3_0(.dout(w_dff_A_eznnZOei5_0),.din(w_dff_A_XhDmHjHt3_0),.clk(gclk));
	jdff dff_A_eznnZOei5_0(.dout(w_dff_A_wXsQ7jNt0_0),.din(w_dff_A_eznnZOei5_0),.clk(gclk));
	jdff dff_A_wXsQ7jNt0_0(.dout(w_dff_A_4uSpfTKP6_0),.din(w_dff_A_wXsQ7jNt0_0),.clk(gclk));
	jdff dff_A_4uSpfTKP6_0(.dout(w_dff_A_tMcjrITX7_0),.din(w_dff_A_4uSpfTKP6_0),.clk(gclk));
	jdff dff_A_tMcjrITX7_0(.dout(G610),.din(w_dff_A_tMcjrITX7_0),.clk(gclk));
	jdff dff_A_1Y5z3GHA5_2(.dout(w_dff_A_6mKFJZtH4_0),.din(w_dff_A_1Y5z3GHA5_2),.clk(gclk));
	jdff dff_A_6mKFJZtH4_0(.dout(w_dff_A_SClSIx3D4_0),.din(w_dff_A_6mKFJZtH4_0),.clk(gclk));
	jdff dff_A_SClSIx3D4_0(.dout(w_dff_A_mO3TAI7N9_0),.din(w_dff_A_SClSIx3D4_0),.clk(gclk));
	jdff dff_A_mO3TAI7N9_0(.dout(w_dff_A_BsXMaR2q6_0),.din(w_dff_A_mO3TAI7N9_0),.clk(gclk));
	jdff dff_A_BsXMaR2q6_0(.dout(w_dff_A_wyyUYXBi0_0),.din(w_dff_A_BsXMaR2q6_0),.clk(gclk));
	jdff dff_A_wyyUYXBi0_0(.dout(w_dff_A_1K3U7Dog4_0),.din(w_dff_A_wyyUYXBi0_0),.clk(gclk));
	jdff dff_A_1K3U7Dog4_0(.dout(w_dff_A_Zkpdexlu9_0),.din(w_dff_A_1K3U7Dog4_0),.clk(gclk));
	jdff dff_A_Zkpdexlu9_0(.dout(w_dff_A_bgTExiT65_0),.din(w_dff_A_Zkpdexlu9_0),.clk(gclk));
	jdff dff_A_bgTExiT65_0(.dout(w_dff_A_39LV0Tle6_0),.din(w_dff_A_bgTExiT65_0),.clk(gclk));
	jdff dff_A_39LV0Tle6_0(.dout(w_dff_A_YAEenahu5_0),.din(w_dff_A_39LV0Tle6_0),.clk(gclk));
	jdff dff_A_YAEenahu5_0(.dout(w_dff_A_QZqQ3MDU8_0),.din(w_dff_A_YAEenahu5_0),.clk(gclk));
	jdff dff_A_QZqQ3MDU8_0(.dout(w_dff_A_ysQvKkY57_0),.din(w_dff_A_QZqQ3MDU8_0),.clk(gclk));
	jdff dff_A_ysQvKkY57_0(.dout(w_dff_A_Qo3YxnXS4_0),.din(w_dff_A_ysQvKkY57_0),.clk(gclk));
	jdff dff_A_Qo3YxnXS4_0(.dout(w_dff_A_rW1A6dMn7_0),.din(w_dff_A_Qo3YxnXS4_0),.clk(gclk));
	jdff dff_A_rW1A6dMn7_0(.dout(w_dff_A_gtzFmx681_0),.din(w_dff_A_rW1A6dMn7_0),.clk(gclk));
	jdff dff_A_gtzFmx681_0(.dout(w_dff_A_fe9XJN7P3_0),.din(w_dff_A_gtzFmx681_0),.clk(gclk));
	jdff dff_A_fe9XJN7P3_0(.dout(G588),.din(w_dff_A_fe9XJN7P3_0),.clk(gclk));
	jdff dff_A_1RVBZJEC9_2(.dout(w_dff_A_lg3O4dSr0_0),.din(w_dff_A_1RVBZJEC9_2),.clk(gclk));
	jdff dff_A_lg3O4dSr0_0(.dout(w_dff_A_PyMsVnxY7_0),.din(w_dff_A_lg3O4dSr0_0),.clk(gclk));
	jdff dff_A_PyMsVnxY7_0(.dout(w_dff_A_tjNuhyl60_0),.din(w_dff_A_PyMsVnxY7_0),.clk(gclk));
	jdff dff_A_tjNuhyl60_0(.dout(w_dff_A_Bc6Pi9S97_0),.din(w_dff_A_tjNuhyl60_0),.clk(gclk));
	jdff dff_A_Bc6Pi9S97_0(.dout(w_dff_A_DHpRZK6A6_0),.din(w_dff_A_Bc6Pi9S97_0),.clk(gclk));
	jdff dff_A_DHpRZK6A6_0(.dout(w_dff_A_8VtVH8Zc9_0),.din(w_dff_A_DHpRZK6A6_0),.clk(gclk));
	jdff dff_A_8VtVH8Zc9_0(.dout(w_dff_A_tMm9O2NF4_0),.din(w_dff_A_8VtVH8Zc9_0),.clk(gclk));
	jdff dff_A_tMm9O2NF4_0(.dout(w_dff_A_tk5gZflL7_0),.din(w_dff_A_tMm9O2NF4_0),.clk(gclk));
	jdff dff_A_tk5gZflL7_0(.dout(w_dff_A_zMzcfgqZ6_0),.din(w_dff_A_tk5gZflL7_0),.clk(gclk));
	jdff dff_A_zMzcfgqZ6_0(.dout(w_dff_A_g6DLGaA93_0),.din(w_dff_A_zMzcfgqZ6_0),.clk(gclk));
	jdff dff_A_g6DLGaA93_0(.dout(w_dff_A_9zgSJVXK9_0),.din(w_dff_A_g6DLGaA93_0),.clk(gclk));
	jdff dff_A_9zgSJVXK9_0(.dout(w_dff_A_y11EIFcp0_0),.din(w_dff_A_9zgSJVXK9_0),.clk(gclk));
	jdff dff_A_y11EIFcp0_0(.dout(w_dff_A_gW4fRWOh3_0),.din(w_dff_A_y11EIFcp0_0),.clk(gclk));
	jdff dff_A_gW4fRWOh3_0(.dout(w_dff_A_eo7xhwDm5_0),.din(w_dff_A_gW4fRWOh3_0),.clk(gclk));
	jdff dff_A_eo7xhwDm5_0(.dout(w_dff_A_S1PPWCCf4_0),.din(w_dff_A_eo7xhwDm5_0),.clk(gclk));
	jdff dff_A_S1PPWCCf4_0(.dout(w_dff_A_OqjykQxo0_0),.din(w_dff_A_S1PPWCCf4_0),.clk(gclk));
	jdff dff_A_OqjykQxo0_0(.dout(w_dff_A_Ix4GRr790_0),.din(w_dff_A_OqjykQxo0_0),.clk(gclk));
	jdff dff_A_Ix4GRr790_0(.dout(G615),.din(w_dff_A_Ix4GRr790_0),.clk(gclk));
	jdff dff_A_6f5g0anK1_2(.dout(w_dff_A_38CuFKku4_0),.din(w_dff_A_6f5g0anK1_2),.clk(gclk));
	jdff dff_A_38CuFKku4_0(.dout(w_dff_A_SzKK9Fja5_0),.din(w_dff_A_38CuFKku4_0),.clk(gclk));
	jdff dff_A_SzKK9Fja5_0(.dout(w_dff_A_mmkQvEi36_0),.din(w_dff_A_SzKK9Fja5_0),.clk(gclk));
	jdff dff_A_mmkQvEi36_0(.dout(w_dff_A_rqeZYy1E6_0),.din(w_dff_A_mmkQvEi36_0),.clk(gclk));
	jdff dff_A_rqeZYy1E6_0(.dout(w_dff_A_T099VD2t0_0),.din(w_dff_A_rqeZYy1E6_0),.clk(gclk));
	jdff dff_A_T099VD2t0_0(.dout(w_dff_A_TWZOUUEW6_0),.din(w_dff_A_T099VD2t0_0),.clk(gclk));
	jdff dff_A_TWZOUUEW6_0(.dout(w_dff_A_fJZqshVa5_0),.din(w_dff_A_TWZOUUEW6_0),.clk(gclk));
	jdff dff_A_fJZqshVa5_0(.dout(w_dff_A_MwaSSTyt6_0),.din(w_dff_A_fJZqshVa5_0),.clk(gclk));
	jdff dff_A_MwaSSTyt6_0(.dout(w_dff_A_KLBo8KOs1_0),.din(w_dff_A_MwaSSTyt6_0),.clk(gclk));
	jdff dff_A_KLBo8KOs1_0(.dout(w_dff_A_tGUpexzz3_0),.din(w_dff_A_KLBo8KOs1_0),.clk(gclk));
	jdff dff_A_tGUpexzz3_0(.dout(w_dff_A_c8KBWf9d8_0),.din(w_dff_A_tGUpexzz3_0),.clk(gclk));
	jdff dff_A_c8KBWf9d8_0(.dout(w_dff_A_tFSk4fLO9_0),.din(w_dff_A_c8KBWf9d8_0),.clk(gclk));
	jdff dff_A_tFSk4fLO9_0(.dout(w_dff_A_uVeofMBM9_0),.din(w_dff_A_tFSk4fLO9_0),.clk(gclk));
	jdff dff_A_uVeofMBM9_0(.dout(w_dff_A_iJPTT4OC1_0),.din(w_dff_A_uVeofMBM9_0),.clk(gclk));
	jdff dff_A_iJPTT4OC1_0(.dout(w_dff_A_KugvriIB1_0),.din(w_dff_A_iJPTT4OC1_0),.clk(gclk));
	jdff dff_A_KugvriIB1_0(.dout(w_dff_A_NUMpbhzy4_0),.din(w_dff_A_KugvriIB1_0),.clk(gclk));
	jdff dff_A_NUMpbhzy4_0(.dout(w_dff_A_Wdrk0HfE8_0),.din(w_dff_A_NUMpbhzy4_0),.clk(gclk));
	jdff dff_A_Wdrk0HfE8_0(.dout(G626),.din(w_dff_A_Wdrk0HfE8_0),.clk(gclk));
	jdff dff_A_gMde8Pq87_2(.dout(w_dff_A_mUELzTNT7_0),.din(w_dff_A_gMde8Pq87_2),.clk(gclk));
	jdff dff_A_mUELzTNT7_0(.dout(w_dff_A_EEbaj8fe6_0),.din(w_dff_A_mUELzTNT7_0),.clk(gclk));
	jdff dff_A_EEbaj8fe6_0(.dout(w_dff_A_lbS2m6tv1_0),.din(w_dff_A_EEbaj8fe6_0),.clk(gclk));
	jdff dff_A_lbS2m6tv1_0(.dout(w_dff_A_yjByoIOU9_0),.din(w_dff_A_lbS2m6tv1_0),.clk(gclk));
	jdff dff_A_yjByoIOU9_0(.dout(w_dff_A_tmQ5SDGO2_0),.din(w_dff_A_yjByoIOU9_0),.clk(gclk));
	jdff dff_A_tmQ5SDGO2_0(.dout(w_dff_A_M7a6ZIA49_0),.din(w_dff_A_tmQ5SDGO2_0),.clk(gclk));
	jdff dff_A_M7a6ZIA49_0(.dout(w_dff_A_aCwq3sVQ4_0),.din(w_dff_A_M7a6ZIA49_0),.clk(gclk));
	jdff dff_A_aCwq3sVQ4_0(.dout(w_dff_A_6gz6ynCf5_0),.din(w_dff_A_aCwq3sVQ4_0),.clk(gclk));
	jdff dff_A_6gz6ynCf5_0(.dout(w_dff_A_MUyoWCGW4_0),.din(w_dff_A_6gz6ynCf5_0),.clk(gclk));
	jdff dff_A_MUyoWCGW4_0(.dout(w_dff_A_ba10qmmZ2_0),.din(w_dff_A_MUyoWCGW4_0),.clk(gclk));
	jdff dff_A_ba10qmmZ2_0(.dout(w_dff_A_lvd94Pe93_0),.din(w_dff_A_ba10qmmZ2_0),.clk(gclk));
	jdff dff_A_lvd94Pe93_0(.dout(w_dff_A_misKMs3Y2_0),.din(w_dff_A_lvd94Pe93_0),.clk(gclk));
	jdff dff_A_misKMs3Y2_0(.dout(w_dff_A_NYuERfdE4_0),.din(w_dff_A_misKMs3Y2_0),.clk(gclk));
	jdff dff_A_NYuERfdE4_0(.dout(w_dff_A_xm2H86XY3_0),.din(w_dff_A_NYuERfdE4_0),.clk(gclk));
	jdff dff_A_xm2H86XY3_0(.dout(w_dff_A_jdEkR0ve4_0),.din(w_dff_A_xm2H86XY3_0),.clk(gclk));
	jdff dff_A_jdEkR0ve4_0(.dout(w_dff_A_snxzDqXo5_0),.din(w_dff_A_jdEkR0ve4_0),.clk(gclk));
	jdff dff_A_snxzDqXo5_0(.dout(G632),.din(w_dff_A_snxzDqXo5_0),.clk(gclk));
	jdff dff_A_jl9DVvEN6_1(.dout(w_dff_A_zmXuPf7S1_0),.din(w_dff_A_jl9DVvEN6_1),.clk(gclk));
	jdff dff_A_zmXuPf7S1_0(.dout(w_dff_A_B9T7G3PS5_0),.din(w_dff_A_zmXuPf7S1_0),.clk(gclk));
	jdff dff_A_B9T7G3PS5_0(.dout(w_dff_A_eiicRrsq4_0),.din(w_dff_A_B9T7G3PS5_0),.clk(gclk));
	jdff dff_A_eiicRrsq4_0(.dout(w_dff_A_AXlfZhwq4_0),.din(w_dff_A_eiicRrsq4_0),.clk(gclk));
	jdff dff_A_AXlfZhwq4_0(.dout(w_dff_A_vUYvSS6t9_0),.din(w_dff_A_AXlfZhwq4_0),.clk(gclk));
	jdff dff_A_vUYvSS6t9_0(.dout(w_dff_A_xD0wl7nN6_0),.din(w_dff_A_vUYvSS6t9_0),.clk(gclk));
	jdff dff_A_xD0wl7nN6_0(.dout(w_dff_A_jluNa5RS8_0),.din(w_dff_A_xD0wl7nN6_0),.clk(gclk));
	jdff dff_A_jluNa5RS8_0(.dout(w_dff_A_6WXl4seo8_0),.din(w_dff_A_jluNa5RS8_0),.clk(gclk));
	jdff dff_A_6WXl4seo8_0(.dout(w_dff_A_TIM5BsFK4_0),.din(w_dff_A_6WXl4seo8_0),.clk(gclk));
	jdff dff_A_TIM5BsFK4_0(.dout(w_dff_A_lu6Xl9b30_0),.din(w_dff_A_TIM5BsFK4_0),.clk(gclk));
	jdff dff_A_lu6Xl9b30_0(.dout(w_dff_A_ddVIOdPE8_0),.din(w_dff_A_lu6Xl9b30_0),.clk(gclk));
	jdff dff_A_ddVIOdPE8_0(.dout(w_dff_A_oZ1LAy2l3_0),.din(w_dff_A_ddVIOdPE8_0),.clk(gclk));
	jdff dff_A_oZ1LAy2l3_0(.dout(w_dff_A_NxvexjAB3_0),.din(w_dff_A_oZ1LAy2l3_0),.clk(gclk));
	jdff dff_A_NxvexjAB3_0(.dout(w_dff_A_2Dx8xmxM2_0),.din(w_dff_A_NxvexjAB3_0),.clk(gclk));
	jdff dff_A_2Dx8xmxM2_0(.dout(w_dff_A_OLFFV1fO6_0),.din(w_dff_A_2Dx8xmxM2_0),.clk(gclk));
	jdff dff_A_OLFFV1fO6_0(.dout(w_dff_A_MagLAuyn3_0),.din(w_dff_A_OLFFV1fO6_0),.clk(gclk));
	jdff dff_A_MagLAuyn3_0(.dout(w_dff_A_i04Fd4Iv1_0),.din(w_dff_A_MagLAuyn3_0),.clk(gclk));
	jdff dff_A_i04Fd4Iv1_0(.dout(w_dff_A_hFhS8SEb8_0),.din(w_dff_A_i04Fd4Iv1_0),.clk(gclk));
	jdff dff_A_hFhS8SEb8_0(.dout(w_dff_A_vMBXWVcX1_0),.din(w_dff_A_hFhS8SEb8_0),.clk(gclk));
	jdff dff_A_vMBXWVcX1_0(.dout(w_dff_A_sw7Bi2oV4_0),.din(w_dff_A_vMBXWVcX1_0),.clk(gclk));
	jdff dff_A_sw7Bi2oV4_0(.dout(w_dff_A_vYiPlc5d7_0),.din(w_dff_A_sw7Bi2oV4_0),.clk(gclk));
	jdff dff_A_vYiPlc5d7_0(.dout(w_dff_A_YqVRDqit3_0),.din(w_dff_A_vYiPlc5d7_0),.clk(gclk));
	jdff dff_A_YqVRDqit3_0(.dout(G1002),.din(w_dff_A_YqVRDqit3_0),.clk(gclk));
	jdff dff_A_9BfOiUdX0_1(.dout(w_dff_A_svXeqnba4_0),.din(w_dff_A_9BfOiUdX0_1),.clk(gclk));
	jdff dff_A_svXeqnba4_0(.dout(w_dff_A_XsK7Yd838_0),.din(w_dff_A_svXeqnba4_0),.clk(gclk));
	jdff dff_A_XsK7Yd838_0(.dout(w_dff_A_pexPtVeX2_0),.din(w_dff_A_XsK7Yd838_0),.clk(gclk));
	jdff dff_A_pexPtVeX2_0(.dout(w_dff_A_Bz761Y1V6_0),.din(w_dff_A_pexPtVeX2_0),.clk(gclk));
	jdff dff_A_Bz761Y1V6_0(.dout(w_dff_A_0nTzUGia5_0),.din(w_dff_A_Bz761Y1V6_0),.clk(gclk));
	jdff dff_A_0nTzUGia5_0(.dout(w_dff_A_Z34NABgk1_0),.din(w_dff_A_0nTzUGia5_0),.clk(gclk));
	jdff dff_A_Z34NABgk1_0(.dout(w_dff_A_20tJYRad7_0),.din(w_dff_A_Z34NABgk1_0),.clk(gclk));
	jdff dff_A_20tJYRad7_0(.dout(w_dff_A_ghTPUouy1_0),.din(w_dff_A_20tJYRad7_0),.clk(gclk));
	jdff dff_A_ghTPUouy1_0(.dout(w_dff_A_iOmxQnJb5_0),.din(w_dff_A_ghTPUouy1_0),.clk(gclk));
	jdff dff_A_iOmxQnJb5_0(.dout(w_dff_A_Vnydl0Od7_0),.din(w_dff_A_iOmxQnJb5_0),.clk(gclk));
	jdff dff_A_Vnydl0Od7_0(.dout(w_dff_A_bmTpO0vX7_0),.din(w_dff_A_Vnydl0Od7_0),.clk(gclk));
	jdff dff_A_bmTpO0vX7_0(.dout(w_dff_A_mfa69Sig2_0),.din(w_dff_A_bmTpO0vX7_0),.clk(gclk));
	jdff dff_A_mfa69Sig2_0(.dout(w_dff_A_EUFshqh56_0),.din(w_dff_A_mfa69Sig2_0),.clk(gclk));
	jdff dff_A_EUFshqh56_0(.dout(w_dff_A_7VTg7RxP4_0),.din(w_dff_A_EUFshqh56_0),.clk(gclk));
	jdff dff_A_7VTg7RxP4_0(.dout(w_dff_A_gv9A0ZLZ1_0),.din(w_dff_A_7VTg7RxP4_0),.clk(gclk));
	jdff dff_A_gv9A0ZLZ1_0(.dout(w_dff_A_3Yth2iJE9_0),.din(w_dff_A_gv9A0ZLZ1_0),.clk(gclk));
	jdff dff_A_3Yth2iJE9_0(.dout(w_dff_A_c9c0t3Hh7_0),.din(w_dff_A_3Yth2iJE9_0),.clk(gclk));
	jdff dff_A_c9c0t3Hh7_0(.dout(w_dff_A_D9F6MfN13_0),.din(w_dff_A_c9c0t3Hh7_0),.clk(gclk));
	jdff dff_A_D9F6MfN13_0(.dout(w_dff_A_VFbQQQC16_0),.din(w_dff_A_D9F6MfN13_0),.clk(gclk));
	jdff dff_A_VFbQQQC16_0(.dout(w_dff_A_PDpvrrDB6_0),.din(w_dff_A_VFbQQQC16_0),.clk(gclk));
	jdff dff_A_PDpvrrDB6_0(.dout(w_dff_A_iUwMaq9k0_0),.din(w_dff_A_PDpvrrDB6_0),.clk(gclk));
	jdff dff_A_iUwMaq9k0_0(.dout(w_dff_A_nNBaGDLA8_0),.din(w_dff_A_iUwMaq9k0_0),.clk(gclk));
	jdff dff_A_nNBaGDLA8_0(.dout(G1004),.din(w_dff_A_nNBaGDLA8_0),.clk(gclk));
	jdff dff_A_SAvAS5ac4_2(.dout(w_dff_A_0ZmKSFZq0_0),.din(w_dff_A_SAvAS5ac4_2),.clk(gclk));
	jdff dff_A_0ZmKSFZq0_0(.dout(w_dff_A_Su4B4ZxA6_0),.din(w_dff_A_0ZmKSFZq0_0),.clk(gclk));
	jdff dff_A_Su4B4ZxA6_0(.dout(w_dff_A_tEpm2T1x9_0),.din(w_dff_A_Su4B4ZxA6_0),.clk(gclk));
	jdff dff_A_tEpm2T1x9_0(.dout(w_dff_A_yaQLeFVI3_0),.din(w_dff_A_tEpm2T1x9_0),.clk(gclk));
	jdff dff_A_yaQLeFVI3_0(.dout(w_dff_A_SgJ4JHkq2_0),.din(w_dff_A_yaQLeFVI3_0),.clk(gclk));
	jdff dff_A_SgJ4JHkq2_0(.dout(w_dff_A_qmvuXtsa6_0),.din(w_dff_A_SgJ4JHkq2_0),.clk(gclk));
	jdff dff_A_qmvuXtsa6_0(.dout(w_dff_A_uAOCnff88_0),.din(w_dff_A_qmvuXtsa6_0),.clk(gclk));
	jdff dff_A_uAOCnff88_0(.dout(w_dff_A_e7AYugUu0_0),.din(w_dff_A_uAOCnff88_0),.clk(gclk));
	jdff dff_A_e7AYugUu0_0(.dout(w_dff_A_bELKA3yD0_0),.din(w_dff_A_e7AYugUu0_0),.clk(gclk));
	jdff dff_A_bELKA3yD0_0(.dout(w_dff_A_xYqzNEyw7_0),.din(w_dff_A_bELKA3yD0_0),.clk(gclk));
	jdff dff_A_xYqzNEyw7_0(.dout(w_dff_A_LqrRWkdQ1_0),.din(w_dff_A_xYqzNEyw7_0),.clk(gclk));
	jdff dff_A_LqrRWkdQ1_0(.dout(w_dff_A_v4tDnsaq1_0),.din(w_dff_A_LqrRWkdQ1_0),.clk(gclk));
	jdff dff_A_v4tDnsaq1_0(.dout(w_dff_A_1lamenRD4_0),.din(w_dff_A_v4tDnsaq1_0),.clk(gclk));
	jdff dff_A_1lamenRD4_0(.dout(G591),.din(w_dff_A_1lamenRD4_0),.clk(gclk));
	jdff dff_A_GkJoW1s90_2(.dout(w_dff_A_kHHxi3Eg5_0),.din(w_dff_A_GkJoW1s90_2),.clk(gclk));
	jdff dff_A_kHHxi3Eg5_0(.dout(w_dff_A_tWAHHwad8_0),.din(w_dff_A_kHHxi3Eg5_0),.clk(gclk));
	jdff dff_A_tWAHHwad8_0(.dout(w_dff_A_yRaoE6ub6_0),.din(w_dff_A_tWAHHwad8_0),.clk(gclk));
	jdff dff_A_yRaoE6ub6_0(.dout(w_dff_A_QSB2vzVF0_0),.din(w_dff_A_yRaoE6ub6_0),.clk(gclk));
	jdff dff_A_QSB2vzVF0_0(.dout(w_dff_A_CR2oVjbp0_0),.din(w_dff_A_QSB2vzVF0_0),.clk(gclk));
	jdff dff_A_CR2oVjbp0_0(.dout(w_dff_A_pqyknbbY7_0),.din(w_dff_A_CR2oVjbp0_0),.clk(gclk));
	jdff dff_A_pqyknbbY7_0(.dout(w_dff_A_AMzYwiJV6_0),.din(w_dff_A_pqyknbbY7_0),.clk(gclk));
	jdff dff_A_AMzYwiJV6_0(.dout(w_dff_A_RnIMg0oD0_0),.din(w_dff_A_AMzYwiJV6_0),.clk(gclk));
	jdff dff_A_RnIMg0oD0_0(.dout(w_dff_A_95iPqvg70_0),.din(w_dff_A_RnIMg0oD0_0),.clk(gclk));
	jdff dff_A_95iPqvg70_0(.dout(w_dff_A_zNjTUnoR9_0),.din(w_dff_A_95iPqvg70_0),.clk(gclk));
	jdff dff_A_zNjTUnoR9_0(.dout(w_dff_A_vrUoWyx38_0),.din(w_dff_A_zNjTUnoR9_0),.clk(gclk));
	jdff dff_A_vrUoWyx38_0(.dout(w_dff_A_r8nApT5A3_0),.din(w_dff_A_vrUoWyx38_0),.clk(gclk));
	jdff dff_A_r8nApT5A3_0(.dout(w_dff_A_Np0KkK0m3_0),.din(w_dff_A_r8nApT5A3_0),.clk(gclk));
	jdff dff_A_Np0KkK0m3_0(.dout(w_dff_A_lGedkKfI9_0),.din(w_dff_A_Np0KkK0m3_0),.clk(gclk));
	jdff dff_A_lGedkKfI9_0(.dout(G618),.din(w_dff_A_lGedkKfI9_0),.clk(gclk));
	jdff dff_A_SEr1vClL9_2(.dout(w_dff_A_lD8JTnvG5_0),.din(w_dff_A_SEr1vClL9_2),.clk(gclk));
	jdff dff_A_lD8JTnvG5_0(.dout(w_dff_A_sCHPlANe3_0),.din(w_dff_A_lD8JTnvG5_0),.clk(gclk));
	jdff dff_A_sCHPlANe3_0(.dout(w_dff_A_iYkt8Cqv1_0),.din(w_dff_A_sCHPlANe3_0),.clk(gclk));
	jdff dff_A_iYkt8Cqv1_0(.dout(w_dff_A_cMRybDRq1_0),.din(w_dff_A_iYkt8Cqv1_0),.clk(gclk));
	jdff dff_A_cMRybDRq1_0(.dout(w_dff_A_2X7E52Sn6_0),.din(w_dff_A_cMRybDRq1_0),.clk(gclk));
	jdff dff_A_2X7E52Sn6_0(.dout(w_dff_A_a0qmWvzK5_0),.din(w_dff_A_2X7E52Sn6_0),.clk(gclk));
	jdff dff_A_a0qmWvzK5_0(.dout(w_dff_A_mbANAgzG8_0),.din(w_dff_A_a0qmWvzK5_0),.clk(gclk));
	jdff dff_A_mbANAgzG8_0(.dout(w_dff_A_ICFyReGj3_0),.din(w_dff_A_mbANAgzG8_0),.clk(gclk));
	jdff dff_A_ICFyReGj3_0(.dout(w_dff_A_rsWZvl7p4_0),.din(w_dff_A_ICFyReGj3_0),.clk(gclk));
	jdff dff_A_rsWZvl7p4_0(.dout(w_dff_A_1obtUJJx0_0),.din(w_dff_A_rsWZvl7p4_0),.clk(gclk));
	jdff dff_A_1obtUJJx0_0(.dout(w_dff_A_UyrFTC8R9_0),.din(w_dff_A_1obtUJJx0_0),.clk(gclk));
	jdff dff_A_UyrFTC8R9_0(.dout(w_dff_A_egFEADV73_0),.din(w_dff_A_UyrFTC8R9_0),.clk(gclk));
	jdff dff_A_egFEADV73_0(.dout(w_dff_A_tWd3LFVg6_0),.din(w_dff_A_egFEADV73_0),.clk(gclk));
	jdff dff_A_tWd3LFVg6_0(.dout(G621),.din(w_dff_A_tWd3LFVg6_0),.clk(gclk));
	jdff dff_A_FP0rTFvM2_2(.dout(w_dff_A_FCe3qd0e1_0),.din(w_dff_A_FP0rTFvM2_2),.clk(gclk));
	jdff dff_A_FCe3qd0e1_0(.dout(w_dff_A_eRd5USvR9_0),.din(w_dff_A_FCe3qd0e1_0),.clk(gclk));
	jdff dff_A_eRd5USvR9_0(.dout(w_dff_A_E8eSqdeW2_0),.din(w_dff_A_eRd5USvR9_0),.clk(gclk));
	jdff dff_A_E8eSqdeW2_0(.dout(w_dff_A_kGiw5Vi43_0),.din(w_dff_A_E8eSqdeW2_0),.clk(gclk));
	jdff dff_A_kGiw5Vi43_0(.dout(w_dff_A_Gh4X3QHl7_0),.din(w_dff_A_kGiw5Vi43_0),.clk(gclk));
	jdff dff_A_Gh4X3QHl7_0(.dout(w_dff_A_ZzrmXXHP1_0),.din(w_dff_A_Gh4X3QHl7_0),.clk(gclk));
	jdff dff_A_ZzrmXXHP1_0(.dout(w_dff_A_uBmhPkcc7_0),.din(w_dff_A_ZzrmXXHP1_0),.clk(gclk));
	jdff dff_A_uBmhPkcc7_0(.dout(w_dff_A_PgWNlTPo2_0),.din(w_dff_A_uBmhPkcc7_0),.clk(gclk));
	jdff dff_A_PgWNlTPo2_0(.dout(w_dff_A_ik9mDEgu2_0),.din(w_dff_A_PgWNlTPo2_0),.clk(gclk));
	jdff dff_A_ik9mDEgu2_0(.dout(w_dff_A_AZEL8e0W7_0),.din(w_dff_A_ik9mDEgu2_0),.clk(gclk));
	jdff dff_A_AZEL8e0W7_0(.dout(w_dff_A_SQfEEdu85_0),.din(w_dff_A_AZEL8e0W7_0),.clk(gclk));
	jdff dff_A_SQfEEdu85_0(.dout(w_dff_A_0UCpNHT47_0),.din(w_dff_A_SQfEEdu85_0),.clk(gclk));
	jdff dff_A_0UCpNHT47_0(.dout(w_dff_A_rfYQQaAQ3_0),.din(w_dff_A_0UCpNHT47_0),.clk(gclk));
	jdff dff_A_rfYQQaAQ3_0(.dout(w_dff_A_y6aTy7GM3_0),.din(w_dff_A_rfYQQaAQ3_0),.clk(gclk));
	jdff dff_A_y6aTy7GM3_0(.dout(G629),.din(w_dff_A_y6aTy7GM3_0),.clk(gclk));
	jdff dff_A_VYShTGcq8_1(.dout(w_dff_A_xyW8xbEx9_0),.din(w_dff_A_VYShTGcq8_1),.clk(gclk));
	jdff dff_A_xyW8xbEx9_0(.dout(w_dff_A_WCff8LI80_0),.din(w_dff_A_xyW8xbEx9_0),.clk(gclk));
	jdff dff_A_WCff8LI80_0(.dout(w_dff_A_Fw1PBLGG1_0),.din(w_dff_A_WCff8LI80_0),.clk(gclk));
	jdff dff_A_Fw1PBLGG1_0(.dout(w_dff_A_40glEXYn3_0),.din(w_dff_A_Fw1PBLGG1_0),.clk(gclk));
	jdff dff_A_40glEXYn3_0(.dout(w_dff_A_EUyf9Bfa4_0),.din(w_dff_A_40glEXYn3_0),.clk(gclk));
	jdff dff_A_EUyf9Bfa4_0(.dout(w_dff_A_4EGNw5dr6_0),.din(w_dff_A_EUyf9Bfa4_0),.clk(gclk));
	jdff dff_A_4EGNw5dr6_0(.dout(w_dff_A_7n38dQYW1_0),.din(w_dff_A_4EGNw5dr6_0),.clk(gclk));
	jdff dff_A_7n38dQYW1_0(.dout(w_dff_A_xxKOFpVR4_0),.din(w_dff_A_7n38dQYW1_0),.clk(gclk));
	jdff dff_A_xxKOFpVR4_0(.dout(w_dff_A_K0lIoeYy9_0),.din(w_dff_A_xxKOFpVR4_0),.clk(gclk));
	jdff dff_A_K0lIoeYy9_0(.dout(w_dff_A_IWT87sXT8_0),.din(w_dff_A_K0lIoeYy9_0),.clk(gclk));
	jdff dff_A_IWT87sXT8_0(.dout(w_dff_A_nKDkwGaY3_0),.din(w_dff_A_IWT87sXT8_0),.clk(gclk));
	jdff dff_A_nKDkwGaY3_0(.dout(w_dff_A_zCMl7dFs7_0),.din(w_dff_A_nKDkwGaY3_0),.clk(gclk));
	jdff dff_A_zCMl7dFs7_0(.dout(w_dff_A_OC11v3q14_0),.din(w_dff_A_zCMl7dFs7_0),.clk(gclk));
	jdff dff_A_OC11v3q14_0(.dout(w_dff_A_Jr3knpH14_0),.din(w_dff_A_OC11v3q14_0),.clk(gclk));
	jdff dff_A_Jr3knpH14_0(.dout(w_dff_A_uiFkqbSb7_0),.din(w_dff_A_Jr3knpH14_0),.clk(gclk));
	jdff dff_A_uiFkqbSb7_0(.dout(w_dff_A_e8F93ljk0_0),.din(w_dff_A_uiFkqbSb7_0),.clk(gclk));
	jdff dff_A_e8F93ljk0_0(.dout(w_dff_A_OdXzH4895_0),.din(w_dff_A_e8F93ljk0_0),.clk(gclk));
	jdff dff_A_OdXzH4895_0(.dout(w_dff_A_bMx2MXwA4_0),.din(w_dff_A_OdXzH4895_0),.clk(gclk));
	jdff dff_A_bMx2MXwA4_0(.dout(w_dff_A_GsjzM8tQ4_0),.din(w_dff_A_bMx2MXwA4_0),.clk(gclk));
	jdff dff_A_GsjzM8tQ4_0(.dout(G822),.din(w_dff_A_GsjzM8tQ4_0),.clk(gclk));
	jdff dff_A_UAv8zeNK0_1(.dout(w_dff_A_ls6mhGSr5_0),.din(w_dff_A_UAv8zeNK0_1),.clk(gclk));
	jdff dff_A_ls6mhGSr5_0(.dout(w_dff_A_4ocDkuqr3_0),.din(w_dff_A_ls6mhGSr5_0),.clk(gclk));
	jdff dff_A_4ocDkuqr3_0(.dout(w_dff_A_bUbhWxaa5_0),.din(w_dff_A_4ocDkuqr3_0),.clk(gclk));
	jdff dff_A_bUbhWxaa5_0(.dout(w_dff_A_ESFZwOak5_0),.din(w_dff_A_bUbhWxaa5_0),.clk(gclk));
	jdff dff_A_ESFZwOak5_0(.dout(w_dff_A_evMm0Wyl8_0),.din(w_dff_A_ESFZwOak5_0),.clk(gclk));
	jdff dff_A_evMm0Wyl8_0(.dout(w_dff_A_cqcqpeiv9_0),.din(w_dff_A_evMm0Wyl8_0),.clk(gclk));
	jdff dff_A_cqcqpeiv9_0(.dout(w_dff_A_3dtCgJOa6_0),.din(w_dff_A_cqcqpeiv9_0),.clk(gclk));
	jdff dff_A_3dtCgJOa6_0(.dout(w_dff_A_hLjg8dKo5_0),.din(w_dff_A_3dtCgJOa6_0),.clk(gclk));
	jdff dff_A_hLjg8dKo5_0(.dout(w_dff_A_xFTgryao0_0),.din(w_dff_A_hLjg8dKo5_0),.clk(gclk));
	jdff dff_A_xFTgryao0_0(.dout(w_dff_A_htkS74VD0_0),.din(w_dff_A_xFTgryao0_0),.clk(gclk));
	jdff dff_A_htkS74VD0_0(.dout(w_dff_A_RvdXaJ2C8_0),.din(w_dff_A_htkS74VD0_0),.clk(gclk));
	jdff dff_A_RvdXaJ2C8_0(.dout(w_dff_A_fNsojorH1_0),.din(w_dff_A_RvdXaJ2C8_0),.clk(gclk));
	jdff dff_A_fNsojorH1_0(.dout(w_dff_A_zjiM5xx56_0),.din(w_dff_A_fNsojorH1_0),.clk(gclk));
	jdff dff_A_zjiM5xx56_0(.dout(w_dff_A_nRxtJe0P7_0),.din(w_dff_A_zjiM5xx56_0),.clk(gclk));
	jdff dff_A_nRxtJe0P7_0(.dout(G838),.din(w_dff_A_nRxtJe0P7_0),.clk(gclk));
	jdff dff_A_IgwmqSnl4_1(.dout(w_dff_A_CVw9f9ZQ0_0),.din(w_dff_A_IgwmqSnl4_1),.clk(gclk));
	jdff dff_A_CVw9f9ZQ0_0(.dout(w_dff_A_kgvT1LDn1_0),.din(w_dff_A_CVw9f9ZQ0_0),.clk(gclk));
	jdff dff_A_kgvT1LDn1_0(.dout(w_dff_A_QsJHV1aW7_0),.din(w_dff_A_kgvT1LDn1_0),.clk(gclk));
	jdff dff_A_QsJHV1aW7_0(.dout(w_dff_A_aWkJYRAU2_0),.din(w_dff_A_QsJHV1aW7_0),.clk(gclk));
	jdff dff_A_aWkJYRAU2_0(.dout(w_dff_A_eC2gi2Dt8_0),.din(w_dff_A_aWkJYRAU2_0),.clk(gclk));
	jdff dff_A_eC2gi2Dt8_0(.dout(w_dff_A_s59l3sbf2_0),.din(w_dff_A_eC2gi2Dt8_0),.clk(gclk));
	jdff dff_A_s59l3sbf2_0(.dout(w_dff_A_DRdD1hxp6_0),.din(w_dff_A_s59l3sbf2_0),.clk(gclk));
	jdff dff_A_DRdD1hxp6_0(.dout(w_dff_A_6XBHXxyY9_0),.din(w_dff_A_DRdD1hxp6_0),.clk(gclk));
	jdff dff_A_6XBHXxyY9_0(.dout(w_dff_A_zWnInFWt9_0),.din(w_dff_A_6XBHXxyY9_0),.clk(gclk));
	jdff dff_A_zWnInFWt9_0(.dout(w_dff_A_cJmTzp6k2_0),.din(w_dff_A_zWnInFWt9_0),.clk(gclk));
	jdff dff_A_cJmTzp6k2_0(.dout(w_dff_A_v9fxuwNP4_0),.din(w_dff_A_cJmTzp6k2_0),.clk(gclk));
	jdff dff_A_v9fxuwNP4_0(.dout(w_dff_A_TagAa3n83_0),.din(w_dff_A_v9fxuwNP4_0),.clk(gclk));
	jdff dff_A_TagAa3n83_0(.dout(w_dff_A_texKzv0j4_0),.din(w_dff_A_TagAa3n83_0),.clk(gclk));
	jdff dff_A_texKzv0j4_0(.dout(w_dff_A_jsGW8a3P6_0),.din(w_dff_A_texKzv0j4_0),.clk(gclk));
	jdff dff_A_jsGW8a3P6_0(.dout(w_dff_A_rRSyD1XI1_0),.din(w_dff_A_jsGW8a3P6_0),.clk(gclk));
	jdff dff_A_rRSyD1XI1_0(.dout(w_dff_A_K4sjGOlI5_0),.din(w_dff_A_rRSyD1XI1_0),.clk(gclk));
	jdff dff_A_K4sjGOlI5_0(.dout(w_dff_A_elshjJ2a6_0),.din(w_dff_A_K4sjGOlI5_0),.clk(gclk));
	jdff dff_A_elshjJ2a6_0(.dout(G861),.din(w_dff_A_elshjJ2a6_0),.clk(gclk));
	jdff dff_A_b7Uj8T3n5_1(.dout(w_dff_A_Q5Bl4VHM5_0),.din(w_dff_A_b7Uj8T3n5_1),.clk(gclk));
	jdff dff_A_Q5Bl4VHM5_0(.dout(w_dff_A_F6Fyb4PK9_0),.din(w_dff_A_Q5Bl4VHM5_0),.clk(gclk));
	jdff dff_A_F6Fyb4PK9_0(.dout(w_dff_A_ORhDGbi24_0),.din(w_dff_A_F6Fyb4PK9_0),.clk(gclk));
	jdff dff_A_ORhDGbi24_0(.dout(w_dff_A_yIg9xb0S5_0),.din(w_dff_A_ORhDGbi24_0),.clk(gclk));
	jdff dff_A_yIg9xb0S5_0(.dout(w_dff_A_VuKjo45b0_0),.din(w_dff_A_yIg9xb0S5_0),.clk(gclk));
	jdff dff_A_VuKjo45b0_0(.dout(w_dff_A_aFvmcpgY1_0),.din(w_dff_A_VuKjo45b0_0),.clk(gclk));
	jdff dff_A_aFvmcpgY1_0(.dout(w_dff_A_RrmLO3lS0_0),.din(w_dff_A_aFvmcpgY1_0),.clk(gclk));
	jdff dff_A_RrmLO3lS0_0(.dout(w_dff_A_FbwFgVBz2_0),.din(w_dff_A_RrmLO3lS0_0),.clk(gclk));
	jdff dff_A_FbwFgVBz2_0(.dout(w_dff_A_B8YhUJlE8_0),.din(w_dff_A_FbwFgVBz2_0),.clk(gclk));
	jdff dff_A_B8YhUJlE8_0(.dout(G623),.din(w_dff_A_B8YhUJlE8_0),.clk(gclk));
	jdff dff_A_O7wYAVdt7_2(.dout(w_dff_A_cJ1xjnVx9_0),.din(w_dff_A_O7wYAVdt7_2),.clk(gclk));
	jdff dff_A_cJ1xjnVx9_0(.dout(w_dff_A_O5aBwdkq7_0),.din(w_dff_A_cJ1xjnVx9_0),.clk(gclk));
	jdff dff_A_O5aBwdkq7_0(.dout(w_dff_A_MUpUZpCL0_0),.din(w_dff_A_O5aBwdkq7_0),.clk(gclk));
	jdff dff_A_MUpUZpCL0_0(.dout(w_dff_A_melqquDJ0_0),.din(w_dff_A_MUpUZpCL0_0),.clk(gclk));
	jdff dff_A_melqquDJ0_0(.dout(w_dff_A_k0NN3Ywp3_0),.din(w_dff_A_melqquDJ0_0),.clk(gclk));
	jdff dff_A_k0NN3Ywp3_0(.dout(w_dff_A_G7tl7YLo8_0),.din(w_dff_A_k0NN3Ywp3_0),.clk(gclk));
	jdff dff_A_G7tl7YLo8_0(.dout(w_dff_A_Bkgeuktz1_0),.din(w_dff_A_G7tl7YLo8_0),.clk(gclk));
	jdff dff_A_Bkgeuktz1_0(.dout(w_dff_A_t2lJX0nL8_0),.din(w_dff_A_Bkgeuktz1_0),.clk(gclk));
	jdff dff_A_t2lJX0nL8_0(.dout(w_dff_A_dKmiRRz30_0),.din(w_dff_A_t2lJX0nL8_0),.clk(gclk));
	jdff dff_A_dKmiRRz30_0(.dout(w_dff_A_6SCb69Xz2_0),.din(w_dff_A_dKmiRRz30_0),.clk(gclk));
	jdff dff_A_6SCb69Xz2_0(.dout(w_dff_A_Ryq8wyXX4_0),.din(w_dff_A_6SCb69Xz2_0),.clk(gclk));
	jdff dff_A_Ryq8wyXX4_0(.dout(w_dff_A_UNqPTvZZ1_0),.din(w_dff_A_Ryq8wyXX4_0),.clk(gclk));
	jdff dff_A_UNqPTvZZ1_0(.dout(w_dff_A_8AKhhv408_0),.din(w_dff_A_UNqPTvZZ1_0),.clk(gclk));
	jdff dff_A_8AKhhv408_0(.dout(G722),.din(w_dff_A_8AKhhv408_0),.clk(gclk));
	jdff dff_A_TjtWKR5k2_1(.dout(w_dff_A_6O1ncbqr8_0),.din(w_dff_A_TjtWKR5k2_1),.clk(gclk));
	jdff dff_A_6O1ncbqr8_0(.dout(w_dff_A_Z8S8p4Et6_0),.din(w_dff_A_6O1ncbqr8_0),.clk(gclk));
	jdff dff_A_Z8S8p4Et6_0(.dout(w_dff_A_C8sX4F7e2_0),.din(w_dff_A_Z8S8p4Et6_0),.clk(gclk));
	jdff dff_A_C8sX4F7e2_0(.dout(w_dff_A_AbcY5CPb6_0),.din(w_dff_A_C8sX4F7e2_0),.clk(gclk));
	jdff dff_A_AbcY5CPb6_0(.dout(w_dff_A_cXmOX0607_0),.din(w_dff_A_AbcY5CPb6_0),.clk(gclk));
	jdff dff_A_cXmOX0607_0(.dout(w_dff_A_1mje5fvU4_0),.din(w_dff_A_cXmOX0607_0),.clk(gclk));
	jdff dff_A_1mje5fvU4_0(.dout(w_dff_A_7OsreSFE6_0),.din(w_dff_A_1mje5fvU4_0),.clk(gclk));
	jdff dff_A_7OsreSFE6_0(.dout(w_dff_A_DG1LGQhe9_0),.din(w_dff_A_7OsreSFE6_0),.clk(gclk));
	jdff dff_A_DG1LGQhe9_0(.dout(w_dff_A_4jxs10DW8_0),.din(w_dff_A_DG1LGQhe9_0),.clk(gclk));
	jdff dff_A_4jxs10DW8_0(.dout(w_dff_A_EKGmmqRE8_0),.din(w_dff_A_4jxs10DW8_0),.clk(gclk));
	jdff dff_A_EKGmmqRE8_0(.dout(w_dff_A_H3Ie7GYo3_0),.din(w_dff_A_EKGmmqRE8_0),.clk(gclk));
	jdff dff_A_H3Ie7GYo3_0(.dout(w_dff_A_5v8gAEv80_0),.din(w_dff_A_H3Ie7GYo3_0),.clk(gclk));
	jdff dff_A_5v8gAEv80_0(.dout(G832),.din(w_dff_A_5v8gAEv80_0),.clk(gclk));
	jdff dff_A_ICQfSecU6_1(.dout(w_dff_A_HBq5g8BD2_0),.din(w_dff_A_ICQfSecU6_1),.clk(gclk));
	jdff dff_A_HBq5g8BD2_0(.dout(w_dff_A_UurNwGC50_0),.din(w_dff_A_HBq5g8BD2_0),.clk(gclk));
	jdff dff_A_UurNwGC50_0(.dout(w_dff_A_BMfZRL0S7_0),.din(w_dff_A_UurNwGC50_0),.clk(gclk));
	jdff dff_A_BMfZRL0S7_0(.dout(w_dff_A_zXAtMbVa4_0),.din(w_dff_A_BMfZRL0S7_0),.clk(gclk));
	jdff dff_A_zXAtMbVa4_0(.dout(w_dff_A_lNRIbo8S5_0),.din(w_dff_A_zXAtMbVa4_0),.clk(gclk));
	jdff dff_A_lNRIbo8S5_0(.dout(w_dff_A_mLd0LmI91_0),.din(w_dff_A_lNRIbo8S5_0),.clk(gclk));
	jdff dff_A_mLd0LmI91_0(.dout(w_dff_A_G7go82SA9_0),.din(w_dff_A_mLd0LmI91_0),.clk(gclk));
	jdff dff_A_G7go82SA9_0(.dout(w_dff_A_XMX7SZIL3_0),.din(w_dff_A_G7go82SA9_0),.clk(gclk));
	jdff dff_A_XMX7SZIL3_0(.dout(w_dff_A_bfLltZk06_0),.din(w_dff_A_XMX7SZIL3_0),.clk(gclk));
	jdff dff_A_bfLltZk06_0(.dout(w_dff_A_eWJlX53v9_0),.din(w_dff_A_bfLltZk06_0),.clk(gclk));
	jdff dff_A_eWJlX53v9_0(.dout(w_dff_A_VCaEGqlS3_0),.din(w_dff_A_eWJlX53v9_0),.clk(gclk));
	jdff dff_A_VCaEGqlS3_0(.dout(w_dff_A_R1gMeFM25_0),.din(w_dff_A_VCaEGqlS3_0),.clk(gclk));
	jdff dff_A_R1gMeFM25_0(.dout(w_dff_A_VpNYpXeO6_0),.din(w_dff_A_R1gMeFM25_0),.clk(gclk));
	jdff dff_A_VpNYpXeO6_0(.dout(G834),.din(w_dff_A_VpNYpXeO6_0),.clk(gclk));
	jdff dff_A_DX7YKSnO2_1(.dout(w_dff_A_V1ipFKI50_0),.din(w_dff_A_DX7YKSnO2_1),.clk(gclk));
	jdff dff_A_V1ipFKI50_0(.dout(w_dff_A_71wCERyd5_0),.din(w_dff_A_V1ipFKI50_0),.clk(gclk));
	jdff dff_A_71wCERyd5_0(.dout(w_dff_A_Qk0UTxZ88_0),.din(w_dff_A_71wCERyd5_0),.clk(gclk));
	jdff dff_A_Qk0UTxZ88_0(.dout(w_dff_A_bKMqDHhF2_0),.din(w_dff_A_Qk0UTxZ88_0),.clk(gclk));
	jdff dff_A_bKMqDHhF2_0(.dout(w_dff_A_9JDT9cUL6_0),.din(w_dff_A_bKMqDHhF2_0),.clk(gclk));
	jdff dff_A_9JDT9cUL6_0(.dout(w_dff_A_733b8GSb6_0),.din(w_dff_A_9JDT9cUL6_0),.clk(gclk));
	jdff dff_A_733b8GSb6_0(.dout(w_dff_A_5MfQFAFV6_0),.din(w_dff_A_733b8GSb6_0),.clk(gclk));
	jdff dff_A_5MfQFAFV6_0(.dout(w_dff_A_ZfBiNJ3K1_0),.din(w_dff_A_5MfQFAFV6_0),.clk(gclk));
	jdff dff_A_ZfBiNJ3K1_0(.dout(w_dff_A_ifCqtWTi1_0),.din(w_dff_A_ZfBiNJ3K1_0),.clk(gclk));
	jdff dff_A_ifCqtWTi1_0(.dout(w_dff_A_mpvxJe0J1_0),.din(w_dff_A_ifCqtWTi1_0),.clk(gclk));
	jdff dff_A_mpvxJe0J1_0(.dout(w_dff_A_T6zbLVaV4_0),.din(w_dff_A_mpvxJe0J1_0),.clk(gclk));
	jdff dff_A_T6zbLVaV4_0(.dout(w_dff_A_xH5JX65S8_0),.din(w_dff_A_T6zbLVaV4_0),.clk(gclk));
	jdff dff_A_xH5JX65S8_0(.dout(w_dff_A_XOZeyNdL8_0),.din(w_dff_A_xH5JX65S8_0),.clk(gclk));
	jdff dff_A_XOZeyNdL8_0(.dout(w_dff_A_h8iynxhB5_0),.din(w_dff_A_XOZeyNdL8_0),.clk(gclk));
	jdff dff_A_h8iynxhB5_0(.dout(w_dff_A_bVecHrRU9_0),.din(w_dff_A_h8iynxhB5_0),.clk(gclk));
	jdff dff_A_bVecHrRU9_0(.dout(G836),.din(w_dff_A_bVecHrRU9_0),.clk(gclk));
	jdff dff_A_YcIv6Ant5_2(.dout(w_dff_A_LvCLKEHe6_0),.din(w_dff_A_YcIv6Ant5_2),.clk(gclk));
	jdff dff_A_LvCLKEHe6_0(.dout(w_dff_A_p7Vu2e9s1_0),.din(w_dff_A_LvCLKEHe6_0),.clk(gclk));
	jdff dff_A_p7Vu2e9s1_0(.dout(w_dff_A_LCsMit8Q6_0),.din(w_dff_A_p7Vu2e9s1_0),.clk(gclk));
	jdff dff_A_LCsMit8Q6_0(.dout(w_dff_A_GjJmMtvB5_0),.din(w_dff_A_LCsMit8Q6_0),.clk(gclk));
	jdff dff_A_GjJmMtvB5_0(.dout(w_dff_A_1AE6zYd27_0),.din(w_dff_A_GjJmMtvB5_0),.clk(gclk));
	jdff dff_A_1AE6zYd27_0(.dout(w_dff_A_hvEwHQYS9_0),.din(w_dff_A_1AE6zYd27_0),.clk(gclk));
	jdff dff_A_hvEwHQYS9_0(.dout(w_dff_A_2uN7VHXT1_0),.din(w_dff_A_hvEwHQYS9_0),.clk(gclk));
	jdff dff_A_2uN7VHXT1_0(.dout(w_dff_A_gla9WPjz3_0),.din(w_dff_A_2uN7VHXT1_0),.clk(gclk));
	jdff dff_A_gla9WPjz3_0(.dout(w_dff_A_tfKgofmr3_0),.din(w_dff_A_gla9WPjz3_0),.clk(gclk));
	jdff dff_A_tfKgofmr3_0(.dout(w_dff_A_HdoQgVSL0_0),.din(w_dff_A_tfKgofmr3_0),.clk(gclk));
	jdff dff_A_HdoQgVSL0_0(.dout(w_dff_A_IckMEeNR6_0),.din(w_dff_A_HdoQgVSL0_0),.clk(gclk));
	jdff dff_A_IckMEeNR6_0(.dout(w_dff_A_YYKl1Pk89_0),.din(w_dff_A_IckMEeNR6_0),.clk(gclk));
	jdff dff_A_YYKl1Pk89_0(.dout(w_dff_A_8s3ojIhh0_0),.din(w_dff_A_YYKl1Pk89_0),.clk(gclk));
	jdff dff_A_8s3ojIhh0_0(.dout(G859),.din(w_dff_A_8s3ojIhh0_0),.clk(gclk));
	jdff dff_A_zejxgGKu4_1(.dout(w_dff_A_Swr7ePZR6_0),.din(w_dff_A_zejxgGKu4_1),.clk(gclk));
	jdff dff_A_Swr7ePZR6_0(.dout(w_dff_A_lxhTkNBZ7_0),.din(w_dff_A_Swr7ePZR6_0),.clk(gclk));
	jdff dff_A_lxhTkNBZ7_0(.dout(w_dff_A_7LmGl7iO2_0),.din(w_dff_A_lxhTkNBZ7_0),.clk(gclk));
	jdff dff_A_7LmGl7iO2_0(.dout(w_dff_A_3kEi4fWn7_0),.din(w_dff_A_7LmGl7iO2_0),.clk(gclk));
	jdff dff_A_3kEi4fWn7_0(.dout(w_dff_A_NqsgGsBB6_0),.din(w_dff_A_3kEi4fWn7_0),.clk(gclk));
	jdff dff_A_NqsgGsBB6_0(.dout(w_dff_A_vKsavxpf8_0),.din(w_dff_A_NqsgGsBB6_0),.clk(gclk));
	jdff dff_A_vKsavxpf8_0(.dout(w_dff_A_cC5lB1vs8_0),.din(w_dff_A_vKsavxpf8_0),.clk(gclk));
	jdff dff_A_cC5lB1vs8_0(.dout(w_dff_A_YZ7eOhAK6_0),.din(w_dff_A_cC5lB1vs8_0),.clk(gclk));
	jdff dff_A_YZ7eOhAK6_0(.dout(w_dff_A_CdxDHFtJ8_0),.din(w_dff_A_YZ7eOhAK6_0),.clk(gclk));
	jdff dff_A_CdxDHFtJ8_0(.dout(w_dff_A_pD1sp2v62_0),.din(w_dff_A_CdxDHFtJ8_0),.clk(gclk));
	jdff dff_A_pD1sp2v62_0(.dout(w_dff_A_T9d2ZPJ94_0),.din(w_dff_A_pD1sp2v62_0),.clk(gclk));
	jdff dff_A_T9d2ZPJ94_0(.dout(w_dff_A_ToOisfaa0_0),.din(w_dff_A_T9d2ZPJ94_0),.clk(gclk));
	jdff dff_A_ToOisfaa0_0(.dout(G871),.din(w_dff_A_ToOisfaa0_0),.clk(gclk));
	jdff dff_A_GJ5SWN8q8_1(.dout(w_dff_A_BAhmKwth2_0),.din(w_dff_A_GJ5SWN8q8_1),.clk(gclk));
	jdff dff_A_BAhmKwth2_0(.dout(w_dff_A_GiN9TrU71_0),.din(w_dff_A_BAhmKwth2_0),.clk(gclk));
	jdff dff_A_GiN9TrU71_0(.dout(w_dff_A_uzZ4rg3E6_0),.din(w_dff_A_GiN9TrU71_0),.clk(gclk));
	jdff dff_A_uzZ4rg3E6_0(.dout(w_dff_A_n2wEUx6e6_0),.din(w_dff_A_uzZ4rg3E6_0),.clk(gclk));
	jdff dff_A_n2wEUx6e6_0(.dout(w_dff_A_oikmc1Of0_0),.din(w_dff_A_n2wEUx6e6_0),.clk(gclk));
	jdff dff_A_oikmc1Of0_0(.dout(w_dff_A_LtPMtd7i4_0),.din(w_dff_A_oikmc1Of0_0),.clk(gclk));
	jdff dff_A_LtPMtd7i4_0(.dout(w_dff_A_ilgVdTpA3_0),.din(w_dff_A_LtPMtd7i4_0),.clk(gclk));
	jdff dff_A_ilgVdTpA3_0(.dout(w_dff_A_Q79gbO417_0),.din(w_dff_A_ilgVdTpA3_0),.clk(gclk));
	jdff dff_A_Q79gbO417_0(.dout(w_dff_A_tnGp9QKG4_0),.din(w_dff_A_Q79gbO417_0),.clk(gclk));
	jdff dff_A_tnGp9QKG4_0(.dout(w_dff_A_dCZ14Seu2_0),.din(w_dff_A_tnGp9QKG4_0),.clk(gclk));
	jdff dff_A_dCZ14Seu2_0(.dout(w_dff_A_tyhJ43JA8_0),.din(w_dff_A_dCZ14Seu2_0),.clk(gclk));
	jdff dff_A_tyhJ43JA8_0(.dout(w_dff_A_N9Y2z3J89_0),.din(w_dff_A_tyhJ43JA8_0),.clk(gclk));
	jdff dff_A_N9Y2z3J89_0(.dout(w_dff_A_Lm0zIVvd0_0),.din(w_dff_A_N9Y2z3J89_0),.clk(gclk));
	jdff dff_A_Lm0zIVvd0_0(.dout(w_dff_A_Tr4PIag82_0),.din(w_dff_A_Lm0zIVvd0_0),.clk(gclk));
	jdff dff_A_Tr4PIag82_0(.dout(G873),.din(w_dff_A_Tr4PIag82_0),.clk(gclk));
	jdff dff_A_Mw7p5bZZ9_1(.dout(w_dff_A_riPvdVm94_0),.din(w_dff_A_Mw7p5bZZ9_1),.clk(gclk));
	jdff dff_A_riPvdVm94_0(.dout(w_dff_A_96hsr8m75_0),.din(w_dff_A_riPvdVm94_0),.clk(gclk));
	jdff dff_A_96hsr8m75_0(.dout(w_dff_A_UDPQ0TMp0_0),.din(w_dff_A_96hsr8m75_0),.clk(gclk));
	jdff dff_A_UDPQ0TMp0_0(.dout(w_dff_A_NVelT6201_0),.din(w_dff_A_UDPQ0TMp0_0),.clk(gclk));
	jdff dff_A_NVelT6201_0(.dout(w_dff_A_zNyBUt6x9_0),.din(w_dff_A_NVelT6201_0),.clk(gclk));
	jdff dff_A_zNyBUt6x9_0(.dout(w_dff_A_QZloL7CX6_0),.din(w_dff_A_zNyBUt6x9_0),.clk(gclk));
	jdff dff_A_QZloL7CX6_0(.dout(w_dff_A_kIMkhQaN1_0),.din(w_dff_A_QZloL7CX6_0),.clk(gclk));
	jdff dff_A_kIMkhQaN1_0(.dout(w_dff_A_rOJqvXHS1_0),.din(w_dff_A_kIMkhQaN1_0),.clk(gclk));
	jdff dff_A_rOJqvXHS1_0(.dout(w_dff_A_Jx62Wi8y3_0),.din(w_dff_A_rOJqvXHS1_0),.clk(gclk));
	jdff dff_A_Jx62Wi8y3_0(.dout(w_dff_A_kyo4D9q72_0),.din(w_dff_A_Jx62Wi8y3_0),.clk(gclk));
	jdff dff_A_kyo4D9q72_0(.dout(w_dff_A_Xd1Dq2hO6_0),.din(w_dff_A_kyo4D9q72_0),.clk(gclk));
	jdff dff_A_Xd1Dq2hO6_0(.dout(w_dff_A_bU2asTuS1_0),.din(w_dff_A_Xd1Dq2hO6_0),.clk(gclk));
	jdff dff_A_bU2asTuS1_0(.dout(w_dff_A_EL2eZkGB1_0),.din(w_dff_A_bU2asTuS1_0),.clk(gclk));
	jdff dff_A_EL2eZkGB1_0(.dout(w_dff_A_0W3XIyY75_0),.din(w_dff_A_EL2eZkGB1_0),.clk(gclk));
	jdff dff_A_0W3XIyY75_0(.dout(w_dff_A_Cbga3JiT6_0),.din(w_dff_A_0W3XIyY75_0),.clk(gclk));
	jdff dff_A_Cbga3JiT6_0(.dout(G875),.din(w_dff_A_Cbga3JiT6_0),.clk(gclk));
	jdff dff_A_tYluNs5U4_1(.dout(w_dff_A_AkfcQQ514_0),.din(w_dff_A_tYluNs5U4_1),.clk(gclk));
	jdff dff_A_AkfcQQ514_0(.dout(w_dff_A_VOK4Vf6D5_0),.din(w_dff_A_AkfcQQ514_0),.clk(gclk));
	jdff dff_A_VOK4Vf6D5_0(.dout(w_dff_A_UfUGh8qC2_0),.din(w_dff_A_VOK4Vf6D5_0),.clk(gclk));
	jdff dff_A_UfUGh8qC2_0(.dout(w_dff_A_lfufGkjl8_0),.din(w_dff_A_UfUGh8qC2_0),.clk(gclk));
	jdff dff_A_lfufGkjl8_0(.dout(w_dff_A_k1MVLzG81_0),.din(w_dff_A_lfufGkjl8_0),.clk(gclk));
	jdff dff_A_k1MVLzG81_0(.dout(w_dff_A_ZDMPVXmH9_0),.din(w_dff_A_k1MVLzG81_0),.clk(gclk));
	jdff dff_A_ZDMPVXmH9_0(.dout(w_dff_A_Z18riH2b9_0),.din(w_dff_A_ZDMPVXmH9_0),.clk(gclk));
	jdff dff_A_Z18riH2b9_0(.dout(w_dff_A_bxd1OX6V3_0),.din(w_dff_A_Z18riH2b9_0),.clk(gclk));
	jdff dff_A_bxd1OX6V3_0(.dout(w_dff_A_A7s0WCXi5_0),.din(w_dff_A_bxd1OX6V3_0),.clk(gclk));
	jdff dff_A_A7s0WCXi5_0(.dout(w_dff_A_1hb5tI9c0_0),.din(w_dff_A_A7s0WCXi5_0),.clk(gclk));
	jdff dff_A_1hb5tI9c0_0(.dout(w_dff_A_WruQ7unO2_0),.din(w_dff_A_1hb5tI9c0_0),.clk(gclk));
	jdff dff_A_WruQ7unO2_0(.dout(w_dff_A_AG1Yefvt4_0),.din(w_dff_A_WruQ7unO2_0),.clk(gclk));
	jdff dff_A_AG1Yefvt4_0(.dout(w_dff_A_Js2Iwlbi9_0),.din(w_dff_A_AG1Yefvt4_0),.clk(gclk));
	jdff dff_A_Js2Iwlbi9_0(.dout(w_dff_A_SDeLTR803_0),.din(w_dff_A_Js2Iwlbi9_0),.clk(gclk));
	jdff dff_A_SDeLTR803_0(.dout(w_dff_A_lxbpSUFO1_0),.din(w_dff_A_SDeLTR803_0),.clk(gclk));
	jdff dff_A_lxbpSUFO1_0(.dout(w_dff_A_VZhTkJ8A9_0),.din(w_dff_A_lxbpSUFO1_0),.clk(gclk));
	jdff dff_A_VZhTkJ8A9_0(.dout(G877),.din(w_dff_A_VZhTkJ8A9_0),.clk(gclk));
	jdff dff_A_VCOqhx971_1(.dout(w_dff_A_DSsVtlGx1_0),.din(w_dff_A_VCOqhx971_1),.clk(gclk));
	jdff dff_A_DSsVtlGx1_0(.dout(w_dff_A_bvgUWODH4_0),.din(w_dff_A_DSsVtlGx1_0),.clk(gclk));
	jdff dff_A_bvgUWODH4_0(.dout(w_dff_A_wx7f1ws41_0),.din(w_dff_A_bvgUWODH4_0),.clk(gclk));
	jdff dff_A_wx7f1ws41_0(.dout(w_dff_A_lll9M0gF2_0),.din(w_dff_A_wx7f1ws41_0),.clk(gclk));
	jdff dff_A_lll9M0gF2_0(.dout(w_dff_A_VDnvuVfq4_0),.din(w_dff_A_lll9M0gF2_0),.clk(gclk));
	jdff dff_A_VDnvuVfq4_0(.dout(w_dff_A_B7n5shkg1_0),.din(w_dff_A_VDnvuVfq4_0),.clk(gclk));
	jdff dff_A_B7n5shkg1_0(.dout(w_dff_A_rIVw8x059_0),.din(w_dff_A_B7n5shkg1_0),.clk(gclk));
	jdff dff_A_rIVw8x059_0(.dout(w_dff_A_kc5eWfPe8_0),.din(w_dff_A_rIVw8x059_0),.clk(gclk));
	jdff dff_A_kc5eWfPe8_0(.dout(w_dff_A_GruaQll22_0),.din(w_dff_A_kc5eWfPe8_0),.clk(gclk));
	jdff dff_A_GruaQll22_0(.dout(w_dff_A_GomFKmbj6_0),.din(w_dff_A_GruaQll22_0),.clk(gclk));
	jdff dff_A_GomFKmbj6_0(.dout(w_dff_A_nIofH8gm5_0),.din(w_dff_A_GomFKmbj6_0),.clk(gclk));
	jdff dff_A_nIofH8gm5_0(.dout(w_dff_A_Qkga69BT1_0),.din(w_dff_A_nIofH8gm5_0),.clk(gclk));
	jdff dff_A_Qkga69BT1_0(.dout(w_dff_A_Zs6yYYrq1_0),.din(w_dff_A_Qkga69BT1_0),.clk(gclk));
	jdff dff_A_Zs6yYYrq1_0(.dout(w_dff_A_6mdw8nKD8_0),.din(w_dff_A_Zs6yYYrq1_0),.clk(gclk));
	jdff dff_A_6mdw8nKD8_0(.dout(w_dff_A_zjPEDVJY6_0),.din(w_dff_A_6mdw8nKD8_0),.clk(gclk));
	jdff dff_A_zjPEDVJY6_0(.dout(w_dff_A_gisvbRPS4_0),.din(w_dff_A_zjPEDVJY6_0),.clk(gclk));
	jdff dff_A_gisvbRPS4_0(.dout(w_dff_A_wMQj2HOW1_0),.din(w_dff_A_gisvbRPS4_0),.clk(gclk));
	jdff dff_A_wMQj2HOW1_0(.dout(w_dff_A_ZeDwIcdB4_0),.din(w_dff_A_wMQj2HOW1_0),.clk(gclk));
	jdff dff_A_ZeDwIcdB4_0(.dout(w_dff_A_w5QIYCX30_0),.din(w_dff_A_ZeDwIcdB4_0),.clk(gclk));
	jdff dff_A_w5QIYCX30_0(.dout(G998),.din(w_dff_A_w5QIYCX30_0),.clk(gclk));
	jdff dff_A_LwGy0wKt8_1(.dout(w_dff_A_UMWbK1I59_0),.din(w_dff_A_LwGy0wKt8_1),.clk(gclk));
	jdff dff_A_UMWbK1I59_0(.dout(w_dff_A_wOpQxbba9_0),.din(w_dff_A_UMWbK1I59_0),.clk(gclk));
	jdff dff_A_wOpQxbba9_0(.dout(w_dff_A_H628PjGa7_0),.din(w_dff_A_wOpQxbba9_0),.clk(gclk));
	jdff dff_A_H628PjGa7_0(.dout(w_dff_A_5dcQwNL23_0),.din(w_dff_A_H628PjGa7_0),.clk(gclk));
	jdff dff_A_5dcQwNL23_0(.dout(w_dff_A_RI9xOgm12_0),.din(w_dff_A_5dcQwNL23_0),.clk(gclk));
	jdff dff_A_RI9xOgm12_0(.dout(w_dff_A_6mZPKRnS4_0),.din(w_dff_A_RI9xOgm12_0),.clk(gclk));
	jdff dff_A_6mZPKRnS4_0(.dout(w_dff_A_byCsdSYY1_0),.din(w_dff_A_6mZPKRnS4_0),.clk(gclk));
	jdff dff_A_byCsdSYY1_0(.dout(w_dff_A_RE8xx5Y86_0),.din(w_dff_A_byCsdSYY1_0),.clk(gclk));
	jdff dff_A_RE8xx5Y86_0(.dout(w_dff_A_Gz7OPc0w6_0),.din(w_dff_A_RE8xx5Y86_0),.clk(gclk));
	jdff dff_A_Gz7OPc0w6_0(.dout(w_dff_A_Ey6ZTc9l3_0),.din(w_dff_A_Gz7OPc0w6_0),.clk(gclk));
	jdff dff_A_Ey6ZTc9l3_0(.dout(w_dff_A_5pYGop5e6_0),.din(w_dff_A_Ey6ZTc9l3_0),.clk(gclk));
	jdff dff_A_5pYGop5e6_0(.dout(w_dff_A_USPkTnw22_0),.din(w_dff_A_5pYGop5e6_0),.clk(gclk));
	jdff dff_A_USPkTnw22_0(.dout(w_dff_A_8hLPYmK71_0),.din(w_dff_A_USPkTnw22_0),.clk(gclk));
	jdff dff_A_8hLPYmK71_0(.dout(w_dff_A_qNgihvDH8_0),.din(w_dff_A_8hLPYmK71_0),.clk(gclk));
	jdff dff_A_qNgihvDH8_0(.dout(w_dff_A_Xjdwz6K91_0),.din(w_dff_A_qNgihvDH8_0),.clk(gclk));
	jdff dff_A_Xjdwz6K91_0(.dout(w_dff_A_3OgcdmYG1_0),.din(w_dff_A_Xjdwz6K91_0),.clk(gclk));
	jdff dff_A_3OgcdmYG1_0(.dout(w_dff_A_PYPhHZgk5_0),.din(w_dff_A_3OgcdmYG1_0),.clk(gclk));
	jdff dff_A_PYPhHZgk5_0(.dout(w_dff_A_42ToleIv4_0),.din(w_dff_A_PYPhHZgk5_0),.clk(gclk));
	jdff dff_A_42ToleIv4_0(.dout(G1000),.din(w_dff_A_42ToleIv4_0),.clk(gclk));
	jdff dff_A_FSDJereM4_2(.dout(w_dff_A_HHiqvebf1_0),.din(w_dff_A_FSDJereM4_2),.clk(gclk));
	jdff dff_A_HHiqvebf1_0(.dout(w_dff_A_dJUBUOwU3_0),.din(w_dff_A_HHiqvebf1_0),.clk(gclk));
	jdff dff_A_dJUBUOwU3_0(.dout(w_dff_A_lub9GHR85_0),.din(w_dff_A_dJUBUOwU3_0),.clk(gclk));
	jdff dff_A_lub9GHR85_0(.dout(w_dff_A_JOpDG86Z1_0),.din(w_dff_A_lub9GHR85_0),.clk(gclk));
	jdff dff_A_JOpDG86Z1_0(.dout(w_dff_A_dLcHtqtE8_0),.din(w_dff_A_JOpDG86Z1_0),.clk(gclk));
	jdff dff_A_dLcHtqtE8_0(.dout(w_dff_A_R51BVZxY1_0),.din(w_dff_A_dLcHtqtE8_0),.clk(gclk));
	jdff dff_A_R51BVZxY1_0(.dout(w_dff_A_WF5LyqbK8_0),.din(w_dff_A_R51BVZxY1_0),.clk(gclk));
	jdff dff_A_WF5LyqbK8_0(.dout(G575),.din(w_dff_A_WF5LyqbK8_0),.clk(gclk));
	jdff dff_A_5ltDjXuT8_2(.dout(w_dff_A_9elRzTD92_0),.din(w_dff_A_5ltDjXuT8_2),.clk(gclk));
	jdff dff_A_9elRzTD92_0(.dout(w_dff_A_13r5drHY0_0),.din(w_dff_A_9elRzTD92_0),.clk(gclk));
	jdff dff_A_13r5drHY0_0(.dout(w_dff_A_tKUZ6f0L6_0),.din(w_dff_A_13r5drHY0_0),.clk(gclk));
	jdff dff_A_tKUZ6f0L6_0(.dout(w_dff_A_ShtN6qJE5_0),.din(w_dff_A_tKUZ6f0L6_0),.clk(gclk));
	jdff dff_A_ShtN6qJE5_0(.dout(w_dff_A_u0euAwMQ6_0),.din(w_dff_A_ShtN6qJE5_0),.clk(gclk));
	jdff dff_A_u0euAwMQ6_0(.dout(w_dff_A_nB7mZ6QU1_0),.din(w_dff_A_u0euAwMQ6_0),.clk(gclk));
	jdff dff_A_nB7mZ6QU1_0(.dout(G585),.din(w_dff_A_nB7mZ6QU1_0),.clk(gclk));
	jdff dff_A_09IHvNaL4_2(.dout(w_dff_A_0z5KShPv8_0),.din(w_dff_A_09IHvNaL4_2),.clk(gclk));
	jdff dff_A_0z5KShPv8_0(.dout(w_dff_A_wdlBjPRD8_0),.din(w_dff_A_0z5KShPv8_0),.clk(gclk));
	jdff dff_A_wdlBjPRD8_0(.dout(w_dff_A_avpExcFZ4_0),.din(w_dff_A_wdlBjPRD8_0),.clk(gclk));
	jdff dff_A_avpExcFZ4_0(.dout(w_dff_A_ZRN1OL2a7_0),.din(w_dff_A_avpExcFZ4_0),.clk(gclk));
	jdff dff_A_ZRN1OL2a7_0(.dout(w_dff_A_jzCJoAw88_0),.din(w_dff_A_ZRN1OL2a7_0),.clk(gclk));
	jdff dff_A_jzCJoAw88_0(.dout(w_dff_A_9kWVhh6m3_0),.din(w_dff_A_jzCJoAw88_0),.clk(gclk));
	jdff dff_A_9kWVhh6m3_0(.dout(w_dff_A_rfuAabCB2_0),.din(w_dff_A_9kWVhh6m3_0),.clk(gclk));
	jdff dff_A_rfuAabCB2_0(.dout(w_dff_A_iPLSuyM16_0),.din(w_dff_A_rfuAabCB2_0),.clk(gclk));
	jdff dff_A_iPLSuyM16_0(.dout(w_dff_A_I5lE0ZMI8_0),.din(w_dff_A_iPLSuyM16_0),.clk(gclk));
	jdff dff_A_I5lE0ZMI8_0(.dout(w_dff_A_jId4hxGS5_0),.din(w_dff_A_I5lE0ZMI8_0),.clk(gclk));
	jdff dff_A_jId4hxGS5_0(.dout(w_dff_A_GD0IxNRl0_0),.din(w_dff_A_jId4hxGS5_0),.clk(gclk));
	jdff dff_A_GD0IxNRl0_0(.dout(G661),.din(w_dff_A_GD0IxNRl0_0),.clk(gclk));
	jdff dff_A_SWMAgAUJ9_2(.dout(w_dff_A_X8hPznN83_0),.din(w_dff_A_SWMAgAUJ9_2),.clk(gclk));
	jdff dff_A_X8hPznN83_0(.dout(w_dff_A_t7Y1YB2L2_0),.din(w_dff_A_X8hPznN83_0),.clk(gclk));
	jdff dff_A_t7Y1YB2L2_0(.dout(w_dff_A_gRc20hDv8_0),.din(w_dff_A_t7Y1YB2L2_0),.clk(gclk));
	jdff dff_A_gRc20hDv8_0(.dout(w_dff_A_ZqvBhCuH3_0),.din(w_dff_A_gRc20hDv8_0),.clk(gclk));
	jdff dff_A_ZqvBhCuH3_0(.dout(w_dff_A_jjchhgrc3_0),.din(w_dff_A_ZqvBhCuH3_0),.clk(gclk));
	jdff dff_A_jjchhgrc3_0(.dout(w_dff_A_2Df1oeOe4_0),.din(w_dff_A_jjchhgrc3_0),.clk(gclk));
	jdff dff_A_2Df1oeOe4_0(.dout(w_dff_A_0X8yqpJ23_0),.din(w_dff_A_2Df1oeOe4_0),.clk(gclk));
	jdff dff_A_0X8yqpJ23_0(.dout(w_dff_A_JglzB5JZ1_0),.din(w_dff_A_0X8yqpJ23_0),.clk(gclk));
	jdff dff_A_JglzB5JZ1_0(.dout(w_dff_A_vtKLSkfV0_0),.din(w_dff_A_JglzB5JZ1_0),.clk(gclk));
	jdff dff_A_vtKLSkfV0_0(.dout(w_dff_A_iAdslHC67_0),.din(w_dff_A_vtKLSkfV0_0),.clk(gclk));
	jdff dff_A_iAdslHC67_0(.dout(w_dff_A_Vs5YWyeM5_0),.din(w_dff_A_iAdslHC67_0),.clk(gclk));
	jdff dff_A_Vs5YWyeM5_0(.dout(G693),.din(w_dff_A_Vs5YWyeM5_0),.clk(gclk));
	jdff dff_A_Z13qQidg2_2(.dout(w_dff_A_iaw37lKi0_0),.din(w_dff_A_Z13qQidg2_2),.clk(gclk));
	jdff dff_A_iaw37lKi0_0(.dout(w_dff_A_PJIlZVhL5_0),.din(w_dff_A_iaw37lKi0_0),.clk(gclk));
	jdff dff_A_PJIlZVhL5_0(.dout(w_dff_A_nPVp7hgW5_0),.din(w_dff_A_PJIlZVhL5_0),.clk(gclk));
	jdff dff_A_nPVp7hgW5_0(.dout(w_dff_A_Msx2FQCk2_0),.din(w_dff_A_nPVp7hgW5_0),.clk(gclk));
	jdff dff_A_Msx2FQCk2_0(.dout(w_dff_A_OnEzG93A8_0),.din(w_dff_A_Msx2FQCk2_0),.clk(gclk));
	jdff dff_A_OnEzG93A8_0(.dout(w_dff_A_686Kjme78_0),.din(w_dff_A_OnEzG93A8_0),.clk(gclk));
	jdff dff_A_686Kjme78_0(.dout(w_dff_A_zC53FGcG8_0),.din(w_dff_A_686Kjme78_0),.clk(gclk));
	jdff dff_A_zC53FGcG8_0(.dout(G747),.din(w_dff_A_zC53FGcG8_0),.clk(gclk));
	jdff dff_A_NZTKntos3_2(.dout(w_dff_A_E6caPdRQ5_0),.din(w_dff_A_NZTKntos3_2),.clk(gclk));
	jdff dff_A_E6caPdRQ5_0(.dout(w_dff_A_UFV7DIaL8_0),.din(w_dff_A_E6caPdRQ5_0),.clk(gclk));
	jdff dff_A_UFV7DIaL8_0(.dout(w_dff_A_1TEYMkQF2_0),.din(w_dff_A_UFV7DIaL8_0),.clk(gclk));
	jdff dff_A_1TEYMkQF2_0(.dout(w_dff_A_jshwYzZa9_0),.din(w_dff_A_1TEYMkQF2_0),.clk(gclk));
	jdff dff_A_jshwYzZa9_0(.dout(w_dff_A_h08DBtkS3_0),.din(w_dff_A_jshwYzZa9_0),.clk(gclk));
	jdff dff_A_h08DBtkS3_0(.dout(w_dff_A_HJmdpaXa5_0),.din(w_dff_A_h08DBtkS3_0),.clk(gclk));
	jdff dff_A_HJmdpaXa5_0(.dout(w_dff_A_aZfPtXqN0_0),.din(w_dff_A_HJmdpaXa5_0),.clk(gclk));
	jdff dff_A_aZfPtXqN0_0(.dout(w_dff_A_daZ8IuUb1_0),.din(w_dff_A_aZfPtXqN0_0),.clk(gclk));
	jdff dff_A_daZ8IuUb1_0(.dout(G752),.din(w_dff_A_daZ8IuUb1_0),.clk(gclk));
	jdff dff_A_qtJUbwCW9_2(.dout(w_dff_A_OQdHWbEG0_0),.din(w_dff_A_qtJUbwCW9_2),.clk(gclk));
	jdff dff_A_OQdHWbEG0_0(.dout(w_dff_A_ld4v8GRD8_0),.din(w_dff_A_OQdHWbEG0_0),.clk(gclk));
	jdff dff_A_ld4v8GRD8_0(.dout(w_dff_A_BvsGC0n13_0),.din(w_dff_A_ld4v8GRD8_0),.clk(gclk));
	jdff dff_A_BvsGC0n13_0(.dout(w_dff_A_v46Juft24_0),.din(w_dff_A_BvsGC0n13_0),.clk(gclk));
	jdff dff_A_v46Juft24_0(.dout(w_dff_A_jv2rH8Mi2_0),.din(w_dff_A_v46Juft24_0),.clk(gclk));
	jdff dff_A_jv2rH8Mi2_0(.dout(w_dff_A_ZEUcR0DH0_0),.din(w_dff_A_jv2rH8Mi2_0),.clk(gclk));
	jdff dff_A_ZEUcR0DH0_0(.dout(w_dff_A_vksXmgQj2_0),.din(w_dff_A_ZEUcR0DH0_0),.clk(gclk));
	jdff dff_A_vksXmgQj2_0(.dout(w_dff_A_XeOilhG90_0),.din(w_dff_A_vksXmgQj2_0),.clk(gclk));
	jdff dff_A_XeOilhG90_0(.dout(w_dff_A_gjWOBSJW8_0),.din(w_dff_A_XeOilhG90_0),.clk(gclk));
	jdff dff_A_gjWOBSJW8_0(.dout(w_dff_A_8sHvb8cP2_0),.din(w_dff_A_gjWOBSJW8_0),.clk(gclk));
	jdff dff_A_8sHvb8cP2_0(.dout(G757),.din(w_dff_A_8sHvb8cP2_0),.clk(gclk));
	jdff dff_A_0IUNpq9e5_2(.dout(w_dff_A_qjBO1FYl0_0),.din(w_dff_A_0IUNpq9e5_2),.clk(gclk));
	jdff dff_A_qjBO1FYl0_0(.dout(w_dff_A_lyixb6jW9_0),.din(w_dff_A_qjBO1FYl0_0),.clk(gclk));
	jdff dff_A_lyixb6jW9_0(.dout(w_dff_A_BEnYyW0t0_0),.din(w_dff_A_lyixb6jW9_0),.clk(gclk));
	jdff dff_A_BEnYyW0t0_0(.dout(w_dff_A_MV8PkqOu3_0),.din(w_dff_A_BEnYyW0t0_0),.clk(gclk));
	jdff dff_A_MV8PkqOu3_0(.dout(w_dff_A_ALKN8NLc6_0),.din(w_dff_A_MV8PkqOu3_0),.clk(gclk));
	jdff dff_A_ALKN8NLc6_0(.dout(w_dff_A_J35WFDl26_0),.din(w_dff_A_ALKN8NLc6_0),.clk(gclk));
	jdff dff_A_J35WFDl26_0(.dout(w_dff_A_9Y82Ca4a4_0),.din(w_dff_A_J35WFDl26_0),.clk(gclk));
	jdff dff_A_9Y82Ca4a4_0(.dout(w_dff_A_pfcEfYFX1_0),.din(w_dff_A_9Y82Ca4a4_0),.clk(gclk));
	jdff dff_A_pfcEfYFX1_0(.dout(w_dff_A_hxEKEWhE7_0),.din(w_dff_A_pfcEfYFX1_0),.clk(gclk));
	jdff dff_A_hxEKEWhE7_0(.dout(G762),.din(w_dff_A_hxEKEWhE7_0),.clk(gclk));
	jdff dff_A_7okTC8Yv1_2(.dout(w_dff_A_UdOHfssJ2_0),.din(w_dff_A_7okTC8Yv1_2),.clk(gclk));
	jdff dff_A_UdOHfssJ2_0(.dout(w_dff_A_wUyKTX7H2_0),.din(w_dff_A_UdOHfssJ2_0),.clk(gclk));
	jdff dff_A_wUyKTX7H2_0(.dout(w_dff_A_136G7pCc2_0),.din(w_dff_A_wUyKTX7H2_0),.clk(gclk));
	jdff dff_A_136G7pCc2_0(.dout(w_dff_A_6xN0F4Ky9_0),.din(w_dff_A_136G7pCc2_0),.clk(gclk));
	jdff dff_A_6xN0F4Ky9_0(.dout(w_dff_A_El1yBSPs2_0),.din(w_dff_A_6xN0F4Ky9_0),.clk(gclk));
	jdff dff_A_El1yBSPs2_0(.dout(w_dff_A_jc0Nd6Ch7_0),.din(w_dff_A_El1yBSPs2_0),.clk(gclk));
	jdff dff_A_jc0Nd6Ch7_0(.dout(w_dff_A_N7VnJMEt4_0),.din(w_dff_A_jc0Nd6Ch7_0),.clk(gclk));
	jdff dff_A_N7VnJMEt4_0(.dout(G787),.din(w_dff_A_N7VnJMEt4_0),.clk(gclk));
	jdff dff_A_la5HpM0d0_2(.dout(w_dff_A_uhU1qVvX1_0),.din(w_dff_A_la5HpM0d0_2),.clk(gclk));
	jdff dff_A_uhU1qVvX1_0(.dout(w_dff_A_ld8Okegi0_0),.din(w_dff_A_uhU1qVvX1_0),.clk(gclk));
	jdff dff_A_ld8Okegi0_0(.dout(w_dff_A_rwPsz4Vu7_0),.din(w_dff_A_ld8Okegi0_0),.clk(gclk));
	jdff dff_A_rwPsz4Vu7_0(.dout(w_dff_A_MvUyKAxC6_0),.din(w_dff_A_rwPsz4Vu7_0),.clk(gclk));
	jdff dff_A_MvUyKAxC6_0(.dout(w_dff_A_b47ixkoL5_0),.din(w_dff_A_MvUyKAxC6_0),.clk(gclk));
	jdff dff_A_b47ixkoL5_0(.dout(w_dff_A_x6MDbt6g2_0),.din(w_dff_A_b47ixkoL5_0),.clk(gclk));
	jdff dff_A_x6MDbt6g2_0(.dout(w_dff_A_d4v70wGJ5_0),.din(w_dff_A_x6MDbt6g2_0),.clk(gclk));
	jdff dff_A_d4v70wGJ5_0(.dout(w_dff_A_TZiQctQs4_0),.din(w_dff_A_d4v70wGJ5_0),.clk(gclk));
	jdff dff_A_TZiQctQs4_0(.dout(G792),.din(w_dff_A_TZiQctQs4_0),.clk(gclk));
	jdff dff_A_K4sCI48D9_2(.dout(w_dff_A_uK49aPco9_0),.din(w_dff_A_K4sCI48D9_2),.clk(gclk));
	jdff dff_A_uK49aPco9_0(.dout(w_dff_A_bPgwSsLQ7_0),.din(w_dff_A_uK49aPco9_0),.clk(gclk));
	jdff dff_A_bPgwSsLQ7_0(.dout(w_dff_A_4DRn44Wr6_0),.din(w_dff_A_bPgwSsLQ7_0),.clk(gclk));
	jdff dff_A_4DRn44Wr6_0(.dout(w_dff_A_zp1xJMM23_0),.din(w_dff_A_4DRn44Wr6_0),.clk(gclk));
	jdff dff_A_zp1xJMM23_0(.dout(w_dff_A_1MHXBTZU7_0),.din(w_dff_A_zp1xJMM23_0),.clk(gclk));
	jdff dff_A_1MHXBTZU7_0(.dout(w_dff_A_xTISa4Gm6_0),.din(w_dff_A_1MHXBTZU7_0),.clk(gclk));
	jdff dff_A_xTISa4Gm6_0(.dout(w_dff_A_pEwuXo406_0),.din(w_dff_A_xTISa4Gm6_0),.clk(gclk));
	jdff dff_A_pEwuXo406_0(.dout(w_dff_A_rrLmQzxn5_0),.din(w_dff_A_pEwuXo406_0),.clk(gclk));
	jdff dff_A_rrLmQzxn5_0(.dout(w_dff_A_Lf5p5ICS0_0),.din(w_dff_A_rrLmQzxn5_0),.clk(gclk));
	jdff dff_A_Lf5p5ICS0_0(.dout(w_dff_A_mzwdSda61_0),.din(w_dff_A_Lf5p5ICS0_0),.clk(gclk));
	jdff dff_A_mzwdSda61_0(.dout(G797),.din(w_dff_A_mzwdSda61_0),.clk(gclk));
	jdff dff_A_aqlIY8yf5_2(.dout(w_dff_A_DFSNL7144_0),.din(w_dff_A_aqlIY8yf5_2),.clk(gclk));
	jdff dff_A_DFSNL7144_0(.dout(w_dff_A_rmPsxOxx1_0),.din(w_dff_A_DFSNL7144_0),.clk(gclk));
	jdff dff_A_rmPsxOxx1_0(.dout(w_dff_A_amVKJrEN7_0),.din(w_dff_A_rmPsxOxx1_0),.clk(gclk));
	jdff dff_A_amVKJrEN7_0(.dout(w_dff_A_oxQn4gGd5_0),.din(w_dff_A_amVKJrEN7_0),.clk(gclk));
	jdff dff_A_oxQn4gGd5_0(.dout(w_dff_A_7eb8C3BA7_0),.din(w_dff_A_oxQn4gGd5_0),.clk(gclk));
	jdff dff_A_7eb8C3BA7_0(.dout(w_dff_A_t4oGr6SV6_0),.din(w_dff_A_7eb8C3BA7_0),.clk(gclk));
	jdff dff_A_t4oGr6SV6_0(.dout(w_dff_A_xRwmHPoW1_0),.din(w_dff_A_t4oGr6SV6_0),.clk(gclk));
	jdff dff_A_xRwmHPoW1_0(.dout(w_dff_A_bNr40E0a0_0),.din(w_dff_A_xRwmHPoW1_0),.clk(gclk));
	jdff dff_A_bNr40E0a0_0(.dout(w_dff_A_ZOWXptlU5_0),.din(w_dff_A_bNr40E0a0_0),.clk(gclk));
	jdff dff_A_ZOWXptlU5_0(.dout(G802),.din(w_dff_A_ZOWXptlU5_0),.clk(gclk));
	jdff dff_A_eXtTYCE04_2(.dout(w_dff_A_vLQhPHQD5_0),.din(w_dff_A_eXtTYCE04_2),.clk(gclk));
	jdff dff_A_vLQhPHQD5_0(.dout(w_dff_A_MscugdSa8_0),.din(w_dff_A_vLQhPHQD5_0),.clk(gclk));
	jdff dff_A_MscugdSa8_0(.dout(w_dff_A_NLAFOEsr3_0),.din(w_dff_A_MscugdSa8_0),.clk(gclk));
	jdff dff_A_NLAFOEsr3_0(.dout(w_dff_A_84gJBveH0_0),.din(w_dff_A_NLAFOEsr3_0),.clk(gclk));
	jdff dff_A_84gJBveH0_0(.dout(w_dff_A_loWyxih61_0),.din(w_dff_A_84gJBveH0_0),.clk(gclk));
	jdff dff_A_loWyxih61_0(.dout(w_dff_A_DPlg8d4j7_0),.din(w_dff_A_loWyxih61_0),.clk(gclk));
	jdff dff_A_DPlg8d4j7_0(.dout(G642),.din(w_dff_A_DPlg8d4j7_0),.clk(gclk));
	jdff dff_A_vEcDfA282_2(.dout(w_dff_A_hjGNh0Ov3_0),.din(w_dff_A_vEcDfA282_2),.clk(gclk));
	jdff dff_A_hjGNh0Ov3_0(.dout(w_dff_A_yICnxMbu7_0),.din(w_dff_A_hjGNh0Ov3_0),.clk(gclk));
	jdff dff_A_yICnxMbu7_0(.dout(w_dff_A_J4t0CWys9_0),.din(w_dff_A_yICnxMbu7_0),.clk(gclk));
	jdff dff_A_J4t0CWys9_0(.dout(w_dff_A_85X6aOHD4_0),.din(w_dff_A_J4t0CWys9_0),.clk(gclk));
	jdff dff_A_85X6aOHD4_0(.dout(w_dff_A_q0fHmOFP9_0),.din(w_dff_A_85X6aOHD4_0),.clk(gclk));
	jdff dff_A_q0fHmOFP9_0(.dout(w_dff_A_hh8VPUhr5_0),.din(w_dff_A_q0fHmOFP9_0),.clk(gclk));
	jdff dff_A_hh8VPUhr5_0(.dout(w_dff_A_zd9X5JB64_0),.din(w_dff_A_hh8VPUhr5_0),.clk(gclk));
	jdff dff_A_zd9X5JB64_0(.dout(w_dff_A_82lGhO7J4_0),.din(w_dff_A_zd9X5JB64_0),.clk(gclk));
	jdff dff_A_82lGhO7J4_0(.dout(w_dff_A_DN1txea69_0),.din(w_dff_A_82lGhO7J4_0),.clk(gclk));
	jdff dff_A_DN1txea69_0(.dout(G664),.din(w_dff_A_DN1txea69_0),.clk(gclk));
	jdff dff_A_b47UtnYZ5_2(.dout(w_dff_A_RNg2sWhJ3_0),.din(w_dff_A_b47UtnYZ5_2),.clk(gclk));
	jdff dff_A_RNg2sWhJ3_0(.dout(w_dff_A_bTnVNkDb6_0),.din(w_dff_A_RNg2sWhJ3_0),.clk(gclk));
	jdff dff_A_bTnVNkDb6_0(.dout(w_dff_A_PRX7tc082_0),.din(w_dff_A_bTnVNkDb6_0),.clk(gclk));
	jdff dff_A_PRX7tc082_0(.dout(w_dff_A_L689P2z35_0),.din(w_dff_A_PRX7tc082_0),.clk(gclk));
	jdff dff_A_L689P2z35_0(.dout(w_dff_A_6LTlPDZi0_0),.din(w_dff_A_L689P2z35_0),.clk(gclk));
	jdff dff_A_6LTlPDZi0_0(.dout(w_dff_A_xBqalnDu3_0),.din(w_dff_A_6LTlPDZi0_0),.clk(gclk));
	jdff dff_A_xBqalnDu3_0(.dout(w_dff_A_Jtl3DNmx6_0),.din(w_dff_A_xBqalnDu3_0),.clk(gclk));
	jdff dff_A_Jtl3DNmx6_0(.dout(w_dff_A_W5aAhiir0_0),.din(w_dff_A_Jtl3DNmx6_0),.clk(gclk));
	jdff dff_A_W5aAhiir0_0(.dout(w_dff_A_XwjwO0SP4_0),.din(w_dff_A_W5aAhiir0_0),.clk(gclk));
	jdff dff_A_XwjwO0SP4_0(.dout(G667),.din(w_dff_A_XwjwO0SP4_0),.clk(gclk));
	jdff dff_A_TjGCcada8_2(.dout(w_dff_A_lNidFfVa1_0),.din(w_dff_A_TjGCcada8_2),.clk(gclk));
	jdff dff_A_lNidFfVa1_0(.dout(w_dff_A_HnHEaCUI1_0),.din(w_dff_A_lNidFfVa1_0),.clk(gclk));
	jdff dff_A_HnHEaCUI1_0(.dout(w_dff_A_XwUVbQzP7_0),.din(w_dff_A_HnHEaCUI1_0),.clk(gclk));
	jdff dff_A_XwUVbQzP7_0(.dout(w_dff_A_CnVd3AWM2_0),.din(w_dff_A_XwUVbQzP7_0),.clk(gclk));
	jdff dff_A_CnVd3AWM2_0(.dout(w_dff_A_3sCpdZ7t4_0),.din(w_dff_A_CnVd3AWM2_0),.clk(gclk));
	jdff dff_A_3sCpdZ7t4_0(.dout(w_dff_A_EwaKgt3w8_0),.din(w_dff_A_3sCpdZ7t4_0),.clk(gclk));
	jdff dff_A_EwaKgt3w8_0(.dout(w_dff_A_4JjTPkhD2_0),.din(w_dff_A_EwaKgt3w8_0),.clk(gclk));
	jdff dff_A_4JjTPkhD2_0(.dout(w_dff_A_r0clN1f40_0),.din(w_dff_A_4JjTPkhD2_0),.clk(gclk));
	jdff dff_A_r0clN1f40_0(.dout(G670),.din(w_dff_A_r0clN1f40_0),.clk(gclk));
	jdff dff_A_CNem8CWd3_2(.dout(w_dff_A_On70pndX7_0),.din(w_dff_A_CNem8CWd3_2),.clk(gclk));
	jdff dff_A_On70pndX7_0(.dout(w_dff_A_hrWcbxEX9_0),.din(w_dff_A_On70pndX7_0),.clk(gclk));
	jdff dff_A_hrWcbxEX9_0(.dout(w_dff_A_D6qH2stF1_0),.din(w_dff_A_hrWcbxEX9_0),.clk(gclk));
	jdff dff_A_D6qH2stF1_0(.dout(w_dff_A_uGb9sllM2_0),.din(w_dff_A_D6qH2stF1_0),.clk(gclk));
	jdff dff_A_uGb9sllM2_0(.dout(w_dff_A_r64SKWGI5_0),.din(w_dff_A_uGb9sllM2_0),.clk(gclk));
	jdff dff_A_r64SKWGI5_0(.dout(G676),.din(w_dff_A_r64SKWGI5_0),.clk(gclk));
	jdff dff_A_rqUWwm8M5_2(.dout(w_dff_A_RVgwCXR00_0),.din(w_dff_A_rqUWwm8M5_2),.clk(gclk));
	jdff dff_A_RVgwCXR00_0(.dout(w_dff_A_7YlJ9mEM7_0),.din(w_dff_A_RVgwCXR00_0),.clk(gclk));
	jdff dff_A_7YlJ9mEM7_0(.dout(w_dff_A_eKUg72am9_0),.din(w_dff_A_7YlJ9mEM7_0),.clk(gclk));
	jdff dff_A_eKUg72am9_0(.dout(w_dff_A_5YzybX6G4_0),.din(w_dff_A_eKUg72am9_0),.clk(gclk));
	jdff dff_A_5YzybX6G4_0(.dout(w_dff_A_YANTPxk09_0),.din(w_dff_A_5YzybX6G4_0),.clk(gclk));
	jdff dff_A_YANTPxk09_0(.dout(w_dff_A_tYg2fACr8_0),.din(w_dff_A_YANTPxk09_0),.clk(gclk));
	jdff dff_A_tYg2fACr8_0(.dout(w_dff_A_GNYJi9ud8_0),.din(w_dff_A_tYg2fACr8_0),.clk(gclk));
	jdff dff_A_GNYJi9ud8_0(.dout(w_dff_A_73A43DHf0_0),.din(w_dff_A_GNYJi9ud8_0),.clk(gclk));
	jdff dff_A_73A43DHf0_0(.dout(w_dff_A_AdDZzCPb6_0),.din(w_dff_A_73A43DHf0_0),.clk(gclk));
	jdff dff_A_AdDZzCPb6_0(.dout(G696),.din(w_dff_A_AdDZzCPb6_0),.clk(gclk));
	jdff dff_A_Wj8inUZF4_2(.dout(w_dff_A_m1ysEKYC5_0),.din(w_dff_A_Wj8inUZF4_2),.clk(gclk));
	jdff dff_A_m1ysEKYC5_0(.dout(w_dff_A_TerU8ija8_0),.din(w_dff_A_m1ysEKYC5_0),.clk(gclk));
	jdff dff_A_TerU8ija8_0(.dout(w_dff_A_fSESxPlQ3_0),.din(w_dff_A_TerU8ija8_0),.clk(gclk));
	jdff dff_A_fSESxPlQ3_0(.dout(w_dff_A_hAhKblHz6_0),.din(w_dff_A_fSESxPlQ3_0),.clk(gclk));
	jdff dff_A_hAhKblHz6_0(.dout(w_dff_A_YhryUOm46_0),.din(w_dff_A_hAhKblHz6_0),.clk(gclk));
	jdff dff_A_YhryUOm46_0(.dout(w_dff_A_rakfXR4h6_0),.din(w_dff_A_YhryUOm46_0),.clk(gclk));
	jdff dff_A_rakfXR4h6_0(.dout(w_dff_A_89qsdqi22_0),.din(w_dff_A_rakfXR4h6_0),.clk(gclk));
	jdff dff_A_89qsdqi22_0(.dout(w_dff_A_bH1RFDNj6_0),.din(w_dff_A_89qsdqi22_0),.clk(gclk));
	jdff dff_A_bH1RFDNj6_0(.dout(w_dff_A_HnHM054f8_0),.din(w_dff_A_bH1RFDNj6_0),.clk(gclk));
	jdff dff_A_HnHM054f8_0(.dout(G699),.din(w_dff_A_HnHM054f8_0),.clk(gclk));
	jdff dff_A_8GjDZDev4_2(.dout(w_dff_A_OUJpiErG8_0),.din(w_dff_A_8GjDZDev4_2),.clk(gclk));
	jdff dff_A_OUJpiErG8_0(.dout(w_dff_A_eK4G8LO80_0),.din(w_dff_A_OUJpiErG8_0),.clk(gclk));
	jdff dff_A_eK4G8LO80_0(.dout(w_dff_A_iHvmmtZ78_0),.din(w_dff_A_eK4G8LO80_0),.clk(gclk));
	jdff dff_A_iHvmmtZ78_0(.dout(w_dff_A_PmvazPgh1_0),.din(w_dff_A_iHvmmtZ78_0),.clk(gclk));
	jdff dff_A_PmvazPgh1_0(.dout(w_dff_A_6CL4psut4_0),.din(w_dff_A_PmvazPgh1_0),.clk(gclk));
	jdff dff_A_6CL4psut4_0(.dout(w_dff_A_ugJeT2CF6_0),.din(w_dff_A_6CL4psut4_0),.clk(gclk));
	jdff dff_A_ugJeT2CF6_0(.dout(w_dff_A_UEELVarc9_0),.din(w_dff_A_ugJeT2CF6_0),.clk(gclk));
	jdff dff_A_UEELVarc9_0(.dout(w_dff_A_nV8OGsFS9_0),.din(w_dff_A_UEELVarc9_0),.clk(gclk));
	jdff dff_A_nV8OGsFS9_0(.dout(G702),.din(w_dff_A_nV8OGsFS9_0),.clk(gclk));
	jdff dff_A_TaBL4Brs2_2(.dout(w_dff_A_aX8uaQA84_0),.din(w_dff_A_TaBL4Brs2_2),.clk(gclk));
	jdff dff_A_aX8uaQA84_0(.dout(w_dff_A_hGewjCFE3_0),.din(w_dff_A_aX8uaQA84_0),.clk(gclk));
	jdff dff_A_hGewjCFE3_0(.dout(w_dff_A_RUnnaiW58_0),.din(w_dff_A_hGewjCFE3_0),.clk(gclk));
	jdff dff_A_RUnnaiW58_0(.dout(w_dff_A_t3nFALht1_0),.din(w_dff_A_RUnnaiW58_0),.clk(gclk));
	jdff dff_A_t3nFALht1_0(.dout(w_dff_A_YoPMJSqe7_0),.din(w_dff_A_t3nFALht1_0),.clk(gclk));
	jdff dff_A_YoPMJSqe7_0(.dout(w_dff_A_l25XVDb49_0),.din(w_dff_A_YoPMJSqe7_0),.clk(gclk));
	jdff dff_A_l25XVDb49_0(.dout(G818),.din(w_dff_A_l25XVDb49_0),.clk(gclk));
	jdff dff_A_8tn0NyFO1_2(.dout(w_dff_A_i4HuO8CL5_0),.din(w_dff_A_8tn0NyFO1_2),.clk(gclk));
	jdff dff_A_i4HuO8CL5_0(.dout(w_dff_A_n3XQRd0k8_0),.din(w_dff_A_i4HuO8CL5_0),.clk(gclk));
	jdff dff_A_n3XQRd0k8_0(.dout(w_dff_A_27NPS7526_0),.din(w_dff_A_n3XQRd0k8_0),.clk(gclk));
	jdff dff_A_27NPS7526_0(.dout(w_dff_A_R4cvzddh6_0),.din(w_dff_A_27NPS7526_0),.clk(gclk));
	jdff dff_A_R4cvzddh6_0(.dout(w_dff_A_g50MpUcu0_0),.din(w_dff_A_R4cvzddh6_0),.clk(gclk));
	jdff dff_A_g50MpUcu0_0(.dout(w_dff_A_p0MuONXz7_0),.din(w_dff_A_g50MpUcu0_0),.clk(gclk));
	jdff dff_A_p0MuONXz7_0(.dout(w_dff_A_lngJ7pm18_0),.din(w_dff_A_p0MuONXz7_0),.clk(gclk));
	jdff dff_A_lngJ7pm18_0(.dout(w_dff_A_wsb8YRE63_0),.din(w_dff_A_lngJ7pm18_0),.clk(gclk));
	jdff dff_A_wsb8YRE63_0(.dout(w_dff_A_04KwKPAI3_0),.din(w_dff_A_wsb8YRE63_0),.clk(gclk));
	jdff dff_A_04KwKPAI3_0(.dout(G813),.din(w_dff_A_04KwKPAI3_0),.clk(gclk));
	jdff dff_A_qGyy1NWt1_1(.dout(w_dff_A_9udiq8sW3_0),.din(w_dff_A_qGyy1NWt1_1),.clk(gclk));
	jdff dff_A_9udiq8sW3_0(.dout(w_dff_A_TeoSuiwr3_0),.din(w_dff_A_9udiq8sW3_0),.clk(gclk));
	jdff dff_A_TeoSuiwr3_0(.dout(w_dff_A_ThNxRt8K2_0),.din(w_dff_A_TeoSuiwr3_0),.clk(gclk));
	jdff dff_A_ThNxRt8K2_0(.dout(w_dff_A_QN73JLJy3_0),.din(w_dff_A_ThNxRt8K2_0),.clk(gclk));
	jdff dff_A_QN73JLJy3_0(.dout(w_dff_A_IUXEYW0j0_0),.din(w_dff_A_QN73JLJy3_0),.clk(gclk));
	jdff dff_A_IUXEYW0j0_0(.dout(w_dff_A_AUdd2RtT1_0),.din(w_dff_A_IUXEYW0j0_0),.clk(gclk));
	jdff dff_A_AUdd2RtT1_0(.dout(G824),.din(w_dff_A_AUdd2RtT1_0),.clk(gclk));
	jdff dff_A_EVE9Od673_1(.dout(w_dff_A_IBGsDboQ8_0),.din(w_dff_A_EVE9Od673_1),.clk(gclk));
	jdff dff_A_IBGsDboQ8_0(.dout(w_dff_A_V5Kd3ZdL7_0),.din(w_dff_A_IBGsDboQ8_0),.clk(gclk));
	jdff dff_A_V5Kd3ZdL7_0(.dout(w_dff_A_P6oYNQt77_0),.din(w_dff_A_V5Kd3ZdL7_0),.clk(gclk));
	jdff dff_A_P6oYNQt77_0(.dout(w_dff_A_WAYN5J1M7_0),.din(w_dff_A_P6oYNQt77_0),.clk(gclk));
	jdff dff_A_WAYN5J1M7_0(.dout(w_dff_A_EIHCPb6O5_0),.din(w_dff_A_WAYN5J1M7_0),.clk(gclk));
	jdff dff_A_EIHCPb6O5_0(.dout(w_dff_A_n8bX5quK9_0),.din(w_dff_A_EIHCPb6O5_0),.clk(gclk));
	jdff dff_A_n8bX5quK9_0(.dout(w_dff_A_D04dZ3iq8_0),.din(w_dff_A_n8bX5quK9_0),.clk(gclk));
	jdff dff_A_D04dZ3iq8_0(.dout(G826),.din(w_dff_A_D04dZ3iq8_0),.clk(gclk));
	jdff dff_A_vpYvFGV21_1(.dout(w_dff_A_7d1GtTVh1_0),.din(w_dff_A_vpYvFGV21_1),.clk(gclk));
	jdff dff_A_7d1GtTVh1_0(.dout(w_dff_A_g1BN4ShE0_0),.din(w_dff_A_7d1GtTVh1_0),.clk(gclk));
	jdff dff_A_g1BN4ShE0_0(.dout(w_dff_A_mHCZCoet1_0),.din(w_dff_A_g1BN4ShE0_0),.clk(gclk));
	jdff dff_A_mHCZCoet1_0(.dout(w_dff_A_hR5TQsUY8_0),.din(w_dff_A_mHCZCoet1_0),.clk(gclk));
	jdff dff_A_hR5TQsUY8_0(.dout(w_dff_A_YszCFn920_0),.din(w_dff_A_hR5TQsUY8_0),.clk(gclk));
	jdff dff_A_YszCFn920_0(.dout(w_dff_A_UsZQS2zR0_0),.din(w_dff_A_YszCFn920_0),.clk(gclk));
	jdff dff_A_UsZQS2zR0_0(.dout(G828),.din(w_dff_A_UsZQS2zR0_0),.clk(gclk));
	jdff dff_A_CpoHOeGU4_1(.dout(w_dff_A_40UM4Gm46_0),.din(w_dff_A_CpoHOeGU4_1),.clk(gclk));
	jdff dff_A_40UM4Gm46_0(.dout(w_dff_A_Gn1N5gGs0_0),.din(w_dff_A_40UM4Gm46_0),.clk(gclk));
	jdff dff_A_Gn1N5gGs0_0(.dout(w_dff_A_aTlV2qug6_0),.din(w_dff_A_Gn1N5gGs0_0),.clk(gclk));
	jdff dff_A_aTlV2qug6_0(.dout(w_dff_A_6LA6kV310_0),.din(w_dff_A_aTlV2qug6_0),.clk(gclk));
	jdff dff_A_6LA6kV310_0(.dout(w_dff_A_vIdbinNX7_0),.din(w_dff_A_6LA6kV310_0),.clk(gclk));
	jdff dff_A_vIdbinNX7_0(.dout(w_dff_A_Y0LvZxw86_0),.din(w_dff_A_vIdbinNX7_0),.clk(gclk));
	jdff dff_A_Y0LvZxw86_0(.dout(w_dff_A_og5PqnC33_0),.din(w_dff_A_Y0LvZxw86_0),.clk(gclk));
	jdff dff_A_og5PqnC33_0(.dout(w_dff_A_tquKRHqe5_0),.din(w_dff_A_og5PqnC33_0),.clk(gclk));
	jdff dff_A_tquKRHqe5_0(.dout(w_dff_A_7AvzbBGl1_0),.din(w_dff_A_tquKRHqe5_0),.clk(gclk));
	jdff dff_A_7AvzbBGl1_0(.dout(w_dff_A_NrDadm585_0),.din(w_dff_A_7AvzbBGl1_0),.clk(gclk));
	jdff dff_A_NrDadm585_0(.dout(w_dff_A_zEMcQFle9_0),.din(w_dff_A_NrDadm585_0),.clk(gclk));
	jdff dff_A_zEMcQFle9_0(.dout(G830),.din(w_dff_A_zEMcQFle9_0),.clk(gclk));
	jdff dff_A_HFgIIjdN5_2(.dout(w_dff_A_ooiQQtaX5_0),.din(w_dff_A_HFgIIjdN5_2),.clk(gclk));
	jdff dff_A_ooiQQtaX5_0(.dout(w_dff_A_1qbW3D1c9_0),.din(w_dff_A_ooiQQtaX5_0),.clk(gclk));
	jdff dff_A_1qbW3D1c9_0(.dout(w_dff_A_G3PhFWIu5_0),.din(w_dff_A_1qbW3D1c9_0),.clk(gclk));
	jdff dff_A_G3PhFWIu5_0(.dout(w_dff_A_cG5ObuCm2_0),.din(w_dff_A_G3PhFWIu5_0),.clk(gclk));
	jdff dff_A_cG5ObuCm2_0(.dout(w_dff_A_v6BqUteU5_0),.din(w_dff_A_cG5ObuCm2_0),.clk(gclk));
	jdff dff_A_v6BqUteU5_0(.dout(w_dff_A_kiQ5mfNK6_0),.din(w_dff_A_v6BqUteU5_0),.clk(gclk));
	jdff dff_A_kiQ5mfNK6_0(.dout(w_dff_A_NQN3EwPf8_0),.din(w_dff_A_kiQ5mfNK6_0),.clk(gclk));
	jdff dff_A_NQN3EwPf8_0(.dout(w_dff_A_WsOyHbMF3_0),.din(w_dff_A_NQN3EwPf8_0),.clk(gclk));
	jdff dff_A_WsOyHbMF3_0(.dout(w_dff_A_lEq7x3RI4_0),.din(w_dff_A_WsOyHbMF3_0),.clk(gclk));
	jdff dff_A_lEq7x3RI4_0(.dout(w_dff_A_coaJiB730_0),.din(w_dff_A_lEq7x3RI4_0),.clk(gclk));
	jdff dff_A_coaJiB730_0(.dout(w_dff_A_e1piiQAt9_0),.din(w_dff_A_coaJiB730_0),.clk(gclk));
	jdff dff_A_e1piiQAt9_0(.dout(w_dff_A_G3wm3Dk56_0),.din(w_dff_A_e1piiQAt9_0),.clk(gclk));
	jdff dff_A_G3wm3Dk56_0(.dout(w_dff_A_iXpnZ5X21_0),.din(w_dff_A_G3wm3Dk56_0),.clk(gclk));
	jdff dff_A_iXpnZ5X21_0(.dout(w_dff_A_cq8gQ2nO1_0),.din(w_dff_A_iXpnZ5X21_0),.clk(gclk));
	jdff dff_A_cq8gQ2nO1_0(.dout(w_dff_A_pwfMFyjE5_0),.din(w_dff_A_cq8gQ2nO1_0),.clk(gclk));
	jdff dff_A_pwfMFyjE5_0(.dout(w_dff_A_bz3TO0ZZ9_0),.din(w_dff_A_pwfMFyjE5_0),.clk(gclk));
	jdff dff_A_bz3TO0ZZ9_0(.dout(G854),.din(w_dff_A_bz3TO0ZZ9_0),.clk(gclk));
	jdff dff_A_TarUmmSU2_1(.dout(w_dff_A_LCwyfpbh4_0),.din(w_dff_A_TarUmmSU2_1),.clk(gclk));
	jdff dff_A_LCwyfpbh4_0(.dout(w_dff_A_BbQD3Zps0_0),.din(w_dff_A_LCwyfpbh4_0),.clk(gclk));
	jdff dff_A_BbQD3Zps0_0(.dout(w_dff_A_GRlkehMQ9_0),.din(w_dff_A_BbQD3Zps0_0),.clk(gclk));
	jdff dff_A_GRlkehMQ9_0(.dout(w_dff_A_YfJci39l0_0),.din(w_dff_A_GRlkehMQ9_0),.clk(gclk));
	jdff dff_A_YfJci39l0_0(.dout(w_dff_A_FGag6nlK5_0),.din(w_dff_A_YfJci39l0_0),.clk(gclk));
	jdff dff_A_FGag6nlK5_0(.dout(G863),.din(w_dff_A_FGag6nlK5_0),.clk(gclk));
	jdff dff_A_bx1a0Rhg8_1(.dout(w_dff_A_qDFT43pG4_0),.din(w_dff_A_bx1a0Rhg8_1),.clk(gclk));
	jdff dff_A_qDFT43pG4_0(.dout(w_dff_A_4gLWta1w7_0),.din(w_dff_A_qDFT43pG4_0),.clk(gclk));
	jdff dff_A_4gLWta1w7_0(.dout(w_dff_A_K2ccRX827_0),.din(w_dff_A_4gLWta1w7_0),.clk(gclk));
	jdff dff_A_K2ccRX827_0(.dout(w_dff_A_quagDw2X3_0),.din(w_dff_A_K2ccRX827_0),.clk(gclk));
	jdff dff_A_quagDw2X3_0(.dout(w_dff_A_YQJEdmnT2_0),.din(w_dff_A_quagDw2X3_0),.clk(gclk));
	jdff dff_A_YQJEdmnT2_0(.dout(w_dff_A_ax7oc2fh9_0),.din(w_dff_A_YQJEdmnT2_0),.clk(gclk));
	jdff dff_A_ax7oc2fh9_0(.dout(w_dff_A_XNWDjkFu4_0),.din(w_dff_A_ax7oc2fh9_0),.clk(gclk));
	jdff dff_A_XNWDjkFu4_0(.dout(w_dff_A_jlqeiFKW9_0),.din(w_dff_A_XNWDjkFu4_0),.clk(gclk));
	jdff dff_A_jlqeiFKW9_0(.dout(G865),.din(w_dff_A_jlqeiFKW9_0),.clk(gclk));
	jdff dff_A_mmpAPBTa5_1(.dout(w_dff_A_0KVkXGpU7_0),.din(w_dff_A_mmpAPBTa5_1),.clk(gclk));
	jdff dff_A_0KVkXGpU7_0(.dout(w_dff_A_cciaEVbv3_0),.din(w_dff_A_0KVkXGpU7_0),.clk(gclk));
	jdff dff_A_cciaEVbv3_0(.dout(w_dff_A_ujBfOO7C9_0),.din(w_dff_A_cciaEVbv3_0),.clk(gclk));
	jdff dff_A_ujBfOO7C9_0(.dout(w_dff_A_yNfjHOCH1_0),.din(w_dff_A_ujBfOO7C9_0),.clk(gclk));
	jdff dff_A_yNfjHOCH1_0(.dout(w_dff_A_p4NjGlo98_0),.din(w_dff_A_yNfjHOCH1_0),.clk(gclk));
	jdff dff_A_p4NjGlo98_0(.dout(w_dff_A_phV0KFNN6_0),.din(w_dff_A_p4NjGlo98_0),.clk(gclk));
	jdff dff_A_phV0KFNN6_0(.dout(G867),.din(w_dff_A_phV0KFNN6_0),.clk(gclk));
	jdff dff_A_2o5mNUNN0_1(.dout(w_dff_A_xbvKmbTE9_0),.din(w_dff_A_2o5mNUNN0_1),.clk(gclk));
	jdff dff_A_xbvKmbTE9_0(.dout(w_dff_A_f6RXQBsj0_0),.din(w_dff_A_xbvKmbTE9_0),.clk(gclk));
	jdff dff_A_f6RXQBsj0_0(.dout(w_dff_A_7i8SECPA4_0),.din(w_dff_A_f6RXQBsj0_0),.clk(gclk));
	jdff dff_A_7i8SECPA4_0(.dout(w_dff_A_fLEa04VA1_0),.din(w_dff_A_7i8SECPA4_0),.clk(gclk));
	jdff dff_A_fLEa04VA1_0(.dout(w_dff_A_U9mEhFMP1_0),.din(w_dff_A_fLEa04VA1_0),.clk(gclk));
	jdff dff_A_U9mEhFMP1_0(.dout(w_dff_A_SiaW7h2d5_0),.din(w_dff_A_U9mEhFMP1_0),.clk(gclk));
	jdff dff_A_SiaW7h2d5_0(.dout(w_dff_A_LIXYn4HD6_0),.din(w_dff_A_SiaW7h2d5_0),.clk(gclk));
	jdff dff_A_LIXYn4HD6_0(.dout(w_dff_A_d8ELLy8O1_0),.din(w_dff_A_LIXYn4HD6_0),.clk(gclk));
	jdff dff_A_d8ELLy8O1_0(.dout(w_dff_A_dkTqBuXF4_0),.din(w_dff_A_d8ELLy8O1_0),.clk(gclk));
	jdff dff_A_dkTqBuXF4_0(.dout(G869),.din(w_dff_A_dkTqBuXF4_0),.clk(gclk));
	jdff dff_A_dkFs5zUM9_2(.dout(w_dff_A_9KNRyLUd4_0),.din(w_dff_A_dkFs5zUM9_2),.clk(gclk));
	jdff dff_A_9KNRyLUd4_0(.dout(w_dff_A_06QcdIBx6_0),.din(w_dff_A_9KNRyLUd4_0),.clk(gclk));
	jdff dff_A_06QcdIBx6_0(.dout(w_dff_A_GsRwyzkb8_0),.din(w_dff_A_06QcdIBx6_0),.clk(gclk));
	jdff dff_A_GsRwyzkb8_0(.dout(G712),.din(w_dff_A_GsRwyzkb8_0),.clk(gclk));
	jdff dff_A_xn8VXQlt9_2(.dout(w_dff_A_rMDzb1GG3_0),.din(w_dff_A_xn8VXQlt9_2),.clk(gclk));
	jdff dff_A_rMDzb1GG3_0(.dout(w_dff_A_QLjD2Cn63_0),.din(w_dff_A_rMDzb1GG3_0),.clk(gclk));
	jdff dff_A_QLjD2Cn63_0(.dout(G727),.din(w_dff_A_QLjD2Cn63_0),.clk(gclk));
	jdff dff_A_ThgarqCR8_2(.dout(w_dff_A_qysuLA4i7_0),.din(w_dff_A_ThgarqCR8_2),.clk(gclk));
	jdff dff_A_qysuLA4i7_0(.dout(w_dff_A_yDzih88r6_0),.din(w_dff_A_qysuLA4i7_0),.clk(gclk));
	jdff dff_A_yDzih88r6_0(.dout(w_dff_A_FcZtCV8G2_0),.din(w_dff_A_yDzih88r6_0),.clk(gclk));
	jdff dff_A_FcZtCV8G2_0(.dout(G732),.din(w_dff_A_FcZtCV8G2_0),.clk(gclk));
	jdff dff_A_iLcxeVf72_2(.dout(w_dff_A_f5FTN0vF7_0),.din(w_dff_A_iLcxeVf72_2),.clk(gclk));
	jdff dff_A_f5FTN0vF7_0(.dout(w_dff_A_tQEcwiIb0_0),.din(w_dff_A_f5FTN0vF7_0),.clk(gclk));
	jdff dff_A_tQEcwiIb0_0(.dout(w_dff_A_B8Yf720Y3_0),.din(w_dff_A_tQEcwiIb0_0),.clk(gclk));
	jdff dff_A_B8Yf720Y3_0(.dout(G737),.din(w_dff_A_B8Yf720Y3_0),.clk(gclk));
	jdff dff_A_VciU7eAY5_2(.dout(w_dff_A_T84PciTu9_0),.din(w_dff_A_VciU7eAY5_2),.clk(gclk));
	jdff dff_A_T84PciTu9_0(.dout(w_dff_A_9JuzTgrz0_0),.din(w_dff_A_T84PciTu9_0),.clk(gclk));
	jdff dff_A_9JuzTgrz0_0(.dout(w_dff_A_9NOqxWAq6_0),.din(w_dff_A_9JuzTgrz0_0),.clk(gclk));
	jdff dff_A_9NOqxWAq6_0(.dout(w_dff_A_VaDNWgO74_0),.din(w_dff_A_9NOqxWAq6_0),.clk(gclk));
	jdff dff_A_VaDNWgO74_0(.dout(G742),.din(w_dff_A_VaDNWgO74_0),.clk(gclk));
	jdff dff_A_iVCTOc7f1_2(.dout(w_dff_A_EIppLBGv6_0),.din(w_dff_A_iVCTOc7f1_2),.clk(gclk));
	jdff dff_A_EIppLBGv6_0(.dout(w_dff_A_tG2R1g567_0),.din(w_dff_A_EIppLBGv6_0),.clk(gclk));
	jdff dff_A_tG2R1g567_0(.dout(w_dff_A_Hb80b2Iz1_0),.din(w_dff_A_tG2R1g567_0),.clk(gclk));
	jdff dff_A_Hb80b2Iz1_0(.dout(G772),.din(w_dff_A_Hb80b2Iz1_0),.clk(gclk));
	jdff dff_A_QaYaxUiX3_2(.dout(w_dff_A_3MJ5qlH03_0),.din(w_dff_A_QaYaxUiX3_2),.clk(gclk));
	jdff dff_A_3MJ5qlH03_0(.dout(w_dff_A_faciHVZ36_0),.din(w_dff_A_3MJ5qlH03_0),.clk(gclk));
	jdff dff_A_faciHVZ36_0(.dout(w_dff_A_db1yODmM4_0),.din(w_dff_A_faciHVZ36_0),.clk(gclk));
	jdff dff_A_db1yODmM4_0(.dout(G777),.din(w_dff_A_db1yODmM4_0),.clk(gclk));
	jdff dff_A_ukNOl0VY4_2(.dout(w_dff_A_7YO21lXD0_0),.din(w_dff_A_ukNOl0VY4_2),.clk(gclk));
	jdff dff_A_7YO21lXD0_0(.dout(w_dff_A_ubVsCTJd9_0),.din(w_dff_A_7YO21lXD0_0),.clk(gclk));
	jdff dff_A_ubVsCTJd9_0(.dout(w_dff_A_cdz5R05I0_0),.din(w_dff_A_ubVsCTJd9_0),.clk(gclk));
	jdff dff_A_cdz5R05I0_0(.dout(w_dff_A_zJeWIyi92_0),.din(w_dff_A_cdz5R05I0_0),.clk(gclk));
	jdff dff_A_zJeWIyi92_0(.dout(G782),.din(w_dff_A_zJeWIyi92_0),.clk(gclk));
	jdff dff_A_OlaI97sX7_2(.dout(w_dff_A_S58ioXd06_0),.din(w_dff_A_OlaI97sX7_2),.clk(gclk));
	jdff dff_A_S58ioXd06_0(.dout(w_dff_A_7JwnNXlg0_0),.din(w_dff_A_S58ioXd06_0),.clk(gclk));
	jdff dff_A_7JwnNXlg0_0(.dout(w_dff_A_hA4dvUqD0_0),.din(w_dff_A_7JwnNXlg0_0),.clk(gclk));
	jdff dff_A_hA4dvUqD0_0(.dout(G645),.din(w_dff_A_hA4dvUqD0_0),.clk(gclk));
	jdff dff_A_TBsLnPUK2_2(.dout(w_dff_A_RgdYOw2L6_0),.din(w_dff_A_TBsLnPUK2_2),.clk(gclk));
	jdff dff_A_RgdYOw2L6_0(.dout(w_dff_A_iCXl4u621_0),.din(w_dff_A_RgdYOw2L6_0),.clk(gclk));
	jdff dff_A_iCXl4u621_0(.dout(G648),.din(w_dff_A_iCXl4u621_0),.clk(gclk));
	jdff dff_A_dzvMNPTC6_2(.dout(w_dff_A_B3NYq2Fm8_0),.din(w_dff_A_dzvMNPTC6_2),.clk(gclk));
	jdff dff_A_B3NYq2Fm8_0(.dout(w_dff_A_cTWeL9db5_0),.din(w_dff_A_B3NYq2Fm8_0),.clk(gclk));
	jdff dff_A_cTWeL9db5_0(.dout(G651),.din(w_dff_A_cTWeL9db5_0),.clk(gclk));
	jdff dff_A_NOl4MacD3_2(.dout(w_dff_A_MbvSoAG75_0),.din(w_dff_A_NOl4MacD3_2),.clk(gclk));
	jdff dff_A_MbvSoAG75_0(.dout(G654),.din(w_dff_A_MbvSoAG75_0),.clk(gclk));
	jdff dff_A_Udi9HLES1_2(.dout(w_dff_A_WL61JqNm2_0),.din(w_dff_A_Udi9HLES1_2),.clk(gclk));
	jdff dff_A_WL61JqNm2_0(.dout(w_dff_A_UrviIedY4_0),.din(w_dff_A_WL61JqNm2_0),.clk(gclk));
	jdff dff_A_UrviIedY4_0(.dout(w_dff_A_rrSdEsv22_0),.din(w_dff_A_UrviIedY4_0),.clk(gclk));
	jdff dff_A_rrSdEsv22_0(.dout(G679),.din(w_dff_A_rrSdEsv22_0),.clk(gclk));
	jdff dff_A_CXlZvC9V9_2(.dout(w_dff_A_ig96CRdK0_0),.din(w_dff_A_CXlZvC9V9_2),.clk(gclk));
	jdff dff_A_ig96CRdK0_0(.dout(w_dff_A_SWrQAXbD7_0),.din(w_dff_A_ig96CRdK0_0),.clk(gclk));
	jdff dff_A_SWrQAXbD7_0(.dout(G682),.din(w_dff_A_SWrQAXbD7_0),.clk(gclk));
	jdff dff_A_jSG9y9fp6_2(.dout(w_dff_A_59OFn7UG6_0),.din(w_dff_A_jSG9y9fp6_2),.clk(gclk));
	jdff dff_A_59OFn7UG6_0(.dout(w_dff_A_FIXTm6cC6_0),.din(w_dff_A_59OFn7UG6_0),.clk(gclk));
	jdff dff_A_FIXTm6cC6_0(.dout(G685),.din(w_dff_A_FIXTm6cC6_0),.clk(gclk));
	jdff dff_A_xHbVfs0P9_2(.dout(w_dff_A_WA0UNGcW0_0),.din(w_dff_A_xHbVfs0P9_2),.clk(gclk));
	jdff dff_A_WA0UNGcW0_0(.dout(w_dff_A_2QiH6WY53_0),.din(w_dff_A_WA0UNGcW0_0),.clk(gclk));
	jdff dff_A_2QiH6WY53_0(.dout(G688),.din(w_dff_A_2QiH6WY53_0),.clk(gclk));
	jdff dff_A_YSK6IrZh6_2(.dout(w_dff_A_JLlRlcw25_0),.din(w_dff_A_YSK6IrZh6_2),.clk(gclk));
	jdff dff_A_JLlRlcw25_0(.dout(w_dff_A_cr7Vl9ua8_0),.din(w_dff_A_JLlRlcw25_0),.clk(gclk));
	jdff dff_A_cr7Vl9ua8_0(.dout(w_dff_A_iMYy5M7z7_0),.din(w_dff_A_cr7Vl9ua8_0),.clk(gclk));
	jdff dff_A_iMYy5M7z7_0(.dout(w_dff_A_75L5Xd0x9_0),.din(w_dff_A_iMYy5M7z7_0),.clk(gclk));
	jdff dff_A_75L5Xd0x9_0(.dout(w_dff_A_FsBNdA3J3_0),.din(w_dff_A_75L5Xd0x9_0),.clk(gclk));
	jdff dff_A_FsBNdA3J3_0(.dout(G843),.din(w_dff_A_FsBNdA3J3_0),.clk(gclk));
	jdff dff_A_vmfcvb7t4_2(.dout(w_dff_A_ZQ3ej7MJ4_0),.din(w_dff_A_vmfcvb7t4_2),.clk(gclk));
	jdff dff_A_ZQ3ej7MJ4_0(.dout(w_dff_A_m9uFebf27_0),.din(w_dff_A_ZQ3ej7MJ4_0),.clk(gclk));
	jdff dff_A_m9uFebf27_0(.dout(w_dff_A_8opvLAEc3_0),.din(w_dff_A_m9uFebf27_0),.clk(gclk));
	jdff dff_A_8opvLAEc3_0(.dout(w_dff_A_CzW6VcWB6_0),.din(w_dff_A_8opvLAEc3_0),.clk(gclk));
	jdff dff_A_CzW6VcWB6_0(.dout(w_dff_A_8ZbA5KkE6_0),.din(w_dff_A_CzW6VcWB6_0),.clk(gclk));
	jdff dff_A_8ZbA5KkE6_0(.dout(G882),.din(w_dff_A_8ZbA5KkE6_0),.clk(gclk));
	jdff dff_A_RE0tB8YO4_2(.dout(G767),.din(w_dff_A_RE0tB8YO4_2),.clk(gclk));
	jdff dff_A_pwFU8BN14_2(.dout(G807),.din(w_dff_A_pwFU8BN14_2),.clk(gclk));
endmodule

