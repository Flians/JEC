/*

c432:
	jxor: 1
	jspl: 84
	jspl3: 48
	jnot: 47
	jdff: 340
	jand: 104
	jor: 104

Summary:
	jxor: 1
	jspl: 84
	jspl3: 48
	jnot: 47
	jdff: 340
	jand: 104
	jor: 104

The maximum logic level gap of any gate:
	c432: 7
*/

module gf_c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n43;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G4gat_0;
	wire[2:0] w_G8gat_0;
	wire[2:0] w_G11gat_0;
	wire[2:0] w_G14gat_0;
	wire[2:0] w_G17gat_0;
	wire[2:0] w_G21gat_0;
	wire[2:0] w_G24gat_0;
	wire[1:0] w_G27gat_0;
	wire[2:0] w_G30gat_0;
	wire[2:0] w_G34gat_0;
	wire[1:0] w_G40gat_0;
	wire[1:0] w_G43gat_0;
	wire[2:0] w_G47gat_0;
	wire[1:0] w_G50gat_0;
	wire[1:0] w_G53gat_0;
	wire[2:0] w_G56gat_0;
	wire[1:0] w_G56gat_1;
	wire[1:0] w_G60gat_0;
	wire[2:0] w_G63gat_0;
	wire[2:0] w_G66gat_0;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G73gat_0;
	wire[2:0] w_G76gat_0;
	wire[1:0] w_G79gat_0;
	wire[2:0] w_G82gat_0;
	wire[2:0] w_G86gat_0;
	wire[2:0] w_G89gat_0;
	wire[2:0] w_G92gat_0;
	wire[2:0] w_G95gat_0;
	wire[2:0] w_G99gat_0;
	wire[1:0] w_G102gat_0;
	wire[1:0] w_G105gat_0;
	wire[2:0] w_G108gat_0;
	wire[2:0] w_G112gat_0;
	wire[1:0] w_G115gat_0;
	wire[2:0] w_G223gat_0;
	wire[2:0] w_G223gat_1;
	wire[2:0] w_G223gat_2;
	wire[2:0] w_G223gat_3;
	wire w_G223gat_4;
	wire G223gat_fa_;
	wire[2:0] w_G329gat_0;
	wire[2:0] w_G329gat_1;
	wire[2:0] w_G329gat_2;
	wire[2:0] w_G329gat_3;
	wire w_G329gat_4;
	wire G329gat_fa_;
	wire[2:0] w_G370gat_0;
	wire[1:0] w_G370gat_1;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire[1:0] w_n43_0;
	wire[1:0] w_n44_0;
	wire[1:0] w_n45_0;
	wire[2:0] w_n46_0;
	wire[1:0] w_n47_0;
	wire[1:0] w_n49_0;
	wire[1:0] w_n51_0;
	wire[1:0] w_n54_0;
	wire[1:0] w_n57_0;
	wire[1:0] w_n60_0;
	wire[1:0] w_n62_0;
	wire[1:0] w_n64_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n73_0;
	wire[1:0] w_n75_0;
	wire[1:0] w_n78_0;
	wire[1:0] w_n80_0;
	wire[1:0] w_n81_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[1:0] w_n88_0;
	wire[2:0] w_n93_0;
	wire[2:0] w_n93_1;
	wire[2:0] w_n93_2;
	wire[2:0] w_n93_3;
	wire[1:0] w_n95_0;
	wire[1:0] w_n102_0;
	wire[1:0] w_n104_0;
	wire[1:0] w_n106_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n111_0;
	wire[1:0] w_n113_0;
	wire[1:0] w_n117_0;
	wire[2:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[1:0] w_n121_0;
	wire[1:0] w_n123_0;
	wire[1:0] w_n125_0;
	wire[1:0] w_n127_0;
	wire[2:0] w_n131_0;
	wire[1:0] w_n138_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n141_0;
	wire[1:0] w_n144_0;
	wire[1:0] w_n145_0;
	wire[1:0] w_n147_0;
	wire[1:0] w_n149_0;
	wire[1:0] w_n151_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n159_0;
	wire[1:0] w_n164_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n173_0;
	wire[2:0] w_n181_0;
	wire[2:0] w_n181_1;
	wire[2:0] w_n181_2;
	wire[1:0] w_n183_0;
	wire[1:0] w_n185_0;
	wire[1:0] w_n200_0;
	wire[1:0] w_n202_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n209_0;
	wire[1:0] w_n211_0;
	wire[1:0] w_n222_0;
	wire[1:0] w_n227_0;
	wire[1:0] w_n230_0;
	wire[2:0] w_n246_0;
	wire[2:0] w_n246_1;
	wire[2:0] w_n246_2;
	wire[1:0] w_n248_0;
	wire[1:0] w_n250_0;
	wire[1:0] w_n251_0;
	wire[1:0] w_n253_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n257_0;
	wire[1:0] w_n264_0;
	wire[1:0] w_n265_0;
	wire[1:0] w_n269_0;
	wire[1:0] w_n271_0;
	wire[1:0] w_n281_0;
	wire[1:0] w_n288_0;
	wire[1:0] w_n290_0;
	wire w_dff_B_TUGn5viz4_0;
	wire w_dff_B_tG6glVm67_0;
	wire w_dff_B_VHlRVsXk8_0;
	wire w_dff_B_3PqJqlKa2_0;
	wire w_dff_B_5mbO5f7u4_0;
	wire w_dff_B_RHpznR979_0;
	wire w_dff_B_gfFb8n1K8_0;
	wire w_dff_B_djEVmgys0_0;
	wire w_dff_B_haVkYUuq3_0;
	wire w_dff_B_3sV01tN74_2;
	wire w_dff_A_UHkQgKLo7_0;
	wire w_dff_B_FlrqaWjo7_2;
	wire w_dff_A_4ZGDBSoA9_1;
	wire w_dff_B_93W8t1sd2_1;
	wire w_dff_B_JqKvAV603_1;
	wire w_dff_B_AfVnNhxM8_1;
	wire w_dff_B_nwJrN7zD5_1;
	wire w_dff_B_jGLnkveQ9_1;
	wire w_dff_B_kXx7g4k74_1;
	wire w_dff_B_nSLP0dXm0_1;
	wire w_dff_B_XljKjWDk9_1;
	wire w_dff_B_qv6pQL5z4_1;
	wire w_dff_B_Dz4jzG8q1_1;
	wire w_dff_B_5MUvVNGe7_1;
	wire w_dff_B_5opjKqlz4_1;
	wire w_dff_B_Chl8E2SN0_1;
	wire w_dff_B_0b0j6Mz34_1;
	wire w_dff_B_3552XGda2_1;
	wire w_dff_B_6dsNo7H12_1;
	wire w_dff_B_dSzDWF9f1_1;
	wire w_dff_B_ZYhtOIYc2_1;
	wire w_dff_B_BsagiSh45_1;
	wire w_dff_B_3682yVZD5_1;
	wire w_dff_B_00FgM2Us0_1;
	wire w_dff_B_X0KPIGTs9_1;
	wire w_dff_B_0vHgPdV99_1;
	wire w_dff_B_OjPKiWFI0_1;
	wire w_dff_B_sD7gCxad0_2;
	wire w_dff_A_vHQ7tY2m1_0;
	wire w_dff_A_OWCEaoKo1_0;
	wire w_dff_A_kXafuMAw3_0;
	wire w_dff_B_aiwcWzfd6_1;
	wire w_dff_A_rF4bOhRf9_0;
	wire w_dff_A_OU0O9T7b6_0;
	wire w_dff_A_28gX06vb9_0;
	wire w_dff_A_fl6lqKnc0_0;
	wire w_dff_A_yCH6Anye4_0;
	wire w_dff_A_vcKH6jI99_0;
	wire w_dff_B_xSd0xNja4_1;
	wire w_dff_B_vdGQaMzM1_1;
	wire w_dff_B_fD9aqSh78_1;
	wire w_dff_B_Pgl1Z3jn0_1;
	wire w_dff_B_X6jdc4lQ9_1;
	wire w_dff_B_TpjrsyKd5_1;
	wire w_dff_B_lXsBvo7M9_1;
	wire w_dff_B_yHMnvESC0_0;
	wire w_dff_B_zsKn8oIK0_0;
	wire w_dff_B_j9aclB070_0;
	wire w_dff_B_MJ3zYHxJ4_0;
	wire w_dff_A_TBysbvAN3_1;
	wire w_dff_A_EkcHTEVP3_1;
	wire w_dff_A_f6EYMW6q4_1;
	wire w_dff_A_uKSJ0XJD1_1;
	wire w_dff_A_YeVc5UOD3_1;
	wire w_dff_B_lwXOQWpt6_1;
	wire w_dff_B_QP2GGXYy0_0;
	wire w_dff_A_u0cATR1T7_0;
	wire w_dff_A_ImyC5g2F8_0;
	wire w_dff_A_vMrf8DEo2_0;
	wire w_dff_A_UUKWveyy9_0;
	wire w_dff_A_k72FSdyG6_0;
	wire w_dff_A_yja1jA0G3_0;
	wire w_dff_A_xpBVrZqa7_0;
	wire w_dff_A_9Oa7IXWv2_0;
	wire w_dff_A_oYOZjsMc3_0;
	wire w_dff_A_3BB9E95F3_0;
	wire w_dff_A_UiOlqUe47_0;
	wire w_dff_B_oB8hc8ck0_2;
	wire w_dff_B_EnUAYsxq2_2;
	wire w_dff_B_RCcX7fqy0_2;
	wire w_dff_B_JSIR8IyY8_2;
	wire w_dff_B_oyNdbX3W0_2;
	wire w_dff_B_FhvYs9X27_2;
	wire w_dff_B_j2r1NXJu1_2;
	wire w_dff_B_MUJwKZYJ3_2;
	wire w_dff_B_0W3BZIxm2_2;
	wire w_dff_B_RW7WA03W4_2;
	wire w_dff_B_RIqo5qxR1_2;
	wire w_dff_B_nG7Wb0xO8_2;
	wire w_dff_B_sDsCO4mc0_2;
	wire w_dff_B_6RajPZ225_2;
	wire w_dff_A_QQWtvWjU9_0;
	wire w_dff_A_wByZYIIs9_0;
	wire w_dff_A_TPdwe9sJ7_0;
	wire w_dff_A_QdplOECX8_0;
	wire w_dff_A_iK6c3yTo1_0;
	wire w_dff_A_vZXliEu80_0;
	wire w_dff_A_nfzWIevA8_0;
	wire w_dff_A_Gt0gk1ij9_0;
	wire w_dff_A_v25vqoHc5_0;
	wire w_dff_A_jyvsJMA14_0;
	wire w_dff_A_OYZRaIO26_0;
	wire w_dff_B_9SOwJs438_2;
	wire w_dff_B_4pVfDyK01_2;
	wire w_dff_B_LYcO2Dkx2_2;
	wire w_dff_B_jskmvLJw5_2;
	wire w_dff_B_mkvCYlCP0_2;
	wire w_dff_B_b28DU7yA4_2;
	wire w_dff_B_44SDUm2A6_2;
	wire w_dff_B_fH9OvtBY1_2;
	wire w_dff_B_jDSVQKhW6_2;
	wire w_dff_B_2FL64ZH11_2;
	wire w_dff_B_YDsxh9a20_2;
	wire w_dff_B_If33qaQs2_2;
	wire w_dff_B_SPDZuxGI7_2;
	wire w_dff_B_Wbgx3rRy1_2;
	wire w_dff_B_6wTHl1Ox4_1;
	wire w_dff_B_rR2VyiWp9_1;
	wire w_dff_B_JGmtUXc49_1;
	wire w_dff_B_NLmdutY57_1;
	wire w_dff_B_vEVx6HVV3_1;
	wire w_dff_B_gPz9X9k84_1;
	wire w_dff_B_C87uUjoD4_1;
	wire w_dff_B_cOB7HS469_1;
	wire w_dff_B_HHhJVLGv9_1;
	wire w_dff_B_MUwpo5Z39_1;
	wire w_dff_B_oJRZRVc22_1;
	wire w_dff_B_Ye824Mux6_1;
	wire w_dff_B_eYelOqLP8_1;
	wire w_dff_B_ba0Ln3Us5_1;
	wire w_dff_B_YjHmnK9K0_1;
	wire w_dff_B_sIB6d5EG7_1;
	wire w_dff_B_vwMLsJ4L1_1;
	wire w_dff_B_83viOYOt7_1;
	wire w_dff_B_Mkb0lWqA0_1;
	wire w_dff_B_9Pr8HhzR3_1;
	wire w_dff_B_uCHmCYaJ6_1;
	wire w_dff_B_i6f3iihH5_1;
	wire w_dff_B_BFMrnTK47_1;
	wire w_dff_B_r3aWFr4W3_1;
	wire w_dff_B_PrGcamn13_1;
	wire w_dff_B_MUbeO81a9_1;
	wire w_dff_B_kkv2ItSd5_1;
	wire w_dff_B_qspT91km1_1;
	wire w_dff_A_PWdLB2rj7_0;
	wire w_dff_A_a91x22Jj1_0;
	wire w_dff_A_AkvgC7Sw9_0;
	wire w_dff_A_4gXPYZx31_0;
	wire w_dff_A_odEaCUEE8_0;
	wire w_dff_B_d4lvTgFq6_2;
	wire w_dff_B_nEgizuqm5_2;
	wire w_dff_B_eLgSdFBi3_2;
	wire w_dff_B_RNKea2g00_2;
	wire w_dff_B_SLgAIdx72_2;
	wire w_dff_B_bFYxaDpP3_2;
	wire w_dff_B_PLBUo2M06_2;
	wire w_dff_B_FcCrHuge5_2;
	wire w_dff_B_yQ9uAffr2_2;
	wire w_dff_B_gEIczuo23_2;
	wire w_dff_B_EVwBVohv4_2;
	wire w_dff_B_pbP9fPTx8_2;
	wire w_dff_B_13lMLyaC0_2;
	wire w_dff_B_SS5Ks74t8_2;
	wire w_dff_B_qVZ41wor8_2;
	wire w_dff_A_B2Z8rNqE5_0;
	wire w_dff_A_4p99zO6p2_0;
	wire w_dff_A_qCrNttSH4_0;
	wire w_dff_A_GUdBd9mu6_0;
	wire w_dff_A_nuSDMEPB6_0;
	wire w_dff_B_rCZn44ug3_2;
	wire w_dff_B_UBOJ8tzV7_2;
	wire w_dff_B_Ivo7Af3v1_2;
	wire w_dff_B_GHIdF3Hc5_2;
	wire w_dff_B_bn2DgXrP1_2;
	wire w_dff_B_mFyrlaSO8_2;
	wire w_dff_B_5RLFVkOf8_2;
	wire w_dff_B_qrsygGXs1_2;
	wire w_dff_B_eTK4Z6O22_2;
	wire w_dff_B_07mkwv4R7_2;
	wire w_dff_B_Ob73atk08_2;
	wire w_dff_B_tEEgs9xm5_2;
	wire w_dff_B_prjuiRUh1_2;
	wire w_dff_B_NBVsFsuc1_2;
	wire w_dff_A_oR4OMqBV7_0;
	wire w_dff_A_3IivIiSm3_0;
	wire w_dff_A_gOR6YDZr9_0;
	wire w_dff_A_ChFNvTk20_0;
	wire w_dff_A_pGeBBPKK0_0;
	wire w_dff_A_maON4xc73_0;
	wire w_dff_A_HY831AbW1_0;
	wire w_dff_A_YT86EpGx6_0;
	wire w_dff_A_qhDd3nSX7_0;
	wire w_dff_B_BSaj4DT15_1;
	wire w_dff_B_I2UqC6LA6_0;
	wire w_dff_A_XrUML48z4_0;
	wire w_dff_A_M5UfqVuK0_0;
	wire w_dff_A_N8AXmMWc8_0;
	wire w_dff_A_MOH7kBoI3_0;
	wire w_dff_A_Z6GXP7BJ3_0;
	wire w_dff_A_ynRIomY82_0;
	wire w_dff_A_ayfftHHh7_0;
	wire w_dff_A_P3ID5Ro71_0;
	wire w_dff_A_2pu4Shy09_0;
	wire w_dff_A_nD7T96vq3_0;
	wire w_dff_A_hve5nfuh0_0;
	wire w_dff_A_r3X03Ksn2_0;
	wire w_dff_B_rXmzRcqG0_1;
	wire w_dff_B_8WQo3Ph79_1;
	wire w_dff_B_2Eq2SDi60_1;
	wire w_dff_B_A74Dl4Lh8_1;
	wire w_dff_B_BjofQXO58_1;
	wire w_dff_A_odnU3JUb8_1;
	wire w_dff_B_LLRggoRx9_0;
	wire w_dff_B_y4l3xiDs4_0;
	wire w_dff_B_42Pvyqep0_0;
	wire w_dff_B_qUCQ2tVg4_0;
	wire w_dff_B_ZGg3Kssf1_0;
	wire w_dff_B_semhg0XA5_0;
	wire w_dff_A_Izc7gCgG6_0;
	wire w_dff_A_szyTS6Oa8_0;
	wire w_dff_A_51DMl5vl0_0;
	wire w_dff_A_CT5UaxRu8_0;
	wire w_dff_A_364EBhxd6_0;
	wire w_dff_A_63oZoyoF8_0;
	wire w_dff_B_XlN4GTGu6_2;
	wire w_dff_B_GI47OmJT5_2;
	wire w_dff_B_TS1nPMOJ9_2;
	wire w_dff_B_xiAKdumT6_2;
	wire w_dff_B_h4k8gdO21_2;
	wire w_dff_B_xKEzMDkM2_2;
	wire w_dff_B_3JvXLvY50_2;
	wire w_dff_B_JzZmHrNh0_2;
	wire w_dff_B_kx7Iet5W7_2;
	wire w_dff_B_BgT0exiJ8_2;
	wire w_dff_B_59OVdDxG3_2;
	wire w_dff_B_AtgwB8iE9_2;
	wire w_dff_B_lddyxjpx2_2;
	wire w_dff_B_YtIYVhHE4_2;
	wire w_dff_A_sKoCC3zh9_0;
	wire w_dff_A_NrIqP14M4_0;
	wire w_dff_A_2KzzHUxH0_0;
	wire w_dff_A_BpFrD0KW4_0;
	wire w_dff_A_1bTNjptD8_0;
	wire w_dff_A_gYVfYYle3_0;
	wire w_dff_B_0zfirOu97_1;
	wire w_dff_B_o9ZLIsAW3_1;
	wire w_dff_A_4uHBuKwJ9_0;
	wire w_dff_A_Zydon2Kb9_0;
	wire w_dff_A_RP8PBlkw9_0;
	wire w_dff_A_q3qz3Tvs6_0;
	wire w_dff_A_jJaiJ6vH3_0;
	wire w_dff_A_DnX4lryc8_0;
	wire w_dff_A_EIG2JM9W2_0;
	wire w_dff_A_4E7vCqTU1_0;
	wire w_dff_A_vAOwm7wp0_0;
	wire w_dff_A_l5z1HdZr0_0;
	wire w_dff_A_f6I0oko83_0;
	wire w_dff_A_to77wHFK6_0;
	wire w_dff_B_Lz8LZPOU1_1;
	wire w_dff_B_E5NdmgxO1_0;
	wire w_dff_A_bSXelBOE6_0;
	wire w_dff_A_wGzVZ1eT5_0;
	wire w_dff_A_YD51Llv40_0;
	wire w_dff_A_S54NF0lG5_0;
	wire w_dff_A_wM5s8YQ61_0;
	wire w_dff_A_jBN2c32x7_0;
	wire w_dff_B_KZlWoY7g0_1;
	wire w_dff_B_umaKUS525_1;
	wire w_dff_B_dTnArEg17_1;
	wire w_dff_B_9duBFX6L7_1;
	wire w_dff_B_85G61gFE4_1;
	wire w_dff_B_bgBLIMi30_1;
	wire w_dff_A_gBtP3tnQ1_0;
	wire w_dff_A_yu0xCXRO9_0;
	wire w_dff_A_ia1CDLVJ7_0;
	wire w_dff_A_xdUMVmIc8_0;
	wire w_dff_A_CxuA7Qma4_0;
	wire w_dff_A_3fldbpnW8_0;
	wire w_dff_A_4k5SSRp42_0;
	wire w_dff_A_VfBKlTKA0_0;
	wire w_dff_A_MJUiek4X8_0;
	wire w_dff_A_DIKNDfFh7_0;
	wire w_dff_A_Uic0RTvi3_0;
	wire w_dff_A_HKPFXnOD2_0;
	wire w_dff_A_WWUwobV88_1;
	wire w_dff_A_SapwMk784_1;
	wire w_dff_A_3zICCvER9_1;
	wire w_dff_A_KKlfiE8u7_1;
	wire w_dff_A_jGi9B9Xj8_1;
	wire w_dff_A_yYIsqFhH3_1;
	wire w_dff_A_XZ4IyHh82_0;
	wire w_dff_A_tr7D1iqO5_0;
	wire w_dff_A_zErVdf3p5_0;
	wire w_dff_A_xR8dBdnR1_0;
	wire w_dff_A_bc4wkJP60_0;
	wire w_dff_A_9BNznCqm5_0;
	wire w_dff_A_toHHMGld8_1;
	wire w_dff_A_hMAXkXG39_0;
	wire w_dff_A_JjcMM0Nf4_0;
	wire w_dff_A_eYdukx852_0;
	wire w_dff_A_ndOpu0aO1_0;
	wire w_dff_A_uABBfnFD9_0;
	wire w_dff_A_qKXRGcob8_0;
	wire w_dff_A_zdN3M1Yr4_0;
	wire w_dff_A_zGn1J7RA6_0;
	wire w_dff_A_UfIpb2WJ6_0;
	wire w_dff_A_iGMr5L8y5_0;
	wire w_dff_A_Q8mnEBbA1_0;
	wire w_dff_A_Ud3K8bkm7_0;
	wire w_dff_A_62ZBuxpt8_0;
	wire w_dff_A_YcS3E57m0_0;
	wire w_dff_A_oSvDBZ9y5_0;
	wire w_dff_A_jnphPJQq4_0;
	wire w_dff_A_e9UdxjJX2_0;
	wire w_dff_A_pVghKH8V0_0;
	wire w_dff_A_kyqh7XdT3_0;
	wire w_dff_A_I9c9A40x6_0;
	wire w_dff_A_HtwnrXEd7_1;
	wire w_dff_A_bnOtvpbk1_0;
	wire w_dff_A_nKAG9DvF0_0;
	wire w_dff_A_p6GH5ayH4_0;
	wire w_dff_A_yTinfqHI7_0;
	wire w_dff_A_PxgQhShx3_0;
	wire w_dff_A_Ju0kYDkb4_0;
	wire w_dff_A_KjOYL2s89_0;
	wire w_dff_A_FG5twln81_0;
	wire w_dff_A_Q9QrCNcM2_0;
	wire w_dff_A_Y8y80gZX3_0;
	wire w_dff_A_zUNyRLWq9_0;
	wire w_dff_A_M4nRc6jE1_0;
	wire w_dff_A_wVczK4xJ1_0;
	wire w_dff_A_CQ7xasqQ2_2;
	wire w_dff_A_QMiACvvH1_0;
	wire w_dff_A_MdlvTLdw8_0;
	wire w_dff_A_RM0lo1XM4_0;
	wire w_dff_A_0hA5HcLW0_0;
	wire w_dff_A_WRDgAVWl6_0;
	wire w_dff_A_nTSprNPu2_0;
	wire w_dff_A_Gk1ONaMb3_1;
	wire w_dff_A_ScGCnjWl0_0;
	jnot g000(.din(w_G102gat_0[1]),.dout(n43),.clk(gclk));
	jand g001(.dina(w_G108gat_0[2]),.dinb(w_n43_0[1]),.dout(n44),.clk(gclk));
	jnot g002(.din(w_G43gat_0[1]),.dout(n45),.clk(gclk));
	jor g003(.dina(w_n45_0[1]),.dinb(G37gat),.dout(n46),.clk(gclk));
	jnot g004(.din(w_n46_0[2]),.dout(n47),.clk(gclk));
	jor g005(.dina(w_n47_0[1]),.dinb(w_n44_0[1]),.dout(n48),.clk(gclk));
	jnot g006(.din(w_G63gat_0[2]),.dout(n49),.clk(gclk));
	jand g007(.dina(w_G69gat_0[2]),.dinb(w_n49_0[1]),.dout(n50),.clk(gclk));
	jnot g008(.din(w_G11gat_0[2]),.dout(n51),.clk(gclk));
	jand g009(.dina(w_G17gat_0[2]),.dinb(w_n51_0[1]),.dout(n52),.clk(gclk));
	jor g010(.dina(n52),.dinb(n50),.dout(n53),.clk(gclk));
	jnot g011(.din(w_G24gat_0[2]),.dout(n54),.clk(gclk));
	jand g012(.dina(w_G30gat_0[2]),.dinb(w_n54_0[1]),.dout(n55),.clk(gclk));
	jnot g013(.din(w_G50gat_0[1]),.dout(n56),.clk(gclk));
	jand g014(.dina(w_G56gat_1[1]),.dinb(n56),.dout(n57),.clk(gclk));
	jor g015(.dina(w_n57_0[1]),.dinb(n55),.dout(n58),.clk(gclk));
	jor g016(.dina(n58),.dinb(n53),.dout(n59),.clk(gclk));
	jnot g017(.din(w_G1gat_0[2]),.dout(n60),.clk(gclk));
	jand g018(.dina(w_G4gat_0[2]),.dinb(w_n60_0[1]),.dout(n61),.clk(gclk));
	jnot g019(.din(w_G89gat_0[2]),.dout(n62),.clk(gclk));
	jand g020(.dina(w_G95gat_0[2]),.dinb(w_n62_0[1]),.dout(n63),.clk(gclk));
	jnot g021(.din(w_G76gat_0[2]),.dout(n64),.clk(gclk));
	jand g022(.dina(w_G82gat_0[2]),.dinb(w_n64_0[1]),.dout(n65),.clk(gclk));
	jor g023(.dina(n65),.dinb(n63),.dout(n66),.clk(gclk));
	jor g024(.dina(n66),.dinb(n61),.dout(n67),.clk(gclk));
	jor g025(.dina(n67),.dinb(n59),.dout(n68),.clk(gclk));
	jor g026(.dina(n68),.dinb(n48),.dout(G223gat_fa_),.clk(gclk));
	jnot g027(.din(w_G21gat_0[2]),.dout(n70),.clk(gclk));
	jnot g028(.din(w_n44_0[0]),.dout(n71),.clk(gclk));
	jand g029(.dina(w_n46_0[1]),.dinb(n71),.dout(n72),.clk(gclk));
	jnot g030(.din(w_G69gat_0[1]),.dout(n73),.clk(gclk));
	jor g031(.dina(w_n73_0[1]),.dinb(w_G63gat_0[1]),.dout(n74),.clk(gclk));
	jnot g032(.din(w_G17gat_0[1]),.dout(n75),.clk(gclk));
	jor g033(.dina(w_n75_0[1]),.dinb(w_G11gat_0[1]),.dout(n76),.clk(gclk));
	jand g034(.dina(n76),.dinb(n74),.dout(n77),.clk(gclk));
	jnot g035(.din(w_G30gat_0[1]),.dout(n78),.clk(gclk));
	jor g036(.dina(w_n78_0[1]),.dinb(w_G24gat_0[1]),.dout(n79),.clk(gclk));
	jnot g037(.din(w_G56gat_1[0]),.dout(n80),.clk(gclk));
	jor g038(.dina(w_n80_0[1]),.dinb(w_G50gat_0[0]),.dout(n81),.clk(gclk));
	jand g039(.dina(w_n81_0[1]),.dinb(n79),.dout(n82),.clk(gclk));
	jand g040(.dina(n82),.dinb(n77),.dout(n83),.clk(gclk));
	jnot g041(.din(w_G4gat_0[1]),.dout(n84),.clk(gclk));
	jor g042(.dina(w_n84_0[1]),.dinb(w_G1gat_0[1]),.dout(n85),.clk(gclk));
	jnot g043(.din(w_G95gat_0[1]),.dout(n86),.clk(gclk));
	jor g044(.dina(w_n86_0[1]),.dinb(w_G89gat_0[1]),.dout(n87),.clk(gclk));
	jnot g045(.din(w_G82gat_0[1]),.dout(n88),.clk(gclk));
	jor g046(.dina(w_n88_0[1]),.dinb(w_G76gat_0[1]),.dout(n89),.clk(gclk));
	jand g047(.dina(n89),.dinb(n87),.dout(n90),.clk(gclk));
	jand g048(.dina(n90),.dinb(n85),.dout(n91),.clk(gclk));
	jand g049(.dina(n91),.dinb(n83),.dout(n92),.clk(gclk));
	jand g050(.dina(n92),.dinb(n72),.dout(n93),.clk(gclk));
	jor g051(.dina(w_n93_3[2]),.dinb(w_n51_0[0]),.dout(n94),.clk(gclk));
	jand g052(.dina(n94),.dinb(w_G17gat_0[0]),.dout(n95),.clk(gclk));
	jand g053(.dina(w_n95_0[1]),.dinb(w_n70_0[1]),.dout(n96),.clk(gclk));
	jnot g054(.din(w_G99gat_0[2]),.dout(n97),.clk(gclk));
	jor g055(.dina(w_n93_3[1]),.dinb(w_n62_0[0]),.dout(n98),.clk(gclk));
	jand g056(.dina(n98),.dinb(w_G95gat_0[0]),.dout(n99),.clk(gclk));
	jand g057(.dina(n99),.dinb(n97),.dout(n100),.clk(gclk));
	jor g058(.dina(n100),.dinb(n96),.dout(n101),.clk(gclk));
	jnot g059(.din(w_G73gat_0[2]),.dout(n102),.clk(gclk));
	jor g060(.dina(w_n93_3[0]),.dinb(w_n49_0[0]),.dout(n103),.clk(gclk));
	jand g061(.dina(n103),.dinb(w_G69gat_0[0]),.dout(n104),.clk(gclk));
	jand g062(.dina(w_n104_0[1]),.dinb(w_n102_0[1]),.dout(n105),.clk(gclk));
	jnot g063(.din(w_G34gat_0[2]),.dout(n106),.clk(gclk));
	jor g064(.dina(w_n93_2[2]),.dinb(w_n54_0[0]),.dout(n107),.clk(gclk));
	jand g065(.dina(n107),.dinb(w_G30gat_0[0]),.dout(n108),.clk(gclk));
	jand g066(.dina(w_n108_0[1]),.dinb(w_n106_0[1]),.dout(n109),.clk(gclk));
	jor g067(.dina(n109),.dinb(n105),.dout(n110),.clk(gclk));
	jnot g068(.din(w_G112gat_0[2]),.dout(n111),.clk(gclk));
	jor g069(.dina(w_n93_2[1]),.dinb(w_n43_0[0]),.dout(n112),.clk(gclk));
	jand g070(.dina(n112),.dinb(w_G108gat_0[1]),.dout(n113),.clk(gclk));
	jand g071(.dina(w_n113_0[1]),.dinb(w_n111_0[1]),.dout(n114),.clk(gclk));
	jor g072(.dina(n114),.dinb(n110),.dout(n115),.clk(gclk));
	jor g073(.dina(n115),.dinb(n101),.dout(n116),.clk(gclk));
	jnot g074(.din(w_G60gat_0[1]),.dout(n117),.clk(gclk));
	jxor g075(.dina(w_n93_2[0]),.dinb(w_n57_0[0]),.dout(n118),.clk(gclk));
	jand g076(.dina(n118),.dinb(w_G56gat_0[2]),.dout(n119),.clk(gclk));
	jand g077(.dina(w_n119_0[2]),.dinb(w_n117_0[1]),.dout(n120),.clk(gclk));
	jnot g078(.din(w_G86gat_0[2]),.dout(n121),.clk(gclk));
	jor g079(.dina(w_n93_1[2]),.dinb(w_n64_0[0]),.dout(n122),.clk(gclk));
	jand g080(.dina(n122),.dinb(w_G82gat_0[0]),.dout(n123),.clk(gclk));
	jand g081(.dina(w_n123_0[1]),.dinb(w_n121_0[1]),.dout(n124),.clk(gclk));
	jnot g082(.din(w_G8gat_0[2]),.dout(n125),.clk(gclk));
	jor g083(.dina(w_n93_1[1]),.dinb(w_n60_0[0]),.dout(n126),.clk(gclk));
	jand g084(.dina(n126),.dinb(w_G4gat_0[0]),.dout(n127),.clk(gclk));
	jand g085(.dina(w_n127_0[1]),.dinb(w_n125_0[1]),.dout(n128),.clk(gclk));
	jnot g086(.din(w_G47gat_0[2]),.dout(n129),.clk(gclk));
	jor g087(.dina(w_n93_1[0]),.dinb(w_n47_0[0]),.dout(n130),.clk(gclk));
	jand g088(.dina(n130),.dinb(w_G43gat_0[0]),.dout(n131),.clk(gclk));
	jand g089(.dina(w_n131_0[2]),.dinb(n129),.dout(n132),.clk(gclk));
	jor g090(.dina(n132),.dinb(n128),.dout(n133),.clk(gclk));
	jor g091(.dina(n133),.dinb(n124),.dout(n134),.clk(gclk));
	jor g092(.dina(n134),.dinb(w_n120_0[1]),.dout(n135),.clk(gclk));
	jor g093(.dina(n135),.dinb(n116),.dout(G329gat_fa_),.clk(gclk));
	jand g094(.dina(w_G223gat_4),.dinb(w_G89gat_0[0]),.dout(n137),.clk(gclk));
	jor g095(.dina(n137),.dinb(w_n86_0[0]),.dout(n138),.clk(gclk));
	jand g096(.dina(w_G329gat_4),.dinb(w_G99gat_0[1]),.dout(n139),.clk(gclk));
	jor g097(.dina(n139),.dinb(w_n138_0[1]),.dout(n140),.clk(gclk));
	jor g098(.dina(w_n140_0[1]),.dinb(w_G105gat_0[1]),.dout(n141),.clk(gclk));
	jnot g099(.din(w_n141_0[1]),.dout(n142),.clk(gclk));
	jand g100(.dina(w_G329gat_3[2]),.dinb(w_G47gat_0[1]),.dout(n143),.clk(gclk));
	jnot g101(.din(n143),.dout(n144),.clk(gclk));
	jnot g102(.din(w_G53gat_0[1]),.dout(n145),.clk(gclk));
	jand g103(.dina(w_n131_0[1]),.dinb(w_n145_0[1]),.dout(n146),.clk(gclk));
	jand g104(.dina(w_dff_B_semhg0XA5_0),.dinb(w_n144_0[1]),.dout(n147),.clk(gclk));
	jor g105(.dina(w_n147_0[1]),.dinb(n142),.dout(n148),.clk(gclk));
	jnot g106(.din(w_G40gat_0[1]),.dout(n149),.clk(gclk));
	jand g107(.dina(w_G223gat_3[2]),.dinb(w_G11gat_0[0]),.dout(n150),.clk(gclk));
	jor g108(.dina(n150),.dinb(w_n75_0[0]),.dout(n151),.clk(gclk));
	jor g109(.dina(w_n151_0[1]),.dinb(w_G21gat_0[1]),.dout(n152),.clk(gclk));
	jor g110(.dina(w_n138_0[0]),.dinb(w_G99gat_0[0]),.dout(n153),.clk(gclk));
	jand g111(.dina(n153),.dinb(n152),.dout(n154),.clk(gclk));
	jand g112(.dina(w_G223gat_3[1]),.dinb(w_G63gat_0[0]),.dout(n155),.clk(gclk));
	jor g113(.dina(n155),.dinb(w_n73_0[0]),.dout(n156),.clk(gclk));
	jor g114(.dina(w_n156_0[1]),.dinb(w_G73gat_0[1]),.dout(n157),.clk(gclk));
	jand g115(.dina(w_G223gat_3[0]),.dinb(w_G24gat_0[0]),.dout(n158),.clk(gclk));
	jor g116(.dina(n158),.dinb(w_n78_0[0]),.dout(n159),.clk(gclk));
	jor g117(.dina(w_n159_0[1]),.dinb(w_G34gat_0[1]),.dout(n160),.clk(gclk));
	jand g118(.dina(n160),.dinb(n157),.dout(n161),.clk(gclk));
	jnot g119(.din(w_G108gat_0[0]),.dout(n162),.clk(gclk));
	jand g120(.dina(w_G223gat_2[2]),.dinb(w_G102gat_0[0]),.dout(n163),.clk(gclk));
	jor g121(.dina(n163),.dinb(w_dff_B_bgBLIMi30_1),.dout(n164),.clk(gclk));
	jor g122(.dina(w_n164_0[1]),.dinb(w_G112gat_0[1]),.dout(n165),.clk(gclk));
	jand g123(.dina(w_dff_B_E5NdmgxO1_0),.dinb(n161),.dout(n166),.clk(gclk));
	jand g124(.dina(n166),.dinb(w_dff_B_Lz8LZPOU1_1),.dout(n167),.clk(gclk));
	jnot g125(.din(w_n120_0[0]),.dout(n168),.clk(gclk));
	jand g126(.dina(w_G223gat_2[1]),.dinb(w_G76gat_0[0]),.dout(n169),.clk(gclk));
	jor g127(.dina(n169),.dinb(w_n88_0[0]),.dout(n170),.clk(gclk));
	jor g128(.dina(w_n170_0[1]),.dinb(w_G86gat_0[1]),.dout(n171),.clk(gclk));
	jand g129(.dina(w_G223gat_2[0]),.dinb(w_G1gat_0[0]),.dout(n172),.clk(gclk));
	jor g130(.dina(n172),.dinb(w_n84_0[0]),.dout(n173),.clk(gclk));
	jor g131(.dina(w_n173_0[1]),.dinb(w_G8gat_0[1]),.dout(n174),.clk(gclk));
	jand g132(.dina(w_G223gat_1[2]),.dinb(w_n46_0[0]),.dout(n175),.clk(gclk));
	jor g133(.dina(n175),.dinb(w_n45_0[0]),.dout(n176),.clk(gclk));
	jor g134(.dina(n176),.dinb(w_G47gat_0[0]),.dout(n177),.clk(gclk));
	jand g135(.dina(n177),.dinb(n174),.dout(n178),.clk(gclk));
	jand g136(.dina(n178),.dinb(w_dff_B_o9ZLIsAW3_1),.dout(n179),.clk(gclk));
	jand g137(.dina(n179),.dinb(w_dff_B_0zfirOu97_1),.dout(n180),.clk(gclk));
	jand g138(.dina(n180),.dinb(n167),.dout(n181),.clk(gclk));
	jor g139(.dina(w_n181_2[2]),.dinb(w_n106_0[0]),.dout(n182),.clk(gclk));
	jand g140(.dina(n182),.dinb(w_n108_0[0]),.dout(n183),.clk(gclk));
	jand g141(.dina(w_n183_0[1]),.dinb(w_n149_0[1]),.dout(n184),.clk(gclk));
	jnot g142(.din(w_G66gat_0[2]),.dout(n185),.clk(gclk));
	jor g143(.dina(w_n181_2[1]),.dinb(w_n117_0[0]),.dout(n186),.clk(gclk));
	jand g144(.dina(n186),.dinb(w_n119_0[1]),.dout(n187),.clk(gclk));
	jand g145(.dina(n187),.dinb(w_n185_0[1]),.dout(n188),.clk(gclk));
	jor g146(.dina(n188),.dinb(n184),.dout(n189),.clk(gclk));
	jnot g147(.din(w_G14gat_0[2]),.dout(n190),.clk(gclk));
	jor g148(.dina(w_n181_2[0]),.dinb(w_n125_0[0]),.dout(n191),.clk(gclk));
	jand g149(.dina(n191),.dinb(w_n127_0[0]),.dout(n192),.clk(gclk));
	jand g150(.dina(n192),.dinb(w_dff_B_qspT91km1_1),.dout(n193),.clk(gclk));
	jnot g151(.din(w_G92gat_0[2]),.dout(n194),.clk(gclk));
	jor g152(.dina(w_n181_1[2]),.dinb(w_n121_0[0]),.dout(n195),.clk(gclk));
	jand g153(.dina(n195),.dinb(w_n123_0[0]),.dout(n196),.clk(gclk));
	jand g154(.dina(n196),.dinb(w_dff_B_ba0Ln3Us5_1),.dout(n197),.clk(gclk));
	jor g155(.dina(n197),.dinb(n193),.dout(n198),.clk(gclk));
	jor g156(.dina(n198),.dinb(n189),.dout(n199),.clk(gclk));
	jnot g157(.din(w_G79gat_0[1]),.dout(n200),.clk(gclk));
	jor g158(.dina(w_n181_1[1]),.dinb(w_n102_0[0]),.dout(n201),.clk(gclk));
	jand g159(.dina(n201),.dinb(w_n104_0[0]),.dout(n202),.clk(gclk));
	jand g160(.dina(w_n202_0[1]),.dinb(w_n200_0[1]),.dout(n203),.clk(gclk));
	jnot g161(.din(w_G115gat_0[1]),.dout(n204),.clk(gclk));
	jor g162(.dina(w_n181_1[0]),.dinb(w_n111_0[0]),.dout(n205),.clk(gclk));
	jand g163(.dina(n205),.dinb(w_n113_0[0]),.dout(n206),.clk(gclk));
	jand g164(.dina(w_n206_0[1]),.dinb(w_n204_0[1]),.dout(n207),.clk(gclk));
	jor g165(.dina(n207),.dinb(n203),.dout(n208),.clk(gclk));
	jnot g166(.din(w_G27gat_0[1]),.dout(n209),.clk(gclk));
	jor g167(.dina(w_n181_0[2]),.dinb(w_n70_0[0]),.dout(n210),.clk(gclk));
	jand g168(.dina(n210),.dinb(w_n95_0[0]),.dout(n211),.clk(gclk));
	jand g169(.dina(w_n211_0[1]),.dinb(w_n209_0[1]),.dout(n212),.clk(gclk));
	jor g170(.dina(w_dff_B_QP2GGXYy0_0),.dinb(n208),.dout(n213),.clk(gclk));
	jor g171(.dina(n213),.dinb(n199),.dout(n214),.clk(gclk));
	jor g172(.dina(n214),.dinb(w_dff_B_lwXOQWpt6_1),.dout(G370gat_fa_),.clk(gclk));
	jnot g173(.din(w_n147_0[0]),.dout(n216),.clk(gclk));
	jand g174(.dina(n216),.dinb(w_n141_0[0]),.dout(n217),.clk(gclk));
	jand g175(.dina(w_G329gat_3[1]),.dinb(w_G34gat_0[0]),.dout(n218),.clk(gclk));
	jor g176(.dina(n218),.dinb(w_n159_0[0]),.dout(n219),.clk(gclk));
	jor g177(.dina(n219),.dinb(w_G40gat_0[0]),.dout(n220),.clk(gclk));
	jnot g178(.din(w_n119_0[0]),.dout(n221),.clk(gclk));
	jand g179(.dina(w_G329gat_3[0]),.dinb(w_G60gat_0[0]),.dout(n222),.clk(gclk));
	jor g180(.dina(w_n222_0[1]),.dinb(w_dff_B_BjofQXO58_1),.dout(n223),.clk(gclk));
	jor g181(.dina(n223),.dinb(w_G66gat_0[1]),.dout(n224),.clk(gclk));
	jand g182(.dina(n224),.dinb(n220),.dout(n225),.clk(gclk));
	jand g183(.dina(w_G329gat_2[2]),.dinb(w_G8gat_0[0]),.dout(n226),.clk(gclk));
	jor g184(.dina(n226),.dinb(w_n173_0[0]),.dout(n227),.clk(gclk));
	jor g185(.dina(w_n227_0[1]),.dinb(w_G14gat_0[1]),.dout(n228),.clk(gclk));
	jand g186(.dina(w_G329gat_2[1]),.dinb(w_G86gat_0[0]),.dout(n229),.clk(gclk));
	jor g187(.dina(n229),.dinb(w_n170_0[0]),.dout(n230),.clk(gclk));
	jor g188(.dina(w_n230_0[1]),.dinb(w_G92gat_0[1]),.dout(n231),.clk(gclk));
	jand g189(.dina(n231),.dinb(n228),.dout(n232),.clk(gclk));
	jand g190(.dina(n232),.dinb(n225),.dout(n233),.clk(gclk));
	jand g191(.dina(w_G329gat_2[0]),.dinb(w_G73gat_0[0]),.dout(n234),.clk(gclk));
	jor g192(.dina(n234),.dinb(w_n156_0[0]),.dout(n235),.clk(gclk));
	jor g193(.dina(n235),.dinb(w_G79gat_0[0]),.dout(n236),.clk(gclk));
	jand g194(.dina(w_G329gat_1[2]),.dinb(w_G112gat_0[0]),.dout(n237),.clk(gclk));
	jor g195(.dina(n237),.dinb(w_n164_0[0]),.dout(n238),.clk(gclk));
	jor g196(.dina(n238),.dinb(w_G115gat_0[0]),.dout(n239),.clk(gclk));
	jand g197(.dina(n239),.dinb(n236),.dout(n240),.clk(gclk));
	jand g198(.dina(w_G329gat_1[1]),.dinb(w_G21gat_0[0]),.dout(n241),.clk(gclk));
	jor g199(.dina(n241),.dinb(w_n151_0[0]),.dout(n242),.clk(gclk));
	jor g200(.dina(n242),.dinb(w_G27gat_0[0]),.dout(n243),.clk(gclk));
	jand g201(.dina(w_dff_B_I2UqC6LA6_0),.dinb(n240),.dout(n244),.clk(gclk));
	jand g202(.dina(n244),.dinb(n233),.dout(n245),.clk(gclk));
	jand g203(.dina(n245),.dinb(w_dff_B_BSaj4DT15_1),.dout(n246),.clk(gclk));
	jor g204(.dina(w_n246_2[2]),.dinb(w_n209_0[0]),.dout(n247),.clk(gclk));
	jand g205(.dina(n247),.dinb(w_n211_0[0]),.dout(n248),.clk(gclk));
	jor g206(.dina(w_n246_2[1]),.dinb(w_n149_0[0]),.dout(n249),.clk(gclk));
	jand g207(.dina(n249),.dinb(w_n183_0[0]),.dout(n250),.clk(gclk));
	jor g208(.dina(w_n250_0[1]),.dinb(w_n248_0[1]),.dout(n251),.clk(gclk));
	jor g209(.dina(w_n246_2[0]),.dinb(w_n145_0[0]),.dout(n252),.clk(gclk));
	jand g210(.dina(w_n144_0[0]),.dinb(w_n131_0[0]),.dout(n253),.clk(gclk));
	jand g211(.dina(w_n253_0[1]),.dinb(n252),.dout(n254),.clk(gclk));
	jor g212(.dina(w_n246_1[2]),.dinb(w_n185_0[0]),.dout(n255),.clk(gclk));
	jand g213(.dina(w_G223gat_1[1]),.dinb(w_n81_0[0]),.dout(n256),.clk(gclk));
	jor g214(.dina(w_n222_0[0]),.dinb(w_dff_B_lXsBvo7M9_1),.dout(n257),.clk(gclk));
	jnot g215(.din(w_n257_0[1]),.dout(n258),.clk(gclk));
	jand g216(.dina(w_dff_B_haVkYUuq3_0),.dinb(n255),.dout(n259),.clk(gclk));
	jand g217(.dina(n259),.dinb(w_G56gat_0[1]),.dout(n260),.clk(gclk));
	jor g218(.dina(n260),.dinb(w_n254_0[1]),.dout(n261),.clk(gclk));
	jor g219(.dina(n261),.dinb(w_n251_0[1]),.dout(G430gat_fa_),.clk(gclk));
	jand g220(.dina(w_G370gat_1[1]),.dinb(w_G92gat_0[0]),.dout(n263),.clk(gclk));
	jor g221(.dina(n263),.dinb(w_n230_0[0]),.dout(n264),.clk(gclk));
	jnot g222(.din(w_n264_0[1]),.dout(n265),.clk(gclk));
	jnot g223(.din(w_n140_0[0]),.dout(n266),.clk(gclk));
	jnot g224(.din(w_G105gat_0[0]),.dout(n267),.clk(gclk));
	jor g225(.dina(w_n246_1[1]),.dinb(w_dff_B_OjPKiWFI0_1),.dout(n268),.clk(gclk));
	jand g226(.dina(n268),.dinb(w_dff_B_jGLnkveQ9_1),.dout(n269),.clk(gclk));
	jor g227(.dina(w_n246_1[0]),.dinb(w_n200_0[0]),.dout(n270),.clk(gclk));
	jand g228(.dina(n270),.dinb(w_n202_0[0]),.dout(n271),.clk(gclk));
	jor g229(.dina(w_n246_0[2]),.dinb(w_n204_0[0]),.dout(n272),.clk(gclk));
	jand g230(.dina(n272),.dinb(w_n206_0[0]),.dout(n273),.clk(gclk));
	jor g231(.dina(n273),.dinb(w_n271_0[1]),.dout(n274),.clk(gclk));
	jor g232(.dina(n274),.dinb(w_n269_0[1]),.dout(n275),.clk(gclk));
	jor g233(.dina(n275),.dinb(w_n265_0[1]),.dout(n276),.clk(gclk));
	jor g234(.dina(n276),.dinb(w_G430gat_0),.dout(n277),.clk(gclk));
	jand g235(.dina(w_G370gat_1[0]),.dinb(w_G14gat_0[0]),.dout(n278),.clk(gclk));
	jor g236(.dina(n278),.dinb(w_n227_0[0]),.dout(n279),.clk(gclk));
	jand g237(.dina(w_dff_B_3PqJqlKa2_0),.dinb(n277),.dout(G421gat),.clk(gclk));
	jnot g238(.din(w_n250_0[0]),.dout(n281),.clk(gclk));
	jand g239(.dina(w_G370gat_0[2]),.dinb(w_G53gat_0[0]),.dout(n282),.clk(gclk));
	jnot g240(.din(w_n253_0[0]),.dout(n283),.clk(gclk));
	jor g241(.dina(w_dff_B_MJ3zYHxJ4_0),.dinb(n282),.dout(n284),.clk(gclk));
	jand g242(.dina(w_G370gat_0[1]),.dinb(w_G66gat_0[0]),.dout(n285),.clk(gclk));
	jor g243(.dina(w_n257_0[0]),.dinb(n285),.dout(n286),.clk(gclk));
	jor g244(.dina(n286),.dinb(w_n80_0[0]),.dout(n287),.clk(gclk));
	jand g245(.dina(n287),.dinb(w_dff_B_aiwcWzfd6_1),.dout(n288),.clk(gclk));
	jand g246(.dina(w_n288_0[1]),.dinb(w_n281_0[1]),.dout(n289),.clk(gclk));
	jand g247(.dina(n289),.dinb(w_n271_0[0]),.dout(n290),.clk(gclk));
	jand g248(.dina(w_n265_0[0]),.dinb(w_n288_0[0]),.dout(n291),.clk(gclk));
	jor g249(.dina(n291),.dinb(w_n251_0[0]),.dout(n292),.clk(gclk));
	jor g250(.dina(n292),.dinb(w_n290_0[1]),.dout(G431gat),.clk(gclk));
	jand g251(.dina(w_n269_0[0]),.dinb(w_n264_0[0]),.dout(n294),.clk(gclk));
	jor g252(.dina(n294),.dinb(w_n254_0[0]),.dout(n295),.clk(gclk));
	jand g253(.dina(n295),.dinb(w_n281_0[0]),.dout(n296),.clk(gclk));
	jor g254(.dina(n296),.dinb(w_n248_0[0]),.dout(n297),.clk(gclk));
	jor g255(.dina(n297),.dinb(w_n290_0[0]),.dout(G432gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_G4gat_0[0]),.doutb(w_G4gat_0[1]),.doutc(w_G4gat_0[2]),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G11gat_0(.douta(w_G11gat_0[0]),.doutb(w_G11gat_0[1]),.doutc(w_G11gat_0[2]),.din(G11gat));
	jspl3 jspl3_w_G14gat_0(.douta(w_G14gat_0[0]),.doutb(w_G14gat_0[1]),.doutc(w_G14gat_0[2]),.din(G14gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_G21gat_0[0]),.doutb(w_G21gat_0[1]),.doutc(w_G21gat_0[2]),.din(G21gat));
	jspl3 jspl3_w_G24gat_0(.douta(w_G24gat_0[0]),.doutb(w_G24gat_0[1]),.doutc(w_G24gat_0[2]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_G27gat_0[0]),.doutb(w_G27gat_0[1]),.din(G27gat));
	jspl3 jspl3_w_G30gat_0(.douta(w_G30gat_0[0]),.doutb(w_G30gat_0[1]),.doutc(w_G30gat_0[2]),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_G34gat_0[0]),.doutb(w_G34gat_0[1]),.doutc(w_G34gat_0[2]),.din(G34gat));
	jspl jspl_w_G40gat_0(.douta(w_G40gat_0[0]),.doutb(w_G40gat_0[1]),.din(G40gat));
	jspl jspl_w_G43gat_0(.douta(w_G43gat_0[0]),.doutb(w_G43gat_0[1]),.din(G43gat));
	jspl3 jspl3_w_G47gat_0(.douta(w_G47gat_0[0]),.doutb(w_G47gat_0[1]),.doutc(w_G47gat_0[2]),.din(G47gat));
	jspl jspl_w_G50gat_0(.douta(w_G50gat_0[0]),.doutb(w_G50gat_0[1]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_G53gat_0[0]),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_G56gat_0[0]),.doutb(w_G56gat_0[1]),.doutc(w_G56gat_0[2]),.din(G56gat));
	jspl jspl_w_G56gat_1(.douta(w_G56gat_1[0]),.doutb(w_G56gat_1[1]),.din(w_G56gat_0[0]));
	jspl jspl_w_G60gat_0(.douta(w_G60gat_0[0]),.doutb(w_G60gat_0[1]),.din(G60gat));
	jspl3 jspl3_w_G63gat_0(.douta(w_G63gat_0[0]),.doutb(w_G63gat_0[1]),.doutc(w_G63gat_0[2]),.din(G63gat));
	jspl3 jspl3_w_G66gat_0(.douta(w_G66gat_0[0]),.doutb(w_G66gat_0[1]),.doutc(w_G66gat_0[2]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G73gat_0(.douta(w_G73gat_0[0]),.doutb(w_G73gat_0[1]),.doutc(w_G73gat_0[2]),.din(G73gat));
	jspl3 jspl3_w_G76gat_0(.douta(w_G76gat_0[0]),.doutb(w_G76gat_0[1]),.doutc(w_G76gat_0[2]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_G79gat_0[0]),.doutb(w_G79gat_0[1]),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_G82gat_0[0]),.doutb(w_G82gat_0[1]),.doutc(w_G82gat_0[2]),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G89gat_0(.douta(w_G89gat_0[0]),.doutb(w_G89gat_0[1]),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_G92gat_0[0]),.doutb(w_G92gat_0[1]),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_G95gat_0[0]),.doutb(w_G95gat_0[1]),.doutc(w_G95gat_0[2]),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_G99gat_0[0]),.doutb(w_G99gat_0[1]),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl jspl_w_G102gat_0(.douta(w_G102gat_0[0]),.doutb(w_G102gat_0[1]),.din(G102gat));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_G105gat_0[1]),.din(G105gat));
	jspl3 jspl3_w_G108gat_0(.douta(w_G108gat_0[0]),.doutb(w_G108gat_0[1]),.doutc(w_G108gat_0[2]),.din(G108gat));
	jspl3 jspl3_w_G112gat_0(.douta(w_G112gat_0[0]),.doutb(w_G112gat_0[1]),.doutc(w_G112gat_0[2]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_G115gat_0[0]),.doutb(w_G115gat_0[1]),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(w_G223gat_3[2]),.din(w_G223gat_0[2]));
	jspl jspl_w_G223gat_4(.douta(w_G223gat_4),.doutb(w_dff_A_toHHMGld8_1),.din(w_G223gat_1[0]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl jspl_w_G329gat_4(.douta(w_G329gat_4),.doutb(w_dff_A_HtwnrXEd7_1),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_dff_A_CQ7xasqQ2_2),.din(w_G370gat_0[0]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(w_dff_A_Gk1ONaMb3_1),.din(G430gat_fa_));
	jspl jspl_w_n43_0(.douta(w_n43_0[0]),.doutb(w_n43_0[1]),.din(n43));
	jspl jspl_w_n44_0(.douta(w_n44_0[0]),.doutb(w_n44_0[1]),.din(n44));
	jspl jspl_w_n45_0(.douta(w_n45_0[0]),.doutb(w_n45_0[1]),.din(n45));
	jspl3 jspl3_w_n46_0(.douta(w_n46_0[0]),.doutb(w_n46_0[1]),.doutc(w_n46_0[2]),.din(n46));
	jspl jspl_w_n47_0(.douta(w_n47_0[0]),.doutb(w_n47_0[1]),.din(n47));
	jspl jspl_w_n49_0(.douta(w_n49_0[0]),.doutb(w_n49_0[1]),.din(n49));
	jspl jspl_w_n51_0(.douta(w_n51_0[0]),.doutb(w_n51_0[1]),.din(n51));
	jspl jspl_w_n54_0(.douta(w_n54_0[0]),.doutb(w_n54_0[1]),.din(n54));
	jspl jspl_w_n57_0(.douta(w_n57_0[0]),.doutb(w_n57_0[1]),.din(n57));
	jspl jspl_w_n60_0(.douta(w_n60_0[0]),.doutb(w_n60_0[1]),.din(n60));
	jspl jspl_w_n62_0(.douta(w_n62_0[0]),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n64_0(.douta(w_n64_0[0]),.doutb(w_n64_0[1]),.din(n64));
	jspl jspl_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.din(n80));
	jspl jspl_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.din(n81));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl3 jspl3_w_n93_1(.douta(w_n93_1[0]),.doutb(w_n93_1[1]),.doutc(w_n93_1[2]),.din(w_n93_0[0]));
	jspl3 jspl3_w_n93_2(.douta(w_n93_2[0]),.doutb(w_n93_2[1]),.doutc(w_n93_2[2]),.din(w_n93_0[1]));
	jspl3 jspl3_w_n93_3(.douta(w_n93_3[0]),.doutb(w_n93_3[1]),.doutc(w_n93_3[2]),.din(w_n93_0[2]));
	jspl jspl_w_n95_0(.douta(w_n95_0[0]),.doutb(w_n95_0[1]),.din(n95));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n106_0(.douta(w_n106_0[0]),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.din(n113));
	jspl jspl_w_n117_0(.douta(w_n117_0[0]),.doutb(w_n117_0[1]),.din(n117));
	jspl3 jspl3_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.doutc(w_n119_0[2]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl3 jspl3_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.doutc(w_n131_0[2]),.din(n131));
	jspl jspl_w_n138_0(.douta(w_n138_0[0]),.doutb(w_dff_A_yYIsqFhH3_1),.din(n138));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n141_0(.douta(w_dff_A_Izc7gCgG6_0),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(n144));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_dff_A_odnU3JUb8_1),.din(n147));
	jspl jspl_w_n149_0(.douta(w_dff_A_nuSDMEPB6_0),.doutb(w_n149_0[1]),.din(w_dff_B_NBVsFsuc1_2));
	jspl jspl_w_n151_0(.douta(w_dff_A_9BNznCqm5_0),.doutb(w_n151_0[1]),.din(n151));
	jspl jspl_w_n156_0(.douta(w_dff_A_HKPFXnOD2_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n159_0(.douta(w_dff_A_3fldbpnW8_0),.doutb(w_n159_0[1]),.din(n159));
	jspl jspl_w_n164_0(.douta(w_dff_A_jBN2c32x7_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n170_0(.douta(w_dff_A_to77wHFK6_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n173_0(.douta(w_dff_A_DnX4lryc8_0),.doutb(w_n173_0[1]),.din(n173));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n181_2(.douta(w_n181_2[0]),.doutb(w_n181_2[1]),.doutc(w_n181_2[2]),.din(w_n181_0[1]));
	jspl jspl_w_n183_0(.douta(w_dff_A_maON4xc73_0),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n185_0(.douta(w_dff_A_odEaCUEE8_0),.doutb(w_n185_0[1]),.din(w_dff_B_SS5Ks74t8_2));
	jspl jspl_w_n200_0(.douta(w_dff_A_63oZoyoF8_0),.doutb(w_n200_0[1]),.din(w_dff_B_YtIYVhHE4_2));
	jspl jspl_w_n202_0(.douta(w_dff_A_gYVfYYle3_0),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n204_0(.douta(w_dff_A_OYZRaIO26_0),.doutb(w_n204_0[1]),.din(w_dff_B_Wbgx3rRy1_2));
	jspl jspl_w_n206_0(.douta(w_dff_A_vZXliEu80_0),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n209_0(.douta(w_dff_A_UiOlqUe47_0),.doutb(w_n209_0[1]),.din(w_dff_B_6RajPZ225_2));
	jspl jspl_w_n211_0(.douta(w_dff_A_yja1jA0G3_0),.doutb(w_n211_0[1]),.din(n211));
	jspl jspl_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n227_0(.douta(w_dff_A_r3X03Ksn2_0),.doutb(w_n227_0[1]),.din(n227));
	jspl jspl_w_n230_0(.douta(w_dff_A_ynRIomY82_0),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl3 jspl3_w_n246_1(.douta(w_n246_1[0]),.doutb(w_n246_1[1]),.doutc(w_n246_1[2]),.din(w_n246_0[0]));
	jspl3 jspl3_w_n246_2(.douta(w_n246_2[0]),.doutb(w_n246_2[1]),.doutc(w_n246_2[2]),.din(w_n246_0[1]));
	jspl jspl_w_n248_0(.douta(w_dff_A_kXafuMAw3_0),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_dff_A_UHkQgKLo7_0),.doutb(w_n251_0[1]),.din(w_dff_B_FlrqaWjo7_2));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_dff_A_YeVc5UOD3_1),.din(n253));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(w_dff_B_sD7gCxad0_2));
	jspl jspl_w_n257_0(.douta(w_dff_A_vcKH6jI99_0),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(w_dff_B_3sV01tN74_2));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_dff_A_4ZGDBSoA9_1),.din(n269));
	jspl jspl_w_n271_0(.douta(w_dff_A_qhDd3nSX7_0),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.din(w_dff_B_qVZ41wor8_2));
	jspl jspl_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.din(n288));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(n290));
	jdff dff_B_TUGn5viz4_0(.din(n279),.dout(w_dff_B_TUGn5viz4_0),.clk(gclk));
	jdff dff_B_tG6glVm67_0(.din(w_dff_B_TUGn5viz4_0),.dout(w_dff_B_tG6glVm67_0),.clk(gclk));
	jdff dff_B_VHlRVsXk8_0(.din(w_dff_B_tG6glVm67_0),.dout(w_dff_B_VHlRVsXk8_0),.clk(gclk));
	jdff dff_B_3PqJqlKa2_0(.din(w_dff_B_VHlRVsXk8_0),.dout(w_dff_B_3PqJqlKa2_0),.clk(gclk));
	jdff dff_B_5mbO5f7u4_0(.din(n258),.dout(w_dff_B_5mbO5f7u4_0),.clk(gclk));
	jdff dff_B_RHpznR979_0(.din(w_dff_B_5mbO5f7u4_0),.dout(w_dff_B_RHpznR979_0),.clk(gclk));
	jdff dff_B_gfFb8n1K8_0(.din(w_dff_B_RHpznR979_0),.dout(w_dff_B_gfFb8n1K8_0),.clk(gclk));
	jdff dff_B_djEVmgys0_0(.din(w_dff_B_gfFb8n1K8_0),.dout(w_dff_B_djEVmgys0_0),.clk(gclk));
	jdff dff_B_haVkYUuq3_0(.din(w_dff_B_djEVmgys0_0),.dout(w_dff_B_haVkYUuq3_0),.clk(gclk));
	jdff dff_B_3sV01tN74_2(.din(n265),.dout(w_dff_B_3sV01tN74_2),.clk(gclk));
	jdff dff_A_UHkQgKLo7_0(.dout(w_n251_0[0]),.din(w_dff_A_UHkQgKLo7_0),.clk(gclk));
	jdff dff_B_FlrqaWjo7_2(.din(n251),.dout(w_dff_B_FlrqaWjo7_2),.clk(gclk));
	jdff dff_A_4ZGDBSoA9_1(.dout(w_n269_0[1]),.din(w_dff_A_4ZGDBSoA9_1),.clk(gclk));
	jdff dff_B_93W8t1sd2_1(.din(n266),.dout(w_dff_B_93W8t1sd2_1),.clk(gclk));
	jdff dff_B_JqKvAV603_1(.din(w_dff_B_93W8t1sd2_1),.dout(w_dff_B_JqKvAV603_1),.clk(gclk));
	jdff dff_B_AfVnNhxM8_1(.din(w_dff_B_JqKvAV603_1),.dout(w_dff_B_AfVnNhxM8_1),.clk(gclk));
	jdff dff_B_nwJrN7zD5_1(.din(w_dff_B_AfVnNhxM8_1),.dout(w_dff_B_nwJrN7zD5_1),.clk(gclk));
	jdff dff_B_jGLnkveQ9_1(.din(w_dff_B_nwJrN7zD5_1),.dout(w_dff_B_jGLnkveQ9_1),.clk(gclk));
	jdff dff_B_kXx7g4k74_1(.din(n267),.dout(w_dff_B_kXx7g4k74_1),.clk(gclk));
	jdff dff_B_nSLP0dXm0_1(.din(w_dff_B_kXx7g4k74_1),.dout(w_dff_B_nSLP0dXm0_1),.clk(gclk));
	jdff dff_B_XljKjWDk9_1(.din(w_dff_B_nSLP0dXm0_1),.dout(w_dff_B_XljKjWDk9_1),.clk(gclk));
	jdff dff_B_qv6pQL5z4_1(.din(w_dff_B_XljKjWDk9_1),.dout(w_dff_B_qv6pQL5z4_1),.clk(gclk));
	jdff dff_B_Dz4jzG8q1_1(.din(w_dff_B_qv6pQL5z4_1),.dout(w_dff_B_Dz4jzG8q1_1),.clk(gclk));
	jdff dff_B_5MUvVNGe7_1(.din(w_dff_B_Dz4jzG8q1_1),.dout(w_dff_B_5MUvVNGe7_1),.clk(gclk));
	jdff dff_B_5opjKqlz4_1(.din(w_dff_B_5MUvVNGe7_1),.dout(w_dff_B_5opjKqlz4_1),.clk(gclk));
	jdff dff_B_Chl8E2SN0_1(.din(w_dff_B_5opjKqlz4_1),.dout(w_dff_B_Chl8E2SN0_1),.clk(gclk));
	jdff dff_B_0b0j6Mz34_1(.din(w_dff_B_Chl8E2SN0_1),.dout(w_dff_B_0b0j6Mz34_1),.clk(gclk));
	jdff dff_B_3552XGda2_1(.din(w_dff_B_0b0j6Mz34_1),.dout(w_dff_B_3552XGda2_1),.clk(gclk));
	jdff dff_B_6dsNo7H12_1(.din(w_dff_B_3552XGda2_1),.dout(w_dff_B_6dsNo7H12_1),.clk(gclk));
	jdff dff_B_dSzDWF9f1_1(.din(w_dff_B_6dsNo7H12_1),.dout(w_dff_B_dSzDWF9f1_1),.clk(gclk));
	jdff dff_B_ZYhtOIYc2_1(.din(w_dff_B_dSzDWF9f1_1),.dout(w_dff_B_ZYhtOIYc2_1),.clk(gclk));
	jdff dff_B_BsagiSh45_1(.din(w_dff_B_ZYhtOIYc2_1),.dout(w_dff_B_BsagiSh45_1),.clk(gclk));
	jdff dff_B_3682yVZD5_1(.din(w_dff_B_BsagiSh45_1),.dout(w_dff_B_3682yVZD5_1),.clk(gclk));
	jdff dff_B_00FgM2Us0_1(.din(w_dff_B_3682yVZD5_1),.dout(w_dff_B_00FgM2Us0_1),.clk(gclk));
	jdff dff_B_X0KPIGTs9_1(.din(w_dff_B_00FgM2Us0_1),.dout(w_dff_B_X0KPIGTs9_1),.clk(gclk));
	jdff dff_B_0vHgPdV99_1(.din(w_dff_B_X0KPIGTs9_1),.dout(w_dff_B_0vHgPdV99_1),.clk(gclk));
	jdff dff_B_OjPKiWFI0_1(.din(w_dff_B_0vHgPdV99_1),.dout(w_dff_B_OjPKiWFI0_1),.clk(gclk));
	jdff dff_B_sD7gCxad0_2(.din(n254),.dout(w_dff_B_sD7gCxad0_2),.clk(gclk));
	jdff dff_A_vHQ7tY2m1_0(.dout(w_n248_0[0]),.din(w_dff_A_vHQ7tY2m1_0),.clk(gclk));
	jdff dff_A_OWCEaoKo1_0(.dout(w_dff_A_vHQ7tY2m1_0),.din(w_dff_A_OWCEaoKo1_0),.clk(gclk));
	jdff dff_A_kXafuMAw3_0(.dout(w_dff_A_OWCEaoKo1_0),.din(w_dff_A_kXafuMAw3_0),.clk(gclk));
	jdff dff_B_aiwcWzfd6_1(.din(n284),.dout(w_dff_B_aiwcWzfd6_1),.clk(gclk));
	jdff dff_A_rF4bOhRf9_0(.dout(w_n257_0[0]),.din(w_dff_A_rF4bOhRf9_0),.clk(gclk));
	jdff dff_A_OU0O9T7b6_0(.dout(w_dff_A_rF4bOhRf9_0),.din(w_dff_A_OU0O9T7b6_0),.clk(gclk));
	jdff dff_A_28gX06vb9_0(.dout(w_dff_A_OU0O9T7b6_0),.din(w_dff_A_28gX06vb9_0),.clk(gclk));
	jdff dff_A_fl6lqKnc0_0(.dout(w_dff_A_28gX06vb9_0),.din(w_dff_A_fl6lqKnc0_0),.clk(gclk));
	jdff dff_A_yCH6Anye4_0(.dout(w_dff_A_fl6lqKnc0_0),.din(w_dff_A_yCH6Anye4_0),.clk(gclk));
	jdff dff_A_vcKH6jI99_0(.dout(w_dff_A_yCH6Anye4_0),.din(w_dff_A_vcKH6jI99_0),.clk(gclk));
	jdff dff_B_xSd0xNja4_1(.din(n256),.dout(w_dff_B_xSd0xNja4_1),.clk(gclk));
	jdff dff_B_vdGQaMzM1_1(.din(w_dff_B_xSd0xNja4_1),.dout(w_dff_B_vdGQaMzM1_1),.clk(gclk));
	jdff dff_B_fD9aqSh78_1(.din(w_dff_B_vdGQaMzM1_1),.dout(w_dff_B_fD9aqSh78_1),.clk(gclk));
	jdff dff_B_Pgl1Z3jn0_1(.din(w_dff_B_fD9aqSh78_1),.dout(w_dff_B_Pgl1Z3jn0_1),.clk(gclk));
	jdff dff_B_X6jdc4lQ9_1(.din(w_dff_B_Pgl1Z3jn0_1),.dout(w_dff_B_X6jdc4lQ9_1),.clk(gclk));
	jdff dff_B_TpjrsyKd5_1(.din(w_dff_B_X6jdc4lQ9_1),.dout(w_dff_B_TpjrsyKd5_1),.clk(gclk));
	jdff dff_B_lXsBvo7M9_1(.din(w_dff_B_TpjrsyKd5_1),.dout(w_dff_B_lXsBvo7M9_1),.clk(gclk));
	jdff dff_B_yHMnvESC0_0(.din(n283),.dout(w_dff_B_yHMnvESC0_0),.clk(gclk));
	jdff dff_B_zsKn8oIK0_0(.din(w_dff_B_yHMnvESC0_0),.dout(w_dff_B_zsKn8oIK0_0),.clk(gclk));
	jdff dff_B_j9aclB070_0(.din(w_dff_B_zsKn8oIK0_0),.dout(w_dff_B_j9aclB070_0),.clk(gclk));
	jdff dff_B_MJ3zYHxJ4_0(.din(w_dff_B_j9aclB070_0),.dout(w_dff_B_MJ3zYHxJ4_0),.clk(gclk));
	jdff dff_A_TBysbvAN3_1(.dout(w_n253_0[1]),.din(w_dff_A_TBysbvAN3_1),.clk(gclk));
	jdff dff_A_EkcHTEVP3_1(.dout(w_dff_A_TBysbvAN3_1),.din(w_dff_A_EkcHTEVP3_1),.clk(gclk));
	jdff dff_A_f6EYMW6q4_1(.dout(w_dff_A_EkcHTEVP3_1),.din(w_dff_A_f6EYMW6q4_1),.clk(gclk));
	jdff dff_A_uKSJ0XJD1_1(.dout(w_dff_A_f6EYMW6q4_1),.din(w_dff_A_uKSJ0XJD1_1),.clk(gclk));
	jdff dff_A_YeVc5UOD3_1(.dout(w_dff_A_uKSJ0XJD1_1),.din(w_dff_A_YeVc5UOD3_1),.clk(gclk));
	jdff dff_B_lwXOQWpt6_1(.din(n148),.dout(w_dff_B_lwXOQWpt6_1),.clk(gclk));
	jdff dff_B_QP2GGXYy0_0(.din(n212),.dout(w_dff_B_QP2GGXYy0_0),.clk(gclk));
	jdff dff_A_u0cATR1T7_0(.dout(w_n211_0[0]),.din(w_dff_A_u0cATR1T7_0),.clk(gclk));
	jdff dff_A_ImyC5g2F8_0(.dout(w_dff_A_u0cATR1T7_0),.din(w_dff_A_ImyC5g2F8_0),.clk(gclk));
	jdff dff_A_vMrf8DEo2_0(.dout(w_dff_A_ImyC5g2F8_0),.din(w_dff_A_vMrf8DEo2_0),.clk(gclk));
	jdff dff_A_UUKWveyy9_0(.dout(w_dff_A_vMrf8DEo2_0),.din(w_dff_A_UUKWveyy9_0),.clk(gclk));
	jdff dff_A_k72FSdyG6_0(.dout(w_dff_A_UUKWveyy9_0),.din(w_dff_A_k72FSdyG6_0),.clk(gclk));
	jdff dff_A_yja1jA0G3_0(.dout(w_dff_A_k72FSdyG6_0),.din(w_dff_A_yja1jA0G3_0),.clk(gclk));
	jdff dff_A_xpBVrZqa7_0(.dout(w_n209_0[0]),.din(w_dff_A_xpBVrZqa7_0),.clk(gclk));
	jdff dff_A_9Oa7IXWv2_0(.dout(w_dff_A_xpBVrZqa7_0),.din(w_dff_A_9Oa7IXWv2_0),.clk(gclk));
	jdff dff_A_oYOZjsMc3_0(.dout(w_dff_A_9Oa7IXWv2_0),.din(w_dff_A_oYOZjsMc3_0),.clk(gclk));
	jdff dff_A_3BB9E95F3_0(.dout(w_dff_A_oYOZjsMc3_0),.din(w_dff_A_3BB9E95F3_0),.clk(gclk));
	jdff dff_A_UiOlqUe47_0(.dout(w_dff_A_3BB9E95F3_0),.din(w_dff_A_UiOlqUe47_0),.clk(gclk));
	jdff dff_B_oB8hc8ck0_2(.din(n209),.dout(w_dff_B_oB8hc8ck0_2),.clk(gclk));
	jdff dff_B_EnUAYsxq2_2(.din(w_dff_B_oB8hc8ck0_2),.dout(w_dff_B_EnUAYsxq2_2),.clk(gclk));
	jdff dff_B_RCcX7fqy0_2(.din(w_dff_B_EnUAYsxq2_2),.dout(w_dff_B_RCcX7fqy0_2),.clk(gclk));
	jdff dff_B_JSIR8IyY8_2(.din(w_dff_B_RCcX7fqy0_2),.dout(w_dff_B_JSIR8IyY8_2),.clk(gclk));
	jdff dff_B_oyNdbX3W0_2(.din(w_dff_B_JSIR8IyY8_2),.dout(w_dff_B_oyNdbX3W0_2),.clk(gclk));
	jdff dff_B_FhvYs9X27_2(.din(w_dff_B_oyNdbX3W0_2),.dout(w_dff_B_FhvYs9X27_2),.clk(gclk));
	jdff dff_B_j2r1NXJu1_2(.din(w_dff_B_FhvYs9X27_2),.dout(w_dff_B_j2r1NXJu1_2),.clk(gclk));
	jdff dff_B_MUJwKZYJ3_2(.din(w_dff_B_j2r1NXJu1_2),.dout(w_dff_B_MUJwKZYJ3_2),.clk(gclk));
	jdff dff_B_0W3BZIxm2_2(.din(w_dff_B_MUJwKZYJ3_2),.dout(w_dff_B_0W3BZIxm2_2),.clk(gclk));
	jdff dff_B_RW7WA03W4_2(.din(w_dff_B_0W3BZIxm2_2),.dout(w_dff_B_RW7WA03W4_2),.clk(gclk));
	jdff dff_B_RIqo5qxR1_2(.din(w_dff_B_RW7WA03W4_2),.dout(w_dff_B_RIqo5qxR1_2),.clk(gclk));
	jdff dff_B_nG7Wb0xO8_2(.din(w_dff_B_RIqo5qxR1_2),.dout(w_dff_B_nG7Wb0xO8_2),.clk(gclk));
	jdff dff_B_sDsCO4mc0_2(.din(w_dff_B_nG7Wb0xO8_2),.dout(w_dff_B_sDsCO4mc0_2),.clk(gclk));
	jdff dff_B_6RajPZ225_2(.din(w_dff_B_sDsCO4mc0_2),.dout(w_dff_B_6RajPZ225_2),.clk(gclk));
	jdff dff_A_QQWtvWjU9_0(.dout(w_n206_0[0]),.din(w_dff_A_QQWtvWjU9_0),.clk(gclk));
	jdff dff_A_wByZYIIs9_0(.dout(w_dff_A_QQWtvWjU9_0),.din(w_dff_A_wByZYIIs9_0),.clk(gclk));
	jdff dff_A_TPdwe9sJ7_0(.dout(w_dff_A_wByZYIIs9_0),.din(w_dff_A_TPdwe9sJ7_0),.clk(gclk));
	jdff dff_A_QdplOECX8_0(.dout(w_dff_A_TPdwe9sJ7_0),.din(w_dff_A_QdplOECX8_0),.clk(gclk));
	jdff dff_A_iK6c3yTo1_0(.dout(w_dff_A_QdplOECX8_0),.din(w_dff_A_iK6c3yTo1_0),.clk(gclk));
	jdff dff_A_vZXliEu80_0(.dout(w_dff_A_iK6c3yTo1_0),.din(w_dff_A_vZXliEu80_0),.clk(gclk));
	jdff dff_A_nfzWIevA8_0(.dout(w_n204_0[0]),.din(w_dff_A_nfzWIevA8_0),.clk(gclk));
	jdff dff_A_Gt0gk1ij9_0(.dout(w_dff_A_nfzWIevA8_0),.din(w_dff_A_Gt0gk1ij9_0),.clk(gclk));
	jdff dff_A_v25vqoHc5_0(.dout(w_dff_A_Gt0gk1ij9_0),.din(w_dff_A_v25vqoHc5_0),.clk(gclk));
	jdff dff_A_jyvsJMA14_0(.dout(w_dff_A_v25vqoHc5_0),.din(w_dff_A_jyvsJMA14_0),.clk(gclk));
	jdff dff_A_OYZRaIO26_0(.dout(w_dff_A_jyvsJMA14_0),.din(w_dff_A_OYZRaIO26_0),.clk(gclk));
	jdff dff_B_9SOwJs438_2(.din(n204),.dout(w_dff_B_9SOwJs438_2),.clk(gclk));
	jdff dff_B_4pVfDyK01_2(.din(w_dff_B_9SOwJs438_2),.dout(w_dff_B_4pVfDyK01_2),.clk(gclk));
	jdff dff_B_LYcO2Dkx2_2(.din(w_dff_B_4pVfDyK01_2),.dout(w_dff_B_LYcO2Dkx2_2),.clk(gclk));
	jdff dff_B_jskmvLJw5_2(.din(w_dff_B_LYcO2Dkx2_2),.dout(w_dff_B_jskmvLJw5_2),.clk(gclk));
	jdff dff_B_mkvCYlCP0_2(.din(w_dff_B_jskmvLJw5_2),.dout(w_dff_B_mkvCYlCP0_2),.clk(gclk));
	jdff dff_B_b28DU7yA4_2(.din(w_dff_B_mkvCYlCP0_2),.dout(w_dff_B_b28DU7yA4_2),.clk(gclk));
	jdff dff_B_44SDUm2A6_2(.din(w_dff_B_b28DU7yA4_2),.dout(w_dff_B_44SDUm2A6_2),.clk(gclk));
	jdff dff_B_fH9OvtBY1_2(.din(w_dff_B_44SDUm2A6_2),.dout(w_dff_B_fH9OvtBY1_2),.clk(gclk));
	jdff dff_B_jDSVQKhW6_2(.din(w_dff_B_fH9OvtBY1_2),.dout(w_dff_B_jDSVQKhW6_2),.clk(gclk));
	jdff dff_B_2FL64ZH11_2(.din(w_dff_B_jDSVQKhW6_2),.dout(w_dff_B_2FL64ZH11_2),.clk(gclk));
	jdff dff_B_YDsxh9a20_2(.din(w_dff_B_2FL64ZH11_2),.dout(w_dff_B_YDsxh9a20_2),.clk(gclk));
	jdff dff_B_If33qaQs2_2(.din(w_dff_B_YDsxh9a20_2),.dout(w_dff_B_If33qaQs2_2),.clk(gclk));
	jdff dff_B_SPDZuxGI7_2(.din(w_dff_B_If33qaQs2_2),.dout(w_dff_B_SPDZuxGI7_2),.clk(gclk));
	jdff dff_B_Wbgx3rRy1_2(.din(w_dff_B_SPDZuxGI7_2),.dout(w_dff_B_Wbgx3rRy1_2),.clk(gclk));
	jdff dff_B_6wTHl1Ox4_1(.din(n194),.dout(w_dff_B_6wTHl1Ox4_1),.clk(gclk));
	jdff dff_B_rR2VyiWp9_1(.din(w_dff_B_6wTHl1Ox4_1),.dout(w_dff_B_rR2VyiWp9_1),.clk(gclk));
	jdff dff_B_JGmtUXc49_1(.din(w_dff_B_rR2VyiWp9_1),.dout(w_dff_B_JGmtUXc49_1),.clk(gclk));
	jdff dff_B_NLmdutY57_1(.din(w_dff_B_JGmtUXc49_1),.dout(w_dff_B_NLmdutY57_1),.clk(gclk));
	jdff dff_B_vEVx6HVV3_1(.din(w_dff_B_NLmdutY57_1),.dout(w_dff_B_vEVx6HVV3_1),.clk(gclk));
	jdff dff_B_gPz9X9k84_1(.din(w_dff_B_vEVx6HVV3_1),.dout(w_dff_B_gPz9X9k84_1),.clk(gclk));
	jdff dff_B_C87uUjoD4_1(.din(w_dff_B_gPz9X9k84_1),.dout(w_dff_B_C87uUjoD4_1),.clk(gclk));
	jdff dff_B_cOB7HS469_1(.din(w_dff_B_C87uUjoD4_1),.dout(w_dff_B_cOB7HS469_1),.clk(gclk));
	jdff dff_B_HHhJVLGv9_1(.din(w_dff_B_cOB7HS469_1),.dout(w_dff_B_HHhJVLGv9_1),.clk(gclk));
	jdff dff_B_MUwpo5Z39_1(.din(w_dff_B_HHhJVLGv9_1),.dout(w_dff_B_MUwpo5Z39_1),.clk(gclk));
	jdff dff_B_oJRZRVc22_1(.din(w_dff_B_MUwpo5Z39_1),.dout(w_dff_B_oJRZRVc22_1),.clk(gclk));
	jdff dff_B_Ye824Mux6_1(.din(w_dff_B_oJRZRVc22_1),.dout(w_dff_B_Ye824Mux6_1),.clk(gclk));
	jdff dff_B_eYelOqLP8_1(.din(w_dff_B_Ye824Mux6_1),.dout(w_dff_B_eYelOqLP8_1),.clk(gclk));
	jdff dff_B_ba0Ln3Us5_1(.din(w_dff_B_eYelOqLP8_1),.dout(w_dff_B_ba0Ln3Us5_1),.clk(gclk));
	jdff dff_B_YjHmnK9K0_1(.din(n190),.dout(w_dff_B_YjHmnK9K0_1),.clk(gclk));
	jdff dff_B_sIB6d5EG7_1(.din(w_dff_B_YjHmnK9K0_1),.dout(w_dff_B_sIB6d5EG7_1),.clk(gclk));
	jdff dff_B_vwMLsJ4L1_1(.din(w_dff_B_sIB6d5EG7_1),.dout(w_dff_B_vwMLsJ4L1_1),.clk(gclk));
	jdff dff_B_83viOYOt7_1(.din(w_dff_B_vwMLsJ4L1_1),.dout(w_dff_B_83viOYOt7_1),.clk(gclk));
	jdff dff_B_Mkb0lWqA0_1(.din(w_dff_B_83viOYOt7_1),.dout(w_dff_B_Mkb0lWqA0_1),.clk(gclk));
	jdff dff_B_9Pr8HhzR3_1(.din(w_dff_B_Mkb0lWqA0_1),.dout(w_dff_B_9Pr8HhzR3_1),.clk(gclk));
	jdff dff_B_uCHmCYaJ6_1(.din(w_dff_B_9Pr8HhzR3_1),.dout(w_dff_B_uCHmCYaJ6_1),.clk(gclk));
	jdff dff_B_i6f3iihH5_1(.din(w_dff_B_uCHmCYaJ6_1),.dout(w_dff_B_i6f3iihH5_1),.clk(gclk));
	jdff dff_B_BFMrnTK47_1(.din(w_dff_B_i6f3iihH5_1),.dout(w_dff_B_BFMrnTK47_1),.clk(gclk));
	jdff dff_B_r3aWFr4W3_1(.din(w_dff_B_BFMrnTK47_1),.dout(w_dff_B_r3aWFr4W3_1),.clk(gclk));
	jdff dff_B_PrGcamn13_1(.din(w_dff_B_r3aWFr4W3_1),.dout(w_dff_B_PrGcamn13_1),.clk(gclk));
	jdff dff_B_MUbeO81a9_1(.din(w_dff_B_PrGcamn13_1),.dout(w_dff_B_MUbeO81a9_1),.clk(gclk));
	jdff dff_B_kkv2ItSd5_1(.din(w_dff_B_MUbeO81a9_1),.dout(w_dff_B_kkv2ItSd5_1),.clk(gclk));
	jdff dff_B_qspT91km1_1(.din(w_dff_B_kkv2ItSd5_1),.dout(w_dff_B_qspT91km1_1),.clk(gclk));
	jdff dff_A_PWdLB2rj7_0(.dout(w_n185_0[0]),.din(w_dff_A_PWdLB2rj7_0),.clk(gclk));
	jdff dff_A_a91x22Jj1_0(.dout(w_dff_A_PWdLB2rj7_0),.din(w_dff_A_a91x22Jj1_0),.clk(gclk));
	jdff dff_A_AkvgC7Sw9_0(.dout(w_dff_A_a91x22Jj1_0),.din(w_dff_A_AkvgC7Sw9_0),.clk(gclk));
	jdff dff_A_4gXPYZx31_0(.dout(w_dff_A_AkvgC7Sw9_0),.din(w_dff_A_4gXPYZx31_0),.clk(gclk));
	jdff dff_A_odEaCUEE8_0(.dout(w_dff_A_4gXPYZx31_0),.din(w_dff_A_odEaCUEE8_0),.clk(gclk));
	jdff dff_B_d4lvTgFq6_2(.din(n185),.dout(w_dff_B_d4lvTgFq6_2),.clk(gclk));
	jdff dff_B_nEgizuqm5_2(.din(w_dff_B_d4lvTgFq6_2),.dout(w_dff_B_nEgizuqm5_2),.clk(gclk));
	jdff dff_B_eLgSdFBi3_2(.din(w_dff_B_nEgizuqm5_2),.dout(w_dff_B_eLgSdFBi3_2),.clk(gclk));
	jdff dff_B_RNKea2g00_2(.din(w_dff_B_eLgSdFBi3_2),.dout(w_dff_B_RNKea2g00_2),.clk(gclk));
	jdff dff_B_SLgAIdx72_2(.din(w_dff_B_RNKea2g00_2),.dout(w_dff_B_SLgAIdx72_2),.clk(gclk));
	jdff dff_B_bFYxaDpP3_2(.din(w_dff_B_SLgAIdx72_2),.dout(w_dff_B_bFYxaDpP3_2),.clk(gclk));
	jdff dff_B_PLBUo2M06_2(.din(w_dff_B_bFYxaDpP3_2),.dout(w_dff_B_PLBUo2M06_2),.clk(gclk));
	jdff dff_B_FcCrHuge5_2(.din(w_dff_B_PLBUo2M06_2),.dout(w_dff_B_FcCrHuge5_2),.clk(gclk));
	jdff dff_B_yQ9uAffr2_2(.din(w_dff_B_FcCrHuge5_2),.dout(w_dff_B_yQ9uAffr2_2),.clk(gclk));
	jdff dff_B_gEIczuo23_2(.din(w_dff_B_yQ9uAffr2_2),.dout(w_dff_B_gEIczuo23_2),.clk(gclk));
	jdff dff_B_EVwBVohv4_2(.din(w_dff_B_gEIczuo23_2),.dout(w_dff_B_EVwBVohv4_2),.clk(gclk));
	jdff dff_B_pbP9fPTx8_2(.din(w_dff_B_EVwBVohv4_2),.dout(w_dff_B_pbP9fPTx8_2),.clk(gclk));
	jdff dff_B_13lMLyaC0_2(.din(w_dff_B_pbP9fPTx8_2),.dout(w_dff_B_13lMLyaC0_2),.clk(gclk));
	jdff dff_B_SS5Ks74t8_2(.din(w_dff_B_13lMLyaC0_2),.dout(w_dff_B_SS5Ks74t8_2),.clk(gclk));
	jdff dff_B_qVZ41wor8_2(.din(n281),.dout(w_dff_B_qVZ41wor8_2),.clk(gclk));
	jdff dff_A_B2Z8rNqE5_0(.dout(w_n149_0[0]),.din(w_dff_A_B2Z8rNqE5_0),.clk(gclk));
	jdff dff_A_4p99zO6p2_0(.dout(w_dff_A_B2Z8rNqE5_0),.din(w_dff_A_4p99zO6p2_0),.clk(gclk));
	jdff dff_A_qCrNttSH4_0(.dout(w_dff_A_4p99zO6p2_0),.din(w_dff_A_qCrNttSH4_0),.clk(gclk));
	jdff dff_A_GUdBd9mu6_0(.dout(w_dff_A_qCrNttSH4_0),.din(w_dff_A_GUdBd9mu6_0),.clk(gclk));
	jdff dff_A_nuSDMEPB6_0(.dout(w_dff_A_GUdBd9mu6_0),.din(w_dff_A_nuSDMEPB6_0),.clk(gclk));
	jdff dff_B_rCZn44ug3_2(.din(n149),.dout(w_dff_B_rCZn44ug3_2),.clk(gclk));
	jdff dff_B_UBOJ8tzV7_2(.din(w_dff_B_rCZn44ug3_2),.dout(w_dff_B_UBOJ8tzV7_2),.clk(gclk));
	jdff dff_B_Ivo7Af3v1_2(.din(w_dff_B_UBOJ8tzV7_2),.dout(w_dff_B_Ivo7Af3v1_2),.clk(gclk));
	jdff dff_B_GHIdF3Hc5_2(.din(w_dff_B_Ivo7Af3v1_2),.dout(w_dff_B_GHIdF3Hc5_2),.clk(gclk));
	jdff dff_B_bn2DgXrP1_2(.din(w_dff_B_GHIdF3Hc5_2),.dout(w_dff_B_bn2DgXrP1_2),.clk(gclk));
	jdff dff_B_mFyrlaSO8_2(.din(w_dff_B_bn2DgXrP1_2),.dout(w_dff_B_mFyrlaSO8_2),.clk(gclk));
	jdff dff_B_5RLFVkOf8_2(.din(w_dff_B_mFyrlaSO8_2),.dout(w_dff_B_5RLFVkOf8_2),.clk(gclk));
	jdff dff_B_qrsygGXs1_2(.din(w_dff_B_5RLFVkOf8_2),.dout(w_dff_B_qrsygGXs1_2),.clk(gclk));
	jdff dff_B_eTK4Z6O22_2(.din(w_dff_B_qrsygGXs1_2),.dout(w_dff_B_eTK4Z6O22_2),.clk(gclk));
	jdff dff_B_07mkwv4R7_2(.din(w_dff_B_eTK4Z6O22_2),.dout(w_dff_B_07mkwv4R7_2),.clk(gclk));
	jdff dff_B_Ob73atk08_2(.din(w_dff_B_07mkwv4R7_2),.dout(w_dff_B_Ob73atk08_2),.clk(gclk));
	jdff dff_B_tEEgs9xm5_2(.din(w_dff_B_Ob73atk08_2),.dout(w_dff_B_tEEgs9xm5_2),.clk(gclk));
	jdff dff_B_prjuiRUh1_2(.din(w_dff_B_tEEgs9xm5_2),.dout(w_dff_B_prjuiRUh1_2),.clk(gclk));
	jdff dff_B_NBVsFsuc1_2(.din(w_dff_B_prjuiRUh1_2),.dout(w_dff_B_NBVsFsuc1_2),.clk(gclk));
	jdff dff_A_oR4OMqBV7_0(.dout(w_n183_0[0]),.din(w_dff_A_oR4OMqBV7_0),.clk(gclk));
	jdff dff_A_3IivIiSm3_0(.dout(w_dff_A_oR4OMqBV7_0),.din(w_dff_A_3IivIiSm3_0),.clk(gclk));
	jdff dff_A_gOR6YDZr9_0(.dout(w_dff_A_3IivIiSm3_0),.din(w_dff_A_gOR6YDZr9_0),.clk(gclk));
	jdff dff_A_ChFNvTk20_0(.dout(w_dff_A_gOR6YDZr9_0),.din(w_dff_A_ChFNvTk20_0),.clk(gclk));
	jdff dff_A_pGeBBPKK0_0(.dout(w_dff_A_ChFNvTk20_0),.din(w_dff_A_pGeBBPKK0_0),.clk(gclk));
	jdff dff_A_maON4xc73_0(.dout(w_dff_A_pGeBBPKK0_0),.din(w_dff_A_maON4xc73_0),.clk(gclk));
	jdff dff_A_HY831AbW1_0(.dout(w_n271_0[0]),.din(w_dff_A_HY831AbW1_0),.clk(gclk));
	jdff dff_A_YT86EpGx6_0(.dout(w_dff_A_HY831AbW1_0),.din(w_dff_A_YT86EpGx6_0),.clk(gclk));
	jdff dff_A_qhDd3nSX7_0(.dout(w_dff_A_YT86EpGx6_0),.din(w_dff_A_qhDd3nSX7_0),.clk(gclk));
	jdff dff_B_BSaj4DT15_1(.din(n217),.dout(w_dff_B_BSaj4DT15_1),.clk(gclk));
	jdff dff_B_I2UqC6LA6_0(.din(n243),.dout(w_dff_B_I2UqC6LA6_0),.clk(gclk));
	jdff dff_A_XrUML48z4_0(.dout(w_n230_0[0]),.din(w_dff_A_XrUML48z4_0),.clk(gclk));
	jdff dff_A_M5UfqVuK0_0(.dout(w_dff_A_XrUML48z4_0),.din(w_dff_A_M5UfqVuK0_0),.clk(gclk));
	jdff dff_A_N8AXmMWc8_0(.dout(w_dff_A_M5UfqVuK0_0),.din(w_dff_A_N8AXmMWc8_0),.clk(gclk));
	jdff dff_A_MOH7kBoI3_0(.dout(w_dff_A_N8AXmMWc8_0),.din(w_dff_A_MOH7kBoI3_0),.clk(gclk));
	jdff dff_A_Z6GXP7BJ3_0(.dout(w_dff_A_MOH7kBoI3_0),.din(w_dff_A_Z6GXP7BJ3_0),.clk(gclk));
	jdff dff_A_ynRIomY82_0(.dout(w_dff_A_Z6GXP7BJ3_0),.din(w_dff_A_ynRIomY82_0),.clk(gclk));
	jdff dff_A_ayfftHHh7_0(.dout(w_n227_0[0]),.din(w_dff_A_ayfftHHh7_0),.clk(gclk));
	jdff dff_A_P3ID5Ro71_0(.dout(w_dff_A_ayfftHHh7_0),.din(w_dff_A_P3ID5Ro71_0),.clk(gclk));
	jdff dff_A_2pu4Shy09_0(.dout(w_dff_A_P3ID5Ro71_0),.din(w_dff_A_2pu4Shy09_0),.clk(gclk));
	jdff dff_A_nD7T96vq3_0(.dout(w_dff_A_2pu4Shy09_0),.din(w_dff_A_nD7T96vq3_0),.clk(gclk));
	jdff dff_A_hve5nfuh0_0(.dout(w_dff_A_nD7T96vq3_0),.din(w_dff_A_hve5nfuh0_0),.clk(gclk));
	jdff dff_A_r3X03Ksn2_0(.dout(w_dff_A_hve5nfuh0_0),.din(w_dff_A_r3X03Ksn2_0),.clk(gclk));
	jdff dff_B_rXmzRcqG0_1(.din(n221),.dout(w_dff_B_rXmzRcqG0_1),.clk(gclk));
	jdff dff_B_8WQo3Ph79_1(.din(w_dff_B_rXmzRcqG0_1),.dout(w_dff_B_8WQo3Ph79_1),.clk(gclk));
	jdff dff_B_2Eq2SDi60_1(.din(w_dff_B_8WQo3Ph79_1),.dout(w_dff_B_2Eq2SDi60_1),.clk(gclk));
	jdff dff_B_A74Dl4Lh8_1(.din(w_dff_B_2Eq2SDi60_1),.dout(w_dff_B_A74Dl4Lh8_1),.clk(gclk));
	jdff dff_B_BjofQXO58_1(.din(w_dff_B_A74Dl4Lh8_1),.dout(w_dff_B_BjofQXO58_1),.clk(gclk));
	jdff dff_A_odnU3JUb8_1(.dout(w_n147_0[1]),.din(w_dff_A_odnU3JUb8_1),.clk(gclk));
	jdff dff_B_LLRggoRx9_0(.din(n146),.dout(w_dff_B_LLRggoRx9_0),.clk(gclk));
	jdff dff_B_y4l3xiDs4_0(.din(w_dff_B_LLRggoRx9_0),.dout(w_dff_B_y4l3xiDs4_0),.clk(gclk));
	jdff dff_B_42Pvyqep0_0(.din(w_dff_B_y4l3xiDs4_0),.dout(w_dff_B_42Pvyqep0_0),.clk(gclk));
	jdff dff_B_qUCQ2tVg4_0(.din(w_dff_B_42Pvyqep0_0),.dout(w_dff_B_qUCQ2tVg4_0),.clk(gclk));
	jdff dff_B_ZGg3Kssf1_0(.din(w_dff_B_qUCQ2tVg4_0),.dout(w_dff_B_ZGg3Kssf1_0),.clk(gclk));
	jdff dff_B_semhg0XA5_0(.din(w_dff_B_ZGg3Kssf1_0),.dout(w_dff_B_semhg0XA5_0),.clk(gclk));
	jdff dff_A_Izc7gCgG6_0(.dout(w_n141_0[0]),.din(w_dff_A_Izc7gCgG6_0),.clk(gclk));
	jdff dff_A_szyTS6Oa8_0(.dout(w_n200_0[0]),.din(w_dff_A_szyTS6Oa8_0),.clk(gclk));
	jdff dff_A_51DMl5vl0_0(.dout(w_dff_A_szyTS6Oa8_0),.din(w_dff_A_51DMl5vl0_0),.clk(gclk));
	jdff dff_A_CT5UaxRu8_0(.dout(w_dff_A_51DMl5vl0_0),.din(w_dff_A_CT5UaxRu8_0),.clk(gclk));
	jdff dff_A_364EBhxd6_0(.dout(w_dff_A_CT5UaxRu8_0),.din(w_dff_A_364EBhxd6_0),.clk(gclk));
	jdff dff_A_63oZoyoF8_0(.dout(w_dff_A_364EBhxd6_0),.din(w_dff_A_63oZoyoF8_0),.clk(gclk));
	jdff dff_B_XlN4GTGu6_2(.din(n200),.dout(w_dff_B_XlN4GTGu6_2),.clk(gclk));
	jdff dff_B_GI47OmJT5_2(.din(w_dff_B_XlN4GTGu6_2),.dout(w_dff_B_GI47OmJT5_2),.clk(gclk));
	jdff dff_B_TS1nPMOJ9_2(.din(w_dff_B_GI47OmJT5_2),.dout(w_dff_B_TS1nPMOJ9_2),.clk(gclk));
	jdff dff_B_xiAKdumT6_2(.din(w_dff_B_TS1nPMOJ9_2),.dout(w_dff_B_xiAKdumT6_2),.clk(gclk));
	jdff dff_B_h4k8gdO21_2(.din(w_dff_B_xiAKdumT6_2),.dout(w_dff_B_h4k8gdO21_2),.clk(gclk));
	jdff dff_B_xKEzMDkM2_2(.din(w_dff_B_h4k8gdO21_2),.dout(w_dff_B_xKEzMDkM2_2),.clk(gclk));
	jdff dff_B_3JvXLvY50_2(.din(w_dff_B_xKEzMDkM2_2),.dout(w_dff_B_3JvXLvY50_2),.clk(gclk));
	jdff dff_B_JzZmHrNh0_2(.din(w_dff_B_3JvXLvY50_2),.dout(w_dff_B_JzZmHrNh0_2),.clk(gclk));
	jdff dff_B_kx7Iet5W7_2(.din(w_dff_B_JzZmHrNh0_2),.dout(w_dff_B_kx7Iet5W7_2),.clk(gclk));
	jdff dff_B_BgT0exiJ8_2(.din(w_dff_B_kx7Iet5W7_2),.dout(w_dff_B_BgT0exiJ8_2),.clk(gclk));
	jdff dff_B_59OVdDxG3_2(.din(w_dff_B_BgT0exiJ8_2),.dout(w_dff_B_59OVdDxG3_2),.clk(gclk));
	jdff dff_B_AtgwB8iE9_2(.din(w_dff_B_59OVdDxG3_2),.dout(w_dff_B_AtgwB8iE9_2),.clk(gclk));
	jdff dff_B_lddyxjpx2_2(.din(w_dff_B_AtgwB8iE9_2),.dout(w_dff_B_lddyxjpx2_2),.clk(gclk));
	jdff dff_B_YtIYVhHE4_2(.din(w_dff_B_lddyxjpx2_2),.dout(w_dff_B_YtIYVhHE4_2),.clk(gclk));
	jdff dff_A_sKoCC3zh9_0(.dout(w_n202_0[0]),.din(w_dff_A_sKoCC3zh9_0),.clk(gclk));
	jdff dff_A_NrIqP14M4_0(.dout(w_dff_A_sKoCC3zh9_0),.din(w_dff_A_NrIqP14M4_0),.clk(gclk));
	jdff dff_A_2KzzHUxH0_0(.dout(w_dff_A_NrIqP14M4_0),.din(w_dff_A_2KzzHUxH0_0),.clk(gclk));
	jdff dff_A_BpFrD0KW4_0(.dout(w_dff_A_2KzzHUxH0_0),.din(w_dff_A_BpFrD0KW4_0),.clk(gclk));
	jdff dff_A_1bTNjptD8_0(.dout(w_dff_A_BpFrD0KW4_0),.din(w_dff_A_1bTNjptD8_0),.clk(gclk));
	jdff dff_A_gYVfYYle3_0(.dout(w_dff_A_1bTNjptD8_0),.din(w_dff_A_gYVfYYle3_0),.clk(gclk));
	jdff dff_B_0zfirOu97_1(.din(n168),.dout(w_dff_B_0zfirOu97_1),.clk(gclk));
	jdff dff_B_o9ZLIsAW3_1(.din(n171),.dout(w_dff_B_o9ZLIsAW3_1),.clk(gclk));
	jdff dff_A_4uHBuKwJ9_0(.dout(w_n173_0[0]),.din(w_dff_A_4uHBuKwJ9_0),.clk(gclk));
	jdff dff_A_Zydon2Kb9_0(.dout(w_dff_A_4uHBuKwJ9_0),.din(w_dff_A_Zydon2Kb9_0),.clk(gclk));
	jdff dff_A_RP8PBlkw9_0(.dout(w_dff_A_Zydon2Kb9_0),.din(w_dff_A_RP8PBlkw9_0),.clk(gclk));
	jdff dff_A_q3qz3Tvs6_0(.dout(w_dff_A_RP8PBlkw9_0),.din(w_dff_A_q3qz3Tvs6_0),.clk(gclk));
	jdff dff_A_jJaiJ6vH3_0(.dout(w_dff_A_q3qz3Tvs6_0),.din(w_dff_A_jJaiJ6vH3_0),.clk(gclk));
	jdff dff_A_DnX4lryc8_0(.dout(w_dff_A_jJaiJ6vH3_0),.din(w_dff_A_DnX4lryc8_0),.clk(gclk));
	jdff dff_A_EIG2JM9W2_0(.dout(w_n170_0[0]),.din(w_dff_A_EIG2JM9W2_0),.clk(gclk));
	jdff dff_A_4E7vCqTU1_0(.dout(w_dff_A_EIG2JM9W2_0),.din(w_dff_A_4E7vCqTU1_0),.clk(gclk));
	jdff dff_A_vAOwm7wp0_0(.dout(w_dff_A_4E7vCqTU1_0),.din(w_dff_A_vAOwm7wp0_0),.clk(gclk));
	jdff dff_A_l5z1HdZr0_0(.dout(w_dff_A_vAOwm7wp0_0),.din(w_dff_A_l5z1HdZr0_0),.clk(gclk));
	jdff dff_A_f6I0oko83_0(.dout(w_dff_A_l5z1HdZr0_0),.din(w_dff_A_f6I0oko83_0),.clk(gclk));
	jdff dff_A_to77wHFK6_0(.dout(w_dff_A_f6I0oko83_0),.din(w_dff_A_to77wHFK6_0),.clk(gclk));
	jdff dff_B_Lz8LZPOU1_1(.din(n154),.dout(w_dff_B_Lz8LZPOU1_1),.clk(gclk));
	jdff dff_B_E5NdmgxO1_0(.din(n165),.dout(w_dff_B_E5NdmgxO1_0),.clk(gclk));
	jdff dff_A_bSXelBOE6_0(.dout(w_n164_0[0]),.din(w_dff_A_bSXelBOE6_0),.clk(gclk));
	jdff dff_A_wGzVZ1eT5_0(.dout(w_dff_A_bSXelBOE6_0),.din(w_dff_A_wGzVZ1eT5_0),.clk(gclk));
	jdff dff_A_YD51Llv40_0(.dout(w_dff_A_wGzVZ1eT5_0),.din(w_dff_A_YD51Llv40_0),.clk(gclk));
	jdff dff_A_S54NF0lG5_0(.dout(w_dff_A_YD51Llv40_0),.din(w_dff_A_S54NF0lG5_0),.clk(gclk));
	jdff dff_A_wM5s8YQ61_0(.dout(w_dff_A_S54NF0lG5_0),.din(w_dff_A_wM5s8YQ61_0),.clk(gclk));
	jdff dff_A_jBN2c32x7_0(.dout(w_dff_A_wM5s8YQ61_0),.din(w_dff_A_jBN2c32x7_0),.clk(gclk));
	jdff dff_B_KZlWoY7g0_1(.din(n162),.dout(w_dff_B_KZlWoY7g0_1),.clk(gclk));
	jdff dff_B_umaKUS525_1(.din(w_dff_B_KZlWoY7g0_1),.dout(w_dff_B_umaKUS525_1),.clk(gclk));
	jdff dff_B_dTnArEg17_1(.din(w_dff_B_umaKUS525_1),.dout(w_dff_B_dTnArEg17_1),.clk(gclk));
	jdff dff_B_9duBFX6L7_1(.din(w_dff_B_dTnArEg17_1),.dout(w_dff_B_9duBFX6L7_1),.clk(gclk));
	jdff dff_B_85G61gFE4_1(.din(w_dff_B_9duBFX6L7_1),.dout(w_dff_B_85G61gFE4_1),.clk(gclk));
	jdff dff_B_bgBLIMi30_1(.din(w_dff_B_85G61gFE4_1),.dout(w_dff_B_bgBLIMi30_1),.clk(gclk));
	jdff dff_A_gBtP3tnQ1_0(.dout(w_n159_0[0]),.din(w_dff_A_gBtP3tnQ1_0),.clk(gclk));
	jdff dff_A_yu0xCXRO9_0(.dout(w_dff_A_gBtP3tnQ1_0),.din(w_dff_A_yu0xCXRO9_0),.clk(gclk));
	jdff dff_A_ia1CDLVJ7_0(.dout(w_dff_A_yu0xCXRO9_0),.din(w_dff_A_ia1CDLVJ7_0),.clk(gclk));
	jdff dff_A_xdUMVmIc8_0(.dout(w_dff_A_ia1CDLVJ7_0),.din(w_dff_A_xdUMVmIc8_0),.clk(gclk));
	jdff dff_A_CxuA7Qma4_0(.dout(w_dff_A_xdUMVmIc8_0),.din(w_dff_A_CxuA7Qma4_0),.clk(gclk));
	jdff dff_A_3fldbpnW8_0(.dout(w_dff_A_CxuA7Qma4_0),.din(w_dff_A_3fldbpnW8_0),.clk(gclk));
	jdff dff_A_4k5SSRp42_0(.dout(w_n156_0[0]),.din(w_dff_A_4k5SSRp42_0),.clk(gclk));
	jdff dff_A_VfBKlTKA0_0(.dout(w_dff_A_4k5SSRp42_0),.din(w_dff_A_VfBKlTKA0_0),.clk(gclk));
	jdff dff_A_MJUiek4X8_0(.dout(w_dff_A_VfBKlTKA0_0),.din(w_dff_A_MJUiek4X8_0),.clk(gclk));
	jdff dff_A_DIKNDfFh7_0(.dout(w_dff_A_MJUiek4X8_0),.din(w_dff_A_DIKNDfFh7_0),.clk(gclk));
	jdff dff_A_Uic0RTvi3_0(.dout(w_dff_A_DIKNDfFh7_0),.din(w_dff_A_Uic0RTvi3_0),.clk(gclk));
	jdff dff_A_HKPFXnOD2_0(.dout(w_dff_A_Uic0RTvi3_0),.din(w_dff_A_HKPFXnOD2_0),.clk(gclk));
	jdff dff_A_WWUwobV88_1(.dout(w_n138_0[1]),.din(w_dff_A_WWUwobV88_1),.clk(gclk));
	jdff dff_A_SapwMk784_1(.dout(w_dff_A_WWUwobV88_1),.din(w_dff_A_SapwMk784_1),.clk(gclk));
	jdff dff_A_3zICCvER9_1(.dout(w_dff_A_SapwMk784_1),.din(w_dff_A_3zICCvER9_1),.clk(gclk));
	jdff dff_A_KKlfiE8u7_1(.dout(w_dff_A_3zICCvER9_1),.din(w_dff_A_KKlfiE8u7_1),.clk(gclk));
	jdff dff_A_jGi9B9Xj8_1(.dout(w_dff_A_KKlfiE8u7_1),.din(w_dff_A_jGi9B9Xj8_1),.clk(gclk));
	jdff dff_A_yYIsqFhH3_1(.dout(w_dff_A_jGi9B9Xj8_1),.din(w_dff_A_yYIsqFhH3_1),.clk(gclk));
	jdff dff_A_XZ4IyHh82_0(.dout(w_n151_0[0]),.din(w_dff_A_XZ4IyHh82_0),.clk(gclk));
	jdff dff_A_tr7D1iqO5_0(.dout(w_dff_A_XZ4IyHh82_0),.din(w_dff_A_tr7D1iqO5_0),.clk(gclk));
	jdff dff_A_zErVdf3p5_0(.dout(w_dff_A_tr7D1iqO5_0),.din(w_dff_A_zErVdf3p5_0),.clk(gclk));
	jdff dff_A_xR8dBdnR1_0(.dout(w_dff_A_zErVdf3p5_0),.din(w_dff_A_xR8dBdnR1_0),.clk(gclk));
	jdff dff_A_bc4wkJP60_0(.dout(w_dff_A_xR8dBdnR1_0),.din(w_dff_A_bc4wkJP60_0),.clk(gclk));
	jdff dff_A_9BNznCqm5_0(.dout(w_dff_A_bc4wkJP60_0),.din(w_dff_A_9BNznCqm5_0),.clk(gclk));
	jdff dff_A_toHHMGld8_1(.dout(w_dff_A_hMAXkXG39_0),.din(w_dff_A_toHHMGld8_1),.clk(gclk));
	jdff dff_A_hMAXkXG39_0(.dout(w_dff_A_JjcMM0Nf4_0),.din(w_dff_A_hMAXkXG39_0),.clk(gclk));
	jdff dff_A_JjcMM0Nf4_0(.dout(w_dff_A_eYdukx852_0),.din(w_dff_A_JjcMM0Nf4_0),.clk(gclk));
	jdff dff_A_eYdukx852_0(.dout(w_dff_A_ndOpu0aO1_0),.din(w_dff_A_eYdukx852_0),.clk(gclk));
	jdff dff_A_ndOpu0aO1_0(.dout(w_dff_A_uABBfnFD9_0),.din(w_dff_A_ndOpu0aO1_0),.clk(gclk));
	jdff dff_A_uABBfnFD9_0(.dout(w_dff_A_qKXRGcob8_0),.din(w_dff_A_uABBfnFD9_0),.clk(gclk));
	jdff dff_A_qKXRGcob8_0(.dout(w_dff_A_zdN3M1Yr4_0),.din(w_dff_A_qKXRGcob8_0),.clk(gclk));
	jdff dff_A_zdN3M1Yr4_0(.dout(w_dff_A_zGn1J7RA6_0),.din(w_dff_A_zdN3M1Yr4_0),.clk(gclk));
	jdff dff_A_zGn1J7RA6_0(.dout(w_dff_A_UfIpb2WJ6_0),.din(w_dff_A_zGn1J7RA6_0),.clk(gclk));
	jdff dff_A_UfIpb2WJ6_0(.dout(w_dff_A_iGMr5L8y5_0),.din(w_dff_A_UfIpb2WJ6_0),.clk(gclk));
	jdff dff_A_iGMr5L8y5_0(.dout(w_dff_A_Q8mnEBbA1_0),.din(w_dff_A_iGMr5L8y5_0),.clk(gclk));
	jdff dff_A_Q8mnEBbA1_0(.dout(w_dff_A_Ud3K8bkm7_0),.din(w_dff_A_Q8mnEBbA1_0),.clk(gclk));
	jdff dff_A_Ud3K8bkm7_0(.dout(w_dff_A_62ZBuxpt8_0),.din(w_dff_A_Ud3K8bkm7_0),.clk(gclk));
	jdff dff_A_62ZBuxpt8_0(.dout(w_dff_A_YcS3E57m0_0),.din(w_dff_A_62ZBuxpt8_0),.clk(gclk));
	jdff dff_A_YcS3E57m0_0(.dout(w_dff_A_oSvDBZ9y5_0),.din(w_dff_A_YcS3E57m0_0),.clk(gclk));
	jdff dff_A_oSvDBZ9y5_0(.dout(w_dff_A_jnphPJQq4_0),.din(w_dff_A_oSvDBZ9y5_0),.clk(gclk));
	jdff dff_A_jnphPJQq4_0(.dout(w_dff_A_e9UdxjJX2_0),.din(w_dff_A_jnphPJQq4_0),.clk(gclk));
	jdff dff_A_e9UdxjJX2_0(.dout(w_dff_A_pVghKH8V0_0),.din(w_dff_A_e9UdxjJX2_0),.clk(gclk));
	jdff dff_A_pVghKH8V0_0(.dout(w_dff_A_kyqh7XdT3_0),.din(w_dff_A_pVghKH8V0_0),.clk(gclk));
	jdff dff_A_kyqh7XdT3_0(.dout(w_dff_A_I9c9A40x6_0),.din(w_dff_A_kyqh7XdT3_0),.clk(gclk));
	jdff dff_A_I9c9A40x6_0(.dout(G223gat),.din(w_dff_A_I9c9A40x6_0),.clk(gclk));
	jdff dff_A_HtwnrXEd7_1(.dout(w_dff_A_bnOtvpbk1_0),.din(w_dff_A_HtwnrXEd7_1),.clk(gclk));
	jdff dff_A_bnOtvpbk1_0(.dout(w_dff_A_nKAG9DvF0_0),.din(w_dff_A_bnOtvpbk1_0),.clk(gclk));
	jdff dff_A_nKAG9DvF0_0(.dout(w_dff_A_p6GH5ayH4_0),.din(w_dff_A_nKAG9DvF0_0),.clk(gclk));
	jdff dff_A_p6GH5ayH4_0(.dout(w_dff_A_yTinfqHI7_0),.din(w_dff_A_p6GH5ayH4_0),.clk(gclk));
	jdff dff_A_yTinfqHI7_0(.dout(w_dff_A_PxgQhShx3_0),.din(w_dff_A_yTinfqHI7_0),.clk(gclk));
	jdff dff_A_PxgQhShx3_0(.dout(w_dff_A_Ju0kYDkb4_0),.din(w_dff_A_PxgQhShx3_0),.clk(gclk));
	jdff dff_A_Ju0kYDkb4_0(.dout(w_dff_A_KjOYL2s89_0),.din(w_dff_A_Ju0kYDkb4_0),.clk(gclk));
	jdff dff_A_KjOYL2s89_0(.dout(w_dff_A_FG5twln81_0),.din(w_dff_A_KjOYL2s89_0),.clk(gclk));
	jdff dff_A_FG5twln81_0(.dout(w_dff_A_Q9QrCNcM2_0),.din(w_dff_A_FG5twln81_0),.clk(gclk));
	jdff dff_A_Q9QrCNcM2_0(.dout(w_dff_A_Y8y80gZX3_0),.din(w_dff_A_Q9QrCNcM2_0),.clk(gclk));
	jdff dff_A_Y8y80gZX3_0(.dout(w_dff_A_zUNyRLWq9_0),.din(w_dff_A_Y8y80gZX3_0),.clk(gclk));
	jdff dff_A_zUNyRLWq9_0(.dout(w_dff_A_M4nRc6jE1_0),.din(w_dff_A_zUNyRLWq9_0),.clk(gclk));
	jdff dff_A_M4nRc6jE1_0(.dout(w_dff_A_wVczK4xJ1_0),.din(w_dff_A_M4nRc6jE1_0),.clk(gclk));
	jdff dff_A_wVczK4xJ1_0(.dout(G329gat),.din(w_dff_A_wVczK4xJ1_0),.clk(gclk));
	jdff dff_A_CQ7xasqQ2_2(.dout(w_dff_A_QMiACvvH1_0),.din(w_dff_A_CQ7xasqQ2_2),.clk(gclk));
	jdff dff_A_QMiACvvH1_0(.dout(w_dff_A_MdlvTLdw8_0),.din(w_dff_A_QMiACvvH1_0),.clk(gclk));
	jdff dff_A_MdlvTLdw8_0(.dout(w_dff_A_RM0lo1XM4_0),.din(w_dff_A_MdlvTLdw8_0),.clk(gclk));
	jdff dff_A_RM0lo1XM4_0(.dout(w_dff_A_0hA5HcLW0_0),.din(w_dff_A_RM0lo1XM4_0),.clk(gclk));
	jdff dff_A_0hA5HcLW0_0(.dout(w_dff_A_WRDgAVWl6_0),.din(w_dff_A_0hA5HcLW0_0),.clk(gclk));
	jdff dff_A_WRDgAVWl6_0(.dout(w_dff_A_nTSprNPu2_0),.din(w_dff_A_WRDgAVWl6_0),.clk(gclk));
	jdff dff_A_nTSprNPu2_0(.dout(G370gat),.din(w_dff_A_nTSprNPu2_0),.clk(gclk));
	jdff dff_A_Gk1ONaMb3_1(.dout(w_dff_A_ScGCnjWl0_0),.din(w_dff_A_Gk1ONaMb3_1),.clk(gclk));
	jdff dff_A_ScGCnjWl0_0(.dout(G430gat),.din(w_dff_A_ScGCnjWl0_0),.clk(gclk));
endmodule

