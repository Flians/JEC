/*
rf_c3540:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jdff: 1943
	jand: 535
	jor: 374

Summary:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jdff: 1943
	jand: 535
	jor: 374

The maximum logic level gap of any gate:
	rf_c3540: 26
*/

module rf_c3540(gclk, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402);
	input gclk;
	input G1;
	input G13;
	input G20;
	input G33;
	input G41;
	input G45;
	input G50;
	input G58;
	input G68;
	input G77;
	input G87;
	input G97;
	input G107;
	input G116;
	input G124;
	input G125;
	input G128;
	input G132;
	input G137;
	input G143;
	input G150;
	input G159;
	input G169;
	input G179;
	input G190;
	input G200;
	input G213;
	input G222;
	input G223;
	input G226;
	input G232;
	input G238;
	input G244;
	input G250;
	input G257;
	input G264;
	input G270;
	input G274;
	input G283;
	input G294;
	input G303;
	input G311;
	input G317;
	input G322;
	input G326;
	input G329;
	input G330;
	input G343;
	input G1698;
	input G2897;
	output G353;
	output G355;
	output G361;
	output G358;
	output G351;
	output G372;
	output G369;
	output G399;
	output G364;
	output G396;
	output G384;
	output G367;
	output G387;
	output G393;
	output G390;
	output G378;
	output G375;
	output G381;
	output G407;
	output G409;
	output G405;
	output G402;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [2:0] w_G1_2;
	wire [1:0] w_G1_3;
	wire [2:0] w_G13_0;
	wire [1:0] w_G13_1;
	wire [2:0] w_G20_0;
	wire [2:0] w_G20_1;
	wire [2:0] w_G20_2;
	wire [2:0] w_G20_3;
	wire [2:0] w_G20_4;
	wire [2:0] w_G20_5;
	wire [2:0] w_G20_6;
	wire [1:0] w_G20_7;
	wire [2:0] w_G33_0;
	wire [2:0] w_G33_1;
	wire [2:0] w_G33_2;
	wire [2:0] w_G33_3;
	wire [2:0] w_G33_4;
	wire [2:0] w_G33_5;
	wire [2:0] w_G33_6;
	wire [2:0] w_G33_7;
	wire [2:0] w_G33_8;
	wire [2:0] w_G33_9;
	wire [2:0] w_G33_10;
	wire [2:0] w_G33_11;
	wire [2:0] w_G41_0;
	wire [1:0] w_G41_1;
	wire [2:0] w_G45_0;
	wire [2:0] w_G45_1;
	wire [2:0] w_G50_0;
	wire [2:0] w_G50_1;
	wire [2:0] w_G50_2;
	wire [2:0] w_G50_3;
	wire [2:0] w_G50_4;
	wire [2:0] w_G50_5;
	wire [2:0] w_G58_0;
	wire [2:0] w_G58_1;
	wire [2:0] w_G58_2;
	wire [2:0] w_G58_3;
	wire [2:0] w_G58_4;
	wire [1:0] w_G58_5;
	wire [2:0] w_G68_0;
	wire [2:0] w_G68_1;
	wire [2:0] w_G68_2;
	wire [2:0] w_G68_3;
	wire [2:0] w_G68_4;
	wire [1:0] w_G68_5;
	wire [2:0] w_G77_0;
	wire [2:0] w_G77_1;
	wire [2:0] w_G77_2;
	wire [2:0] w_G77_3;
	wire [2:0] w_G77_4;
	wire [1:0] w_G77_5;
	wire [2:0] w_G87_0;
	wire [2:0] w_G87_1;
	wire [2:0] w_G87_2;
	wire [2:0] w_G87_3;
	wire [2:0] w_G97_0;
	wire [2:0] w_G97_1;
	wire [2:0] w_G97_2;
	wire [2:0] w_G97_3;
	wire [2:0] w_G97_4;
	wire [1:0] w_G97_5;
	wire [2:0] w_G107_0;
	wire [2:0] w_G107_1;
	wire [2:0] w_G107_2;
	wire [2:0] w_G107_3;
	wire [2:0] w_G107_4;
	wire [1:0] w_G107_5;
	wire [2:0] w_G116_0;
	wire [2:0] w_G116_1;
	wire [2:0] w_G116_2;
	wire [2:0] w_G116_3;
	wire [2:0] w_G116_4;
	wire [1:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [2:0] w_G132_0;
	wire [1:0] w_G132_1;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G143_0;
	wire [2:0] w_G143_1;
	wire [1:0] w_G143_2;
	wire [2:0] w_G150_0;
	wire [2:0] w_G150_1;
	wire [2:0] w_G150_2;
	wire [1:0] w_G150_3;
	wire [2:0] w_G159_0;
	wire [2:0] w_G159_1;
	wire [2:0] w_G159_2;
	wire [2:0] w_G159_3;
	wire [2:0] w_G169_0;
	wire [1:0] w_G169_1;
	wire [2:0] w_G179_0;
	wire [2:0] w_G179_1;
	wire [2:0] w_G179_2;
	wire [2:0] w_G190_0;
	wire [2:0] w_G190_1;
	wire [2:0] w_G190_2;
	wire [2:0] w_G190_3;
	wire [1:0] w_G190_4;
	wire [2:0] w_G200_0;
	wire [2:0] w_G200_1;
	wire [2:0] w_G200_2;
	wire [2:0] w_G200_3;
	wire [2:0] w_G200_4;
	wire [2:0] w_G213_0;
	wire [1:0] w_G223_0;
	wire [2:0] w_G226_0;
	wire [1:0] w_G226_1;
	wire [2:0] w_G232_0;
	wire [2:0] w_G232_1;
	wire [2:0] w_G238_0;
	wire [2:0] w_G238_1;
	wire [2:0] w_G244_0;
	wire [2:0] w_G244_1;
	wire [2:0] w_G250_0;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [2:0] w_G264_0;
	wire [1:0] w_G264_1;
	wire [2:0] w_G270_0;
	wire [2:0] w_G274_0;
	wire [2:0] w_G283_0;
	wire [2:0] w_G283_1;
	wire [2:0] w_G283_2;
	wire [2:0] w_G283_3;
	wire [2:0] w_G294_0;
	wire [2:0] w_G294_1;
	wire [2:0] w_G294_2;
	wire [1:0] w_G294_3;
	wire [2:0] w_G303_0;
	wire [2:0] w_G303_1;
	wire [2:0] w_G303_2;
	wire [2:0] w_G311_0;
	wire [2:0] w_G311_1;
	wire [2:0] w_G317_0;
	wire [1:0] w_G317_1;
	wire [2:0] w_G322_0;
	wire [1:0] w_G326_0;
	wire [1:0] w_G330_0;
	wire [1:0] w_G343_0;
	wire [2:0] w_G1698_0;
	wire w_G355_0;
	wire G355_fa_;
	wire [1:0] w_G396_0;
	wire G396_fa_;
	wire w_G384_0;
	wire G384_fa_;
	wire [1:0] w_G387_0;
	wire G387_fa_;
	wire [2:0] w_n72_0;
	wire [1:0] w_n72_1;
	wire [2:0] w_n73_0;
	wire [2:0] w_n73_1;
	wire [2:0] w_n73_2;
	wire [2:0] w_n74_0;
	wire [1:0] w_n74_1;
	wire [2:0] w_n75_0;
	wire [1:0] w_n75_1;
	wire [1:0] w_n76_0;
	wire [1:0] w_n77_0;
	wire [2:0] w_n79_0;
	wire [2:0] w_n80_0;
	wire [1:0] w_n80_1;
	wire [2:0] w_n81_0;
	wire [2:0] w_n85_0;
	wire [1:0] w_n86_0;
	wire [2:0] w_n88_0;
	wire [1:0] w_n88_1;
	wire [2:0] w_n91_0;
	wire [2:0] w_n91_1;
	wire [1:0] w_n93_0;
	wire [2:0] w_n97_0;
	wire [2:0] w_n97_1;
	wire [1:0] w_n97_2;
	wire [2:0] w_n98_0;
	wire [2:0] w_n98_1;
	wire [1:0] w_n98_2;
	wire [2:0] w_n103_0;
	wire [2:0] w_n105_0;
	wire [2:0] w_n105_1;
	wire [1:0] w_n105_2;
	wire [1:0] w_n106_0;
	wire [2:0] w_n112_0;
	wire [2:0] w_n112_1;
	wire [2:0] w_n112_2;
	wire [2:0] w_n112_3;
	wire [2:0] w_n112_4;
	wire [2:0] w_n112_5;
	wire [2:0] w_n113_0;
	wire [2:0] w_n113_1;
	wire [2:0] w_n113_2;
	wire [1:0] w_n113_3;
	wire [2:0] w_n114_0;
	wire [2:0] w_n114_1;
	wire [2:0] w_n115_0;
	wire [1:0] w_n115_1;
	wire [1:0] w_n116_0;
	wire [2:0] w_n118_0;
	wire [2:0] w_n121_0;
	wire [2:0] w_n122_0;
	wire [1:0] w_n122_1;
	wire [2:0] w_n123_0;
	wire [2:0] w_n123_1;
	wire [1:0] w_n131_0;
	wire [1:0] w_n135_0;
	wire [2:0] w_n137_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n144_0;
	wire [2:0] w_n146_0;
	wire [2:0] w_n146_1;
	wire [2:0] w_n146_2;
	wire [2:0] w_n146_3;
	wire [2:0] w_n147_0;
	wire [2:0] w_n148_0;
	wire [2:0] w_n148_1;
	wire [2:0] w_n148_2;
	wire [2:0] w_n148_3;
	wire [2:0] w_n148_4;
	wire [2:0] w_n148_5;
	wire [2:0] w_n148_6;
	wire [2:0] w_n148_7;
	wire [2:0] w_n148_8;
	wire [2:0] w_n148_9;
	wire [2:0] w_n149_0;
	wire [2:0] w_n149_1;
	wire [1:0] w_n149_2;
	wire [2:0] w_n151_0;
	wire [2:0] w_n151_1;
	wire [2:0] w_n151_2;
	wire [2:0] w_n151_3;
	wire [2:0] w_n151_4;
	wire [2:0] w_n152_0;
	wire [2:0] w_n152_1;
	wire [2:0] w_n152_2;
	wire [1:0] w_n152_3;
	wire [1:0] w_n154_0;
	wire [2:0] w_n155_0;
	wire [2:0] w_n155_1;
	wire [2:0] w_n155_2;
	wire [1:0] w_n155_3;
	wire [2:0] w_n157_0;
	wire [2:0] w_n161_0;
	wire [1:0] w_n161_1;
	wire [2:0] w_n162_0;
	wire [1:0] w_n163_0;
	wire [2:0] w_n166_0;
	wire [2:0] w_n166_1;
	wire [2:0] w_n166_2;
	wire [1:0] w_n166_3;
	wire [2:0] w_n170_0;
	wire [1:0] w_n172_0;
	wire [2:0] w_n179_0;
	wire [2:0] w_n179_1;
	wire [1:0] w_n180_0;
	wire [2:0] w_n185_0;
	wire [2:0] w_n185_1;
	wire [2:0] w_n185_2;
	wire [2:0] w_n185_3;
	wire [2:0] w_n189_0;
	wire [2:0] w_n189_1;
	wire [1:0] w_n189_2;
	wire [2:0] w_n190_0;
	wire [2:0] w_n190_1;
	wire [2:0] w_n191_0;
	wire [1:0] w_n195_0;
	wire [2:0] w_n196_0;
	wire [2:0] w_n196_1;
	wire [2:0] w_n196_2;
	wire [2:0] w_n197_0;
	wire [1:0] w_n197_1;
	wire [2:0] w_n199_0;
	wire [1:0] w_n199_1;
	wire [1:0] w_n201_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n206_0;
	wire [2:0] w_n210_0;
	wire [1:0] w_n213_0;
	wire [1:0] w_n214_0;
	wire [1:0] w_n218_0;
	wire [1:0] w_n219_0;
	wire [2:0] w_n221_0;
	wire [1:0] w_n228_0;
	wire [2:0] w_n229_0;
	wire [1:0] w_n230_0;
	wire [2:0] w_n231_0;
	wire [2:0] w_n234_0;
	wire [1:0] w_n241_0;
	wire [2:0] w_n242_0;
	wire [2:0] w_n243_0;
	wire [2:0] w_n246_0;
	wire [1:0] w_n246_1;
	wire [1:0] w_n249_0;
	wire [1:0] w_n255_0;
	wire [1:0] w_n257_0;
	wire [1:0] w_n259_0;
	wire [1:0] w_n261_0;
	wire [1:0] w_n262_0;
	wire [2:0] w_n269_0;
	wire [2:0] w_n269_1;
	wire [1:0] w_n270_0;
	wire [2:0] w_n271_0;
	wire [2:0] w_n271_1;
	wire [2:0] w_n274_0;
	wire [1:0] w_n278_0;
	wire [1:0] w_n279_0;
	wire [1:0] w_n281_0;
	wire [2:0] w_n288_0;
	wire [1:0] w_n288_1;
	wire [1:0] w_n296_0;
	wire [1:0] w_n298_0;
	wire [1:0] w_n300_0;
	wire [1:0] w_n303_0;
	wire [2:0] w_n312_0;
	wire [1:0] w_n312_1;
	wire [1:0] w_n315_0;
	wire [1:0] w_n320_0;
	wire [1:0] w_n324_0;
	wire [1:0] w_n328_0;
	wire [1:0] w_n334_0;
	wire [1:0] w_n339_0;
	wire [2:0] w_n346_0;
	wire [1:0] w_n346_1;
	wire [2:0] w_n355_0;
	wire [1:0] w_n355_1;
	wire [1:0] w_n362_0;
	wire [2:0] w_n367_0;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n374_0;
	wire [1:0] w_n381_0;
	wire [2:0] w_n382_0;
	wire [1:0] w_n382_1;
	wire [2:0] w_n385_0;
	wire [1:0] w_n385_1;
	wire [2:0] w_n387_0;
	wire [1:0] w_n387_1;
	wire [1:0] w_n390_0;
	wire [2:0] w_n401_0;
	wire [2:0] w_n404_0;
	wire [1:0] w_n405_0;
	wire [2:0] w_n407_0;
	wire [2:0] w_n407_1;
	wire [1:0] w_n407_2;
	wire [1:0] w_n412_0;
	wire [2:0] w_n420_0;
	wire [1:0] w_n420_1;
	wire [2:0] w_n425_0;
	wire [2:0] w_n425_1;
	wire [1:0] w_n426_0;
	wire [1:0] w_n430_0;
	wire [2:0] w_n436_0;
	wire [2:0] w_n439_0;
	wire [1:0] w_n439_1;
	wire [1:0] w_n445_0;
	wire [1:0] w_n446_0;
	wire [2:0] w_n455_0;
	wire [2:0] w_n462_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n474_0;
	wire [1:0] w_n475_0;
	wire [1:0] w_n478_0;
	wire [1:0] w_n479_0;
	wire [1:0] w_n483_0;
	wire [1:0] w_n484_0;
	wire [2:0] w_n492_0;
	wire [1:0] w_n507_0;
	wire [1:0] w_n508_0;
	wire [1:0] w_n511_0;
	wire [1:0] w_n512_0;
	wire [1:0] w_n516_0;
	wire [1:0] w_n517_0;
	wire [2:0] w_n519_0;
	wire [2:0] w_n519_1;
	wire [1:0] w_n523_0;
	wire [1:0] w_n524_0;
	wire [1:0] w_n528_0;
	wire [1:0] w_n532_0;
	wire [1:0] w_n534_0;
	wire [2:0] w_n536_0;
	wire [1:0] w_n539_0;
	wire [1:0] w_n541_0;
	wire [2:0] w_n542_0;
	wire [1:0] w_n543_0;
	wire [2:0] w_n548_0;
	wire [1:0] w_n550_0;
	wire [2:0] w_n552_0;
	wire [1:0] w_n552_1;
	wire [2:0] w_n553_0;
	wire [2:0] w_n553_1;
	wire [2:0] w_n553_2;
	wire [2:0] w_n554_0;
	wire [2:0] w_n554_1;
	wire [2:0] w_n554_2;
	wire [2:0] w_n554_3;
	wire [1:0] w_n556_0;
	wire [1:0] w_n557_0;
	wire [2:0] w_n561_0;
	wire [2:0] w_n563_0;
	wire [1:0] w_n564_0;
	wire [1:0] w_n565_0;
	wire [1:0] w_n567_0;
	wire [2:0] w_n571_0;
	wire [2:0] w_n572_0;
	wire [2:0] w_n573_0;
	wire [2:0] w_n576_0;
	wire [1:0] w_n576_1;
	wire [2:0] w_n588_0;
	wire [1:0] w_n588_1;
	wire [2:0] w_n589_0;
	wire [2:0] w_n589_1;
	wire [2:0] w_n591_0;
	wire [1:0] w_n591_1;
	wire [2:0] w_n592_0;
	wire [2:0] w_n592_1;
	wire [1:0] w_n592_2;
	wire [2:0] w_n593_0;
	wire [1:0] w_n602_0;
	wire [2:0] w_n603_0;
	wire [2:0] w_n603_1;
	wire [1:0] w_n603_2;
	wire [2:0] w_n604_0;
	wire [2:0] w_n604_1;
	wire [1:0] w_n604_2;
	wire [2:0] w_n605_0;
	wire [2:0] w_n605_1;
	wire [2:0] w_n608_0;
	wire [2:0] w_n608_1;
	wire [2:0] w_n612_0;
	wire [2:0] w_n612_1;
	wire [2:0] w_n612_2;
	wire [2:0] w_n612_3;
	wire [1:0] w_n612_4;
	wire [2:0] w_n613_0;
	wire [1:0] w_n613_1;
	wire [1:0] w_n615_0;
	wire [1:0] w_n616_0;
	wire [2:0] w_n617_0;
	wire [2:0] w_n617_1;
	wire [2:0] w_n617_2;
	wire [2:0] w_n617_3;
	wire [2:0] w_n617_4;
	wire [2:0] w_n617_5;
	wire [1:0] w_n617_6;
	wire [1:0] w_n619_0;
	wire [1:0] w_n622_0;
	wire [2:0] w_n623_0;
	wire [2:0] w_n623_1;
	wire [2:0] w_n623_2;
	wire [2:0] w_n623_3;
	wire [2:0] w_n623_4;
	wire [1:0] w_n623_5;
	wire [1:0] w_n626_0;
	wire [2:0] w_n627_0;
	wire [2:0] w_n627_1;
	wire [2:0] w_n627_2;
	wire [2:0] w_n627_3;
	wire [2:0] w_n627_4;
	wire [2:0] w_n627_5;
	wire [2:0] w_n627_6;
	wire [1:0] w_n627_7;
	wire [2:0] w_n631_0;
	wire [2:0] w_n631_1;
	wire [2:0] w_n631_2;
	wire [2:0] w_n631_3;
	wire [2:0] w_n631_4;
	wire [2:0] w_n631_5;
	wire [2:0] w_n631_6;
	wire [1:0] w_n631_7;
	wire [2:0] w_n634_0;
	wire [2:0] w_n634_1;
	wire [2:0] w_n634_2;
	wire [2:0] w_n634_3;
	wire [1:0] w_n634_4;
	wire [2:0] w_n636_0;
	wire [2:0] w_n636_1;
	wire [2:0] w_n636_2;
	wire [2:0] w_n636_3;
	wire [2:0] w_n636_4;
	wire [2:0] w_n636_5;
	wire [2:0] w_n636_6;
	wire [1:0] w_n636_7;
	wire [1:0] w_n639_0;
	wire [2:0] w_n640_0;
	wire [2:0] w_n640_1;
	wire [2:0] w_n640_2;
	wire [2:0] w_n640_3;
	wire [2:0] w_n640_4;
	wire [2:0] w_n640_5;
	wire [2:0] w_n640_6;
	wire [1:0] w_n640_7;
	wire [2:0] w_n642_0;
	wire [2:0] w_n642_1;
	wire [2:0] w_n642_2;
	wire [2:0] w_n642_3;
	wire [2:0] w_n642_4;
	wire [2:0] w_n642_5;
	wire [2:0] w_n642_6;
	wire [1:0] w_n642_7;
	wire [1:0] w_n654_0;
	wire [1:0] w_n657_0;
	wire [1:0] w_n661_0;
	wire [2:0] w_n672_0;
	wire [1:0] w_n672_1;
	wire [2:0] w_n675_0;
	wire [1:0] w_n676_0;
	wire [1:0] w_n680_0;
	wire [1:0] w_n692_0;
	wire [2:0] w_n696_0;
	wire [2:0] w_n696_1;
	wire [1:0] w_n717_0;
	wire [1:0] w_n728_0;
	wire [2:0] w_n743_0;
	wire [1:0] w_n743_1;
	wire [1:0] w_n750_0;
	wire [1:0] w_n754_0;
	wire [2:0] w_n758_0;
	wire [1:0] w_n758_1;
	wire [1:0] w_n759_0;
	wire [1:0] w_n760_0;
	wire [2:0] w_n764_0;
	wire [2:0] w_n764_1;
	wire [1:0] w_n769_0;
	wire [2:0] w_n771_0;
	wire [1:0] w_n779_0;
	wire [1:0] w_n797_0;
	wire [1:0] w_n801_0;
	wire [1:0] w_n816_0;
	wire [1:0] w_n823_0;
	wire [1:0] w_n825_0;
	wire [2:0] w_n853_0;
	wire [2:0] w_n855_0;
	wire [2:0] w_n861_0;
	wire [1:0] w_n861_1;
	wire [1:0] w_n863_0;
	wire [1:0] w_n864_0;
	wire [1:0] w_n899_0;
	wire [1:0] w_n909_0;
	wire [2:0] w_n937_0;
	wire [1:0] w_n940_0;
	wire [1:0] w_n962_0;
	wire [2:0] w_n988_0;
	wire [1:0] w_n990_0;
	wire [2:0] w_n991_0;
	wire [1:0] w_n992_0;
	wire [2:0] w_n994_0;
	wire [2:0] w_n996_0;
	wire [1:0] w_n999_0;
	wire [2:0] w_n1001_0;
	wire [2:0] w_n1002_0;
	wire [1:0] w_n1003_0;
	wire [2:0] w_n1049_0;
	wire [1:0] w_n1052_0;
	wire [1:0] w_n1057_0;
	wire [1:0] w_n1059_0;
	wire [1:0] w_n1088_0;
	wire [2:0] w_n1114_0;
	wire [2:0] w_n1162_0;
	wire [1:0] w_n1164_0;
	wire [1:0] w_n1172_0;
	wire [1:0] w_n1175_0;
	wire [1:0] w_n1183_0;
	wire [1:0] w_n1184_0;
	wire [1:0] w_n1187_0;
	wire w_dff_B_ZbIvEJMZ1_1;
	wire w_dff_B_RKYEFx1F2_0;
	wire w_dff_B_XAQHaUNc9_0;
	wire w_dff_A_35iZO2qL7_1;
	wire w_dff_A_vGw5cjWo7_1;
	wire w_dff_A_QFqMBReo8_0;
	wire w_dff_B_TiI7vb9P6_1;
	wire w_dff_B_57HSYb0W9_0;
	wire w_dff_B_gqmF82y40_0;
	wire w_dff_B_FqyPStGC8_0;
	wire w_dff_B_bR07qUFD3_0;
	wire w_dff_B_fekINiU85_0;
	wire w_dff_B_FfPOBCUt9_0;
	wire w_dff_B_Txu07bCc5_0;
	wire w_dff_B_oyBfdrSg1_0;
	wire w_dff_B_pnhV1Ahu7_0;
	wire w_dff_B_aW8cQsyk1_0;
	wire w_dff_B_30hQyZDl3_0;
	wire w_dff_B_z4aZpyvY0_0;
	wire w_dff_B_r7GeDUeT2_0;
	wire w_dff_B_eRMJhjTK0_0;
	wire w_dff_B_zRFfzQZT1_0;
	wire w_dff_B_GrKdLDr06_0;
	wire w_dff_B_wUJghsZH9_0;
	wire w_dff_B_KIZG7nLE8_0;
	wire w_dff_B_F9VlwxNV5_0;
	wire w_dff_B_0prqLHRs9_0;
	wire w_dff_B_3vzv6ll53_0;
	wire w_dff_B_1o8dJWyL5_0;
	wire w_dff_B_iS3n88y91_0;
	wire w_dff_B_gRaPGDVy3_0;
	wire w_dff_B_3ciAPUTD0_0;
	wire w_dff_B_abRt2R1v3_0;
	wire w_dff_B_7uld260A0_0;
	wire w_dff_B_iHgZDsFN1_0;
	wire w_dff_B_S17TyMTG2_1;
	wire w_dff_B_ucJF10Ej6_0;
	wire w_dff_B_oaMhJkbn7_0;
	wire w_dff_B_bgnk8CN45_0;
	wire w_dff_B_DiO322YL7_0;
	wire w_dff_B_QSAAz7sD6_0;
	wire w_dff_B_2phjyk4W1_0;
	wire w_dff_B_HKKGKKBb7_0;
	wire w_dff_B_slILIBFh7_0;
	wire w_dff_B_GnEZZa5h6_0;
	wire w_dff_B_2XRZcm3V8_0;
	wire w_dff_B_EFk3Y9Tt1_0;
	wire w_dff_B_zseAXeDE6_0;
	wire w_dff_B_9IuZgE8F7_0;
	wire w_dff_B_MpSWbReq4_0;
	wire w_dff_B_alibiwfi3_0;
	wire w_dff_B_L8rAT8m70_0;
	wire w_dff_B_39uXXub01_0;
	wire w_dff_B_bLDCNedl5_0;
	wire w_dff_B_Q1LIwqe58_0;
	wire w_dff_A_pq1kqkUf9_1;
	wire w_dff_A_76i7BKoX5_1;
	wire w_dff_B_INXKO3Aj0_0;
	wire w_dff_A_3ErFUkCU3_0;
	wire w_dff_B_ismogaiY2_1;
	wire w_dff_A_Tqa4XRTQ6_0;
	wire w_dff_B_1lyPjolQ8_1;
	wire w_dff_B_STSgn9S99_1;
	wire w_dff_B_ksuYp0Ct0_1;
	wire w_dff_B_cUnlXmVH2_1;
	wire w_dff_B_7xWKsNru0_1;
	wire w_dff_B_OLwqOrq20_1;
	wire w_dff_B_j5kNHohR6_1;
	wire w_dff_B_av9rlSH53_1;
	wire w_dff_B_CQ4RFwI08_1;
	wire w_dff_B_EP064UMY9_1;
	wire w_dff_B_6wGLHJU34_1;
	wire w_dff_B_vckcHnIO7_1;
	wire w_dff_B_FYYw2jGJ6_1;
	wire w_dff_B_bIzB3b574_1;
	wire w_dff_B_GYgaBrU91_1;
	wire w_dff_B_m8yHHaLW0_1;
	wire w_dff_B_9dBhZNRm2_1;
	wire w_dff_B_ABL8aGuQ4_1;
	wire w_dff_B_oD7sEuKY4_1;
	wire w_dff_B_0cGMx41z6_1;
	wire w_dff_B_e8nhOBiv9_1;
	wire w_dff_B_7lWRFK0D9_1;
	wire w_dff_B_M7PXAHRb5_1;
	wire w_dff_B_PtNcMZnx7_1;
	wire w_dff_B_fVe4i1GS5_1;
	wire w_dff_B_Dkas4rHc5_1;
	wire w_dff_A_1gHWTp1M2_0;
	wire w_dff_B_d1iaAPKo4_1;
	wire w_dff_B_F6HiktET4_1;
	wire w_dff_B_Itre6EaQ7_1;
	wire w_dff_B_WPTFmLO94_1;
	wire w_dff_B_0KnA5P1y8_1;
	wire w_dff_B_qKV9czAu7_1;
	wire w_dff_B_S7POIotw4_1;
	wire w_dff_B_KGURSiXD8_1;
	wire w_dff_B_71sAdNul4_1;
	wire w_dff_B_oMD68yai7_1;
	wire w_dff_B_ow1ivQgc4_1;
	wire w_dff_B_Yw4TcDea7_1;
	wire w_dff_B_xRYm96vM2_1;
	wire w_dff_B_eUB6iv2E4_1;
	wire w_dff_B_cEsRtduB3_1;
	wire w_dff_B_8nXiF0Vw6_1;
	wire w_dff_B_srSpfLWX5_1;
	wire w_dff_B_aaCjEMMh1_1;
	wire w_dff_B_3XkVdb4L2_1;
	wire w_dff_B_haZlQY2K5_1;
	wire w_dff_B_eHtJxHqZ6_1;
	wire w_dff_B_atyYGVVP2_1;
	wire w_dff_B_GBCDlgHM7_1;
	wire w_dff_B_PNjCKbEy0_1;
	wire w_dff_B_nNzt09gq4_1;
	wire w_dff_B_nr9EUWKf8_1;
	wire w_dff_B_HoUtMLY20_1;
	wire w_dff_B_Tn5Dfvsh7_1;
	wire w_dff_A_FkrEWMOn2_0;
	wire w_dff_A_i13Nxk1d4_0;
	wire w_dff_A_wMshBjsY8_0;
	wire w_dff_A_elJ3kVjw5_0;
	wire w_dff_A_LXcfYMdX0_0;
	wire w_dff_A_0OlSHuzH1_0;
	wire w_dff_A_8XzyIIqw3_0;
	wire w_dff_A_7aIAM5uW5_0;
	wire w_dff_A_JX7QnrZu6_0;
	wire w_dff_A_YYX4gCcC9_0;
	wire w_dff_A_ezIhfjT26_0;
	wire w_dff_A_EinBL5jg3_0;
	wire w_dff_A_fWezhZQK1_0;
	wire w_dff_A_pyHyVM520_0;
	wire w_dff_A_uTB02lxm3_0;
	wire w_dff_A_Czfwup3U9_0;
	wire w_dff_A_s2qmCIG71_0;
	wire w_dff_A_fLRtkNEI5_0;
	wire w_dff_A_QiWqXZtD8_0;
	wire w_dff_A_hlIfiqL39_0;
	wire w_dff_A_wZ6b6fHU0_0;
	wire w_dff_A_0WDg3HZv0_0;
	wire w_dff_A_ED2r026o9_0;
	wire w_dff_A_2gFj4f353_0;
	wire w_dff_A_CUINI1G20_1;
	wire w_dff_A_qG5g4Kdt6_1;
	wire w_dff_A_VKYtCPlx4_1;
	wire w_dff_A_KWqK4jsg9_1;
	wire w_dff_A_fSoq5eSk9_1;
	wire w_dff_A_2RZGnjge1_1;
	wire w_dff_A_jlR3c4od4_1;
	wire w_dff_A_YbRQWkiM0_1;
	wire w_dff_A_LpgbsOwJ3_1;
	wire w_dff_A_HkHWyVHQ7_1;
	wire w_dff_A_bPrk78ai6_1;
	wire w_dff_A_RwyT5Put4_1;
	wire w_dff_A_BSkzwkY28_1;
	wire w_dff_A_GYfWShQb6_1;
	wire w_dff_A_9sO4ZTmB4_1;
	wire w_dff_A_EAUOJHMP3_1;
	wire w_dff_A_hjlqjJGa8_1;
	wire w_dff_A_WW1YB6Nx9_1;
	wire w_dff_A_6kQ4PVCa9_1;
	wire w_dff_A_UnE89SV35_1;
	wire w_dff_A_TwVIFBZk6_1;
	wire w_dff_A_BVhJRhXi2_1;
	wire w_dff_A_2P7m60Fo7_1;
	wire w_dff_A_TkG7pfVH7_1;
	wire w_dff_A_PBO6IMgf3_1;
	wire w_dff_A_75qdFNfU4_0;
	wire w_dff_B_DVFnj4U50_1;
	wire w_dff_B_kjZczfGZ9_0;
	wire w_dff_B_z9x0sSSx3_0;
	wire w_dff_B_mueMJx3S2_0;
	wire w_dff_B_krCILoBk6_0;
	wire w_dff_B_7VYOSbKx5_0;
	wire w_dff_B_H8cVUlWX9_0;
	wire w_dff_B_KyoqtR4A7_0;
	wire w_dff_B_92gJze930_0;
	wire w_dff_B_8BSMLYpj6_0;
	wire w_dff_B_9ILQ2W4v2_0;
	wire w_dff_B_S2QAhHBW2_0;
	wire w_dff_B_uRmScwGU2_0;
	wire w_dff_B_fS9LehUH7_0;
	wire w_dff_B_wBzgC1T75_0;
	wire w_dff_B_ROu9VDUx5_0;
	wire w_dff_B_2cDIwnZe2_1;
	wire w_dff_B_oF2J7WMc8_1;
	wire w_dff_B_SsjTCZ8P9_1;
	wire w_dff_B_bhAskbXh4_1;
	wire w_dff_B_BtmoNtxU2_1;
	wire w_dff_B_x9p7lb4a7_1;
	wire w_dff_B_IP1rCXvj1_1;
	wire w_dff_B_PeH7jio82_1;
	wire w_dff_B_VB52pyBY9_1;
	wire w_dff_B_qrhrT4zO7_0;
	wire w_dff_B_MQBvZFPF6_0;
	wire w_dff_B_LIftqJ252_0;
	wire w_dff_B_71J1ASuV1_0;
	wire w_dff_B_wH6kjyXK3_0;
	wire w_dff_B_snN3B2LV6_0;
	wire w_dff_B_LYXjIAr02_0;
	wire w_dff_B_7iHYmG9Z8_0;
	wire w_dff_B_l64JFMp40_1;
	wire w_dff_B_gLKpy3Be3_1;
	wire w_dff_B_NepKsP0S7_1;
	wire w_dff_B_hNlRGnM00_0;
	wire w_dff_B_W0sNcPpq6_0;
	wire w_dff_B_j0Bgs2dV7_0;
	wire w_dff_B_5S8Al6CO4_0;
	wire w_dff_B_NtJjTnVt0_1;
	wire w_dff_B_YsUganJu0_1;
	wire w_dff_B_HVAqcWer1_0;
	wire w_dff_B_TFXDdaWy7_1;
	wire w_dff_B_SFjiaPKT8_1;
	wire w_dff_B_ggGMsJUX2_1;
	wire w_dff_B_eJtHe2Jq2_1;
	wire w_dff_B_10xCu5ic8_1;
	wire w_dff_B_9YDK52XL0_1;
	wire w_dff_B_vnVczlSn4_1;
	wire w_dff_B_EG6ARHJv1_1;
	wire w_dff_B_dYravbQS3_0;
	wire w_dff_B_7XdmRs1Y7_0;
	wire w_dff_B_AVUazYlt7_0;
	wire w_dff_B_dtJPXaif5_0;
	wire w_dff_B_9uif3c2I5_1;
	wire w_dff_B_qMUJgFx84_1;
	wire w_dff_B_MqphnD900_1;
	wire w_dff_B_XlWbM8QL0_1;
	wire w_dff_B_d1NIOL8X8_1;
	wire w_dff_A_RZtshrj92_1;
	wire w_dff_A_Xxqvm21W1_1;
	wire w_dff_A_j760mmVa3_1;
	wire w_dff_A_6aGBmUHX2_1;
	wire w_dff_A_gRcrxL502_1;
	wire w_dff_A_qQrMKb5R0_0;
	wire w_dff_B_1vL66lyp4_1;
	wire w_dff_B_C7ktbf3h3_1;
	wire w_dff_B_cRQJmgxW2_1;
	wire w_dff_B_66AscVry2_1;
	wire w_dff_B_tqzWkzFC0_1;
	wire w_dff_B_vGoV2cZb0_1;
	wire w_dff_A_5Tgp0F3a0_1;
	wire w_dff_A_kExtFxnH9_1;
	wire w_dff_A_XQEGH7Fg5_1;
	wire w_dff_B_tAnG3rFH9_0;
	wire w_dff_B_ROk0rJVR8_0;
	wire w_dff_B_sGAdXcQK9_0;
	wire w_dff_B_u9jzawup9_0;
	wire w_dff_B_ttQFE8Zp5_0;
	wire w_dff_B_OFsKvyEN6_0;
	wire w_dff_B_lsqKqCwg4_0;
	wire w_dff_B_Au4qUoU05_0;
	wire w_dff_A_WJXeNyEx8_0;
	wire w_dff_A_pbWzgCyS4_0;
	wire w_dff_A_pSs0Kn2T5_1;
	wire w_dff_A_qpemC9y70_1;
	wire w_dff_B_SWbG8yOW4_0;
	wire w_dff_B_Nrqi0ynE4_0;
	wire w_dff_B_tjgyHJ106_0;
	wire w_dff_B_DjOAi9Nd9_0;
	wire w_dff_B_QcnaCo5a3_0;
	wire w_dff_B_eAU6ZNs84_0;
	wire w_dff_B_VwXBFnol2_0;
	wire w_dff_B_2ViURvvM0_0;
	wire w_dff_B_v7qJ2qFU7_0;
	wire w_dff_B_l6gt4ru40_0;
	wire w_dff_B_LwLodLqI6_0;
	wire w_dff_B_Af0sdr0X2_1;
	wire w_dff_B_vXFnbtG86_1;
	wire w_dff_B_TQP1YUm59_1;
	wire w_dff_B_RP8VEQR27_1;
	wire w_dff_B_86zZpgHb2_1;
	wire w_dff_B_M3Zz5C7m8_0;
	wire w_dff_B_RFjhdhla7_1;
	wire w_dff_B_yGPfwFgA3_1;
	wire w_dff_B_wFxVZoM59_1;
	wire w_dff_B_0MkERJX76_1;
	wire w_dff_B_fUpwtMpE7_1;
	wire w_dff_B_UOaAKzrk5_0;
	wire w_dff_A_xsEWv84P2_1;
	wire w_dff_B_HHCElp5e4_2;
	wire w_dff_B_G86RNpOp3_2;
	wire w_dff_B_p5Pr9xfC7_2;
	wire w_dff_A_slKm5Ewo6_1;
	wire w_dff_A_7FpSlnU95_1;
	wire w_dff_A_wMvQFKzl8_0;
	wire w_dff_A_hOWFdUb55_1;
	wire w_dff_A_MmctwkeV4_1;
	wire w_dff_A_qmBZvkLz6_1;
	wire w_dff_A_7ay8bsDi0_0;
	wire w_dff_B_BXD6qlQV4_0;
	wire w_dff_B_WgF3nB0b5_0;
	wire w_dff_B_gPf7eztG3_0;
	wire w_dff_B_YDYslqhf5_0;
	wire w_dff_A_pnr9ZWDy8_2;
	wire w_dff_A_FQjyNBXB6_2;
	wire w_dff_A_mU4FV3g02_1;
	wire w_dff_B_3exNftqn2_1;
	wire w_dff_B_mMffx1gt7_1;
	wire w_dff_B_sSNfvP074_1;
	wire w_dff_B_V1j9SyVP8_1;
	wire w_dff_B_nePEl5Xx0_1;
	wire w_dff_A_Cy2pFh2x2_0;
	wire w_dff_A_fyeVzkVI3_0;
	wire w_dff_A_O5BkJj945_1;
	wire w_dff_B_Cx17UkaA4_0;
	wire w_dff_B_fRdCpgyv1_0;
	wire w_dff_B_c6pRVtlX6_0;
	wire w_dff_B_2JuQXva06_0;
	wire w_dff_B_n3TuTuIJ8_0;
	wire w_dff_B_aNkwzhXz0_0;
	wire w_dff_B_M8nSWbet7_0;
	wire w_dff_B_rDa61NF65_0;
	wire w_dff_B_0avh9kPH0_1;
	wire w_dff_B_XvEe2tqO0_1;
	wire w_dff_B_Lb7neYNf5_0;
	wire w_dff_A_jQ6iCYFb7_2;
	wire w_dff_B_C5qcIsB09_2;
	wire w_dff_B_MvjVfA9W0_1;
	wire w_dff_B_ywj6lkni5_1;
	wire w_dff_B_whVeXqgD6_1;
	wire w_dff_B_WnjYk9sv3_1;
	wire w_dff_B_q2pNGgEz9_0;
	wire w_dff_A_PQFRbtVo2_0;
	wire w_dff_A_qQppqKnn2_2;
	wire w_dff_A_hfLMMskf5_1;
	wire w_dff_A_WWK0B2oo7_1;
	wire w_dff_A_FEpwPMUa3_1;
	wire w_dff_A_sVwYQHnY4_1;
	wire w_dff_A_mp6aKalC4_2;
	wire w_dff_A_gdXVBH7B5_2;
	wire w_dff_A_acilBIRd4_2;
	wire w_dff_A_yjpnAqiE4_2;
	wire w_dff_B_QnFifl5M3_0;
	wire w_dff_A_snOCCsqR1_1;
	wire w_dff_B_HzyL4HYi9_1;
	wire w_dff_B_OhcYGMIq1_1;
	wire w_dff_B_ByV9zlj97_1;
	wire w_dff_B_VJfuxWIR1_0;
	wire w_dff_B_AOeF9rv66_1;
	wire w_dff_B_8j7u9TlS3_0;
	wire w_dff_A_lgUsyUaz7_0;
	wire w_dff_A_Qfqo2AYs7_0;
	wire w_dff_A_P4ZigKiT8_0;
	wire w_dff_B_FStJrMIY0_1;
	wire w_dff_B_NmMHFuky2_1;
	wire w_dff_B_sHP7iWLK0_1;
	wire w_dff_B_Un1tSFFn9_1;
	wire w_dff_B_sdMd6HLu4_1;
	wire w_dff_B_eRk8zz767_1;
	wire w_dff_B_YYMkNhYA5_0;
	wire w_dff_B_roZoaxUK5_0;
	wire w_dff_B_6Fz6g5cU3_1;
	wire w_dff_B_xvuZQWgj8_1;
	wire w_dff_B_9rSm278z7_1;
	wire w_dff_B_Iti47Lbc7_1;
	wire w_dff_B_84D6kbgx2_1;
	wire w_dff_B_8swdFZdK9_1;
	wire w_dff_A_dgcepEnl3_1;
	wire w_dff_A_RyHrEmPo5_1;
	wire w_dff_A_rwQYYhjr9_2;
	wire w_dff_A_R0rFJcId8_2;
	wire w_dff_B_2jr7qtF45_0;
	wire w_dff_B_ZbbISUN88_0;
	wire w_dff_B_Sq1nVs155_0;
	wire w_dff_B_WuxO66pk5_0;
	wire w_dff_A_vBAbKGaa3_1;
	wire w_dff_A_phdcRowx4_1;
	wire w_dff_A_6IF8HUCr3_2;
	wire w_dff_A_qh0ueVTK0_2;
	wire w_dff_B_OEX3IkGW5_1;
	wire w_dff_B_O1xqApWe3_1;
	wire w_dff_B_76bfDyqF7_1;
	wire w_dff_B_mxVotttX4_0;
	wire w_dff_B_vakdpU0h4_0;
	wire w_dff_B_waiU3iPW9_0;
	wire w_dff_B_8GtkNEO43_0;
	wire w_dff_B_0dxtSe3b5_0;
	wire w_dff_B_XK9Rr1Md4_0;
	wire w_dff_B_HGegVXfg3_1;
	wire w_dff_B_EkAG2G5A5_1;
	wire w_dff_B_cNBDWlkf7_0;
	wire w_dff_A_6vLKW1ti3_0;
	wire w_dff_B_dBwvH5b50_1;
	wire w_dff_B_ZsphsNXi2_1;
	wire w_dff_B_9EpyEEZg7_1;
	wire w_dff_B_tafiDLO83_1;
	wire w_dff_B_E9q2u0Q57_1;
	wire w_dff_B_l1n21D5a6_1;
	wire w_dff_B_KfVTBMJA0_1;
	wire w_dff_B_GOaq4DFZ9_1;
	wire w_dff_B_Xkqgtt0R2_1;
	wire w_dff_B_qpC0aZAa8_1;
	wire w_dff_B_kG1WRgHS8_1;
	wire w_dff_B_TTOk1bak3_1;
	wire w_dff_B_LAJJ92v23_1;
	wire w_dff_B_liQ1UMAM7_1;
	wire w_dff_B_5f1pzdeI0_0;
	wire w_dff_A_bwpleDz36_2;
	wire w_dff_A_TdwTkyIG6_0;
	wire w_dff_A_eYQCiEqf0_0;
	wire w_dff_A_LTfKkiCi8_0;
	wire w_dff_A_4UiU7fNk1_0;
	wire w_dff_B_N4HDd12h4_0;
	wire w_dff_B_O0aVY1Bz7_0;
	wire w_dff_A_JPVkXb1c2_0;
	wire w_dff_B_SiD7b9u99_0;
	wire w_dff_B_afRYyTAp2_0;
	wire w_dff_B_VXjngd2T1_0;
	wire w_dff_B_ZNbBFqDO1_0;
	wire w_dff_B_Nw4q9f9k2_0;
	wire w_dff_B_lUDGU5Tm8_1;
	wire w_dff_B_l03SnlX31_1;
	wire w_dff_B_qd4Dr2xX7_1;
	wire w_dff_B_YfOZGs5a8_1;
	wire w_dff_B_1EorlipC6_1;
	wire w_dff_A_6VDFVZtn3_1;
	wire w_dff_A_Eux4reDN6_1;
	wire w_dff_B_hpJU5pAe0_1;
	wire w_dff_B_y8ZMZmyl1_1;
	wire w_dff_B_dTs5iTOn6_1;
	wire w_dff_B_40pmEBcG8_1;
	wire w_dff_B_ywfEaQGJ9_1;
	wire w_dff_A_Atnr6eaZ2_0;
	wire w_dff_A_u6lMMEG02_1;
	wire w_dff_A_JEUNizrH2_1;
	wire w_dff_A_uiOC0J294_1;
	wire w_dff_A_f2WoVYay3_2;
	wire w_dff_A_4ndtRwkk5_2;
	wire w_dff_A_YzKwCjno0_2;
	wire w_dff_A_6KVDIPDC3_2;
	wire w_dff_A_UaieZtxF1_1;
	wire w_dff_B_fkrlfE7F9_0;
	wire w_dff_A_rBK6NEAD6_0;
	wire w_dff_A_n8CIkRW42_0;
	wire w_dff_A_05j5Fhvw0_2;
	wire w_dff_A_JtTPq6K41_2;
	wire w_dff_B_s3dYIOLe0_1;
	wire w_dff_B_t8HqBvIk0_1;
	wire w_dff_B_ijOsRv3d3_0;
	wire w_dff_B_oAB1G1BA4_0;
	wire w_dff_A_nFcxiCu25_1;
	wire w_dff_A_Ig1MTnX10_2;
	wire w_dff_B_C8F25GoX1_1;
	wire w_dff_B_ArWb2Guz8_0;
	wire w_dff_A_KSVncrO02_0;
	wire w_dff_A_cOYiOvKk8_1;
	wire w_dff_A_XSZpSyWq1_1;
	wire w_dff_B_GWUvgwss7_1;
	wire w_dff_B_CQS8NZev0_1;
	wire w_dff_A_TtFrPdwf5_0;
	wire w_dff_A_4OJKC0OR5_0;
	wire w_dff_A_0YiUR0Ss4_0;
	wire w_dff_A_PXFsuTRE2_0;
	wire w_dff_A_8VaEDlcY7_0;
	wire w_dff_A_Iq24XGYr3_1;
	wire w_dff_B_SYCE2BTn7_0;
	wire w_dff_B_IQmQYXWB0_0;
	wire w_dff_B_q1yVKbPA9_2;
	wire w_dff_B_6XuEDFwA5_2;
	wire w_dff_A_lRlMu4sD7_0;
	wire w_dff_A_M0tghYyO0_0;
	wire w_dff_A_i1S5ziKV7_0;
	wire w_dff_B_Ks7agVIe9_0;
	wire w_dff_B_pbid71fM7_0;
	wire w_dff_B_t2vIVQ5S6_0;
	wire w_dff_B_ijCClu5V1_0;
	wire w_dff_B_TgwTAz0T8_1;
	wire w_dff_B_PrSaw47k1_1;
	wire w_dff_B_wnaAccVc0_2;
	wire w_dff_B_tSC1lAtp1_1;
	wire w_dff_B_q8O96NZW0_1;
	wire w_dff_B_aPhNAm609_0;
	wire w_dff_A_Hu6cMehe4_1;
	wire w_dff_A_lbvI5AZX7_1;
	wire w_dff_A_7SeFFzao1_1;
	wire w_dff_A_DMFkWSl72_2;
	wire w_dff_A_ndWtT0954_2;
	wire w_dff_A_s4K4jVzF7_2;
	wire w_dff_B_WR5Qgovz9_1;
	wire w_dff_B_SollERH45_1;
	wire w_dff_B_DUUwAbIW3_1;
	wire w_dff_B_JOmrejZn1_1;
	wire w_dff_B_NFw4p7kh4_1;
	wire w_dff_B_cnEI5OKQ2_1;
	wire w_dff_B_fNJBprkP0_0;
	wire w_dff_B_zytjr5lS4_1;
	wire w_dff_B_YeRo1S9M1_1;
	wire w_dff_B_xbbZLR3d2_0;
	wire w_dff_A_WorGWE6A7_0;
	wire w_dff_B_A1KkwWH95_3;
	wire w_dff_B_3ApFXNkh1_3;
	wire w_dff_B_shLEtSI70_3;
	wire w_dff_A_U500Ob7a2_0;
	wire w_dff_B_8nMucfrd1_2;
	wire w_dff_B_GGu0UJGT6_2;
	wire w_dff_B_uJt7CJLp2_2;
	wire w_dff_B_HZGkihJZ2_0;
	wire w_dff_B_gx73yGy73_1;
	wire w_dff_B_HFEHj2gJ7_1;
	wire w_dff_B_ovBAT9NH3_1;
	wire w_dff_B_g3sqqxTD0_1;
	wire w_dff_A_zvJHdfOq5_1;
	wire w_dff_A_9QZE4nlL5_1;
	wire w_dff_A_Z4ls5wLR7_1;
	wire w_dff_A_dJDGDyOs2_2;
	wire w_dff_A_TLWREQpl6_2;
	wire w_dff_B_vPKyQSuR3_1;
	wire w_dff_B_luZy6lJH8_0;
	wire w_dff_A_2rrUxUIP9_0;
	wire w_dff_B_u0neskAZ0_3;
	wire w_dff_B_bUL5dkCT3_3;
	wire w_dff_B_cWNoaYa40_3;
	wire w_dff_A_zP6meR3B7_1;
	wire w_dff_A_SvGabuyZ0_1;
	wire w_dff_A_v4aMslTG5_1;
	wire w_dff_A_mEvHV7Qt0_1;
	wire w_dff_A_fO1gaAU48_1;
	wire w_dff_A_pq2AYniU8_1;
	wire w_dff_A_tmTvCkbU6_1;
	wire w_dff_A_fKgJXFjY1_1;
	wire w_dff_A_YCzhrQoY5_0;
	wire w_dff_A_oHrPOyqK9_0;
	wire w_dff_A_D8WSjl5f6_0;
	wire w_dff_A_Pp5xVGwQ0_0;
	wire w_dff_A_SCHK0TrY7_0;
	wire w_dff_A_DEZNKbo81_0;
	wire w_dff_A_nBl04f0e9_0;
	wire w_dff_A_B0I6oQeg1_0;
	wire w_dff_A_w0rZFdYh7_0;
	wire w_dff_A_mLqKf1by0_0;
	wire w_dff_A_TGBdpbH83_0;
	wire w_dff_A_OSUnoYmz9_2;
	wire w_dff_A_dtUhY7JZ5_2;
	wire w_dff_A_tVr9P22h8_2;
	wire w_dff_A_6vPwiSX80_2;
	wire w_dff_A_iRk3bfpv5_2;
	wire w_dff_A_hO7d4Kf21_2;
	wire w_dff_A_gqzlGGGV6_2;
	wire w_dff_A_yKOyCE6l8_2;
	wire w_dff_A_zOV6tKue4_2;
	wire w_dff_A_duMeiHOw2_2;
	wire w_dff_A_VPwrvW8B8_2;
	wire w_dff_A_hmxa8FcC1_1;
	wire w_dff_A_vuWhESbr7_1;
	wire w_dff_A_9ANYxGzJ0_1;
	wire w_dff_A_4tFhnOGS8_1;
	wire w_dff_A_83D1z8j85_1;
	wire w_dff_A_qUKP8lz83_1;
	wire w_dff_A_DmbFSuqA3_1;
	wire w_dff_A_cZg4qVCH0_1;
	wire w_dff_A_Bgh0kV3x6_1;
	wire w_dff_A_Gs6Q1S7n4_1;
	wire w_dff_A_NoSDn8eT1_1;
	wire w_dff_A_C14hPYGJ7_2;
	wire w_dff_A_z19pZXV52_2;
	wire w_dff_A_hAhtHYXq4_2;
	wire w_dff_A_un2wKVAb1_2;
	wire w_dff_A_ym5MLrHo3_2;
	wire w_dff_A_38imtwwk0_2;
	wire w_dff_A_sCNAwjks1_2;
	wire w_dff_A_yXDZaVji8_2;
	wire w_dff_A_gzFbaoh53_2;
	wire w_dff_A_8VT3rPAv2_2;
	wire w_dff_A_BxA3UUOd6_2;
	wire w_dff_B_5JTB6iA73_0;
	wire w_dff_B_7Q94a7311_0;
	wire w_dff_B_ppoLYKA67_0;
	wire w_dff_B_jMsEwQnn4_0;
	wire w_dff_B_15lHvnoi4_0;
	wire w_dff_A_Z6UpHq8j9_0;
	wire w_dff_A_cJa5wY6U9_0;
	wire w_dff_A_zxUPhaMp4_1;
	wire w_dff_A_kgYENZ1Q6_1;
	wire w_dff_A_TXHv3qj30_1;
	wire w_dff_A_mqDiXdHA4_2;
	wire w_dff_A_bzLkRZRK6_2;
	wire w_dff_A_YFww9s9J9_2;
	wire w_dff_B_nX47N2lT6_2;
	wire w_dff_B_14nPjPx62_2;
	wire w_dff_B_DL4bW3ni6_2;
	wire w_dff_B_MAKAai9F3_2;
	wire w_dff_B_czCQDN6x0_2;
	wire w_dff_B_RNkarPww9_2;
	wire w_dff_B_habat80T5_2;
	wire w_dff_B_KsGKK0G76_2;
	wire w_dff_B_ZSSh2JVA7_2;
	wire w_dff_B_VDRNsdvG6_2;
	wire w_dff_B_AdqVhlJ89_2;
	wire w_dff_B_WXIz7OC84_2;
	wire w_dff_B_9D8UaAZR2_2;
	wire w_dff_A_5O7iKcwa2_1;
	wire w_dff_B_ozhs6JXt9_0;
	wire w_dff_B_CJNgHhWI8_0;
	wire w_dff_B_hsTIU0Cm3_0;
	wire w_dff_B_szGITtq51_0;
	wire w_dff_B_yb2WQYBS8_0;
	wire w_dff_B_J0Qggegj6_0;
	wire w_dff_B_kl4sFjwJ4_0;
	wire w_dff_B_Vkys7uUa8_0;
	wire w_dff_B_rHfN2sbM6_0;
	wire w_dff_B_fGBXe76r0_0;
	wire w_dff_B_QWgYZoqw4_0;
	wire w_dff_B_l531TE5W7_1;
	wire w_dff_B_gNhm7Jq30_1;
	wire w_dff_B_Vg4DbODl7_1;
	wire w_dff_B_txrUvoTl4_1;
	wire w_dff_A_aDjpHZsX8_1;
	wire w_dff_A_mKI2h6GU8_1;
	wire w_dff_A_d7F1LZsA6_2;
	wire w_dff_A_WKomwQt33_1;
	wire w_dff_A_pTgtjDkw0_1;
	wire w_dff_A_Jfle1PDM7_1;
	wire w_dff_A_qIt7Kmcb5_1;
	wire w_dff_A_UUP4SJzO6_2;
	wire w_dff_A_mHDmsGcR5_2;
	wire w_dff_A_sZ8z3e048_2;
	wire w_dff_A_4vBQYFhr8_2;
	wire w_dff_A_0gSbFn020_1;
	wire w_dff_A_KEt89Ekc1_0;
	wire w_dff_A_x3Kkhbnz1_0;
	wire w_dff_A_ih6rqG6O8_0;
	wire w_dff_A_U58CLjyT4_0;
	wire w_dff_A_2wQ2Iwbd5_2;
	wire w_dff_A_h94jdN7j6_2;
	wire w_dff_A_bvHmkObR7_2;
	wire w_dff_A_TtR7O4zu8_1;
	wire w_dff_B_tY6y2k0Q3_1;
	wire w_dff_B_2SeKlOP91_1;
	wire w_dff_B_Qnxe6shB7_1;
	wire w_dff_B_0c9EyVMM9_0;
	wire w_dff_A_pOidVMvc1_1;
	wire w_dff_A_oQWicbQb0_2;
	wire w_dff_A_SMHDbw023_0;
	wire w_dff_B_PFjQ1lNL0_3;
	wire w_dff_B_ZdBjMDb04_3;
	wire w_dff_B_RnScCPeN8_3;
	wire w_dff_B_WXlW6o9w3_1;
	wire w_dff_B_fMJ8Nppx0_0;
	wire w_dff_A_sSARz3Q60_0;
	wire w_dff_A_zBlBIKOh8_1;
	wire w_dff_A_ApvMYCUy9_1;
	wire w_dff_A_CEa41W7O4_1;
	wire w_dff_A_hhva3E7w0_1;
	wire w_dff_A_NBZcib8g9_1;
	wire w_dff_A_kLq6bmX15_1;
	wire w_dff_A_qpAvnoHG2_1;
	wire w_dff_A_zVexCDq21_1;
	wire w_dff_A_ImVemRGn4_2;
	wire w_dff_A_Lohcljm11_2;
	wire w_dff_B_lTVgmxFJ7_0;
	wire w_dff_B_HkOfbMn44_0;
	wire w_dff_B_2kSKJuTH6_0;
	wire w_dff_B_0Jc9uF4g1_0;
	wire w_dff_A_3xcn83Zx7_0;
	wire w_dff_B_YExEAZQO6_0;
	wire w_dff_B_u4VORMBn5_0;
	wire w_dff_B_qKnH7FET3_0;
	wire w_dff_B_B7L1Bb4k5_0;
	wire w_dff_B_9Lpsubch3_0;
	wire w_dff_A_fzv4lvqZ5_2;
	wire w_dff_A_ObJL9Qaa6_1;
	wire w_dff_A_Qbg4QAcq7_1;
	wire w_dff_A_6kHp5xAf2_2;
	wire w_dff_A_tidmV6Lo7_2;
	wire w_dff_A_fjKKoOcc0_0;
	wire w_dff_A_ZCBBHjxo5_1;
	wire w_dff_A_RpbsJLj51_1;
	wire w_dff_A_bVqstwWx0_1;
	wire w_dff_A_Czkz7sXW1_1;
	wire w_dff_B_Z7Hernbb6_1;
	wire w_dff_B_ubAYFKGy2_1;
	wire w_dff_A_2IVlRPjg5_1;
	wire w_dff_B_3aaOt5mu4_1;
	wire w_dff_B_aqXTkkMr3_0;
	wire w_dff_B_VgwORNHx7_0;
	wire w_dff_B_Hn1TlILC1_0;
	wire w_dff_B_kXyk0Mo37_1;
	wire w_dff_A_0y4SqIvc2_0;
	wire w_dff_A_z5vuix598_0;
	wire w_dff_B_Y6P4RbDG7_1;
	wire w_dff_B_tU88pgl64_1;
	wire w_dff_A_Mr7Yxxtc5_0;
	wire w_dff_A_Kv3wMfzj6_0;
	wire w_dff_B_mjwAJ0fu9_0;
	wire w_dff_B_pJ9vBfb10_1;
	wire w_dff_B_QBUlf6Y68_1;
	wire w_dff_B_fFkLKxll7_1;
	wire w_dff_B_E3nHGAMP2_1;
	wire w_dff_B_d1fElbSb7_0;
	wire w_dff_B_Qwl99s273_0;
	wire w_dff_B_Do6o7OWl5_1;
	wire w_dff_B_qsInAYaB2_1;
	wire w_dff_B_YL6HbYWE5_1;
	wire w_dff_A_iiFMhJsK0_1;
	wire w_dff_A_H2zRB4zY0_1;
	wire w_dff_B_ZtZugRSf2_1;
	wire w_dff_B_CaBe6qHK8_1;
	wire w_dff_A_yHGBWbls2_0;
	wire w_dff_A_JChnqbdl4_0;
	wire w_dff_A_kl66bIPt4_0;
	wire w_dff_A_OF2BZT4e7_0;
	wire w_dff_B_GpNB0XTN4_0;
	wire w_dff_A_eCFQ9eAD7_1;
	wire w_dff_A_khPh2FFN8_1;
	wire w_dff_A_z5f1lVWD4_2;
	wire w_dff_A_6eS5xXQT3_2;
	wire w_dff_A_xE7CJdnU0_2;
	wire w_dff_A_K5vSNaX49_2;
	wire w_dff_B_PusZ0kJy6_1;
	wire w_dff_B_Nv2GfN377_1;
	wire w_dff_B_ymDCuxVv0_1;
	wire w_dff_A_JFeIDYY74_0;
	wire w_dff_B_C0Fl309u4_2;
	wire w_dff_A_TiB3qEKA3_1;
	wire w_dff_A_UVDxzX8X4_1;
	wire w_dff_A_O31Yevz94_1;
	wire w_dff_B_ZA4Xncnc2_2;
	wire w_dff_B_3TZf6n5G1_2;
	wire w_dff_B_5ysRGQcf9_1;
	wire w_dff_B_3Teu5xFQ4_1;
	wire w_dff_B_7vdPgLY42_1;
	wire w_dff_B_jWr6xEqu8_0;
	wire w_dff_B_7SgsIywN8_0;
	wire w_dff_A_Nwsjq0xo4_2;
	wire w_dff_B_oW9LfIcp4_1;
	wire w_dff_B_3fcaVetG8_1;
	wire w_dff_B_6GLiXLf15_1;
	wire w_dff_A_OY2GCQl84_1;
	wire w_dff_A_iJX6d4KT1_1;
	wire w_dff_A_h1U14QZ20_1;
	wire w_dff_A_cQXYitet4_2;
	wire w_dff_A_nBSbsODQ5_2;
	wire w_dff_A_sPbkiv5R3_2;
	wire w_dff_A_MwT9xHbC5_2;
	wire w_dff_A_45ig0oRf4_1;
	wire w_dff_A_XNuT9Fvx8_1;
	wire w_dff_A_tPqs1ct78_1;
	wire w_dff_A_JEStj55Q1_2;
	wire w_dff_A_efvVhaa88_2;
	wire w_dff_A_DwRq8D7V4_0;
	wire w_dff_A_OzhMKkGv7_0;
	wire w_dff_A_PVARDvkW4_2;
	wire w_dff_A_puSTSz594_2;
	wire w_dff_A_EL2YGJlr6_2;
	wire w_dff_A_y6OI6irt9_2;
	wire w_dff_A_ayd9RTX27_1;
	wire w_dff_A_0UwmGFFC3_1;
	wire w_dff_A_dc4sKXuE5_1;
	wire w_dff_A_pJ3juYXa6_0;
	wire w_dff_A_UyoE6NVP6_0;
	wire w_dff_A_AEGITx9G9_1;
	wire w_dff_A_n01tZAbE4_0;
	wire w_dff_A_scg5wolC8_2;
	wire w_dff_A_8FLMUrlX5_2;
	wire w_dff_A_0dGGcx4t0_2;
	wire w_dff_A_sQxHYeYf6_2;
	wire w_dff_A_zwqU6G3F3_0;
	wire w_dff_A_ndypIZMF9_0;
	wire w_dff_A_Jz517UPj8_0;
	wire w_dff_A_cIUoVB911_0;
	wire w_dff_B_6Uzw4xNH4_0;
	wire w_dff_B_Oz0vXoYE2_0;
	wire w_dff_B_SfEUcmPy1_0;
	wire w_dff_B_3Tn9GTCJ1_0;
	wire w_dff_B_fwNpmsjn6_0;
	wire w_dff_B_ddHmRJrI4_0;
	wire w_dff_B_QLeR7zmG1_0;
	wire w_dff_B_kW1l0wiA6_0;
	wire w_dff_B_huqK92bP3_0;
	wire w_dff_A_kdtt9xD15_2;
	wire w_dff_A_sjnLsLoA7_2;
	wire w_dff_A_G4bUzfxV5_2;
	wire w_dff_A_SCpKaUiZ8_2;
	wire w_dff_A_W39ACTMm9_2;
	wire w_dff_A_AtOJHKKB4_2;
	wire w_dff_A_VIUQCjfj6_2;
	wire w_dff_A_a5wMNEEO6_2;
	wire w_dff_A_ZJcudOfX8_0;
	wire w_dff_A_OJPfcFCa2_0;
	wire w_dff_A_2EEPRluq6_0;
	wire w_dff_A_kKrqoSoW7_0;
	wire w_dff_B_3h42XZni7_1;
	wire w_dff_B_kltxwDtL7_1;
	wire w_dff_B_aEOYgQuj1_1;
	wire w_dff_B_iyLyyVWW7_1;
	wire w_dff_B_ZxTVggiG3_1;
	wire w_dff_B_ZNVwHKRe3_0;
	wire w_dff_A_dWwjfL9n6_0;
	wire w_dff_A_HaSaHwL92_0;
	wire w_dff_A_Au7l3aAv2_0;
	wire w_dff_A_gbf3SjqU5_0;
	wire w_dff_A_oXNKXIQd4_2;
	wire w_dff_A_RRAZWhbs1_2;
	wire w_dff_A_nByLp5Ye4_0;
	wire w_dff_A_vlp8hzqz8_2;
	wire w_dff_A_8G95VIjC4_2;
	wire w_dff_B_IAYrVm0P9_1;
	wire w_dff_B_kbc6CHlm6_0;
	wire w_dff_A_Rbqv7i2E2_1;
	wire w_dff_B_3Zls9Asu0_3;
	wire w_dff_B_UKTj6RAy9_3;
	wire w_dff_B_mqa966gy6_3;
	wire w_dff_B_0Qpqs9IT5_1;
	wire w_dff_B_qOHNn4DT0_1;
	wire w_dff_B_mA1TS2tU5_1;
	wire w_dff_B_2WoV4lU33_1;
	wire w_dff_A_gYiziej66_1;
	wire w_dff_A_EuaQOspZ3_1;
	wire w_dff_A_2pHJVp7l8_1;
	wire w_dff_A_jZRrQYj11_2;
	wire w_dff_A_9JmFPU7u0_2;
	wire w_dff_A_36uqRPDS7_1;
	wire w_dff_B_aHADKo1m3_3;
	wire w_dff_B_BfoOu98b4_3;
	wire w_dff_B_a8BNTn3r7_3;
	wire w_dff_B_HTpOZOSe8_3;
	wire w_dff_B_e3iksa357_3;
	wire w_dff_B_9juV44ph8_3;
	wire w_dff_A_ZKbKDlC72_0;
	wire w_dff_A_hvwHxbc04_1;
	wire w_dff_A_Jkc8FQ2x6_1;
	wire w_dff_A_ML8Wsi7R7_0;
	wire w_dff_A_VmKgOIih9_0;
	wire w_dff_A_QZZj3G500_1;
	wire w_dff_B_qkfBigxd2_3;
	wire w_dff_B_CuiEmr8G7_3;
	wire w_dff_A_SktWqd4B6_1;
	wire w_dff_A_ngQMY0wi1_1;
	wire w_dff_A_pnXBJf900_1;
	wire w_dff_A_HraerFyz3_1;
	wire w_dff_A_CAXAfBzv5_1;
	wire w_dff_A_qthwE6YC3_2;
	wire w_dff_A_sGBZWvyE2_2;
	wire w_dff_A_eSlwqHHA1_2;
	wire w_dff_A_X6IwQgEE1_2;
	wire w_dff_A_pNsegoOF1_2;
	wire w_dff_A_rPHqTFGY3_0;
	wire w_dff_A_QROsBE3b5_0;
	wire w_dff_A_o3YWIpC56_0;
	wire w_dff_A_Babz9X3p5_2;
	wire w_dff_A_Y3f56pMO3_2;
	wire w_dff_A_xOecG1PY4_2;
	wire w_dff_A_r1HWMIYL7_2;
	wire w_dff_A_3Dlfw6DB4_1;
	wire w_dff_A_8RbOiNs66_1;
	wire w_dff_A_ZukS50L22_1;
	wire w_dff_A_DHGzt0N55_0;
	wire w_dff_A_RppjfKcu5_0;
	wire w_dff_A_hEyGmNLP2_0;
	wire w_dff_A_RACd9pjg9_0;
	wire w_dff_A_4PgoHSVp7_1;
	wire w_dff_A_oDlAgc7P2_1;
	wire w_dff_A_ybsNGNwS9_1;
	wire w_dff_A_uXXzrEnG6_1;
	wire w_dff_A_JkA8zOvk6_1;
	wire w_dff_B_y90EBVFx6_1;
	wire w_dff_B_h2dKfwho3_0;
	wire w_dff_A_aPGmUDHU2_0;
	wire w_dff_A_5v8xR5wt0_0;
	wire w_dff_A_wgMpoDW27_0;
	wire w_dff_A_otD5R4BN9_0;
	wire w_dff_A_yX6ndfia3_0;
	wire w_dff_A_NQlKKxwd2_0;
	wire w_dff_A_NkwA5IIM6_1;
	wire w_dff_A_8Xx64vZW0_1;
	wire w_dff_A_UpKDQn5S3_1;
	wire w_dff_A_r5Tudtj48_0;
	wire w_dff_A_Rn3uLTyX2_1;
	wire w_dff_A_O0F2LtgJ8_1;
	wire w_dff_A_IlhzGVfX4_1;
	wire w_dff_A_WbvVSi4P5_1;
	wire w_dff_A_p9A7aHDN9_1;
	wire w_dff_A_U7BP3JGa3_1;
	wire w_dff_A_qmAdwVV27_1;
	wire w_dff_A_mz2Ma50S4_1;
	wire w_dff_A_3g9wCvOT0_1;
	wire w_dff_A_im6BpvSm3_2;
	wire w_dff_A_37RYzBOf2_2;
	wire w_dff_A_Cd5N8OoT3_2;
	wire w_dff_A_ImJQOAUL9_2;
	wire w_dff_A_b7z7NBeM2_2;
	wire w_dff_A_vZuHoIeq9_2;
	wire w_dff_A_UHz0db1u2_2;
	wire w_dff_A_V3ymdB0E2_0;
	wire w_dff_A_Zn9s1wEB5_0;
	wire w_dff_A_QvwrTc9j0_1;
	wire w_dff_A_ZwLwUUqu8_1;
	wire w_dff_A_BmJHWTNA3_1;
	wire w_dff_B_koyEFjA78_3;
	wire w_dff_B_vdjU1Jx73_3;
	wire w_dff_B_9BanF2Hg6_3;
	wire w_dff_A_jXoD36EM4_0;
	wire w_dff_A_MJe5nHEv3_0;
	wire w_dff_A_z3nenk1G6_0;
	wire w_dff_A_b59GNd0f5_0;
	wire w_dff_A_x9e5xlAp3_0;
	wire w_dff_A_lTvxQf551_0;
	wire w_dff_A_y2vQ4Fxq2_0;
	wire w_dff_A_rVInVeyA9_0;
	wire w_dff_A_bOjiu0b69_0;
	wire w_dff_A_orL5Xhbm1_2;
	wire w_dff_A_6LUEUNu30_2;
	wire w_dff_A_p8SEAqju9_2;
	wire w_dff_A_A7y32vC20_2;
	wire w_dff_A_CWC3RigB3_2;
	wire w_dff_A_5arkXnx99_2;
	wire w_dff_A_Ul0QIhXY5_2;
	wire w_dff_A_O9EwWugZ5_2;
	wire w_dff_A_dBm7to3B0_2;
	wire w_dff_A_T7vBhMUj8_1;
	wire w_dff_A_aK57UsaL5_1;
	wire w_dff_A_9AWkHB5g3_1;
	wire w_dff_A_olxTOttA6_1;
	wire w_dff_A_gtx9BhxV3_1;
	wire w_dff_A_BwpN446w0_1;
	wire w_dff_A_UZVNZD1m5_1;
	wire w_dff_A_MfMg31SE1_1;
	wire w_dff_A_KVSAQB6x9_1;
	wire w_dff_A_wcuik72z9_1;
	wire w_dff_A_GWnmYwJh7_1;
	wire w_dff_A_lAyJxtep3_1;
	wire w_dff_A_pyxeLgzK9_1;
	wire w_dff_A_REnI5YUr6_2;
	wire w_dff_A_wCBDH8kw1_2;
	wire w_dff_A_7cPEC6TA0_2;
	wire w_dff_A_Q2HUV31o5_2;
	wire w_dff_A_yCjTMs0C2_2;
	wire w_dff_A_o0x1YyjQ7_2;
	wire w_dff_A_QFjLQ9A31_0;
	wire w_dff_A_Qj78QzEa8_0;
	wire w_dff_A_yz5Me03f0_0;
	wire w_dff_A_lo2DMc579_0;
	wire w_dff_A_pZgIn6Mn2_0;
	wire w_dff_A_9lcQDSgC5_0;
	wire w_dff_A_Y3zWFNcr3_0;
	wire w_dff_A_Q3jL4xQ95_0;
	wire w_dff_A_6y2D3p9b0_0;
	wire w_dff_A_YLSA4Nci2_0;
	wire w_dff_A_qyCW8pT93_0;
	wire w_dff_A_1rrweAxJ5_0;
	wire w_dff_A_U1nsvXFK9_0;
	wire w_dff_A_QlUl0lp24_1;
	wire w_dff_A_bir5F7eH1_1;
	wire w_dff_A_5sMzEO2c4_1;
	wire w_dff_A_EAuUh3eM7_1;
	wire w_dff_A_F2iBFrld3_1;
	wire w_dff_A_sfCHYGZB6_1;
	wire w_dff_A_HgWHZUp25_1;
	wire w_dff_A_BbBgQ5tH3_1;
	wire w_dff_A_x4Ctfyb41_1;
	wire w_dff_A_xW3tbapP7_1;
	wire w_dff_A_EoSQQ67C1_1;
	wire w_dff_A_frGaIkcL7_1;
	wire w_dff_A_01HEKiPv4_1;
	wire w_dff_A_apbNwcZG3_1;
	wire w_dff_A_bnQIZaMM6_1;
	wire w_dff_A_Iu4eF7L16_1;
	wire w_dff_A_gFnsGjdN1_1;
	wire w_dff_A_q46AWpcw8_1;
	wire w_dff_A_MZzf122x5_1;
	wire w_dff_A_3CMLQwKD1_1;
	wire w_dff_A_VmAgNmDG8_1;
	wire w_dff_A_fQNzXRoa0_1;
	wire w_dff_A_VYsKwuZb0_1;
	wire w_dff_A_xKz9M7fS3_1;
	wire w_dff_A_ubaIKEJ61_1;
	wire w_dff_A_juqvY5ge5_1;
	wire w_dff_A_Ieevp0XE1_2;
	wire w_dff_A_mcVKIyD40_2;
	wire w_dff_A_CL60yoVR8_2;
	wire w_dff_A_5yu8exKE4_2;
	wire w_dff_A_Uv0Xm1Bb8_2;
	wire w_dff_A_SX3EYtG92_2;
	wire w_dff_A_gfvpNFiO8_2;
	wire w_dff_A_7Y2f3YIX2_2;
	wire w_dff_A_6vzYT7Q89_2;
	wire w_dff_A_WXjVGyeo0_2;
	wire w_dff_A_icESleKK9_2;
	wire w_dff_A_9mB63LIe3_2;
	wire w_dff_A_Srm5kXMA6_2;
	wire w_dff_A_O64eRFnd9_0;
	wire w_dff_A_Zgm7zyNm4_0;
	wire w_dff_A_MY5eYnyZ8_0;
	wire w_dff_A_jQb7DLmM0_0;
	wire w_dff_A_wbPRxEi36_1;
	wire w_dff_A_BYuIiKA37_1;
	wire w_dff_B_ToFRmcGQ2_0;
	wire w_dff_A_2YbzKGby8_0;
	wire w_dff_A_i5Ds5bN29_0;
	wire w_dff_A_F0VobcyN5_2;
	wire w_dff_A_vjNhp4wO4_2;
	wire w_dff_A_f46lkmuH0_2;
	wire w_dff_A_LupTeA0c5_2;
	wire w_dff_A_BkhVbplY0_2;
	wire w_dff_A_ZEPqOYZy9_2;
	wire w_dff_A_cf21gQDV6_2;
	wire w_dff_A_OSkJvifp7_2;
	wire w_dff_A_igeVjMAd9_0;
	wire w_dff_A_DHZW8wk15_0;
	wire w_dff_A_wM0pIoMX7_2;
	wire w_dff_A_9f9VqMzN8_2;
	wire w_dff_A_RDucMg3G7_0;
	wire w_dff_A_8a8GQP3p1_0;
	wire w_dff_A_ZHy6qTz98_0;
	wire w_dff_A_eGnqnVtQ8_0;
	wire w_dff_A_MU4ralJA4_0;
	wire w_dff_A_xPo6llk43_0;
	wire w_dff_A_sitLDePJ2_0;
	wire w_dff_A_3HYZCYkx5_0;
	wire w_dff_A_0a75YB7r5_0;
	wire w_dff_A_yVn1imyF0_0;
	wire w_dff_A_UeTQRlg70_0;
	wire w_dff_A_qUiSdLMH8_0;
	wire w_dff_A_fpbiBcSI7_0;
	wire w_dff_A_tKvRylP32_0;
	wire w_dff_A_QcUlEmmC5_0;
	wire w_dff_A_ExKlLBAI1_0;
	wire w_dff_A_3ntxPuHO3_0;
	wire w_dff_A_8TwwIrNO1_0;
	wire w_dff_A_XSZ6sDf47_0;
	wire w_dff_A_f96h5L4Q5_0;
	wire w_dff_A_hr5bMELX1_0;
	wire w_dff_A_9B9zPNJo4_0;
	wire w_dff_A_OnG5Egny5_0;
	wire w_dff_A_67LEQ4PA8_0;
	wire w_dff_A_4RRiHoEs0_0;
	wire w_dff_A_hrOe6sHs6_2;
	wire w_dff_A_izinCztL5_2;
	wire w_dff_A_dh3MLIUd3_2;
	wire w_dff_A_mfRb8nQY3_2;
	wire w_dff_A_VqJR3Y8P5_2;
	wire w_dff_A_NQkrsk995_2;
	wire w_dff_A_h2SzWK0d5_2;
	wire w_dff_A_7cqMFiTh1_2;
	wire w_dff_A_4WHxmVZT4_2;
	wire w_dff_A_2RlqY59s8_2;
	wire w_dff_A_dzuvx9Vi0_2;
	wire w_dff_A_2eAAhsCk3_2;
	wire w_dff_A_NMzqwxXi2_2;
	wire w_dff_A_2KKKMxEO2_0;
	wire w_dff_A_kklXdGwp8_0;
	wire w_dff_A_kSUrakpl0_0;
	wire w_dff_A_Ze8pyVHu9_0;
	wire w_dff_A_Raxmyxn51_0;
	wire w_dff_A_uZI1uxxm9_0;
	wire w_dff_A_00EfuHWr5_0;
	wire w_dff_A_GMZfWSSF1_0;
	wire w_dff_A_ZdbF9i3h5_0;
	wire w_dff_A_TlThXpMa5_0;
	wire w_dff_A_IogcAiqi6_0;
	wire w_dff_A_KkVA1EWI4_0;
	wire w_dff_A_xqHPYubh0_0;
	wire w_dff_A_eZKsSnD04_0;
	wire w_dff_A_gETiBfap9_0;
	wire w_dff_A_bqP0hXwQ1_0;
	wire w_dff_A_hhWxJAtF1_0;
	wire w_dff_A_qJzcbsiQ5_0;
	wire w_dff_A_fm3xRMa22_0;
	wire w_dff_A_Bzdl7SUk7_0;
	wire w_dff_A_60nDHZ7A3_0;
	wire w_dff_A_r1a9DKN97_0;
	wire w_dff_A_twgUN3sy1_0;
	wire w_dff_A_EjT8DoTg4_0;
	wire w_dff_A_kC8sCidG6_0;
	wire w_dff_A_4EBPQli13_0;
	wire w_dff_A_w1Dw10HK4_0;
	wire w_dff_A_6X0v1u8U8_0;
	wire w_dff_A_8j4ASYBC0_0;
	wire w_dff_A_KNHB5mhX4_0;
	wire w_dff_A_tTRGCba08_2;
	wire w_dff_A_9XtKLYwL2_2;
	wire w_dff_A_mVGq03yY8_2;
	wire w_dff_A_l0g4ARMN5_2;
	wire w_dff_A_v63deK9y4_2;
	wire w_dff_A_sNeVUY8j4_2;
	wire w_dff_A_g4AOfy8l0_2;
	wire w_dff_A_vzpxu5bz9_2;
	wire w_dff_A_zifp6hnE8_2;
	wire w_dff_A_NM5hwlAr7_2;
	wire w_dff_A_bKRGQ5hY0_2;
	wire w_dff_A_3tXTZQie8_2;
	wire w_dff_A_8RFzvmkn8_2;
	wire w_dff_A_ImjYv5sH8_2;
	wire w_dff_A_vEtMHDQE6_2;
	wire w_dff_A_pbO59dpv8_2;
	wire w_dff_A_hXaqpHIU1_1;
	wire w_dff_A_q6PhK3IL6_1;
	wire w_dff_A_5XEw9YYy7_1;
	wire w_dff_A_ZuZ08gKE8_1;
	wire w_dff_A_QVJ07exF8_1;
	wire w_dff_A_0oqXYBeD5_1;
	wire w_dff_A_5QKhZG5x9_1;
	wire w_dff_A_rbymtoR63_1;
	wire w_dff_A_aVB2aesx0_1;
	wire w_dff_A_S5mYsdfC6_1;
	wire w_dff_A_kzp80mkF1_1;
	wire w_dff_A_ekH6s8rA2_1;
	wire w_dff_A_7UXBHXrr8_1;
	wire w_dff_A_hMqIvqxr9_1;
	wire w_dff_A_P99KkVrv0_1;
	wire w_dff_A_QdsBB7La3_2;
	wire w_dff_A_USn8cusi8_2;
	wire w_dff_A_aIuZPe2o1_2;
	wire w_dff_A_mH5eGrmt9_2;
	wire w_dff_A_319wHlOC7_2;
	wire w_dff_A_dz3mmXd33_2;
	wire w_dff_A_vDtdNpEu0_2;
	wire w_dff_A_msf1W9BA9_2;
	wire w_dff_A_gEkg5rZd3_2;
	wire w_dff_A_hcecLVZx0_2;
	wire w_dff_A_J7f9aLGS7_2;
	wire w_dff_A_FFiuvnBX3_2;
	wire w_dff_A_OcLCl1li7_2;
	wire w_dff_A_wOa8UGtJ2_2;
	wire w_dff_A_7Mf11hn86_2;
	wire w_dff_A_9oa9JSFi3_2;
	wire w_dff_A_o8jC3wy89_0;
	wire w_dff_B_q5AGVv120_1;
	wire w_dff_A_FCrx7MFn5_0;
	wire w_dff_A_LzAARKpC1_2;
	wire w_dff_A_TBk7QCdd1_1;
	wire w_dff_A_Im8C63OO4_1;
	wire w_dff_B_cMsoc7sh1_2;
	wire w_dff_B_0IyZh3r87_1;
	wire w_dff_B_Ja2zN20d8_1;
	wire w_dff_A_QPOjnUF42_1;
	wire w_dff_A_CiMjb1I22_1;
	wire w_dff_A_e41t7c4X0_1;
	wire w_dff_A_fRyBsshg1_1;
	wire w_dff_A_RGq7ptNu3_1;
	wire w_dff_A_rM0bwNhF2_1;
	wire w_dff_A_iI3BAws32_2;
	wire w_dff_A_NuGbAMwL1_1;
	wire w_dff_B_ZH0hIGre5_1;
	wire w_dff_B_w8aVsJPu0_1;
	wire w_dff_B_7aS6B6hN6_1;
	wire w_dff_B_dP8ERMqf7_1;
	wire w_dff_B_AFu2vZVl4_0;
	wire w_dff_B_7Nb557uG9_0;
	wire w_dff_A_FZiDhw6C1_1;
	wire w_dff_A_GqESV7yA9_1;
	wire w_dff_A_S2bmOonB3_1;
	wire w_dff_A_vLREaknN6_2;
	wire w_dff_A_FKNrCzj53_2;
	wire w_dff_B_I3nt5hgZ5_0;
	wire w_dff_A_xzFq9UPv6_0;
	wire w_dff_A_XCiI2xG81_0;
	wire w_dff_A_i59xcJY51_1;
	wire w_dff_A_63v7l7Vq9_1;
	wire w_dff_A_QWWqCtkg0_0;
	wire w_dff_A_Mjh3b7UO7_1;
	wire w_dff_A_6m0bHzbb6_0;
	wire w_dff_A_PrZhEze71_2;
	wire w_dff_A_Xg3pnDtJ4_2;
	wire w_dff_A_BtUpt0110_2;
	wire w_dff_A_pR8uKgO07_2;
	wire w_dff_A_i85muIC40_1;
	wire w_dff_A_vHIhuok02_2;
	wire w_dff_A_V3pXokVU0_2;
	wire w_dff_A_cxfkScNB3_2;
	wire w_dff_A_Jgno6nkh7_1;
	wire w_dff_A_igQewKez1_2;
	wire w_dff_A_7sF9HlrM6_2;
	wire w_dff_B_NU60nkyg4_2;
	wire w_dff_B_MPLAYylK2_2;
	wire w_dff_A_yVgeO5789_0;
	wire w_dff_A_F2nHkO901_0;
	wire w_dff_A_pZJDfEC69_0;
	wire w_dff_A_aVsadp7V2_0;
	wire w_dff_A_470PHLTQ0_1;
	wire w_dff_A_qq2etdfU1_1;
	wire w_dff_A_wcSOMHkc7_1;
	wire w_dff_A_rGYIVoJs5_1;
	wire w_dff_A_UY8yXUs39_1;
	wire w_dff_A_nhFB6Wdy6_1;
	wire w_dff_B_v9vq1SUv1_1;
	wire w_dff_A_qLHi8o0E6_0;
	wire w_dff_A_2sF6EAVe2_0;
	wire w_dff_A_lwoF2VS19_1;
	wire w_dff_A_3fRE8kKZ3_1;
	wire w_dff_A_PDBLOkoQ0_1;
	wire w_dff_A_rwJfIo3F3_1;
	wire w_dff_A_CZISefcV8_1;
	wire w_dff_A_dfXod0py9_2;
	wire w_dff_A_wZ3zF3iC5_2;
	wire w_dff_B_Yea19fe24_0;
	wire w_dff_A_lrS1MQPf1_1;
	wire w_dff_B_LzLWH8KM7_1;
	wire w_dff_A_IHmCwTyd5_1;
	wire w_dff_A_Uky4l53N4_0;
	wire w_dff_A_AdDCGg8T0_2;
	wire w_dff_A_ufRxWv6b1_2;
	wire w_dff_B_Ao6zYikO0_0;
	wire w_dff_B_2iHUmqcd2_1;
	wire w_dff_B_KdKHTE9v4_1;
	wire w_dff_A_bXVRJXjo6_1;
	wire w_dff_A_lE9FDNoY9_2;
	wire w_dff_A_SsxPyY0o6_2;
	wire w_dff_A_5zizEvxm1_2;
	wire w_dff_A_irrr2R7R5_2;
	wire w_dff_A_4iVzRieL8_2;
	wire w_dff_A_NINKWWWh6_0;
	wire w_dff_A_3ISqDeBM3_0;
	wire w_dff_A_P8mMtLYv0_0;
	wire w_dff_A_jwSb8tfs3_1;
	wire w_dff_A_hMeOEyx59_1;
	wire w_dff_B_URPYmcRE4_3;
	wire w_dff_B_4euaslRD6_3;
	wire w_dff_A_Ym3uFM6E0_0;
	wire w_dff_A_t7bUeRsk7_0;
	wire w_dff_A_xJcSlXtV9_0;
	wire w_dff_A_QZyOovr08_0;
	wire w_dff_A_Nai817tk0_0;
	wire w_dff_A_Ai49wWVh2_0;
	wire w_dff_A_Vbndpgai8_0;
	wire w_dff_A_pl2QGNfM2_0;
	wire w_dff_A_e30Kr4GF0_0;
	wire w_dff_A_dozsGobe8_0;
	wire w_dff_A_0JOd5oEu3_0;
	wire w_dff_A_L9d9XzyQ5_0;
	wire w_dff_A_slHywqOc0_0;
	wire w_dff_A_FGocdD9N7_0;
	wire w_dff_A_A7wXq5rE3_0;
	wire w_dff_A_D6sZjnq76_0;
	wire w_dff_A_3cS0A53x5_0;
	wire w_dff_A_26Dzk5OR2_0;
	wire w_dff_A_82IQy6tX3_0;
	wire w_dff_A_96QSHZBZ9_0;
	wire w_dff_A_XTPuqfGv3_0;
	wire w_dff_A_1IoTyaGF1_0;
	wire w_dff_A_cuxQ11mA4_1;
	wire w_dff_A_fLATu3s21_1;
	wire w_dff_A_I1W9SNlC3_1;
	wire w_dff_A_LpwxVUGw7_1;
	wire w_dff_A_SgKpglzj9_1;
	wire w_dff_A_qcuyOwu73_0;
	wire w_dff_A_Nzq8A0ba9_0;
	wire w_dff_A_oRBHHkxw3_0;
	wire w_dff_A_TEJfY3zX3_0;
	wire w_dff_A_0yt1rV2I1_2;
	wire w_dff_A_sejDLEvb2_2;
	wire w_dff_A_jReJ0Rc02_2;
	wire w_dff_A_KbtCw2Be9_2;
	wire w_dff_A_uDb9li524_2;
	wire w_dff_A_sHrhhkQJ2_2;
	wire w_dff_A_CL3hdu101_1;
	wire w_dff_A_Uzp6K9k27_1;
	wire w_dff_A_ghBuExEe4_1;
	wire w_dff_A_P1pQTy2S6_1;
	wire w_dff_A_GfNU974E0_1;
	wire w_dff_A_G0TcI57k1_1;
	wire w_dff_A_YGVxfLki0_1;
	wire w_dff_A_VlSN2j3M8_2;
	wire w_dff_A_T0u8ZC016_2;
	wire w_dff_A_qZ6PRYIe3_2;
	wire w_dff_A_wYlX2dmG9_2;
	wire w_dff_A_KOyNZY7v0_2;
	wire w_dff_A_c7UUtwWp8_2;
	wire w_dff_A_q1KHmSbO4_2;
	wire w_dff_A_nj5ryxbi9_0;
	wire w_dff_A_06UoBpWW4_2;
	wire w_dff_A_G2iJTLxm5_0;
	wire w_dff_A_CoFQTjdU4_0;
	wire w_dff_A_0FsblvdM4_1;
	wire w_dff_A_awiYCCAm5_1;
	wire w_dff_A_DvqUdaea1_1;
	wire w_dff_A_IVfs17j22_1;
	wire w_dff_A_L7dgG65K4_1;
	wire w_dff_A_yESD0x6O4_1;
	wire w_dff_A_275NIoSS5_1;
	wire w_dff_A_rhmi6y775_1;
	wire w_dff_A_Ihnghm883_1;
	wire w_dff_A_sjoCCasm5_1;
	wire w_dff_A_Q7ura78J7_1;
	wire w_dff_A_92H3T4840_1;
	wire w_dff_A_uDYQkja50_1;
	wire w_dff_A_umE1GkFi4_1;
	wire w_dff_A_BFcuhVbu6_1;
	wire w_dff_A_k97hcDSh2_1;
	wire w_dff_A_aunUDTkh1_1;
	wire w_dff_A_Su7s7ao33_1;
	wire w_dff_A_OLc4brm52_1;
	wire w_dff_B_nuHoV5pA2_0;
	wire w_dff_B_Dh2jux470_1;
	wire w_dff_B_0LuljrnG7_1;
	wire w_dff_A_c2WzAXFN8_0;
	wire w_dff_A_S9HSg5NO7_0;
	wire w_dff_A_7Og8lSIe5_0;
	wire w_dff_A_Bn0WMGDC3_0;
	wire w_dff_A_mMUfU7md6_0;
	wire w_dff_A_GsTMAoUY0_0;
	wire w_dff_A_pnpF4iId6_0;
	wire w_dff_A_fjjXIW3l0_0;
	wire w_dff_A_IwzbsjN37_0;
	wire w_dff_A_J5Js87zm5_1;
	wire w_dff_A_5N0sKK5d5_1;
	wire w_dff_A_KiT15BBB8_1;
	wire w_dff_A_pH3RywLK4_0;
	wire w_dff_A_mgJE9RLR9_1;
	wire w_dff_B_xrpfOxV02_0;
	wire w_dff_A_i2aqhp5d0_0;
	wire w_dff_A_luOPKde94_0;
	wire w_dff_B_UDmTyMk91_0;
	wire w_dff_A_p2P0Q2Iy0_0;
	wire w_dff_A_HoFi2L3R1_1;
	wire w_dff_B_MNYOayjY1_0;
	wire w_dff_B_WMEaKdvL2_1;
	wire w_dff_A_PYEzkkyH2_1;
	wire w_dff_A_yvxDBaBU2_1;
	wire w_dff_A_SZozDlnA3_1;
	wire w_dff_A_5HCXgE3r5_1;
	wire w_dff_A_FDG7s6lR2_1;
	wire w_dff_A_C3p8AZF36_1;
	wire w_dff_A_XHC4JfNo2_1;
	wire w_dff_A_Jks76VVu9_2;
	wire w_dff_A_JpmrROEI9_2;
	wire w_dff_A_htK27Vyk1_2;
	wire w_dff_A_MFiCQyL13_2;
	wire w_dff_A_mdaEY9wk8_2;
	wire w_dff_A_FpXd7hDV2_2;
	wire w_dff_A_59Z4Cv8n6_2;
	wire w_dff_B_igReF1fn0_0;
	wire w_dff_B_IpaO9w8W7_1;
	wire w_dff_A_kyk90hop2_1;
	wire w_dff_B_xzNoOxiA6_1;
	wire w_dff_A_v5uxyzdr9_0;
	wire w_dff_A_HZLZcV8W5_0;
	wire w_dff_A_kgIT8jEI1_0;
	wire w_dff_A_YG7pT8e90_1;
	wire w_dff_A_9jxpiqiL7_1;
	wire w_dff_A_Q14htJgy1_1;
	wire w_dff_A_UANVtvih1_2;
	wire w_dff_A_oSJIeN5g9_1;
	wire w_dff_A_0HjbQwMa6_2;
	wire w_dff_A_O5qOvHQS3_1;
	wire w_dff_A_8bu2HjsL3_1;
	wire w_dff_A_stTYGT9I3_0;
	wire w_dff_A_gFIWSjUS3_0;
	wire w_dff_A_mo8oFZxj4_1;
	wire w_dff_A_jBWtepp39_1;
	wire w_dff_A_0cZKzsvq7_0;
	wire w_dff_A_1Sn75JW53_2;
	wire w_dff_A_GzRYhqYM5_0;
	wire w_dff_A_3zW65Z0I5_0;
	wire w_dff_A_uDH37AKn4_0;
	wire w_dff_A_ubeslu0t4_2;
	wire w_dff_A_iFfqgdzM0_2;
	wire w_dff_A_BWR7BzNB9_2;
	wire w_dff_A_KXGCIGqG1_0;
	wire w_dff_A_zOSz57x41_1;
	wire w_dff_A_JBeus7uJ0_1;
	wire w_dff_A_7SAmofy49_1;
	wire w_dff_A_13G9R5bH5_1;
	wire w_dff_A_BAlsuDBm7_1;
	wire w_dff_A_jfWcgGkF8_0;
	wire w_dff_A_hTVxTAEg9_0;
	wire w_dff_A_zgFStbQ32_0;
	wire w_dff_A_DyEtyjAH1_1;
	wire w_dff_A_Y612Y2Iu4_1;
	wire w_dff_A_ccuwuU1G7_1;
	wire w_dff_A_fhN7CvxK0_0;
	wire w_dff_A_5tAOFhHm9_0;
	wire w_dff_A_wltsfTSv8_0;
	wire w_dff_A_vbCK6CD48_0;
	wire w_dff_B_TqeE9gwh0_1;
	wire w_dff_A_mVRfsAVZ1_1;
	wire w_dff_A_1Aer3cB25_1;
	wire w_dff_A_fsN6Eq2c3_0;
	wire w_dff_A_HmsmWUc61_0;
	wire w_dff_A_aqNT9f7j3_0;
	wire w_dff_A_xeeYnU4x7_1;
	wire w_dff_A_xhzSbQc21_1;
	wire w_dff_A_x85Fx5Bk9_1;
	wire w_dff_A_pNIHpZ1O9_1;
	wire w_dff_A_anOMJ07M0_0;
	wire w_dff_A_6Rvvtwnz2_0;
	wire w_dff_A_JSgvNSVS9_0;
	wire w_dff_A_9pmlRJzT8_2;
	wire w_dff_A_I7DHatgn6_2;
	wire w_dff_A_AWdAOljJ4_2;
	wire w_dff_A_bKPcwFxw3_2;
	wire w_dff_A_x2ult2f57_1;
	wire w_dff_A_BcTVejTc8_1;
	wire w_dff_A_h14eZX9o8_1;
	wire w_dff_A_MmzHCcUA0_1;
	wire w_dff_A_nuy12LkE4_2;
	wire w_dff_A_iinwmgc79_2;
	wire w_dff_B_E1mUxj7c0_1;
	wire w_dff_A_Wl9EksWk0_1;
	wire w_dff_A_g5LRjXiN1_0;
	wire w_dff_B_SP53AS286_2;
	wire w_dff_A_KlMvPo997_0;
	wire w_dff_A_qbX6Uqo06_0;
	wire w_dff_A_lAM3NFgD3_0;
	wire w_dff_A_TxZONEDW8_0;
	wire w_dff_A_5pCyFonK3_1;
	wire w_dff_A_VJNwAm6t4_0;
	wire w_dff_A_HhEUSmbu4_0;
	wire w_dff_A_ic6VYL2s1_0;
	wire w_dff_A_nxOb1jX52_1;
	wire w_dff_B_sT0q3vOJ5_0;
	wire w_dff_B_wdu0KqcM0_1;
	wire w_dff_A_AribFjuc2_0;
	wire w_dff_A_EJ8QD03f7_0;
	wire w_dff_A_v7wVNXzV8_0;
	wire w_dff_A_Esk9FLPn0_0;
	wire w_dff_A_DIxhcRxu7_1;
	wire w_dff_A_dfSf8Hys6_0;
	wire w_dff_A_ByuNwsEG1_0;
	wire w_dff_A_pllA2Bln3_2;
	wire w_dff_A_7RCLjyTf9_2;
	wire w_dff_A_oAMkPFud9_2;
	wire w_dff_A_WUSlaZ817_2;
	wire w_dff_B_bwUjs0ls1_2;
	wire w_dff_B_ZgjgcbpT5_2;
	wire w_dff_A_xsnjI4353_0;
	wire w_dff_A_FREIkpu59_0;
	wire w_dff_A_iaCFZwZi5_0;
	wire w_dff_A_uORXY95T9_0;
	wire w_dff_A_wQjxCHQ43_0;
	wire w_dff_A_oJvYPEnJ3_0;
	wire w_dff_A_PfzZNePP1_0;
	wire w_dff_B_HzC0cx2C7_1;
	wire w_dff_B_pauv6il10_1;
	wire w_dff_A_MjqUp2IV7_0;
	wire w_dff_A_eLh1wXtP2_0;
	wire w_dff_A_HOvEmfsF0_0;
	wire w_dff_A_rT4nJnsx9_1;
	wire w_dff_A_H6Myhpd09_1;
	wire w_dff_A_Mc4qclDQ7_0;
	wire w_dff_A_VcdHeGSe5_0;
	wire w_dff_A_QS6hAFmE7_0;
	wire w_dff_A_PsGS15dS5_1;
	wire w_dff_A_FROdvvJx1_0;
	wire w_dff_A_OEyQfNX14_0;
	wire w_dff_A_llzU1GyE4_0;
	wire w_dff_A_EcODS1TM6_0;
	wire w_dff_A_TfyK3HW66_1;
	wire w_dff_A_B60DKuWp4_1;
	wire w_dff_A_l4Toek0g7_1;
	wire w_dff_A_IbB9Taz62_2;
	wire w_dff_A_irs9bHBr5_2;
	wire w_dff_A_DtA0yE6o6_1;
	wire w_dff_A_udrKFxna6_0;
	wire w_dff_A_3xRNxzVm0_0;
	wire w_dff_A_wFYZV4pb7_1;
	wire w_dff_A_zzM06KLE7_1;
	wire w_dff_A_e6fQA4aB6_0;
	wire w_dff_A_JnrTIHvl0_0;
	wire w_dff_A_8GO6iolU1_0;
	wire w_dff_A_KPDjnYZZ5_1;
	wire w_dff_A_G3VZeg0G8_1;
	wire w_dff_A_RndfyFv52_1;
	wire w_dff_A_U3y76x5D0_1;
	wire w_dff_A_vc88hoFt9_0;
	wire w_dff_A_m64AZkit3_0;
	wire w_dff_A_REC5uBRg6_0;
	wire w_dff_A_32enTWEY8_1;
	wire w_dff_A_M3EiS25C9_1;
	wire w_dff_A_zlfUFNxN7_1;
	wire w_dff_A_EhSyXoq93_2;
	wire w_dff_B_suPl964r6_1;
	wire w_dff_A_8yi5hHaE5_0;
	wire w_dff_A_26xsE9xa2_0;
	wire w_dff_A_lt9IHk169_0;
	wire w_dff_A_4CpzGqHi7_0;
	wire w_dff_A_mWcYaPyM8_0;
	wire w_dff_A_3FKnpT776_0;
	wire w_dff_A_bGE5KNDJ7_0;
	wire w_dff_A_2pTMC7fh9_1;
	wire w_dff_A_2nITGxT72_2;
	wire w_dff_A_I4W3GC0P2_2;
	wire w_dff_A_bN7ldxU20_2;
	wire w_dff_A_LPUcDJBS2_2;
	wire w_dff_A_sMpOPvSM9_2;
	wire w_dff_A_4Il5uod24_2;
	wire w_dff_A_mJWlEdhi3_2;
	wire w_dff_A_qayL26XG4_0;
	wire w_dff_A_wAzwG5NF6_0;
	wire w_dff_A_eeXcb0LK1_0;
	wire w_dff_A_7rw9GJCL1_0;
	wire w_dff_A_tkwBkKGg1_0;
	wire w_dff_A_MToV3uQi0_0;
	wire w_dff_A_dVvesc1C1_0;
	wire w_dff_A_Ac1t2Z0B9_1;
	wire w_dff_A_F0YiJfRp5_1;
	wire w_dff_A_wCBPIBH18_1;
	wire w_dff_A_4kFVSjYh8_1;
	wire w_dff_A_0M59mrjU1_1;
	wire w_dff_A_hz48tvZj2_0;
	wire w_dff_A_PbvQEbvw8_0;
	wire w_dff_B_6KcOzGgC9_2;
	wire w_dff_A_mVCFVMyS7_0;
	wire w_dff_A_uzO5xhyl4_2;
	wire w_dff_A_6k8eSR7l3_1;
	wire w_dff_A_PWuV5Axc5_0;
	wire w_dff_A_VCFA39Bw3_1;
	wire w_dff_A_ZTcFboHJ9_0;
	wire w_dff_A_JFjoZqRm7_2;
	wire w_dff_B_T99fJxNq5_3;
	wire w_dff_B_HskBRdxc1_3;
	wire w_dff_B_uYtT4eQu5_3;
	wire w_dff_B_vNKcW1C49_3;
	wire w_dff_B_kIJv506o1_3;
	wire w_dff_A_xCs0uLOj3_0;
	wire w_dff_A_XKSjJ5hH1_0;
	wire w_dff_A_e7tTGEca3_0;
	wire w_dff_A_DE7AwlLp0_0;
	wire w_dff_A_Ks2d8K442_0;
	wire w_dff_A_Fqlu81ZI1_0;
	wire w_dff_A_suGe9WPO6_0;
	wire w_dff_A_DLUYiEM47_1;
	wire w_dff_A_hJM2TBQB1_1;
	wire w_dff_A_q7JbCo8W6_1;
	wire w_dff_A_QzUOOnDj6_1;
	wire w_dff_A_q1vMp6Xt8_1;
	wire w_dff_A_7k4l7qt24_1;
	wire w_dff_A_J1ih0qTn6_1;
	wire w_dff_A_lF4JxzxQ2_0;
	wire w_dff_A_4SFMbZqQ6_0;
	wire w_dff_A_ZUQtZJlv5_0;
	wire w_dff_A_WJoMVyUr7_0;
	wire w_dff_A_NS9sNu3e4_0;
	wire w_dff_A_f208jTEV9_0;
	wire w_dff_A_Dr0dLoVk1_0;
	wire w_dff_B_CTKC3q9z3_0;
	wire w_dff_A_BhaIHiIi3_1;
	wire w_dff_A_NTvaMBSR8_0;
	wire w_dff_A_bYTrrIyV4_0;
	wire w_dff_A_ObhdSrtI1_2;
	wire w_dff_A_tijpbY7D0_0;
	wire w_dff_A_65zy7shZ0_0;
	wire w_dff_A_UAB7M2MC5_2;
	wire w_dff_A_bDTE1pCU5_2;
	wire w_dff_A_VyS28cge1_2;
	wire w_dff_A_HZd2GatY8_2;
	wire w_dff_A_tnr0FCP54_0;
	wire w_dff_A_J9rY81dQ7_1;
	wire w_dff_A_gHYXEe3V2_1;
	wire w_dff_A_sasnW2SN5_1;
	wire w_dff_A_ffrbgNc21_1;
	wire w_dff_A_6luVzNKG7_2;
	wire w_dff_A_mnmkF3jC1_2;
	wire w_dff_A_lqG2rG0X8_2;
	wire w_dff_A_Ilu1AmxG0_2;
	wire w_dff_A_h6lmthOs1_2;
	wire w_dff_A_NY5FChnJ6_2;
	wire w_dff_A_dmDIpHXg8_2;
	wire w_dff_A_O1jHvSWP8_2;
	wire w_dff_A_31bST4RG1_1;
	wire w_dff_A_pd9Unxrj0_1;
	wire w_dff_A_FTkE7pQJ2_1;
	wire w_dff_A_tsI1dVCL6_2;
	wire w_dff_A_fWt6MUaE7_2;
	wire w_dff_A_pw1EcozM1_2;
	wire w_dff_A_W52wfV0H7_0;
	wire w_dff_A_vIXjKMLs5_0;
	wire w_dff_A_GViDkCJD7_0;
	wire w_dff_A_AZl59P653_1;
	wire w_dff_A_swqtA9sL9_0;
	wire w_dff_A_001aC8LN9_0;
	wire w_dff_A_ZsQLVsqs3_2;
	wire w_dff_A_oGYHcEpi4_2;
	wire w_dff_A_c7vPv7cN1_2;
	wire w_dff_A_3AMTUf409_0;
	wire w_dff_A_vI1MDHPb8_0;
	wire w_dff_A_yTyBwOZq2_0;
	wire w_dff_A_w42ZATqo8_1;
	wire w_dff_A_jPwCkNEH8_1;
	wire w_dff_A_Vmkku8fN4_2;
	wire w_dff_A_F7j5jKl69_2;
	wire w_dff_A_VSlHQ9P36_2;
	wire w_dff_A_Madlfysn3_1;
	wire w_dff_A_8wMjJHIG7_0;
	wire w_dff_A_PJNWczpa1_1;
	wire w_dff_A_0corOKVj7_0;
	wire w_dff_A_DxGsPXO13_2;
	wire w_dff_A_0ztcYfpW6_2;
	wire w_dff_A_h2tkC4do5_2;
	wire w_dff_A_aD3bYPsb3_2;
	wire w_dff_A_si08ltWt9_2;
	wire w_dff_A_1cQcbg208_1;
	wire w_dff_A_1hQTGFhM4_0;
	wire w_dff_A_Ekx2lsgO5_2;
	wire w_dff_A_nOj7S6af6_0;
	wire w_dff_B_dhtP6ddm7_2;
	wire w_dff_B_mCDef9Oe5_2;
	wire w_dff_A_iGp4QjM17_0;
	wire w_dff_A_VF4oUAvq4_0;
	wire w_dff_A_uB9kAt2B0_0;
	wire w_dff_A_Afu5Kpga3_2;
	wire w_dff_A_MERfyLJc9_2;
	wire w_dff_A_6TTriCEI5_2;
	wire w_dff_A_9oPM0F8E6_2;
	wire w_dff_A_b8Aotwq21_1;
	wire w_dff_A_ALhdn8qc6_1;
	wire w_dff_A_C9em7tj81_1;
	wire w_dff_A_8qEqV5IG1_2;
	wire w_dff_A_fxc072rn5_0;
	wire w_dff_A_uZz1fQBT7_1;
	wire w_dff_A_4Ouj8ThX9_0;
	wire w_dff_B_2Q9ieLS33_0;
	wire w_dff_A_PoliPYxD4_0;
	wire w_dff_A_YQsvCYYk7_0;
	wire w_dff_A_coUzNFjU0_0;
	wire w_dff_A_0eV7BkGz8_2;
	wire w_dff_A_5BzSVzfU8_2;
	wire w_dff_A_UAPhG3Vn9_0;
	wire w_dff_B_WYnzbP1T3_0;
	wire w_dff_A_vtqn6Ngn9_2;
	wire w_dff_A_NG8iqZFU6_0;
	wire w_dff_A_FoBBaqwL2_1;
	wire w_dff_A_hTYt0Sei3_0;
	wire w_dff_A_USztoXLK7_2;
	wire w_dff_A_Xy8ZZeI59_2;
	wire w_dff_A_pIExNAhw0_2;
	wire w_dff_A_ZxELQh9I5_0;
	wire w_dff_A_CO9EWdaC6_0;
	wire w_dff_A_GFDKQ38K5_1;
	wire w_dff_A_tEVBWGW62_1;
	wire w_dff_A_qrTS6Gwh7_1;
	wire w_dff_A_yQTxWFRA1_1;
	wire w_dff_A_bV0VerXU7_2;
	wire w_dff_A_TRFGqDUJ8_2;
	wire w_dff_A_UYUfUEAd4_2;
	wire w_dff_A_hEPKzEzv3_0;
	wire w_dff_A_KVIzA3Ct9_1;
	wire w_dff_A_LFyYcmB27_0;
	wire w_dff_A_0Dr2K6jL4_0;
	wire w_dff_A_rZmdm5qG0_1;
	wire w_dff_A_c67gaj6g8_1;
	wire w_dff_B_GRNElknY8_1;
	wire w_dff_A_9ww3VlH63_0;
	wire w_dff_A_GHAbKBh17_0;
	wire w_dff_A_DQKieqpc6_2;
	wire w_dff_A_tcKA3BhQ5_2;
	wire w_dff_A_ydHFQ62C3_1;
	wire w_dff_A_WHghHJm77_1;
	wire w_dff_A_raVhjKGT5_1;
	wire w_dff_A_ktoydHJt5_2;
	wire w_dff_A_Ar3Xl1TE6_2;
	wire w_dff_A_pzus6SVP7_2;
	wire w_dff_A_fglkHkid8_1;
	wire w_dff_A_UpmNlgzu2_1;
	wire w_dff_A_6sEZr79Z9_1;
	wire w_dff_A_JUzIhdWg1_2;
	wire w_dff_A_TBnhXvjT5_0;
	wire w_dff_A_303rdBsU8_0;
	wire w_dff_A_hukRPu1H1_1;
	wire w_dff_A_f3QAmBdV4_1;
	wire w_dff_A_XCrtveZf8_1;
	wire w_dff_A_pJc5Nymd0_1;
	wire w_dff_A_zPI9h0pG0_2;
	wire w_dff_A_9N91VHxD5_2;
	wire w_dff_A_Mlfa3Jcp5_2;
	wire w_dff_A_Z0cjFDHq7_0;
	wire w_dff_A_oHNNeNEI2_0;
	wire w_dff_A_06D0wKbJ5_1;
	wire w_dff_A_6nObsZ5H3_1;
	wire w_dff_A_lJ3aMjpq8_1;
	wire w_dff_A_iaPOG52y2_1;
	wire w_dff_A_4o0p8slk3_2;
	wire w_dff_A_bj6XxWiH2_2;
	wire w_dff_A_ppGTzq2G7_2;
	wire w_dff_A_upYG8lUr4_2;
	wire w_dff_A_rYRdCdk93_1;
	wire w_dff_A_kDyzheB88_1;
	wire w_dff_A_eRcHLr176_2;
	wire w_dff_A_EWytyrHp6_2;
	wire w_dff_A_FJazkNfU9_1;
	wire w_dff_A_bZl15ToZ9_1;
	wire w_dff_A_sgKsKajD0_0;
	wire w_dff_A_eheZoAGo8_1;
	wire w_dff_A_HgYY2dUb4_2;
	wire w_dff_A_AH0KJFDU0_2;
	wire w_dff_A_a3mhyjEm2_2;
	wire w_dff_A_inB6gsfz0_2;
	wire w_dff_A_ogfXx8KF4_2;
	wire w_dff_A_a59X2VON1_2;
	wire w_dff_A_8qgATIe62_2;
	wire w_dff_A_KPWEOBb32_0;
	wire w_dff_A_slPEs5cW2_1;
	wire w_dff_A_PQfOk9nx5_2;
	wire w_dff_A_pLbnh99t5_1;
	wire w_dff_A_4bLfR68l3_2;
	wire w_dff_A_0eRuYOQO3_2;
	wire w_dff_A_3nvoBC4Z2_0;
	wire w_dff_A_O3PSfUPA3_2;
	wire w_dff_A_iAdXw7Hj8_0;
	wire w_dff_A_YK0gGx2Z1_1;
	wire w_dff_A_EA9FYDxy9_1;
	wire w_dff_A_l0bbccIh9_1;
	wire w_dff_A_quvSuv8u5_1;
	wire w_dff_A_xsBHwhZ30_1;
	wire w_dff_A_m8wv256D9_1;
	wire w_dff_A_UBBdH3Pi7_2;
	wire w_dff_A_awll7jxE2_2;
	wire w_dff_A_PpQpP64P8_2;
	wire w_dff_A_VsF606or9_2;
	wire w_dff_A_9tTkdQcL6_2;
	wire w_dff_A_fLtmlSke3_2;
	wire w_dff_A_SDNStn4c4_0;
	wire w_dff_A_GM2LTRIx2_0;
	wire w_dff_A_sLGr2W334_0;
	wire w_dff_A_hdZFUim10_0;
	wire w_dff_A_6ZgD6zws4_0;
	wire w_dff_A_Hn2rZI4c7_0;
	wire w_dff_A_G6PyO8im8_0;
	wire w_dff_A_BTJJSqX32_1;
	wire w_dff_A_76qXpSFo4_1;
	wire w_dff_A_SXKzKZXg9_1;
	wire w_dff_A_gcq7ZLJ48_1;
	wire w_dff_A_5YOTw2ai0_1;
	wire w_dff_A_cNWazVGD3_1;
	wire w_dff_A_73xXv1qJ4_1;
	wire w_dff_A_jZlf7qoN7_2;
	wire w_dff_A_FLMG89st7_2;
	wire w_dff_A_6mrcnqob9_2;
	wire w_dff_A_myXmhWVs2_2;
	wire w_dff_A_PWB9Dwhw3_2;
	wire w_dff_A_YxIiNnCT8_2;
	wire w_dff_A_QuWBZkPP5_2;
	wire w_dff_A_jDDyjmOM9_2;
	wire w_dff_A_oCeIctIc4_0;
	wire w_dff_A_yTGtcVRg0_0;
	wire w_dff_A_8JwgpaaC9_0;
	wire w_dff_A_bPrcsCRS4_0;
	wire w_dff_A_XEUnkOtK1_0;
	wire w_dff_A_04jcxYzU7_0;
	wire w_dff_A_ou87bcHz4_0;
	wire w_dff_A_qtcryspU0_0;
	wire w_dff_A_ja7F6qH94_0;
	wire w_dff_A_FE7Sq7Tl2_0;
	wire w_dff_A_Vdc5lXXl2_0;
	wire w_dff_A_0TUAKMoS1_0;
	wire w_dff_A_sO0ezfUK2_0;
	wire w_dff_A_Py8YTI9G5_0;
	wire w_dff_A_XHUR7MiC5_0;
	wire w_dff_A_W46RsyYx0_0;
	wire w_dff_A_NbxblaA19_0;
	wire w_dff_A_MQoacw8Q9_0;
	wire w_dff_A_LAqLvMI30_0;
	wire w_dff_A_mkE7Z8ts0_0;
	wire w_dff_A_46Ybfo041_0;
	wire w_dff_A_HGzp22941_0;
	wire w_dff_A_PFGQIOju3_0;
	wire w_dff_A_ihUofMly6_0;
	wire w_dff_A_b4JJi3Xo9_1;
	wire w_dff_A_3D80Yf1i6_0;
	wire w_dff_A_5nhhep6d9_0;
	wire w_dff_A_0thdKQix0_0;
	wire w_dff_A_4ge9LgrV4_0;
	wire w_dff_A_wKJWkuGj9_0;
	wire w_dff_A_aI3kkDP84_0;
	wire w_dff_A_XA72lHkS1_0;
	wire w_dff_A_jsIA8eKB8_0;
	wire w_dff_A_c60NlIbj0_0;
	wire w_dff_A_2ewcdiOT9_0;
	wire w_dff_A_2VzzZEfu5_0;
	wire w_dff_A_XSxjnDbD9_0;
	wire w_dff_A_mzsI8NCp0_0;
	wire w_dff_A_uxR2QE8v0_0;
	wire w_dff_A_A9gopoxK0_0;
	wire w_dff_A_mHTJaAdx4_0;
	wire w_dff_A_GCl3sPpe3_0;
	wire w_dff_A_Hl1KhlD93_0;
	wire w_dff_A_k5zRfPFm4_0;
	wire w_dff_A_JyflBbLh1_0;
	wire w_dff_A_oyZYblEz3_0;
	wire w_dff_A_gWKpw2w06_0;
	wire w_dff_A_yunia8tt0_0;
	wire w_dff_A_yu2mnwg27_2;
	wire w_dff_A_bPEi8vwn8_0;
	wire w_dff_A_lGzCx7Df2_0;
	wire w_dff_A_mCSCtIhU9_0;
	wire w_dff_A_sMl3qcMf6_0;
	wire w_dff_A_ypir7DjH3_0;
	wire w_dff_A_rPmcsS9X7_0;
	wire w_dff_A_eFcD9XJe2_0;
	wire w_dff_A_fLrCvENM3_0;
	wire w_dff_A_gqOq2OKz3_0;
	wire w_dff_A_LSXYNV9I7_0;
	wire w_dff_A_GgQZkZ8N0_0;
	wire w_dff_A_MUil1Pu22_0;
	wire w_dff_A_F7PTQD1p0_0;
	wire w_dff_A_LCwPXFQN8_0;
	wire w_dff_A_igeNho1x0_0;
	wire w_dff_A_2j63eibE7_0;
	wire w_dff_A_6z13bnug1_0;
	wire w_dff_A_h1nEpwY53_0;
	wire w_dff_A_CLRBlX9P2_0;
	wire w_dff_A_hyFJq4Tp4_0;
	wire w_dff_A_KxktjB0M1_2;
	wire w_dff_A_ETfMRraI8_0;
	wire w_dff_A_i5LiCjT30_0;
	wire w_dff_A_b7GGSp3J5_0;
	wire w_dff_A_YLwcEg3v9_0;
	wire w_dff_A_S8gd0K6y9_0;
	wire w_dff_A_AJsGT4HC7_0;
	wire w_dff_A_M1uryMSr8_0;
	wire w_dff_A_kbFLxLLY1_0;
	wire w_dff_A_7xcccwWZ0_0;
	wire w_dff_A_PSGaGukk8_0;
	wire w_dff_A_Aw3cQnog9_0;
	wire w_dff_A_9JTme08A5_0;
	wire w_dff_A_JxT0K3Sj4_0;
	wire w_dff_A_XwkblzX26_0;
	wire w_dff_A_PrdI3O528_0;
	wire w_dff_A_GJc1JsfS1_0;
	wire w_dff_A_f7inSK2C2_0;
	wire w_dff_A_oglXmj6O5_0;
	wire w_dff_A_nyPwmjWf0_0;
	wire w_dff_A_dFuDFUHC4_0;
	wire w_dff_A_OcB7E4FS6_0;
	wire w_dff_A_fOdpVXOa1_0;
	wire w_dff_A_KNTDztRT6_0;
	wire w_dff_A_hm8XpUoB1_2;
	wire w_dff_A_N4XF6Hnn0_0;
	wire w_dff_A_u2pQx0fr2_0;
	wire w_dff_A_f4p5mze87_0;
	wire w_dff_A_V7ZJnNfe1_0;
	wire w_dff_A_cBFbio7O4_0;
	wire w_dff_A_vXZQ5h5j9_0;
	wire w_dff_A_2S85BXrz9_0;
	wire w_dff_A_egVfUnC77_0;
	wire w_dff_A_mgfaHL9H3_0;
	wire w_dff_A_TOneLI254_0;
	wire w_dff_A_k1fWSuVW4_0;
	wire w_dff_A_o6u0Nn5F9_0;
	wire w_dff_A_xyL8Gekh9_0;
	wire w_dff_A_Il4rDvRK9_0;
	wire w_dff_A_bl42ncSb2_0;
	wire w_dff_A_eAyqwCzZ6_0;
	wire w_dff_A_OC9iKQH58_0;
	wire w_dff_A_2w8vXaEC5_0;
	wire w_dff_A_hqzYHSbg0_0;
	wire w_dff_A_VK5lhS117_0;
	wire w_dff_A_kqRTBoj71_0;
	wire w_dff_A_dnWPRKXl7_0;
	wire w_dff_A_XBN2pRht0_0;
	wire w_dff_A_Fo7AjoZB3_2;
	wire w_dff_A_3SRJIUlD6_0;
	wire w_dff_A_d1Py6wvc5_0;
	wire w_dff_A_qyS5Wz0A7_0;
	wire w_dff_A_XnUb4Zlr3_0;
	wire w_dff_A_issZT9NH3_0;
	wire w_dff_A_CHVGcIuR9_0;
	wire w_dff_A_lMKux7055_0;
	wire w_dff_A_UU5ENAX71_0;
	wire w_dff_A_cAUmK5Mm7_0;
	wire w_dff_A_zrjxHRTb1_0;
	wire w_dff_A_vj5vTeuW9_0;
	wire w_dff_A_rPyJpGr71_0;
	wire w_dff_A_swsvL5td8_0;
	wire w_dff_A_yKE6Pi2p6_2;
	wire w_dff_A_ILl5k9cI5_0;
	wire w_dff_A_VOcmU1MJ3_0;
	wire w_dff_A_NE5UXxOC0_0;
	wire w_dff_A_LPvpTHiz2_0;
	wire w_dff_A_Q5jFwPwD3_0;
	wire w_dff_A_ohcL0so56_0;
	wire w_dff_A_EpvJVHbi5_0;
	wire w_dff_A_Hsa47J9Y2_0;
	wire w_dff_A_On5sCEYo3_0;
	wire w_dff_A_Y7PXSUVf4_0;
	wire w_dff_A_SyK2xPPD8_0;
	wire w_dff_A_TMIQp7yB0_2;
	wire w_dff_A_40r01Umj8_0;
	wire w_dff_A_sZTAlPqr8_0;
	wire w_dff_A_dC2RTqVH5_0;
	wire w_dff_A_oYxdiuPb2_0;
	wire w_dff_A_bUqrFaCj4_0;
	wire w_dff_A_IBhUu7Qm6_0;
	wire w_dff_A_wzJh5yps6_0;
	wire w_dff_A_kYLZHSdZ3_0;
	wire w_dff_A_hwO46wRc7_0;
	wire w_dff_A_E7jguRXM1_0;
	wire w_dff_A_0WVEvPGS5_2;
	wire w_dff_A_bjZscRO61_0;
	wire w_dff_A_ipYufpMg8_0;
	wire w_dff_A_nfIuEa7O8_0;
	wire w_dff_A_WIolRQIE1_0;
	wire w_dff_A_04fPKSR12_0;
	wire w_dff_A_hblpjV0x7_0;
	wire w_dff_A_iCJiOi5u8_0;
	wire w_dff_A_j3MvBzGw5_0;
	wire w_dff_A_x0zfNS5s1_0;
	wire w_dff_A_eJhMTvLA1_0;
	wire w_dff_A_JvhgudXb7_2;
	wire w_dff_A_7jU79r5T3_0;
	wire w_dff_A_zJMLiDnG9_0;
	wire w_dff_A_fgn35j2M0_0;
	wire w_dff_A_LtUMQUBu0_0;
	wire w_dff_A_hI41J0ac3_0;
	wire w_dff_A_KTddD5ff1_0;
	wire w_dff_A_idLnCTGo6_0;
	wire w_dff_A_o6sNFGwq7_0;
	wire w_dff_A_yQqCGAVL5_0;
	wire w_dff_A_SdWRPurT6_0;
	wire w_dff_A_MK7puvqH4_1;
	wire w_dff_A_T3sTSkls0_0;
	wire w_dff_A_8GJ6RkPC8_0;
	wire w_dff_A_pZuEXSwI3_0;
	wire w_dff_A_Dz2LoSbI3_0;
	wire w_dff_A_qeYaqAiR2_0;
	wire w_dff_A_KfbbFbyt7_0;
	wire w_dff_A_dwFfx8zJ1_0;
	wire w_dff_A_OjXgsc6F9_2;
	wire w_dff_A_kItvCpdm3_0;
	wire w_dff_A_NuQSjE8t0_0;
	wire w_dff_A_VkvuCOeX2_0;
	wire w_dff_A_1OsQOe6J0_0;
	wire w_dff_A_gMbPIbhZ9_2;
	wire w_dff_A_pePACUYr0_0;
	wire w_dff_A_J8CYK0z98_0;
	wire w_dff_A_lh9HrNeF8_0;
	wire w_dff_A_C6v6yx9W8_0;
	wire w_dff_A_6AG3SgwF9_1;
	wire w_dff_A_1wa6scRT4_0;
	wire w_dff_A_EZIh7BOM0_0;
	wire w_dff_A_QDHzbLAS4_0;
	wire w_dff_A_7B7YrEgs1_0;
	wire w_dff_A_lGrXPsPf5_0;
	wire w_dff_A_63rnxrt66_0;
	wire w_dff_A_zmyyTuog8_1;
	wire w_dff_A_h8B1FVzK0_0;
	wire w_dff_A_OSUarnG38_0;
	wire w_dff_A_PDseqAHC6_0;
	wire w_dff_A_Ev65jC9w8_0;
	wire w_dff_A_aUQ6yJFl6_0;
	wire w_dff_A_ywGiTRig5_1;
	wire w_dff_A_hCj3951Q9_0;
	wire w_dff_A_Y34FfsEq6_0;
	wire w_dff_A_KbweROGQ1_0;
	wire w_dff_A_RAOIGzOa2_0;
	wire w_dff_A_ULxsSlua0_1;
	wire w_dff_A_CB5hT0D90_0;
	wire w_dff_A_VKLgk1X27_0;
	wire w_dff_A_BEk3hAnd8_1;
	wire w_dff_A_OYV2J0ds3_0;
	wire w_dff_A_Sp6VE8id9_0;
	wire w_dff_A_FoPg98jD2_0;
	wire w_dff_A_UJV9lTxp4_0;
	wire w_dff_A_jCISqWYT9_1;
	wire w_dff_A_ysFzlHig4_2;
	jnot g0000(.din(w_G77_5[1]),.dout(n72),.clk(gclk));
	jnot g0001(.din(w_G50_5[2]),.dout(n73),.clk(gclk));
	jnot g0002(.din(w_G58_5[1]),.dout(n74),.clk(gclk));
	jnot g0003(.din(w_G68_5[1]),.dout(n75),.clk(gclk));
	jand g0004(.dina(w_n75_1[1]),.dinb(w_n74_1[1]),.dout(n76),.clk(gclk));
	jand g0005(.dina(w_n76_0[1]),.dinb(w_n73_2[2]),.dout(n77),.clk(gclk));
	jand g0006(.dina(w_n77_0[1]),.dinb(w_n72_1[1]),.dout(w_dff_A_jDDyjmOM9_2),.clk(gclk));
	jnot g0007(.din(w_G97_5[1]),.dout(n79),.clk(gclk));
	jnot g0008(.din(w_G107_5[1]),.dout(n80),.clk(gclk));
	jand g0009(.dina(w_n80_1[1]),.dinb(w_n79_0[2]),.dout(n81),.clk(gclk));
	jnot g0010(.din(w_n81_0[2]),.dout(n82),.clk(gclk));
	jand g0011(.dina(n82),.dinb(w_G87_3[2]),.dout(n83),.clk(gclk));
	jnot g0012(.din(n83),.dout(G355_fa_),.clk(gclk));
	jand g0013(.dina(w_G20_7[1]),.dinb(w_G1_3[1]),.dout(n85),.clk(gclk));
	jnot g0014(.din(w_G226_1[1]),.dout(n86),.clk(gclk));
	jor g0015(.dina(w_n86_0[1]),.dinb(w_n73_2[1]),.dout(n87),.clk(gclk));
	jnot g0016(.din(w_G264_1[1]),.dout(n88),.clk(gclk));
	jor g0017(.dina(w_n88_1[1]),.dinb(w_n80_1[0]),.dout(n89),.clk(gclk));
	jand g0018(.dina(n89),.dinb(n87),.dout(n90),.clk(gclk));
	jnot g0019(.din(w_G257_1[2]),.dout(n91),.clk(gclk));
	jor g0020(.dina(w_n91_1[2]),.dinb(w_n79_0[1]),.dout(n92),.clk(gclk));
	jnot g0021(.din(w_G238_1[2]),.dout(n93),.clk(gclk));
	jor g0022(.dina(w_n93_0[1]),.dinb(w_n75_1[0]),.dout(n94),.clk(gclk));
	jand g0023(.dina(n94),.dinb(n92),.dout(n95),.clk(gclk));
	jand g0024(.dina(n95),.dinb(n90),.dout(n96),.clk(gclk));
	jnot g0025(.din(w_G87_3[1]),.dout(n97),.clk(gclk));
	jnot g0026(.din(w_G250_0[2]),.dout(n98),.clk(gclk));
	jor g0027(.dina(w_n98_2[1]),.dinb(w_n97_2[1]),.dout(n99),.clk(gclk));
	jnot g0028(.din(w_G232_1[2]),.dout(n100),.clk(gclk));
	jor g0029(.dina(n100),.dinb(w_n74_1[0]),.dout(n101),.clk(gclk));
	jand g0030(.dina(n101),.dinb(n99),.dout(n102),.clk(gclk));
	jnot g0031(.din(w_G244_1[2]),.dout(n103),.clk(gclk));
	jor g0032(.dina(w_n103_0[2]),.dinb(w_n72_1[0]),.dout(n104),.clk(gclk));
	jnot g0033(.din(w_G116_4[2]),.dout(n105),.clk(gclk));
	jnot g0034(.din(w_G270_0[2]),.dout(n106),.clk(gclk));
	jor g0035(.dina(w_n106_0[1]),.dinb(w_n105_2[1]),.dout(n107),.clk(gclk));
	jand g0036(.dina(n107),.dinb(n104),.dout(n108),.clk(gclk));
	jand g0037(.dina(n108),.dinb(n102),.dout(n109),.clk(gclk));
	jand g0038(.dina(n109),.dinb(n96),.dout(n110),.clk(gclk));
	jor g0039(.dina(n110),.dinb(w_n85_0[2]),.dout(n111),.clk(gclk));
	jnot g0040(.din(w_G20_7[0]),.dout(n112),.clk(gclk));
	jnot g0041(.din(w_G1_3[0]),.dout(n113),.clk(gclk));
	jnot g0042(.din(w_G13_1[1]),.dout(n114),.clk(gclk));
	jor g0043(.dina(w_n114_1[2]),.dinb(w_n113_3[1]),.dout(n115),.clk(gclk));
	jor g0044(.dina(w_n115_1[1]),.dinb(w_n112_5[2]),.dout(n116),.clk(gclk));
	jnot g0045(.din(w_n76_0[0]),.dout(n117),.clk(gclk));
	jand g0046(.dina(n117),.dinb(w_G50_5[1]),.dout(n118),.clk(gclk));
	jnot g0047(.din(w_n118_0[2]),.dout(n119),.clk(gclk));
	jor g0048(.dina(n119),.dinb(w_n116_0[1]),.dout(n120),.clk(gclk));
	jand g0049(.dina(w_n114_1[1]),.dinb(w_G1_2[2]),.dout(n121),.clk(gclk));
	jand g0050(.dina(w_n121_0[2]),.dinb(w_G20_6[2]),.dout(n122),.clk(gclk));
	jnot g0051(.din(w_n122_1[1]),.dout(n123),.clk(gclk));
	jand g0052(.dina(w_n88_1[0]),.dinb(w_n91_1[1]),.dout(n124),.clk(gclk));
	jor g0053(.dina(n124),.dinb(w_n98_2[0]),.dout(n125),.clk(gclk));
	jor g0054(.dina(w_dff_B_XAQHaUNc9_0),.dinb(w_n123_1[2]),.dout(n126),.clk(gclk));
	jand g0055(.dina(w_dff_B_RKYEFx1F2_0),.dinb(n120),.dout(n127),.clk(gclk));
	jand g0056(.dina(n127),.dinb(w_dff_B_ZbIvEJMZ1_1),.dout(w_dff_A_yu2mnwg27_2),.clk(gclk));
	jxor g0057(.dina(w_G270_0[1]),.dinb(w_G264_1[0]),.dout(n129),.clk(gclk));
	jxor g0058(.dina(w_G257_1[1]),.dinb(w_n98_1[2]),.dout(n130),.clk(gclk));
	jxor g0059(.dina(n130),.dinb(w_dff_B_dBwvH5b50_1),.dout(n131),.clk(gclk));
	jnot g0060(.din(w_n131_0[1]),.dout(n132),.clk(gclk));
	jxor g0061(.dina(w_G244_1[1]),.dinb(w_G238_1[1]),.dout(n133),.clk(gclk));
	jxor g0062(.dina(w_G232_1[1]),.dinb(w_n86_0[0]),.dout(n134),.clk(gclk));
	jxor g0063(.dina(n134),.dinb(w_dff_B_hpJU5pAe0_1),.dout(n135),.clk(gclk));
	jxor g0064(.dina(w_n135_0[1]),.dinb(n132),.dout(w_dff_A_KxktjB0M1_2),.clk(gclk));
	jxor g0065(.dina(w_G68_5[0]),.dinb(w_G58_5[0]),.dout(n137),.clk(gclk));
	jnot g0066(.din(w_n137_0[2]),.dout(n138),.clk(gclk));
	jxor g0067(.dina(w_G77_5[0]),.dinb(w_G50_5[0]),.dout(n139),.clk(gclk));
	jxor g0068(.dina(w_dff_B_aPhNAm609_0),.dinb(n138),.dout(n140),.clk(gclk));
	jnot g0069(.din(w_n140_0[1]),.dout(n141),.clk(gclk));
	jxor g0070(.dina(w_G116_4[1]),.dinb(w_G107_5[0]),.dout(n142),.clk(gclk));
	jxor g0071(.dina(w_G97_5[0]),.dinb(w_n97_2[0]),.dout(n143),.clk(gclk));
	jxor g0072(.dina(n143),.dinb(w_dff_B_MvjVfA9W0_1),.dout(n144),.clk(gclk));
	jxor g0073(.dina(w_n144_0[1]),.dinb(n141),.dout(w_dff_A_hm8XpUoB1_2),.clk(gclk));
	jnot g0074(.din(w_G169_1[1]),.dout(n146),.clk(gclk));
	jand g0075(.dina(w_G13_1[0]),.dinb(w_G1_2[1]),.dout(n147),.clk(gclk));
	jnot g0076(.din(w_G33_11[2]),.dout(n148),.clk(gclk));
	jnot g0077(.din(w_G41_1[1]),.dout(n149),.clk(gclk));
	jor g0078(.dina(w_n149_2[1]),.dinb(w_n148_9[2]),.dout(n150),.clk(gclk));
	jand g0079(.dina(n150),.dinb(w_n147_0[2]),.dout(n151),.clk(gclk));
	jand g0080(.dina(w_G1698_0[2]),.dinb(w_n148_9[1]),.dout(n152),.clk(gclk));
	jand g0081(.dina(w_n152_3[1]),.dinb(w_G244_1[0]),.dout(n153),.clk(gclk));
	jnot g0082(.din(w_G1698_0[1]),.dout(n154),.clk(gclk));
	jand g0083(.dina(w_n154_0[1]),.dinb(w_n148_9[0]),.dout(n155),.clk(gclk));
	jand g0084(.dina(w_n155_3[1]),.dinb(w_G238_1[0]),.dout(n156),.clk(gclk));
	jand g0085(.dina(w_G116_4[0]),.dinb(w_G33_11[1]),.dout(n157),.clk(gclk));
	jor g0086(.dina(w_n157_0[2]),.dinb(n156),.dout(n158),.clk(gclk));
	jor g0087(.dina(n158),.dinb(w_dff_B_GRNElknY8_1),.dout(n159),.clk(gclk));
	jand g0088(.dina(n159),.dinb(w_n151_4[2]),.dout(n160),.clk(gclk));
	jnot g0089(.din(w_G45_1[2]),.dout(n161),.clk(gclk));
	jor g0090(.dina(w_n161_1[1]),.dinb(w_G1_2[0]),.dout(n162),.clk(gclk));
	jand g0091(.dina(w_n162_0[2]),.dinb(w_n98_1[1]),.dout(n163),.clk(gclk));
	jnot g0092(.din(w_n163_0[1]),.dout(n164),.clk(gclk));
	jand g0093(.dina(w_G41_1[0]),.dinb(w_G33_11[0]),.dout(n165),.clk(gclk));
	jor g0094(.dina(w_dff_B_WYnzbP1T3_0),.dinb(w_n115_1[0]),.dout(n166),.clk(gclk));
	jor g0095(.dina(w_n162_0[1]),.dinb(w_G274_0[2]),.dout(n167),.clk(gclk));
	jand g0096(.dina(n167),.dinb(w_n166_3[1]),.dout(n168),.clk(gclk));
	jand g0097(.dina(n168),.dinb(n164),.dout(n169),.clk(gclk));
	jor g0098(.dina(w_dff_B_2Q9ieLS33_0),.dinb(n160),.dout(n170),.clk(gclk));
	jand g0099(.dina(w_n170_0[2]),.dinb(w_n146_3[2]),.dout(n171),.clk(gclk));
	jand g0100(.dina(w_G97_4[2]),.dinb(w_G33_10[2]),.dout(n172),.clk(gclk));
	jand g0101(.dina(w_G68_4[2]),.dinb(w_n148_8[2]),.dout(n173),.clk(gclk));
	jor g0102(.dina(n173),.dinb(w_G20_6[1]),.dout(n174),.clk(gclk));
	jor g0103(.dina(n174),.dinb(w_n172_0[1]),.dout(n175),.clk(gclk));
	jnot g0104(.din(n175),.dout(n176),.clk(gclk));
	jor g0105(.dina(w_n112_5[1]),.dinb(w_n113_3[0]),.dout(n177),.clk(gclk));
	jor g0106(.dina(n177),.dinb(w_n148_8[1]),.dout(n178),.clk(gclk));
	jand g0107(.dina(n178),.dinb(w_n115_0[2]),.dout(n179),.clk(gclk));
	jand g0108(.dina(w_n81_0[1]),.dinb(w_n97_1[2]),.dout(n180),.clk(gclk));
	jand g0109(.dina(w_n180_0[1]),.dinb(w_G20_6[0]),.dout(n181),.clk(gclk));
	jor g0110(.dina(n181),.dinb(w_n179_1[2]),.dout(n182),.clk(gclk));
	jor g0111(.dina(n182),.dinb(n176),.dout(n183),.clk(gclk));
	jand g0112(.dina(w_G20_5[2]),.dinb(w_n113_2[2]),.dout(n184),.clk(gclk));
	jand g0113(.dina(n184),.dinb(w_G13_0[2]),.dout(n185),.clk(gclk));
	jand g0114(.dina(w_n185_3[2]),.dinb(w_n97_1[1]),.dout(n186),.clk(gclk));
	jnot g0115(.din(n186),.dout(n187),.clk(gclk));
	jand g0116(.dina(w_n85_0[1]),.dinb(w_G33_10[1]),.dout(n188),.clk(gclk));
	jor g0117(.dina(n188),.dinb(w_n147_0[1]),.dout(n189),.clk(gclk));
	jor g0118(.dina(w_n185_3[1]),.dinb(w_n189_2[1]),.dout(n190),.clk(gclk));
	jand g0119(.dina(w_G33_10[0]),.dinb(w_n113_2[1]),.dout(n191),.clk(gclk));
	jor g0120(.dina(w_n191_0[2]),.dinb(w_n97_1[0]),.dout(n192),.clk(gclk));
	jor g0121(.dina(w_dff_B_CTKC3q9z3_0),.dinb(w_n190_1[2]),.dout(n193),.clk(gclk));
	jand g0122(.dina(n193),.dinb(n187),.dout(n194),.clk(gclk));
	jand g0123(.dina(n194),.dinb(n183),.dout(n195),.clk(gclk));
	jnot g0124(.din(w_G179_2[2]),.dout(n196),.clk(gclk));
	jor g0125(.dina(w_n154_0[0]),.dinb(w_G33_9[2]),.dout(n197),.clk(gclk));
	jor g0126(.dina(w_n197_1[1]),.dinb(w_n103_0[1]),.dout(n198),.clk(gclk));
	jor g0127(.dina(w_G1698_0[0]),.dinb(w_G33_9[1]),.dout(n199),.clk(gclk));
	jor g0128(.dina(w_n199_1[1]),.dinb(w_n93_0[0]),.dout(n200),.clk(gclk));
	jnot g0129(.din(w_n157_0[1]),.dout(n201),.clk(gclk));
	jand g0130(.dina(w_n201_0[1]),.dinb(n200),.dout(n202),.clk(gclk));
	jand g0131(.dina(n202),.dinb(n198),.dout(n203),.clk(gclk));
	jor g0132(.dina(n203),.dinb(w_n166_3[0]),.dout(n204),.clk(gclk));
	jnot g0133(.din(w_G274_0[1]),.dout(n205),.clk(gclk));
	jand g0134(.dina(w_G45_1[1]),.dinb(w_n113_2[0]),.dout(n206),.clk(gclk));
	jand g0135(.dina(w_n206_0[1]),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jor g0136(.dina(n207),.dinb(w_n151_4[1]),.dout(n208),.clk(gclk));
	jor g0137(.dina(n208),.dinb(w_n163_0[0]),.dout(n209),.clk(gclk));
	jand g0138(.dina(n209),.dinb(n204),.dout(n210),.clk(gclk));
	jand g0139(.dina(w_n210_0[2]),.dinb(w_n196_2[2]),.dout(n211),.clk(gclk));
	jor g0140(.dina(n211),.dinb(w_n195_0[1]),.dout(n212),.clk(gclk));
	jor g0141(.dina(n212),.dinb(n171),.dout(n213),.clk(gclk));
	jnot g0142(.din(w_n195_0[0]),.dout(n214),.clk(gclk));
	jand g0143(.dina(w_n210_0[1]),.dinb(w_G190_4[1]),.dout(n215),.clk(gclk));
	jand g0144(.dina(w_n170_0[1]),.dinb(w_G200_4[2]),.dout(n216),.clk(gclk));
	jor g0145(.dina(n216),.dinb(w_dff_B_suPl964r6_1),.dout(n217),.clk(gclk));
	jor g0146(.dina(n217),.dinb(w_n214_0[1]),.dout(n218),.clk(gclk));
	jand g0147(.dina(w_n218_0[1]),.dinb(w_n213_0[1]),.dout(n219),.clk(gclk));
	jor g0148(.dina(w_n197_1[0]),.dinb(w_n98_1[0]),.dout(n220),.clk(gclk));
	jand g0149(.dina(w_G283_3[2]),.dinb(w_G33_9[0]),.dout(n221),.clk(gclk));
	jnot g0150(.din(w_n221_0[2]),.dout(n222),.clk(gclk));
	jor g0151(.dina(w_n199_1[0]),.dinb(w_n103_0[0]),.dout(n223),.clk(gclk));
	jand g0152(.dina(n223),.dinb(n222),.dout(n224),.clk(gclk));
	jand g0153(.dina(n224),.dinb(n220),.dout(n225),.clk(gclk));
	jor g0154(.dina(n225),.dinb(w_n166_2[2]),.dout(n226),.clk(gclk));
	jor g0155(.dina(w_n151_4[0]),.dinb(w_n205_0[0]),.dout(n227),.clk(gclk));
	jor g0156(.dina(w_n162_0[0]),.dinb(w_G41_0[2]),.dout(n228),.clk(gclk));
	jor g0157(.dina(w_n228_0[1]),.dinb(n227),.dout(n229),.clk(gclk));
	jand g0158(.dina(w_n206_0[0]),.dinb(w_n149_2[0]),.dout(n230),.clk(gclk));
	jor g0159(.dina(w_n230_0[1]),.dinb(w_n151_3[2]),.dout(n231),.clk(gclk));
	jor g0160(.dina(w_n231_0[2]),.dinb(w_n91_1[0]),.dout(n232),.clk(gclk));
	jand g0161(.dina(n232),.dinb(w_n229_0[2]),.dout(n233),.clk(gclk));
	jand g0162(.dina(n233),.dinb(w_dff_B_pauv6il10_1),.dout(n234),.clk(gclk));
	jor g0163(.dina(w_n234_0[2]),.dinb(w_n146_3[1]),.dout(n235),.clk(gclk));
	jand g0164(.dina(w_n152_3[0]),.dinb(w_G250_0[1]),.dout(n236),.clk(gclk));
	jand g0165(.dina(w_n155_3[0]),.dinb(w_G244_0[2]),.dout(n237),.clk(gclk));
	jor g0166(.dina(n237),.dinb(w_n221_0[1]),.dout(n238),.clk(gclk));
	jor g0167(.dina(n238),.dinb(w_dff_B_HzC0cx2C7_1),.dout(n239),.clk(gclk));
	jand g0168(.dina(n239),.dinb(w_n151_3[1]),.dout(n240),.clk(gclk));
	jand g0169(.dina(w_n166_2[1]),.dinb(w_G274_0[0]),.dout(n241),.clk(gclk));
	jand g0170(.dina(w_n230_0[0]),.dinb(w_n241_0[1]),.dout(n242),.clk(gclk));
	jand g0171(.dina(w_n228_0[0]),.dinb(w_n166_2[0]),.dout(n243),.clk(gclk));
	jand g0172(.dina(w_n243_0[2]),.dinb(w_G257_1[0]),.dout(n244),.clk(gclk));
	jor g0173(.dina(n244),.dinb(w_n242_0[2]),.dout(n245),.clk(gclk));
	jor g0174(.dina(n245),.dinb(n240),.dout(n246),.clk(gclk));
	jor g0175(.dina(w_n246_1[1]),.dinb(w_n196_2[1]),.dout(n247),.clk(gclk));
	jand g0176(.dina(n247),.dinb(n235),.dout(n248),.clk(gclk));
	jand g0177(.dina(w_G107_4[2]),.dinb(w_G33_8[2]),.dout(n249),.clk(gclk));
	jand g0178(.dina(w_G77_4[2]),.dinb(w_n148_8[0]),.dout(n250),.clk(gclk));
	jor g0179(.dina(n250),.dinb(w_G20_5[1]),.dout(n251),.clk(gclk));
	jor g0180(.dina(n251),.dinb(w_n249_0[1]),.dout(n252),.clk(gclk));
	jand g0181(.dina(w_G107_4[1]),.dinb(w_G97_4[1]),.dout(n253),.clk(gclk));
	jor g0182(.dina(n253),.dinb(w_n112_5[0]),.dout(n254),.clk(gclk));
	jor g0183(.dina(n254),.dinb(w_n81_0[0]),.dout(n255),.clk(gclk));
	jand g0184(.dina(w_n255_0[1]),.dinb(n252),.dout(n256),.clk(gclk));
	jand g0185(.dina(n256),.dinb(w_n189_2[0]),.dout(n257),.clk(gclk));
	jnot g0186(.din(w_n257_0[1]),.dout(n258),.clk(gclk));
	jand g0187(.dina(w_n185_3[0]),.dinb(w_n79_0[0]),.dout(n259),.clk(gclk));
	jnot g0188(.din(w_n259_0[1]),.dout(n260),.clk(gclk));
	jnot g0189(.din(w_n191_0[1]),.dout(n261),.clk(gclk));
	jand g0190(.dina(w_n261_0[1]),.dinb(w_G97_4[0]),.dout(n262),.clk(gclk));
	jnot g0191(.din(w_n262_0[1]),.dout(n263),.clk(gclk));
	jor g0192(.dina(n263),.dinb(w_n190_1[1]),.dout(n264),.clk(gclk));
	jand g0193(.dina(n264),.dinb(w_dff_B_wdu0KqcM0_1),.dout(n265),.clk(gclk));
	jand g0194(.dina(n265),.dinb(n258),.dout(n266),.clk(gclk));
	jor g0195(.dina(w_dff_B_sT0q3vOJ5_0),.dinb(n248),.dout(n267),.clk(gclk));
	jand g0196(.dina(w_n246_1[0]),.dinb(w_G200_4[1]),.dout(n268),.clk(gclk));
	jor g0197(.dina(w_n112_4[2]),.dinb(w_G1_1[2]),.dout(n269),.clk(gclk));
	jor g0198(.dina(w_n269_1[2]),.dinb(w_n114_1[0]),.dout(n270),.clk(gclk));
	jand g0199(.dina(w_n270_0[1]),.dinb(w_n179_1[1]),.dout(n271),.clk(gclk));
	jand g0200(.dina(w_n262_0[0]),.dinb(w_n271_1[2]),.dout(n272),.clk(gclk));
	jor g0201(.dina(n272),.dinb(w_n259_0[0]),.dout(n273),.clk(gclk));
	jor g0202(.dina(n273),.dinb(w_n257_0[0]),.dout(n274),.clk(gclk));
	jand g0203(.dina(w_n234_0[1]),.dinb(w_G190_4[0]),.dout(n275),.clk(gclk));
	jor g0204(.dina(n275),.dinb(w_n274_0[2]),.dout(n276),.clk(gclk));
	jor g0205(.dina(n276),.dinb(w_dff_B_E1mUxj7c0_1),.dout(n277),.clk(gclk));
	jand g0206(.dina(n277),.dinb(n267),.dout(n278),.clk(gclk));
	jand g0207(.dina(w_n278_0[1]),.dinb(w_n219_0[1]),.dout(n279),.clk(gclk));
	jand g0208(.dina(w_n152_2[2]),.dinb(w_G264_0[2]),.dout(n280),.clk(gclk));
	jand g0209(.dina(w_G303_2[2]),.dinb(w_G33_8[1]),.dout(n281),.clk(gclk));
	jand g0210(.dina(w_n155_2[2]),.dinb(w_G257_0[2]),.dout(n282),.clk(gclk));
	jor g0211(.dina(n282),.dinb(w_n281_0[1]),.dout(n283),.clk(gclk));
	jor g0212(.dina(n283),.dinb(w_dff_B_TqeE9gwh0_1),.dout(n284),.clk(gclk));
	jand g0213(.dina(n284),.dinb(w_n151_3[0]),.dout(n285),.clk(gclk));
	jand g0214(.dina(w_n243_0[1]),.dinb(w_G270_0[0]),.dout(n286),.clk(gclk));
	jor g0215(.dina(n286),.dinb(w_n242_0[1]),.dout(n287),.clk(gclk));
	jor g0216(.dina(n287),.dinb(n285),.dout(n288),.clk(gclk));
	jand g0217(.dina(w_n288_1[1]),.dinb(w_n146_3[0]),.dout(n289),.clk(gclk));
	jand g0218(.dina(w_G97_3[2]),.dinb(w_n148_7[2]),.dout(n290),.clk(gclk));
	jor g0219(.dina(n290),.dinb(w_G20_5[0]),.dout(n291),.clk(gclk));
	jor g0220(.dina(n291),.dinb(w_n221_0[0]),.dout(n292),.clk(gclk));
	jand g0221(.dina(w_n105_2[0]),.dinb(w_G20_4[2]),.dout(n293),.clk(gclk));
	jnot g0222(.din(n293),.dout(n294),.clk(gclk));
	jand g0223(.dina(n294),.dinb(w_n189_1[2]),.dout(n295),.clk(gclk));
	jand g0224(.dina(n295),.dinb(n292),.dout(n296),.clk(gclk));
	jnot g0225(.din(w_n296_0[1]),.dout(n297),.clk(gclk));
	jand g0226(.dina(w_n185_2[2]),.dinb(w_n105_1[2]),.dout(n298),.clk(gclk));
	jnot g0227(.din(w_n298_0[1]),.dout(n299),.clk(gclk));
	jor g0228(.dina(w_n191_0[0]),.dinb(w_n105_1[1]),.dout(n300),.clk(gclk));
	jor g0229(.dina(w_n300_0[1]),.dinb(w_n190_1[0]),.dout(n301),.clk(gclk));
	jand g0230(.dina(n301),.dinb(n299),.dout(n302),.clk(gclk));
	jand g0231(.dina(n302),.dinb(n297),.dout(n303),.clk(gclk));
	jor g0232(.dina(w_n197_0[2]),.dinb(w_n88_0[2]),.dout(n304),.clk(gclk));
	jnot g0233(.din(w_n281_0[0]),.dout(n305),.clk(gclk));
	jor g0234(.dina(w_n199_0[2]),.dinb(w_n91_0[2]),.dout(n306),.clk(gclk));
	jand g0235(.dina(n306),.dinb(n305),.dout(n307),.clk(gclk));
	jand g0236(.dina(n307),.dinb(n304),.dout(n308),.clk(gclk));
	jor g0237(.dina(n308),.dinb(w_n166_1[2]),.dout(n309),.clk(gclk));
	jor g0238(.dina(w_n231_0[1]),.dinb(w_n106_0[0]),.dout(n310),.clk(gclk));
	jand g0239(.dina(n310),.dinb(w_n229_0[1]),.dout(n311),.clk(gclk));
	jand g0240(.dina(n311),.dinb(w_dff_B_xzNoOxiA6_1),.dout(n312),.clk(gclk));
	jand g0241(.dina(w_n312_1[1]),.dinb(w_n196_2[0]),.dout(n313),.clk(gclk));
	jor g0242(.dina(n313),.dinb(w_n303_0[1]),.dout(n314),.clk(gclk));
	jor g0243(.dina(n314),.dinb(w_dff_B_IpaO9w8W7_1),.dout(n315),.clk(gclk));
	jand g0244(.dina(w_n288_1[0]),.dinb(w_G200_4[0]),.dout(n316),.clk(gclk));
	jnot g0245(.din(w_n300_0[0]),.dout(n317),.clk(gclk));
	jand g0246(.dina(w_dff_B_igReF1fn0_0),.dinb(w_n271_1[1]),.dout(n318),.clk(gclk));
	jor g0247(.dina(n318),.dinb(w_n298_0[0]),.dout(n319),.clk(gclk));
	jor g0248(.dina(n319),.dinb(w_n296_0[0]),.dout(n320),.clk(gclk));
	jand g0249(.dina(w_n312_1[0]),.dinb(w_G190_3[2]),.dout(n321),.clk(gclk));
	jor g0250(.dina(n321),.dinb(w_n320_0[1]),.dout(n322),.clk(gclk));
	jor g0251(.dina(n322),.dinb(w_dff_B_WMEaKdvL2_1),.dout(n323),.clk(gclk));
	jand g0252(.dina(n323),.dinb(w_n315_0[1]),.dout(n324),.clk(gclk));
	jor g0253(.dina(w_n97_0[2]),.dinb(w_G33_8[0]),.dout(n325),.clk(gclk));
	jand g0254(.dina(n325),.dinb(w_n112_4[1]),.dout(n326),.clk(gclk));
	jand g0255(.dina(n326),.dinb(w_n201_0[0]),.dout(n327),.clk(gclk));
	jor g0256(.dina(n327),.dinb(w_n179_1[0]),.dout(n328),.clk(gclk));
	jor g0257(.dina(w_n328_0[1]),.dinb(w_G20_4[1]),.dout(n329),.clk(gclk));
	jand g0258(.dina(n329),.dinb(w_G107_4[0]),.dout(n330),.clk(gclk));
	jand g0259(.dina(w_n328_0[0]),.dinb(w_n270_0[0]),.dout(n331),.clk(gclk));
	jor g0260(.dina(w_dff_B_MNYOayjY1_0),.dinb(n330),.dout(n332),.clk(gclk));
	jand g0261(.dina(w_n261_0[0]),.dinb(w_G107_3[2]),.dout(n333),.clk(gclk));
	jand g0262(.dina(w_dff_B_UDmTyMk91_0),.dinb(w_n271_1[0]),.dout(n334),.clk(gclk));
	jnot g0263(.din(w_n334_0[1]),.dout(n335),.clk(gclk));
	jand g0264(.dina(w_dff_B_xrpfOxV02_0),.dinb(n332),.dout(n336),.clk(gclk));
	jor g0265(.dina(w_n197_0[1]),.dinb(w_n91_0[1]),.dout(n337),.clk(gclk));
	jor g0266(.dina(w_n199_0[1]),.dinb(w_n98_0[2]),.dout(n338),.clk(gclk));
	jand g0267(.dina(w_G294_3[1]),.dinb(w_G33_7[2]),.dout(n339),.clk(gclk));
	jnot g0268(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jand g0269(.dina(n340),.dinb(n338),.dout(n341),.clk(gclk));
	jand g0270(.dina(n341),.dinb(n337),.dout(n342),.clk(gclk));
	jor g0271(.dina(n342),.dinb(w_n166_1[1]),.dout(n343),.clk(gclk));
	jor g0272(.dina(w_n231_0[0]),.dinb(w_n88_0[1]),.dout(n344),.clk(gclk));
	jand g0273(.dina(n344),.dinb(w_n229_0[0]),.dout(n345),.clk(gclk));
	jand g0274(.dina(n345),.dinb(w_dff_B_0LuljrnG7_1),.dout(n346),.clk(gclk));
	jand g0275(.dina(w_n346_1[1]),.dinb(w_n196_1[2]),.dout(n347),.clk(gclk));
	jand g0276(.dina(w_n152_2[1]),.dinb(w_G257_0[1]),.dout(n348),.clk(gclk));
	jand g0277(.dina(w_n155_2[1]),.dinb(w_G250_0[0]),.dout(n349),.clk(gclk));
	jor g0278(.dina(w_n339_0[0]),.dinb(n349),.dout(n350),.clk(gclk));
	jor g0279(.dina(n350),.dinb(w_dff_B_Dh2jux470_1),.dout(n351),.clk(gclk));
	jand g0280(.dina(n351),.dinb(w_n151_2[2]),.dout(n352),.clk(gclk));
	jand g0281(.dina(w_n243_0[0]),.dinb(w_G264_0[1]),.dout(n353),.clk(gclk));
	jor g0282(.dina(n353),.dinb(w_n242_0[0]),.dout(n354),.clk(gclk));
	jor g0283(.dina(n354),.dinb(n352),.dout(n355),.clk(gclk));
	jand g0284(.dina(w_n355_1[1]),.dinb(w_n146_2[2]),.dout(n356),.clk(gclk));
	jor g0285(.dina(n356),.dinb(n347),.dout(n357),.clk(gclk));
	jor g0286(.dina(n357),.dinb(n336),.dout(n358),.clk(gclk));
	jand g0287(.dina(w_G87_3[0]),.dinb(w_n148_7[1]),.dout(n359),.clk(gclk));
	jor g0288(.dina(n359),.dinb(w_G20_4[0]),.dout(n360),.clk(gclk));
	jor g0289(.dina(n360),.dinb(w_n157_0[0]),.dout(n361),.clk(gclk));
	jand g0290(.dina(n361),.dinb(w_n189_1[1]),.dout(n362),.clk(gclk));
	jand g0291(.dina(w_n362_0[1]),.dinb(w_n112_4[0]),.dout(n363),.clk(gclk));
	jor g0292(.dina(n363),.dinb(w_n80_0[2]),.dout(n364),.clk(gclk));
	jor g0293(.dina(w_n362_0[0]),.dinb(w_n185_2[1]),.dout(n365),.clk(gclk));
	jand g0294(.dina(w_dff_B_nuHoV5pA2_0),.dinb(n364),.dout(n366),.clk(gclk));
	jor g0295(.dina(w_n334_0[0]),.dinb(n366),.dout(n367),.clk(gclk));
	jor g0296(.dina(w_n355_1[0]),.dinb(w_G190_3[1]),.dout(n368),.clk(gclk));
	jor g0297(.dina(w_n346_1[0]),.dinb(w_G200_3[2]),.dout(n369),.clk(gclk));
	jand g0298(.dina(n369),.dinb(n368),.dout(n370),.clk(gclk));
	jor g0299(.dina(n370),.dinb(w_n367_0[2]),.dout(n371),.clk(gclk));
	jand g0300(.dina(w_n371_0[1]),.dinb(n358),.dout(n372),.clk(gclk));
	jand g0301(.dina(w_n372_0[1]),.dinb(w_n324_0[1]),.dout(n373),.clk(gclk));
	jand g0302(.dina(n373),.dinb(w_n279_0[1]),.dout(n374),.clk(gclk));
	jand g0303(.dina(w_n155_2[0]),.dinb(w_G232_1[0]),.dout(n375),.clk(gclk));
	jand g0304(.dina(w_n152_2[0]),.dinb(w_G238_0[2]),.dout(n376),.clk(gclk));
	jor g0305(.dina(n376),.dinb(w_n249_0[0]),.dout(n377),.clk(gclk));
	jor g0306(.dina(n377),.dinb(w_dff_B_v9vq1SUv1_1),.dout(n378),.clk(gclk));
	jand g0307(.dina(n378),.dinb(w_n151_2[1]),.dout(n379),.clk(gclk));
	jand g0308(.dina(w_n161_1[0]),.dinb(w_n149_1[2]),.dout(n380),.clk(gclk));
	jor g0309(.dina(n380),.dinb(w_G1_1[1]),.dout(n381),.clk(gclk));
	jand g0310(.dina(w_n381_0[1]),.dinb(w_n166_1[0]),.dout(n382),.clk(gclk));
	jand g0311(.dina(w_n382_1[1]),.dinb(w_G244_0[1]),.dout(n383),.clk(gclk));
	jnot g0312(.din(w_n381_0[0]),.dout(n384),.clk(gclk));
	jand g0313(.dina(n384),.dinb(w_n241_0[0]),.dout(n385),.clk(gclk));
	jor g0314(.dina(w_n385_1[1]),.dinb(n383),.dout(n386),.clk(gclk));
	jor g0315(.dina(n386),.dinb(n379),.dout(n387),.clk(gclk));
	jand g0316(.dina(w_n387_1[1]),.dinb(w_n146_2[1]),.dout(n388),.clk(gclk));
	jnot g0317(.din(n388),.dout(n389),.clk(gclk));
	jand g0318(.dina(w_G87_2[2]),.dinb(w_G33_7[1]),.dout(n390),.clk(gclk));
	jand g0319(.dina(w_G58_4[2]),.dinb(w_n148_7[0]),.dout(n391),.clk(gclk));
	jor g0320(.dina(n391),.dinb(w_G20_3[2]),.dout(n392),.clk(gclk));
	jor g0321(.dina(n392),.dinb(w_n390_0[1]),.dout(n393),.clk(gclk));
	jor g0322(.dina(w_G77_4[1]),.dinb(w_n112_3[2]),.dout(n394),.clk(gclk));
	jand g0323(.dina(w_dff_B_I3nt5hgZ5_0),.dinb(w_n189_1[0]),.dout(n395),.clk(gclk));
	jand g0324(.dina(n395),.dinb(n393),.dout(n396),.clk(gclk));
	jand g0325(.dina(w_n185_2[0]),.dinb(w_n72_0[2]),.dout(n397),.clk(gclk));
	jand g0326(.dina(w_n269_1[1]),.dinb(w_G77_4[0]),.dout(n398),.clk(gclk));
	jand g0327(.dina(w_dff_B_7Nb557uG9_0),.dinb(w_n271_0[2]),.dout(n399),.clk(gclk));
	jor g0328(.dina(n399),.dinb(w_dff_B_dP8ERMqf7_1),.dout(n400),.clk(gclk));
	jor g0329(.dina(n400),.dinb(w_dff_B_w8aVsJPu0_1),.dout(n401),.clk(gclk));
	jor g0330(.dina(w_n387_1[0]),.dinb(w_G179_2[1]),.dout(n402),.clk(gclk));
	jand g0331(.dina(n402),.dinb(w_n401_0[2]),.dout(n403),.clk(gclk));
	jand g0332(.dina(n403),.dinb(n389),.dout(n404),.clk(gclk));
	jnot g0333(.din(w_n404_0[2]),.dout(n405),.clk(gclk));
	jand g0334(.dina(w_n387_0[2]),.dinb(w_G200_3[1]),.dout(n406),.clk(gclk));
	jnot g0335(.din(w_G190_3[0]),.dout(n407),.clk(gclk));
	jor g0336(.dina(w_n387_0[1]),.dinb(w_n407_2[1]),.dout(n408),.clk(gclk));
	jnot g0337(.din(n408),.dout(n409),.clk(gclk));
	jor g0338(.dina(n409),.dinb(w_n401_0[1]),.dout(n410),.clk(gclk));
	jor g0339(.dina(n410),.dinb(w_dff_B_Ja2zN20d8_1),.dout(n411),.clk(gclk));
	jand g0340(.dina(n411),.dinb(w_n405_0[1]),.dout(n412),.clk(gclk));
	jand g0341(.dina(w_n155_1[2]),.dinb(w_G226_1[0]),.dout(n413),.clk(gclk));
	jand g0342(.dina(w_n152_1[2]),.dinb(w_G232_0[2]),.dout(n414),.clk(gclk));
	jor g0343(.dina(n414),.dinb(w_n172_0[0]),.dout(n415),.clk(gclk));
	jor g0344(.dina(n415),.dinb(w_dff_B_kXyk0Mo37_1),.dout(n416),.clk(gclk));
	jand g0345(.dina(n416),.dinb(w_n151_2[0]),.dout(n417),.clk(gclk));
	jand g0346(.dina(w_n382_1[0]),.dinb(w_G238_0[1]),.dout(n418),.clk(gclk));
	jor g0347(.dina(n418),.dinb(w_n385_1[0]),.dout(n419),.clk(gclk));
	jor g0348(.dina(n419),.dinb(n417),.dout(n420),.clk(gclk));
	jand g0349(.dina(w_n420_1[1]),.dinb(w_n146_2[0]),.dout(n421),.clk(gclk));
	jnot g0350(.din(n421),.dout(n422),.clk(gclk));
	jand g0351(.dina(w_n269_1[0]),.dinb(w_G68_4[1]),.dout(n423),.clk(gclk));
	jand g0352(.dina(w_dff_B_Hn1TlILC1_0),.dinb(w_n271_0[1]),.dout(n424),.clk(gclk));
	jand g0353(.dina(w_n148_6[2]),.dinb(w_n114_0[2]),.dout(n425),.clk(gclk));
	jnot g0354(.din(w_n425_1[2]),.dout(n426),.clk(gclk));
	jand g0355(.dina(w_n426_0[1]),.dinb(w_n85_0[0]),.dout(n427),.clk(gclk));
	jor g0356(.dina(n427),.dinb(w_n185_1[2]),.dout(n428),.clk(gclk));
	jand g0357(.dina(n428),.dinb(w_n75_0[2]),.dout(n429),.clk(gclk));
	jand g0358(.dina(w_G77_3[2]),.dinb(w_G33_7[0]),.dout(n430),.clk(gclk));
	jand g0359(.dina(w_G50_4[2]),.dinb(w_n148_6[1]),.dout(n431),.clk(gclk));
	jor g0360(.dina(n431),.dinb(w_n430_0[1]),.dout(n432),.clk(gclk));
	jand g0361(.dina(n432),.dinb(w_n112_3[1]),.dout(n433),.clk(gclk));
	jand g0362(.dina(n433),.dinb(w_n189_0[2]),.dout(n434),.clk(gclk));
	jor g0363(.dina(w_dff_B_aqXTkkMr3_0),.dinb(n429),.dout(n435),.clk(gclk));
	jor g0364(.dina(n435),.dinb(w_dff_B_3aaOt5mu4_1),.dout(n436),.clk(gclk));
	jor g0365(.dina(w_n420_1[0]),.dinb(w_G179_2[0]),.dout(n437),.clk(gclk));
	jand g0366(.dina(n437),.dinb(w_n436_0[2]),.dout(n438),.clk(gclk));
	jand g0367(.dina(n438),.dinb(n422),.dout(n439),.clk(gclk));
	jnot g0368(.din(w_n439_1[1]),.dout(n440),.clk(gclk));
	jand g0369(.dina(w_n420_0[2]),.dinb(w_G200_3[0]),.dout(n441),.clk(gclk));
	jor g0370(.dina(w_n420_0[1]),.dinb(w_n407_2[0]),.dout(n442),.clk(gclk));
	jnot g0371(.din(n442),.dout(n443),.clk(gclk));
	jor g0372(.dina(n443),.dinb(w_n436_0[1]),.dout(n444),.clk(gclk));
	jor g0373(.dina(n444),.dinb(w_dff_B_ubAYFKGy2_1),.dout(n445),.clk(gclk));
	jand g0374(.dina(w_n445_0[1]),.dinb(n440),.dout(n446),.clk(gclk));
	jand g0375(.dina(w_n446_0[1]),.dinb(w_n412_0[1]),.dout(n447),.clk(gclk));
	jand g0376(.dina(w_n152_1[1]),.dinb(w_G223_0[1]),.dout(n448),.clk(gclk));
	jand g0377(.dina(w_n155_1[1]),.dinb(w_dff_B_ymDCuxVv0_1),.dout(n449),.clk(gclk));
	jor g0378(.dina(n449),.dinb(w_n430_0[0]),.dout(n450),.clk(gclk));
	jor g0379(.dina(n450),.dinb(w_dff_B_PusZ0kJy6_1),.dout(n451),.clk(gclk));
	jand g0380(.dina(n451),.dinb(w_n151_1[2]),.dout(n452),.clk(gclk));
	jand g0381(.dina(w_n382_0[2]),.dinb(w_G226_0[2]),.dout(n453),.clk(gclk));
	jor g0382(.dina(n453),.dinb(w_n385_0[2]),.dout(n454),.clk(gclk));
	jor g0383(.dina(n454),.dinb(n452),.dout(n455),.clk(gclk));
	jand g0384(.dina(w_n455_0[2]),.dinb(w_n146_1[2]),.dout(n456),.clk(gclk));
	jand g0385(.dina(w_n269_0[2]),.dinb(w_G50_4[1]),.dout(n457),.clk(gclk));
	jnot g0386(.din(n457),.dout(n458),.clk(gclk));
	jor g0387(.dina(n458),.dinb(w_n190_0[2]),.dout(n459),.clk(gclk));
	jor g0388(.dina(w_n77_0[0]),.dinb(w_n112_3[0]),.dout(n460),.clk(gclk));
	jnot g0389(.din(w_G150_3[1]),.dout(n461),.clk(gclk));
	jand g0390(.dina(w_n148_6[0]),.dinb(w_n112_2[2]),.dout(n462),.clk(gclk));
	jnot g0391(.din(w_n462_0[2]),.dout(n463),.clk(gclk));
	jor g0392(.dina(n463),.dinb(w_dff_B_6GLiXLf15_1),.dout(n464),.clk(gclk));
	jand g0393(.dina(w_G33_6[2]),.dinb(w_n112_2[1]),.dout(n465),.clk(gclk));
	jand g0394(.dina(w_n465_0[1]),.dinb(w_G58_4[1]),.dout(n466),.clk(gclk));
	jnot g0395(.din(n466),.dout(n467),.clk(gclk));
	jand g0396(.dina(n467),.dinb(n464),.dout(n468),.clk(gclk));
	jand g0397(.dina(n468),.dinb(w_dff_B_oW9LfIcp4_1),.dout(n469),.clk(gclk));
	jor g0398(.dina(n469),.dinb(w_n179_0[2]),.dout(n470),.clk(gclk));
	jand g0399(.dina(w_n185_1[1]),.dinb(w_n73_2[0]),.dout(n471),.clk(gclk));
	jnot g0400(.din(n471),.dout(n472),.clk(gclk));
	jand g0401(.dina(w_dff_B_7SgsIywN8_0),.dinb(n470),.dout(n473),.clk(gclk));
	jand g0402(.dina(n473),.dinb(w_dff_B_7vdPgLY42_1),.dout(n474),.clk(gclk));
	jnot g0403(.din(w_n455_0[1]),.dout(n475),.clk(gclk));
	jand g0404(.dina(w_n475_0[1]),.dinb(w_n196_1[1]),.dout(n476),.clk(gclk));
	jor g0405(.dina(n476),.dinb(w_n474_0[1]),.dout(n477),.clk(gclk));
	jor g0406(.dina(n477),.dinb(w_dff_B_CaBe6qHK8_1),.dout(n478),.clk(gclk));
	jnot g0407(.din(w_n474_0[0]),.dout(n479),.clk(gclk));
	jand g0408(.dina(w_n475_0[0]),.dinb(w_G190_2[2]),.dout(n480),.clk(gclk));
	jand g0409(.dina(w_n455_0[0]),.dinb(w_G200_2[2]),.dout(n481),.clk(gclk));
	jor g0410(.dina(w_dff_B_GpNB0XTN4_0),.dinb(n480),.dout(n482),.clk(gclk));
	jor g0411(.dina(n482),.dinb(w_n479_0[1]),.dout(n483),.clk(gclk));
	jand g0412(.dina(w_n483_0[1]),.dinb(w_n478_0[1]),.dout(n484),.clk(gclk));
	jand g0413(.dina(w_n152_1[0]),.dinb(w_G226_0[1]),.dout(n485),.clk(gclk));
	jand g0414(.dina(w_n155_1[0]),.dinb(w_G223_0[0]),.dout(n486),.clk(gclk));
	jor g0415(.dina(n486),.dinb(w_n390_0[0]),.dout(n487),.clk(gclk));
	jor g0416(.dina(n487),.dinb(w_dff_B_pJ9vBfb10_1),.dout(n488),.clk(gclk));
	jand g0417(.dina(n488),.dinb(w_n151_1[1]),.dout(n489),.clk(gclk));
	jand g0418(.dina(w_n382_0[1]),.dinb(w_G232_0[1]),.dout(n490),.clk(gclk));
	jor g0419(.dina(n490),.dinb(w_n385_0[1]),.dout(n491),.clk(gclk));
	jor g0420(.dina(n491),.dinb(n489),.dout(n492),.clk(gclk));
	jand g0421(.dina(w_n492_0[2]),.dinb(w_n146_1[1]),.dout(n493),.clk(gclk));
	jand g0422(.dina(w_n269_0[1]),.dinb(w_G58_4[0]),.dout(n494),.clk(gclk));
	jnot g0423(.din(n494),.dout(n495),.clk(gclk));
	jor g0424(.dina(n495),.dinb(w_n190_0[1]),.dout(n496),.clk(gclk));
	jor g0425(.dina(w_n137_0[1]),.dinb(w_n112_2[0]),.dout(n497),.clk(gclk));
	jand g0426(.dina(w_n462_0[1]),.dinb(w_G159_3[2]),.dout(n498),.clk(gclk));
	jand g0427(.dina(w_n465_0[0]),.dinb(w_G68_4[0]),.dout(n499),.clk(gclk));
	jor g0428(.dina(n499),.dinb(n498),.dout(n500),.clk(gclk));
	jnot g0429(.din(n500),.dout(n501),.clk(gclk));
	jand g0430(.dina(n501),.dinb(w_dff_B_YL6HbYWE5_1),.dout(n502),.clk(gclk));
	jor g0431(.dina(n502),.dinb(w_n179_0[1]),.dout(n503),.clk(gclk));
	jand g0432(.dina(w_n185_1[0]),.dinb(w_n74_0[2]),.dout(n504),.clk(gclk));
	jnot g0433(.din(n504),.dout(n505),.clk(gclk));
	jand g0434(.dina(w_dff_B_Qwl99s273_0),.dinb(n503),.dout(n506),.clk(gclk));
	jand g0435(.dina(n506),.dinb(w_dff_B_E3nHGAMP2_1),.dout(n507),.clk(gclk));
	jnot g0436(.din(w_n492_0[1]),.dout(n508),.clk(gclk));
	jand g0437(.dina(w_n508_0[1]),.dinb(w_n196_1[0]),.dout(n509),.clk(gclk));
	jor g0438(.dina(n509),.dinb(w_n507_0[1]),.dout(n510),.clk(gclk));
	jor g0439(.dina(n510),.dinb(w_dff_B_tU88pgl64_1),.dout(n511),.clk(gclk));
	jnot g0440(.din(w_n507_0[0]),.dout(n512),.clk(gclk));
	jand g0441(.dina(w_n508_0[0]),.dinb(w_G190_2[1]),.dout(n513),.clk(gclk));
	jand g0442(.dina(w_n492_0[0]),.dinb(w_G200_2[1]),.dout(n514),.clk(gclk));
	jor g0443(.dina(w_dff_B_mjwAJ0fu9_0),.dinb(n513),.dout(n515),.clk(gclk));
	jor g0444(.dina(n515),.dinb(w_n512_0[1]),.dout(n516),.clk(gclk));
	jand g0445(.dina(w_n516_0[1]),.dinb(w_n511_0[1]),.dout(n517),.clk(gclk));
	jand g0446(.dina(w_n517_0[1]),.dinb(w_n484_0[1]),.dout(n518),.clk(gclk));
	jand g0447(.dina(n518),.dinb(n447),.dout(n519),.clk(gclk));
	jand g0448(.dina(w_n519_1[2]),.dinb(w_n374_0[1]),.dout(w_dff_A_Fo7AjoZB3_2),.clk(gclk));
	jor g0449(.dina(w_n355_0[2]),.dinb(w_G179_1[2]),.dout(n521),.clk(gclk));
	jor g0450(.dina(w_n346_0[2]),.dinb(w_G169_1[0]),.dout(n522),.clk(gclk));
	jand g0451(.dina(n522),.dinb(n521),.dout(n523),.clk(gclk));
	jand g0452(.dina(w_n523_0[1]),.dinb(w_n367_0[1]),.dout(n524),.clk(gclk));
	jor g0453(.dina(w_n312_0[2]),.dinb(w_G169_0[2]),.dout(n525),.clk(gclk));
	jor g0454(.dina(w_n288_0[2]),.dinb(w_G179_1[1]),.dout(n526),.clk(gclk));
	jand g0455(.dina(n526),.dinb(w_n320_0[0]),.dout(n527),.clk(gclk));
	jand g0456(.dina(n527),.dinb(w_dff_B_LzLWH8KM7_1),.dout(n528),.clk(gclk));
	jand g0457(.dina(w_n371_0[0]),.dinb(w_n528_0[1]),.dout(n529),.clk(gclk));
	jor g0458(.dina(n529),.dinb(w_n524_0[1]),.dout(n530),.clk(gclk));
	jand g0459(.dina(n530),.dinb(w_n279_0[0]),.dout(n531),.clk(gclk));
	jnot g0460(.din(w_n213_0[0]),.dout(n532),.clk(gclk));
	jand g0461(.dina(w_n246_0[2]),.dinb(w_G169_0[1]),.dout(n533),.clk(gclk));
	jand g0462(.dina(w_n234_0[0]),.dinb(w_G179_1[0]),.dout(n534),.clk(gclk));
	jor g0463(.dina(w_n534_0[1]),.dinb(n533),.dout(n535),.clk(gclk));
	jand g0464(.dina(w_n274_0[1]),.dinb(n535),.dout(n536),.clk(gclk));
	jand g0465(.dina(w_n536_0[2]),.dinb(w_n218_0[0]),.dout(n537),.clk(gclk));
	jor g0466(.dina(n537),.dinb(w_n532_0[1]),.dout(n538),.clk(gclk));
	jor g0467(.dina(w_dff_B_Yea19fe24_0),.dinb(n531),.dout(n539),.clk(gclk));
	jand g0468(.dina(w_n539_0[1]),.dinb(w_n519_1[1]),.dout(n540),.clk(gclk));
	jnot g0469(.din(w_n478_0[0]),.dout(n541),.clk(gclk));
	jnot g0470(.din(w_n511_0[0]),.dout(n542),.clk(gclk));
	jor g0471(.dina(w_n439_1[0]),.dinb(w_n404_0[1]),.dout(n543),.clk(gclk));
	jand g0472(.dina(w_n543_0[1]),.dinb(w_n445_0[0]),.dout(n544),.clk(gclk));
	jor g0473(.dina(n544),.dinb(w_n542_0[2]),.dout(n545),.clk(gclk));
	jand g0474(.dina(n545),.dinb(w_n516_0[0]),.dout(n546),.clk(gclk));
	jor g0475(.dina(n546),.dinb(w_n541_0[1]),.dout(n547),.clk(gclk));
	jand g0476(.dina(n547),.dinb(w_n483_0[0]),.dout(n548),.clk(gclk));
	jor g0477(.dina(w_n548_0[2]),.dinb(w_dff_B_TiI7vb9P6_1),.dout(w_dff_A_yKE6Pi2p6_2),.clk(gclk));
	jand g0478(.dina(w_n112_1[2]),.dinb(w_G13_0[1]),.dout(n550),.clk(gclk));
	jand g0479(.dina(w_G213_0[2]),.dinb(w_n113_1[2]),.dout(n551),.clk(gclk));
	jand g0480(.dina(n551),.dinb(w_n550_0[1]),.dout(n552),.clk(gclk));
	jand g0481(.dina(w_n552_1[1]),.dinb(w_G343_0[1]),.dout(n553),.clk(gclk));
	jnot g0482(.din(w_n553_2[2]),.dout(n554),.clk(gclk));
	jand g0483(.dina(w_n554_3[2]),.dinb(w_n524_0[0]),.dout(n555),.clk(gclk));
	jand g0484(.dina(w_n554_3[1]),.dinb(w_n528_0[0]),.dout(n556),.clk(gclk));
	jand g0485(.dina(w_n553_2[1]),.dinb(w_n367_0[0]),.dout(n557),.clk(gclk));
	jnot g0486(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jand g0487(.dina(n558),.dinb(w_n372_0[0]),.dout(n559),.clk(gclk));
	jand g0488(.dina(w_n557_0[0]),.dinb(w_n523_0[0]),.dout(n560),.clk(gclk));
	jor g0489(.dina(w_dff_B_IQmQYXWB0_0),.dinb(n559),.dout(n561),.clk(gclk));
	jand g0490(.dina(w_n561_0[2]),.dinb(w_n556_0[1]),.dout(n562),.clk(gclk));
	jor g0491(.dina(n562),.dinb(w_dff_B_76bfDyqF7_1),.dout(n563),.clk(gclk));
	jnot g0492(.din(w_n561_0[1]),.dout(n564),.clk(gclk));
	jnot g0493(.din(w_G330_0[1]),.dout(n565),.clk(gclk));
	jnot g0494(.din(w_n324_0[0]),.dout(n566),.clk(gclk));
	jor g0495(.dina(w_n554_3[0]),.dinb(w_n303_0[0]),.dout(n567),.clk(gclk));
	jnot g0496(.din(w_n567_0[1]),.dout(n568),.clk(gclk));
	jor g0497(.dina(w_dff_B_15lHvnoi4_0),.dinb(n566),.dout(n569),.clk(gclk));
	jor g0498(.dina(w_n567_0[0]),.dinb(w_n315_0[0]),.dout(n570),.clk(gclk));
	jand g0499(.dina(w_dff_B_7Q94a7311_0),.dinb(n569),.dout(n571),.clk(gclk));
	jor g0500(.dina(w_n571_0[2]),.dinb(w_n565_0[1]),.dout(n572),.clk(gclk));
	jor g0501(.dina(w_n572_0[2]),.dinb(w_n564_0[1]),.dout(n573),.clk(gclk));
	jnot g0502(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jor g0503(.dina(n574),.dinb(w_n563_0[2]),.dout(w_dff_A_TMIQp7yB0_2),.clk(gclk));
	jand g0504(.dina(w_n554_2[2]),.dinb(w_n539_0[0]),.dout(n576),.clk(gclk));
	jor g0505(.dina(w_n553_2[0]),.dinb(w_n374_0[0]),.dout(n577),.clk(gclk));
	jand g0506(.dina(w_n346_0[1]),.dinb(w_n210_0[0]),.dout(n578),.clk(gclk));
	jand g0507(.dina(n578),.dinb(w_n312_0[1]),.dout(n579),.clk(gclk));
	jand g0508(.dina(n579),.dinb(w_n534_0[0]),.dout(n580),.clk(gclk));
	jand g0509(.dina(w_n288_0[1]),.dinb(w_n196_0[2]),.dout(n581),.clk(gclk));
	jand g0510(.dina(w_n355_0[1]),.dinb(w_n246_0[1]),.dout(n582),.clk(gclk));
	jand g0511(.dina(n582),.dinb(w_n170_0[0]),.dout(n583),.clk(gclk));
	jand g0512(.dina(n583),.dinb(w_dff_B_KdKHTE9v4_1),.dout(n584),.clk(gclk));
	jor g0513(.dina(n584),.dinb(w_n554_2[1]),.dout(n585),.clk(gclk));
	jor g0514(.dina(n585),.dinb(w_dff_B_2iHUmqcd2_1),.dout(n586),.clk(gclk));
	jand g0515(.dina(n586),.dinb(w_G330_0[0]),.dout(n587),.clk(gclk));
	jand g0516(.dina(w_dff_B_Ao6zYikO0_0),.dinb(n577),.dout(n588),.clk(gclk));
	jor g0517(.dina(w_n588_1[1]),.dinb(w_n576_1[1]),.dout(n589),.clk(gclk));
	jand g0518(.dina(w_n589_1[2]),.dinb(w_n113_1[1]),.dout(n590),.clk(gclk));
	jand g0519(.dina(w_n122_1[0]),.dinb(w_n149_1[1]),.dout(n591),.clk(gclk));
	jnot g0520(.din(w_n591_1[1]),.dout(n592),.clk(gclk));
	jand g0521(.dina(w_n180_0[0]),.dinb(w_n105_1[0]),.dout(n593),.clk(gclk));
	jand g0522(.dina(w_n593_0[2]),.dinb(w_G1_1[0]),.dout(n594),.clk(gclk));
	jand g0523(.dina(n594),.dinb(w_n592_2[1]),.dout(n595),.clk(gclk));
	jand g0524(.dina(w_n591_1[0]),.dinb(w_n118_0[1]),.dout(n596),.clk(gclk));
	jor g0525(.dina(w_dff_B_30hQyZDl3_0),.dinb(n595),.dout(n597),.clk(gclk));
	jor g0526(.dina(w_dff_B_aW8cQsyk1_0),.dinb(n590),.dout(w_dff_A_0WVEvPGS5_2),.clk(gclk));
	jand g0527(.dina(w_n571_0[1]),.dinb(w_n565_0[0]),.dout(n599),.clk(gclk));
	jnot g0528(.din(n599),.dout(n600),.clk(gclk));
	jand g0529(.dina(w_n550_0[0]),.dinb(w_G45_1[0]),.dout(n601),.clk(gclk));
	jor g0530(.dina(n601),.dinb(w_n113_1[0]),.dout(n602),.clk(gclk));
	jnot g0531(.din(w_n602_0[1]),.dout(n603),.clk(gclk));
	jand g0532(.dina(w_n603_2[1]),.dinb(w_n592_2[0]),.dout(n604),.clk(gclk));
	jnot g0533(.din(w_n604_2[1]),.dout(n605),.clk(gclk));
	jand g0534(.dina(w_n605_1[2]),.dinb(w_n572_0[1]),.dout(n606),.clk(gclk));
	jand g0535(.dina(n606),.dinb(n600),.dout(n607),.clk(gclk));
	jand g0536(.dina(w_n462_0[0]),.dinb(w_n114_0[1]),.dout(n608),.clk(gclk));
	jand g0537(.dina(w_n608_1[2]),.dinb(w_n571_0[0]),.dout(n609),.clk(gclk));
	jnot g0538(.din(n609),.dout(n610),.clk(gclk));
	jand g0539(.dina(w_n146_1[0]),.dinb(w_G20_3[1]),.dout(n611),.clk(gclk));
	jor g0540(.dina(n611),.dinb(w_n115_0[1]),.dout(n612),.clk(gclk));
	jand g0541(.dina(w_G179_0[2]),.dinb(w_G20_3[0]),.dout(n613),.clk(gclk));
	jnot g0542(.din(w_n613_1[1]),.dout(n614),.clk(gclk));
	jand g0543(.dina(w_G200_2[0]),.dinb(w_G20_2[2]),.dout(n615),.clk(gclk));
	jand g0544(.dina(w_n615_0[1]),.dinb(n614),.dout(n616),.clk(gclk));
	jand g0545(.dina(w_n616_0[1]),.dinb(w_G190_2[0]),.dout(n617),.clk(gclk));
	jand g0546(.dina(w_n617_6[1]),.dinb(w_G303_2[1]),.dout(n618),.clk(gclk));
	jand g0547(.dina(w_n407_1[2]),.dinb(w_G20_2[1]),.dout(n619),.clk(gclk));
	jnot g0548(.din(w_n619_0[1]),.dout(n620),.clk(gclk));
	jor g0549(.dina(w_n615_0[0]),.dinb(w_n613_1[0]),.dout(n621),.clk(gclk));
	jnot g0550(.din(n621),.dout(n622),.clk(gclk));
	jand g0551(.dina(w_n622_0[1]),.dinb(n620),.dout(n623),.clk(gclk));
	jand g0552(.dina(w_n623_5[1]),.dinb(w_G294_3[0]),.dout(n624),.clk(gclk));
	jnot g0553(.din(w_G200_1[2]),.dout(n625),.clk(gclk));
	jand g0554(.dina(w_n613_0[2]),.dinb(n625),.dout(n626),.clk(gclk));
	jand g0555(.dina(w_n626_0[1]),.dinb(w_G190_1[2]),.dout(n627),.clk(gclk));
	jand g0556(.dina(w_n627_7[1]),.dinb(w_G322_0[2]),.dout(n628),.clk(gclk));
	jor g0557(.dina(w_dff_B_luZy6lJH8_0),.dinb(n624),.dout(n629),.clk(gclk));
	jor g0558(.dina(n629),.dinb(w_dff_B_vPKyQSuR3_1),.dout(n630),.clk(gclk));
	jand g0559(.dina(w_n622_0[0]),.dinb(w_n619_0[0]),.dout(n631),.clk(gclk));
	jand g0560(.dina(w_n631_7[1]),.dinb(w_dff_B_g3sqqxTD0_1),.dout(n632),.clk(gclk));
	jor g0561(.dina(n632),.dinb(w_n148_5[2]),.dout(n633),.clk(gclk));
	jand g0562(.dina(w_n616_0[0]),.dinb(w_n407_1[1]),.dout(n634),.clk(gclk));
	jand g0563(.dina(w_n634_4[1]),.dinb(w_G283_3[1]),.dout(n635),.clk(gclk));
	jand g0564(.dina(w_n626_0[0]),.dinb(w_n407_1[0]),.dout(n636),.clk(gclk));
	jand g0565(.dina(w_n636_7[1]),.dinb(w_G311_1[2]),.dout(n637),.clk(gclk));
	jor g0566(.dina(w_dff_B_HZGkihJZ2_0),.dinb(n635),.dout(n638),.clk(gclk));
	jand g0567(.dina(w_n613_0[1]),.dinb(w_G200_1[1]),.dout(n639),.clk(gclk));
	jand g0568(.dina(w_n639_0[1]),.dinb(w_G190_1[1]),.dout(n640),.clk(gclk));
	jand g0569(.dina(w_n640_7[1]),.dinb(w_G326_0[1]),.dout(n641),.clk(gclk));
	jand g0570(.dina(w_n639_0[0]),.dinb(w_n407_0[2]),.dout(n642),.clk(gclk));
	jand g0571(.dina(w_n642_7[1]),.dinb(w_G317_1[1]),.dout(n643),.clk(gclk));
	jor g0572(.dina(n643),.dinb(n641),.dout(n644),.clk(gclk));
	jor g0573(.dina(w_dff_B_xbbZLR3d2_0),.dinb(n638),.dout(n645),.clk(gclk));
	jor g0574(.dina(n645),.dinb(w_dff_B_YeRo1S9M1_1),.dout(n646),.clk(gclk));
	jor g0575(.dina(n646),.dinb(w_dff_B_zytjr5lS4_1),.dout(n647),.clk(gclk));
	jand g0576(.dina(w_n631_7[0]),.dinb(w_G159_3[1]),.dout(n648),.clk(gclk));
	jand g0577(.dina(w_n640_7[0]),.dinb(w_G50_4[0]),.dout(n649),.clk(gclk));
	jand g0578(.dina(w_n642_7[0]),.dinb(w_G68_3[2]),.dout(n650),.clk(gclk));
	jor g0579(.dina(n650),.dinb(n649),.dout(n651),.clk(gclk));
	jor g0580(.dina(n651),.dinb(n648),.dout(n652),.clk(gclk));
	jnot g0581(.din(n652),.dout(n653),.clk(gclk));
	jand g0582(.dina(w_n617_6[0]),.dinb(w_G87_2[1]),.dout(n654),.clk(gclk));
	jnot g0583(.din(w_n654_0[1]),.dout(n655),.clk(gclk));
	jand g0584(.dina(n655),.dinb(w_n148_5[1]),.dout(n656),.clk(gclk));
	jand g0585(.dina(w_n634_4[0]),.dinb(w_G107_3[1]),.dout(n657),.clk(gclk));
	jand g0586(.dina(w_n636_7[0]),.dinb(w_G77_3[1]),.dout(n658),.clk(gclk));
	jor g0587(.dina(w_dff_B_fNJBprkP0_0),.dinb(w_n657_0[1]),.dout(n659),.clk(gclk));
	jand g0588(.dina(w_n627_7[0]),.dinb(w_G58_3[2]),.dout(n660),.clk(gclk));
	jand g0589(.dina(w_n623_5[0]),.dinb(w_G97_3[1]),.dout(n661),.clk(gclk));
	jor g0590(.dina(w_n661_0[1]),.dinb(w_dff_B_cnEI5OKQ2_1),.dout(n662),.clk(gclk));
	jor g0591(.dina(n662),.dinb(n659),.dout(n663),.clk(gclk));
	jnot g0592(.din(n663),.dout(n664),.clk(gclk));
	jand g0593(.dina(n664),.dinb(w_dff_B_NFw4p7kh4_1),.dout(n665),.clk(gclk));
	jand g0594(.dina(n665),.dinb(w_dff_B_JOmrejZn1_1),.dout(n666),.clk(gclk));
	jnot g0595(.din(n666),.dout(n667),.clk(gclk));
	jand g0596(.dina(n667),.dinb(w_dff_B_SollERH45_1),.dout(n668),.clk(gclk));
	jor g0597(.dina(n668),.dinb(w_n612_4[1]),.dout(n669),.clk(gclk));
	jnot g0598(.din(w_n608_1[1]),.dout(n670),.clk(gclk));
	jand g0599(.dina(w_n612_4[0]),.dinb(n670),.dout(n671),.clk(gclk));
	jnot g0600(.din(n671),.dout(n672),.clk(gclk));
	jand g0601(.dina(w_n140_0[0]),.dinb(w_G45_0[2]),.dout(n673),.clk(gclk));
	jand g0602(.dina(w_n118_0[0]),.dinb(w_n161_0[2]),.dout(n674),.clk(gclk));
	jand g0603(.dina(w_n122_0[2]),.dinb(w_G33_6[1]),.dout(n675),.clk(gclk));
	jnot g0604(.din(w_n675_0[2]),.dout(n676),.clk(gclk));
	jor g0605(.dina(w_n676_0[1]),.dinb(n674),.dout(n677),.clk(gclk));
	jor g0606(.dina(n677),.dinb(w_dff_B_q8O96NZW0_1),.dout(n678),.clk(gclk));
	jand g0607(.dina(w_n123_1[1]),.dinb(w_n105_0[2]),.dout(n679),.clk(gclk));
	jand g0608(.dina(w_n122_0[1]),.dinb(w_n148_5[0]),.dout(n680),.clk(gclk));
	jand g0609(.dina(w_n680_0[1]),.dinb(w_G355_0),.dout(n681),.clk(gclk));
	jor g0610(.dina(n681),.dinb(w_dff_B_PrSaw47k1_1),.dout(n682),.clk(gclk));
	jnot g0611(.din(n682),.dout(n683),.clk(gclk));
	jand g0612(.dina(n683),.dinb(w_dff_B_TgwTAz0T8_1),.dout(n684),.clk(gclk));
	jor g0613(.dina(n684),.dinb(w_n672_1[1]),.dout(n685),.clk(gclk));
	jand g0614(.dina(n685),.dinb(w_n604_2[0]),.dout(n686),.clk(gclk));
	jand g0615(.dina(w_dff_B_ijCClu5V1_0),.dinb(n669),.dout(n687),.clk(gclk));
	jand g0616(.dina(w_dff_B_pbid71fM7_0),.dinb(n610),.dout(n688),.clk(gclk));
	jor g0617(.dina(n688),.dinb(n607),.dout(G396_fa_),.clk(gclk));
	jnot g0618(.din(w_n588_1[0]),.dout(n690),.clk(gclk));
	jnot g0619(.din(w_n401_0[0]),.dout(n691),.clk(gclk));
	jor g0620(.dina(w_n554_2[0]),.dinb(n691),.dout(n692),.clk(gclk));
	jand g0621(.dina(w_n692_0[1]),.dinb(w_n412_0[0]),.dout(n693),.clk(gclk));
	jor g0622(.dina(w_n692_0[0]),.dinb(w_n405_0[0]),.dout(n694),.clk(gclk));
	jnot g0623(.din(n694),.dout(n695),.clk(gclk));
	jor g0624(.dina(n695),.dinb(n693),.dout(n696),.clk(gclk));
	jxor g0625(.dina(w_n696_1[2]),.dinb(w_n576_1[0]),.dout(n697),.clk(gclk));
	jnot g0626(.din(n697),.dout(n698),.clk(gclk));
	jand g0627(.dina(n698),.dinb(w_dff_B_q5AGVv120_1),.dout(n699),.clk(gclk));
	jor g0628(.dina(w_n991_0[2]),.dinb(w_n604_1[2]),.dout(n701),.clk(gclk));
	jor g0629(.dina(w_dff_B_ToFRmcGQ2_0),.dinb(n699),.dout(n702),.clk(gclk));
	jnot g0630(.din(w_n696_1[1]),.dout(n703),.clk(gclk));
	jand g0631(.dina(n703),.dinb(w_n425_1[1]),.dout(n704),.clk(gclk));
	jnot g0632(.din(n704),.dout(n705),.clk(gclk));
	jand g0633(.dina(w_n631_6[2]),.dinb(w_G132_1[1]),.dout(n706),.clk(gclk));
	jand g0634(.dina(w_n623_4[2]),.dinb(w_G58_3[1]),.dout(n707),.clk(gclk));
	jand g0635(.dina(w_n642_6[2]),.dinb(w_G150_3[0]),.dout(n708),.clk(gclk));
	jor g0636(.dina(w_dff_B_h2dKfwho3_0),.dinb(n707),.dout(n709),.clk(gclk));
	jor g0637(.dina(n709),.dinb(w_dff_B_y90EBVFx6_1),.dout(n710),.clk(gclk));
	jand g0638(.dina(w_n617_5[2]),.dinb(w_G50_3[2]),.dout(n711),.clk(gclk));
	jor g0639(.dina(n711),.dinb(w_G33_6[0]),.dout(n712),.clk(gclk));
	jand g0640(.dina(w_n636_6[2]),.dinb(w_G159_3[0]),.dout(n713),.clk(gclk));
	jand g0641(.dina(w_n627_6[2]),.dinb(w_G143_2[1]),.dout(n714),.clk(gclk));
	jor g0642(.dina(n714),.dinb(n713),.dout(n715),.clk(gclk));
	jand g0643(.dina(w_n640_6[2]),.dinb(w_G137_1[2]),.dout(n716),.clk(gclk));
	jand g0644(.dina(w_n634_3[2]),.dinb(w_G68_3[1]),.dout(n717),.clk(gclk));
	jor g0645(.dina(w_n717_0[1]),.dinb(w_dff_B_2WoV4lU33_1),.dout(n718),.clk(gclk));
	jor g0646(.dina(n718),.dinb(w_dff_B_mA1TS2tU5_1),.dout(n719),.clk(gclk));
	jor g0647(.dina(n719),.dinb(w_dff_B_qOHNn4DT0_1),.dout(n720),.clk(gclk));
	jor g0648(.dina(n720),.dinb(w_dff_B_0Qpqs9IT5_1),.dout(n721),.clk(gclk));
	jand g0649(.dina(w_n631_6[1]),.dinb(w_G311_1[1]),.dout(n722),.clk(gclk));
	jand g0650(.dina(w_n617_5[1]),.dinb(w_G107_3[0]),.dout(n723),.clk(gclk));
	jand g0651(.dina(w_n642_6[1]),.dinb(w_G283_3[0]),.dout(n724),.clk(gclk));
	jor g0652(.dina(w_dff_B_kbc6CHlm6_0),.dinb(n723),.dout(n725),.clk(gclk));
	jor g0653(.dina(n725),.dinb(w_dff_B_IAYrVm0P9_1),.dout(n726),.clk(gclk));
	jnot g0654(.din(n726),.dout(n727),.clk(gclk));
	jand g0655(.dina(w_n634_3[1]),.dinb(w_G87_2[0]),.dout(n728),.clk(gclk));
	jnot g0656(.din(w_n728_0[1]),.dout(n729),.clk(gclk));
	jand g0657(.dina(n729),.dinb(w_G33_5[2]),.dout(n730),.clk(gclk));
	jand g0658(.dina(w_n636_6[1]),.dinb(w_G116_3[2]),.dout(n731),.clk(gclk));
	jand g0659(.dina(w_n627_6[1]),.dinb(w_G294_2[2]),.dout(n732),.clk(gclk));
	jor g0660(.dina(n732),.dinb(n731),.dout(n733),.clk(gclk));
	jand g0661(.dina(w_n640_6[1]),.dinb(w_G303_2[0]),.dout(n734),.clk(gclk));
	jor g0662(.dina(w_dff_B_ZNVwHKRe3_0),.dinb(w_n661_0[0]),.dout(n735),.clk(gclk));
	jor g0663(.dina(n735),.dinb(w_dff_B_ZxTVggiG3_1),.dout(n736),.clk(gclk));
	jnot g0664(.din(n736),.dout(n737),.clk(gclk));
	jand g0665(.dina(n737),.dinb(w_dff_B_iyLyyVWW7_1),.dout(n738),.clk(gclk));
	jand g0666(.dina(n738),.dinb(w_dff_B_aEOYgQuj1_1),.dout(n739),.clk(gclk));
	jnot g0667(.din(n739),.dout(n740),.clk(gclk));
	jand g0668(.dina(n740),.dinb(w_dff_B_kltxwDtL7_1),.dout(n741),.clk(gclk));
	jor g0669(.dina(n741),.dinb(w_n612_3[2]),.dout(n742),.clk(gclk));
	jand g0670(.dina(w_n612_3[1]),.dinb(w_n426_0[0]),.dout(n743),.clk(gclk));
	jand g0671(.dina(w_n743_1[1]),.dinb(w_n72_0[1]),.dout(n744),.clk(gclk));
	jor g0672(.dina(w_dff_B_huqK92bP3_0),.dinb(w_n605_1[1]),.dout(n745),.clk(gclk));
	jnot g0673(.din(n745),.dout(n746),.clk(gclk));
	jand g0674(.dina(w_dff_B_QLeR7zmG1_0),.dinb(n742),.dout(n747),.clk(gclk));
	jand g0675(.dina(w_dff_B_SfEUcmPy1_0),.dinb(n705),.dout(n748),.clk(gclk));
	jnot g0676(.din(n748),.dout(n749),.clk(gclk));
	jand g0677(.dina(n749),.dinb(n702),.dout(n750),.clk(gclk));
	jnot g0678(.din(w_n750_0[1]),.dout(G384_fa_),.clk(gclk));
	jnot g0679(.din(w_n552_1[0]),.dout(n752),.clk(gclk));
	jand g0680(.dina(w_dff_B_Au4qUoU05_0),.dinb(w_n542_0[1]),.dout(n753),.clk(gclk));
	jand g0681(.dina(w_n552_0[2]),.dinb(w_n512_0[0]),.dout(n754),.clk(gclk));
	jnot g0682(.din(w_n754_0[1]),.dout(n755),.clk(gclk));
	jand g0683(.dina(n755),.dinb(w_n517_0[0]),.dout(n756),.clk(gclk));
	jand g0684(.dina(w_n754_0[0]),.dinb(w_n542_0[0]),.dout(n757),.clk(gclk));
	jor g0685(.dina(n757),.dinb(n756),.dout(n758),.clk(gclk));
	jand g0686(.dina(w_n696_1[0]),.dinb(w_n576_0[2]),.dout(n759),.clk(gclk));
	jand g0687(.dina(w_n553_1[2]),.dinb(w_n436_0[0]),.dout(n760),.clk(gclk));
	jnot g0688(.din(w_n760_0[1]),.dout(n761),.clk(gclk));
	jand g0689(.dina(w_dff_B_0Jc9uF4g1_0),.dinb(w_n446_0[0]),.dout(n762),.clk(gclk));
	jand g0690(.dina(w_n760_0[0]),.dinb(w_n439_0[2]),.dout(n763),.clk(gclk));
	jor g0691(.dina(w_dff_B_HkOfbMn44_0),.dinb(n762),.dout(n764),.clk(gclk));
	jand g0692(.dina(w_n764_1[2]),.dinb(w_n759_0[1]),.dout(n765),.clk(gclk));
	jor g0693(.dina(w_n764_1[1]),.dinb(w_n439_0[1]),.dout(n766),.clk(gclk));
	jand g0694(.dina(w_n554_1[2]),.dinb(w_n543_0[0]),.dout(n767),.clk(gclk));
	jand g0695(.dina(w_dff_B_YDYslqhf5_0),.dinb(n766),.dout(n768),.clk(gclk));
	jor g0696(.dina(w_dff_B_BXD6qlQV4_0),.dinb(n765),.dout(n769),.clk(gclk));
	jand g0697(.dina(w_n769_0[1]),.dinb(w_n758_1[1]),.dout(n770),.clk(gclk));
	jor g0698(.dina(n770),.dinb(w_dff_B_vGoV2cZb0_1),.dout(n771),.clk(gclk));
	jnot g0699(.din(w_n771_0[2]),.dout(n772),.clk(gclk));
	jand g0700(.dina(w_n576_0[1]),.dinb(w_n519_1[0]),.dout(n773),.clk(gclk));
	jor g0701(.dina(n773),.dinb(w_n548_0[1]),.dout(n774),.clk(gclk));
	jand g0702(.dina(w_n764_1[0]),.dinb(w_n696_0[2]),.dout(n775),.clk(gclk));
	jand g0703(.dina(n775),.dinb(w_n758_1[0]),.dout(n776),.clk(gclk));
	jxor g0704(.dina(n776),.dinb(w_n519_0[2]),.dout(n777),.clk(gclk));
	jand g0705(.dina(n777),.dinb(w_n588_0[2]),.dout(n778),.clk(gclk));
	jxor g0706(.dina(n778),.dinb(w_dff_B_ismogaiY2_1),.dout(n779),.clk(gclk));
	jnot g0707(.din(w_n779_0[1]),.dout(n780),.clk(gclk));
	jor g0708(.dina(w_dff_B_INXKO3Aj0_0),.dinb(n772),.dout(n781),.clk(gclk));
	jor g0709(.dina(w_n779_0[0]),.dinb(w_n771_0[1]),.dout(n782),.clk(gclk));
	jnot g0710(.din(w_n121_0[1]),.dout(n783),.clk(gclk));
	jand g0711(.dina(n783),.dinb(w_n116_0[0]),.dout(n784),.clk(gclk));
	jand g0712(.dina(w_dff_B_Q1LIwqe58_0),.dinb(n782),.dout(n785),.clk(gclk));
	jand g0713(.dina(n785),.dinb(n781),.dout(n786),.clk(gclk));
	jand g0714(.dina(w_G77_3[0]),.dinb(w_G50_3[1]),.dout(n787),.clk(gclk));
	jand g0715(.dina(n787),.dinb(w_n137_0[0]),.dout(n788),.clk(gclk));
	jand g0716(.dina(w_G68_3[0]),.dinb(w_n73_1[2]),.dout(n789),.clk(gclk));
	jor g0717(.dina(n789),.dinb(n788),.dout(n790),.clk(gclk));
	jand g0718(.dina(n790),.dinb(w_n121_0[0]),.dout(n791),.clk(gclk));
	jnot g0719(.din(w_n255_0[0]),.dout(n792),.clk(gclk));
	jand g0720(.dina(w_n147_0[0]),.dinb(w_G116_3[1]),.dout(n793),.clk(gclk));
	jand g0721(.dina(w_dff_B_oaMhJkbn7_0),.dinb(n792),.dout(n794),.clk(gclk));
	jor g0722(.dina(n794),.dinb(w_dff_B_S17TyMTG2_1),.dout(n795),.clk(gclk));
	jor g0723(.dina(w_dff_B_iHgZDsFN1_0),.dinb(n786),.dout(w_dff_A_OjXgsc6F9_2),.clk(gclk));
	jand g0724(.dina(w_n553_1[1]),.dinb(w_n214_0[0]),.dout(n797),.clk(gclk));
	jnot g0725(.din(w_n797_0[1]),.dout(n798),.clk(gclk));
	jand g0726(.dina(w_dff_B_O0aVY1Bz7_0),.dinb(w_n219_0[0]),.dout(n799),.clk(gclk));
	jand g0727(.dina(w_n797_0[0]),.dinb(w_n532_0[0]),.dout(n800),.clk(gclk));
	jor g0728(.dina(w_dff_B_N4HDd12h4_0),.dinb(n799),.dout(n801),.clk(gclk));
	jnot g0729(.din(w_n801_0[1]),.dout(n802),.clk(gclk));
	jand g0730(.dina(n802),.dinb(w_n608_1[0]),.dout(n803),.clk(gclk));
	jnot g0731(.din(n803),.dout(n804),.clk(gclk));
	jand g0732(.dina(w_n631_6[0]),.dinb(w_G317_1[0]),.dout(n805),.clk(gclk));
	jand g0733(.dina(w_n623_4[1]),.dinb(w_G107_2[2]),.dout(n806),.clk(gclk));
	jand g0734(.dina(w_n642_6[0]),.dinb(w_G294_2[1]),.dout(n807),.clk(gclk));
	jor g0735(.dina(w_dff_B_5f1pzdeI0_0),.dinb(n806),.dout(n808),.clk(gclk));
	jor g0736(.dina(n808),.dinb(w_dff_B_liQ1UMAM7_1),.dout(n809),.clk(gclk));
	jand g0737(.dina(w_n617_5[0]),.dinb(w_G116_3[0]),.dout(n810),.clk(gclk));
	jor g0738(.dina(n810),.dinb(w_n148_4[2]),.dout(n811),.clk(gclk));
	jand g0739(.dina(w_n636_6[0]),.dinb(w_G283_2[2]),.dout(n812),.clk(gclk));
	jand g0740(.dina(w_n627_6[0]),.dinb(w_G303_1[2]),.dout(n813),.clk(gclk));
	jor g0741(.dina(n813),.dinb(n812),.dout(n814),.clk(gclk));
	jand g0742(.dina(w_n640_6[0]),.dinb(w_G311_1[0]),.dout(n815),.clk(gclk));
	jand g0743(.dina(w_n634_3[0]),.dinb(w_G97_3[0]),.dout(n816),.clk(gclk));
	jor g0744(.dina(w_n816_0[1]),.dinb(w_dff_B_LAJJ92v23_1),.dout(n817),.clk(gclk));
	jor g0745(.dina(n817),.dinb(w_dff_B_TTOk1bak3_1),.dout(n818),.clk(gclk));
	jor g0746(.dina(n818),.dinb(w_dff_B_kG1WRgHS8_1),.dout(n819),.clk(gclk));
	jor g0747(.dina(n819),.dinb(w_dff_B_qpC0aZAa8_1),.dout(n820),.clk(gclk));
	jand g0748(.dina(w_n631_5[2]),.dinb(w_G137_1[1]),.dout(n821),.clk(gclk));
	jnot g0749(.din(n821),.dout(n822),.clk(gclk));
	jand g0750(.dina(w_n623_4[0]),.dinb(w_G68_2[2]),.dout(n823),.clk(gclk));
	jnot g0751(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jand g0752(.dina(w_n634_2[2]),.dinb(w_G77_2[2]),.dout(n825),.clk(gclk));
	jnot g0753(.din(w_n825_0[1]),.dout(n826),.clk(gclk));
	jand g0754(.dina(n826),.dinb(n824),.dout(n827),.clk(gclk));
	jand g0755(.dina(n827),.dinb(w_dff_B_Xkqgtt0R2_1),.dout(n828),.clk(gclk));
	jand g0756(.dina(w_n642_5[2]),.dinb(w_G159_2[2]),.dout(n829),.clk(gclk));
	jor g0757(.dina(n829),.dinb(w_G33_5[1]),.dout(n830),.clk(gclk));
	jand g0758(.dina(w_n640_5[2]),.dinb(w_G143_2[0]),.dout(n831),.clk(gclk));
	jand g0759(.dina(w_n627_5[2]),.dinb(w_G150_2[2]),.dout(n832),.clk(gclk));
	jor g0760(.dina(n832),.dinb(n831),.dout(n833),.clk(gclk));
	jand g0761(.dina(w_n636_5[2]),.dinb(w_G50_3[0]),.dout(n834),.clk(gclk));
	jand g0762(.dina(w_n617_4[2]),.dinb(w_G58_3[0]),.dout(n835),.clk(gclk));
	jor g0763(.dina(n835),.dinb(w_dff_B_GOaq4DFZ9_1),.dout(n836),.clk(gclk));
	jor g0764(.dina(n836),.dinb(w_dff_B_KfVTBMJA0_1),.dout(n837),.clk(gclk));
	jor g0765(.dina(n837),.dinb(w_dff_B_l1n21D5a6_1),.dout(n838),.clk(gclk));
	jnot g0766(.din(n838),.dout(n839),.clk(gclk));
	jand g0767(.dina(n839),.dinb(w_dff_B_tafiDLO83_1),.dout(n840),.clk(gclk));
	jnot g0768(.din(n840),.dout(n841),.clk(gclk));
	jand g0769(.dina(n841),.dinb(w_dff_B_9EpyEEZg7_1),.dout(n842),.clk(gclk));
	jor g0770(.dina(n842),.dinb(w_n612_3[0]),.dout(n843),.clk(gclk));
	jand g0771(.dina(w_n675_0[1]),.dinb(w_n131_0[0]),.dout(n844),.clk(gclk));
	jand g0772(.dina(w_n123_1[0]),.dinb(w_G87_1[2]),.dout(n845),.clk(gclk));
	jor g0773(.dina(w_dff_B_cNBDWlkf7_0),.dinb(w_n672_1[0]),.dout(n846),.clk(gclk));
	jor g0774(.dina(n846),.dinb(w_dff_B_EkAG2G5A5_1),.dout(n847),.clk(gclk));
	jand g0775(.dina(n847),.dinb(w_n604_1[1]),.dout(n848),.clk(gclk));
	jand g0776(.dina(w_dff_B_XK9Rr1Md4_0),.dinb(n843),.dout(n849),.clk(gclk));
	jand g0777(.dina(w_dff_B_vakdpU0h4_0),.dinb(n804),.dout(n850),.clk(gclk));
	jnot g0778(.din(w_n589_1[1]),.dout(n851),.clk(gclk));
	jxor g0779(.dina(w_n561_0[0]),.dinb(w_n556_0[0]),.dout(n852),.clk(gclk));
	jxor g0780(.dina(w_dff_B_SYCE2BTn7_0),.dinb(w_n572_0[0]),.dout(n853),.clk(gclk));
	jnot g0781(.din(w_n853_0[2]),.dout(n854),.clk(gclk));
	jand g0782(.dina(n854),.dinb(n851),.dout(n855),.clk(gclk));
	jnot g0783(.din(w_n278_0[0]),.dout(n856),.clk(gclk));
	jand g0784(.dina(w_n553_1[0]),.dinb(w_n274_0[0]),.dout(n857),.clk(gclk));
	jor g0785(.dina(w_dff_B_WuxO66pk5_0),.dinb(n856),.dout(n858),.clk(gclk));
	jand g0786(.dina(w_n553_0[2]),.dinb(w_n536_0[1]),.dout(n859),.clk(gclk));
	jnot g0787(.din(n859),.dout(n860),.clk(gclk));
	jand g0788(.dina(w_dff_B_2jr7qtF45_0),.dinb(n858),.dout(n861),.clk(gclk));
	jxor g0789(.dina(w_n861_1[1]),.dinb(w_n573_0[1]),.dout(n862),.clk(gclk));
	jxor g0790(.dina(n862),.dinb(w_n563_0[1]),.dout(n863),.clk(gclk));
	jand g0791(.dina(w_n863_0[1]),.dinb(w_n855_0[2]),.dout(n864),.clk(gclk));
	jor g0792(.dina(w_n864_0[1]),.dinb(w_n589_1[0]),.dout(n865),.clk(gclk));
	jand g0793(.dina(n865),.dinb(w_n591_0[2]),.dout(n866),.clk(gclk));
	jor g0794(.dina(n866),.dinb(w_n602_0[0]),.dout(n867),.clk(gclk));
	jand g0795(.dina(w_n554_1[1]),.dinb(w_n536_0[0]),.dout(n868),.clk(gclk));
	jnot g0796(.din(w_n861_1[0]),.dout(n869),.clk(gclk));
	jand g0797(.dina(n869),.dinb(w_n563_0[0]),.dout(n870),.clk(gclk));
	jor g0798(.dina(n870),.dinb(w_dff_B_8swdFZdK9_1),.dout(n871),.clk(gclk));
	jor g0799(.dina(w_n861_0[2]),.dinb(w_n573_0[0]),.dout(n872),.clk(gclk));
	jxor g0800(.dina(n872),.dinb(w_n801_0[0]),.dout(n873),.clk(gclk));
	jxor g0801(.dina(n873),.dinb(w_dff_B_6Fz6g5cU3_1),.dout(n874),.clk(gclk));
	jnot g0802(.din(n874),.dout(n875),.clk(gclk));
	jand g0803(.dina(w_dff_B_roZoaxUK5_0),.dinb(n867),.dout(n876),.clk(gclk));
	jor g0804(.dina(n876),.dinb(w_dff_B_eRk8zz767_1),.dout(G387_fa_),.clk(gclk));
	jand g0805(.dina(w_n853_0[1]),.dinb(w_n589_0[2]),.dout(n878),.clk(gclk));
	jor g0806(.dina(w_n855_0[1]),.dinb(w_n592_1[2]),.dout(n879),.clk(gclk));
	jor g0807(.dina(n879),.dinb(w_dff_B_CQS8NZev0_1),.dout(n880),.clk(gclk));
	jor g0808(.dina(w_n853_0[0]),.dinb(w_n603_2[0]),.dout(n881),.clk(gclk));
	jand g0809(.dina(w_n608_0[2]),.dinb(w_n564_0[0]),.dout(n882),.clk(gclk));
	jand g0810(.dina(w_n631_5[1]),.dinb(w_G326_0[0]),.dout(n883),.clk(gclk));
	jand g0811(.dina(w_n623_3[2]),.dinb(w_G283_2[1]),.dout(n884),.clk(gclk));
	jand g0812(.dina(w_n627_5[1]),.dinb(w_G317_0[2]),.dout(n885),.clk(gclk));
	jor g0813(.dina(w_dff_B_ArWb2Guz8_0),.dinb(n884),.dout(n886),.clk(gclk));
	jor g0814(.dina(n886),.dinb(w_dff_B_C8F25GoX1_1),.dout(n887),.clk(gclk));
	jand g0815(.dina(w_n617_4[1]),.dinb(w_G294_2[0]),.dout(n888),.clk(gclk));
	jor g0816(.dina(n888),.dinb(w_n148_4[1]),.dout(n889),.clk(gclk));
	jand g0817(.dina(w_n634_2[1]),.dinb(w_G116_2[2]),.dout(n890),.clk(gclk));
	jand g0818(.dina(w_n636_5[1]),.dinb(w_G303_1[1]),.dout(n891),.clk(gclk));
	jor g0819(.dina(w_dff_B_oAB1G1BA4_0),.dinb(n890),.dout(n892),.clk(gclk));
	jand g0820(.dina(w_n640_5[1]),.dinb(w_G322_0[1]),.dout(n893),.clk(gclk));
	jand g0821(.dina(w_n642_5[1]),.dinb(w_G311_0[2]),.dout(n894),.clk(gclk));
	jor g0822(.dina(n894),.dinb(n893),.dout(n895),.clk(gclk));
	jor g0823(.dina(w_dff_B_ijOsRv3d3_0),.dinb(n892),.dout(n896),.clk(gclk));
	jor g0824(.dina(n896),.dinb(w_dff_B_t8HqBvIk0_1),.dout(n897),.clk(gclk));
	jor g0825(.dina(n897),.dinb(w_dff_B_s3dYIOLe0_1),.dout(n898),.clk(gclk));
	jand g0826(.dina(w_n623_3[1]),.dinb(w_G87_1[1]),.dout(n899),.clk(gclk));
	jand g0827(.dina(w_n642_5[0]),.dinb(w_G58_2[2]),.dout(n900),.clk(gclk));
	jor g0828(.dina(w_dff_B_fkrlfE7F9_0),.dinb(w_n816_0[0]),.dout(n901),.clk(gclk));
	jor g0829(.dina(n901),.dinb(w_n899_0[1]),.dout(n902),.clk(gclk));
	jand g0830(.dina(w_n631_5[0]),.dinb(w_G150_2[1]),.dout(n903),.clk(gclk));
	jor g0831(.dina(n903),.dinb(w_G33_5[0]),.dout(n904),.clk(gclk));
	jand g0832(.dina(w_n640_5[0]),.dinb(w_G159_2[1]),.dout(n905),.clk(gclk));
	jand g0833(.dina(w_n636_5[0]),.dinb(w_G68_2[1]),.dout(n906),.clk(gclk));
	jor g0834(.dina(n906),.dinb(n905),.dout(n907),.clk(gclk));
	jand g0835(.dina(w_n627_5[0]),.dinb(w_G50_2[2]),.dout(n908),.clk(gclk));
	jand g0836(.dina(w_n617_4[0]),.dinb(w_G77_2[1]),.dout(n909),.clk(gclk));
	jor g0837(.dina(w_n909_0[1]),.dinb(w_dff_B_ywfEaQGJ9_1),.dout(n910),.clk(gclk));
	jor g0838(.dina(n910),.dinb(w_dff_B_40pmEBcG8_1),.dout(n911),.clk(gclk));
	jor g0839(.dina(n911),.dinb(w_dff_B_dTs5iTOn6_1),.dout(n912),.clk(gclk));
	jor g0840(.dina(n912),.dinb(w_dff_B_y8ZMZmyl1_1),.dout(n913),.clk(gclk));
	jand g0841(.dina(n913),.dinb(n898),.dout(n914),.clk(gclk));
	jor g0842(.dina(n914),.dinb(w_n612_2[2]),.dout(n915),.clk(gclk));
	jand g0843(.dina(w_n135_0[0]),.dinb(w_G45_0[1]),.dout(n916),.clk(gclk));
	jand g0844(.dina(w_G77_2[0]),.dinb(w_G68_2[0]),.dout(n917),.clk(gclk));
	jnot g0845(.din(n917),.dout(n918),.clk(gclk));
	jand g0846(.dina(w_G58_2[1]),.dinb(w_n161_0[1]),.dout(n919),.clk(gclk));
	jand g0847(.dina(n919),.dinb(w_n73_1[1]),.dout(n920),.clk(gclk));
	jand g0848(.dina(n920),.dinb(w_dff_B_1EorlipC6_1),.dout(n921),.clk(gclk));
	jand g0849(.dina(n921),.dinb(w_n593_0[1]),.dout(n922),.clk(gclk));
	jor g0850(.dina(n922),.dinb(w_n676_0[0]),.dout(n923),.clk(gclk));
	jor g0851(.dina(n923),.dinb(w_dff_B_YfOZGs5a8_1),.dout(n924),.clk(gclk));
	jand g0852(.dina(w_n123_0[2]),.dinb(w_n80_0[1]),.dout(n925),.clk(gclk));
	jnot g0853(.din(w_n593_0[0]),.dout(n926),.clk(gclk));
	jand g0854(.dina(w_n680_0[0]),.dinb(n926),.dout(n927),.clk(gclk));
	jor g0855(.dina(n927),.dinb(w_dff_B_l03SnlX31_1),.dout(n928),.clk(gclk));
	jnot g0856(.din(n928),.dout(n929),.clk(gclk));
	jand g0857(.dina(n929),.dinb(w_dff_B_lUDGU5Tm8_1),.dout(n930),.clk(gclk));
	jor g0858(.dina(n930),.dinb(w_n672_0[2]),.dout(n931),.clk(gclk));
	jand g0859(.dina(n931),.dinb(w_n604_1[0]),.dout(n932),.clk(gclk));
	jand g0860(.dina(n932),.dinb(n915),.dout(n933),.clk(gclk));
	jnot g0861(.din(n933),.dout(n934),.clk(gclk));
	jor g0862(.dina(w_dff_B_Nw4q9f9k2_0),.dinb(n882),.dout(n935),.clk(gclk));
	jand g0863(.dina(w_dff_B_VXjngd2T1_0),.dinb(n881),.dout(n936),.clk(gclk));
	jand g0864(.dina(w_dff_B_afRYyTAp2_0),.dinb(n880),.dout(n937),.clk(gclk));
	jnot g0865(.din(w_n937_0[2]),.dout(w_dff_A_6AG3SgwF9_1),.clk(gclk));
	jnot g0866(.din(w_n855_0[0]),.dout(n939),.clk(gclk));
	jnot g0867(.din(w_n863_0[0]),.dout(n940),.clk(gclk));
	jand g0868(.dina(w_n940_0[1]),.dinb(n939),.dout(n941),.clk(gclk));
	jor g0869(.dina(w_n864_0[0]),.dinb(w_n592_1[1]),.dout(n942),.clk(gclk));
	jor g0870(.dina(n942),.dinb(n941),.dout(n943),.clk(gclk));
	jor g0871(.dina(w_n940_0[0]),.dinb(w_n603_1[2]),.dout(n944),.clk(gclk));
	jand g0872(.dina(w_n861_0[1]),.dinb(w_n608_0[1]),.dout(n945),.clk(gclk));
	jnot g0873(.din(n945),.dout(n946),.clk(gclk));
	jand g0874(.dina(w_n623_3[0]),.dinb(w_G116_2[1]),.dout(n947),.clk(gclk));
	jand g0875(.dina(w_n617_3[2]),.dinb(w_G283_2[0]),.dout(n948),.clk(gclk));
	jand g0876(.dina(w_n642_4[2]),.dinb(w_G303_1[0]),.dout(n949),.clk(gclk));
	jor g0877(.dina(w_dff_B_8j7u9TlS3_0),.dinb(n948),.dout(n950),.clk(gclk));
	jor g0878(.dina(n950),.dinb(w_dff_B_AOeF9rv66_1),.dout(n951),.clk(gclk));
	jand g0879(.dina(w_n631_4[2]),.dinb(w_G322_0[0]),.dout(n952),.clk(gclk));
	jor g0880(.dina(n952),.dinb(w_n148_4[0]),.dout(n953),.clk(gclk));
	jand g0881(.dina(w_n636_4[2]),.dinb(w_G294_1[2]),.dout(n954),.clk(gclk));
	jand g0882(.dina(w_n627_4[2]),.dinb(w_G311_0[1]),.dout(n955),.clk(gclk));
	jor g0883(.dina(n955),.dinb(n954),.dout(n956),.clk(gclk));
	jand g0884(.dina(w_n640_4[2]),.dinb(w_G317_0[1]),.dout(n957),.clk(gclk));
	jor g0885(.dina(w_dff_B_VJfuxWIR1_0),.dinb(w_n657_0[0]),.dout(n958),.clk(gclk));
	jor g0886(.dina(n958),.dinb(w_dff_B_ByV9zlj97_1),.dout(n959),.clk(gclk));
	jor g0887(.dina(n959),.dinb(w_dff_B_OhcYGMIq1_1),.dout(n960),.clk(gclk));
	jor g0888(.dina(n960),.dinb(w_dff_B_HzyL4HYi9_1),.dout(n961),.clk(gclk));
	jand g0889(.dina(w_n623_2[2]),.dinb(w_G77_1[2]),.dout(n962),.clk(gclk));
	jand g0890(.dina(w_n617_3[1]),.dinb(w_G68_1[2]),.dout(n963),.clk(gclk));
	jand g0891(.dina(w_n642_4[1]),.dinb(w_G50_2[1]),.dout(n964),.clk(gclk));
	jor g0892(.dina(w_dff_B_QnFifl5M3_0),.dinb(n963),.dout(n965),.clk(gclk));
	jor g0893(.dina(n965),.dinb(w_n962_0[1]),.dout(n966),.clk(gclk));
	jand g0894(.dina(w_n631_4[1]),.dinb(w_G143_1[2]),.dout(n967),.clk(gclk));
	jor g0895(.dina(n967),.dinb(w_G33_4[2]),.dout(n968),.clk(gclk));
	jand g0896(.dina(w_n636_4[1]),.dinb(w_G58_2[0]),.dout(n969),.clk(gclk));
	jand g0897(.dina(w_n627_4[1]),.dinb(w_G159_2[0]),.dout(n970),.clk(gclk));
	jor g0898(.dina(n970),.dinb(n969),.dout(n971),.clk(gclk));
	jand g0899(.dina(w_n640_4[1]),.dinb(w_G150_2[0]),.dout(n972),.clk(gclk));
	jor g0900(.dina(w_dff_B_q2pNGgEz9_0),.dinb(w_n728_0[0]),.dout(n973),.clk(gclk));
	jor g0901(.dina(n973),.dinb(w_dff_B_WnjYk9sv3_1),.dout(n974),.clk(gclk));
	jor g0902(.dina(n974),.dinb(w_dff_B_whVeXqgD6_1),.dout(n975),.clk(gclk));
	jor g0903(.dina(n975),.dinb(w_dff_B_ywj6lkni5_1),.dout(n976),.clk(gclk));
	jand g0904(.dina(n976),.dinb(n961),.dout(n977),.clk(gclk));
	jor g0905(.dina(n977),.dinb(w_n612_2[1]),.dout(n978),.clk(gclk));
	jand g0906(.dina(w_n675_0[0]),.dinb(w_n144_0[0]),.dout(n979),.clk(gclk));
	jand g0907(.dina(w_n123_0[1]),.dinb(w_G97_2[2]),.dout(n980),.clk(gclk));
	jor g0908(.dina(w_dff_B_Lb7neYNf5_0),.dinb(w_n672_0[1]),.dout(n981),.clk(gclk));
	jor g0909(.dina(n981),.dinb(w_dff_B_XvEe2tqO0_1),.dout(n982),.clk(gclk));
	jand g0910(.dina(n982),.dinb(w_n604_0[2]),.dout(n983),.clk(gclk));
	jand g0911(.dina(w_dff_B_rDa61NF65_0),.dinb(n978),.dout(n984),.clk(gclk));
	jand g0912(.dina(w_dff_B_aNkwzhXz0_0),.dinb(n946),.dout(n985),.clk(gclk));
	jnot g0913(.din(n985),.dout(n986),.clk(gclk));
	jand g0914(.dina(w_dff_B_fRdCpgyv1_0),.dinb(n944),.dout(n987),.clk(gclk));
	jand g0915(.dina(n987),.dinb(n943),.dout(n988),.clk(gclk));
	jnot g0916(.din(w_n988_0[2]),.dout(w_dff_A_zmyyTuog8_1),.clk(gclk));
	jnot g0917(.din(w_n758_0[2]),.dout(n990),.clk(gclk));
	jand g0918(.dina(w_n696_0[1]),.dinb(w_n588_0[1]),.dout(n991),.clk(gclk));
	jand g0919(.dina(w_n991_0[1]),.dinb(w_n764_0[2]),.dout(n992),.clk(gclk));
	jxor g0920(.dina(w_n992_0[1]),.dinb(w_n990_0[1]),.dout(n993),.clk(gclk));
	jxor g0921(.dina(n993),.dinb(w_n769_0[0]),.dout(n994),.clk(gclk));
	jand g0922(.dina(w_n589_0[1]),.dinb(w_n519_0[1]),.dout(n995),.clk(gclk));
	jor g0923(.dina(n995),.dinb(w_n548_0[0]),.dout(n996),.clk(gclk));
	jand g0924(.dina(w_n554_1[0]),.dinb(w_n404_0[0]),.dout(n997),.clk(gclk));
	jor g0925(.dina(w_dff_B_9Lpsubch3_0),.dinb(w_n759_0[0]),.dout(n998),.clk(gclk));
	jnot g0926(.din(w_n764_0[1]),.dout(n999),.clk(gclk));
	jxor g0927(.dina(w_n991_0[0]),.dinb(w_n999_0[1]),.dout(n1000),.clk(gclk));
	jxor g0928(.dina(n1000),.dinb(n998),.dout(n1001),.clk(gclk));
	jor g0929(.dina(w_n1001_0[2]),.dinb(w_n996_0[2]),.dout(n1002),.clk(gclk));
	jor g0930(.dina(w_n1002_0[2]),.dinb(w_n994_0[2]),.dout(n1003),.clk(gclk));
	jnot g0931(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jand g0932(.dina(w_n1002_0[1]),.dinb(w_n994_0[1]),.dout(n1005),.clk(gclk));
	jor g0933(.dina(n1005),.dinb(w_n592_1[0]),.dout(n1006),.clk(gclk));
	jor g0934(.dina(n1006),.dinb(n1004),.dout(n1007),.clk(gclk));
	jor g0935(.dina(w_n994_0[0]),.dinb(w_n603_1[1]),.dout(n1008),.clk(gclk));
	jand g0936(.dina(w_n990_0[0]),.dinb(w_n425_1[0]),.dout(n1009),.clk(gclk));
	jnot g0937(.din(n1009),.dout(n1010),.clk(gclk));
	jand g0938(.dina(w_n631_4[0]),.dinb(w_G125_0[1]),.dout(n1011),.clk(gclk));
	jand g0939(.dina(w_n623_2[1]),.dinb(w_G159_1[2]),.dout(n1012),.clk(gclk));
	jand g0940(.dina(w_n642_4[0]),.dinb(w_G137_1[0]),.dout(n1013),.clk(gclk));
	jor g0941(.dina(w_dff_B_UOaAKzrk5_0),.dinb(n1012),.dout(n1014),.clk(gclk));
	jor g0942(.dina(n1014),.dinb(w_dff_B_fUpwtMpE7_1),.dout(n1015),.clk(gclk));
	jand g0943(.dina(w_n617_3[0]),.dinb(w_G150_1[2]),.dout(n1016),.clk(gclk));
	jor g0944(.dina(n1016),.dinb(w_G33_4[1]),.dout(n1017),.clk(gclk));
	jand g0945(.dina(w_n636_4[0]),.dinb(w_G143_1[1]),.dout(n1018),.clk(gclk));
	jand g0946(.dina(w_n627_4[0]),.dinb(w_G132_1[0]),.dout(n1019),.clk(gclk));
	jor g0947(.dina(n1019),.dinb(n1018),.dout(n1020),.clk(gclk));
	jand g0948(.dina(w_n640_4[0]),.dinb(w_G128_0[2]),.dout(n1021),.clk(gclk));
	jand g0949(.dina(w_n634_2[0]),.dinb(w_G50_2[0]),.dout(n1022),.clk(gclk));
	jor g0950(.dina(n1022),.dinb(w_dff_B_0MkERJX76_1),.dout(n1023),.clk(gclk));
	jor g0951(.dina(n1023),.dinb(w_dff_B_wFxVZoM59_1),.dout(n1024),.clk(gclk));
	jor g0952(.dina(n1024),.dinb(w_dff_B_yGPfwFgA3_1),.dout(n1025),.clk(gclk));
	jor g0953(.dina(n1025),.dinb(w_dff_B_RFjhdhla7_1),.dout(n1026),.clk(gclk));
	jand g0954(.dina(w_n631_3[2]),.dinb(w_G294_1[1]),.dout(n1027),.clk(gclk));
	jand g0955(.dina(w_n642_3[2]),.dinb(w_G107_2[1]),.dout(n1028),.clk(gclk));
	jor g0956(.dina(w_dff_B_M3Zz5C7m8_0),.dinb(w_n962_0[0]),.dout(n1029),.clk(gclk));
	jor g0957(.dina(n1029),.dinb(w_dff_B_86zZpgHb2_1),.dout(n1030),.clk(gclk));
	jand g0958(.dina(w_n640_3[2]),.dinb(w_G283_1[2]),.dout(n1031),.clk(gclk));
	jor g0959(.dina(n1031),.dinb(w_n148_3[2]),.dout(n1032),.clk(gclk));
	jand g0960(.dina(w_n636_3[2]),.dinb(w_G97_2[1]),.dout(n1033),.clk(gclk));
	jand g0961(.dina(w_n627_3[2]),.dinb(w_G116_2[0]),.dout(n1034),.clk(gclk));
	jor g0962(.dina(n1034),.dinb(n1033),.dout(n1035),.clk(gclk));
	jor g0963(.dina(w_n717_0[0]),.dinb(w_n654_0[0]),.dout(n1036),.clk(gclk));
	jor g0964(.dina(n1036),.dinb(w_dff_B_RP8VEQR27_1),.dout(n1037),.clk(gclk));
	jor g0965(.dina(n1037),.dinb(w_dff_B_TQP1YUm59_1),.dout(n1038),.clk(gclk));
	jor g0966(.dina(n1038),.dinb(w_dff_B_Af0sdr0X2_1),.dout(n1039),.clk(gclk));
	jand g0967(.dina(n1039),.dinb(n1026),.dout(n1040),.clk(gclk));
	jor g0968(.dina(n1040),.dinb(w_n612_2[0]),.dout(n1041),.clk(gclk));
	jand g0969(.dina(w_n743_1[0]),.dinb(w_n74_0[1]),.dout(n1042),.clk(gclk));
	jor g0970(.dina(w_dff_B_LwLodLqI6_0),.dinb(w_n605_1[0]),.dout(n1043),.clk(gclk));
	jnot g0971(.din(n1043),.dout(n1044),.clk(gclk));
	jand g0972(.dina(w_dff_B_v7qJ2qFU7_0),.dinb(n1041),.dout(n1045),.clk(gclk));
	jand g0973(.dina(w_dff_B_VwXBFnol2_0),.dinb(n1010),.dout(n1046),.clk(gclk));
	jnot g0974(.din(n1046),.dout(n1047),.clk(gclk));
	jand g0975(.dina(w_dff_B_Nrqi0ynE4_0),.dinb(n1008),.dout(n1048),.clk(gclk));
	jand g0976(.dina(w_dff_B_SWbG8yOW4_0),.dinb(n1007),.dout(n1049),.clk(gclk));
	jnot g0977(.din(w_n1049_0[2]),.dout(w_dff_A_ywGiTRig5_1),.clk(gclk));
	jand g0978(.dina(w_n992_0[0]),.dinb(w_n758_0[1]),.dout(n1051),.clk(gclk));
	jand g0979(.dina(w_n552_0[1]),.dinb(w_n479_0[0]),.dout(n1052),.clk(gclk));
	jnot g0980(.din(w_n1052_0[1]),.dout(n1053),.clk(gclk));
	jand g0981(.dina(n1053),.dinb(w_n484_0[0]),.dout(n1054),.clk(gclk));
	jand g0982(.dina(w_n1052_0[0]),.dinb(w_n541_0[0]),.dout(n1055),.clk(gclk));
	jor g0983(.dina(n1055),.dinb(n1054),.dout(n1056),.clk(gclk));
	jnot g0984(.din(n1056),.dout(n1057),.clk(gclk));
	jxor g0985(.dina(w_n1057_0[1]),.dinb(w_n771_0[0]),.dout(n1058),.clk(gclk));
	jxor g0986(.dina(n1058),.dinb(w_dff_B_d1NIOL8X8_1),.dout(n1059),.clk(gclk));
	jor g0987(.dina(w_n1059_0[1]),.dinb(w_n603_1[0]),.dout(n1060),.clk(gclk));
	jnot g0988(.din(w_n996_0[1]),.dout(n1061),.clk(gclk));
	jand g0989(.dina(w_n1003_0[0]),.dinb(w_dff_B_qMUJgFx84_1),.dout(n1062),.clk(gclk));
	jor g0990(.dina(n1062),.dinb(w_n592_0[2]),.dout(n1063),.clk(gclk));
	jor g0991(.dina(n1063),.dinb(w_n1059_0[0]),.dout(n1064),.clk(gclk));
	jand g0992(.dina(w_n1057_0[0]),.dinb(w_n425_0[2]),.dout(n1065),.clk(gclk));
	jnot g0993(.din(w_n612_1[2]),.dout(n1066),.clk(gclk));
	jand g0994(.dina(w_n642_3[1]),.dinb(w_G132_0[2]),.dout(n1067),.clk(gclk));
	jand g0995(.dina(w_n627_3[1]),.dinb(w_G128_0[1]),.dout(n1068),.clk(gclk));
	jand g0996(.dina(w_n636_3[1]),.dinb(w_G137_0[2]),.dout(n1069),.clk(gclk));
	jor g0997(.dina(n1069),.dinb(n1068),.dout(n1070),.clk(gclk));
	jor g0998(.dina(n1070),.dinb(w_dff_B_9uif3c2I5_1),.dout(n1071),.clk(gclk));
	jnot g0999(.din(n1071),.dout(n1072),.clk(gclk));
	jand g1000(.dina(w_n623_2[0]),.dinb(w_G150_1[1]),.dout(n1073),.clk(gclk));
	jnot g1001(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1002(.dina(w_n149_1[0]),.dinb(w_n148_3[1]),.dout(n1075),.clk(gclk));
	jand g1003(.dina(w_dff_B_dtJPXaif5_0),.dinb(n1074),.dout(n1076),.clk(gclk));
	jand g1004(.dina(w_n640_3[1]),.dinb(w_G125_0[0]),.dout(n1077),.clk(gclk));
	jand g1005(.dina(w_n617_2[2]),.dinb(w_G143_1[0]),.dout(n1078),.clk(gclk));
	jor g1006(.dina(n1078),.dinb(w_dff_B_EG6ARHJv1_1),.dout(n1079),.clk(gclk));
	jand g1007(.dina(w_n631_3[1]),.dinb(w_dff_B_vnVczlSn4_1),.dout(n1080),.clk(gclk));
	jand g1008(.dina(w_n634_1[2]),.dinb(w_G159_1[1]),.dout(n1081),.clk(gclk));
	jor g1009(.dina(n1081),.dinb(n1080),.dout(n1082),.clk(gclk));
	jor g1010(.dina(n1082),.dinb(n1079),.dout(n1083),.clk(gclk));
	jnot g1011(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1012(.dina(n1084),.dinb(w_dff_B_ggGMsJUX2_1),.dout(n1085),.clk(gclk));
	jand g1013(.dina(n1085),.dinb(w_dff_B_SFjiaPKT8_1),.dout(n1086),.clk(gclk));
	jand g1014(.dina(w_n627_3[0]),.dinb(w_G107_2[0]),.dout(n1087),.clk(gclk));
	jand g1015(.dina(w_n634_1[1]),.dinb(w_G58_1[2]),.dout(n1088),.clk(gclk));
	jand g1016(.dina(w_n636_3[0]),.dinb(w_G87_1[0]),.dout(n1089),.clk(gclk));
	jor g1017(.dina(w_dff_B_HVAqcWer1_0),.dinb(w_n1088_0[1]),.dout(n1090),.clk(gclk));
	jor g1018(.dina(n1090),.dinb(w_dff_B_YsUganJu0_1),.dout(n1091),.clk(gclk));
	jnot g1019(.din(n1091),.dout(n1092),.clk(gclk));
	jand g1020(.dina(w_n642_3[0]),.dinb(w_G97_2[0]),.dout(n1093),.clk(gclk));
	jnot g1021(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1022(.dina(w_n149_0[2]),.dinb(w_G33_4[0]),.dout(n1095),.clk(gclk));
	jand g1023(.dina(w_dff_B_5S8Al6CO4_0),.dinb(n1094),.dout(n1096),.clk(gclk));
	jand g1024(.dina(w_n631_3[0]),.dinb(w_G283_1[1]),.dout(n1097),.clk(gclk));
	jor g1025(.dina(n1097),.dinb(w_n823_0[0]),.dout(n1098),.clk(gclk));
	jand g1026(.dina(w_n640_3[0]),.dinb(w_G116_1[2]),.dout(n1099),.clk(gclk));
	jor g1027(.dina(w_dff_B_hNlRGnM00_0),.dinb(w_n909_0[0]),.dout(n1100),.clk(gclk));
	jor g1028(.dina(n1100),.dinb(n1098),.dout(n1101),.clk(gclk));
	jnot g1029(.din(n1101),.dout(n1102),.clk(gclk));
	jand g1030(.dina(n1102),.dinb(w_dff_B_NepKsP0S7_1),.dout(n1103),.clk(gclk));
	jand g1031(.dina(n1103),.dinb(w_dff_B_l64JFMp40_1),.dout(n1104),.clk(gclk));
	jand g1032(.dina(w_n73_1[0]),.dinb(w_G41_0[1]),.dout(n1105),.clk(gclk));
	jor g1033(.dina(w_dff_B_7iHYmG9Z8_0),.dinb(n1104),.dout(n1106),.clk(gclk));
	jor g1034(.dina(n1106),.dinb(w_dff_B_VB52pyBY9_1),.dout(n1107),.clk(gclk));
	jand g1035(.dina(n1107),.dinb(w_dff_B_PeH7jio82_1),.dout(n1108),.clk(gclk));
	jand g1036(.dina(w_n743_0[2]),.dinb(w_n73_0[2]),.dout(n1109),.clk(gclk));
	jor g1037(.dina(w_dff_B_ROu9VDUx5_0),.dinb(w_n605_0[2]),.dout(n1110),.clk(gclk));
	jor g1038(.dina(w_dff_B_fS9LehUH7_0),.dinb(n1108),.dout(n1111),.clk(gclk));
	jor g1039(.dina(w_dff_B_92gJze930_0),.dinb(n1065),.dout(n1112),.clk(gclk));
	jand g1040(.dina(w_dff_B_H8cVUlWX9_0),.dinb(n1064),.dout(n1113),.clk(gclk));
	jand g1041(.dina(n1113),.dinb(w_dff_B_DVFnj4U50_1),.dout(n1114),.clk(gclk));
	jnot g1042(.din(w_n1114_0[2]),.dout(w_dff_A_ULxsSlua0_1),.clk(gclk));
	jand g1043(.dina(w_n1001_0[1]),.dinb(w_n996_0[0]),.dout(n1116),.clk(gclk));
	jnot g1044(.din(n1116),.dout(n1117),.clk(gclk));
	jand g1045(.dina(w_n1002_0[0]),.dinb(w_n591_0[1]),.dout(n1118),.clk(gclk));
	jand g1046(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jnot g1047(.din(n1119),.dout(n1120),.clk(gclk));
	jor g1048(.dina(w_n1001_0[0]),.dinb(w_n603_0[2]),.dout(n1121),.clk(gclk));
	jand g1049(.dina(w_n999_0[0]),.dinb(w_n425_0[1]),.dout(n1122),.clk(gclk));
	jnot g1050(.din(n1122),.dout(n1123),.clk(gclk));
	jand g1051(.dina(w_n623_1[2]),.dinb(w_G50_1[2]),.dout(n1124),.clk(gclk));
	jand g1052(.dina(w_n617_2[1]),.dinb(w_G159_1[0]),.dout(n1125),.clk(gclk));
	jand g1053(.dina(w_n642_2[2]),.dinb(w_G143_0[2]),.dout(n1126),.clk(gclk));
	jor g1054(.dina(w_dff_B_fMJ8Nppx0_0),.dinb(n1125),.dout(n1127),.clk(gclk));
	jor g1055(.dina(n1127),.dinb(w_dff_B_WXlW6o9w3_1),.dout(n1128),.clk(gclk));
	jand g1056(.dina(w_n631_2[2]),.dinb(w_G128_0[0]),.dout(n1129),.clk(gclk));
	jor g1057(.dina(n1129),.dinb(w_G33_3[2]),.dout(n1130),.clk(gclk));
	jand g1058(.dina(w_n636_2[2]),.dinb(w_G150_1[0]),.dout(n1131),.clk(gclk));
	jand g1059(.dina(w_n627_2[2]),.dinb(w_G137_0[1]),.dout(n1132),.clk(gclk));
	jor g1060(.dina(n1132),.dinb(n1131),.dout(n1133),.clk(gclk));
	jand g1061(.dina(w_n640_2[2]),.dinb(w_G132_0[1]),.dout(n1134),.clk(gclk));
	jor g1062(.dina(w_dff_B_0c9EyVMM9_0),.dinb(w_n1088_0[0]),.dout(n1135),.clk(gclk));
	jor g1063(.dina(n1135),.dinb(w_dff_B_Qnxe6shB7_1),.dout(n1136),.clk(gclk));
	jor g1064(.dina(n1136),.dinb(w_dff_B_2SeKlOP91_1),.dout(n1137),.clk(gclk));
	jor g1065(.dina(n1137),.dinb(w_dff_B_tY6y2k0Q3_1),.dout(n1138),.clk(gclk));
	jand g1066(.dina(w_n617_2[0]),.dinb(w_G97_1[2]),.dout(n1139),.clk(gclk));
	jand g1067(.dina(w_n640_2[1]),.dinb(w_G294_1[0]),.dout(n1140),.clk(gclk));
	jand g1068(.dina(w_n642_2[1]),.dinb(w_G116_1[1]),.dout(n1141),.clk(gclk));
	jor g1069(.dina(n1141),.dinb(n1140),.dout(n1142),.clk(gclk));
	jor g1070(.dina(n1142),.dinb(n1139),.dout(n1143),.clk(gclk));
	jand g1071(.dina(w_n631_2[1]),.dinb(w_G303_0[2]),.dout(n1144),.clk(gclk));
	jor g1072(.dina(n1144),.dinb(w_n148_3[0]),.dout(n1145),.clk(gclk));
	jand g1073(.dina(w_n636_2[1]),.dinb(w_G107_1[2]),.dout(n1146),.clk(gclk));
	jand g1074(.dina(w_n627_2[1]),.dinb(w_G283_1[0]),.dout(n1147),.clk(gclk));
	jor g1075(.dina(n1147),.dinb(n1146),.dout(n1148),.clk(gclk));
	jor g1076(.dina(w_n899_0[0]),.dinb(w_n825_0[0]),.dout(n1149),.clk(gclk));
	jor g1077(.dina(n1149),.dinb(w_dff_B_txrUvoTl4_1),.dout(n1150),.clk(gclk));
	jor g1078(.dina(n1150),.dinb(w_dff_B_Vg4DbODl7_1),.dout(n1151),.clk(gclk));
	jor g1079(.dina(n1151),.dinb(w_dff_B_gNhm7Jq30_1),.dout(n1152),.clk(gclk));
	jand g1080(.dina(n1152),.dinb(n1138),.dout(n1153),.clk(gclk));
	jor g1081(.dina(n1153),.dinb(w_n612_1[1]),.dout(n1154),.clk(gclk));
	jand g1082(.dina(w_n743_0[1]),.dinb(w_n75_0[1]),.dout(n1155),.clk(gclk));
	jor g1083(.dina(w_dff_B_QWgYZoqw4_0),.dinb(w_n605_0[1]),.dout(n1156),.clk(gclk));
	jnot g1084(.din(n1156),.dout(n1157),.clk(gclk));
	jand g1085(.dina(w_dff_B_rHfN2sbM6_0),.dinb(n1154),.dout(n1158),.clk(gclk));
	jand g1086(.dina(w_dff_B_kl4sFjwJ4_0),.dinb(n1123),.dout(n1159),.clk(gclk));
	jnot g1087(.din(n1159),.dout(n1160),.clk(gclk));
	jand g1088(.dina(n1160),.dinb(n1121),.dout(n1161),.clk(gclk));
	jand g1089(.dina(w_dff_B_CJNgHhWI8_0),.dinb(n1120),.dout(n1162),.clk(gclk));
	jnot g1090(.din(w_n1162_0[2]),.dout(w_dff_A_BEk3hAnd8_1),.clk(gclk));
	jand g1091(.dina(w_n1114_0[1]),.dinb(w_n1049_0[1]),.dout(n1164),.clk(gclk));
	jnot g1092(.din(w_G387_0[1]),.dout(n1165),.clk(gclk));
	jnot g1093(.din(w_G396_0[1]),.dout(n1166),.clk(gclk));
	jand g1094(.dina(w_n937_0[1]),.dinb(w_dff_B_F6HiktET4_1),.dout(n1167),.clk(gclk));
	jand g1095(.dina(n1167),.dinb(w_n750_0[0]),.dout(n1168),.clk(gclk));
	jand g1096(.dina(n1168),.dinb(w_n988_0[1]),.dout(n1169),.clk(gclk));
	jand g1097(.dina(n1169),.dinb(w_n1162_0[1]),.dout(n1170),.clk(gclk));
	jand g1098(.dina(n1170),.dinb(n1165),.dout(n1171),.clk(gclk));
	jand g1099(.dina(n1171),.dinb(w_n1164_0[1]),.dout(n1172),.clk(gclk));
	jnot g1100(.din(w_n1172_0[1]),.dout(w_dff_A_jCISqWYT9_1),.clk(gclk));
	jnot g1101(.din(w_G213_0[1]),.dout(n1174),.clk(gclk));
	jnot g1102(.din(w_G343_0[0]),.dout(n1175),.clk(gclk));
	jand g1103(.dina(w_n1164_0[0]),.dinb(w_n1175_0[1]),.dout(n1176),.clk(gclk));
	jor g1104(.dina(n1176),.dinb(w_dff_B_Dkas4rHc5_1),.dout(n1177),.clk(gclk));
	jor g1105(.dina(n1177),.dinb(w_n1172_0[0]),.dout(G409),.clk(gclk));
	jxor g1106(.dina(w_n1162_0[0]),.dinb(w_G384_0),.dout(n1179),.clk(gclk));
	jxor g1107(.dina(w_n937_0[0]),.dinb(w_G396_0[0]),.dout(n1180),.clk(gclk));
	jxor g1108(.dina(w_n988_0[0]),.dinb(w_G387_0[0]),.dout(n1181),.clk(gclk));
	jxor g1109(.dina(n1181),.dinb(w_dff_B_nePEl5Xx0_1),.dout(n1182),.clk(gclk));
	jxor g1110(.dina(n1182),.dinb(w_dff_B_mMffx1gt7_1),.dout(n1183),.clk(gclk));
	jand g1111(.dina(w_n1175_0[0]),.dinb(w_G213_0[0]),.dout(n1184),.clk(gclk));
	jnot g1112(.din(w_n1184_0[1]),.dout(n1185),.clk(gclk));
	jor g1113(.dina(n1185),.dinb(w_dff_B_Tn5Dfvsh7_1),.dout(n1186),.clk(gclk));
	jxor g1114(.dina(w_n1114_0[0]),.dinb(w_n1049_0[0]),.dout(n1187),.clk(gclk));
	jor g1115(.dina(w_n1187_0[1]),.dinb(w_n1184_0[0]),.dout(n1188),.clk(gclk));
	jand g1116(.dina(n1188),.dinb(w_dff_B_nNzt09gq4_1),.dout(n1189),.clk(gclk));
	jxor g1117(.dina(n1189),.dinb(w_n1183_0[1]),.dout(G405),.clk(gclk));
	jxor g1118(.dina(w_n1187_0[0]),.dinb(w_n1183_0[0]),.dout(w_dff_A_ysFzlHig4_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_dff_A_iAdXw7Hj8_0),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_dff_A_ic6VYL2s1_0),.doutb(w_dff_A_nxOb1jX52_1),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G1_2(.douta(w_dff_A_3nvoBC4Z2_0),.doutb(w_G1_2[1]),.doutc(w_dff_A_O3PSfUPA3_2),.din(w_G1_0[1]));
	jspl jspl_w_G1_3(.douta(w_G1_3[0]),.doutb(w_G1_3[1]),.din(w_G1_0[2]));
	jspl3 jspl3_w_G13_0(.douta(w_G13_0[0]),.doutb(w_dff_A_pLbnh99t5_1),.doutc(w_dff_A_0eRuYOQO3_2),.din(G13));
	jspl jspl_w_G13_1(.douta(w_G13_1[0]),.doutb(w_G13_1[1]),.din(w_G13_0[0]));
	jspl3 jspl3_w_G20_0(.douta(w_dff_A_nOj7S6af6_0),.doutb(w_G20_0[1]),.doutc(w_G20_0[2]),.din(G20));
	jspl3 jspl3_w_G20_1(.douta(w_G20_1[0]),.doutb(w_G20_1[1]),.doutc(w_dff_A_Ekx2lsgO5_2),.din(w_G20_0[0]));
	jspl3 jspl3_w_G20_2(.douta(w_G20_2[0]),.doutb(w_dff_A_Madlfysn3_1),.doutc(w_G20_2[2]),.din(w_G20_0[1]));
	jspl3 jspl3_w_G20_3(.douta(w_G20_3[0]),.doutb(w_dff_A_Jgno6nkh7_1),.doutc(w_dff_A_7sF9HlrM6_2),.din(w_G20_0[2]));
	jspl3 jspl3_w_G20_4(.douta(w_dff_A_KXGCIGqG1_0),.doutb(w_dff_A_13G9R5bH5_1),.doutc(w_G20_4[2]),.din(w_G20_1[0]));
	jspl3 jspl3_w_G20_5(.douta(w_dff_A_tnr0FCP54_0),.doutb(w_dff_A_J9rY81dQ7_1),.doutc(w_G20_5[2]),.din(w_G20_1[1]));
	jspl3 jspl3_w_G20_6(.douta(w_dff_A_1hQTGFhM4_0),.doutb(w_G20_6[1]),.doutc(w_G20_6[2]),.din(w_G20_1[2]));
	jspl jspl_w_G20_7(.douta(w_G20_7[0]),.doutb(w_G20_7[1]),.din(w_G20_2[0]));
	jspl3 jspl3_w_G33_0(.douta(w_dff_A_KPWEOBb32_0),.doutb(w_G33_0[1]),.doutc(w_G33_0[2]),.din(G33));
	jspl3 jspl3_w_G33_1(.douta(w_G33_1[0]),.doutb(w_dff_A_JkA8zOvk6_1),.doutc(w_G33_1[2]),.din(w_G33_0[0]));
	jspl3 jspl3_w_G33_2(.douta(w_G33_2[0]),.doutb(w_G33_2[1]),.doutc(w_G33_2[2]),.din(w_G33_0[1]));
	jspl3 jspl3_w_G33_3(.douta(w_G33_3[0]),.doutb(w_G33_3[1]),.doutc(w_dff_A_8qgATIe62_2),.din(w_G33_0[2]));
	jspl3 jspl3_w_G33_4(.douta(w_G33_4[0]),.doutb(w_dff_A_sVwYQHnY4_1),.doutc(w_dff_A_yjpnAqiE4_2),.din(w_G33_1[0]));
	jspl3 jspl3_w_G33_5(.douta(w_dff_A_nByLp5Ye4_0),.doutb(w_G33_5[1]),.doutc(w_dff_A_8G95VIjC4_2),.din(w_G33_1[1]));
	jspl3 jspl3_w_G33_6(.douta(w_dff_A_RACd9pjg9_0),.doutb(w_dff_A_oDlAgc7P2_1),.doutc(w_G33_6[2]),.din(w_G33_1[2]));
	jspl3 jspl3_w_G33_7(.douta(w_G33_7[0]),.doutb(w_G33_7[1]),.doutc(w_G33_7[2]),.din(w_G33_2[0]));
	jspl3 jspl3_w_G33_8(.douta(w_dff_A_PfzZNePP1_0),.doutb(w_G33_8[1]),.doutc(w_G33_8[2]),.din(w_G33_2[1]));
	jspl3 jspl3_w_G33_9(.douta(w_G33_9[0]),.doutb(w_G33_9[1]),.doutc(w_dff_A_uzO5xhyl4_2),.din(w_G33_2[2]));
	jspl3 jspl3_w_G33_10(.douta(w_dff_A_fxc072rn5_0),.doutb(w_dff_A_uZz1fQBT7_1),.doutc(w_G33_10[2]),.din(w_G33_3[0]));
	jspl3 jspl3_w_G33_11(.douta(w_G33_11[0]),.doutb(w_G33_11[1]),.doutc(w_G33_11[2]),.din(w_G33_3[1]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_dff_A_eheZoAGo8_1),.doutc(w_dff_A_AH0KJFDU0_2),.din(G41));
	jspl jspl_w_G41_1(.douta(w_G41_1[0]),.doutb(w_G41_1[1]),.din(w_G41_0[0]));
	jspl3 jspl3_w_G45_0(.douta(w_G45_0[0]),.doutb(w_dff_A_yQTxWFRA1_1),.doutc(w_dff_A_UYUfUEAd4_2),.din(G45));
	jspl3 jspl3_w_G45_1(.douta(w_dff_A_CO9EWdaC6_0),.doutb(w_dff_A_GFDKQ38K5_1),.doutc(w_G45_1[2]),.din(w_G45_0[0]));
	jspl3 jspl3_w_G50_0(.douta(w_G50_0[0]),.doutb(w_dff_A_ZukS50L22_1),.doutc(w_G50_0[2]),.din(G50));
	jspl3 jspl3_w_G50_1(.douta(w_dff_A_n01tZAbE4_0),.doutb(w_G50_1[1]),.doutc(w_dff_A_sQxHYeYf6_2),.din(w_G50_0[0]));
	jspl3 jspl3_w_G50_2(.douta(w_dff_A_Atnr6eaZ2_0),.doutb(w_G50_2[1]),.doutc(w_G50_2[2]),.din(w_G50_0[1]));
	jspl3 jspl3_w_G50_3(.douta(w_dff_A_o3YWIpC56_0),.doutb(w_G50_3[1]),.doutc(w_dff_A_r1HWMIYL7_2),.din(w_G50_0[2]));
	jspl3 jspl3_w_G50_4(.douta(w_dff_A_UyoE6NVP6_0),.doutb(w_dff_A_AEGITx9G9_1),.doutc(w_G50_4[2]),.din(w_G50_1[0]));
	jspl3 jspl3_w_G50_5(.douta(w_G50_5[0]),.doutb(w_dff_A_dc4sKXuE5_1),.doutc(w_G50_5[2]),.din(w_G50_1[1]));
	jspl3 jspl3_w_G58_0(.douta(w_G58_0[0]),.doutb(w_dff_A_i85muIC40_1),.doutc(w_dff_A_cxfkScNB3_2),.din(G58));
	jspl3 jspl3_w_G58_1(.douta(w_dff_A_6m0bHzbb6_0),.doutb(w_G58_1[1]),.doutc(w_dff_A_pR8uKgO07_2),.din(w_G58_0[0]));
	jspl3 jspl3_w_G58_2(.douta(w_dff_A_n8CIkRW42_0),.doutb(w_G58_2[1]),.doutc(w_dff_A_JtTPq6K41_2),.din(w_G58_0[1]));
	jspl3 jspl3_w_G58_3(.douta(w_dff_A_r5Tudtj48_0),.doutb(w_dff_A_Rn3uLTyX2_1),.doutc(w_G58_3[2]),.din(w_G58_0[2]));
	jspl3 jspl3_w_G58_4(.douta(w_dff_A_QWWqCtkg0_0),.doutb(w_dff_A_Mjh3b7UO7_1),.doutc(w_G58_4[2]),.din(w_G58_1[0]));
	jspl jspl_w_G58_5(.douta(w_G58_5[0]),.doutb(w_G58_5[1]),.din(w_G58_1[1]));
	jspl3 jspl3_w_G68_0(.douta(w_G68_0[0]),.doutb(w_G68_0[1]),.doutc(w_dff_A_si08ltWt9_2),.din(G68));
	jspl3 jspl3_w_G68_1(.douta(w_dff_A_0corOKVj7_0),.doutb(w_G68_1[1]),.doutc(w_dff_A_aD3bYPsb3_2),.din(w_G68_0[0]));
	jspl3 jspl3_w_G68_2(.douta(w_G68_2[0]),.doutb(w_dff_A_uiOC0J294_1),.doutc(w_dff_A_6KVDIPDC3_2),.din(w_G68_0[1]));
	jspl3 jspl3_w_G68_3(.douta(w_G68_3[0]),.doutb(w_dff_A_2pHJVp7l8_1),.doutc(w_dff_A_9JmFPU7u0_2),.din(w_G68_0[2]));
	jspl3 jspl3_w_G68_4(.douta(w_dff_A_8wMjJHIG7_0),.doutb(w_dff_A_PJNWczpa1_1),.doutc(w_G68_4[2]),.din(w_G68_1[0]));
	jspl jspl_w_G68_5(.douta(w_G68_5[0]),.doutb(w_G68_5[1]),.din(w_G68_1[1]));
	jspl3 jspl3_w_G77_0(.douta(w_G77_0[0]),.doutb(w_G77_0[1]),.doutc(w_G77_0[2]),.din(G77));
	jspl3 jspl3_w_G77_1(.douta(w_dff_A_ByuNwsEG1_0),.doutb(w_G77_1[1]),.doutc(w_dff_A_WUSlaZ817_2),.din(w_G77_0[0]));
	jspl3 jspl3_w_G77_2(.douta(w_G77_2[0]),.doutb(w_dff_A_qIt7Kmcb5_1),.doutc(w_dff_A_4vBQYFhr8_2),.din(w_G77_0[1]));
	jspl3 jspl3_w_G77_3(.douta(w_G77_3[0]),.doutb(w_dff_A_O31Yevz94_1),.doutc(w_G77_3[2]),.din(w_G77_0[2]));
	jspl3 jspl3_w_G77_4(.douta(w_dff_A_dfSf8Hys6_0),.doutb(w_G77_4[1]),.doutc(w_G77_4[2]),.din(w_G77_1[0]));
	jspl jspl_w_G77_5(.douta(w_G77_5[0]),.doutb(w_G77_5[1]),.din(w_G77_1[1]));
	jspl3 jspl3_w_G87_0(.douta(w_dff_A_yTyBwOZq2_0),.doutb(w_G87_0[1]),.doutc(w_G87_0[2]),.din(G87));
	jspl3 jspl3_w_G87_1(.douta(w_G87_1[0]),.doutb(w_dff_A_mKI2h6GU8_1),.doutc(w_dff_A_d7F1LZsA6_2),.din(w_G87_0[0]));
	jspl3 jspl3_w_G87_2(.douta(w_dff_A_aVsadp7V2_0),.doutb(w_dff_A_rGYIVoJs5_1),.doutc(w_G87_2[2]),.din(w_G87_0[1]));
	jspl3 jspl3_w_G87_3(.douta(w_dff_A_001aC8LN9_0),.doutb(w_G87_3[1]),.doutc(w_dff_A_c7vPv7cN1_2),.din(w_G87_0[2]));
	jspl3 jspl3_w_G97_0(.douta(w_G97_0[0]),.doutb(w_dff_A_C9em7tj81_1),.doutc(w_dff_A_8qEqV5IG1_2),.din(G97));
	jspl3 jspl3_w_G97_1(.douta(w_G97_1[0]),.doutb(w_G97_1[1]),.doutc(w_dff_A_9oPM0F8E6_2),.din(w_G97_0[0]));
	jspl3 jspl3_w_G97_2(.douta(w_G97_2[0]),.doutb(w_G97_2[1]),.doutc(w_dff_A_jQ6iCYFb7_2),.din(w_G97_0[1]));
	jspl3 jspl3_w_G97_3(.douta(w_dff_A_zgFStbQ32_0),.doutb(w_dff_A_ccuwuU1G7_1),.doutc(w_G97_3[2]),.din(w_G97_0[2]));
	jspl3 jspl3_w_G97_4(.douta(w_dff_A_uB9kAt2B0_0),.doutb(w_G97_4[1]),.doutc(w_G97_4[2]),.din(w_G97_1[0]));
	jspl jspl_w_G97_5(.douta(w_dff_A_GViDkCJD7_0),.doutb(w_G97_5[1]),.din(w_G97_1[1]));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_dff_A_FTkE7pQJ2_1),.doutc(w_dff_A_pw1EcozM1_2),.din(G107));
	jspl3 jspl3_w_G107_1(.douta(w_G107_1[0]),.doutb(w_G107_1[1]),.doutc(w_dff_A_O1jHvSWP8_2),.din(w_G107_0[0]));
	jspl3 jspl3_w_G107_2(.douta(w_G107_2[0]),.doutb(w_G107_2[1]),.doutc(w_dff_A_bwpleDz36_2),.din(w_G107_0[1]));
	jspl3 jspl3_w_G107_3(.douta(w_dff_A_p2P0Q2Iy0_0),.doutb(w_dff_A_HoFi2L3R1_1),.doutc(w_G107_3[2]),.din(w_G107_0[2]));
	jspl3 jspl3_w_G107_4(.douta(w_dff_A_oJvYPEnJ3_0),.doutb(w_G107_4[1]),.doutc(w_G107_4[2]),.din(w_G107_1[0]));
	jspl jspl_w_G107_5(.douta(w_G107_5[0]),.doutb(w_G107_5[1]),.din(w_G107_1[1]));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_dff_A_6sEZr79Z9_1),.doutc(w_dff_A_JUzIhdWg1_2),.din(G116));
	jspl3 jspl3_w_G116_1(.douta(w_G116_1[0]),.doutb(w_dff_A_raVhjKGT5_1),.doutc(w_dff_A_pzus6SVP7_2),.din(w_G116_0[0]));
	jspl3 jspl3_w_G116_2(.douta(w_G116_2[0]),.doutb(w_dff_A_nFcxiCu25_1),.doutc(w_dff_A_Ig1MTnX10_2),.din(w_G116_0[1]));
	jspl3 jspl3_w_G116_3(.douta(w_dff_A_gbf3SjqU5_0),.doutb(w_G116_3[1]),.doutc(w_dff_A_RRAZWhbs1_2),.din(w_G116_0[2]));
	jspl3 jspl3_w_G116_4(.douta(w_G116_4[0]),.doutb(w_G116_4[1]),.doutc(w_G116_4[2]),.din(w_G116_1[0]));
	jspl jspl_w_G125_0(.douta(w_G125_0[0]),.doutb(w_dff_A_xsEWv84P2_1),.din(w_dff_B_p5Pr9xfC7_2));
	jspl3 jspl3_w_G128_0(.douta(w_dff_A_SMHDbw023_0),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(w_dff_B_RnScCPeN8_3));
	jspl3 jspl3_w_G132_0(.douta(w_G132_0[0]),.doutb(w_G132_0[1]),.doutc(w_G132_0[2]),.din(w_dff_B_9BanF2Hg6_3));
	jspl jspl_w_G132_1(.douta(w_G132_1[0]),.doutb(w_dff_A_BmJHWTNA3_1),.din(w_G132_0[0]));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(w_dff_B_a8BNTn3r7_3));
	jspl3 jspl3_w_G137_1(.douta(w_G137_1[0]),.doutb(w_dff_A_36uqRPDS7_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(w_dff_B_9juV44ph8_3));
	jspl3 jspl3_w_G143_1(.douta(w_dff_A_PQFRbtVo2_0),.doutb(w_G143_1[1]),.doutc(w_dff_A_qQppqKnn2_2),.din(w_G143_0[0]));
	jspl jspl_w_G143_2(.douta(w_G143_2[0]),.doutb(w_G143_2[1]),.din(w_G143_0[1]));
	jspl3 jspl3_w_G150_0(.douta(w_dff_A_NQlKKxwd2_0),.doutb(w_dff_A_UpKDQn5S3_1),.doutc(w_G150_0[2]),.din(G150));
	jspl3 jspl3_w_G150_1(.douta(w_G150_1[0]),.doutb(w_dff_A_pOidVMvc1_1),.doutc(w_dff_A_oQWicbQb0_2),.din(w_G150_0[0]));
	jspl3 jspl3_w_G150_2(.douta(w_G150_2[0]),.doutb(w_dff_A_UaieZtxF1_1),.doutc(w_G150_2[2]),.din(w_G150_0[1]));
	jspl jspl_w_G150_3(.douta(w_dff_A_wgMpoDW27_0),.doutb(w_G150_3[1]),.din(w_G150_0[2]));
	jspl3 jspl3_w_G159_0(.douta(w_dff_A_VmKgOIih9_0),.doutb(w_dff_A_QZZj3G500_1),.doutc(w_G159_0[2]),.din(w_dff_B_CuiEmr8G7_3));
	jspl3 jspl3_w_G159_1(.douta(w_G159_1[0]),.doutb(w_G159_1[1]),.doutc(w_G159_1[2]),.din(w_G159_0[0]));
	jspl3 jspl3_w_G159_2(.douta(w_G159_2[0]),.doutb(w_G159_2[1]),.doutc(w_G159_2[2]),.din(w_G159_0[1]));
	jspl3 jspl3_w_G159_3(.douta(w_dff_A_ZKbKDlC72_0),.doutb(w_dff_A_Jkc8FQ2x6_1),.doutc(w_G159_3[2]),.din(w_G159_0[2]));
	jspl3 jspl3_w_G169_0(.douta(w_G169_0[0]),.doutb(w_dff_A_73xXv1qJ4_1),.doutc(w_dff_A_QuWBZkPP5_2),.din(G169));
	jspl jspl_w_G169_1(.douta(w_dff_A_G6PyO8im8_0),.doutb(w_G169_1[1]),.din(w_G169_0[0]));
	jspl3 jspl3_w_G179_0(.douta(w_dff_A_Dr0dLoVk1_0),.doutb(w_G179_0[1]),.doutc(w_G179_0[2]),.din(G179));
	jspl3 jspl3_w_G179_1(.douta(w_G179_1[0]),.doutb(w_G179_1[1]),.doutc(w_G179_1[2]),.din(w_G179_0[0]));
	jspl3 jspl3_w_G179_2(.douta(w_dff_A_suGe9WPO6_0),.doutb(w_dff_A_J1ih0qTn6_1),.doutc(w_G179_2[2]),.din(w_G179_0[1]));
	jspl3 jspl3_w_G190_0(.douta(w_dff_A_dVvesc1C1_0),.doutb(w_dff_A_wCBPIBH18_1),.doutc(w_G190_0[2]),.din(G190));
	jspl3 jspl3_w_G190_1(.douta(w_dff_A_tkwBkKGg1_0),.doutb(w_G190_1[1]),.doutc(w_G190_1[2]),.din(w_G190_0[0]));
	jspl3 jspl3_w_G190_2(.douta(w_G190_2[0]),.doutb(w_dff_A_CAXAfBzv5_1),.doutc(w_dff_A_pNsegoOF1_2),.din(w_G190_0[1]));
	jspl3 jspl3_w_G190_3(.douta(w_G190_3[0]),.doutb(w_dff_A_XHC4JfNo2_1),.doutc(w_dff_A_59Z4Cv8n6_2),.din(w_G190_0[2]));
	jspl jspl_w_G190_4(.douta(w_dff_A_qayL26XG4_0),.doutb(w_G190_4[1]),.din(w_G190_1[0]));
	jspl3 jspl3_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.doutc(w_dff_A_mJWlEdhi3_2),.din(G200));
	jspl3 jspl3_w_G200_1(.douta(w_dff_A_bGE5KNDJ7_0),.doutb(w_dff_A_2pTMC7fh9_1),.doutc(w_G200_1[2]),.din(w_G200_0[0]));
	jspl3 jspl3_w_G200_2(.douta(w_G200_2[0]),.doutb(w_dff_A_3g9wCvOT0_1),.doutc(w_dff_A_UHz0db1u2_2),.din(w_G200_0[1]));
	jspl3 jspl3_w_G200_3(.douta(w_G200_3[0]),.doutb(w_G200_3[1]),.doutc(w_G200_3[2]),.din(w_G200_0[2]));
	jspl3 jspl3_w_G200_4(.douta(w_G200_4[0]),.doutb(w_G200_4[1]),.doutc(w_G200_4[2]),.din(w_G200_1[0]));
	jspl3 jspl3_w_G213_0(.douta(w_dff_A_nj5ryxbi9_0),.doutb(w_G213_0[1]),.doutc(w_dff_A_06UoBpWW4_2),.din(G213));
	jspl jspl_w_G223_0(.douta(w_G223_0[0]),.doutb(w_G223_0[1]),.din(w_dff_B_3TZf6n5G1_2));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_dff_A_khPh2FFN8_1),.doutc(w_dff_A_K5vSNaX49_2),.din(G226));
	jspl jspl_w_G226_1(.douta(w_dff_A_z5vuix598_0),.doutb(w_G226_1[1]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G232_0(.douta(w_G232_0[0]),.doutb(w_dff_A_CZISefcV8_1),.doutc(w_dff_A_wZ3zF3iC5_2),.din(G232));
	jspl3 jspl3_w_G232_1(.douta(w_dff_A_2sF6EAVe2_0),.doutb(w_dff_A_lwoF2VS19_1),.doutc(w_G232_1[2]),.din(w_G232_0[0]));
	jspl3 jspl3_w_G238_0(.douta(w_G238_0[0]),.doutb(w_dff_A_pJc5Nymd0_1),.doutc(w_dff_A_9N91VHxD5_2),.din(G238));
	jspl3 jspl3_w_G238_1(.douta(w_dff_A_303rdBsU8_0),.doutb(w_G238_1[1]),.doutc(w_G238_1[2]),.din(w_G238_0[0]));
	jspl3 jspl3_w_G244_0(.douta(w_G244_0[0]),.doutb(w_dff_A_iaPOG52y2_1),.doutc(w_dff_A_bj6XxWiH2_2),.din(G244));
	jspl3 jspl3_w_G244_1(.douta(w_dff_A_oHNNeNEI2_0),.doutb(w_G244_1[1]),.doutc(w_G244_1[2]),.din(w_G244_0[0]));
	jspl3 jspl3_w_G250_0(.douta(w_dff_A_0Dr2K6jL4_0),.doutb(w_dff_A_c67gaj6g8_1),.doutc(w_G250_0[2]),.din(G250));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_dff_A_l4Toek0g7_1),.doutc(w_dff_A_irs9bHBr5_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_EcODS1TM6_0),.doutb(w_dff_A_TfyK3HW66_1),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G264_0(.douta(w_G264_0[0]),.doutb(w_dff_A_MmzHCcUA0_1),.doutc(w_dff_A_iinwmgc79_2),.din(G264));
	jspl jspl_w_G264_1(.douta(w_G264_1[0]),.doutb(w_G264_1[1]),.din(w_G264_0[0]));
	jspl3 jspl3_w_G270_0(.douta(w_dff_A_vbCK6CD48_0),.doutb(w_G270_0[1]),.doutc(w_G270_0[2]),.din(G270));
	jspl3 jspl3_w_G274_0(.douta(w_dff_A_coUzNFjU0_0),.doutb(w_G274_0[1]),.doutc(w_dff_A_5BzSVzfU8_2),.din(G274));
	jspl3 jspl3_w_G283_0(.douta(w_dff_A_REC5uBRg6_0),.doutb(w_dff_A_zlfUFNxN7_1),.doutc(w_G283_0[2]),.din(G283));
	jspl3 jspl3_w_G283_1(.douta(w_G283_1[0]),.doutb(w_dff_A_0gSbFn020_1),.doutc(w_G283_1[2]),.din(w_G283_0[0]));
	jspl3 jspl3_w_G283_2(.douta(w_dff_A_KSVncrO02_0),.doutb(w_dff_A_cOYiOvKk8_1),.doutc(w_G283_2[2]),.din(w_G283_0[1]));
	jspl3 jspl3_w_G283_3(.douta(w_dff_A_8GO6iolU1_0),.doutb(w_dff_A_U3y76x5D0_1),.doutc(w_G283_3[2]),.din(w_G283_0[2]));
	jspl3 jspl3_w_G294_0(.douta(w_dff_A_IwzbsjN37_0),.doutb(w_dff_A_KiT15BBB8_1),.doutc(w_G294_0[2]),.din(G294));
	jspl3 jspl3_w_G294_1(.douta(w_G294_1[0]),.doutb(w_dff_A_TtR7O4zu8_1),.doutc(w_G294_1[2]),.din(w_G294_0[0]));
	jspl3 jspl3_w_G294_2(.douta(w_dff_A_dWwjfL9n6_0),.doutb(w_G294_2[1]),.doutc(w_G294_2[2]),.din(w_G294_0[1]));
	jspl jspl_w_G294_3(.douta(w_dff_A_GsTMAoUY0_0),.doutb(w_G294_3[1]),.din(w_G294_0[2]));
	jspl3 jspl3_w_G303_0(.douta(w_dff_A_JSgvNSVS9_0),.doutb(w_G303_0[1]),.doutc(w_dff_A_bKPcwFxw3_2),.din(G303));
	jspl3 jspl3_w_G303_1(.douta(w_G303_1[0]),.doutb(w_G303_1[1]),.doutc(w_G303_1[2]),.din(w_G303_0[0]));
	jspl3 jspl3_w_G303_2(.douta(w_dff_A_aqNT9f7j3_0),.doutb(w_dff_A_pNIHpZ1O9_1),.doutc(w_G303_2[2]),.din(w_G303_0[1]));
	jspl3 jspl3_w_G311_0(.douta(w_G311_0[0]),.doutb(w_G311_0[1]),.doutc(w_G311_0[2]),.din(w_dff_B_mqa966gy6_3));
	jspl3 jspl3_w_G311_1(.douta(w_G311_1[0]),.doutb(w_dff_A_Rbqv7i2E2_1),.doutc(w_G311_1[2]),.din(w_G311_0[0]));
	jspl3 jspl3_w_G317_0(.douta(w_G317_0[0]),.doutb(w_G317_0[1]),.doutc(w_G317_0[2]),.din(w_dff_B_shLEtSI70_3));
	jspl jspl_w_G317_1(.douta(w_dff_A_WorGWE6A7_0),.doutb(w_G317_1[1]),.din(w_G317_0[0]));
	jspl3 jspl3_w_G322_0(.douta(w_dff_A_2rrUxUIP9_0),.doutb(w_G322_0[1]),.doutc(w_G322_0[2]),.din(w_dff_B_cWNoaYa40_3));
	jspl jspl_w_G326_0(.douta(w_dff_A_U500Ob7a2_0),.doutb(w_G326_0[1]),.din(w_dff_B_uJt7CJLp2_2));
	jspl jspl_w_G330_0(.douta(w_dff_A_slHywqOc0_0),.doutb(w_G330_0[1]),.din(G330));
	jspl jspl_w_G343_0(.douta(w_G343_0[0]),.doutb(w_dff_A_Su7s7ao33_1),.din(G343));
	jspl3 jspl3_w_G1698_0(.douta(w_G1698_0[0]),.doutb(w_G1698_0[1]),.doutc(w_dff_A_Mlfa3Jcp5_2),.din(G1698));
	jspl jspl_w_G355_0(.douta(w_G355_0),.doutb(w_dff_A_b4JJi3Xo9_1),.din(G355_fa_));
	jspl3 jspl3_w_G396_0(.douta(w_dff_A_i1S5ziKV7_0),.doutb(w_G396_0[1]),.doutc(w_dff_A_JvhgudXb7_2),.din(G396_fa_));
	jspl jspl_w_G384_0(.douta(w_dff_A_ndypIZMF9_0),.doutb(w_dff_A_MK7puvqH4_1),.din(G384_fa_));
	jspl3 jspl3_w_G387_0(.douta(w_G387_0[0]),.doutb(w_G387_0[1]),.doutc(w_dff_A_gMbPIbhZ9_2),.din(G387_fa_));
	jspl3 jspl3_w_n72_0(.douta(w_n72_0[0]),.doutb(w_dff_A_S2bmOonB3_1),.doutc(w_dff_A_FKNrCzj53_2),.din(n72));
	jspl jspl_w_n72_1(.douta(w_n72_1[0]),.doutb(w_dff_A_vGw5cjWo7_1),.din(w_n72_0[0]));
	jspl3 jspl3_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.doutc(w_dff_A_y6OI6irt9_2),.din(n73));
	jspl3 jspl3_w_n73_1(.douta(w_n73_1[0]),.doutb(w_dff_A_6VDFVZtn3_1),.doutc(w_n73_1[2]),.din(w_n73_0[0]));
	jspl3 jspl3_w_n73_2(.douta(w_dff_A_OzhMKkGv7_0),.doutb(w_n73_2[1]),.doutc(w_dff_A_PVARDvkW4_2),.din(w_n73_0[1]));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_dff_A_tPqs1ct78_1),.doutc(w_dff_A_efvVhaa88_2),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_dff_A_h1U14QZ20_1),.doutc(w_dff_A_MwT9xHbC5_2),.din(n75));
	jspl jspl_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.din(w_n75_0[0]));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.din(n76));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl3 jspl3_w_n79_0(.douta(w_dff_A_vIXjKMLs5_0),.doutb(w_n79_0[1]),.doutc(w_n79_0[2]),.din(n79));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_dff_A_ffrbgNc21_1),.doutc(w_dff_A_h6lmthOs1_2),.din(n80));
	jspl jspl_w_n80_1(.douta(w_n80_1[0]),.doutb(w_n80_1[1]),.din(w_n80_0[0]));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_65zy7shZ0_0),.doutb(w_n85_0[1]),.doutc(w_dff_A_HZd2GatY8_2),.din(n85));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n88_0(.douta(w_n88_0[0]),.doutb(w_dff_A_Q14htJgy1_1),.doutc(w_dff_A_UANVtvih1_2),.din(n88));
	jspl jspl_w_n88_1(.douta(w_n88_1[0]),.doutb(w_n88_1[1]),.din(w_n88_0[0]));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_dff_A_PsGS15dS5_1),.doutc(w_n91_0[2]),.din(n91));
	jspl3 jspl3_w_n91_1(.douta(w_dff_A_QS6hAFmE7_0),.doutb(w_n91_1[1]),.doutc(w_n91_1[2]),.din(w_n91_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n97_0(.douta(w_dff_A_swqtA9sL9_0),.doutb(w_n97_0[1]),.doutc(w_n97_0[2]),.din(n97));
	jspl3 jspl3_w_n97_1(.douta(w_n97_1[0]),.doutb(w_dff_A_AZl59P653_1),.doutc(w_n97_1[2]),.din(w_n97_0[0]));
	jspl jspl_w_n97_2(.douta(w_n97_2[0]),.doutb(w_n97_2[1]),.din(w_n97_0[1]));
	jspl3 jspl3_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.doutc(w_n98_0[2]),.din(n98));
	jspl3 jspl3_w_n98_1(.douta(w_dff_A_hEPKzEzv3_0),.doutb(w_dff_A_KVIzA3Ct9_1),.doutc(w_n98_1[2]),.din(w_n98_0[0]));
	jspl jspl_w_n98_2(.douta(w_dff_A_QFqMBReo8_0),.doutb(w_n98_2[1]),.din(w_n98_0[1]));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_6k8eSR7l3_1),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n105_0(.douta(w_dff_A_uDH37AKn4_0),.doutb(w_n105_0[1]),.doutc(w_dff_A_BWR7BzNB9_2),.din(n105));
	jspl3 jspl3_w_n105_1(.douta(w_dff_A_0cZKzsvq7_0),.doutb(w_n105_1[1]),.doutc(w_dff_A_1Sn75JW53_2),.din(w_n105_0[0]));
	jspl jspl_w_n105_2(.douta(w_n105_2[0]),.doutb(w_n105_2[1]),.din(w_n105_0[1]));
	jspl jspl_w_n106_0(.douta(w_dff_A_kgIT8jEI1_0),.doutb(w_n106_0[1]),.din(n106));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl3 jspl3_w_n112_3(.douta(w_dff_A_XCiI2xG81_0),.doutb(w_dff_A_63v7l7Vq9_1),.doutc(w_n112_3[2]),.din(w_n112_0[2]));
	jspl3 jspl3_w_n112_4(.douta(w_dff_A_TxZONEDW8_0),.doutb(w_dff_A_5pCyFonK3_1),.doutc(w_n112_4[2]),.din(w_n112_1[0]));
	jspl3 jspl3_w_n112_5(.douta(w_n112_5[0]),.doutb(w_n112_5[1]),.doutc(w_dff_A_VSlHQ9P36_2),.din(w_n112_1[1]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.doutc(w_n113_0[2]),.din(n113));
	jspl3 jspl3_w_n113_1(.douta(w_dff_A_CoFQTjdU4_0),.doutb(w_dff_A_BFcuhVbu6_1),.doutc(w_n113_1[2]),.din(w_n113_0[0]));
	jspl3 jspl3_w_n113_2(.douta(w_n113_2[0]),.doutb(w_n113_2[1]),.doutc(w_n113_2[2]),.din(w_n113_0[1]));
	jspl jspl_w_n113_3(.douta(w_n113_3[0]),.doutb(w_n113_3[1]),.din(w_n113_0[2]));
	jspl3 jspl3_w_n114_0(.douta(w_n114_0[0]),.doutb(w_dff_A_FoBBaqwL2_1),.doutc(w_n114_0[2]),.din(n114));
	jspl3 jspl3_w_n114_1(.douta(w_dff_A_NG8iqZFU6_0),.doutb(w_n114_1[1]),.doutc(w_n114_1[2]),.din(w_n114_0[0]));
	jspl3 jspl3_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.doutc(w_dff_A_vtqn6Ngn9_2),.din(n115));
	jspl jspl_w_n115_1(.douta(w_n115_1[0]),.doutb(w_n115_1[1]),.din(w_n115_0[0]));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_dff_A_76i7BKoX5_1),.din(n116));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl3 jspl3_w_n121_0(.douta(w_dff_A_o8jC3wy89_0),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.doutc(w_n122_0[2]),.din(n122));
	jspl jspl_w_n122_1(.douta(w_n122_1[0]),.doutb(w_n122_1[1]),.din(w_n122_0[0]));
	jspl3 jspl3_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.doutc(w_n123_0[2]),.din(n123));
	jspl3 jspl3_w_n123_1(.douta(w_n123_1[0]),.doutb(w_n123_1[1]),.doutc(w_n123_1[2]),.din(w_n123_0[0]));
	jspl jspl_w_n131_0(.douta(w_dff_A_6vLKW1ti3_0),.doutb(w_n131_0[1]),.din(n131));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_dff_A_Eux4reDN6_1),.din(n135));
	jspl3 jspl3_w_n137_0(.douta(w_n137_0[0]),.doutb(w_n137_0[1]),.doutc(w_n137_0[2]),.din(n137));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(w_dff_B_C5qcIsB09_2));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_m8wv256D9_1),.doutc(w_dff_A_fLtmlSke3_2),.din(n146));
	jspl3 jspl3_w_n146_1(.douta(w_n146_1[0]),.doutb(w_dff_A_pyxeLgzK9_1),.doutc(w_dff_A_o0x1YyjQ7_2),.din(w_n146_0[0]));
	jspl3 jspl3_w_n146_2(.douta(w_n146_2[0]),.doutb(w_n146_2[1]),.doutc(w_n146_2[2]),.din(w_n146_0[1]));
	jspl3 jspl3_w_n146_3(.douta(w_n146_3[0]),.doutb(w_n146_3[1]),.doutc(w_n146_3[2]),.din(w_n146_0[2]));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_dff_A_slPEs5cW2_1),.doutc(w_dff_A_PQfOk9nx5_2),.din(n147));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_dff_A_jQb7DLmM0_0),.doutb(w_dff_A_BYuIiKA37_1),.doutc(w_n148_1[2]),.din(w_n148_0[0]));
	jspl3 jspl3_w_n148_2(.douta(w_n148_2[0]),.doutb(w_n148_2[1]),.doutc(w_n148_2[2]),.din(w_n148_0[1]));
	jspl3 jspl3_w_n148_3(.douta(w_dff_A_U58CLjyT4_0),.doutb(w_n148_3[1]),.doutc(w_dff_A_bvHmkObR7_2),.din(w_n148_0[2]));
	jspl3 jspl3_w_n148_4(.douta(w_n148_4[0]),.doutb(w_n148_4[1]),.doutc(w_n148_4[2]),.din(w_n148_1[0]));
	jspl3 jspl3_w_n148_5(.douta(w_n148_5[0]),.doutb(w_dff_A_Z4ls5wLR7_1),.doutc(w_dff_A_TLWREQpl6_2),.din(w_n148_1[1]));
	jspl3 jspl3_w_n148_6(.douta(w_n148_6[0]),.doutb(w_n148_6[1]),.doutc(w_n148_6[2]),.din(w_n148_1[2]));
	jspl3 jspl3_w_n148_7(.douta(w_n148_7[0]),.doutb(w_n148_7[1]),.doutc(w_n148_7[2]),.din(w_n148_2[0]));
	jspl3 jspl3_w_n148_8(.douta(w_n148_8[0]),.doutb(w_dff_A_1cQcbg208_1),.doutc(w_n148_8[2]),.din(w_n148_2[1]));
	jspl3 jspl3_w_n148_9(.douta(w_n148_9[0]),.doutb(w_n148_9[1]),.doutc(w_n148_9[2]),.din(w_n148_2[2]));
	jspl3 jspl3_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.doutc(w_n149_0[2]),.din(n149));
	jspl3 jspl3_w_n149_1(.douta(w_n149_1[0]),.doutb(w_dff_A_nhFB6Wdy6_1),.doutc(w_n149_1[2]),.din(w_n149_0[0]));
	jspl jspl_w_n149_2(.douta(w_dff_A_sgKsKajD0_0),.doutb(w_n149_2[1]),.din(w_n149_0[1]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_bZl15ToZ9_1),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_dff_A_kDyzheB88_1),.doutc(w_dff_A_EWytyrHp6_2),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_n151_2[0]),.doutb(w_n151_2[1]),.doutc(w_n151_2[2]),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_dff_A_HOvEmfsF0_0),.doutb(w_dff_A_H6Myhpd09_1),.doutc(w_n151_3[2]),.din(w_n151_0[2]));
	jspl3 jspl3_w_n151_4(.douta(w_n151_4[0]),.doutb(w_n151_4[1]),.doutc(w_dff_A_upYG8lUr4_2),.din(w_n151_1[0]));
	jspl3 jspl3_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.doutc(w_n152_0[2]),.din(n152));
	jspl3 jspl3_w_n152_1(.douta(w_n152_1[0]),.doutb(w_n152_1[1]),.doutc(w_n152_1[2]),.din(w_n152_0[0]));
	jspl3 jspl3_w_n152_2(.douta(w_n152_2[0]),.doutb(w_n152_2[1]),.doutc(w_n152_2[2]),.din(w_n152_0[1]));
	jspl jspl_w_n152_3(.douta(w_n152_3[0]),.doutb(w_n152_3[1]),.din(w_n152_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(n154));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl3 jspl3_w_n155_1(.douta(w_n155_1[0]),.doutb(w_n155_1[1]),.doutc(w_n155_1[2]),.din(w_n155_0[0]));
	jspl3 jspl3_w_n155_2(.douta(w_n155_2[0]),.doutb(w_n155_2[1]),.doutc(w_n155_2[2]),.din(w_n155_0[1]));
	jspl jspl_w_n155_3(.douta(w_n155_3[0]),.doutb(w_n155_3[1]),.din(w_n155_0[2]));
	jspl3 jspl3_w_n157_0(.douta(w_dff_A_GHAbKBh17_0),.doutb(w_n157_0[1]),.doutc(w_dff_A_tcKA3BhQ5_2),.din(n157));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_dff_A_pIExNAhw0_2),.din(n161));
	jspl jspl_w_n161_1(.douta(w_n161_1[0]),.doutb(w_n161_1[1]),.din(w_n161_0[0]));
	jspl3 jspl3_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.doutc(w_n162_0[2]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_dff_A_hTYt0Sei3_0),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_dff_A_oSJIeN5g9_1),.doutc(w_dff_A_0HjbQwMa6_2),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_dff_A_EhSyXoq93_2),.din(w_n166_0[1]));
	jspl jspl_w_n166_3(.douta(w_dff_A_UAPhG3Vn9_0),.doutb(w_n166_3[1]),.din(w_n166_0[2]));
	jspl3 jspl3_w_n170_0(.douta(w_dff_A_4Ouj8ThX9_0),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(w_dff_B_mCDef9Oe5_2));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_dff_A_jPwCkNEH8_1),.doutc(w_dff_A_F7j5jKl69_2),.din(n179));
	jspl3 jspl3_w_n179_1(.douta(w_n179_1[0]),.doutb(w_n179_1[1]),.doutc(w_n179_1[2]),.din(w_n179_0[0]));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.doutc(w_n185_0[2]),.din(n185));
	jspl3 jspl3_w_n185_1(.douta(w_n185_1[0]),.doutb(w_n185_1[1]),.doutc(w_dff_A_Nwsjq0xo4_2),.din(w_n185_0[0]));
	jspl3 jspl3_w_n185_2(.douta(w_n185_2[0]),.doutb(w_dff_A_jBWtepp39_1),.doutc(w_n185_2[2]),.din(w_n185_0[1]));
	jspl3 jspl3_w_n185_3(.douta(w_n185_3[0]),.doutb(w_n185_3[1]),.doutc(w_n185_3[2]),.din(w_n185_0[2]));
	jspl3 jspl3_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.doutc(w_dff_A_ObhdSrtI1_2),.din(n189));
	jspl3 jspl3_w_n189_1(.douta(w_n189_1[0]),.doutb(w_dff_A_BAlsuDBm7_1),.doutc(w_n189_1[2]),.din(w_n189_0[0]));
	jspl jspl_w_n189_2(.douta(w_dff_A_bYTrrIyV4_0),.doutb(w_n189_2[1]),.din(w_n189_0[1]));
	jspl3 jspl3_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.doutc(w_n190_0[2]),.din(n190));
	jspl3 jspl3_w_n190_1(.douta(w_n190_1[0]),.doutb(w_dff_A_BhaIHiIi3_1),.doutc(w_n190_1[2]),.din(w_n190_0[0]));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_dff_A_ZTcFboHJ9_0),.doutb(w_n196_0[1]),.doutc(w_dff_A_JFjoZqRm7_2),.din(w_dff_B_kIJv506o1_3));
	jspl3 jspl3_w_n196_1(.douta(w_dff_A_pH3RywLK4_0),.doutb(w_dff_A_mgJE9RLR9_1),.doutc(w_n196_1[2]),.din(w_n196_0[0]));
	jspl3 jspl3_w_n196_2(.douta(w_dff_A_PWuV5Axc5_0),.doutb(w_dff_A_VCFA39Bw3_1),.doutc(w_n196_2[2]),.din(w_n196_0[1]));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_n197_1[0]),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n199_1(.douta(w_n199_1[0]),.doutb(w_n199_1[1]),.din(w_n199_0[0]));
	jspl jspl_w_n201_0(.douta(w_dff_A_mVCFVMyS7_0),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n205_0(.douta(w_dff_A_PbvQEbvw8_0),.doutb(w_n205_0[1]),.din(w_dff_B_6KcOzGgC9_2));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl3 jspl3_w_n210_0(.douta(w_dff_A_hz48tvZj2_0),.doutb(w_n210_0[1]),.doutc(w_n210_0[2]),.din(n210));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_dff_A_0M59mrjU1_1),.din(n213));
	jspl jspl_w_n214_0(.douta(w_n214_0[0]),.doutb(w_dff_A_4kFVSjYh8_1),.din(n214));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl3 jspl3_w_n221_0(.douta(w_dff_A_3xRNxzVm0_0),.doutb(w_dff_A_zzM06KLE7_1),.doutc(w_n221_0[2]),.din(n221));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_dff_A_DtA0yE6o6_1),.din(n228));
	jspl3 jspl3_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.doutc(w_n229_0[2]),.din(n229));
	jspl jspl_w_n230_0(.douta(w_dff_A_MjqUp2IV7_0),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.doutc(w_n231_0[2]),.din(n231));
	jspl3 jspl3_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.doutc(w_n234_0[2]),.din(n234));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(n241));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl jspl_w_n246_1(.douta(w_n246_1[0]),.doutb(w_n246_1[1]),.din(w_n246_0[0]));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_ZgjgcbpT5_2));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_dff_A_DIxhcRxu7_1),.din(n255));
	jspl jspl_w_n257_0(.douta(w_dff_A_Esk9FLPn0_0),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n259_0(.douta(w_dff_A_v7wVNXzV8_0),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n262_0(.douta(w_dff_A_AribFjuc2_0),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.doutc(w_n269_1[2]),.din(w_n269_0[0]));
	jspl jspl_w_n270_0(.douta(w_dff_A_g5LRjXiN1_0),.doutb(w_n270_0[1]),.din(w_dff_B_SP53AS286_2));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_n271_1[0]),.doutb(w_n271_1[1]),.doutc(w_n271_1[2]),.din(w_n271_0[0]));
	jspl3 jspl3_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_Wl9EksWk0_1),.doutc(w_n274_0[2]),.din(n274));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(n278));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(n279));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_dff_A_1Aer3cB25_1),.din(n281));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n288_1(.douta(w_n288_1[0]),.doutb(w_n288_1[1]),.din(w_n288_0[0]));
	jspl jspl_w_n296_0(.douta(w_dff_A_3zW65Z0I5_0),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n298_0(.douta(w_dff_A_gFIWSjUS3_0),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_dff_A_8bu2HjsL3_1),.din(n300));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_O5qOvHQS3_1),.din(n303));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_dff_A_kyk90hop2_1),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n334_0(.douta(w_dff_A_luOPKde94_0),.doutb(w_n334_0[1]),.din(n334));
	jspl jspl_w_n339_0(.douta(w_dff_A_S9HSg5NO7_0),.doutb(w_n339_0[1]),.din(n339));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl jspl_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.din(w_n355_0[0]));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_dff_A_OLc4brm52_1),.din(n374));
	jspl jspl_w_n381_0(.douta(w_n381_0[0]),.doutb(w_n381_0[1]),.din(n381));
	jspl3 jspl3_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.doutc(w_n382_0[2]),.din(n382));
	jspl jspl_w_n382_1(.douta(w_n382_1[0]),.doutb(w_n382_1[1]),.din(w_n382_0[0]));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl jspl_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(w_dff_B_MPLAYylK2_2));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_dff_A_NuGbAMwL1_1),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n407_0(.douta(w_n407_0[0]),.doutb(w_dff_A_rM0bwNhF2_1),.doutc(w_dff_A_iI3BAws32_2),.din(n407));
	jspl3 jspl3_w_n407_1(.douta(w_dff_A_Zn9s1wEB5_0),.doutb(w_dff_A_ZwLwUUqu8_1),.doutc(w_n407_1[2]),.din(w_n407_0[0]));
	jspl jspl_w_n407_2(.douta(w_n407_2[0]),.doutb(w_n407_2[1]),.din(w_n407_0[1]));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(n412));
	jspl3 jspl3_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jspl jspl_w_n420_1(.douta(w_n420_1[0]),.doutb(w_n420_1[1]),.din(w_n420_0[0]));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_dff_A_juqvY5ge5_1),.doutc(w_dff_A_Srm5kXMA6_2),.din(n425));
	jspl3 jspl3_w_n425_1(.douta(w_dff_A_U1nsvXFK9_0),.doutb(w_dff_A_01HEKiPv4_1),.doutc(w_n425_1[2]),.din(w_n425_0[0]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl jspl_w_n430_0(.douta(w_dff_A_JFeIDYY74_0),.doutb(w_n430_0[1]),.din(w_dff_B_C0Fl309u4_2));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_dff_A_2IVlRPjg5_1),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_dff_A_Czkz7sXW1_1),.doutc(w_n439_0[2]),.din(n439));
	jspl jspl_w_n439_1(.douta(w_n439_1[0]),.doutb(w_n439_1[1]),.din(w_n439_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl3 jspl3_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.doutc(w_n455_0[2]),.din(n455));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(n474));
	jspl jspl_w_n475_0(.douta(w_n475_0[0]),.doutb(w_n475_0[1]),.din(n475));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(n479));
	jspl jspl_w_n483_0(.douta(w_dff_A_OF2BZT4e7_0),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl3 jspl3_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.doutc(w_n492_0[2]),.din(n492));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n516_0(.douta(w_dff_A_Kv3wMfzj6_0),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n519_0(.douta(w_n519_0[0]),.doutb(w_dff_A_Qbg4QAcq7_1),.doutc(w_dff_A_tidmV6Lo7_2),.din(n519));
	jspl3 jspl3_w_n519_1(.douta(w_dff_A_Tqa4XRTQ6_0),.doutb(w_n519_1[1]),.doutc(w_n519_1[2]),.din(w_n519_0[0]));
	jspl jspl_w_n523_0(.douta(w_dff_A_Uky4l53N4_0),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_dff_A_IHmCwTyd5_1),.din(n524));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_dff_A_lrS1MQPf1_1),.din(n532));
	jspl jspl_w_n534_0(.douta(w_dff_A_Ym3uFM6E0_0),.doutb(w_n534_0[1]),.din(n534));
	jspl3 jspl3_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.doutc(w_n536_0[2]),.din(n536));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_dff_A_H2zRB4zY0_1),.din(n541));
	jspl3 jspl3_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.doutc(w_n542_0[2]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n548_0(.douta(w_dff_A_fjKKoOcc0_0),.doutb(w_n548_0[1]),.doutc(w_n548_0[2]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl3 jspl3_w_n552_0(.douta(w_n552_0[0]),.doutb(w_dff_A_YGVxfLki0_1),.doutc(w_dff_A_q1KHmSbO4_2),.din(n552));
	jspl jspl_w_n552_1(.douta(w_n552_1[0]),.doutb(w_n552_1[1]),.din(w_n552_0[0]));
	jspl3 jspl3_w_n553_0(.douta(w_dff_A_TEJfY3zX3_0),.doutb(w_n553_0[1]),.doutc(w_dff_A_sHrhhkQJ2_2),.din(n553));
	jspl3 jspl3_w_n553_1(.douta(w_n553_1[0]),.doutb(w_n553_1[1]),.doutc(w_n553_1[2]),.din(w_n553_0[0]));
	jspl3 jspl3_w_n553_2(.douta(w_dff_A_1IoTyaGF1_0),.doutb(w_dff_A_SgKpglzj9_1),.doutc(w_n553_2[2]),.din(w_n553_0[1]));
	jspl3 jspl3_w_n554_0(.douta(w_dff_A_P8mMtLYv0_0),.doutb(w_dff_A_hMeOEyx59_1),.doutc(w_n554_0[2]),.din(w_dff_B_4euaslRD6_3));
	jspl3 jspl3_w_n554_1(.douta(w_n554_1[0]),.doutb(w_n554_1[1]),.doutc(w_dff_A_fzv4lvqZ5_2),.din(w_n554_0[0]));
	jspl3 jspl3_w_n554_2(.douta(w_n554_2[0]),.doutb(w_dff_A_bXVRJXjo6_1),.doutc(w_dff_A_4iVzRieL8_2),.din(w_n554_0[1]));
	jspl3 jspl3_w_n554_3(.douta(w_n554_3[0]),.doutb(w_dff_A_TXHv3qj30_1),.doutc(w_dff_A_YFww9s9J9_2),.din(w_n554_0[2]));
	jspl jspl_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.din(w_dff_B_6XuEDFwA5_2));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl3 jspl3_w_n563_0(.douta(w_n563_0[0]),.doutb(w_dff_A_phdcRowx4_1),.doutc(w_dff_A_qh0ueVTK0_2),.din(n563));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_XSZpSyWq1_1),.din(n564));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(w_dff_B_9D8UaAZR2_2));
	jspl jspl_w_n567_0(.douta(w_dff_A_cJa5wY6U9_0),.doutb(w_n567_0[1]),.din(n567));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_n571_0[2]),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n576_1(.douta(w_n576_1[0]),.doutb(w_n576_1[1]),.din(w_n576_0[0]));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_dff_A_ufRxWv6b1_2),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n589_0(.douta(w_n589_0[0]),.doutb(w_n589_0[1]),.doutc(w_n589_0[2]),.din(n589));
	jspl3 jspl3_w_n589_1(.douta(w_dff_A_0YiUR0Ss4_0),.doutb(w_n589_1[1]),.doutc(w_n589_1[2]),.din(w_n589_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_dff_A_P99KkVrv0_1),.doutc(w_dff_A_9oa9JSFi3_2),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_dff_A_KNHB5mhX4_0),.doutb(w_n592_0[1]),.doutc(w_dff_A_pbO59dpv8_2),.din(n592));
	jspl3 jspl3_w_n592_1(.douta(w_dff_A_8VaEDlcY7_0),.doutb(w_dff_A_Iq24XGYr3_1),.doutc(w_n592_1[2]),.din(w_n592_0[0]));
	jspl jspl_w_n592_2(.douta(w_n592_2[0]),.doutb(w_n592_2[1]),.din(w_n592_0[1]));
	jspl3 jspl3_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.doutc(w_n593_0[2]),.din(n593));
	jspl jspl_w_n602_0(.douta(w_dff_A_hhWxJAtF1_0),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n603_0(.douta(w_dff_A_4RRiHoEs0_0),.doutb(w_n603_0[1]),.doutc(w_dff_A_NMzqwxXi2_2),.din(n603));
	jspl3 jspl3_w_n603_1(.douta(w_dff_A_P4ZigKiT8_0),.doutb(w_n603_1[1]),.doutc(w_n603_1[2]),.din(w_n603_0[0]));
	jspl jspl_w_n603_2(.douta(w_dff_A_UeTQRlg70_0),.doutb(w_n603_2[1]),.din(w_n603_0[1]));
	jspl3 jspl3_w_n604_0(.douta(w_dff_A_DHZW8wk15_0),.doutb(w_n604_0[1]),.doutc(w_dff_A_9f9VqMzN8_2),.din(n604));
	jspl3 jspl3_w_n604_1(.douta(w_dff_A_i5Ds5bN29_0),.doutb(w_n604_1[1]),.doutc(w_dff_A_OSkJvifp7_2),.din(w_n604_0[0]));
	jspl jspl_w_n604_2(.douta(w_dff_A_kKrqoSoW7_0),.doutb(w_n604_2[1]),.din(w_n604_0[1]));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_dff_A_a5wMNEEO6_2),.din(w_n605_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_dff_A_NoSDn8eT1_1),.doutc(w_dff_A_BxA3UUOd6_2),.din(n608));
	jspl3 jspl3_w_n608_1(.douta(w_dff_A_TGBdpbH83_0),.doutb(w_n608_1[1]),.doutc(w_dff_A_VPwrvW8B8_2),.din(w_n608_0[0]));
	jspl3 jspl3_w_n612_0(.douta(w_n612_0[0]),.doutb(w_dff_A_UZVNZD1m5_1),.doutc(w_n612_0[2]),.din(n612));
	jspl3 jspl3_w_n612_1(.douta(w_dff_A_sSARz3Q60_0),.doutb(w_dff_A_qpAvnoHG2_1),.doutc(w_n612_1[2]),.din(w_n612_0[0]));
	jspl3 jspl3_w_n612_2(.douta(w_n612_2[0]),.doutb(w_n612_2[1]),.doutc(w_n612_2[2]),.din(w_n612_0[1]));
	jspl3 jspl3_w_n612_3(.douta(w_dff_A_bOjiu0b69_0),.doutb(w_n612_3[1]),.doutc(w_dff_A_dBm7to3B0_2),.din(w_n612_0[2]));
	jspl jspl_w_n612_4(.douta(w_n612_4[0]),.doutb(w_dff_A_fKgJXFjY1_1),.din(w_n612_1[0]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl jspl_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.din(w_n613_0[0]));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_dff_A_O0F2LtgJ8_1),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl3 jspl3_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.doutc(w_n617_1[2]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n617_2(.douta(w_n617_2[0]),.doutb(w_n617_2[1]),.doutc(w_n617_2[2]),.din(w_n617_0[1]));
	jspl3 jspl3_w_n617_3(.douta(w_n617_3[0]),.doutb(w_n617_3[1]),.doutc(w_n617_3[2]),.din(w_n617_0[2]));
	jspl3 jspl3_w_n617_4(.douta(w_n617_4[0]),.doutb(w_n617_4[1]),.doutc(w_n617_4[2]),.din(w_n617_1[0]));
	jspl3 jspl3_w_n617_5(.douta(w_n617_5[0]),.doutb(w_n617_5[1]),.doutc(w_n617_5[2]),.din(w_n617_1[1]));
	jspl jspl_w_n617_6(.douta(w_n617_6[0]),.doutb(w_n617_6[1]),.din(w_n617_1[2]));
	jspl jspl_w_n619_0(.douta(w_dff_A_V3ymdB0E2_0),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl3 jspl3_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.doutc(w_n623_0[2]),.din(n623));
	jspl3 jspl3_w_n623_1(.douta(w_n623_1[0]),.doutb(w_n623_1[1]),.doutc(w_n623_1[2]),.din(w_n623_0[0]));
	jspl3 jspl3_w_n623_2(.douta(w_n623_2[0]),.doutb(w_n623_2[1]),.doutc(w_n623_2[2]),.din(w_n623_0[1]));
	jspl3 jspl3_w_n623_3(.douta(w_n623_3[0]),.doutb(w_n623_3[1]),.doutc(w_n623_3[2]),.din(w_n623_0[2]));
	jspl3 jspl3_w_n623_4(.douta(w_n623_4[0]),.doutb(w_n623_4[1]),.doutc(w_n623_4[2]),.din(w_n623_1[0]));
	jspl jspl_w_n623_5(.douta(w_n623_5[0]),.doutb(w_n623_5[1]),.din(w_n623_1[1]));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(n626));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl3 jspl3_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.doutc(w_n627_1[2]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n627_2(.douta(w_n627_2[0]),.doutb(w_n627_2[1]),.doutc(w_n627_2[2]),.din(w_n627_0[1]));
	jspl3 jspl3_w_n627_3(.douta(w_n627_3[0]),.doutb(w_n627_3[1]),.doutc(w_n627_3[2]),.din(w_n627_0[2]));
	jspl3 jspl3_w_n627_4(.douta(w_n627_4[0]),.doutb(w_n627_4[1]),.doutc(w_n627_4[2]),.din(w_n627_1[0]));
	jspl3 jspl3_w_n627_5(.douta(w_n627_5[0]),.doutb(w_n627_5[1]),.doutc(w_n627_5[2]),.din(w_n627_1[1]));
	jspl3 jspl3_w_n627_6(.douta(w_n627_6[0]),.doutb(w_n627_6[1]),.doutc(w_n627_6[2]),.din(w_n627_1[2]));
	jspl jspl_w_n627_7(.douta(w_n627_7[0]),.doutb(w_n627_7[1]),.din(w_n627_2[0]));
	jspl3 jspl3_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.doutc(w_n631_0[2]),.din(n631));
	jspl3 jspl3_w_n631_1(.douta(w_n631_1[0]),.doutb(w_n631_1[1]),.doutc(w_n631_1[2]),.din(w_n631_0[0]));
	jspl3 jspl3_w_n631_2(.douta(w_n631_2[0]),.doutb(w_n631_2[1]),.doutc(w_n631_2[2]),.din(w_n631_0[1]));
	jspl3 jspl3_w_n631_3(.douta(w_n631_3[0]),.doutb(w_n631_3[1]),.doutc(w_n631_3[2]),.din(w_n631_0[2]));
	jspl3 jspl3_w_n631_4(.douta(w_n631_4[0]),.doutb(w_n631_4[1]),.doutc(w_n631_4[2]),.din(w_n631_1[0]));
	jspl3 jspl3_w_n631_5(.douta(w_n631_5[0]),.doutb(w_n631_5[1]),.doutc(w_n631_5[2]),.din(w_n631_1[1]));
	jspl3 jspl3_w_n631_6(.douta(w_n631_6[0]),.doutb(w_n631_6[1]),.doutc(w_n631_6[2]),.din(w_n631_1[2]));
	jspl jspl_w_n631_7(.douta(w_n631_7[0]),.doutb(w_n631_7[1]),.din(w_n631_2[0]));
	jspl3 jspl3_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.doutc(w_n634_0[2]),.din(n634));
	jspl3 jspl3_w_n634_1(.douta(w_n634_1[0]),.doutb(w_n634_1[1]),.doutc(w_n634_1[2]),.din(w_n634_0[0]));
	jspl3 jspl3_w_n634_2(.douta(w_n634_2[0]),.doutb(w_n634_2[1]),.doutc(w_n634_2[2]),.din(w_n634_0[1]));
	jspl3 jspl3_w_n634_3(.douta(w_n634_3[0]),.doutb(w_n634_3[1]),.doutc(w_n634_3[2]),.din(w_n634_0[2]));
	jspl jspl_w_n634_4(.douta(w_n634_4[0]),.doutb(w_n634_4[1]),.din(w_n634_1[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n636_1(.douta(w_n636_1[0]),.doutb(w_n636_1[1]),.doutc(w_n636_1[2]),.din(w_n636_0[0]));
	jspl3 jspl3_w_n636_2(.douta(w_n636_2[0]),.doutb(w_n636_2[1]),.doutc(w_n636_2[2]),.din(w_n636_0[1]));
	jspl3 jspl3_w_n636_3(.douta(w_n636_3[0]),.doutb(w_n636_3[1]),.doutc(w_n636_3[2]),.din(w_n636_0[2]));
	jspl3 jspl3_w_n636_4(.douta(w_n636_4[0]),.doutb(w_n636_4[1]),.doutc(w_n636_4[2]),.din(w_n636_1[0]));
	jspl3 jspl3_w_n636_5(.douta(w_n636_5[0]),.doutb(w_n636_5[1]),.doutc(w_n636_5[2]),.din(w_n636_1[1]));
	jspl3 jspl3_w_n636_6(.douta(w_n636_6[0]),.doutb(w_n636_6[1]),.doutc(w_n636_6[2]),.din(w_n636_1[2]));
	jspl jspl_w_n636_7(.douta(w_n636_7[0]),.doutb(w_n636_7[1]),.din(w_n636_2[0]));
	jspl jspl_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.din(n639));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl3 jspl3_w_n640_2(.douta(w_n640_2[0]),.doutb(w_n640_2[1]),.doutc(w_n640_2[2]),.din(w_n640_0[1]));
	jspl3 jspl3_w_n640_3(.douta(w_n640_3[0]),.doutb(w_n640_3[1]),.doutc(w_n640_3[2]),.din(w_n640_0[2]));
	jspl3 jspl3_w_n640_4(.douta(w_n640_4[0]),.doutb(w_n640_4[1]),.doutc(w_n640_4[2]),.din(w_n640_1[0]));
	jspl3 jspl3_w_n640_5(.douta(w_n640_5[0]),.doutb(w_n640_5[1]),.doutc(w_n640_5[2]),.din(w_n640_1[1]));
	jspl3 jspl3_w_n640_6(.douta(w_n640_6[0]),.doutb(w_n640_6[1]),.doutc(w_n640_6[2]),.din(w_n640_1[2]));
	jspl jspl_w_n640_7(.douta(w_n640_7[0]),.doutb(w_n640_7[1]),.din(w_n640_2[0]));
	jspl3 jspl3_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.doutc(w_n642_0[2]),.din(n642));
	jspl3 jspl3_w_n642_1(.douta(w_n642_1[0]),.doutb(w_n642_1[1]),.doutc(w_n642_1[2]),.din(w_n642_0[0]));
	jspl3 jspl3_w_n642_2(.douta(w_n642_2[0]),.doutb(w_n642_2[1]),.doutc(w_n642_2[2]),.din(w_n642_0[1]));
	jspl3 jspl3_w_n642_3(.douta(w_n642_3[0]),.doutb(w_n642_3[1]),.doutc(w_n642_3[2]),.din(w_n642_0[2]));
	jspl3 jspl3_w_n642_4(.douta(w_n642_4[0]),.doutb(w_n642_4[1]),.doutc(w_n642_4[2]),.din(w_n642_1[0]));
	jspl3 jspl3_w_n642_5(.douta(w_n642_5[0]),.doutb(w_n642_5[1]),.doutc(w_n642_5[2]),.din(w_n642_1[1]));
	jspl3 jspl3_w_n642_6(.douta(w_n642_6[0]),.doutb(w_n642_6[1]),.doutc(w_n642_6[2]),.din(w_n642_1[2]));
	jspl jspl_w_n642_7(.douta(w_n642_7[0]),.doutb(w_n642_7[1]),.din(w_n642_2[0]));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(n654));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl3 jspl3_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.doutc(w_dff_A_s4K4jVzF7_2),.din(n672));
	jspl jspl_w_n672_1(.douta(w_n672_1[0]),.doutb(w_dff_A_7SeFFzao1_1),.din(w_n672_0[0]));
	jspl3 jspl3_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.doutc(w_n675_0[2]),.din(n675));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(w_dff_B_wnaAccVc0_2));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_dff_A_Im8C63OO4_1),.din(w_dff_B_cMsoc7sh1_2));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_dff_A_TBk7QCdd1_1),.doutc(w_n696_0[2]),.din(n696));
	jspl3 jspl3_w_n696_1(.douta(w_dff_A_FCrx7MFn5_0),.doutb(w_n696_1[1]),.doutc(w_dff_A_LzAARKpC1_2),.din(w_n696_0[0]));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.doutc(w_n743_0[2]),.din(n743));
	jspl jspl_w_n743_1(.douta(w_n743_1[0]),.doutb(w_n743_1[1]),.din(w_n743_0[0]));
	jspl jspl_w_n750_0(.douta(w_dff_A_cIUoVB911_0),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n754_0(.douta(w_dff_A_7ay8bsDi0_0),.doutb(w_n754_0[1]),.din(n754));
	jspl3 jspl3_w_n758_0(.douta(w_dff_A_wMvQFKzl8_0),.doutb(w_dff_A_qmBZvkLz6_1),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n758_1(.douta(w_n758_1[0]),.doutb(w_dff_A_XQEGH7Fg5_1),.din(w_n758_0[0]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_dff_A_3xcn83Zx7_0),.doutb(w_n760_0[1]),.din(n760));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_dff_A_Lohcljm11_2),.din(n764));
	jspl3 jspl3_w_n764_1(.douta(w_n764_1[0]),.doutb(w_n764_1[1]),.doutc(w_dff_A_FQjyNBXB6_2),.din(w_n764_0[0]));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_n771_0[2]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_dff_A_3ErFUkCU3_0),.doutb(w_n779_0[1]),.din(n779));
	jspl jspl_w_n797_0(.douta(w_dff_A_JPVkXb1c2_0),.doutb(w_n797_0[1]),.din(n797));
	jspl jspl_w_n801_0(.douta(w_dff_A_4UiU7fNk1_0),.doutb(w_n801_0[1]),.din(n801));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl3 jspl3_w_n853_0(.douta(w_n853_0[0]),.doutb(w_n853_0[1]),.doutc(w_n853_0[2]),.din(n853));
	jspl3 jspl3_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.doutc(w_n855_0[2]),.din(n855));
	jspl3 jspl3_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.doutc(w_dff_A_R0rFJcId8_2),.din(n861));
	jspl jspl_w_n861_1(.douta(w_n861_1[0]),.doutb(w_dff_A_RyHrEmPo5_1),.din(w_n861_0[0]));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.din(n863));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_dff_A_aDjpHZsX8_1),.din(n899));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl3 jspl3_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.doutc(w_n937_0[2]),.din(n937));
	jspl jspl_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.din(n940));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_dff_A_snOCCsqR1_1),.din(n962));
	jspl3 jspl3_w_n988_0(.douta(w_dff_A_fyeVzkVI3_0),.doutb(w_dff_A_O5BkJj945_1),.doutc(w_n988_0[2]),.din(n988));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_dff_A_7FpSlnU95_1),.din(n990));
	jspl3 jspl3_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.doutc(w_n991_0[2]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_dff_A_zVexCDq21_1),.din(n999));
	jspl3 jspl3_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.doutc(w_n1001_0[2]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.doutc(w_n1002_0[2]),.din(n1002));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl3 jspl3_w_n1049_0(.douta(w_dff_A_pbWzgCyS4_0),.doutb(w_dff_A_qpemC9y70_1),.doutc(w_n1049_0[2]),.din(n1049));
	jspl jspl_w_n1052_0(.douta(w_dff_A_qQrMKb5R0_0),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_dff_A_gRcrxL502_1),.din(n1057));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(n1059));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl3 jspl3_w_n1162_0(.douta(w_n1162_0[0]),.doutb(w_dff_A_5O7iKcwa2_1),.doutc(w_n1162_0[2]),.din(n1162));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(n1164));
	jspl jspl_w_n1172_0(.douta(w_dff_A_1gHWTp1M2_0),.doutb(w_n1172_0[1]),.din(n1172));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_dff_A_PBO6IMgf3_1),.din(n1175));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_dff_A_mU4FV3g02_1),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_dff_A_2gFj4f353_0),.doutb(w_n1184_0[1]),.din(n1184));
	jspl jspl_w_n1187_0(.douta(w_dff_A_75qdFNfU4_0),.doutb(w_n1187_0[1]),.din(n1187));
	jdff dff_B_ZbIvEJMZ1_1(.din(n111),.dout(w_dff_B_ZbIvEJMZ1_1),.clk(gclk));
	jdff dff_B_RKYEFx1F2_0(.din(n126),.dout(w_dff_B_RKYEFx1F2_0),.clk(gclk));
	jdff dff_B_XAQHaUNc9_0(.din(n125),.dout(w_dff_B_XAQHaUNc9_0),.clk(gclk));
	jdff dff_A_35iZO2qL7_1(.dout(w_n72_1[1]),.din(w_dff_A_35iZO2qL7_1),.clk(gclk));
	jdff dff_A_vGw5cjWo7_1(.dout(w_dff_A_35iZO2qL7_1),.din(w_dff_A_vGw5cjWo7_1),.clk(gclk));
	jdff dff_A_QFqMBReo8_0(.dout(w_n98_2[0]),.din(w_dff_A_QFqMBReo8_0),.clk(gclk));
	jdff dff_B_TiI7vb9P6_1(.din(n540),.dout(w_dff_B_TiI7vb9P6_1),.clk(gclk));
	jdff dff_B_57HSYb0W9_0(.din(n597),.dout(w_dff_B_57HSYb0W9_0),.clk(gclk));
	jdff dff_B_gqmF82y40_0(.din(w_dff_B_57HSYb0W9_0),.dout(w_dff_B_gqmF82y40_0),.clk(gclk));
	jdff dff_B_FqyPStGC8_0(.din(w_dff_B_gqmF82y40_0),.dout(w_dff_B_FqyPStGC8_0),.clk(gclk));
	jdff dff_B_bR07qUFD3_0(.din(w_dff_B_FqyPStGC8_0),.dout(w_dff_B_bR07qUFD3_0),.clk(gclk));
	jdff dff_B_fekINiU85_0(.din(w_dff_B_bR07qUFD3_0),.dout(w_dff_B_fekINiU85_0),.clk(gclk));
	jdff dff_B_FfPOBCUt9_0(.din(w_dff_B_fekINiU85_0),.dout(w_dff_B_FfPOBCUt9_0),.clk(gclk));
	jdff dff_B_Txu07bCc5_0(.din(w_dff_B_FfPOBCUt9_0),.dout(w_dff_B_Txu07bCc5_0),.clk(gclk));
	jdff dff_B_oyBfdrSg1_0(.din(w_dff_B_Txu07bCc5_0),.dout(w_dff_B_oyBfdrSg1_0),.clk(gclk));
	jdff dff_B_pnhV1Ahu7_0(.din(w_dff_B_oyBfdrSg1_0),.dout(w_dff_B_pnhV1Ahu7_0),.clk(gclk));
	jdff dff_B_aW8cQsyk1_0(.din(w_dff_B_pnhV1Ahu7_0),.dout(w_dff_B_aW8cQsyk1_0),.clk(gclk));
	jdff dff_B_30hQyZDl3_0(.din(n596),.dout(w_dff_B_30hQyZDl3_0),.clk(gclk));
	jdff dff_B_z4aZpyvY0_0(.din(n795),.dout(w_dff_B_z4aZpyvY0_0),.clk(gclk));
	jdff dff_B_r7GeDUeT2_0(.din(w_dff_B_z4aZpyvY0_0),.dout(w_dff_B_r7GeDUeT2_0),.clk(gclk));
	jdff dff_B_eRMJhjTK0_0(.din(w_dff_B_r7GeDUeT2_0),.dout(w_dff_B_eRMJhjTK0_0),.clk(gclk));
	jdff dff_B_zRFfzQZT1_0(.din(w_dff_B_eRMJhjTK0_0),.dout(w_dff_B_zRFfzQZT1_0),.clk(gclk));
	jdff dff_B_GrKdLDr06_0(.din(w_dff_B_zRFfzQZT1_0),.dout(w_dff_B_GrKdLDr06_0),.clk(gclk));
	jdff dff_B_wUJghsZH9_0(.din(w_dff_B_GrKdLDr06_0),.dout(w_dff_B_wUJghsZH9_0),.clk(gclk));
	jdff dff_B_KIZG7nLE8_0(.din(w_dff_B_wUJghsZH9_0),.dout(w_dff_B_KIZG7nLE8_0),.clk(gclk));
	jdff dff_B_F9VlwxNV5_0(.din(w_dff_B_KIZG7nLE8_0),.dout(w_dff_B_F9VlwxNV5_0),.clk(gclk));
	jdff dff_B_0prqLHRs9_0(.din(w_dff_B_F9VlwxNV5_0),.dout(w_dff_B_0prqLHRs9_0),.clk(gclk));
	jdff dff_B_3vzv6ll53_0(.din(w_dff_B_0prqLHRs9_0),.dout(w_dff_B_3vzv6ll53_0),.clk(gclk));
	jdff dff_B_1o8dJWyL5_0(.din(w_dff_B_3vzv6ll53_0),.dout(w_dff_B_1o8dJWyL5_0),.clk(gclk));
	jdff dff_B_iS3n88y91_0(.din(w_dff_B_1o8dJWyL5_0),.dout(w_dff_B_iS3n88y91_0),.clk(gclk));
	jdff dff_B_gRaPGDVy3_0(.din(w_dff_B_iS3n88y91_0),.dout(w_dff_B_gRaPGDVy3_0),.clk(gclk));
	jdff dff_B_3ciAPUTD0_0(.din(w_dff_B_gRaPGDVy3_0),.dout(w_dff_B_3ciAPUTD0_0),.clk(gclk));
	jdff dff_B_abRt2R1v3_0(.din(w_dff_B_3ciAPUTD0_0),.dout(w_dff_B_abRt2R1v3_0),.clk(gclk));
	jdff dff_B_7uld260A0_0(.din(w_dff_B_abRt2R1v3_0),.dout(w_dff_B_7uld260A0_0),.clk(gclk));
	jdff dff_B_iHgZDsFN1_0(.din(w_dff_B_7uld260A0_0),.dout(w_dff_B_iHgZDsFN1_0),.clk(gclk));
	jdff dff_B_S17TyMTG2_1(.din(n791),.dout(w_dff_B_S17TyMTG2_1),.clk(gclk));
	jdff dff_B_ucJF10Ej6_0(.din(n793),.dout(w_dff_B_ucJF10Ej6_0),.clk(gclk));
	jdff dff_B_oaMhJkbn7_0(.din(w_dff_B_ucJF10Ej6_0),.dout(w_dff_B_oaMhJkbn7_0),.clk(gclk));
	jdff dff_B_bgnk8CN45_0(.din(n784),.dout(w_dff_B_bgnk8CN45_0),.clk(gclk));
	jdff dff_B_DiO322YL7_0(.din(w_dff_B_bgnk8CN45_0),.dout(w_dff_B_DiO322YL7_0),.clk(gclk));
	jdff dff_B_QSAAz7sD6_0(.din(w_dff_B_DiO322YL7_0),.dout(w_dff_B_QSAAz7sD6_0),.clk(gclk));
	jdff dff_B_2phjyk4W1_0(.din(w_dff_B_QSAAz7sD6_0),.dout(w_dff_B_2phjyk4W1_0),.clk(gclk));
	jdff dff_B_HKKGKKBb7_0(.din(w_dff_B_2phjyk4W1_0),.dout(w_dff_B_HKKGKKBb7_0),.clk(gclk));
	jdff dff_B_slILIBFh7_0(.din(w_dff_B_HKKGKKBb7_0),.dout(w_dff_B_slILIBFh7_0),.clk(gclk));
	jdff dff_B_GnEZZa5h6_0(.din(w_dff_B_slILIBFh7_0),.dout(w_dff_B_GnEZZa5h6_0),.clk(gclk));
	jdff dff_B_2XRZcm3V8_0(.din(w_dff_B_GnEZZa5h6_0),.dout(w_dff_B_2XRZcm3V8_0),.clk(gclk));
	jdff dff_B_EFk3Y9Tt1_0(.din(w_dff_B_2XRZcm3V8_0),.dout(w_dff_B_EFk3Y9Tt1_0),.clk(gclk));
	jdff dff_B_zseAXeDE6_0(.din(w_dff_B_EFk3Y9Tt1_0),.dout(w_dff_B_zseAXeDE6_0),.clk(gclk));
	jdff dff_B_9IuZgE8F7_0(.din(w_dff_B_zseAXeDE6_0),.dout(w_dff_B_9IuZgE8F7_0),.clk(gclk));
	jdff dff_B_MpSWbReq4_0(.din(w_dff_B_9IuZgE8F7_0),.dout(w_dff_B_MpSWbReq4_0),.clk(gclk));
	jdff dff_B_alibiwfi3_0(.din(w_dff_B_MpSWbReq4_0),.dout(w_dff_B_alibiwfi3_0),.clk(gclk));
	jdff dff_B_L8rAT8m70_0(.din(w_dff_B_alibiwfi3_0),.dout(w_dff_B_L8rAT8m70_0),.clk(gclk));
	jdff dff_B_39uXXub01_0(.din(w_dff_B_L8rAT8m70_0),.dout(w_dff_B_39uXXub01_0),.clk(gclk));
	jdff dff_B_bLDCNedl5_0(.din(w_dff_B_39uXXub01_0),.dout(w_dff_B_bLDCNedl5_0),.clk(gclk));
	jdff dff_B_Q1LIwqe58_0(.din(w_dff_B_bLDCNedl5_0),.dout(w_dff_B_Q1LIwqe58_0),.clk(gclk));
	jdff dff_A_pq1kqkUf9_1(.dout(w_n116_0[1]),.din(w_dff_A_pq1kqkUf9_1),.clk(gclk));
	jdff dff_A_76i7BKoX5_1(.dout(w_dff_A_pq1kqkUf9_1),.din(w_dff_A_76i7BKoX5_1),.clk(gclk));
	jdff dff_B_INXKO3Aj0_0(.din(n780),.dout(w_dff_B_INXKO3Aj0_0),.clk(gclk));
	jdff dff_A_3ErFUkCU3_0(.dout(w_n779_0[0]),.din(w_dff_A_3ErFUkCU3_0),.clk(gclk));
	jdff dff_B_ismogaiY2_1(.din(n774),.dout(w_dff_B_ismogaiY2_1),.clk(gclk));
	jdff dff_A_Tqa4XRTQ6_0(.dout(w_n519_1[0]),.din(w_dff_A_Tqa4XRTQ6_0),.clk(gclk));
	jdff dff_B_1lyPjolQ8_1(.din(n1174),.dout(w_dff_B_1lyPjolQ8_1),.clk(gclk));
	jdff dff_B_STSgn9S99_1(.din(w_dff_B_1lyPjolQ8_1),.dout(w_dff_B_STSgn9S99_1),.clk(gclk));
	jdff dff_B_ksuYp0Ct0_1(.din(w_dff_B_STSgn9S99_1),.dout(w_dff_B_ksuYp0Ct0_1),.clk(gclk));
	jdff dff_B_cUnlXmVH2_1(.din(w_dff_B_ksuYp0Ct0_1),.dout(w_dff_B_cUnlXmVH2_1),.clk(gclk));
	jdff dff_B_7xWKsNru0_1(.din(w_dff_B_cUnlXmVH2_1),.dout(w_dff_B_7xWKsNru0_1),.clk(gclk));
	jdff dff_B_OLwqOrq20_1(.din(w_dff_B_7xWKsNru0_1),.dout(w_dff_B_OLwqOrq20_1),.clk(gclk));
	jdff dff_B_j5kNHohR6_1(.din(w_dff_B_OLwqOrq20_1),.dout(w_dff_B_j5kNHohR6_1),.clk(gclk));
	jdff dff_B_av9rlSH53_1(.din(w_dff_B_j5kNHohR6_1),.dout(w_dff_B_av9rlSH53_1),.clk(gclk));
	jdff dff_B_CQ4RFwI08_1(.din(w_dff_B_av9rlSH53_1),.dout(w_dff_B_CQ4RFwI08_1),.clk(gclk));
	jdff dff_B_EP064UMY9_1(.din(w_dff_B_CQ4RFwI08_1),.dout(w_dff_B_EP064UMY9_1),.clk(gclk));
	jdff dff_B_6wGLHJU34_1(.din(w_dff_B_EP064UMY9_1),.dout(w_dff_B_6wGLHJU34_1),.clk(gclk));
	jdff dff_B_vckcHnIO7_1(.din(w_dff_B_6wGLHJU34_1),.dout(w_dff_B_vckcHnIO7_1),.clk(gclk));
	jdff dff_B_FYYw2jGJ6_1(.din(w_dff_B_vckcHnIO7_1),.dout(w_dff_B_FYYw2jGJ6_1),.clk(gclk));
	jdff dff_B_bIzB3b574_1(.din(w_dff_B_FYYw2jGJ6_1),.dout(w_dff_B_bIzB3b574_1),.clk(gclk));
	jdff dff_B_GYgaBrU91_1(.din(w_dff_B_bIzB3b574_1),.dout(w_dff_B_GYgaBrU91_1),.clk(gclk));
	jdff dff_B_m8yHHaLW0_1(.din(w_dff_B_GYgaBrU91_1),.dout(w_dff_B_m8yHHaLW0_1),.clk(gclk));
	jdff dff_B_9dBhZNRm2_1(.din(w_dff_B_m8yHHaLW0_1),.dout(w_dff_B_9dBhZNRm2_1),.clk(gclk));
	jdff dff_B_ABL8aGuQ4_1(.din(w_dff_B_9dBhZNRm2_1),.dout(w_dff_B_ABL8aGuQ4_1),.clk(gclk));
	jdff dff_B_oD7sEuKY4_1(.din(w_dff_B_ABL8aGuQ4_1),.dout(w_dff_B_oD7sEuKY4_1),.clk(gclk));
	jdff dff_B_0cGMx41z6_1(.din(w_dff_B_oD7sEuKY4_1),.dout(w_dff_B_0cGMx41z6_1),.clk(gclk));
	jdff dff_B_e8nhOBiv9_1(.din(w_dff_B_0cGMx41z6_1),.dout(w_dff_B_e8nhOBiv9_1),.clk(gclk));
	jdff dff_B_7lWRFK0D9_1(.din(w_dff_B_e8nhOBiv9_1),.dout(w_dff_B_7lWRFK0D9_1),.clk(gclk));
	jdff dff_B_M7PXAHRb5_1(.din(w_dff_B_7lWRFK0D9_1),.dout(w_dff_B_M7PXAHRb5_1),.clk(gclk));
	jdff dff_B_PtNcMZnx7_1(.din(w_dff_B_M7PXAHRb5_1),.dout(w_dff_B_PtNcMZnx7_1),.clk(gclk));
	jdff dff_B_fVe4i1GS5_1(.din(w_dff_B_PtNcMZnx7_1),.dout(w_dff_B_fVe4i1GS5_1),.clk(gclk));
	jdff dff_B_Dkas4rHc5_1(.din(w_dff_B_fVe4i1GS5_1),.dout(w_dff_B_Dkas4rHc5_1),.clk(gclk));
	jdff dff_A_1gHWTp1M2_0(.dout(w_n1172_0[0]),.din(w_dff_A_1gHWTp1M2_0),.clk(gclk));
	jdff dff_B_d1iaAPKo4_1(.din(n1166),.dout(w_dff_B_d1iaAPKo4_1),.clk(gclk));
	jdff dff_B_F6HiktET4_1(.din(w_dff_B_d1iaAPKo4_1),.dout(w_dff_B_F6HiktET4_1),.clk(gclk));
	jdff dff_B_Itre6EaQ7_1(.din(n1186),.dout(w_dff_B_Itre6EaQ7_1),.clk(gclk));
	jdff dff_B_WPTFmLO94_1(.din(w_dff_B_Itre6EaQ7_1),.dout(w_dff_B_WPTFmLO94_1),.clk(gclk));
	jdff dff_B_0KnA5P1y8_1(.din(w_dff_B_WPTFmLO94_1),.dout(w_dff_B_0KnA5P1y8_1),.clk(gclk));
	jdff dff_B_qKV9czAu7_1(.din(w_dff_B_0KnA5P1y8_1),.dout(w_dff_B_qKV9czAu7_1),.clk(gclk));
	jdff dff_B_S7POIotw4_1(.din(w_dff_B_qKV9czAu7_1),.dout(w_dff_B_S7POIotw4_1),.clk(gclk));
	jdff dff_B_KGURSiXD8_1(.din(w_dff_B_S7POIotw4_1),.dout(w_dff_B_KGURSiXD8_1),.clk(gclk));
	jdff dff_B_71sAdNul4_1(.din(w_dff_B_KGURSiXD8_1),.dout(w_dff_B_71sAdNul4_1),.clk(gclk));
	jdff dff_B_oMD68yai7_1(.din(w_dff_B_71sAdNul4_1),.dout(w_dff_B_oMD68yai7_1),.clk(gclk));
	jdff dff_B_ow1ivQgc4_1(.din(w_dff_B_oMD68yai7_1),.dout(w_dff_B_ow1ivQgc4_1),.clk(gclk));
	jdff dff_B_Yw4TcDea7_1(.din(w_dff_B_ow1ivQgc4_1),.dout(w_dff_B_Yw4TcDea7_1),.clk(gclk));
	jdff dff_B_xRYm96vM2_1(.din(w_dff_B_Yw4TcDea7_1),.dout(w_dff_B_xRYm96vM2_1),.clk(gclk));
	jdff dff_B_eUB6iv2E4_1(.din(w_dff_B_xRYm96vM2_1),.dout(w_dff_B_eUB6iv2E4_1),.clk(gclk));
	jdff dff_B_cEsRtduB3_1(.din(w_dff_B_eUB6iv2E4_1),.dout(w_dff_B_cEsRtduB3_1),.clk(gclk));
	jdff dff_B_8nXiF0Vw6_1(.din(w_dff_B_cEsRtduB3_1),.dout(w_dff_B_8nXiF0Vw6_1),.clk(gclk));
	jdff dff_B_srSpfLWX5_1(.din(w_dff_B_8nXiF0Vw6_1),.dout(w_dff_B_srSpfLWX5_1),.clk(gclk));
	jdff dff_B_aaCjEMMh1_1(.din(w_dff_B_srSpfLWX5_1),.dout(w_dff_B_aaCjEMMh1_1),.clk(gclk));
	jdff dff_B_3XkVdb4L2_1(.din(w_dff_B_aaCjEMMh1_1),.dout(w_dff_B_3XkVdb4L2_1),.clk(gclk));
	jdff dff_B_haZlQY2K5_1(.din(w_dff_B_3XkVdb4L2_1),.dout(w_dff_B_haZlQY2K5_1),.clk(gclk));
	jdff dff_B_eHtJxHqZ6_1(.din(w_dff_B_haZlQY2K5_1),.dout(w_dff_B_eHtJxHqZ6_1),.clk(gclk));
	jdff dff_B_atyYGVVP2_1(.din(w_dff_B_eHtJxHqZ6_1),.dout(w_dff_B_atyYGVVP2_1),.clk(gclk));
	jdff dff_B_GBCDlgHM7_1(.din(w_dff_B_atyYGVVP2_1),.dout(w_dff_B_GBCDlgHM7_1),.clk(gclk));
	jdff dff_B_PNjCKbEy0_1(.din(w_dff_B_GBCDlgHM7_1),.dout(w_dff_B_PNjCKbEy0_1),.clk(gclk));
	jdff dff_B_nNzt09gq4_1(.din(w_dff_B_PNjCKbEy0_1),.dout(w_dff_B_nNzt09gq4_1),.clk(gclk));
	jdff dff_B_nr9EUWKf8_1(.din(G2897),.dout(w_dff_B_nr9EUWKf8_1),.clk(gclk));
	jdff dff_B_HoUtMLY20_1(.din(w_dff_B_nr9EUWKf8_1),.dout(w_dff_B_HoUtMLY20_1),.clk(gclk));
	jdff dff_B_Tn5Dfvsh7_1(.din(w_dff_B_HoUtMLY20_1),.dout(w_dff_B_Tn5Dfvsh7_1),.clk(gclk));
	jdff dff_A_FkrEWMOn2_0(.dout(w_n1184_0[0]),.din(w_dff_A_FkrEWMOn2_0),.clk(gclk));
	jdff dff_A_i13Nxk1d4_0(.dout(w_dff_A_FkrEWMOn2_0),.din(w_dff_A_i13Nxk1d4_0),.clk(gclk));
	jdff dff_A_wMshBjsY8_0(.dout(w_dff_A_i13Nxk1d4_0),.din(w_dff_A_wMshBjsY8_0),.clk(gclk));
	jdff dff_A_elJ3kVjw5_0(.dout(w_dff_A_wMshBjsY8_0),.din(w_dff_A_elJ3kVjw5_0),.clk(gclk));
	jdff dff_A_LXcfYMdX0_0(.dout(w_dff_A_elJ3kVjw5_0),.din(w_dff_A_LXcfYMdX0_0),.clk(gclk));
	jdff dff_A_0OlSHuzH1_0(.dout(w_dff_A_LXcfYMdX0_0),.din(w_dff_A_0OlSHuzH1_0),.clk(gclk));
	jdff dff_A_8XzyIIqw3_0(.dout(w_dff_A_0OlSHuzH1_0),.din(w_dff_A_8XzyIIqw3_0),.clk(gclk));
	jdff dff_A_7aIAM5uW5_0(.dout(w_dff_A_8XzyIIqw3_0),.din(w_dff_A_7aIAM5uW5_0),.clk(gclk));
	jdff dff_A_JX7QnrZu6_0(.dout(w_dff_A_7aIAM5uW5_0),.din(w_dff_A_JX7QnrZu6_0),.clk(gclk));
	jdff dff_A_YYX4gCcC9_0(.dout(w_dff_A_JX7QnrZu6_0),.din(w_dff_A_YYX4gCcC9_0),.clk(gclk));
	jdff dff_A_ezIhfjT26_0(.dout(w_dff_A_YYX4gCcC9_0),.din(w_dff_A_ezIhfjT26_0),.clk(gclk));
	jdff dff_A_EinBL5jg3_0(.dout(w_dff_A_ezIhfjT26_0),.din(w_dff_A_EinBL5jg3_0),.clk(gclk));
	jdff dff_A_fWezhZQK1_0(.dout(w_dff_A_EinBL5jg3_0),.din(w_dff_A_fWezhZQK1_0),.clk(gclk));
	jdff dff_A_pyHyVM520_0(.dout(w_dff_A_fWezhZQK1_0),.din(w_dff_A_pyHyVM520_0),.clk(gclk));
	jdff dff_A_uTB02lxm3_0(.dout(w_dff_A_pyHyVM520_0),.din(w_dff_A_uTB02lxm3_0),.clk(gclk));
	jdff dff_A_Czfwup3U9_0(.dout(w_dff_A_uTB02lxm3_0),.din(w_dff_A_Czfwup3U9_0),.clk(gclk));
	jdff dff_A_s2qmCIG71_0(.dout(w_dff_A_Czfwup3U9_0),.din(w_dff_A_s2qmCIG71_0),.clk(gclk));
	jdff dff_A_fLRtkNEI5_0(.dout(w_dff_A_s2qmCIG71_0),.din(w_dff_A_fLRtkNEI5_0),.clk(gclk));
	jdff dff_A_QiWqXZtD8_0(.dout(w_dff_A_fLRtkNEI5_0),.din(w_dff_A_QiWqXZtD8_0),.clk(gclk));
	jdff dff_A_hlIfiqL39_0(.dout(w_dff_A_QiWqXZtD8_0),.din(w_dff_A_hlIfiqL39_0),.clk(gclk));
	jdff dff_A_wZ6b6fHU0_0(.dout(w_dff_A_hlIfiqL39_0),.din(w_dff_A_wZ6b6fHU0_0),.clk(gclk));
	jdff dff_A_0WDg3HZv0_0(.dout(w_dff_A_wZ6b6fHU0_0),.din(w_dff_A_0WDg3HZv0_0),.clk(gclk));
	jdff dff_A_ED2r026o9_0(.dout(w_dff_A_0WDg3HZv0_0),.din(w_dff_A_ED2r026o9_0),.clk(gclk));
	jdff dff_A_2gFj4f353_0(.dout(w_dff_A_ED2r026o9_0),.din(w_dff_A_2gFj4f353_0),.clk(gclk));
	jdff dff_A_CUINI1G20_1(.dout(w_n1175_0[1]),.din(w_dff_A_CUINI1G20_1),.clk(gclk));
	jdff dff_A_qG5g4Kdt6_1(.dout(w_dff_A_CUINI1G20_1),.din(w_dff_A_qG5g4Kdt6_1),.clk(gclk));
	jdff dff_A_VKYtCPlx4_1(.dout(w_dff_A_qG5g4Kdt6_1),.din(w_dff_A_VKYtCPlx4_1),.clk(gclk));
	jdff dff_A_KWqK4jsg9_1(.dout(w_dff_A_VKYtCPlx4_1),.din(w_dff_A_KWqK4jsg9_1),.clk(gclk));
	jdff dff_A_fSoq5eSk9_1(.dout(w_dff_A_KWqK4jsg9_1),.din(w_dff_A_fSoq5eSk9_1),.clk(gclk));
	jdff dff_A_2RZGnjge1_1(.dout(w_dff_A_fSoq5eSk9_1),.din(w_dff_A_2RZGnjge1_1),.clk(gclk));
	jdff dff_A_jlR3c4od4_1(.dout(w_dff_A_2RZGnjge1_1),.din(w_dff_A_jlR3c4od4_1),.clk(gclk));
	jdff dff_A_YbRQWkiM0_1(.dout(w_dff_A_jlR3c4od4_1),.din(w_dff_A_YbRQWkiM0_1),.clk(gclk));
	jdff dff_A_LpgbsOwJ3_1(.dout(w_dff_A_YbRQWkiM0_1),.din(w_dff_A_LpgbsOwJ3_1),.clk(gclk));
	jdff dff_A_HkHWyVHQ7_1(.dout(w_dff_A_LpgbsOwJ3_1),.din(w_dff_A_HkHWyVHQ7_1),.clk(gclk));
	jdff dff_A_bPrk78ai6_1(.dout(w_dff_A_HkHWyVHQ7_1),.din(w_dff_A_bPrk78ai6_1),.clk(gclk));
	jdff dff_A_RwyT5Put4_1(.dout(w_dff_A_bPrk78ai6_1),.din(w_dff_A_RwyT5Put4_1),.clk(gclk));
	jdff dff_A_BSkzwkY28_1(.dout(w_dff_A_RwyT5Put4_1),.din(w_dff_A_BSkzwkY28_1),.clk(gclk));
	jdff dff_A_GYfWShQb6_1(.dout(w_dff_A_BSkzwkY28_1),.din(w_dff_A_GYfWShQb6_1),.clk(gclk));
	jdff dff_A_9sO4ZTmB4_1(.dout(w_dff_A_GYfWShQb6_1),.din(w_dff_A_9sO4ZTmB4_1),.clk(gclk));
	jdff dff_A_EAUOJHMP3_1(.dout(w_dff_A_9sO4ZTmB4_1),.din(w_dff_A_EAUOJHMP3_1),.clk(gclk));
	jdff dff_A_hjlqjJGa8_1(.dout(w_dff_A_EAUOJHMP3_1),.din(w_dff_A_hjlqjJGa8_1),.clk(gclk));
	jdff dff_A_WW1YB6Nx9_1(.dout(w_dff_A_hjlqjJGa8_1),.din(w_dff_A_WW1YB6Nx9_1),.clk(gclk));
	jdff dff_A_6kQ4PVCa9_1(.dout(w_dff_A_WW1YB6Nx9_1),.din(w_dff_A_6kQ4PVCa9_1),.clk(gclk));
	jdff dff_A_UnE89SV35_1(.dout(w_dff_A_6kQ4PVCa9_1),.din(w_dff_A_UnE89SV35_1),.clk(gclk));
	jdff dff_A_TwVIFBZk6_1(.dout(w_dff_A_UnE89SV35_1),.din(w_dff_A_TwVIFBZk6_1),.clk(gclk));
	jdff dff_A_BVhJRhXi2_1(.dout(w_dff_A_TwVIFBZk6_1),.din(w_dff_A_BVhJRhXi2_1),.clk(gclk));
	jdff dff_A_2P7m60Fo7_1(.dout(w_dff_A_BVhJRhXi2_1),.din(w_dff_A_2P7m60Fo7_1),.clk(gclk));
	jdff dff_A_TkG7pfVH7_1(.dout(w_dff_A_2P7m60Fo7_1),.din(w_dff_A_TkG7pfVH7_1),.clk(gclk));
	jdff dff_A_PBO6IMgf3_1(.dout(w_dff_A_TkG7pfVH7_1),.din(w_dff_A_PBO6IMgf3_1),.clk(gclk));
	jdff dff_A_75qdFNfU4_0(.dout(w_n1187_0[0]),.din(w_dff_A_75qdFNfU4_0),.clk(gclk));
	jdff dff_B_DVFnj4U50_1(.din(n1060),.dout(w_dff_B_DVFnj4U50_1),.clk(gclk));
	jdff dff_B_kjZczfGZ9_0(.din(n1112),.dout(w_dff_B_kjZczfGZ9_0),.clk(gclk));
	jdff dff_B_z9x0sSSx3_0(.din(w_dff_B_kjZczfGZ9_0),.dout(w_dff_B_z9x0sSSx3_0),.clk(gclk));
	jdff dff_B_mueMJx3S2_0(.din(w_dff_B_z9x0sSSx3_0),.dout(w_dff_B_mueMJx3S2_0),.clk(gclk));
	jdff dff_B_krCILoBk6_0(.din(w_dff_B_mueMJx3S2_0),.dout(w_dff_B_krCILoBk6_0),.clk(gclk));
	jdff dff_B_7VYOSbKx5_0(.din(w_dff_B_krCILoBk6_0),.dout(w_dff_B_7VYOSbKx5_0),.clk(gclk));
	jdff dff_B_H8cVUlWX9_0(.din(w_dff_B_7VYOSbKx5_0),.dout(w_dff_B_H8cVUlWX9_0),.clk(gclk));
	jdff dff_B_KyoqtR4A7_0(.din(n1111),.dout(w_dff_B_KyoqtR4A7_0),.clk(gclk));
	jdff dff_B_92gJze930_0(.din(w_dff_B_KyoqtR4A7_0),.dout(w_dff_B_92gJze930_0),.clk(gclk));
	jdff dff_B_8BSMLYpj6_0(.din(n1110),.dout(w_dff_B_8BSMLYpj6_0),.clk(gclk));
	jdff dff_B_9ILQ2W4v2_0(.din(w_dff_B_8BSMLYpj6_0),.dout(w_dff_B_9ILQ2W4v2_0),.clk(gclk));
	jdff dff_B_S2QAhHBW2_0(.din(w_dff_B_9ILQ2W4v2_0),.dout(w_dff_B_S2QAhHBW2_0),.clk(gclk));
	jdff dff_B_uRmScwGU2_0(.din(w_dff_B_S2QAhHBW2_0),.dout(w_dff_B_uRmScwGU2_0),.clk(gclk));
	jdff dff_B_fS9LehUH7_0(.din(w_dff_B_uRmScwGU2_0),.dout(w_dff_B_fS9LehUH7_0),.clk(gclk));
	jdff dff_B_wBzgC1T75_0(.din(n1109),.dout(w_dff_B_wBzgC1T75_0),.clk(gclk));
	jdff dff_B_ROu9VDUx5_0(.din(w_dff_B_wBzgC1T75_0),.dout(w_dff_B_ROu9VDUx5_0),.clk(gclk));
	jdff dff_B_2cDIwnZe2_1(.din(n1066),.dout(w_dff_B_2cDIwnZe2_1),.clk(gclk));
	jdff dff_B_oF2J7WMc8_1(.din(w_dff_B_2cDIwnZe2_1),.dout(w_dff_B_oF2J7WMc8_1),.clk(gclk));
	jdff dff_B_SsjTCZ8P9_1(.din(w_dff_B_oF2J7WMc8_1),.dout(w_dff_B_SsjTCZ8P9_1),.clk(gclk));
	jdff dff_B_bhAskbXh4_1(.din(w_dff_B_SsjTCZ8P9_1),.dout(w_dff_B_bhAskbXh4_1),.clk(gclk));
	jdff dff_B_BtmoNtxU2_1(.din(w_dff_B_bhAskbXh4_1),.dout(w_dff_B_BtmoNtxU2_1),.clk(gclk));
	jdff dff_B_x9p7lb4a7_1(.din(w_dff_B_BtmoNtxU2_1),.dout(w_dff_B_x9p7lb4a7_1),.clk(gclk));
	jdff dff_B_IP1rCXvj1_1(.din(w_dff_B_x9p7lb4a7_1),.dout(w_dff_B_IP1rCXvj1_1),.clk(gclk));
	jdff dff_B_PeH7jio82_1(.din(w_dff_B_IP1rCXvj1_1),.dout(w_dff_B_PeH7jio82_1),.clk(gclk));
	jdff dff_B_VB52pyBY9_1(.din(n1086),.dout(w_dff_B_VB52pyBY9_1),.clk(gclk));
	jdff dff_B_qrhrT4zO7_0(.din(n1105),.dout(w_dff_B_qrhrT4zO7_0),.clk(gclk));
	jdff dff_B_MQBvZFPF6_0(.din(w_dff_B_qrhrT4zO7_0),.dout(w_dff_B_MQBvZFPF6_0),.clk(gclk));
	jdff dff_B_LIftqJ252_0(.din(w_dff_B_MQBvZFPF6_0),.dout(w_dff_B_LIftqJ252_0),.clk(gclk));
	jdff dff_B_71J1ASuV1_0(.din(w_dff_B_LIftqJ252_0),.dout(w_dff_B_71J1ASuV1_0),.clk(gclk));
	jdff dff_B_wH6kjyXK3_0(.din(w_dff_B_71J1ASuV1_0),.dout(w_dff_B_wH6kjyXK3_0),.clk(gclk));
	jdff dff_B_snN3B2LV6_0(.din(w_dff_B_wH6kjyXK3_0),.dout(w_dff_B_snN3B2LV6_0),.clk(gclk));
	jdff dff_B_LYXjIAr02_0(.din(w_dff_B_snN3B2LV6_0),.dout(w_dff_B_LYXjIAr02_0),.clk(gclk));
	jdff dff_B_7iHYmG9Z8_0(.din(w_dff_B_LYXjIAr02_0),.dout(w_dff_B_7iHYmG9Z8_0),.clk(gclk));
	jdff dff_B_l64JFMp40_1(.din(n1092),.dout(w_dff_B_l64JFMp40_1),.clk(gclk));
	jdff dff_B_gLKpy3Be3_1(.din(n1096),.dout(w_dff_B_gLKpy3Be3_1),.clk(gclk));
	jdff dff_B_NepKsP0S7_1(.din(w_dff_B_gLKpy3Be3_1),.dout(w_dff_B_NepKsP0S7_1),.clk(gclk));
	jdff dff_B_hNlRGnM00_0(.din(n1099),.dout(w_dff_B_hNlRGnM00_0),.clk(gclk));
	jdff dff_B_W0sNcPpq6_0(.din(n1095),.dout(w_dff_B_W0sNcPpq6_0),.clk(gclk));
	jdff dff_B_j0Bgs2dV7_0(.din(w_dff_B_W0sNcPpq6_0),.dout(w_dff_B_j0Bgs2dV7_0),.clk(gclk));
	jdff dff_B_5S8Al6CO4_0(.din(w_dff_B_j0Bgs2dV7_0),.dout(w_dff_B_5S8Al6CO4_0),.clk(gclk));
	jdff dff_B_NtJjTnVt0_1(.din(n1087),.dout(w_dff_B_NtJjTnVt0_1),.clk(gclk));
	jdff dff_B_YsUganJu0_1(.din(w_dff_B_NtJjTnVt0_1),.dout(w_dff_B_YsUganJu0_1),.clk(gclk));
	jdff dff_B_HVAqcWer1_0(.din(n1089),.dout(w_dff_B_HVAqcWer1_0),.clk(gclk));
	jdff dff_B_TFXDdaWy7_1(.din(n1072),.dout(w_dff_B_TFXDdaWy7_1),.clk(gclk));
	jdff dff_B_SFjiaPKT8_1(.din(w_dff_B_TFXDdaWy7_1),.dout(w_dff_B_SFjiaPKT8_1),.clk(gclk));
	jdff dff_B_ggGMsJUX2_1(.din(n1076),.dout(w_dff_B_ggGMsJUX2_1),.clk(gclk));
	jdff dff_B_eJtHe2Jq2_1(.din(G124),.dout(w_dff_B_eJtHe2Jq2_1),.clk(gclk));
	jdff dff_B_10xCu5ic8_1(.din(w_dff_B_eJtHe2Jq2_1),.dout(w_dff_B_10xCu5ic8_1),.clk(gclk));
	jdff dff_B_9YDK52XL0_1(.din(w_dff_B_10xCu5ic8_1),.dout(w_dff_B_9YDK52XL0_1),.clk(gclk));
	jdff dff_B_vnVczlSn4_1(.din(w_dff_B_9YDK52XL0_1),.dout(w_dff_B_vnVczlSn4_1),.clk(gclk));
	jdff dff_B_EG6ARHJv1_1(.din(n1077),.dout(w_dff_B_EG6ARHJv1_1),.clk(gclk));
	jdff dff_B_dYravbQS3_0(.din(n1075),.dout(w_dff_B_dYravbQS3_0),.clk(gclk));
	jdff dff_B_7XdmRs1Y7_0(.din(w_dff_B_dYravbQS3_0),.dout(w_dff_B_7XdmRs1Y7_0),.clk(gclk));
	jdff dff_B_AVUazYlt7_0(.din(w_dff_B_7XdmRs1Y7_0),.dout(w_dff_B_AVUazYlt7_0),.clk(gclk));
	jdff dff_B_dtJPXaif5_0(.din(w_dff_B_AVUazYlt7_0),.dout(w_dff_B_dtJPXaif5_0),.clk(gclk));
	jdff dff_B_9uif3c2I5_1(.din(n1067),.dout(w_dff_B_9uif3c2I5_1),.clk(gclk));
	jdff dff_B_qMUJgFx84_1(.din(n1061),.dout(w_dff_B_qMUJgFx84_1),.clk(gclk));
	jdff dff_B_MqphnD900_1(.din(n1051),.dout(w_dff_B_MqphnD900_1),.clk(gclk));
	jdff dff_B_XlWbM8QL0_1(.din(w_dff_B_MqphnD900_1),.dout(w_dff_B_XlWbM8QL0_1),.clk(gclk));
	jdff dff_B_d1NIOL8X8_1(.din(w_dff_B_XlWbM8QL0_1),.dout(w_dff_B_d1NIOL8X8_1),.clk(gclk));
	jdff dff_A_RZtshrj92_1(.dout(w_n1057_0[1]),.din(w_dff_A_RZtshrj92_1),.clk(gclk));
	jdff dff_A_Xxqvm21W1_1(.dout(w_dff_A_RZtshrj92_1),.din(w_dff_A_Xxqvm21W1_1),.clk(gclk));
	jdff dff_A_j760mmVa3_1(.dout(w_dff_A_Xxqvm21W1_1),.din(w_dff_A_j760mmVa3_1),.clk(gclk));
	jdff dff_A_6aGBmUHX2_1(.dout(w_dff_A_j760mmVa3_1),.din(w_dff_A_6aGBmUHX2_1),.clk(gclk));
	jdff dff_A_gRcrxL502_1(.dout(w_dff_A_6aGBmUHX2_1),.din(w_dff_A_gRcrxL502_1),.clk(gclk));
	jdff dff_A_qQrMKb5R0_0(.dout(w_n1052_0[0]),.din(w_dff_A_qQrMKb5R0_0),.clk(gclk));
	jdff dff_B_1vL66lyp4_1(.din(n753),.dout(w_dff_B_1vL66lyp4_1),.clk(gclk));
	jdff dff_B_C7ktbf3h3_1(.din(w_dff_B_1vL66lyp4_1),.dout(w_dff_B_C7ktbf3h3_1),.clk(gclk));
	jdff dff_B_cRQJmgxW2_1(.din(w_dff_B_C7ktbf3h3_1),.dout(w_dff_B_cRQJmgxW2_1),.clk(gclk));
	jdff dff_B_66AscVry2_1(.din(w_dff_B_cRQJmgxW2_1),.dout(w_dff_B_66AscVry2_1),.clk(gclk));
	jdff dff_B_tqzWkzFC0_1(.din(w_dff_B_66AscVry2_1),.dout(w_dff_B_tqzWkzFC0_1),.clk(gclk));
	jdff dff_B_vGoV2cZb0_1(.din(w_dff_B_tqzWkzFC0_1),.dout(w_dff_B_vGoV2cZb0_1),.clk(gclk));
	jdff dff_A_5Tgp0F3a0_1(.dout(w_n758_1[1]),.din(w_dff_A_5Tgp0F3a0_1),.clk(gclk));
	jdff dff_A_kExtFxnH9_1(.dout(w_dff_A_5Tgp0F3a0_1),.din(w_dff_A_kExtFxnH9_1),.clk(gclk));
	jdff dff_A_XQEGH7Fg5_1(.dout(w_dff_A_kExtFxnH9_1),.din(w_dff_A_XQEGH7Fg5_1),.clk(gclk));
	jdff dff_B_tAnG3rFH9_0(.din(n752),.dout(w_dff_B_tAnG3rFH9_0),.clk(gclk));
	jdff dff_B_ROk0rJVR8_0(.din(w_dff_B_tAnG3rFH9_0),.dout(w_dff_B_ROk0rJVR8_0),.clk(gclk));
	jdff dff_B_sGAdXcQK9_0(.din(w_dff_B_ROk0rJVR8_0),.dout(w_dff_B_sGAdXcQK9_0),.clk(gclk));
	jdff dff_B_u9jzawup9_0(.din(w_dff_B_sGAdXcQK9_0),.dout(w_dff_B_u9jzawup9_0),.clk(gclk));
	jdff dff_B_ttQFE8Zp5_0(.din(w_dff_B_u9jzawup9_0),.dout(w_dff_B_ttQFE8Zp5_0),.clk(gclk));
	jdff dff_B_OFsKvyEN6_0(.din(w_dff_B_ttQFE8Zp5_0),.dout(w_dff_B_OFsKvyEN6_0),.clk(gclk));
	jdff dff_B_lsqKqCwg4_0(.din(w_dff_B_OFsKvyEN6_0),.dout(w_dff_B_lsqKqCwg4_0),.clk(gclk));
	jdff dff_B_Au4qUoU05_0(.din(w_dff_B_lsqKqCwg4_0),.dout(w_dff_B_Au4qUoU05_0),.clk(gclk));
	jdff dff_A_WJXeNyEx8_0(.dout(w_n1049_0[0]),.din(w_dff_A_WJXeNyEx8_0),.clk(gclk));
	jdff dff_A_pbWzgCyS4_0(.dout(w_dff_A_WJXeNyEx8_0),.din(w_dff_A_pbWzgCyS4_0),.clk(gclk));
	jdff dff_A_pSs0Kn2T5_1(.dout(w_n1049_0[1]),.din(w_dff_A_pSs0Kn2T5_1),.clk(gclk));
	jdff dff_A_qpemC9y70_1(.dout(w_dff_A_pSs0Kn2T5_1),.din(w_dff_A_qpemC9y70_1),.clk(gclk));
	jdff dff_B_SWbG8yOW4_0(.din(n1048),.dout(w_dff_B_SWbG8yOW4_0),.clk(gclk));
	jdff dff_B_Nrqi0ynE4_0(.din(n1047),.dout(w_dff_B_Nrqi0ynE4_0),.clk(gclk));
	jdff dff_B_tjgyHJ106_0(.din(n1045),.dout(w_dff_B_tjgyHJ106_0),.clk(gclk));
	jdff dff_B_DjOAi9Nd9_0(.din(w_dff_B_tjgyHJ106_0),.dout(w_dff_B_DjOAi9Nd9_0),.clk(gclk));
	jdff dff_B_QcnaCo5a3_0(.din(w_dff_B_DjOAi9Nd9_0),.dout(w_dff_B_QcnaCo5a3_0),.clk(gclk));
	jdff dff_B_eAU6ZNs84_0(.din(w_dff_B_QcnaCo5a3_0),.dout(w_dff_B_eAU6ZNs84_0),.clk(gclk));
	jdff dff_B_VwXBFnol2_0(.din(w_dff_B_eAU6ZNs84_0),.dout(w_dff_B_VwXBFnol2_0),.clk(gclk));
	jdff dff_B_2ViURvvM0_0(.din(n1044),.dout(w_dff_B_2ViURvvM0_0),.clk(gclk));
	jdff dff_B_v7qJ2qFU7_0(.din(w_dff_B_2ViURvvM0_0),.dout(w_dff_B_v7qJ2qFU7_0),.clk(gclk));
	jdff dff_B_l6gt4ru40_0(.din(n1042),.dout(w_dff_B_l6gt4ru40_0),.clk(gclk));
	jdff dff_B_LwLodLqI6_0(.din(w_dff_B_l6gt4ru40_0),.dout(w_dff_B_LwLodLqI6_0),.clk(gclk));
	jdff dff_B_Af0sdr0X2_1(.din(n1030),.dout(w_dff_B_Af0sdr0X2_1),.clk(gclk));
	jdff dff_B_vXFnbtG86_1(.din(n1032),.dout(w_dff_B_vXFnbtG86_1),.clk(gclk));
	jdff dff_B_TQP1YUm59_1(.din(w_dff_B_vXFnbtG86_1),.dout(w_dff_B_TQP1YUm59_1),.clk(gclk));
	jdff dff_B_RP8VEQR27_1(.din(n1035),.dout(w_dff_B_RP8VEQR27_1),.clk(gclk));
	jdff dff_B_86zZpgHb2_1(.din(n1027),.dout(w_dff_B_86zZpgHb2_1),.clk(gclk));
	jdff dff_B_M3Zz5C7m8_0(.din(n1028),.dout(w_dff_B_M3Zz5C7m8_0),.clk(gclk));
	jdff dff_B_RFjhdhla7_1(.din(n1015),.dout(w_dff_B_RFjhdhla7_1),.clk(gclk));
	jdff dff_B_yGPfwFgA3_1(.din(n1017),.dout(w_dff_B_yGPfwFgA3_1),.clk(gclk));
	jdff dff_B_wFxVZoM59_1(.din(n1020),.dout(w_dff_B_wFxVZoM59_1),.clk(gclk));
	jdff dff_B_0MkERJX76_1(.din(n1021),.dout(w_dff_B_0MkERJX76_1),.clk(gclk));
	jdff dff_B_fUpwtMpE7_1(.din(n1011),.dout(w_dff_B_fUpwtMpE7_1),.clk(gclk));
	jdff dff_B_UOaAKzrk5_0(.din(n1013),.dout(w_dff_B_UOaAKzrk5_0),.clk(gclk));
	jdff dff_A_xsEWv84P2_1(.dout(w_G125_0[1]),.din(w_dff_A_xsEWv84P2_1),.clk(gclk));
	jdff dff_B_HHCElp5e4_2(.din(G125),.dout(w_dff_B_HHCElp5e4_2),.clk(gclk));
	jdff dff_B_G86RNpOp3_2(.din(w_dff_B_HHCElp5e4_2),.dout(w_dff_B_G86RNpOp3_2),.clk(gclk));
	jdff dff_B_p5Pr9xfC7_2(.din(w_dff_B_G86RNpOp3_2),.dout(w_dff_B_p5Pr9xfC7_2),.clk(gclk));
	jdff dff_A_slKm5Ewo6_1(.dout(w_n990_0[1]),.din(w_dff_A_slKm5Ewo6_1),.clk(gclk));
	jdff dff_A_7FpSlnU95_1(.dout(w_dff_A_slKm5Ewo6_1),.din(w_dff_A_7FpSlnU95_1),.clk(gclk));
	jdff dff_A_wMvQFKzl8_0(.dout(w_n758_0[0]),.din(w_dff_A_wMvQFKzl8_0),.clk(gclk));
	jdff dff_A_hOWFdUb55_1(.dout(w_n758_0[1]),.din(w_dff_A_hOWFdUb55_1),.clk(gclk));
	jdff dff_A_MmctwkeV4_1(.dout(w_dff_A_hOWFdUb55_1),.din(w_dff_A_MmctwkeV4_1),.clk(gclk));
	jdff dff_A_qmBZvkLz6_1(.dout(w_dff_A_MmctwkeV4_1),.din(w_dff_A_qmBZvkLz6_1),.clk(gclk));
	jdff dff_A_7ay8bsDi0_0(.dout(w_n754_0[0]),.din(w_dff_A_7ay8bsDi0_0),.clk(gclk));
	jdff dff_B_BXD6qlQV4_0(.din(n768),.dout(w_dff_B_BXD6qlQV4_0),.clk(gclk));
	jdff dff_B_WgF3nB0b5_0(.din(n767),.dout(w_dff_B_WgF3nB0b5_0),.clk(gclk));
	jdff dff_B_gPf7eztG3_0(.din(w_dff_B_WgF3nB0b5_0),.dout(w_dff_B_gPf7eztG3_0),.clk(gclk));
	jdff dff_B_YDYslqhf5_0(.din(w_dff_B_gPf7eztG3_0),.dout(w_dff_B_YDYslqhf5_0),.clk(gclk));
	jdff dff_A_pnr9ZWDy8_2(.dout(w_n764_1[2]),.din(w_dff_A_pnr9ZWDy8_2),.clk(gclk));
	jdff dff_A_FQjyNBXB6_2(.dout(w_dff_A_pnr9ZWDy8_2),.din(w_dff_A_FQjyNBXB6_2),.clk(gclk));
	jdff dff_A_mU4FV3g02_1(.dout(w_n1183_0[1]),.din(w_dff_A_mU4FV3g02_1),.clk(gclk));
	jdff dff_B_3exNftqn2_1(.din(n1179),.dout(w_dff_B_3exNftqn2_1),.clk(gclk));
	jdff dff_B_mMffx1gt7_1(.din(w_dff_B_3exNftqn2_1),.dout(w_dff_B_mMffx1gt7_1),.clk(gclk));
	jdff dff_B_sSNfvP074_1(.din(n1180),.dout(w_dff_B_sSNfvP074_1),.clk(gclk));
	jdff dff_B_V1j9SyVP8_1(.din(w_dff_B_sSNfvP074_1),.dout(w_dff_B_V1j9SyVP8_1),.clk(gclk));
	jdff dff_B_nePEl5Xx0_1(.din(w_dff_B_V1j9SyVP8_1),.dout(w_dff_B_nePEl5Xx0_1),.clk(gclk));
	jdff dff_A_Cy2pFh2x2_0(.dout(w_n988_0[0]),.din(w_dff_A_Cy2pFh2x2_0),.clk(gclk));
	jdff dff_A_fyeVzkVI3_0(.dout(w_dff_A_Cy2pFh2x2_0),.din(w_dff_A_fyeVzkVI3_0),.clk(gclk));
	jdff dff_A_O5BkJj945_1(.dout(w_n988_0[1]),.din(w_dff_A_O5BkJj945_1),.clk(gclk));
	jdff dff_B_Cx17UkaA4_0(.din(n986),.dout(w_dff_B_Cx17UkaA4_0),.clk(gclk));
	jdff dff_B_fRdCpgyv1_0(.din(w_dff_B_Cx17UkaA4_0),.dout(w_dff_B_fRdCpgyv1_0),.clk(gclk));
	jdff dff_B_c6pRVtlX6_0(.din(n984),.dout(w_dff_B_c6pRVtlX6_0),.clk(gclk));
	jdff dff_B_2JuQXva06_0(.din(w_dff_B_c6pRVtlX6_0),.dout(w_dff_B_2JuQXva06_0),.clk(gclk));
	jdff dff_B_n3TuTuIJ8_0(.din(w_dff_B_2JuQXva06_0),.dout(w_dff_B_n3TuTuIJ8_0),.clk(gclk));
	jdff dff_B_aNkwzhXz0_0(.din(w_dff_B_n3TuTuIJ8_0),.dout(w_dff_B_aNkwzhXz0_0),.clk(gclk));
	jdff dff_B_M8nSWbet7_0(.din(n983),.dout(w_dff_B_M8nSWbet7_0),.clk(gclk));
	jdff dff_B_rDa61NF65_0(.din(w_dff_B_M8nSWbet7_0),.dout(w_dff_B_rDa61NF65_0),.clk(gclk));
	jdff dff_B_0avh9kPH0_1(.din(n979),.dout(w_dff_B_0avh9kPH0_1),.clk(gclk));
	jdff dff_B_XvEe2tqO0_1(.din(w_dff_B_0avh9kPH0_1),.dout(w_dff_B_XvEe2tqO0_1),.clk(gclk));
	jdff dff_B_Lb7neYNf5_0(.din(n980),.dout(w_dff_B_Lb7neYNf5_0),.clk(gclk));
	jdff dff_A_jQ6iCYFb7_2(.dout(w_G97_2[2]),.din(w_dff_A_jQ6iCYFb7_2),.clk(gclk));
	jdff dff_B_C5qcIsB09_2(.din(n144),.dout(w_dff_B_C5qcIsB09_2),.clk(gclk));
	jdff dff_B_MvjVfA9W0_1(.din(n142),.dout(w_dff_B_MvjVfA9W0_1),.clk(gclk));
	jdff dff_B_ywj6lkni5_1(.din(n966),.dout(w_dff_B_ywj6lkni5_1),.clk(gclk));
	jdff dff_B_whVeXqgD6_1(.din(n968),.dout(w_dff_B_whVeXqgD6_1),.clk(gclk));
	jdff dff_B_WnjYk9sv3_1(.din(n971),.dout(w_dff_B_WnjYk9sv3_1),.clk(gclk));
	jdff dff_B_q2pNGgEz9_0(.din(n972),.dout(w_dff_B_q2pNGgEz9_0),.clk(gclk));
	jdff dff_A_PQFRbtVo2_0(.dout(w_G143_1[0]),.din(w_dff_A_PQFRbtVo2_0),.clk(gclk));
	jdff dff_A_qQppqKnn2_2(.dout(w_G143_1[2]),.din(w_dff_A_qQppqKnn2_2),.clk(gclk));
	jdff dff_A_hfLMMskf5_1(.dout(w_G33_4[1]),.din(w_dff_A_hfLMMskf5_1),.clk(gclk));
	jdff dff_A_WWK0B2oo7_1(.dout(w_dff_A_hfLMMskf5_1),.din(w_dff_A_WWK0B2oo7_1),.clk(gclk));
	jdff dff_A_FEpwPMUa3_1(.dout(w_dff_A_WWK0B2oo7_1),.din(w_dff_A_FEpwPMUa3_1),.clk(gclk));
	jdff dff_A_sVwYQHnY4_1(.dout(w_dff_A_FEpwPMUa3_1),.din(w_dff_A_sVwYQHnY4_1),.clk(gclk));
	jdff dff_A_mp6aKalC4_2(.dout(w_G33_4[2]),.din(w_dff_A_mp6aKalC4_2),.clk(gclk));
	jdff dff_A_gdXVBH7B5_2(.dout(w_dff_A_mp6aKalC4_2),.din(w_dff_A_gdXVBH7B5_2),.clk(gclk));
	jdff dff_A_acilBIRd4_2(.dout(w_dff_A_gdXVBH7B5_2),.din(w_dff_A_acilBIRd4_2),.clk(gclk));
	jdff dff_A_yjpnAqiE4_2(.dout(w_dff_A_acilBIRd4_2),.din(w_dff_A_yjpnAqiE4_2),.clk(gclk));
	jdff dff_B_QnFifl5M3_0(.din(n964),.dout(w_dff_B_QnFifl5M3_0),.clk(gclk));
	jdff dff_A_snOCCsqR1_1(.dout(w_n962_0[1]),.din(w_dff_A_snOCCsqR1_1),.clk(gclk));
	jdff dff_B_HzyL4HYi9_1(.din(n951),.dout(w_dff_B_HzyL4HYi9_1),.clk(gclk));
	jdff dff_B_OhcYGMIq1_1(.din(n953),.dout(w_dff_B_OhcYGMIq1_1),.clk(gclk));
	jdff dff_B_ByV9zlj97_1(.din(n956),.dout(w_dff_B_ByV9zlj97_1),.clk(gclk));
	jdff dff_B_VJfuxWIR1_0(.din(n957),.dout(w_dff_B_VJfuxWIR1_0),.clk(gclk));
	jdff dff_B_AOeF9rv66_1(.din(n947),.dout(w_dff_B_AOeF9rv66_1),.clk(gclk));
	jdff dff_B_8j7u9TlS3_0(.din(n949),.dout(w_dff_B_8j7u9TlS3_0),.clk(gclk));
	jdff dff_A_lgUsyUaz7_0(.dout(w_n603_1[0]),.din(w_dff_A_lgUsyUaz7_0),.clk(gclk));
	jdff dff_A_Qfqo2AYs7_0(.dout(w_dff_A_lgUsyUaz7_0),.din(w_dff_A_Qfqo2AYs7_0),.clk(gclk));
	jdff dff_A_P4ZigKiT8_0(.dout(w_dff_A_Qfqo2AYs7_0),.din(w_dff_A_P4ZigKiT8_0),.clk(gclk));
	jdff dff_B_FStJrMIY0_1(.din(n850),.dout(w_dff_B_FStJrMIY0_1),.clk(gclk));
	jdff dff_B_NmMHFuky2_1(.din(w_dff_B_FStJrMIY0_1),.dout(w_dff_B_NmMHFuky2_1),.clk(gclk));
	jdff dff_B_sHP7iWLK0_1(.din(w_dff_B_NmMHFuky2_1),.dout(w_dff_B_sHP7iWLK0_1),.clk(gclk));
	jdff dff_B_Un1tSFFn9_1(.din(w_dff_B_sHP7iWLK0_1),.dout(w_dff_B_Un1tSFFn9_1),.clk(gclk));
	jdff dff_B_sdMd6HLu4_1(.din(w_dff_B_Un1tSFFn9_1),.dout(w_dff_B_sdMd6HLu4_1),.clk(gclk));
	jdff dff_B_eRk8zz767_1(.din(w_dff_B_sdMd6HLu4_1),.dout(w_dff_B_eRk8zz767_1),.clk(gclk));
	jdff dff_B_YYMkNhYA5_0(.din(n875),.dout(w_dff_B_YYMkNhYA5_0),.clk(gclk));
	jdff dff_B_roZoaxUK5_0(.din(w_dff_B_YYMkNhYA5_0),.dout(w_dff_B_roZoaxUK5_0),.clk(gclk));
	jdff dff_B_6Fz6g5cU3_1(.din(n871),.dout(w_dff_B_6Fz6g5cU3_1),.clk(gclk));
	jdff dff_B_xvuZQWgj8_1(.din(n868),.dout(w_dff_B_xvuZQWgj8_1),.clk(gclk));
	jdff dff_B_9rSm278z7_1(.din(w_dff_B_xvuZQWgj8_1),.dout(w_dff_B_9rSm278z7_1),.clk(gclk));
	jdff dff_B_Iti47Lbc7_1(.din(w_dff_B_9rSm278z7_1),.dout(w_dff_B_Iti47Lbc7_1),.clk(gclk));
	jdff dff_B_84D6kbgx2_1(.din(w_dff_B_Iti47Lbc7_1),.dout(w_dff_B_84D6kbgx2_1),.clk(gclk));
	jdff dff_B_8swdFZdK9_1(.din(w_dff_B_84D6kbgx2_1),.dout(w_dff_B_8swdFZdK9_1),.clk(gclk));
	jdff dff_A_dgcepEnl3_1(.dout(w_n861_1[1]),.din(w_dff_A_dgcepEnl3_1),.clk(gclk));
	jdff dff_A_RyHrEmPo5_1(.dout(w_dff_A_dgcepEnl3_1),.din(w_dff_A_RyHrEmPo5_1),.clk(gclk));
	jdff dff_A_rwQYYhjr9_2(.dout(w_n861_0[2]),.din(w_dff_A_rwQYYhjr9_2),.clk(gclk));
	jdff dff_A_R0rFJcId8_2(.dout(w_dff_A_rwQYYhjr9_2),.din(w_dff_A_R0rFJcId8_2),.clk(gclk));
	jdff dff_B_2jr7qtF45_0(.din(n860),.dout(w_dff_B_2jr7qtF45_0),.clk(gclk));
	jdff dff_B_ZbbISUN88_0(.din(n857),.dout(w_dff_B_ZbbISUN88_0),.clk(gclk));
	jdff dff_B_Sq1nVs155_0(.din(w_dff_B_ZbbISUN88_0),.dout(w_dff_B_Sq1nVs155_0),.clk(gclk));
	jdff dff_B_WuxO66pk5_0(.din(w_dff_B_Sq1nVs155_0),.dout(w_dff_B_WuxO66pk5_0),.clk(gclk));
	jdff dff_A_vBAbKGaa3_1(.dout(w_n563_0[1]),.din(w_dff_A_vBAbKGaa3_1),.clk(gclk));
	jdff dff_A_phdcRowx4_1(.dout(w_dff_A_vBAbKGaa3_1),.din(w_dff_A_phdcRowx4_1),.clk(gclk));
	jdff dff_A_6IF8HUCr3_2(.dout(w_n563_0[2]),.din(w_dff_A_6IF8HUCr3_2),.clk(gclk));
	jdff dff_A_qh0ueVTK0_2(.dout(w_dff_A_6IF8HUCr3_2),.din(w_dff_A_qh0ueVTK0_2),.clk(gclk));
	jdff dff_B_OEX3IkGW5_1(.din(n555),.dout(w_dff_B_OEX3IkGW5_1),.clk(gclk));
	jdff dff_B_O1xqApWe3_1(.din(w_dff_B_OEX3IkGW5_1),.dout(w_dff_B_O1xqApWe3_1),.clk(gclk));
	jdff dff_B_76bfDyqF7_1(.din(w_dff_B_O1xqApWe3_1),.dout(w_dff_B_76bfDyqF7_1),.clk(gclk));
	jdff dff_B_mxVotttX4_0(.din(n849),.dout(w_dff_B_mxVotttX4_0),.clk(gclk));
	jdff dff_B_vakdpU0h4_0(.din(w_dff_B_mxVotttX4_0),.dout(w_dff_B_vakdpU0h4_0),.clk(gclk));
	jdff dff_B_waiU3iPW9_0(.din(n848),.dout(w_dff_B_waiU3iPW9_0),.clk(gclk));
	jdff dff_B_8GtkNEO43_0(.din(w_dff_B_waiU3iPW9_0),.dout(w_dff_B_8GtkNEO43_0),.clk(gclk));
	jdff dff_B_0dxtSe3b5_0(.din(w_dff_B_8GtkNEO43_0),.dout(w_dff_B_0dxtSe3b5_0),.clk(gclk));
	jdff dff_B_XK9Rr1Md4_0(.din(w_dff_B_0dxtSe3b5_0),.dout(w_dff_B_XK9Rr1Md4_0),.clk(gclk));
	jdff dff_B_HGegVXfg3_1(.din(n844),.dout(w_dff_B_HGegVXfg3_1),.clk(gclk));
	jdff dff_B_EkAG2G5A5_1(.din(w_dff_B_HGegVXfg3_1),.dout(w_dff_B_EkAG2G5A5_1),.clk(gclk));
	jdff dff_B_cNBDWlkf7_0(.din(n845),.dout(w_dff_B_cNBDWlkf7_0),.clk(gclk));
	jdff dff_A_6vLKW1ti3_0(.dout(w_n131_0[0]),.din(w_dff_A_6vLKW1ti3_0),.clk(gclk));
	jdff dff_B_dBwvH5b50_1(.din(n129),.dout(w_dff_B_dBwvH5b50_1),.clk(gclk));
	jdff dff_B_ZsphsNXi2_1(.din(n820),.dout(w_dff_B_ZsphsNXi2_1),.clk(gclk));
	jdff dff_B_9EpyEEZg7_1(.din(w_dff_B_ZsphsNXi2_1),.dout(w_dff_B_9EpyEEZg7_1),.clk(gclk));
	jdff dff_B_tafiDLO83_1(.din(n828),.dout(w_dff_B_tafiDLO83_1),.clk(gclk));
	jdff dff_B_E9q2u0Q57_1(.din(n830),.dout(w_dff_B_E9q2u0Q57_1),.clk(gclk));
	jdff dff_B_l1n21D5a6_1(.din(w_dff_B_E9q2u0Q57_1),.dout(w_dff_B_l1n21D5a6_1),.clk(gclk));
	jdff dff_B_KfVTBMJA0_1(.din(n833),.dout(w_dff_B_KfVTBMJA0_1),.clk(gclk));
	jdff dff_B_GOaq4DFZ9_1(.din(n834),.dout(w_dff_B_GOaq4DFZ9_1),.clk(gclk));
	jdff dff_B_Xkqgtt0R2_1(.din(n822),.dout(w_dff_B_Xkqgtt0R2_1),.clk(gclk));
	jdff dff_B_qpC0aZAa8_1(.din(n809),.dout(w_dff_B_qpC0aZAa8_1),.clk(gclk));
	jdff dff_B_kG1WRgHS8_1(.din(n811),.dout(w_dff_B_kG1WRgHS8_1),.clk(gclk));
	jdff dff_B_TTOk1bak3_1(.din(n814),.dout(w_dff_B_TTOk1bak3_1),.clk(gclk));
	jdff dff_B_LAJJ92v23_1(.din(n815),.dout(w_dff_B_LAJJ92v23_1),.clk(gclk));
	jdff dff_B_liQ1UMAM7_1(.din(n805),.dout(w_dff_B_liQ1UMAM7_1),.clk(gclk));
	jdff dff_B_5f1pzdeI0_0(.din(n807),.dout(w_dff_B_5f1pzdeI0_0),.clk(gclk));
	jdff dff_A_bwpleDz36_2(.dout(w_G107_2[2]),.din(w_dff_A_bwpleDz36_2),.clk(gclk));
	jdff dff_A_TdwTkyIG6_0(.dout(w_n801_0[0]),.din(w_dff_A_TdwTkyIG6_0),.clk(gclk));
	jdff dff_A_eYQCiEqf0_0(.dout(w_dff_A_TdwTkyIG6_0),.din(w_dff_A_eYQCiEqf0_0),.clk(gclk));
	jdff dff_A_LTfKkiCi8_0(.dout(w_dff_A_eYQCiEqf0_0),.din(w_dff_A_LTfKkiCi8_0),.clk(gclk));
	jdff dff_A_4UiU7fNk1_0(.dout(w_dff_A_LTfKkiCi8_0),.din(w_dff_A_4UiU7fNk1_0),.clk(gclk));
	jdff dff_B_N4HDd12h4_0(.din(n800),.dout(w_dff_B_N4HDd12h4_0),.clk(gclk));
	jdff dff_B_O0aVY1Bz7_0(.din(n798),.dout(w_dff_B_O0aVY1Bz7_0),.clk(gclk));
	jdff dff_A_JPVkXb1c2_0(.dout(w_n797_0[0]),.din(w_dff_A_JPVkXb1c2_0),.clk(gclk));
	jdff dff_B_SiD7b9u99_0(.din(n936),.dout(w_dff_B_SiD7b9u99_0),.clk(gclk));
	jdff dff_B_afRYyTAp2_0(.din(w_dff_B_SiD7b9u99_0),.dout(w_dff_B_afRYyTAp2_0),.clk(gclk));
	jdff dff_B_VXjngd2T1_0(.din(n935),.dout(w_dff_B_VXjngd2T1_0),.clk(gclk));
	jdff dff_B_ZNbBFqDO1_0(.din(n934),.dout(w_dff_B_ZNbBFqDO1_0),.clk(gclk));
	jdff dff_B_Nw4q9f9k2_0(.din(w_dff_B_ZNbBFqDO1_0),.dout(w_dff_B_Nw4q9f9k2_0),.clk(gclk));
	jdff dff_B_lUDGU5Tm8_1(.din(n924),.dout(w_dff_B_lUDGU5Tm8_1),.clk(gclk));
	jdff dff_B_l03SnlX31_1(.din(n925),.dout(w_dff_B_l03SnlX31_1),.clk(gclk));
	jdff dff_B_qd4Dr2xX7_1(.din(n916),.dout(w_dff_B_qd4Dr2xX7_1),.clk(gclk));
	jdff dff_B_YfOZGs5a8_1(.din(w_dff_B_qd4Dr2xX7_1),.dout(w_dff_B_YfOZGs5a8_1),.clk(gclk));
	jdff dff_B_1EorlipC6_1(.din(n918),.dout(w_dff_B_1EorlipC6_1),.clk(gclk));
	jdff dff_A_6VDFVZtn3_1(.dout(w_n73_1[1]),.din(w_dff_A_6VDFVZtn3_1),.clk(gclk));
	jdff dff_A_Eux4reDN6_1(.dout(w_n135_0[1]),.din(w_dff_A_Eux4reDN6_1),.clk(gclk));
	jdff dff_B_hpJU5pAe0_1(.din(n133),.dout(w_dff_B_hpJU5pAe0_1),.clk(gclk));
	jdff dff_B_y8ZMZmyl1_1(.din(n902),.dout(w_dff_B_y8ZMZmyl1_1),.clk(gclk));
	jdff dff_B_dTs5iTOn6_1(.din(n904),.dout(w_dff_B_dTs5iTOn6_1),.clk(gclk));
	jdff dff_B_40pmEBcG8_1(.din(n907),.dout(w_dff_B_40pmEBcG8_1),.clk(gclk));
	jdff dff_B_ywfEaQGJ9_1(.din(n908),.dout(w_dff_B_ywfEaQGJ9_1),.clk(gclk));
	jdff dff_A_Atnr6eaZ2_0(.dout(w_G50_2[0]),.din(w_dff_A_Atnr6eaZ2_0),.clk(gclk));
	jdff dff_A_u6lMMEG02_1(.dout(w_G68_2[1]),.din(w_dff_A_u6lMMEG02_1),.clk(gclk));
	jdff dff_A_JEUNizrH2_1(.dout(w_dff_A_u6lMMEG02_1),.din(w_dff_A_JEUNizrH2_1),.clk(gclk));
	jdff dff_A_uiOC0J294_1(.dout(w_dff_A_JEUNizrH2_1),.din(w_dff_A_uiOC0J294_1),.clk(gclk));
	jdff dff_A_f2WoVYay3_2(.dout(w_G68_2[2]),.din(w_dff_A_f2WoVYay3_2),.clk(gclk));
	jdff dff_A_4ndtRwkk5_2(.dout(w_dff_A_f2WoVYay3_2),.din(w_dff_A_4ndtRwkk5_2),.clk(gclk));
	jdff dff_A_YzKwCjno0_2(.dout(w_dff_A_4ndtRwkk5_2),.din(w_dff_A_YzKwCjno0_2),.clk(gclk));
	jdff dff_A_6KVDIPDC3_2(.dout(w_dff_A_YzKwCjno0_2),.din(w_dff_A_6KVDIPDC3_2),.clk(gclk));
	jdff dff_A_UaieZtxF1_1(.dout(w_G150_2[1]),.din(w_dff_A_UaieZtxF1_1),.clk(gclk));
	jdff dff_B_fkrlfE7F9_0(.din(n900),.dout(w_dff_B_fkrlfE7F9_0),.clk(gclk));
	jdff dff_A_rBK6NEAD6_0(.dout(w_G58_2[0]),.din(w_dff_A_rBK6NEAD6_0),.clk(gclk));
	jdff dff_A_n8CIkRW42_0(.dout(w_dff_A_rBK6NEAD6_0),.din(w_dff_A_n8CIkRW42_0),.clk(gclk));
	jdff dff_A_05j5Fhvw0_2(.dout(w_G58_2[2]),.din(w_dff_A_05j5Fhvw0_2),.clk(gclk));
	jdff dff_A_JtTPq6K41_2(.dout(w_dff_A_05j5Fhvw0_2),.din(w_dff_A_JtTPq6K41_2),.clk(gclk));
	jdff dff_B_s3dYIOLe0_1(.din(n887),.dout(w_dff_B_s3dYIOLe0_1),.clk(gclk));
	jdff dff_B_t8HqBvIk0_1(.din(n889),.dout(w_dff_B_t8HqBvIk0_1),.clk(gclk));
	jdff dff_B_ijOsRv3d3_0(.din(n895),.dout(w_dff_B_ijOsRv3d3_0),.clk(gclk));
	jdff dff_B_oAB1G1BA4_0(.din(n891),.dout(w_dff_B_oAB1G1BA4_0),.clk(gclk));
	jdff dff_A_nFcxiCu25_1(.dout(w_G116_2[1]),.din(w_dff_A_nFcxiCu25_1),.clk(gclk));
	jdff dff_A_Ig1MTnX10_2(.dout(w_G116_2[2]),.din(w_dff_A_Ig1MTnX10_2),.clk(gclk));
	jdff dff_B_C8F25GoX1_1(.din(n883),.dout(w_dff_B_C8F25GoX1_1),.clk(gclk));
	jdff dff_B_ArWb2Guz8_0(.din(n885),.dout(w_dff_B_ArWb2Guz8_0),.clk(gclk));
	jdff dff_A_KSVncrO02_0(.dout(w_G283_2[0]),.din(w_dff_A_KSVncrO02_0),.clk(gclk));
	jdff dff_A_cOYiOvKk8_1(.dout(w_G283_2[1]),.din(w_dff_A_cOYiOvKk8_1),.clk(gclk));
	jdff dff_A_XSZpSyWq1_1(.dout(w_n564_0[1]),.din(w_dff_A_XSZpSyWq1_1),.clk(gclk));
	jdff dff_B_GWUvgwss7_1(.din(n878),.dout(w_dff_B_GWUvgwss7_1),.clk(gclk));
	jdff dff_B_CQS8NZev0_1(.din(w_dff_B_GWUvgwss7_1),.dout(w_dff_B_CQS8NZev0_1),.clk(gclk));
	jdff dff_A_TtFrPdwf5_0(.dout(w_n589_1[0]),.din(w_dff_A_TtFrPdwf5_0),.clk(gclk));
	jdff dff_A_4OJKC0OR5_0(.dout(w_dff_A_TtFrPdwf5_0),.din(w_dff_A_4OJKC0OR5_0),.clk(gclk));
	jdff dff_A_0YiUR0Ss4_0(.dout(w_dff_A_4OJKC0OR5_0),.din(w_dff_A_0YiUR0Ss4_0),.clk(gclk));
	jdff dff_A_PXFsuTRE2_0(.dout(w_n592_1[0]),.din(w_dff_A_PXFsuTRE2_0),.clk(gclk));
	jdff dff_A_8VaEDlcY7_0(.dout(w_dff_A_PXFsuTRE2_0),.din(w_dff_A_8VaEDlcY7_0),.clk(gclk));
	jdff dff_A_Iq24XGYr3_1(.dout(w_n592_1[1]),.din(w_dff_A_Iq24XGYr3_1),.clk(gclk));
	jdff dff_B_SYCE2BTn7_0(.din(n852),.dout(w_dff_B_SYCE2BTn7_0),.clk(gclk));
	jdff dff_B_IQmQYXWB0_0(.din(n560),.dout(w_dff_B_IQmQYXWB0_0),.clk(gclk));
	jdff dff_B_q1yVKbPA9_2(.din(n556),.dout(w_dff_B_q1yVKbPA9_2),.clk(gclk));
	jdff dff_B_6XuEDFwA5_2(.din(w_dff_B_q1yVKbPA9_2),.dout(w_dff_B_6XuEDFwA5_2),.clk(gclk));
	jdff dff_A_lRlMu4sD7_0(.dout(w_G396_0[0]),.din(w_dff_A_lRlMu4sD7_0),.clk(gclk));
	jdff dff_A_M0tghYyO0_0(.dout(w_dff_A_lRlMu4sD7_0),.din(w_dff_A_M0tghYyO0_0),.clk(gclk));
	jdff dff_A_i1S5ziKV7_0(.dout(w_dff_A_M0tghYyO0_0),.din(w_dff_A_i1S5ziKV7_0),.clk(gclk));
	jdff dff_B_Ks7agVIe9_0(.din(n687),.dout(w_dff_B_Ks7agVIe9_0),.clk(gclk));
	jdff dff_B_pbid71fM7_0(.din(w_dff_B_Ks7agVIe9_0),.dout(w_dff_B_pbid71fM7_0),.clk(gclk));
	jdff dff_B_t2vIVQ5S6_0(.din(n686),.dout(w_dff_B_t2vIVQ5S6_0),.clk(gclk));
	jdff dff_B_ijCClu5V1_0(.din(w_dff_B_t2vIVQ5S6_0),.dout(w_dff_B_ijCClu5V1_0),.clk(gclk));
	jdff dff_B_TgwTAz0T8_1(.din(n678),.dout(w_dff_B_TgwTAz0T8_1),.clk(gclk));
	jdff dff_B_PrSaw47k1_1(.din(n679),.dout(w_dff_B_PrSaw47k1_1),.clk(gclk));
	jdff dff_B_wnaAccVc0_2(.din(n680),.dout(w_dff_B_wnaAccVc0_2),.clk(gclk));
	jdff dff_B_tSC1lAtp1_1(.din(n673),.dout(w_dff_B_tSC1lAtp1_1),.clk(gclk));
	jdff dff_B_q8O96NZW0_1(.din(w_dff_B_tSC1lAtp1_1),.dout(w_dff_B_q8O96NZW0_1),.clk(gclk));
	jdff dff_B_aPhNAm609_0(.din(n139),.dout(w_dff_B_aPhNAm609_0),.clk(gclk));
	jdff dff_A_Hu6cMehe4_1(.dout(w_n672_1[1]),.din(w_dff_A_Hu6cMehe4_1),.clk(gclk));
	jdff dff_A_lbvI5AZX7_1(.dout(w_dff_A_Hu6cMehe4_1),.din(w_dff_A_lbvI5AZX7_1),.clk(gclk));
	jdff dff_A_7SeFFzao1_1(.dout(w_dff_A_lbvI5AZX7_1),.din(w_dff_A_7SeFFzao1_1),.clk(gclk));
	jdff dff_A_DMFkWSl72_2(.dout(w_n672_0[2]),.din(w_dff_A_DMFkWSl72_2),.clk(gclk));
	jdff dff_A_ndWtT0954_2(.dout(w_dff_A_DMFkWSl72_2),.din(w_dff_A_ndWtT0954_2),.clk(gclk));
	jdff dff_A_s4K4jVzF7_2(.dout(w_dff_A_ndWtT0954_2),.din(w_dff_A_s4K4jVzF7_2),.clk(gclk));
	jdff dff_B_WR5Qgovz9_1(.din(n647),.dout(w_dff_B_WR5Qgovz9_1),.clk(gclk));
	jdff dff_B_SollERH45_1(.din(w_dff_B_WR5Qgovz9_1),.dout(w_dff_B_SollERH45_1),.clk(gclk));
	jdff dff_B_DUUwAbIW3_1(.din(n653),.dout(w_dff_B_DUUwAbIW3_1),.clk(gclk));
	jdff dff_B_JOmrejZn1_1(.din(w_dff_B_DUUwAbIW3_1),.dout(w_dff_B_JOmrejZn1_1),.clk(gclk));
	jdff dff_B_NFw4p7kh4_1(.din(n656),.dout(w_dff_B_NFw4p7kh4_1),.clk(gclk));
	jdff dff_B_cnEI5OKQ2_1(.din(n660),.dout(w_dff_B_cnEI5OKQ2_1),.clk(gclk));
	jdff dff_B_fNJBprkP0_0(.din(n658),.dout(w_dff_B_fNJBprkP0_0),.clk(gclk));
	jdff dff_B_zytjr5lS4_1(.din(n630),.dout(w_dff_B_zytjr5lS4_1),.clk(gclk));
	jdff dff_B_YeRo1S9M1_1(.din(n633),.dout(w_dff_B_YeRo1S9M1_1),.clk(gclk));
	jdff dff_B_xbbZLR3d2_0(.din(n644),.dout(w_dff_B_xbbZLR3d2_0),.clk(gclk));
	jdff dff_A_WorGWE6A7_0(.dout(w_G317_1[0]),.din(w_dff_A_WorGWE6A7_0),.clk(gclk));
	jdff dff_B_A1KkwWH95_3(.din(G317),.dout(w_dff_B_A1KkwWH95_3),.clk(gclk));
	jdff dff_B_3ApFXNkh1_3(.din(w_dff_B_A1KkwWH95_3),.dout(w_dff_B_3ApFXNkh1_3),.clk(gclk));
	jdff dff_B_shLEtSI70_3(.din(w_dff_B_3ApFXNkh1_3),.dout(w_dff_B_shLEtSI70_3),.clk(gclk));
	jdff dff_A_U500Ob7a2_0(.dout(w_G326_0[0]),.din(w_dff_A_U500Ob7a2_0),.clk(gclk));
	jdff dff_B_8nMucfrd1_2(.din(G326),.dout(w_dff_B_8nMucfrd1_2),.clk(gclk));
	jdff dff_B_GGu0UJGT6_2(.din(w_dff_B_8nMucfrd1_2),.dout(w_dff_B_GGu0UJGT6_2),.clk(gclk));
	jdff dff_B_uJt7CJLp2_2(.din(w_dff_B_GGu0UJGT6_2),.dout(w_dff_B_uJt7CJLp2_2),.clk(gclk));
	jdff dff_B_HZGkihJZ2_0(.din(n637),.dout(w_dff_B_HZGkihJZ2_0),.clk(gclk));
	jdff dff_B_gx73yGy73_1(.din(G329),.dout(w_dff_B_gx73yGy73_1),.clk(gclk));
	jdff dff_B_HFEHj2gJ7_1(.din(w_dff_B_gx73yGy73_1),.dout(w_dff_B_HFEHj2gJ7_1),.clk(gclk));
	jdff dff_B_ovBAT9NH3_1(.din(w_dff_B_HFEHj2gJ7_1),.dout(w_dff_B_ovBAT9NH3_1),.clk(gclk));
	jdff dff_B_g3sqqxTD0_1(.din(w_dff_B_ovBAT9NH3_1),.dout(w_dff_B_g3sqqxTD0_1),.clk(gclk));
	jdff dff_A_zvJHdfOq5_1(.dout(w_n148_5[1]),.din(w_dff_A_zvJHdfOq5_1),.clk(gclk));
	jdff dff_A_9QZE4nlL5_1(.dout(w_dff_A_zvJHdfOq5_1),.din(w_dff_A_9QZE4nlL5_1),.clk(gclk));
	jdff dff_A_Z4ls5wLR7_1(.dout(w_dff_A_9QZE4nlL5_1),.din(w_dff_A_Z4ls5wLR7_1),.clk(gclk));
	jdff dff_A_dJDGDyOs2_2(.dout(w_n148_5[2]),.din(w_dff_A_dJDGDyOs2_2),.clk(gclk));
	jdff dff_A_TLWREQpl6_2(.dout(w_dff_A_dJDGDyOs2_2),.din(w_dff_A_TLWREQpl6_2),.clk(gclk));
	jdff dff_B_vPKyQSuR3_1(.din(n618),.dout(w_dff_B_vPKyQSuR3_1),.clk(gclk));
	jdff dff_B_luZy6lJH8_0(.din(n628),.dout(w_dff_B_luZy6lJH8_0),.clk(gclk));
	jdff dff_A_2rrUxUIP9_0(.dout(w_G322_0[0]),.din(w_dff_A_2rrUxUIP9_0),.clk(gclk));
	jdff dff_B_u0neskAZ0_3(.din(G322),.dout(w_dff_B_u0neskAZ0_3),.clk(gclk));
	jdff dff_B_bUL5dkCT3_3(.din(w_dff_B_u0neskAZ0_3),.dout(w_dff_B_bUL5dkCT3_3),.clk(gclk));
	jdff dff_B_cWNoaYa40_3(.din(w_dff_B_bUL5dkCT3_3),.dout(w_dff_B_cWNoaYa40_3),.clk(gclk));
	jdff dff_A_zP6meR3B7_1(.dout(w_n612_4[1]),.din(w_dff_A_zP6meR3B7_1),.clk(gclk));
	jdff dff_A_SvGabuyZ0_1(.dout(w_dff_A_zP6meR3B7_1),.din(w_dff_A_SvGabuyZ0_1),.clk(gclk));
	jdff dff_A_v4aMslTG5_1(.dout(w_dff_A_SvGabuyZ0_1),.din(w_dff_A_v4aMslTG5_1),.clk(gclk));
	jdff dff_A_mEvHV7Qt0_1(.dout(w_dff_A_v4aMslTG5_1),.din(w_dff_A_mEvHV7Qt0_1),.clk(gclk));
	jdff dff_A_fO1gaAU48_1(.dout(w_dff_A_mEvHV7Qt0_1),.din(w_dff_A_fO1gaAU48_1),.clk(gclk));
	jdff dff_A_pq2AYniU8_1(.dout(w_dff_A_fO1gaAU48_1),.din(w_dff_A_pq2AYniU8_1),.clk(gclk));
	jdff dff_A_tmTvCkbU6_1(.dout(w_dff_A_pq2AYniU8_1),.din(w_dff_A_tmTvCkbU6_1),.clk(gclk));
	jdff dff_A_fKgJXFjY1_1(.dout(w_dff_A_tmTvCkbU6_1),.din(w_dff_A_fKgJXFjY1_1),.clk(gclk));
	jdff dff_A_YCzhrQoY5_0(.dout(w_n608_1[0]),.din(w_dff_A_YCzhrQoY5_0),.clk(gclk));
	jdff dff_A_oHrPOyqK9_0(.dout(w_dff_A_YCzhrQoY5_0),.din(w_dff_A_oHrPOyqK9_0),.clk(gclk));
	jdff dff_A_D8WSjl5f6_0(.dout(w_dff_A_oHrPOyqK9_0),.din(w_dff_A_D8WSjl5f6_0),.clk(gclk));
	jdff dff_A_Pp5xVGwQ0_0(.dout(w_dff_A_D8WSjl5f6_0),.din(w_dff_A_Pp5xVGwQ0_0),.clk(gclk));
	jdff dff_A_SCHK0TrY7_0(.dout(w_dff_A_Pp5xVGwQ0_0),.din(w_dff_A_SCHK0TrY7_0),.clk(gclk));
	jdff dff_A_DEZNKbo81_0(.dout(w_dff_A_SCHK0TrY7_0),.din(w_dff_A_DEZNKbo81_0),.clk(gclk));
	jdff dff_A_nBl04f0e9_0(.dout(w_dff_A_DEZNKbo81_0),.din(w_dff_A_nBl04f0e9_0),.clk(gclk));
	jdff dff_A_B0I6oQeg1_0(.dout(w_dff_A_nBl04f0e9_0),.din(w_dff_A_B0I6oQeg1_0),.clk(gclk));
	jdff dff_A_w0rZFdYh7_0(.dout(w_dff_A_B0I6oQeg1_0),.din(w_dff_A_w0rZFdYh7_0),.clk(gclk));
	jdff dff_A_mLqKf1by0_0(.dout(w_dff_A_w0rZFdYh7_0),.din(w_dff_A_mLqKf1by0_0),.clk(gclk));
	jdff dff_A_TGBdpbH83_0(.dout(w_dff_A_mLqKf1by0_0),.din(w_dff_A_TGBdpbH83_0),.clk(gclk));
	jdff dff_A_OSUnoYmz9_2(.dout(w_n608_1[2]),.din(w_dff_A_OSUnoYmz9_2),.clk(gclk));
	jdff dff_A_dtUhY7JZ5_2(.dout(w_dff_A_OSUnoYmz9_2),.din(w_dff_A_dtUhY7JZ5_2),.clk(gclk));
	jdff dff_A_tVr9P22h8_2(.dout(w_dff_A_dtUhY7JZ5_2),.din(w_dff_A_tVr9P22h8_2),.clk(gclk));
	jdff dff_A_6vPwiSX80_2(.dout(w_dff_A_tVr9P22h8_2),.din(w_dff_A_6vPwiSX80_2),.clk(gclk));
	jdff dff_A_iRk3bfpv5_2(.dout(w_dff_A_6vPwiSX80_2),.din(w_dff_A_iRk3bfpv5_2),.clk(gclk));
	jdff dff_A_hO7d4Kf21_2(.dout(w_dff_A_iRk3bfpv5_2),.din(w_dff_A_hO7d4Kf21_2),.clk(gclk));
	jdff dff_A_gqzlGGGV6_2(.dout(w_dff_A_hO7d4Kf21_2),.din(w_dff_A_gqzlGGGV6_2),.clk(gclk));
	jdff dff_A_yKOyCE6l8_2(.dout(w_dff_A_gqzlGGGV6_2),.din(w_dff_A_yKOyCE6l8_2),.clk(gclk));
	jdff dff_A_zOV6tKue4_2(.dout(w_dff_A_yKOyCE6l8_2),.din(w_dff_A_zOV6tKue4_2),.clk(gclk));
	jdff dff_A_duMeiHOw2_2(.dout(w_dff_A_zOV6tKue4_2),.din(w_dff_A_duMeiHOw2_2),.clk(gclk));
	jdff dff_A_VPwrvW8B8_2(.dout(w_dff_A_duMeiHOw2_2),.din(w_dff_A_VPwrvW8B8_2),.clk(gclk));
	jdff dff_A_hmxa8FcC1_1(.dout(w_n608_0[1]),.din(w_dff_A_hmxa8FcC1_1),.clk(gclk));
	jdff dff_A_vuWhESbr7_1(.dout(w_dff_A_hmxa8FcC1_1),.din(w_dff_A_vuWhESbr7_1),.clk(gclk));
	jdff dff_A_9ANYxGzJ0_1(.dout(w_dff_A_vuWhESbr7_1),.din(w_dff_A_9ANYxGzJ0_1),.clk(gclk));
	jdff dff_A_4tFhnOGS8_1(.dout(w_dff_A_9ANYxGzJ0_1),.din(w_dff_A_4tFhnOGS8_1),.clk(gclk));
	jdff dff_A_83D1z8j85_1(.dout(w_dff_A_4tFhnOGS8_1),.din(w_dff_A_83D1z8j85_1),.clk(gclk));
	jdff dff_A_qUKP8lz83_1(.dout(w_dff_A_83D1z8j85_1),.din(w_dff_A_qUKP8lz83_1),.clk(gclk));
	jdff dff_A_DmbFSuqA3_1(.dout(w_dff_A_qUKP8lz83_1),.din(w_dff_A_DmbFSuqA3_1),.clk(gclk));
	jdff dff_A_cZg4qVCH0_1(.dout(w_dff_A_DmbFSuqA3_1),.din(w_dff_A_cZg4qVCH0_1),.clk(gclk));
	jdff dff_A_Bgh0kV3x6_1(.dout(w_dff_A_cZg4qVCH0_1),.din(w_dff_A_Bgh0kV3x6_1),.clk(gclk));
	jdff dff_A_Gs6Q1S7n4_1(.dout(w_dff_A_Bgh0kV3x6_1),.din(w_dff_A_Gs6Q1S7n4_1),.clk(gclk));
	jdff dff_A_NoSDn8eT1_1(.dout(w_dff_A_Gs6Q1S7n4_1),.din(w_dff_A_NoSDn8eT1_1),.clk(gclk));
	jdff dff_A_C14hPYGJ7_2(.dout(w_n608_0[2]),.din(w_dff_A_C14hPYGJ7_2),.clk(gclk));
	jdff dff_A_z19pZXV52_2(.dout(w_dff_A_C14hPYGJ7_2),.din(w_dff_A_z19pZXV52_2),.clk(gclk));
	jdff dff_A_hAhtHYXq4_2(.dout(w_dff_A_z19pZXV52_2),.din(w_dff_A_hAhtHYXq4_2),.clk(gclk));
	jdff dff_A_un2wKVAb1_2(.dout(w_dff_A_hAhtHYXq4_2),.din(w_dff_A_un2wKVAb1_2),.clk(gclk));
	jdff dff_A_ym5MLrHo3_2(.dout(w_dff_A_un2wKVAb1_2),.din(w_dff_A_ym5MLrHo3_2),.clk(gclk));
	jdff dff_A_38imtwwk0_2(.dout(w_dff_A_ym5MLrHo3_2),.din(w_dff_A_38imtwwk0_2),.clk(gclk));
	jdff dff_A_sCNAwjks1_2(.dout(w_dff_A_38imtwwk0_2),.din(w_dff_A_sCNAwjks1_2),.clk(gclk));
	jdff dff_A_yXDZaVji8_2(.dout(w_dff_A_sCNAwjks1_2),.din(w_dff_A_yXDZaVji8_2),.clk(gclk));
	jdff dff_A_gzFbaoh53_2(.dout(w_dff_A_yXDZaVji8_2),.din(w_dff_A_gzFbaoh53_2),.clk(gclk));
	jdff dff_A_8VT3rPAv2_2(.dout(w_dff_A_gzFbaoh53_2),.din(w_dff_A_8VT3rPAv2_2),.clk(gclk));
	jdff dff_A_BxA3UUOd6_2(.dout(w_dff_A_8VT3rPAv2_2),.din(w_dff_A_BxA3UUOd6_2),.clk(gclk));
	jdff dff_B_5JTB6iA73_0(.din(n570),.dout(w_dff_B_5JTB6iA73_0),.clk(gclk));
	jdff dff_B_7Q94a7311_0(.din(w_dff_B_5JTB6iA73_0),.dout(w_dff_B_7Q94a7311_0),.clk(gclk));
	jdff dff_B_ppoLYKA67_0(.din(n568),.dout(w_dff_B_ppoLYKA67_0),.clk(gclk));
	jdff dff_B_jMsEwQnn4_0(.din(w_dff_B_ppoLYKA67_0),.dout(w_dff_B_jMsEwQnn4_0),.clk(gclk));
	jdff dff_B_15lHvnoi4_0(.din(w_dff_B_jMsEwQnn4_0),.dout(w_dff_B_15lHvnoi4_0),.clk(gclk));
	jdff dff_A_Z6UpHq8j9_0(.dout(w_n567_0[0]),.din(w_dff_A_Z6UpHq8j9_0),.clk(gclk));
	jdff dff_A_cJa5wY6U9_0(.dout(w_dff_A_Z6UpHq8j9_0),.din(w_dff_A_cJa5wY6U9_0),.clk(gclk));
	jdff dff_A_zxUPhaMp4_1(.dout(w_n554_3[1]),.din(w_dff_A_zxUPhaMp4_1),.clk(gclk));
	jdff dff_A_kgYENZ1Q6_1(.dout(w_dff_A_zxUPhaMp4_1),.din(w_dff_A_kgYENZ1Q6_1),.clk(gclk));
	jdff dff_A_TXHv3qj30_1(.dout(w_dff_A_kgYENZ1Q6_1),.din(w_dff_A_TXHv3qj30_1),.clk(gclk));
	jdff dff_A_mqDiXdHA4_2(.dout(w_n554_3[2]),.din(w_dff_A_mqDiXdHA4_2),.clk(gclk));
	jdff dff_A_bzLkRZRK6_2(.dout(w_dff_A_mqDiXdHA4_2),.din(w_dff_A_bzLkRZRK6_2),.clk(gclk));
	jdff dff_A_YFww9s9J9_2(.dout(w_dff_A_bzLkRZRK6_2),.din(w_dff_A_YFww9s9J9_2),.clk(gclk));
	jdff dff_B_nX47N2lT6_2(.din(n565),.dout(w_dff_B_nX47N2lT6_2),.clk(gclk));
	jdff dff_B_14nPjPx62_2(.din(w_dff_B_nX47N2lT6_2),.dout(w_dff_B_14nPjPx62_2),.clk(gclk));
	jdff dff_B_DL4bW3ni6_2(.din(w_dff_B_14nPjPx62_2),.dout(w_dff_B_DL4bW3ni6_2),.clk(gclk));
	jdff dff_B_MAKAai9F3_2(.din(w_dff_B_DL4bW3ni6_2),.dout(w_dff_B_MAKAai9F3_2),.clk(gclk));
	jdff dff_B_czCQDN6x0_2(.din(w_dff_B_MAKAai9F3_2),.dout(w_dff_B_czCQDN6x0_2),.clk(gclk));
	jdff dff_B_RNkarPww9_2(.din(w_dff_B_czCQDN6x0_2),.dout(w_dff_B_RNkarPww9_2),.clk(gclk));
	jdff dff_B_habat80T5_2(.din(w_dff_B_RNkarPww9_2),.dout(w_dff_B_habat80T5_2),.clk(gclk));
	jdff dff_B_KsGKK0G76_2(.din(w_dff_B_habat80T5_2),.dout(w_dff_B_KsGKK0G76_2),.clk(gclk));
	jdff dff_B_ZSSh2JVA7_2(.din(w_dff_B_KsGKK0G76_2),.dout(w_dff_B_ZSSh2JVA7_2),.clk(gclk));
	jdff dff_B_VDRNsdvG6_2(.din(w_dff_B_ZSSh2JVA7_2),.dout(w_dff_B_VDRNsdvG6_2),.clk(gclk));
	jdff dff_B_AdqVhlJ89_2(.din(w_dff_B_VDRNsdvG6_2),.dout(w_dff_B_AdqVhlJ89_2),.clk(gclk));
	jdff dff_B_WXIz7OC84_2(.din(w_dff_B_AdqVhlJ89_2),.dout(w_dff_B_WXIz7OC84_2),.clk(gclk));
	jdff dff_B_9D8UaAZR2_2(.din(w_dff_B_WXIz7OC84_2),.dout(w_dff_B_9D8UaAZR2_2),.clk(gclk));
	jdff dff_A_5O7iKcwa2_1(.dout(w_n1162_0[1]),.din(w_dff_A_5O7iKcwa2_1),.clk(gclk));
	jdff dff_B_ozhs6JXt9_0(.din(n1161),.dout(w_dff_B_ozhs6JXt9_0),.clk(gclk));
	jdff dff_B_CJNgHhWI8_0(.din(w_dff_B_ozhs6JXt9_0),.dout(w_dff_B_CJNgHhWI8_0),.clk(gclk));
	jdff dff_B_hsTIU0Cm3_0(.din(n1158),.dout(w_dff_B_hsTIU0Cm3_0),.clk(gclk));
	jdff dff_B_szGITtq51_0(.din(w_dff_B_hsTIU0Cm3_0),.dout(w_dff_B_szGITtq51_0),.clk(gclk));
	jdff dff_B_yb2WQYBS8_0(.din(w_dff_B_szGITtq51_0),.dout(w_dff_B_yb2WQYBS8_0),.clk(gclk));
	jdff dff_B_J0Qggegj6_0(.din(w_dff_B_yb2WQYBS8_0),.dout(w_dff_B_J0Qggegj6_0),.clk(gclk));
	jdff dff_B_kl4sFjwJ4_0(.din(w_dff_B_J0Qggegj6_0),.dout(w_dff_B_kl4sFjwJ4_0),.clk(gclk));
	jdff dff_B_Vkys7uUa8_0(.din(n1157),.dout(w_dff_B_Vkys7uUa8_0),.clk(gclk));
	jdff dff_B_rHfN2sbM6_0(.din(w_dff_B_Vkys7uUa8_0),.dout(w_dff_B_rHfN2sbM6_0),.clk(gclk));
	jdff dff_B_fGBXe76r0_0(.din(n1155),.dout(w_dff_B_fGBXe76r0_0),.clk(gclk));
	jdff dff_B_QWgYZoqw4_0(.din(w_dff_B_fGBXe76r0_0),.dout(w_dff_B_QWgYZoqw4_0),.clk(gclk));
	jdff dff_B_l531TE5W7_1(.din(n1143),.dout(w_dff_B_l531TE5W7_1),.clk(gclk));
	jdff dff_B_gNhm7Jq30_1(.din(w_dff_B_l531TE5W7_1),.dout(w_dff_B_gNhm7Jq30_1),.clk(gclk));
	jdff dff_B_Vg4DbODl7_1(.din(n1145),.dout(w_dff_B_Vg4DbODl7_1),.clk(gclk));
	jdff dff_B_txrUvoTl4_1(.din(n1148),.dout(w_dff_B_txrUvoTl4_1),.clk(gclk));
	jdff dff_A_aDjpHZsX8_1(.dout(w_n899_0[1]),.din(w_dff_A_aDjpHZsX8_1),.clk(gclk));
	jdff dff_A_mKI2h6GU8_1(.dout(w_G87_1[1]),.din(w_dff_A_mKI2h6GU8_1),.clk(gclk));
	jdff dff_A_d7F1LZsA6_2(.dout(w_G87_1[2]),.din(w_dff_A_d7F1LZsA6_2),.clk(gclk));
	jdff dff_A_WKomwQt33_1(.dout(w_G77_2[1]),.din(w_dff_A_WKomwQt33_1),.clk(gclk));
	jdff dff_A_pTgtjDkw0_1(.dout(w_dff_A_WKomwQt33_1),.din(w_dff_A_pTgtjDkw0_1),.clk(gclk));
	jdff dff_A_Jfle1PDM7_1(.dout(w_dff_A_pTgtjDkw0_1),.din(w_dff_A_Jfle1PDM7_1),.clk(gclk));
	jdff dff_A_qIt7Kmcb5_1(.dout(w_dff_A_Jfle1PDM7_1),.din(w_dff_A_qIt7Kmcb5_1),.clk(gclk));
	jdff dff_A_UUP4SJzO6_2(.dout(w_G77_2[2]),.din(w_dff_A_UUP4SJzO6_2),.clk(gclk));
	jdff dff_A_mHDmsGcR5_2(.dout(w_dff_A_UUP4SJzO6_2),.din(w_dff_A_mHDmsGcR5_2),.clk(gclk));
	jdff dff_A_sZ8z3e048_2(.dout(w_dff_A_mHDmsGcR5_2),.din(w_dff_A_sZ8z3e048_2),.clk(gclk));
	jdff dff_A_4vBQYFhr8_2(.dout(w_dff_A_sZ8z3e048_2),.din(w_dff_A_4vBQYFhr8_2),.clk(gclk));
	jdff dff_A_0gSbFn020_1(.dout(w_G283_1[1]),.din(w_dff_A_0gSbFn020_1),.clk(gclk));
	jdff dff_A_KEt89Ekc1_0(.dout(w_n148_3[0]),.din(w_dff_A_KEt89Ekc1_0),.clk(gclk));
	jdff dff_A_x3Kkhbnz1_0(.dout(w_dff_A_KEt89Ekc1_0),.din(w_dff_A_x3Kkhbnz1_0),.clk(gclk));
	jdff dff_A_ih6rqG6O8_0(.dout(w_dff_A_x3Kkhbnz1_0),.din(w_dff_A_ih6rqG6O8_0),.clk(gclk));
	jdff dff_A_U58CLjyT4_0(.dout(w_dff_A_ih6rqG6O8_0),.din(w_dff_A_U58CLjyT4_0),.clk(gclk));
	jdff dff_A_2wQ2Iwbd5_2(.dout(w_n148_3[2]),.din(w_dff_A_2wQ2Iwbd5_2),.clk(gclk));
	jdff dff_A_h94jdN7j6_2(.dout(w_dff_A_2wQ2Iwbd5_2),.din(w_dff_A_h94jdN7j6_2),.clk(gclk));
	jdff dff_A_bvHmkObR7_2(.dout(w_dff_A_h94jdN7j6_2),.din(w_dff_A_bvHmkObR7_2),.clk(gclk));
	jdff dff_A_TtR7O4zu8_1(.dout(w_G294_1[1]),.din(w_dff_A_TtR7O4zu8_1),.clk(gclk));
	jdff dff_B_tY6y2k0Q3_1(.din(n1128),.dout(w_dff_B_tY6y2k0Q3_1),.clk(gclk));
	jdff dff_B_2SeKlOP91_1(.din(n1130),.dout(w_dff_B_2SeKlOP91_1),.clk(gclk));
	jdff dff_B_Qnxe6shB7_1(.din(n1133),.dout(w_dff_B_Qnxe6shB7_1),.clk(gclk));
	jdff dff_B_0c9EyVMM9_0(.din(n1134),.dout(w_dff_B_0c9EyVMM9_0),.clk(gclk));
	jdff dff_A_pOidVMvc1_1(.dout(w_G150_1[1]),.din(w_dff_A_pOidVMvc1_1),.clk(gclk));
	jdff dff_A_oQWicbQb0_2(.dout(w_G150_1[2]),.din(w_dff_A_oQWicbQb0_2),.clk(gclk));
	jdff dff_A_SMHDbw023_0(.dout(w_G128_0[0]),.din(w_dff_A_SMHDbw023_0),.clk(gclk));
	jdff dff_B_PFjQ1lNL0_3(.din(G128),.dout(w_dff_B_PFjQ1lNL0_3),.clk(gclk));
	jdff dff_B_ZdBjMDb04_3(.din(w_dff_B_PFjQ1lNL0_3),.dout(w_dff_B_ZdBjMDb04_3),.clk(gclk));
	jdff dff_B_RnScCPeN8_3(.din(w_dff_B_ZdBjMDb04_3),.dout(w_dff_B_RnScCPeN8_3),.clk(gclk));
	jdff dff_B_WXlW6o9w3_1(.din(n1124),.dout(w_dff_B_WXlW6o9w3_1),.clk(gclk));
	jdff dff_B_fMJ8Nppx0_0(.din(n1126),.dout(w_dff_B_fMJ8Nppx0_0),.clk(gclk));
	jdff dff_A_sSARz3Q60_0(.dout(w_n612_1[0]),.din(w_dff_A_sSARz3Q60_0),.clk(gclk));
	jdff dff_A_zBlBIKOh8_1(.dout(w_n612_1[1]),.din(w_dff_A_zBlBIKOh8_1),.clk(gclk));
	jdff dff_A_ApvMYCUy9_1(.dout(w_dff_A_zBlBIKOh8_1),.din(w_dff_A_ApvMYCUy9_1),.clk(gclk));
	jdff dff_A_CEa41W7O4_1(.dout(w_dff_A_ApvMYCUy9_1),.din(w_dff_A_CEa41W7O4_1),.clk(gclk));
	jdff dff_A_hhva3E7w0_1(.dout(w_dff_A_CEa41W7O4_1),.din(w_dff_A_hhva3E7w0_1),.clk(gclk));
	jdff dff_A_NBZcib8g9_1(.dout(w_dff_A_hhva3E7w0_1),.din(w_dff_A_NBZcib8g9_1),.clk(gclk));
	jdff dff_A_kLq6bmX15_1(.dout(w_dff_A_NBZcib8g9_1),.din(w_dff_A_kLq6bmX15_1),.clk(gclk));
	jdff dff_A_qpAvnoHG2_1(.dout(w_dff_A_kLq6bmX15_1),.din(w_dff_A_qpAvnoHG2_1),.clk(gclk));
	jdff dff_A_zVexCDq21_1(.dout(w_n999_0[1]),.din(w_dff_A_zVexCDq21_1),.clk(gclk));
	jdff dff_A_ImVemRGn4_2(.dout(w_n764_0[2]),.din(w_dff_A_ImVemRGn4_2),.clk(gclk));
	jdff dff_A_Lohcljm11_2(.dout(w_dff_A_ImVemRGn4_2),.din(w_dff_A_Lohcljm11_2),.clk(gclk));
	jdff dff_B_lTVgmxFJ7_0(.din(n763),.dout(w_dff_B_lTVgmxFJ7_0),.clk(gclk));
	jdff dff_B_HkOfbMn44_0(.din(w_dff_B_lTVgmxFJ7_0),.dout(w_dff_B_HkOfbMn44_0),.clk(gclk));
	jdff dff_B_2kSKJuTH6_0(.din(n761),.dout(w_dff_B_2kSKJuTH6_0),.clk(gclk));
	jdff dff_B_0Jc9uF4g1_0(.din(w_dff_B_2kSKJuTH6_0),.dout(w_dff_B_0Jc9uF4g1_0),.clk(gclk));
	jdff dff_A_3xcn83Zx7_0(.dout(w_n760_0[0]),.din(w_dff_A_3xcn83Zx7_0),.clk(gclk));
	jdff dff_B_YExEAZQO6_0(.din(n997),.dout(w_dff_B_YExEAZQO6_0),.clk(gclk));
	jdff dff_B_u4VORMBn5_0(.din(w_dff_B_YExEAZQO6_0),.dout(w_dff_B_u4VORMBn5_0),.clk(gclk));
	jdff dff_B_qKnH7FET3_0(.din(w_dff_B_u4VORMBn5_0),.dout(w_dff_B_qKnH7FET3_0),.clk(gclk));
	jdff dff_B_B7L1Bb4k5_0(.din(w_dff_B_qKnH7FET3_0),.dout(w_dff_B_B7L1Bb4k5_0),.clk(gclk));
	jdff dff_B_9Lpsubch3_0(.din(w_dff_B_B7L1Bb4k5_0),.dout(w_dff_B_9Lpsubch3_0),.clk(gclk));
	jdff dff_A_fzv4lvqZ5_2(.dout(w_n554_1[2]),.din(w_dff_A_fzv4lvqZ5_2),.clk(gclk));
	jdff dff_A_ObJL9Qaa6_1(.dout(w_n519_0[1]),.din(w_dff_A_ObJL9Qaa6_1),.clk(gclk));
	jdff dff_A_Qbg4QAcq7_1(.dout(w_dff_A_ObJL9Qaa6_1),.din(w_dff_A_Qbg4QAcq7_1),.clk(gclk));
	jdff dff_A_6kHp5xAf2_2(.dout(w_n519_0[2]),.din(w_dff_A_6kHp5xAf2_2),.clk(gclk));
	jdff dff_A_tidmV6Lo7_2(.dout(w_dff_A_6kHp5xAf2_2),.din(w_dff_A_tidmV6Lo7_2),.clk(gclk));
	jdff dff_A_fjKKoOcc0_0(.dout(w_n548_0[0]),.din(w_dff_A_fjKKoOcc0_0),.clk(gclk));
	jdff dff_A_ZCBBHjxo5_1(.dout(w_n439_0[1]),.din(w_dff_A_ZCBBHjxo5_1),.clk(gclk));
	jdff dff_A_RpbsJLj51_1(.dout(w_dff_A_ZCBBHjxo5_1),.din(w_dff_A_RpbsJLj51_1),.clk(gclk));
	jdff dff_A_bVqstwWx0_1(.dout(w_dff_A_RpbsJLj51_1),.din(w_dff_A_bVqstwWx0_1),.clk(gclk));
	jdff dff_A_Czkz7sXW1_1(.dout(w_dff_A_bVqstwWx0_1),.din(w_dff_A_Czkz7sXW1_1),.clk(gclk));
	jdff dff_B_Z7Hernbb6_1(.din(n441),.dout(w_dff_B_Z7Hernbb6_1),.clk(gclk));
	jdff dff_B_ubAYFKGy2_1(.din(w_dff_B_Z7Hernbb6_1),.dout(w_dff_B_ubAYFKGy2_1),.clk(gclk));
	jdff dff_A_2IVlRPjg5_1(.dout(w_n436_0[1]),.din(w_dff_A_2IVlRPjg5_1),.clk(gclk));
	jdff dff_B_3aaOt5mu4_1(.din(n424),.dout(w_dff_B_3aaOt5mu4_1),.clk(gclk));
	jdff dff_B_aqXTkkMr3_0(.din(n434),.dout(w_dff_B_aqXTkkMr3_0),.clk(gclk));
	jdff dff_B_VgwORNHx7_0(.din(n423),.dout(w_dff_B_VgwORNHx7_0),.clk(gclk));
	jdff dff_B_Hn1TlILC1_0(.din(w_dff_B_VgwORNHx7_0),.dout(w_dff_B_Hn1TlILC1_0),.clk(gclk));
	jdff dff_B_kXyk0Mo37_1(.din(n413),.dout(w_dff_B_kXyk0Mo37_1),.clk(gclk));
	jdff dff_A_0y4SqIvc2_0(.dout(w_G226_1[0]),.din(w_dff_A_0y4SqIvc2_0),.clk(gclk));
	jdff dff_A_z5vuix598_0(.dout(w_dff_A_0y4SqIvc2_0),.din(w_dff_A_z5vuix598_0),.clk(gclk));
	jdff dff_B_Y6P4RbDG7_1(.din(n493),.dout(w_dff_B_Y6P4RbDG7_1),.clk(gclk));
	jdff dff_B_tU88pgl64_1(.din(w_dff_B_Y6P4RbDG7_1),.dout(w_dff_B_tU88pgl64_1),.clk(gclk));
	jdff dff_A_Mr7Yxxtc5_0(.dout(w_n516_0[0]),.din(w_dff_A_Mr7Yxxtc5_0),.clk(gclk));
	jdff dff_A_Kv3wMfzj6_0(.dout(w_dff_A_Mr7Yxxtc5_0),.din(w_dff_A_Kv3wMfzj6_0),.clk(gclk));
	jdff dff_B_mjwAJ0fu9_0(.din(n514),.dout(w_dff_B_mjwAJ0fu9_0),.clk(gclk));
	jdff dff_B_pJ9vBfb10_1(.din(n485),.dout(w_dff_B_pJ9vBfb10_1),.clk(gclk));
	jdff dff_B_QBUlf6Y68_1(.din(n496),.dout(w_dff_B_QBUlf6Y68_1),.clk(gclk));
	jdff dff_B_fFkLKxll7_1(.din(w_dff_B_QBUlf6Y68_1),.dout(w_dff_B_fFkLKxll7_1),.clk(gclk));
	jdff dff_B_E3nHGAMP2_1(.din(w_dff_B_fFkLKxll7_1),.dout(w_dff_B_E3nHGAMP2_1),.clk(gclk));
	jdff dff_B_d1fElbSb7_0(.din(n505),.dout(w_dff_B_d1fElbSb7_0),.clk(gclk));
	jdff dff_B_Qwl99s273_0(.din(w_dff_B_d1fElbSb7_0),.dout(w_dff_B_Qwl99s273_0),.clk(gclk));
	jdff dff_B_Do6o7OWl5_1(.din(n497),.dout(w_dff_B_Do6o7OWl5_1),.clk(gclk));
	jdff dff_B_qsInAYaB2_1(.din(w_dff_B_Do6o7OWl5_1),.dout(w_dff_B_qsInAYaB2_1),.clk(gclk));
	jdff dff_B_YL6HbYWE5_1(.din(w_dff_B_qsInAYaB2_1),.dout(w_dff_B_YL6HbYWE5_1),.clk(gclk));
	jdff dff_A_iiFMhJsK0_1(.dout(w_n541_0[1]),.din(w_dff_A_iiFMhJsK0_1),.clk(gclk));
	jdff dff_A_H2zRB4zY0_1(.dout(w_dff_A_iiFMhJsK0_1),.din(w_dff_A_H2zRB4zY0_1),.clk(gclk));
	jdff dff_B_ZtZugRSf2_1(.din(n456),.dout(w_dff_B_ZtZugRSf2_1),.clk(gclk));
	jdff dff_B_CaBe6qHK8_1(.din(w_dff_B_ZtZugRSf2_1),.dout(w_dff_B_CaBe6qHK8_1),.clk(gclk));
	jdff dff_A_yHGBWbls2_0(.dout(w_n483_0[0]),.din(w_dff_A_yHGBWbls2_0),.clk(gclk));
	jdff dff_A_JChnqbdl4_0(.dout(w_dff_A_yHGBWbls2_0),.din(w_dff_A_JChnqbdl4_0),.clk(gclk));
	jdff dff_A_kl66bIPt4_0(.dout(w_dff_A_JChnqbdl4_0),.din(w_dff_A_kl66bIPt4_0),.clk(gclk));
	jdff dff_A_OF2BZT4e7_0(.dout(w_dff_A_kl66bIPt4_0),.din(w_dff_A_OF2BZT4e7_0),.clk(gclk));
	jdff dff_B_GpNB0XTN4_0(.din(n481),.dout(w_dff_B_GpNB0XTN4_0),.clk(gclk));
	jdff dff_A_eCFQ9eAD7_1(.dout(w_G226_0[1]),.din(w_dff_A_eCFQ9eAD7_1),.clk(gclk));
	jdff dff_A_khPh2FFN8_1(.dout(w_dff_A_eCFQ9eAD7_1),.din(w_dff_A_khPh2FFN8_1),.clk(gclk));
	jdff dff_A_z5f1lVWD4_2(.dout(w_G226_0[2]),.din(w_dff_A_z5f1lVWD4_2),.clk(gclk));
	jdff dff_A_6eS5xXQT3_2(.dout(w_dff_A_z5f1lVWD4_2),.din(w_dff_A_6eS5xXQT3_2),.clk(gclk));
	jdff dff_A_xE7CJdnU0_2(.dout(w_dff_A_6eS5xXQT3_2),.din(w_dff_A_xE7CJdnU0_2),.clk(gclk));
	jdff dff_A_K5vSNaX49_2(.dout(w_dff_A_xE7CJdnU0_2),.din(w_dff_A_K5vSNaX49_2),.clk(gclk));
	jdff dff_B_PusZ0kJy6_1(.din(n448),.dout(w_dff_B_PusZ0kJy6_1),.clk(gclk));
	jdff dff_B_Nv2GfN377_1(.din(G222),.dout(w_dff_B_Nv2GfN377_1),.clk(gclk));
	jdff dff_B_ymDCuxVv0_1(.din(w_dff_B_Nv2GfN377_1),.dout(w_dff_B_ymDCuxVv0_1),.clk(gclk));
	jdff dff_A_JFeIDYY74_0(.dout(w_n430_0[0]),.din(w_dff_A_JFeIDYY74_0),.clk(gclk));
	jdff dff_B_C0Fl309u4_2(.din(n430),.dout(w_dff_B_C0Fl309u4_2),.clk(gclk));
	jdff dff_A_TiB3qEKA3_1(.dout(w_G77_3[1]),.din(w_dff_A_TiB3qEKA3_1),.clk(gclk));
	jdff dff_A_UVDxzX8X4_1(.dout(w_dff_A_TiB3qEKA3_1),.din(w_dff_A_UVDxzX8X4_1),.clk(gclk));
	jdff dff_A_O31Yevz94_1(.dout(w_dff_A_UVDxzX8X4_1),.din(w_dff_A_O31Yevz94_1),.clk(gclk));
	jdff dff_B_ZA4Xncnc2_2(.din(G223),.dout(w_dff_B_ZA4Xncnc2_2),.clk(gclk));
	jdff dff_B_3TZf6n5G1_2(.din(w_dff_B_ZA4Xncnc2_2),.dout(w_dff_B_3TZf6n5G1_2),.clk(gclk));
	jdff dff_B_5ysRGQcf9_1(.din(n459),.dout(w_dff_B_5ysRGQcf9_1),.clk(gclk));
	jdff dff_B_3Teu5xFQ4_1(.din(w_dff_B_5ysRGQcf9_1),.dout(w_dff_B_3Teu5xFQ4_1),.clk(gclk));
	jdff dff_B_7vdPgLY42_1(.din(w_dff_B_3Teu5xFQ4_1),.dout(w_dff_B_7vdPgLY42_1),.clk(gclk));
	jdff dff_B_jWr6xEqu8_0(.din(n472),.dout(w_dff_B_jWr6xEqu8_0),.clk(gclk));
	jdff dff_B_7SgsIywN8_0(.din(w_dff_B_jWr6xEqu8_0),.dout(w_dff_B_7SgsIywN8_0),.clk(gclk));
	jdff dff_A_Nwsjq0xo4_2(.dout(w_n185_1[2]),.din(w_dff_A_Nwsjq0xo4_2),.clk(gclk));
	jdff dff_B_oW9LfIcp4_1(.din(n460),.dout(w_dff_B_oW9LfIcp4_1),.clk(gclk));
	jdff dff_B_3fcaVetG8_1(.din(n461),.dout(w_dff_B_3fcaVetG8_1),.clk(gclk));
	jdff dff_B_6GLiXLf15_1(.din(w_dff_B_3fcaVetG8_1),.dout(w_dff_B_6GLiXLf15_1),.clk(gclk));
	jdff dff_A_OY2GCQl84_1(.dout(w_n75_0[1]),.din(w_dff_A_OY2GCQl84_1),.clk(gclk));
	jdff dff_A_iJX6d4KT1_1(.dout(w_dff_A_OY2GCQl84_1),.din(w_dff_A_iJX6d4KT1_1),.clk(gclk));
	jdff dff_A_h1U14QZ20_1(.dout(w_dff_A_iJX6d4KT1_1),.din(w_dff_A_h1U14QZ20_1),.clk(gclk));
	jdff dff_A_cQXYitet4_2(.dout(w_n75_0[2]),.din(w_dff_A_cQXYitet4_2),.clk(gclk));
	jdff dff_A_nBSbsODQ5_2(.dout(w_dff_A_cQXYitet4_2),.din(w_dff_A_nBSbsODQ5_2),.clk(gclk));
	jdff dff_A_sPbkiv5R3_2(.dout(w_dff_A_nBSbsODQ5_2),.din(w_dff_A_sPbkiv5R3_2),.clk(gclk));
	jdff dff_A_MwT9xHbC5_2(.dout(w_dff_A_sPbkiv5R3_2),.din(w_dff_A_MwT9xHbC5_2),.clk(gclk));
	jdff dff_A_45ig0oRf4_1(.dout(w_n74_0[1]),.din(w_dff_A_45ig0oRf4_1),.clk(gclk));
	jdff dff_A_XNuT9Fvx8_1(.dout(w_dff_A_45ig0oRf4_1),.din(w_dff_A_XNuT9Fvx8_1),.clk(gclk));
	jdff dff_A_tPqs1ct78_1(.dout(w_dff_A_XNuT9Fvx8_1),.din(w_dff_A_tPqs1ct78_1),.clk(gclk));
	jdff dff_A_JEStj55Q1_2(.dout(w_n74_0[2]),.din(w_dff_A_JEStj55Q1_2),.clk(gclk));
	jdff dff_A_efvVhaa88_2(.dout(w_dff_A_JEStj55Q1_2),.din(w_dff_A_efvVhaa88_2),.clk(gclk));
	jdff dff_A_DwRq8D7V4_0(.dout(w_n73_2[0]),.din(w_dff_A_DwRq8D7V4_0),.clk(gclk));
	jdff dff_A_OzhMKkGv7_0(.dout(w_dff_A_DwRq8D7V4_0),.din(w_dff_A_OzhMKkGv7_0),.clk(gclk));
	jdff dff_A_PVARDvkW4_2(.dout(w_n73_2[2]),.din(w_dff_A_PVARDvkW4_2),.clk(gclk));
	jdff dff_A_puSTSz594_2(.dout(w_n73_0[2]),.din(w_dff_A_puSTSz594_2),.clk(gclk));
	jdff dff_A_EL2YGJlr6_2(.dout(w_dff_A_puSTSz594_2),.din(w_dff_A_EL2YGJlr6_2),.clk(gclk));
	jdff dff_A_y6OI6irt9_2(.dout(w_dff_A_EL2YGJlr6_2),.din(w_dff_A_y6OI6irt9_2),.clk(gclk));
	jdff dff_A_ayd9RTX27_1(.dout(w_G50_5[1]),.din(w_dff_A_ayd9RTX27_1),.clk(gclk));
	jdff dff_A_0UwmGFFC3_1(.dout(w_dff_A_ayd9RTX27_1),.din(w_dff_A_0UwmGFFC3_1),.clk(gclk));
	jdff dff_A_dc4sKXuE5_1(.dout(w_dff_A_0UwmGFFC3_1),.din(w_dff_A_dc4sKXuE5_1),.clk(gclk));
	jdff dff_A_pJ3juYXa6_0(.dout(w_G50_4[0]),.din(w_dff_A_pJ3juYXa6_0),.clk(gclk));
	jdff dff_A_UyoE6NVP6_0(.dout(w_dff_A_pJ3juYXa6_0),.din(w_dff_A_UyoE6NVP6_0),.clk(gclk));
	jdff dff_A_AEGITx9G9_1(.dout(w_G50_4[1]),.din(w_dff_A_AEGITx9G9_1),.clk(gclk));
	jdff dff_A_n01tZAbE4_0(.dout(w_G50_1[0]),.din(w_dff_A_n01tZAbE4_0),.clk(gclk));
	jdff dff_A_scg5wolC8_2(.dout(w_G50_1[2]),.din(w_dff_A_scg5wolC8_2),.clk(gclk));
	jdff dff_A_8FLMUrlX5_2(.dout(w_dff_A_scg5wolC8_2),.din(w_dff_A_8FLMUrlX5_2),.clk(gclk));
	jdff dff_A_0dGGcx4t0_2(.dout(w_dff_A_8FLMUrlX5_2),.din(w_dff_A_0dGGcx4t0_2),.clk(gclk));
	jdff dff_A_sQxHYeYf6_2(.dout(w_dff_A_0dGGcx4t0_2),.din(w_dff_A_sQxHYeYf6_2),.clk(gclk));
	jdff dff_A_zwqU6G3F3_0(.dout(w_G384_0),.din(w_dff_A_zwqU6G3F3_0),.clk(gclk));
	jdff dff_A_ndypIZMF9_0(.dout(w_dff_A_zwqU6G3F3_0),.din(w_dff_A_ndypIZMF9_0),.clk(gclk));
	jdff dff_A_Jz517UPj8_0(.dout(w_n750_0[0]),.din(w_dff_A_Jz517UPj8_0),.clk(gclk));
	jdff dff_A_cIUoVB911_0(.dout(w_dff_A_Jz517UPj8_0),.din(w_dff_A_cIUoVB911_0),.clk(gclk));
	jdff dff_B_6Uzw4xNH4_0(.din(n747),.dout(w_dff_B_6Uzw4xNH4_0),.clk(gclk));
	jdff dff_B_Oz0vXoYE2_0(.din(w_dff_B_6Uzw4xNH4_0),.dout(w_dff_B_Oz0vXoYE2_0),.clk(gclk));
	jdff dff_B_SfEUcmPy1_0(.din(w_dff_B_Oz0vXoYE2_0),.dout(w_dff_B_SfEUcmPy1_0),.clk(gclk));
	jdff dff_B_3Tn9GTCJ1_0(.din(n746),.dout(w_dff_B_3Tn9GTCJ1_0),.clk(gclk));
	jdff dff_B_fwNpmsjn6_0(.din(w_dff_B_3Tn9GTCJ1_0),.dout(w_dff_B_fwNpmsjn6_0),.clk(gclk));
	jdff dff_B_ddHmRJrI4_0(.din(w_dff_B_fwNpmsjn6_0),.dout(w_dff_B_ddHmRJrI4_0),.clk(gclk));
	jdff dff_B_QLeR7zmG1_0(.din(w_dff_B_ddHmRJrI4_0),.dout(w_dff_B_QLeR7zmG1_0),.clk(gclk));
	jdff dff_B_kW1l0wiA6_0(.din(n744),.dout(w_dff_B_kW1l0wiA6_0),.clk(gclk));
	jdff dff_B_huqK92bP3_0(.din(w_dff_B_kW1l0wiA6_0),.dout(w_dff_B_huqK92bP3_0),.clk(gclk));
	jdff dff_A_kdtt9xD15_2(.dout(w_n605_1[2]),.din(w_dff_A_kdtt9xD15_2),.clk(gclk));
	jdff dff_A_sjnLsLoA7_2(.dout(w_dff_A_kdtt9xD15_2),.din(w_dff_A_sjnLsLoA7_2),.clk(gclk));
	jdff dff_A_G4bUzfxV5_2(.dout(w_dff_A_sjnLsLoA7_2),.din(w_dff_A_G4bUzfxV5_2),.clk(gclk));
	jdff dff_A_SCpKaUiZ8_2(.dout(w_dff_A_G4bUzfxV5_2),.din(w_dff_A_SCpKaUiZ8_2),.clk(gclk));
	jdff dff_A_W39ACTMm9_2(.dout(w_dff_A_SCpKaUiZ8_2),.din(w_dff_A_W39ACTMm9_2),.clk(gclk));
	jdff dff_A_AtOJHKKB4_2(.dout(w_dff_A_W39ACTMm9_2),.din(w_dff_A_AtOJHKKB4_2),.clk(gclk));
	jdff dff_A_VIUQCjfj6_2(.dout(w_dff_A_AtOJHKKB4_2),.din(w_dff_A_VIUQCjfj6_2),.clk(gclk));
	jdff dff_A_a5wMNEEO6_2(.dout(w_dff_A_VIUQCjfj6_2),.din(w_dff_A_a5wMNEEO6_2),.clk(gclk));
	jdff dff_A_ZJcudOfX8_0(.dout(w_n604_2[0]),.din(w_dff_A_ZJcudOfX8_0),.clk(gclk));
	jdff dff_A_OJPfcFCa2_0(.dout(w_dff_A_ZJcudOfX8_0),.din(w_dff_A_OJPfcFCa2_0),.clk(gclk));
	jdff dff_A_2EEPRluq6_0(.dout(w_dff_A_OJPfcFCa2_0),.din(w_dff_A_2EEPRluq6_0),.clk(gclk));
	jdff dff_A_kKrqoSoW7_0(.dout(w_dff_A_2EEPRluq6_0),.din(w_dff_A_kKrqoSoW7_0),.clk(gclk));
	jdff dff_B_3h42XZni7_1(.din(n721),.dout(w_dff_B_3h42XZni7_1),.clk(gclk));
	jdff dff_B_kltxwDtL7_1(.din(w_dff_B_3h42XZni7_1),.dout(w_dff_B_kltxwDtL7_1),.clk(gclk));
	jdff dff_B_aEOYgQuj1_1(.din(n727),.dout(w_dff_B_aEOYgQuj1_1),.clk(gclk));
	jdff dff_B_iyLyyVWW7_1(.din(n730),.dout(w_dff_B_iyLyyVWW7_1),.clk(gclk));
	jdff dff_B_ZxTVggiG3_1(.din(n733),.dout(w_dff_B_ZxTVggiG3_1),.clk(gclk));
	jdff dff_B_ZNVwHKRe3_0(.din(n734),.dout(w_dff_B_ZNVwHKRe3_0),.clk(gclk));
	jdff dff_A_dWwjfL9n6_0(.dout(w_G294_2[0]),.din(w_dff_A_dWwjfL9n6_0),.clk(gclk));
	jdff dff_A_HaSaHwL92_0(.dout(w_G116_3[0]),.din(w_dff_A_HaSaHwL92_0),.clk(gclk));
	jdff dff_A_Au7l3aAv2_0(.dout(w_dff_A_HaSaHwL92_0),.din(w_dff_A_Au7l3aAv2_0),.clk(gclk));
	jdff dff_A_gbf3SjqU5_0(.dout(w_dff_A_Au7l3aAv2_0),.din(w_dff_A_gbf3SjqU5_0),.clk(gclk));
	jdff dff_A_oXNKXIQd4_2(.dout(w_G116_3[2]),.din(w_dff_A_oXNKXIQd4_2),.clk(gclk));
	jdff dff_A_RRAZWhbs1_2(.dout(w_dff_A_oXNKXIQd4_2),.din(w_dff_A_RRAZWhbs1_2),.clk(gclk));
	jdff dff_A_nByLp5Ye4_0(.dout(w_G33_5[0]),.din(w_dff_A_nByLp5Ye4_0),.clk(gclk));
	jdff dff_A_vlp8hzqz8_2(.dout(w_G33_5[2]),.din(w_dff_A_vlp8hzqz8_2),.clk(gclk));
	jdff dff_A_8G95VIjC4_2(.dout(w_dff_A_vlp8hzqz8_2),.din(w_dff_A_8G95VIjC4_2),.clk(gclk));
	jdff dff_B_IAYrVm0P9_1(.din(n722),.dout(w_dff_B_IAYrVm0P9_1),.clk(gclk));
	jdff dff_B_kbc6CHlm6_0(.din(n724),.dout(w_dff_B_kbc6CHlm6_0),.clk(gclk));
	jdff dff_A_Rbqv7i2E2_1(.dout(w_G311_1[1]),.din(w_dff_A_Rbqv7i2E2_1),.clk(gclk));
	jdff dff_B_3Zls9Asu0_3(.din(G311),.dout(w_dff_B_3Zls9Asu0_3),.clk(gclk));
	jdff dff_B_UKTj6RAy9_3(.din(w_dff_B_3Zls9Asu0_3),.dout(w_dff_B_UKTj6RAy9_3),.clk(gclk));
	jdff dff_B_mqa966gy6_3(.din(w_dff_B_UKTj6RAy9_3),.dout(w_dff_B_mqa966gy6_3),.clk(gclk));
	jdff dff_B_0Qpqs9IT5_1(.din(n710),.dout(w_dff_B_0Qpqs9IT5_1),.clk(gclk));
	jdff dff_B_qOHNn4DT0_1(.din(n712),.dout(w_dff_B_qOHNn4DT0_1),.clk(gclk));
	jdff dff_B_mA1TS2tU5_1(.din(n715),.dout(w_dff_B_mA1TS2tU5_1),.clk(gclk));
	jdff dff_B_2WoV4lU33_1(.din(n716),.dout(w_dff_B_2WoV4lU33_1),.clk(gclk));
	jdff dff_A_gYiziej66_1(.dout(w_G68_3[1]),.din(w_dff_A_gYiziej66_1),.clk(gclk));
	jdff dff_A_EuaQOspZ3_1(.dout(w_dff_A_gYiziej66_1),.din(w_dff_A_EuaQOspZ3_1),.clk(gclk));
	jdff dff_A_2pHJVp7l8_1(.dout(w_dff_A_EuaQOspZ3_1),.din(w_dff_A_2pHJVp7l8_1),.clk(gclk));
	jdff dff_A_jZRrQYj11_2(.dout(w_G68_3[2]),.din(w_dff_A_jZRrQYj11_2),.clk(gclk));
	jdff dff_A_9JmFPU7u0_2(.dout(w_dff_A_jZRrQYj11_2),.din(w_dff_A_9JmFPU7u0_2),.clk(gclk));
	jdff dff_A_36uqRPDS7_1(.dout(w_G137_1[1]),.din(w_dff_A_36uqRPDS7_1),.clk(gclk));
	jdff dff_B_aHADKo1m3_3(.din(G137),.dout(w_dff_B_aHADKo1m3_3),.clk(gclk));
	jdff dff_B_BfoOu98b4_3(.din(w_dff_B_aHADKo1m3_3),.dout(w_dff_B_BfoOu98b4_3),.clk(gclk));
	jdff dff_B_a8BNTn3r7_3(.din(w_dff_B_BfoOu98b4_3),.dout(w_dff_B_a8BNTn3r7_3),.clk(gclk));
	jdff dff_B_HTpOZOSe8_3(.din(G143),.dout(w_dff_B_HTpOZOSe8_3),.clk(gclk));
	jdff dff_B_e3iksa357_3(.din(w_dff_B_HTpOZOSe8_3),.dout(w_dff_B_e3iksa357_3),.clk(gclk));
	jdff dff_B_9juV44ph8_3(.din(w_dff_B_e3iksa357_3),.dout(w_dff_B_9juV44ph8_3),.clk(gclk));
	jdff dff_A_ZKbKDlC72_0(.dout(w_G159_3[0]),.din(w_dff_A_ZKbKDlC72_0),.clk(gclk));
	jdff dff_A_hvwHxbc04_1(.dout(w_G159_3[1]),.din(w_dff_A_hvwHxbc04_1),.clk(gclk));
	jdff dff_A_Jkc8FQ2x6_1(.dout(w_dff_A_hvwHxbc04_1),.din(w_dff_A_Jkc8FQ2x6_1),.clk(gclk));
	jdff dff_A_ML8Wsi7R7_0(.dout(w_G159_0[0]),.din(w_dff_A_ML8Wsi7R7_0),.clk(gclk));
	jdff dff_A_VmKgOIih9_0(.dout(w_dff_A_ML8Wsi7R7_0),.din(w_dff_A_VmKgOIih9_0),.clk(gclk));
	jdff dff_A_QZZj3G500_1(.dout(w_G159_0[1]),.din(w_dff_A_QZZj3G500_1),.clk(gclk));
	jdff dff_B_qkfBigxd2_3(.din(G159),.dout(w_dff_B_qkfBigxd2_3),.clk(gclk));
	jdff dff_B_CuiEmr8G7_3(.din(w_dff_B_qkfBigxd2_3),.dout(w_dff_B_CuiEmr8G7_3),.clk(gclk));
	jdff dff_A_SktWqd4B6_1(.dout(w_G190_2[1]),.din(w_dff_A_SktWqd4B6_1),.clk(gclk));
	jdff dff_A_ngQMY0wi1_1(.dout(w_dff_A_SktWqd4B6_1),.din(w_dff_A_ngQMY0wi1_1),.clk(gclk));
	jdff dff_A_pnXBJf900_1(.dout(w_dff_A_ngQMY0wi1_1),.din(w_dff_A_pnXBJf900_1),.clk(gclk));
	jdff dff_A_HraerFyz3_1(.dout(w_dff_A_pnXBJf900_1),.din(w_dff_A_HraerFyz3_1),.clk(gclk));
	jdff dff_A_CAXAfBzv5_1(.dout(w_dff_A_HraerFyz3_1),.din(w_dff_A_CAXAfBzv5_1),.clk(gclk));
	jdff dff_A_qthwE6YC3_2(.dout(w_G190_2[2]),.din(w_dff_A_qthwE6YC3_2),.clk(gclk));
	jdff dff_A_sGBZWvyE2_2(.dout(w_dff_A_qthwE6YC3_2),.din(w_dff_A_sGBZWvyE2_2),.clk(gclk));
	jdff dff_A_eSlwqHHA1_2(.dout(w_dff_A_sGBZWvyE2_2),.din(w_dff_A_eSlwqHHA1_2),.clk(gclk));
	jdff dff_A_X6IwQgEE1_2(.dout(w_dff_A_eSlwqHHA1_2),.din(w_dff_A_X6IwQgEE1_2),.clk(gclk));
	jdff dff_A_pNsegoOF1_2(.dout(w_dff_A_X6IwQgEE1_2),.din(w_dff_A_pNsegoOF1_2),.clk(gclk));
	jdff dff_A_rPHqTFGY3_0(.dout(w_G50_3[0]),.din(w_dff_A_rPHqTFGY3_0),.clk(gclk));
	jdff dff_A_QROsBE3b5_0(.dout(w_dff_A_rPHqTFGY3_0),.din(w_dff_A_QROsBE3b5_0),.clk(gclk));
	jdff dff_A_o3YWIpC56_0(.dout(w_dff_A_QROsBE3b5_0),.din(w_dff_A_o3YWIpC56_0),.clk(gclk));
	jdff dff_A_Babz9X3p5_2(.dout(w_G50_3[2]),.din(w_dff_A_Babz9X3p5_2),.clk(gclk));
	jdff dff_A_Y3f56pMO3_2(.dout(w_dff_A_Babz9X3p5_2),.din(w_dff_A_Y3f56pMO3_2),.clk(gclk));
	jdff dff_A_xOecG1PY4_2(.dout(w_dff_A_Y3f56pMO3_2),.din(w_dff_A_xOecG1PY4_2),.clk(gclk));
	jdff dff_A_r1HWMIYL7_2(.dout(w_dff_A_xOecG1PY4_2),.din(w_dff_A_r1HWMIYL7_2),.clk(gclk));
	jdff dff_A_3Dlfw6DB4_1(.dout(w_G50_0[1]),.din(w_dff_A_3Dlfw6DB4_1),.clk(gclk));
	jdff dff_A_8RbOiNs66_1(.dout(w_dff_A_3Dlfw6DB4_1),.din(w_dff_A_8RbOiNs66_1),.clk(gclk));
	jdff dff_A_ZukS50L22_1(.dout(w_dff_A_8RbOiNs66_1),.din(w_dff_A_ZukS50L22_1),.clk(gclk));
	jdff dff_A_DHGzt0N55_0(.dout(w_G33_6[0]),.din(w_dff_A_DHGzt0N55_0),.clk(gclk));
	jdff dff_A_RppjfKcu5_0(.dout(w_dff_A_DHGzt0N55_0),.din(w_dff_A_RppjfKcu5_0),.clk(gclk));
	jdff dff_A_hEyGmNLP2_0(.dout(w_dff_A_RppjfKcu5_0),.din(w_dff_A_hEyGmNLP2_0),.clk(gclk));
	jdff dff_A_RACd9pjg9_0(.dout(w_dff_A_hEyGmNLP2_0),.din(w_dff_A_RACd9pjg9_0),.clk(gclk));
	jdff dff_A_4PgoHSVp7_1(.dout(w_G33_6[1]),.din(w_dff_A_4PgoHSVp7_1),.clk(gclk));
	jdff dff_A_oDlAgc7P2_1(.dout(w_dff_A_4PgoHSVp7_1),.din(w_dff_A_oDlAgc7P2_1),.clk(gclk));
	jdff dff_A_ybsNGNwS9_1(.dout(w_G33_1[1]),.din(w_dff_A_ybsNGNwS9_1),.clk(gclk));
	jdff dff_A_uXXzrEnG6_1(.dout(w_dff_A_ybsNGNwS9_1),.din(w_dff_A_uXXzrEnG6_1),.clk(gclk));
	jdff dff_A_JkA8zOvk6_1(.dout(w_dff_A_uXXzrEnG6_1),.din(w_dff_A_JkA8zOvk6_1),.clk(gclk));
	jdff dff_B_y90EBVFx6_1(.din(n706),.dout(w_dff_B_y90EBVFx6_1),.clk(gclk));
	jdff dff_B_h2dKfwho3_0(.din(n708),.dout(w_dff_B_h2dKfwho3_0),.clk(gclk));
	jdff dff_A_aPGmUDHU2_0(.dout(w_G150_3[0]),.din(w_dff_A_aPGmUDHU2_0),.clk(gclk));
	jdff dff_A_5v8xR5wt0_0(.dout(w_dff_A_aPGmUDHU2_0),.din(w_dff_A_5v8xR5wt0_0),.clk(gclk));
	jdff dff_A_wgMpoDW27_0(.dout(w_dff_A_5v8xR5wt0_0),.din(w_dff_A_wgMpoDW27_0),.clk(gclk));
	jdff dff_A_otD5R4BN9_0(.dout(w_G150_0[0]),.din(w_dff_A_otD5R4BN9_0),.clk(gclk));
	jdff dff_A_yX6ndfia3_0(.dout(w_dff_A_otD5R4BN9_0),.din(w_dff_A_yX6ndfia3_0),.clk(gclk));
	jdff dff_A_NQlKKxwd2_0(.dout(w_dff_A_yX6ndfia3_0),.din(w_dff_A_NQlKKxwd2_0),.clk(gclk));
	jdff dff_A_NkwA5IIM6_1(.dout(w_G150_0[1]),.din(w_dff_A_NkwA5IIM6_1),.clk(gclk));
	jdff dff_A_8Xx64vZW0_1(.dout(w_dff_A_NkwA5IIM6_1),.din(w_dff_A_8Xx64vZW0_1),.clk(gclk));
	jdff dff_A_UpKDQn5S3_1(.dout(w_dff_A_8Xx64vZW0_1),.din(w_dff_A_UpKDQn5S3_1),.clk(gclk));
	jdff dff_A_r5Tudtj48_0(.dout(w_G58_3[0]),.din(w_dff_A_r5Tudtj48_0),.clk(gclk));
	jdff dff_A_Rn3uLTyX2_1(.dout(w_G58_3[1]),.din(w_dff_A_Rn3uLTyX2_1),.clk(gclk));
	jdff dff_A_O0F2LtgJ8_1(.dout(w_n615_0[1]),.din(w_dff_A_O0F2LtgJ8_1),.clk(gclk));
	jdff dff_A_IlhzGVfX4_1(.dout(w_G200_2[1]),.din(w_dff_A_IlhzGVfX4_1),.clk(gclk));
	jdff dff_A_WbvVSi4P5_1(.dout(w_dff_A_IlhzGVfX4_1),.din(w_dff_A_WbvVSi4P5_1),.clk(gclk));
	jdff dff_A_p9A7aHDN9_1(.dout(w_dff_A_WbvVSi4P5_1),.din(w_dff_A_p9A7aHDN9_1),.clk(gclk));
	jdff dff_A_U7BP3JGa3_1(.dout(w_dff_A_p9A7aHDN9_1),.din(w_dff_A_U7BP3JGa3_1),.clk(gclk));
	jdff dff_A_qmAdwVV27_1(.dout(w_dff_A_U7BP3JGa3_1),.din(w_dff_A_qmAdwVV27_1),.clk(gclk));
	jdff dff_A_mz2Ma50S4_1(.dout(w_dff_A_qmAdwVV27_1),.din(w_dff_A_mz2Ma50S4_1),.clk(gclk));
	jdff dff_A_3g9wCvOT0_1(.dout(w_dff_A_mz2Ma50S4_1),.din(w_dff_A_3g9wCvOT0_1),.clk(gclk));
	jdff dff_A_im6BpvSm3_2(.dout(w_G200_2[2]),.din(w_dff_A_im6BpvSm3_2),.clk(gclk));
	jdff dff_A_37RYzBOf2_2(.dout(w_dff_A_im6BpvSm3_2),.din(w_dff_A_37RYzBOf2_2),.clk(gclk));
	jdff dff_A_Cd5N8OoT3_2(.dout(w_dff_A_37RYzBOf2_2),.din(w_dff_A_Cd5N8OoT3_2),.clk(gclk));
	jdff dff_A_ImJQOAUL9_2(.dout(w_dff_A_Cd5N8OoT3_2),.din(w_dff_A_ImJQOAUL9_2),.clk(gclk));
	jdff dff_A_b7z7NBeM2_2(.dout(w_dff_A_ImJQOAUL9_2),.din(w_dff_A_b7z7NBeM2_2),.clk(gclk));
	jdff dff_A_vZuHoIeq9_2(.dout(w_dff_A_b7z7NBeM2_2),.din(w_dff_A_vZuHoIeq9_2),.clk(gclk));
	jdff dff_A_UHz0db1u2_2(.dout(w_dff_A_vZuHoIeq9_2),.din(w_dff_A_UHz0db1u2_2),.clk(gclk));
	jdff dff_A_V3ymdB0E2_0(.dout(w_n619_0[0]),.din(w_dff_A_V3ymdB0E2_0),.clk(gclk));
	jdff dff_A_Zn9s1wEB5_0(.dout(w_n407_1[0]),.din(w_dff_A_Zn9s1wEB5_0),.clk(gclk));
	jdff dff_A_QvwrTc9j0_1(.dout(w_n407_1[1]),.din(w_dff_A_QvwrTc9j0_1),.clk(gclk));
	jdff dff_A_ZwLwUUqu8_1(.dout(w_dff_A_QvwrTc9j0_1),.din(w_dff_A_ZwLwUUqu8_1),.clk(gclk));
	jdff dff_A_BmJHWTNA3_1(.dout(w_G132_1[1]),.din(w_dff_A_BmJHWTNA3_1),.clk(gclk));
	jdff dff_B_koyEFjA78_3(.din(G132),.dout(w_dff_B_koyEFjA78_3),.clk(gclk));
	jdff dff_B_vdjU1Jx73_3(.din(w_dff_B_koyEFjA78_3),.dout(w_dff_B_vdjU1Jx73_3),.clk(gclk));
	jdff dff_B_9BanF2Hg6_3(.din(w_dff_B_vdjU1Jx73_3),.dout(w_dff_B_9BanF2Hg6_3),.clk(gclk));
	jdff dff_A_jXoD36EM4_0(.dout(w_n612_3[0]),.din(w_dff_A_jXoD36EM4_0),.clk(gclk));
	jdff dff_A_MJe5nHEv3_0(.dout(w_dff_A_jXoD36EM4_0),.din(w_dff_A_MJe5nHEv3_0),.clk(gclk));
	jdff dff_A_z3nenk1G6_0(.dout(w_dff_A_MJe5nHEv3_0),.din(w_dff_A_z3nenk1G6_0),.clk(gclk));
	jdff dff_A_b59GNd0f5_0(.dout(w_dff_A_z3nenk1G6_0),.din(w_dff_A_b59GNd0f5_0),.clk(gclk));
	jdff dff_A_x9e5xlAp3_0(.dout(w_dff_A_b59GNd0f5_0),.din(w_dff_A_x9e5xlAp3_0),.clk(gclk));
	jdff dff_A_lTvxQf551_0(.dout(w_dff_A_x9e5xlAp3_0),.din(w_dff_A_lTvxQf551_0),.clk(gclk));
	jdff dff_A_y2vQ4Fxq2_0(.dout(w_dff_A_lTvxQf551_0),.din(w_dff_A_y2vQ4Fxq2_0),.clk(gclk));
	jdff dff_A_rVInVeyA9_0(.dout(w_dff_A_y2vQ4Fxq2_0),.din(w_dff_A_rVInVeyA9_0),.clk(gclk));
	jdff dff_A_bOjiu0b69_0(.dout(w_dff_A_rVInVeyA9_0),.din(w_dff_A_bOjiu0b69_0),.clk(gclk));
	jdff dff_A_orL5Xhbm1_2(.dout(w_n612_3[2]),.din(w_dff_A_orL5Xhbm1_2),.clk(gclk));
	jdff dff_A_6LUEUNu30_2(.dout(w_dff_A_orL5Xhbm1_2),.din(w_dff_A_6LUEUNu30_2),.clk(gclk));
	jdff dff_A_p8SEAqju9_2(.dout(w_dff_A_6LUEUNu30_2),.din(w_dff_A_p8SEAqju9_2),.clk(gclk));
	jdff dff_A_A7y32vC20_2(.dout(w_dff_A_p8SEAqju9_2),.din(w_dff_A_A7y32vC20_2),.clk(gclk));
	jdff dff_A_CWC3RigB3_2(.dout(w_dff_A_A7y32vC20_2),.din(w_dff_A_CWC3RigB3_2),.clk(gclk));
	jdff dff_A_5arkXnx99_2(.dout(w_dff_A_CWC3RigB3_2),.din(w_dff_A_5arkXnx99_2),.clk(gclk));
	jdff dff_A_Ul0QIhXY5_2(.dout(w_dff_A_5arkXnx99_2),.din(w_dff_A_Ul0QIhXY5_2),.clk(gclk));
	jdff dff_A_O9EwWugZ5_2(.dout(w_dff_A_Ul0QIhXY5_2),.din(w_dff_A_O9EwWugZ5_2),.clk(gclk));
	jdff dff_A_dBm7to3B0_2(.dout(w_dff_A_O9EwWugZ5_2),.din(w_dff_A_dBm7to3B0_2),.clk(gclk));
	jdff dff_A_T7vBhMUj8_1(.dout(w_n612_0[1]),.din(w_dff_A_T7vBhMUj8_1),.clk(gclk));
	jdff dff_A_aK57UsaL5_1(.dout(w_dff_A_T7vBhMUj8_1),.din(w_dff_A_aK57UsaL5_1),.clk(gclk));
	jdff dff_A_9AWkHB5g3_1(.dout(w_dff_A_aK57UsaL5_1),.din(w_dff_A_9AWkHB5g3_1),.clk(gclk));
	jdff dff_A_olxTOttA6_1(.dout(w_dff_A_9AWkHB5g3_1),.din(w_dff_A_olxTOttA6_1),.clk(gclk));
	jdff dff_A_gtx9BhxV3_1(.dout(w_dff_A_olxTOttA6_1),.din(w_dff_A_gtx9BhxV3_1),.clk(gclk));
	jdff dff_A_BwpN446w0_1(.dout(w_dff_A_gtx9BhxV3_1),.din(w_dff_A_BwpN446w0_1),.clk(gclk));
	jdff dff_A_UZVNZD1m5_1(.dout(w_dff_A_BwpN446w0_1),.din(w_dff_A_UZVNZD1m5_1),.clk(gclk));
	jdff dff_A_MfMg31SE1_1(.dout(w_n146_1[1]),.din(w_dff_A_MfMg31SE1_1),.clk(gclk));
	jdff dff_A_KVSAQB6x9_1(.dout(w_dff_A_MfMg31SE1_1),.din(w_dff_A_KVSAQB6x9_1),.clk(gclk));
	jdff dff_A_wcuik72z9_1(.dout(w_dff_A_KVSAQB6x9_1),.din(w_dff_A_wcuik72z9_1),.clk(gclk));
	jdff dff_A_GWnmYwJh7_1(.dout(w_dff_A_wcuik72z9_1),.din(w_dff_A_GWnmYwJh7_1),.clk(gclk));
	jdff dff_A_lAyJxtep3_1(.dout(w_dff_A_GWnmYwJh7_1),.din(w_dff_A_lAyJxtep3_1),.clk(gclk));
	jdff dff_A_pyxeLgzK9_1(.dout(w_dff_A_lAyJxtep3_1),.din(w_dff_A_pyxeLgzK9_1),.clk(gclk));
	jdff dff_A_REnI5YUr6_2(.dout(w_n146_1[2]),.din(w_dff_A_REnI5YUr6_2),.clk(gclk));
	jdff dff_A_wCBDH8kw1_2(.dout(w_dff_A_REnI5YUr6_2),.din(w_dff_A_wCBDH8kw1_2),.clk(gclk));
	jdff dff_A_7cPEC6TA0_2(.dout(w_dff_A_wCBDH8kw1_2),.din(w_dff_A_7cPEC6TA0_2),.clk(gclk));
	jdff dff_A_Q2HUV31o5_2(.dout(w_dff_A_7cPEC6TA0_2),.din(w_dff_A_Q2HUV31o5_2),.clk(gclk));
	jdff dff_A_yCjTMs0C2_2(.dout(w_dff_A_Q2HUV31o5_2),.din(w_dff_A_yCjTMs0C2_2),.clk(gclk));
	jdff dff_A_o0x1YyjQ7_2(.dout(w_dff_A_yCjTMs0C2_2),.din(w_dff_A_o0x1YyjQ7_2),.clk(gclk));
	jdff dff_A_QFjLQ9A31_0(.dout(w_n425_1[0]),.din(w_dff_A_QFjLQ9A31_0),.clk(gclk));
	jdff dff_A_Qj78QzEa8_0(.dout(w_dff_A_QFjLQ9A31_0),.din(w_dff_A_Qj78QzEa8_0),.clk(gclk));
	jdff dff_A_yz5Me03f0_0(.dout(w_dff_A_Qj78QzEa8_0),.din(w_dff_A_yz5Me03f0_0),.clk(gclk));
	jdff dff_A_lo2DMc579_0(.dout(w_dff_A_yz5Me03f0_0),.din(w_dff_A_lo2DMc579_0),.clk(gclk));
	jdff dff_A_pZgIn6Mn2_0(.dout(w_dff_A_lo2DMc579_0),.din(w_dff_A_pZgIn6Mn2_0),.clk(gclk));
	jdff dff_A_9lcQDSgC5_0(.dout(w_dff_A_pZgIn6Mn2_0),.din(w_dff_A_9lcQDSgC5_0),.clk(gclk));
	jdff dff_A_Y3zWFNcr3_0(.dout(w_dff_A_9lcQDSgC5_0),.din(w_dff_A_Y3zWFNcr3_0),.clk(gclk));
	jdff dff_A_Q3jL4xQ95_0(.dout(w_dff_A_Y3zWFNcr3_0),.din(w_dff_A_Q3jL4xQ95_0),.clk(gclk));
	jdff dff_A_6y2D3p9b0_0(.dout(w_dff_A_Q3jL4xQ95_0),.din(w_dff_A_6y2D3p9b0_0),.clk(gclk));
	jdff dff_A_YLSA4Nci2_0(.dout(w_dff_A_6y2D3p9b0_0),.din(w_dff_A_YLSA4Nci2_0),.clk(gclk));
	jdff dff_A_qyCW8pT93_0(.dout(w_dff_A_YLSA4Nci2_0),.din(w_dff_A_qyCW8pT93_0),.clk(gclk));
	jdff dff_A_1rrweAxJ5_0(.dout(w_dff_A_qyCW8pT93_0),.din(w_dff_A_1rrweAxJ5_0),.clk(gclk));
	jdff dff_A_U1nsvXFK9_0(.dout(w_dff_A_1rrweAxJ5_0),.din(w_dff_A_U1nsvXFK9_0),.clk(gclk));
	jdff dff_A_QlUl0lp24_1(.dout(w_n425_1[1]),.din(w_dff_A_QlUl0lp24_1),.clk(gclk));
	jdff dff_A_bir5F7eH1_1(.dout(w_dff_A_QlUl0lp24_1),.din(w_dff_A_bir5F7eH1_1),.clk(gclk));
	jdff dff_A_5sMzEO2c4_1(.dout(w_dff_A_bir5F7eH1_1),.din(w_dff_A_5sMzEO2c4_1),.clk(gclk));
	jdff dff_A_EAuUh3eM7_1(.dout(w_dff_A_5sMzEO2c4_1),.din(w_dff_A_EAuUh3eM7_1),.clk(gclk));
	jdff dff_A_F2iBFrld3_1(.dout(w_dff_A_EAuUh3eM7_1),.din(w_dff_A_F2iBFrld3_1),.clk(gclk));
	jdff dff_A_sfCHYGZB6_1(.dout(w_dff_A_F2iBFrld3_1),.din(w_dff_A_sfCHYGZB6_1),.clk(gclk));
	jdff dff_A_HgWHZUp25_1(.dout(w_dff_A_sfCHYGZB6_1),.din(w_dff_A_HgWHZUp25_1),.clk(gclk));
	jdff dff_A_BbBgQ5tH3_1(.dout(w_dff_A_HgWHZUp25_1),.din(w_dff_A_BbBgQ5tH3_1),.clk(gclk));
	jdff dff_A_x4Ctfyb41_1(.dout(w_dff_A_BbBgQ5tH3_1),.din(w_dff_A_x4Ctfyb41_1),.clk(gclk));
	jdff dff_A_xW3tbapP7_1(.dout(w_dff_A_x4Ctfyb41_1),.din(w_dff_A_xW3tbapP7_1),.clk(gclk));
	jdff dff_A_EoSQQ67C1_1(.dout(w_dff_A_xW3tbapP7_1),.din(w_dff_A_EoSQQ67C1_1),.clk(gclk));
	jdff dff_A_frGaIkcL7_1(.dout(w_dff_A_EoSQQ67C1_1),.din(w_dff_A_frGaIkcL7_1),.clk(gclk));
	jdff dff_A_01HEKiPv4_1(.dout(w_dff_A_frGaIkcL7_1),.din(w_dff_A_01HEKiPv4_1),.clk(gclk));
	jdff dff_A_apbNwcZG3_1(.dout(w_n425_0[1]),.din(w_dff_A_apbNwcZG3_1),.clk(gclk));
	jdff dff_A_bnQIZaMM6_1(.dout(w_dff_A_apbNwcZG3_1),.din(w_dff_A_bnQIZaMM6_1),.clk(gclk));
	jdff dff_A_Iu4eF7L16_1(.dout(w_dff_A_bnQIZaMM6_1),.din(w_dff_A_Iu4eF7L16_1),.clk(gclk));
	jdff dff_A_gFnsGjdN1_1(.dout(w_dff_A_Iu4eF7L16_1),.din(w_dff_A_gFnsGjdN1_1),.clk(gclk));
	jdff dff_A_q46AWpcw8_1(.dout(w_dff_A_gFnsGjdN1_1),.din(w_dff_A_q46AWpcw8_1),.clk(gclk));
	jdff dff_A_MZzf122x5_1(.dout(w_dff_A_q46AWpcw8_1),.din(w_dff_A_MZzf122x5_1),.clk(gclk));
	jdff dff_A_3CMLQwKD1_1(.dout(w_dff_A_MZzf122x5_1),.din(w_dff_A_3CMLQwKD1_1),.clk(gclk));
	jdff dff_A_VmAgNmDG8_1(.dout(w_dff_A_3CMLQwKD1_1),.din(w_dff_A_VmAgNmDG8_1),.clk(gclk));
	jdff dff_A_fQNzXRoa0_1(.dout(w_dff_A_VmAgNmDG8_1),.din(w_dff_A_fQNzXRoa0_1),.clk(gclk));
	jdff dff_A_VYsKwuZb0_1(.dout(w_dff_A_fQNzXRoa0_1),.din(w_dff_A_VYsKwuZb0_1),.clk(gclk));
	jdff dff_A_xKz9M7fS3_1(.dout(w_dff_A_VYsKwuZb0_1),.din(w_dff_A_xKz9M7fS3_1),.clk(gclk));
	jdff dff_A_ubaIKEJ61_1(.dout(w_dff_A_xKz9M7fS3_1),.din(w_dff_A_ubaIKEJ61_1),.clk(gclk));
	jdff dff_A_juqvY5ge5_1(.dout(w_dff_A_ubaIKEJ61_1),.din(w_dff_A_juqvY5ge5_1),.clk(gclk));
	jdff dff_A_Ieevp0XE1_2(.dout(w_n425_0[2]),.din(w_dff_A_Ieevp0XE1_2),.clk(gclk));
	jdff dff_A_mcVKIyD40_2(.dout(w_dff_A_Ieevp0XE1_2),.din(w_dff_A_mcVKIyD40_2),.clk(gclk));
	jdff dff_A_CL60yoVR8_2(.dout(w_dff_A_mcVKIyD40_2),.din(w_dff_A_CL60yoVR8_2),.clk(gclk));
	jdff dff_A_5yu8exKE4_2(.dout(w_dff_A_CL60yoVR8_2),.din(w_dff_A_5yu8exKE4_2),.clk(gclk));
	jdff dff_A_Uv0Xm1Bb8_2(.dout(w_dff_A_5yu8exKE4_2),.din(w_dff_A_Uv0Xm1Bb8_2),.clk(gclk));
	jdff dff_A_SX3EYtG92_2(.dout(w_dff_A_Uv0Xm1Bb8_2),.din(w_dff_A_SX3EYtG92_2),.clk(gclk));
	jdff dff_A_gfvpNFiO8_2(.dout(w_dff_A_SX3EYtG92_2),.din(w_dff_A_gfvpNFiO8_2),.clk(gclk));
	jdff dff_A_7Y2f3YIX2_2(.dout(w_dff_A_gfvpNFiO8_2),.din(w_dff_A_7Y2f3YIX2_2),.clk(gclk));
	jdff dff_A_6vzYT7Q89_2(.dout(w_dff_A_7Y2f3YIX2_2),.din(w_dff_A_6vzYT7Q89_2),.clk(gclk));
	jdff dff_A_WXjVGyeo0_2(.dout(w_dff_A_6vzYT7Q89_2),.din(w_dff_A_WXjVGyeo0_2),.clk(gclk));
	jdff dff_A_icESleKK9_2(.dout(w_dff_A_WXjVGyeo0_2),.din(w_dff_A_icESleKK9_2),.clk(gclk));
	jdff dff_A_9mB63LIe3_2(.dout(w_dff_A_icESleKK9_2),.din(w_dff_A_9mB63LIe3_2),.clk(gclk));
	jdff dff_A_Srm5kXMA6_2(.dout(w_dff_A_9mB63LIe3_2),.din(w_dff_A_Srm5kXMA6_2),.clk(gclk));
	jdff dff_A_O64eRFnd9_0(.dout(w_n148_1[0]),.din(w_dff_A_O64eRFnd9_0),.clk(gclk));
	jdff dff_A_Zgm7zyNm4_0(.dout(w_dff_A_O64eRFnd9_0),.din(w_dff_A_Zgm7zyNm4_0),.clk(gclk));
	jdff dff_A_MY5eYnyZ8_0(.dout(w_dff_A_Zgm7zyNm4_0),.din(w_dff_A_MY5eYnyZ8_0),.clk(gclk));
	jdff dff_A_jQb7DLmM0_0(.dout(w_dff_A_MY5eYnyZ8_0),.din(w_dff_A_jQb7DLmM0_0),.clk(gclk));
	jdff dff_A_wbPRxEi36_1(.dout(w_n148_1[1]),.din(w_dff_A_wbPRxEi36_1),.clk(gclk));
	jdff dff_A_BYuIiKA37_1(.dout(w_dff_A_wbPRxEi36_1),.din(w_dff_A_BYuIiKA37_1),.clk(gclk));
	jdff dff_B_ToFRmcGQ2_0(.din(n701),.dout(w_dff_B_ToFRmcGQ2_0),.clk(gclk));
	jdff dff_A_2YbzKGby8_0(.dout(w_n604_1[0]),.din(w_dff_A_2YbzKGby8_0),.clk(gclk));
	jdff dff_A_i5Ds5bN29_0(.dout(w_dff_A_2YbzKGby8_0),.din(w_dff_A_i5Ds5bN29_0),.clk(gclk));
	jdff dff_A_F0VobcyN5_2(.dout(w_n604_1[2]),.din(w_dff_A_F0VobcyN5_2),.clk(gclk));
	jdff dff_A_vjNhp4wO4_2(.dout(w_dff_A_F0VobcyN5_2),.din(w_dff_A_vjNhp4wO4_2),.clk(gclk));
	jdff dff_A_f46lkmuH0_2(.dout(w_dff_A_vjNhp4wO4_2),.din(w_dff_A_f46lkmuH0_2),.clk(gclk));
	jdff dff_A_LupTeA0c5_2(.dout(w_dff_A_f46lkmuH0_2),.din(w_dff_A_LupTeA0c5_2),.clk(gclk));
	jdff dff_A_BkhVbplY0_2(.dout(w_dff_A_LupTeA0c5_2),.din(w_dff_A_BkhVbplY0_2),.clk(gclk));
	jdff dff_A_ZEPqOYZy9_2(.dout(w_dff_A_BkhVbplY0_2),.din(w_dff_A_ZEPqOYZy9_2),.clk(gclk));
	jdff dff_A_cf21gQDV6_2(.dout(w_dff_A_ZEPqOYZy9_2),.din(w_dff_A_cf21gQDV6_2),.clk(gclk));
	jdff dff_A_OSkJvifp7_2(.dout(w_dff_A_cf21gQDV6_2),.din(w_dff_A_OSkJvifp7_2),.clk(gclk));
	jdff dff_A_igeVjMAd9_0(.dout(w_n604_0[0]),.din(w_dff_A_igeVjMAd9_0),.clk(gclk));
	jdff dff_A_DHZW8wk15_0(.dout(w_dff_A_igeVjMAd9_0),.din(w_dff_A_DHZW8wk15_0),.clk(gclk));
	jdff dff_A_wM0pIoMX7_2(.dout(w_n604_0[2]),.din(w_dff_A_wM0pIoMX7_2),.clk(gclk));
	jdff dff_A_9f9VqMzN8_2(.dout(w_dff_A_wM0pIoMX7_2),.din(w_dff_A_9f9VqMzN8_2),.clk(gclk));
	jdff dff_A_RDucMg3G7_0(.dout(w_n603_2[0]),.din(w_dff_A_RDucMg3G7_0),.clk(gclk));
	jdff dff_A_8a8GQP3p1_0(.dout(w_dff_A_RDucMg3G7_0),.din(w_dff_A_8a8GQP3p1_0),.clk(gclk));
	jdff dff_A_ZHy6qTz98_0(.dout(w_dff_A_8a8GQP3p1_0),.din(w_dff_A_ZHy6qTz98_0),.clk(gclk));
	jdff dff_A_eGnqnVtQ8_0(.dout(w_dff_A_ZHy6qTz98_0),.din(w_dff_A_eGnqnVtQ8_0),.clk(gclk));
	jdff dff_A_MU4ralJA4_0(.dout(w_dff_A_eGnqnVtQ8_0),.din(w_dff_A_MU4ralJA4_0),.clk(gclk));
	jdff dff_A_xPo6llk43_0(.dout(w_dff_A_MU4ralJA4_0),.din(w_dff_A_xPo6llk43_0),.clk(gclk));
	jdff dff_A_sitLDePJ2_0(.dout(w_dff_A_xPo6llk43_0),.din(w_dff_A_sitLDePJ2_0),.clk(gclk));
	jdff dff_A_3HYZCYkx5_0(.dout(w_dff_A_sitLDePJ2_0),.din(w_dff_A_3HYZCYkx5_0),.clk(gclk));
	jdff dff_A_0a75YB7r5_0(.dout(w_dff_A_3HYZCYkx5_0),.din(w_dff_A_0a75YB7r5_0),.clk(gclk));
	jdff dff_A_yVn1imyF0_0(.dout(w_dff_A_0a75YB7r5_0),.din(w_dff_A_yVn1imyF0_0),.clk(gclk));
	jdff dff_A_UeTQRlg70_0(.dout(w_dff_A_yVn1imyF0_0),.din(w_dff_A_UeTQRlg70_0),.clk(gclk));
	jdff dff_A_qUiSdLMH8_0(.dout(w_n603_0[0]),.din(w_dff_A_qUiSdLMH8_0),.clk(gclk));
	jdff dff_A_fpbiBcSI7_0(.dout(w_dff_A_qUiSdLMH8_0),.din(w_dff_A_fpbiBcSI7_0),.clk(gclk));
	jdff dff_A_tKvRylP32_0(.dout(w_dff_A_fpbiBcSI7_0),.din(w_dff_A_tKvRylP32_0),.clk(gclk));
	jdff dff_A_QcUlEmmC5_0(.dout(w_dff_A_tKvRylP32_0),.din(w_dff_A_QcUlEmmC5_0),.clk(gclk));
	jdff dff_A_ExKlLBAI1_0(.dout(w_dff_A_QcUlEmmC5_0),.din(w_dff_A_ExKlLBAI1_0),.clk(gclk));
	jdff dff_A_3ntxPuHO3_0(.dout(w_dff_A_ExKlLBAI1_0),.din(w_dff_A_3ntxPuHO3_0),.clk(gclk));
	jdff dff_A_8TwwIrNO1_0(.dout(w_dff_A_3ntxPuHO3_0),.din(w_dff_A_8TwwIrNO1_0),.clk(gclk));
	jdff dff_A_XSZ6sDf47_0(.dout(w_dff_A_8TwwIrNO1_0),.din(w_dff_A_XSZ6sDf47_0),.clk(gclk));
	jdff dff_A_f96h5L4Q5_0(.dout(w_dff_A_XSZ6sDf47_0),.din(w_dff_A_f96h5L4Q5_0),.clk(gclk));
	jdff dff_A_hr5bMELX1_0(.dout(w_dff_A_f96h5L4Q5_0),.din(w_dff_A_hr5bMELX1_0),.clk(gclk));
	jdff dff_A_9B9zPNJo4_0(.dout(w_dff_A_hr5bMELX1_0),.din(w_dff_A_9B9zPNJo4_0),.clk(gclk));
	jdff dff_A_OnG5Egny5_0(.dout(w_dff_A_9B9zPNJo4_0),.din(w_dff_A_OnG5Egny5_0),.clk(gclk));
	jdff dff_A_67LEQ4PA8_0(.dout(w_dff_A_OnG5Egny5_0),.din(w_dff_A_67LEQ4PA8_0),.clk(gclk));
	jdff dff_A_4RRiHoEs0_0(.dout(w_dff_A_67LEQ4PA8_0),.din(w_dff_A_4RRiHoEs0_0),.clk(gclk));
	jdff dff_A_hrOe6sHs6_2(.dout(w_n603_0[2]),.din(w_dff_A_hrOe6sHs6_2),.clk(gclk));
	jdff dff_A_izinCztL5_2(.dout(w_dff_A_hrOe6sHs6_2),.din(w_dff_A_izinCztL5_2),.clk(gclk));
	jdff dff_A_dh3MLIUd3_2(.dout(w_dff_A_izinCztL5_2),.din(w_dff_A_dh3MLIUd3_2),.clk(gclk));
	jdff dff_A_mfRb8nQY3_2(.dout(w_dff_A_dh3MLIUd3_2),.din(w_dff_A_mfRb8nQY3_2),.clk(gclk));
	jdff dff_A_VqJR3Y8P5_2(.dout(w_dff_A_mfRb8nQY3_2),.din(w_dff_A_VqJR3Y8P5_2),.clk(gclk));
	jdff dff_A_NQkrsk995_2(.dout(w_dff_A_VqJR3Y8P5_2),.din(w_dff_A_NQkrsk995_2),.clk(gclk));
	jdff dff_A_h2SzWK0d5_2(.dout(w_dff_A_NQkrsk995_2),.din(w_dff_A_h2SzWK0d5_2),.clk(gclk));
	jdff dff_A_7cqMFiTh1_2(.dout(w_dff_A_h2SzWK0d5_2),.din(w_dff_A_7cqMFiTh1_2),.clk(gclk));
	jdff dff_A_4WHxmVZT4_2(.dout(w_dff_A_7cqMFiTh1_2),.din(w_dff_A_4WHxmVZT4_2),.clk(gclk));
	jdff dff_A_2RlqY59s8_2(.dout(w_dff_A_4WHxmVZT4_2),.din(w_dff_A_2RlqY59s8_2),.clk(gclk));
	jdff dff_A_dzuvx9Vi0_2(.dout(w_dff_A_2RlqY59s8_2),.din(w_dff_A_dzuvx9Vi0_2),.clk(gclk));
	jdff dff_A_2eAAhsCk3_2(.dout(w_dff_A_dzuvx9Vi0_2),.din(w_dff_A_2eAAhsCk3_2),.clk(gclk));
	jdff dff_A_NMzqwxXi2_2(.dout(w_dff_A_2eAAhsCk3_2),.din(w_dff_A_NMzqwxXi2_2),.clk(gclk));
	jdff dff_A_2KKKMxEO2_0(.dout(w_n602_0[0]),.din(w_dff_A_2KKKMxEO2_0),.clk(gclk));
	jdff dff_A_kklXdGwp8_0(.dout(w_dff_A_2KKKMxEO2_0),.din(w_dff_A_kklXdGwp8_0),.clk(gclk));
	jdff dff_A_kSUrakpl0_0(.dout(w_dff_A_kklXdGwp8_0),.din(w_dff_A_kSUrakpl0_0),.clk(gclk));
	jdff dff_A_Ze8pyVHu9_0(.dout(w_dff_A_kSUrakpl0_0),.din(w_dff_A_Ze8pyVHu9_0),.clk(gclk));
	jdff dff_A_Raxmyxn51_0(.dout(w_dff_A_Ze8pyVHu9_0),.din(w_dff_A_Raxmyxn51_0),.clk(gclk));
	jdff dff_A_uZI1uxxm9_0(.dout(w_dff_A_Raxmyxn51_0),.din(w_dff_A_uZI1uxxm9_0),.clk(gclk));
	jdff dff_A_00EfuHWr5_0(.dout(w_dff_A_uZI1uxxm9_0),.din(w_dff_A_00EfuHWr5_0),.clk(gclk));
	jdff dff_A_GMZfWSSF1_0(.dout(w_dff_A_00EfuHWr5_0),.din(w_dff_A_GMZfWSSF1_0),.clk(gclk));
	jdff dff_A_ZdbF9i3h5_0(.dout(w_dff_A_GMZfWSSF1_0),.din(w_dff_A_ZdbF9i3h5_0),.clk(gclk));
	jdff dff_A_TlThXpMa5_0(.dout(w_dff_A_ZdbF9i3h5_0),.din(w_dff_A_TlThXpMa5_0),.clk(gclk));
	jdff dff_A_IogcAiqi6_0(.dout(w_dff_A_TlThXpMa5_0),.din(w_dff_A_IogcAiqi6_0),.clk(gclk));
	jdff dff_A_KkVA1EWI4_0(.dout(w_dff_A_IogcAiqi6_0),.din(w_dff_A_KkVA1EWI4_0),.clk(gclk));
	jdff dff_A_xqHPYubh0_0(.dout(w_dff_A_KkVA1EWI4_0),.din(w_dff_A_xqHPYubh0_0),.clk(gclk));
	jdff dff_A_eZKsSnD04_0(.dout(w_dff_A_xqHPYubh0_0),.din(w_dff_A_eZKsSnD04_0),.clk(gclk));
	jdff dff_A_gETiBfap9_0(.dout(w_dff_A_eZKsSnD04_0),.din(w_dff_A_gETiBfap9_0),.clk(gclk));
	jdff dff_A_bqP0hXwQ1_0(.dout(w_dff_A_gETiBfap9_0),.din(w_dff_A_bqP0hXwQ1_0),.clk(gclk));
	jdff dff_A_hhWxJAtF1_0(.dout(w_dff_A_bqP0hXwQ1_0),.din(w_dff_A_hhWxJAtF1_0),.clk(gclk));
	jdff dff_A_qJzcbsiQ5_0(.dout(w_n592_0[0]),.din(w_dff_A_qJzcbsiQ5_0),.clk(gclk));
	jdff dff_A_fm3xRMa22_0(.dout(w_dff_A_qJzcbsiQ5_0),.din(w_dff_A_fm3xRMa22_0),.clk(gclk));
	jdff dff_A_Bzdl7SUk7_0(.dout(w_dff_A_fm3xRMa22_0),.din(w_dff_A_Bzdl7SUk7_0),.clk(gclk));
	jdff dff_A_60nDHZ7A3_0(.dout(w_dff_A_Bzdl7SUk7_0),.din(w_dff_A_60nDHZ7A3_0),.clk(gclk));
	jdff dff_A_r1a9DKN97_0(.dout(w_dff_A_60nDHZ7A3_0),.din(w_dff_A_r1a9DKN97_0),.clk(gclk));
	jdff dff_A_twgUN3sy1_0(.dout(w_dff_A_r1a9DKN97_0),.din(w_dff_A_twgUN3sy1_0),.clk(gclk));
	jdff dff_A_EjT8DoTg4_0(.dout(w_dff_A_twgUN3sy1_0),.din(w_dff_A_EjT8DoTg4_0),.clk(gclk));
	jdff dff_A_kC8sCidG6_0(.dout(w_dff_A_EjT8DoTg4_0),.din(w_dff_A_kC8sCidG6_0),.clk(gclk));
	jdff dff_A_4EBPQli13_0(.dout(w_dff_A_kC8sCidG6_0),.din(w_dff_A_4EBPQli13_0),.clk(gclk));
	jdff dff_A_w1Dw10HK4_0(.dout(w_dff_A_4EBPQli13_0),.din(w_dff_A_w1Dw10HK4_0),.clk(gclk));
	jdff dff_A_6X0v1u8U8_0(.dout(w_dff_A_w1Dw10HK4_0),.din(w_dff_A_6X0v1u8U8_0),.clk(gclk));
	jdff dff_A_8j4ASYBC0_0(.dout(w_dff_A_6X0v1u8U8_0),.din(w_dff_A_8j4ASYBC0_0),.clk(gclk));
	jdff dff_A_KNHB5mhX4_0(.dout(w_dff_A_8j4ASYBC0_0),.din(w_dff_A_KNHB5mhX4_0),.clk(gclk));
	jdff dff_A_tTRGCba08_2(.dout(w_n592_0[2]),.din(w_dff_A_tTRGCba08_2),.clk(gclk));
	jdff dff_A_9XtKLYwL2_2(.dout(w_dff_A_tTRGCba08_2),.din(w_dff_A_9XtKLYwL2_2),.clk(gclk));
	jdff dff_A_mVGq03yY8_2(.dout(w_dff_A_9XtKLYwL2_2),.din(w_dff_A_mVGq03yY8_2),.clk(gclk));
	jdff dff_A_l0g4ARMN5_2(.dout(w_dff_A_mVGq03yY8_2),.din(w_dff_A_l0g4ARMN5_2),.clk(gclk));
	jdff dff_A_v63deK9y4_2(.dout(w_dff_A_l0g4ARMN5_2),.din(w_dff_A_v63deK9y4_2),.clk(gclk));
	jdff dff_A_sNeVUY8j4_2(.dout(w_dff_A_v63deK9y4_2),.din(w_dff_A_sNeVUY8j4_2),.clk(gclk));
	jdff dff_A_g4AOfy8l0_2(.dout(w_dff_A_sNeVUY8j4_2),.din(w_dff_A_g4AOfy8l0_2),.clk(gclk));
	jdff dff_A_vzpxu5bz9_2(.dout(w_dff_A_g4AOfy8l0_2),.din(w_dff_A_vzpxu5bz9_2),.clk(gclk));
	jdff dff_A_zifp6hnE8_2(.dout(w_dff_A_vzpxu5bz9_2),.din(w_dff_A_zifp6hnE8_2),.clk(gclk));
	jdff dff_A_NM5hwlAr7_2(.dout(w_dff_A_zifp6hnE8_2),.din(w_dff_A_NM5hwlAr7_2),.clk(gclk));
	jdff dff_A_bKRGQ5hY0_2(.dout(w_dff_A_NM5hwlAr7_2),.din(w_dff_A_bKRGQ5hY0_2),.clk(gclk));
	jdff dff_A_3tXTZQie8_2(.dout(w_dff_A_bKRGQ5hY0_2),.din(w_dff_A_3tXTZQie8_2),.clk(gclk));
	jdff dff_A_8RFzvmkn8_2(.dout(w_dff_A_3tXTZQie8_2),.din(w_dff_A_8RFzvmkn8_2),.clk(gclk));
	jdff dff_A_ImjYv5sH8_2(.dout(w_dff_A_8RFzvmkn8_2),.din(w_dff_A_ImjYv5sH8_2),.clk(gclk));
	jdff dff_A_vEtMHDQE6_2(.dout(w_dff_A_ImjYv5sH8_2),.din(w_dff_A_vEtMHDQE6_2),.clk(gclk));
	jdff dff_A_pbO59dpv8_2(.dout(w_dff_A_vEtMHDQE6_2),.din(w_dff_A_pbO59dpv8_2),.clk(gclk));
	jdff dff_A_hXaqpHIU1_1(.dout(w_n591_0[1]),.din(w_dff_A_hXaqpHIU1_1),.clk(gclk));
	jdff dff_A_q6PhK3IL6_1(.dout(w_dff_A_hXaqpHIU1_1),.din(w_dff_A_q6PhK3IL6_1),.clk(gclk));
	jdff dff_A_5XEw9YYy7_1(.dout(w_dff_A_q6PhK3IL6_1),.din(w_dff_A_5XEw9YYy7_1),.clk(gclk));
	jdff dff_A_ZuZ08gKE8_1(.dout(w_dff_A_5XEw9YYy7_1),.din(w_dff_A_ZuZ08gKE8_1),.clk(gclk));
	jdff dff_A_QVJ07exF8_1(.dout(w_dff_A_ZuZ08gKE8_1),.din(w_dff_A_QVJ07exF8_1),.clk(gclk));
	jdff dff_A_0oqXYBeD5_1(.dout(w_dff_A_QVJ07exF8_1),.din(w_dff_A_0oqXYBeD5_1),.clk(gclk));
	jdff dff_A_5QKhZG5x9_1(.dout(w_dff_A_0oqXYBeD5_1),.din(w_dff_A_5QKhZG5x9_1),.clk(gclk));
	jdff dff_A_rbymtoR63_1(.dout(w_dff_A_5QKhZG5x9_1),.din(w_dff_A_rbymtoR63_1),.clk(gclk));
	jdff dff_A_aVB2aesx0_1(.dout(w_dff_A_rbymtoR63_1),.din(w_dff_A_aVB2aesx0_1),.clk(gclk));
	jdff dff_A_S5mYsdfC6_1(.dout(w_dff_A_aVB2aesx0_1),.din(w_dff_A_S5mYsdfC6_1),.clk(gclk));
	jdff dff_A_kzp80mkF1_1(.dout(w_dff_A_S5mYsdfC6_1),.din(w_dff_A_kzp80mkF1_1),.clk(gclk));
	jdff dff_A_ekH6s8rA2_1(.dout(w_dff_A_kzp80mkF1_1),.din(w_dff_A_ekH6s8rA2_1),.clk(gclk));
	jdff dff_A_7UXBHXrr8_1(.dout(w_dff_A_ekH6s8rA2_1),.din(w_dff_A_7UXBHXrr8_1),.clk(gclk));
	jdff dff_A_hMqIvqxr9_1(.dout(w_dff_A_7UXBHXrr8_1),.din(w_dff_A_hMqIvqxr9_1),.clk(gclk));
	jdff dff_A_P99KkVrv0_1(.dout(w_dff_A_hMqIvqxr9_1),.din(w_dff_A_P99KkVrv0_1),.clk(gclk));
	jdff dff_A_QdsBB7La3_2(.dout(w_n591_0[2]),.din(w_dff_A_QdsBB7La3_2),.clk(gclk));
	jdff dff_A_USn8cusi8_2(.dout(w_dff_A_QdsBB7La3_2),.din(w_dff_A_USn8cusi8_2),.clk(gclk));
	jdff dff_A_aIuZPe2o1_2(.dout(w_dff_A_USn8cusi8_2),.din(w_dff_A_aIuZPe2o1_2),.clk(gclk));
	jdff dff_A_mH5eGrmt9_2(.dout(w_dff_A_aIuZPe2o1_2),.din(w_dff_A_mH5eGrmt9_2),.clk(gclk));
	jdff dff_A_319wHlOC7_2(.dout(w_dff_A_mH5eGrmt9_2),.din(w_dff_A_319wHlOC7_2),.clk(gclk));
	jdff dff_A_dz3mmXd33_2(.dout(w_dff_A_319wHlOC7_2),.din(w_dff_A_dz3mmXd33_2),.clk(gclk));
	jdff dff_A_vDtdNpEu0_2(.dout(w_dff_A_dz3mmXd33_2),.din(w_dff_A_vDtdNpEu0_2),.clk(gclk));
	jdff dff_A_msf1W9BA9_2(.dout(w_dff_A_vDtdNpEu0_2),.din(w_dff_A_msf1W9BA9_2),.clk(gclk));
	jdff dff_A_gEkg5rZd3_2(.dout(w_dff_A_msf1W9BA9_2),.din(w_dff_A_gEkg5rZd3_2),.clk(gclk));
	jdff dff_A_hcecLVZx0_2(.dout(w_dff_A_gEkg5rZd3_2),.din(w_dff_A_hcecLVZx0_2),.clk(gclk));
	jdff dff_A_J7f9aLGS7_2(.dout(w_dff_A_hcecLVZx0_2),.din(w_dff_A_J7f9aLGS7_2),.clk(gclk));
	jdff dff_A_FFiuvnBX3_2(.dout(w_dff_A_J7f9aLGS7_2),.din(w_dff_A_FFiuvnBX3_2),.clk(gclk));
	jdff dff_A_OcLCl1li7_2(.dout(w_dff_A_FFiuvnBX3_2),.din(w_dff_A_OcLCl1li7_2),.clk(gclk));
	jdff dff_A_wOa8UGtJ2_2(.dout(w_dff_A_OcLCl1li7_2),.din(w_dff_A_wOa8UGtJ2_2),.clk(gclk));
	jdff dff_A_7Mf11hn86_2(.dout(w_dff_A_wOa8UGtJ2_2),.din(w_dff_A_7Mf11hn86_2),.clk(gclk));
	jdff dff_A_9oa9JSFi3_2(.dout(w_dff_A_7Mf11hn86_2),.din(w_dff_A_9oa9JSFi3_2),.clk(gclk));
	jdff dff_A_o8jC3wy89_0(.dout(w_n121_0[0]),.din(w_dff_A_o8jC3wy89_0),.clk(gclk));
	jdff dff_B_q5AGVv120_1(.din(n690),.dout(w_dff_B_q5AGVv120_1),.clk(gclk));
	jdff dff_A_FCrx7MFn5_0(.dout(w_n696_1[0]),.din(w_dff_A_FCrx7MFn5_0),.clk(gclk));
	jdff dff_A_LzAARKpC1_2(.dout(w_n696_1[2]),.din(w_dff_A_LzAARKpC1_2),.clk(gclk));
	jdff dff_A_TBk7QCdd1_1(.dout(w_n696_0[1]),.din(w_dff_A_TBk7QCdd1_1),.clk(gclk));
	jdff dff_A_Im8C63OO4_1(.dout(w_n692_0[1]),.din(w_dff_A_Im8C63OO4_1),.clk(gclk));
	jdff dff_B_cMsoc7sh1_2(.din(n692),.dout(w_dff_B_cMsoc7sh1_2),.clk(gclk));
	jdff dff_B_0IyZh3r87_1(.din(n406),.dout(w_dff_B_0IyZh3r87_1),.clk(gclk));
	jdff dff_B_Ja2zN20d8_1(.din(w_dff_B_0IyZh3r87_1),.dout(w_dff_B_Ja2zN20d8_1),.clk(gclk));
	jdff dff_A_QPOjnUF42_1(.dout(w_n407_0[1]),.din(w_dff_A_QPOjnUF42_1),.clk(gclk));
	jdff dff_A_CiMjb1I22_1(.dout(w_dff_A_QPOjnUF42_1),.din(w_dff_A_CiMjb1I22_1),.clk(gclk));
	jdff dff_A_e41t7c4X0_1(.dout(w_dff_A_CiMjb1I22_1),.din(w_dff_A_e41t7c4X0_1),.clk(gclk));
	jdff dff_A_fRyBsshg1_1(.dout(w_dff_A_e41t7c4X0_1),.din(w_dff_A_fRyBsshg1_1),.clk(gclk));
	jdff dff_A_RGq7ptNu3_1(.dout(w_dff_A_fRyBsshg1_1),.din(w_dff_A_RGq7ptNu3_1),.clk(gclk));
	jdff dff_A_rM0bwNhF2_1(.dout(w_dff_A_RGq7ptNu3_1),.din(w_dff_A_rM0bwNhF2_1),.clk(gclk));
	jdff dff_A_iI3BAws32_2(.dout(w_n407_0[2]),.din(w_dff_A_iI3BAws32_2),.clk(gclk));
	jdff dff_A_NuGbAMwL1_1(.dout(w_n401_0[1]),.din(w_dff_A_NuGbAMwL1_1),.clk(gclk));
	jdff dff_B_ZH0hIGre5_1(.din(n396),.dout(w_dff_B_ZH0hIGre5_1),.clk(gclk));
	jdff dff_B_w8aVsJPu0_1(.din(w_dff_B_ZH0hIGre5_1),.dout(w_dff_B_w8aVsJPu0_1),.clk(gclk));
	jdff dff_B_7aS6B6hN6_1(.din(n397),.dout(w_dff_B_7aS6B6hN6_1),.clk(gclk));
	jdff dff_B_dP8ERMqf7_1(.din(w_dff_B_7aS6B6hN6_1),.dout(w_dff_B_dP8ERMqf7_1),.clk(gclk));
	jdff dff_B_AFu2vZVl4_0(.din(n398),.dout(w_dff_B_AFu2vZVl4_0),.clk(gclk));
	jdff dff_B_7Nb557uG9_0(.din(w_dff_B_AFu2vZVl4_0),.dout(w_dff_B_7Nb557uG9_0),.clk(gclk));
	jdff dff_A_FZiDhw6C1_1(.dout(w_n72_0[1]),.din(w_dff_A_FZiDhw6C1_1),.clk(gclk));
	jdff dff_A_GqESV7yA9_1(.dout(w_dff_A_FZiDhw6C1_1),.din(w_dff_A_GqESV7yA9_1),.clk(gclk));
	jdff dff_A_S2bmOonB3_1(.dout(w_dff_A_GqESV7yA9_1),.din(w_dff_A_S2bmOonB3_1),.clk(gclk));
	jdff dff_A_vLREaknN6_2(.dout(w_n72_0[2]),.din(w_dff_A_vLREaknN6_2),.clk(gclk));
	jdff dff_A_FKNrCzj53_2(.dout(w_dff_A_vLREaknN6_2),.din(w_dff_A_FKNrCzj53_2),.clk(gclk));
	jdff dff_B_I3nt5hgZ5_0(.din(n394),.dout(w_dff_B_I3nt5hgZ5_0),.clk(gclk));
	jdff dff_A_xzFq9UPv6_0(.dout(w_n112_3[0]),.din(w_dff_A_xzFq9UPv6_0),.clk(gclk));
	jdff dff_A_XCiI2xG81_0(.dout(w_dff_A_xzFq9UPv6_0),.din(w_dff_A_XCiI2xG81_0),.clk(gclk));
	jdff dff_A_i59xcJY51_1(.dout(w_n112_3[1]),.din(w_dff_A_i59xcJY51_1),.clk(gclk));
	jdff dff_A_63v7l7Vq9_1(.dout(w_dff_A_i59xcJY51_1),.din(w_dff_A_63v7l7Vq9_1),.clk(gclk));
	jdff dff_A_QWWqCtkg0_0(.dout(w_G58_4[0]),.din(w_dff_A_QWWqCtkg0_0),.clk(gclk));
	jdff dff_A_Mjh3b7UO7_1(.dout(w_G58_4[1]),.din(w_dff_A_Mjh3b7UO7_1),.clk(gclk));
	jdff dff_A_6m0bHzbb6_0(.dout(w_G58_1[0]),.din(w_dff_A_6m0bHzbb6_0),.clk(gclk));
	jdff dff_A_PrZhEze71_2(.dout(w_G58_1[2]),.din(w_dff_A_PrZhEze71_2),.clk(gclk));
	jdff dff_A_Xg3pnDtJ4_2(.dout(w_dff_A_PrZhEze71_2),.din(w_dff_A_Xg3pnDtJ4_2),.clk(gclk));
	jdff dff_A_BtUpt0110_2(.dout(w_dff_A_Xg3pnDtJ4_2),.din(w_dff_A_BtUpt0110_2),.clk(gclk));
	jdff dff_A_pR8uKgO07_2(.dout(w_dff_A_BtUpt0110_2),.din(w_dff_A_pR8uKgO07_2),.clk(gclk));
	jdff dff_A_i85muIC40_1(.dout(w_G58_0[1]),.din(w_dff_A_i85muIC40_1),.clk(gclk));
	jdff dff_A_vHIhuok02_2(.dout(w_G58_0[2]),.din(w_dff_A_vHIhuok02_2),.clk(gclk));
	jdff dff_A_V3pXokVU0_2(.dout(w_dff_A_vHIhuok02_2),.din(w_dff_A_V3pXokVU0_2),.clk(gclk));
	jdff dff_A_cxfkScNB3_2(.dout(w_dff_A_V3pXokVU0_2),.din(w_dff_A_cxfkScNB3_2),.clk(gclk));
	jdff dff_A_Jgno6nkh7_1(.dout(w_G20_3[1]),.din(w_dff_A_Jgno6nkh7_1),.clk(gclk));
	jdff dff_A_igQewKez1_2(.dout(w_G20_3[2]),.din(w_dff_A_igQewKez1_2),.clk(gclk));
	jdff dff_A_7sF9HlrM6_2(.dout(w_dff_A_igQewKez1_2),.din(w_dff_A_7sF9HlrM6_2),.clk(gclk));
	jdff dff_B_NU60nkyg4_2(.din(n390),.dout(w_dff_B_NU60nkyg4_2),.clk(gclk));
	jdff dff_B_MPLAYylK2_2(.din(w_dff_B_NU60nkyg4_2),.dout(w_dff_B_MPLAYylK2_2),.clk(gclk));
	jdff dff_A_yVgeO5789_0(.dout(w_G87_2[0]),.din(w_dff_A_yVgeO5789_0),.clk(gclk));
	jdff dff_A_F2nHkO901_0(.dout(w_dff_A_yVgeO5789_0),.din(w_dff_A_F2nHkO901_0),.clk(gclk));
	jdff dff_A_pZJDfEC69_0(.dout(w_dff_A_F2nHkO901_0),.din(w_dff_A_pZJDfEC69_0),.clk(gclk));
	jdff dff_A_aVsadp7V2_0(.dout(w_dff_A_pZJDfEC69_0),.din(w_dff_A_aVsadp7V2_0),.clk(gclk));
	jdff dff_A_470PHLTQ0_1(.dout(w_G87_2[1]),.din(w_dff_A_470PHLTQ0_1),.clk(gclk));
	jdff dff_A_qq2etdfU1_1(.dout(w_dff_A_470PHLTQ0_1),.din(w_dff_A_qq2etdfU1_1),.clk(gclk));
	jdff dff_A_wcSOMHkc7_1(.dout(w_dff_A_qq2etdfU1_1),.din(w_dff_A_wcSOMHkc7_1),.clk(gclk));
	jdff dff_A_rGYIVoJs5_1(.dout(w_dff_A_wcSOMHkc7_1),.din(w_dff_A_rGYIVoJs5_1),.clk(gclk));
	jdff dff_A_UY8yXUs39_1(.dout(w_n149_1[1]),.din(w_dff_A_UY8yXUs39_1),.clk(gclk));
	jdff dff_A_nhFB6Wdy6_1(.dout(w_dff_A_UY8yXUs39_1),.din(w_dff_A_nhFB6Wdy6_1),.clk(gclk));
	jdff dff_B_v9vq1SUv1_1(.din(n375),.dout(w_dff_B_v9vq1SUv1_1),.clk(gclk));
	jdff dff_A_qLHi8o0E6_0(.dout(w_G232_1[0]),.din(w_dff_A_qLHi8o0E6_0),.clk(gclk));
	jdff dff_A_2sF6EAVe2_0(.dout(w_dff_A_qLHi8o0E6_0),.din(w_dff_A_2sF6EAVe2_0),.clk(gclk));
	jdff dff_A_lwoF2VS19_1(.dout(w_G232_1[1]),.din(w_dff_A_lwoF2VS19_1),.clk(gclk));
	jdff dff_A_3fRE8kKZ3_1(.dout(w_G232_0[1]),.din(w_dff_A_3fRE8kKZ3_1),.clk(gclk));
	jdff dff_A_PDBLOkoQ0_1(.dout(w_dff_A_3fRE8kKZ3_1),.din(w_dff_A_PDBLOkoQ0_1),.clk(gclk));
	jdff dff_A_rwJfIo3F3_1(.dout(w_dff_A_PDBLOkoQ0_1),.din(w_dff_A_rwJfIo3F3_1),.clk(gclk));
	jdff dff_A_CZISefcV8_1(.dout(w_dff_A_rwJfIo3F3_1),.din(w_dff_A_CZISefcV8_1),.clk(gclk));
	jdff dff_A_dfXod0py9_2(.dout(w_G232_0[2]),.din(w_dff_A_dfXod0py9_2),.clk(gclk));
	jdff dff_A_wZ3zF3iC5_2(.dout(w_dff_A_dfXod0py9_2),.din(w_dff_A_wZ3zF3iC5_2),.clk(gclk));
	jdff dff_B_Yea19fe24_0(.din(n538),.dout(w_dff_B_Yea19fe24_0),.clk(gclk));
	jdff dff_A_lrS1MQPf1_1(.dout(w_n532_0[1]),.din(w_dff_A_lrS1MQPf1_1),.clk(gclk));
	jdff dff_B_LzLWH8KM7_1(.din(n525),.dout(w_dff_B_LzLWH8KM7_1),.clk(gclk));
	jdff dff_A_IHmCwTyd5_1(.dout(w_n524_0[1]),.din(w_dff_A_IHmCwTyd5_1),.clk(gclk));
	jdff dff_A_Uky4l53N4_0(.dout(w_n523_0[0]),.din(w_dff_A_Uky4l53N4_0),.clk(gclk));
	jdff dff_A_AdDCGg8T0_2(.dout(w_n588_0[2]),.din(w_dff_A_AdDCGg8T0_2),.clk(gclk));
	jdff dff_A_ufRxWv6b1_2(.dout(w_dff_A_AdDCGg8T0_2),.din(w_dff_A_ufRxWv6b1_2),.clk(gclk));
	jdff dff_B_Ao6zYikO0_0(.din(n587),.dout(w_dff_B_Ao6zYikO0_0),.clk(gclk));
	jdff dff_B_2iHUmqcd2_1(.din(n580),.dout(w_dff_B_2iHUmqcd2_1),.clk(gclk));
	jdff dff_B_KdKHTE9v4_1(.din(n581),.dout(w_dff_B_KdKHTE9v4_1),.clk(gclk));
	jdff dff_A_bXVRJXjo6_1(.dout(w_n554_2[1]),.din(w_dff_A_bXVRJXjo6_1),.clk(gclk));
	jdff dff_A_lE9FDNoY9_2(.dout(w_n554_2[2]),.din(w_dff_A_lE9FDNoY9_2),.clk(gclk));
	jdff dff_A_SsxPyY0o6_2(.dout(w_dff_A_lE9FDNoY9_2),.din(w_dff_A_SsxPyY0o6_2),.clk(gclk));
	jdff dff_A_5zizEvxm1_2(.dout(w_dff_A_SsxPyY0o6_2),.din(w_dff_A_5zizEvxm1_2),.clk(gclk));
	jdff dff_A_irrr2R7R5_2(.dout(w_dff_A_5zizEvxm1_2),.din(w_dff_A_irrr2R7R5_2),.clk(gclk));
	jdff dff_A_4iVzRieL8_2(.dout(w_dff_A_irrr2R7R5_2),.din(w_dff_A_4iVzRieL8_2),.clk(gclk));
	jdff dff_A_NINKWWWh6_0(.dout(w_n554_0[0]),.din(w_dff_A_NINKWWWh6_0),.clk(gclk));
	jdff dff_A_3ISqDeBM3_0(.dout(w_dff_A_NINKWWWh6_0),.din(w_dff_A_3ISqDeBM3_0),.clk(gclk));
	jdff dff_A_P8mMtLYv0_0(.dout(w_dff_A_3ISqDeBM3_0),.din(w_dff_A_P8mMtLYv0_0),.clk(gclk));
	jdff dff_A_jwSb8tfs3_1(.dout(w_n554_0[1]),.din(w_dff_A_jwSb8tfs3_1),.clk(gclk));
	jdff dff_A_hMeOEyx59_1(.dout(w_dff_A_jwSb8tfs3_1),.din(w_dff_A_hMeOEyx59_1),.clk(gclk));
	jdff dff_B_URPYmcRE4_3(.din(n554),.dout(w_dff_B_URPYmcRE4_3),.clk(gclk));
	jdff dff_B_4euaslRD6_3(.din(w_dff_B_URPYmcRE4_3),.dout(w_dff_B_4euaslRD6_3),.clk(gclk));
	jdff dff_A_Ym3uFM6E0_0(.dout(w_n534_0[0]),.din(w_dff_A_Ym3uFM6E0_0),.clk(gclk));
	jdff dff_A_t7bUeRsk7_0(.dout(w_G330_0[0]),.din(w_dff_A_t7bUeRsk7_0),.clk(gclk));
	jdff dff_A_xJcSlXtV9_0(.dout(w_dff_A_t7bUeRsk7_0),.din(w_dff_A_xJcSlXtV9_0),.clk(gclk));
	jdff dff_A_QZyOovr08_0(.dout(w_dff_A_xJcSlXtV9_0),.din(w_dff_A_QZyOovr08_0),.clk(gclk));
	jdff dff_A_Nai817tk0_0(.dout(w_dff_A_QZyOovr08_0),.din(w_dff_A_Nai817tk0_0),.clk(gclk));
	jdff dff_A_Ai49wWVh2_0(.dout(w_dff_A_Nai817tk0_0),.din(w_dff_A_Ai49wWVh2_0),.clk(gclk));
	jdff dff_A_Vbndpgai8_0(.dout(w_dff_A_Ai49wWVh2_0),.din(w_dff_A_Vbndpgai8_0),.clk(gclk));
	jdff dff_A_pl2QGNfM2_0(.dout(w_dff_A_Vbndpgai8_0),.din(w_dff_A_pl2QGNfM2_0),.clk(gclk));
	jdff dff_A_e30Kr4GF0_0(.dout(w_dff_A_pl2QGNfM2_0),.din(w_dff_A_e30Kr4GF0_0),.clk(gclk));
	jdff dff_A_dozsGobe8_0(.dout(w_dff_A_e30Kr4GF0_0),.din(w_dff_A_dozsGobe8_0),.clk(gclk));
	jdff dff_A_0JOd5oEu3_0(.dout(w_dff_A_dozsGobe8_0),.din(w_dff_A_0JOd5oEu3_0),.clk(gclk));
	jdff dff_A_L9d9XzyQ5_0(.dout(w_dff_A_0JOd5oEu3_0),.din(w_dff_A_L9d9XzyQ5_0),.clk(gclk));
	jdff dff_A_slHywqOc0_0(.dout(w_dff_A_L9d9XzyQ5_0),.din(w_dff_A_slHywqOc0_0),.clk(gclk));
	jdff dff_A_FGocdD9N7_0(.dout(w_n553_2[0]),.din(w_dff_A_FGocdD9N7_0),.clk(gclk));
	jdff dff_A_A7wXq5rE3_0(.dout(w_dff_A_FGocdD9N7_0),.din(w_dff_A_A7wXq5rE3_0),.clk(gclk));
	jdff dff_A_D6sZjnq76_0(.dout(w_dff_A_A7wXq5rE3_0),.din(w_dff_A_D6sZjnq76_0),.clk(gclk));
	jdff dff_A_3cS0A53x5_0(.dout(w_dff_A_D6sZjnq76_0),.din(w_dff_A_3cS0A53x5_0),.clk(gclk));
	jdff dff_A_26Dzk5OR2_0(.dout(w_dff_A_3cS0A53x5_0),.din(w_dff_A_26Dzk5OR2_0),.clk(gclk));
	jdff dff_A_82IQy6tX3_0(.dout(w_dff_A_26Dzk5OR2_0),.din(w_dff_A_82IQy6tX3_0),.clk(gclk));
	jdff dff_A_96QSHZBZ9_0(.dout(w_dff_A_82IQy6tX3_0),.din(w_dff_A_96QSHZBZ9_0),.clk(gclk));
	jdff dff_A_XTPuqfGv3_0(.dout(w_dff_A_96QSHZBZ9_0),.din(w_dff_A_XTPuqfGv3_0),.clk(gclk));
	jdff dff_A_1IoTyaGF1_0(.dout(w_dff_A_XTPuqfGv3_0),.din(w_dff_A_1IoTyaGF1_0),.clk(gclk));
	jdff dff_A_cuxQ11mA4_1(.dout(w_n553_2[1]),.din(w_dff_A_cuxQ11mA4_1),.clk(gclk));
	jdff dff_A_fLATu3s21_1(.dout(w_dff_A_cuxQ11mA4_1),.din(w_dff_A_fLATu3s21_1),.clk(gclk));
	jdff dff_A_I1W9SNlC3_1(.dout(w_dff_A_fLATu3s21_1),.din(w_dff_A_I1W9SNlC3_1),.clk(gclk));
	jdff dff_A_LpwxVUGw7_1(.dout(w_dff_A_I1W9SNlC3_1),.din(w_dff_A_LpwxVUGw7_1),.clk(gclk));
	jdff dff_A_SgKpglzj9_1(.dout(w_dff_A_LpwxVUGw7_1),.din(w_dff_A_SgKpglzj9_1),.clk(gclk));
	jdff dff_A_qcuyOwu73_0(.dout(w_n553_0[0]),.din(w_dff_A_qcuyOwu73_0),.clk(gclk));
	jdff dff_A_Nzq8A0ba9_0(.dout(w_dff_A_qcuyOwu73_0),.din(w_dff_A_Nzq8A0ba9_0),.clk(gclk));
	jdff dff_A_oRBHHkxw3_0(.dout(w_dff_A_Nzq8A0ba9_0),.din(w_dff_A_oRBHHkxw3_0),.clk(gclk));
	jdff dff_A_TEJfY3zX3_0(.dout(w_dff_A_oRBHHkxw3_0),.din(w_dff_A_TEJfY3zX3_0),.clk(gclk));
	jdff dff_A_0yt1rV2I1_2(.dout(w_n553_0[2]),.din(w_dff_A_0yt1rV2I1_2),.clk(gclk));
	jdff dff_A_sejDLEvb2_2(.dout(w_dff_A_0yt1rV2I1_2),.din(w_dff_A_sejDLEvb2_2),.clk(gclk));
	jdff dff_A_jReJ0Rc02_2(.dout(w_dff_A_sejDLEvb2_2),.din(w_dff_A_jReJ0Rc02_2),.clk(gclk));
	jdff dff_A_KbtCw2Be9_2(.dout(w_dff_A_jReJ0Rc02_2),.din(w_dff_A_KbtCw2Be9_2),.clk(gclk));
	jdff dff_A_uDb9li524_2(.dout(w_dff_A_KbtCw2Be9_2),.din(w_dff_A_uDb9li524_2),.clk(gclk));
	jdff dff_A_sHrhhkQJ2_2(.dout(w_dff_A_uDb9li524_2),.din(w_dff_A_sHrhhkQJ2_2),.clk(gclk));
	jdff dff_A_CL3hdu101_1(.dout(w_n552_0[1]),.din(w_dff_A_CL3hdu101_1),.clk(gclk));
	jdff dff_A_Uzp6K9k27_1(.dout(w_dff_A_CL3hdu101_1),.din(w_dff_A_Uzp6K9k27_1),.clk(gclk));
	jdff dff_A_ghBuExEe4_1(.dout(w_dff_A_Uzp6K9k27_1),.din(w_dff_A_ghBuExEe4_1),.clk(gclk));
	jdff dff_A_P1pQTy2S6_1(.dout(w_dff_A_ghBuExEe4_1),.din(w_dff_A_P1pQTy2S6_1),.clk(gclk));
	jdff dff_A_GfNU974E0_1(.dout(w_dff_A_P1pQTy2S6_1),.din(w_dff_A_GfNU974E0_1),.clk(gclk));
	jdff dff_A_G0TcI57k1_1(.dout(w_dff_A_GfNU974E0_1),.din(w_dff_A_G0TcI57k1_1),.clk(gclk));
	jdff dff_A_YGVxfLki0_1(.dout(w_dff_A_G0TcI57k1_1),.din(w_dff_A_YGVxfLki0_1),.clk(gclk));
	jdff dff_A_VlSN2j3M8_2(.dout(w_n552_0[2]),.din(w_dff_A_VlSN2j3M8_2),.clk(gclk));
	jdff dff_A_T0u8ZC016_2(.dout(w_dff_A_VlSN2j3M8_2),.din(w_dff_A_T0u8ZC016_2),.clk(gclk));
	jdff dff_A_qZ6PRYIe3_2(.dout(w_dff_A_T0u8ZC016_2),.din(w_dff_A_qZ6PRYIe3_2),.clk(gclk));
	jdff dff_A_wYlX2dmG9_2(.dout(w_dff_A_qZ6PRYIe3_2),.din(w_dff_A_wYlX2dmG9_2),.clk(gclk));
	jdff dff_A_KOyNZY7v0_2(.dout(w_dff_A_wYlX2dmG9_2),.din(w_dff_A_KOyNZY7v0_2),.clk(gclk));
	jdff dff_A_c7UUtwWp8_2(.dout(w_dff_A_KOyNZY7v0_2),.din(w_dff_A_c7UUtwWp8_2),.clk(gclk));
	jdff dff_A_q1KHmSbO4_2(.dout(w_dff_A_c7UUtwWp8_2),.din(w_dff_A_q1KHmSbO4_2),.clk(gclk));
	jdff dff_A_nj5ryxbi9_0(.dout(w_G213_0[0]),.din(w_dff_A_nj5ryxbi9_0),.clk(gclk));
	jdff dff_A_06UoBpWW4_2(.dout(w_G213_0[2]),.din(w_dff_A_06UoBpWW4_2),.clk(gclk));
	jdff dff_A_G2iJTLxm5_0(.dout(w_n113_1[0]),.din(w_dff_A_G2iJTLxm5_0),.clk(gclk));
	jdff dff_A_CoFQTjdU4_0(.dout(w_dff_A_G2iJTLxm5_0),.din(w_dff_A_CoFQTjdU4_0),.clk(gclk));
	jdff dff_A_0FsblvdM4_1(.dout(w_n113_1[1]),.din(w_dff_A_0FsblvdM4_1),.clk(gclk));
	jdff dff_A_awiYCCAm5_1(.dout(w_dff_A_0FsblvdM4_1),.din(w_dff_A_awiYCCAm5_1),.clk(gclk));
	jdff dff_A_DvqUdaea1_1(.dout(w_dff_A_awiYCCAm5_1),.din(w_dff_A_DvqUdaea1_1),.clk(gclk));
	jdff dff_A_IVfs17j22_1(.dout(w_dff_A_DvqUdaea1_1),.din(w_dff_A_IVfs17j22_1),.clk(gclk));
	jdff dff_A_L7dgG65K4_1(.dout(w_dff_A_IVfs17j22_1),.din(w_dff_A_L7dgG65K4_1),.clk(gclk));
	jdff dff_A_yESD0x6O4_1(.dout(w_dff_A_L7dgG65K4_1),.din(w_dff_A_yESD0x6O4_1),.clk(gclk));
	jdff dff_A_275NIoSS5_1(.dout(w_dff_A_yESD0x6O4_1),.din(w_dff_A_275NIoSS5_1),.clk(gclk));
	jdff dff_A_rhmi6y775_1(.dout(w_dff_A_275NIoSS5_1),.din(w_dff_A_rhmi6y775_1),.clk(gclk));
	jdff dff_A_Ihnghm883_1(.dout(w_dff_A_rhmi6y775_1),.din(w_dff_A_Ihnghm883_1),.clk(gclk));
	jdff dff_A_sjoCCasm5_1(.dout(w_dff_A_Ihnghm883_1),.din(w_dff_A_sjoCCasm5_1),.clk(gclk));
	jdff dff_A_Q7ura78J7_1(.dout(w_dff_A_sjoCCasm5_1),.din(w_dff_A_Q7ura78J7_1),.clk(gclk));
	jdff dff_A_92H3T4840_1(.dout(w_dff_A_Q7ura78J7_1),.din(w_dff_A_92H3T4840_1),.clk(gclk));
	jdff dff_A_uDYQkja50_1(.dout(w_dff_A_92H3T4840_1),.din(w_dff_A_uDYQkja50_1),.clk(gclk));
	jdff dff_A_umE1GkFi4_1(.dout(w_dff_A_uDYQkja50_1),.din(w_dff_A_umE1GkFi4_1),.clk(gclk));
	jdff dff_A_BFcuhVbu6_1(.dout(w_dff_A_umE1GkFi4_1),.din(w_dff_A_BFcuhVbu6_1),.clk(gclk));
	jdff dff_A_k97hcDSh2_1(.dout(w_G343_0[1]),.din(w_dff_A_k97hcDSh2_1),.clk(gclk));
	jdff dff_A_aunUDTkh1_1(.dout(w_dff_A_k97hcDSh2_1),.din(w_dff_A_aunUDTkh1_1),.clk(gclk));
	jdff dff_A_Su7s7ao33_1(.dout(w_dff_A_aunUDTkh1_1),.din(w_dff_A_Su7s7ao33_1),.clk(gclk));
	jdff dff_A_OLc4brm52_1(.dout(w_n374_0[1]),.din(w_dff_A_OLc4brm52_1),.clk(gclk));
	jdff dff_B_nuHoV5pA2_0(.din(n365),.dout(w_dff_B_nuHoV5pA2_0),.clk(gclk));
	jdff dff_B_Dh2jux470_1(.din(n348),.dout(w_dff_B_Dh2jux470_1),.clk(gclk));
	jdff dff_B_0LuljrnG7_1(.din(n343),.dout(w_dff_B_0LuljrnG7_1),.clk(gclk));
	jdff dff_A_c2WzAXFN8_0(.dout(w_n339_0[0]),.din(w_dff_A_c2WzAXFN8_0),.clk(gclk));
	jdff dff_A_S9HSg5NO7_0(.dout(w_dff_A_c2WzAXFN8_0),.din(w_dff_A_S9HSg5NO7_0),.clk(gclk));
	jdff dff_A_7Og8lSIe5_0(.dout(w_G294_3[0]),.din(w_dff_A_7Og8lSIe5_0),.clk(gclk));
	jdff dff_A_Bn0WMGDC3_0(.dout(w_dff_A_7Og8lSIe5_0),.din(w_dff_A_Bn0WMGDC3_0),.clk(gclk));
	jdff dff_A_mMUfU7md6_0(.dout(w_dff_A_Bn0WMGDC3_0),.din(w_dff_A_mMUfU7md6_0),.clk(gclk));
	jdff dff_A_GsTMAoUY0_0(.dout(w_dff_A_mMUfU7md6_0),.din(w_dff_A_GsTMAoUY0_0),.clk(gclk));
	jdff dff_A_pnpF4iId6_0(.dout(w_G294_0[0]),.din(w_dff_A_pnpF4iId6_0),.clk(gclk));
	jdff dff_A_fjjXIW3l0_0(.dout(w_dff_A_pnpF4iId6_0),.din(w_dff_A_fjjXIW3l0_0),.clk(gclk));
	jdff dff_A_IwzbsjN37_0(.dout(w_dff_A_fjjXIW3l0_0),.din(w_dff_A_IwzbsjN37_0),.clk(gclk));
	jdff dff_A_J5Js87zm5_1(.dout(w_G294_0[1]),.din(w_dff_A_J5Js87zm5_1),.clk(gclk));
	jdff dff_A_5N0sKK5d5_1(.dout(w_dff_A_J5Js87zm5_1),.din(w_dff_A_5N0sKK5d5_1),.clk(gclk));
	jdff dff_A_KiT15BBB8_1(.dout(w_dff_A_5N0sKK5d5_1),.din(w_dff_A_KiT15BBB8_1),.clk(gclk));
	jdff dff_A_pH3RywLK4_0(.dout(w_n196_1[0]),.din(w_dff_A_pH3RywLK4_0),.clk(gclk));
	jdff dff_A_mgJE9RLR9_1(.dout(w_n196_1[1]),.din(w_dff_A_mgJE9RLR9_1),.clk(gclk));
	jdff dff_B_xrpfOxV02_0(.din(n335),.dout(w_dff_B_xrpfOxV02_0),.clk(gclk));
	jdff dff_A_i2aqhp5d0_0(.dout(w_n334_0[0]),.din(w_dff_A_i2aqhp5d0_0),.clk(gclk));
	jdff dff_A_luOPKde94_0(.dout(w_dff_A_i2aqhp5d0_0),.din(w_dff_A_luOPKde94_0),.clk(gclk));
	jdff dff_B_UDmTyMk91_0(.din(n333),.dout(w_dff_B_UDmTyMk91_0),.clk(gclk));
	jdff dff_A_p2P0Q2Iy0_0(.dout(w_G107_3[0]),.din(w_dff_A_p2P0Q2Iy0_0),.clk(gclk));
	jdff dff_A_HoFi2L3R1_1(.dout(w_G107_3[1]),.din(w_dff_A_HoFi2L3R1_1),.clk(gclk));
	jdff dff_B_MNYOayjY1_0(.din(n331),.dout(w_dff_B_MNYOayjY1_0),.clk(gclk));
	jdff dff_B_WMEaKdvL2_1(.din(n316),.dout(w_dff_B_WMEaKdvL2_1),.clk(gclk));
	jdff dff_A_PYEzkkyH2_1(.dout(w_G190_3[1]),.din(w_dff_A_PYEzkkyH2_1),.clk(gclk));
	jdff dff_A_yvxDBaBU2_1(.dout(w_dff_A_PYEzkkyH2_1),.din(w_dff_A_yvxDBaBU2_1),.clk(gclk));
	jdff dff_A_SZozDlnA3_1(.dout(w_dff_A_yvxDBaBU2_1),.din(w_dff_A_SZozDlnA3_1),.clk(gclk));
	jdff dff_A_5HCXgE3r5_1(.dout(w_dff_A_SZozDlnA3_1),.din(w_dff_A_5HCXgE3r5_1),.clk(gclk));
	jdff dff_A_FDG7s6lR2_1(.dout(w_dff_A_5HCXgE3r5_1),.din(w_dff_A_FDG7s6lR2_1),.clk(gclk));
	jdff dff_A_C3p8AZF36_1(.dout(w_dff_A_FDG7s6lR2_1),.din(w_dff_A_C3p8AZF36_1),.clk(gclk));
	jdff dff_A_XHC4JfNo2_1(.dout(w_dff_A_C3p8AZF36_1),.din(w_dff_A_XHC4JfNo2_1),.clk(gclk));
	jdff dff_A_Jks76VVu9_2(.dout(w_G190_3[2]),.din(w_dff_A_Jks76VVu9_2),.clk(gclk));
	jdff dff_A_JpmrROEI9_2(.dout(w_dff_A_Jks76VVu9_2),.din(w_dff_A_JpmrROEI9_2),.clk(gclk));
	jdff dff_A_htK27Vyk1_2(.dout(w_dff_A_JpmrROEI9_2),.din(w_dff_A_htK27Vyk1_2),.clk(gclk));
	jdff dff_A_MFiCQyL13_2(.dout(w_dff_A_htK27Vyk1_2),.din(w_dff_A_MFiCQyL13_2),.clk(gclk));
	jdff dff_A_mdaEY9wk8_2(.dout(w_dff_A_MFiCQyL13_2),.din(w_dff_A_mdaEY9wk8_2),.clk(gclk));
	jdff dff_A_FpXd7hDV2_2(.dout(w_dff_A_mdaEY9wk8_2),.din(w_dff_A_FpXd7hDV2_2),.clk(gclk));
	jdff dff_A_59Z4Cv8n6_2(.dout(w_dff_A_FpXd7hDV2_2),.din(w_dff_A_59Z4Cv8n6_2),.clk(gclk));
	jdff dff_B_igReF1fn0_0(.din(n317),.dout(w_dff_B_igReF1fn0_0),.clk(gclk));
	jdff dff_B_IpaO9w8W7_1(.din(n289),.dout(w_dff_B_IpaO9w8W7_1),.clk(gclk));
	jdff dff_A_kyk90hop2_1(.dout(w_n312_0[1]),.din(w_dff_A_kyk90hop2_1),.clk(gclk));
	jdff dff_B_xzNoOxiA6_1(.din(n309),.dout(w_dff_B_xzNoOxiA6_1),.clk(gclk));
	jdff dff_A_v5uxyzdr9_0(.dout(w_n106_0[0]),.din(w_dff_A_v5uxyzdr9_0),.clk(gclk));
	jdff dff_A_HZLZcV8W5_0(.dout(w_dff_A_v5uxyzdr9_0),.din(w_dff_A_HZLZcV8W5_0),.clk(gclk));
	jdff dff_A_kgIT8jEI1_0(.dout(w_dff_A_HZLZcV8W5_0),.din(w_dff_A_kgIT8jEI1_0),.clk(gclk));
	jdff dff_A_YG7pT8e90_1(.dout(w_n88_0[1]),.din(w_dff_A_YG7pT8e90_1),.clk(gclk));
	jdff dff_A_9jxpiqiL7_1(.dout(w_dff_A_YG7pT8e90_1),.din(w_dff_A_9jxpiqiL7_1),.clk(gclk));
	jdff dff_A_Q14htJgy1_1(.dout(w_dff_A_9jxpiqiL7_1),.din(w_dff_A_Q14htJgy1_1),.clk(gclk));
	jdff dff_A_UANVtvih1_2(.dout(w_n88_0[2]),.din(w_dff_A_UANVtvih1_2),.clk(gclk));
	jdff dff_A_oSJIeN5g9_1(.dout(w_n166_1[1]),.din(w_dff_A_oSJIeN5g9_1),.clk(gclk));
	jdff dff_A_0HjbQwMa6_2(.dout(w_n166_1[2]),.din(w_dff_A_0HjbQwMa6_2),.clk(gclk));
	jdff dff_A_O5qOvHQS3_1(.dout(w_n303_0[1]),.din(w_dff_A_O5qOvHQS3_1),.clk(gclk));
	jdff dff_A_8bu2HjsL3_1(.dout(w_n300_0[1]),.din(w_dff_A_8bu2HjsL3_1),.clk(gclk));
	jdff dff_A_stTYGT9I3_0(.dout(w_n298_0[0]),.din(w_dff_A_stTYGT9I3_0),.clk(gclk));
	jdff dff_A_gFIWSjUS3_0(.dout(w_dff_A_stTYGT9I3_0),.din(w_dff_A_gFIWSjUS3_0),.clk(gclk));
	jdff dff_A_mo8oFZxj4_1(.dout(w_n185_2[1]),.din(w_dff_A_mo8oFZxj4_1),.clk(gclk));
	jdff dff_A_jBWtepp39_1(.dout(w_dff_A_mo8oFZxj4_1),.din(w_dff_A_jBWtepp39_1),.clk(gclk));
	jdff dff_A_0cZKzsvq7_0(.dout(w_n105_1[0]),.din(w_dff_A_0cZKzsvq7_0),.clk(gclk));
	jdff dff_A_1Sn75JW53_2(.dout(w_n105_1[2]),.din(w_dff_A_1Sn75JW53_2),.clk(gclk));
	jdff dff_A_GzRYhqYM5_0(.dout(w_n296_0[0]),.din(w_dff_A_GzRYhqYM5_0),.clk(gclk));
	jdff dff_A_3zW65Z0I5_0(.dout(w_dff_A_GzRYhqYM5_0),.din(w_dff_A_3zW65Z0I5_0),.clk(gclk));
	jdff dff_A_uDH37AKn4_0(.dout(w_n105_0[0]),.din(w_dff_A_uDH37AKn4_0),.clk(gclk));
	jdff dff_A_ubeslu0t4_2(.dout(w_n105_0[2]),.din(w_dff_A_ubeslu0t4_2),.clk(gclk));
	jdff dff_A_iFfqgdzM0_2(.dout(w_dff_A_ubeslu0t4_2),.din(w_dff_A_iFfqgdzM0_2),.clk(gclk));
	jdff dff_A_BWR7BzNB9_2(.dout(w_dff_A_iFfqgdzM0_2),.din(w_dff_A_BWR7BzNB9_2),.clk(gclk));
	jdff dff_A_KXGCIGqG1_0(.dout(w_G20_4[0]),.din(w_dff_A_KXGCIGqG1_0),.clk(gclk));
	jdff dff_A_zOSz57x41_1(.dout(w_G20_4[1]),.din(w_dff_A_zOSz57x41_1),.clk(gclk));
	jdff dff_A_JBeus7uJ0_1(.dout(w_dff_A_zOSz57x41_1),.din(w_dff_A_JBeus7uJ0_1),.clk(gclk));
	jdff dff_A_7SAmofy49_1(.dout(w_dff_A_JBeus7uJ0_1),.din(w_dff_A_7SAmofy49_1),.clk(gclk));
	jdff dff_A_13G9R5bH5_1(.dout(w_dff_A_7SAmofy49_1),.din(w_dff_A_13G9R5bH5_1),.clk(gclk));
	jdff dff_A_BAlsuDBm7_1(.dout(w_n189_1[1]),.din(w_dff_A_BAlsuDBm7_1),.clk(gclk));
	jdff dff_A_jfWcgGkF8_0(.dout(w_G97_3[0]),.din(w_dff_A_jfWcgGkF8_0),.clk(gclk));
	jdff dff_A_hTVxTAEg9_0(.dout(w_dff_A_jfWcgGkF8_0),.din(w_dff_A_hTVxTAEg9_0),.clk(gclk));
	jdff dff_A_zgFStbQ32_0(.dout(w_dff_A_hTVxTAEg9_0),.din(w_dff_A_zgFStbQ32_0),.clk(gclk));
	jdff dff_A_DyEtyjAH1_1(.dout(w_G97_3[1]),.din(w_dff_A_DyEtyjAH1_1),.clk(gclk));
	jdff dff_A_Y612Y2Iu4_1(.dout(w_dff_A_DyEtyjAH1_1),.din(w_dff_A_Y612Y2Iu4_1),.clk(gclk));
	jdff dff_A_ccuwuU1G7_1(.dout(w_dff_A_Y612Y2Iu4_1),.din(w_dff_A_ccuwuU1G7_1),.clk(gclk));
	jdff dff_A_fhN7CvxK0_0(.dout(w_G270_0[0]),.din(w_dff_A_fhN7CvxK0_0),.clk(gclk));
	jdff dff_A_5tAOFhHm9_0(.dout(w_dff_A_fhN7CvxK0_0),.din(w_dff_A_5tAOFhHm9_0),.clk(gclk));
	jdff dff_A_wltsfTSv8_0(.dout(w_dff_A_5tAOFhHm9_0),.din(w_dff_A_wltsfTSv8_0),.clk(gclk));
	jdff dff_A_vbCK6CD48_0(.dout(w_dff_A_wltsfTSv8_0),.din(w_dff_A_vbCK6CD48_0),.clk(gclk));
	jdff dff_B_TqeE9gwh0_1(.din(n280),.dout(w_dff_B_TqeE9gwh0_1),.clk(gclk));
	jdff dff_A_mVRfsAVZ1_1(.dout(w_n281_0[1]),.din(w_dff_A_mVRfsAVZ1_1),.clk(gclk));
	jdff dff_A_1Aer3cB25_1(.dout(w_dff_A_mVRfsAVZ1_1),.din(w_dff_A_1Aer3cB25_1),.clk(gclk));
	jdff dff_A_fsN6Eq2c3_0(.dout(w_G303_2[0]),.din(w_dff_A_fsN6Eq2c3_0),.clk(gclk));
	jdff dff_A_HmsmWUc61_0(.dout(w_dff_A_fsN6Eq2c3_0),.din(w_dff_A_HmsmWUc61_0),.clk(gclk));
	jdff dff_A_aqNT9f7j3_0(.dout(w_dff_A_HmsmWUc61_0),.din(w_dff_A_aqNT9f7j3_0),.clk(gclk));
	jdff dff_A_xeeYnU4x7_1(.dout(w_G303_2[1]),.din(w_dff_A_xeeYnU4x7_1),.clk(gclk));
	jdff dff_A_xhzSbQc21_1(.dout(w_dff_A_xeeYnU4x7_1),.din(w_dff_A_xhzSbQc21_1),.clk(gclk));
	jdff dff_A_x85Fx5Bk9_1(.dout(w_dff_A_xhzSbQc21_1),.din(w_dff_A_x85Fx5Bk9_1),.clk(gclk));
	jdff dff_A_pNIHpZ1O9_1(.dout(w_dff_A_x85Fx5Bk9_1),.din(w_dff_A_pNIHpZ1O9_1),.clk(gclk));
	jdff dff_A_anOMJ07M0_0(.dout(w_G303_0[0]),.din(w_dff_A_anOMJ07M0_0),.clk(gclk));
	jdff dff_A_6Rvvtwnz2_0(.dout(w_dff_A_anOMJ07M0_0),.din(w_dff_A_6Rvvtwnz2_0),.clk(gclk));
	jdff dff_A_JSgvNSVS9_0(.dout(w_dff_A_6Rvvtwnz2_0),.din(w_dff_A_JSgvNSVS9_0),.clk(gclk));
	jdff dff_A_9pmlRJzT8_2(.dout(w_G303_0[2]),.din(w_dff_A_9pmlRJzT8_2),.clk(gclk));
	jdff dff_A_I7DHatgn6_2(.dout(w_dff_A_9pmlRJzT8_2),.din(w_dff_A_I7DHatgn6_2),.clk(gclk));
	jdff dff_A_AWdAOljJ4_2(.dout(w_dff_A_I7DHatgn6_2),.din(w_dff_A_AWdAOljJ4_2),.clk(gclk));
	jdff dff_A_bKPcwFxw3_2(.dout(w_dff_A_AWdAOljJ4_2),.din(w_dff_A_bKPcwFxw3_2),.clk(gclk));
	jdff dff_A_x2ult2f57_1(.dout(w_G264_0[1]),.din(w_dff_A_x2ult2f57_1),.clk(gclk));
	jdff dff_A_BcTVejTc8_1(.dout(w_dff_A_x2ult2f57_1),.din(w_dff_A_BcTVejTc8_1),.clk(gclk));
	jdff dff_A_h14eZX9o8_1(.dout(w_dff_A_BcTVejTc8_1),.din(w_dff_A_h14eZX9o8_1),.clk(gclk));
	jdff dff_A_MmzHCcUA0_1(.dout(w_dff_A_h14eZX9o8_1),.din(w_dff_A_MmzHCcUA0_1),.clk(gclk));
	jdff dff_A_nuy12LkE4_2(.dout(w_G264_0[2]),.din(w_dff_A_nuy12LkE4_2),.clk(gclk));
	jdff dff_A_iinwmgc79_2(.dout(w_dff_A_nuy12LkE4_2),.din(w_dff_A_iinwmgc79_2),.clk(gclk));
	jdff dff_B_E1mUxj7c0_1(.din(n268),.dout(w_dff_B_E1mUxj7c0_1),.clk(gclk));
	jdff dff_A_Wl9EksWk0_1(.dout(w_n274_0[1]),.din(w_dff_A_Wl9EksWk0_1),.clk(gclk));
	jdff dff_A_g5LRjXiN1_0(.dout(w_n270_0[0]),.din(w_dff_A_g5LRjXiN1_0),.clk(gclk));
	jdff dff_B_SP53AS286_2(.din(n270),.dout(w_dff_B_SP53AS286_2),.clk(gclk));
	jdff dff_A_KlMvPo997_0(.dout(w_n112_4[0]),.din(w_dff_A_KlMvPo997_0),.clk(gclk));
	jdff dff_A_qbX6Uqo06_0(.dout(w_dff_A_KlMvPo997_0),.din(w_dff_A_qbX6Uqo06_0),.clk(gclk));
	jdff dff_A_lAM3NFgD3_0(.dout(w_dff_A_qbX6Uqo06_0),.din(w_dff_A_lAM3NFgD3_0),.clk(gclk));
	jdff dff_A_TxZONEDW8_0(.dout(w_dff_A_lAM3NFgD3_0),.din(w_dff_A_TxZONEDW8_0),.clk(gclk));
	jdff dff_A_5pCyFonK3_1(.dout(w_n112_4[1]),.din(w_dff_A_5pCyFonK3_1),.clk(gclk));
	jdff dff_A_VJNwAm6t4_0(.dout(w_G1_1[0]),.din(w_dff_A_VJNwAm6t4_0),.clk(gclk));
	jdff dff_A_HhEUSmbu4_0(.dout(w_dff_A_VJNwAm6t4_0),.din(w_dff_A_HhEUSmbu4_0),.clk(gclk));
	jdff dff_A_ic6VYL2s1_0(.dout(w_dff_A_HhEUSmbu4_0),.din(w_dff_A_ic6VYL2s1_0),.clk(gclk));
	jdff dff_A_nxOb1jX52_1(.dout(w_G1_1[1]),.din(w_dff_A_nxOb1jX52_1),.clk(gclk));
	jdff dff_B_sT0q3vOJ5_0(.din(n266),.dout(w_dff_B_sT0q3vOJ5_0),.clk(gclk));
	jdff dff_B_wdu0KqcM0_1(.din(n260),.dout(w_dff_B_wdu0KqcM0_1),.clk(gclk));
	jdff dff_A_AribFjuc2_0(.dout(w_n262_0[0]),.din(w_dff_A_AribFjuc2_0),.clk(gclk));
	jdff dff_A_EJ8QD03f7_0(.dout(w_n259_0[0]),.din(w_dff_A_EJ8QD03f7_0),.clk(gclk));
	jdff dff_A_v7wVNXzV8_0(.dout(w_dff_A_EJ8QD03f7_0),.din(w_dff_A_v7wVNXzV8_0),.clk(gclk));
	jdff dff_A_Esk9FLPn0_0(.dout(w_n257_0[0]),.din(w_dff_A_Esk9FLPn0_0),.clk(gclk));
	jdff dff_A_DIxhcRxu7_1(.dout(w_n255_0[1]),.din(w_dff_A_DIxhcRxu7_1),.clk(gclk));
	jdff dff_A_dfSf8Hys6_0(.dout(w_G77_4[0]),.din(w_dff_A_dfSf8Hys6_0),.clk(gclk));
	jdff dff_A_ByuNwsEG1_0(.dout(w_G77_1[0]),.din(w_dff_A_ByuNwsEG1_0),.clk(gclk));
	jdff dff_A_pllA2Bln3_2(.dout(w_G77_1[2]),.din(w_dff_A_pllA2Bln3_2),.clk(gclk));
	jdff dff_A_7RCLjyTf9_2(.dout(w_dff_A_pllA2Bln3_2),.din(w_dff_A_7RCLjyTf9_2),.clk(gclk));
	jdff dff_A_oAMkPFud9_2(.dout(w_dff_A_7RCLjyTf9_2),.din(w_dff_A_oAMkPFud9_2),.clk(gclk));
	jdff dff_A_WUSlaZ817_2(.dout(w_dff_A_oAMkPFud9_2),.din(w_dff_A_WUSlaZ817_2),.clk(gclk));
	jdff dff_B_bwUjs0ls1_2(.din(n249),.dout(w_dff_B_bwUjs0ls1_2),.clk(gclk));
	jdff dff_B_ZgjgcbpT5_2(.din(w_dff_B_bwUjs0ls1_2),.dout(w_dff_B_ZgjgcbpT5_2),.clk(gclk));
	jdff dff_A_xsnjI4353_0(.dout(w_G107_4[0]),.din(w_dff_A_xsnjI4353_0),.clk(gclk));
	jdff dff_A_FREIkpu59_0(.dout(w_dff_A_xsnjI4353_0),.din(w_dff_A_FREIkpu59_0),.clk(gclk));
	jdff dff_A_iaCFZwZi5_0(.dout(w_dff_A_FREIkpu59_0),.din(w_dff_A_iaCFZwZi5_0),.clk(gclk));
	jdff dff_A_uORXY95T9_0(.dout(w_dff_A_iaCFZwZi5_0),.din(w_dff_A_uORXY95T9_0),.clk(gclk));
	jdff dff_A_wQjxCHQ43_0(.dout(w_dff_A_uORXY95T9_0),.din(w_dff_A_wQjxCHQ43_0),.clk(gclk));
	jdff dff_A_oJvYPEnJ3_0(.dout(w_dff_A_wQjxCHQ43_0),.din(w_dff_A_oJvYPEnJ3_0),.clk(gclk));
	jdff dff_A_PfzZNePP1_0(.dout(w_G33_8[0]),.din(w_dff_A_PfzZNePP1_0),.clk(gclk));
	jdff dff_B_HzC0cx2C7_1(.din(n236),.dout(w_dff_B_HzC0cx2C7_1),.clk(gclk));
	jdff dff_B_pauv6il10_1(.din(n226),.dout(w_dff_B_pauv6il10_1),.clk(gclk));
	jdff dff_A_MjqUp2IV7_0(.dout(w_n230_0[0]),.din(w_dff_A_MjqUp2IV7_0),.clk(gclk));
	jdff dff_A_eLh1wXtP2_0(.dout(w_n151_3[0]),.din(w_dff_A_eLh1wXtP2_0),.clk(gclk));
	jdff dff_A_HOvEmfsF0_0(.dout(w_dff_A_eLh1wXtP2_0),.din(w_dff_A_HOvEmfsF0_0),.clk(gclk));
	jdff dff_A_rT4nJnsx9_1(.dout(w_n151_3[1]),.din(w_dff_A_rT4nJnsx9_1),.clk(gclk));
	jdff dff_A_H6Myhpd09_1(.dout(w_dff_A_rT4nJnsx9_1),.din(w_dff_A_H6Myhpd09_1),.clk(gclk));
	jdff dff_A_Mc4qclDQ7_0(.dout(w_n91_1[0]),.din(w_dff_A_Mc4qclDQ7_0),.clk(gclk));
	jdff dff_A_VcdHeGSe5_0(.dout(w_dff_A_Mc4qclDQ7_0),.din(w_dff_A_VcdHeGSe5_0),.clk(gclk));
	jdff dff_A_QS6hAFmE7_0(.dout(w_dff_A_VcdHeGSe5_0),.din(w_dff_A_QS6hAFmE7_0),.clk(gclk));
	jdff dff_A_PsGS15dS5_1(.dout(w_n91_0[1]),.din(w_dff_A_PsGS15dS5_1),.clk(gclk));
	jdff dff_A_FROdvvJx1_0(.dout(w_G257_1[0]),.din(w_dff_A_FROdvvJx1_0),.clk(gclk));
	jdff dff_A_OEyQfNX14_0(.dout(w_dff_A_FROdvvJx1_0),.din(w_dff_A_OEyQfNX14_0),.clk(gclk));
	jdff dff_A_llzU1GyE4_0(.dout(w_dff_A_OEyQfNX14_0),.din(w_dff_A_llzU1GyE4_0),.clk(gclk));
	jdff dff_A_EcODS1TM6_0(.dout(w_dff_A_llzU1GyE4_0),.din(w_dff_A_EcODS1TM6_0),.clk(gclk));
	jdff dff_A_TfyK3HW66_1(.dout(w_G257_1[1]),.din(w_dff_A_TfyK3HW66_1),.clk(gclk));
	jdff dff_A_B60DKuWp4_1(.dout(w_G257_0[1]),.din(w_dff_A_B60DKuWp4_1),.clk(gclk));
	jdff dff_A_l4Toek0g7_1(.dout(w_dff_A_B60DKuWp4_1),.din(w_dff_A_l4Toek0g7_1),.clk(gclk));
	jdff dff_A_IbB9Taz62_2(.dout(w_G257_0[2]),.din(w_dff_A_IbB9Taz62_2),.clk(gclk));
	jdff dff_A_irs9bHBr5_2(.dout(w_dff_A_IbB9Taz62_2),.din(w_dff_A_irs9bHBr5_2),.clk(gclk));
	jdff dff_A_DtA0yE6o6_1(.dout(w_n228_0[1]),.din(w_dff_A_DtA0yE6o6_1),.clk(gclk));
	jdff dff_A_udrKFxna6_0(.dout(w_n221_0[0]),.din(w_dff_A_udrKFxna6_0),.clk(gclk));
	jdff dff_A_3xRNxzVm0_0(.dout(w_dff_A_udrKFxna6_0),.din(w_dff_A_3xRNxzVm0_0),.clk(gclk));
	jdff dff_A_wFYZV4pb7_1(.dout(w_n221_0[1]),.din(w_dff_A_wFYZV4pb7_1),.clk(gclk));
	jdff dff_A_zzM06KLE7_1(.dout(w_dff_A_wFYZV4pb7_1),.din(w_dff_A_zzM06KLE7_1),.clk(gclk));
	jdff dff_A_e6fQA4aB6_0(.dout(w_G283_3[0]),.din(w_dff_A_e6fQA4aB6_0),.clk(gclk));
	jdff dff_A_JnrTIHvl0_0(.dout(w_dff_A_e6fQA4aB6_0),.din(w_dff_A_JnrTIHvl0_0),.clk(gclk));
	jdff dff_A_8GO6iolU1_0(.dout(w_dff_A_JnrTIHvl0_0),.din(w_dff_A_8GO6iolU1_0),.clk(gclk));
	jdff dff_A_KPDjnYZZ5_1(.dout(w_G283_3[1]),.din(w_dff_A_KPDjnYZZ5_1),.clk(gclk));
	jdff dff_A_G3VZeg0G8_1(.dout(w_dff_A_KPDjnYZZ5_1),.din(w_dff_A_G3VZeg0G8_1),.clk(gclk));
	jdff dff_A_RndfyFv52_1(.dout(w_dff_A_G3VZeg0G8_1),.din(w_dff_A_RndfyFv52_1),.clk(gclk));
	jdff dff_A_U3y76x5D0_1(.dout(w_dff_A_RndfyFv52_1),.din(w_dff_A_U3y76x5D0_1),.clk(gclk));
	jdff dff_A_vc88hoFt9_0(.dout(w_G283_0[0]),.din(w_dff_A_vc88hoFt9_0),.clk(gclk));
	jdff dff_A_m64AZkit3_0(.dout(w_dff_A_vc88hoFt9_0),.din(w_dff_A_m64AZkit3_0),.clk(gclk));
	jdff dff_A_REC5uBRg6_0(.dout(w_dff_A_m64AZkit3_0),.din(w_dff_A_REC5uBRg6_0),.clk(gclk));
	jdff dff_A_32enTWEY8_1(.dout(w_G283_0[1]),.din(w_dff_A_32enTWEY8_1),.clk(gclk));
	jdff dff_A_M3EiS25C9_1(.dout(w_dff_A_32enTWEY8_1),.din(w_dff_A_M3EiS25C9_1),.clk(gclk));
	jdff dff_A_zlfUFNxN7_1(.dout(w_dff_A_M3EiS25C9_1),.din(w_dff_A_zlfUFNxN7_1),.clk(gclk));
	jdff dff_A_EhSyXoq93_2(.dout(w_n166_2[2]),.din(w_dff_A_EhSyXoq93_2),.clk(gclk));
	jdff dff_B_suPl964r6_1(.din(n215),.dout(w_dff_B_suPl964r6_1),.clk(gclk));
	jdff dff_A_8yi5hHaE5_0(.dout(w_G200_1[0]),.din(w_dff_A_8yi5hHaE5_0),.clk(gclk));
	jdff dff_A_26xsE9xa2_0(.dout(w_dff_A_8yi5hHaE5_0),.din(w_dff_A_26xsE9xa2_0),.clk(gclk));
	jdff dff_A_lt9IHk169_0(.dout(w_dff_A_26xsE9xa2_0),.din(w_dff_A_lt9IHk169_0),.clk(gclk));
	jdff dff_A_4CpzGqHi7_0(.dout(w_dff_A_lt9IHk169_0),.din(w_dff_A_4CpzGqHi7_0),.clk(gclk));
	jdff dff_A_mWcYaPyM8_0(.dout(w_dff_A_4CpzGqHi7_0),.din(w_dff_A_mWcYaPyM8_0),.clk(gclk));
	jdff dff_A_3FKnpT776_0(.dout(w_dff_A_mWcYaPyM8_0),.din(w_dff_A_3FKnpT776_0),.clk(gclk));
	jdff dff_A_bGE5KNDJ7_0(.dout(w_dff_A_3FKnpT776_0),.din(w_dff_A_bGE5KNDJ7_0),.clk(gclk));
	jdff dff_A_2pTMC7fh9_1(.dout(w_G200_1[1]),.din(w_dff_A_2pTMC7fh9_1),.clk(gclk));
	jdff dff_A_2nITGxT72_2(.dout(w_G200_0[2]),.din(w_dff_A_2nITGxT72_2),.clk(gclk));
	jdff dff_A_I4W3GC0P2_2(.dout(w_dff_A_2nITGxT72_2),.din(w_dff_A_I4W3GC0P2_2),.clk(gclk));
	jdff dff_A_bN7ldxU20_2(.dout(w_dff_A_I4W3GC0P2_2),.din(w_dff_A_bN7ldxU20_2),.clk(gclk));
	jdff dff_A_LPUcDJBS2_2(.dout(w_dff_A_bN7ldxU20_2),.din(w_dff_A_LPUcDJBS2_2),.clk(gclk));
	jdff dff_A_sMpOPvSM9_2(.dout(w_dff_A_LPUcDJBS2_2),.din(w_dff_A_sMpOPvSM9_2),.clk(gclk));
	jdff dff_A_4Il5uod24_2(.dout(w_dff_A_sMpOPvSM9_2),.din(w_dff_A_4Il5uod24_2),.clk(gclk));
	jdff dff_A_mJWlEdhi3_2(.dout(w_dff_A_4Il5uod24_2),.din(w_dff_A_mJWlEdhi3_2),.clk(gclk));
	jdff dff_A_qayL26XG4_0(.dout(w_G190_4[0]),.din(w_dff_A_qayL26XG4_0),.clk(gclk));
	jdff dff_A_wAzwG5NF6_0(.dout(w_G190_1[0]),.din(w_dff_A_wAzwG5NF6_0),.clk(gclk));
	jdff dff_A_eeXcb0LK1_0(.dout(w_dff_A_wAzwG5NF6_0),.din(w_dff_A_eeXcb0LK1_0),.clk(gclk));
	jdff dff_A_7rw9GJCL1_0(.dout(w_dff_A_eeXcb0LK1_0),.din(w_dff_A_7rw9GJCL1_0),.clk(gclk));
	jdff dff_A_tkwBkKGg1_0(.dout(w_dff_A_7rw9GJCL1_0),.din(w_dff_A_tkwBkKGg1_0),.clk(gclk));
	jdff dff_A_MToV3uQi0_0(.dout(w_G190_0[0]),.din(w_dff_A_MToV3uQi0_0),.clk(gclk));
	jdff dff_A_dVvesc1C1_0(.dout(w_dff_A_MToV3uQi0_0),.din(w_dff_A_dVvesc1C1_0),.clk(gclk));
	jdff dff_A_Ac1t2Z0B9_1(.dout(w_G190_0[1]),.din(w_dff_A_Ac1t2Z0B9_1),.clk(gclk));
	jdff dff_A_F0YiJfRp5_1(.dout(w_dff_A_Ac1t2Z0B9_1),.din(w_dff_A_F0YiJfRp5_1),.clk(gclk));
	jdff dff_A_wCBPIBH18_1(.dout(w_dff_A_F0YiJfRp5_1),.din(w_dff_A_wCBPIBH18_1),.clk(gclk));
	jdff dff_A_4kFVSjYh8_1(.dout(w_n214_0[1]),.din(w_dff_A_4kFVSjYh8_1),.clk(gclk));
	jdff dff_A_0M59mrjU1_1(.dout(w_n213_0[1]),.din(w_dff_A_0M59mrjU1_1),.clk(gclk));
	jdff dff_A_hz48tvZj2_0(.dout(w_n210_0[0]),.din(w_dff_A_hz48tvZj2_0),.clk(gclk));
	jdff dff_A_PbvQEbvw8_0(.dout(w_n205_0[0]),.din(w_dff_A_PbvQEbvw8_0),.clk(gclk));
	jdff dff_B_6KcOzGgC9_2(.din(n205),.dout(w_dff_B_6KcOzGgC9_2),.clk(gclk));
	jdff dff_A_mVCFVMyS7_0(.dout(w_n201_0[0]),.din(w_dff_A_mVCFVMyS7_0),.clk(gclk));
	jdff dff_A_uzO5xhyl4_2(.dout(w_G33_9[2]),.din(w_dff_A_uzO5xhyl4_2),.clk(gclk));
	jdff dff_A_6k8eSR7l3_1(.dout(w_n103_0[1]),.din(w_dff_A_6k8eSR7l3_1),.clk(gclk));
	jdff dff_A_PWuV5Axc5_0(.dout(w_n196_2[0]),.din(w_dff_A_PWuV5Axc5_0),.clk(gclk));
	jdff dff_A_VCFA39Bw3_1(.dout(w_n196_2[1]),.din(w_dff_A_VCFA39Bw3_1),.clk(gclk));
	jdff dff_A_ZTcFboHJ9_0(.dout(w_n196_0[0]),.din(w_dff_A_ZTcFboHJ9_0),.clk(gclk));
	jdff dff_A_JFjoZqRm7_2(.dout(w_n196_0[2]),.din(w_dff_A_JFjoZqRm7_2),.clk(gclk));
	jdff dff_B_T99fJxNq5_3(.din(n196),.dout(w_dff_B_T99fJxNq5_3),.clk(gclk));
	jdff dff_B_HskBRdxc1_3(.din(w_dff_B_T99fJxNq5_3),.dout(w_dff_B_HskBRdxc1_3),.clk(gclk));
	jdff dff_B_uYtT4eQu5_3(.din(w_dff_B_HskBRdxc1_3),.dout(w_dff_B_uYtT4eQu5_3),.clk(gclk));
	jdff dff_B_vNKcW1C49_3(.din(w_dff_B_uYtT4eQu5_3),.dout(w_dff_B_vNKcW1C49_3),.clk(gclk));
	jdff dff_B_kIJv506o1_3(.din(w_dff_B_vNKcW1C49_3),.dout(w_dff_B_kIJv506o1_3),.clk(gclk));
	jdff dff_A_xCs0uLOj3_0(.dout(w_G179_2[0]),.din(w_dff_A_xCs0uLOj3_0),.clk(gclk));
	jdff dff_A_XKSjJ5hH1_0(.dout(w_dff_A_xCs0uLOj3_0),.din(w_dff_A_XKSjJ5hH1_0),.clk(gclk));
	jdff dff_A_e7tTGEca3_0(.dout(w_dff_A_XKSjJ5hH1_0),.din(w_dff_A_e7tTGEca3_0),.clk(gclk));
	jdff dff_A_DE7AwlLp0_0(.dout(w_dff_A_e7tTGEca3_0),.din(w_dff_A_DE7AwlLp0_0),.clk(gclk));
	jdff dff_A_Ks2d8K442_0(.dout(w_dff_A_DE7AwlLp0_0),.din(w_dff_A_Ks2d8K442_0),.clk(gclk));
	jdff dff_A_Fqlu81ZI1_0(.dout(w_dff_A_Ks2d8K442_0),.din(w_dff_A_Fqlu81ZI1_0),.clk(gclk));
	jdff dff_A_suGe9WPO6_0(.dout(w_dff_A_Fqlu81ZI1_0),.din(w_dff_A_suGe9WPO6_0),.clk(gclk));
	jdff dff_A_DLUYiEM47_1(.dout(w_G179_2[1]),.din(w_dff_A_DLUYiEM47_1),.clk(gclk));
	jdff dff_A_hJM2TBQB1_1(.dout(w_dff_A_DLUYiEM47_1),.din(w_dff_A_hJM2TBQB1_1),.clk(gclk));
	jdff dff_A_q7JbCo8W6_1(.dout(w_dff_A_hJM2TBQB1_1),.din(w_dff_A_q7JbCo8W6_1),.clk(gclk));
	jdff dff_A_QzUOOnDj6_1(.dout(w_dff_A_q7JbCo8W6_1),.din(w_dff_A_QzUOOnDj6_1),.clk(gclk));
	jdff dff_A_q1vMp6Xt8_1(.dout(w_dff_A_QzUOOnDj6_1),.din(w_dff_A_q1vMp6Xt8_1),.clk(gclk));
	jdff dff_A_7k4l7qt24_1(.dout(w_dff_A_q1vMp6Xt8_1),.din(w_dff_A_7k4l7qt24_1),.clk(gclk));
	jdff dff_A_J1ih0qTn6_1(.dout(w_dff_A_7k4l7qt24_1),.din(w_dff_A_J1ih0qTn6_1),.clk(gclk));
	jdff dff_A_lF4JxzxQ2_0(.dout(w_G179_0[0]),.din(w_dff_A_lF4JxzxQ2_0),.clk(gclk));
	jdff dff_A_4SFMbZqQ6_0(.dout(w_dff_A_lF4JxzxQ2_0),.din(w_dff_A_4SFMbZqQ6_0),.clk(gclk));
	jdff dff_A_ZUQtZJlv5_0(.dout(w_dff_A_4SFMbZqQ6_0),.din(w_dff_A_ZUQtZJlv5_0),.clk(gclk));
	jdff dff_A_WJoMVyUr7_0(.dout(w_dff_A_ZUQtZJlv5_0),.din(w_dff_A_WJoMVyUr7_0),.clk(gclk));
	jdff dff_A_NS9sNu3e4_0(.dout(w_dff_A_WJoMVyUr7_0),.din(w_dff_A_NS9sNu3e4_0),.clk(gclk));
	jdff dff_A_f208jTEV9_0(.dout(w_dff_A_NS9sNu3e4_0),.din(w_dff_A_f208jTEV9_0),.clk(gclk));
	jdff dff_A_Dr0dLoVk1_0(.dout(w_dff_A_f208jTEV9_0),.din(w_dff_A_Dr0dLoVk1_0),.clk(gclk));
	jdff dff_B_CTKC3q9z3_0(.din(n192),.dout(w_dff_B_CTKC3q9z3_0),.clk(gclk));
	jdff dff_A_BhaIHiIi3_1(.dout(w_n190_1[1]),.din(w_dff_A_BhaIHiIi3_1),.clk(gclk));
	jdff dff_A_NTvaMBSR8_0(.dout(w_n189_2[0]),.din(w_dff_A_NTvaMBSR8_0),.clk(gclk));
	jdff dff_A_bYTrrIyV4_0(.dout(w_dff_A_NTvaMBSR8_0),.din(w_dff_A_bYTrrIyV4_0),.clk(gclk));
	jdff dff_A_ObhdSrtI1_2(.dout(w_n189_0[2]),.din(w_dff_A_ObhdSrtI1_2),.clk(gclk));
	jdff dff_A_tijpbY7D0_0(.dout(w_n85_0[0]),.din(w_dff_A_tijpbY7D0_0),.clk(gclk));
	jdff dff_A_65zy7shZ0_0(.dout(w_dff_A_tijpbY7D0_0),.din(w_dff_A_65zy7shZ0_0),.clk(gclk));
	jdff dff_A_UAB7M2MC5_2(.dout(w_n85_0[2]),.din(w_dff_A_UAB7M2MC5_2),.clk(gclk));
	jdff dff_A_bDTE1pCU5_2(.dout(w_dff_A_UAB7M2MC5_2),.din(w_dff_A_bDTE1pCU5_2),.clk(gclk));
	jdff dff_A_VyS28cge1_2(.dout(w_dff_A_bDTE1pCU5_2),.din(w_dff_A_VyS28cge1_2),.clk(gclk));
	jdff dff_A_HZd2GatY8_2(.dout(w_dff_A_VyS28cge1_2),.din(w_dff_A_HZd2GatY8_2),.clk(gclk));
	jdff dff_A_tnr0FCP54_0(.dout(w_G20_5[0]),.din(w_dff_A_tnr0FCP54_0),.clk(gclk));
	jdff dff_A_J9rY81dQ7_1(.dout(w_G20_5[1]),.din(w_dff_A_J9rY81dQ7_1),.clk(gclk));
	jdff dff_A_gHYXEe3V2_1(.dout(w_n80_0[1]),.din(w_dff_A_gHYXEe3V2_1),.clk(gclk));
	jdff dff_A_sasnW2SN5_1(.dout(w_dff_A_gHYXEe3V2_1),.din(w_dff_A_sasnW2SN5_1),.clk(gclk));
	jdff dff_A_ffrbgNc21_1(.dout(w_dff_A_sasnW2SN5_1),.din(w_dff_A_ffrbgNc21_1),.clk(gclk));
	jdff dff_A_6luVzNKG7_2(.dout(w_n80_0[2]),.din(w_dff_A_6luVzNKG7_2),.clk(gclk));
	jdff dff_A_mnmkF3jC1_2(.dout(w_dff_A_6luVzNKG7_2),.din(w_dff_A_mnmkF3jC1_2),.clk(gclk));
	jdff dff_A_lqG2rG0X8_2(.dout(w_dff_A_mnmkF3jC1_2),.din(w_dff_A_lqG2rG0X8_2),.clk(gclk));
	jdff dff_A_Ilu1AmxG0_2(.dout(w_dff_A_lqG2rG0X8_2),.din(w_dff_A_Ilu1AmxG0_2),.clk(gclk));
	jdff dff_A_h6lmthOs1_2(.dout(w_dff_A_Ilu1AmxG0_2),.din(w_dff_A_h6lmthOs1_2),.clk(gclk));
	jdff dff_A_NY5FChnJ6_2(.dout(w_G107_1[2]),.din(w_dff_A_NY5FChnJ6_2),.clk(gclk));
	jdff dff_A_dmDIpHXg8_2(.dout(w_dff_A_NY5FChnJ6_2),.din(w_dff_A_dmDIpHXg8_2),.clk(gclk));
	jdff dff_A_O1jHvSWP8_2(.dout(w_dff_A_dmDIpHXg8_2),.din(w_dff_A_O1jHvSWP8_2),.clk(gclk));
	jdff dff_A_31bST4RG1_1(.dout(w_G107_0[1]),.din(w_dff_A_31bST4RG1_1),.clk(gclk));
	jdff dff_A_pd9Unxrj0_1(.dout(w_dff_A_31bST4RG1_1),.din(w_dff_A_pd9Unxrj0_1),.clk(gclk));
	jdff dff_A_FTkE7pQJ2_1(.dout(w_dff_A_pd9Unxrj0_1),.din(w_dff_A_FTkE7pQJ2_1),.clk(gclk));
	jdff dff_A_tsI1dVCL6_2(.dout(w_G107_0[2]),.din(w_dff_A_tsI1dVCL6_2),.clk(gclk));
	jdff dff_A_fWt6MUaE7_2(.dout(w_dff_A_tsI1dVCL6_2),.din(w_dff_A_fWt6MUaE7_2),.clk(gclk));
	jdff dff_A_pw1EcozM1_2(.dout(w_dff_A_fWt6MUaE7_2),.din(w_dff_A_pw1EcozM1_2),.clk(gclk));
	jdff dff_A_W52wfV0H7_0(.dout(w_n79_0[0]),.din(w_dff_A_W52wfV0H7_0),.clk(gclk));
	jdff dff_A_vIXjKMLs5_0(.dout(w_dff_A_W52wfV0H7_0),.din(w_dff_A_vIXjKMLs5_0),.clk(gclk));
	jdff dff_A_GViDkCJD7_0(.dout(w_G97_5[0]),.din(w_dff_A_GViDkCJD7_0),.clk(gclk));
	jdff dff_A_AZl59P653_1(.dout(w_n97_1[1]),.din(w_dff_A_AZl59P653_1),.clk(gclk));
	jdff dff_A_swqtA9sL9_0(.dout(w_n97_0[0]),.din(w_dff_A_swqtA9sL9_0),.clk(gclk));
	jdff dff_A_001aC8LN9_0(.dout(w_G87_3[0]),.din(w_dff_A_001aC8LN9_0),.clk(gclk));
	jdff dff_A_ZsQLVsqs3_2(.dout(w_G87_3[2]),.din(w_dff_A_ZsQLVsqs3_2),.clk(gclk));
	jdff dff_A_oGYHcEpi4_2(.dout(w_dff_A_ZsQLVsqs3_2),.din(w_dff_A_oGYHcEpi4_2),.clk(gclk));
	jdff dff_A_c7vPv7cN1_2(.dout(w_dff_A_oGYHcEpi4_2),.din(w_dff_A_c7vPv7cN1_2),.clk(gclk));
	jdff dff_A_3AMTUf409_0(.dout(w_G87_0[0]),.din(w_dff_A_3AMTUf409_0),.clk(gclk));
	jdff dff_A_vI1MDHPb8_0(.dout(w_dff_A_3AMTUf409_0),.din(w_dff_A_vI1MDHPb8_0),.clk(gclk));
	jdff dff_A_yTyBwOZq2_0(.dout(w_dff_A_vI1MDHPb8_0),.din(w_dff_A_yTyBwOZq2_0),.clk(gclk));
	jdff dff_A_w42ZATqo8_1(.dout(w_n179_0[1]),.din(w_dff_A_w42ZATqo8_1),.clk(gclk));
	jdff dff_A_jPwCkNEH8_1(.dout(w_dff_A_w42ZATqo8_1),.din(w_dff_A_jPwCkNEH8_1),.clk(gclk));
	jdff dff_A_Vmkku8fN4_2(.dout(w_n179_0[2]),.din(w_dff_A_Vmkku8fN4_2),.clk(gclk));
	jdff dff_A_F7j5jKl69_2(.dout(w_dff_A_Vmkku8fN4_2),.din(w_dff_A_F7j5jKl69_2),.clk(gclk));
	jdff dff_A_VSlHQ9P36_2(.dout(w_n112_5[2]),.din(w_dff_A_VSlHQ9P36_2),.clk(gclk));
	jdff dff_A_Madlfysn3_1(.dout(w_G20_2[1]),.din(w_dff_A_Madlfysn3_1),.clk(gclk));
	jdff dff_A_8wMjJHIG7_0(.dout(w_G68_4[0]),.din(w_dff_A_8wMjJHIG7_0),.clk(gclk));
	jdff dff_A_PJNWczpa1_1(.dout(w_G68_4[1]),.din(w_dff_A_PJNWczpa1_1),.clk(gclk));
	jdff dff_A_0corOKVj7_0(.dout(w_G68_1[0]),.din(w_dff_A_0corOKVj7_0),.clk(gclk));
	jdff dff_A_DxGsPXO13_2(.dout(w_G68_1[2]),.din(w_dff_A_DxGsPXO13_2),.clk(gclk));
	jdff dff_A_0ztcYfpW6_2(.dout(w_dff_A_DxGsPXO13_2),.din(w_dff_A_0ztcYfpW6_2),.clk(gclk));
	jdff dff_A_h2tkC4do5_2(.dout(w_dff_A_0ztcYfpW6_2),.din(w_dff_A_h2tkC4do5_2),.clk(gclk));
	jdff dff_A_aD3bYPsb3_2(.dout(w_dff_A_h2tkC4do5_2),.din(w_dff_A_aD3bYPsb3_2),.clk(gclk));
	jdff dff_A_si08ltWt9_2(.dout(w_G68_0[2]),.din(w_dff_A_si08ltWt9_2),.clk(gclk));
	jdff dff_A_1cQcbg208_1(.dout(w_n148_8[1]),.din(w_dff_A_1cQcbg208_1),.clk(gclk));
	jdff dff_A_1hQTGFhM4_0(.dout(w_G20_6[0]),.din(w_dff_A_1hQTGFhM4_0),.clk(gclk));
	jdff dff_A_Ekx2lsgO5_2(.dout(w_G20_1[2]),.din(w_dff_A_Ekx2lsgO5_2),.clk(gclk));
	jdff dff_A_nOj7S6af6_0(.dout(w_G20_0[0]),.din(w_dff_A_nOj7S6af6_0),.clk(gclk));
	jdff dff_B_dhtP6ddm7_2(.din(n172),.dout(w_dff_B_dhtP6ddm7_2),.clk(gclk));
	jdff dff_B_mCDef9Oe5_2(.din(w_dff_B_dhtP6ddm7_2),.dout(w_dff_B_mCDef9Oe5_2),.clk(gclk));
	jdff dff_A_iGp4QjM17_0(.dout(w_G97_4[0]),.din(w_dff_A_iGp4QjM17_0),.clk(gclk));
	jdff dff_A_VF4oUAvq4_0(.dout(w_dff_A_iGp4QjM17_0),.din(w_dff_A_VF4oUAvq4_0),.clk(gclk));
	jdff dff_A_uB9kAt2B0_0(.dout(w_dff_A_VF4oUAvq4_0),.din(w_dff_A_uB9kAt2B0_0),.clk(gclk));
	jdff dff_A_Afu5Kpga3_2(.dout(w_G97_1[2]),.din(w_dff_A_Afu5Kpga3_2),.clk(gclk));
	jdff dff_A_MERfyLJc9_2(.dout(w_dff_A_Afu5Kpga3_2),.din(w_dff_A_MERfyLJc9_2),.clk(gclk));
	jdff dff_A_6TTriCEI5_2(.dout(w_dff_A_MERfyLJc9_2),.din(w_dff_A_6TTriCEI5_2),.clk(gclk));
	jdff dff_A_9oPM0F8E6_2(.dout(w_dff_A_6TTriCEI5_2),.din(w_dff_A_9oPM0F8E6_2),.clk(gclk));
	jdff dff_A_b8Aotwq21_1(.dout(w_G97_0[1]),.din(w_dff_A_b8Aotwq21_1),.clk(gclk));
	jdff dff_A_ALhdn8qc6_1(.dout(w_dff_A_b8Aotwq21_1),.din(w_dff_A_ALhdn8qc6_1),.clk(gclk));
	jdff dff_A_C9em7tj81_1(.dout(w_dff_A_ALhdn8qc6_1),.din(w_dff_A_C9em7tj81_1),.clk(gclk));
	jdff dff_A_8qEqV5IG1_2(.dout(w_G97_0[2]),.din(w_dff_A_8qEqV5IG1_2),.clk(gclk));
	jdff dff_A_fxc072rn5_0(.dout(w_G33_10[0]),.din(w_dff_A_fxc072rn5_0),.clk(gclk));
	jdff dff_A_uZz1fQBT7_1(.dout(w_G33_10[1]),.din(w_dff_A_uZz1fQBT7_1),.clk(gclk));
	jdff dff_A_4Ouj8ThX9_0(.dout(w_n170_0[0]),.din(w_dff_A_4Ouj8ThX9_0),.clk(gclk));
	jdff dff_B_2Q9ieLS33_0(.din(n169),.dout(w_dff_B_2Q9ieLS33_0),.clk(gclk));
	jdff dff_A_PoliPYxD4_0(.dout(w_G274_0[0]),.din(w_dff_A_PoliPYxD4_0),.clk(gclk));
	jdff dff_A_YQsvCYYk7_0(.dout(w_dff_A_PoliPYxD4_0),.din(w_dff_A_YQsvCYYk7_0),.clk(gclk));
	jdff dff_A_coUzNFjU0_0(.dout(w_dff_A_YQsvCYYk7_0),.din(w_dff_A_coUzNFjU0_0),.clk(gclk));
	jdff dff_A_0eV7BkGz8_2(.dout(w_G274_0[2]),.din(w_dff_A_0eV7BkGz8_2),.clk(gclk));
	jdff dff_A_5BzSVzfU8_2(.dout(w_dff_A_0eV7BkGz8_2),.din(w_dff_A_5BzSVzfU8_2),.clk(gclk));
	jdff dff_A_UAPhG3Vn9_0(.dout(w_n166_3[0]),.din(w_dff_A_UAPhG3Vn9_0),.clk(gclk));
	jdff dff_B_WYnzbP1T3_0(.din(n165),.dout(w_dff_B_WYnzbP1T3_0),.clk(gclk));
	jdff dff_A_vtqn6Ngn9_2(.dout(w_n115_0[2]),.din(w_dff_A_vtqn6Ngn9_2),.clk(gclk));
	jdff dff_A_NG8iqZFU6_0(.dout(w_n114_1[0]),.din(w_dff_A_NG8iqZFU6_0),.clk(gclk));
	jdff dff_A_FoBBaqwL2_1(.dout(w_n114_0[1]),.din(w_dff_A_FoBBaqwL2_1),.clk(gclk));
	jdff dff_A_hTYt0Sei3_0(.dout(w_n163_0[0]),.din(w_dff_A_hTYt0Sei3_0),.clk(gclk));
	jdff dff_A_USztoXLK7_2(.dout(w_n161_0[2]),.din(w_dff_A_USztoXLK7_2),.clk(gclk));
	jdff dff_A_Xy8ZZeI59_2(.dout(w_dff_A_USztoXLK7_2),.din(w_dff_A_Xy8ZZeI59_2),.clk(gclk));
	jdff dff_A_pIExNAhw0_2(.dout(w_dff_A_Xy8ZZeI59_2),.din(w_dff_A_pIExNAhw0_2),.clk(gclk));
	jdff dff_A_ZxELQh9I5_0(.dout(w_G45_1[0]),.din(w_dff_A_ZxELQh9I5_0),.clk(gclk));
	jdff dff_A_CO9EWdaC6_0(.dout(w_dff_A_ZxELQh9I5_0),.din(w_dff_A_CO9EWdaC6_0),.clk(gclk));
	jdff dff_A_GFDKQ38K5_1(.dout(w_G45_1[1]),.din(w_dff_A_GFDKQ38K5_1),.clk(gclk));
	jdff dff_A_tEVBWGW62_1(.dout(w_G45_0[1]),.din(w_dff_A_tEVBWGW62_1),.clk(gclk));
	jdff dff_A_qrTS6Gwh7_1(.dout(w_dff_A_tEVBWGW62_1),.din(w_dff_A_qrTS6Gwh7_1),.clk(gclk));
	jdff dff_A_yQTxWFRA1_1(.dout(w_dff_A_qrTS6Gwh7_1),.din(w_dff_A_yQTxWFRA1_1),.clk(gclk));
	jdff dff_A_bV0VerXU7_2(.dout(w_G45_0[2]),.din(w_dff_A_bV0VerXU7_2),.clk(gclk));
	jdff dff_A_TRFGqDUJ8_2(.dout(w_dff_A_bV0VerXU7_2),.din(w_dff_A_TRFGqDUJ8_2),.clk(gclk));
	jdff dff_A_UYUfUEAd4_2(.dout(w_dff_A_TRFGqDUJ8_2),.din(w_dff_A_UYUfUEAd4_2),.clk(gclk));
	jdff dff_A_hEPKzEzv3_0(.dout(w_n98_1[0]),.din(w_dff_A_hEPKzEzv3_0),.clk(gclk));
	jdff dff_A_KVIzA3Ct9_1(.dout(w_n98_1[1]),.din(w_dff_A_KVIzA3Ct9_1),.clk(gclk));
	jdff dff_A_LFyYcmB27_0(.dout(w_G250_0[0]),.din(w_dff_A_LFyYcmB27_0),.clk(gclk));
	jdff dff_A_0Dr2K6jL4_0(.dout(w_dff_A_LFyYcmB27_0),.din(w_dff_A_0Dr2K6jL4_0),.clk(gclk));
	jdff dff_A_rZmdm5qG0_1(.dout(w_G250_0[1]),.din(w_dff_A_rZmdm5qG0_1),.clk(gclk));
	jdff dff_A_c67gaj6g8_1(.dout(w_dff_A_rZmdm5qG0_1),.din(w_dff_A_c67gaj6g8_1),.clk(gclk));
	jdff dff_B_GRNElknY8_1(.din(n153),.dout(w_dff_B_GRNElknY8_1),.clk(gclk));
	jdff dff_A_9ww3VlH63_0(.dout(w_n157_0[0]),.din(w_dff_A_9ww3VlH63_0),.clk(gclk));
	jdff dff_A_GHAbKBh17_0(.dout(w_dff_A_9ww3VlH63_0),.din(w_dff_A_GHAbKBh17_0),.clk(gclk));
	jdff dff_A_DQKieqpc6_2(.dout(w_n157_0[2]),.din(w_dff_A_DQKieqpc6_2),.clk(gclk));
	jdff dff_A_tcKA3BhQ5_2(.dout(w_dff_A_DQKieqpc6_2),.din(w_dff_A_tcKA3BhQ5_2),.clk(gclk));
	jdff dff_A_ydHFQ62C3_1(.dout(w_G116_1[1]),.din(w_dff_A_ydHFQ62C3_1),.clk(gclk));
	jdff dff_A_WHghHJm77_1(.dout(w_dff_A_ydHFQ62C3_1),.din(w_dff_A_WHghHJm77_1),.clk(gclk));
	jdff dff_A_raVhjKGT5_1(.dout(w_dff_A_WHghHJm77_1),.din(w_dff_A_raVhjKGT5_1),.clk(gclk));
	jdff dff_A_ktoydHJt5_2(.dout(w_G116_1[2]),.din(w_dff_A_ktoydHJt5_2),.clk(gclk));
	jdff dff_A_Ar3Xl1TE6_2(.dout(w_dff_A_ktoydHJt5_2),.din(w_dff_A_Ar3Xl1TE6_2),.clk(gclk));
	jdff dff_A_pzus6SVP7_2(.dout(w_dff_A_Ar3Xl1TE6_2),.din(w_dff_A_pzus6SVP7_2),.clk(gclk));
	jdff dff_A_fglkHkid8_1(.dout(w_G116_0[1]),.din(w_dff_A_fglkHkid8_1),.clk(gclk));
	jdff dff_A_UpmNlgzu2_1(.dout(w_dff_A_fglkHkid8_1),.din(w_dff_A_UpmNlgzu2_1),.clk(gclk));
	jdff dff_A_6sEZr79Z9_1(.dout(w_dff_A_UpmNlgzu2_1),.din(w_dff_A_6sEZr79Z9_1),.clk(gclk));
	jdff dff_A_JUzIhdWg1_2(.dout(w_G116_0[2]),.din(w_dff_A_JUzIhdWg1_2),.clk(gclk));
	jdff dff_A_TBnhXvjT5_0(.dout(w_G238_1[0]),.din(w_dff_A_TBnhXvjT5_0),.clk(gclk));
	jdff dff_A_303rdBsU8_0(.dout(w_dff_A_TBnhXvjT5_0),.din(w_dff_A_303rdBsU8_0),.clk(gclk));
	jdff dff_A_hukRPu1H1_1(.dout(w_G238_0[1]),.din(w_dff_A_hukRPu1H1_1),.clk(gclk));
	jdff dff_A_f3QAmBdV4_1(.dout(w_dff_A_hukRPu1H1_1),.din(w_dff_A_f3QAmBdV4_1),.clk(gclk));
	jdff dff_A_XCrtveZf8_1(.dout(w_dff_A_f3QAmBdV4_1),.din(w_dff_A_XCrtveZf8_1),.clk(gclk));
	jdff dff_A_pJc5Nymd0_1(.dout(w_dff_A_XCrtveZf8_1),.din(w_dff_A_pJc5Nymd0_1),.clk(gclk));
	jdff dff_A_zPI9h0pG0_2(.dout(w_G238_0[2]),.din(w_dff_A_zPI9h0pG0_2),.clk(gclk));
	jdff dff_A_9N91VHxD5_2(.dout(w_dff_A_zPI9h0pG0_2),.din(w_dff_A_9N91VHxD5_2),.clk(gclk));
	jdff dff_A_Mlfa3Jcp5_2(.dout(w_G1698_0[2]),.din(w_dff_A_Mlfa3Jcp5_2),.clk(gclk));
	jdff dff_A_Z0cjFDHq7_0(.dout(w_G244_1[0]),.din(w_dff_A_Z0cjFDHq7_0),.clk(gclk));
	jdff dff_A_oHNNeNEI2_0(.dout(w_dff_A_Z0cjFDHq7_0),.din(w_dff_A_oHNNeNEI2_0),.clk(gclk));
	jdff dff_A_06D0wKbJ5_1(.dout(w_G244_0[1]),.din(w_dff_A_06D0wKbJ5_1),.clk(gclk));
	jdff dff_A_6nObsZ5H3_1(.dout(w_dff_A_06D0wKbJ5_1),.din(w_dff_A_6nObsZ5H3_1),.clk(gclk));
	jdff dff_A_lJ3aMjpq8_1(.dout(w_dff_A_6nObsZ5H3_1),.din(w_dff_A_lJ3aMjpq8_1),.clk(gclk));
	jdff dff_A_iaPOG52y2_1(.dout(w_dff_A_lJ3aMjpq8_1),.din(w_dff_A_iaPOG52y2_1),.clk(gclk));
	jdff dff_A_4o0p8slk3_2(.dout(w_G244_0[2]),.din(w_dff_A_4o0p8slk3_2),.clk(gclk));
	jdff dff_A_bj6XxWiH2_2(.dout(w_dff_A_4o0p8slk3_2),.din(w_dff_A_bj6XxWiH2_2),.clk(gclk));
	jdff dff_A_ppGTzq2G7_2(.dout(w_n151_4[2]),.din(w_dff_A_ppGTzq2G7_2),.clk(gclk));
	jdff dff_A_upYG8lUr4_2(.dout(w_dff_A_ppGTzq2G7_2),.din(w_dff_A_upYG8lUr4_2),.clk(gclk));
	jdff dff_A_rYRdCdk93_1(.dout(w_n151_1[1]),.din(w_dff_A_rYRdCdk93_1),.clk(gclk));
	jdff dff_A_kDyzheB88_1(.dout(w_dff_A_rYRdCdk93_1),.din(w_dff_A_kDyzheB88_1),.clk(gclk));
	jdff dff_A_eRcHLr176_2(.dout(w_n151_1[2]),.din(w_dff_A_eRcHLr176_2),.clk(gclk));
	jdff dff_A_EWytyrHp6_2(.dout(w_dff_A_eRcHLr176_2),.din(w_dff_A_EWytyrHp6_2),.clk(gclk));
	jdff dff_A_FJazkNfU9_1(.dout(w_n151_0[1]),.din(w_dff_A_FJazkNfU9_1),.clk(gclk));
	jdff dff_A_bZl15ToZ9_1(.dout(w_dff_A_FJazkNfU9_1),.din(w_dff_A_bZl15ToZ9_1),.clk(gclk));
	jdff dff_A_sgKsKajD0_0(.dout(w_n149_2[0]),.din(w_dff_A_sgKsKajD0_0),.clk(gclk));
	jdff dff_A_eheZoAGo8_1(.dout(w_G41_0[1]),.din(w_dff_A_eheZoAGo8_1),.clk(gclk));
	jdff dff_A_HgYY2dUb4_2(.dout(w_G41_0[2]),.din(w_dff_A_HgYY2dUb4_2),.clk(gclk));
	jdff dff_A_AH0KJFDU0_2(.dout(w_dff_A_HgYY2dUb4_2),.din(w_dff_A_AH0KJFDU0_2),.clk(gclk));
	jdff dff_A_a3mhyjEm2_2(.dout(w_G33_3[2]),.din(w_dff_A_a3mhyjEm2_2),.clk(gclk));
	jdff dff_A_inB6gsfz0_2(.dout(w_dff_A_a3mhyjEm2_2),.din(w_dff_A_inB6gsfz0_2),.clk(gclk));
	jdff dff_A_ogfXx8KF4_2(.dout(w_dff_A_inB6gsfz0_2),.din(w_dff_A_ogfXx8KF4_2),.clk(gclk));
	jdff dff_A_a59X2VON1_2(.dout(w_dff_A_ogfXx8KF4_2),.din(w_dff_A_a59X2VON1_2),.clk(gclk));
	jdff dff_A_8qgATIe62_2(.dout(w_dff_A_a59X2VON1_2),.din(w_dff_A_8qgATIe62_2),.clk(gclk));
	jdff dff_A_KPWEOBb32_0(.dout(w_G33_0[0]),.din(w_dff_A_KPWEOBb32_0),.clk(gclk));
	jdff dff_A_slPEs5cW2_1(.dout(w_n147_0[1]),.din(w_dff_A_slPEs5cW2_1),.clk(gclk));
	jdff dff_A_PQfOk9nx5_2(.dout(w_n147_0[2]),.din(w_dff_A_PQfOk9nx5_2),.clk(gclk));
	jdff dff_A_pLbnh99t5_1(.dout(w_G13_0[1]),.din(w_dff_A_pLbnh99t5_1),.clk(gclk));
	jdff dff_A_4bLfR68l3_2(.dout(w_G13_0[2]),.din(w_dff_A_4bLfR68l3_2),.clk(gclk));
	jdff dff_A_0eRuYOQO3_2(.dout(w_dff_A_4bLfR68l3_2),.din(w_dff_A_0eRuYOQO3_2),.clk(gclk));
	jdff dff_A_3nvoBC4Z2_0(.dout(w_G1_2[0]),.din(w_dff_A_3nvoBC4Z2_0),.clk(gclk));
	jdff dff_A_O3PSfUPA3_2(.dout(w_G1_2[2]),.din(w_dff_A_O3PSfUPA3_2),.clk(gclk));
	jdff dff_A_iAdXw7Hj8_0(.dout(w_G1_0[0]),.din(w_dff_A_iAdXw7Hj8_0),.clk(gclk));
	jdff dff_A_YK0gGx2Z1_1(.dout(w_n146_0[1]),.din(w_dff_A_YK0gGx2Z1_1),.clk(gclk));
	jdff dff_A_EA9FYDxy9_1(.dout(w_dff_A_YK0gGx2Z1_1),.din(w_dff_A_EA9FYDxy9_1),.clk(gclk));
	jdff dff_A_l0bbccIh9_1(.dout(w_dff_A_EA9FYDxy9_1),.din(w_dff_A_l0bbccIh9_1),.clk(gclk));
	jdff dff_A_quvSuv8u5_1(.dout(w_dff_A_l0bbccIh9_1),.din(w_dff_A_quvSuv8u5_1),.clk(gclk));
	jdff dff_A_xsBHwhZ30_1(.dout(w_dff_A_quvSuv8u5_1),.din(w_dff_A_xsBHwhZ30_1),.clk(gclk));
	jdff dff_A_m8wv256D9_1(.dout(w_dff_A_xsBHwhZ30_1),.din(w_dff_A_m8wv256D9_1),.clk(gclk));
	jdff dff_A_UBBdH3Pi7_2(.dout(w_n146_0[2]),.din(w_dff_A_UBBdH3Pi7_2),.clk(gclk));
	jdff dff_A_awll7jxE2_2(.dout(w_dff_A_UBBdH3Pi7_2),.din(w_dff_A_awll7jxE2_2),.clk(gclk));
	jdff dff_A_PpQpP64P8_2(.dout(w_dff_A_awll7jxE2_2),.din(w_dff_A_PpQpP64P8_2),.clk(gclk));
	jdff dff_A_VsF606or9_2(.dout(w_dff_A_PpQpP64P8_2),.din(w_dff_A_VsF606or9_2),.clk(gclk));
	jdff dff_A_9tTkdQcL6_2(.dout(w_dff_A_VsF606or9_2),.din(w_dff_A_9tTkdQcL6_2),.clk(gclk));
	jdff dff_A_fLtmlSke3_2(.dout(w_dff_A_9tTkdQcL6_2),.din(w_dff_A_fLtmlSke3_2),.clk(gclk));
	jdff dff_A_SDNStn4c4_0(.dout(w_G169_1[0]),.din(w_dff_A_SDNStn4c4_0),.clk(gclk));
	jdff dff_A_GM2LTRIx2_0(.dout(w_dff_A_SDNStn4c4_0),.din(w_dff_A_GM2LTRIx2_0),.clk(gclk));
	jdff dff_A_sLGr2W334_0(.dout(w_dff_A_GM2LTRIx2_0),.din(w_dff_A_sLGr2W334_0),.clk(gclk));
	jdff dff_A_hdZFUim10_0(.dout(w_dff_A_sLGr2W334_0),.din(w_dff_A_hdZFUim10_0),.clk(gclk));
	jdff dff_A_6ZgD6zws4_0(.dout(w_dff_A_hdZFUim10_0),.din(w_dff_A_6ZgD6zws4_0),.clk(gclk));
	jdff dff_A_Hn2rZI4c7_0(.dout(w_dff_A_6ZgD6zws4_0),.din(w_dff_A_Hn2rZI4c7_0),.clk(gclk));
	jdff dff_A_G6PyO8im8_0(.dout(w_dff_A_Hn2rZI4c7_0),.din(w_dff_A_G6PyO8im8_0),.clk(gclk));
	jdff dff_A_BTJJSqX32_1(.dout(w_G169_0[1]),.din(w_dff_A_BTJJSqX32_1),.clk(gclk));
	jdff dff_A_76qXpSFo4_1(.dout(w_dff_A_BTJJSqX32_1),.din(w_dff_A_76qXpSFo4_1),.clk(gclk));
	jdff dff_A_SXKzKZXg9_1(.dout(w_dff_A_76qXpSFo4_1),.din(w_dff_A_SXKzKZXg9_1),.clk(gclk));
	jdff dff_A_gcq7ZLJ48_1(.dout(w_dff_A_SXKzKZXg9_1),.din(w_dff_A_gcq7ZLJ48_1),.clk(gclk));
	jdff dff_A_5YOTw2ai0_1(.dout(w_dff_A_gcq7ZLJ48_1),.din(w_dff_A_5YOTw2ai0_1),.clk(gclk));
	jdff dff_A_cNWazVGD3_1(.dout(w_dff_A_5YOTw2ai0_1),.din(w_dff_A_cNWazVGD3_1),.clk(gclk));
	jdff dff_A_73xXv1qJ4_1(.dout(w_dff_A_cNWazVGD3_1),.din(w_dff_A_73xXv1qJ4_1),.clk(gclk));
	jdff dff_A_jZlf7qoN7_2(.dout(w_G169_0[2]),.din(w_dff_A_jZlf7qoN7_2),.clk(gclk));
	jdff dff_A_FLMG89st7_2(.dout(w_dff_A_jZlf7qoN7_2),.din(w_dff_A_FLMG89st7_2),.clk(gclk));
	jdff dff_A_6mrcnqob9_2(.dout(w_dff_A_FLMG89st7_2),.din(w_dff_A_6mrcnqob9_2),.clk(gclk));
	jdff dff_A_myXmhWVs2_2(.dout(w_dff_A_6mrcnqob9_2),.din(w_dff_A_myXmhWVs2_2),.clk(gclk));
	jdff dff_A_PWB9Dwhw3_2(.dout(w_dff_A_myXmhWVs2_2),.din(w_dff_A_PWB9Dwhw3_2),.clk(gclk));
	jdff dff_A_YxIiNnCT8_2(.dout(w_dff_A_PWB9Dwhw3_2),.din(w_dff_A_YxIiNnCT8_2),.clk(gclk));
	jdff dff_A_QuWBZkPP5_2(.dout(w_dff_A_YxIiNnCT8_2),.din(w_dff_A_QuWBZkPP5_2),.clk(gclk));
	jdff dff_A_jDDyjmOM9_2(.dout(w_dff_A_oCeIctIc4_0),.din(w_dff_A_jDDyjmOM9_2),.clk(gclk));
	jdff dff_A_oCeIctIc4_0(.dout(w_dff_A_yTGtcVRg0_0),.din(w_dff_A_oCeIctIc4_0),.clk(gclk));
	jdff dff_A_yTGtcVRg0_0(.dout(w_dff_A_8JwgpaaC9_0),.din(w_dff_A_yTGtcVRg0_0),.clk(gclk));
	jdff dff_A_8JwgpaaC9_0(.dout(w_dff_A_bPrcsCRS4_0),.din(w_dff_A_8JwgpaaC9_0),.clk(gclk));
	jdff dff_A_bPrcsCRS4_0(.dout(w_dff_A_XEUnkOtK1_0),.din(w_dff_A_bPrcsCRS4_0),.clk(gclk));
	jdff dff_A_XEUnkOtK1_0(.dout(w_dff_A_04jcxYzU7_0),.din(w_dff_A_XEUnkOtK1_0),.clk(gclk));
	jdff dff_A_04jcxYzU7_0(.dout(w_dff_A_ou87bcHz4_0),.din(w_dff_A_04jcxYzU7_0),.clk(gclk));
	jdff dff_A_ou87bcHz4_0(.dout(w_dff_A_qtcryspU0_0),.din(w_dff_A_ou87bcHz4_0),.clk(gclk));
	jdff dff_A_qtcryspU0_0(.dout(w_dff_A_ja7F6qH94_0),.din(w_dff_A_qtcryspU0_0),.clk(gclk));
	jdff dff_A_ja7F6qH94_0(.dout(w_dff_A_FE7Sq7Tl2_0),.din(w_dff_A_ja7F6qH94_0),.clk(gclk));
	jdff dff_A_FE7Sq7Tl2_0(.dout(w_dff_A_Vdc5lXXl2_0),.din(w_dff_A_FE7Sq7Tl2_0),.clk(gclk));
	jdff dff_A_Vdc5lXXl2_0(.dout(w_dff_A_0TUAKMoS1_0),.din(w_dff_A_Vdc5lXXl2_0),.clk(gclk));
	jdff dff_A_0TUAKMoS1_0(.dout(w_dff_A_sO0ezfUK2_0),.din(w_dff_A_0TUAKMoS1_0),.clk(gclk));
	jdff dff_A_sO0ezfUK2_0(.dout(w_dff_A_Py8YTI9G5_0),.din(w_dff_A_sO0ezfUK2_0),.clk(gclk));
	jdff dff_A_Py8YTI9G5_0(.dout(w_dff_A_XHUR7MiC5_0),.din(w_dff_A_Py8YTI9G5_0),.clk(gclk));
	jdff dff_A_XHUR7MiC5_0(.dout(w_dff_A_W46RsyYx0_0),.din(w_dff_A_XHUR7MiC5_0),.clk(gclk));
	jdff dff_A_W46RsyYx0_0(.dout(w_dff_A_NbxblaA19_0),.din(w_dff_A_W46RsyYx0_0),.clk(gclk));
	jdff dff_A_NbxblaA19_0(.dout(w_dff_A_MQoacw8Q9_0),.din(w_dff_A_NbxblaA19_0),.clk(gclk));
	jdff dff_A_MQoacw8Q9_0(.dout(w_dff_A_LAqLvMI30_0),.din(w_dff_A_MQoacw8Q9_0),.clk(gclk));
	jdff dff_A_LAqLvMI30_0(.dout(w_dff_A_mkE7Z8ts0_0),.din(w_dff_A_LAqLvMI30_0),.clk(gclk));
	jdff dff_A_mkE7Z8ts0_0(.dout(w_dff_A_46Ybfo041_0),.din(w_dff_A_mkE7Z8ts0_0),.clk(gclk));
	jdff dff_A_46Ybfo041_0(.dout(w_dff_A_HGzp22941_0),.din(w_dff_A_46Ybfo041_0),.clk(gclk));
	jdff dff_A_HGzp22941_0(.dout(w_dff_A_PFGQIOju3_0),.din(w_dff_A_HGzp22941_0),.clk(gclk));
	jdff dff_A_PFGQIOju3_0(.dout(w_dff_A_ihUofMly6_0),.din(w_dff_A_PFGQIOju3_0),.clk(gclk));
	jdff dff_A_ihUofMly6_0(.dout(G353),.din(w_dff_A_ihUofMly6_0),.clk(gclk));
	jdff dff_A_b4JJi3Xo9_1(.dout(w_dff_A_3D80Yf1i6_0),.din(w_dff_A_b4JJi3Xo9_1),.clk(gclk));
	jdff dff_A_3D80Yf1i6_0(.dout(w_dff_A_5nhhep6d9_0),.din(w_dff_A_3D80Yf1i6_0),.clk(gclk));
	jdff dff_A_5nhhep6d9_0(.dout(w_dff_A_0thdKQix0_0),.din(w_dff_A_5nhhep6d9_0),.clk(gclk));
	jdff dff_A_0thdKQix0_0(.dout(w_dff_A_4ge9LgrV4_0),.din(w_dff_A_0thdKQix0_0),.clk(gclk));
	jdff dff_A_4ge9LgrV4_0(.dout(w_dff_A_wKJWkuGj9_0),.din(w_dff_A_4ge9LgrV4_0),.clk(gclk));
	jdff dff_A_wKJWkuGj9_0(.dout(w_dff_A_aI3kkDP84_0),.din(w_dff_A_wKJWkuGj9_0),.clk(gclk));
	jdff dff_A_aI3kkDP84_0(.dout(w_dff_A_XA72lHkS1_0),.din(w_dff_A_aI3kkDP84_0),.clk(gclk));
	jdff dff_A_XA72lHkS1_0(.dout(w_dff_A_jsIA8eKB8_0),.din(w_dff_A_XA72lHkS1_0),.clk(gclk));
	jdff dff_A_jsIA8eKB8_0(.dout(w_dff_A_c60NlIbj0_0),.din(w_dff_A_jsIA8eKB8_0),.clk(gclk));
	jdff dff_A_c60NlIbj0_0(.dout(w_dff_A_2ewcdiOT9_0),.din(w_dff_A_c60NlIbj0_0),.clk(gclk));
	jdff dff_A_2ewcdiOT9_0(.dout(w_dff_A_2VzzZEfu5_0),.din(w_dff_A_2ewcdiOT9_0),.clk(gclk));
	jdff dff_A_2VzzZEfu5_0(.dout(w_dff_A_XSxjnDbD9_0),.din(w_dff_A_2VzzZEfu5_0),.clk(gclk));
	jdff dff_A_XSxjnDbD9_0(.dout(w_dff_A_mzsI8NCp0_0),.din(w_dff_A_XSxjnDbD9_0),.clk(gclk));
	jdff dff_A_mzsI8NCp0_0(.dout(w_dff_A_uxR2QE8v0_0),.din(w_dff_A_mzsI8NCp0_0),.clk(gclk));
	jdff dff_A_uxR2QE8v0_0(.dout(w_dff_A_A9gopoxK0_0),.din(w_dff_A_uxR2QE8v0_0),.clk(gclk));
	jdff dff_A_A9gopoxK0_0(.dout(w_dff_A_mHTJaAdx4_0),.din(w_dff_A_A9gopoxK0_0),.clk(gclk));
	jdff dff_A_mHTJaAdx4_0(.dout(w_dff_A_GCl3sPpe3_0),.din(w_dff_A_mHTJaAdx4_0),.clk(gclk));
	jdff dff_A_GCl3sPpe3_0(.dout(w_dff_A_Hl1KhlD93_0),.din(w_dff_A_GCl3sPpe3_0),.clk(gclk));
	jdff dff_A_Hl1KhlD93_0(.dout(w_dff_A_k5zRfPFm4_0),.din(w_dff_A_Hl1KhlD93_0),.clk(gclk));
	jdff dff_A_k5zRfPFm4_0(.dout(w_dff_A_JyflBbLh1_0),.din(w_dff_A_k5zRfPFm4_0),.clk(gclk));
	jdff dff_A_JyflBbLh1_0(.dout(w_dff_A_oyZYblEz3_0),.din(w_dff_A_JyflBbLh1_0),.clk(gclk));
	jdff dff_A_oyZYblEz3_0(.dout(w_dff_A_gWKpw2w06_0),.din(w_dff_A_oyZYblEz3_0),.clk(gclk));
	jdff dff_A_gWKpw2w06_0(.dout(w_dff_A_yunia8tt0_0),.din(w_dff_A_gWKpw2w06_0),.clk(gclk));
	jdff dff_A_yunia8tt0_0(.dout(G355),.din(w_dff_A_yunia8tt0_0),.clk(gclk));
	jdff dff_A_yu2mnwg27_2(.dout(w_dff_A_bPEi8vwn8_0),.din(w_dff_A_yu2mnwg27_2),.clk(gclk));
	jdff dff_A_bPEi8vwn8_0(.dout(w_dff_A_lGzCx7Df2_0),.din(w_dff_A_bPEi8vwn8_0),.clk(gclk));
	jdff dff_A_lGzCx7Df2_0(.dout(w_dff_A_mCSCtIhU9_0),.din(w_dff_A_lGzCx7Df2_0),.clk(gclk));
	jdff dff_A_mCSCtIhU9_0(.dout(w_dff_A_sMl3qcMf6_0),.din(w_dff_A_mCSCtIhU9_0),.clk(gclk));
	jdff dff_A_sMl3qcMf6_0(.dout(w_dff_A_ypir7DjH3_0),.din(w_dff_A_sMl3qcMf6_0),.clk(gclk));
	jdff dff_A_ypir7DjH3_0(.dout(w_dff_A_rPmcsS9X7_0),.din(w_dff_A_ypir7DjH3_0),.clk(gclk));
	jdff dff_A_rPmcsS9X7_0(.dout(w_dff_A_eFcD9XJe2_0),.din(w_dff_A_rPmcsS9X7_0),.clk(gclk));
	jdff dff_A_eFcD9XJe2_0(.dout(w_dff_A_fLrCvENM3_0),.din(w_dff_A_eFcD9XJe2_0),.clk(gclk));
	jdff dff_A_fLrCvENM3_0(.dout(w_dff_A_gqOq2OKz3_0),.din(w_dff_A_fLrCvENM3_0),.clk(gclk));
	jdff dff_A_gqOq2OKz3_0(.dout(w_dff_A_LSXYNV9I7_0),.din(w_dff_A_gqOq2OKz3_0),.clk(gclk));
	jdff dff_A_LSXYNV9I7_0(.dout(w_dff_A_GgQZkZ8N0_0),.din(w_dff_A_LSXYNV9I7_0),.clk(gclk));
	jdff dff_A_GgQZkZ8N0_0(.dout(w_dff_A_MUil1Pu22_0),.din(w_dff_A_GgQZkZ8N0_0),.clk(gclk));
	jdff dff_A_MUil1Pu22_0(.dout(w_dff_A_F7PTQD1p0_0),.din(w_dff_A_MUil1Pu22_0),.clk(gclk));
	jdff dff_A_F7PTQD1p0_0(.dout(w_dff_A_LCwPXFQN8_0),.din(w_dff_A_F7PTQD1p0_0),.clk(gclk));
	jdff dff_A_LCwPXFQN8_0(.dout(w_dff_A_igeNho1x0_0),.din(w_dff_A_LCwPXFQN8_0),.clk(gclk));
	jdff dff_A_igeNho1x0_0(.dout(w_dff_A_2j63eibE7_0),.din(w_dff_A_igeNho1x0_0),.clk(gclk));
	jdff dff_A_2j63eibE7_0(.dout(w_dff_A_6z13bnug1_0),.din(w_dff_A_2j63eibE7_0),.clk(gclk));
	jdff dff_A_6z13bnug1_0(.dout(w_dff_A_h1nEpwY53_0),.din(w_dff_A_6z13bnug1_0),.clk(gclk));
	jdff dff_A_h1nEpwY53_0(.dout(w_dff_A_CLRBlX9P2_0),.din(w_dff_A_h1nEpwY53_0),.clk(gclk));
	jdff dff_A_CLRBlX9P2_0(.dout(w_dff_A_hyFJq4Tp4_0),.din(w_dff_A_CLRBlX9P2_0),.clk(gclk));
	jdff dff_A_hyFJq4Tp4_0(.dout(G361),.din(w_dff_A_hyFJq4Tp4_0),.clk(gclk));
	jdff dff_A_KxktjB0M1_2(.dout(w_dff_A_ETfMRraI8_0),.din(w_dff_A_KxktjB0M1_2),.clk(gclk));
	jdff dff_A_ETfMRraI8_0(.dout(w_dff_A_i5LiCjT30_0),.din(w_dff_A_ETfMRraI8_0),.clk(gclk));
	jdff dff_A_i5LiCjT30_0(.dout(w_dff_A_b7GGSp3J5_0),.din(w_dff_A_i5LiCjT30_0),.clk(gclk));
	jdff dff_A_b7GGSp3J5_0(.dout(w_dff_A_YLwcEg3v9_0),.din(w_dff_A_b7GGSp3J5_0),.clk(gclk));
	jdff dff_A_YLwcEg3v9_0(.dout(w_dff_A_S8gd0K6y9_0),.din(w_dff_A_YLwcEg3v9_0),.clk(gclk));
	jdff dff_A_S8gd0K6y9_0(.dout(w_dff_A_AJsGT4HC7_0),.din(w_dff_A_S8gd0K6y9_0),.clk(gclk));
	jdff dff_A_AJsGT4HC7_0(.dout(w_dff_A_M1uryMSr8_0),.din(w_dff_A_AJsGT4HC7_0),.clk(gclk));
	jdff dff_A_M1uryMSr8_0(.dout(w_dff_A_kbFLxLLY1_0),.din(w_dff_A_M1uryMSr8_0),.clk(gclk));
	jdff dff_A_kbFLxLLY1_0(.dout(w_dff_A_7xcccwWZ0_0),.din(w_dff_A_kbFLxLLY1_0),.clk(gclk));
	jdff dff_A_7xcccwWZ0_0(.dout(w_dff_A_PSGaGukk8_0),.din(w_dff_A_7xcccwWZ0_0),.clk(gclk));
	jdff dff_A_PSGaGukk8_0(.dout(w_dff_A_Aw3cQnog9_0),.din(w_dff_A_PSGaGukk8_0),.clk(gclk));
	jdff dff_A_Aw3cQnog9_0(.dout(w_dff_A_9JTme08A5_0),.din(w_dff_A_Aw3cQnog9_0),.clk(gclk));
	jdff dff_A_9JTme08A5_0(.dout(w_dff_A_JxT0K3Sj4_0),.din(w_dff_A_9JTme08A5_0),.clk(gclk));
	jdff dff_A_JxT0K3Sj4_0(.dout(w_dff_A_XwkblzX26_0),.din(w_dff_A_JxT0K3Sj4_0),.clk(gclk));
	jdff dff_A_XwkblzX26_0(.dout(w_dff_A_PrdI3O528_0),.din(w_dff_A_XwkblzX26_0),.clk(gclk));
	jdff dff_A_PrdI3O528_0(.dout(w_dff_A_GJc1JsfS1_0),.din(w_dff_A_PrdI3O528_0),.clk(gclk));
	jdff dff_A_GJc1JsfS1_0(.dout(w_dff_A_f7inSK2C2_0),.din(w_dff_A_GJc1JsfS1_0),.clk(gclk));
	jdff dff_A_f7inSK2C2_0(.dout(w_dff_A_oglXmj6O5_0),.din(w_dff_A_f7inSK2C2_0),.clk(gclk));
	jdff dff_A_oglXmj6O5_0(.dout(w_dff_A_nyPwmjWf0_0),.din(w_dff_A_oglXmj6O5_0),.clk(gclk));
	jdff dff_A_nyPwmjWf0_0(.dout(w_dff_A_dFuDFUHC4_0),.din(w_dff_A_nyPwmjWf0_0),.clk(gclk));
	jdff dff_A_dFuDFUHC4_0(.dout(w_dff_A_OcB7E4FS6_0),.din(w_dff_A_dFuDFUHC4_0),.clk(gclk));
	jdff dff_A_OcB7E4FS6_0(.dout(w_dff_A_fOdpVXOa1_0),.din(w_dff_A_OcB7E4FS6_0),.clk(gclk));
	jdff dff_A_fOdpVXOa1_0(.dout(w_dff_A_KNTDztRT6_0),.din(w_dff_A_fOdpVXOa1_0),.clk(gclk));
	jdff dff_A_KNTDztRT6_0(.dout(G358),.din(w_dff_A_KNTDztRT6_0),.clk(gclk));
	jdff dff_A_hm8XpUoB1_2(.dout(w_dff_A_N4XF6Hnn0_0),.din(w_dff_A_hm8XpUoB1_2),.clk(gclk));
	jdff dff_A_N4XF6Hnn0_0(.dout(w_dff_A_u2pQx0fr2_0),.din(w_dff_A_N4XF6Hnn0_0),.clk(gclk));
	jdff dff_A_u2pQx0fr2_0(.dout(w_dff_A_f4p5mze87_0),.din(w_dff_A_u2pQx0fr2_0),.clk(gclk));
	jdff dff_A_f4p5mze87_0(.dout(w_dff_A_V7ZJnNfe1_0),.din(w_dff_A_f4p5mze87_0),.clk(gclk));
	jdff dff_A_V7ZJnNfe1_0(.dout(w_dff_A_cBFbio7O4_0),.din(w_dff_A_V7ZJnNfe1_0),.clk(gclk));
	jdff dff_A_cBFbio7O4_0(.dout(w_dff_A_vXZQ5h5j9_0),.din(w_dff_A_cBFbio7O4_0),.clk(gclk));
	jdff dff_A_vXZQ5h5j9_0(.dout(w_dff_A_2S85BXrz9_0),.din(w_dff_A_vXZQ5h5j9_0),.clk(gclk));
	jdff dff_A_2S85BXrz9_0(.dout(w_dff_A_egVfUnC77_0),.din(w_dff_A_2S85BXrz9_0),.clk(gclk));
	jdff dff_A_egVfUnC77_0(.dout(w_dff_A_mgfaHL9H3_0),.din(w_dff_A_egVfUnC77_0),.clk(gclk));
	jdff dff_A_mgfaHL9H3_0(.dout(w_dff_A_TOneLI254_0),.din(w_dff_A_mgfaHL9H3_0),.clk(gclk));
	jdff dff_A_TOneLI254_0(.dout(w_dff_A_k1fWSuVW4_0),.din(w_dff_A_TOneLI254_0),.clk(gclk));
	jdff dff_A_k1fWSuVW4_0(.dout(w_dff_A_o6u0Nn5F9_0),.din(w_dff_A_k1fWSuVW4_0),.clk(gclk));
	jdff dff_A_o6u0Nn5F9_0(.dout(w_dff_A_xyL8Gekh9_0),.din(w_dff_A_o6u0Nn5F9_0),.clk(gclk));
	jdff dff_A_xyL8Gekh9_0(.dout(w_dff_A_Il4rDvRK9_0),.din(w_dff_A_xyL8Gekh9_0),.clk(gclk));
	jdff dff_A_Il4rDvRK9_0(.dout(w_dff_A_bl42ncSb2_0),.din(w_dff_A_Il4rDvRK9_0),.clk(gclk));
	jdff dff_A_bl42ncSb2_0(.dout(w_dff_A_eAyqwCzZ6_0),.din(w_dff_A_bl42ncSb2_0),.clk(gclk));
	jdff dff_A_eAyqwCzZ6_0(.dout(w_dff_A_OC9iKQH58_0),.din(w_dff_A_eAyqwCzZ6_0),.clk(gclk));
	jdff dff_A_OC9iKQH58_0(.dout(w_dff_A_2w8vXaEC5_0),.din(w_dff_A_OC9iKQH58_0),.clk(gclk));
	jdff dff_A_2w8vXaEC5_0(.dout(w_dff_A_hqzYHSbg0_0),.din(w_dff_A_2w8vXaEC5_0),.clk(gclk));
	jdff dff_A_hqzYHSbg0_0(.dout(w_dff_A_VK5lhS117_0),.din(w_dff_A_hqzYHSbg0_0),.clk(gclk));
	jdff dff_A_VK5lhS117_0(.dout(w_dff_A_kqRTBoj71_0),.din(w_dff_A_VK5lhS117_0),.clk(gclk));
	jdff dff_A_kqRTBoj71_0(.dout(w_dff_A_dnWPRKXl7_0),.din(w_dff_A_kqRTBoj71_0),.clk(gclk));
	jdff dff_A_dnWPRKXl7_0(.dout(w_dff_A_XBN2pRht0_0),.din(w_dff_A_dnWPRKXl7_0),.clk(gclk));
	jdff dff_A_XBN2pRht0_0(.dout(G351),.din(w_dff_A_XBN2pRht0_0),.clk(gclk));
	jdff dff_A_Fo7AjoZB3_2(.dout(w_dff_A_3SRJIUlD6_0),.din(w_dff_A_Fo7AjoZB3_2),.clk(gclk));
	jdff dff_A_3SRJIUlD6_0(.dout(w_dff_A_d1Py6wvc5_0),.din(w_dff_A_3SRJIUlD6_0),.clk(gclk));
	jdff dff_A_d1Py6wvc5_0(.dout(w_dff_A_qyS5Wz0A7_0),.din(w_dff_A_d1Py6wvc5_0),.clk(gclk));
	jdff dff_A_qyS5Wz0A7_0(.dout(w_dff_A_XnUb4Zlr3_0),.din(w_dff_A_qyS5Wz0A7_0),.clk(gclk));
	jdff dff_A_XnUb4Zlr3_0(.dout(w_dff_A_issZT9NH3_0),.din(w_dff_A_XnUb4Zlr3_0),.clk(gclk));
	jdff dff_A_issZT9NH3_0(.dout(w_dff_A_CHVGcIuR9_0),.din(w_dff_A_issZT9NH3_0),.clk(gclk));
	jdff dff_A_CHVGcIuR9_0(.dout(w_dff_A_lMKux7055_0),.din(w_dff_A_CHVGcIuR9_0),.clk(gclk));
	jdff dff_A_lMKux7055_0(.dout(w_dff_A_UU5ENAX71_0),.din(w_dff_A_lMKux7055_0),.clk(gclk));
	jdff dff_A_UU5ENAX71_0(.dout(w_dff_A_cAUmK5Mm7_0),.din(w_dff_A_UU5ENAX71_0),.clk(gclk));
	jdff dff_A_cAUmK5Mm7_0(.dout(w_dff_A_zrjxHRTb1_0),.din(w_dff_A_cAUmK5Mm7_0),.clk(gclk));
	jdff dff_A_zrjxHRTb1_0(.dout(w_dff_A_vj5vTeuW9_0),.din(w_dff_A_zrjxHRTb1_0),.clk(gclk));
	jdff dff_A_vj5vTeuW9_0(.dout(w_dff_A_rPyJpGr71_0),.din(w_dff_A_vj5vTeuW9_0),.clk(gclk));
	jdff dff_A_rPyJpGr71_0(.dout(w_dff_A_swsvL5td8_0),.din(w_dff_A_rPyJpGr71_0),.clk(gclk));
	jdff dff_A_swsvL5td8_0(.dout(G372),.din(w_dff_A_swsvL5td8_0),.clk(gclk));
	jdff dff_A_yKE6Pi2p6_2(.dout(w_dff_A_ILl5k9cI5_0),.din(w_dff_A_yKE6Pi2p6_2),.clk(gclk));
	jdff dff_A_ILl5k9cI5_0(.dout(w_dff_A_VOcmU1MJ3_0),.din(w_dff_A_ILl5k9cI5_0),.clk(gclk));
	jdff dff_A_VOcmU1MJ3_0(.dout(w_dff_A_NE5UXxOC0_0),.din(w_dff_A_VOcmU1MJ3_0),.clk(gclk));
	jdff dff_A_NE5UXxOC0_0(.dout(w_dff_A_LPvpTHiz2_0),.din(w_dff_A_NE5UXxOC0_0),.clk(gclk));
	jdff dff_A_LPvpTHiz2_0(.dout(w_dff_A_Q5jFwPwD3_0),.din(w_dff_A_LPvpTHiz2_0),.clk(gclk));
	jdff dff_A_Q5jFwPwD3_0(.dout(w_dff_A_ohcL0so56_0),.din(w_dff_A_Q5jFwPwD3_0),.clk(gclk));
	jdff dff_A_ohcL0so56_0(.dout(w_dff_A_EpvJVHbi5_0),.din(w_dff_A_ohcL0so56_0),.clk(gclk));
	jdff dff_A_EpvJVHbi5_0(.dout(w_dff_A_Hsa47J9Y2_0),.din(w_dff_A_EpvJVHbi5_0),.clk(gclk));
	jdff dff_A_Hsa47J9Y2_0(.dout(w_dff_A_On5sCEYo3_0),.din(w_dff_A_Hsa47J9Y2_0),.clk(gclk));
	jdff dff_A_On5sCEYo3_0(.dout(w_dff_A_Y7PXSUVf4_0),.din(w_dff_A_On5sCEYo3_0),.clk(gclk));
	jdff dff_A_Y7PXSUVf4_0(.dout(w_dff_A_SyK2xPPD8_0),.din(w_dff_A_Y7PXSUVf4_0),.clk(gclk));
	jdff dff_A_SyK2xPPD8_0(.dout(G369),.din(w_dff_A_SyK2xPPD8_0),.clk(gclk));
	jdff dff_A_TMIQp7yB0_2(.dout(w_dff_A_40r01Umj8_0),.din(w_dff_A_TMIQp7yB0_2),.clk(gclk));
	jdff dff_A_40r01Umj8_0(.dout(w_dff_A_sZTAlPqr8_0),.din(w_dff_A_40r01Umj8_0),.clk(gclk));
	jdff dff_A_sZTAlPqr8_0(.dout(w_dff_A_dC2RTqVH5_0),.din(w_dff_A_sZTAlPqr8_0),.clk(gclk));
	jdff dff_A_dC2RTqVH5_0(.dout(w_dff_A_oYxdiuPb2_0),.din(w_dff_A_dC2RTqVH5_0),.clk(gclk));
	jdff dff_A_oYxdiuPb2_0(.dout(w_dff_A_bUqrFaCj4_0),.din(w_dff_A_oYxdiuPb2_0),.clk(gclk));
	jdff dff_A_bUqrFaCj4_0(.dout(w_dff_A_IBhUu7Qm6_0),.din(w_dff_A_bUqrFaCj4_0),.clk(gclk));
	jdff dff_A_IBhUu7Qm6_0(.dout(w_dff_A_wzJh5yps6_0),.din(w_dff_A_IBhUu7Qm6_0),.clk(gclk));
	jdff dff_A_wzJh5yps6_0(.dout(w_dff_A_kYLZHSdZ3_0),.din(w_dff_A_wzJh5yps6_0),.clk(gclk));
	jdff dff_A_kYLZHSdZ3_0(.dout(w_dff_A_hwO46wRc7_0),.din(w_dff_A_kYLZHSdZ3_0),.clk(gclk));
	jdff dff_A_hwO46wRc7_0(.dout(w_dff_A_E7jguRXM1_0),.din(w_dff_A_hwO46wRc7_0),.clk(gclk));
	jdff dff_A_E7jguRXM1_0(.dout(G399),.din(w_dff_A_E7jguRXM1_0),.clk(gclk));
	jdff dff_A_0WVEvPGS5_2(.dout(w_dff_A_bjZscRO61_0),.din(w_dff_A_0WVEvPGS5_2),.clk(gclk));
	jdff dff_A_bjZscRO61_0(.dout(w_dff_A_ipYufpMg8_0),.din(w_dff_A_bjZscRO61_0),.clk(gclk));
	jdff dff_A_ipYufpMg8_0(.dout(w_dff_A_nfIuEa7O8_0),.din(w_dff_A_ipYufpMg8_0),.clk(gclk));
	jdff dff_A_nfIuEa7O8_0(.dout(w_dff_A_WIolRQIE1_0),.din(w_dff_A_nfIuEa7O8_0),.clk(gclk));
	jdff dff_A_WIolRQIE1_0(.dout(w_dff_A_04fPKSR12_0),.din(w_dff_A_WIolRQIE1_0),.clk(gclk));
	jdff dff_A_04fPKSR12_0(.dout(w_dff_A_hblpjV0x7_0),.din(w_dff_A_04fPKSR12_0),.clk(gclk));
	jdff dff_A_hblpjV0x7_0(.dout(w_dff_A_iCJiOi5u8_0),.din(w_dff_A_hblpjV0x7_0),.clk(gclk));
	jdff dff_A_iCJiOi5u8_0(.dout(w_dff_A_j3MvBzGw5_0),.din(w_dff_A_iCJiOi5u8_0),.clk(gclk));
	jdff dff_A_j3MvBzGw5_0(.dout(w_dff_A_x0zfNS5s1_0),.din(w_dff_A_j3MvBzGw5_0),.clk(gclk));
	jdff dff_A_x0zfNS5s1_0(.dout(w_dff_A_eJhMTvLA1_0),.din(w_dff_A_x0zfNS5s1_0),.clk(gclk));
	jdff dff_A_eJhMTvLA1_0(.dout(G364),.din(w_dff_A_eJhMTvLA1_0),.clk(gclk));
	jdff dff_A_JvhgudXb7_2(.dout(w_dff_A_7jU79r5T3_0),.din(w_dff_A_JvhgudXb7_2),.clk(gclk));
	jdff dff_A_7jU79r5T3_0(.dout(w_dff_A_zJMLiDnG9_0),.din(w_dff_A_7jU79r5T3_0),.clk(gclk));
	jdff dff_A_zJMLiDnG9_0(.dout(w_dff_A_fgn35j2M0_0),.din(w_dff_A_zJMLiDnG9_0),.clk(gclk));
	jdff dff_A_fgn35j2M0_0(.dout(w_dff_A_LtUMQUBu0_0),.din(w_dff_A_fgn35j2M0_0),.clk(gclk));
	jdff dff_A_LtUMQUBu0_0(.dout(w_dff_A_hI41J0ac3_0),.din(w_dff_A_LtUMQUBu0_0),.clk(gclk));
	jdff dff_A_hI41J0ac3_0(.dout(w_dff_A_KTddD5ff1_0),.din(w_dff_A_hI41J0ac3_0),.clk(gclk));
	jdff dff_A_KTddD5ff1_0(.dout(w_dff_A_idLnCTGo6_0),.din(w_dff_A_KTddD5ff1_0),.clk(gclk));
	jdff dff_A_idLnCTGo6_0(.dout(w_dff_A_o6sNFGwq7_0),.din(w_dff_A_idLnCTGo6_0),.clk(gclk));
	jdff dff_A_o6sNFGwq7_0(.dout(w_dff_A_yQqCGAVL5_0),.din(w_dff_A_o6sNFGwq7_0),.clk(gclk));
	jdff dff_A_yQqCGAVL5_0(.dout(w_dff_A_SdWRPurT6_0),.din(w_dff_A_yQqCGAVL5_0),.clk(gclk));
	jdff dff_A_SdWRPurT6_0(.dout(G396),.din(w_dff_A_SdWRPurT6_0),.clk(gclk));
	jdff dff_A_MK7puvqH4_1(.dout(w_dff_A_T3sTSkls0_0),.din(w_dff_A_MK7puvqH4_1),.clk(gclk));
	jdff dff_A_T3sTSkls0_0(.dout(w_dff_A_8GJ6RkPC8_0),.din(w_dff_A_T3sTSkls0_0),.clk(gclk));
	jdff dff_A_8GJ6RkPC8_0(.dout(w_dff_A_pZuEXSwI3_0),.din(w_dff_A_8GJ6RkPC8_0),.clk(gclk));
	jdff dff_A_pZuEXSwI3_0(.dout(w_dff_A_Dz2LoSbI3_0),.din(w_dff_A_pZuEXSwI3_0),.clk(gclk));
	jdff dff_A_Dz2LoSbI3_0(.dout(w_dff_A_qeYaqAiR2_0),.din(w_dff_A_Dz2LoSbI3_0),.clk(gclk));
	jdff dff_A_qeYaqAiR2_0(.dout(w_dff_A_KfbbFbyt7_0),.din(w_dff_A_qeYaqAiR2_0),.clk(gclk));
	jdff dff_A_KfbbFbyt7_0(.dout(w_dff_A_dwFfx8zJ1_0),.din(w_dff_A_KfbbFbyt7_0),.clk(gclk));
	jdff dff_A_dwFfx8zJ1_0(.dout(G384),.din(w_dff_A_dwFfx8zJ1_0),.clk(gclk));
	jdff dff_A_OjXgsc6F9_2(.dout(w_dff_A_kItvCpdm3_0),.din(w_dff_A_OjXgsc6F9_2),.clk(gclk));
	jdff dff_A_kItvCpdm3_0(.dout(w_dff_A_NuQSjE8t0_0),.din(w_dff_A_kItvCpdm3_0),.clk(gclk));
	jdff dff_A_NuQSjE8t0_0(.dout(w_dff_A_VkvuCOeX2_0),.din(w_dff_A_NuQSjE8t0_0),.clk(gclk));
	jdff dff_A_VkvuCOeX2_0(.dout(w_dff_A_1OsQOe6J0_0),.din(w_dff_A_VkvuCOeX2_0),.clk(gclk));
	jdff dff_A_1OsQOe6J0_0(.dout(G367),.din(w_dff_A_1OsQOe6J0_0),.clk(gclk));
	jdff dff_A_gMbPIbhZ9_2(.dout(w_dff_A_pePACUYr0_0),.din(w_dff_A_gMbPIbhZ9_2),.clk(gclk));
	jdff dff_A_pePACUYr0_0(.dout(w_dff_A_J8CYK0z98_0),.din(w_dff_A_pePACUYr0_0),.clk(gclk));
	jdff dff_A_J8CYK0z98_0(.dout(w_dff_A_lh9HrNeF8_0),.din(w_dff_A_J8CYK0z98_0),.clk(gclk));
	jdff dff_A_lh9HrNeF8_0(.dout(w_dff_A_C6v6yx9W8_0),.din(w_dff_A_lh9HrNeF8_0),.clk(gclk));
	jdff dff_A_C6v6yx9W8_0(.dout(G387),.din(w_dff_A_C6v6yx9W8_0),.clk(gclk));
	jdff dff_A_6AG3SgwF9_1(.dout(w_dff_A_1wa6scRT4_0),.din(w_dff_A_6AG3SgwF9_1),.clk(gclk));
	jdff dff_A_1wa6scRT4_0(.dout(w_dff_A_EZIh7BOM0_0),.din(w_dff_A_1wa6scRT4_0),.clk(gclk));
	jdff dff_A_EZIh7BOM0_0(.dout(w_dff_A_QDHzbLAS4_0),.din(w_dff_A_EZIh7BOM0_0),.clk(gclk));
	jdff dff_A_QDHzbLAS4_0(.dout(w_dff_A_7B7YrEgs1_0),.din(w_dff_A_QDHzbLAS4_0),.clk(gclk));
	jdff dff_A_7B7YrEgs1_0(.dout(w_dff_A_lGrXPsPf5_0),.din(w_dff_A_7B7YrEgs1_0),.clk(gclk));
	jdff dff_A_lGrXPsPf5_0(.dout(w_dff_A_63rnxrt66_0),.din(w_dff_A_lGrXPsPf5_0),.clk(gclk));
	jdff dff_A_63rnxrt66_0(.dout(G393),.din(w_dff_A_63rnxrt66_0),.clk(gclk));
	jdff dff_A_zmyyTuog8_1(.dout(w_dff_A_h8B1FVzK0_0),.din(w_dff_A_zmyyTuog8_1),.clk(gclk));
	jdff dff_A_h8B1FVzK0_0(.dout(w_dff_A_OSUarnG38_0),.din(w_dff_A_h8B1FVzK0_0),.clk(gclk));
	jdff dff_A_OSUarnG38_0(.dout(w_dff_A_PDseqAHC6_0),.din(w_dff_A_OSUarnG38_0),.clk(gclk));
	jdff dff_A_PDseqAHC6_0(.dout(w_dff_A_Ev65jC9w8_0),.din(w_dff_A_PDseqAHC6_0),.clk(gclk));
	jdff dff_A_Ev65jC9w8_0(.dout(w_dff_A_aUQ6yJFl6_0),.din(w_dff_A_Ev65jC9w8_0),.clk(gclk));
	jdff dff_A_aUQ6yJFl6_0(.dout(G390),.din(w_dff_A_aUQ6yJFl6_0),.clk(gclk));
	jdff dff_A_ywGiTRig5_1(.dout(w_dff_A_hCj3951Q9_0),.din(w_dff_A_ywGiTRig5_1),.clk(gclk));
	jdff dff_A_hCj3951Q9_0(.dout(w_dff_A_Y34FfsEq6_0),.din(w_dff_A_hCj3951Q9_0),.clk(gclk));
	jdff dff_A_Y34FfsEq6_0(.dout(w_dff_A_KbweROGQ1_0),.din(w_dff_A_Y34FfsEq6_0),.clk(gclk));
	jdff dff_A_KbweROGQ1_0(.dout(w_dff_A_RAOIGzOa2_0),.din(w_dff_A_KbweROGQ1_0),.clk(gclk));
	jdff dff_A_RAOIGzOa2_0(.dout(G378),.din(w_dff_A_RAOIGzOa2_0),.clk(gclk));
	jdff dff_A_ULxsSlua0_1(.dout(w_dff_A_CB5hT0D90_0),.din(w_dff_A_ULxsSlua0_1),.clk(gclk));
	jdff dff_A_CB5hT0D90_0(.dout(w_dff_A_VKLgk1X27_0),.din(w_dff_A_CB5hT0D90_0),.clk(gclk));
	jdff dff_A_VKLgk1X27_0(.dout(G375),.din(w_dff_A_VKLgk1X27_0),.clk(gclk));
	jdff dff_A_BEk3hAnd8_1(.dout(w_dff_A_OYV2J0ds3_0),.din(w_dff_A_BEk3hAnd8_1),.clk(gclk));
	jdff dff_A_OYV2J0ds3_0(.dout(w_dff_A_Sp6VE8id9_0),.din(w_dff_A_OYV2J0ds3_0),.clk(gclk));
	jdff dff_A_Sp6VE8id9_0(.dout(w_dff_A_FoPg98jD2_0),.din(w_dff_A_Sp6VE8id9_0),.clk(gclk));
	jdff dff_A_FoPg98jD2_0(.dout(w_dff_A_UJV9lTxp4_0),.din(w_dff_A_FoPg98jD2_0),.clk(gclk));
	jdff dff_A_UJV9lTxp4_0(.dout(G381),.din(w_dff_A_UJV9lTxp4_0),.clk(gclk));
	jdff dff_A_jCISqWYT9_1(.dout(G407),.din(w_dff_A_jCISqWYT9_1),.clk(gclk));
	jdff dff_A_ysFzlHig4_2(.dout(G402),.din(w_dff_A_ysFzlHig4_2),.clk(gclk));
endmodule

