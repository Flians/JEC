/*
gf_c1908:
	jxor: 78
	jspl: 105
	jspl3: 86
	jnot: 30
	jdff: 969
	jor: 87
	jand: 120

Summary:
	jxor: 78
	jspl: 105
	jspl3: 86
	jnot: 30
	jdff: 969
	jor: 87
	jand: 120

The maximum logic level gap of any gate:
	gf_c1908: 17
*/

module gf_c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n173;
	wire n174;
	wire n175;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n201;
	wire n203;
	wire n204;
	wire n206;
	wire n207;
	wire n208;
	wire n210;
	wire n211;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n220;
	wire n222;
	wire n223;
	wire n224;
	wire n226;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n270;
	wire n271;
	wire n272;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n348;
	wire n349;
	wire n350;
	wire n352;
	wire n353;
	wire n354;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n369;
	wire n370;
	wire n371;
	wire [2:0] w_G101_0;
	wire [2:0] w_G104_0;
	wire [2:0] w_G107_0;
	wire [2:0] w_G110_0;
	wire [2:0] w_G113_0;
	wire [2:0] w_G116_0;
	wire [2:0] w_G119_0;
	wire [2:0] w_G122_0;
	wire [1:0] w_G122_1;
	wire [2:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [2:0] w_G131_0;
	wire [2:0] w_G134_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G140_0;
	wire [2:0] w_G143_0;
	wire [2:0] w_G146_0;
	wire [2:0] w_G210_0;
	wire [1:0] w_G214_0;
	wire [2:0] w_G217_0;
	wire [1:0] w_G221_0;
	wire [1:0] w_G224_0;
	wire [1:0] w_G227_0;
	wire [2:0] w_G234_0;
	wire [1:0] w_G234_1;
	wire [2:0] w_G237_0;
	wire [2:0] w_G469_0;
	wire [2:0] w_G472_0;
	wire [2:0] w_G475_0;
	wire [2:0] w_G478_0;
	wire [1:0] w_G898_0;
	wire [1:0] w_G900_0;
	wire [2:0] w_G902_0;
	wire [2:0] w_G902_1;
	wire [2:0] w_G902_2;
	wire [2:0] w_G902_3;
	wire [2:0] w_G952_0;
	wire [2:0] w_G953_0;
	wire [2:0] w_G953_1;
	wire [1:0] w_G953_2;
	wire [2:0] w_n58_0;
	wire [2:0] w_n58_1;
	wire [2:0] w_n58_2;
	wire [1:0] w_n63_0;
	wire [1:0] w_n66_0;
	wire [1:0] w_n67_0;
	wire [1:0] w_n70_0;
	wire [1:0] w_n71_0;
	wire [1:0] w_n73_0;
	wire [1:0] w_n74_0;
	wire [2:0] w_n76_0;
	wire [2:0] w_n76_1;
	wire [1:0] w_n77_0;
	wire [1:0] w_n78_0;
	wire [2:0] w_n81_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n86_0;
	wire [1:0] w_n90_0;
	wire [1:0] w_n91_0;
	wire [2:0] w_n92_0;
	wire [1:0] w_n92_1;
	wire [2:0] w_n93_0;
	wire [1:0] w_n93_1;
	wire [1:0] w_n94_0;
	wire [2:0] w_n95_0;
	wire [1:0] w_n95_1;
	wire [2:0] w_n96_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n102_0;
	wire [2:0] w_n103_0;
	wire [2:0] w_n103_1;
	wire [2:0] w_n103_2;
	wire [2:0] w_n103_3;
	wire [1:0] w_n107_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n109_0;
	wire [1:0] w_n110_0;
	wire [1:0] w_n111_0;
	wire [2:0] w_n112_0;
	wire [1:0] w_n112_1;
	wire [2:0] w_n113_0;
	wire [1:0] w_n118_0;
	wire [1:0] w_n119_0;
	wire [1:0] w_n120_0;
	wire [1:0] w_n121_0;
	wire [2:0] w_n122_0;
	wire [1:0] w_n122_1;
	wire [1:0] w_n124_0;
	wire [1:0] w_n126_0;
	wire [1:0] w_n127_0;
	wire [2:0] w_n130_0;
	wire [1:0] w_n130_1;
	wire [2:0] w_n131_0;
	wire [2:0] w_n131_1;
	wire [1:0] w_n139_0;
	wire [1:0] w_n140_0;
	wire [2:0] w_n141_0;
	wire [1:0] w_n141_1;
	wire [2:0] w_n151_0;
	wire [1:0] w_n152_0;
	wire [2:0] w_n153_0;
	wire [1:0] w_n153_1;
	wire [2:0] w_n154_0;
	wire [1:0] w_n154_1;
	wire [1:0] w_n155_0;
	wire [1:0] w_n156_0;
	wire [1:0] w_n157_0;
	wire [2:0] w_n160_0;
	wire [2:0] w_n160_1;
	wire [2:0] w_n161_0;
	wire [1:0] w_n161_1;
	wire [1:0] w_n162_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n163_1;
	wire [1:0] w_n164_0;
	wire [2:0] w_n165_0;
	wire [1:0] w_n166_0;
	wire [2:0] w_n168_0;
	wire [1:0] w_n168_1;
	wire [1:0] w_n169_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n171_0;
	wire [2:0] w_n173_0;
	wire [1:0] w_n173_1;
	wire [1:0] w_n174_0;
	wire [1:0] w_n175_0;
	wire [2:0] w_n177_0;
	wire [1:0] w_n178_0;
	wire [1:0] w_n180_0;
	wire [2:0] w_n182_0;
	wire [2:0] w_n182_1;
	wire [2:0] w_n183_0;
	wire [1:0] w_n184_0;
	wire [1:0] w_n186_0;
	wire [1:0] w_n189_0;
	wire [2:0] w_n191_0;
	wire [2:0] w_n192_0;
	wire [2:0] w_n195_0;
	wire [2:0] w_n197_0;
	wire [1:0] w_n197_1;
	wire [1:0] w_n198_0;
	wire [2:0] w_n199_0;
	wire [1:0] w_n201_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n206_0;
	wire [1:0] w_n208_0;
	wire [1:0] w_n210_0;
	wire [1:0] w_n211_0;
	wire [2:0] w_n214_0;
	wire [2:0] w_n216_0;
	wire [1:0] w_n216_1;
	wire [1:0] w_n217_0;
	wire [1:0] w_n218_0;
	wire [1:0] w_n220_0;
	wire [1:0] w_n224_0;
	wire [1:0] w_n226_0;
	wire [2:0] w_n242_0;
	wire [2:0] w_n242_1;
	wire [2:0] w_n242_2;
	wire [1:0] w_n243_0;
	wire [1:0] w_n249_0;
	wire [2:0] w_n258_0;
	wire [2:0] w_n265_0;
	wire [2:0] w_n265_1;
	wire [1:0] w_n265_2;
	wire [1:0] w_n274_0;
	wire [2:0] w_n278_0;
	wire [1:0] w_n279_0;
	wire [1:0] w_n280_0;
	wire [2:0] w_n282_0;
	wire [1:0] w_n282_1;
	wire [1:0] w_n286_0;
	wire [2:0] w_n287_0;
	wire [1:0] w_n287_1;
	wire [1:0] w_n288_0;
	wire [2:0] w_n291_0;
	wire [1:0] w_n291_1;
	wire [1:0] w_n292_0;
	wire [1:0] w_n293_0;
	wire [1:0] w_n294_0;
	wire [1:0] w_n297_0;
	wire [1:0] w_n303_0;
	wire [2:0] w_n307_0;
	wire [1:0] w_n313_0;
	wire [2:0] w_n316_0;
	wire [2:0] w_n317_0;
	wire [1:0] w_n322_0;
	wire [1:0] w_n323_0;
	wire [1:0] w_n327_0;
	wire [1:0] w_n329_0;
	wire [1:0] w_n341_0;
	wire w_dff_B_KUG64qFo9_0;
	wire w_dff_B_394Fxekk6_0;
	wire w_dff_B_alWpnuZ68_0;
	wire w_dff_B_flIMqsTO9_0;
	wire w_dff_B_X1XwYjW90_0;
	wire w_dff_B_oCKmzzRJ2_0;
	wire w_dff_B_HucuwSJG9_0;
	wire w_dff_B_eggdHZDG6_0;
	wire w_dff_A_IG0CL64y6_0;
	wire w_dff_A_v3ni466f3_0;
	wire w_dff_B_k5gOsM257_0;
	wire w_dff_B_JBz7l3hc8_0;
	wire w_dff_B_hT1JvqQo9_0;
	wire w_dff_B_QTJGx9Zi8_0;
	wire w_dff_B_E3zHyqyO6_0;
	wire w_dff_B_8UVV9BKq0_1;
	wire w_dff_B_Lvpku14t8_1;
	wire w_dff_B_dvRgyTWL3_1;
	wire w_dff_B_f3V5GFWe6_1;
	wire w_dff_B_w1ZBE5So9_1;
	wire w_dff_B_D6vUSOhQ9_1;
	wire w_dff_B_wo1dfjjy0_1;
	wire w_dff_B_HxB01BHw8_1;
	wire w_dff_B_LP0n0gDD2_1;
	wire w_dff_B_j5g1Z4K63_1;
	wire w_dff_B_nOi7yzSc6_1;
	wire w_dff_B_XY4RlwRU3_1;
	wire w_dff_B_oVS34vDx7_0;
	wire w_dff_B_s2iS1UZf1_0;
	wire w_dff_B_Km60sTcO5_0;
	wire w_dff_B_7cITet7p8_0;
	wire w_dff_B_aJLU51O03_0;
	wire w_dff_B_8yblqgjN8_0;
	wire w_dff_B_GPNNfbOx8_0;
	wire w_dff_B_h0NNqSV74_0;
	wire w_dff_B_FmKeF8Sd9_0;
	wire w_dff_B_A9yugYQe2_0;
	wire w_dff_B_CNdE24Io0_0;
	wire w_dff_B_9UvZ2llQ9_0;
	wire w_dff_B_f547bRLo4_0;
	wire w_dff_B_U4qzGoUC9_0;
	wire w_dff_A_XxGbtZY94_1;
	wire w_dff_A_I3PxFMEP5_1;
	wire w_dff_A_TGFYP5zS4_1;
	wire w_dff_A_2ZW7aQZH7_1;
	wire w_dff_A_pLuSHK438_1;
	wire w_dff_A_crK3MAGE6_1;
	wire w_dff_A_QKwrXAwl5_1;
	wire w_dff_A_kmB8DmzN6_1;
	wire w_dff_A_X7vahN7m6_1;
	wire w_dff_A_aohLhlQ79_1;
	wire w_dff_A_RYgo71xN7_1;
	wire w_dff_A_DGTpZgc44_1;
	wire w_dff_A_k12CDglC2_1;
	wire w_dff_A_l53IoIuA6_1;
	wire w_dff_A_gLLZy1pU5_1;
	wire w_dff_A_syXOUwlA2_1;
	wire w_dff_A_vuuSfQjb4_1;
	wire w_dff_A_z7TEBZSF4_1;
	wire w_dff_A_p3pKopkY3_1;
	wire w_dff_A_FGhfCPHc4_1;
	wire w_dff_A_dp7rQfin0_1;
	wire w_dff_A_pHGEWigZ7_1;
	wire w_dff_A_A9Mpn6Mo7_1;
	wire w_dff_A_vEDHGsRF1_1;
	wire w_dff_A_wke8CEi98_1;
	wire w_dff_A_Hi8O8vN88_1;
	wire w_dff_A_kt91S0nH0_1;
	wire w_dff_A_mFka8xG79_1;
	wire w_dff_A_GmsY3EdE6_1;
	wire w_dff_A_AXsYIj0G3_1;
	wire w_dff_A_QVseP5Xn5_1;
	wire w_dff_A_TYWhiCcb1_1;
	wire w_dff_A_iGmSLGYQ0_2;
	wire w_dff_A_JNDw6oqa7_2;
	wire w_dff_A_F7AUvBLO4_2;
	wire w_dff_A_v3Az2e4l6_2;
	wire w_dff_A_ShRa6vIr0_2;
	wire w_dff_A_7ucS4sL53_2;
	wire w_dff_A_YPE5SCWC0_2;
	wire w_dff_A_QzBMqiCV4_2;
	wire w_dff_A_zOufd4Aa8_2;
	wire w_dff_A_T2uI2d8G1_2;
	wire w_dff_A_ayxp7PCQ1_2;
	wire w_dff_A_2KVwM7VM7_2;
	wire w_dff_A_GnsqHrad7_2;
	wire w_dff_A_ToUJgmBh8_2;
	wire w_dff_A_5YD3cgRK2_2;
	wire w_dff_A_mDqaywDU7_2;
	wire w_dff_A_WXr3mAOY7_2;
	wire w_dff_A_fX4U4ovf9_0;
	wire w_dff_A_cMFoa89n8_1;
	wire w_dff_B_hGOzfkvM9_1;
	wire w_dff_B_YURzaCoG9_1;
	wire w_dff_B_5LsUcDqb1_1;
	wire w_dff_B_lWogwtJi2_1;
	wire w_dff_B_8Hz62FqG2_1;
	wire w_dff_B_vFUmr7hp3_1;
	wire w_dff_B_J5luUa8b5_1;
	wire w_dff_B_drqsJAl31_1;
	wire w_dff_B_aiC7ouoZ6_1;
	wire w_dff_B_WNGVCYfI7_1;
	wire w_dff_B_0XerGWij3_1;
	wire w_dff_B_8QhtpKir0_1;
	wire w_dff_B_UX1OY6Gb2_0;
	wire w_dff_B_QpE7LmeA5_0;
	wire w_dff_B_FbnBAdS51_0;
	wire w_dff_B_w35X5nWO4_0;
	wire w_dff_B_w41uq7435_0;
	wire w_dff_B_3mQRfDGC9_0;
	wire w_dff_B_86QDvtdV9_0;
	wire w_dff_B_HeISs4qd9_0;
	wire w_dff_B_YxJ0zRfD3_0;
	wire w_dff_B_vvhr6LsZ4_0;
	wire w_dff_B_240jvMa60_0;
	wire w_dff_B_HAqUgjKD2_0;
	wire w_dff_B_0o4YFTJ35_0;
	wire w_dff_B_uSiNie2K1_0;
	wire w_dff_B_xxqWYu090_1;
	wire w_dff_B_gJdEHobR1_1;
	wire w_dff_B_o1k8CBxA6_1;
	wire w_dff_B_BvqV64tH2_1;
	wire w_dff_B_i6qCSWfC6_2;
	wire w_dff_A_ABtNJUFx6_1;
	wire w_dff_B_K6u4Fd705_2;
	wire w_dff_A_DoAoh6qP1_2;
	wire w_dff_A_bGwVcjBD4_2;
	wire w_dff_B_OqorBsIl3_3;
	wire w_dff_B_sb9iZ8bG2_3;
	wire w_dff_B_VkBUUOFb5_0;
	wire w_dff_B_wIc1UPH12_0;
	wire w_dff_B_VQ2fVj6Q2_0;
	wire w_dff_B_z823ZQ8i2_0;
	wire w_dff_B_CKP56xHB2_0;
	wire w_dff_B_Xx7E4TlV7_0;
	wire w_dff_B_mHbSeaVo7_0;
	wire w_dff_B_PygfWZwp8_0;
	wire w_dff_B_eh4kMKeL8_0;
	wire w_dff_B_WZiz5vdx3_0;
	wire w_dff_B_G6Pc5LI60_0;
	wire w_dff_B_WGDz4yIs8_0;
	wire w_dff_B_lXOg0ONp7_0;
	wire w_dff_B_vBaRG9Ml8_0;
	wire w_dff_B_C5LRueNP1_0;
	wire w_dff_B_d6aTAMLa3_0;
	wire w_dff_B_Jho5Yf9L0_0;
	wire w_dff_B_jrfgMv3B0_0;
	wire w_dff_B_M7QJVnjF3_0;
	wire w_dff_B_rWpQweSu9_0;
	wire w_dff_B_9a3Fue1j0_0;
	wire w_dff_B_Mklt5Ah61_0;
	wire w_dff_B_PuUswaoM0_0;
	wire w_dff_B_bHWz2Acr8_0;
	wire w_dff_B_WPzS1h6Y7_0;
	wire w_dff_B_ai9z8Ib93_0;
	wire w_dff_B_l8DfnSgd7_1;
	wire w_dff_B_slj6ZFIj6_1;
	wire w_dff_B_JQNBt3Tw0_1;
	wire w_dff_A_AlG92Tz52_1;
	wire w_dff_A_WANtlcxU1_2;
	wire w_dff_A_nJmoAc6P5_1;
	wire w_dff_A_Mfurm3pw8_1;
	wire w_dff_A_1yr2Fkib6_1;
	wire w_dff_A_FPGOcCb08_2;
	wire w_dff_A_82Ol37eH4_1;
	wire w_dff_A_3sTCNM3y5_0;
	wire w_dff_A_aVPtgSo02_2;
	wire w_dff_A_Hp3hdCfF5_0;
	wire w_dff_A_lGq66MbF9_1;
	wire w_dff_B_hFGawRW00_2;
	wire w_dff_A_33pc2Raq6_0;
	wire w_dff_A_wTKLKhEd4_2;
	wire w_dff_A_gmOYxxun3_0;
	wire w_dff_A_WSLk10X92_2;
	wire w_dff_B_YpyyUZvx8_3;
	wire w_dff_B_6OB8wPMk2_3;
	wire w_dff_A_cCQcj4iH3_1;
	wire w_dff_A_2sTvlTIs9_2;
	wire w_dff_B_9j5Z6XY35_0;
	wire w_dff_B_To039hLW4_0;
	wire w_dff_B_qS0RVbv06_0;
	wire w_dff_B_QMmS2fVF6_0;
	wire w_dff_B_XWojwD808_0;
	wire w_dff_B_wRxdAre98_0;
	wire w_dff_B_1bIDSDbp4_0;
	wire w_dff_B_z32MSyet2_0;
	wire w_dff_B_toAuobQO5_0;
	wire w_dff_B_nTDLVa0Y5_0;
	wire w_dff_B_C2Wt8arC7_0;
	wire w_dff_B_jPLi9S8P9_0;
	wire w_dff_B_jzpWERoA1_0;
	wire w_dff_B_o3xNFRU61_0;
	wire w_dff_B_GVXrhrtJ9_0;
	wire w_dff_A_cxbLVBeD5_1;
	wire w_dff_A_HVcZbEPt6_1;
	wire w_dff_A_uD3aOx0V1_1;
	wire w_dff_A_mOpspPGk4_1;
	wire w_dff_A_WqcpWQGw2_1;
	wire w_dff_A_10g0eqLL5_1;
	wire w_dff_A_mNwDuFKi5_1;
	wire w_dff_A_6qXO61xc4_1;
	wire w_dff_A_fpPIGJVJ4_1;
	wire w_dff_A_ntxM5n5S8_1;
	wire w_dff_A_6kRSMX3n4_1;
	wire w_dff_A_GShpcJh22_1;
	wire w_dff_A_NJQ70hQm1_1;
	wire w_dff_A_OgvA04eG7_1;
	wire w_dff_A_pQFwUsRx7_1;
	wire w_dff_A_9JcezBKN5_1;
	wire w_dff_A_eveR7xjG5_1;
	wire w_dff_A_R0P7A7Oe4_2;
	wire w_dff_A_doPstua32_2;
	wire w_dff_A_IaklNWCl1_2;
	wire w_dff_A_vl8SOYU20_2;
	wire w_dff_A_OOXBT9eP7_2;
	wire w_dff_A_LSOiE9oF1_2;
	wire w_dff_A_0UcrAbvE0_2;
	wire w_dff_A_ULUrvKIz6_2;
	wire w_dff_A_XUxngNkg4_2;
	wire w_dff_A_Sj6X3e9V5_2;
	wire w_dff_A_Xg6o16VL7_2;
	wire w_dff_A_YDDeoh0r5_2;
	wire w_dff_A_VtmdS7t47_2;
	wire w_dff_A_fIZEEFDX0_2;
	wire w_dff_A_SkIp3MHM6_2;
	wire w_dff_A_C32Ed3NP0_2;
	wire w_dff_A_9vXg7p2U9_2;
	wire w_dff_B_RqHLDa1b8_1;
	wire w_dff_B_JC95DaZ65_1;
	wire w_dff_A_1VRB2xs14_0;
	wire w_dff_A_szBFXo8J3_1;
	wire w_dff_A_BsJ2jOKO4_2;
	wire w_dff_A_qvlnoTIO5_0;
	wire w_dff_A_zlZRoQlY1_2;
	wire w_dff_B_PzhPMEus9_0;
	wire w_dff_B_dkcwcKti5_0;
	wire w_dff_B_2muhCsUb1_0;
	wire w_dff_A_ZJtyRA0T1_1;
	wire w_dff_A_CRco7veP1_0;
	wire w_dff_A_dKrVgv1U3_2;
	wire w_dff_A_jElLZGmm8_1;
	wire w_dff_A_3CCsnjzW2_0;
	wire w_dff_A_19G8xX9t3_0;
	wire w_dff_A_EwZWUKIS7_0;
	wire w_dff_A_pmbcomq20_2;
	wire w_dff_A_9S237OTl6_2;
	wire w_dff_A_8pmT6EMg5_2;
	wire w_dff_A_eHRBrCIQ1_2;
	wire w_dff_A_Xv4Re0VA8_0;
	wire w_dff_A_Cpn0gaCa7_1;
	wire w_dff_A_gPnpAazZ3_1;
	wire w_dff_A_ZwXfHhEL8_2;
	wire w_dff_A_WjCKIAiK5_0;
	wire w_dff_A_DTPDCWCH0_1;
	wire w_dff_B_vDF4uLgW4_2;
	wire w_dff_A_yPVhSkGV2_1;
	wire w_dff_A_oqBjpYYL8_1;
	wire w_dff_A_2ypsFFp70_0;
	wire w_dff_B_L2sw5HXi6_2;
	wire w_dff_A_REp22pjD7_2;
	wire w_dff_A_zT089Ygc2_2;
	wire w_dff_A_3b8lsqOb6_2;
	wire w_dff_A_SWInxcw56_2;
	wire w_dff_B_MRaEe7G13_1;
	wire w_dff_B_2bzhOtmf4_1;
	wire w_dff_B_OZ6XhuiB2_1;
	wire w_dff_B_S3yyGRCa6_1;
	wire w_dff_B_4GcJj6UK9_1;
	wire w_dff_A_jeviynMh1_1;
	wire w_dff_A_Goheoi8v6_1;
	wire w_dff_A_UUI63NDL8_1;
	wire w_dff_A_Zo59uV6y7_2;
	wire w_dff_A_dgHihsKT6_0;
	wire w_dff_A_AE1D2ZU45_1;
	wire w_dff_A_znOEPE3t7_2;
	wire w_dff_B_5nsrbSC05_1;
	wire w_dff_B_OPIO8SGq4_1;
	wire w_dff_B_UnXNkBs69_1;
	wire w_dff_B_pkG8ZWhz3_1;
	wire w_dff_B_kbcpQt2j9_1;
	wire w_dff_A_NAtrOi5y4_1;
	wire w_dff_A_6Mu5TVS08_0;
	wire w_dff_A_ESbhtxXb4_1;
	wire w_dff_B_k6APoGJQ8_1;
	wire w_dff_B_DS7aIEQu2_1;
	wire w_dff_B_h9cOKgaC6_1;
	wire w_dff_B_xn4tmahP4_1;
	wire w_dff_B_NsDCSFXi4_1;
	wire w_dff_A_zDABCEQv4_0;
	wire w_dff_A_IwDaN4mS1_0;
	wire w_dff_A_Ep1bIAFe4_0;
	wire w_dff_A_nmWGtdch3_0;
	wire w_dff_A_B7fuyqWW3_0;
	wire w_dff_A_nUzh37dZ2_0;
	wire w_dff_A_EJl3uVnT3_0;
	wire w_dff_A_DyOqZUPQ7_0;
	wire w_dff_A_4kAObYLq2_0;
	wire w_dff_A_1ggNEJ7t1_0;
	wire w_dff_A_U73lyVPM5_0;
	wire w_dff_A_tQh4oj1H7_0;
	wire w_dff_A_tqndhuCu4_0;
	wire w_dff_A_EQkrYTW60_1;
	wire w_dff_A_Nep6uVWh4_0;
	wire w_dff_A_i7U0X4g38_0;
	wire w_dff_A_N29Ib9Xp6_0;
	wire w_dff_A_iatluKOH0_0;
	wire w_dff_A_nxfbMlCP2_0;
	wire w_dff_A_oDForQPh5_0;
	wire w_dff_A_Z6J848JK0_0;
	wire w_dff_A_fpR1vrs22_0;
	wire w_dff_A_jIcyLV9S1_0;
	wire w_dff_A_BDCUAhlO5_0;
	wire w_dff_A_IP1JPemf0_0;
	wire w_dff_A_kDqQp4wh2_0;
	wire w_dff_A_zoEEl4xc9_0;
	wire w_dff_A_MMQqbunt0_0;
	wire w_dff_A_NUweUMAO7_0;
	wire w_dff_A_HvlivWmk0_0;
	wire w_dff_A_r5oBXoY02_2;
	wire w_dff_A_Fe6t2XlX6_2;
	wire w_dff_A_wWIJ0g4Y4_2;
	wire w_dff_A_YmUIaqRu3_2;
	wire w_dff_A_hDwbYA1M4_2;
	wire w_dff_A_ULtBYnlK8_2;
	wire w_dff_A_sjWVkpVN1_1;
	wire w_dff_A_kHyHxSiA5_1;
	wire w_dff_A_HtiQBFxH9_2;
	wire w_dff_A_wQPGfbPQ3_2;
	wire w_dff_A_OU8Ehhts9_1;
	wire w_dff_A_aYi1miGV4_1;
	wire w_dff_A_vI1tui6I2_1;
	wire w_dff_A_tjuDygRx7_2;
	wire w_dff_A_Pe5pLhwT1_2;
	wire w_dff_A_zSeAZakS0_2;
	wire w_dff_A_FLf3qhb67_1;
	wire w_dff_A_XnCSF2Rn3_1;
	wire w_dff_A_9E2EhCul1_1;
	wire w_dff_A_BPSgy5466_1;
	wire w_dff_A_LYnqv5er8_0;
	wire w_dff_A_D7vO2Dl39_0;
	wire w_dff_A_v0qq9xQJ7_0;
	wire w_dff_A_oyVB0b665_0;
	wire w_dff_A_8XfYXIVT6_0;
	wire w_dff_A_FmUb1ebN6_0;
	wire w_dff_A_bOi4UE0B1_0;
	wire w_dff_A_Wj38kN3O5_0;
	wire w_dff_A_kCc9f4Ez3_0;
	wire w_dff_A_ym2UMXSd0_0;
	wire w_dff_A_PkLqv2Px5_0;
	wire w_dff_A_iQSMFodB5_0;
	wire w_dff_A_ASSNhaad5_0;
	wire w_dff_B_aFnTQLtg1_1;
	wire w_dff_A_x4CoadrC8_1;
	wire w_dff_B_mpwLwhvW6_0;
	wire w_dff_B_JxaDq2Ff9_0;
	wire w_dff_A_9dENtCRg6_0;
	wire w_dff_A_TXUsMIO52_1;
	wire w_dff_A_4iQ5PsFD0_1;
	wire w_dff_A_SOb0HfFp1_2;
	wire w_dff_A_DyND0V2T2_2;
	wire w_dff_B_iZSNUWk79_3;
	wire w_dff_B_sq9N4pXi0_3;
	wire w_dff_A_JQVYE69n0_0;
	wire w_dff_A_hZVR3lWF6_0;
	wire w_dff_A_PIaYCAmj5_1;
	wire w_dff_A_wcBhESmt3_1;
	wire w_dff_A_m9EiKjWD6_1;
	wire w_dff_A_geY3g1Pp7_1;
	wire w_dff_A_4hau76MP3_1;
	wire w_dff_A_ZJ1LG8BS8_2;
	wire w_dff_A_Mskq4TCj1_2;
	wire w_dff_A_laEriNyn6_2;
	wire w_dff_A_GrrdG6wv4_2;
	wire w_dff_A_woUgFLQV7_2;
	wire w_dff_A_bZqGKQsJ5_1;
	wire w_dff_A_tUN8qgig9_2;
	wire w_dff_B_SmSmmBJM7_3;
	wire w_dff_B_AYMGgiWa9_1;
	wire w_dff_B_6H4SbxbY6_1;
	wire w_dff_B_yHm5oCLr0_1;
	wire w_dff_B_ZOuoeaeS6_1;
	wire w_dff_B_P7OwcfVU5_1;
	wire w_dff_A_kl9t13r57_0;
	wire w_dff_A_TNj0WbIB7_0;
	wire w_dff_A_U89xG9Vd2_0;
	wire w_dff_A_fuuvUbSH8_0;
	wire w_dff_A_slbVTk6q2_0;
	wire w_dff_A_G9t4kHd51_0;
	wire w_dff_A_2X9bSZv90_0;
	wire w_dff_A_NWg9P04g9_0;
	wire w_dff_A_clhh5mhz1_0;
	wire w_dff_A_qKPCwKQn3_0;
	wire w_dff_A_ruJATUgD2_0;
	wire w_dff_A_tU0QD92Y8_0;
	wire w_dff_A_hB3DFJRv7_0;
	wire w_dff_A_4xVr9j2f6_0;
	wire w_dff_A_mjXoH1J22_0;
	wire w_dff_A_k6Pbvkn38_0;
	wire w_dff_A_SGzMnbvN2_0;
	wire w_dff_A_jwQz4vQy2_0;
	wire w_dff_A_AXm7U6Us4_0;
	wire w_dff_A_zAgb3OdD2_0;
	wire w_dff_A_2V1e7Wgg3_0;
	wire w_dff_A_vYQArisC2_0;
	wire w_dff_A_4blA1VWQ2_0;
	wire w_dff_A_mgyOkLTl1_0;
	wire w_dff_A_JB0utwUz8_0;
	wire w_dff_A_QrAafOiN1_0;
	wire w_dff_A_e7Eaff0f4_0;
	wire w_dff_A_VyrqZWlM8_0;
	wire w_dff_A_2wciar0F4_1;
	wire w_dff_A_eFk3xNBu3_0;
	wire w_dff_A_pXDpby4W7_0;
	wire w_dff_A_W2ztJ7SQ4_0;
	wire w_dff_A_hvYfNHjT3_0;
	wire w_dff_A_5V4Ph5x29_0;
	wire w_dff_A_hH17uga58_0;
	wire w_dff_A_NwXol6hV0_0;
	wire w_dff_A_M5IvXN4M6_0;
	wire w_dff_A_DiOHebvu5_0;
	wire w_dff_A_nHufrf4W8_0;
	wire w_dff_A_tkN9220D2_0;
	wire w_dff_A_5yz7tMgP9_2;
	wire w_dff_A_of9VE2Fz6_2;
	wire w_dff_A_ok4oxW2C4_1;
	wire w_dff_A_jm8LVCm13_1;
	wire w_dff_A_wdagkMWX9_2;
	wire w_dff_A_HL6lsrHG2_2;
	wire w_dff_A_jovm5fYq5_2;
	wire w_dff_A_Ty6DqOdE5_2;
	wire w_dff_A_ux5drhZs3_2;
	wire w_dff_A_7PyvplTS7_2;
	wire w_dff_A_6gxqJhLc9_2;
	wire w_dff_B_4qFwiVGm8_0;
	wire w_dff_A_atZXIHD73_0;
	wire w_dff_A_qpoPMpyG5_0;
	wire w_dff_A_I9CkvksI5_0;
	wire w_dff_A_QHyjIXl35_0;
	wire w_dff_A_3YG4nnEL4_0;
	wire w_dff_A_ene5vLYs2_0;
	wire w_dff_A_GzlSrgQs0_0;
	wire w_dff_A_jnLxujRO1_0;
	wire w_dff_A_0LJTcGe11_0;
	wire w_dff_A_MqlHttQF1_0;
	wire w_dff_A_n7J2kp7O1_0;
	wire w_dff_A_KailyL7u5_0;
	wire w_dff_A_QRFDXzvI1_0;
	wire w_dff_A_iDaGQMjD6_0;
	wire w_dff_A_12fiUFWN7_0;
	wire w_dff_B_r8oAmEr11_0;
	wire w_dff_B_LJSWXHrT7_0;
	wire w_dff_A_Yx99ZoGm0_0;
	wire w_dff_A_1E1OJPCW5_0;
	wire w_dff_A_j7AwUOtD4_0;
	wire w_dff_A_6A9Lev4r5_0;
	wire w_dff_A_v3PehkQg4_0;
	wire w_dff_A_Y5XU4Hfp1_0;
	wire w_dff_A_LTvMCBkk0_0;
	wire w_dff_A_IfLVXqSD8_0;
	wire w_dff_A_qJTHVnl13_0;
	wire w_dff_A_iF4bgQ0X4_0;
	wire w_dff_A_NV5cEZc60_0;
	wire w_dff_B_XiehfK7Z2_0;
	wire w_dff_A_pYCeHdjc8_0;
	wire w_dff_A_iU8Vv90l2_0;
	wire w_dff_A_DDLbsdKx4_0;
	wire w_dff_A_MIOm2Y5d6_0;
	wire w_dff_A_QOpjK0sa1_0;
	wire w_dff_A_SNhItwJm2_0;
	wire w_dff_A_m6rWxWNt5_0;
	wire w_dff_A_kG3Sw8WA6_0;
	wire w_dff_A_tUnhX7UW6_0;
	wire w_dff_A_SFbsM8nx7_0;
	wire w_dff_A_zQr574PS7_0;
	wire w_dff_A_pnVt8Qtv5_2;
	wire w_dff_A_d8mwiH3Y7_0;
	wire w_dff_A_NVAp0T9d8_0;
	wire w_dff_A_KvebgTYX9_0;
	wire w_dff_A_lkrQ8U7C8_0;
	wire w_dff_A_zWtAHudD5_0;
	wire w_dff_A_kl2sIsMx1_0;
	wire w_dff_A_p0tcYRmA8_0;
	wire w_dff_A_frApIrAX3_0;
	wire w_dff_A_YPTbDuYP4_0;
	wire w_dff_A_zwFgS79g3_0;
	wire w_dff_A_VJyD25BW2_0;
	wire w_dff_B_LDZoSPUp5_1;
	wire w_dff_A_rh5X5q869_0;
	wire w_dff_A_uC1SOD1I5_0;
	wire w_dff_A_8kbSZhd42_0;
	wire w_dff_A_UmkrL2Bk1_0;
	wire w_dff_A_XPV2EKVR7_0;
	wire w_dff_A_5HXS80rJ5_0;
	wire w_dff_A_9srne13f0_0;
	wire w_dff_A_IfPdIVTn7_0;
	wire w_dff_A_oFeZ3aKP2_2;
	wire w_dff_A_51Ifwn6Q6_2;
	wire w_dff_A_sdkKZKsZ1_2;
	wire w_dff_A_H9Rx8CDR8_2;
	wire w_dff_A_ksj7tYHN6_0;
	wire w_dff_A_Itc80Ea72_0;
	wire w_dff_A_M39xwuIo0_0;
	wire w_dff_A_vjxMacjW1_2;
	wire w_dff_A_6kFU2oJx0_2;
	wire w_dff_A_I3fxLiWP0_2;
	wire w_dff_A_UuNkoUaZ8_2;
	wire w_dff_A_kdAG6Xfd1_2;
	wire w_dff_A_eGqH9LWf9_1;
	wire w_dff_A_JxLCtbbS1_1;
	wire w_dff_A_lQnAgIGT8_1;
	wire w_dff_A_IHjKN1eP7_1;
	wire w_dff_A_TULZPGgB3_2;
	wire w_dff_A_PXokvH883_2;
	wire w_dff_A_6O1qeEnr7_2;
	wire w_dff_A_ranaXLiv7_2;
	wire w_dff_A_B7FQSY6u3_2;
	wire w_dff_A_lCVW8TrR0_2;
	wire w_dff_A_5UsLVNNZ0_2;
	wire w_dff_A_mf0Nb3ry8_2;
	wire w_dff_A_oEm0Nfpx8_2;
	wire w_dff_A_raUcn9Zs3_0;
	wire w_dff_A_HRi1yhR67_1;
	wire w_dff_A_SipQVlaa6_0;
	wire w_dff_A_lZsDVJ0U6_0;
	wire w_dff_A_zbzxFhuo2_0;
	wire w_dff_A_uI0Twndm0_1;
	wire w_dff_A_ZMcwRGWY9_1;
	wire w_dff_A_0Q9UZn8v8_1;
	wire w_dff_A_tod14Z6Y6_1;
	wire w_dff_A_n8swF2ru4_1;
	wire w_dff_A_zUrRyy1A7_1;
	wire w_dff_A_EAxCJBL25_1;
	wire w_dff_A_QKGNkm4x4_1;
	wire w_dff_A_ZwthStk77_1;
	wire w_dff_A_w9kyeGvU5_1;
	wire w_dff_A_pqYUnlPZ3_1;
	wire w_dff_A_oAl19vRy1_1;
	wire w_dff_B_MznmxNAg2_1;
	wire w_dff_B_Ny6Ilyp92_1;
	wire w_dff_A_IU5JvZM81_0;
	wire w_dff_A_fUlEsfb87_0;
	wire w_dff_A_QoXljbPT5_0;
	wire w_dff_A_DZezbzRa5_0;
	wire w_dff_A_wGEc2Yr71_0;
	wire w_dff_A_QOh7BTgc6_0;
	wire w_dff_A_ooAehbF87_0;
	wire w_dff_A_D6q22Tbe9_0;
	wire w_dff_A_I8DYA9Qv1_0;
	wire w_dff_A_evfcDjfb0_0;
	wire w_dff_A_ttSlfJ5X7_0;
	wire w_dff_A_CzsLeHrX3_2;
	wire w_dff_A_4wyfpWne7_1;
	wire w_dff_A_1s77Wb1L3_1;
	wire w_dff_A_Hri4DIpK9_0;
	wire w_dff_A_i447xYnj1_0;
	wire w_dff_A_keIiaf2X8_0;
	wire w_dff_A_rdWeC6J85_0;
	wire w_dff_A_BDE4x2dQ5_0;
	wire w_dff_A_h0zXj6WS3_0;
	wire w_dff_A_voyEWAbT6_0;
	wire w_dff_A_THTWZ5bi7_0;
	wire w_dff_A_To3tX07H9_0;
	wire w_dff_A_e4q1WrRp3_0;
	wire w_dff_A_LpAuHaD96_0;
	wire w_dff_A_FVrwDWEu1_0;
	wire w_dff_A_tg2iyD9N2_0;
	wire w_dff_A_muDEwOhg9_0;
	wire w_dff_A_ZPd97mhW6_1;
	wire w_dff_A_cXjJ8Opy8_0;
	wire w_dff_A_7ke4v4vb5_0;
	wire w_dff_A_rD8LgLhk2_0;
	wire w_dff_A_z2yKjB7S3_0;
	wire w_dff_A_bx9JhTvo5_0;
	wire w_dff_A_tMyZlCyb5_0;
	wire w_dff_A_szBWCZSm2_0;
	wire w_dff_A_2S0qgKkv2_0;
	wire w_dff_A_zZLvdgRX9_0;
	wire w_dff_A_LcBNfvQP6_0;
	wire w_dff_A_tFgBrtCK8_0;
	wire w_dff_A_0z7d7R0o8_1;
	wire w_dff_A_5e6SVyaf6_1;
	wire w_dff_A_oSJkky0K2_0;
	wire w_dff_A_MigrqXIy2_0;
	wire w_dff_A_51TVHLii9_0;
	wire w_dff_A_qTNc97ON5_0;
	wire w_dff_A_TSwgDWBk9_0;
	wire w_dff_A_UmJmSd2S3_0;
	wire w_dff_A_ZFmGawyg9_0;
	wire w_dff_A_5VP60dUO9_0;
	wire w_dff_A_sNAq7mdA3_0;
	wire w_dff_A_DX3jurAJ6_0;
	wire w_dff_B_QYOxYyQh7_3;
	wire w_dff_A_q10kKYis6_0;
	wire w_dff_A_xIbWc7Ky0_0;
	wire w_dff_A_gWk1F5el2_0;
	wire w_dff_A_mk8zZIpv4_0;
	wire w_dff_A_bpPjve709_0;
	wire w_dff_A_HFEBdRvo1_0;
	wire w_dff_A_T3f7AEBb4_0;
	wire w_dff_A_x38dOZzJ8_0;
	wire w_dff_A_QAexxTV21_0;
	wire w_dff_A_AYKDvV884_0;
	wire w_dff_A_NWJHmVeC7_0;
	wire w_dff_A_O6x76RM51_0;
	wire w_dff_A_b90dULUd8_0;
	wire w_dff_A_w4W009VD0_0;
	wire w_dff_A_UzgZewKc1_0;
	wire w_dff_A_BTydVxyW5_0;
	wire w_dff_A_8JAonBZg2_0;
	wire w_dff_A_ttCS3nBG4_0;
	wire w_dff_A_1mz5hszx0_0;
	wire w_dff_A_2FjiCEY75_0;
	wire w_dff_A_f6iP0Ym57_0;
	wire w_dff_A_FBAHzrOq1_0;
	wire w_dff_A_eUbbvWIE2_1;
	wire w_dff_A_gxkjBzf02_1;
	wire w_dff_A_ZliZVfE29_1;
	wire w_dff_A_RMrCSklw6_1;
	wire w_dff_A_RjTJWRhP6_1;
	wire w_dff_A_wrzlxhLN1_1;
	wire w_dff_A_kUu1Mzls8_1;
	wire w_dff_A_xUoOSNcT2_0;
	wire w_dff_A_mcS7BPxg3_0;
	wire w_dff_A_YwwUhA365_0;
	wire w_dff_A_Qja3vFFE1_0;
	wire w_dff_A_hgcMTnVZ5_0;
	wire w_dff_A_oF4bRuhQ9_0;
	wire w_dff_A_9PowGjIE1_0;
	wire w_dff_A_VvIYXqj79_0;
	wire w_dff_A_2vxRWCz35_0;
	wire w_dff_A_1xla2iDB4_0;
	wire w_dff_A_5YYL5PxY7_0;
	wire w_dff_A_6MTAriep6_0;
	wire w_dff_A_POImPkBN8_0;
	wire w_dff_B_rSeBfPmu5_1;
	wire w_dff_B_CN858ycW5_1;
	wire w_dff_B_bm62cSlV3_0;
	wire w_dff_A_IJjrdxt81_1;
	wire w_dff_A_Y3wHbrTA3_1;
	wire w_dff_A_MQYJhE4y9_1;
	wire w_dff_A_EQX7NdHE4_1;
	wire w_dff_A_VBLw9gIW4_1;
	wire w_dff_A_uHo0OgwD3_1;
	wire w_dff_A_8E6CQeG16_1;
	wire w_dff_A_6Z6ifrbO5_1;
	wire w_dff_A_dSleeQiT2_1;
	wire w_dff_A_MFjApbeP1_1;
	wire w_dff_A_i3wbb3jA9_1;
	wire w_dff_A_68C1tYLB7_1;
	wire w_dff_A_nga2Iew62_0;
	wire w_dff_A_Prbkge5E7_0;
	wire w_dff_A_nyqnGPiK0_0;
	wire w_dff_A_g30tdJAs5_0;
	wire w_dff_A_57r37bCg9_0;
	wire w_dff_A_RnaV8Cpi8_0;
	wire w_dff_A_3wMrxpah6_0;
	wire w_dff_A_TiER8Ba95_0;
	wire w_dff_A_0bVYrvQ19_0;
	wire w_dff_A_N5DlPHLb0_0;
	wire w_dff_A_NLyaARlw7_0;
	wire w_dff_A_49YsQQxQ0_0;
	wire w_dff_A_8p83rKFq1_0;
	wire w_dff_A_iUkqLGaB4_0;
	wire w_dff_A_yRgsuM321_0;
	wire w_dff_A_vVB9dRLj0_0;
	wire w_dff_A_2zdQqUdi1_0;
	wire w_dff_A_qtxv1z6j6_0;
	wire w_dff_A_9oU8Yl8g4_0;
	wire w_dff_A_rh4Mc7Np3_0;
	wire w_dff_A_yuS9hSMZ4_0;
	wire w_dff_A_CesXBU2u2_0;
	wire w_dff_A_6FeGUKFN4_1;
	wire w_dff_A_bly7LfRR9_2;
	wire w_dff_A_kfr5z0gz9_2;
	wire w_dff_A_XAwPxIpV3_1;
	wire w_dff_A_AaRWqBMq8_0;
	wire w_dff_A_9P4CbAt02_0;
	wire w_dff_A_dcESeOtO4_0;
	wire w_dff_A_pDr1Ffty0_0;
	wire w_dff_A_1XeUmfh58_0;
	wire w_dff_A_UN32hoSG4_0;
	wire w_dff_A_hSTybxa97_0;
	wire w_dff_A_gY1PkqQ66_0;
	wire w_dff_A_zKFyXN3O9_0;
	wire w_dff_A_P0HFjRp93_0;
	wire w_dff_A_oTlpMXOD9_0;
	wire w_dff_A_AjRwY4x19_0;
	wire w_dff_A_sI67HIFr7_0;
	wire w_dff_A_mYZjQoQo4_0;
	wire w_dff_A_JcBqaPAX3_2;
	wire w_dff_B_oh5QZlDJ4_3;
	wire w_dff_B_M3j6QPic7_3;
	wire w_dff_A_DcTb4TUm5_0;
	wire w_dff_A_fSoIHhZ60_0;
	wire w_dff_A_UFQDDTAz1_0;
	wire w_dff_A_tqndewNR1_0;
	wire w_dff_A_msk2iWml3_0;
	wire w_dff_A_g6NQHAoh9_0;
	wire w_dff_A_Q03tJHuo7_0;
	wire w_dff_A_zS251Rh04_0;
	wire w_dff_A_eAuW7okS4_0;
	wire w_dff_A_PAAYFXB99_0;
	wire w_dff_A_ryEwEkan5_0;
	wire w_dff_A_dmHWo8dH3_1;
	wire w_dff_A_1Zt6HHmR4_0;
	wire w_dff_A_2OvaMXge7_0;
	wire w_dff_A_hHsEpiOP6_0;
	wire w_dff_A_naPrRy4H7_0;
	wire w_dff_A_6RwbPwZM9_0;
	wire w_dff_A_fnWTvjgw0_0;
	wire w_dff_A_oszF1gkS2_0;
	wire w_dff_A_lEWY4w7D6_0;
	wire w_dff_A_bpc1Pi4f8_0;
	wire w_dff_A_4U4Dn5B10_0;
	wire w_dff_A_7dghcLrw1_0;
	wire w_dff_A_4MXdOiW35_0;
	wire w_dff_A_699554VJ5_0;
	wire w_dff_A_WciAu2Qa8_0;
	wire w_dff_A_N7BOy3hJ9_0;
	wire w_dff_A_3mtpfrEd9_0;
	wire w_dff_A_INH41D6U6_0;
	wire w_dff_A_PzPKDana9_0;
	wire w_dff_A_ZO63gEjH1_0;
	wire w_dff_A_rnKEsWx37_0;
	wire w_dff_A_NDNan9j49_0;
	wire w_dff_A_7gLeVlQI2_0;
	wire w_dff_A_XcRayItl7_1;
	wire w_dff_A_i9Og0RTD8_0;
	wire w_dff_A_yEqPEles3_0;
	wire w_dff_A_cVYZLGLT9_0;
	wire w_dff_A_lPlN46Zi2_0;
	wire w_dff_A_rA1iVUIV8_2;
	wire w_dff_A_lqjD7w6a1_2;
	wire w_dff_A_6vZRGKSU4_2;
	wire w_dff_A_z0LuLn477_2;
	wire w_dff_A_1yJTqHgw8_0;
	wire w_dff_A_ekZdutAZ2_0;
	wire w_dff_A_v6I2KH7f2_0;
	wire w_dff_A_JzvUZGg29_0;
	wire w_dff_A_azIfX3Y38_0;
	wire w_dff_A_DmcJJByz4_0;
	wire w_dff_A_DQ4NMHGq0_0;
	wire w_dff_A_g7pf2V5u6_0;
	wire w_dff_A_po0E5KME4_0;
	wire w_dff_A_sSABVEBM1_0;
	wire w_dff_A_wSa2KBbh5_0;
	wire w_dff_A_UwQepUMf0_0;
	wire w_dff_A_zjJnu9ml6_0;
	wire w_dff_A_53XppaRC8_0;
	wire w_dff_A_N1vGFIui8_0;
	wire w_dff_A_A3mIpxqX5_0;
	wire w_dff_A_Pb6hprQj1_0;
	wire w_dff_A_H4EUOxXu5_0;
	wire w_dff_A_z11SiYkI1_1;
	wire w_dff_A_u17sdarp3_1;
	wire w_dff_A_uejkKqTt8_1;
	wire w_dff_A_ErbHBAEZ7_1;
	wire w_dff_A_EBDUmzyk5_1;
	wire w_dff_A_bF80AltB1_1;
	wire w_dff_A_apHLc5GV3_1;
	wire w_dff_B_FkmzQT5x0_3;
	wire w_dff_B_sdL8uqzI8_3;
	wire w_dff_B_glo3kX217_3;
	wire w_dff_B_jqo5RMfB2_3;
	wire w_dff_B_3i79ASGC1_3;
	wire w_dff_B_orduQgoF1_3;
	wire w_dff_B_mKTavY603_3;
	wire w_dff_B_YiyA7Xno4_3;
	wire w_dff_B_JwMiTnx43_3;
	wire w_dff_B_5oOo1v0z3_3;
	wire w_dff_B_JDfv641l3_3;
	wire w_dff_B_ZOBIZjc95_3;
	wire w_dff_B_aM2RjltO6_3;
	wire w_dff_B_QKUuJj6k5_3;
	wire w_dff_B_PhKd6gim7_3;
	wire w_dff_B_ABthXCsD1_3;
	wire w_dff_A_zpocZClW1_0;
	wire w_dff_A_kzb2hd9g2_0;
	wire w_dff_A_tPvQ50N17_0;
	wire w_dff_A_0iwGuBup5_0;
	wire w_dff_A_1JkvPatN8_0;
	wire w_dff_A_dnb0bL5J6_0;
	wire w_dff_A_noxCN2xs0_0;
	wire w_dff_A_cmziJ8rH0_0;
	wire w_dff_A_PTOOPFEP7_0;
	wire w_dff_A_5uLjN7M02_0;
	wire w_dff_A_U89RAlI01_0;
	wire w_dff_A_jZCOVcyN5_0;
	wire w_dff_A_EUiMTc6g9_0;
	wire w_dff_A_3qGi0CTf2_0;
	wire w_dff_A_j20f81iP6_0;
	wire w_dff_A_dsLaRl0i4_1;
	wire w_dff_A_JPs7umaD0_1;
	wire w_dff_A_QPQ4pMGT8_1;
	wire w_dff_A_boM86YGm1_1;
	wire w_dff_A_essMvL466_1;
	wire w_dff_A_TMAstcUh7_1;
	wire w_dff_A_NAHX9de54_1;
	wire w_dff_A_Bi0O1SEm3_1;
	wire w_dff_A_kyiRyx2l1_1;
	wire w_dff_A_BVOeA0sq0_1;
	wire w_dff_A_wUT6urke0_1;
	wire w_dff_A_6Rsph3Hg4_1;
	wire w_dff_A_8MQaLwTx7_2;
	wire w_dff_A_bbIVZ2GE6_2;
	wire w_dff_A_BLAfd50W6_2;
	wire w_dff_A_6a1B3lW21_2;
	wire w_dff_A_lF46ez6K4_2;
	wire w_dff_A_CtgLOVyt6_2;
	wire w_dff_A_NVQNUgLU8_2;
	wire w_dff_A_41mZbeXE9_2;
	wire w_dff_A_i8Bpewt29_2;
	wire w_dff_A_KObVYEQX8_2;
	wire w_dff_A_QKLFT9Vj5_2;
	wire w_dff_A_9q7KrHWp5_2;
	wire w_dff_A_lFjUfkaK7_2;
	wire w_dff_A_BnUQP51w1_2;
	wire w_dff_A_TcigiV841_2;
	wire w_dff_A_eJ8WeTly5_1;
	wire w_dff_A_kB4SSVFo8_1;
	wire w_dff_A_q5XNO7724_1;
	wire w_dff_A_KbNwem6D8_1;
	wire w_dff_A_Bcs8i3FC8_1;
	wire w_dff_A_L04gicix8_1;
	wire w_dff_A_oxWsyVxS3_1;
	wire w_dff_A_rBR9K8g67_1;
	wire w_dff_A_PE3lYjSi0_1;
	wire w_dff_A_DNaSOExD5_1;
	wire w_dff_A_lqCeg8BL0_1;
	wire w_dff_A_56Wg1G6r6_1;
	wire w_dff_A_dI8Hm2Kf7_1;
	wire w_dff_A_xR0wmvLR0_1;
	wire w_dff_A_Y3lDFskQ4_1;
	wire w_dff_A_fyg1Pvi90_1;
	wire w_dff_A_9rtk9RnC4_2;
	wire w_dff_B_rfC0uYMu3_3;
	wire w_dff_A_MwqRsx0w6_2;
	wire w_dff_A_SMnVsTUa9_0;
	wire w_dff_A_fve125FU0_0;
	wire w_dff_A_OQIf7Pgw2_0;
	wire w_dff_A_dpkeVIAL3_0;
	wire w_dff_A_GI9QouZV0_0;
	wire w_dff_A_ujBRfDho2_0;
	wire w_dff_A_bHBPXyAM6_0;
	wire w_dff_A_y0S1Air87_2;
	wire w_dff_A_XU688eYr5_0;
	wire w_dff_A_8USHUJhp6_0;
	wire w_dff_A_987J6CRB3_0;
	wire w_dff_A_Eq74QE4D7_0;
	wire w_dff_A_KyyL9Txj4_0;
	wire w_dff_A_0YMYoiDk5_0;
	wire w_dff_A_d4RSwXSv6_0;
	wire w_dff_A_N02qW1yA7_2;
	wire w_dff_A_EiKuOHs69_0;
	wire w_dff_A_k0UDo0I42_0;
	wire w_dff_A_e86XZncz6_0;
	wire w_dff_A_he6nAg600_0;
	wire w_dff_A_UtqTR2KL3_0;
	wire w_dff_A_6uNN18sl4_0;
	wire w_dff_A_TRxK1wIw3_0;
	wire w_dff_A_DlpRYtCa6_2;
	wire w_dff_A_HEvIMrhO8_0;
	wire w_dff_A_z5QkHR330_0;
	wire w_dff_A_BWrBfszh5_0;
	wire w_dff_A_7arxUe0W1_0;
	wire w_dff_A_1vEWcUA41_0;
	wire w_dff_A_odBtbIM31_0;
	wire w_dff_A_q9vckpvG5_0;
	wire w_dff_A_apRAkZg53_2;
	wire w_dff_A_uHEe57WI6_0;
	wire w_dff_A_FBgM1fRJ7_0;
	wire w_dff_A_W1YKKNVp8_0;
	wire w_dff_A_46LN5FKU6_0;
	wire w_dff_A_L0YRChQu4_0;
	wire w_dff_A_7jMzdGF19_0;
	wire w_dff_A_APq4wjnn3_0;
	wire w_dff_A_R0NrbBNi0_2;
	wire w_dff_A_0CGTH1bS1_0;
	wire w_dff_A_MiuQvP6e8_0;
	wire w_dff_A_Z6zVLBMN3_0;
	wire w_dff_A_zV37IviQ9_0;
	wire w_dff_A_XCrhnlh61_0;
	wire w_dff_A_srCUVw1T3_0;
	wire w_dff_A_BhoUwC8V8_0;
	wire w_dff_A_CDdRnRdY1_2;
	wire w_dff_A_TwZMTknQ6_0;
	wire w_dff_A_r50859xe3_0;
	wire w_dff_A_duzyz5qb1_0;
	wire w_dff_A_Y4lLNQqh1_0;
	wire w_dff_A_KXNZUKy93_0;
	wire w_dff_A_rH4t5jcW6_0;
	wire w_dff_A_B8RMUIgp3_0;
	wire w_dff_A_E06fr8vG6_2;
	wire w_dff_A_sXNTBL0W1_0;
	wire w_dff_A_jQHsaafC8_0;
	wire w_dff_A_sjmTYC5l1_0;
	wire w_dff_A_Zuo1Q2Tg7_0;
	wire w_dff_A_8IxNtXV07_0;
	wire w_dff_A_pXdMvCaZ5_0;
	wire w_dff_A_rSjKCHNd3_0;
	wire w_dff_A_YMIk41gS8_2;
	wire w_dff_A_4MA2UY1h2_0;
	wire w_dff_A_DzfdTRno5_0;
	wire w_dff_A_3gpJ598J6_0;
	wire w_dff_A_5a5NmolD0_0;
	wire w_dff_A_LNaBgbuO0_0;
	wire w_dff_A_KptFUmx34_0;
	wire w_dff_A_YLO0uwsg6_0;
	wire w_dff_A_s8rXBoX56_2;
	wire w_dff_A_ZZdXydGm6_0;
	wire w_dff_A_QqLKm64w6_0;
	wire w_dff_A_eJCCopJa8_0;
	wire w_dff_A_z5WKZ6gX1_0;
	wire w_dff_A_QfYmXPBM9_0;
	wire w_dff_A_dVTLmbqY8_0;
	wire w_dff_A_Woh6OdVs2_0;
	wire w_dff_A_48L5gWb59_2;
	wire w_dff_A_pFBbqCNZ4_0;
	wire w_dff_A_FEyCJMKm5_0;
	wire w_dff_A_KoVzu7q37_0;
	wire w_dff_A_O11JJmVx6_0;
	wire w_dff_A_65Oxlssu0_0;
	wire w_dff_A_fvL8DYi59_0;
	wire w_dff_A_ve0cAdrm6_2;
	wire w_dff_A_RkFR6puO5_0;
	wire w_dff_A_hrAlhNAm1_0;
	wire w_dff_A_5WpE3FLY3_0;
	wire w_dff_A_q0ckrtDo0_0;
	wire w_dff_A_jaUi27hL0_0;
	wire w_dff_A_3exUiFpL3_0;
	wire w_dff_A_UjaTMIZF1_0;
	wire w_dff_A_pvSnXxJb3_2;
	wire w_dff_A_BURVCN1F8_0;
	wire w_dff_A_4AI7CPcV2_0;
	wire w_dff_A_cFslUK5m3_0;
	wire w_dff_A_bnlqfMaz2_0;
	wire w_dff_A_66F1CsVM0_0;
	wire w_dff_A_iY3FJa145_0;
	wire w_dff_A_2uHjnuT57_0;
	wire w_dff_A_9hMXUQKg7_2;
	wire w_dff_A_uOSfjerm5_0;
	wire w_dff_A_S2Tp7smu0_0;
	wire w_dff_A_HinQTAFs2_0;
	wire w_dff_A_WZS4Vqqr7_0;
	wire w_dff_A_8KdmLDuJ5_0;
	wire w_dff_A_6hExMG0z6_0;
	wire w_dff_A_9S8T0T9S2_0;
	wire w_dff_A_H0wbY1Ub8_2;
	wire w_dff_A_5Bs10Pmm9_0;
	wire w_dff_A_xevfPlMV8_0;
	wire w_dff_A_gCTlPJdx7_0;
	wire w_dff_A_pQ3YMCOW1_0;
	wire w_dff_A_s3ze39kW7_0;
	wire w_dff_A_yvSMQFQ96_0;
	wire w_dff_A_qGGumymi0_0;
	wire w_dff_A_K9N8MOyh8_2;
	wire w_dff_A_vxdStgLY0_0;
	wire w_dff_A_gIDHvzis8_0;
	wire w_dff_A_gAgSSfCd1_0;
	wire w_dff_A_C5lsZQZP3_0;
	wire w_dff_A_KIFz7CH72_0;
	wire w_dff_A_tGRE1uAg3_0;
	wire w_dff_A_ADq0GnWf3_0;
	wire w_dff_A_NWXt4Snf1_2;
	wire w_dff_A_jrsgWhlw6_2;
	wire w_dff_A_FggnYhHZ2_0;
	wire w_dff_A_bfIBpwvT2_2;
	wire w_dff_A_Xaaac5Zg9_0;
	wire w_dff_A_CR8MmAXU9_2;
	jnot g000(.din(w_G902_3[2]),.dout(n58),.clk(gclk));
	jnot g001(.din(w_G221_0[1]),.dout(n59),.clk(gclk));
	jnot g002(.din(w_G234_1[1]),.dout(n60),.clk(gclk));
	jor g003(.dina(w_G953_2[1]),.dinb(n60),.dout(n61),.clk(gclk));
	jor g004(.dina(n61),.dinb(w_dff_B_LDZoSPUp5_1),.dout(n62),.clk(gclk));
	jnot g005(.din(w_G110_0[2]),.dout(n63),.clk(gclk));
	jxor g006(.dina(w_G119_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jxor g007(.dina(w_dff_B_XiehfK7Z2_0),.dinb(n62),.dout(n65),.clk(gclk));
	jxor g008(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n66),.clk(gclk));
	jxor g009(.dina(w_n66_0[1]),.dinb(w_G146_0[2]),.dout(n67),.clk(gclk));
	jxor g010(.dina(w_G137_0[2]),.dinb(w_G128_0[2]),.dout(n68),.clk(gclk));
	jxor g011(.dina(w_dff_B_LJSWXHrT7_0),.dinb(w_n67_0[1]),.dout(n69),.clk(gclk));
	jxor g012(.dina(w_dff_B_r8oAmEr11_0),.dinb(n65),.dout(n70),.clk(gclk));
	jand g013(.dina(w_n70_0[1]),.dinb(w_n58_2[2]),.dout(n71),.clk(gclk));
	jand g014(.dina(w_n58_2[1]),.dinb(w_G234_1[0]),.dout(n72),.clk(gclk));
	jnot g015(.din(n72),.dout(n73),.clk(gclk));
	jand g016(.dina(w_n73_0[1]),.dinb(w_G217_0[2]),.dout(n74),.clk(gclk));
	jnot g017(.din(w_n74_0[1]),.dout(n75),.clk(gclk));
	jxor g018(.dina(w_dff_B_4qFwiVGm8_0),.dinb(w_n71_0[1]),.dout(n76),.clk(gclk));
	jxor g019(.dina(w_G143_0[2]),.dinb(w_G128_0[1]),.dout(n77),.clk(gclk));
	jxor g020(.dina(w_n77_0[1]),.dinb(w_G146_0[1]),.dout(n78),.clk(gclk));
	jxor g021(.dina(w_G137_0[1]),.dinb(w_G134_0[2]),.dout(n79),.clk(gclk));
	jxor g022(.dina(n79),.dinb(w_G131_0[2]),.dout(n80),.clk(gclk));
	jxor g023(.dina(n80),.dinb(w_n78_0[1]),.dout(n81),.clk(gclk));
	jnot g024(.din(w_G113_0[2]),.dout(n82),.clk(gclk));
	jxor g025(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g026(.dina(n83),.dinb(n82),.dout(n84),.clk(gclk));
	jnot g027(.din(w_G210_0[2]),.dout(n85),.clk(gclk));
	jor g028(.dina(w_G953_2[0]),.dinb(w_G237_0[2]),.dout(n86),.clk(gclk));
	jor g029(.dina(w_n86_0[1]),.dinb(n85),.dout(n87),.clk(gclk));
	jxor g030(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g031(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g032(.dina(n89),.dinb(w_n81_0[2]),.dout(n90),.clk(gclk));
	jand g033(.dina(w_n90_0[1]),.dinb(w_n58_2[0]),.dout(n91),.clk(gclk));
	jxor g034(.dina(w_n91_0[1]),.dinb(w_G472_0[2]),.dout(n92),.clk(gclk));
	jand g035(.dina(w_n92_1[1]),.dinb(w_n76_1[2]),.dout(n93),.clk(gclk));
	jor g036(.dina(w_G902_3[1]),.dinb(w_G237_0[1]),.dout(n94),.clk(gclk));
	jand g037(.dina(w_n94_0[1]),.dinb(w_G214_0[1]),.dout(n95),.clk(gclk));
	jnot g038(.din(w_n95_1[1]),.dout(n96),.clk(gclk));
	jnot g039(.din(w_G101_0[1]),.dout(n97),.clk(gclk));
	jxor g040(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n98),.clk(gclk));
	jxor g041(.dina(n98),.dinb(n97),.dout(n99),.clk(gclk));
	jxor g042(.dina(w_n99_0[1]),.dinb(w_n84_0[0]),.dout(n100),.clk(gclk));
	jxor g043(.dina(w_G122_1[1]),.dinb(w_G110_0[1]),.dout(n101),.clk(gclk));
	jxor g044(.dina(w_dff_B_JxaDq2Ff9_0),.dinb(n100),.dout(n102),.clk(gclk));
	jnot g045(.din(w_G953_1[2]),.dout(n103),.clk(gclk));
	jand g046(.dina(w_n103_3[2]),.dinb(w_G224_0[1]),.dout(n104),.clk(gclk));
	jxor g047(.dina(w_n78_0[0]),.dinb(w_G125_0[1]),.dout(n105),.clk(gclk));
	jxor g048(.dina(n105),.dinb(w_dff_B_aFnTQLtg1_1),.dout(n106),.clk(gclk));
	jxor g049(.dina(n106),.dinb(w_n102_0[1]),.dout(n107),.clk(gclk));
	jand g050(.dina(w_n107_0[1]),.dinb(w_n58_1[2]),.dout(n108),.clk(gclk));
	jand g051(.dina(w_n94_0[0]),.dinb(w_G210_0[1]),.dout(n109),.clk(gclk));
	jxor g052(.dina(w_n109_0[1]),.dinb(w_n108_0[1]),.dout(n110),.clk(gclk));
	jand g053(.dina(w_n110_0[1]),.dinb(w_n96_0[2]),.dout(n111),.clk(gclk));
	jand g054(.dina(w_n73_0[0]),.dinb(w_G221_0[0]),.dout(n112),.clk(gclk));
	jnot g055(.din(w_n112_1[1]),.dout(n113),.clk(gclk));
	jand g056(.dina(w_n103_3[1]),.dinb(w_G227_0[1]),.dout(n114),.clk(gclk));
	jxor g057(.dina(w_G140_0[1]),.dinb(w_n63_0[0]),.dout(n115),.clk(gclk));
	jxor g058(.dina(n115),.dinb(n114),.dout(n116),.clk(gclk));
	jxor g059(.dina(n116),.dinb(w_n99_0[0]),.dout(n117),.clk(gclk));
	jxor g060(.dina(n117),.dinb(w_n81_0[1]),.dout(n118),.clk(gclk));
	jand g061(.dina(w_n118_0[1]),.dinb(w_n58_1[1]),.dout(n119),.clk(gclk));
	jxor g062(.dina(w_n119_0[1]),.dinb(w_G469_0[2]),.dout(n120),.clk(gclk));
	jand g063(.dina(w_n120_0[1]),.dinb(w_n113_0[2]),.dout(n121),.clk(gclk));
	jand g064(.dina(w_n121_0[1]),.dinb(w_n111_0[1]),.dout(n122),.clk(gclk));
	jor g065(.dina(w_n103_3[0]),.dinb(w_G898_0[1]),.dout(n123),.clk(gclk));
	jnot g066(.din(n123),.dout(n124),.clk(gclk));
	jand g067(.dina(w_G237_0[0]),.dinb(w_G234_0[2]),.dout(n125),.clk(gclk));
	jnot g068(.din(n125),.dout(n126),.clk(gclk));
	jand g069(.dina(w_n126_0[1]),.dinb(w_G902_3[0]),.dout(n127),.clk(gclk));
	jand g070(.dina(w_n127_0[1]),.dinb(w_n124_0[1]),.dout(n128),.clk(gclk));
	jand g071(.dina(w_n126_0[0]),.dinb(w_G952_0[2]),.dout(n129),.clk(gclk));
	jand g072(.dina(n129),.dinb(w_n103_2[2]),.dout(n130),.clk(gclk));
	jor g073(.dina(w_n130_1[1]),.dinb(n128),.dout(n131),.clk(gclk));
	jnot g074(.din(w_G478_0[2]),.dout(n132),.clk(gclk));
	jxor g075(.dina(w_n77_0[0]),.dinb(w_G134_0[1]),.dout(n133),.clk(gclk));
	jand g076(.dina(w_n103_2[1]),.dinb(w_G234_0[1]),.dout(n134),.clk(gclk));
	jand g077(.dina(n134),.dinb(w_G217_0[1]),.dout(n135),.clk(gclk));
	jxor g078(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n136),.clk(gclk));
	jxor g079(.dina(n136),.dinb(w_G107_0[1]),.dout(n137),.clk(gclk));
	jxor g080(.dina(w_dff_B_bm62cSlV3_0),.dinb(n135),.dout(n138),.clk(gclk));
	jxor g081(.dina(n138),.dinb(w_dff_B_CN858ycW5_1),.dout(n139),.clk(gclk));
	jand g082(.dina(w_n139_0[1]),.dinb(w_n58_1[0]),.dout(n140),.clk(gclk));
	jxor g083(.dina(w_n140_0[1]),.dinb(w_dff_B_kbcpQt2j9_1),.dout(n141),.clk(gclk));
	jnot g084(.din(w_G475_0[2]),.dout(n142),.clk(gclk));
	jxor g085(.dina(w_G122_0[2]),.dinb(w_G113_0[1]),.dout(n143),.clk(gclk));
	jxor g086(.dina(n143),.dinb(w_G104_0[1]),.dout(n144),.clk(gclk));
	jnot g087(.din(w_G214_0[0]),.dout(n145),.clk(gclk));
	jor g088(.dina(w_n86_0[0]),.dinb(n145),.dout(n146),.clk(gclk));
	jnot g089(.din(w_G131_0[1]),.dout(n147),.clk(gclk));
	jxor g090(.dina(w_G143_0[1]),.dinb(n147),.dout(n148),.clk(gclk));
	jxor g091(.dina(n148),.dinb(n146),.dout(n149),.clk(gclk));
	jxor g092(.dina(n149),.dinb(w_n67_0[0]),.dout(n150),.clk(gclk));
	jxor g093(.dina(n150),.dinb(w_dff_B_Ny6Ilyp92_1),.dout(n151),.clk(gclk));
	jand g094(.dina(w_n151_0[2]),.dinb(w_n58_0[2]),.dout(n152),.clk(gclk));
	jxor g095(.dina(w_n152_0[1]),.dinb(w_dff_B_4GcJj6UK9_1),.dout(n153),.clk(gclk));
	jand g096(.dina(w_n153_1[1]),.dinb(w_n141_1[1]),.dout(n154),.clk(gclk));
	jand g097(.dina(w_n154_1[1]),.dinb(w_n131_1[2]),.dout(n155),.clk(gclk));
	jand g098(.dina(w_n155_0[1]),.dinb(w_n122_1[1]),.dout(n156),.clk(gclk));
	jand g099(.dina(w_n156_0[1]),.dinb(w_n93_1[1]),.dout(n157),.clk(gclk));
	jxor g100(.dina(w_n157_0[1]),.dinb(w_G101_0[0]),.dout(w_dff_A_MwqRsx0w6_2),.clk(gclk));
	jnot g101(.din(w_G472_0[1]),.dout(n159),.clk(gclk));
	jxor g102(.dina(w_n91_0[0]),.dinb(w_dff_B_P7OwcfVU5_1),.dout(n160),.clk(gclk));
	jand g103(.dina(w_n160_1[2]),.dinb(w_n76_1[1]),.dout(n161),.clk(gclk));
	jand g104(.dina(w_n161_1[1]),.dinb(w_n122_1[0]),.dout(n162),.clk(gclk));
	jxor g105(.dina(w_n152_0[0]),.dinb(w_G475_0[1]),.dout(n163),.clk(gclk));
	jand g106(.dina(w_n163_1[1]),.dinb(w_n141_1[0]),.dout(n164),.clk(gclk));
	jand g107(.dina(w_n164_0[1]),.dinb(w_n131_1[1]),.dout(n165),.clk(gclk));
	jand g108(.dina(w_n165_0[2]),.dinb(w_n162_0[1]),.dout(n166),.clk(gclk));
	jxor g109(.dina(w_n166_0[1]),.dinb(w_G104_0[0]),.dout(w_dff_A_y0S1Air87_2),.clk(gclk));
	jxor g110(.dina(w_n140_0[0]),.dinb(w_G478_0[1]),.dout(n168),.clk(gclk));
	jand g111(.dina(w_n153_1[0]),.dinb(w_n168_1[1]),.dout(n169),.clk(gclk));
	jand g112(.dina(w_n169_0[1]),.dinb(w_n131_1[0]),.dout(n170),.clk(gclk));
	jand g113(.dina(w_n170_0[1]),.dinb(w_n162_0[0]),.dout(n171),.clk(gclk));
	jxor g114(.dina(w_n171_0[1]),.dinb(w_G107_0[0]),.dout(w_dff_A_N02qW1yA7_2),.clk(gclk));
	jxor g115(.dina(w_n74_0[0]),.dinb(w_n71_0[0]),.dout(n173),.clk(gclk));
	jand g116(.dina(w_n160_1[1]),.dinb(w_n173_1[1]),.dout(n174),.clk(gclk));
	jand g117(.dina(w_n174_0[1]),.dinb(w_n156_0[0]),.dout(n175),.clk(gclk));
	jxor g118(.dina(w_n175_0[1]),.dinb(w_G110_0[0]),.dout(w_dff_A_DlpRYtCa6_2),.clk(gclk));
	jand g119(.dina(w_n92_1[0]),.dinb(w_n173_1[0]),.dout(n177),.clk(gclk));
	jand g120(.dina(w_n177_0[2]),.dinb(w_n122_0[2]),.dout(n178),.clk(gclk));
	jor g121(.dina(w_n103_2[0]),.dinb(w_G900_0[1]),.dout(n179),.clk(gclk));
	jnot g122(.din(n179),.dout(n180),.clk(gclk));
	jand g123(.dina(w_n180_0[1]),.dinb(w_n127_0[0]),.dout(n181),.clk(gclk));
	jor g124(.dina(n181),.dinb(w_n130_1[0]),.dout(n182),.clk(gclk));
	jand g125(.dina(w_n182_1[2]),.dinb(w_n169_0[0]),.dout(n183),.clk(gclk));
	jand g126(.dina(w_n183_0[2]),.dinb(w_n178_0[1]),.dout(n184),.clk(gclk));
	jxor g127(.dina(w_n184_0[1]),.dinb(w_G128_0[0]),.dout(w_dff_A_apRAkZg53_2),.clk(gclk));
	jand g128(.dina(w_n163_1[0]),.dinb(w_n168_1[0]),.dout(n186),.clk(gclk));
	jand g129(.dina(w_n186_0[1]),.dinb(w_n93_1[0]),.dout(n187),.clk(gclk));
	jand g130(.dina(n187),.dinb(w_n182_1[1]),.dout(n188),.clk(gclk));
	jand g131(.dina(n188),.dinb(w_n122_0[1]),.dout(n189),.clk(gclk));
	jxor g132(.dina(w_n189_0[1]),.dinb(w_G143_0[0]),.dout(w_dff_A_R0NrbBNi0_2),.clk(gclk));
	jand g133(.dina(w_n182_1[0]),.dinb(w_n164_0[0]),.dout(n191),.clk(gclk));
	jand g134(.dina(w_n191_0[2]),.dinb(w_n178_0[0]),.dout(n192),.clk(gclk));
	jxor g135(.dina(w_n192_0[2]),.dinb(w_G146_0[0]),.dout(w_dff_A_CDdRnRdY1_2),.clk(gclk));
	jnot g136(.din(w_G469_0[1]),.dout(n194),.clk(gclk));
	jxor g137(.dina(w_n119_0[0]),.dinb(w_dff_B_NsDCSFXi4_1),.dout(n195),.clk(gclk));
	jand g138(.dina(w_n195_0[2]),.dinb(w_n113_0[1]),.dout(n196),.clk(gclk));
	jand g139(.dina(n196),.dinb(w_n111_0[0]),.dout(n197),.clk(gclk));
	jand g140(.dina(w_n197_1[1]),.dinb(w_n93_0[2]),.dout(n198),.clk(gclk));
	jand g141(.dina(w_n198_0[1]),.dinb(w_n165_0[1]),.dout(n199),.clk(gclk));
	jxor g142(.dina(w_n199_0[2]),.dinb(w_G113_0[0]),.dout(w_dff_A_E06fr8vG6_2),.clk(gclk));
	jand g143(.dina(w_n198_0[0]),.dinb(w_n170_0[0]),.dout(n201),.clk(gclk));
	jxor g144(.dina(w_n201_0[1]),.dinb(w_G116_0[0]),.dout(w_dff_A_YMIk41gS8_2),.clk(gclk));
	jand g145(.dina(w_n177_0[1]),.dinb(w_n155_0[0]),.dout(n203),.clk(gclk));
	jand g146(.dina(n203),.dinb(w_n197_1[0]),.dout(n204),.clk(gclk));
	jxor g147(.dina(w_n204_0[1]),.dinb(w_G119_0[0]),.dout(w_dff_A_s8rXBoX56_2),.clk(gclk));
	jand g148(.dina(w_n197_0[2]),.dinb(w_n161_1[0]),.dout(n206),.clk(gclk));
	jand g149(.dina(w_n206_0[1]),.dinb(w_n131_0[2]),.dout(n207),.clk(gclk));
	jand g150(.dina(n207),.dinb(w_n186_0[0]),.dout(n208),.clk(gclk));
	jxor g151(.dina(w_n208_0[1]),.dinb(w_G122_0[1]),.dout(w_dff_A_48L5gWb59_2),.clk(gclk));
	jand g152(.dina(w_n191_0[1]),.dinb(w_n174_0[0]),.dout(n210),.clk(gclk));
	jand g153(.dina(w_n210_0[1]),.dinb(w_n197_0[1]),.dout(n211),.clk(gclk));
	jxor g154(.dina(w_n211_0[1]),.dinb(w_G125_0[0]),.dout(w_dff_A_ve0cAdrm6_2),.clk(gclk));
	jnot g155(.din(w_n109_0[0]),.dout(n213),.clk(gclk));
	jxor g156(.dina(w_dff_B_2muhCsUb1_0),.dinb(w_n108_0[0]),.dout(n214),.clk(gclk));
	jand g157(.dina(w_n214_0[2]),.dinb(w_n96_0[1]),.dout(n215),.clk(gclk));
	jand g158(.dina(n215),.dinb(w_n121_0[0]),.dout(n216),.clk(gclk));
	jand g159(.dina(w_n216_1[1]),.dinb(w_n93_0[1]),.dout(n217),.clk(gclk));
	jand g160(.dina(w_n217_0[1]),.dinb(w_n191_0[0]),.dout(n218),.clk(gclk));
	jxor g161(.dina(w_n218_0[1]),.dinb(w_G131_0[0]),.dout(w_dff_A_pvSnXxJb3_2),.clk(gclk));
	jand g162(.dina(w_n217_0[0]),.dinb(w_n183_0[1]),.dout(n220),.clk(gclk));
	jxor g163(.dina(w_n220_0[1]),.dinb(w_G134_0[0]),.dout(w_dff_A_9hMXUQKg7_2),.clk(gclk));
	jand g164(.dina(w_n177_0[0]),.dinb(w_n154_1[0]),.dout(n222),.clk(gclk));
	jand g165(.dina(n222),.dinb(w_n182_0[2]),.dout(n223),.clk(gclk));
	jand g166(.dina(n223),.dinb(w_n216_1[0]),.dout(n224),.clk(gclk));
	jxor g167(.dina(w_n224_0[1]),.dinb(w_G137_0[0]),.dout(w_dff_A_H0wbY1Ub8_2),.clk(gclk));
	jand g168(.dina(w_n216_0[2]),.dinb(w_n210_0[0]),.dout(n226),.clk(gclk));
	jxor g169(.dina(w_n226_0[1]),.dinb(w_G140_0[0]),.dout(w_dff_A_K9N8MOyh8_2),.clk(gclk));
	jor g170(.dina(w_n171_0[0]),.dinb(w_n157_0[0]),.dout(n228),.clk(gclk));
	jor g171(.dina(n228),.dinb(w_n166_0[0]),.dout(n229),.clk(gclk));
	jor g172(.dina(n229),.dinb(w_n208_0[0]),.dout(n230),.clk(gclk));
	jor g173(.dina(w_n204_0[0]),.dinb(w_n201_0[0]),.dout(n231),.clk(gclk));
	jor g174(.dina(n231),.dinb(w_n175_0[0]),.dout(n232),.clk(gclk));
	jor g175(.dina(n232),.dinb(w_n199_0[1]),.dout(n233),.clk(gclk));
	jor g176(.dina(n233),.dinb(n230),.dout(n234),.clk(gclk));
	jor g177(.dina(w_n226_0[0]),.dinb(w_n224_0[0]),.dout(n235),.clk(gclk));
	jor g178(.dina(n235),.dinb(w_n192_0[1]),.dout(n236),.clk(gclk));
	jor g179(.dina(w_n220_0[0]),.dinb(w_n218_0[0]),.dout(n237),.clk(gclk));
	jor g180(.dina(w_n211_0[0]),.dinb(w_n189_0[0]),.dout(n238),.clk(gclk));
	jor g181(.dina(n238),.dinb(w_n184_0[0]),.dout(n239),.clk(gclk));
	jor g182(.dina(n239),.dinb(w_dff_B_JC95DaZ65_1),.dout(n240),.clk(gclk));
	jor g183(.dina(n240),.dinb(w_dff_B_RqHLDa1b8_1),.dout(n241),.clk(gclk));
	jor g184(.dina(n241),.dinb(n234),.dout(n242),.clk(gclk));
	jand g185(.dina(w_n195_0[1]),.dinb(w_n214_0[1]),.dout(n243),.clk(gclk));
	jxor g186(.dina(w_n112_1[0]),.dinb(w_n95_1[0]),.dout(n244),.clk(gclk));
	jand g187(.dina(w_dff_B_E3zHyqyO6_0),.dinb(w_n243_0[1]),.dout(n245),.clk(gclk));
	jor g188(.dina(n245),.dinb(w_n216_0[1]),.dout(n246),.clk(gclk));
	jand g189(.dina(n246),.dinb(w_n161_0[2]),.dout(n247),.clk(gclk));
	jand g190(.dina(w_n113_0[0]),.dinb(w_n96_0[0]),.dout(n248),.clk(gclk));
	jand g191(.dina(w_dff_B_JBz7l3hc8_0),.dinb(w_n243_0[0]),.dout(n249),.clk(gclk));
	jxor g192(.dina(w_n160_1[0]),.dinb(w_n76_1[0]),.dout(n250),.clk(gclk));
	jand g193(.dina(w_dff_B_eggdHZDG6_0),.dinb(w_n249_0[1]),.dout(n251),.clk(gclk));
	jor g194(.dina(n251),.dinb(w_n206_0[0]),.dout(n252),.clk(gclk));
	jor g195(.dina(n252),.dinb(n247),.dout(n253),.clk(gclk));
	jand g196(.dina(n253),.dinb(w_n154_0[2]),.dout(n254),.clk(gclk));
	jand g197(.dina(n254),.dinb(w_n130_0[2]),.dout(n255),.clk(gclk));
	jor g198(.dina(w_dff_B_HucuwSJG9_0),.dinb(w_n242_2[2]),.dout(n256),.clk(gclk));
	jand g199(.dina(n256),.dinb(w_G952_0[1]),.dout(n257),.clk(gclk));
	jor g200(.dina(w_n153_0[2]),.dinb(w_n141_0[2]),.dout(n258),.clk(gclk));
	jor g201(.dina(w_n154_0[1]),.dinb(w_n130_0[1]),.dout(n259),.clk(gclk));
	jand g202(.dina(n259),.dinb(w_n258_0[2]),.dout(n260),.clk(gclk));
	jand g203(.dina(n260),.dinb(w_n161_0[1]),.dout(n261),.clk(gclk));
	jand g204(.dina(n261),.dinb(w_n249_0[0]),.dout(n262),.clk(gclk));
	jor g205(.dina(n262),.dinb(w_G953_1[1]),.dout(n263),.clk(gclk));
	jor g206(.dina(w_dff_B_X1XwYjW90_0),.dinb(n257),.dout(w_dff_A_NWXt4Snf1_2),.clk(gclk));
	jor g207(.dina(w_n103_1[2]),.dinb(w_G952_0[0]),.dout(n265),.clk(gclk));
	jand g208(.dina(w_n242_2[1]),.dinb(w_G210_0[0]),.dout(n266),.clk(gclk));
	jand g209(.dina(n266),.dinb(w_G902_2[2]),.dout(n267),.clk(gclk));
	jxor g210(.dina(n267),.dinb(w_n107_0[0]),.dout(n268),.clk(gclk));
	jand g211(.dina(n268),.dinb(w_n265_2[1]),.dout(G51),.clk(gclk));
	jand g212(.dina(w_n242_2[0]),.dinb(w_G469_0[0]),.dout(n270),.clk(gclk));
	jand g213(.dina(n270),.dinb(w_G902_2[1]),.dout(n271),.clk(gclk));
	jxor g214(.dina(n271),.dinb(w_n118_0[0]),.dout(n272),.clk(gclk));
	jand g215(.dina(n272),.dinb(w_n265_2[0]),.dout(G54),.clk(gclk));
	jand g216(.dina(w_G902_2[0]),.dinb(w_G475_0[0]),.dout(n274),.clk(gclk));
	jand g217(.dina(w_n274_0[1]),.dinb(w_n242_1[2]),.dout(n275),.clk(gclk));
	jor g218(.dina(n275),.dinb(w_n151_0[1]),.dout(n276),.clk(gclk));
	jnot g219(.din(w_n151_0[0]),.dout(n277),.clk(gclk));
	jnot g220(.din(w_n131_0[1]),.dout(n278),.clk(gclk));
	jor g221(.dina(w_n92_0[2]),.dinb(w_n173_0[2]),.dout(n279),.clk(gclk));
	jor g222(.dina(w_n214_0[0]),.dinb(w_n95_0[2]),.dout(n280),.clk(gclk));
	jor g223(.dina(w_n120_0[0]),.dinb(w_n112_0[2]),.dout(n281),.clk(gclk));
	jor g224(.dina(n281),.dinb(w_n280_0[1]),.dout(n282),.clk(gclk));
	jor g225(.dina(w_n282_1[1]),.dinb(w_n279_0[1]),.dout(n283),.clk(gclk));
	jor g226(.dina(n283),.dinb(w_n278_0[2]),.dout(n284),.clk(gclk));
	jor g227(.dina(n284),.dinb(w_n258_0[1]),.dout(n285),.clk(gclk));
	jor g228(.dina(w_n195_0[0]),.dinb(w_n112_0[1]),.dout(n286),.clk(gclk));
	jor g229(.dina(w_n286_0[1]),.dinb(w_n280_0[0]),.dout(n287),.clk(gclk));
	jor g230(.dina(w_n279_0[0]),.dinb(w_n287_1[1]),.dout(n288),.clk(gclk));
	jnot g231(.din(w_n165_0[0]),.dout(n289),.clk(gclk));
	jor g232(.dina(n289),.dinb(w_n288_0[1]),.dout(n290),.clk(gclk));
	jor g233(.dina(w_n160_0[2]),.dinb(w_n173_0[1]),.dout(n291),.clk(gclk));
	jor g234(.dina(w_n163_0[2]),.dinb(w_n168_0[2]),.dout(n292),.clk(gclk));
	jor g235(.dina(w_n292_0[1]),.dinb(w_n278_0[1]),.dout(n293),.clk(gclk));
	jor g236(.dina(w_n293_0[1]),.dinb(w_n287_1[0]),.dout(n294),.clk(gclk));
	jor g237(.dina(w_n294_0[1]),.dinb(w_n291_1[1]),.dout(n295),.clk(gclk));
	jor g238(.dina(w_n163_0[1]),.dinb(w_n141_0[1]),.dout(n296),.clk(gclk));
	jor g239(.dina(n296),.dinb(w_n278_0[0]),.dout(n297),.clk(gclk));
	jor g240(.dina(w_n297_0[1]),.dinb(w_n288_0[0]),.dout(n298),.clk(gclk));
	jand g241(.dina(n298),.dinb(n295),.dout(n299),.clk(gclk));
	jand g242(.dina(n299),.dinb(w_dff_B_BvqV64tH2_1),.dout(n300),.clk(gclk));
	jand g243(.dina(n300),.dinb(w_dff_B_o1k8CBxA6_1),.dout(n301),.clk(gclk));
	jnot g244(.din(w_n199_0[0]),.dout(n302),.clk(gclk));
	jor g245(.dina(w_n92_0[1]),.dinb(w_n76_0[2]),.dout(n303),.clk(gclk));
	jor g246(.dina(w_n303_0[1]),.dinb(w_n294_0[0]),.dout(n304),.clk(gclk));
	jor g247(.dina(w_n282_1[0]),.dinb(w_n291_1[0]),.dout(n305),.clk(gclk));
	jor g248(.dina(n305),.dinb(w_n297_0[0]),.dout(n306),.clk(gclk));
	jor g249(.dina(w_n160_0[1]),.dinb(w_n76_0[1]),.dout(n307),.clk(gclk));
	jor g250(.dina(w_n307_0[2]),.dinb(w_n293_0[0]),.dout(n308),.clk(gclk));
	jor g251(.dina(n308),.dinb(w_n282_0[2]),.dout(n309),.clk(gclk));
	jand g252(.dina(n309),.dinb(n306),.dout(n310),.clk(gclk));
	jand g253(.dina(n310),.dinb(w_dff_B_gJdEHobR1_1),.dout(n311),.clk(gclk));
	jand g254(.dina(n311),.dinb(w_dff_B_xxqWYu090_1),.dout(n312),.clk(gclk));
	jand g255(.dina(n312),.dinb(n301),.dout(n313),.clk(gclk));
	jnot g256(.din(w_n192_0[0]),.dout(n314),.clk(gclk));
	jor g257(.dina(w_n110_0[0]),.dinb(w_n95_0[1]),.dout(n315),.clk(gclk));
	jor g258(.dina(n315),.dinb(w_n286_0[0]),.dout(n316),.clk(gclk));
	jnot g259(.din(w_n182_0[1]),.dout(n317),.clk(gclk));
	jor g260(.dina(w_n307_0[1]),.dinb(w_n292_0[0]),.dout(n318),.clk(gclk));
	jor g261(.dina(n318),.dinb(w_n317_0[2]),.dout(n319),.clk(gclk));
	jor g262(.dina(n319),.dinb(w_n316_0[2]),.dout(n320),.clk(gclk));
	jor g263(.dina(w_n153_0[1]),.dinb(w_n168_0[1]),.dout(n321),.clk(gclk));
	jor g264(.dina(w_n317_0[1]),.dinb(n321),.dout(n322),.clk(gclk));
	jor g265(.dina(w_n322_0[1]),.dinb(w_n303_0[0]),.dout(n323),.clk(gclk));
	jor g266(.dina(w_n316_0[1]),.dinb(w_n323_0[1]),.dout(n324),.clk(gclk));
	jand g267(.dina(n324),.dinb(n320),.dout(n325),.clk(gclk));
	jand g268(.dina(n325),.dinb(n314),.dout(n326),.clk(gclk));
	jor g269(.dina(w_n316_0[0]),.dinb(w_n291_0[2]),.dout(n327),.clk(gclk));
	jor g270(.dina(w_n327_0[1]),.dinb(w_n322_0[0]),.dout(n328),.clk(gclk));
	jnot g271(.din(w_n183_0[0]),.dout(n329),.clk(gclk));
	jor g272(.dina(w_n327_0[0]),.dinb(w_n329_0[1]),.dout(n330),.clk(gclk));
	jand g273(.dina(n330),.dinb(n328),.dout(n331),.clk(gclk));
	jor g274(.dina(w_n307_0[0]),.dinb(w_n287_0[2]),.dout(n332),.clk(gclk));
	jor g275(.dina(w_n329_0[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jor g276(.dina(w_n258_0[0]),.dinb(w_n291_0[1]),.dout(n334),.clk(gclk));
	jor g277(.dina(n334),.dinb(w_n317_0[0]),.dout(n335),.clk(gclk));
	jor g278(.dina(n335),.dinb(w_n287_0[1]),.dout(n336),.clk(gclk));
	jor g279(.dina(w_n323_0[0]),.dinb(w_n282_0[1]),.dout(n337),.clk(gclk));
	jand g280(.dina(n337),.dinb(n336),.dout(n338),.clk(gclk));
	jand g281(.dina(n338),.dinb(w_dff_B_JQNBt3Tw0_1),.dout(n339),.clk(gclk));
	jand g282(.dina(n339),.dinb(w_dff_B_slj6ZFIj6_1),.dout(n340),.clk(gclk));
	jand g283(.dina(n340),.dinb(w_dff_B_l8DfnSgd7_1),.dout(n341),.clk(gclk));
	jand g284(.dina(w_n341_0[1]),.dinb(w_n313_0[1]),.dout(n342),.clk(gclk));
	jnot g285(.din(w_n274_0[0]),.dout(n343),.clk(gclk));
	jor g286(.dina(w_dff_B_U4qzGoUC9_0),.dinb(n342),.dout(n344),.clk(gclk));
	jor g287(.dina(n344),.dinb(w_dff_B_XY4RlwRU3_1),.dout(n345),.clk(gclk));
	jand g288(.dina(n345),.dinb(w_n265_1[2]),.dout(n346),.clk(gclk));
	jand g289(.dina(n346),.dinb(w_dff_B_8UVV9BKq0_1),.dout(G60),.clk(gclk));
	jand g290(.dina(w_n242_1[1]),.dinb(w_G478_0[0]),.dout(n348),.clk(gclk));
	jand g291(.dina(n348),.dinb(w_G902_1[2]),.dout(n349),.clk(gclk));
	jxor g292(.dina(n349),.dinb(w_n139_0[0]),.dout(n350),.clk(gclk));
	jand g293(.dina(n350),.dinb(w_n265_1[1]),.dout(G63),.clk(gclk));
	jand g294(.dina(w_n242_1[0]),.dinb(w_G217_0[0]),.dout(n352),.clk(gclk));
	jand g295(.dina(n352),.dinb(w_G902_1[1]),.dout(n353),.clk(gclk));
	jxor g296(.dina(n353),.dinb(w_n70_0[0]),.dout(n354),.clk(gclk));
	jand g297(.dina(n354),.dinb(w_n265_1[0]),.dout(G66),.clk(gclk));
	jor g298(.dina(w_n124_0[0]),.dinb(w_n102_0[0]),.dout(n356),.clk(gclk));
	jor g299(.dina(w_n313_0[0]),.dinb(w_G953_1[0]),.dout(n357),.clk(gclk));
	jand g300(.dina(w_G898_0[0]),.dinb(w_G224_0[0]),.dout(n358),.clk(gclk));
	jor g301(.dina(n358),.dinb(w_n103_1[1]),.dout(n359),.clk(gclk));
	jand g302(.dina(w_dff_B_uSiNie2K1_0),.dinb(n357),.dout(n360),.clk(gclk));
	jxor g303(.dina(n360),.dinb(w_dff_B_8QhtpKir0_1),.dout(w_dff_A_jrsgWhlw6_2),.clk(gclk));
	jor g304(.dina(w_n341_0[0]),.dinb(w_G953_0[2]),.dout(n362),.clk(gclk));
	jand g305(.dina(w_G900_0[0]),.dinb(w_G227_0[0]),.dout(n363),.clk(gclk));
	jor g306(.dina(n363),.dinb(w_n103_1[0]),.dout(n364),.clk(gclk));
	jand g307(.dina(w_dff_B_ai9z8Ib93_0),.dinb(n362),.dout(n365),.clk(gclk));
	jxor g308(.dina(w_n81_0[0]),.dinb(w_n66_0[0]),.dout(n366),.clk(gclk));
	jor g309(.dina(n366),.dinb(w_n180_0[0]),.dout(n367),.clk(gclk));
	jxor g310(.dina(w_dff_B_WGDz4yIs8_0),.dinb(n365),.dout(w_dff_A_bfIBpwvT2_2),.clk(gclk));
	jand g311(.dina(w_G902_1[0]),.dinb(w_G472_0[0]),.dout(n369),.clk(gclk));
	jand g312(.dina(w_dff_B_GVXrhrtJ9_0),.dinb(w_n242_0[2]),.dout(n370),.clk(gclk));
	jxor g313(.dina(n370),.dinb(w_n90_0[0]),.dout(n371),.clk(gclk));
	jand g314(.dina(n371),.dinb(w_n265_0[2]),.dout(w_dff_A_CR8MmAXU9_2),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_dff_A_tkN9220D2_0),.doutb(w_G101_0[1]),.doutc(w_dff_A_of9VE2Fz6_2),.din(G101));
	jspl3 jspl3_w_G104_0(.douta(w_dff_A_FBAHzrOq1_0),.doutb(w_dff_A_eUbbvWIE2_1),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_dff_A_CesXBU2u2_0),.doutb(w_dff_A_6FeGUKFN4_1),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_dff_A_VJyD25BW2_0),.doutb(w_G110_0[1]),.doutc(w_G110_0[2]),.din(G110));
	jspl3 jspl3_w_G113_0(.douta(w_dff_A_NWJHmVeC7_0),.doutb(w_G113_0[1]),.doutc(w_G113_0[2]),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_dff_A_NLyaARlw7_0),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_dff_A_zQr574PS7_0),.doutb(w_G119_0[1]),.doutc(w_dff_A_pnVt8Qtv5_2),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_dff_A_68C1tYLB7_1),.doutc(w_G122_0[2]),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_G122_1[1]),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_dff_A_tFgBrtCK8_0),.doutb(w_dff_A_5e6SVyaf6_1),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_dff_A_7dghcLrw1_0),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(G128));
	jspl3 jspl3_w_G131_0(.douta(w_dff_A_ttSlfJ5X7_0),.doutb(w_G131_0[1]),.doutc(w_dff_A_CzsLeHrX3_2),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_dff_A_7gLeVlQI2_0),.doutb(w_dff_A_XcRayItl7_1),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_NV5cEZc60_0),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G140_0(.douta(w_dff_A_muDEwOhg9_0),.doutb(w_dff_A_ZPd97mhW6_1),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_dff_A_ryEwEkan5_0),.doutb(w_dff_A_dmHWo8dH3_1),.doutc(w_G143_0[2]),.din(G143));
	jspl3 jspl3_w_G146_0(.douta(w_dff_A_DX3jurAJ6_0),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(w_dff_B_QYOxYyQh7_3));
	jspl3 jspl3_w_G210_0(.douta(w_dff_A_VyrqZWlM8_0),.doutb(w_dff_A_2wciar0F4_1),.doutc(w_G210_0[2]),.din(G210));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_dff_A_1s77Wb1L3_1),.din(G214));
	jspl3 jspl3_w_G217_0(.douta(w_dff_A_mYZjQoQo4_0),.doutb(w_G217_0[1]),.doutc(w_dff_A_JcBqaPAX3_2),.din(w_dff_B_M3j6QPic7_3));
	jspl jspl_w_G221_0(.douta(w_dff_A_UmkrL2Bk1_0),.doutb(w_G221_0[1]),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_dff_A_x4CoadrC8_1),.din(G224));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_dff_A_EQkrYTW60_1),.din(G227));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_dff_A_XAwPxIpV3_1),.doutc(w_G234_0[2]),.din(G234));
	jspl jspl_w_G234_1(.douta(w_dff_A_rh5X5q869_0),.doutb(w_G234_1[1]),.din(w_G234_0[0]));
	jspl3 jspl3_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.doutc(w_G237_0[2]),.din(G237));
	jspl3 jspl3_w_G469_0(.douta(w_dff_A_HvlivWmk0_0),.doutb(w_G469_0[1]),.doutc(w_dff_A_ULtBYnlK8_2),.din(G469));
	jspl3 jspl3_w_G472_0(.douta(w_G472_0[0]),.doutb(w_G472_0[1]),.doutc(w_dff_A_6gxqJhLc9_2),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_dff_A_kUu1Mzls8_1),.doutc(w_G475_0[2]),.din(G475));
	jspl3 jspl3_w_G478_0(.douta(w_dff_A_H4EUOxXu5_0),.doutb(w_dff_A_bF80AltB1_1),.doutc(w_G478_0[2]),.din(G478));
	jspl jspl_w_G898_0(.douta(w_G898_0[0]),.doutb(w_dff_A_HRi1yhR67_1),.din(G898));
	jspl jspl_w_G900_0(.douta(w_G900_0[0]),.doutb(w_dff_A_Cpn0gaCa7_1),.din(G900));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_G902_0[2]),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_dff_A_eveR7xjG5_1),.doutc(w_dff_A_9vXg7p2U9_2),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_dff_A_TYWhiCcb1_1),.doutc(w_dff_A_WXr3mAOY7_2),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_dff_A_ekZdutAZ2_0),.doutb(w_G902_3[1]),.doutc(w_G902_3[2]),.din(w_G902_0[2]));
	jspl3 jspl3_w_G952_0(.douta(w_G952_0[0]),.doutb(w_dff_A_fyg1Pvi90_1),.doutc(w_dff_A_9rtk9RnC4_2),.din(w_dff_B_rfC0uYMu3_3));
	jspl3 jspl3_w_G953_0(.douta(w_G953_0[0]),.doutb(w_G953_0[1]),.doutc(w_dff_A_TcigiV841_2),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_dff_A_j20f81iP6_0),.doutb(w_dff_A_6Rsph3Hg4_1),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl jspl_w_G953_2(.douta(w_G953_2[0]),.doutb(w_dff_A_4wyfpWne7_1),.din(w_G953_0[1]));
	jspl3 jspl3_w_n58_0(.douta(w_dff_A_lPlN46Zi2_0),.doutb(w_n58_0[1]),.doutc(w_dff_A_z0LuLn477_2),.din(n58));
	jspl3 jspl3_w_n58_1(.douta(w_n58_1[0]),.doutb(w_n58_1[1]),.doutc(w_n58_1[2]),.din(w_n58_0[0]));
	jspl3 jspl3_w_n58_2(.douta(w_dff_A_IfPdIVTn7_0),.doutb(w_n58_2[1]),.doutc(w_dff_A_H9Rx8CDR8_2),.din(w_n58_0[1]));
	jspl jspl_w_n63_0(.douta(w_n63_0[0]),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n66_0(.douta(w_dff_A_keIiaf2X8_0),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_dff_A_Hri4DIpK9_0),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n70_0(.douta(w_dff_A_12fiUFWN7_0),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n74_0(.douta(w_dff_A_qpoPMpyG5_0),.doutb(w_n74_0[1]),.din(n74));
	jspl3 jspl3_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.doutc(w_n76_0[2]),.din(n76));
	jspl3 jspl3_w_n76_1(.douta(w_n76_1[0]),.doutb(w_n76_1[1]),.doutc(w_n76_1[2]),.din(w_n76_0[0]));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_dff_A_jm8LVCm13_1),.doutc(w_dff_A_wdagkMWX9_2),.din(n81));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_dff_A_ok4oxW2C4_1),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n90_0(.douta(w_dff_A_tU0QD92Y8_0),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.din(n91));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n92_1(.douta(w_n92_1[0]),.doutb(w_n92_1[1]),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_dff_A_UUI63NDL8_1),.doutc(w_dff_A_Zo59uV6y7_2),.din(n93));
	jspl jspl_w_n93_1(.douta(w_n93_1[0]),.doutb(w_dff_A_Goheoi8v6_1),.din(w_n93_0[0]));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n95_0(.douta(w_n95_0[0]),.doutb(w_dff_A_4hau76MP3_1),.doutc(w_dff_A_woUgFLQV7_2),.din(n95));
	jspl jspl_w_n95_1(.douta(w_dff_A_hZVR3lWF6_0),.doutb(w_n95_1[1]),.din(w_n95_0[0]));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_dff_A_4iQ5PsFD0_1),.doutc(w_dff_A_DyND0V2T2_2),.din(w_dff_B_sq9N4pXi0_3));
	jspl jspl_w_n99_0(.douta(w_dff_A_9dENtCRg6_0),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n103_1(.douta(w_n103_1[0]),.doutb(w_n103_1[1]),.doutc(w_n103_1[2]),.din(w_n103_0[0]));
	jspl3 jspl3_w_n103_2(.douta(w_n103_2[0]),.doutb(w_n103_2[1]),.doutc(w_dff_A_kfr5z0gz9_2),.din(w_n103_0[1]));
	jspl3 jspl3_w_n103_3(.douta(w_n103_3[0]),.doutb(w_n103_3[1]),.doutc(w_n103_3[2]),.din(w_n103_0[2]));
	jspl jspl_w_n107_0(.douta(w_dff_A_ASSNhaad5_0),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_dff_A_BPSgy5466_1),.din(n109));
	jspl jspl_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.din(n110));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_dff_A_vI1tui6I2_1),.doutc(w_dff_A_zSeAZakS0_2),.din(n112));
	jspl jspl_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_dff_A_kHyHxSiA5_1),.doutc(w_dff_A_wQPGfbPQ3_2),.din(n113));
	jspl jspl_w_n118_0(.douta(w_dff_A_tqndhuCu4_0),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_dff_A_NAtrOi5y4_1),.doutc(w_n122_0[2]),.din(n122));
	jspl jspl_w_n122_1(.douta(w_n122_1[0]),.doutb(w_n122_1[1]),.din(w_n122_0[0]));
	jspl jspl_w_n124_0(.douta(w_dff_A_raUcn9Zs3_0),.doutb(w_n124_0[1]),.din(n124));
	jspl jspl_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.din(n126));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl3 jspl3_w_n130_0(.douta(w_n130_0[0]),.doutb(w_dff_A_IHjKN1eP7_1),.doutc(w_dff_A_oEm0Nfpx8_2),.din(n130));
	jspl jspl_w_n130_1(.douta(w_n130_1[0]),.doutb(w_n130_1[1]),.din(w_n130_0[0]));
	jspl3 jspl3_w_n131_0(.douta(w_dff_A_M39xwuIo0_0),.doutb(w_n131_0[1]),.doutc(w_dff_A_kdAG6Xfd1_2),.din(n131));
	jspl3 jspl3_w_n131_1(.douta(w_n131_1[0]),.doutb(w_n131_1[1]),.doutc(w_n131_1[2]),.din(w_n131_0[0]));
	jspl jspl_w_n139_0(.douta(w_dff_A_POImPkBN8_0),.doutb(w_n139_0[1]),.din(n139));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n141_1(.douta(w_n141_1[0]),.doutb(w_n141_1[1]),.din(w_n141_0[0]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_oAl19vRy1_1),.doutc(w_n151_0[2]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl jspl_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_dff_A_SWInxcw56_2),.din(n154));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl3 jspl3_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.doutc(w_n160_0[2]),.din(n160));
	jspl3 jspl3_w_n160_1(.douta(w_n160_1[0]),.doutb(w_n160_1[1]),.doutc(w_n160_1[2]),.din(w_n160_0[0]));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_dff_A_bZqGKQsJ5_1),.doutc(w_dff_A_tUN8qgig9_2),.din(w_dff_B_SmSmmBJM7_3));
	jspl jspl_w_n161_1(.douta(w_n161_1[0]),.doutb(w_n161_1[1]),.din(w_n161_0[0]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_n163_0[2]),.din(n163));
	jspl jspl_w_n163_1(.douta(w_n163_1[0]),.doutb(w_n163_1[1]),.din(w_n163_0[0]));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_AE1D2ZU45_1),.doutc(w_dff_A_znOEPE3t7_2),.din(n165));
	jspl jspl_w_n166_0(.douta(w_dff_A_dgHihsKT6_0),.doutb(w_n166_0[1]),.din(n166));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl jspl_w_n168_1(.douta(w_n168_1[0]),.doutb(w_n168_1[1]),.din(w_n168_0[0]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(w_dff_B_L2sw5HXi6_2));
	jspl jspl_w_n171_0(.douta(w_n171_0[0]),.doutb(w_n171_0[1]),.din(n171));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl jspl_w_n173_1(.douta(w_n173_1[0]),.doutb(w_n173_1[1]),.din(w_n173_0[0]));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_dff_A_DTPDCWCH0_1),.din(w_dff_B_vDF4uLgW4_2));
	jspl jspl_w_n175_0(.douta(w_dff_A_WjCKIAiK5_0),.doutb(w_n175_0[1]),.din(n175));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_dff_A_gPnpAazZ3_1),.doutc(w_dff_A_ZwXfHhEL8_2),.din(n177));
	jspl jspl_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.din(n178));
	jspl jspl_w_n180_0(.douta(w_dff_A_Xv4Re0VA8_0),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n182_0(.douta(w_dff_A_EwZWUKIS7_0),.doutb(w_n182_0[1]),.doutc(w_dff_A_eHRBrCIQ1_2),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_dff_A_jElLZGmm8_1),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n183_0(.douta(w_n183_0[0]),.doutb(w_dff_A_szBFXo8J3_1),.doutc(w_dff_A_BsJ2jOKO4_2),.din(n183));
	jspl jspl_w_n184_0(.douta(w_dff_A_1VRB2xs14_0),.doutb(w_n184_0[1]),.din(n184));
	jspl jspl_w_n186_0(.douta(w_dff_A_zbzxFhuo2_0),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n191_0(.douta(w_dff_A_CRco7veP1_0),.doutb(w_n191_0[1]),.doutc(w_dff_A_dKrVgv1U3_2),.din(n191));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_dff_A_ZJtyRA0T1_1),.doutc(w_n192_0[2]),.din(n192));
	jspl3 jspl3_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.doutc(w_n195_0[2]),.din(n195));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_dff_A_ESbhtxXb4_1),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_dff_A_2ypsFFp70_0),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_dff_A_oqBjpYYL8_1),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n208_0(.douta(w_dff_A_6Mu5TVS08_0),.doutb(w_n208_0[1]),.din(n208));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.din(n211));
	jspl3 jspl3_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.doutc(w_n214_0[2]),.din(n214));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.doutc(w_dff_A_zlZRoQlY1_2),.din(n216));
	jspl jspl_w_n216_1(.douta(w_dff_A_qvlnoTIO5_0),.doutb(w_n216_1[1]),.din(w_n216_0[0]));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl3 jspl3_w_n242_1(.douta(w_n242_1[0]),.doutb(w_n242_1[1]),.doutc(w_n242_1[2]),.din(w_n242_0[0]));
	jspl3 jspl3_w_n242_2(.douta(w_n242_2[0]),.doutb(w_n242_2[1]),.doutc(w_n242_2[2]),.din(w_n242_0[1]));
	jspl jspl_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.din(n243));
	jspl jspl_w_n249_0(.douta(w_dff_A_v3ni466f3_0),.doutb(w_n249_0[1]),.din(n249));
	jspl3 jspl3_w_n258_0(.douta(w_n258_0[0]),.doutb(w_dff_A_1yr2Fkib6_1),.doutc(w_dff_A_FPGOcCb08_2),.din(n258));
	jspl3 jspl3_w_n265_0(.douta(w_n265_0[0]),.doutb(w_dff_A_apHLc5GV3_1),.doutc(w_n265_0[2]),.din(w_dff_B_ABthXCsD1_3));
	jspl3 jspl3_w_n265_1(.douta(w_dff_A_fX4U4ovf9_0),.doutb(w_dff_A_cMFoa89n8_1),.doutc(w_n265_1[2]),.din(w_n265_0[0]));
	jspl jspl_w_n265_2(.douta(w_n265_2[0]),.doutb(w_n265_2[1]),.din(w_n265_0[1]));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_gLLZy1pU5_1),.din(n274));
	jspl3 jspl3_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.doutc(w_dff_A_bGwVcjBD4_2),.din(w_dff_B_sb9iZ8bG2_3));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(w_dff_B_K6u4Fd705_2));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n282_0(.douta(w_n282_0[0]),.doutb(w_dff_A_AlG92Tz52_1),.doutc(w_dff_A_WANtlcxU1_2),.din(n282));
	jspl jspl_w_n282_1(.douta(w_n282_1[0]),.doutb(w_n282_1[1]),.din(w_n282_0[0]));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(n286));
	jspl3 jspl3_w_n287_0(.douta(w_n287_0[0]),.doutb(w_dff_A_82Ol37eH4_1),.doutc(w_n287_0[2]),.din(n287));
	jspl jspl_w_n287_1(.douta(w_n287_1[0]),.doutb(w_n287_1[1]),.din(w_n287_0[0]));
	jspl jspl_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.din(n288));
	jspl3 jspl3_w_n291_0(.douta(w_dff_A_3sTCNM3y5_0),.doutb(w_n291_0[1]),.doutc(w_dff_A_aVPtgSo02_2),.din(n291));
	jspl jspl_w_n291_1(.douta(w_n291_1[0]),.doutb(w_dff_A_ABtNJUFx6_1),.din(w_n291_0[0]));
	jspl jspl_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.din(n292));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n294_0(.douta(w_n294_0[0]),.doutb(w_n294_0[1]),.din(n294));
	jspl jspl_w_n297_0(.douta(w_n297_0[0]),.doutb(w_n297_0[1]),.din(w_dff_B_i6qCSWfC6_2));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_lGq66MbF9_1),.din(w_dff_B_hFGawRW00_2));
	jspl3 jspl3_w_n307_0(.douta(w_dff_A_33pc2Raq6_0),.doutb(w_n307_0[1]),.doutc(w_dff_A_wTKLKhEd4_2),.din(n307));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n316_0(.douta(w_n316_0[0]),.doutb(w_dff_A_cCQcj4iH3_1),.doutc(w_dff_A_2sTvlTIs9_2),.din(n316));
	jspl3 jspl3_w_n317_0(.douta(w_dff_A_gmOYxxun3_0),.doutb(w_n317_0[1]),.doutc(w_dff_A_WSLk10X92_2),.din(w_dff_B_6OB8wPMk2_3));
	jspl jspl_w_n322_0(.douta(w_dff_A_Hp3hdCfF5_0),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(n323));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(n327));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n341_0(.douta(w_n341_0[0]),.doutb(w_n341_0[1]),.din(n341));
	jdff dff_B_KUG64qFo9_0(.din(n263),.dout(w_dff_B_KUG64qFo9_0),.clk(gclk));
	jdff dff_B_394Fxekk6_0(.din(w_dff_B_KUG64qFo9_0),.dout(w_dff_B_394Fxekk6_0),.clk(gclk));
	jdff dff_B_alWpnuZ68_0(.din(w_dff_B_394Fxekk6_0),.dout(w_dff_B_alWpnuZ68_0),.clk(gclk));
	jdff dff_B_flIMqsTO9_0(.din(w_dff_B_alWpnuZ68_0),.dout(w_dff_B_flIMqsTO9_0),.clk(gclk));
	jdff dff_B_X1XwYjW90_0(.din(w_dff_B_flIMqsTO9_0),.dout(w_dff_B_X1XwYjW90_0),.clk(gclk));
	jdff dff_B_oCKmzzRJ2_0(.din(n255),.dout(w_dff_B_oCKmzzRJ2_0),.clk(gclk));
	jdff dff_B_HucuwSJG9_0(.din(w_dff_B_oCKmzzRJ2_0),.dout(w_dff_B_HucuwSJG9_0),.clk(gclk));
	jdff dff_B_eggdHZDG6_0(.din(n250),.dout(w_dff_B_eggdHZDG6_0),.clk(gclk));
	jdff dff_A_IG0CL64y6_0(.dout(w_n249_0[0]),.din(w_dff_A_IG0CL64y6_0),.clk(gclk));
	jdff dff_A_v3ni466f3_0(.dout(w_dff_A_IG0CL64y6_0),.din(w_dff_A_v3ni466f3_0),.clk(gclk));
	jdff dff_B_k5gOsM257_0(.din(n248),.dout(w_dff_B_k5gOsM257_0),.clk(gclk));
	jdff dff_B_JBz7l3hc8_0(.din(w_dff_B_k5gOsM257_0),.dout(w_dff_B_JBz7l3hc8_0),.clk(gclk));
	jdff dff_B_hT1JvqQo9_0(.din(n244),.dout(w_dff_B_hT1JvqQo9_0),.clk(gclk));
	jdff dff_B_QTJGx9Zi8_0(.din(w_dff_B_hT1JvqQo9_0),.dout(w_dff_B_QTJGx9Zi8_0),.clk(gclk));
	jdff dff_B_E3zHyqyO6_0(.din(w_dff_B_QTJGx9Zi8_0),.dout(w_dff_B_E3zHyqyO6_0),.clk(gclk));
	jdff dff_B_8UVV9BKq0_1(.din(n276),.dout(w_dff_B_8UVV9BKq0_1),.clk(gclk));
	jdff dff_B_Lvpku14t8_1(.din(n277),.dout(w_dff_B_Lvpku14t8_1),.clk(gclk));
	jdff dff_B_dvRgyTWL3_1(.din(w_dff_B_Lvpku14t8_1),.dout(w_dff_B_dvRgyTWL3_1),.clk(gclk));
	jdff dff_B_f3V5GFWe6_1(.din(w_dff_B_dvRgyTWL3_1),.dout(w_dff_B_f3V5GFWe6_1),.clk(gclk));
	jdff dff_B_w1ZBE5So9_1(.din(w_dff_B_f3V5GFWe6_1),.dout(w_dff_B_w1ZBE5So9_1),.clk(gclk));
	jdff dff_B_D6vUSOhQ9_1(.din(w_dff_B_w1ZBE5So9_1),.dout(w_dff_B_D6vUSOhQ9_1),.clk(gclk));
	jdff dff_B_wo1dfjjy0_1(.din(w_dff_B_D6vUSOhQ9_1),.dout(w_dff_B_wo1dfjjy0_1),.clk(gclk));
	jdff dff_B_HxB01BHw8_1(.din(w_dff_B_wo1dfjjy0_1),.dout(w_dff_B_HxB01BHw8_1),.clk(gclk));
	jdff dff_B_LP0n0gDD2_1(.din(w_dff_B_HxB01BHw8_1),.dout(w_dff_B_LP0n0gDD2_1),.clk(gclk));
	jdff dff_B_j5g1Z4K63_1(.din(w_dff_B_LP0n0gDD2_1),.dout(w_dff_B_j5g1Z4K63_1),.clk(gclk));
	jdff dff_B_nOi7yzSc6_1(.din(w_dff_B_j5g1Z4K63_1),.dout(w_dff_B_nOi7yzSc6_1),.clk(gclk));
	jdff dff_B_XY4RlwRU3_1(.din(w_dff_B_nOi7yzSc6_1),.dout(w_dff_B_XY4RlwRU3_1),.clk(gclk));
	jdff dff_B_oVS34vDx7_0(.din(n343),.dout(w_dff_B_oVS34vDx7_0),.clk(gclk));
	jdff dff_B_s2iS1UZf1_0(.din(w_dff_B_oVS34vDx7_0),.dout(w_dff_B_s2iS1UZf1_0),.clk(gclk));
	jdff dff_B_Km60sTcO5_0(.din(w_dff_B_s2iS1UZf1_0),.dout(w_dff_B_Km60sTcO5_0),.clk(gclk));
	jdff dff_B_7cITet7p8_0(.din(w_dff_B_Km60sTcO5_0),.dout(w_dff_B_7cITet7p8_0),.clk(gclk));
	jdff dff_B_aJLU51O03_0(.din(w_dff_B_7cITet7p8_0),.dout(w_dff_B_aJLU51O03_0),.clk(gclk));
	jdff dff_B_8yblqgjN8_0(.din(w_dff_B_aJLU51O03_0),.dout(w_dff_B_8yblqgjN8_0),.clk(gclk));
	jdff dff_B_GPNNfbOx8_0(.din(w_dff_B_8yblqgjN8_0),.dout(w_dff_B_GPNNfbOx8_0),.clk(gclk));
	jdff dff_B_h0NNqSV74_0(.din(w_dff_B_GPNNfbOx8_0),.dout(w_dff_B_h0NNqSV74_0),.clk(gclk));
	jdff dff_B_FmKeF8Sd9_0(.din(w_dff_B_h0NNqSV74_0),.dout(w_dff_B_FmKeF8Sd9_0),.clk(gclk));
	jdff dff_B_A9yugYQe2_0(.din(w_dff_B_FmKeF8Sd9_0),.dout(w_dff_B_A9yugYQe2_0),.clk(gclk));
	jdff dff_B_CNdE24Io0_0(.din(w_dff_B_A9yugYQe2_0),.dout(w_dff_B_CNdE24Io0_0),.clk(gclk));
	jdff dff_B_9UvZ2llQ9_0(.din(w_dff_B_CNdE24Io0_0),.dout(w_dff_B_9UvZ2llQ9_0),.clk(gclk));
	jdff dff_B_f547bRLo4_0(.din(w_dff_B_9UvZ2llQ9_0),.dout(w_dff_B_f547bRLo4_0),.clk(gclk));
	jdff dff_B_U4qzGoUC9_0(.din(w_dff_B_f547bRLo4_0),.dout(w_dff_B_U4qzGoUC9_0),.clk(gclk));
	jdff dff_A_XxGbtZY94_1(.dout(w_n274_0[1]),.din(w_dff_A_XxGbtZY94_1),.clk(gclk));
	jdff dff_A_I3PxFMEP5_1(.dout(w_dff_A_XxGbtZY94_1),.din(w_dff_A_I3PxFMEP5_1),.clk(gclk));
	jdff dff_A_TGFYP5zS4_1(.dout(w_dff_A_I3PxFMEP5_1),.din(w_dff_A_TGFYP5zS4_1),.clk(gclk));
	jdff dff_A_2ZW7aQZH7_1(.dout(w_dff_A_TGFYP5zS4_1),.din(w_dff_A_2ZW7aQZH7_1),.clk(gclk));
	jdff dff_A_pLuSHK438_1(.dout(w_dff_A_2ZW7aQZH7_1),.din(w_dff_A_pLuSHK438_1),.clk(gclk));
	jdff dff_A_crK3MAGE6_1(.dout(w_dff_A_pLuSHK438_1),.din(w_dff_A_crK3MAGE6_1),.clk(gclk));
	jdff dff_A_QKwrXAwl5_1(.dout(w_dff_A_crK3MAGE6_1),.din(w_dff_A_QKwrXAwl5_1),.clk(gclk));
	jdff dff_A_kmB8DmzN6_1(.dout(w_dff_A_QKwrXAwl5_1),.din(w_dff_A_kmB8DmzN6_1),.clk(gclk));
	jdff dff_A_X7vahN7m6_1(.dout(w_dff_A_kmB8DmzN6_1),.din(w_dff_A_X7vahN7m6_1),.clk(gclk));
	jdff dff_A_aohLhlQ79_1(.dout(w_dff_A_X7vahN7m6_1),.din(w_dff_A_aohLhlQ79_1),.clk(gclk));
	jdff dff_A_RYgo71xN7_1(.dout(w_dff_A_aohLhlQ79_1),.din(w_dff_A_RYgo71xN7_1),.clk(gclk));
	jdff dff_A_DGTpZgc44_1(.dout(w_dff_A_RYgo71xN7_1),.din(w_dff_A_DGTpZgc44_1),.clk(gclk));
	jdff dff_A_k12CDglC2_1(.dout(w_dff_A_DGTpZgc44_1),.din(w_dff_A_k12CDglC2_1),.clk(gclk));
	jdff dff_A_l53IoIuA6_1(.dout(w_dff_A_k12CDglC2_1),.din(w_dff_A_l53IoIuA6_1),.clk(gclk));
	jdff dff_A_gLLZy1pU5_1(.dout(w_dff_A_l53IoIuA6_1),.din(w_dff_A_gLLZy1pU5_1),.clk(gclk));
	jdff dff_A_syXOUwlA2_1(.dout(w_G902_2[1]),.din(w_dff_A_syXOUwlA2_1),.clk(gclk));
	jdff dff_A_vuuSfQjb4_1(.dout(w_dff_A_syXOUwlA2_1),.din(w_dff_A_vuuSfQjb4_1),.clk(gclk));
	jdff dff_A_z7TEBZSF4_1(.dout(w_dff_A_vuuSfQjb4_1),.din(w_dff_A_z7TEBZSF4_1),.clk(gclk));
	jdff dff_A_p3pKopkY3_1(.dout(w_dff_A_z7TEBZSF4_1),.din(w_dff_A_p3pKopkY3_1),.clk(gclk));
	jdff dff_A_FGhfCPHc4_1(.dout(w_dff_A_p3pKopkY3_1),.din(w_dff_A_FGhfCPHc4_1),.clk(gclk));
	jdff dff_A_dp7rQfin0_1(.dout(w_dff_A_FGhfCPHc4_1),.din(w_dff_A_dp7rQfin0_1),.clk(gclk));
	jdff dff_A_pHGEWigZ7_1(.dout(w_dff_A_dp7rQfin0_1),.din(w_dff_A_pHGEWigZ7_1),.clk(gclk));
	jdff dff_A_A9Mpn6Mo7_1(.dout(w_dff_A_pHGEWigZ7_1),.din(w_dff_A_A9Mpn6Mo7_1),.clk(gclk));
	jdff dff_A_vEDHGsRF1_1(.dout(w_dff_A_A9Mpn6Mo7_1),.din(w_dff_A_vEDHGsRF1_1),.clk(gclk));
	jdff dff_A_wke8CEi98_1(.dout(w_dff_A_vEDHGsRF1_1),.din(w_dff_A_wke8CEi98_1),.clk(gclk));
	jdff dff_A_Hi8O8vN88_1(.dout(w_dff_A_wke8CEi98_1),.din(w_dff_A_Hi8O8vN88_1),.clk(gclk));
	jdff dff_A_kt91S0nH0_1(.dout(w_dff_A_Hi8O8vN88_1),.din(w_dff_A_kt91S0nH0_1),.clk(gclk));
	jdff dff_A_mFka8xG79_1(.dout(w_dff_A_kt91S0nH0_1),.din(w_dff_A_mFka8xG79_1),.clk(gclk));
	jdff dff_A_GmsY3EdE6_1(.dout(w_dff_A_mFka8xG79_1),.din(w_dff_A_GmsY3EdE6_1),.clk(gclk));
	jdff dff_A_AXsYIj0G3_1(.dout(w_dff_A_GmsY3EdE6_1),.din(w_dff_A_AXsYIj0G3_1),.clk(gclk));
	jdff dff_A_QVseP5Xn5_1(.dout(w_dff_A_AXsYIj0G3_1),.din(w_dff_A_QVseP5Xn5_1),.clk(gclk));
	jdff dff_A_TYWhiCcb1_1(.dout(w_dff_A_QVseP5Xn5_1),.din(w_dff_A_TYWhiCcb1_1),.clk(gclk));
	jdff dff_A_iGmSLGYQ0_2(.dout(w_G902_2[2]),.din(w_dff_A_iGmSLGYQ0_2),.clk(gclk));
	jdff dff_A_JNDw6oqa7_2(.dout(w_dff_A_iGmSLGYQ0_2),.din(w_dff_A_JNDw6oqa7_2),.clk(gclk));
	jdff dff_A_F7AUvBLO4_2(.dout(w_dff_A_JNDw6oqa7_2),.din(w_dff_A_F7AUvBLO4_2),.clk(gclk));
	jdff dff_A_v3Az2e4l6_2(.dout(w_dff_A_F7AUvBLO4_2),.din(w_dff_A_v3Az2e4l6_2),.clk(gclk));
	jdff dff_A_ShRa6vIr0_2(.dout(w_dff_A_v3Az2e4l6_2),.din(w_dff_A_ShRa6vIr0_2),.clk(gclk));
	jdff dff_A_7ucS4sL53_2(.dout(w_dff_A_ShRa6vIr0_2),.din(w_dff_A_7ucS4sL53_2),.clk(gclk));
	jdff dff_A_YPE5SCWC0_2(.dout(w_dff_A_7ucS4sL53_2),.din(w_dff_A_YPE5SCWC0_2),.clk(gclk));
	jdff dff_A_QzBMqiCV4_2(.dout(w_dff_A_YPE5SCWC0_2),.din(w_dff_A_QzBMqiCV4_2),.clk(gclk));
	jdff dff_A_zOufd4Aa8_2(.dout(w_dff_A_QzBMqiCV4_2),.din(w_dff_A_zOufd4Aa8_2),.clk(gclk));
	jdff dff_A_T2uI2d8G1_2(.dout(w_dff_A_zOufd4Aa8_2),.din(w_dff_A_T2uI2d8G1_2),.clk(gclk));
	jdff dff_A_ayxp7PCQ1_2(.dout(w_dff_A_T2uI2d8G1_2),.din(w_dff_A_ayxp7PCQ1_2),.clk(gclk));
	jdff dff_A_2KVwM7VM7_2(.dout(w_dff_A_ayxp7PCQ1_2),.din(w_dff_A_2KVwM7VM7_2),.clk(gclk));
	jdff dff_A_GnsqHrad7_2(.dout(w_dff_A_2KVwM7VM7_2),.din(w_dff_A_GnsqHrad7_2),.clk(gclk));
	jdff dff_A_ToUJgmBh8_2(.dout(w_dff_A_GnsqHrad7_2),.din(w_dff_A_ToUJgmBh8_2),.clk(gclk));
	jdff dff_A_5YD3cgRK2_2(.dout(w_dff_A_ToUJgmBh8_2),.din(w_dff_A_5YD3cgRK2_2),.clk(gclk));
	jdff dff_A_mDqaywDU7_2(.dout(w_dff_A_5YD3cgRK2_2),.din(w_dff_A_mDqaywDU7_2),.clk(gclk));
	jdff dff_A_WXr3mAOY7_2(.dout(w_dff_A_mDqaywDU7_2),.din(w_dff_A_WXr3mAOY7_2),.clk(gclk));
	jdff dff_A_fX4U4ovf9_0(.dout(w_n265_1[0]),.din(w_dff_A_fX4U4ovf9_0),.clk(gclk));
	jdff dff_A_cMFoa89n8_1(.dout(w_n265_1[1]),.din(w_dff_A_cMFoa89n8_1),.clk(gclk));
	jdff dff_B_hGOzfkvM9_1(.din(n356),.dout(w_dff_B_hGOzfkvM9_1),.clk(gclk));
	jdff dff_B_YURzaCoG9_1(.din(w_dff_B_hGOzfkvM9_1),.dout(w_dff_B_YURzaCoG9_1),.clk(gclk));
	jdff dff_B_5LsUcDqb1_1(.din(w_dff_B_YURzaCoG9_1),.dout(w_dff_B_5LsUcDqb1_1),.clk(gclk));
	jdff dff_B_lWogwtJi2_1(.din(w_dff_B_5LsUcDqb1_1),.dout(w_dff_B_lWogwtJi2_1),.clk(gclk));
	jdff dff_B_8Hz62FqG2_1(.din(w_dff_B_lWogwtJi2_1),.dout(w_dff_B_8Hz62FqG2_1),.clk(gclk));
	jdff dff_B_vFUmr7hp3_1(.din(w_dff_B_8Hz62FqG2_1),.dout(w_dff_B_vFUmr7hp3_1),.clk(gclk));
	jdff dff_B_J5luUa8b5_1(.din(w_dff_B_vFUmr7hp3_1),.dout(w_dff_B_J5luUa8b5_1),.clk(gclk));
	jdff dff_B_drqsJAl31_1(.din(w_dff_B_J5luUa8b5_1),.dout(w_dff_B_drqsJAl31_1),.clk(gclk));
	jdff dff_B_aiC7ouoZ6_1(.din(w_dff_B_drqsJAl31_1),.dout(w_dff_B_aiC7ouoZ6_1),.clk(gclk));
	jdff dff_B_WNGVCYfI7_1(.din(w_dff_B_aiC7ouoZ6_1),.dout(w_dff_B_WNGVCYfI7_1),.clk(gclk));
	jdff dff_B_0XerGWij3_1(.din(w_dff_B_WNGVCYfI7_1),.dout(w_dff_B_0XerGWij3_1),.clk(gclk));
	jdff dff_B_8QhtpKir0_1(.din(w_dff_B_0XerGWij3_1),.dout(w_dff_B_8QhtpKir0_1),.clk(gclk));
	jdff dff_B_UX1OY6Gb2_0(.din(n359),.dout(w_dff_B_UX1OY6Gb2_0),.clk(gclk));
	jdff dff_B_QpE7LmeA5_0(.din(w_dff_B_UX1OY6Gb2_0),.dout(w_dff_B_QpE7LmeA5_0),.clk(gclk));
	jdff dff_B_FbnBAdS51_0(.din(w_dff_B_QpE7LmeA5_0),.dout(w_dff_B_FbnBAdS51_0),.clk(gclk));
	jdff dff_B_w35X5nWO4_0(.din(w_dff_B_FbnBAdS51_0),.dout(w_dff_B_w35X5nWO4_0),.clk(gclk));
	jdff dff_B_w41uq7435_0(.din(w_dff_B_w35X5nWO4_0),.dout(w_dff_B_w41uq7435_0),.clk(gclk));
	jdff dff_B_3mQRfDGC9_0(.din(w_dff_B_w41uq7435_0),.dout(w_dff_B_3mQRfDGC9_0),.clk(gclk));
	jdff dff_B_86QDvtdV9_0(.din(w_dff_B_3mQRfDGC9_0),.dout(w_dff_B_86QDvtdV9_0),.clk(gclk));
	jdff dff_B_HeISs4qd9_0(.din(w_dff_B_86QDvtdV9_0),.dout(w_dff_B_HeISs4qd9_0),.clk(gclk));
	jdff dff_B_YxJ0zRfD3_0(.din(w_dff_B_HeISs4qd9_0),.dout(w_dff_B_YxJ0zRfD3_0),.clk(gclk));
	jdff dff_B_vvhr6LsZ4_0(.din(w_dff_B_YxJ0zRfD3_0),.dout(w_dff_B_vvhr6LsZ4_0),.clk(gclk));
	jdff dff_B_240jvMa60_0(.din(w_dff_B_vvhr6LsZ4_0),.dout(w_dff_B_240jvMa60_0),.clk(gclk));
	jdff dff_B_HAqUgjKD2_0(.din(w_dff_B_240jvMa60_0),.dout(w_dff_B_HAqUgjKD2_0),.clk(gclk));
	jdff dff_B_0o4YFTJ35_0(.din(w_dff_B_HAqUgjKD2_0),.dout(w_dff_B_0o4YFTJ35_0),.clk(gclk));
	jdff dff_B_uSiNie2K1_0(.din(w_dff_B_0o4YFTJ35_0),.dout(w_dff_B_uSiNie2K1_0),.clk(gclk));
	jdff dff_B_xxqWYu090_1(.din(n302),.dout(w_dff_B_xxqWYu090_1),.clk(gclk));
	jdff dff_B_gJdEHobR1_1(.din(n304),.dout(w_dff_B_gJdEHobR1_1),.clk(gclk));
	jdff dff_B_o1k8CBxA6_1(.din(n285),.dout(w_dff_B_o1k8CBxA6_1),.clk(gclk));
	jdff dff_B_BvqV64tH2_1(.din(n290),.dout(w_dff_B_BvqV64tH2_1),.clk(gclk));
	jdff dff_B_i6qCSWfC6_2(.din(n297),.dout(w_dff_B_i6qCSWfC6_2),.clk(gclk));
	jdff dff_A_ABtNJUFx6_1(.dout(w_n291_1[1]),.din(w_dff_A_ABtNJUFx6_1),.clk(gclk));
	jdff dff_B_K6u4Fd705_2(.din(n279),.dout(w_dff_B_K6u4Fd705_2),.clk(gclk));
	jdff dff_A_DoAoh6qP1_2(.dout(w_n278_0[2]),.din(w_dff_A_DoAoh6qP1_2),.clk(gclk));
	jdff dff_A_bGwVcjBD4_2(.dout(w_dff_A_DoAoh6qP1_2),.din(w_dff_A_bGwVcjBD4_2),.clk(gclk));
	jdff dff_B_OqorBsIl3_3(.din(n278),.dout(w_dff_B_OqorBsIl3_3),.clk(gclk));
	jdff dff_B_sb9iZ8bG2_3(.din(w_dff_B_OqorBsIl3_3),.dout(w_dff_B_sb9iZ8bG2_3),.clk(gclk));
	jdff dff_B_VkBUUOFb5_0(.din(n367),.dout(w_dff_B_VkBUUOFb5_0),.clk(gclk));
	jdff dff_B_wIc1UPH12_0(.din(w_dff_B_VkBUUOFb5_0),.dout(w_dff_B_wIc1UPH12_0),.clk(gclk));
	jdff dff_B_VQ2fVj6Q2_0(.din(w_dff_B_wIc1UPH12_0),.dout(w_dff_B_VQ2fVj6Q2_0),.clk(gclk));
	jdff dff_B_z823ZQ8i2_0(.din(w_dff_B_VQ2fVj6Q2_0),.dout(w_dff_B_z823ZQ8i2_0),.clk(gclk));
	jdff dff_B_CKP56xHB2_0(.din(w_dff_B_z823ZQ8i2_0),.dout(w_dff_B_CKP56xHB2_0),.clk(gclk));
	jdff dff_B_Xx7E4TlV7_0(.din(w_dff_B_CKP56xHB2_0),.dout(w_dff_B_Xx7E4TlV7_0),.clk(gclk));
	jdff dff_B_mHbSeaVo7_0(.din(w_dff_B_Xx7E4TlV7_0),.dout(w_dff_B_mHbSeaVo7_0),.clk(gclk));
	jdff dff_B_PygfWZwp8_0(.din(w_dff_B_mHbSeaVo7_0),.dout(w_dff_B_PygfWZwp8_0),.clk(gclk));
	jdff dff_B_eh4kMKeL8_0(.din(w_dff_B_PygfWZwp8_0),.dout(w_dff_B_eh4kMKeL8_0),.clk(gclk));
	jdff dff_B_WZiz5vdx3_0(.din(w_dff_B_eh4kMKeL8_0),.dout(w_dff_B_WZiz5vdx3_0),.clk(gclk));
	jdff dff_B_G6Pc5LI60_0(.din(w_dff_B_WZiz5vdx3_0),.dout(w_dff_B_G6Pc5LI60_0),.clk(gclk));
	jdff dff_B_WGDz4yIs8_0(.din(w_dff_B_G6Pc5LI60_0),.dout(w_dff_B_WGDz4yIs8_0),.clk(gclk));
	jdff dff_B_lXOg0ONp7_0(.din(n364),.dout(w_dff_B_lXOg0ONp7_0),.clk(gclk));
	jdff dff_B_vBaRG9Ml8_0(.din(w_dff_B_lXOg0ONp7_0),.dout(w_dff_B_vBaRG9Ml8_0),.clk(gclk));
	jdff dff_B_C5LRueNP1_0(.din(w_dff_B_vBaRG9Ml8_0),.dout(w_dff_B_C5LRueNP1_0),.clk(gclk));
	jdff dff_B_d6aTAMLa3_0(.din(w_dff_B_C5LRueNP1_0),.dout(w_dff_B_d6aTAMLa3_0),.clk(gclk));
	jdff dff_B_Jho5Yf9L0_0(.din(w_dff_B_d6aTAMLa3_0),.dout(w_dff_B_Jho5Yf9L0_0),.clk(gclk));
	jdff dff_B_jrfgMv3B0_0(.din(w_dff_B_Jho5Yf9L0_0),.dout(w_dff_B_jrfgMv3B0_0),.clk(gclk));
	jdff dff_B_M7QJVnjF3_0(.din(w_dff_B_jrfgMv3B0_0),.dout(w_dff_B_M7QJVnjF3_0),.clk(gclk));
	jdff dff_B_rWpQweSu9_0(.din(w_dff_B_M7QJVnjF3_0),.dout(w_dff_B_rWpQweSu9_0),.clk(gclk));
	jdff dff_B_9a3Fue1j0_0(.din(w_dff_B_rWpQweSu9_0),.dout(w_dff_B_9a3Fue1j0_0),.clk(gclk));
	jdff dff_B_Mklt5Ah61_0(.din(w_dff_B_9a3Fue1j0_0),.dout(w_dff_B_Mklt5Ah61_0),.clk(gclk));
	jdff dff_B_PuUswaoM0_0(.din(w_dff_B_Mklt5Ah61_0),.dout(w_dff_B_PuUswaoM0_0),.clk(gclk));
	jdff dff_B_bHWz2Acr8_0(.din(w_dff_B_PuUswaoM0_0),.dout(w_dff_B_bHWz2Acr8_0),.clk(gclk));
	jdff dff_B_WPzS1h6Y7_0(.din(w_dff_B_bHWz2Acr8_0),.dout(w_dff_B_WPzS1h6Y7_0),.clk(gclk));
	jdff dff_B_ai9z8Ib93_0(.din(w_dff_B_WPzS1h6Y7_0),.dout(w_dff_B_ai9z8Ib93_0),.clk(gclk));
	jdff dff_B_l8DfnSgd7_1(.din(n326),.dout(w_dff_B_l8DfnSgd7_1),.clk(gclk));
	jdff dff_B_slj6ZFIj6_1(.din(n331),.dout(w_dff_B_slj6ZFIj6_1),.clk(gclk));
	jdff dff_B_JQNBt3Tw0_1(.din(n333),.dout(w_dff_B_JQNBt3Tw0_1),.clk(gclk));
	jdff dff_A_AlG92Tz52_1(.dout(w_n282_0[1]),.din(w_dff_A_AlG92Tz52_1),.clk(gclk));
	jdff dff_A_WANtlcxU1_2(.dout(w_n282_0[2]),.din(w_dff_A_WANtlcxU1_2),.clk(gclk));
	jdff dff_A_nJmoAc6P5_1(.dout(w_n258_0[1]),.din(w_dff_A_nJmoAc6P5_1),.clk(gclk));
	jdff dff_A_Mfurm3pw8_1(.dout(w_dff_A_nJmoAc6P5_1),.din(w_dff_A_Mfurm3pw8_1),.clk(gclk));
	jdff dff_A_1yr2Fkib6_1(.dout(w_dff_A_Mfurm3pw8_1),.din(w_dff_A_1yr2Fkib6_1),.clk(gclk));
	jdff dff_A_FPGOcCb08_2(.dout(w_n258_0[2]),.din(w_dff_A_FPGOcCb08_2),.clk(gclk));
	jdff dff_A_82Ol37eH4_1(.dout(w_n287_0[1]),.din(w_dff_A_82Ol37eH4_1),.clk(gclk));
	jdff dff_A_3sTCNM3y5_0(.dout(w_n291_0[0]),.din(w_dff_A_3sTCNM3y5_0),.clk(gclk));
	jdff dff_A_aVPtgSo02_2(.dout(w_n291_0[2]),.din(w_dff_A_aVPtgSo02_2),.clk(gclk));
	jdff dff_A_Hp3hdCfF5_0(.dout(w_n322_0[0]),.din(w_dff_A_Hp3hdCfF5_0),.clk(gclk));
	jdff dff_A_lGq66MbF9_1(.dout(w_n303_0[1]),.din(w_dff_A_lGq66MbF9_1),.clk(gclk));
	jdff dff_B_hFGawRW00_2(.din(n303),.dout(w_dff_B_hFGawRW00_2),.clk(gclk));
	jdff dff_A_33pc2Raq6_0(.dout(w_n307_0[0]),.din(w_dff_A_33pc2Raq6_0),.clk(gclk));
	jdff dff_A_wTKLKhEd4_2(.dout(w_n307_0[2]),.din(w_dff_A_wTKLKhEd4_2),.clk(gclk));
	jdff dff_A_gmOYxxun3_0(.dout(w_n317_0[0]),.din(w_dff_A_gmOYxxun3_0),.clk(gclk));
	jdff dff_A_WSLk10X92_2(.dout(w_n317_0[2]),.din(w_dff_A_WSLk10X92_2),.clk(gclk));
	jdff dff_B_YpyyUZvx8_3(.din(n317),.dout(w_dff_B_YpyyUZvx8_3),.clk(gclk));
	jdff dff_B_6OB8wPMk2_3(.din(w_dff_B_YpyyUZvx8_3),.dout(w_dff_B_6OB8wPMk2_3),.clk(gclk));
	jdff dff_A_cCQcj4iH3_1(.dout(w_n316_0[1]),.din(w_dff_A_cCQcj4iH3_1),.clk(gclk));
	jdff dff_A_2sTvlTIs9_2(.dout(w_n316_0[2]),.din(w_dff_A_2sTvlTIs9_2),.clk(gclk));
	jdff dff_B_9j5Z6XY35_0(.din(n369),.dout(w_dff_B_9j5Z6XY35_0),.clk(gclk));
	jdff dff_B_To039hLW4_0(.din(w_dff_B_9j5Z6XY35_0),.dout(w_dff_B_To039hLW4_0),.clk(gclk));
	jdff dff_B_qS0RVbv06_0(.din(w_dff_B_To039hLW4_0),.dout(w_dff_B_qS0RVbv06_0),.clk(gclk));
	jdff dff_B_QMmS2fVF6_0(.din(w_dff_B_qS0RVbv06_0),.dout(w_dff_B_QMmS2fVF6_0),.clk(gclk));
	jdff dff_B_XWojwD808_0(.din(w_dff_B_QMmS2fVF6_0),.dout(w_dff_B_XWojwD808_0),.clk(gclk));
	jdff dff_B_wRxdAre98_0(.din(w_dff_B_XWojwD808_0),.dout(w_dff_B_wRxdAre98_0),.clk(gclk));
	jdff dff_B_1bIDSDbp4_0(.din(w_dff_B_wRxdAre98_0),.dout(w_dff_B_1bIDSDbp4_0),.clk(gclk));
	jdff dff_B_z32MSyet2_0(.din(w_dff_B_1bIDSDbp4_0),.dout(w_dff_B_z32MSyet2_0),.clk(gclk));
	jdff dff_B_toAuobQO5_0(.din(w_dff_B_z32MSyet2_0),.dout(w_dff_B_toAuobQO5_0),.clk(gclk));
	jdff dff_B_nTDLVa0Y5_0(.din(w_dff_B_toAuobQO5_0),.dout(w_dff_B_nTDLVa0Y5_0),.clk(gclk));
	jdff dff_B_C2Wt8arC7_0(.din(w_dff_B_nTDLVa0Y5_0),.dout(w_dff_B_C2Wt8arC7_0),.clk(gclk));
	jdff dff_B_jPLi9S8P9_0(.din(w_dff_B_C2Wt8arC7_0),.dout(w_dff_B_jPLi9S8P9_0),.clk(gclk));
	jdff dff_B_jzpWERoA1_0(.din(w_dff_B_jPLi9S8P9_0),.dout(w_dff_B_jzpWERoA1_0),.clk(gclk));
	jdff dff_B_o3xNFRU61_0(.din(w_dff_B_jzpWERoA1_0),.dout(w_dff_B_o3xNFRU61_0),.clk(gclk));
	jdff dff_B_GVXrhrtJ9_0(.din(w_dff_B_o3xNFRU61_0),.dout(w_dff_B_GVXrhrtJ9_0),.clk(gclk));
	jdff dff_A_cxbLVBeD5_1(.dout(w_G902_1[1]),.din(w_dff_A_cxbLVBeD5_1),.clk(gclk));
	jdff dff_A_HVcZbEPt6_1(.dout(w_dff_A_cxbLVBeD5_1),.din(w_dff_A_HVcZbEPt6_1),.clk(gclk));
	jdff dff_A_uD3aOx0V1_1(.dout(w_dff_A_HVcZbEPt6_1),.din(w_dff_A_uD3aOx0V1_1),.clk(gclk));
	jdff dff_A_mOpspPGk4_1(.dout(w_dff_A_uD3aOx0V1_1),.din(w_dff_A_mOpspPGk4_1),.clk(gclk));
	jdff dff_A_WqcpWQGw2_1(.dout(w_dff_A_mOpspPGk4_1),.din(w_dff_A_WqcpWQGw2_1),.clk(gclk));
	jdff dff_A_10g0eqLL5_1(.dout(w_dff_A_WqcpWQGw2_1),.din(w_dff_A_10g0eqLL5_1),.clk(gclk));
	jdff dff_A_mNwDuFKi5_1(.dout(w_dff_A_10g0eqLL5_1),.din(w_dff_A_mNwDuFKi5_1),.clk(gclk));
	jdff dff_A_6qXO61xc4_1(.dout(w_dff_A_mNwDuFKi5_1),.din(w_dff_A_6qXO61xc4_1),.clk(gclk));
	jdff dff_A_fpPIGJVJ4_1(.dout(w_dff_A_6qXO61xc4_1),.din(w_dff_A_fpPIGJVJ4_1),.clk(gclk));
	jdff dff_A_ntxM5n5S8_1(.dout(w_dff_A_fpPIGJVJ4_1),.din(w_dff_A_ntxM5n5S8_1),.clk(gclk));
	jdff dff_A_6kRSMX3n4_1(.dout(w_dff_A_ntxM5n5S8_1),.din(w_dff_A_6kRSMX3n4_1),.clk(gclk));
	jdff dff_A_GShpcJh22_1(.dout(w_dff_A_6kRSMX3n4_1),.din(w_dff_A_GShpcJh22_1),.clk(gclk));
	jdff dff_A_NJQ70hQm1_1(.dout(w_dff_A_GShpcJh22_1),.din(w_dff_A_NJQ70hQm1_1),.clk(gclk));
	jdff dff_A_OgvA04eG7_1(.dout(w_dff_A_NJQ70hQm1_1),.din(w_dff_A_OgvA04eG7_1),.clk(gclk));
	jdff dff_A_pQFwUsRx7_1(.dout(w_dff_A_OgvA04eG7_1),.din(w_dff_A_pQFwUsRx7_1),.clk(gclk));
	jdff dff_A_9JcezBKN5_1(.dout(w_dff_A_pQFwUsRx7_1),.din(w_dff_A_9JcezBKN5_1),.clk(gclk));
	jdff dff_A_eveR7xjG5_1(.dout(w_dff_A_9JcezBKN5_1),.din(w_dff_A_eveR7xjG5_1),.clk(gclk));
	jdff dff_A_R0P7A7Oe4_2(.dout(w_G902_1[2]),.din(w_dff_A_R0P7A7Oe4_2),.clk(gclk));
	jdff dff_A_doPstua32_2(.dout(w_dff_A_R0P7A7Oe4_2),.din(w_dff_A_doPstua32_2),.clk(gclk));
	jdff dff_A_IaklNWCl1_2(.dout(w_dff_A_doPstua32_2),.din(w_dff_A_IaklNWCl1_2),.clk(gclk));
	jdff dff_A_vl8SOYU20_2(.dout(w_dff_A_IaklNWCl1_2),.din(w_dff_A_vl8SOYU20_2),.clk(gclk));
	jdff dff_A_OOXBT9eP7_2(.dout(w_dff_A_vl8SOYU20_2),.din(w_dff_A_OOXBT9eP7_2),.clk(gclk));
	jdff dff_A_LSOiE9oF1_2(.dout(w_dff_A_OOXBT9eP7_2),.din(w_dff_A_LSOiE9oF1_2),.clk(gclk));
	jdff dff_A_0UcrAbvE0_2(.dout(w_dff_A_LSOiE9oF1_2),.din(w_dff_A_0UcrAbvE0_2),.clk(gclk));
	jdff dff_A_ULUrvKIz6_2(.dout(w_dff_A_0UcrAbvE0_2),.din(w_dff_A_ULUrvKIz6_2),.clk(gclk));
	jdff dff_A_XUxngNkg4_2(.dout(w_dff_A_ULUrvKIz6_2),.din(w_dff_A_XUxngNkg4_2),.clk(gclk));
	jdff dff_A_Sj6X3e9V5_2(.dout(w_dff_A_XUxngNkg4_2),.din(w_dff_A_Sj6X3e9V5_2),.clk(gclk));
	jdff dff_A_Xg6o16VL7_2(.dout(w_dff_A_Sj6X3e9V5_2),.din(w_dff_A_Xg6o16VL7_2),.clk(gclk));
	jdff dff_A_YDDeoh0r5_2(.dout(w_dff_A_Xg6o16VL7_2),.din(w_dff_A_YDDeoh0r5_2),.clk(gclk));
	jdff dff_A_VtmdS7t47_2(.dout(w_dff_A_YDDeoh0r5_2),.din(w_dff_A_VtmdS7t47_2),.clk(gclk));
	jdff dff_A_fIZEEFDX0_2(.dout(w_dff_A_VtmdS7t47_2),.din(w_dff_A_fIZEEFDX0_2),.clk(gclk));
	jdff dff_A_SkIp3MHM6_2(.dout(w_dff_A_fIZEEFDX0_2),.din(w_dff_A_SkIp3MHM6_2),.clk(gclk));
	jdff dff_A_C32Ed3NP0_2(.dout(w_dff_A_SkIp3MHM6_2),.din(w_dff_A_C32Ed3NP0_2),.clk(gclk));
	jdff dff_A_9vXg7p2U9_2(.dout(w_dff_A_C32Ed3NP0_2),.din(w_dff_A_9vXg7p2U9_2),.clk(gclk));
	jdff dff_B_RqHLDa1b8_1(.din(n236),.dout(w_dff_B_RqHLDa1b8_1),.clk(gclk));
	jdff dff_B_JC95DaZ65_1(.din(n237),.dout(w_dff_B_JC95DaZ65_1),.clk(gclk));
	jdff dff_A_1VRB2xs14_0(.dout(w_n184_0[0]),.din(w_dff_A_1VRB2xs14_0),.clk(gclk));
	jdff dff_A_szBFXo8J3_1(.dout(w_n183_0[1]),.din(w_dff_A_szBFXo8J3_1),.clk(gclk));
	jdff dff_A_BsJ2jOKO4_2(.dout(w_n183_0[2]),.din(w_dff_A_BsJ2jOKO4_2),.clk(gclk));
	jdff dff_A_qvlnoTIO5_0(.dout(w_n216_1[0]),.din(w_dff_A_qvlnoTIO5_0),.clk(gclk));
	jdff dff_A_zlZRoQlY1_2(.dout(w_n216_0[2]),.din(w_dff_A_zlZRoQlY1_2),.clk(gclk));
	jdff dff_B_PzhPMEus9_0(.din(n213),.dout(w_dff_B_PzhPMEus9_0),.clk(gclk));
	jdff dff_B_dkcwcKti5_0(.din(w_dff_B_PzhPMEus9_0),.dout(w_dff_B_dkcwcKti5_0),.clk(gclk));
	jdff dff_B_2muhCsUb1_0(.din(w_dff_B_dkcwcKti5_0),.dout(w_dff_B_2muhCsUb1_0),.clk(gclk));
	jdff dff_A_ZJtyRA0T1_1(.dout(w_n192_0[1]),.din(w_dff_A_ZJtyRA0T1_1),.clk(gclk));
	jdff dff_A_CRco7veP1_0(.dout(w_n191_0[0]),.din(w_dff_A_CRco7veP1_0),.clk(gclk));
	jdff dff_A_dKrVgv1U3_2(.dout(w_n191_0[2]),.din(w_dff_A_dKrVgv1U3_2),.clk(gclk));
	jdff dff_A_jElLZGmm8_1(.dout(w_n182_1[1]),.din(w_dff_A_jElLZGmm8_1),.clk(gclk));
	jdff dff_A_3CCsnjzW2_0(.dout(w_n182_0[0]),.din(w_dff_A_3CCsnjzW2_0),.clk(gclk));
	jdff dff_A_19G8xX9t3_0(.dout(w_dff_A_3CCsnjzW2_0),.din(w_dff_A_19G8xX9t3_0),.clk(gclk));
	jdff dff_A_EwZWUKIS7_0(.dout(w_dff_A_19G8xX9t3_0),.din(w_dff_A_EwZWUKIS7_0),.clk(gclk));
	jdff dff_A_pmbcomq20_2(.dout(w_n182_0[2]),.din(w_dff_A_pmbcomq20_2),.clk(gclk));
	jdff dff_A_9S237OTl6_2(.dout(w_dff_A_pmbcomq20_2),.din(w_dff_A_9S237OTl6_2),.clk(gclk));
	jdff dff_A_8pmT6EMg5_2(.dout(w_dff_A_9S237OTl6_2),.din(w_dff_A_8pmT6EMg5_2),.clk(gclk));
	jdff dff_A_eHRBrCIQ1_2(.dout(w_dff_A_8pmT6EMg5_2),.din(w_dff_A_eHRBrCIQ1_2),.clk(gclk));
	jdff dff_A_Xv4Re0VA8_0(.dout(w_n180_0[0]),.din(w_dff_A_Xv4Re0VA8_0),.clk(gclk));
	jdff dff_A_Cpn0gaCa7_1(.dout(w_G900_0[1]),.din(w_dff_A_Cpn0gaCa7_1),.clk(gclk));
	jdff dff_A_gPnpAazZ3_1(.dout(w_n177_0[1]),.din(w_dff_A_gPnpAazZ3_1),.clk(gclk));
	jdff dff_A_ZwXfHhEL8_2(.dout(w_n177_0[2]),.din(w_dff_A_ZwXfHhEL8_2),.clk(gclk));
	jdff dff_A_WjCKIAiK5_0(.dout(w_n175_0[0]),.din(w_dff_A_WjCKIAiK5_0),.clk(gclk));
	jdff dff_A_DTPDCWCH0_1(.dout(w_n174_0[1]),.din(w_dff_A_DTPDCWCH0_1),.clk(gclk));
	jdff dff_B_vDF4uLgW4_2(.din(n174),.dout(w_dff_B_vDF4uLgW4_2),.clk(gclk));
	jdff dff_A_yPVhSkGV2_1(.dout(w_n199_0[1]),.din(w_dff_A_yPVhSkGV2_1),.clk(gclk));
	jdff dff_A_oqBjpYYL8_1(.dout(w_dff_A_yPVhSkGV2_1),.din(w_dff_A_oqBjpYYL8_1),.clk(gclk));
	jdff dff_A_2ypsFFp70_0(.dout(w_n197_1[0]),.din(w_dff_A_2ypsFFp70_0),.clk(gclk));
	jdff dff_B_L2sw5HXi6_2(.din(n170),.dout(w_dff_B_L2sw5HXi6_2),.clk(gclk));
	jdff dff_A_REp22pjD7_2(.dout(w_n154_0[2]),.din(w_dff_A_REp22pjD7_2),.clk(gclk));
	jdff dff_A_zT089Ygc2_2(.dout(w_dff_A_REp22pjD7_2),.din(w_dff_A_zT089Ygc2_2),.clk(gclk));
	jdff dff_A_3b8lsqOb6_2(.dout(w_dff_A_zT089Ygc2_2),.din(w_dff_A_3b8lsqOb6_2),.clk(gclk));
	jdff dff_A_SWInxcw56_2(.dout(w_dff_A_3b8lsqOb6_2),.din(w_dff_A_SWInxcw56_2),.clk(gclk));
	jdff dff_B_MRaEe7G13_1(.din(n142),.dout(w_dff_B_MRaEe7G13_1),.clk(gclk));
	jdff dff_B_2bzhOtmf4_1(.din(w_dff_B_MRaEe7G13_1),.dout(w_dff_B_2bzhOtmf4_1),.clk(gclk));
	jdff dff_B_OZ6XhuiB2_1(.din(w_dff_B_2bzhOtmf4_1),.dout(w_dff_B_OZ6XhuiB2_1),.clk(gclk));
	jdff dff_B_S3yyGRCa6_1(.din(w_dff_B_OZ6XhuiB2_1),.dout(w_dff_B_S3yyGRCa6_1),.clk(gclk));
	jdff dff_B_4GcJj6UK9_1(.din(w_dff_B_S3yyGRCa6_1),.dout(w_dff_B_4GcJj6UK9_1),.clk(gclk));
	jdff dff_A_jeviynMh1_1(.dout(w_n93_1[1]),.din(w_dff_A_jeviynMh1_1),.clk(gclk));
	jdff dff_A_Goheoi8v6_1(.dout(w_dff_A_jeviynMh1_1),.din(w_dff_A_Goheoi8v6_1),.clk(gclk));
	jdff dff_A_UUI63NDL8_1(.dout(w_n93_0[1]),.din(w_dff_A_UUI63NDL8_1),.clk(gclk));
	jdff dff_A_Zo59uV6y7_2(.dout(w_n93_0[2]),.din(w_dff_A_Zo59uV6y7_2),.clk(gclk));
	jdff dff_A_dgHihsKT6_0(.dout(w_n166_0[0]),.din(w_dff_A_dgHihsKT6_0),.clk(gclk));
	jdff dff_A_AE1D2ZU45_1(.dout(w_n165_0[1]),.din(w_dff_A_AE1D2ZU45_1),.clk(gclk));
	jdff dff_A_znOEPE3t7_2(.dout(w_n165_0[2]),.din(w_dff_A_znOEPE3t7_2),.clk(gclk));
	jdff dff_B_5nsrbSC05_1(.din(n132),.dout(w_dff_B_5nsrbSC05_1),.clk(gclk));
	jdff dff_B_OPIO8SGq4_1(.din(w_dff_B_5nsrbSC05_1),.dout(w_dff_B_OPIO8SGq4_1),.clk(gclk));
	jdff dff_B_UnXNkBs69_1(.din(w_dff_B_OPIO8SGq4_1),.dout(w_dff_B_UnXNkBs69_1),.clk(gclk));
	jdff dff_B_pkG8ZWhz3_1(.din(w_dff_B_UnXNkBs69_1),.dout(w_dff_B_pkG8ZWhz3_1),.clk(gclk));
	jdff dff_B_kbcpQt2j9_1(.din(w_dff_B_pkG8ZWhz3_1),.dout(w_dff_B_kbcpQt2j9_1),.clk(gclk));
	jdff dff_A_NAtrOi5y4_1(.dout(w_n122_0[1]),.din(w_dff_A_NAtrOi5y4_1),.clk(gclk));
	jdff dff_A_6Mu5TVS08_0(.dout(w_n208_0[0]),.din(w_dff_A_6Mu5TVS08_0),.clk(gclk));
	jdff dff_A_ESbhtxXb4_1(.dout(w_n197_0[1]),.din(w_dff_A_ESbhtxXb4_1),.clk(gclk));
	jdff dff_B_k6APoGJQ8_1(.din(n194),.dout(w_dff_B_k6APoGJQ8_1),.clk(gclk));
	jdff dff_B_DS7aIEQu2_1(.din(w_dff_B_k6APoGJQ8_1),.dout(w_dff_B_DS7aIEQu2_1),.clk(gclk));
	jdff dff_B_h9cOKgaC6_1(.din(w_dff_B_DS7aIEQu2_1),.dout(w_dff_B_h9cOKgaC6_1),.clk(gclk));
	jdff dff_B_xn4tmahP4_1(.din(w_dff_B_h9cOKgaC6_1),.dout(w_dff_B_xn4tmahP4_1),.clk(gclk));
	jdff dff_B_NsDCSFXi4_1(.din(w_dff_B_xn4tmahP4_1),.dout(w_dff_B_NsDCSFXi4_1),.clk(gclk));
	jdff dff_A_zDABCEQv4_0(.dout(w_n118_0[0]),.din(w_dff_A_zDABCEQv4_0),.clk(gclk));
	jdff dff_A_IwDaN4mS1_0(.dout(w_dff_A_zDABCEQv4_0),.din(w_dff_A_IwDaN4mS1_0),.clk(gclk));
	jdff dff_A_Ep1bIAFe4_0(.dout(w_dff_A_IwDaN4mS1_0),.din(w_dff_A_Ep1bIAFe4_0),.clk(gclk));
	jdff dff_A_nmWGtdch3_0(.dout(w_dff_A_Ep1bIAFe4_0),.din(w_dff_A_nmWGtdch3_0),.clk(gclk));
	jdff dff_A_B7fuyqWW3_0(.dout(w_dff_A_nmWGtdch3_0),.din(w_dff_A_B7fuyqWW3_0),.clk(gclk));
	jdff dff_A_nUzh37dZ2_0(.dout(w_dff_A_B7fuyqWW3_0),.din(w_dff_A_nUzh37dZ2_0),.clk(gclk));
	jdff dff_A_EJl3uVnT3_0(.dout(w_dff_A_nUzh37dZ2_0),.din(w_dff_A_EJl3uVnT3_0),.clk(gclk));
	jdff dff_A_DyOqZUPQ7_0(.dout(w_dff_A_EJl3uVnT3_0),.din(w_dff_A_DyOqZUPQ7_0),.clk(gclk));
	jdff dff_A_4kAObYLq2_0(.dout(w_dff_A_DyOqZUPQ7_0),.din(w_dff_A_4kAObYLq2_0),.clk(gclk));
	jdff dff_A_1ggNEJ7t1_0(.dout(w_dff_A_4kAObYLq2_0),.din(w_dff_A_1ggNEJ7t1_0),.clk(gclk));
	jdff dff_A_U73lyVPM5_0(.dout(w_dff_A_1ggNEJ7t1_0),.din(w_dff_A_U73lyVPM5_0),.clk(gclk));
	jdff dff_A_tQh4oj1H7_0(.dout(w_dff_A_U73lyVPM5_0),.din(w_dff_A_tQh4oj1H7_0),.clk(gclk));
	jdff dff_A_tqndhuCu4_0(.dout(w_dff_A_tQh4oj1H7_0),.din(w_dff_A_tqndhuCu4_0),.clk(gclk));
	jdff dff_A_EQkrYTW60_1(.dout(w_G227_0[1]),.din(w_dff_A_EQkrYTW60_1),.clk(gclk));
	jdff dff_A_Nep6uVWh4_0(.dout(w_G469_0[0]),.din(w_dff_A_Nep6uVWh4_0),.clk(gclk));
	jdff dff_A_i7U0X4g38_0(.dout(w_dff_A_Nep6uVWh4_0),.din(w_dff_A_i7U0X4g38_0),.clk(gclk));
	jdff dff_A_N29Ib9Xp6_0(.dout(w_dff_A_i7U0X4g38_0),.din(w_dff_A_N29Ib9Xp6_0),.clk(gclk));
	jdff dff_A_iatluKOH0_0(.dout(w_dff_A_N29Ib9Xp6_0),.din(w_dff_A_iatluKOH0_0),.clk(gclk));
	jdff dff_A_nxfbMlCP2_0(.dout(w_dff_A_iatluKOH0_0),.din(w_dff_A_nxfbMlCP2_0),.clk(gclk));
	jdff dff_A_oDForQPh5_0(.dout(w_dff_A_nxfbMlCP2_0),.din(w_dff_A_oDForQPh5_0),.clk(gclk));
	jdff dff_A_Z6J848JK0_0(.dout(w_dff_A_oDForQPh5_0),.din(w_dff_A_Z6J848JK0_0),.clk(gclk));
	jdff dff_A_fpR1vrs22_0(.dout(w_dff_A_Z6J848JK0_0),.din(w_dff_A_fpR1vrs22_0),.clk(gclk));
	jdff dff_A_jIcyLV9S1_0(.dout(w_dff_A_fpR1vrs22_0),.din(w_dff_A_jIcyLV9S1_0),.clk(gclk));
	jdff dff_A_BDCUAhlO5_0(.dout(w_dff_A_jIcyLV9S1_0),.din(w_dff_A_BDCUAhlO5_0),.clk(gclk));
	jdff dff_A_IP1JPemf0_0(.dout(w_dff_A_BDCUAhlO5_0),.din(w_dff_A_IP1JPemf0_0),.clk(gclk));
	jdff dff_A_kDqQp4wh2_0(.dout(w_dff_A_IP1JPemf0_0),.din(w_dff_A_kDqQp4wh2_0),.clk(gclk));
	jdff dff_A_zoEEl4xc9_0(.dout(w_dff_A_kDqQp4wh2_0),.din(w_dff_A_zoEEl4xc9_0),.clk(gclk));
	jdff dff_A_MMQqbunt0_0(.dout(w_dff_A_zoEEl4xc9_0),.din(w_dff_A_MMQqbunt0_0),.clk(gclk));
	jdff dff_A_NUweUMAO7_0(.dout(w_dff_A_MMQqbunt0_0),.din(w_dff_A_NUweUMAO7_0),.clk(gclk));
	jdff dff_A_HvlivWmk0_0(.dout(w_dff_A_NUweUMAO7_0),.din(w_dff_A_HvlivWmk0_0),.clk(gclk));
	jdff dff_A_r5oBXoY02_2(.dout(w_G469_0[2]),.din(w_dff_A_r5oBXoY02_2),.clk(gclk));
	jdff dff_A_Fe6t2XlX6_2(.dout(w_dff_A_r5oBXoY02_2),.din(w_dff_A_Fe6t2XlX6_2),.clk(gclk));
	jdff dff_A_wWIJ0g4Y4_2(.dout(w_dff_A_Fe6t2XlX6_2),.din(w_dff_A_wWIJ0g4Y4_2),.clk(gclk));
	jdff dff_A_YmUIaqRu3_2(.dout(w_dff_A_wWIJ0g4Y4_2),.din(w_dff_A_YmUIaqRu3_2),.clk(gclk));
	jdff dff_A_hDwbYA1M4_2(.dout(w_dff_A_YmUIaqRu3_2),.din(w_dff_A_hDwbYA1M4_2),.clk(gclk));
	jdff dff_A_ULtBYnlK8_2(.dout(w_dff_A_hDwbYA1M4_2),.din(w_dff_A_ULtBYnlK8_2),.clk(gclk));
	jdff dff_A_sjWVkpVN1_1(.dout(w_n113_0[1]),.din(w_dff_A_sjWVkpVN1_1),.clk(gclk));
	jdff dff_A_kHyHxSiA5_1(.dout(w_dff_A_sjWVkpVN1_1),.din(w_dff_A_kHyHxSiA5_1),.clk(gclk));
	jdff dff_A_HtiQBFxH9_2(.dout(w_n113_0[2]),.din(w_dff_A_HtiQBFxH9_2),.clk(gclk));
	jdff dff_A_wQPGfbPQ3_2(.dout(w_dff_A_HtiQBFxH9_2),.din(w_dff_A_wQPGfbPQ3_2),.clk(gclk));
	jdff dff_A_OU8Ehhts9_1(.dout(w_n112_0[1]),.din(w_dff_A_OU8Ehhts9_1),.clk(gclk));
	jdff dff_A_aYi1miGV4_1(.dout(w_dff_A_OU8Ehhts9_1),.din(w_dff_A_aYi1miGV4_1),.clk(gclk));
	jdff dff_A_vI1tui6I2_1(.dout(w_dff_A_aYi1miGV4_1),.din(w_dff_A_vI1tui6I2_1),.clk(gclk));
	jdff dff_A_tjuDygRx7_2(.dout(w_n112_0[2]),.din(w_dff_A_tjuDygRx7_2),.clk(gclk));
	jdff dff_A_Pe5pLhwT1_2(.dout(w_dff_A_tjuDygRx7_2),.din(w_dff_A_Pe5pLhwT1_2),.clk(gclk));
	jdff dff_A_zSeAZakS0_2(.dout(w_dff_A_Pe5pLhwT1_2),.din(w_dff_A_zSeAZakS0_2),.clk(gclk));
	jdff dff_A_FLf3qhb67_1(.dout(w_n109_0[1]),.din(w_dff_A_FLf3qhb67_1),.clk(gclk));
	jdff dff_A_XnCSF2Rn3_1(.dout(w_dff_A_FLf3qhb67_1),.din(w_dff_A_XnCSF2Rn3_1),.clk(gclk));
	jdff dff_A_9E2EhCul1_1(.dout(w_dff_A_XnCSF2Rn3_1),.din(w_dff_A_9E2EhCul1_1),.clk(gclk));
	jdff dff_A_BPSgy5466_1(.dout(w_dff_A_9E2EhCul1_1),.din(w_dff_A_BPSgy5466_1),.clk(gclk));
	jdff dff_A_LYnqv5er8_0(.dout(w_n107_0[0]),.din(w_dff_A_LYnqv5er8_0),.clk(gclk));
	jdff dff_A_D7vO2Dl39_0(.dout(w_dff_A_LYnqv5er8_0),.din(w_dff_A_D7vO2Dl39_0),.clk(gclk));
	jdff dff_A_v0qq9xQJ7_0(.dout(w_dff_A_D7vO2Dl39_0),.din(w_dff_A_v0qq9xQJ7_0),.clk(gclk));
	jdff dff_A_oyVB0b665_0(.dout(w_dff_A_v0qq9xQJ7_0),.din(w_dff_A_oyVB0b665_0),.clk(gclk));
	jdff dff_A_8XfYXIVT6_0(.dout(w_dff_A_oyVB0b665_0),.din(w_dff_A_8XfYXIVT6_0),.clk(gclk));
	jdff dff_A_FmUb1ebN6_0(.dout(w_dff_A_8XfYXIVT6_0),.din(w_dff_A_FmUb1ebN6_0),.clk(gclk));
	jdff dff_A_bOi4UE0B1_0(.dout(w_dff_A_FmUb1ebN6_0),.din(w_dff_A_bOi4UE0B1_0),.clk(gclk));
	jdff dff_A_Wj38kN3O5_0(.dout(w_dff_A_bOi4UE0B1_0),.din(w_dff_A_Wj38kN3O5_0),.clk(gclk));
	jdff dff_A_kCc9f4Ez3_0(.dout(w_dff_A_Wj38kN3O5_0),.din(w_dff_A_kCc9f4Ez3_0),.clk(gclk));
	jdff dff_A_ym2UMXSd0_0(.dout(w_dff_A_kCc9f4Ez3_0),.din(w_dff_A_ym2UMXSd0_0),.clk(gclk));
	jdff dff_A_PkLqv2Px5_0(.dout(w_dff_A_ym2UMXSd0_0),.din(w_dff_A_PkLqv2Px5_0),.clk(gclk));
	jdff dff_A_iQSMFodB5_0(.dout(w_dff_A_PkLqv2Px5_0),.din(w_dff_A_iQSMFodB5_0),.clk(gclk));
	jdff dff_A_ASSNhaad5_0(.dout(w_dff_A_iQSMFodB5_0),.din(w_dff_A_ASSNhaad5_0),.clk(gclk));
	jdff dff_B_aFnTQLtg1_1(.din(n104),.dout(w_dff_B_aFnTQLtg1_1),.clk(gclk));
	jdff dff_A_x4CoadrC8_1(.dout(w_G224_0[1]),.din(w_dff_A_x4CoadrC8_1),.clk(gclk));
	jdff dff_B_mpwLwhvW6_0(.din(n101),.dout(w_dff_B_mpwLwhvW6_0),.clk(gclk));
	jdff dff_B_JxaDq2Ff9_0(.din(w_dff_B_mpwLwhvW6_0),.dout(w_dff_B_JxaDq2Ff9_0),.clk(gclk));
	jdff dff_A_9dENtCRg6_0(.dout(w_n99_0[0]),.din(w_dff_A_9dENtCRg6_0),.clk(gclk));
	jdff dff_A_TXUsMIO52_1(.dout(w_n96_0[1]),.din(w_dff_A_TXUsMIO52_1),.clk(gclk));
	jdff dff_A_4iQ5PsFD0_1(.dout(w_dff_A_TXUsMIO52_1),.din(w_dff_A_4iQ5PsFD0_1),.clk(gclk));
	jdff dff_A_SOb0HfFp1_2(.dout(w_n96_0[2]),.din(w_dff_A_SOb0HfFp1_2),.clk(gclk));
	jdff dff_A_DyND0V2T2_2(.dout(w_dff_A_SOb0HfFp1_2),.din(w_dff_A_DyND0V2T2_2),.clk(gclk));
	jdff dff_B_iZSNUWk79_3(.din(n96),.dout(w_dff_B_iZSNUWk79_3),.clk(gclk));
	jdff dff_B_sq9N4pXi0_3(.din(w_dff_B_iZSNUWk79_3),.dout(w_dff_B_sq9N4pXi0_3),.clk(gclk));
	jdff dff_A_JQVYE69n0_0(.dout(w_n95_1[0]),.din(w_dff_A_JQVYE69n0_0),.clk(gclk));
	jdff dff_A_hZVR3lWF6_0(.dout(w_dff_A_JQVYE69n0_0),.din(w_dff_A_hZVR3lWF6_0),.clk(gclk));
	jdff dff_A_PIaYCAmj5_1(.dout(w_n95_0[1]),.din(w_dff_A_PIaYCAmj5_1),.clk(gclk));
	jdff dff_A_wcBhESmt3_1(.dout(w_dff_A_PIaYCAmj5_1),.din(w_dff_A_wcBhESmt3_1),.clk(gclk));
	jdff dff_A_m9EiKjWD6_1(.dout(w_dff_A_wcBhESmt3_1),.din(w_dff_A_m9EiKjWD6_1),.clk(gclk));
	jdff dff_A_geY3g1Pp7_1(.dout(w_dff_A_m9EiKjWD6_1),.din(w_dff_A_geY3g1Pp7_1),.clk(gclk));
	jdff dff_A_4hau76MP3_1(.dout(w_dff_A_geY3g1Pp7_1),.din(w_dff_A_4hau76MP3_1),.clk(gclk));
	jdff dff_A_ZJ1LG8BS8_2(.dout(w_n95_0[2]),.din(w_dff_A_ZJ1LG8BS8_2),.clk(gclk));
	jdff dff_A_Mskq4TCj1_2(.dout(w_dff_A_ZJ1LG8BS8_2),.din(w_dff_A_Mskq4TCj1_2),.clk(gclk));
	jdff dff_A_laEriNyn6_2(.dout(w_dff_A_Mskq4TCj1_2),.din(w_dff_A_laEriNyn6_2),.clk(gclk));
	jdff dff_A_GrrdG6wv4_2(.dout(w_dff_A_laEriNyn6_2),.din(w_dff_A_GrrdG6wv4_2),.clk(gclk));
	jdff dff_A_woUgFLQV7_2(.dout(w_dff_A_GrrdG6wv4_2),.din(w_dff_A_woUgFLQV7_2),.clk(gclk));
	jdff dff_A_bZqGKQsJ5_1(.dout(w_n161_0[1]),.din(w_dff_A_bZqGKQsJ5_1),.clk(gclk));
	jdff dff_A_tUN8qgig9_2(.dout(w_n161_0[2]),.din(w_dff_A_tUN8qgig9_2),.clk(gclk));
	jdff dff_B_SmSmmBJM7_3(.din(n161),.dout(w_dff_B_SmSmmBJM7_3),.clk(gclk));
	jdff dff_B_AYMGgiWa9_1(.din(n159),.dout(w_dff_B_AYMGgiWa9_1),.clk(gclk));
	jdff dff_B_6H4SbxbY6_1(.din(w_dff_B_AYMGgiWa9_1),.dout(w_dff_B_6H4SbxbY6_1),.clk(gclk));
	jdff dff_B_yHm5oCLr0_1(.din(w_dff_B_6H4SbxbY6_1),.dout(w_dff_B_yHm5oCLr0_1),.clk(gclk));
	jdff dff_B_ZOuoeaeS6_1(.din(w_dff_B_yHm5oCLr0_1),.dout(w_dff_B_ZOuoeaeS6_1),.clk(gclk));
	jdff dff_B_P7OwcfVU5_1(.din(w_dff_B_ZOuoeaeS6_1),.dout(w_dff_B_P7OwcfVU5_1),.clk(gclk));
	jdff dff_A_kl9t13r57_0(.dout(w_n90_0[0]),.din(w_dff_A_kl9t13r57_0),.clk(gclk));
	jdff dff_A_TNj0WbIB7_0(.dout(w_dff_A_kl9t13r57_0),.din(w_dff_A_TNj0WbIB7_0),.clk(gclk));
	jdff dff_A_U89xG9Vd2_0(.dout(w_dff_A_TNj0WbIB7_0),.din(w_dff_A_U89xG9Vd2_0),.clk(gclk));
	jdff dff_A_fuuvUbSH8_0(.dout(w_dff_A_U89xG9Vd2_0),.din(w_dff_A_fuuvUbSH8_0),.clk(gclk));
	jdff dff_A_slbVTk6q2_0(.dout(w_dff_A_fuuvUbSH8_0),.din(w_dff_A_slbVTk6q2_0),.clk(gclk));
	jdff dff_A_G9t4kHd51_0(.dout(w_dff_A_slbVTk6q2_0),.din(w_dff_A_G9t4kHd51_0),.clk(gclk));
	jdff dff_A_2X9bSZv90_0(.dout(w_dff_A_G9t4kHd51_0),.din(w_dff_A_2X9bSZv90_0),.clk(gclk));
	jdff dff_A_NWg9P04g9_0(.dout(w_dff_A_2X9bSZv90_0),.din(w_dff_A_NWg9P04g9_0),.clk(gclk));
	jdff dff_A_clhh5mhz1_0(.dout(w_dff_A_NWg9P04g9_0),.din(w_dff_A_clhh5mhz1_0),.clk(gclk));
	jdff dff_A_qKPCwKQn3_0(.dout(w_dff_A_clhh5mhz1_0),.din(w_dff_A_qKPCwKQn3_0),.clk(gclk));
	jdff dff_A_ruJATUgD2_0(.dout(w_dff_A_qKPCwKQn3_0),.din(w_dff_A_ruJATUgD2_0),.clk(gclk));
	jdff dff_A_tU0QD92Y8_0(.dout(w_dff_A_ruJATUgD2_0),.din(w_dff_A_tU0QD92Y8_0),.clk(gclk));
	jdff dff_A_hB3DFJRv7_0(.dout(w_G210_0[0]),.din(w_dff_A_hB3DFJRv7_0),.clk(gclk));
	jdff dff_A_4xVr9j2f6_0(.dout(w_dff_A_hB3DFJRv7_0),.din(w_dff_A_4xVr9j2f6_0),.clk(gclk));
	jdff dff_A_mjXoH1J22_0(.dout(w_dff_A_4xVr9j2f6_0),.din(w_dff_A_mjXoH1J22_0),.clk(gclk));
	jdff dff_A_k6Pbvkn38_0(.dout(w_dff_A_mjXoH1J22_0),.din(w_dff_A_k6Pbvkn38_0),.clk(gclk));
	jdff dff_A_SGzMnbvN2_0(.dout(w_dff_A_k6Pbvkn38_0),.din(w_dff_A_SGzMnbvN2_0),.clk(gclk));
	jdff dff_A_jwQz4vQy2_0(.dout(w_dff_A_SGzMnbvN2_0),.din(w_dff_A_jwQz4vQy2_0),.clk(gclk));
	jdff dff_A_AXm7U6Us4_0(.dout(w_dff_A_jwQz4vQy2_0),.din(w_dff_A_AXm7U6Us4_0),.clk(gclk));
	jdff dff_A_zAgb3OdD2_0(.dout(w_dff_A_AXm7U6Us4_0),.din(w_dff_A_zAgb3OdD2_0),.clk(gclk));
	jdff dff_A_2V1e7Wgg3_0(.dout(w_dff_A_zAgb3OdD2_0),.din(w_dff_A_2V1e7Wgg3_0),.clk(gclk));
	jdff dff_A_vYQArisC2_0(.dout(w_dff_A_2V1e7Wgg3_0),.din(w_dff_A_vYQArisC2_0),.clk(gclk));
	jdff dff_A_4blA1VWQ2_0(.dout(w_dff_A_vYQArisC2_0),.din(w_dff_A_4blA1VWQ2_0),.clk(gclk));
	jdff dff_A_mgyOkLTl1_0(.dout(w_dff_A_4blA1VWQ2_0),.din(w_dff_A_mgyOkLTl1_0),.clk(gclk));
	jdff dff_A_JB0utwUz8_0(.dout(w_dff_A_mgyOkLTl1_0),.din(w_dff_A_JB0utwUz8_0),.clk(gclk));
	jdff dff_A_QrAafOiN1_0(.dout(w_dff_A_JB0utwUz8_0),.din(w_dff_A_QrAafOiN1_0),.clk(gclk));
	jdff dff_A_e7Eaff0f4_0(.dout(w_dff_A_QrAafOiN1_0),.din(w_dff_A_e7Eaff0f4_0),.clk(gclk));
	jdff dff_A_VyrqZWlM8_0(.dout(w_dff_A_e7Eaff0f4_0),.din(w_dff_A_VyrqZWlM8_0),.clk(gclk));
	jdff dff_A_2wciar0F4_1(.dout(w_G210_0[1]),.din(w_dff_A_2wciar0F4_1),.clk(gclk));
	jdff dff_A_eFk3xNBu3_0(.dout(w_G101_0[0]),.din(w_dff_A_eFk3xNBu3_0),.clk(gclk));
	jdff dff_A_pXDpby4W7_0(.dout(w_dff_A_eFk3xNBu3_0),.din(w_dff_A_pXDpby4W7_0),.clk(gclk));
	jdff dff_A_W2ztJ7SQ4_0(.dout(w_dff_A_pXDpby4W7_0),.din(w_dff_A_W2ztJ7SQ4_0),.clk(gclk));
	jdff dff_A_hvYfNHjT3_0(.dout(w_dff_A_W2ztJ7SQ4_0),.din(w_dff_A_hvYfNHjT3_0),.clk(gclk));
	jdff dff_A_5V4Ph5x29_0(.dout(w_dff_A_hvYfNHjT3_0),.din(w_dff_A_5V4Ph5x29_0),.clk(gclk));
	jdff dff_A_hH17uga58_0(.dout(w_dff_A_5V4Ph5x29_0),.din(w_dff_A_hH17uga58_0),.clk(gclk));
	jdff dff_A_NwXol6hV0_0(.dout(w_dff_A_hH17uga58_0),.din(w_dff_A_NwXol6hV0_0),.clk(gclk));
	jdff dff_A_M5IvXN4M6_0(.dout(w_dff_A_NwXol6hV0_0),.din(w_dff_A_M5IvXN4M6_0),.clk(gclk));
	jdff dff_A_DiOHebvu5_0(.dout(w_dff_A_M5IvXN4M6_0),.din(w_dff_A_DiOHebvu5_0),.clk(gclk));
	jdff dff_A_nHufrf4W8_0(.dout(w_dff_A_DiOHebvu5_0),.din(w_dff_A_nHufrf4W8_0),.clk(gclk));
	jdff dff_A_tkN9220D2_0(.dout(w_dff_A_nHufrf4W8_0),.din(w_dff_A_tkN9220D2_0),.clk(gclk));
	jdff dff_A_5yz7tMgP9_2(.dout(w_G101_0[2]),.din(w_dff_A_5yz7tMgP9_2),.clk(gclk));
	jdff dff_A_of9VE2Fz6_2(.dout(w_dff_A_5yz7tMgP9_2),.din(w_dff_A_of9VE2Fz6_2),.clk(gclk));
	jdff dff_A_ok4oxW2C4_1(.dout(w_n84_0[1]),.din(w_dff_A_ok4oxW2C4_1),.clk(gclk));
	jdff dff_A_jm8LVCm13_1(.dout(w_n81_0[1]),.din(w_dff_A_jm8LVCm13_1),.clk(gclk));
	jdff dff_A_wdagkMWX9_2(.dout(w_n81_0[2]),.din(w_dff_A_wdagkMWX9_2),.clk(gclk));
	jdff dff_A_HL6lsrHG2_2(.dout(w_G472_0[2]),.din(w_dff_A_HL6lsrHG2_2),.clk(gclk));
	jdff dff_A_jovm5fYq5_2(.dout(w_dff_A_HL6lsrHG2_2),.din(w_dff_A_jovm5fYq5_2),.clk(gclk));
	jdff dff_A_Ty6DqOdE5_2(.dout(w_dff_A_jovm5fYq5_2),.din(w_dff_A_Ty6DqOdE5_2),.clk(gclk));
	jdff dff_A_ux5drhZs3_2(.dout(w_dff_A_Ty6DqOdE5_2),.din(w_dff_A_ux5drhZs3_2),.clk(gclk));
	jdff dff_A_7PyvplTS7_2(.dout(w_dff_A_ux5drhZs3_2),.din(w_dff_A_7PyvplTS7_2),.clk(gclk));
	jdff dff_A_6gxqJhLc9_2(.dout(w_dff_A_7PyvplTS7_2),.din(w_dff_A_6gxqJhLc9_2),.clk(gclk));
	jdff dff_B_4qFwiVGm8_0(.din(n75),.dout(w_dff_B_4qFwiVGm8_0),.clk(gclk));
	jdff dff_A_atZXIHD73_0(.dout(w_n74_0[0]),.din(w_dff_A_atZXIHD73_0),.clk(gclk));
	jdff dff_A_qpoPMpyG5_0(.dout(w_dff_A_atZXIHD73_0),.din(w_dff_A_qpoPMpyG5_0),.clk(gclk));
	jdff dff_A_I9CkvksI5_0(.dout(w_n70_0[0]),.din(w_dff_A_I9CkvksI5_0),.clk(gclk));
	jdff dff_A_QHyjIXl35_0(.dout(w_dff_A_I9CkvksI5_0),.din(w_dff_A_QHyjIXl35_0),.clk(gclk));
	jdff dff_A_3YG4nnEL4_0(.dout(w_dff_A_QHyjIXl35_0),.din(w_dff_A_3YG4nnEL4_0),.clk(gclk));
	jdff dff_A_ene5vLYs2_0(.dout(w_dff_A_3YG4nnEL4_0),.din(w_dff_A_ene5vLYs2_0),.clk(gclk));
	jdff dff_A_GzlSrgQs0_0(.dout(w_dff_A_ene5vLYs2_0),.din(w_dff_A_GzlSrgQs0_0),.clk(gclk));
	jdff dff_A_jnLxujRO1_0(.dout(w_dff_A_GzlSrgQs0_0),.din(w_dff_A_jnLxujRO1_0),.clk(gclk));
	jdff dff_A_0LJTcGe11_0(.dout(w_dff_A_jnLxujRO1_0),.din(w_dff_A_0LJTcGe11_0),.clk(gclk));
	jdff dff_A_MqlHttQF1_0(.dout(w_dff_A_0LJTcGe11_0),.din(w_dff_A_MqlHttQF1_0),.clk(gclk));
	jdff dff_A_n7J2kp7O1_0(.dout(w_dff_A_MqlHttQF1_0),.din(w_dff_A_n7J2kp7O1_0),.clk(gclk));
	jdff dff_A_KailyL7u5_0(.dout(w_dff_A_n7J2kp7O1_0),.din(w_dff_A_KailyL7u5_0),.clk(gclk));
	jdff dff_A_QRFDXzvI1_0(.dout(w_dff_A_KailyL7u5_0),.din(w_dff_A_QRFDXzvI1_0),.clk(gclk));
	jdff dff_A_iDaGQMjD6_0(.dout(w_dff_A_QRFDXzvI1_0),.din(w_dff_A_iDaGQMjD6_0),.clk(gclk));
	jdff dff_A_12fiUFWN7_0(.dout(w_dff_A_iDaGQMjD6_0),.din(w_dff_A_12fiUFWN7_0),.clk(gclk));
	jdff dff_B_r8oAmEr11_0(.din(n69),.dout(w_dff_B_r8oAmEr11_0),.clk(gclk));
	jdff dff_B_LJSWXHrT7_0(.din(n68),.dout(w_dff_B_LJSWXHrT7_0),.clk(gclk));
	jdff dff_A_Yx99ZoGm0_0(.dout(w_G137_0[0]),.din(w_dff_A_Yx99ZoGm0_0),.clk(gclk));
	jdff dff_A_1E1OJPCW5_0(.dout(w_dff_A_Yx99ZoGm0_0),.din(w_dff_A_1E1OJPCW5_0),.clk(gclk));
	jdff dff_A_j7AwUOtD4_0(.dout(w_dff_A_1E1OJPCW5_0),.din(w_dff_A_j7AwUOtD4_0),.clk(gclk));
	jdff dff_A_6A9Lev4r5_0(.dout(w_dff_A_j7AwUOtD4_0),.din(w_dff_A_6A9Lev4r5_0),.clk(gclk));
	jdff dff_A_v3PehkQg4_0(.dout(w_dff_A_6A9Lev4r5_0),.din(w_dff_A_v3PehkQg4_0),.clk(gclk));
	jdff dff_A_Y5XU4Hfp1_0(.dout(w_dff_A_v3PehkQg4_0),.din(w_dff_A_Y5XU4Hfp1_0),.clk(gclk));
	jdff dff_A_LTvMCBkk0_0(.dout(w_dff_A_Y5XU4Hfp1_0),.din(w_dff_A_LTvMCBkk0_0),.clk(gclk));
	jdff dff_A_IfLVXqSD8_0(.dout(w_dff_A_LTvMCBkk0_0),.din(w_dff_A_IfLVXqSD8_0),.clk(gclk));
	jdff dff_A_qJTHVnl13_0(.dout(w_dff_A_IfLVXqSD8_0),.din(w_dff_A_qJTHVnl13_0),.clk(gclk));
	jdff dff_A_iF4bgQ0X4_0(.dout(w_dff_A_qJTHVnl13_0),.din(w_dff_A_iF4bgQ0X4_0),.clk(gclk));
	jdff dff_A_NV5cEZc60_0(.dout(w_dff_A_iF4bgQ0X4_0),.din(w_dff_A_NV5cEZc60_0),.clk(gclk));
	jdff dff_B_XiehfK7Z2_0(.din(n64),.dout(w_dff_B_XiehfK7Z2_0),.clk(gclk));
	jdff dff_A_pYCeHdjc8_0(.dout(w_G119_0[0]),.din(w_dff_A_pYCeHdjc8_0),.clk(gclk));
	jdff dff_A_iU8Vv90l2_0(.dout(w_dff_A_pYCeHdjc8_0),.din(w_dff_A_iU8Vv90l2_0),.clk(gclk));
	jdff dff_A_DDLbsdKx4_0(.dout(w_dff_A_iU8Vv90l2_0),.din(w_dff_A_DDLbsdKx4_0),.clk(gclk));
	jdff dff_A_MIOm2Y5d6_0(.dout(w_dff_A_DDLbsdKx4_0),.din(w_dff_A_MIOm2Y5d6_0),.clk(gclk));
	jdff dff_A_QOpjK0sa1_0(.dout(w_dff_A_MIOm2Y5d6_0),.din(w_dff_A_QOpjK0sa1_0),.clk(gclk));
	jdff dff_A_SNhItwJm2_0(.dout(w_dff_A_QOpjK0sa1_0),.din(w_dff_A_SNhItwJm2_0),.clk(gclk));
	jdff dff_A_m6rWxWNt5_0(.dout(w_dff_A_SNhItwJm2_0),.din(w_dff_A_m6rWxWNt5_0),.clk(gclk));
	jdff dff_A_kG3Sw8WA6_0(.dout(w_dff_A_m6rWxWNt5_0),.din(w_dff_A_kG3Sw8WA6_0),.clk(gclk));
	jdff dff_A_tUnhX7UW6_0(.dout(w_dff_A_kG3Sw8WA6_0),.din(w_dff_A_tUnhX7UW6_0),.clk(gclk));
	jdff dff_A_SFbsM8nx7_0(.dout(w_dff_A_tUnhX7UW6_0),.din(w_dff_A_SFbsM8nx7_0),.clk(gclk));
	jdff dff_A_zQr574PS7_0(.dout(w_dff_A_SFbsM8nx7_0),.din(w_dff_A_zQr574PS7_0),.clk(gclk));
	jdff dff_A_pnVt8Qtv5_2(.dout(w_G119_0[2]),.din(w_dff_A_pnVt8Qtv5_2),.clk(gclk));
	jdff dff_A_d8mwiH3Y7_0(.dout(w_G110_0[0]),.din(w_dff_A_d8mwiH3Y7_0),.clk(gclk));
	jdff dff_A_NVAp0T9d8_0(.dout(w_dff_A_d8mwiH3Y7_0),.din(w_dff_A_NVAp0T9d8_0),.clk(gclk));
	jdff dff_A_KvebgTYX9_0(.dout(w_dff_A_NVAp0T9d8_0),.din(w_dff_A_KvebgTYX9_0),.clk(gclk));
	jdff dff_A_lkrQ8U7C8_0(.dout(w_dff_A_KvebgTYX9_0),.din(w_dff_A_lkrQ8U7C8_0),.clk(gclk));
	jdff dff_A_zWtAHudD5_0(.dout(w_dff_A_lkrQ8U7C8_0),.din(w_dff_A_zWtAHudD5_0),.clk(gclk));
	jdff dff_A_kl2sIsMx1_0(.dout(w_dff_A_zWtAHudD5_0),.din(w_dff_A_kl2sIsMx1_0),.clk(gclk));
	jdff dff_A_p0tcYRmA8_0(.dout(w_dff_A_kl2sIsMx1_0),.din(w_dff_A_p0tcYRmA8_0),.clk(gclk));
	jdff dff_A_frApIrAX3_0(.dout(w_dff_A_p0tcYRmA8_0),.din(w_dff_A_frApIrAX3_0),.clk(gclk));
	jdff dff_A_YPTbDuYP4_0(.dout(w_dff_A_frApIrAX3_0),.din(w_dff_A_YPTbDuYP4_0),.clk(gclk));
	jdff dff_A_zwFgS79g3_0(.dout(w_dff_A_YPTbDuYP4_0),.din(w_dff_A_zwFgS79g3_0),.clk(gclk));
	jdff dff_A_VJyD25BW2_0(.dout(w_dff_A_zwFgS79g3_0),.din(w_dff_A_VJyD25BW2_0),.clk(gclk));
	jdff dff_B_LDZoSPUp5_1(.din(n59),.dout(w_dff_B_LDZoSPUp5_1),.clk(gclk));
	jdff dff_A_rh5X5q869_0(.dout(w_G234_1[0]),.din(w_dff_A_rh5X5q869_0),.clk(gclk));
	jdff dff_A_uC1SOD1I5_0(.dout(w_G221_0[0]),.din(w_dff_A_uC1SOD1I5_0),.clk(gclk));
	jdff dff_A_8kbSZhd42_0(.dout(w_dff_A_uC1SOD1I5_0),.din(w_dff_A_8kbSZhd42_0),.clk(gclk));
	jdff dff_A_UmkrL2Bk1_0(.dout(w_dff_A_8kbSZhd42_0),.din(w_dff_A_UmkrL2Bk1_0),.clk(gclk));
	jdff dff_A_XPV2EKVR7_0(.dout(w_n58_2[0]),.din(w_dff_A_XPV2EKVR7_0),.clk(gclk));
	jdff dff_A_5HXS80rJ5_0(.dout(w_dff_A_XPV2EKVR7_0),.din(w_dff_A_5HXS80rJ5_0),.clk(gclk));
	jdff dff_A_9srne13f0_0(.dout(w_dff_A_5HXS80rJ5_0),.din(w_dff_A_9srne13f0_0),.clk(gclk));
	jdff dff_A_IfPdIVTn7_0(.dout(w_dff_A_9srne13f0_0),.din(w_dff_A_IfPdIVTn7_0),.clk(gclk));
	jdff dff_A_oFeZ3aKP2_2(.dout(w_n58_2[2]),.din(w_dff_A_oFeZ3aKP2_2),.clk(gclk));
	jdff dff_A_51Ifwn6Q6_2(.dout(w_dff_A_oFeZ3aKP2_2),.din(w_dff_A_51Ifwn6Q6_2),.clk(gclk));
	jdff dff_A_sdkKZKsZ1_2(.dout(w_dff_A_51Ifwn6Q6_2),.din(w_dff_A_sdkKZKsZ1_2),.clk(gclk));
	jdff dff_A_H9Rx8CDR8_2(.dout(w_dff_A_sdkKZKsZ1_2),.din(w_dff_A_H9Rx8CDR8_2),.clk(gclk));
	jdff dff_A_ksj7tYHN6_0(.dout(w_n131_0[0]),.din(w_dff_A_ksj7tYHN6_0),.clk(gclk));
	jdff dff_A_Itc80Ea72_0(.dout(w_dff_A_ksj7tYHN6_0),.din(w_dff_A_Itc80Ea72_0),.clk(gclk));
	jdff dff_A_M39xwuIo0_0(.dout(w_dff_A_Itc80Ea72_0),.din(w_dff_A_M39xwuIo0_0),.clk(gclk));
	jdff dff_A_vjxMacjW1_2(.dout(w_n131_0[2]),.din(w_dff_A_vjxMacjW1_2),.clk(gclk));
	jdff dff_A_6kFU2oJx0_2(.dout(w_dff_A_vjxMacjW1_2),.din(w_dff_A_6kFU2oJx0_2),.clk(gclk));
	jdff dff_A_I3fxLiWP0_2(.dout(w_dff_A_6kFU2oJx0_2),.din(w_dff_A_I3fxLiWP0_2),.clk(gclk));
	jdff dff_A_UuNkoUaZ8_2(.dout(w_dff_A_I3fxLiWP0_2),.din(w_dff_A_UuNkoUaZ8_2),.clk(gclk));
	jdff dff_A_kdAG6Xfd1_2(.dout(w_dff_A_UuNkoUaZ8_2),.din(w_dff_A_kdAG6Xfd1_2),.clk(gclk));
	jdff dff_A_eGqH9LWf9_1(.dout(w_n130_0[1]),.din(w_dff_A_eGqH9LWf9_1),.clk(gclk));
	jdff dff_A_JxLCtbbS1_1(.dout(w_dff_A_eGqH9LWf9_1),.din(w_dff_A_JxLCtbbS1_1),.clk(gclk));
	jdff dff_A_lQnAgIGT8_1(.dout(w_dff_A_JxLCtbbS1_1),.din(w_dff_A_lQnAgIGT8_1),.clk(gclk));
	jdff dff_A_IHjKN1eP7_1(.dout(w_dff_A_lQnAgIGT8_1),.din(w_dff_A_IHjKN1eP7_1),.clk(gclk));
	jdff dff_A_TULZPGgB3_2(.dout(w_n130_0[2]),.din(w_dff_A_TULZPGgB3_2),.clk(gclk));
	jdff dff_A_PXokvH883_2(.dout(w_dff_A_TULZPGgB3_2),.din(w_dff_A_PXokvH883_2),.clk(gclk));
	jdff dff_A_6O1qeEnr7_2(.dout(w_dff_A_PXokvH883_2),.din(w_dff_A_6O1qeEnr7_2),.clk(gclk));
	jdff dff_A_ranaXLiv7_2(.dout(w_dff_A_6O1qeEnr7_2),.din(w_dff_A_ranaXLiv7_2),.clk(gclk));
	jdff dff_A_B7FQSY6u3_2(.dout(w_dff_A_ranaXLiv7_2),.din(w_dff_A_B7FQSY6u3_2),.clk(gclk));
	jdff dff_A_lCVW8TrR0_2(.dout(w_dff_A_B7FQSY6u3_2),.din(w_dff_A_lCVW8TrR0_2),.clk(gclk));
	jdff dff_A_5UsLVNNZ0_2(.dout(w_dff_A_lCVW8TrR0_2),.din(w_dff_A_5UsLVNNZ0_2),.clk(gclk));
	jdff dff_A_mf0Nb3ry8_2(.dout(w_dff_A_5UsLVNNZ0_2),.din(w_dff_A_mf0Nb3ry8_2),.clk(gclk));
	jdff dff_A_oEm0Nfpx8_2(.dout(w_dff_A_mf0Nb3ry8_2),.din(w_dff_A_oEm0Nfpx8_2),.clk(gclk));
	jdff dff_A_raUcn9Zs3_0(.dout(w_n124_0[0]),.din(w_dff_A_raUcn9Zs3_0),.clk(gclk));
	jdff dff_A_HRi1yhR67_1(.dout(w_G898_0[1]),.din(w_dff_A_HRi1yhR67_1),.clk(gclk));
	jdff dff_A_SipQVlaa6_0(.dout(w_n186_0[0]),.din(w_dff_A_SipQVlaa6_0),.clk(gclk));
	jdff dff_A_lZsDVJ0U6_0(.dout(w_dff_A_SipQVlaa6_0),.din(w_dff_A_lZsDVJ0U6_0),.clk(gclk));
	jdff dff_A_zbzxFhuo2_0(.dout(w_dff_A_lZsDVJ0U6_0),.din(w_dff_A_zbzxFhuo2_0),.clk(gclk));
	jdff dff_A_uI0Twndm0_1(.dout(w_n151_0[1]),.din(w_dff_A_uI0Twndm0_1),.clk(gclk));
	jdff dff_A_ZMcwRGWY9_1(.dout(w_dff_A_uI0Twndm0_1),.din(w_dff_A_ZMcwRGWY9_1),.clk(gclk));
	jdff dff_A_0Q9UZn8v8_1(.dout(w_dff_A_ZMcwRGWY9_1),.din(w_dff_A_0Q9UZn8v8_1),.clk(gclk));
	jdff dff_A_tod14Z6Y6_1(.dout(w_dff_A_0Q9UZn8v8_1),.din(w_dff_A_tod14Z6Y6_1),.clk(gclk));
	jdff dff_A_n8swF2ru4_1(.dout(w_dff_A_tod14Z6Y6_1),.din(w_dff_A_n8swF2ru4_1),.clk(gclk));
	jdff dff_A_zUrRyy1A7_1(.dout(w_dff_A_n8swF2ru4_1),.din(w_dff_A_zUrRyy1A7_1),.clk(gclk));
	jdff dff_A_EAxCJBL25_1(.dout(w_dff_A_zUrRyy1A7_1),.din(w_dff_A_EAxCJBL25_1),.clk(gclk));
	jdff dff_A_QKGNkm4x4_1(.dout(w_dff_A_EAxCJBL25_1),.din(w_dff_A_QKGNkm4x4_1),.clk(gclk));
	jdff dff_A_ZwthStk77_1(.dout(w_dff_A_QKGNkm4x4_1),.din(w_dff_A_ZwthStk77_1),.clk(gclk));
	jdff dff_A_w9kyeGvU5_1(.dout(w_dff_A_ZwthStk77_1),.din(w_dff_A_w9kyeGvU5_1),.clk(gclk));
	jdff dff_A_pqYUnlPZ3_1(.dout(w_dff_A_w9kyeGvU5_1),.din(w_dff_A_pqYUnlPZ3_1),.clk(gclk));
	jdff dff_A_oAl19vRy1_1(.dout(w_dff_A_pqYUnlPZ3_1),.din(w_dff_A_oAl19vRy1_1),.clk(gclk));
	jdff dff_B_MznmxNAg2_1(.din(n144),.dout(w_dff_B_MznmxNAg2_1),.clk(gclk));
	jdff dff_B_Ny6Ilyp92_1(.din(w_dff_B_MznmxNAg2_1),.dout(w_dff_B_Ny6Ilyp92_1),.clk(gclk));
	jdff dff_A_IU5JvZM81_0(.dout(w_G131_0[0]),.din(w_dff_A_IU5JvZM81_0),.clk(gclk));
	jdff dff_A_fUlEsfb87_0(.dout(w_dff_A_IU5JvZM81_0),.din(w_dff_A_fUlEsfb87_0),.clk(gclk));
	jdff dff_A_QoXljbPT5_0(.dout(w_dff_A_fUlEsfb87_0),.din(w_dff_A_QoXljbPT5_0),.clk(gclk));
	jdff dff_A_DZezbzRa5_0(.dout(w_dff_A_QoXljbPT5_0),.din(w_dff_A_DZezbzRa5_0),.clk(gclk));
	jdff dff_A_wGEc2Yr71_0(.dout(w_dff_A_DZezbzRa5_0),.din(w_dff_A_wGEc2Yr71_0),.clk(gclk));
	jdff dff_A_QOh7BTgc6_0(.dout(w_dff_A_wGEc2Yr71_0),.din(w_dff_A_QOh7BTgc6_0),.clk(gclk));
	jdff dff_A_ooAehbF87_0(.dout(w_dff_A_QOh7BTgc6_0),.din(w_dff_A_ooAehbF87_0),.clk(gclk));
	jdff dff_A_D6q22Tbe9_0(.dout(w_dff_A_ooAehbF87_0),.din(w_dff_A_D6q22Tbe9_0),.clk(gclk));
	jdff dff_A_I8DYA9Qv1_0(.dout(w_dff_A_D6q22Tbe9_0),.din(w_dff_A_I8DYA9Qv1_0),.clk(gclk));
	jdff dff_A_evfcDjfb0_0(.dout(w_dff_A_I8DYA9Qv1_0),.din(w_dff_A_evfcDjfb0_0),.clk(gclk));
	jdff dff_A_ttSlfJ5X7_0(.dout(w_dff_A_evfcDjfb0_0),.din(w_dff_A_ttSlfJ5X7_0),.clk(gclk));
	jdff dff_A_CzsLeHrX3_2(.dout(w_G131_0[2]),.din(w_dff_A_CzsLeHrX3_2),.clk(gclk));
	jdff dff_A_4wyfpWne7_1(.dout(w_G953_2[1]),.din(w_dff_A_4wyfpWne7_1),.clk(gclk));
	jdff dff_A_1s77Wb1L3_1(.dout(w_G214_0[1]),.din(w_dff_A_1s77Wb1L3_1),.clk(gclk));
	jdff dff_A_Hri4DIpK9_0(.dout(w_n67_0[0]),.din(w_dff_A_Hri4DIpK9_0),.clk(gclk));
	jdff dff_A_i447xYnj1_0(.dout(w_n66_0[0]),.din(w_dff_A_i447xYnj1_0),.clk(gclk));
	jdff dff_A_keIiaf2X8_0(.dout(w_dff_A_i447xYnj1_0),.din(w_dff_A_keIiaf2X8_0),.clk(gclk));
	jdff dff_A_rdWeC6J85_0(.dout(w_G140_0[0]),.din(w_dff_A_rdWeC6J85_0),.clk(gclk));
	jdff dff_A_BDE4x2dQ5_0(.dout(w_dff_A_rdWeC6J85_0),.din(w_dff_A_BDE4x2dQ5_0),.clk(gclk));
	jdff dff_A_h0zXj6WS3_0(.dout(w_dff_A_BDE4x2dQ5_0),.din(w_dff_A_h0zXj6WS3_0),.clk(gclk));
	jdff dff_A_voyEWAbT6_0(.dout(w_dff_A_h0zXj6WS3_0),.din(w_dff_A_voyEWAbT6_0),.clk(gclk));
	jdff dff_A_THTWZ5bi7_0(.dout(w_dff_A_voyEWAbT6_0),.din(w_dff_A_THTWZ5bi7_0),.clk(gclk));
	jdff dff_A_To3tX07H9_0(.dout(w_dff_A_THTWZ5bi7_0),.din(w_dff_A_To3tX07H9_0),.clk(gclk));
	jdff dff_A_e4q1WrRp3_0(.dout(w_dff_A_To3tX07H9_0),.din(w_dff_A_e4q1WrRp3_0),.clk(gclk));
	jdff dff_A_LpAuHaD96_0(.dout(w_dff_A_e4q1WrRp3_0),.din(w_dff_A_LpAuHaD96_0),.clk(gclk));
	jdff dff_A_FVrwDWEu1_0(.dout(w_dff_A_LpAuHaD96_0),.din(w_dff_A_FVrwDWEu1_0),.clk(gclk));
	jdff dff_A_tg2iyD9N2_0(.dout(w_dff_A_FVrwDWEu1_0),.din(w_dff_A_tg2iyD9N2_0),.clk(gclk));
	jdff dff_A_muDEwOhg9_0(.dout(w_dff_A_tg2iyD9N2_0),.din(w_dff_A_muDEwOhg9_0),.clk(gclk));
	jdff dff_A_ZPd97mhW6_1(.dout(w_G140_0[1]),.din(w_dff_A_ZPd97mhW6_1),.clk(gclk));
	jdff dff_A_cXjJ8Opy8_0(.dout(w_G125_0[0]),.din(w_dff_A_cXjJ8Opy8_0),.clk(gclk));
	jdff dff_A_7ke4v4vb5_0(.dout(w_dff_A_cXjJ8Opy8_0),.din(w_dff_A_7ke4v4vb5_0),.clk(gclk));
	jdff dff_A_rD8LgLhk2_0(.dout(w_dff_A_7ke4v4vb5_0),.din(w_dff_A_rD8LgLhk2_0),.clk(gclk));
	jdff dff_A_z2yKjB7S3_0(.dout(w_dff_A_rD8LgLhk2_0),.din(w_dff_A_z2yKjB7S3_0),.clk(gclk));
	jdff dff_A_bx9JhTvo5_0(.dout(w_dff_A_z2yKjB7S3_0),.din(w_dff_A_bx9JhTvo5_0),.clk(gclk));
	jdff dff_A_tMyZlCyb5_0(.dout(w_dff_A_bx9JhTvo5_0),.din(w_dff_A_tMyZlCyb5_0),.clk(gclk));
	jdff dff_A_szBWCZSm2_0(.dout(w_dff_A_tMyZlCyb5_0),.din(w_dff_A_szBWCZSm2_0),.clk(gclk));
	jdff dff_A_2S0qgKkv2_0(.dout(w_dff_A_szBWCZSm2_0),.din(w_dff_A_2S0qgKkv2_0),.clk(gclk));
	jdff dff_A_zZLvdgRX9_0(.dout(w_dff_A_2S0qgKkv2_0),.din(w_dff_A_zZLvdgRX9_0),.clk(gclk));
	jdff dff_A_LcBNfvQP6_0(.dout(w_dff_A_zZLvdgRX9_0),.din(w_dff_A_LcBNfvQP6_0),.clk(gclk));
	jdff dff_A_tFgBrtCK8_0(.dout(w_dff_A_LcBNfvQP6_0),.din(w_dff_A_tFgBrtCK8_0),.clk(gclk));
	jdff dff_A_0z7d7R0o8_1(.dout(w_G125_0[1]),.din(w_dff_A_0z7d7R0o8_1),.clk(gclk));
	jdff dff_A_5e6SVyaf6_1(.dout(w_dff_A_0z7d7R0o8_1),.din(w_dff_A_5e6SVyaf6_1),.clk(gclk));
	jdff dff_A_oSJkky0K2_0(.dout(w_G146_0[0]),.din(w_dff_A_oSJkky0K2_0),.clk(gclk));
	jdff dff_A_MigrqXIy2_0(.dout(w_dff_A_oSJkky0K2_0),.din(w_dff_A_MigrqXIy2_0),.clk(gclk));
	jdff dff_A_51TVHLii9_0(.dout(w_dff_A_MigrqXIy2_0),.din(w_dff_A_51TVHLii9_0),.clk(gclk));
	jdff dff_A_qTNc97ON5_0(.dout(w_dff_A_51TVHLii9_0),.din(w_dff_A_qTNc97ON5_0),.clk(gclk));
	jdff dff_A_TSwgDWBk9_0(.dout(w_dff_A_qTNc97ON5_0),.din(w_dff_A_TSwgDWBk9_0),.clk(gclk));
	jdff dff_A_UmJmSd2S3_0(.dout(w_dff_A_TSwgDWBk9_0),.din(w_dff_A_UmJmSd2S3_0),.clk(gclk));
	jdff dff_A_ZFmGawyg9_0(.dout(w_dff_A_UmJmSd2S3_0),.din(w_dff_A_ZFmGawyg9_0),.clk(gclk));
	jdff dff_A_5VP60dUO9_0(.dout(w_dff_A_ZFmGawyg9_0),.din(w_dff_A_5VP60dUO9_0),.clk(gclk));
	jdff dff_A_sNAq7mdA3_0(.dout(w_dff_A_5VP60dUO9_0),.din(w_dff_A_sNAq7mdA3_0),.clk(gclk));
	jdff dff_A_DX3jurAJ6_0(.dout(w_dff_A_sNAq7mdA3_0),.din(w_dff_A_DX3jurAJ6_0),.clk(gclk));
	jdff dff_B_QYOxYyQh7_3(.din(G146),.dout(w_dff_B_QYOxYyQh7_3),.clk(gclk));
	jdff dff_A_q10kKYis6_0(.dout(w_G113_0[0]),.din(w_dff_A_q10kKYis6_0),.clk(gclk));
	jdff dff_A_xIbWc7Ky0_0(.dout(w_dff_A_q10kKYis6_0),.din(w_dff_A_xIbWc7Ky0_0),.clk(gclk));
	jdff dff_A_gWk1F5el2_0(.dout(w_dff_A_xIbWc7Ky0_0),.din(w_dff_A_gWk1F5el2_0),.clk(gclk));
	jdff dff_A_mk8zZIpv4_0(.dout(w_dff_A_gWk1F5el2_0),.din(w_dff_A_mk8zZIpv4_0),.clk(gclk));
	jdff dff_A_bpPjve709_0(.dout(w_dff_A_mk8zZIpv4_0),.din(w_dff_A_bpPjve709_0),.clk(gclk));
	jdff dff_A_HFEBdRvo1_0(.dout(w_dff_A_bpPjve709_0),.din(w_dff_A_HFEBdRvo1_0),.clk(gclk));
	jdff dff_A_T3f7AEBb4_0(.dout(w_dff_A_HFEBdRvo1_0),.din(w_dff_A_T3f7AEBb4_0),.clk(gclk));
	jdff dff_A_x38dOZzJ8_0(.dout(w_dff_A_T3f7AEBb4_0),.din(w_dff_A_x38dOZzJ8_0),.clk(gclk));
	jdff dff_A_QAexxTV21_0(.dout(w_dff_A_x38dOZzJ8_0),.din(w_dff_A_QAexxTV21_0),.clk(gclk));
	jdff dff_A_AYKDvV884_0(.dout(w_dff_A_QAexxTV21_0),.din(w_dff_A_AYKDvV884_0),.clk(gclk));
	jdff dff_A_NWJHmVeC7_0(.dout(w_dff_A_AYKDvV884_0),.din(w_dff_A_NWJHmVeC7_0),.clk(gclk));
	jdff dff_A_O6x76RM51_0(.dout(w_G104_0[0]),.din(w_dff_A_O6x76RM51_0),.clk(gclk));
	jdff dff_A_b90dULUd8_0(.dout(w_dff_A_O6x76RM51_0),.din(w_dff_A_b90dULUd8_0),.clk(gclk));
	jdff dff_A_w4W009VD0_0(.dout(w_dff_A_b90dULUd8_0),.din(w_dff_A_w4W009VD0_0),.clk(gclk));
	jdff dff_A_UzgZewKc1_0(.dout(w_dff_A_w4W009VD0_0),.din(w_dff_A_UzgZewKc1_0),.clk(gclk));
	jdff dff_A_BTydVxyW5_0(.dout(w_dff_A_UzgZewKc1_0),.din(w_dff_A_BTydVxyW5_0),.clk(gclk));
	jdff dff_A_8JAonBZg2_0(.dout(w_dff_A_BTydVxyW5_0),.din(w_dff_A_8JAonBZg2_0),.clk(gclk));
	jdff dff_A_ttCS3nBG4_0(.dout(w_dff_A_8JAonBZg2_0),.din(w_dff_A_ttCS3nBG4_0),.clk(gclk));
	jdff dff_A_1mz5hszx0_0(.dout(w_dff_A_ttCS3nBG4_0),.din(w_dff_A_1mz5hszx0_0),.clk(gclk));
	jdff dff_A_2FjiCEY75_0(.dout(w_dff_A_1mz5hszx0_0),.din(w_dff_A_2FjiCEY75_0),.clk(gclk));
	jdff dff_A_f6iP0Ym57_0(.dout(w_dff_A_2FjiCEY75_0),.din(w_dff_A_f6iP0Ym57_0),.clk(gclk));
	jdff dff_A_FBAHzrOq1_0(.dout(w_dff_A_f6iP0Ym57_0),.din(w_dff_A_FBAHzrOq1_0),.clk(gclk));
	jdff dff_A_eUbbvWIE2_1(.dout(w_G104_0[1]),.din(w_dff_A_eUbbvWIE2_1),.clk(gclk));
	jdff dff_A_gxkjBzf02_1(.dout(w_G475_0[1]),.din(w_dff_A_gxkjBzf02_1),.clk(gclk));
	jdff dff_A_ZliZVfE29_1(.dout(w_dff_A_gxkjBzf02_1),.din(w_dff_A_ZliZVfE29_1),.clk(gclk));
	jdff dff_A_RMrCSklw6_1(.dout(w_dff_A_ZliZVfE29_1),.din(w_dff_A_RMrCSklw6_1),.clk(gclk));
	jdff dff_A_RjTJWRhP6_1(.dout(w_dff_A_RMrCSklw6_1),.din(w_dff_A_RjTJWRhP6_1),.clk(gclk));
	jdff dff_A_wrzlxhLN1_1(.dout(w_dff_A_RjTJWRhP6_1),.din(w_dff_A_wrzlxhLN1_1),.clk(gclk));
	jdff dff_A_kUu1Mzls8_1(.dout(w_dff_A_wrzlxhLN1_1),.din(w_dff_A_kUu1Mzls8_1),.clk(gclk));
	jdff dff_A_xUoOSNcT2_0(.dout(w_n139_0[0]),.din(w_dff_A_xUoOSNcT2_0),.clk(gclk));
	jdff dff_A_mcS7BPxg3_0(.dout(w_dff_A_xUoOSNcT2_0),.din(w_dff_A_mcS7BPxg3_0),.clk(gclk));
	jdff dff_A_YwwUhA365_0(.dout(w_dff_A_mcS7BPxg3_0),.din(w_dff_A_YwwUhA365_0),.clk(gclk));
	jdff dff_A_Qja3vFFE1_0(.dout(w_dff_A_YwwUhA365_0),.din(w_dff_A_Qja3vFFE1_0),.clk(gclk));
	jdff dff_A_hgcMTnVZ5_0(.dout(w_dff_A_Qja3vFFE1_0),.din(w_dff_A_hgcMTnVZ5_0),.clk(gclk));
	jdff dff_A_oF4bRuhQ9_0(.dout(w_dff_A_hgcMTnVZ5_0),.din(w_dff_A_oF4bRuhQ9_0),.clk(gclk));
	jdff dff_A_9PowGjIE1_0(.dout(w_dff_A_oF4bRuhQ9_0),.din(w_dff_A_9PowGjIE1_0),.clk(gclk));
	jdff dff_A_VvIYXqj79_0(.dout(w_dff_A_9PowGjIE1_0),.din(w_dff_A_VvIYXqj79_0),.clk(gclk));
	jdff dff_A_2vxRWCz35_0(.dout(w_dff_A_VvIYXqj79_0),.din(w_dff_A_2vxRWCz35_0),.clk(gclk));
	jdff dff_A_1xla2iDB4_0(.dout(w_dff_A_2vxRWCz35_0),.din(w_dff_A_1xla2iDB4_0),.clk(gclk));
	jdff dff_A_5YYL5PxY7_0(.dout(w_dff_A_1xla2iDB4_0),.din(w_dff_A_5YYL5PxY7_0),.clk(gclk));
	jdff dff_A_6MTAriep6_0(.dout(w_dff_A_5YYL5PxY7_0),.din(w_dff_A_6MTAriep6_0),.clk(gclk));
	jdff dff_A_POImPkBN8_0(.dout(w_dff_A_6MTAriep6_0),.din(w_dff_A_POImPkBN8_0),.clk(gclk));
	jdff dff_B_rSeBfPmu5_1(.din(n133),.dout(w_dff_B_rSeBfPmu5_1),.clk(gclk));
	jdff dff_B_CN858ycW5_1(.din(w_dff_B_rSeBfPmu5_1),.dout(w_dff_B_CN858ycW5_1),.clk(gclk));
	jdff dff_B_bm62cSlV3_0(.din(n137),.dout(w_dff_B_bm62cSlV3_0),.clk(gclk));
	jdff dff_A_IJjrdxt81_1(.dout(w_G122_0[1]),.din(w_dff_A_IJjrdxt81_1),.clk(gclk));
	jdff dff_A_Y3wHbrTA3_1(.dout(w_dff_A_IJjrdxt81_1),.din(w_dff_A_Y3wHbrTA3_1),.clk(gclk));
	jdff dff_A_MQYJhE4y9_1(.dout(w_dff_A_Y3wHbrTA3_1),.din(w_dff_A_MQYJhE4y9_1),.clk(gclk));
	jdff dff_A_EQX7NdHE4_1(.dout(w_dff_A_MQYJhE4y9_1),.din(w_dff_A_EQX7NdHE4_1),.clk(gclk));
	jdff dff_A_VBLw9gIW4_1(.dout(w_dff_A_EQX7NdHE4_1),.din(w_dff_A_VBLw9gIW4_1),.clk(gclk));
	jdff dff_A_uHo0OgwD3_1(.dout(w_dff_A_VBLw9gIW4_1),.din(w_dff_A_uHo0OgwD3_1),.clk(gclk));
	jdff dff_A_8E6CQeG16_1(.dout(w_dff_A_uHo0OgwD3_1),.din(w_dff_A_8E6CQeG16_1),.clk(gclk));
	jdff dff_A_6Z6ifrbO5_1(.dout(w_dff_A_8E6CQeG16_1),.din(w_dff_A_6Z6ifrbO5_1),.clk(gclk));
	jdff dff_A_dSleeQiT2_1(.dout(w_dff_A_6Z6ifrbO5_1),.din(w_dff_A_dSleeQiT2_1),.clk(gclk));
	jdff dff_A_MFjApbeP1_1(.dout(w_dff_A_dSleeQiT2_1),.din(w_dff_A_MFjApbeP1_1),.clk(gclk));
	jdff dff_A_i3wbb3jA9_1(.dout(w_dff_A_MFjApbeP1_1),.din(w_dff_A_i3wbb3jA9_1),.clk(gclk));
	jdff dff_A_68C1tYLB7_1(.dout(w_dff_A_i3wbb3jA9_1),.din(w_dff_A_68C1tYLB7_1),.clk(gclk));
	jdff dff_A_nga2Iew62_0(.dout(w_G116_0[0]),.din(w_dff_A_nga2Iew62_0),.clk(gclk));
	jdff dff_A_Prbkge5E7_0(.dout(w_dff_A_nga2Iew62_0),.din(w_dff_A_Prbkge5E7_0),.clk(gclk));
	jdff dff_A_nyqnGPiK0_0(.dout(w_dff_A_Prbkge5E7_0),.din(w_dff_A_nyqnGPiK0_0),.clk(gclk));
	jdff dff_A_g30tdJAs5_0(.dout(w_dff_A_nyqnGPiK0_0),.din(w_dff_A_g30tdJAs5_0),.clk(gclk));
	jdff dff_A_57r37bCg9_0(.dout(w_dff_A_g30tdJAs5_0),.din(w_dff_A_57r37bCg9_0),.clk(gclk));
	jdff dff_A_RnaV8Cpi8_0(.dout(w_dff_A_57r37bCg9_0),.din(w_dff_A_RnaV8Cpi8_0),.clk(gclk));
	jdff dff_A_3wMrxpah6_0(.dout(w_dff_A_RnaV8Cpi8_0),.din(w_dff_A_3wMrxpah6_0),.clk(gclk));
	jdff dff_A_TiER8Ba95_0(.dout(w_dff_A_3wMrxpah6_0),.din(w_dff_A_TiER8Ba95_0),.clk(gclk));
	jdff dff_A_0bVYrvQ19_0(.dout(w_dff_A_TiER8Ba95_0),.din(w_dff_A_0bVYrvQ19_0),.clk(gclk));
	jdff dff_A_N5DlPHLb0_0(.dout(w_dff_A_0bVYrvQ19_0),.din(w_dff_A_N5DlPHLb0_0),.clk(gclk));
	jdff dff_A_NLyaARlw7_0(.dout(w_dff_A_N5DlPHLb0_0),.din(w_dff_A_NLyaARlw7_0),.clk(gclk));
	jdff dff_A_49YsQQxQ0_0(.dout(w_G107_0[0]),.din(w_dff_A_49YsQQxQ0_0),.clk(gclk));
	jdff dff_A_8p83rKFq1_0(.dout(w_dff_A_49YsQQxQ0_0),.din(w_dff_A_8p83rKFq1_0),.clk(gclk));
	jdff dff_A_iUkqLGaB4_0(.dout(w_dff_A_8p83rKFq1_0),.din(w_dff_A_iUkqLGaB4_0),.clk(gclk));
	jdff dff_A_yRgsuM321_0(.dout(w_dff_A_iUkqLGaB4_0),.din(w_dff_A_yRgsuM321_0),.clk(gclk));
	jdff dff_A_vVB9dRLj0_0(.dout(w_dff_A_yRgsuM321_0),.din(w_dff_A_vVB9dRLj0_0),.clk(gclk));
	jdff dff_A_2zdQqUdi1_0(.dout(w_dff_A_vVB9dRLj0_0),.din(w_dff_A_2zdQqUdi1_0),.clk(gclk));
	jdff dff_A_qtxv1z6j6_0(.dout(w_dff_A_2zdQqUdi1_0),.din(w_dff_A_qtxv1z6j6_0),.clk(gclk));
	jdff dff_A_9oU8Yl8g4_0(.dout(w_dff_A_qtxv1z6j6_0),.din(w_dff_A_9oU8Yl8g4_0),.clk(gclk));
	jdff dff_A_rh4Mc7Np3_0(.dout(w_dff_A_9oU8Yl8g4_0),.din(w_dff_A_rh4Mc7Np3_0),.clk(gclk));
	jdff dff_A_yuS9hSMZ4_0(.dout(w_dff_A_rh4Mc7Np3_0),.din(w_dff_A_yuS9hSMZ4_0),.clk(gclk));
	jdff dff_A_CesXBU2u2_0(.dout(w_dff_A_yuS9hSMZ4_0),.din(w_dff_A_CesXBU2u2_0),.clk(gclk));
	jdff dff_A_6FeGUKFN4_1(.dout(w_G107_0[1]),.din(w_dff_A_6FeGUKFN4_1),.clk(gclk));
	jdff dff_A_bly7LfRR9_2(.dout(w_n103_2[2]),.din(w_dff_A_bly7LfRR9_2),.clk(gclk));
	jdff dff_A_kfr5z0gz9_2(.dout(w_dff_A_bly7LfRR9_2),.din(w_dff_A_kfr5z0gz9_2),.clk(gclk));
	jdff dff_A_XAwPxIpV3_1(.dout(w_G234_0[1]),.din(w_dff_A_XAwPxIpV3_1),.clk(gclk));
	jdff dff_A_AaRWqBMq8_0(.dout(w_G217_0[0]),.din(w_dff_A_AaRWqBMq8_0),.clk(gclk));
	jdff dff_A_9P4CbAt02_0(.dout(w_dff_A_AaRWqBMq8_0),.din(w_dff_A_9P4CbAt02_0),.clk(gclk));
	jdff dff_A_dcESeOtO4_0(.dout(w_dff_A_9P4CbAt02_0),.din(w_dff_A_dcESeOtO4_0),.clk(gclk));
	jdff dff_A_pDr1Ffty0_0(.dout(w_dff_A_dcESeOtO4_0),.din(w_dff_A_pDr1Ffty0_0),.clk(gclk));
	jdff dff_A_1XeUmfh58_0(.dout(w_dff_A_pDr1Ffty0_0),.din(w_dff_A_1XeUmfh58_0),.clk(gclk));
	jdff dff_A_UN32hoSG4_0(.dout(w_dff_A_1XeUmfh58_0),.din(w_dff_A_UN32hoSG4_0),.clk(gclk));
	jdff dff_A_hSTybxa97_0(.dout(w_dff_A_UN32hoSG4_0),.din(w_dff_A_hSTybxa97_0),.clk(gclk));
	jdff dff_A_gY1PkqQ66_0(.dout(w_dff_A_hSTybxa97_0),.din(w_dff_A_gY1PkqQ66_0),.clk(gclk));
	jdff dff_A_zKFyXN3O9_0(.dout(w_dff_A_gY1PkqQ66_0),.din(w_dff_A_zKFyXN3O9_0),.clk(gclk));
	jdff dff_A_P0HFjRp93_0(.dout(w_dff_A_zKFyXN3O9_0),.din(w_dff_A_P0HFjRp93_0),.clk(gclk));
	jdff dff_A_oTlpMXOD9_0(.dout(w_dff_A_P0HFjRp93_0),.din(w_dff_A_oTlpMXOD9_0),.clk(gclk));
	jdff dff_A_AjRwY4x19_0(.dout(w_dff_A_oTlpMXOD9_0),.din(w_dff_A_AjRwY4x19_0),.clk(gclk));
	jdff dff_A_sI67HIFr7_0(.dout(w_dff_A_AjRwY4x19_0),.din(w_dff_A_sI67HIFr7_0),.clk(gclk));
	jdff dff_A_mYZjQoQo4_0(.dout(w_dff_A_sI67HIFr7_0),.din(w_dff_A_mYZjQoQo4_0),.clk(gclk));
	jdff dff_A_JcBqaPAX3_2(.dout(w_G217_0[2]),.din(w_dff_A_JcBqaPAX3_2),.clk(gclk));
	jdff dff_B_oh5QZlDJ4_3(.din(G217),.dout(w_dff_B_oh5QZlDJ4_3),.clk(gclk));
	jdff dff_B_M3j6QPic7_3(.din(w_dff_B_oh5QZlDJ4_3),.dout(w_dff_B_M3j6QPic7_3),.clk(gclk));
	jdff dff_A_DcTb4TUm5_0(.dout(w_G143_0[0]),.din(w_dff_A_DcTb4TUm5_0),.clk(gclk));
	jdff dff_A_fSoIHhZ60_0(.dout(w_dff_A_DcTb4TUm5_0),.din(w_dff_A_fSoIHhZ60_0),.clk(gclk));
	jdff dff_A_UFQDDTAz1_0(.dout(w_dff_A_fSoIHhZ60_0),.din(w_dff_A_UFQDDTAz1_0),.clk(gclk));
	jdff dff_A_tqndewNR1_0(.dout(w_dff_A_UFQDDTAz1_0),.din(w_dff_A_tqndewNR1_0),.clk(gclk));
	jdff dff_A_msk2iWml3_0(.dout(w_dff_A_tqndewNR1_0),.din(w_dff_A_msk2iWml3_0),.clk(gclk));
	jdff dff_A_g6NQHAoh9_0(.dout(w_dff_A_msk2iWml3_0),.din(w_dff_A_g6NQHAoh9_0),.clk(gclk));
	jdff dff_A_Q03tJHuo7_0(.dout(w_dff_A_g6NQHAoh9_0),.din(w_dff_A_Q03tJHuo7_0),.clk(gclk));
	jdff dff_A_zS251Rh04_0(.dout(w_dff_A_Q03tJHuo7_0),.din(w_dff_A_zS251Rh04_0),.clk(gclk));
	jdff dff_A_eAuW7okS4_0(.dout(w_dff_A_zS251Rh04_0),.din(w_dff_A_eAuW7okS4_0),.clk(gclk));
	jdff dff_A_PAAYFXB99_0(.dout(w_dff_A_eAuW7okS4_0),.din(w_dff_A_PAAYFXB99_0),.clk(gclk));
	jdff dff_A_ryEwEkan5_0(.dout(w_dff_A_PAAYFXB99_0),.din(w_dff_A_ryEwEkan5_0),.clk(gclk));
	jdff dff_A_dmHWo8dH3_1(.dout(w_G143_0[1]),.din(w_dff_A_dmHWo8dH3_1),.clk(gclk));
	jdff dff_A_1Zt6HHmR4_0(.dout(w_G128_0[0]),.din(w_dff_A_1Zt6HHmR4_0),.clk(gclk));
	jdff dff_A_2OvaMXge7_0(.dout(w_dff_A_1Zt6HHmR4_0),.din(w_dff_A_2OvaMXge7_0),.clk(gclk));
	jdff dff_A_hHsEpiOP6_0(.dout(w_dff_A_2OvaMXge7_0),.din(w_dff_A_hHsEpiOP6_0),.clk(gclk));
	jdff dff_A_naPrRy4H7_0(.dout(w_dff_A_hHsEpiOP6_0),.din(w_dff_A_naPrRy4H7_0),.clk(gclk));
	jdff dff_A_6RwbPwZM9_0(.dout(w_dff_A_naPrRy4H7_0),.din(w_dff_A_6RwbPwZM9_0),.clk(gclk));
	jdff dff_A_fnWTvjgw0_0(.dout(w_dff_A_6RwbPwZM9_0),.din(w_dff_A_fnWTvjgw0_0),.clk(gclk));
	jdff dff_A_oszF1gkS2_0(.dout(w_dff_A_fnWTvjgw0_0),.din(w_dff_A_oszF1gkS2_0),.clk(gclk));
	jdff dff_A_lEWY4w7D6_0(.dout(w_dff_A_oszF1gkS2_0),.din(w_dff_A_lEWY4w7D6_0),.clk(gclk));
	jdff dff_A_bpc1Pi4f8_0(.dout(w_dff_A_lEWY4w7D6_0),.din(w_dff_A_bpc1Pi4f8_0),.clk(gclk));
	jdff dff_A_4U4Dn5B10_0(.dout(w_dff_A_bpc1Pi4f8_0),.din(w_dff_A_4U4Dn5B10_0),.clk(gclk));
	jdff dff_A_7dghcLrw1_0(.dout(w_dff_A_4U4Dn5B10_0),.din(w_dff_A_7dghcLrw1_0),.clk(gclk));
	jdff dff_A_4MXdOiW35_0(.dout(w_G134_0[0]),.din(w_dff_A_4MXdOiW35_0),.clk(gclk));
	jdff dff_A_699554VJ5_0(.dout(w_dff_A_4MXdOiW35_0),.din(w_dff_A_699554VJ5_0),.clk(gclk));
	jdff dff_A_WciAu2Qa8_0(.dout(w_dff_A_699554VJ5_0),.din(w_dff_A_WciAu2Qa8_0),.clk(gclk));
	jdff dff_A_N7BOy3hJ9_0(.dout(w_dff_A_WciAu2Qa8_0),.din(w_dff_A_N7BOy3hJ9_0),.clk(gclk));
	jdff dff_A_3mtpfrEd9_0(.dout(w_dff_A_N7BOy3hJ9_0),.din(w_dff_A_3mtpfrEd9_0),.clk(gclk));
	jdff dff_A_INH41D6U6_0(.dout(w_dff_A_3mtpfrEd9_0),.din(w_dff_A_INH41D6U6_0),.clk(gclk));
	jdff dff_A_PzPKDana9_0(.dout(w_dff_A_INH41D6U6_0),.din(w_dff_A_PzPKDana9_0),.clk(gclk));
	jdff dff_A_ZO63gEjH1_0(.dout(w_dff_A_PzPKDana9_0),.din(w_dff_A_ZO63gEjH1_0),.clk(gclk));
	jdff dff_A_rnKEsWx37_0(.dout(w_dff_A_ZO63gEjH1_0),.din(w_dff_A_rnKEsWx37_0),.clk(gclk));
	jdff dff_A_NDNan9j49_0(.dout(w_dff_A_rnKEsWx37_0),.din(w_dff_A_NDNan9j49_0),.clk(gclk));
	jdff dff_A_7gLeVlQI2_0(.dout(w_dff_A_NDNan9j49_0),.din(w_dff_A_7gLeVlQI2_0),.clk(gclk));
	jdff dff_A_XcRayItl7_1(.dout(w_G134_0[1]),.din(w_dff_A_XcRayItl7_1),.clk(gclk));
	jdff dff_A_i9Og0RTD8_0(.dout(w_n58_0[0]),.din(w_dff_A_i9Og0RTD8_0),.clk(gclk));
	jdff dff_A_yEqPEles3_0(.dout(w_dff_A_i9Og0RTD8_0),.din(w_dff_A_yEqPEles3_0),.clk(gclk));
	jdff dff_A_cVYZLGLT9_0(.dout(w_dff_A_yEqPEles3_0),.din(w_dff_A_cVYZLGLT9_0),.clk(gclk));
	jdff dff_A_lPlN46Zi2_0(.dout(w_dff_A_cVYZLGLT9_0),.din(w_dff_A_lPlN46Zi2_0),.clk(gclk));
	jdff dff_A_rA1iVUIV8_2(.dout(w_n58_0[2]),.din(w_dff_A_rA1iVUIV8_2),.clk(gclk));
	jdff dff_A_lqjD7w6a1_2(.dout(w_dff_A_rA1iVUIV8_2),.din(w_dff_A_lqjD7w6a1_2),.clk(gclk));
	jdff dff_A_6vZRGKSU4_2(.dout(w_dff_A_lqjD7w6a1_2),.din(w_dff_A_6vZRGKSU4_2),.clk(gclk));
	jdff dff_A_z0LuLn477_2(.dout(w_dff_A_6vZRGKSU4_2),.din(w_dff_A_z0LuLn477_2),.clk(gclk));
	jdff dff_A_1yJTqHgw8_0(.dout(w_G902_3[0]),.din(w_dff_A_1yJTqHgw8_0),.clk(gclk));
	jdff dff_A_ekZdutAZ2_0(.dout(w_dff_A_1yJTqHgw8_0),.din(w_dff_A_ekZdutAZ2_0),.clk(gclk));
	jdff dff_A_v6I2KH7f2_0(.dout(w_G478_0[0]),.din(w_dff_A_v6I2KH7f2_0),.clk(gclk));
	jdff dff_A_JzvUZGg29_0(.dout(w_dff_A_v6I2KH7f2_0),.din(w_dff_A_JzvUZGg29_0),.clk(gclk));
	jdff dff_A_azIfX3Y38_0(.dout(w_dff_A_JzvUZGg29_0),.din(w_dff_A_azIfX3Y38_0),.clk(gclk));
	jdff dff_A_DmcJJByz4_0(.dout(w_dff_A_azIfX3Y38_0),.din(w_dff_A_DmcJJByz4_0),.clk(gclk));
	jdff dff_A_DQ4NMHGq0_0(.dout(w_dff_A_DmcJJByz4_0),.din(w_dff_A_DQ4NMHGq0_0),.clk(gclk));
	jdff dff_A_g7pf2V5u6_0(.dout(w_dff_A_DQ4NMHGq0_0),.din(w_dff_A_g7pf2V5u6_0),.clk(gclk));
	jdff dff_A_po0E5KME4_0(.dout(w_dff_A_g7pf2V5u6_0),.din(w_dff_A_po0E5KME4_0),.clk(gclk));
	jdff dff_A_sSABVEBM1_0(.dout(w_dff_A_po0E5KME4_0),.din(w_dff_A_sSABVEBM1_0),.clk(gclk));
	jdff dff_A_wSa2KBbh5_0(.dout(w_dff_A_sSABVEBM1_0),.din(w_dff_A_wSa2KBbh5_0),.clk(gclk));
	jdff dff_A_UwQepUMf0_0(.dout(w_dff_A_wSa2KBbh5_0),.din(w_dff_A_UwQepUMf0_0),.clk(gclk));
	jdff dff_A_zjJnu9ml6_0(.dout(w_dff_A_UwQepUMf0_0),.din(w_dff_A_zjJnu9ml6_0),.clk(gclk));
	jdff dff_A_53XppaRC8_0(.dout(w_dff_A_zjJnu9ml6_0),.din(w_dff_A_53XppaRC8_0),.clk(gclk));
	jdff dff_A_N1vGFIui8_0(.dout(w_dff_A_53XppaRC8_0),.din(w_dff_A_N1vGFIui8_0),.clk(gclk));
	jdff dff_A_A3mIpxqX5_0(.dout(w_dff_A_N1vGFIui8_0),.din(w_dff_A_A3mIpxqX5_0),.clk(gclk));
	jdff dff_A_Pb6hprQj1_0(.dout(w_dff_A_A3mIpxqX5_0),.din(w_dff_A_Pb6hprQj1_0),.clk(gclk));
	jdff dff_A_H4EUOxXu5_0(.dout(w_dff_A_Pb6hprQj1_0),.din(w_dff_A_H4EUOxXu5_0),.clk(gclk));
	jdff dff_A_z11SiYkI1_1(.dout(w_G478_0[1]),.din(w_dff_A_z11SiYkI1_1),.clk(gclk));
	jdff dff_A_u17sdarp3_1(.dout(w_dff_A_z11SiYkI1_1),.din(w_dff_A_u17sdarp3_1),.clk(gclk));
	jdff dff_A_uejkKqTt8_1(.dout(w_dff_A_u17sdarp3_1),.din(w_dff_A_uejkKqTt8_1),.clk(gclk));
	jdff dff_A_ErbHBAEZ7_1(.dout(w_dff_A_uejkKqTt8_1),.din(w_dff_A_ErbHBAEZ7_1),.clk(gclk));
	jdff dff_A_EBDUmzyk5_1(.dout(w_dff_A_ErbHBAEZ7_1),.din(w_dff_A_EBDUmzyk5_1),.clk(gclk));
	jdff dff_A_bF80AltB1_1(.dout(w_dff_A_EBDUmzyk5_1),.din(w_dff_A_bF80AltB1_1),.clk(gclk));
	jdff dff_A_apHLc5GV3_1(.dout(w_n265_0[1]),.din(w_dff_A_apHLc5GV3_1),.clk(gclk));
	jdff dff_B_FkmzQT5x0_3(.din(n265),.dout(w_dff_B_FkmzQT5x0_3),.clk(gclk));
	jdff dff_B_sdL8uqzI8_3(.din(w_dff_B_FkmzQT5x0_3),.dout(w_dff_B_sdL8uqzI8_3),.clk(gclk));
	jdff dff_B_glo3kX217_3(.din(w_dff_B_sdL8uqzI8_3),.dout(w_dff_B_glo3kX217_3),.clk(gclk));
	jdff dff_B_jqo5RMfB2_3(.din(w_dff_B_glo3kX217_3),.dout(w_dff_B_jqo5RMfB2_3),.clk(gclk));
	jdff dff_B_3i79ASGC1_3(.din(w_dff_B_jqo5RMfB2_3),.dout(w_dff_B_3i79ASGC1_3),.clk(gclk));
	jdff dff_B_orduQgoF1_3(.din(w_dff_B_3i79ASGC1_3),.dout(w_dff_B_orduQgoF1_3),.clk(gclk));
	jdff dff_B_mKTavY603_3(.din(w_dff_B_orduQgoF1_3),.dout(w_dff_B_mKTavY603_3),.clk(gclk));
	jdff dff_B_YiyA7Xno4_3(.din(w_dff_B_mKTavY603_3),.dout(w_dff_B_YiyA7Xno4_3),.clk(gclk));
	jdff dff_B_JwMiTnx43_3(.din(w_dff_B_YiyA7Xno4_3),.dout(w_dff_B_JwMiTnx43_3),.clk(gclk));
	jdff dff_B_5oOo1v0z3_3(.din(w_dff_B_JwMiTnx43_3),.dout(w_dff_B_5oOo1v0z3_3),.clk(gclk));
	jdff dff_B_JDfv641l3_3(.din(w_dff_B_5oOo1v0z3_3),.dout(w_dff_B_JDfv641l3_3),.clk(gclk));
	jdff dff_B_ZOBIZjc95_3(.din(w_dff_B_JDfv641l3_3),.dout(w_dff_B_ZOBIZjc95_3),.clk(gclk));
	jdff dff_B_aM2RjltO6_3(.din(w_dff_B_ZOBIZjc95_3),.dout(w_dff_B_aM2RjltO6_3),.clk(gclk));
	jdff dff_B_QKUuJj6k5_3(.din(w_dff_B_aM2RjltO6_3),.dout(w_dff_B_QKUuJj6k5_3),.clk(gclk));
	jdff dff_B_PhKd6gim7_3(.din(w_dff_B_QKUuJj6k5_3),.dout(w_dff_B_PhKd6gim7_3),.clk(gclk));
	jdff dff_B_ABthXCsD1_3(.din(w_dff_B_PhKd6gim7_3),.dout(w_dff_B_ABthXCsD1_3),.clk(gclk));
	jdff dff_A_zpocZClW1_0(.dout(w_G953_1[0]),.din(w_dff_A_zpocZClW1_0),.clk(gclk));
	jdff dff_A_kzb2hd9g2_0(.dout(w_dff_A_zpocZClW1_0),.din(w_dff_A_kzb2hd9g2_0),.clk(gclk));
	jdff dff_A_tPvQ50N17_0(.dout(w_dff_A_kzb2hd9g2_0),.din(w_dff_A_tPvQ50N17_0),.clk(gclk));
	jdff dff_A_0iwGuBup5_0(.dout(w_dff_A_tPvQ50N17_0),.din(w_dff_A_0iwGuBup5_0),.clk(gclk));
	jdff dff_A_1JkvPatN8_0(.dout(w_dff_A_0iwGuBup5_0),.din(w_dff_A_1JkvPatN8_0),.clk(gclk));
	jdff dff_A_dnb0bL5J6_0(.dout(w_dff_A_1JkvPatN8_0),.din(w_dff_A_dnb0bL5J6_0),.clk(gclk));
	jdff dff_A_noxCN2xs0_0(.dout(w_dff_A_dnb0bL5J6_0),.din(w_dff_A_noxCN2xs0_0),.clk(gclk));
	jdff dff_A_cmziJ8rH0_0(.dout(w_dff_A_noxCN2xs0_0),.din(w_dff_A_cmziJ8rH0_0),.clk(gclk));
	jdff dff_A_PTOOPFEP7_0(.dout(w_dff_A_cmziJ8rH0_0),.din(w_dff_A_PTOOPFEP7_0),.clk(gclk));
	jdff dff_A_5uLjN7M02_0(.dout(w_dff_A_PTOOPFEP7_0),.din(w_dff_A_5uLjN7M02_0),.clk(gclk));
	jdff dff_A_U89RAlI01_0(.dout(w_dff_A_5uLjN7M02_0),.din(w_dff_A_U89RAlI01_0),.clk(gclk));
	jdff dff_A_jZCOVcyN5_0(.dout(w_dff_A_U89RAlI01_0),.din(w_dff_A_jZCOVcyN5_0),.clk(gclk));
	jdff dff_A_EUiMTc6g9_0(.dout(w_dff_A_jZCOVcyN5_0),.din(w_dff_A_EUiMTc6g9_0),.clk(gclk));
	jdff dff_A_3qGi0CTf2_0(.dout(w_dff_A_EUiMTc6g9_0),.din(w_dff_A_3qGi0CTf2_0),.clk(gclk));
	jdff dff_A_j20f81iP6_0(.dout(w_dff_A_3qGi0CTf2_0),.din(w_dff_A_j20f81iP6_0),.clk(gclk));
	jdff dff_A_dsLaRl0i4_1(.dout(w_G953_1[1]),.din(w_dff_A_dsLaRl0i4_1),.clk(gclk));
	jdff dff_A_JPs7umaD0_1(.dout(w_dff_A_dsLaRl0i4_1),.din(w_dff_A_JPs7umaD0_1),.clk(gclk));
	jdff dff_A_QPQ4pMGT8_1(.dout(w_dff_A_JPs7umaD0_1),.din(w_dff_A_QPQ4pMGT8_1),.clk(gclk));
	jdff dff_A_boM86YGm1_1(.dout(w_dff_A_QPQ4pMGT8_1),.din(w_dff_A_boM86YGm1_1),.clk(gclk));
	jdff dff_A_essMvL466_1(.dout(w_dff_A_boM86YGm1_1),.din(w_dff_A_essMvL466_1),.clk(gclk));
	jdff dff_A_TMAstcUh7_1(.dout(w_dff_A_essMvL466_1),.din(w_dff_A_TMAstcUh7_1),.clk(gclk));
	jdff dff_A_NAHX9de54_1(.dout(w_dff_A_TMAstcUh7_1),.din(w_dff_A_NAHX9de54_1),.clk(gclk));
	jdff dff_A_Bi0O1SEm3_1(.dout(w_dff_A_NAHX9de54_1),.din(w_dff_A_Bi0O1SEm3_1),.clk(gclk));
	jdff dff_A_kyiRyx2l1_1(.dout(w_dff_A_Bi0O1SEm3_1),.din(w_dff_A_kyiRyx2l1_1),.clk(gclk));
	jdff dff_A_BVOeA0sq0_1(.dout(w_dff_A_kyiRyx2l1_1),.din(w_dff_A_BVOeA0sq0_1),.clk(gclk));
	jdff dff_A_wUT6urke0_1(.dout(w_dff_A_BVOeA0sq0_1),.din(w_dff_A_wUT6urke0_1),.clk(gclk));
	jdff dff_A_6Rsph3Hg4_1(.dout(w_dff_A_wUT6urke0_1),.din(w_dff_A_6Rsph3Hg4_1),.clk(gclk));
	jdff dff_A_8MQaLwTx7_2(.dout(w_G953_0[2]),.din(w_dff_A_8MQaLwTx7_2),.clk(gclk));
	jdff dff_A_bbIVZ2GE6_2(.dout(w_dff_A_8MQaLwTx7_2),.din(w_dff_A_bbIVZ2GE6_2),.clk(gclk));
	jdff dff_A_BLAfd50W6_2(.dout(w_dff_A_bbIVZ2GE6_2),.din(w_dff_A_BLAfd50W6_2),.clk(gclk));
	jdff dff_A_6a1B3lW21_2(.dout(w_dff_A_BLAfd50W6_2),.din(w_dff_A_6a1B3lW21_2),.clk(gclk));
	jdff dff_A_lF46ez6K4_2(.dout(w_dff_A_6a1B3lW21_2),.din(w_dff_A_lF46ez6K4_2),.clk(gclk));
	jdff dff_A_CtgLOVyt6_2(.dout(w_dff_A_lF46ez6K4_2),.din(w_dff_A_CtgLOVyt6_2),.clk(gclk));
	jdff dff_A_NVQNUgLU8_2(.dout(w_dff_A_CtgLOVyt6_2),.din(w_dff_A_NVQNUgLU8_2),.clk(gclk));
	jdff dff_A_41mZbeXE9_2(.dout(w_dff_A_NVQNUgLU8_2),.din(w_dff_A_41mZbeXE9_2),.clk(gclk));
	jdff dff_A_i8Bpewt29_2(.dout(w_dff_A_41mZbeXE9_2),.din(w_dff_A_i8Bpewt29_2),.clk(gclk));
	jdff dff_A_KObVYEQX8_2(.dout(w_dff_A_i8Bpewt29_2),.din(w_dff_A_KObVYEQX8_2),.clk(gclk));
	jdff dff_A_QKLFT9Vj5_2(.dout(w_dff_A_KObVYEQX8_2),.din(w_dff_A_QKLFT9Vj5_2),.clk(gclk));
	jdff dff_A_9q7KrHWp5_2(.dout(w_dff_A_QKLFT9Vj5_2),.din(w_dff_A_9q7KrHWp5_2),.clk(gclk));
	jdff dff_A_lFjUfkaK7_2(.dout(w_dff_A_9q7KrHWp5_2),.din(w_dff_A_lFjUfkaK7_2),.clk(gclk));
	jdff dff_A_BnUQP51w1_2(.dout(w_dff_A_lFjUfkaK7_2),.din(w_dff_A_BnUQP51w1_2),.clk(gclk));
	jdff dff_A_TcigiV841_2(.dout(w_dff_A_BnUQP51w1_2),.din(w_dff_A_TcigiV841_2),.clk(gclk));
	jdff dff_A_eJ8WeTly5_1(.dout(w_G952_0[1]),.din(w_dff_A_eJ8WeTly5_1),.clk(gclk));
	jdff dff_A_kB4SSVFo8_1(.dout(w_dff_A_eJ8WeTly5_1),.din(w_dff_A_kB4SSVFo8_1),.clk(gclk));
	jdff dff_A_q5XNO7724_1(.dout(w_dff_A_kB4SSVFo8_1),.din(w_dff_A_q5XNO7724_1),.clk(gclk));
	jdff dff_A_KbNwem6D8_1(.dout(w_dff_A_q5XNO7724_1),.din(w_dff_A_KbNwem6D8_1),.clk(gclk));
	jdff dff_A_Bcs8i3FC8_1(.dout(w_dff_A_KbNwem6D8_1),.din(w_dff_A_Bcs8i3FC8_1),.clk(gclk));
	jdff dff_A_L04gicix8_1(.dout(w_dff_A_Bcs8i3FC8_1),.din(w_dff_A_L04gicix8_1),.clk(gclk));
	jdff dff_A_oxWsyVxS3_1(.dout(w_dff_A_L04gicix8_1),.din(w_dff_A_oxWsyVxS3_1),.clk(gclk));
	jdff dff_A_rBR9K8g67_1(.dout(w_dff_A_oxWsyVxS3_1),.din(w_dff_A_rBR9K8g67_1),.clk(gclk));
	jdff dff_A_PE3lYjSi0_1(.dout(w_dff_A_rBR9K8g67_1),.din(w_dff_A_PE3lYjSi0_1),.clk(gclk));
	jdff dff_A_DNaSOExD5_1(.dout(w_dff_A_PE3lYjSi0_1),.din(w_dff_A_DNaSOExD5_1),.clk(gclk));
	jdff dff_A_lqCeg8BL0_1(.dout(w_dff_A_DNaSOExD5_1),.din(w_dff_A_lqCeg8BL0_1),.clk(gclk));
	jdff dff_A_56Wg1G6r6_1(.dout(w_dff_A_lqCeg8BL0_1),.din(w_dff_A_56Wg1G6r6_1),.clk(gclk));
	jdff dff_A_dI8Hm2Kf7_1(.dout(w_dff_A_56Wg1G6r6_1),.din(w_dff_A_dI8Hm2Kf7_1),.clk(gclk));
	jdff dff_A_xR0wmvLR0_1(.dout(w_dff_A_dI8Hm2Kf7_1),.din(w_dff_A_xR0wmvLR0_1),.clk(gclk));
	jdff dff_A_Y3lDFskQ4_1(.dout(w_dff_A_xR0wmvLR0_1),.din(w_dff_A_Y3lDFskQ4_1),.clk(gclk));
	jdff dff_A_fyg1Pvi90_1(.dout(w_dff_A_Y3lDFskQ4_1),.din(w_dff_A_fyg1Pvi90_1),.clk(gclk));
	jdff dff_A_9rtk9RnC4_2(.dout(w_G952_0[2]),.din(w_dff_A_9rtk9RnC4_2),.clk(gclk));
	jdff dff_B_rfC0uYMu3_3(.din(G952),.dout(w_dff_B_rfC0uYMu3_3),.clk(gclk));
	jdff dff_A_MwqRsx0w6_2(.dout(w_dff_A_SMnVsTUa9_0),.din(w_dff_A_MwqRsx0w6_2),.clk(gclk));
	jdff dff_A_SMnVsTUa9_0(.dout(w_dff_A_fve125FU0_0),.din(w_dff_A_SMnVsTUa9_0),.clk(gclk));
	jdff dff_A_fve125FU0_0(.dout(w_dff_A_OQIf7Pgw2_0),.din(w_dff_A_fve125FU0_0),.clk(gclk));
	jdff dff_A_OQIf7Pgw2_0(.dout(w_dff_A_dpkeVIAL3_0),.din(w_dff_A_OQIf7Pgw2_0),.clk(gclk));
	jdff dff_A_dpkeVIAL3_0(.dout(w_dff_A_GI9QouZV0_0),.din(w_dff_A_dpkeVIAL3_0),.clk(gclk));
	jdff dff_A_GI9QouZV0_0(.dout(w_dff_A_ujBRfDho2_0),.din(w_dff_A_GI9QouZV0_0),.clk(gclk));
	jdff dff_A_ujBRfDho2_0(.dout(w_dff_A_bHBPXyAM6_0),.din(w_dff_A_ujBRfDho2_0),.clk(gclk));
	jdff dff_A_bHBPXyAM6_0(.dout(G3),.din(w_dff_A_bHBPXyAM6_0),.clk(gclk));
	jdff dff_A_y0S1Air87_2(.dout(w_dff_A_XU688eYr5_0),.din(w_dff_A_y0S1Air87_2),.clk(gclk));
	jdff dff_A_XU688eYr5_0(.dout(w_dff_A_8USHUJhp6_0),.din(w_dff_A_XU688eYr5_0),.clk(gclk));
	jdff dff_A_8USHUJhp6_0(.dout(w_dff_A_987J6CRB3_0),.din(w_dff_A_8USHUJhp6_0),.clk(gclk));
	jdff dff_A_987J6CRB3_0(.dout(w_dff_A_Eq74QE4D7_0),.din(w_dff_A_987J6CRB3_0),.clk(gclk));
	jdff dff_A_Eq74QE4D7_0(.dout(w_dff_A_KyyL9Txj4_0),.din(w_dff_A_Eq74QE4D7_0),.clk(gclk));
	jdff dff_A_KyyL9Txj4_0(.dout(w_dff_A_0YMYoiDk5_0),.din(w_dff_A_KyyL9Txj4_0),.clk(gclk));
	jdff dff_A_0YMYoiDk5_0(.dout(w_dff_A_d4RSwXSv6_0),.din(w_dff_A_0YMYoiDk5_0),.clk(gclk));
	jdff dff_A_d4RSwXSv6_0(.dout(G6),.din(w_dff_A_d4RSwXSv6_0),.clk(gclk));
	jdff dff_A_N02qW1yA7_2(.dout(w_dff_A_EiKuOHs69_0),.din(w_dff_A_N02qW1yA7_2),.clk(gclk));
	jdff dff_A_EiKuOHs69_0(.dout(w_dff_A_k0UDo0I42_0),.din(w_dff_A_EiKuOHs69_0),.clk(gclk));
	jdff dff_A_k0UDo0I42_0(.dout(w_dff_A_e86XZncz6_0),.din(w_dff_A_k0UDo0I42_0),.clk(gclk));
	jdff dff_A_e86XZncz6_0(.dout(w_dff_A_he6nAg600_0),.din(w_dff_A_e86XZncz6_0),.clk(gclk));
	jdff dff_A_he6nAg600_0(.dout(w_dff_A_UtqTR2KL3_0),.din(w_dff_A_he6nAg600_0),.clk(gclk));
	jdff dff_A_UtqTR2KL3_0(.dout(w_dff_A_6uNN18sl4_0),.din(w_dff_A_UtqTR2KL3_0),.clk(gclk));
	jdff dff_A_6uNN18sl4_0(.dout(w_dff_A_TRxK1wIw3_0),.din(w_dff_A_6uNN18sl4_0),.clk(gclk));
	jdff dff_A_TRxK1wIw3_0(.dout(G9),.din(w_dff_A_TRxK1wIw3_0),.clk(gclk));
	jdff dff_A_DlpRYtCa6_2(.dout(w_dff_A_HEvIMrhO8_0),.din(w_dff_A_DlpRYtCa6_2),.clk(gclk));
	jdff dff_A_HEvIMrhO8_0(.dout(w_dff_A_z5QkHR330_0),.din(w_dff_A_HEvIMrhO8_0),.clk(gclk));
	jdff dff_A_z5QkHR330_0(.dout(w_dff_A_BWrBfszh5_0),.din(w_dff_A_z5QkHR330_0),.clk(gclk));
	jdff dff_A_BWrBfszh5_0(.dout(w_dff_A_7arxUe0W1_0),.din(w_dff_A_BWrBfszh5_0),.clk(gclk));
	jdff dff_A_7arxUe0W1_0(.dout(w_dff_A_1vEWcUA41_0),.din(w_dff_A_7arxUe0W1_0),.clk(gclk));
	jdff dff_A_1vEWcUA41_0(.dout(w_dff_A_odBtbIM31_0),.din(w_dff_A_1vEWcUA41_0),.clk(gclk));
	jdff dff_A_odBtbIM31_0(.dout(w_dff_A_q9vckpvG5_0),.din(w_dff_A_odBtbIM31_0),.clk(gclk));
	jdff dff_A_q9vckpvG5_0(.dout(G12),.din(w_dff_A_q9vckpvG5_0),.clk(gclk));
	jdff dff_A_apRAkZg53_2(.dout(w_dff_A_uHEe57WI6_0),.din(w_dff_A_apRAkZg53_2),.clk(gclk));
	jdff dff_A_uHEe57WI6_0(.dout(w_dff_A_FBgM1fRJ7_0),.din(w_dff_A_uHEe57WI6_0),.clk(gclk));
	jdff dff_A_FBgM1fRJ7_0(.dout(w_dff_A_W1YKKNVp8_0),.din(w_dff_A_FBgM1fRJ7_0),.clk(gclk));
	jdff dff_A_W1YKKNVp8_0(.dout(w_dff_A_46LN5FKU6_0),.din(w_dff_A_W1YKKNVp8_0),.clk(gclk));
	jdff dff_A_46LN5FKU6_0(.dout(w_dff_A_L0YRChQu4_0),.din(w_dff_A_46LN5FKU6_0),.clk(gclk));
	jdff dff_A_L0YRChQu4_0(.dout(w_dff_A_7jMzdGF19_0),.din(w_dff_A_L0YRChQu4_0),.clk(gclk));
	jdff dff_A_7jMzdGF19_0(.dout(w_dff_A_APq4wjnn3_0),.din(w_dff_A_7jMzdGF19_0),.clk(gclk));
	jdff dff_A_APq4wjnn3_0(.dout(G30),.din(w_dff_A_APq4wjnn3_0),.clk(gclk));
	jdff dff_A_R0NrbBNi0_2(.dout(w_dff_A_0CGTH1bS1_0),.din(w_dff_A_R0NrbBNi0_2),.clk(gclk));
	jdff dff_A_0CGTH1bS1_0(.dout(w_dff_A_MiuQvP6e8_0),.din(w_dff_A_0CGTH1bS1_0),.clk(gclk));
	jdff dff_A_MiuQvP6e8_0(.dout(w_dff_A_Z6zVLBMN3_0),.din(w_dff_A_MiuQvP6e8_0),.clk(gclk));
	jdff dff_A_Z6zVLBMN3_0(.dout(w_dff_A_zV37IviQ9_0),.din(w_dff_A_Z6zVLBMN3_0),.clk(gclk));
	jdff dff_A_zV37IviQ9_0(.dout(w_dff_A_XCrhnlh61_0),.din(w_dff_A_zV37IviQ9_0),.clk(gclk));
	jdff dff_A_XCrhnlh61_0(.dout(w_dff_A_srCUVw1T3_0),.din(w_dff_A_XCrhnlh61_0),.clk(gclk));
	jdff dff_A_srCUVw1T3_0(.dout(w_dff_A_BhoUwC8V8_0),.din(w_dff_A_srCUVw1T3_0),.clk(gclk));
	jdff dff_A_BhoUwC8V8_0(.dout(G45),.din(w_dff_A_BhoUwC8V8_0),.clk(gclk));
	jdff dff_A_CDdRnRdY1_2(.dout(w_dff_A_TwZMTknQ6_0),.din(w_dff_A_CDdRnRdY1_2),.clk(gclk));
	jdff dff_A_TwZMTknQ6_0(.dout(w_dff_A_r50859xe3_0),.din(w_dff_A_TwZMTknQ6_0),.clk(gclk));
	jdff dff_A_r50859xe3_0(.dout(w_dff_A_duzyz5qb1_0),.din(w_dff_A_r50859xe3_0),.clk(gclk));
	jdff dff_A_duzyz5qb1_0(.dout(w_dff_A_Y4lLNQqh1_0),.din(w_dff_A_duzyz5qb1_0),.clk(gclk));
	jdff dff_A_Y4lLNQqh1_0(.dout(w_dff_A_KXNZUKy93_0),.din(w_dff_A_Y4lLNQqh1_0),.clk(gclk));
	jdff dff_A_KXNZUKy93_0(.dout(w_dff_A_rH4t5jcW6_0),.din(w_dff_A_KXNZUKy93_0),.clk(gclk));
	jdff dff_A_rH4t5jcW6_0(.dout(w_dff_A_B8RMUIgp3_0),.din(w_dff_A_rH4t5jcW6_0),.clk(gclk));
	jdff dff_A_B8RMUIgp3_0(.dout(G48),.din(w_dff_A_B8RMUIgp3_0),.clk(gclk));
	jdff dff_A_E06fr8vG6_2(.dout(w_dff_A_sXNTBL0W1_0),.din(w_dff_A_E06fr8vG6_2),.clk(gclk));
	jdff dff_A_sXNTBL0W1_0(.dout(w_dff_A_jQHsaafC8_0),.din(w_dff_A_sXNTBL0W1_0),.clk(gclk));
	jdff dff_A_jQHsaafC8_0(.dout(w_dff_A_sjmTYC5l1_0),.din(w_dff_A_jQHsaafC8_0),.clk(gclk));
	jdff dff_A_sjmTYC5l1_0(.dout(w_dff_A_Zuo1Q2Tg7_0),.din(w_dff_A_sjmTYC5l1_0),.clk(gclk));
	jdff dff_A_Zuo1Q2Tg7_0(.dout(w_dff_A_8IxNtXV07_0),.din(w_dff_A_Zuo1Q2Tg7_0),.clk(gclk));
	jdff dff_A_8IxNtXV07_0(.dout(w_dff_A_pXdMvCaZ5_0),.din(w_dff_A_8IxNtXV07_0),.clk(gclk));
	jdff dff_A_pXdMvCaZ5_0(.dout(w_dff_A_rSjKCHNd3_0),.din(w_dff_A_pXdMvCaZ5_0),.clk(gclk));
	jdff dff_A_rSjKCHNd3_0(.dout(G15),.din(w_dff_A_rSjKCHNd3_0),.clk(gclk));
	jdff dff_A_YMIk41gS8_2(.dout(w_dff_A_4MA2UY1h2_0),.din(w_dff_A_YMIk41gS8_2),.clk(gclk));
	jdff dff_A_4MA2UY1h2_0(.dout(w_dff_A_DzfdTRno5_0),.din(w_dff_A_4MA2UY1h2_0),.clk(gclk));
	jdff dff_A_DzfdTRno5_0(.dout(w_dff_A_3gpJ598J6_0),.din(w_dff_A_DzfdTRno5_0),.clk(gclk));
	jdff dff_A_3gpJ598J6_0(.dout(w_dff_A_5a5NmolD0_0),.din(w_dff_A_3gpJ598J6_0),.clk(gclk));
	jdff dff_A_5a5NmolD0_0(.dout(w_dff_A_LNaBgbuO0_0),.din(w_dff_A_5a5NmolD0_0),.clk(gclk));
	jdff dff_A_LNaBgbuO0_0(.dout(w_dff_A_KptFUmx34_0),.din(w_dff_A_LNaBgbuO0_0),.clk(gclk));
	jdff dff_A_KptFUmx34_0(.dout(w_dff_A_YLO0uwsg6_0),.din(w_dff_A_KptFUmx34_0),.clk(gclk));
	jdff dff_A_YLO0uwsg6_0(.dout(G18),.din(w_dff_A_YLO0uwsg6_0),.clk(gclk));
	jdff dff_A_s8rXBoX56_2(.dout(w_dff_A_ZZdXydGm6_0),.din(w_dff_A_s8rXBoX56_2),.clk(gclk));
	jdff dff_A_ZZdXydGm6_0(.dout(w_dff_A_QqLKm64w6_0),.din(w_dff_A_ZZdXydGm6_0),.clk(gclk));
	jdff dff_A_QqLKm64w6_0(.dout(w_dff_A_eJCCopJa8_0),.din(w_dff_A_QqLKm64w6_0),.clk(gclk));
	jdff dff_A_eJCCopJa8_0(.dout(w_dff_A_z5WKZ6gX1_0),.din(w_dff_A_eJCCopJa8_0),.clk(gclk));
	jdff dff_A_z5WKZ6gX1_0(.dout(w_dff_A_QfYmXPBM9_0),.din(w_dff_A_z5WKZ6gX1_0),.clk(gclk));
	jdff dff_A_QfYmXPBM9_0(.dout(w_dff_A_dVTLmbqY8_0),.din(w_dff_A_QfYmXPBM9_0),.clk(gclk));
	jdff dff_A_dVTLmbqY8_0(.dout(w_dff_A_Woh6OdVs2_0),.din(w_dff_A_dVTLmbqY8_0),.clk(gclk));
	jdff dff_A_Woh6OdVs2_0(.dout(G21),.din(w_dff_A_Woh6OdVs2_0),.clk(gclk));
	jdff dff_A_48L5gWb59_2(.dout(w_dff_A_pFBbqCNZ4_0),.din(w_dff_A_48L5gWb59_2),.clk(gclk));
	jdff dff_A_pFBbqCNZ4_0(.dout(w_dff_A_FEyCJMKm5_0),.din(w_dff_A_pFBbqCNZ4_0),.clk(gclk));
	jdff dff_A_FEyCJMKm5_0(.dout(w_dff_A_KoVzu7q37_0),.din(w_dff_A_FEyCJMKm5_0),.clk(gclk));
	jdff dff_A_KoVzu7q37_0(.dout(w_dff_A_O11JJmVx6_0),.din(w_dff_A_KoVzu7q37_0),.clk(gclk));
	jdff dff_A_O11JJmVx6_0(.dout(w_dff_A_65Oxlssu0_0),.din(w_dff_A_O11JJmVx6_0),.clk(gclk));
	jdff dff_A_65Oxlssu0_0(.dout(w_dff_A_fvL8DYi59_0),.din(w_dff_A_65Oxlssu0_0),.clk(gclk));
	jdff dff_A_fvL8DYi59_0(.dout(G24),.din(w_dff_A_fvL8DYi59_0),.clk(gclk));
	jdff dff_A_ve0cAdrm6_2(.dout(w_dff_A_RkFR6puO5_0),.din(w_dff_A_ve0cAdrm6_2),.clk(gclk));
	jdff dff_A_RkFR6puO5_0(.dout(w_dff_A_hrAlhNAm1_0),.din(w_dff_A_RkFR6puO5_0),.clk(gclk));
	jdff dff_A_hrAlhNAm1_0(.dout(w_dff_A_5WpE3FLY3_0),.din(w_dff_A_hrAlhNAm1_0),.clk(gclk));
	jdff dff_A_5WpE3FLY3_0(.dout(w_dff_A_q0ckrtDo0_0),.din(w_dff_A_5WpE3FLY3_0),.clk(gclk));
	jdff dff_A_q0ckrtDo0_0(.dout(w_dff_A_jaUi27hL0_0),.din(w_dff_A_q0ckrtDo0_0),.clk(gclk));
	jdff dff_A_jaUi27hL0_0(.dout(w_dff_A_3exUiFpL3_0),.din(w_dff_A_jaUi27hL0_0),.clk(gclk));
	jdff dff_A_3exUiFpL3_0(.dout(w_dff_A_UjaTMIZF1_0),.din(w_dff_A_3exUiFpL3_0),.clk(gclk));
	jdff dff_A_UjaTMIZF1_0(.dout(G27),.din(w_dff_A_UjaTMIZF1_0),.clk(gclk));
	jdff dff_A_pvSnXxJb3_2(.dout(w_dff_A_BURVCN1F8_0),.din(w_dff_A_pvSnXxJb3_2),.clk(gclk));
	jdff dff_A_BURVCN1F8_0(.dout(w_dff_A_4AI7CPcV2_0),.din(w_dff_A_BURVCN1F8_0),.clk(gclk));
	jdff dff_A_4AI7CPcV2_0(.dout(w_dff_A_cFslUK5m3_0),.din(w_dff_A_4AI7CPcV2_0),.clk(gclk));
	jdff dff_A_cFslUK5m3_0(.dout(w_dff_A_bnlqfMaz2_0),.din(w_dff_A_cFslUK5m3_0),.clk(gclk));
	jdff dff_A_bnlqfMaz2_0(.dout(w_dff_A_66F1CsVM0_0),.din(w_dff_A_bnlqfMaz2_0),.clk(gclk));
	jdff dff_A_66F1CsVM0_0(.dout(w_dff_A_iY3FJa145_0),.din(w_dff_A_66F1CsVM0_0),.clk(gclk));
	jdff dff_A_iY3FJa145_0(.dout(w_dff_A_2uHjnuT57_0),.din(w_dff_A_iY3FJa145_0),.clk(gclk));
	jdff dff_A_2uHjnuT57_0(.dout(G33),.din(w_dff_A_2uHjnuT57_0),.clk(gclk));
	jdff dff_A_9hMXUQKg7_2(.dout(w_dff_A_uOSfjerm5_0),.din(w_dff_A_9hMXUQKg7_2),.clk(gclk));
	jdff dff_A_uOSfjerm5_0(.dout(w_dff_A_S2Tp7smu0_0),.din(w_dff_A_uOSfjerm5_0),.clk(gclk));
	jdff dff_A_S2Tp7smu0_0(.dout(w_dff_A_HinQTAFs2_0),.din(w_dff_A_S2Tp7smu0_0),.clk(gclk));
	jdff dff_A_HinQTAFs2_0(.dout(w_dff_A_WZS4Vqqr7_0),.din(w_dff_A_HinQTAFs2_0),.clk(gclk));
	jdff dff_A_WZS4Vqqr7_0(.dout(w_dff_A_8KdmLDuJ5_0),.din(w_dff_A_WZS4Vqqr7_0),.clk(gclk));
	jdff dff_A_8KdmLDuJ5_0(.dout(w_dff_A_6hExMG0z6_0),.din(w_dff_A_8KdmLDuJ5_0),.clk(gclk));
	jdff dff_A_6hExMG0z6_0(.dout(w_dff_A_9S8T0T9S2_0),.din(w_dff_A_6hExMG0z6_0),.clk(gclk));
	jdff dff_A_9S8T0T9S2_0(.dout(G36),.din(w_dff_A_9S8T0T9S2_0),.clk(gclk));
	jdff dff_A_H0wbY1Ub8_2(.dout(w_dff_A_5Bs10Pmm9_0),.din(w_dff_A_H0wbY1Ub8_2),.clk(gclk));
	jdff dff_A_5Bs10Pmm9_0(.dout(w_dff_A_xevfPlMV8_0),.din(w_dff_A_5Bs10Pmm9_0),.clk(gclk));
	jdff dff_A_xevfPlMV8_0(.dout(w_dff_A_gCTlPJdx7_0),.din(w_dff_A_xevfPlMV8_0),.clk(gclk));
	jdff dff_A_gCTlPJdx7_0(.dout(w_dff_A_pQ3YMCOW1_0),.din(w_dff_A_gCTlPJdx7_0),.clk(gclk));
	jdff dff_A_pQ3YMCOW1_0(.dout(w_dff_A_s3ze39kW7_0),.din(w_dff_A_pQ3YMCOW1_0),.clk(gclk));
	jdff dff_A_s3ze39kW7_0(.dout(w_dff_A_yvSMQFQ96_0),.din(w_dff_A_s3ze39kW7_0),.clk(gclk));
	jdff dff_A_yvSMQFQ96_0(.dout(w_dff_A_qGGumymi0_0),.din(w_dff_A_yvSMQFQ96_0),.clk(gclk));
	jdff dff_A_qGGumymi0_0(.dout(G39),.din(w_dff_A_qGGumymi0_0),.clk(gclk));
	jdff dff_A_K9N8MOyh8_2(.dout(w_dff_A_vxdStgLY0_0),.din(w_dff_A_K9N8MOyh8_2),.clk(gclk));
	jdff dff_A_vxdStgLY0_0(.dout(w_dff_A_gIDHvzis8_0),.din(w_dff_A_vxdStgLY0_0),.clk(gclk));
	jdff dff_A_gIDHvzis8_0(.dout(w_dff_A_gAgSSfCd1_0),.din(w_dff_A_gIDHvzis8_0),.clk(gclk));
	jdff dff_A_gAgSSfCd1_0(.dout(w_dff_A_C5lsZQZP3_0),.din(w_dff_A_gAgSSfCd1_0),.clk(gclk));
	jdff dff_A_C5lsZQZP3_0(.dout(w_dff_A_KIFz7CH72_0),.din(w_dff_A_C5lsZQZP3_0),.clk(gclk));
	jdff dff_A_KIFz7CH72_0(.dout(w_dff_A_tGRE1uAg3_0),.din(w_dff_A_KIFz7CH72_0),.clk(gclk));
	jdff dff_A_tGRE1uAg3_0(.dout(w_dff_A_ADq0GnWf3_0),.din(w_dff_A_tGRE1uAg3_0),.clk(gclk));
	jdff dff_A_ADq0GnWf3_0(.dout(G42),.din(w_dff_A_ADq0GnWf3_0),.clk(gclk));
	jdff dff_A_NWXt4Snf1_2(.dout(G75),.din(w_dff_A_NWXt4Snf1_2),.clk(gclk));
	jdff dff_A_jrsgWhlw6_2(.dout(w_dff_A_FggnYhHZ2_0),.din(w_dff_A_jrsgWhlw6_2),.clk(gclk));
	jdff dff_A_FggnYhHZ2_0(.dout(G69),.din(w_dff_A_FggnYhHZ2_0),.clk(gclk));
	jdff dff_A_bfIBpwvT2_2(.dout(w_dff_A_Xaaac5Zg9_0),.din(w_dff_A_bfIBpwvT2_2),.clk(gclk));
	jdff dff_A_Xaaac5Zg9_0(.dout(G72),.din(w_dff_A_Xaaac5Zg9_0),.clk(gclk));
	jdff dff_A_CR8MmAXU9_2(.dout(G57),.din(w_dff_A_CR8MmAXU9_2),.clk(gclk));
endmodule

