module rf_c1355(G233gat, G228gat, G229gat, G227gat, G218gat, G211gat, G197gat, G50gat, G64gat, G43gat, G232gat, G22gat, G36gat, G127gat, G29gat, G78gat, G230gat, G15gat, G8gat, G71gat, G120gat, G226gat, G162gat, G85gat, G57gat, G92gat, G1gat, G190gat, G148gat, G99gat, G155gat, G106gat, G225gat, G113gat, G134gat, G141gat, G204gat, G169gat, G176gat, G231gat, G183gat, G1353gat, G1355gat, G1335gat, G1338gat, G1334gat, G1332gat, G1340gat, G1354gat, G1331gat, G1329gat, G1350gat, G1352gat, G1328gat, G1327gat, G1336gat, G1326gat, G1341gat, G1344gat, G1333gat, G1325gat, G1343gat, G1330gat, G1339gat, G1337gat, G1342gat, G1324gat, G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1351gat);
    input G233gat, G228gat, G229gat, G227gat, G218gat, G211gat, G197gat, G50gat, G64gat, G43gat, G232gat, G22gat, G36gat, G127gat, G29gat, G78gat, G230gat, G15gat, G8gat, G71gat, G120gat, G226gat, G162gat, G85gat, G57gat, G92gat, G1gat, G190gat, G148gat, G99gat, G155gat, G106gat, G225gat, G113gat, G134gat, G141gat, G204gat, G169gat, G176gat, G231gat, G183gat;
    output G1353gat, G1355gat, G1335gat, G1338gat, G1334gat, G1332gat, G1340gat, G1354gat, G1331gat, G1329gat, G1350gat, G1352gat, G1328gat, G1327gat, G1336gat, G1326gat, G1341gat, G1344gat, G1333gat, G1325gat, G1343gat, G1330gat, G1339gat, G1337gat, G1342gat, G1324gat, G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1351gat;
    wire n76;
    wire n80;
    wire n84;
    wire n88;
    wire n92;
    wire n96;
    wire n100;
    wire n104;
    wire n108;
    wire n112;
    wire n116;
    wire n120;
    wire n124;
    wire n127;
    wire n130;
    wire n134;
    wire n138;
    wire n142;
    wire n145;
    wire n149;
    wire n153;
    wire n157;
    wire n161;
    wire n165;
    wire n169;
    wire n173;
    wire n177;
    wire n181;
    wire n185;
    wire n189;
    wire n193;
    wire n197;
    wire n201;
    wire n204;
    wire n208;
    wire n212;
    wire n216;
    wire n220;
    wire n224;
    wire n228;
    wire n232;
    wire n235;
    wire n239;
    wire n243;
    wire n247;
    wire n251;
    wire n255;
    wire n259;
    wire n263;
    wire n267;
    wire n271;
    wire n275;
    wire n279;
    wire n283;
    wire n287;
    wire n291;
    wire n295;
    wire n299;
    wire n303;
    wire n307;
    wire n311;
    wire n315;
    wire n319;
    wire n323;
    wire n327;
    wire n331;
    wire n335;
    wire n339;
    wire n342;
    wire n346;
    wire n350;
    wire n354;
    wire n358;
    wire n362;
    wire n366;
    wire n370;
    wire n374;
    wire n378;
    wire n382;
    wire n386;
    wire n390;
    wire n394;
    wire n398;
    wire n401;
    wire n405;
    wire n409;
    wire n413;
    wire n417;
    wire n421;
    wire n425;
    wire n429;
    wire n433;
    wire n437;
    wire n441;
    wire n445;
    wire n449;
    wire n453;
    wire n457;
    wire n461;
    wire n465;
    wire n469;
    wire n473;
    wire n481;
    wire n485;
    wire n489;
    wire n493;
    wire n501;
    wire n505;
    wire n509;
    wire n513;
    wire n521;
    wire n525;
    wire n529;
    wire n533;
    wire n541;
    wire n545;
    wire n549;
    wire n552;
    wire n556;
    wire n560;
    wire n564;
    wire n568;
    wire n572;
    wire n576;
    wire n580;
    wire n588;
    wire n596;
    wire n604;
    wire n611;
    wire n615;
    wire n619;
    wire n623;
    wire n627;
    wire n631;
    wire n635;
    wire n639;
    wire n643;
    wire n647;
    wire n651;
    wire n659;
    wire n667;
    wire n675;
    wire n683;
    wire n687;
    wire n691;
    wire n699;
    wire n707;
    wire n715;
    wire n723;
    wire n727;
    wire n731;
    wire n735;
    wire n739;
    wire n743;
    wire n747;
    wire n751;
    wire n755;
    wire n759;
    wire n763;
    wire n767;
    wire n775;
    wire n783;
    wire n791;
    wire n799;
    wire n803;
    wire n807;
    wire n811;
    wire n819;
    wire n827;
    wire n835;
    wire n843;
    wire n847;
    wire n851;
    wire n855;
    wire n863;
    wire n871;
    wire n879;
    wire n887;
    wire n891;
    wire n895;
    wire n903;
    wire n911;
    wire n919;
    wire n1359;
    wire n1362;
    wire n1365;
    wire n1368;
    wire n1371;
    wire n1373;
    wire n1376;
    wire n1379;
    wire n1382;
    wire n1385;
    wire n1388;
    wire n1391;
    wire n1394;
    wire n1397;
    wire n1400;
    wire n1403;
    wire n1406;
    wire n1409;
    wire n1412;
    wire n1415;
    wire n1418;
    wire n1421;
    wire n1424;
    wire n1427;
    wire n1430;
    wire n1433;
    wire n1436;
    wire n1439;
    wire n1442;
    wire n1446;
    wire n1448;
    wire n1451;
    wire n1454;
    wire n1457;
    wire n1460;
    wire n1463;
    wire n1466;
    wire n1469;
    wire n1473;
    wire n1475;
    wire n1478;
    wire n1481;
    wire n1484;
    wire n1487;
    wire n1490;
    wire n1493;
    wire n1496;
    wire n1500;
    wire n1502;
    wire n1505;
    wire n1508;
    wire n1511;
    wire n1514;
    wire n1517;
    wire n1520;
    wire n1523;
    wire n1527;
    wire n1529;
    wire n1532;
    wire n1535;
    wire n1538;
    wire n1541;
    wire n1544;
    wire n1547;
    wire n1550;
    wire n1554;
    wire n1556;
    wire n1559;
    wire n1562;
    wire n1565;
    wire n1568;
    wire n1571;
    wire n1574;
    wire n1577;
    wire n1581;
    wire n1583;
    wire n1586;
    wire n1589;
    wire n1592;
    wire n1595;
    wire n1598;
    wire n1601;
    wire n1604;
    wire n1608;
    wire n1611;
    wire n1613;
    wire n1616;
    wire n1619;
    wire n1622;
    wire n1625;
    wire n1628;
    wire n1631;
    wire n1634;
    wire n1638;
    wire n1640;
    wire n1643;
    wire n1646;
    wire n1649;
    wire n1652;
    wire n1655;
    wire n1658;
    wire n1661;
    wire n1665;
    wire n1667;
    wire n1670;
    wire n1673;
    wire n1676;
    wire n1679;
    wire n1682;
    wire n1685;
    wire n1688;
    wire n1691;
    wire n1694;
    wire n1697;
    wire n1700;
    wire n1703;
    wire n1706;
    wire n1709;
    wire n1712;
    wire n1715;
    wire n1718;
    wire n1721;
    wire n1724;
    wire n1727;
    wire n1730;
    wire n1733;
    wire n1736;
    wire n1739;
    wire n1742;
    wire n1745;
    wire n1748;
    wire n1751;
    wire n1754;
    wire n1757;
    wire n1760;
    wire n1763;
    wire n1766;
    wire n1769;
    wire n1772;
    wire n1775;
    wire n1778;
    wire n1781;
    wire n1784;
    wire n1787;
    wire n1790;
    wire n1793;
    wire n1796;
    wire n1799;
    wire n1802;
    wire n1805;
    wire n1808;
    wire n1811;
    wire n1814;
    wire n1817;
    wire n1820;
    wire n1823;
    wire n1826;
    wire n1829;
    wire n1832;
    wire n1835;
    wire n1838;
    wire n1841;
    wire n1844;
    wire n1847;
    wire n1850;
    wire n1853;
    wire n1856;
    wire n1859;
    wire n1862;
    wire n1865;
    wire n1868;
    wire n1871;
    wire n1874;
    wire n1877;
    wire n1880;
    wire n1883;
    wire n1886;
    wire n1889;
    wire n1892;
    wire n1895;
    wire n1898;
    wire n1901;
    wire n1904;
    wire n1907;
    wire n1910;
    wire n1913;
    wire n1916;
    wire n1919;
    wire n1922;
    wire n1925;
    wire n1928;
    wire n1931;
    wire n1934;
    wire n1937;
    wire n1940;
    wire n1943;
    wire n1946;
    wire n1949;
    wire n1952;
    wire n1955;
    wire n1958;
    wire n1961;
    wire n1964;
    wire n1967;
    wire n1970;
    wire n1973;
    wire n1976;
    wire n1979;
    wire n1982;
    wire n1985;
    wire n1988;
    wire n1991;
    wire n1994;
    wire n1997;
    wire n2000;
    wire n2003;
    wire n2006;
    wire n2009;
    wire n2012;
    wire n2015;
    wire n2018;
    wire n2021;
    wire n2024;
    wire n2027;
    wire n2030;
    wire n2033;
    wire n2036;
    wire n2039;
    wire n2042;
    wire n2045;
    wire n2048;
    wire n2051;
    wire n2054;
    wire n2057;
    wire n2060;
    wire n2063;
    wire n2066;
    wire n2069;
    wire n2072;
    wire n2075;
    wire n2078;
    wire n2081;
    wire n2084;
    wire n2087;
    wire n2090;
    wire n2093;
    wire n2096;
    wire n2099;
    wire n2102;
    wire n2105;
    wire n2108;
    wire n2111;
    wire n2114;
    wire n2117;
    wire n2120;
    wire n2123;
    wire n2126;
    wire n2129;
    wire n2132;
    wire n2135;
    wire n2138;
    wire n2141;
    wire n2144;
    wire n2147;
    wire n2150;
    wire n2153;
    wire n2156;
    wire n2159;
    wire n2162;
    wire n2165;
    wire n2168;
    wire n2171;
    wire n2174;
    wire n2177;
    wire n2180;
    wire n2183;
    wire n2186;
    wire n2189;
    wire n2192;
    wire n2195;
    wire n2198;
    wire n2201;
    wire n2204;
    wire n2207;
    wire n2210;
    wire n2213;
    wire n2216;
    wire n2219;
    wire n2222;
    wire n2225;
    wire n2228;
    wire n2231;
    wire n2234;
    wire n2237;
    wire n2240;
    wire n2243;
    wire n2246;
    wire n2249;
    wire n2252;
    wire n2255;
    wire n2258;
    wire n2261;
    wire n2264;
    wire n2267;
    wire n2270;
    wire n2273;
    wire n2276;
    wire n2279;
    wire n2282;
    wire n2285;
    wire n2288;
    wire n2291;
    wire n2294;
    wire n2297;
    wire n2300;
    wire n2303;
    wire n2306;
    wire n2309;
    wire n2312;
    wire n2315;
    wire n2318;
    wire n2321;
    wire n2324;
    wire n2327;
    wire n2330;
    wire n2333;
    wire n2336;
    wire n2339;
    wire n2342;
    wire n2345;
    wire n2348;
    wire n2351;
    wire n2354;
    wire n2357;
    wire n2360;
    wire n2363;
    wire n2366;
    wire n2369;
    wire n2372;
    wire n2375;
    wire n2378;
    wire n2381;
    wire n2384;
    wire n2387;
    wire n2390;
    wire n2393;
    wire n2396;
    wire n2399;
    wire n2402;
    wire n2405;
    wire n2408;
    wire n2411;
    wire n2414;
    wire n2417;
    wire n2420;
    wire n2423;
    wire n2426;
    wire n2429;
    wire n2432;
    wire n2435;
    wire n2438;
    wire n2441;
    wire n2444;
    wire n2448;
    wire n2450;
    wire n2453;
    wire n2456;
    wire n2459;
    wire n2462;
    wire n2465;
    wire n2468;
    wire n2471;
    wire n2474;
    wire n2477;
    wire n2480;
    wire n2483;
    wire n2486;
    wire n2489;
    wire n2492;
    wire n2495;
    wire n2498;
    wire n2501;
    wire n2504;
    wire n2507;
    wire n2510;
    wire n2513;
    wire n2516;
    wire n2519;
    wire n2522;
    wire n2525;
    wire n2528;
    wire n2531;
    wire n2534;
    wire n2537;
    wire n2540;
    wire n2543;
    wire n2546;
    wire n2549;
    wire n2552;
    wire n2555;
    jand g000(.dinb(G225gat), .dina(G233gat), .dout(n76));
    jxor g001(.dinb(G127gat), .dina(G134gat), .dout(n80));
    jxor g002(.dinb(G113gat), .dina(G120gat), .dout(n84));
    jxor g003(.dinb(n80), .dina(n84), .dout(n88));
    jxor g004(.dinb(n1473), .dina(n88), .dout(n92));
    jxor g005(.dinb(G57gat), .dina(G85gat), .dout(n96));
    jor g006(.dinb(G1gat), .dina(G29gat), .dout(n100));
    jxor g007(.dinb(n96), .dina(n100), .dout(n104));
    jand g008(.dinb(G155gat), .dina(G162gat), .dout(n108));
    jxor g009(.dinb(G141gat), .dina(G148gat), .dout(n112));
    jxor g010(.dinb(n108), .dina(n112), .dout(n116));
    jxor g011(.dinb(n104), .dina(n116), .dout(n120));
    jxor g012(.dinb(n92), .dina(n120), .dout(n124));
    jnot g013(.din(G225gat), .dout(n127));
    jnot g014(.din(G233gat), .dout(n130));
    jor g015(.dinb(n127), .dina(n130), .dout(n134));
    jxor g016(.dinb(n134), .dina(n88), .dout(n138));
    jxor g017(.dinb(n138), .dina(n120), .dout(n142));
    jnot g018(.din(G226gat), .dout(n145));
    jor g019(.dinb(n145), .dina(n130), .dout(n149));
    jxor g020(.dinb(G211gat), .dina(G218gat), .dout(n153));
    jxor g021(.dinb(G197gat), .dina(G204gat), .dout(n157));
    jxor g022(.dinb(n153), .dina(n157), .dout(n161));
    jxor g023(.dinb(n149), .dina(n161), .dout(n165));
    jxor g024(.dinb(G183gat), .dina(G190gat), .dout(n169));
    jxor g025(.dinb(G169gat), .dina(G176gat), .dout(n173));
    jxor g026(.dinb(n169), .dina(n173), .dout(n177));
    jxor g027(.dinb(G64gat), .dina(G92gat), .dout(n181));
    jxor g028(.dinb(G8gat), .dina(G36gat), .dout(n185));
    jxor g029(.dinb(n181), .dina(n185), .dout(n189));
    jxor g030(.dinb(n177), .dina(n189), .dout(n193));
    jxor g031(.dinb(n165), .dina(n193), .dout(n197));
    jxor g032(.dinb(n142), .dina(n197), .dout(n201));
    jnot g033(.din(G227gat), .dout(n204));
    jor g034(.dinb(n204), .dina(n130), .dout(n208));
    jxor g035(.dinb(n88), .dina(n208), .dout(n212));
    jxor g036(.dinb(G71gat), .dina(G99gat), .dout(n216));
    jxor g037(.dinb(G15gat), .dina(G43gat), .dout(n220));
    jxor g038(.dinb(n216), .dina(n220), .dout(n224));
    jxor g039(.dinb(n177), .dina(n224), .dout(n228));
    jxor g040(.dinb(n212), .dina(n228), .dout(n232));
    jnot g041(.din(G228gat), .dout(n235));
    jor g042(.dinb(n235), .dina(n130), .dout(n239));
    jxor g043(.dinb(n116), .dina(n239), .dout(n243));
    jxor g044(.dinb(G78gat), .dina(G106gat), .dout(n247));
    jxor g045(.dinb(G22gat), .dina(G50gat), .dout(n251));
    jxor g046(.dinb(n247), .dina(n251), .dout(n255));
    jxor g047(.dinb(n161), .dina(n255), .dout(n259));
    jxor g048(.dinb(n243), .dina(n259), .dout(n263));
    jand g049(.dinb(n232), .dina(n263), .dout(n267));
    jand g050(.dinb(n201), .dina(n267), .dout(n271));
    jxor g051(.dinb(n232), .dina(n263), .dout(n275));
    jand g052(.dinb(n142), .dina(n197), .dout(n279));
    jand g053(.dinb(n275), .dina(n279), .dout(n283));
    jor g054(.dinb(n271), .dina(n283), .dout(n287));
    jand g055(.dinb(G229gat), .dina(G233gat), .dout(n291));
    jxor g056(.dinb(G43gat), .dina(G50gat), .dout(n295));
    jxor g057(.dinb(G29gat), .dina(G36gat), .dout(n299));
    jxor g058(.dinb(n295), .dina(n299), .dout(n303));
    jxor g059(.dinb(n1554), .dina(n303), .dout(n307));
    jxor g060(.dinb(G15gat), .dina(G22gat), .dout(n311));
    jxor g061(.dinb(G1gat), .dina(G8gat), .dout(n315));
    jxor g062(.dinb(n311), .dina(n315), .dout(n319));
    jxor g063(.dinb(G169gat), .dina(G197gat), .dout(n323));
    jxor g064(.dinb(G113gat), .dina(G141gat), .dout(n327));
    jxor g065(.dinb(n323), .dina(n327), .dout(n331));
    jxor g066(.dinb(n319), .dina(n331), .dout(n335));
    jxor g067(.dinb(n307), .dina(n335), .dout(n339));
    jnot g068(.din(G230gat), .dout(n342));
    jor g069(.dinb(n342), .dina(n130), .dout(n346));
    jxor g070(.dinb(G99gat), .dina(G106gat), .dout(n350));
    jxor g071(.dinb(G85gat), .dina(G92gat), .dout(n354));
    jxor g072(.dinb(n350), .dina(n354), .dout(n358));
    jxor g073(.dinb(n346), .dina(n358), .dout(n362));
    jxor g074(.dinb(G71gat), .dina(G78gat), .dout(n366));
    jxor g075(.dinb(G57gat), .dina(G64gat), .dout(n370));
    jxor g076(.dinb(n366), .dina(n370), .dout(n374));
    jxor g077(.dinb(G176gat), .dina(G204gat), .dout(n378));
    jxor g078(.dinb(G120gat), .dina(G148gat), .dout(n382));
    jxor g079(.dinb(n378), .dina(n382), .dout(n386));
    jxor g080(.dinb(n374), .dina(n386), .dout(n390));
    jxor g081(.dinb(n362), .dina(n390), .dout(n394));
    jand g082(.dinb(n339), .dina(n394), .dout(n398));
    jnot g083(.din(G232gat), .dout(n401));
    jor g084(.dinb(n401), .dina(n130), .dout(n405));
    jxor g085(.dinb(n303), .dina(n405), .dout(n409));
    jxor g086(.dinb(G190gat), .dina(G218gat), .dout(n413));
    jxor g087(.dinb(G134gat), .dina(G162gat), .dout(n417));
    jxor g088(.dinb(n413), .dina(n417), .dout(n421));
    jxor g089(.dinb(n358), .dina(n421), .dout(n425));
    jxor g090(.dinb(n409), .dina(n425), .dout(n429));
    jand g091(.dinb(G231gat), .dina(G233gat), .dout(n433));
    jxor g092(.dinb(n319), .dina(n1608), .dout(n437));
    jxor g093(.dinb(G183gat), .dina(G211gat), .dout(n441));
    jxor g094(.dinb(G127gat), .dina(G155gat), .dout(n445));
    jxor g095(.dinb(n441), .dina(n445), .dout(n449));
    jxor g096(.dinb(n374), .dina(n449), .dout(n453));
    jxor g097(.dinb(n437), .dina(n453), .dout(n457));
    jand g098(.dinb(n429), .dina(n457), .dout(n461));
    jand g099(.dinb(n398), .dina(n461), .dout(n465));
    jand g100(.dinb(n287), .dina(n1359), .dout(n469));
    jand g101(.dinb(n1448), .dina(n469), .dout(n473));
    jxor g102(.dinb(n2126), .dina(n473), .dout(G1324gat));
    jand g103(.dinb(G226gat), .dina(G233gat), .dout(n481));
    jxor g104(.dinb(n1665), .dina(n161), .dout(n485));
    jxor g105(.dinb(n485), .dina(n193), .dout(n489));
    jand g106(.dinb(n1640), .dina(n469), .dout(n493));
    jxor g107(.dinb(n2099), .dina(n493), .dout(G1325gat));
    jand g108(.dinb(G227gat), .dina(G233gat), .dout(n501));
    jxor g109(.dinb(n88), .dina(n1527), .dout(n505));
    jxor g110(.dinb(n505), .dina(n228), .dout(n509));
    jand g111(.dinb(n1502), .dina(n469), .dout(n513));
    jxor g112(.dinb(n2180), .dina(n513), .dout(G1326gat));
    jand g113(.dinb(G228gat), .dina(G233gat), .dout(n521));
    jxor g114(.dinb(n116), .dina(n1638), .dout(n525));
    jxor g115(.dinb(n525), .dina(n259), .dout(n529));
    jand g116(.dinb(n1613), .dina(n469), .dout(n533));
    jxor g117(.dinb(n2153), .dina(n533), .dout(G1327gat));
    jand g118(.dinb(G232gat), .dina(G233gat), .dout(n541));
    jxor g119(.dinb(n303), .dina(n2448), .dout(n545));
    jxor g120(.dinb(n545), .dina(n425), .dout(n549));
    jnot g121(.din(G231gat), .dout(n552));
    jor g122(.dinb(n552), .dina(n130), .dout(n556));
    jxor g123(.dinb(n319), .dina(n556), .dout(n560));
    jxor g124(.dinb(n560), .dina(n453), .dout(n564));
    jand g125(.dinb(n549), .dina(n564), .dout(n568));
    jand g126(.dinb(n398), .dina(n568), .dout(n572));
    jand g127(.dinb(n287), .dina(n1362), .dout(n576));
    jand g128(.dinb(n1448), .dina(n576), .dout(n580));
    jxor g129(.dinb(n2477), .dina(n580), .dout(G1328gat));
    jand g130(.dinb(n1640), .dina(n576), .dout(n588));
    jxor g131(.dinb(n2450), .dina(n588), .dout(G1329gat));
    jand g132(.dinb(n1502), .dina(n576), .dout(n596));
    jxor g133(.dinb(n2531), .dina(n596), .dout(G1330gat));
    jand g134(.dinb(n1613), .dina(n576), .dout(n604));
    jxor g135(.dinb(n2504), .dina(n604), .dout(G1331gat));
    jnot g136(.din(G229gat), .dout(n611));
    jor g137(.dinb(n611), .dina(n130), .dout(n615));
    jxor g138(.dinb(n615), .dina(n303), .dout(n619));
    jxor g139(.dinb(n619), .dina(n335), .dout(n623));
    jand g140(.dinb(G230gat), .dina(G233gat), .dout(n627));
    jxor g141(.dinb(n1581), .dina(n358), .dout(n631));
    jxor g142(.dinb(n631), .dina(n390), .dout(n635));
    jand g143(.dinb(n623), .dina(n635), .dout(n639));
    jand g144(.dinb(n461), .dina(n639), .dout(n643));
    jand g145(.dinb(n287), .dina(n1365), .dout(n647));
    jand g146(.dinb(n1448), .dina(n647), .dout(n651));
    jxor g147(.dinb(n1910), .dina(n651), .dout(G1332gat));
    jand g148(.dinb(n1640), .dina(n647), .dout(n659));
    jxor g149(.dinb(n1883), .dina(n659), .dout(G1333gat));
    jand g150(.dinb(n1502), .dina(n647), .dout(n667));
    jxor g151(.dinb(n1964), .dina(n667), .dout(G1334gat));
    jand g152(.dinb(n1613), .dina(n647), .dout(n675));
    jxor g153(.dinb(n1937), .dina(n675), .dout(G1335gat));
    jand g154(.dinb(n568), .dina(n639), .dout(n683));
    jand g155(.dinb(n287), .dina(n1368), .dout(n687));
    jand g156(.dinb(n1460), .dina(n687), .dout(n691));
    jxor g157(.dinb(n2366), .dina(n691), .dout(G1336gat));
    jand g158(.dinb(n1652), .dina(n687), .dout(n699));
    jxor g159(.dinb(n2339), .dina(n699), .dout(G1337gat));
    jand g160(.dinb(n1514), .dina(n687), .dout(n707));
    jxor g161(.dinb(n2420), .dina(n707), .dout(G1338gat));
    jand g162(.dinb(n1625), .dina(n687), .dout(n715));
    jxor g163(.dinb(n2393), .dina(n715), .dout(G1339gat));
    jxor g164(.dinb(n623), .dina(n394), .dout(n723));
    jand g165(.dinb(n429), .dina(n564), .dout(n727));
    jand g166(.dinb(n723), .dina(n727), .dout(n731));
    jxor g167(.dinb(n429), .dina(n564), .dout(n735));
    jand g168(.dinb(n623), .dina(n394), .dout(n739));
    jand g169(.dinb(n735), .dina(n739), .dout(n743));
    jor g170(.dinb(n731), .dina(n743), .dout(n747));
    jand g171(.dinb(n124), .dina(n197), .dout(n751));
    jand g172(.dinb(n509), .dina(n263), .dout(n755));
    jand g173(.dinb(n751), .dina(n755), .dout(n759));
    jand g174(.dinb(n747), .dina(n1371), .dout(n763));
    jand g175(.dinb(n1385), .dina(n763), .dout(n767));
    jxor g176(.dinb(n2018), .dina(n767), .dout(G1340gat));
    jand g177(.dinb(n1409), .dina(n763), .dout(n775));
    jxor g178(.dinb(n1802), .dina(n775), .dout(G1341gat));
    jand g179(.dinb(n1433), .dina(n763), .dout(n783));
    jxor g180(.dinb(n1694), .dina(n783), .dout(G1342gat));
    jand g181(.dinb(n1487), .dina(n763), .dout(n791));
    jxor g182(.dinb(n2258), .dina(n791), .dout(G1343gat));
    jand g183(.dinb(n232), .dina(n529), .dout(n799));
    jand g184(.dinb(n751), .dina(n799), .dout(n803));
    jand g185(.dinb(n747), .dina(n1446), .dout(n807));
    jand g186(.dinb(n1373), .dina(n807), .dout(n811));
    jxor g187(.dinb(n1991), .dina(n811), .dout(G1344gat));
    jand g188(.dinb(n1397), .dina(n807), .dout(n819));
    jxor g189(.dinb(n1775), .dina(n819), .dout(G1345gat));
    jand g190(.dinb(n1421), .dina(n807), .dout(n827));
    jxor g191(.dinb(n1667), .dina(n827), .dout(G1346gat));
    jand g192(.dinb(n1475), .dina(n807), .dout(n835));
    jxor g193(.dinb(n2231), .dina(n835), .dout(G1347gat));
    jand g194(.dinb(n142), .dina(n489), .dout(n843));
    jand g195(.dinb(n843), .dina(n755), .dout(n847));
    jand g196(.dinb(n747), .dina(n1500), .dout(n851));
    jand g197(.dinb(n1541), .dina(n851), .dout(n855));
    jxor g198(.dinb(n2072), .dina(n855), .dout(G1348gat));
    jand g199(.dinb(n1568), .dina(n851), .dout(n863));
    jxor g200(.dinb(n1856), .dina(n863), .dout(G1349gat));
    jand g201(.dinb(n1595), .dina(n851), .dout(n871));
    jxor g202(.dinb(n1748), .dina(n871), .dout(G1350gat));
    jand g203(.dinb(n2219), .dina(n851), .dout(n879));
    jxor g204(.dinb(n2312), .dina(n879), .dout(G1351gat));
    jand g205(.dinb(n843), .dina(n799), .dout(n887));
    jand g206(.dinb(n747), .dina(n1611), .dout(n891));
    jand g207(.dinb(n1529), .dina(n891), .dout(n895));
    jxor g208(.dinb(n2045), .dina(n895), .dout(G1352gat));
    jand g209(.dinb(n1556), .dina(n891), .dout(n903));
    jxor g210(.dinb(n1829), .dina(n903), .dout(G1353gat));
    jand g211(.dinb(n1583), .dina(n891), .dout(n911));
    jxor g212(.dinb(n1721), .dina(n911), .dout(G1354gat));
    jand g213(.dinb(n2207), .dina(n891), .dout(n919));
    jxor g214(.dinb(n2285), .dina(n919), .dout(G1355gat));
    jdff dff_A_xKU3pu0v3_0(.din(G43gat), .dout(n2555));
    jdff dff_A_k8q9Th0a1_0(.din(n2555), .dout(n2552));
    jdff dff_A_NG0MN6Vm1_0(.din(n2552), .dout(n2549));
    jdff dff_A_njk4skQt3_0(.din(n2549), .dout(n2546));
    jdff dff_A_wUecCoOS2_0(.din(n2546), .dout(n2543));
    jdff dff_A_WCC0cFL53_0(.din(n2543), .dout(n2540));
    jdff dff_A_GyiHDLOW6_0(.din(n2540), .dout(n2537));
    jdff dff_A_oxvNklsq6_0(.din(n2537), .dout(n2534));
    jdff dff_A_bO9vSmLO1_0(.din(n2534), .dout(n2531));
    jdff dff_A_RR314R8Q8_0(.din(G50gat), .dout(n2528));
    jdff dff_A_KXBpupiR4_0(.din(n2528), .dout(n2525));
    jdff dff_A_Sjkfhsm35_0(.din(n2525), .dout(n2522));
    jdff dff_A_Q50Ey19F8_0(.din(n2522), .dout(n2519));
    jdff dff_A_uL8KTwu51_0(.din(n2519), .dout(n2516));
    jdff dff_A_ugiMcQxa3_0(.din(n2516), .dout(n2513));
    jdff dff_A_bWZkvBeN1_0(.din(n2513), .dout(n2510));
    jdff dff_A_W5DfZtcP4_0(.din(n2510), .dout(n2507));
    jdff dff_A_6X0t4seZ7_0(.din(n2507), .dout(n2504));
    jdff dff_A_cwe4JHis7_0(.din(G29gat), .dout(n2501));
    jdff dff_A_aJS7xFsV0_0(.din(n2501), .dout(n2498));
    jdff dff_A_REbsdzBz5_0(.din(n2498), .dout(n2495));
    jdff dff_A_XzCJWUbI6_0(.din(n2495), .dout(n2492));
    jdff dff_A_ZgAydz5F8_0(.din(n2492), .dout(n2489));
    jdff dff_A_pSgbLwqn3_0(.din(n2489), .dout(n2486));
    jdff dff_A_jzKO9Grl4_0(.din(n2486), .dout(n2483));
    jdff dff_A_3PPKnkq55_0(.din(n2483), .dout(n2480));
    jdff dff_A_FNEe5dDD9_0(.din(n2480), .dout(n2477));
    jdff dff_A_Bq3AtPiE4_0(.din(G36gat), .dout(n2474));
    jdff dff_A_h5oOH64b1_0(.din(n2474), .dout(n2471));
    jdff dff_A_yv3XfRkb9_0(.din(n2471), .dout(n2468));
    jdff dff_A_6uovOJ424_0(.din(n2468), .dout(n2465));
    jdff dff_A_Bq3wDqe37_0(.din(n2465), .dout(n2462));
    jdff dff_A_bvFep2sR9_0(.din(n2462), .dout(n2459));
    jdff dff_A_00mIk9F13_0(.din(n2459), .dout(n2456));
    jdff dff_A_thNvn5RW8_0(.din(n2456), .dout(n2453));
    jdff dff_A_INFe41zS8_0(.din(n2453), .dout(n2450));
    jdff dff_B_StKXQ8g44_0(.din(n541), .dout(n2448));
    jdff dff_A_siwNkOmM8_0(.din(G99gat), .dout(n2444));
    jdff dff_A_l2boUcIf2_0(.din(n2444), .dout(n2441));
    jdff dff_A_FeE8XdQL3_0(.din(n2441), .dout(n2438));
    jdff dff_A_zd3SEwj73_0(.din(n2438), .dout(n2435));
    jdff dff_A_ArG5ARoO2_0(.din(n2435), .dout(n2432));
    jdff dff_A_NmdLimZI7_0(.din(n2432), .dout(n2429));
    jdff dff_A_DAAtQVSC8_0(.din(n2429), .dout(n2426));
    jdff dff_A_51tWW32V1_0(.din(n2426), .dout(n2423));
    jdff dff_A_PX5r7NvP6_0(.din(n2423), .dout(n2420));
    jdff dff_A_XCfS0hx17_0(.din(G106gat), .dout(n2417));
    jdff dff_A_dynpNwfe3_0(.din(n2417), .dout(n2414));
    jdff dff_A_TToJqUYF4_0(.din(n2414), .dout(n2411));
    jdff dff_A_zyyQjeAt2_0(.din(n2411), .dout(n2408));
    jdff dff_A_I6QaefDj9_0(.din(n2408), .dout(n2405));
    jdff dff_A_crWaQ2cq3_0(.din(n2405), .dout(n2402));
    jdff dff_A_6qTPif2P2_0(.din(n2402), .dout(n2399));
    jdff dff_A_4eHixGT68_0(.din(n2399), .dout(n2396));
    jdff dff_A_buWYYn1y0_0(.din(n2396), .dout(n2393));
    jdff dff_A_qqXMUHAH8_0(.din(G85gat), .dout(n2390));
    jdff dff_A_ciyPJucu6_0(.din(n2390), .dout(n2387));
    jdff dff_A_wymk9I4W2_0(.din(n2387), .dout(n2384));
    jdff dff_A_bqDveV6s0_0(.din(n2384), .dout(n2381));
    jdff dff_A_AaJ38CYA8_0(.din(n2381), .dout(n2378));
    jdff dff_A_CV0YNSpy6_0(.din(n2378), .dout(n2375));
    jdff dff_A_VaGBzg8D2_0(.din(n2375), .dout(n2372));
    jdff dff_A_p73U7kLS5_0(.din(n2372), .dout(n2369));
    jdff dff_A_3YVO4J6d1_0(.din(n2369), .dout(n2366));
    jdff dff_A_MgJSixOf9_0(.din(G92gat), .dout(n2363));
    jdff dff_A_YkasRRmg7_0(.din(n2363), .dout(n2360));
    jdff dff_A_iL3ahK469_0(.din(n2360), .dout(n2357));
    jdff dff_A_FPizLBuH7_0(.din(n2357), .dout(n2354));
    jdff dff_A_1iZWd9NI6_0(.din(n2354), .dout(n2351));
    jdff dff_A_BG8Rh6ER2_0(.din(n2351), .dout(n2348));
    jdff dff_A_CZZsVKvS6_0(.din(n2348), .dout(n2345));
    jdff dff_A_I0nSna0o1_0(.din(n2345), .dout(n2342));
    jdff dff_A_6itGw0pn0_0(.din(n2342), .dout(n2339));
    jdff dff_A_JEIMwhQW5_0(.din(G190gat), .dout(n2336));
    jdff dff_A_7UGSi87B9_0(.din(n2336), .dout(n2333));
    jdff dff_A_PP33N4080_0(.din(n2333), .dout(n2330));
    jdff dff_A_x3gB2pjg3_0(.din(n2330), .dout(n2327));
    jdff dff_A_5KUmLTA78_0(.din(n2327), .dout(n2324));
    jdff dff_A_EOiqoOtc3_0(.din(n2324), .dout(n2321));
    jdff dff_A_51pjyUVx9_0(.din(n2321), .dout(n2318));
    jdff dff_A_cjvwhBHY6_0(.din(n2318), .dout(n2315));
    jdff dff_A_YNTF4iPM5_0(.din(n2315), .dout(n2312));
    jdff dff_A_NcLcEOHg1_0(.din(G218gat), .dout(n2309));
    jdff dff_A_mHpwGrii5_0(.din(n2309), .dout(n2306));
    jdff dff_A_QfHVVHzW6_0(.din(n2306), .dout(n2303));
    jdff dff_A_ymiFnxrf5_0(.din(n2303), .dout(n2300));
    jdff dff_A_d32iqN4p3_0(.din(n2300), .dout(n2297));
    jdff dff_A_2jYj6XY81_0(.din(n2297), .dout(n2294));
    jdff dff_A_gbnpZSMh1_0(.din(n2294), .dout(n2291));
    jdff dff_A_j6oxsm5g0_0(.din(n2291), .dout(n2288));
    jdff dff_A_Ir1Lm2ql8_0(.din(n2288), .dout(n2285));
    jdff dff_A_LV46z0Yb9_0(.din(G134gat), .dout(n2282));
    jdff dff_A_2bUGb2lA2_0(.din(n2282), .dout(n2279));
    jdff dff_A_mi8R0ghj5_0(.din(n2279), .dout(n2276));
    jdff dff_A_1EynZoWp2_0(.din(n2276), .dout(n2273));
    jdff dff_A_GiAzDwGD5_0(.din(n2273), .dout(n2270));
    jdff dff_A_Wv1kBFym4_0(.din(n2270), .dout(n2267));
    jdff dff_A_4jS374O12_0(.din(n2267), .dout(n2264));
    jdff dff_A_I8LepBhM3_0(.din(n2264), .dout(n2261));
    jdff dff_A_RwZViO987_0(.din(n2261), .dout(n2258));
    jdff dff_A_lho714g69_0(.din(G162gat), .dout(n2255));
    jdff dff_A_xcGV2w2Y5_0(.din(n2255), .dout(n2252));
    jdff dff_A_s7R9cKts4_0(.din(n2252), .dout(n2249));
    jdff dff_A_Mkmn6cWL8_0(.din(n2249), .dout(n2246));
    jdff dff_A_hej3TN7m4_0(.din(n2246), .dout(n2243));
    jdff dff_A_QNHDHS1U9_0(.din(n2243), .dout(n2240));
    jdff dff_A_kOposQS96_0(.din(n2240), .dout(n2237));
    jdff dff_A_4TBTaEsG3_0(.din(n2237), .dout(n2234));
    jdff dff_A_gKIRh3Zf0_0(.din(n2234), .dout(n2231));
    jdff dff_A_oTQfcdLk6_2(.din(n549), .dout(n2228));
    jdff dff_A_5oSzWI7y6_2(.din(n2228), .dout(n2225));
    jdff dff_A_hFRdfaKY8_2(.din(n2225), .dout(n2222));
    jdff dff_A_r2atBBmo2_2(.din(n2222), .dout(n2219));
    jdff dff_A_qCFM8bqx2_1(.din(n549), .dout(n2216));
    jdff dff_A_nQm7JGID0_1(.din(n2216), .dout(n2213));
    jdff dff_A_QnjNCbdY0_1(.din(n2213), .dout(n2210));
    jdff dff_A_bEA0MTWC3_1(.din(n2210), .dout(n2207));
    jdff dff_A_EDrBnOSe6_0(.din(G15gat), .dout(n2204));
    jdff dff_B_cmjL1Rww2_0(.din(n465), .dout(n1359));
    jdff dff_B_FPNRDUFh2_0(.din(n572), .dout(n1362));
    jdff dff_B_g286THfp9_0(.din(n643), .dout(n1365));
    jdff dff_B_UxJlklRE2_0(.din(n683), .dout(n1368));
    jdff dff_B_5k43FNqo0_0(.din(n759), .dout(n1371));
    jdff dff_A_mFUH6Rpw1_0(.din(n1376), .dout(n1373));
    jdff dff_A_R2VCqPBv8_0(.din(n1379), .dout(n1376));
    jdff dff_A_Hna1ykVl2_0(.din(n1382), .dout(n1379));
    jdff dff_A_irQBYKDz3_0(.din(n339), .dout(n1382));
    jdff dff_A_1g7kK9tK4_1(.din(n1388), .dout(n1385));
    jdff dff_A_GOLsOaNx2_1(.din(n1391), .dout(n1388));
    jdff dff_A_7OW44oJ96_1(.din(n1394), .dout(n1391));
    jdff dff_A_swWNifuW6_1(.din(n339), .dout(n1394));
    jdff dff_A_pYo6xBRK3_0(.din(n1400), .dout(n1397));
    jdff dff_A_QJCv7gtD6_0(.din(n1403), .dout(n1400));
    jdff dff_A_uyOg5jBy8_0(.din(n1406), .dout(n1403));
    jdff dff_A_f1IOPfgz3_0(.din(n635), .dout(n1406));
    jdff dff_A_hZZVpgyw8_1(.din(n1412), .dout(n1409));
    jdff dff_A_4f73fiM98_1(.din(n1415), .dout(n1412));
    jdff dff_A_eOwpWdtw9_1(.din(n1418), .dout(n1415));
    jdff dff_A_laGYUiyh0_1(.din(n635), .dout(n1418));
    jdff dff_A_d5GjNnaR7_0(.din(n1424), .dout(n1421));
    jdff dff_A_OHR8r6E66_0(.din(n1427), .dout(n1424));
    jdff dff_A_XJZadxSO5_0(.din(n1430), .dout(n1427));
    jdff dff_A_4JGmJ2Fz5_0(.din(n457), .dout(n1430));
    jdff dff_A_9xjOhnnl7_1(.din(n1436), .dout(n1433));
    jdff dff_A_aMeHXUEl5_1(.din(n1439), .dout(n1436));
    jdff dff_A_V0jtAWDO2_1(.din(n1442), .dout(n1439));
    jdff dff_A_Ec2kHaTl7_1(.din(n457), .dout(n1442));
    jdff dff_B_biXbEgPc5_0(.din(n803), .dout(n1446));
    jdff dff_A_4Lqt83Il2_0(.din(n1451), .dout(n1448));
    jdff dff_A_fgTg1Jv04_0(.din(n1454), .dout(n1451));
    jdff dff_A_ftKzKckB4_0(.din(n1457), .dout(n1454));
    jdff dff_A_6SNxPPGn7_0(.din(n124), .dout(n1457));
    jdff dff_A_XZc7wiqf7_2(.din(n1463), .dout(n1460));
    jdff dff_A_me1o9gFW1_2(.din(n1466), .dout(n1463));
    jdff dff_A_D963d9mA5_2(.din(n1469), .dout(n1466));
    jdff dff_A_165Zc2ta7_2(.din(n124), .dout(n1469));
    jdff dff_B_IF8XNhLk2_1(.din(n76), .dout(n1473));
    jdff dff_A_PAJcn9dT3_0(.din(n1478), .dout(n1475));
    jdff dff_A_VqBWrQdn8_0(.din(n1481), .dout(n1478));
    jdff dff_A_IJOxFvg19_0(.din(n1484), .dout(n1481));
    jdff dff_A_V2mDkN3h6_0(.din(n549), .dout(n1484));
    jdff dff_A_abqZqoc75_1(.din(n1490), .dout(n1487));
    jdff dff_A_QXTdGCFf7_1(.din(n1493), .dout(n1490));
    jdff dff_A_mJ5S5fFs4_1(.din(n1496), .dout(n1493));
    jdff dff_A_Njs0eFGX5_1(.din(n549), .dout(n1496));
    jdff dff_B_DRzoBFus7_0(.din(n847), .dout(n1500));
    jdff dff_A_0RhH9Glg8_0(.din(n1505), .dout(n1502));
    jdff dff_A_NtDdDYei2_0(.din(n1508), .dout(n1505));
    jdff dff_A_uc7vfJD15_0(.din(n1511), .dout(n1508));
    jdff dff_A_8EbPuqGC5_0(.din(n509), .dout(n1511));
    jdff dff_A_g66Jxffp3_2(.din(n1517), .dout(n1514));
    jdff dff_A_qeO68XPG9_2(.din(n1520), .dout(n1517));
    jdff dff_A_uYQYbwqh4_2(.din(n1523), .dout(n1520));
    jdff dff_A_QuzHPo0f3_2(.din(n509), .dout(n1523));
    jdff dff_B_1Q2qLYgP3_0(.din(n501), .dout(n1527));
    jdff dff_A_MkVLpoxD8_1(.din(n1532), .dout(n1529));
    jdff dff_A_KHjVajVe8_1(.din(n1535), .dout(n1532));
    jdff dff_A_s7my0yG65_1(.din(n1538), .dout(n1535));
    jdff dff_A_iLlv5r7Y8_1(.din(n339), .dout(n1538));
    jdff dff_A_azsF21Uc0_2(.din(n1544), .dout(n1541));
    jdff dff_A_kauzdbCg4_2(.din(n1547), .dout(n1544));
    jdff dff_A_uVEwfuyz6_2(.din(n1550), .dout(n1547));
    jdff dff_A_hX7bIuiG4_2(.din(n339), .dout(n1550));
    jdff dff_B_BRWr53yS7_1(.din(n291), .dout(n1554));
    jdff dff_A_abikw74r6_1(.din(n1559), .dout(n1556));
    jdff dff_A_giOeR9S01_1(.din(n1562), .dout(n1559));
    jdff dff_A_JOgxZ2Zw3_1(.din(n1565), .dout(n1562));
    jdff dff_A_qgAEe6qb7_1(.din(n635), .dout(n1565));
    jdff dff_A_dixTxDkx3_2(.din(n1571), .dout(n1568));
    jdff dff_A_h4xnA3OS9_2(.din(n1574), .dout(n1571));
    jdff dff_A_co56YYDn6_2(.din(n1577), .dout(n1574));
    jdff dff_A_tgLwfAf03_2(.din(n635), .dout(n1577));
    jdff dff_B_ATjNhD5D2_1(.din(n627), .dout(n1581));
    jdff dff_A_zZ7hvxAY4_1(.din(n1586), .dout(n1583));
    jdff dff_A_Pkdo9yw89_1(.din(n1589), .dout(n1586));
    jdff dff_A_DRMG70dB8_1(.din(n1592), .dout(n1589));
    jdff dff_A_77XtZlWY0_1(.din(n457), .dout(n1592));
    jdff dff_A_mnnJYR4o3_2(.din(n1598), .dout(n1595));
    jdff dff_A_GHH0v3EJ9_2(.din(n1601), .dout(n1598));
    jdff dff_A_27yxxiUe9_2(.din(n1604), .dout(n1601));
    jdff dff_A_y2eWZ3aC8_2(.din(n457), .dout(n1604));
    jdff dff_B_NgC3zm3L5_0(.din(n433), .dout(n1608));
    jdff dff_B_faDAVPS33_0(.din(n887), .dout(n1611));
    jdff dff_A_xGYgun3O5_0(.din(n1616), .dout(n1613));
    jdff dff_A_4ApfXGwl1_0(.din(n1619), .dout(n1616));
    jdff dff_A_cGPag7kS2_0(.din(n1622), .dout(n1619));
    jdff dff_A_j4t0NFdE4_0(.din(n529), .dout(n1622));
    jdff dff_A_CX6efmZS7_2(.din(n1628), .dout(n1625));
    jdff dff_A_kkqL0wvg5_2(.din(n1631), .dout(n1628));
    jdff dff_A_3Ipy0TkH3_2(.din(n1634), .dout(n1631));
    jdff dff_A_TMTY9bze9_2(.din(n529), .dout(n1634));
    jdff dff_B_OAabkUO34_0(.din(n521), .dout(n1638));
    jdff dff_A_kTHGCwjB2_0(.din(n1643), .dout(n1640));
    jdff dff_A_lkooHMxY2_0(.din(n1646), .dout(n1643));
    jdff dff_A_j5pmguDs0_0(.din(n1649), .dout(n1646));
    jdff dff_A_arhL8J0M3_0(.din(n489), .dout(n1649));
    jdff dff_A_I6id7FMa3_2(.din(n1655), .dout(n1652));
    jdff dff_A_O0U1W0oj3_2(.din(n1658), .dout(n1655));
    jdff dff_A_eEp7lKDS0_2(.din(n1661), .dout(n1658));
    jdff dff_A_vCLGyw233_2(.din(n489), .dout(n1661));
    jdff dff_B_ykS351zP7_1(.din(n481), .dout(n1665));
    jdff dff_A_qB7lAl5k2_0(.din(n1670), .dout(n1667));
    jdff dff_A_tsnQdEWQ9_0(.din(n1673), .dout(n1670));
    jdff dff_A_cFfqxeAv7_0(.din(n1676), .dout(n1673));
    jdff dff_A_u7mCIUKN7_0(.din(n1679), .dout(n1676));
    jdff dff_A_dz5SuS8y2_0(.din(n1682), .dout(n1679));
    jdff dff_A_UPFO3qpa1_0(.din(n1685), .dout(n1682));
    jdff dff_A_VLBhRVle0_0(.din(n1688), .dout(n1685));
    jdff dff_A_65Pb4O9y1_0(.din(n1691), .dout(n1688));
    jdff dff_A_hrABN8PT1_0(.din(G155gat), .dout(n1691));
    jdff dff_A_ia10qDMy8_0(.din(n1697), .dout(n1694));
    jdff dff_A_I1qe7yD00_0(.din(n1700), .dout(n1697));
    jdff dff_A_GR8ZImjs2_0(.din(n1703), .dout(n1700));
    jdff dff_A_d3SJtoYx9_0(.din(n1706), .dout(n1703));
    jdff dff_A_AMSi2Fse8_0(.din(n1709), .dout(n1706));
    jdff dff_A_0SCVanTb8_0(.din(n1712), .dout(n1709));
    jdff dff_A_h25C699D6_0(.din(n1715), .dout(n1712));
    jdff dff_A_yfelzNNV0_0(.din(n1718), .dout(n1715));
    jdff dff_A_HRsRVT7z0_0(.din(G127gat), .dout(n1718));
    jdff dff_A_Rwg9vdXE4_0(.din(n1724), .dout(n1721));
    jdff dff_A_FLD0SfPU1_0(.din(n1727), .dout(n1724));
    jdff dff_A_gWhaXPon8_0(.din(n1730), .dout(n1727));
    jdff dff_A_A1GjUc319_0(.din(n1733), .dout(n1730));
    jdff dff_A_eJutMtdA0_0(.din(n1736), .dout(n1733));
    jdff dff_A_fCKJJ77p3_0(.din(n1739), .dout(n1736));
    jdff dff_A_k34smKwz7_0(.din(n1742), .dout(n1739));
    jdff dff_A_qVcmDyjW5_0(.din(n1745), .dout(n1742));
    jdff dff_A_sMB2Q1pA1_0(.din(G211gat), .dout(n1745));
    jdff dff_A_hoTNidvU7_0(.din(n1751), .dout(n1748));
    jdff dff_A_QzYBpNtl1_0(.din(n1754), .dout(n1751));
    jdff dff_A_0l1LUUss6_0(.din(n1757), .dout(n1754));
    jdff dff_A_JffkO1Z07_0(.din(n1760), .dout(n1757));
    jdff dff_A_6dUhSxgR2_0(.din(n1763), .dout(n1760));
    jdff dff_A_C0UBPp7y8_0(.din(n1766), .dout(n1763));
    jdff dff_A_GFdCUhbD9_0(.din(n1769), .dout(n1766));
    jdff dff_A_QC7lxjzY3_0(.din(n1772), .dout(n1769));
    jdff dff_A_rwdRgPLU9_0(.din(G183gat), .dout(n1772));
    jdff dff_A_TaFhftHr7_0(.din(n1778), .dout(n1775));
    jdff dff_A_9mZ0uv9w9_0(.din(n1781), .dout(n1778));
    jdff dff_A_m2yuHWNk7_0(.din(n1784), .dout(n1781));
    jdff dff_A_gyFTaN8y4_0(.din(n1787), .dout(n1784));
    jdff dff_A_CenpC3O09_0(.din(n1790), .dout(n1787));
    jdff dff_A_zi6lMKHg1_0(.din(n1793), .dout(n1790));
    jdff dff_A_WXyU9Cws3_0(.din(n1796), .dout(n1793));
    jdff dff_A_2wjB0cfK8_0(.din(n1799), .dout(n1796));
    jdff dff_A_knIyEPFb6_0(.din(G148gat), .dout(n1799));
    jdff dff_A_XQ32GqAF1_0(.din(n1805), .dout(n1802));
    jdff dff_A_mpAFsUDW8_0(.din(n1808), .dout(n1805));
    jdff dff_A_AK6hX0HS7_0(.din(n1811), .dout(n1808));
    jdff dff_A_1Terjt2j4_0(.din(n1814), .dout(n1811));
    jdff dff_A_4lJPUN5r6_0(.din(n1817), .dout(n1814));
    jdff dff_A_RSIRMd1s2_0(.din(n1820), .dout(n1817));
    jdff dff_A_pExwET6e6_0(.din(n1823), .dout(n1820));
    jdff dff_A_4MrzNXl71_0(.din(n1826), .dout(n1823));
    jdff dff_A_y2e0MzwA2_0(.din(G120gat), .dout(n1826));
    jdff dff_A_2NQ25OFG8_0(.din(n1832), .dout(n1829));
    jdff dff_A_7zQreJSQ9_0(.din(n1835), .dout(n1832));
    jdff dff_A_SFsbXmIp3_0(.din(n1838), .dout(n1835));
    jdff dff_A_eDkExusl6_0(.din(n1841), .dout(n1838));
    jdff dff_A_zOKPIFGT0_0(.din(n1844), .dout(n1841));
    jdff dff_A_b3AZPMtt0_0(.din(n1847), .dout(n1844));
    jdff dff_A_5TIos0bf5_0(.din(n1850), .dout(n1847));
    jdff dff_A_uxi7vzh40_0(.din(n1853), .dout(n1850));
    jdff dff_A_MvHpnhsP3_0(.din(G204gat), .dout(n1853));
    jdff dff_A_PzE3bIde5_0(.din(n1859), .dout(n1856));
    jdff dff_A_Bo8m3msM2_0(.din(n1862), .dout(n1859));
    jdff dff_A_MaFlRc6b0_0(.din(n1865), .dout(n1862));
    jdff dff_A_7T0qLF1t0_0(.din(n1868), .dout(n1865));
    jdff dff_A_XRxx1xOX2_0(.din(n1871), .dout(n1868));
    jdff dff_A_cbCgttHP2_0(.din(n1874), .dout(n1871));
    jdff dff_A_IJoMRqR09_0(.din(n1877), .dout(n1874));
    jdff dff_A_h1ox0id39_0(.din(n1880), .dout(n1877));
    jdff dff_A_YIRFL45Y3_0(.din(G176gat), .dout(n1880));
    jdff dff_A_7LPMIS6T5_0(.din(n1886), .dout(n1883));
    jdff dff_A_SSlCSCVz4_0(.din(n1889), .dout(n1886));
    jdff dff_A_vfmF4NyB9_0(.din(n1892), .dout(n1889));
    jdff dff_A_LkXr15cg5_0(.din(n1895), .dout(n1892));
    jdff dff_A_iEER2hLt7_0(.din(n1898), .dout(n1895));
    jdff dff_A_Un5U760K9_0(.din(n1901), .dout(n1898));
    jdff dff_A_eujsyPpz6_0(.din(n1904), .dout(n1901));
    jdff dff_A_D9hSKu8z5_0(.din(n1907), .dout(n1904));
    jdff dff_A_PCh4XyPB5_0(.din(G64gat), .dout(n1907));
    jdff dff_A_OBqYfbmd2_0(.din(n1913), .dout(n1910));
    jdff dff_A_MVThQCQA5_0(.din(n1916), .dout(n1913));
    jdff dff_A_CWcUuoNK1_0(.din(n1919), .dout(n1916));
    jdff dff_A_2UtB9Zcd6_0(.din(n1922), .dout(n1919));
    jdff dff_A_CANi5Ovk7_0(.din(n1925), .dout(n1922));
    jdff dff_A_aseJEBhw1_0(.din(n1928), .dout(n1925));
    jdff dff_A_lNHjEzV62_0(.din(n1931), .dout(n1928));
    jdff dff_A_aPrBy7Bg8_0(.din(n1934), .dout(n1931));
    jdff dff_A_1GGE4fA08_0(.din(G57gat), .dout(n1934));
    jdff dff_A_wuYBZTMZ3_0(.din(n1940), .dout(n1937));
    jdff dff_A_pg9F8CUe7_0(.din(n1943), .dout(n1940));
    jdff dff_A_RMfMZ3gQ0_0(.din(n1946), .dout(n1943));
    jdff dff_A_lIc1C1mG9_0(.din(n1949), .dout(n1946));
    jdff dff_A_ym4rWUFL8_0(.din(n1952), .dout(n1949));
    jdff dff_A_iaI64tvM0_0(.din(n1955), .dout(n1952));
    jdff dff_A_1jZkb5BH5_0(.din(n1958), .dout(n1955));
    jdff dff_A_ws9SbgJY5_0(.din(n1961), .dout(n1958));
    jdff dff_A_5H5Qu2fp8_0(.din(G78gat), .dout(n1961));
    jdff dff_A_06RdxNoz1_0(.din(n1967), .dout(n1964));
    jdff dff_A_KXq4lMUl4_0(.din(n1970), .dout(n1967));
    jdff dff_A_mVP3H95v0_0(.din(n1973), .dout(n1970));
    jdff dff_A_bkvL7Zry3_0(.din(n1976), .dout(n1973));
    jdff dff_A_NIVzY5fd2_0(.din(n1979), .dout(n1976));
    jdff dff_A_w4zkEwAy1_0(.din(n1982), .dout(n1979));
    jdff dff_A_dAcgyJP35_0(.din(n1985), .dout(n1982));
    jdff dff_A_ruZ2FblI3_0(.din(n1988), .dout(n1985));
    jdff dff_A_2dZxDKmg0_0(.din(G71gat), .dout(n1988));
    jdff dff_A_bMt68ECE2_0(.din(n1994), .dout(n1991));
    jdff dff_A_ohrVgN8K1_0(.din(n1997), .dout(n1994));
    jdff dff_A_ihmJ1Jyk2_0(.din(n2000), .dout(n1997));
    jdff dff_A_vfgyCCxv5_0(.din(n2003), .dout(n2000));
    jdff dff_A_HHfseiVV0_0(.din(n2006), .dout(n2003));
    jdff dff_A_BCkv0GJW6_0(.din(n2009), .dout(n2006));
    jdff dff_A_pmXJN5zz4_0(.din(n2012), .dout(n2009));
    jdff dff_A_v1EU7C0h5_0(.din(n2015), .dout(n2012));
    jdff dff_A_lpOA4F4J5_0(.din(G141gat), .dout(n2015));
    jdff dff_A_okxgO1ni3_0(.din(n2021), .dout(n2018));
    jdff dff_A_U1xkfmc03_0(.din(n2024), .dout(n2021));
    jdff dff_A_ZwHxMxK22_0(.din(n2027), .dout(n2024));
    jdff dff_A_mb4iWFJr9_0(.din(n2030), .dout(n2027));
    jdff dff_A_oEDoqyTs1_0(.din(n2033), .dout(n2030));
    jdff dff_A_qcdvIQSl2_0(.din(n2036), .dout(n2033));
    jdff dff_A_7tqKszuC9_0(.din(n2039), .dout(n2036));
    jdff dff_A_XOP1tVLg1_0(.din(n2042), .dout(n2039));
    jdff dff_A_XKnK0IpQ6_0(.din(G113gat), .dout(n2042));
    jdff dff_A_M82aSmm46_0(.din(n2048), .dout(n2045));
    jdff dff_A_Bi7oAuZk3_0(.din(n2051), .dout(n2048));
    jdff dff_A_2Tt6bKAx7_0(.din(n2054), .dout(n2051));
    jdff dff_A_0EzhDelN5_0(.din(n2057), .dout(n2054));
    jdff dff_A_lfnwCRGr0_0(.din(n2060), .dout(n2057));
    jdff dff_A_Su8N4dkm6_0(.din(n2063), .dout(n2060));
    jdff dff_A_rA4BjDHP1_0(.din(n2066), .dout(n2063));
    jdff dff_A_xABsGxjL6_0(.din(n2069), .dout(n2066));
    jdff dff_A_zjjB4yPj7_0(.din(G197gat), .dout(n2069));
    jdff dff_A_ITNxiFWO1_0(.din(n2075), .dout(n2072));
    jdff dff_A_0GAmDYEG0_0(.din(n2078), .dout(n2075));
    jdff dff_A_cCLJaDTB5_0(.din(n2081), .dout(n2078));
    jdff dff_A_FKS0Nae47_0(.din(n2084), .dout(n2081));
    jdff dff_A_WLDnIt213_0(.din(n2087), .dout(n2084));
    jdff dff_A_Msrcv5TI8_0(.din(n2090), .dout(n2087));
    jdff dff_A_bfYpLoKM3_0(.din(n2093), .dout(n2090));
    jdff dff_A_Jtm72dm39_0(.din(n2096), .dout(n2093));
    jdff dff_A_qVINdlc98_0(.din(G169gat), .dout(n2096));
    jdff dff_A_g5ucGTYv3_0(.din(n2102), .dout(n2099));
    jdff dff_A_fpguqe7k6_0(.din(n2105), .dout(n2102));
    jdff dff_A_LQumOhCh4_0(.din(n2108), .dout(n2105));
    jdff dff_A_f8xloYDE9_0(.din(n2111), .dout(n2108));
    jdff dff_A_vPsxpE5U0_0(.din(n2114), .dout(n2111));
    jdff dff_A_B6wj2OZ82_0(.din(n2117), .dout(n2114));
    jdff dff_A_bACzojML9_0(.din(n2120), .dout(n2117));
    jdff dff_A_aCkKyiZZ1_0(.din(n2123), .dout(n2120));
    jdff dff_A_Al2kpQAe5_0(.din(G8gat), .dout(n2123));
    jdff dff_A_oafRRrxV5_0(.din(n2129), .dout(n2126));
    jdff dff_A_5Jk1VUSf3_0(.din(n2132), .dout(n2129));
    jdff dff_A_cegwtHUk9_0(.din(n2135), .dout(n2132));
    jdff dff_A_d0X9LXvr2_0(.din(n2138), .dout(n2135));
    jdff dff_A_nH9aCpuJ6_0(.din(n2141), .dout(n2138));
    jdff dff_A_VV1jYwGn7_0(.din(n2144), .dout(n2141));
    jdff dff_A_7DCzvcGn9_0(.din(n2147), .dout(n2144));
    jdff dff_A_hew55QgR0_0(.din(n2150), .dout(n2147));
    jdff dff_A_74XVafv40_0(.din(G1gat), .dout(n2150));
    jdff dff_A_t3N9Lzl06_0(.din(n2156), .dout(n2153));
    jdff dff_A_YtzrjX8m4_0(.din(n2159), .dout(n2156));
    jdff dff_A_2VhIgIbs1_0(.din(n2162), .dout(n2159));
    jdff dff_A_fTqJfZlS1_0(.din(n2165), .dout(n2162));
    jdff dff_A_Zp6V0dhq0_0(.din(n2168), .dout(n2165));
    jdff dff_A_mDXsZaiy8_0(.din(n2171), .dout(n2168));
    jdff dff_A_V8u4KqY41_0(.din(n2174), .dout(n2171));
    jdff dff_A_iOn8XWGc9_0(.din(n2177), .dout(n2174));
    jdff dff_A_IWpObeUi7_0(.din(G22gat), .dout(n2177));
    jdff dff_A_YKtxjwDp5_0(.din(n2183), .dout(n2180));
    jdff dff_A_B2dxem342_0(.din(n2186), .dout(n2183));
    jdff dff_A_SNAnrP8L7_0(.din(n2189), .dout(n2186));
    jdff dff_A_d9jsRY9O0_0(.din(n2192), .dout(n2189));
    jdff dff_A_LkIdX5QS1_0(.din(n2195), .dout(n2192));
    jdff dff_A_bWJxwTdc8_0(.din(n2198), .dout(n2195));
    jdff dff_A_fVrQlfmp4_0(.din(n2201), .dout(n2198));
    jdff dff_A_aPptUyuR1_0(.din(n2204), .dout(n2201));
endmodule

