/*

c880:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jcb: 119
	jdff: 540
	jand: 153

Summary:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jcb: 119
	jdff: 540
	jand: 153
*/

module c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n101;
	wire n102;
	wire n103;
	wire n105;
	wire n106;
	wire n107;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n118;
	wire n119;
	wire n121;
	wire n122;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire [2:0] w_G1gat_0;
	wire [1:0] w_G1gat_1;
	wire [1:0] w_G8gat_0;
	wire [1:0] w_G13gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G17gat_1;
	wire [2:0] w_G17gat_2;
	wire [1:0] w_G26gat_0;
	wire [2:0] w_G29gat_0;
	wire [1:0] w_G36gat_0;
	wire [2:0] w_G42gat_0;
	wire [2:0] w_G42gat_1;
	wire [1:0] w_G42gat_2;
	wire [2:0] w_G51gat_0;
	wire [1:0] w_G51gat_1;
	wire [2:0] w_G55gat_0;
	wire [2:0] w_G59gat_0;
	wire [1:0] w_G59gat_1;
	wire [1:0] w_G68gat_0;
	wire [1:0] w_G75gat_0;
	wire [2:0] w_G80gat_0;
	wire [2:0] w_G91gat_0;
	wire [2:0] w_G96gat_0;
	wire [2:0] w_G101gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G111gat_0;
	wire [2:0] w_G116gat_0;
	wire [2:0] w_G121gat_0;
	wire [1:0] w_G126gat_0;
	wire [1:0] w_G130gat_0;
	wire [2:0] w_G138gat_0;
	wire [1:0] w_G138gat_1;
	wire [1:0] w_G143gat_0;
	wire [1:0] w_G146gat_0;
	wire [1:0] w_G149gat_0;
	wire [2:0] w_G153gat_0;
	wire [1:0] w_G156gat_0;
	wire [2:0] w_G159gat_0;
	wire [2:0] w_G159gat_1;
	wire [1:0] w_G159gat_2;
	wire [2:0] w_G165gat_0;
	wire [2:0] w_G165gat_1;
	wire [1:0] w_G165gat_2;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [1:0] w_G171gat_2;
	wire [2:0] w_G177gat_0;
	wire [2:0] w_G177gat_1;
	wire [1:0] w_G177gat_2;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G183gat_1;
	wire [1:0] w_G183gat_2;
	wire [2:0] w_G189gat_0;
	wire [2:0] w_G189gat_1;
	wire [1:0] w_G189gat_2;
	wire [2:0] w_G195gat_0;
	wire [2:0] w_G195gat_1;
	wire [1:0] w_G195gat_2;
	wire [2:0] w_G201gat_0;
	wire [2:0] w_G201gat_1;
	wire [2:0] w_G201gat_2;
	wire [2:0] w_G210gat_0;
	wire [2:0] w_G210gat_1;
	wire [2:0] w_G210gat_2;
	wire [1:0] w_G210gat_3;
	wire [2:0] w_G219gat_0;
	wire [2:0] w_G219gat_1;
	wire [2:0] w_G219gat_2;
	wire [1:0] w_G219gat_3;
	wire [2:0] w_G228gat_0;
	wire [2:0] w_G228gat_1;
	wire [2:0] w_G228gat_2;
	wire [1:0] w_G228gat_3;
	wire [2:0] w_G237gat_0;
	wire [2:0] w_G237gat_1;
	wire [2:0] w_G237gat_2;
	wire [1:0] w_G237gat_3;
	wire [2:0] w_G246gat_0;
	wire [2:0] w_G246gat_1;
	wire [2:0] w_G246gat_2;
	wire [1:0] w_G246gat_3;
	wire [2:0] w_G255gat_0;
	wire [2:0] w_G261gat_0;
	wire [1:0] w_G268gat_0;
	wire [1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire [2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire [1:0] w_n86_0;
	wire [1:0] w_n88_0;
	wire [2:0] w_n92_0;
	wire [1:0] w_n93_0;
	wire [1:0] w_n96_0;
	wire [1:0] w_n98_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n102_0;
	wire [1:0] w_n106_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n111_0;
	wire [2:0] w_n118_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n143_0;
	wire [1:0] w_n149_0;
	wire [2:0] w_n153_0;
	wire [2:0] w_n153_1;
	wire [2:0] w_n153_2;
	wire [1:0] w_n153_3;
	wire [1:0] w_n154_0;
	wire [1:0] w_n157_0;
	wire [2:0] w_n159_0;
	wire [1:0] w_n159_1;
	wire [1:0] w_n162_0;
	wire [1:0] w_n163_0;
	wire [2:0] w_n165_0;
	wire [2:0] w_n165_1;
	wire [2:0] w_n167_0;
	wire [1:0] w_n167_1;
	wire [2:0] w_n168_0;
	wire [2:0] w_n181_0;
	wire [2:0] w_n181_1;
	wire [2:0] w_n181_2;
	wire [1:0] w_n181_3;
	wire [2:0] w_n193_0;
	wire [1:0] w_n193_1;
	wire [2:0] w_n194_0;
	wire [1:0] w_n196_0;
	wire [1:0] w_n213_0;
	wire [2:0] w_n217_0;
	wire [1:0] w_n217_1;
	wire [1:0] w_n218_0;
	wire [2:0] w_n222_0;
	wire [1:0] w_n222_1;
	wire [1:0] w_n223_0;
	wire [1:0] w_n224_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n230_0;
	wire [1:0] w_n232_0;
	wire [2:0] w_n236_0;
	wire [1:0] w_n238_0;
	wire [2:0] w_n252_0;
	wire [1:0] w_n255_0;
	wire [2:0] w_n273_0;
	wire [2:0] w_n292_0;
	wire [1:0] w_n292_1;
	wire [2:0] w_n296_0;
	wire [1:0] w_n296_1;
	wire [2:0] w_n299_0;
	wire [1:0] w_n299_1;
	wire [1:0] w_n302_0;
	wire [1:0] w_n303_0;
	wire [2:0] w_n305_0;
	wire [1:0] w_n305_1;
	wire [2:0] w_n312_0;
	wire [1:0] w_n312_1;
	wire [1:0] w_n315_0;
	wire [2:0] w_n321_0;
	wire [1:0] w_n321_1;
	wire [1:0] w_n322_0;
	wire [2:0] w_n328_0;
	wire [1:0] w_n328_1;
	wire [2:0] w_n329_0;
	wire [2:0] w_n330_0;
	wire [1:0] w_n331_0;
	wire [2:0] w_n335_0;
	wire [2:0] w_n337_0;
	wire [1:0] w_n339_0;
	wire [1:0] w_n340_0;
	wire [2:0] w_n346_0;
	wire [1:0] w_n346_1;
	wire [2:0] w_n347_0;
	wire [2:0] w_n367_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n405_0;
	wire w_dff_A_CCj0la7k5_1;
	wire w_dff_A_rDQOP6sh4_0;
	wire w_dff_B_LJ2LtJgT0_0;
	wire w_dff_B_C3ikhOSA3_1;
	wire w_dff_B_vrtHSlZA2_0;
	wire w_dff_B_J83LNMHI6_1;
	wire w_dff_B_JeFLVpOz7_0;
	wire w_dff_B_rxMu0aUu8_0;
	wire w_dff_B_FK76auAP9_1;
	wire w_dff_B_ngv4l5OW7_0;
	wire w_dff_B_1vBf8jKj0_2;
	wire w_dff_B_xAVV3AjK3_0;
	wire w_dff_B_2xbdBfGN0_0;
	wire w_dff_B_ftLDdwzc9_0;
	wire w_dff_B_szDRvvjH5_0;
	wire w_dff_B_Clg6Up0v0_0;
	wire w_dff_B_n7iFbRDd4_0;
	wire w_dff_B_PC7QqtZB8_0;
	wire w_dff_B_NUiyhTX28_0;
	wire w_dff_B_FUh0rxZd4_0;
	wire w_dff_B_EmdG73Tw1_0;
	wire w_dff_B_dUrOWA1l6_0;
	wire w_dff_A_S8dJ1eao0_1;
	wire w_dff_A_lEctacaT4_1;
	wire w_dff_A_ldmCPNlp5_1;
	wire w_dff_A_5oV02g2c4_1;
	wire w_dff_A_BrG7DVJx9_1;
	wire w_dff_B_jAkB14bt6_0;
	wire w_dff_B_ZDVyxVTw8_0;
	wire w_dff_B_RmpHZQsp4_0;
	wire w_dff_B_sNNyOCMb6_0;
	wire w_dff_B_vOp2ltun6_0;
	wire w_dff_B_6JdlWv7H4_0;
	wire w_dff_B_lurEB3A76_0;
	wire w_dff_B_PLP1zwJM5_0;
	wire w_dff_B_IBnFkczI7_0;
	wire w_dff_B_MQWdLDRe1_0;
	wire w_dff_B_jlwOerqR1_0;
	wire w_dff_B_Lan5YEWw0_0;
	wire w_dff_B_Xjh5BrIx2_0;
	wire w_dff_B_HXyGwlXN3_0;
	wire w_dff_B_lZn1Q91d1_0;
	wire w_dff_B_51qpWO1A7_0;
	wire w_dff_A_IGR0uvxD3_0;
	wire w_dff_B_2zxUmpFN8_1;
	wire w_dff_B_Z6LMu0yv2_1;
	wire w_dff_B_0x0VDcFI8_1;
	wire w_dff_A_fRiY1ZxT2_1;
	wire w_dff_A_wfXCmYf12_0;
	wire w_dff_A_iY15mJi56_0;
	wire w_dff_A_HkLKhpge1_0;
	wire w_dff_A_BdOGBBQ45_0;
	wire w_dff_A_sppNk25w3_0;
	wire w_dff_B_q2wRB0Pm0_0;
	wire w_dff_B_66Si8Cst7_0;
	wire w_dff_B_x4SaXGzy3_0;
	wire w_dff_B_vq8MgUIk5_0;
	wire w_dff_B_rVJolAeM7_0;
	wire w_dff_B_u835j7zb2_0;
	wire w_dff_B_L2msWCfY5_0;
	wire w_dff_B_3CbSHFDQ2_0;
	wire w_dff_B_IYYquxY82_0;
	wire w_dff_B_wFk9ZHSg1_0;
	wire w_dff_B_8wj4ljoW5_0;
	wire w_dff_B_zB26315c0_0;
	wire w_dff_B_wrSngEM43_1;
	wire w_dff_A_ZIMMHt8I0_1;
	wire w_dff_B_q30TG8ee0_0;
	wire w_dff_B_y3vZdYAA7_0;
	wire w_dff_B_yUedXOTY3_0;
	wire w_dff_B_JLXh2En21_0;
	wire w_dff_B_d6WLqoVw0_0;
	wire w_dff_B_sIA58gZx8_0;
	wire w_dff_B_wX6ngeO32_0;
	wire w_dff_B_wMtcj9Wr3_0;
	wire w_dff_B_XFXdJ0H04_0;
	wire w_dff_B_YoxmnRGE2_0;
	wire w_dff_B_lWefJEvt2_0;
	wire w_dff_B_lojKx3UP5_0;
	wire w_dff_B_aaMXyf4Z4_0;
	wire w_dff_B_hYgvfGge0_0;
	wire w_dff_B_Tw52TlZY2_0;
	wire w_dff_B_jwevzxdE7_0;
	wire w_dff_B_d236LyET3_0;
	wire w_dff_B_DaR8gZ0e4_1;
	wire w_dff_B_GOIu13tQ6_1;
	wire w_dff_B_udC7DLF52_1;
	wire w_dff_B_Twib4wUK2_1;
	wire w_dff_B_wNHj402n7_1;
	wire w_dff_B_hW3SXoDk1_1;
	wire w_dff_B_8HssfsbQ3_1;
	wire w_dff_B_gJILkU1J6_1;
	wire w_dff_B_WNOlCCmX6_1;
	wire w_dff_B_OK4sCdpZ2_1;
	wire w_dff_A_krnsjryp8_0;
	wire w_dff_A_LNLuCyBO1_0;
	wire w_dff_A_0QBMoMtA3_0;
	wire w_dff_A_Qis3FsmZ9_0;
	wire w_dff_A_bs0iN9e84_0;
	wire w_dff_B_DInSCSrx2_0;
	wire w_dff_B_aAzmz2sh9_0;
	wire w_dff_B_cuMCaWMG5_0;
	wire w_dff_B_Sz9vkcB09_0;
	wire w_dff_B_s1xDcGTx5_0;
	wire w_dff_B_pQWVkC0d7_0;
	wire w_dff_B_IfZGlIgN7_0;
	wire w_dff_B_Rb809NdJ9_0;
	wire w_dff_B_plBa4Teo8_0;
	wire w_dff_B_nEEZhE1q7_0;
	wire w_dff_B_ILRiZsNh5_0;
	wire w_dff_B_tFldBsGg2_0;
	wire w_dff_B_n42kkEU89_0;
	wire w_dff_B_KnECL4Uk8_0;
	wire w_dff_B_wM7xfgte6_0;
	wire w_dff_B_mVkx3Uhu7_0;
	wire w_dff_B_tv4rNENE0_0;
	wire w_dff_A_a9YVctBP1_0;
	wire w_dff_A_TDbxvCBp3_0;
	wire w_dff_A_BfEzzLk66_2;
	wire w_dff_B_XLilWEjK9_0;
	wire w_dff_B_lHIcKZeN7_0;
	wire w_dff_B_yVRaUIFk9_0;
	wire w_dff_B_QXa92kVt9_0;
	wire w_dff_A_xZkURrot5_1;
	wire w_dff_A_JHrFwDUc3_1;
	wire w_dff_B_B0T2Q3Bw1_0;
	wire w_dff_B_CHonst4n9_0;
	wire w_dff_B_pgUV00sw9_0;
	wire w_dff_B_Emc52eko9_0;
	wire w_dff_B_7PfSUxZl2_0;
	wire w_dff_B_NhgaEgBY1_0;
	wire w_dff_B_P7BHgjtN7_0;
	wire w_dff_B_U3LbnHYo6_0;
	wire w_dff_B_nCR9WiLN1_0;
	wire w_dff_B_3e0Ei4UV6_0;
	wire w_dff_B_OLlmtcHD2_0;
	wire w_dff_B_In2TtRBe7_0;
	wire w_dff_B_LUMsYR5l2_0;
	wire w_dff_B_bO7wV32L2_0;
	wire w_dff_B_Gqut33oe7_0;
	wire w_dff_B_ZoVfNSFA5_0;
	wire w_dff_B_iXQUVTDT3_0;
	wire w_dff_A_xdJBDRS58_1;
	wire w_dff_B_wLgqbGeo6_0;
	wire w_dff_B_KM37Jo824_0;
	wire w_dff_B_cr0COvcA3_0;
	wire w_dff_B_9Zomai555_0;
	wire w_dff_B_dQ8I0KMw6_0;
	wire w_dff_A_2dSaeeMX2_1;
	wire w_dff_A_SvWCnciy3_1;
	wire w_dff_A_gq5DHJoV3_1;
	wire w_dff_A_bdFAh50x8_1;
	wire w_dff_B_eVBAz78o7_0;
	wire w_dff_B_XZ64hbkZ4_1;
	wire w_dff_B_T0dq7uGJ3_1;
	wire w_dff_B_xhUBfYWX6_1;
	wire w_dff_A_Ij6H6NcE8_1;
	wire w_dff_A_dmDOKtie0_1;
	wire w_dff_A_CVDJVjub8_1;
	wire w_dff_A_JaA2xSVq2_1;
	wire w_dff_A_A7tapQ5o7_1;
	wire w_dff_A_9mTDFcAW3_2;
	wire w_dff_A_gTPJyhz25_2;
	wire w_dff_A_MvHYnNG52_2;
	wire w_dff_A_Ecd11qi83_2;
	wire w_dff_A_lTFbYbgh7_2;
	wire w_dff_A_FWdANqlu2_2;
	wire w_dff_A_e72YSGre0_2;
	wire w_dff_A_PonThVdN3_2;
	wire w_dff_A_BeJcpQUe1_2;
	wire w_dff_B_2VIeRZWQ7_0;
	wire w_dff_A_xhaf7J6J9_1;
	wire w_dff_B_e37gPooD5_1;
	wire w_dff_B_fwDGZ7am9_1;
	wire w_dff_B_7qR9MaT48_1;
	wire w_dff_B_lS967LtZ3_0;
	wire w_dff_B_m7gNxFhF7_1;
	wire w_dff_B_5ZRBshz49_1;
	wire w_dff_B_IfKNjEif3_1;
	wire w_dff_B_ESHZQwp54_1;
	wire w_dff_B_W8XVATZZ4_1;
	wire w_dff_B_55b2vjm40_0;
	wire w_dff_B_shj27mWZ2_0;
	wire w_dff_B_dKUX8KWL8_0;
	wire w_dff_B_WDvzYpgM8_0;
	wire w_dff_B_KPucb13f2_0;
	wire w_dff_B_DvaqvEzh1_0;
	wire w_dff_B_fXLA1Kwg5_0;
	wire w_dff_B_uGceBSXD1_0;
	wire w_dff_B_JR4jmXGn9_0;
	wire w_dff_B_yXmJwQZz2_0;
	wire w_dff_B_S9knLuoz8_0;
	wire w_dff_B_gJI4gtky3_0;
	wire w_dff_A_VMdr5KKs9_1;
	wire w_dff_A_cGuV4qg22_1;
	wire w_dff_A_yw5pB7ZU7_1;
	wire w_dff_A_pL6PNmqM0_1;
	wire w_dff_B_QJdRNliO0_0;
	wire w_dff_B_TCeDcF568_0;
	wire w_dff_B_OuzKgyVk5_0;
	wire w_dff_B_zUO9LkF29_0;
	wire w_dff_B_aFNtfmEe2_0;
	wire w_dff_B_IFk6j4hx5_0;
	wire w_dff_B_t7OGI33X9_1;
	wire w_dff_B_NFjd6RZw2_1;
	wire w_dff_B_AWWx6la81_1;
	wire w_dff_B_UHBdicTG1_1;
	wire w_dff_B_OmVkDI6T6_1;
	wire w_dff_B_bCXKeL3Q5_1;
	wire w_dff_B_8lLe8bRO6_1;
	wire w_dff_B_FS4S2gvY5_1;
	wire w_dff_B_VXZhZo694_0;
	wire w_dff_B_1rxVpd3B8_0;
	wire w_dff_B_TNE1fgSQ0_0;
	wire w_dff_B_Q7tIZrvg0_0;
	wire w_dff_A_F26RWqfw3_0;
	wire w_dff_A_w6cCnhXf2_0;
	wire w_dff_A_tP72KhmC0_2;
	wire w_dff_A_LR4Lx2Rl6_2;
	wire w_dff_A_DQ2OP5lH2_0;
	wire w_dff_A_jXjURwr55_0;
	wire w_dff_A_1eFlQMwc5_2;
	wire w_dff_B_hdsHP5x36_1;
	wire w_dff_A_OrTZDfrS0_0;
	wire w_dff_A_0NPLWfx13_0;
	wire w_dff_A_1uYTxSc76_0;
	wire w_dff_A_GroTSMkX2_0;
	wire w_dff_A_hqLRdRXR7_0;
	wire w_dff_A_4QdAKl7x2_0;
	wire w_dff_A_Toq34Ftp1_1;
	wire w_dff_A_u0MbFUW69_1;
	wire w_dff_A_26T9gUqU7_1;
	wire w_dff_B_EBdouLYV6_0;
	wire w_dff_B_hG7FzfcC7_0;
	wire w_dff_B_26EsKGKc5_0;
	wire w_dff_B_8hh0wXRo8_0;
	wire w_dff_A_kde8KbWV6_1;
	wire w_dff_A_IYTe57Ow2_1;
	wire w_dff_A_NEqkcji58_1;
	wire w_dff_A_7fLYM1J14_1;
	wire w_dff_A_nRO6zlfJ6_1;
	wire w_dff_A_kkTtHLAr6_2;
	wire w_dff_A_dcmf4uhW4_2;
	wire w_dff_A_avPUcebe7_2;
	wire w_dff_A_Tuh0rk8I1_2;
	wire w_dff_A_xpiXnAg21_2;
	wire w_dff_A_hrMTLzGq3_2;
	wire w_dff_A_ZqPDn6VT1_2;
	wire w_dff_A_fS6lAHk55_2;
	wire w_dff_A_UlOMJKSX8_2;
	wire w_dff_B_IUIDNKMu1_0;
	wire w_dff_B_UGlBo0xK1_0;
	wire w_dff_B_TNUumohk1_0;
	wire w_dff_B_EMxNHy8h2_0;
	wire w_dff_B_hm1XeEtH1_0;
	wire w_dff_B_SLMKw8mj6_0;
	wire w_dff_B_cu1HmymM7_0;
	wire w_dff_B_gxFDA8u96_0;
	wire w_dff_B_OHzfU9DY0_0;
	wire w_dff_B_bqNuC5lG2_0;
	wire w_dff_B_qDcTqQTy0_0;
	wire w_dff_B_E01akAsv8_0;
	wire w_dff_A_xFuZkLqu4_1;
	wire w_dff_A_eeNuPG999_1;
	wire w_dff_A_exMt7xXh8_1;
	wire w_dff_A_OoE4TLiA8_1;
	wire w_dff_B_bTk1evDX6_1;
	wire w_dff_A_rroH0NRy0_0;
	wire w_dff_A_iJ7ti8ja8_0;
	wire w_dff_B_rQ53D53U7_0;
	wire w_dff_B_bstnPsQi3_0;
	wire w_dff_B_URpqphkC3_0;
	wire w_dff_B_LH0q07pu1_0;
	wire w_dff_B_EDrNy9Qv7_3;
	wire w_dff_B_I197bpcy1_3;
	wire w_dff_B_cB3UcaAg3_3;
	wire w_dff_B_gHPIPODr6_3;
	wire w_dff_B_FXZdrSVc9_3;
	wire w_dff_B_Y2SJCPfc4_3;
	wire w_dff_B_2e29grpO7_3;
	wire w_dff_B_QRYtAD1m5_0;
	wire w_dff_B_IynLEhcC6_0;
	wire w_dff_A_oaewuqkV7_2;
	wire w_dff_A_3fbe5yX90_0;
	wire w_dff_A_Yhi45xwW4_0;
	wire w_dff_A_4ENWc2UQ5_0;
	wire w_dff_B_3dvAC20P0_3;
	wire w_dff_B_JJ8quy0X9_3;
	wire w_dff_B_7IxA7YG45_3;
	wire w_dff_B_8AfPiWn38_3;
	wire w_dff_B_LynXWjTt5_3;
	wire w_dff_B_pxyp9p9L1_3;
	wire w_dff_B_Trd5Tr939_1;
	wire w_dff_B_MwRscJ6z0_1;
	wire w_dff_B_UgSJfTAn9_1;
	wire w_dff_B_CqbQpbKg4_1;
	wire w_dff_B_rXqprOXe5_1;
	wire w_dff_B_Lk9n5vFc8_1;
	wire w_dff_B_IWlkaJ328_1;
	wire w_dff_B_vgmAWVGe2_1;
	wire w_dff_B_1vPFDyg56_1;
	wire w_dff_B_EuNeFiDO4_0;
	wire w_dff_B_yWqxq0RV0_0;
	wire w_dff_B_Wkn7JBwa7_0;
	wire w_dff_B_mDSeZK8l5_0;
	wire w_dff_B_83uWI9Ei6_0;
	wire w_dff_A_meshnIlr3_0;
	wire w_dff_A_o8ZADDjP9_0;
	wire w_dff_A_EfEh2nT13_0;
	wire w_dff_A_AqKNoOu96_0;
	wire w_dff_A_AR0qnh854_0;
	wire w_dff_A_jhnaDi6Q5_0;
	wire w_dff_A_0ruHWeOA0_0;
	wire w_dff_A_tSi1udYA9_0;
	wire w_dff_B_Y21dHlA20_1;
	wire w_dff_B_lFQHA1xg4_1;
	wire w_dff_B_F7k906ye5_1;
	wire w_dff_B_6Wsnj20d7_1;
	wire w_dff_B_mnDYvqjb1_1;
	wire w_dff_B_nL8RapGL9_1;
	wire w_dff_B_narWwQcN6_1;
	wire w_dff_B_aHVTPXgO2_0;
	wire w_dff_B_Trua98Zs7_1;
	wire w_dff_A_V8hvUBDX6_0;
	wire w_dff_A_Cv2sEDgY6_1;
	wire w_dff_A_apuwql6P9_1;
	wire w_dff_A_hgx5JAxi9_1;
	wire w_dff_A_rcEbG1DU5_1;
	wire w_dff_A_PEiE3VZj4_1;
	wire w_dff_A_ZwhRxtqS7_2;
	wire w_dff_A_I2fEbQkG9_2;
	wire w_dff_A_7IM0uEVl7_2;
	wire w_dff_A_OXLvQ9607_2;
	wire w_dff_A_MAcl6UMd6_2;
	wire w_dff_A_fUtHtfC04_1;
	wire w_dff_A_EMXOtX4A2_1;
	wire w_dff_A_IWsJA5zo2_1;
	wire w_dff_A_9eTEvFFl6_1;
	wire w_dff_A_shIFNGEE6_1;
	wire w_dff_A_aSZ1xRXd1_2;
	wire w_dff_A_Z8WyBcoU9_2;
	wire w_dff_A_sGhJTLmD8_2;
	wire w_dff_A_0GZ52bW43_2;
	wire w_dff_A_xVuBfEC40_2;
	wire w_dff_B_61OrHqTo4_0;
	wire w_dff_B_AL7EJi0i1_0;
	wire w_dff_A_PNKwbeGg8_0;
	wire w_dff_A_fwagVIfq9_0;
	wire w_dff_A_9YJutSWW9_0;
	wire w_dff_A_RinIkOCv8_0;
	wire w_dff_A_lavV9sd30_0;
	wire w_dff_A_ozYhWeqW5_0;
	wire w_dff_A_smbCcj5w4_0;
	wire w_dff_A_xQO5tiDz8_0;
	wire w_dff_A_EiDKGSNC4_0;
	wire w_dff_A_cckamYwI8_0;
	wire w_dff_A_ROfnJ5Yt5_2;
	wire w_dff_A_YeruOvK76_2;
	wire w_dff_A_BQ90wCFA9_2;
	wire w_dff_A_SjwLYvEt5_2;
	wire w_dff_A_XbNcbaxR3_0;
	wire w_dff_A_tvGuVQJn9_1;
	wire w_dff_A_Jgz18uXf7_1;
	wire w_dff_A_F5XMcJzC9_1;
	wire w_dff_A_CimypAnj1_1;
	wire w_dff_B_vyXG6hTQ3_2;
	wire w_dff_B_E2MeZ04I1_2;
	wire w_dff_B_9EYRklc78_2;
	wire w_dff_B_zbrf4LS31_2;
	wire w_dff_A_xYCSH7WV4_0;
	wire w_dff_A_BfioD60e7_0;
	wire w_dff_A_GzkKLqZq9_0;
	wire w_dff_A_lV2ZbfwP1_0;
	wire w_dff_A_RvVo3Sl95_0;
	wire w_dff_A_Mwx6w1xR2_2;
	wire w_dff_A_ZYLUP0gu4_2;
	wire w_dff_A_hGaAqTP40_2;
	wire w_dff_A_fNGl3RZk3_2;
	wire w_dff_B_UPcoI7sI3_1;
	wire w_dff_B_kwGqkp5m8_1;
	wire w_dff_B_0XRj0AEU8_1;
	wire w_dff_B_nB9njjf62_1;
	wire w_dff_B_LRtxNgy08_1;
	wire w_dff_B_YR9TAPNw9_1;
	wire w_dff_B_uZ4htwsd5_1;
	wire w_dff_B_fsrMkPh27_1;
	wire w_dff_B_0eKCEbDJ8_1;
	wire w_dff_B_Wv37bgjK0_1;
	wire w_dff_B_O6XjXY0V3_1;
	wire w_dff_A_2UdM7RhN4_1;
	wire w_dff_A_OICYdldO3_0;
	wire w_dff_B_00vgoY1g7_2;
	wire w_dff_B_U1KzZo9Y5_2;
	wire w_dff_B_LYo6SleD5_2;
	wire w_dff_B_hqW6uudj2_2;
	wire w_dff_B_S3J6TAuL5_2;
	wire w_dff_B_rqeHkNQs4_2;
	wire w_dff_A_uWkGS9cc4_0;
	wire w_dff_A_VN7NTbAY7_0;
	wire w_dff_A_wOJn1mwW2_0;
	wire w_dff_A_sYJNZTGl0_0;
	wire w_dff_A_EvZfo1l24_0;
	wire w_dff_A_hyshpDJ33_1;
	wire w_dff_A_FzZXfQwl5_1;
	wire w_dff_A_ZCtu9FJf5_1;
	wire w_dff_A_rELLcDRh6_1;
	wire w_dff_A_W0PampPv6_1;
	wire w_dff_A_nlLGuuQ96_1;
	wire w_dff_A_IelfkTM72_0;
	wire w_dff_A_efxspf6Y1_0;
	wire w_dff_A_c65xE3uH0_0;
	wire w_dff_A_lf6NpmqY2_0;
	wire w_dff_A_uUVRCGzd9_1;
	wire w_dff_A_iyjeknyI0_1;
	wire w_dff_A_I4iK7PvG7_1;
	wire w_dff_A_vTf2BcLL8_1;
	wire w_dff_A_umEvOaAC1_1;
	wire w_dff_A_0HQrlmgz6_2;
	wire w_dff_A_dtkCYSJt1_2;
	wire w_dff_A_dwTOpPhS0_2;
	wire w_dff_A_1Ilctpke0_2;
	wire w_dff_A_ak03yzzv9_2;
	wire w_dff_A_HBMqRywl4_2;
	wire w_dff_A_NH9NBmG28_2;
	wire w_dff_A_1lz8NpTd1_2;
	wire w_dff_A_PdBieuzD8_2;
	wire w_dff_A_yW1cWfIT3_1;
	wire w_dff_A_zL7JR5nd9_1;
	wire w_dff_A_CWcQXXlt9_1;
	wire w_dff_A_fq5Nvc0t6_1;
	wire w_dff_A_1bNLhzwk4_1;
	wire w_dff_A_KVWEHmL78_1;
	wire w_dff_A_i8kZMIhV1_1;
	wire w_dff_A_NzuKRQ147_1;
	wire w_dff_A_u0OO4cb02_1;
	wire w_dff_A_BY2TtJ9M2_2;
	wire w_dff_A_LjJcmoBW0_1;
	wire w_dff_A_fgfiDB7k9_2;
	wire w_dff_B_y2uImBIK9_0;
	wire w_dff_A_5w84HB3h2_0;
	wire w_dff_A_diRpe3DD4_0;
	wire w_dff_A_h23fIEli9_0;
	wire w_dff_B_0qKh4jwL3_2;
	wire w_dff_B_hkQR92ex7_2;
	wire w_dff_B_HRJctjGL9_2;
	wire w_dff_B_jZrZfJia1_2;
	wire w_dff_A_J27AVUAR9_0;
	wire w_dff_A_OvJAZY9D2_0;
	wire w_dff_A_ShPg6NR06_0;
	wire w_dff_A_TuwgX4D81_0;
	wire w_dff_A_29NPMiPM0_0;
	wire w_dff_A_UJ5DfTng2_1;
	wire w_dff_A_Cq9cKhTU2_1;
	wire w_dff_A_zKbzkcZs4_1;
	wire w_dff_A_B6XSKzLl1_1;
	wire w_dff_A_t31raUJ22_2;
	wire w_dff_A_UFZ17GAg2_2;
	wire w_dff_A_JbebVzyX0_2;
	wire w_dff_A_gb44LIHt8_2;
	wire w_dff_A_AWuuuy1O1_2;
	wire w_dff_A_mv9Ijic62_0;
	wire w_dff_A_7mrNzY6F7_0;
	wire w_dff_A_HLFM1v4Q5_0;
	wire w_dff_B_XINNHBO48_0;
	wire w_dff_B_dcKwdGaG9_0;
	wire w_dff_B_t95ur5B18_0;
	wire w_dff_B_SLajnLwI2_0;
	wire w_dff_A_BjRnuQXE3_0;
	wire w_dff_A_NTncug3v0_0;
	wire w_dff_A_bsnBVwCy1_0;
	wire w_dff_A_XwzX1IZ20_0;
	wire w_dff_A_ub3SxmpZ7_2;
	wire w_dff_A_S2iu9R9u6_2;
	wire w_dff_A_HKtZAJux6_2;
	wire w_dff_A_rlkd52HL6_2;
	wire w_dff_A_1sazUBmb2_0;
	wire w_dff_A_9Tfmcu5G7_0;
	wire w_dff_A_hef7QGLh9_0;
	wire w_dff_A_GbRvA3zS6_0;
	wire w_dff_A_KDGTZ9aa0_1;
	wire w_dff_A_lbnqP6Tt5_1;
	wire w_dff_A_Lsj4Xj5k0_1;
	wire w_dff_A_MCWmQIrb5_1;
	wire w_dff_A_QekXYpaX6_1;
	wire w_dff_A_g41BBauG7_2;
	wire w_dff_A_SDZjQGG05_2;
	wire w_dff_A_de0TFssx3_2;
	wire w_dff_A_JGXvROUQ1_2;
	wire w_dff_A_2g5bkTSe1_2;
	wire w_dff_A_YoYoaWoM3_2;
	wire w_dff_A_dSGpSOxS7_2;
	wire w_dff_A_iQWTMBlT9_2;
	wire w_dff_A_lK7Kh6sK2_2;
	wire w_dff_A_T6w0xhap3_1;
	wire w_dff_A_Z2WIqNpL3_1;
	wire w_dff_A_hZVUsbC05_1;
	wire w_dff_B_csxKrAiS0_0;
	wire w_dff_B_gsxFArij2_0;
	wire w_dff_B_9cGXaGUD9_0;
	wire w_dff_B_eZOCjBFj3_0;
	wire w_dff_B_adY790d46_0;
	wire w_dff_A_TQAuJOTq3_0;
	wire w_dff_A_19gmqj0u0_2;
	wire w_dff_A_0saY8HNr4_2;
	wire w_dff_A_Wwlk23wm8_2;
	wire w_dff_A_kSgMlmBC1_0;
	wire w_dff_A_i5nDzkmp4_2;
	wire w_dff_B_zgDD9V7H8_0;
	wire w_dff_A_5jSJjxvG8_0;
	wire w_dff_A_RizNux0Q9_0;
	wire w_dff_A_9yJbgLEK7_0;
	wire w_dff_A_NikhT9437_1;
	wire w_dff_B_mt5ssUfw0_2;
	wire w_dff_B_KTo6driW8_2;
	wire w_dff_B_ApiLYihH5_2;
	wire w_dff_B_l7oNFS4D0_2;
	wire w_dff_B_mHbV2ANM1_0;
	wire w_dff_B_nBrgfEWu0_0;
	wire w_dff_A_A8Hsb4HS4_1;
	wire w_dff_A_pbatWKxq6_1;
	wire w_dff_A_Uz76hR5G2_1;
	wire w_dff_A_0XKpT3Ew1_1;
	wire w_dff_A_QGe30xk99_1;
	wire w_dff_A_swdxVTFa7_1;
	wire w_dff_A_VRGvpubH9_1;
	wire w_dff_A_s6aV5ion3_1;
	wire w_dff_A_n3EUFogI7_1;
	wire w_dff_A_sV31scwQ2_1;
	wire w_dff_A_PoH7qbrr6_1;
	wire w_dff_A_chaatoJs8_1;
	wire w_dff_A_pdHOZErm1_1;
	wire w_dff_A_E1ZocGjz7_2;
	wire w_dff_A_Z6xMvZQA4_2;
	wire w_dff_A_ZYIVTPXM7_2;
	wire w_dff_A_lV20OZUB2_2;
	wire w_dff_A_qLVc8urX8_2;
	wire w_dff_A_setf41397_2;
	wire w_dff_A_l0tJHxvQ6_2;
	wire w_dff_A_PHjBPaZv9_2;
	wire w_dff_A_oD1Gvndw5_2;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(G388gat),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(G389gat),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(G391gat),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_G17gat_2[2]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_n92_0[2]),.dout(G418gat),.clk(gclk));
	jnot g009(.din(w_n93_0[0]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G1gat_1[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G26gat_0[1]),.dout(n97),.clk(gclk));
	jcb g012(.dina(n97),.dinb(w_n96_0[1]),.dout(n98));
	jcb g013(.dina(w_n98_0[1]),.dinb(n95),.dout(n99));
	jcb g014(.dina(w_n99_0[1]),.dinb(w_G390gat_0[1]),.dout(G419gat));
	jnot g015(.din(w_G80gat_0[1]),.dout(n101),.clk(gclk));
	jand g016(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n102),.clk(gclk));
	jnot g017(.din(w_n102_0[1]),.dout(n103),.clk(gclk));
	jcb g018(.dina(n103),.dinb(w_n101_0[1]),.dout(G420gat));
	jnot g019(.din(w_G36gat_0[0]),.dout(n105),.clk(gclk));
	jnot g020(.din(w_G59gat_1[0]),.dout(n106),.clk(gclk));
	jcb g021(.dina(w_n106_0[1]),.dinb(n105),.dout(n107));
	jcb g022(.dina(w_n107_0[1]),.dinb(w_n101_0[0]),.dout(G421gat));
	jnot g023(.din(w_G42gat_1[2]),.dout(n109),.clk(gclk));
	jcb g024(.dina(w_n107_0[0]),.dinb(n109),.dout(G422gat));
	jcb g025(.dina(G88gat),.dinb(G87gat),.dout(n111));
	jand g026(.dina(w_n111_0[1]),.dinb(G90gat),.dout(G423gat),.clk(gclk));
	jnot g027(.din(w_G390gat_0[0]),.dout(n113),.clk(gclk));
	jcb g028(.dina(w_n99_0[0]),.dinb(n113),.dout(G446gat));
	jand g029(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n115),.clk(gclk));
	jand g030(.dina(n115),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g031(.dina(w_G55gat_0[2]),.dinb(w_G13gat_0[0]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_n92_0[1]),.dout(n118),.clk(gclk));
	jand g033(.dina(w_G68gat_0[1]),.dinb(w_G29gat_0[0]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_dff_B_LJ2LtJgT0_0),.dinb(w_n118_0[2]),.dout(G448gat),.clk(gclk));
	jand g035(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n121),.clk(gclk));
	jand g036(.dina(w_n121_0[1]),.dinb(w_dff_B_C3ikhOSA3_1),.dout(n122),.clk(gclk));
	jand g037(.dina(n122),.dinb(w_n118_0[1]),.dout(G449gat),.clk(gclk));
	jand g038(.dina(w_n111_0[0]),.dinb(G89gat),.dout(G450gat),.clk(gclk));
	jxor g039(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n125),.clk(gclk));
	jxor g040(.dina(n125),.dinb(w_G130gat_0[1]),.dout(n126),.clk(gclk));
	jxor g041(.dina(w_G126gat_0[1]),.dinb(w_G121gat_0[2]),.dout(n127),.clk(gclk));
	jxor g042(.dina(w_dff_B_JeFLVpOz7_0),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g043(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n129),.clk(gclk));
	jxor g044(.dina(n129),.dinb(w_dff_B_J83LNMHI6_1),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(w_dff_B_vrtHSlZA2_0),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n128),.dout(G767gat),.clk(gclk));
	jxor g048(.dina(w_G165gat_2[1]),.dinb(w_G159gat_2[1]),.dout(n134),.clk(gclk));
	jxor g049(.dina(n134),.dinb(w_G130gat_0[0]),.dout(n135),.clk(gclk));
	jxor g050(.dina(w_G201gat_2[2]),.dinb(w_G195gat_2[1]),.dout(n136),.clk(gclk));
	jxor g051(.dina(w_dff_B_ngv4l5OW7_0),.dinb(n135),.dout(n137),.clk(gclk));
	jxor g052(.dina(w_G189gat_2[1]),.dinb(w_G183gat_2[1]),.dout(n138),.clk(gclk));
	jxor g053(.dina(n138),.dinb(w_dff_B_FK76auAP9_1),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G177gat_2[1]),.dinb(w_G171gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(w_dff_B_rxMu0aUu8_0),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n137),.dout(G768gat),.clk(gclk));
	jnot g057(.din(w_G261gat_0[2]),.dout(n143),.clk(gclk));
	jand g058(.dina(w_n102_0[0]),.dinb(w_G42gat_1[1]),.dout(n144),.clk(gclk));
	jnot g059(.din(n144),.dout(n145),.clk(gclk));
	jand g060(.dina(w_G51gat_1[0]),.dinb(w_G17gat_2[1]),.dout(n146),.clk(gclk));
	jand g061(.dina(n146),.dinb(w_n92_0[0]),.dout(n147),.clk(gclk));
	jand g062(.dina(w_dff_B_nBrgfEWu0_0),.dinb(n145),.dout(n148),.clk(gclk));
	jand g063(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n149),.clk(gclk));
	jxor g064(.dina(w_G42gat_1[0]),.dinb(w_G17gat_2[0]),.dout(n150),.clk(gclk));
	jand g065(.dina(n150),.dinb(w_n149_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(n151),.dinb(w_G447gat_1),.dout(n152),.clk(gclk));
	jcb g067(.dina(w_dff_B_mHbV2ANM1_0),.dinb(n148),.dout(n153));
	jand g068(.dina(w_n153_3[1]),.dinb(w_G126gat_0[0]),.dout(n154),.clk(gclk));
	jnot g069(.din(w_G156gat_0[0]),.dout(n155),.clk(gclk));
	jcb g070(.dina(n155),.dinb(w_n106_0[0]),.dout(n156));
	jand g071(.dina(w_dff_B_zgDD9V7H8_0),.dinb(w_G447gat_0[2]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n157_0[1]),.dinb(w_G17gat_1[2]),.dout(n158),.clk(gclk));
	jcb g073(.dina(n158),.dinb(w_n96_0[0]),.dout(n159));
	jand g074(.dina(w_n159_1[1]),.dinb(w_G153gat_0[2]),.dout(n160),.clk(gclk));
	jand g075(.dina(w_n86_0[0]),.dinb(w_G80gat_0[0]),.dout(n161),.clk(gclk));
	jand g076(.dina(n161),.dinb(w_G447gat_0[1]),.dout(n162),.clk(gclk));
	jnot g077(.din(w_G268gat_0[1]),.dout(n163),.clk(gclk));
	jand g078(.dina(w_n163_0[1]),.dinb(w_G55gat_0[1]),.dout(n164),.clk(gclk));
	jand g079(.dina(w_dff_B_y2uImBIK9_0),.dinb(w_n162_0[1]),.dout(n165),.clk(gclk));
	jcb g080(.dina(w_n165_1[2]),.dinb(n160),.dout(n166));
	jcb g081(.dina(n166),.dinb(w_n154_0[1]),.dout(n167));
	jxor g082(.dina(w_n167_1[1]),.dinb(w_G201gat_2[1]),.dout(n168),.clk(gclk));
	jnot g083(.din(w_n168_0[2]),.dout(n169),.clk(gclk));
	jcb g084(.dina(n169),.dinb(w_n143_0[1]),.dout(n170));
	jcb g085(.dina(w_n168_0[1]),.dinb(w_G261gat_0[1]),.dout(n171));
	jand g086(.dina(n171),.dinb(w_G219gat_3[1]),.dout(n172),.clk(gclk));
	jand g087(.dina(n172),.dinb(n170),.dout(n173),.clk(gclk));
	jand g088(.dina(w_n168_0[0]),.dinb(w_G228gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_G237gat_3[1]),.dinb(w_G201gat_2[0]),.dout(n175),.clk(gclk));
	jcb g090(.dina(n175),.dinb(w_G246gat_3[1]),.dout(n176));
	jand g091(.dina(w_dff_B_dUrOWA1l6_0),.dinb(w_n167_1[0]),.dout(n177),.clk(gclk));
	jand g092(.dina(G72gat),.dinb(w_G42gat_0[2]),.dout(n178),.clk(gclk));
	jand g093(.dina(n178),.dinb(w_dff_B_bTk1evDX6_1),.dout(n179),.clk(gclk));
	jand g094(.dina(n179),.dinb(w_n121_0[0]),.dout(n180),.clk(gclk));
	jand g095(.dina(n180),.dinb(w_n118_0[0]),.dout(n181),.clk(gclk));
	jand g096(.dina(w_n181_3[1]),.dinb(w_G201gat_1[2]),.dout(n182),.clk(gclk));
	jand g097(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n183),.clk(gclk));
	jand g098(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n184),.clk(gclk));
	jcb g099(.dina(n184),.dinb(n183),.dout(n185));
	jcb g100(.dina(w_dff_B_PC7QqtZB8_0),.dinb(n182),.dout(n186));
	jcb g101(.dina(w_dff_B_ftLDdwzc9_0),.dinb(n177),.dout(n187));
	jcb g102(.dina(w_dff_B_2xbdBfGN0_0),.dinb(n174),.dout(n188));
	jcb g103(.dina(w_dff_B_xAVV3AjK3_0),.dinb(n173),.dout(G850gat));
	jand g104(.dina(w_n159_1[0]),.dinb(w_G143gat_0[1]),.dout(n190),.clk(gclk));
	jand g105(.dina(w_n153_3[0]),.dinb(w_G111gat_0[1]),.dout(n191),.clk(gclk));
	jcb g106(.dina(n191),.dinb(w_n165_1[1]),.dout(n192));
	jcb g107(.dina(n192),.dinb(n190),.dout(n193));
	jxor g108(.dina(w_n193_1[1]),.dinb(w_G183gat_2[0]),.dout(n194),.clk(gclk));
	jnot g109(.din(w_n194_0[2]),.dout(n195),.clk(gclk));
	jand g110(.dina(w_n167_0[2]),.dinb(w_G201gat_1[1]),.dout(n196),.clk(gclk));
	jnot g111(.din(w_n196_0[1]),.dout(n197),.clk(gclk));
	jnot g112(.din(w_G201gat_1[0]),.dout(n198),.clk(gclk));
	jnot g113(.din(w_n154_0[0]),.dout(n199),.clk(gclk));
	jnot g114(.din(w_G153gat_0[1]),.dout(n200),.clk(gclk));
	jnot g115(.din(w_G17gat_1[1]),.dout(n201),.clk(gclk));
	jnot g116(.din(w_G51gat_0[2]),.dout(n202),.clk(gclk));
	jcb g117(.dina(w_n98_0[0]),.dinb(n202),.dout(n203));
	jcb g118(.dina(w_n149_0[0]),.dinb(n203),.dout(n204));
	jcb g119(.dina(n204),.dinb(n201),.dout(n205));
	jand g120(.dina(n205),.dinb(w_G1gat_0[1]),.dout(n206),.clk(gclk));
	jcb g121(.dina(n206),.dinb(w_dff_B_O6XjXY0V3_1),.dout(n207));
	jnot g122(.din(w_n165_1[0]),.dout(n208),.clk(gclk));
	jand g123(.dina(n208),.dinb(w_dff_B_Wv37bgjK0_1),.dout(n209),.clk(gclk));
	jand g124(.dina(n209),.dinb(n199),.dout(n210),.clk(gclk));
	jand g125(.dina(n210),.dinb(w_dff_B_uZ4htwsd5_1),.dout(n211),.clk(gclk));
	jcb g126(.dina(n211),.dinb(w_n143_0[0]),.dout(n212));
	jand g127(.dina(n212),.dinb(w_dff_B_UPcoI7sI3_1),.dout(n213),.clk(gclk));
	jand g128(.dina(w_n159_0[2]),.dinb(w_G146gat_0[1]),.dout(n214),.clk(gclk));
	jand g129(.dina(w_n153_2[2]),.dinb(w_G116gat_0[1]),.dout(n215),.clk(gclk));
	jcb g130(.dina(n215),.dinb(w_n165_0[2]),.dout(n216));
	jcb g131(.dina(n216),.dinb(n214),.dout(n217));
	jcb g132(.dina(w_n217_1[1]),.dinb(w_G189gat_2[0]),.dout(n218));
	jand g133(.dina(w_n159_0[1]),.dinb(w_G149gat_0[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n153_2[1]),.dinb(w_G121gat_0[0]),.dout(n220),.clk(gclk));
	jcb g135(.dina(n220),.dinb(w_n165_0[1]),.dout(n221));
	jcb g136(.dina(n221),.dinb(n219),.dout(n222));
	jcb g137(.dina(w_n222_1[1]),.dinb(w_G195gat_2[0]),.dout(n223));
	jand g138(.dina(w_n223_0[1]),.dinb(w_n218_0[1]),.dout(n224),.clk(gclk));
	jnot g139(.din(w_n224_0[1]),.dout(n225),.clk(gclk));
	jcb g140(.dina(w_dff_B_AL7EJi0i1_0),.dinb(w_n213_0[1]),.dout(n226));
	jand g141(.dina(w_n217_1[0]),.dinb(w_G189gat_1[2]),.dout(n227),.clk(gclk));
	jand g142(.dina(w_n222_1[0]),.dinb(w_G195gat_1[2]),.dout(n228),.clk(gclk));
	jand g143(.dina(w_n228_0[1]),.dinb(w_n218_0[0]),.dout(n229),.clk(gclk));
	jcb g144(.dina(n229),.dinb(w_dff_B_Trua98Zs7_1),.dout(n230));
	jnot g145(.din(w_n230_0[1]),.dout(n231),.clk(gclk));
	jand g146(.dina(w_dff_B_aHVTPXgO2_0),.dinb(n226),.dout(n232),.clk(gclk));
	jcb g147(.dina(w_n232_0[1]),.dinb(w_dff_B_0x0VDcFI8_1),.dout(n233));
	jcb g148(.dina(w_n167_0[1]),.dinb(w_G201gat_0[2]),.dout(n234));
	jand g149(.dina(n234),.dinb(w_G261gat_0[0]),.dout(n235),.clk(gclk));
	jcb g150(.dina(n235),.dinb(w_n196_0[0]),.dout(n236));
	jand g151(.dina(w_n224_0[0]),.dinb(w_n236_0[2]),.dout(n237),.clk(gclk));
	jcb g152(.dina(w_n230_0[0]),.dinb(n237),.dout(n238));
	jcb g153(.dina(w_n238_0[1]),.dinb(w_n194_0[1]),.dout(n239));
	jand g154(.dina(n239),.dinb(w_G219gat_3[0]),.dout(n240),.clk(gclk));
	jand g155(.dina(w_dff_B_51qpWO1A7_0),.dinb(n233),.dout(n241),.clk(gclk));
	jand g156(.dina(w_n194_0[0]),.dinb(w_G228gat_3[0]),.dout(n242),.clk(gclk));
	jand g157(.dina(w_G237gat_3[0]),.dinb(w_G183gat_1[2]),.dout(n243),.clk(gclk));
	jcb g158(.dina(n243),.dinb(w_G246gat_3[0]),.dout(n244));
	jand g159(.dina(w_dff_B_HXyGwlXN3_0),.dinb(w_n193_1[0]),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n181_3[0]),.dinb(w_G183gat_1[1]),.dout(n246),.clk(gclk));
	jand g161(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n247),.clk(gclk));
	jcb g162(.dina(w_dff_B_MQWdLDRe1_0),.dinb(n246),.dout(n248));
	jcb g163(.dina(w_dff_B_6JdlWv7H4_0),.dinb(n245),.dout(n249));
	jcb g164(.dina(w_dff_B_vOp2ltun6_0),.dinb(n242),.dout(n250));
	jcb g165(.dina(w_dff_B_sNNyOCMb6_0),.dinb(n241),.dout(G863gat));
	jxor g166(.dina(w_n217_0[2]),.dinb(w_G189gat_1[1]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n252_0[2]),.dout(n253),.clk(gclk));
	jand g168(.dina(w_n223_0[0]),.dinb(w_n236_0[1]),.dout(n254),.clk(gclk));
	jcb g169(.dina(n254),.dinb(w_n228_0[0]),.dout(n255));
	jnot g170(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jcb g171(.dina(n256),.dinb(w_dff_B_wrSngEM43_1),.dout(n257));
	jcb g172(.dina(w_n255_0[0]),.dinb(w_n252_0[1]),.dout(n258));
	jand g173(.dina(n258),.dinb(w_G219gat_2[2]),.dout(n259),.clk(gclk));
	jand g174(.dina(n259),.dinb(n257),.dout(n260),.clk(gclk));
	jand g175(.dina(w_n252_0[0]),.dinb(w_G228gat_2[2]),.dout(n261),.clk(gclk));
	jand g176(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n262),.clk(gclk));
	jcb g177(.dina(n262),.dinb(w_G246gat_2[2]),.dout(n263));
	jand g178(.dina(w_dff_B_zB26315c0_0),.dinb(w_n217_0[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(w_n181_2[2]),.dinb(w_G189gat_0[2]),.dout(n265),.clk(gclk));
	jand g180(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n266),.clk(gclk));
	jand g181(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n267),.clk(gclk));
	jcb g182(.dina(n267),.dinb(n266),.dout(n268));
	jcb g183(.dina(w_dff_B_3CbSHFDQ2_0),.dinb(n265),.dout(n269));
	jcb g184(.dina(w_dff_B_vq8MgUIk5_0),.dinb(n264),.dout(n270));
	jcb g185(.dina(w_dff_B_x4SaXGzy3_0),.dinb(n261),.dout(n271));
	jcb g186(.dina(w_dff_B_66Si8Cst7_0),.dinb(n260),.dout(G864gat));
	jxor g187(.dina(w_n222_0[2]),.dinb(w_G195gat_1[1]),.dout(n273),.clk(gclk));
	jnot g188(.din(w_n273_0[2]),.dout(n274),.clk(gclk));
	jcb g189(.dina(w_dff_B_d236LyET3_0),.dinb(w_n213_0[0]),.dout(n275));
	jcb g190(.dina(w_n273_0[1]),.dinb(w_n236_0[0]),.dout(n276));
	jand g191(.dina(n276),.dinb(w_G219gat_2[1]),.dout(n277),.clk(gclk));
	jand g192(.dina(w_dff_B_Tw52TlZY2_0),.dinb(n275),.dout(n278),.clk(gclk));
	jand g193(.dina(w_n273_0[0]),.dinb(w_G228gat_2[1]),.dout(n279),.clk(gclk));
	jand g194(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n280),.clk(gclk));
	jcb g195(.dina(n280),.dinb(w_G246gat_2[1]),.dout(n281));
	jand g196(.dina(w_dff_B_aaMXyf4Z4_0),.dinb(w_n222_0[1]),.dout(n282),.clk(gclk));
	jand g197(.dina(w_n181_2[1]),.dinb(w_G195gat_0[2]),.dout(n283),.clk(gclk));
	jand g198(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n284),.clk(gclk));
	jand g199(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n285),.clk(gclk));
	jcb g200(.dina(n285),.dinb(n284),.dout(n286));
	jcb g201(.dina(w_dff_B_XFXdJ0H04_0),.dinb(n283),.dout(n287));
	jcb g202(.dina(w_dff_B_d6WLqoVw0_0),.dinb(n282),.dout(n288));
	jcb g203(.dina(w_dff_B_JLXh2En21_0),.dinb(n279),.dout(n289));
	jcb g204(.dina(w_dff_B_yUedXOTY3_0),.dinb(n278),.dout(G865gat));
	jand g205(.dina(w_n153_2[0]),.dinb(w_G91gat_0[1]),.dout(n291),.clk(gclk));
	jand g206(.dina(w_n157_0[0]),.dinb(w_G55gat_0[0]),.dout(n292),.clk(gclk));
	jand g207(.dina(w_n292_1[1]),.dinb(w_G143gat_0[0]),.dout(n293),.clk(gclk));
	jand g208(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n294),.clk(gclk));
	jand g209(.dina(w_n163_0[0]),.dinb(w_G17gat_1[0]),.dout(n295),.clk(gclk));
	jand g210(.dina(w_dff_B_adY790d46_0),.dinb(w_n162_0[0]),.dout(n296),.clk(gclk));
	jcb g211(.dina(w_n296_1[1]),.dinb(w_dff_B_xhUBfYWX6_1),.dout(n297));
	jcb g212(.dina(w_dff_B_eVBAz78o7_0),.dinb(n293),.dout(n298));
	jcb g213(.dina(n298),.dinb(n291),.dout(n299));
	jand g214(.dina(w_n299_1[1]),.dinb(w_G159gat_2[0]),.dout(n300),.clk(gclk));
	jcb g215(.dina(w_n299_1[0]),.dinb(w_G159gat_1[2]),.dout(n301));
	jand g216(.dina(w_n193_0[2]),.dinb(w_G183gat_1[0]),.dout(n302),.clk(gclk));
	jcb g217(.dina(w_n193_0[1]),.dinb(w_G183gat_0[2]),.dout(n303));
	jand g218(.dina(w_n238_0[0]),.dinb(w_n303_0[1]),.dout(n304),.clk(gclk));
	jcb g219(.dina(n304),.dinb(w_n302_0[1]),.dout(n305));
	jnot g220(.din(w_G165gat_2[0]),.dout(n306),.clk(gclk));
	jand g221(.dina(w_n153_1[2]),.dinb(w_G96gat_0[1]),.dout(n307),.clk(gclk));
	jand g222(.dina(w_n292_1[0]),.dinb(w_G146gat_0[0]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n309),.clk(gclk));
	jcb g224(.dina(w_dff_B_8hh0wXRo8_0),.dinb(w_n296_1[0]),.dout(n310));
	jcb g225(.dina(w_dff_B_EBdouLYV6_0),.dinb(n308),.dout(n311));
	jcb g226(.dina(n311),.dinb(n307),.dout(n312));
	jnot g227(.din(w_n312_1[1]),.dout(n313),.clk(gclk));
	jand g228(.dina(n313),.dinb(w_dff_B_W8XVATZZ4_1),.dout(n314),.clk(gclk));
	jnot g229(.din(n314),.dout(n315),.clk(gclk));
	jand g230(.dina(w_n153_1[1]),.dinb(w_G101gat_0[1]),.dout(n316),.clk(gclk));
	jand g231(.dina(w_n292_0[2]),.dinb(w_G149gat_0[0]),.dout(n317),.clk(gclk));
	jand g232(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n318),.clk(gclk));
	jcb g233(.dina(w_dff_B_eZOCjBFj3_0),.dinb(w_n296_0[2]),.dout(n319));
	jcb g234(.dina(w_dff_B_csxKrAiS0_0),.dinb(n317),.dout(n320));
	jcb g235(.dina(n320),.dinb(n316),.dout(n321));
	jcb g236(.dina(w_n321_1[1]),.dinb(w_G171gat_2[0]),.dout(n322));
	jand g237(.dina(w_n153_1[0]),.dinb(w_G106gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_n292_0[1]),.dinb(w_G153gat_0[0]),.dout(n324),.clk(gclk));
	jand g239(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n325),.clk(gclk));
	jcb g240(.dina(w_dff_B_SLajnLwI2_0),.dinb(w_n296_0[1]),.dout(n326));
	jcb g241(.dina(w_dff_B_XINNHBO48_0),.dinb(n324),.dout(n327));
	jcb g242(.dina(n327),.dinb(n323),.dout(n328));
	jcb g243(.dina(w_n328_1[1]),.dinb(w_G177gat_2[0]),.dout(n329));
	jand g244(.dina(w_n329_0[2]),.dinb(w_n322_0[1]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n330_0[2]),.dinb(w_n315_0[1]),.dout(n331),.clk(gclk));
	jand g246(.dina(w_n331_0[1]),.dinb(w_n305_1[1]),.dout(n332),.clk(gclk));
	jand g247(.dina(w_n312_1[0]),.dinb(w_G165gat_1[2]),.dout(n333),.clk(gclk));
	jand g248(.dina(w_n321_1[0]),.dinb(w_G171gat_1[2]),.dout(n334),.clk(gclk));
	jand g249(.dina(w_n328_1[0]),.dinb(w_G177gat_1[2]),.dout(n335),.clk(gclk));
	jand g250(.dina(w_n335_0[2]),.dinb(w_n322_0[0]),.dout(n336),.clk(gclk));
	jcb g251(.dina(n336),.dinb(w_dff_B_hdsHP5x36_1),.dout(n337));
	jand g252(.dina(w_n337_0[2]),.dinb(w_n315_0[0]),.dout(n338),.clk(gclk));
	jcb g253(.dina(n338),.dinb(w_dff_B_7qR9MaT48_1),.dout(n339));
	jcb g254(.dina(w_n339_0[1]),.dinb(n332),.dout(n340));
	jand g255(.dina(w_n340_0[1]),.dinb(w_dff_B_OK4sCdpZ2_1),.dout(n341),.clk(gclk));
	jcb g256(.dina(n341),.dinb(w_dff_B_wNHj402n7_1),.dout(G866gat));
	jnot g257(.din(w_n302_0[0]),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n303_0[0]),.dout(n344),.clk(gclk));
	jcb g259(.dina(w_n232_0[0]),.dinb(w_dff_B_narWwQcN6_1),.dout(n345));
	jand g260(.dina(n345),.dinb(w_dff_B_F7k906ye5_1),.dout(n346),.clk(gclk));
	jxor g261(.dina(w_n328_0[2]),.dinb(w_G177gat_1[1]),.dout(n347),.clk(gclk));
	jnot g262(.din(w_n347_0[2]),.dout(n348),.clk(gclk));
	jcb g263(.dina(w_dff_B_QXa92kVt9_0),.dinb(w_n346_1[1]),.dout(n349));
	jcb g264(.dina(w_n347_0[1]),.dinb(w_n305_1[0]),.dout(n350));
	jand g265(.dina(n350),.dinb(w_G219gat_2[0]),.dout(n351),.clk(gclk));
	jand g266(.dina(w_dff_B_tv4rNENE0_0),.dinb(n349),.dout(n352),.clk(gclk));
	jand g267(.dina(w_n347_0[0]),.dinb(w_G228gat_2[0]),.dout(n353),.clk(gclk));
	jand g268(.dina(w_G237gat_2[0]),.dinb(w_G177gat_1[0]),.dout(n354),.clk(gclk));
	jcb g269(.dina(n354),.dinb(w_G246gat_2[0]),.dout(n355));
	jand g270(.dina(w_dff_B_wM7xfgte6_0),.dinb(w_n328_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n181_2[0]),.dinb(w_G177gat_0[2]),.dout(n357),.clk(gclk));
	jand g272(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n358),.clk(gclk));
	jcb g273(.dina(w_dff_B_ILRiZsNh5_0),.dinb(n357),.dout(n359));
	jcb g274(.dina(w_dff_B_IfZGlIgN7_0),.dinb(n356),.dout(n360));
	jcb g275(.dina(w_dff_B_pQWVkC0d7_0),.dinb(n353),.dout(n361));
	jcb g276(.dina(w_dff_B_s1xDcGTx5_0),.dinb(n352),.dout(G874gat));
	jnot g277(.din(w_n331_0[0]),.dout(n363),.clk(gclk));
	jcb g278(.dina(w_dff_B_lS967LtZ3_0),.dinb(w_n346_1[0]),.dout(n364));
	jnot g279(.din(w_n339_0[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_dff_B_2VIeRZWQ7_0),.dinb(n364),.dout(n366),.clk(gclk));
	jxor g281(.dina(w_n299_0[2]),.dinb(w_G159gat_1[1]),.dout(n367),.clk(gclk));
	jnot g282(.din(w_n367_0[2]),.dout(n368),.clk(gclk));
	jcb g283(.dina(w_dff_B_dQ8I0KMw6_0),.dinb(n366),.dout(n369));
	jcb g284(.dina(w_n367_0[1]),.dinb(w_n340_0[0]),.dout(n370));
	jand g285(.dina(n370),.dinb(w_G219gat_1[2]),.dout(n371),.clk(gclk));
	jand g286(.dina(w_dff_B_iXQUVTDT3_0),.dinb(n369),.dout(n372),.clk(gclk));
	jand g287(.dina(w_n367_0[0]),.dinb(w_G228gat_1[2]),.dout(n373),.clk(gclk));
	jand g288(.dina(w_G237gat_1[2]),.dinb(w_G159gat_1[0]),.dout(n374),.clk(gclk));
	jcb g289(.dina(n374),.dinb(w_G246gat_1[2]),.dout(n375));
	jand g290(.dina(w_dff_B_ZoVfNSFA5_0),.dinb(w_n299_0[1]),.dout(n376),.clk(gclk));
	jand g291(.dina(w_n181_1[2]),.dinb(w_G159gat_0[2]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n378),.clk(gclk));
	jcb g293(.dina(w_dff_B_In2TtRBe7_0),.dinb(n377),.dout(n379));
	jcb g294(.dina(w_dff_B_U3LbnHYo6_0),.dinb(n376),.dout(n380));
	jcb g295(.dina(w_dff_B_P7BHgjtN7_0),.dinb(n373),.dout(n381));
	jcb g296(.dina(w_dff_B_NhgaEgBY1_0),.dinb(n372),.dout(G878gat));
	jxor g297(.dina(w_n312_0[2]),.dinb(w_G165gat_1[1]),.dout(n383),.clk(gclk));
	jnot g298(.din(w_n383_0[2]),.dout(n384),.clk(gclk));
	jnot g299(.din(w_n337_0[1]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n330_0[1]),.dout(n386),.clk(gclk));
	jcb g301(.dina(w_dff_B_Q7tIZrvg0_0),.dinb(w_n346_0[2]),.dout(n387));
	jand g302(.dina(n387),.dinb(w_dff_B_FS4S2gvY5_1),.dout(n388),.clk(gclk));
	jcb g303(.dina(n388),.dinb(w_dff_B_OmVkDI6T6_1),.dout(n389));
	jand g304(.dina(w_n330_0[0]),.dinb(w_n305_0[2]),.dout(n390),.clk(gclk));
	jcb g305(.dina(n390),.dinb(w_n337_0[0]),.dout(n391));
	jcb g306(.dina(n391),.dinb(w_n383_0[1]),.dout(n392));
	jand g307(.dina(n392),.dinb(w_G219gat_1[1]),.dout(n393),.clk(gclk));
	jand g308(.dina(w_dff_B_IFk6j4hx5_0),.dinb(n389),.dout(n394),.clk(gclk));
	jand g309(.dina(w_n383_0[0]),.dinb(w_G228gat_1[1]),.dout(n395),.clk(gclk));
	jand g310(.dina(w_G237gat_1[1]),.dinb(w_G165gat_1[0]),.dout(n396),.clk(gclk));
	jcb g311(.dina(n396),.dinb(w_G246gat_1[1]),.dout(n397));
	jand g312(.dina(w_dff_B_zUO9LkF29_0),.dinb(w_n312_0[1]),.dout(n398),.clk(gclk));
	jand g313(.dina(w_n181_1[1]),.dinb(w_G165gat_0[2]),.dout(n399),.clk(gclk));
	jand g314(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n400),.clk(gclk));
	jcb g315(.dina(w_dff_B_gJI4gtky3_0),.dinb(n399),.dout(n401));
	jcb g316(.dina(w_dff_B_uGceBSXD1_0),.dinb(n398),.dout(n402));
	jcb g317(.dina(w_dff_B_fXLA1Kwg5_0),.dinb(n395),.dout(n403));
	jcb g318(.dina(w_dff_B_DvaqvEzh1_0),.dinb(n394),.dout(G879gat));
	jxor g319(.dina(w_n321_0[2]),.dinb(w_G171gat_1[1]),.dout(n405),.clk(gclk));
	jnot g320(.din(w_n405_0[2]),.dout(n406),.clk(gclk));
	jnot g321(.din(w_n335_0[1]),.dout(n407),.clk(gclk));
	jnot g322(.din(w_n329_0[1]),.dout(n408),.clk(gclk));
	jcb g323(.dina(w_dff_B_83uWI9Ei6_0),.dinb(w_n346_0[1]),.dout(n409));
	jand g324(.dina(n409),.dinb(w_dff_B_1vPFDyg56_1),.dout(n410),.clk(gclk));
	jcb g325(.dina(n410),.dinb(w_dff_B_rXqprOXe5_1),.dout(n411));
	jand g326(.dina(w_n329_0[0]),.dinb(w_n305_0[1]),.dout(n412),.clk(gclk));
	jcb g327(.dina(n412),.dinb(w_n335_0[0]),.dout(n413));
	jcb g328(.dina(n413),.dinb(w_n405_0[1]),.dout(n414));
	jand g329(.dina(n414),.dinb(w_G219gat_1[0]),.dout(n415),.clk(gclk));
	jand g330(.dina(w_dff_B_IynLEhcC6_0),.dinb(n411),.dout(n416),.clk(gclk));
	jand g331(.dina(w_n405_0[0]),.dinb(w_G228gat_1[0]),.dout(n417),.clk(gclk));
	jand g332(.dina(w_G237gat_1[0]),.dinb(w_G171gat_1[0]),.dout(n418),.clk(gclk));
	jcb g333(.dina(n418),.dinb(w_G246gat_1[0]),.dout(n419));
	jand g334(.dina(w_dff_B_LH0q07pu1_0),.dinb(w_n321_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n181_1[0]),.dinb(w_G171gat_0[2]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jcb g337(.dina(w_dff_B_E01akAsv8_0),.dinb(n421),.dout(n423));
	jcb g338(.dina(w_dff_B_gxFDA8u96_0),.dinb(n420),.dout(n424));
	jcb g339(.dina(w_dff_B_cu1HmymM7_0),.dinb(n417),.dout(n425));
	jcb g340(.dina(w_dff_B_SLMKw8mj6_0),.dinb(n416),.dout(G880gat));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_dff_A_pbatWKxq6_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_G13gat_0[1]),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_dff_A_TQAuJOTq3_0),.doutb(w_G17gat_1[1]),.doutc(w_dff_A_Wwlk23wm8_2),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_G17gat_2[2]),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_G29gat_0[0]),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_dff_A_0XKpT3Ew1_1),.doutc(w_G42gat_0[2]),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_G42gat_1[0]),.doutb(w_dff_A_Uz76hR5G2_1),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_dff_A_A8Hsb4HS4_1),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_dff_A_9yJbgLEK7_0),.doutb(w_dff_A_NikhT9437_1),.doutc(w_G55gat_0[2]),.din(G55gat));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_G68gat_0[1]),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_dff_A_kSgMlmBC1_0),.doutb(w_G80gat_0[1]),.doutc(w_dff_A_i5nDzkmp4_2),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_dff_A_pL6PNmqM0_1),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_dff_A_OoE4TLiA8_1),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_dff_A_s6aV5ion3_1),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_GbRvA3zS6_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_dff_A_NzuKRQ147_1),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_dff_A_CimypAnj1_1),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_dff_A_lavV9sd30_0),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl jspl_w_G126gat_0(.douta(w_dff_A_lf6NpmqY2_0),.doutb(w_G126gat_0[1]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_G130gat_0[1]),.din(w_dff_B_1vBf8jKj0_2));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_G143gat_0[1]),.din(w_dff_B_jZrZfJia1_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_G146gat_0[1]),.din(w_dff_B_zbrf4LS31_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_G149gat_0[1]),.din(w_dff_B_l7oNFS4D0_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_dff_A_XwzX1IZ20_0),.doutb(w_G153gat_0[1]),.doutc(w_dff_A_rlkd52HL6_2),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_G159gat_0[1]),.doutc(w_dff_A_BeJcpQUe1_2),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_G159gat_1[0]),.doutb(w_dff_A_A7tapQ5o7_1),.doutc(w_dff_A_lTFbYbgh7_2),.din(w_G159gat_0[0]));
	jspl jspl_w_G159gat_2(.douta(w_dff_A_bs0iN9e84_0),.doutb(w_G159gat_2[1]),.din(w_G159gat_0[1]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_G165gat_0[1]),.doutc(w_dff_A_UlOMJKSX8_2),.din(G165gat));
	jspl3 jspl3_w_G165gat_1(.douta(w_G165gat_1[0]),.doutb(w_dff_A_nRO6zlfJ6_1),.doutc(w_dff_A_xpiXnAg21_2),.din(w_G165gat_0[0]));
	jspl jspl_w_G165gat_2(.douta(w_G165gat_2[0]),.doutb(w_G165gat_2[1]),.din(w_G165gat_0[1]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_dff_A_oD1Gvndw5_2),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_dff_A_pdHOZErm1_1),.doutc(w_dff_A_qLVc8urX8_2),.din(w_G171gat_0[0]));
	jspl jspl_w_G171gat_2(.douta(w_dff_A_4QdAKl7x2_0),.doutb(w_G171gat_2[1]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_G177gat_0[1]),.doutc(w_dff_A_lK7Kh6sK2_2),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_dff_A_QekXYpaX6_1),.doutc(w_dff_A_2g5bkTSe1_2),.din(w_G177gat_0[0]));
	jspl jspl_w_G177gat_2(.douta(w_dff_A_tSi1udYA9_0),.doutb(w_G177gat_2[1]),.din(w_G177gat_0[1]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_dff_A_AWuuuy1O1_2),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_dff_A_29NPMiPM0_0),.doutb(w_dff_A_B6XSKzLl1_1),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl jspl_w_G183gat_2(.douta(w_dff_A_sppNk25w3_0),.doutb(w_G183gat_2[1]),.din(w_G183gat_0[1]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_dff_A_fNGl3RZk3_2),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_dff_A_shIFNGEE6_1),.doutc(w_dff_A_xVuBfEC40_2),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_dff_A_RvVo3Sl95_0),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_dff_A_SjwLYvEt5_2),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_dff_A_PEiE3VZj4_1),.doutc(w_dff_A_MAcl6UMd6_2),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_dff_A_cckamYwI8_0),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_G201gat_0[1]),.doutc(w_dff_A_PdBieuzD8_2),.din(G201gat));
	jspl3 jspl3_w_G201gat_1(.douta(w_G201gat_1[0]),.doutb(w_dff_A_umEvOaAC1_1),.doutc(w_dff_A_1Ilctpke0_2),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G201gat_2(.douta(w_G201gat_2[0]),.doutb(w_dff_A_BrG7DVJx9_1),.doutc(w_G201gat_2[2]),.din(w_G201gat_0[1]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_4ENWc2UQ5_0),.doutb(w_G219gat_0[1]),.doutc(w_G219gat_0[2]),.din(w_dff_B_pxyp9p9L1_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_G219gat_1[0]),.doutb(w_G219gat_1[1]),.doutc(w_dff_A_oaewuqkV7_2),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_TDbxvCBp3_0),.doutb(w_G219gat_2[1]),.doutc(w_dff_A_BfEzzLk66_2),.din(w_G219gat_0[1]));
	jspl jspl_w_G219gat_3(.douta(w_dff_A_IGR0uvxD3_0),.doutb(w_G219gat_3[1]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_G228gat_0[0]),.doutb(w_G228gat_0[1]),.doutc(w_G228gat_0[2]),.din(w_dff_B_2e29grpO7_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_G228gat_2[0]),.doutb(w_G228gat_2[1]),.doutc(w_G228gat_2[2]),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_G228gat_3[1]),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_G237gat_0[0]),.doutb(w_G237gat_0[1]),.doutc(w_G237gat_0[2]),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_G237gat_2[0]),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_G237gat_3[1]),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_G246gat_0[0]),.doutb(w_G246gat_0[1]),.doutc(w_G246gat_0[2]),.din(w_dff_B_EDrNy9Qv7_3));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_G246gat_2[0]),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_G246gat_3[1]),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_dff_A_EvZfo1l24_0),.doutb(w_dff_A_nlLGuuQ96_1),.doutc(w_G261gat_0[2]),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_G390gat_0[1]),.doutc(G390gat),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_G447gat_0[2]),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(G447gat),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n96_0(.douta(w_dff_A_h23fIEli9_0),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_dff_A_2UdM7RhN4_1),.din(n98));
	jspl jspl_w_n99_0(.douta(w_dff_A_rDQOP6sh4_0),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_dff_A_CCj0la7k5_1),.din(n101));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl jspl_w_n106_0(.douta(w_n106_0[0]),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n118_0(.douta(w_dff_A_iJ7ti8ja8_0),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl jspl_w_n121_0(.douta(w_dff_A_rroH0NRy0_0),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n143_0(.douta(w_dff_A_OICYdldO3_0),.doutb(w_n143_0[1]),.din(w_dff_B_rqeHkNQs4_2));
	jspl jspl_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.din(n149));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.doutc(w_n153_1[2]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n153_2(.douta(w_n153_2[0]),.doutb(w_n153_2[1]),.doutc(w_n153_2[2]),.din(w_n153_0[1]));
	jspl jspl_w_n153_3(.douta(w_n153_3[0]),.doutb(w_n153_3[1]),.din(w_n153_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(n154));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_LjJcmoBW0_1),.doutc(w_dff_A_fgfiDB7k9_2),.din(n165));
	jspl3 jspl3_w_n165_1(.douta(w_n165_1[0]),.doutb(w_dff_A_u0OO4cb02_1),.doutc(w_dff_A_BY2TtJ9M2_2),.din(w_n165_0[0]));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.doutc(w_n167_0[2]),.din(n167));
	jspl jspl_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n181_2(.douta(w_n181_2[0]),.doutb(w_n181_2[1]),.doutc(w_n181_2[2]),.din(w_n181_0[1]));
	jspl jspl_w_n181_3(.douta(w_n181_3[0]),.doutb(w_n181_3[1]),.din(w_n181_0[2]));
	jspl3 jspl3_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.doutc(w_n193_0[2]),.din(n193));
	jspl jspl_w_n193_1(.douta(w_n193_1[0]),.doutb(w_n193_1[1]),.din(w_n193_0[0]));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_dff_A_fRiY1ZxT2_1),.doutc(w_n194_0[2]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.din(n196));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl jspl_w_n217_1(.douta(w_n217_1[0]),.doutb(w_n217_1[1]),.din(w_n217_0[0]));
	jspl jspl_w_n218_0(.douta(w_dff_A_XbNcbaxR3_0),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.doutc(w_n222_0[2]),.din(n222));
	jspl jspl_w_n222_1(.douta(w_n222_1[0]),.doutb(w_n222_1[1]),.din(w_n222_0[0]));
	jspl jspl_w_n223_0(.douta(w_dff_A_PNKwbeGg8_0),.doutb(w_n223_0[1]),.din(n223));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n228_0(.douta(w_dff_A_V8hvUBDX6_0),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.din(n230));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.doutc(w_n236_0[2]),.din(n236));
	jspl jspl_w_n238_0(.douta(w_n238_0[0]),.doutb(w_n238_0[1]),.din(n238));
	jspl3 jspl3_w_n252_0(.douta(w_n252_0[0]),.doutb(w_dff_A_ZIMMHt8I0_1),.doutc(w_n252_0[2]),.din(n252));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.doutc(w_n273_0[2]),.din(n273));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl jspl_w_n292_1(.douta(w_n292_1[0]),.doutb(w_n292_1[1]),.din(w_n292_0[0]));
	jspl3 jspl3_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.doutc(w_n296_0[2]),.din(n296));
	jspl jspl_w_n296_1(.douta(w_n296_1[0]),.doutb(w_n296_1[1]),.din(w_n296_0[0]));
	jspl3 jspl3_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.doutc(w_n299_0[2]),.din(n299));
	jspl jspl_w_n299_1(.douta(w_n299_1[0]),.doutb(w_n299_1[1]),.din(w_n299_0[0]));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_dff_A_fq5Nvc0t6_1),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_zL7JR5nd9_1),.din(n303));
	jspl3 jspl3_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.doutc(w_n305_0[2]),.din(n305));
	jspl jspl_w_n305_1(.douta(w_n305_1[0]),.doutb(w_dff_A_xdJBDRS58_1),.din(w_n305_0[0]));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl3 jspl3_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.doutc(w_n321_0[2]),.din(n321));
	jspl jspl_w_n321_1(.douta(w_n321_1[0]),.doutb(w_n321_1[1]),.din(w_n321_0[0]));
	jspl jspl_w_n322_0(.douta(w_dff_A_OrTZDfrS0_0),.doutb(w_n322_0[1]),.din(n322));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n328_1(.douta(w_n328_1[0]),.doutb(w_n328_1[1]),.din(w_n328_0[0]));
	jspl3 jspl3_w_n329_0(.douta(w_dff_A_EfEh2nT13_0),.doutb(w_n329_0[1]),.doutc(w_n329_0[2]),.din(n329));
	jspl3 jspl3_w_n330_0(.douta(w_dff_A_w6cCnhXf2_0),.doutb(w_n330_0[1]),.doutc(w_dff_A_LR4Lx2Rl6_2),.din(n330));
	jspl jspl_w_n331_0(.douta(w_n331_0[0]),.doutb(w_n331_0[1]),.din(n331));
	jspl3 jspl3_w_n335_0(.douta(w_dff_A_HLFM1v4Q5_0),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n337_0(.douta(w_dff_A_jXjURwr55_0),.doutb(w_n337_0[1]),.doutc(w_dff_A_1eFlQMwc5_2),.din(n337));
	jspl jspl_w_n339_0(.douta(w_n339_0[0]),.doutb(w_dff_A_xhaf7J6J9_1),.din(n339));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n347_0(.douta(w_n347_0[0]),.doutb(w_dff_A_JHrFwDUc3_1),.doutc(w_n347_0[2]),.din(n347));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_dff_A_bdFAh50x8_1),.doutc(w_n367_0[2]),.din(n367));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_dff_A_26T9gUqU7_1),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_dff_A_hZVUsbC05_1),.doutc(w_n405_0[2]),.din(n405));
	jdff dff_A_CCj0la7k5_1(.dout(w_n101_0[1]),.din(w_dff_A_CCj0la7k5_1),.clk(gclk));
	jdff dff_A_rDQOP6sh4_0(.dout(w_n99_0[0]),.din(w_dff_A_rDQOP6sh4_0),.clk(gclk));
	jdff dff_B_LJ2LtJgT0_0(.din(n119),.dout(w_dff_B_LJ2LtJgT0_0),.clk(gclk));
	jdff dff_B_C3ikhOSA3_1(.din(G74gat),.dout(w_dff_B_C3ikhOSA3_1),.clk(gclk));
	jdff dff_B_vrtHSlZA2_0(.din(n131),.dout(w_dff_B_vrtHSlZA2_0),.clk(gclk));
	jdff dff_B_J83LNMHI6_1(.din(G135gat),.dout(w_dff_B_J83LNMHI6_1),.clk(gclk));
	jdff dff_B_JeFLVpOz7_0(.din(n127),.dout(w_dff_B_JeFLVpOz7_0),.clk(gclk));
	jdff dff_B_rxMu0aUu8_0(.din(n140),.dout(w_dff_B_rxMu0aUu8_0),.clk(gclk));
	jdff dff_B_FK76auAP9_1(.din(G207gat),.dout(w_dff_B_FK76auAP9_1),.clk(gclk));
	jdff dff_B_ngv4l5OW7_0(.din(n136),.dout(w_dff_B_ngv4l5OW7_0),.clk(gclk));
	jdff dff_B_1vBf8jKj0_2(.din(G130gat),.dout(w_dff_B_1vBf8jKj0_2),.clk(gclk));
	jdff dff_B_xAVV3AjK3_0(.din(n188),.dout(w_dff_B_xAVV3AjK3_0),.clk(gclk));
	jdff dff_B_2xbdBfGN0_0(.din(n187),.dout(w_dff_B_2xbdBfGN0_0),.clk(gclk));
	jdff dff_B_ftLDdwzc9_0(.din(n186),.dout(w_dff_B_ftLDdwzc9_0),.clk(gclk));
	jdff dff_B_szDRvvjH5_0(.din(n185),.dout(w_dff_B_szDRvvjH5_0),.clk(gclk));
	jdff dff_B_Clg6Up0v0_0(.din(w_dff_B_szDRvvjH5_0),.dout(w_dff_B_Clg6Up0v0_0),.clk(gclk));
	jdff dff_B_n7iFbRDd4_0(.din(w_dff_B_Clg6Up0v0_0),.dout(w_dff_B_n7iFbRDd4_0),.clk(gclk));
	jdff dff_B_PC7QqtZB8_0(.din(w_dff_B_n7iFbRDd4_0),.dout(w_dff_B_PC7QqtZB8_0),.clk(gclk));
	jdff dff_B_NUiyhTX28_0(.din(n176),.dout(w_dff_B_NUiyhTX28_0),.clk(gclk));
	jdff dff_B_FUh0rxZd4_0(.din(w_dff_B_NUiyhTX28_0),.dout(w_dff_B_FUh0rxZd4_0),.clk(gclk));
	jdff dff_B_EmdG73Tw1_0(.din(w_dff_B_FUh0rxZd4_0),.dout(w_dff_B_EmdG73Tw1_0),.clk(gclk));
	jdff dff_B_dUrOWA1l6_0(.din(w_dff_B_EmdG73Tw1_0),.dout(w_dff_B_dUrOWA1l6_0),.clk(gclk));
	jdff dff_A_S8dJ1eao0_1(.dout(w_G201gat_2[1]),.din(w_dff_A_S8dJ1eao0_1),.clk(gclk));
	jdff dff_A_lEctacaT4_1(.dout(w_dff_A_S8dJ1eao0_1),.din(w_dff_A_lEctacaT4_1),.clk(gclk));
	jdff dff_A_ldmCPNlp5_1(.dout(w_dff_A_lEctacaT4_1),.din(w_dff_A_ldmCPNlp5_1),.clk(gclk));
	jdff dff_A_5oV02g2c4_1(.dout(w_dff_A_ldmCPNlp5_1),.din(w_dff_A_5oV02g2c4_1),.clk(gclk));
	jdff dff_A_BrG7DVJx9_1(.dout(w_dff_A_5oV02g2c4_1),.din(w_dff_A_BrG7DVJx9_1),.clk(gclk));
	jdff dff_B_jAkB14bt6_0(.din(n250),.dout(w_dff_B_jAkB14bt6_0),.clk(gclk));
	jdff dff_B_ZDVyxVTw8_0(.din(w_dff_B_jAkB14bt6_0),.dout(w_dff_B_ZDVyxVTw8_0),.clk(gclk));
	jdff dff_B_RmpHZQsp4_0(.din(w_dff_B_ZDVyxVTw8_0),.dout(w_dff_B_RmpHZQsp4_0),.clk(gclk));
	jdff dff_B_sNNyOCMb6_0(.din(w_dff_B_RmpHZQsp4_0),.dout(w_dff_B_sNNyOCMb6_0),.clk(gclk));
	jdff dff_B_vOp2ltun6_0(.din(n249),.dout(w_dff_B_vOp2ltun6_0),.clk(gclk));
	jdff dff_B_6JdlWv7H4_0(.din(n248),.dout(w_dff_B_6JdlWv7H4_0),.clk(gclk));
	jdff dff_B_lurEB3A76_0(.din(n247),.dout(w_dff_B_lurEB3A76_0),.clk(gclk));
	jdff dff_B_PLP1zwJM5_0(.din(w_dff_B_lurEB3A76_0),.dout(w_dff_B_PLP1zwJM5_0),.clk(gclk));
	jdff dff_B_IBnFkczI7_0(.din(w_dff_B_PLP1zwJM5_0),.dout(w_dff_B_IBnFkczI7_0),.clk(gclk));
	jdff dff_B_MQWdLDRe1_0(.din(w_dff_B_IBnFkczI7_0),.dout(w_dff_B_MQWdLDRe1_0),.clk(gclk));
	jdff dff_B_jlwOerqR1_0(.din(n244),.dout(w_dff_B_jlwOerqR1_0),.clk(gclk));
	jdff dff_B_Lan5YEWw0_0(.din(w_dff_B_jlwOerqR1_0),.dout(w_dff_B_Lan5YEWw0_0),.clk(gclk));
	jdff dff_B_Xjh5BrIx2_0(.din(w_dff_B_Lan5YEWw0_0),.dout(w_dff_B_Xjh5BrIx2_0),.clk(gclk));
	jdff dff_B_HXyGwlXN3_0(.din(w_dff_B_Xjh5BrIx2_0),.dout(w_dff_B_HXyGwlXN3_0),.clk(gclk));
	jdff dff_B_lZn1Q91d1_0(.din(n240),.dout(w_dff_B_lZn1Q91d1_0),.clk(gclk));
	jdff dff_B_51qpWO1A7_0(.din(w_dff_B_lZn1Q91d1_0),.dout(w_dff_B_51qpWO1A7_0),.clk(gclk));
	jdff dff_A_IGR0uvxD3_0(.dout(w_G219gat_3[0]),.din(w_dff_A_IGR0uvxD3_0),.clk(gclk));
	jdff dff_B_2zxUmpFN8_1(.din(n195),.dout(w_dff_B_2zxUmpFN8_1),.clk(gclk));
	jdff dff_B_Z6LMu0yv2_1(.din(w_dff_B_2zxUmpFN8_1),.dout(w_dff_B_Z6LMu0yv2_1),.clk(gclk));
	jdff dff_B_0x0VDcFI8_1(.din(w_dff_B_Z6LMu0yv2_1),.dout(w_dff_B_0x0VDcFI8_1),.clk(gclk));
	jdff dff_A_fRiY1ZxT2_1(.dout(w_n194_0[1]),.din(w_dff_A_fRiY1ZxT2_1),.clk(gclk));
	jdff dff_A_wfXCmYf12_0(.dout(w_G183gat_2[0]),.din(w_dff_A_wfXCmYf12_0),.clk(gclk));
	jdff dff_A_iY15mJi56_0(.dout(w_dff_A_wfXCmYf12_0),.din(w_dff_A_iY15mJi56_0),.clk(gclk));
	jdff dff_A_HkLKhpge1_0(.dout(w_dff_A_iY15mJi56_0),.din(w_dff_A_HkLKhpge1_0),.clk(gclk));
	jdff dff_A_BdOGBBQ45_0(.dout(w_dff_A_HkLKhpge1_0),.din(w_dff_A_BdOGBBQ45_0),.clk(gclk));
	jdff dff_A_sppNk25w3_0(.dout(w_dff_A_BdOGBBQ45_0),.din(w_dff_A_sppNk25w3_0),.clk(gclk));
	jdff dff_B_q2wRB0Pm0_0(.din(n271),.dout(w_dff_B_q2wRB0Pm0_0),.clk(gclk));
	jdff dff_B_66Si8Cst7_0(.din(w_dff_B_q2wRB0Pm0_0),.dout(w_dff_B_66Si8Cst7_0),.clk(gclk));
	jdff dff_B_x4SaXGzy3_0(.din(n270),.dout(w_dff_B_x4SaXGzy3_0),.clk(gclk));
	jdff dff_B_vq8MgUIk5_0(.din(n269),.dout(w_dff_B_vq8MgUIk5_0),.clk(gclk));
	jdff dff_B_rVJolAeM7_0(.din(n268),.dout(w_dff_B_rVJolAeM7_0),.clk(gclk));
	jdff dff_B_u835j7zb2_0(.din(w_dff_B_rVJolAeM7_0),.dout(w_dff_B_u835j7zb2_0),.clk(gclk));
	jdff dff_B_L2msWCfY5_0(.din(w_dff_B_u835j7zb2_0),.dout(w_dff_B_L2msWCfY5_0),.clk(gclk));
	jdff dff_B_3CbSHFDQ2_0(.din(w_dff_B_L2msWCfY5_0),.dout(w_dff_B_3CbSHFDQ2_0),.clk(gclk));
	jdff dff_B_IYYquxY82_0(.din(n263),.dout(w_dff_B_IYYquxY82_0),.clk(gclk));
	jdff dff_B_wFk9ZHSg1_0(.din(w_dff_B_IYYquxY82_0),.dout(w_dff_B_wFk9ZHSg1_0),.clk(gclk));
	jdff dff_B_8wj4ljoW5_0(.din(w_dff_B_wFk9ZHSg1_0),.dout(w_dff_B_8wj4ljoW5_0),.clk(gclk));
	jdff dff_B_zB26315c0_0(.din(w_dff_B_8wj4ljoW5_0),.dout(w_dff_B_zB26315c0_0),.clk(gclk));
	jdff dff_B_wrSngEM43_1(.din(n253),.dout(w_dff_B_wrSngEM43_1),.clk(gclk));
	jdff dff_A_ZIMMHt8I0_1(.dout(w_n252_0[1]),.din(w_dff_A_ZIMMHt8I0_1),.clk(gclk));
	jdff dff_B_q30TG8ee0_0(.din(n289),.dout(w_dff_B_q30TG8ee0_0),.clk(gclk));
	jdff dff_B_y3vZdYAA7_0(.din(w_dff_B_q30TG8ee0_0),.dout(w_dff_B_y3vZdYAA7_0),.clk(gclk));
	jdff dff_B_yUedXOTY3_0(.din(w_dff_B_y3vZdYAA7_0),.dout(w_dff_B_yUedXOTY3_0),.clk(gclk));
	jdff dff_B_JLXh2En21_0(.din(n288),.dout(w_dff_B_JLXh2En21_0),.clk(gclk));
	jdff dff_B_d6WLqoVw0_0(.din(n287),.dout(w_dff_B_d6WLqoVw0_0),.clk(gclk));
	jdff dff_B_sIA58gZx8_0(.din(n286),.dout(w_dff_B_sIA58gZx8_0),.clk(gclk));
	jdff dff_B_wX6ngeO32_0(.din(w_dff_B_sIA58gZx8_0),.dout(w_dff_B_wX6ngeO32_0),.clk(gclk));
	jdff dff_B_wMtcj9Wr3_0(.din(w_dff_B_wX6ngeO32_0),.dout(w_dff_B_wMtcj9Wr3_0),.clk(gclk));
	jdff dff_B_XFXdJ0H04_0(.din(w_dff_B_wMtcj9Wr3_0),.dout(w_dff_B_XFXdJ0H04_0),.clk(gclk));
	jdff dff_B_YoxmnRGE2_0(.din(n281),.dout(w_dff_B_YoxmnRGE2_0),.clk(gclk));
	jdff dff_B_lWefJEvt2_0(.din(w_dff_B_YoxmnRGE2_0),.dout(w_dff_B_lWefJEvt2_0),.clk(gclk));
	jdff dff_B_lojKx3UP5_0(.din(w_dff_B_lWefJEvt2_0),.dout(w_dff_B_lojKx3UP5_0),.clk(gclk));
	jdff dff_B_aaMXyf4Z4_0(.din(w_dff_B_lojKx3UP5_0),.dout(w_dff_B_aaMXyf4Z4_0),.clk(gclk));
	jdff dff_B_hYgvfGge0_0(.din(n277),.dout(w_dff_B_hYgvfGge0_0),.clk(gclk));
	jdff dff_B_Tw52TlZY2_0(.din(w_dff_B_hYgvfGge0_0),.dout(w_dff_B_Tw52TlZY2_0),.clk(gclk));
	jdff dff_B_jwevzxdE7_0(.din(n274),.dout(w_dff_B_jwevzxdE7_0),.clk(gclk));
	jdff dff_B_d236LyET3_0(.din(w_dff_B_jwevzxdE7_0),.dout(w_dff_B_d236LyET3_0),.clk(gclk));
	jdff dff_B_DaR8gZ0e4_1(.din(n300),.dout(w_dff_B_DaR8gZ0e4_1),.clk(gclk));
	jdff dff_B_GOIu13tQ6_1(.din(w_dff_B_DaR8gZ0e4_1),.dout(w_dff_B_GOIu13tQ6_1),.clk(gclk));
	jdff dff_B_udC7DLF52_1(.din(w_dff_B_GOIu13tQ6_1),.dout(w_dff_B_udC7DLF52_1),.clk(gclk));
	jdff dff_B_Twib4wUK2_1(.din(w_dff_B_udC7DLF52_1),.dout(w_dff_B_Twib4wUK2_1),.clk(gclk));
	jdff dff_B_wNHj402n7_1(.din(w_dff_B_Twib4wUK2_1),.dout(w_dff_B_wNHj402n7_1),.clk(gclk));
	jdff dff_B_hW3SXoDk1_1(.din(n301),.dout(w_dff_B_hW3SXoDk1_1),.clk(gclk));
	jdff dff_B_8HssfsbQ3_1(.din(w_dff_B_hW3SXoDk1_1),.dout(w_dff_B_8HssfsbQ3_1),.clk(gclk));
	jdff dff_B_gJILkU1J6_1(.din(w_dff_B_8HssfsbQ3_1),.dout(w_dff_B_gJILkU1J6_1),.clk(gclk));
	jdff dff_B_WNOlCCmX6_1(.din(w_dff_B_gJILkU1J6_1),.dout(w_dff_B_WNOlCCmX6_1),.clk(gclk));
	jdff dff_B_OK4sCdpZ2_1(.din(w_dff_B_WNOlCCmX6_1),.dout(w_dff_B_OK4sCdpZ2_1),.clk(gclk));
	jdff dff_A_krnsjryp8_0(.dout(w_G159gat_2[0]),.din(w_dff_A_krnsjryp8_0),.clk(gclk));
	jdff dff_A_LNLuCyBO1_0(.dout(w_dff_A_krnsjryp8_0),.din(w_dff_A_LNLuCyBO1_0),.clk(gclk));
	jdff dff_A_0QBMoMtA3_0(.dout(w_dff_A_LNLuCyBO1_0),.din(w_dff_A_0QBMoMtA3_0),.clk(gclk));
	jdff dff_A_Qis3FsmZ9_0(.dout(w_dff_A_0QBMoMtA3_0),.din(w_dff_A_Qis3FsmZ9_0),.clk(gclk));
	jdff dff_A_bs0iN9e84_0(.dout(w_dff_A_Qis3FsmZ9_0),.din(w_dff_A_bs0iN9e84_0),.clk(gclk));
	jdff dff_B_DInSCSrx2_0(.din(n361),.dout(w_dff_B_DInSCSrx2_0),.clk(gclk));
	jdff dff_B_aAzmz2sh9_0(.din(w_dff_B_DInSCSrx2_0),.dout(w_dff_B_aAzmz2sh9_0),.clk(gclk));
	jdff dff_B_cuMCaWMG5_0(.din(w_dff_B_aAzmz2sh9_0),.dout(w_dff_B_cuMCaWMG5_0),.clk(gclk));
	jdff dff_B_Sz9vkcB09_0(.din(w_dff_B_cuMCaWMG5_0),.dout(w_dff_B_Sz9vkcB09_0),.clk(gclk));
	jdff dff_B_s1xDcGTx5_0(.din(w_dff_B_Sz9vkcB09_0),.dout(w_dff_B_s1xDcGTx5_0),.clk(gclk));
	jdff dff_B_pQWVkC0d7_0(.din(n360),.dout(w_dff_B_pQWVkC0d7_0),.clk(gclk));
	jdff dff_B_IfZGlIgN7_0(.din(n359),.dout(w_dff_B_IfZGlIgN7_0),.clk(gclk));
	jdff dff_B_Rb809NdJ9_0(.din(n358),.dout(w_dff_B_Rb809NdJ9_0),.clk(gclk));
	jdff dff_B_plBa4Teo8_0(.din(w_dff_B_Rb809NdJ9_0),.dout(w_dff_B_plBa4Teo8_0),.clk(gclk));
	jdff dff_B_nEEZhE1q7_0(.din(w_dff_B_plBa4Teo8_0),.dout(w_dff_B_nEEZhE1q7_0),.clk(gclk));
	jdff dff_B_ILRiZsNh5_0(.din(w_dff_B_nEEZhE1q7_0),.dout(w_dff_B_ILRiZsNh5_0),.clk(gclk));
	jdff dff_B_tFldBsGg2_0(.din(n355),.dout(w_dff_B_tFldBsGg2_0),.clk(gclk));
	jdff dff_B_n42kkEU89_0(.din(w_dff_B_tFldBsGg2_0),.dout(w_dff_B_n42kkEU89_0),.clk(gclk));
	jdff dff_B_KnECL4Uk8_0(.din(w_dff_B_n42kkEU89_0),.dout(w_dff_B_KnECL4Uk8_0),.clk(gclk));
	jdff dff_B_wM7xfgte6_0(.din(w_dff_B_KnECL4Uk8_0),.dout(w_dff_B_wM7xfgte6_0),.clk(gclk));
	jdff dff_B_mVkx3Uhu7_0(.din(n351),.dout(w_dff_B_mVkx3Uhu7_0),.clk(gclk));
	jdff dff_B_tv4rNENE0_0(.din(w_dff_B_mVkx3Uhu7_0),.dout(w_dff_B_tv4rNENE0_0),.clk(gclk));
	jdff dff_A_a9YVctBP1_0(.dout(w_G219gat_2[0]),.din(w_dff_A_a9YVctBP1_0),.clk(gclk));
	jdff dff_A_TDbxvCBp3_0(.dout(w_dff_A_a9YVctBP1_0),.din(w_dff_A_TDbxvCBp3_0),.clk(gclk));
	jdff dff_A_BfEzzLk66_2(.dout(w_G219gat_2[2]),.din(w_dff_A_BfEzzLk66_2),.clk(gclk));
	jdff dff_B_XLilWEjK9_0(.din(n348),.dout(w_dff_B_XLilWEjK9_0),.clk(gclk));
	jdff dff_B_lHIcKZeN7_0(.din(w_dff_B_XLilWEjK9_0),.dout(w_dff_B_lHIcKZeN7_0),.clk(gclk));
	jdff dff_B_yVRaUIFk9_0(.din(w_dff_B_lHIcKZeN7_0),.dout(w_dff_B_yVRaUIFk9_0),.clk(gclk));
	jdff dff_B_QXa92kVt9_0(.din(w_dff_B_yVRaUIFk9_0),.dout(w_dff_B_QXa92kVt9_0),.clk(gclk));
	jdff dff_A_xZkURrot5_1(.dout(w_n347_0[1]),.din(w_dff_A_xZkURrot5_1),.clk(gclk));
	jdff dff_A_JHrFwDUc3_1(.dout(w_dff_A_xZkURrot5_1),.din(w_dff_A_JHrFwDUc3_1),.clk(gclk));
	jdff dff_B_B0T2Q3Bw1_0(.din(n381),.dout(w_dff_B_B0T2Q3Bw1_0),.clk(gclk));
	jdff dff_B_CHonst4n9_0(.din(w_dff_B_B0T2Q3Bw1_0),.dout(w_dff_B_CHonst4n9_0),.clk(gclk));
	jdff dff_B_pgUV00sw9_0(.din(w_dff_B_CHonst4n9_0),.dout(w_dff_B_pgUV00sw9_0),.clk(gclk));
	jdff dff_B_Emc52eko9_0(.din(w_dff_B_pgUV00sw9_0),.dout(w_dff_B_Emc52eko9_0),.clk(gclk));
	jdff dff_B_7PfSUxZl2_0(.din(w_dff_B_Emc52eko9_0),.dout(w_dff_B_7PfSUxZl2_0),.clk(gclk));
	jdff dff_B_NhgaEgBY1_0(.din(w_dff_B_7PfSUxZl2_0),.dout(w_dff_B_NhgaEgBY1_0),.clk(gclk));
	jdff dff_B_P7BHgjtN7_0(.din(n380),.dout(w_dff_B_P7BHgjtN7_0),.clk(gclk));
	jdff dff_B_U3LbnHYo6_0(.din(n379),.dout(w_dff_B_U3LbnHYo6_0),.clk(gclk));
	jdff dff_B_nCR9WiLN1_0(.din(n378),.dout(w_dff_B_nCR9WiLN1_0),.clk(gclk));
	jdff dff_B_3e0Ei4UV6_0(.din(w_dff_B_nCR9WiLN1_0),.dout(w_dff_B_3e0Ei4UV6_0),.clk(gclk));
	jdff dff_B_OLlmtcHD2_0(.din(w_dff_B_3e0Ei4UV6_0),.dout(w_dff_B_OLlmtcHD2_0),.clk(gclk));
	jdff dff_B_In2TtRBe7_0(.din(w_dff_B_OLlmtcHD2_0),.dout(w_dff_B_In2TtRBe7_0),.clk(gclk));
	jdff dff_B_LUMsYR5l2_0(.din(n375),.dout(w_dff_B_LUMsYR5l2_0),.clk(gclk));
	jdff dff_B_bO7wV32L2_0(.din(w_dff_B_LUMsYR5l2_0),.dout(w_dff_B_bO7wV32L2_0),.clk(gclk));
	jdff dff_B_Gqut33oe7_0(.din(w_dff_B_bO7wV32L2_0),.dout(w_dff_B_Gqut33oe7_0),.clk(gclk));
	jdff dff_B_ZoVfNSFA5_0(.din(w_dff_B_Gqut33oe7_0),.dout(w_dff_B_ZoVfNSFA5_0),.clk(gclk));
	jdff dff_B_iXQUVTDT3_0(.din(n371),.dout(w_dff_B_iXQUVTDT3_0),.clk(gclk));
	jdff dff_A_xdJBDRS58_1(.dout(w_n305_1[1]),.din(w_dff_A_xdJBDRS58_1),.clk(gclk));
	jdff dff_B_wLgqbGeo6_0(.din(n368),.dout(w_dff_B_wLgqbGeo6_0),.clk(gclk));
	jdff dff_B_KM37Jo824_0(.din(w_dff_B_wLgqbGeo6_0),.dout(w_dff_B_KM37Jo824_0),.clk(gclk));
	jdff dff_B_cr0COvcA3_0(.din(w_dff_B_KM37Jo824_0),.dout(w_dff_B_cr0COvcA3_0),.clk(gclk));
	jdff dff_B_9Zomai555_0(.din(w_dff_B_cr0COvcA3_0),.dout(w_dff_B_9Zomai555_0),.clk(gclk));
	jdff dff_B_dQ8I0KMw6_0(.din(w_dff_B_9Zomai555_0),.dout(w_dff_B_dQ8I0KMw6_0),.clk(gclk));
	jdff dff_A_2dSaeeMX2_1(.dout(w_n367_0[1]),.din(w_dff_A_2dSaeeMX2_1),.clk(gclk));
	jdff dff_A_SvWCnciy3_1(.dout(w_dff_A_2dSaeeMX2_1),.din(w_dff_A_SvWCnciy3_1),.clk(gclk));
	jdff dff_A_gq5DHJoV3_1(.dout(w_dff_A_SvWCnciy3_1),.din(w_dff_A_gq5DHJoV3_1),.clk(gclk));
	jdff dff_A_bdFAh50x8_1(.dout(w_dff_A_gq5DHJoV3_1),.din(w_dff_A_bdFAh50x8_1),.clk(gclk));
	jdff dff_B_eVBAz78o7_0(.din(n297),.dout(w_dff_B_eVBAz78o7_0),.clk(gclk));
	jdff dff_B_XZ64hbkZ4_1(.din(n294),.dout(w_dff_B_XZ64hbkZ4_1),.clk(gclk));
	jdff dff_B_T0dq7uGJ3_1(.din(w_dff_B_XZ64hbkZ4_1),.dout(w_dff_B_T0dq7uGJ3_1),.clk(gclk));
	jdff dff_B_xhUBfYWX6_1(.din(w_dff_B_T0dq7uGJ3_1),.dout(w_dff_B_xhUBfYWX6_1),.clk(gclk));
	jdff dff_A_Ij6H6NcE8_1(.dout(w_G159gat_1[1]),.din(w_dff_A_Ij6H6NcE8_1),.clk(gclk));
	jdff dff_A_dmDOKtie0_1(.dout(w_dff_A_Ij6H6NcE8_1),.din(w_dff_A_dmDOKtie0_1),.clk(gclk));
	jdff dff_A_CVDJVjub8_1(.dout(w_dff_A_dmDOKtie0_1),.din(w_dff_A_CVDJVjub8_1),.clk(gclk));
	jdff dff_A_JaA2xSVq2_1(.dout(w_dff_A_CVDJVjub8_1),.din(w_dff_A_JaA2xSVq2_1),.clk(gclk));
	jdff dff_A_A7tapQ5o7_1(.dout(w_dff_A_JaA2xSVq2_1),.din(w_dff_A_A7tapQ5o7_1),.clk(gclk));
	jdff dff_A_9mTDFcAW3_2(.dout(w_G159gat_1[2]),.din(w_dff_A_9mTDFcAW3_2),.clk(gclk));
	jdff dff_A_gTPJyhz25_2(.dout(w_dff_A_9mTDFcAW3_2),.din(w_dff_A_gTPJyhz25_2),.clk(gclk));
	jdff dff_A_MvHYnNG52_2(.dout(w_dff_A_gTPJyhz25_2),.din(w_dff_A_MvHYnNG52_2),.clk(gclk));
	jdff dff_A_Ecd11qi83_2(.dout(w_dff_A_MvHYnNG52_2),.din(w_dff_A_Ecd11qi83_2),.clk(gclk));
	jdff dff_A_lTFbYbgh7_2(.dout(w_dff_A_Ecd11qi83_2),.din(w_dff_A_lTFbYbgh7_2),.clk(gclk));
	jdff dff_A_FWdANqlu2_2(.dout(w_G159gat_0[2]),.din(w_dff_A_FWdANqlu2_2),.clk(gclk));
	jdff dff_A_e72YSGre0_2(.dout(w_dff_A_FWdANqlu2_2),.din(w_dff_A_e72YSGre0_2),.clk(gclk));
	jdff dff_A_PonThVdN3_2(.dout(w_dff_A_e72YSGre0_2),.din(w_dff_A_PonThVdN3_2),.clk(gclk));
	jdff dff_A_BeJcpQUe1_2(.dout(w_dff_A_PonThVdN3_2),.din(w_dff_A_BeJcpQUe1_2),.clk(gclk));
	jdff dff_B_2VIeRZWQ7_0(.din(n365),.dout(w_dff_B_2VIeRZWQ7_0),.clk(gclk));
	jdff dff_A_xhaf7J6J9_1(.dout(w_n339_0[1]),.din(w_dff_A_xhaf7J6J9_1),.clk(gclk));
	jdff dff_B_e37gPooD5_1(.din(n333),.dout(w_dff_B_e37gPooD5_1),.clk(gclk));
	jdff dff_B_fwDGZ7am9_1(.din(w_dff_B_e37gPooD5_1),.dout(w_dff_B_fwDGZ7am9_1),.clk(gclk));
	jdff dff_B_7qR9MaT48_1(.din(w_dff_B_fwDGZ7am9_1),.dout(w_dff_B_7qR9MaT48_1),.clk(gclk));
	jdff dff_B_lS967LtZ3_0(.din(n363),.dout(w_dff_B_lS967LtZ3_0),.clk(gclk));
	jdff dff_B_m7gNxFhF7_1(.din(n306),.dout(w_dff_B_m7gNxFhF7_1),.clk(gclk));
	jdff dff_B_5ZRBshz49_1(.din(w_dff_B_m7gNxFhF7_1),.dout(w_dff_B_5ZRBshz49_1),.clk(gclk));
	jdff dff_B_IfKNjEif3_1(.din(w_dff_B_5ZRBshz49_1),.dout(w_dff_B_IfKNjEif3_1),.clk(gclk));
	jdff dff_B_ESHZQwp54_1(.din(w_dff_B_IfKNjEif3_1),.dout(w_dff_B_ESHZQwp54_1),.clk(gclk));
	jdff dff_B_W8XVATZZ4_1(.din(w_dff_B_ESHZQwp54_1),.dout(w_dff_B_W8XVATZZ4_1),.clk(gclk));
	jdff dff_B_55b2vjm40_0(.din(n403),.dout(w_dff_B_55b2vjm40_0),.clk(gclk));
	jdff dff_B_shj27mWZ2_0(.din(w_dff_B_55b2vjm40_0),.dout(w_dff_B_shj27mWZ2_0),.clk(gclk));
	jdff dff_B_dKUX8KWL8_0(.din(w_dff_B_shj27mWZ2_0),.dout(w_dff_B_dKUX8KWL8_0),.clk(gclk));
	jdff dff_B_WDvzYpgM8_0(.din(w_dff_B_dKUX8KWL8_0),.dout(w_dff_B_WDvzYpgM8_0),.clk(gclk));
	jdff dff_B_KPucb13f2_0(.din(w_dff_B_WDvzYpgM8_0),.dout(w_dff_B_KPucb13f2_0),.clk(gclk));
	jdff dff_B_DvaqvEzh1_0(.din(w_dff_B_KPucb13f2_0),.dout(w_dff_B_DvaqvEzh1_0),.clk(gclk));
	jdff dff_B_fXLA1Kwg5_0(.din(n402),.dout(w_dff_B_fXLA1Kwg5_0),.clk(gclk));
	jdff dff_B_uGceBSXD1_0(.din(n401),.dout(w_dff_B_uGceBSXD1_0),.clk(gclk));
	jdff dff_B_JR4jmXGn9_0(.din(n400),.dout(w_dff_B_JR4jmXGn9_0),.clk(gclk));
	jdff dff_B_yXmJwQZz2_0(.din(w_dff_B_JR4jmXGn9_0),.dout(w_dff_B_yXmJwQZz2_0),.clk(gclk));
	jdff dff_B_S9knLuoz8_0(.din(w_dff_B_yXmJwQZz2_0),.dout(w_dff_B_S9knLuoz8_0),.clk(gclk));
	jdff dff_B_gJI4gtky3_0(.din(w_dff_B_S9knLuoz8_0),.dout(w_dff_B_gJI4gtky3_0),.clk(gclk));
	jdff dff_A_VMdr5KKs9_1(.dout(w_G91gat_0[1]),.din(w_dff_A_VMdr5KKs9_1),.clk(gclk));
	jdff dff_A_cGuV4qg22_1(.dout(w_dff_A_VMdr5KKs9_1),.din(w_dff_A_cGuV4qg22_1),.clk(gclk));
	jdff dff_A_yw5pB7ZU7_1(.dout(w_dff_A_cGuV4qg22_1),.din(w_dff_A_yw5pB7ZU7_1),.clk(gclk));
	jdff dff_A_pL6PNmqM0_1(.dout(w_dff_A_yw5pB7ZU7_1),.din(w_dff_A_pL6PNmqM0_1),.clk(gclk));
	jdff dff_B_QJdRNliO0_0(.din(n397),.dout(w_dff_B_QJdRNliO0_0),.clk(gclk));
	jdff dff_B_TCeDcF568_0(.din(w_dff_B_QJdRNliO0_0),.dout(w_dff_B_TCeDcF568_0),.clk(gclk));
	jdff dff_B_OuzKgyVk5_0(.din(w_dff_B_TCeDcF568_0),.dout(w_dff_B_OuzKgyVk5_0),.clk(gclk));
	jdff dff_B_zUO9LkF29_0(.din(w_dff_B_OuzKgyVk5_0),.dout(w_dff_B_zUO9LkF29_0),.clk(gclk));
	jdff dff_B_aFNtfmEe2_0(.din(n393),.dout(w_dff_B_aFNtfmEe2_0),.clk(gclk));
	jdff dff_B_IFk6j4hx5_0(.din(w_dff_B_aFNtfmEe2_0),.dout(w_dff_B_IFk6j4hx5_0),.clk(gclk));
	jdff dff_B_t7OGI33X9_1(.din(n384),.dout(w_dff_B_t7OGI33X9_1),.clk(gclk));
	jdff dff_B_NFjd6RZw2_1(.din(w_dff_B_t7OGI33X9_1),.dout(w_dff_B_NFjd6RZw2_1),.clk(gclk));
	jdff dff_B_AWWx6la81_1(.din(w_dff_B_NFjd6RZw2_1),.dout(w_dff_B_AWWx6la81_1),.clk(gclk));
	jdff dff_B_UHBdicTG1_1(.din(w_dff_B_AWWx6la81_1),.dout(w_dff_B_UHBdicTG1_1),.clk(gclk));
	jdff dff_B_OmVkDI6T6_1(.din(w_dff_B_UHBdicTG1_1),.dout(w_dff_B_OmVkDI6T6_1),.clk(gclk));
	jdff dff_B_bCXKeL3Q5_1(.din(n385),.dout(w_dff_B_bCXKeL3Q5_1),.clk(gclk));
	jdff dff_B_8lLe8bRO6_1(.din(w_dff_B_bCXKeL3Q5_1),.dout(w_dff_B_8lLe8bRO6_1),.clk(gclk));
	jdff dff_B_FS4S2gvY5_1(.din(w_dff_B_8lLe8bRO6_1),.dout(w_dff_B_FS4S2gvY5_1),.clk(gclk));
	jdff dff_B_VXZhZo694_0(.din(n386),.dout(w_dff_B_VXZhZo694_0),.clk(gclk));
	jdff dff_B_1rxVpd3B8_0(.din(w_dff_B_VXZhZo694_0),.dout(w_dff_B_1rxVpd3B8_0),.clk(gclk));
	jdff dff_B_TNE1fgSQ0_0(.din(w_dff_B_1rxVpd3B8_0),.dout(w_dff_B_TNE1fgSQ0_0),.clk(gclk));
	jdff dff_B_Q7tIZrvg0_0(.din(w_dff_B_TNE1fgSQ0_0),.dout(w_dff_B_Q7tIZrvg0_0),.clk(gclk));
	jdff dff_A_F26RWqfw3_0(.dout(w_n330_0[0]),.din(w_dff_A_F26RWqfw3_0),.clk(gclk));
	jdff dff_A_w6cCnhXf2_0(.dout(w_dff_A_F26RWqfw3_0),.din(w_dff_A_w6cCnhXf2_0),.clk(gclk));
	jdff dff_A_tP72KhmC0_2(.dout(w_n330_0[2]),.din(w_dff_A_tP72KhmC0_2),.clk(gclk));
	jdff dff_A_LR4Lx2Rl6_2(.dout(w_dff_A_tP72KhmC0_2),.din(w_dff_A_LR4Lx2Rl6_2),.clk(gclk));
	jdff dff_A_DQ2OP5lH2_0(.dout(w_n337_0[0]),.din(w_dff_A_DQ2OP5lH2_0),.clk(gclk));
	jdff dff_A_jXjURwr55_0(.dout(w_dff_A_DQ2OP5lH2_0),.din(w_dff_A_jXjURwr55_0),.clk(gclk));
	jdff dff_A_1eFlQMwc5_2(.dout(w_n337_0[2]),.din(w_dff_A_1eFlQMwc5_2),.clk(gclk));
	jdff dff_B_hdsHP5x36_1(.din(n334),.dout(w_dff_B_hdsHP5x36_1),.clk(gclk));
	jdff dff_A_OrTZDfrS0_0(.dout(w_n322_0[0]),.din(w_dff_A_OrTZDfrS0_0),.clk(gclk));
	jdff dff_A_0NPLWfx13_0(.dout(w_G171gat_2[0]),.din(w_dff_A_0NPLWfx13_0),.clk(gclk));
	jdff dff_A_1uYTxSc76_0(.dout(w_dff_A_0NPLWfx13_0),.din(w_dff_A_1uYTxSc76_0),.clk(gclk));
	jdff dff_A_GroTSMkX2_0(.dout(w_dff_A_1uYTxSc76_0),.din(w_dff_A_GroTSMkX2_0),.clk(gclk));
	jdff dff_A_hqLRdRXR7_0(.dout(w_dff_A_GroTSMkX2_0),.din(w_dff_A_hqLRdRXR7_0),.clk(gclk));
	jdff dff_A_4QdAKl7x2_0(.dout(w_dff_A_hqLRdRXR7_0),.din(w_dff_A_4QdAKl7x2_0),.clk(gclk));
	jdff dff_A_Toq34Ftp1_1(.dout(w_n383_0[1]),.din(w_dff_A_Toq34Ftp1_1),.clk(gclk));
	jdff dff_A_u0MbFUW69_1(.dout(w_dff_A_Toq34Ftp1_1),.din(w_dff_A_u0MbFUW69_1),.clk(gclk));
	jdff dff_A_26T9gUqU7_1(.dout(w_dff_A_u0MbFUW69_1),.din(w_dff_A_26T9gUqU7_1),.clk(gclk));
	jdff dff_B_EBdouLYV6_0(.din(n310),.dout(w_dff_B_EBdouLYV6_0),.clk(gclk));
	jdff dff_B_hG7FzfcC7_0(.din(n309),.dout(w_dff_B_hG7FzfcC7_0),.clk(gclk));
	jdff dff_B_26EsKGKc5_0(.din(w_dff_B_hG7FzfcC7_0),.dout(w_dff_B_26EsKGKc5_0),.clk(gclk));
	jdff dff_B_8hh0wXRo8_0(.din(w_dff_B_26EsKGKc5_0),.dout(w_dff_B_8hh0wXRo8_0),.clk(gclk));
	jdff dff_A_kde8KbWV6_1(.dout(w_G165gat_1[1]),.din(w_dff_A_kde8KbWV6_1),.clk(gclk));
	jdff dff_A_IYTe57Ow2_1(.dout(w_dff_A_kde8KbWV6_1),.din(w_dff_A_IYTe57Ow2_1),.clk(gclk));
	jdff dff_A_NEqkcji58_1(.dout(w_dff_A_IYTe57Ow2_1),.din(w_dff_A_NEqkcji58_1),.clk(gclk));
	jdff dff_A_7fLYM1J14_1(.dout(w_dff_A_NEqkcji58_1),.din(w_dff_A_7fLYM1J14_1),.clk(gclk));
	jdff dff_A_nRO6zlfJ6_1(.dout(w_dff_A_7fLYM1J14_1),.din(w_dff_A_nRO6zlfJ6_1),.clk(gclk));
	jdff dff_A_kkTtHLAr6_2(.dout(w_G165gat_1[2]),.din(w_dff_A_kkTtHLAr6_2),.clk(gclk));
	jdff dff_A_dcmf4uhW4_2(.dout(w_dff_A_kkTtHLAr6_2),.din(w_dff_A_dcmf4uhW4_2),.clk(gclk));
	jdff dff_A_avPUcebe7_2(.dout(w_dff_A_dcmf4uhW4_2),.din(w_dff_A_avPUcebe7_2),.clk(gclk));
	jdff dff_A_Tuh0rk8I1_2(.dout(w_dff_A_avPUcebe7_2),.din(w_dff_A_Tuh0rk8I1_2),.clk(gclk));
	jdff dff_A_xpiXnAg21_2(.dout(w_dff_A_Tuh0rk8I1_2),.din(w_dff_A_xpiXnAg21_2),.clk(gclk));
	jdff dff_A_hrMTLzGq3_2(.dout(w_G165gat_0[2]),.din(w_dff_A_hrMTLzGq3_2),.clk(gclk));
	jdff dff_A_ZqPDn6VT1_2(.dout(w_dff_A_hrMTLzGq3_2),.din(w_dff_A_ZqPDn6VT1_2),.clk(gclk));
	jdff dff_A_fS6lAHk55_2(.dout(w_dff_A_ZqPDn6VT1_2),.din(w_dff_A_fS6lAHk55_2),.clk(gclk));
	jdff dff_A_UlOMJKSX8_2(.dout(w_dff_A_fS6lAHk55_2),.din(w_dff_A_UlOMJKSX8_2),.clk(gclk));
	jdff dff_B_IUIDNKMu1_0(.din(n425),.dout(w_dff_B_IUIDNKMu1_0),.clk(gclk));
	jdff dff_B_UGlBo0xK1_0(.din(w_dff_B_IUIDNKMu1_0),.dout(w_dff_B_UGlBo0xK1_0),.clk(gclk));
	jdff dff_B_TNUumohk1_0(.din(w_dff_B_UGlBo0xK1_0),.dout(w_dff_B_TNUumohk1_0),.clk(gclk));
	jdff dff_B_EMxNHy8h2_0(.din(w_dff_B_TNUumohk1_0),.dout(w_dff_B_EMxNHy8h2_0),.clk(gclk));
	jdff dff_B_hm1XeEtH1_0(.din(w_dff_B_EMxNHy8h2_0),.dout(w_dff_B_hm1XeEtH1_0),.clk(gclk));
	jdff dff_B_SLMKw8mj6_0(.din(w_dff_B_hm1XeEtH1_0),.dout(w_dff_B_SLMKw8mj6_0),.clk(gclk));
	jdff dff_B_cu1HmymM7_0(.din(n424),.dout(w_dff_B_cu1HmymM7_0),.clk(gclk));
	jdff dff_B_gxFDA8u96_0(.din(n423),.dout(w_dff_B_gxFDA8u96_0),.clk(gclk));
	jdff dff_B_OHzfU9DY0_0(.din(n422),.dout(w_dff_B_OHzfU9DY0_0),.clk(gclk));
	jdff dff_B_bqNuC5lG2_0(.din(w_dff_B_OHzfU9DY0_0),.dout(w_dff_B_bqNuC5lG2_0),.clk(gclk));
	jdff dff_B_qDcTqQTy0_0(.din(w_dff_B_bqNuC5lG2_0),.dout(w_dff_B_qDcTqQTy0_0),.clk(gclk));
	jdff dff_B_E01akAsv8_0(.din(w_dff_B_qDcTqQTy0_0),.dout(w_dff_B_E01akAsv8_0),.clk(gclk));
	jdff dff_A_xFuZkLqu4_1(.dout(w_G96gat_0[1]),.din(w_dff_A_xFuZkLqu4_1),.clk(gclk));
	jdff dff_A_eeNuPG999_1(.dout(w_dff_A_xFuZkLqu4_1),.din(w_dff_A_eeNuPG999_1),.clk(gclk));
	jdff dff_A_exMt7xXh8_1(.dout(w_dff_A_eeNuPG999_1),.din(w_dff_A_exMt7xXh8_1),.clk(gclk));
	jdff dff_A_OoE4TLiA8_1(.dout(w_dff_A_exMt7xXh8_1),.din(w_dff_A_OoE4TLiA8_1),.clk(gclk));
	jdff dff_B_bTk1evDX6_1(.din(G73gat),.dout(w_dff_B_bTk1evDX6_1),.clk(gclk));
	jdff dff_A_rroH0NRy0_0(.dout(w_n121_0[0]),.din(w_dff_A_rroH0NRy0_0),.clk(gclk));
	jdff dff_A_iJ7ti8ja8_0(.dout(w_n118_0[0]),.din(w_dff_A_iJ7ti8ja8_0),.clk(gclk));
	jdff dff_B_rQ53D53U7_0(.din(n419),.dout(w_dff_B_rQ53D53U7_0),.clk(gclk));
	jdff dff_B_bstnPsQi3_0(.din(w_dff_B_rQ53D53U7_0),.dout(w_dff_B_bstnPsQi3_0),.clk(gclk));
	jdff dff_B_URpqphkC3_0(.din(w_dff_B_bstnPsQi3_0),.dout(w_dff_B_URpqphkC3_0),.clk(gclk));
	jdff dff_B_LH0q07pu1_0(.din(w_dff_B_URpqphkC3_0),.dout(w_dff_B_LH0q07pu1_0),.clk(gclk));
	jdff dff_B_EDrNy9Qv7_3(.din(G246gat),.dout(w_dff_B_EDrNy9Qv7_3),.clk(gclk));
	jdff dff_B_I197bpcy1_3(.din(G228gat),.dout(w_dff_B_I197bpcy1_3),.clk(gclk));
	jdff dff_B_cB3UcaAg3_3(.din(w_dff_B_I197bpcy1_3),.dout(w_dff_B_cB3UcaAg3_3),.clk(gclk));
	jdff dff_B_gHPIPODr6_3(.din(w_dff_B_cB3UcaAg3_3),.dout(w_dff_B_gHPIPODr6_3),.clk(gclk));
	jdff dff_B_FXZdrSVc9_3(.din(w_dff_B_gHPIPODr6_3),.dout(w_dff_B_FXZdrSVc9_3),.clk(gclk));
	jdff dff_B_Y2SJCPfc4_3(.din(w_dff_B_FXZdrSVc9_3),.dout(w_dff_B_Y2SJCPfc4_3),.clk(gclk));
	jdff dff_B_2e29grpO7_3(.din(w_dff_B_Y2SJCPfc4_3),.dout(w_dff_B_2e29grpO7_3),.clk(gclk));
	jdff dff_B_QRYtAD1m5_0(.din(n415),.dout(w_dff_B_QRYtAD1m5_0),.clk(gclk));
	jdff dff_B_IynLEhcC6_0(.din(w_dff_B_QRYtAD1m5_0),.dout(w_dff_B_IynLEhcC6_0),.clk(gclk));
	jdff dff_A_oaewuqkV7_2(.dout(w_G219gat_1[2]),.din(w_dff_A_oaewuqkV7_2),.clk(gclk));
	jdff dff_A_3fbe5yX90_0(.dout(w_G219gat_0[0]),.din(w_dff_A_3fbe5yX90_0),.clk(gclk));
	jdff dff_A_Yhi45xwW4_0(.dout(w_dff_A_3fbe5yX90_0),.din(w_dff_A_Yhi45xwW4_0),.clk(gclk));
	jdff dff_A_4ENWc2UQ5_0(.dout(w_dff_A_Yhi45xwW4_0),.din(w_dff_A_4ENWc2UQ5_0),.clk(gclk));
	jdff dff_B_3dvAC20P0_3(.din(G219gat),.dout(w_dff_B_3dvAC20P0_3),.clk(gclk));
	jdff dff_B_JJ8quy0X9_3(.din(w_dff_B_3dvAC20P0_3),.dout(w_dff_B_JJ8quy0X9_3),.clk(gclk));
	jdff dff_B_7IxA7YG45_3(.din(w_dff_B_JJ8quy0X9_3),.dout(w_dff_B_7IxA7YG45_3),.clk(gclk));
	jdff dff_B_8AfPiWn38_3(.din(w_dff_B_7IxA7YG45_3),.dout(w_dff_B_8AfPiWn38_3),.clk(gclk));
	jdff dff_B_LynXWjTt5_3(.din(w_dff_B_8AfPiWn38_3),.dout(w_dff_B_LynXWjTt5_3),.clk(gclk));
	jdff dff_B_pxyp9p9L1_3(.din(w_dff_B_LynXWjTt5_3),.dout(w_dff_B_pxyp9p9L1_3),.clk(gclk));
	jdff dff_B_Trd5Tr939_1(.din(n406),.dout(w_dff_B_Trd5Tr939_1),.clk(gclk));
	jdff dff_B_MwRscJ6z0_1(.din(w_dff_B_Trd5Tr939_1),.dout(w_dff_B_MwRscJ6z0_1),.clk(gclk));
	jdff dff_B_UgSJfTAn9_1(.din(w_dff_B_MwRscJ6z0_1),.dout(w_dff_B_UgSJfTAn9_1),.clk(gclk));
	jdff dff_B_CqbQpbKg4_1(.din(w_dff_B_UgSJfTAn9_1),.dout(w_dff_B_CqbQpbKg4_1),.clk(gclk));
	jdff dff_B_rXqprOXe5_1(.din(w_dff_B_CqbQpbKg4_1),.dout(w_dff_B_rXqprOXe5_1),.clk(gclk));
	jdff dff_B_Lk9n5vFc8_1(.din(n407),.dout(w_dff_B_Lk9n5vFc8_1),.clk(gclk));
	jdff dff_B_IWlkaJ328_1(.din(w_dff_B_Lk9n5vFc8_1),.dout(w_dff_B_IWlkaJ328_1),.clk(gclk));
	jdff dff_B_vgmAWVGe2_1(.din(w_dff_B_IWlkaJ328_1),.dout(w_dff_B_vgmAWVGe2_1),.clk(gclk));
	jdff dff_B_1vPFDyg56_1(.din(w_dff_B_vgmAWVGe2_1),.dout(w_dff_B_1vPFDyg56_1),.clk(gclk));
	jdff dff_B_EuNeFiDO4_0(.din(n408),.dout(w_dff_B_EuNeFiDO4_0),.clk(gclk));
	jdff dff_B_yWqxq0RV0_0(.din(w_dff_B_EuNeFiDO4_0),.dout(w_dff_B_yWqxq0RV0_0),.clk(gclk));
	jdff dff_B_Wkn7JBwa7_0(.din(w_dff_B_yWqxq0RV0_0),.dout(w_dff_B_Wkn7JBwa7_0),.clk(gclk));
	jdff dff_B_mDSeZK8l5_0(.din(w_dff_B_Wkn7JBwa7_0),.dout(w_dff_B_mDSeZK8l5_0),.clk(gclk));
	jdff dff_B_83uWI9Ei6_0(.din(w_dff_B_mDSeZK8l5_0),.dout(w_dff_B_83uWI9Ei6_0),.clk(gclk));
	jdff dff_A_meshnIlr3_0(.dout(w_n329_0[0]),.din(w_dff_A_meshnIlr3_0),.clk(gclk));
	jdff dff_A_o8ZADDjP9_0(.dout(w_dff_A_meshnIlr3_0),.din(w_dff_A_o8ZADDjP9_0),.clk(gclk));
	jdff dff_A_EfEh2nT13_0(.dout(w_dff_A_o8ZADDjP9_0),.din(w_dff_A_EfEh2nT13_0),.clk(gclk));
	jdff dff_A_AqKNoOu96_0(.dout(w_G177gat_2[0]),.din(w_dff_A_AqKNoOu96_0),.clk(gclk));
	jdff dff_A_AR0qnh854_0(.dout(w_dff_A_AqKNoOu96_0),.din(w_dff_A_AR0qnh854_0),.clk(gclk));
	jdff dff_A_jhnaDi6Q5_0(.dout(w_dff_A_AR0qnh854_0),.din(w_dff_A_jhnaDi6Q5_0),.clk(gclk));
	jdff dff_A_0ruHWeOA0_0(.dout(w_dff_A_jhnaDi6Q5_0),.din(w_dff_A_0ruHWeOA0_0),.clk(gclk));
	jdff dff_A_tSi1udYA9_0(.dout(w_dff_A_0ruHWeOA0_0),.din(w_dff_A_tSi1udYA9_0),.clk(gclk));
	jdff dff_B_Y21dHlA20_1(.din(n343),.dout(w_dff_B_Y21dHlA20_1),.clk(gclk));
	jdff dff_B_lFQHA1xg4_1(.din(w_dff_B_Y21dHlA20_1),.dout(w_dff_B_lFQHA1xg4_1),.clk(gclk));
	jdff dff_B_F7k906ye5_1(.din(w_dff_B_lFQHA1xg4_1),.dout(w_dff_B_F7k906ye5_1),.clk(gclk));
	jdff dff_B_6Wsnj20d7_1(.din(n344),.dout(w_dff_B_6Wsnj20d7_1),.clk(gclk));
	jdff dff_B_mnDYvqjb1_1(.din(w_dff_B_6Wsnj20d7_1),.dout(w_dff_B_mnDYvqjb1_1),.clk(gclk));
	jdff dff_B_nL8RapGL9_1(.din(w_dff_B_mnDYvqjb1_1),.dout(w_dff_B_nL8RapGL9_1),.clk(gclk));
	jdff dff_B_narWwQcN6_1(.din(w_dff_B_nL8RapGL9_1),.dout(w_dff_B_narWwQcN6_1),.clk(gclk));
	jdff dff_B_aHVTPXgO2_0(.din(n231),.dout(w_dff_B_aHVTPXgO2_0),.clk(gclk));
	jdff dff_B_Trua98Zs7_1(.din(n227),.dout(w_dff_B_Trua98Zs7_1),.clk(gclk));
	jdff dff_A_V8hvUBDX6_0(.dout(w_n228_0[0]),.din(w_dff_A_V8hvUBDX6_0),.clk(gclk));
	jdff dff_A_Cv2sEDgY6_1(.dout(w_G195gat_1[1]),.din(w_dff_A_Cv2sEDgY6_1),.clk(gclk));
	jdff dff_A_apuwql6P9_1(.dout(w_dff_A_Cv2sEDgY6_1),.din(w_dff_A_apuwql6P9_1),.clk(gclk));
	jdff dff_A_hgx5JAxi9_1(.dout(w_dff_A_apuwql6P9_1),.din(w_dff_A_hgx5JAxi9_1),.clk(gclk));
	jdff dff_A_rcEbG1DU5_1(.dout(w_dff_A_hgx5JAxi9_1),.din(w_dff_A_rcEbG1DU5_1),.clk(gclk));
	jdff dff_A_PEiE3VZj4_1(.dout(w_dff_A_rcEbG1DU5_1),.din(w_dff_A_PEiE3VZj4_1),.clk(gclk));
	jdff dff_A_ZwhRxtqS7_2(.dout(w_G195gat_1[2]),.din(w_dff_A_ZwhRxtqS7_2),.clk(gclk));
	jdff dff_A_I2fEbQkG9_2(.dout(w_dff_A_ZwhRxtqS7_2),.din(w_dff_A_I2fEbQkG9_2),.clk(gclk));
	jdff dff_A_7IM0uEVl7_2(.dout(w_dff_A_I2fEbQkG9_2),.din(w_dff_A_7IM0uEVl7_2),.clk(gclk));
	jdff dff_A_OXLvQ9607_2(.dout(w_dff_A_7IM0uEVl7_2),.din(w_dff_A_OXLvQ9607_2),.clk(gclk));
	jdff dff_A_MAcl6UMd6_2(.dout(w_dff_A_OXLvQ9607_2),.din(w_dff_A_MAcl6UMd6_2),.clk(gclk));
	jdff dff_A_fUtHtfC04_1(.dout(w_G189gat_1[1]),.din(w_dff_A_fUtHtfC04_1),.clk(gclk));
	jdff dff_A_EMXOtX4A2_1(.dout(w_dff_A_fUtHtfC04_1),.din(w_dff_A_EMXOtX4A2_1),.clk(gclk));
	jdff dff_A_IWsJA5zo2_1(.dout(w_dff_A_EMXOtX4A2_1),.din(w_dff_A_IWsJA5zo2_1),.clk(gclk));
	jdff dff_A_9eTEvFFl6_1(.dout(w_dff_A_IWsJA5zo2_1),.din(w_dff_A_9eTEvFFl6_1),.clk(gclk));
	jdff dff_A_shIFNGEE6_1(.dout(w_dff_A_9eTEvFFl6_1),.din(w_dff_A_shIFNGEE6_1),.clk(gclk));
	jdff dff_A_aSZ1xRXd1_2(.dout(w_G189gat_1[2]),.din(w_dff_A_aSZ1xRXd1_2),.clk(gclk));
	jdff dff_A_Z8WyBcoU9_2(.dout(w_dff_A_aSZ1xRXd1_2),.din(w_dff_A_Z8WyBcoU9_2),.clk(gclk));
	jdff dff_A_sGhJTLmD8_2(.dout(w_dff_A_Z8WyBcoU9_2),.din(w_dff_A_sGhJTLmD8_2),.clk(gclk));
	jdff dff_A_0GZ52bW43_2(.dout(w_dff_A_sGhJTLmD8_2),.din(w_dff_A_0GZ52bW43_2),.clk(gclk));
	jdff dff_A_xVuBfEC40_2(.dout(w_dff_A_0GZ52bW43_2),.din(w_dff_A_xVuBfEC40_2),.clk(gclk));
	jdff dff_B_61OrHqTo4_0(.din(n225),.dout(w_dff_B_61OrHqTo4_0),.clk(gclk));
	jdff dff_B_AL7EJi0i1_0(.din(w_dff_B_61OrHqTo4_0),.dout(w_dff_B_AL7EJi0i1_0),.clk(gclk));
	jdff dff_A_PNKwbeGg8_0(.dout(w_n223_0[0]),.din(w_dff_A_PNKwbeGg8_0),.clk(gclk));
	jdff dff_A_fwagVIfq9_0(.dout(w_G121gat_0[0]),.din(w_dff_A_fwagVIfq9_0),.clk(gclk));
	jdff dff_A_9YJutSWW9_0(.dout(w_dff_A_fwagVIfq9_0),.din(w_dff_A_9YJutSWW9_0),.clk(gclk));
	jdff dff_A_RinIkOCv8_0(.dout(w_dff_A_9YJutSWW9_0),.din(w_dff_A_RinIkOCv8_0),.clk(gclk));
	jdff dff_A_lavV9sd30_0(.dout(w_dff_A_RinIkOCv8_0),.din(w_dff_A_lavV9sd30_0),.clk(gclk));
	jdff dff_A_ozYhWeqW5_0(.dout(w_G195gat_2[0]),.din(w_dff_A_ozYhWeqW5_0),.clk(gclk));
	jdff dff_A_smbCcj5w4_0(.dout(w_dff_A_ozYhWeqW5_0),.din(w_dff_A_smbCcj5w4_0),.clk(gclk));
	jdff dff_A_xQO5tiDz8_0(.dout(w_dff_A_smbCcj5w4_0),.din(w_dff_A_xQO5tiDz8_0),.clk(gclk));
	jdff dff_A_EiDKGSNC4_0(.dout(w_dff_A_xQO5tiDz8_0),.din(w_dff_A_EiDKGSNC4_0),.clk(gclk));
	jdff dff_A_cckamYwI8_0(.dout(w_dff_A_EiDKGSNC4_0),.din(w_dff_A_cckamYwI8_0),.clk(gclk));
	jdff dff_A_ROfnJ5Yt5_2(.dout(w_G195gat_0[2]),.din(w_dff_A_ROfnJ5Yt5_2),.clk(gclk));
	jdff dff_A_YeruOvK76_2(.dout(w_dff_A_ROfnJ5Yt5_2),.din(w_dff_A_YeruOvK76_2),.clk(gclk));
	jdff dff_A_BQ90wCFA9_2(.dout(w_dff_A_YeruOvK76_2),.din(w_dff_A_BQ90wCFA9_2),.clk(gclk));
	jdff dff_A_SjwLYvEt5_2(.dout(w_dff_A_BQ90wCFA9_2),.din(w_dff_A_SjwLYvEt5_2),.clk(gclk));
	jdff dff_A_XbNcbaxR3_0(.dout(w_n218_0[0]),.din(w_dff_A_XbNcbaxR3_0),.clk(gclk));
	jdff dff_A_tvGuVQJn9_1(.dout(w_G116gat_0[1]),.din(w_dff_A_tvGuVQJn9_1),.clk(gclk));
	jdff dff_A_Jgz18uXf7_1(.dout(w_dff_A_tvGuVQJn9_1),.din(w_dff_A_Jgz18uXf7_1),.clk(gclk));
	jdff dff_A_F5XMcJzC9_1(.dout(w_dff_A_Jgz18uXf7_1),.din(w_dff_A_F5XMcJzC9_1),.clk(gclk));
	jdff dff_A_CimypAnj1_1(.dout(w_dff_A_F5XMcJzC9_1),.din(w_dff_A_CimypAnj1_1),.clk(gclk));
	jdff dff_B_vyXG6hTQ3_2(.din(G146gat),.dout(w_dff_B_vyXG6hTQ3_2),.clk(gclk));
	jdff dff_B_E2MeZ04I1_2(.din(w_dff_B_vyXG6hTQ3_2),.dout(w_dff_B_E2MeZ04I1_2),.clk(gclk));
	jdff dff_B_9EYRklc78_2(.din(w_dff_B_E2MeZ04I1_2),.dout(w_dff_B_9EYRklc78_2),.clk(gclk));
	jdff dff_B_zbrf4LS31_2(.din(w_dff_B_9EYRklc78_2),.dout(w_dff_B_zbrf4LS31_2),.clk(gclk));
	jdff dff_A_xYCSH7WV4_0(.dout(w_G189gat_2[0]),.din(w_dff_A_xYCSH7WV4_0),.clk(gclk));
	jdff dff_A_BfioD60e7_0(.dout(w_dff_A_xYCSH7WV4_0),.din(w_dff_A_BfioD60e7_0),.clk(gclk));
	jdff dff_A_GzkKLqZq9_0(.dout(w_dff_A_BfioD60e7_0),.din(w_dff_A_GzkKLqZq9_0),.clk(gclk));
	jdff dff_A_lV2ZbfwP1_0(.dout(w_dff_A_GzkKLqZq9_0),.din(w_dff_A_lV2ZbfwP1_0),.clk(gclk));
	jdff dff_A_RvVo3Sl95_0(.dout(w_dff_A_lV2ZbfwP1_0),.din(w_dff_A_RvVo3Sl95_0),.clk(gclk));
	jdff dff_A_Mwx6w1xR2_2(.dout(w_G189gat_0[2]),.din(w_dff_A_Mwx6w1xR2_2),.clk(gclk));
	jdff dff_A_ZYLUP0gu4_2(.dout(w_dff_A_Mwx6w1xR2_2),.din(w_dff_A_ZYLUP0gu4_2),.clk(gclk));
	jdff dff_A_hGaAqTP40_2(.dout(w_dff_A_ZYLUP0gu4_2),.din(w_dff_A_hGaAqTP40_2),.clk(gclk));
	jdff dff_A_fNGl3RZk3_2(.dout(w_dff_A_hGaAqTP40_2),.din(w_dff_A_fNGl3RZk3_2),.clk(gclk));
	jdff dff_B_UPcoI7sI3_1(.din(n197),.dout(w_dff_B_UPcoI7sI3_1),.clk(gclk));
	jdff dff_B_kwGqkp5m8_1(.din(n198),.dout(w_dff_B_kwGqkp5m8_1),.clk(gclk));
	jdff dff_B_0XRj0AEU8_1(.din(w_dff_B_kwGqkp5m8_1),.dout(w_dff_B_0XRj0AEU8_1),.clk(gclk));
	jdff dff_B_nB9njjf62_1(.din(w_dff_B_0XRj0AEU8_1),.dout(w_dff_B_nB9njjf62_1),.clk(gclk));
	jdff dff_B_LRtxNgy08_1(.din(w_dff_B_nB9njjf62_1),.dout(w_dff_B_LRtxNgy08_1),.clk(gclk));
	jdff dff_B_YR9TAPNw9_1(.din(w_dff_B_LRtxNgy08_1),.dout(w_dff_B_YR9TAPNw9_1),.clk(gclk));
	jdff dff_B_uZ4htwsd5_1(.din(w_dff_B_YR9TAPNw9_1),.dout(w_dff_B_uZ4htwsd5_1),.clk(gclk));
	jdff dff_B_fsrMkPh27_1(.din(n207),.dout(w_dff_B_fsrMkPh27_1),.clk(gclk));
	jdff dff_B_0eKCEbDJ8_1(.din(w_dff_B_fsrMkPh27_1),.dout(w_dff_B_0eKCEbDJ8_1),.clk(gclk));
	jdff dff_B_Wv37bgjK0_1(.din(w_dff_B_0eKCEbDJ8_1),.dout(w_dff_B_Wv37bgjK0_1),.clk(gclk));
	jdff dff_B_O6XjXY0V3_1(.din(n200),.dout(w_dff_B_O6XjXY0V3_1),.clk(gclk));
	jdff dff_A_2UdM7RhN4_1(.dout(w_n98_0[1]),.din(w_dff_A_2UdM7RhN4_1),.clk(gclk));
	jdff dff_A_OICYdldO3_0(.dout(w_n143_0[0]),.din(w_dff_A_OICYdldO3_0),.clk(gclk));
	jdff dff_B_00vgoY1g7_2(.din(n143),.dout(w_dff_B_00vgoY1g7_2),.clk(gclk));
	jdff dff_B_U1KzZo9Y5_2(.din(w_dff_B_00vgoY1g7_2),.dout(w_dff_B_U1KzZo9Y5_2),.clk(gclk));
	jdff dff_B_LYo6SleD5_2(.din(w_dff_B_U1KzZo9Y5_2),.dout(w_dff_B_LYo6SleD5_2),.clk(gclk));
	jdff dff_B_hqW6uudj2_2(.din(w_dff_B_LYo6SleD5_2),.dout(w_dff_B_hqW6uudj2_2),.clk(gclk));
	jdff dff_B_S3J6TAuL5_2(.din(w_dff_B_hqW6uudj2_2),.dout(w_dff_B_S3J6TAuL5_2),.clk(gclk));
	jdff dff_B_rqeHkNQs4_2(.din(w_dff_B_S3J6TAuL5_2),.dout(w_dff_B_rqeHkNQs4_2),.clk(gclk));
	jdff dff_A_uWkGS9cc4_0(.dout(w_G261gat_0[0]),.din(w_dff_A_uWkGS9cc4_0),.clk(gclk));
	jdff dff_A_VN7NTbAY7_0(.dout(w_dff_A_uWkGS9cc4_0),.din(w_dff_A_VN7NTbAY7_0),.clk(gclk));
	jdff dff_A_wOJn1mwW2_0(.dout(w_dff_A_VN7NTbAY7_0),.din(w_dff_A_wOJn1mwW2_0),.clk(gclk));
	jdff dff_A_sYJNZTGl0_0(.dout(w_dff_A_wOJn1mwW2_0),.din(w_dff_A_sYJNZTGl0_0),.clk(gclk));
	jdff dff_A_EvZfo1l24_0(.dout(w_dff_A_sYJNZTGl0_0),.din(w_dff_A_EvZfo1l24_0),.clk(gclk));
	jdff dff_A_hyshpDJ33_1(.dout(w_G261gat_0[1]),.din(w_dff_A_hyshpDJ33_1),.clk(gclk));
	jdff dff_A_FzZXfQwl5_1(.dout(w_dff_A_hyshpDJ33_1),.din(w_dff_A_FzZXfQwl5_1),.clk(gclk));
	jdff dff_A_ZCtu9FJf5_1(.dout(w_dff_A_FzZXfQwl5_1),.din(w_dff_A_ZCtu9FJf5_1),.clk(gclk));
	jdff dff_A_rELLcDRh6_1(.dout(w_dff_A_ZCtu9FJf5_1),.din(w_dff_A_rELLcDRh6_1),.clk(gclk));
	jdff dff_A_W0PampPv6_1(.dout(w_dff_A_rELLcDRh6_1),.din(w_dff_A_W0PampPv6_1),.clk(gclk));
	jdff dff_A_nlLGuuQ96_1(.dout(w_dff_A_W0PampPv6_1),.din(w_dff_A_nlLGuuQ96_1),.clk(gclk));
	jdff dff_A_IelfkTM72_0(.dout(w_G126gat_0[0]),.din(w_dff_A_IelfkTM72_0),.clk(gclk));
	jdff dff_A_efxspf6Y1_0(.dout(w_dff_A_IelfkTM72_0),.din(w_dff_A_efxspf6Y1_0),.clk(gclk));
	jdff dff_A_c65xE3uH0_0(.dout(w_dff_A_efxspf6Y1_0),.din(w_dff_A_c65xE3uH0_0),.clk(gclk));
	jdff dff_A_lf6NpmqY2_0(.dout(w_dff_A_c65xE3uH0_0),.din(w_dff_A_lf6NpmqY2_0),.clk(gclk));
	jdff dff_A_uUVRCGzd9_1(.dout(w_G201gat_1[1]),.din(w_dff_A_uUVRCGzd9_1),.clk(gclk));
	jdff dff_A_iyjeknyI0_1(.dout(w_dff_A_uUVRCGzd9_1),.din(w_dff_A_iyjeknyI0_1),.clk(gclk));
	jdff dff_A_I4iK7PvG7_1(.dout(w_dff_A_iyjeknyI0_1),.din(w_dff_A_I4iK7PvG7_1),.clk(gclk));
	jdff dff_A_vTf2BcLL8_1(.dout(w_dff_A_I4iK7PvG7_1),.din(w_dff_A_vTf2BcLL8_1),.clk(gclk));
	jdff dff_A_umEvOaAC1_1(.dout(w_dff_A_vTf2BcLL8_1),.din(w_dff_A_umEvOaAC1_1),.clk(gclk));
	jdff dff_A_0HQrlmgz6_2(.dout(w_G201gat_1[2]),.din(w_dff_A_0HQrlmgz6_2),.clk(gclk));
	jdff dff_A_dtkCYSJt1_2(.dout(w_dff_A_0HQrlmgz6_2),.din(w_dff_A_dtkCYSJt1_2),.clk(gclk));
	jdff dff_A_dwTOpPhS0_2(.dout(w_dff_A_dtkCYSJt1_2),.din(w_dff_A_dwTOpPhS0_2),.clk(gclk));
	jdff dff_A_1Ilctpke0_2(.dout(w_dff_A_dwTOpPhS0_2),.din(w_dff_A_1Ilctpke0_2),.clk(gclk));
	jdff dff_A_ak03yzzv9_2(.dout(w_G201gat_0[2]),.din(w_dff_A_ak03yzzv9_2),.clk(gclk));
	jdff dff_A_HBMqRywl4_2(.dout(w_dff_A_ak03yzzv9_2),.din(w_dff_A_HBMqRywl4_2),.clk(gclk));
	jdff dff_A_NH9NBmG28_2(.dout(w_dff_A_HBMqRywl4_2),.din(w_dff_A_NH9NBmG28_2),.clk(gclk));
	jdff dff_A_1lz8NpTd1_2(.dout(w_dff_A_NH9NBmG28_2),.din(w_dff_A_1lz8NpTd1_2),.clk(gclk));
	jdff dff_A_PdBieuzD8_2(.dout(w_dff_A_1lz8NpTd1_2),.din(w_dff_A_PdBieuzD8_2),.clk(gclk));
	jdff dff_A_yW1cWfIT3_1(.dout(w_n303_0[1]),.din(w_dff_A_yW1cWfIT3_1),.clk(gclk));
	jdff dff_A_zL7JR5nd9_1(.dout(w_dff_A_yW1cWfIT3_1),.din(w_dff_A_zL7JR5nd9_1),.clk(gclk));
	jdff dff_A_CWcQXXlt9_1(.dout(w_n302_0[1]),.din(w_dff_A_CWcQXXlt9_1),.clk(gclk));
	jdff dff_A_fq5Nvc0t6_1(.dout(w_dff_A_CWcQXXlt9_1),.din(w_dff_A_fq5Nvc0t6_1),.clk(gclk));
	jdff dff_A_1bNLhzwk4_1(.dout(w_G111gat_0[1]),.din(w_dff_A_1bNLhzwk4_1),.clk(gclk));
	jdff dff_A_KVWEHmL78_1(.dout(w_dff_A_1bNLhzwk4_1),.din(w_dff_A_KVWEHmL78_1),.clk(gclk));
	jdff dff_A_i8kZMIhV1_1(.dout(w_dff_A_KVWEHmL78_1),.din(w_dff_A_i8kZMIhV1_1),.clk(gclk));
	jdff dff_A_NzuKRQ147_1(.dout(w_dff_A_i8kZMIhV1_1),.din(w_dff_A_NzuKRQ147_1),.clk(gclk));
	jdff dff_A_u0OO4cb02_1(.dout(w_n165_1[1]),.din(w_dff_A_u0OO4cb02_1),.clk(gclk));
	jdff dff_A_BY2TtJ9M2_2(.dout(w_n165_1[2]),.din(w_dff_A_BY2TtJ9M2_2),.clk(gclk));
	jdff dff_A_LjJcmoBW0_1(.dout(w_n165_0[1]),.din(w_dff_A_LjJcmoBW0_1),.clk(gclk));
	jdff dff_A_fgfiDB7k9_2(.dout(w_n165_0[2]),.din(w_dff_A_fgfiDB7k9_2),.clk(gclk));
	jdff dff_B_y2uImBIK9_0(.din(n164),.dout(w_dff_B_y2uImBIK9_0),.clk(gclk));
	jdff dff_A_5w84HB3h2_0(.dout(w_n96_0[0]),.din(w_dff_A_5w84HB3h2_0),.clk(gclk));
	jdff dff_A_diRpe3DD4_0(.dout(w_dff_A_5w84HB3h2_0),.din(w_dff_A_diRpe3DD4_0),.clk(gclk));
	jdff dff_A_h23fIEli9_0(.dout(w_dff_A_diRpe3DD4_0),.din(w_dff_A_h23fIEli9_0),.clk(gclk));
	jdff dff_B_0qKh4jwL3_2(.din(G143gat),.dout(w_dff_B_0qKh4jwL3_2),.clk(gclk));
	jdff dff_B_hkQR92ex7_2(.din(w_dff_B_0qKh4jwL3_2),.dout(w_dff_B_hkQR92ex7_2),.clk(gclk));
	jdff dff_B_HRJctjGL9_2(.din(w_dff_B_hkQR92ex7_2),.dout(w_dff_B_HRJctjGL9_2),.clk(gclk));
	jdff dff_B_jZrZfJia1_2(.din(w_dff_B_HRJctjGL9_2),.dout(w_dff_B_jZrZfJia1_2),.clk(gclk));
	jdff dff_A_J27AVUAR9_0(.dout(w_G183gat_1[0]),.din(w_dff_A_J27AVUAR9_0),.clk(gclk));
	jdff dff_A_OvJAZY9D2_0(.dout(w_dff_A_J27AVUAR9_0),.din(w_dff_A_OvJAZY9D2_0),.clk(gclk));
	jdff dff_A_ShPg6NR06_0(.dout(w_dff_A_OvJAZY9D2_0),.din(w_dff_A_ShPg6NR06_0),.clk(gclk));
	jdff dff_A_TuwgX4D81_0(.dout(w_dff_A_ShPg6NR06_0),.din(w_dff_A_TuwgX4D81_0),.clk(gclk));
	jdff dff_A_29NPMiPM0_0(.dout(w_dff_A_TuwgX4D81_0),.din(w_dff_A_29NPMiPM0_0),.clk(gclk));
	jdff dff_A_UJ5DfTng2_1(.dout(w_G183gat_1[1]),.din(w_dff_A_UJ5DfTng2_1),.clk(gclk));
	jdff dff_A_Cq9cKhTU2_1(.dout(w_dff_A_UJ5DfTng2_1),.din(w_dff_A_Cq9cKhTU2_1),.clk(gclk));
	jdff dff_A_zKbzkcZs4_1(.dout(w_dff_A_Cq9cKhTU2_1),.din(w_dff_A_zKbzkcZs4_1),.clk(gclk));
	jdff dff_A_B6XSKzLl1_1(.dout(w_dff_A_zKbzkcZs4_1),.din(w_dff_A_B6XSKzLl1_1),.clk(gclk));
	jdff dff_A_t31raUJ22_2(.dout(w_G183gat_0[2]),.din(w_dff_A_t31raUJ22_2),.clk(gclk));
	jdff dff_A_UFZ17GAg2_2(.dout(w_dff_A_t31raUJ22_2),.din(w_dff_A_UFZ17GAg2_2),.clk(gclk));
	jdff dff_A_JbebVzyX0_2(.dout(w_dff_A_UFZ17GAg2_2),.din(w_dff_A_JbebVzyX0_2),.clk(gclk));
	jdff dff_A_gb44LIHt8_2(.dout(w_dff_A_JbebVzyX0_2),.din(w_dff_A_gb44LIHt8_2),.clk(gclk));
	jdff dff_A_AWuuuy1O1_2(.dout(w_dff_A_gb44LIHt8_2),.din(w_dff_A_AWuuuy1O1_2),.clk(gclk));
	jdff dff_A_mv9Ijic62_0(.dout(w_n335_0[0]),.din(w_dff_A_mv9Ijic62_0),.clk(gclk));
	jdff dff_A_7mrNzY6F7_0(.dout(w_dff_A_mv9Ijic62_0),.din(w_dff_A_7mrNzY6F7_0),.clk(gclk));
	jdff dff_A_HLFM1v4Q5_0(.dout(w_dff_A_7mrNzY6F7_0),.din(w_dff_A_HLFM1v4Q5_0),.clk(gclk));
	jdff dff_B_XINNHBO48_0(.din(n326),.dout(w_dff_B_XINNHBO48_0),.clk(gclk));
	jdff dff_B_dcKwdGaG9_0(.din(n325),.dout(w_dff_B_dcKwdGaG9_0),.clk(gclk));
	jdff dff_B_t95ur5B18_0(.din(w_dff_B_dcKwdGaG9_0),.dout(w_dff_B_t95ur5B18_0),.clk(gclk));
	jdff dff_B_SLajnLwI2_0(.din(w_dff_B_t95ur5B18_0),.dout(w_dff_B_SLajnLwI2_0),.clk(gclk));
	jdff dff_A_BjRnuQXE3_0(.dout(w_G153gat_0[0]),.din(w_dff_A_BjRnuQXE3_0),.clk(gclk));
	jdff dff_A_NTncug3v0_0(.dout(w_dff_A_BjRnuQXE3_0),.din(w_dff_A_NTncug3v0_0),.clk(gclk));
	jdff dff_A_bsnBVwCy1_0(.dout(w_dff_A_NTncug3v0_0),.din(w_dff_A_bsnBVwCy1_0),.clk(gclk));
	jdff dff_A_XwzX1IZ20_0(.dout(w_dff_A_bsnBVwCy1_0),.din(w_dff_A_XwzX1IZ20_0),.clk(gclk));
	jdff dff_A_ub3SxmpZ7_2(.dout(w_G153gat_0[2]),.din(w_dff_A_ub3SxmpZ7_2),.clk(gclk));
	jdff dff_A_S2iu9R9u6_2(.dout(w_dff_A_ub3SxmpZ7_2),.din(w_dff_A_S2iu9R9u6_2),.clk(gclk));
	jdff dff_A_HKtZAJux6_2(.dout(w_dff_A_S2iu9R9u6_2),.din(w_dff_A_HKtZAJux6_2),.clk(gclk));
	jdff dff_A_rlkd52HL6_2(.dout(w_dff_A_HKtZAJux6_2),.din(w_dff_A_rlkd52HL6_2),.clk(gclk));
	jdff dff_A_1sazUBmb2_0(.dout(w_G106gat_0[0]),.din(w_dff_A_1sazUBmb2_0),.clk(gclk));
	jdff dff_A_9Tfmcu5G7_0(.dout(w_dff_A_1sazUBmb2_0),.din(w_dff_A_9Tfmcu5G7_0),.clk(gclk));
	jdff dff_A_hef7QGLh9_0(.dout(w_dff_A_9Tfmcu5G7_0),.din(w_dff_A_hef7QGLh9_0),.clk(gclk));
	jdff dff_A_GbRvA3zS6_0(.dout(w_dff_A_hef7QGLh9_0),.din(w_dff_A_GbRvA3zS6_0),.clk(gclk));
	jdff dff_A_KDGTZ9aa0_1(.dout(w_G177gat_1[1]),.din(w_dff_A_KDGTZ9aa0_1),.clk(gclk));
	jdff dff_A_lbnqP6Tt5_1(.dout(w_dff_A_KDGTZ9aa0_1),.din(w_dff_A_lbnqP6Tt5_1),.clk(gclk));
	jdff dff_A_Lsj4Xj5k0_1(.dout(w_dff_A_lbnqP6Tt5_1),.din(w_dff_A_Lsj4Xj5k0_1),.clk(gclk));
	jdff dff_A_MCWmQIrb5_1(.dout(w_dff_A_Lsj4Xj5k0_1),.din(w_dff_A_MCWmQIrb5_1),.clk(gclk));
	jdff dff_A_QekXYpaX6_1(.dout(w_dff_A_MCWmQIrb5_1),.din(w_dff_A_QekXYpaX6_1),.clk(gclk));
	jdff dff_A_g41BBauG7_2(.dout(w_G177gat_1[2]),.din(w_dff_A_g41BBauG7_2),.clk(gclk));
	jdff dff_A_SDZjQGG05_2(.dout(w_dff_A_g41BBauG7_2),.din(w_dff_A_SDZjQGG05_2),.clk(gclk));
	jdff dff_A_de0TFssx3_2(.dout(w_dff_A_SDZjQGG05_2),.din(w_dff_A_de0TFssx3_2),.clk(gclk));
	jdff dff_A_JGXvROUQ1_2(.dout(w_dff_A_de0TFssx3_2),.din(w_dff_A_JGXvROUQ1_2),.clk(gclk));
	jdff dff_A_2g5bkTSe1_2(.dout(w_dff_A_JGXvROUQ1_2),.din(w_dff_A_2g5bkTSe1_2),.clk(gclk));
	jdff dff_A_YoYoaWoM3_2(.dout(w_G177gat_0[2]),.din(w_dff_A_YoYoaWoM3_2),.clk(gclk));
	jdff dff_A_dSGpSOxS7_2(.dout(w_dff_A_YoYoaWoM3_2),.din(w_dff_A_dSGpSOxS7_2),.clk(gclk));
	jdff dff_A_iQWTMBlT9_2(.dout(w_dff_A_dSGpSOxS7_2),.din(w_dff_A_iQWTMBlT9_2),.clk(gclk));
	jdff dff_A_lK7Kh6sK2_2(.dout(w_dff_A_iQWTMBlT9_2),.din(w_dff_A_lK7Kh6sK2_2),.clk(gclk));
	jdff dff_A_T6w0xhap3_1(.dout(w_n405_0[1]),.din(w_dff_A_T6w0xhap3_1),.clk(gclk));
	jdff dff_A_Z2WIqNpL3_1(.dout(w_dff_A_T6w0xhap3_1),.din(w_dff_A_Z2WIqNpL3_1),.clk(gclk));
	jdff dff_A_hZVUsbC05_1(.dout(w_dff_A_Z2WIqNpL3_1),.din(w_dff_A_hZVUsbC05_1),.clk(gclk));
	jdff dff_B_csxKrAiS0_0(.din(n319),.dout(w_dff_B_csxKrAiS0_0),.clk(gclk));
	jdff dff_B_gsxFArij2_0(.din(n318),.dout(w_dff_B_gsxFArij2_0),.clk(gclk));
	jdff dff_B_9cGXaGUD9_0(.din(w_dff_B_gsxFArij2_0),.dout(w_dff_B_9cGXaGUD9_0),.clk(gclk));
	jdff dff_B_eZOCjBFj3_0(.din(w_dff_B_9cGXaGUD9_0),.dout(w_dff_B_eZOCjBFj3_0),.clk(gclk));
	jdff dff_B_adY790d46_0(.din(n295),.dout(w_dff_B_adY790d46_0),.clk(gclk));
	jdff dff_A_TQAuJOTq3_0(.dout(w_G17gat_1[0]),.din(w_dff_A_TQAuJOTq3_0),.clk(gclk));
	jdff dff_A_19gmqj0u0_2(.dout(w_G17gat_1[2]),.din(w_dff_A_19gmqj0u0_2),.clk(gclk));
	jdff dff_A_0saY8HNr4_2(.dout(w_dff_A_19gmqj0u0_2),.din(w_dff_A_0saY8HNr4_2),.clk(gclk));
	jdff dff_A_Wwlk23wm8_2(.dout(w_dff_A_0saY8HNr4_2),.din(w_dff_A_Wwlk23wm8_2),.clk(gclk));
	jdff dff_A_kSgMlmBC1_0(.dout(w_G80gat_0[0]),.din(w_dff_A_kSgMlmBC1_0),.clk(gclk));
	jdff dff_A_i5nDzkmp4_2(.dout(w_G80gat_0[2]),.din(w_dff_A_i5nDzkmp4_2),.clk(gclk));
	jdff dff_B_zgDD9V7H8_0(.din(n156),.dout(w_dff_B_zgDD9V7H8_0),.clk(gclk));
	jdff dff_A_5jSJjxvG8_0(.dout(w_G55gat_0[0]),.din(w_dff_A_5jSJjxvG8_0),.clk(gclk));
	jdff dff_A_RizNux0Q9_0(.dout(w_dff_A_5jSJjxvG8_0),.din(w_dff_A_RizNux0Q9_0),.clk(gclk));
	jdff dff_A_9yJbgLEK7_0(.dout(w_dff_A_RizNux0Q9_0),.din(w_dff_A_9yJbgLEK7_0),.clk(gclk));
	jdff dff_A_NikhT9437_1(.dout(w_G55gat_0[1]),.din(w_dff_A_NikhT9437_1),.clk(gclk));
	jdff dff_B_mt5ssUfw0_2(.din(G149gat),.dout(w_dff_B_mt5ssUfw0_2),.clk(gclk));
	jdff dff_B_KTo6driW8_2(.din(w_dff_B_mt5ssUfw0_2),.dout(w_dff_B_KTo6driW8_2),.clk(gclk));
	jdff dff_B_ApiLYihH5_2(.din(w_dff_B_KTo6driW8_2),.dout(w_dff_B_ApiLYihH5_2),.clk(gclk));
	jdff dff_B_l7oNFS4D0_2(.din(w_dff_B_ApiLYihH5_2),.dout(w_dff_B_l7oNFS4D0_2),.clk(gclk));
	jdff dff_B_mHbV2ANM1_0(.din(n152),.dout(w_dff_B_mHbV2ANM1_0),.clk(gclk));
	jdff dff_B_nBrgfEWu0_0(.din(n147),.dout(w_dff_B_nBrgfEWu0_0),.clk(gclk));
	jdff dff_A_A8Hsb4HS4_1(.dout(w_G51gat_1[1]),.din(w_dff_A_A8Hsb4HS4_1),.clk(gclk));
	jdff dff_A_pbatWKxq6_1(.dout(w_G1gat_0[1]),.din(w_dff_A_pbatWKxq6_1),.clk(gclk));
	jdff dff_A_Uz76hR5G2_1(.dout(w_G42gat_1[1]),.din(w_dff_A_Uz76hR5G2_1),.clk(gclk));
	jdff dff_A_0XKpT3Ew1_1(.dout(w_G42gat_0[1]),.din(w_dff_A_0XKpT3Ew1_1),.clk(gclk));
	jdff dff_A_QGe30xk99_1(.dout(w_G101gat_0[1]),.din(w_dff_A_QGe30xk99_1),.clk(gclk));
	jdff dff_A_swdxVTFa7_1(.dout(w_dff_A_QGe30xk99_1),.din(w_dff_A_swdxVTFa7_1),.clk(gclk));
	jdff dff_A_VRGvpubH9_1(.dout(w_dff_A_swdxVTFa7_1),.din(w_dff_A_VRGvpubH9_1),.clk(gclk));
	jdff dff_A_s6aV5ion3_1(.dout(w_dff_A_VRGvpubH9_1),.din(w_dff_A_s6aV5ion3_1),.clk(gclk));
	jdff dff_A_n3EUFogI7_1(.dout(w_G171gat_1[1]),.din(w_dff_A_n3EUFogI7_1),.clk(gclk));
	jdff dff_A_sV31scwQ2_1(.dout(w_dff_A_n3EUFogI7_1),.din(w_dff_A_sV31scwQ2_1),.clk(gclk));
	jdff dff_A_PoH7qbrr6_1(.dout(w_dff_A_sV31scwQ2_1),.din(w_dff_A_PoH7qbrr6_1),.clk(gclk));
	jdff dff_A_chaatoJs8_1(.dout(w_dff_A_PoH7qbrr6_1),.din(w_dff_A_chaatoJs8_1),.clk(gclk));
	jdff dff_A_pdHOZErm1_1(.dout(w_dff_A_chaatoJs8_1),.din(w_dff_A_pdHOZErm1_1),.clk(gclk));
	jdff dff_A_E1ZocGjz7_2(.dout(w_G171gat_1[2]),.din(w_dff_A_E1ZocGjz7_2),.clk(gclk));
	jdff dff_A_Z6xMvZQA4_2(.dout(w_dff_A_E1ZocGjz7_2),.din(w_dff_A_Z6xMvZQA4_2),.clk(gclk));
	jdff dff_A_ZYIVTPXM7_2(.dout(w_dff_A_Z6xMvZQA4_2),.din(w_dff_A_ZYIVTPXM7_2),.clk(gclk));
	jdff dff_A_lV20OZUB2_2(.dout(w_dff_A_ZYIVTPXM7_2),.din(w_dff_A_lV20OZUB2_2),.clk(gclk));
	jdff dff_A_qLVc8urX8_2(.dout(w_dff_A_lV20OZUB2_2),.din(w_dff_A_qLVc8urX8_2),.clk(gclk));
	jdff dff_A_setf41397_2(.dout(w_G171gat_0[2]),.din(w_dff_A_setf41397_2),.clk(gclk));
	jdff dff_A_l0tJHxvQ6_2(.dout(w_dff_A_setf41397_2),.din(w_dff_A_l0tJHxvQ6_2),.clk(gclk));
	jdff dff_A_PHjBPaZv9_2(.dout(w_dff_A_l0tJHxvQ6_2),.din(w_dff_A_PHjBPaZv9_2),.clk(gclk));
	jdff dff_A_oD1Gvndw5_2(.dout(w_dff_A_PHjBPaZv9_2),.din(w_dff_A_oD1Gvndw5_2),.clk(gclk));
endmodule

